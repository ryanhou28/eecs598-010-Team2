
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  n2491_lo,
  n2575_lo,
  n2587_lo,
  n2599_lo,
  n2611_lo,
  n2623_lo,
  n2635_lo,
  n2647_lo,
  n2659_lo,
  n2671_lo,
  n2683_lo,
  n2734_lo,
  n2746_lo,
  n2758_lo,
  n2770_lo,
  n2782_lo,
  n2785_lo,
  n2794_lo,
  n2797_lo,
  n2806_lo,
  n2809_lo,
  n2818_lo,
  n2821_lo,
  n2830_lo,
  n2833_lo,
  n2836_lo,
  n2839_lo,
  n2842_lo,
  n2845_lo,
  n2848_lo,
  n2851_lo,
  n2854_lo,
  n2857_lo,
  n2860_lo,
  n2863_lo,
  n4871_o2,
  n4893_o2,
  n4938_o2,
  n5056_o2,
  n5100_o2,
  n5122_o2,
  n5254_o2,
  n5276_o2,
  n5316_o2,
  n5434_o2,
  n5473_o2,
  n5494_o2,
  n5620_o2,
  n5643_o2,
  n5682_o2,
  n5798_o2,
  n5839_o2,
  n5867_o2,
  n6052_o2,
  n6087_o2,
  n6153_o2,
  n6408_o2,
  n6454_o2,
  n6509_o2,
  n6775_o2,
  n6818_o2,
  n6892_o2,
  n5779_o2,
  n5780_o2,
  n7156_o2,
  n5792_o2,
  n7205_o2,
  n5842_o2,
  n5863_o2,
  n7263_o2,
  n5881_o2,
  n5930_o2,
  n5959_o2,
  n5981_o2,
  n6042_o2,
  n6075_o2,
  n6103_o2,
  n7610_o2,
  n6169_o2,
  n7665_o2,
  n6205_o2,
  n6239_o2,
  n7788_o2,
  n6309_o2,
  n6461_o2,
  n6476_o2,
  n325_inv,
  n6545_o2,
  G578_o2,
  G5106_o2,
  n6713_o2,
  G5164_o2,
  n343_inv,
  n6810_o2,
  n6973_o2,
  n352_inv,
  n7053_o2,
  G581_o2,
  G5467_o2,
  n7231_o2,
  G5527_o2,
  n370_inv,
  n7304_o2,
  n7530_o2,
  n379_inv,
  n7653_o2,
  G584_o2,
  G5820_o2,
  n7148_o2,
  n7149_o2,
  n7224_o2,
  n7916_o2,
  G5868_o2,
  n406_inv,
  n7280_o2,
  n7313_o2,
  n8056_o2,
  n7323_o2,
  n7398_o2,
  n7459_o2,
  n7501_o2,
  n7518_o2,
  G563_o2,
  n7606_o2,
  n439_inv,
  n7675_o2,
  G3410_o2,
  n7722_o2,
  n7747_o2,
  n7835_o2,
  G587_o2,
  G6046_o2,
  n7909_o2,
  G566_o2,
  G6070_o2,
  n472_inv,
  n8086_o2,
  n8093_o2,
  G3752_o2,
  n484_inv,
  n8199_o2,
  n2800_lo_buf_o2,
  G548_o2,
  n496_inv,
  G569_o2,
  G1761_o2,
  n505_inv,
  G4101_o2,
  G551_o2,
  n514_inv,
  G4743_o2,
  G5271_o2,
  G5790_o2,
  G6122_o2,
  G2082_o2,
  n2812_lo_buf_o2,
  n2668_lo_buf_o2,
  n2680_lo_buf_o2,
  G572_o2,
  G6125_o2,
  n547_inv,
  n2656_lo_buf_o2,
  G554_o2,
  G4452_o2,
  n559_inv,
  n2644_lo_buf_o2,
  G2410_o2,
  n2632_lo_buf_o2,
  n2620_lo_buf_o2,
  G6131_o2,
  G4693_o2,
  G5209_o2,
  G5741_o2,
  G6082_o2,
  G6119_o2,
  n2608_lo_buf_o2,
  n2596_lo_buf_o2,
  n2584_lo_buf_o2,
  n2572_lo_buf_o2,
  n2704_lo_buf_o2,
  G557_o2,
  G5936_o2,
  G5442_o2,
  G4926_o2,
  G6134_o2,
  G3929_o2,
  G4425_o2,
  G4947_o2,
  n2764_lo_buf_o2,
  n634_inv,
  n2560_lo_buf_o2,
  n2824_lo_buf_o2,
  G575_o2,
  G2740_o2,
  n649_inv,
  n2548_lo_buf_o2,
  n2536_lo_buf_o2,
  n2524_lo_buf_o2,
  G875_o2,
  G1064_o2,
  G1253_o2,
  G6140_o2,
  G5151_o2,
  G5686_o2,
  G6061_o2,
  G4803_o2,
  G5332_o2,
  G5844_o2,
  G6114_o2,
  G4806_o2,
  G3881_o2,
  G4370_o2,
  G4896_o2,
  G5001_o2,
  G3121_o2,
  n2512_lo_buf_o2,
  G4085_o2,
  G4605_o2,
  G5118_o2,
  G4997_o2,
  n2500_lo_buf_o2,
  n2716_lo_buf_o2,
  G560_o2,
  G1895_o2,
  G3064_o2,
  G3269_o2,
  G3569_o2,
  n748_inv,
  G1196_o2,
  G1007_o2,
  G818_o2,
  G674_o2,
  G5041_o2,
  G5562_o2,
  G6005_o2,
  G5214_o2,
  G5746_o2,
  G6087_o2,
  G6086_o2,
  G5745_o2,
  G5213_o2,
  G5893_o2,
  G5391_o2,
  G4864_o2,
  G6143_o2,
  G6008_o2,
  G5565_o2,
  G5044_o2,
  G3813_o2,
  G4325_o2,
  G4834_o2,
  G4993_o2,
  G3989_o2,
  G4490_o2,
  G5011_o2,
  G5112_o2,
  n2776_lo_buf_o2,
  G3298_o2,
  G3073_o2,
  G3265_o2,
  G3624_o2,
  G1642_o2,
  G1980_o2,
  n2488_lo_buf_o2,
  G626_o2,
  G1139_o2,
  G950_o2,
  G707_o2,
  G545_o2,
  G4217_o2,
  G4716_o2,
  G5244_o2,
  G3136_o2,
  G3499_o2,
  G3885_o2,
  G5243_o2,
  G3886_o2,
  G4375_o2,
  G4901_o2,
  G5054_o2,
  G4374_o2,
  G4900_o2,
  G5053_o2,
  G5242_o2,
  G4034_o2,
  G4556_o2,
  G5064_o2,
  G5172_o2,
  G2030_o2,
  G3016_o2,
  G3520_o2,
  G3261_o2,
  G3620_o2,
  G4220_o2,
  G4719_o2,
  G5247_o2,
  G5109_o2,
  G1638_o2,
  G1976_o2,
  G3560_o2,
  G3205_o2,
  G3193_o2,
  G3367_o2,
  G3670_o2,
  n979_inv,
  G1280_o2,
  G902_o2,
  G659_o2,
  G983_o2,
  G740_o2,
  G2917_o2,
  G3391_o2,
  G3494_o2,
  G1512_o2,
  G1854_o2,
  G2203_o2,
  G3493_o2,
  G3069_o2,
  G3574_o2,
  G3319_o2,
  G3667_o2,
  G3068_o2,
  G3573_o2,
  G3666_o2,
  G3318_o2,
  G3492_o2,
  G3241_o2,
  G3722_o2,
  G3422_o2,
  G1445_o2,
  G3257_o2,
  G3616_o2,
  G1634_o2,
  G1972_o2,
  G2256_o2,
  G3394_o2,
  G3557_o2,
  G3364_o2,
  G3719_o2,
  G2253_o2,
  G1583_o2,
  G1917_o2,
  G1727_o2,
  G2061_o2,
  G935_o2,
  G692_o2,
  G2136_o2,
  G1507_o2,
  G1849_o2,
  G2198_o2,
  G2197_o2,
  G1848_o2,
  G1689_o2,
  G2016_o2,
  G2314_o2,
  G2313_o2,
  G1688_o2,
  G2015_o2,
  G1847_o2,
  G2196_o2,
  G2118_o2,
  G1777_o2,
  G1630_o2,
  G1968_o2,
  G2309_o2,
  G2139_o2,
  G1580_o2,
  G2250_o2,
  G1914_o2,
  G1724_o2,
  G2058_o2,
  n2728_lo_buf_o2,
  G6257,
  G6258,
  G6259,
  G6260,
  G6261,
  G6262,
  G6263,
  G6264,
  G6265,
  G6266,
  G6267,
  G6268,
  G6269,
  G6270,
  G6271,
  G6272,
  G6273,
  G6274,
  G6275,
  G6276,
  G6277,
  G6278,
  G6279,
  G6280,
  G6281,
  G6282,
  G6283,
  G6284,
  G6285,
  G6286,
  G6287,
  G6288,
  n2491_li,
  n2575_li,
  n2587_li,
  n2599_li,
  n2611_li,
  n2623_li,
  n2635_li,
  n2647_li,
  n2659_li,
  n2671_li,
  n2683_li,
  n2734_li,
  n2746_li,
  n2758_li,
  n2770_li,
  n2782_li,
  n2785_li,
  n2794_li,
  n2797_li,
  n2806_li,
  n2809_li,
  n2818_li,
  n2821_li,
  n2830_li,
  n2833_li,
  n2836_li,
  n2839_li,
  n2842_li,
  n2845_li,
  n2848_li,
  n2851_li,
  n2854_li,
  n2857_li,
  n2860_li,
  n2863_li,
  n4871_i2,
  n4893_i2,
  n4938_i2,
  n5056_i2,
  n5100_i2,
  n5122_i2,
  n5254_i2,
  n5276_i2,
  n5316_i2,
  n5434_i2,
  n5473_i2,
  n5494_i2,
  n5620_i2,
  n5643_i2,
  n5682_i2,
  n5798_i2,
  n5839_i2,
  n5867_i2,
  n6052_i2,
  n6087_i2,
  n6153_i2,
  n6408_i2,
  n6454_i2,
  n6509_i2,
  n6775_i2,
  n6818_i2,
  n6892_i2,
  n5779_i2,
  n5780_i2,
  n7156_i2,
  n5792_i2,
  n7205_i2,
  n5842_i2,
  n5863_i2,
  n7263_i2,
  n5881_i2,
  n5930_i2,
  n5959_i2,
  n5981_i2,
  n6042_i2,
  n6075_i2,
  n6103_i2,
  n7610_i2,
  n6169_i2,
  n7665_i2,
  n6205_i2,
  n6239_i2,
  n7788_i2,
  n6309_i2,
  n6461_i2,
  n6476_i2,
  n6521_i2,
  n6545_i2,
  G578_i2,
  G5106_i2,
  n6713_i2,
  G5164_i2,
  n6771_i2,
  n6810_i2,
  n6973_i2,
  n6995_i2,
  n7053_i2,
  G581_i2,
  G5467_i2,
  n7231_i2,
  G5527_i2,
  n7277_i2,
  n7304_i2,
  n7530_i2,
  n7595_i2,
  n7653_i2,
  G584_i2,
  G5820_i2,
  n7148_i2,
  n7149_i2,
  n7224_i2,
  n7916_i2,
  G5868_i2,
  n7958_i2,
  n7280_i2,
  n7313_i2,
  n8056_i2,
  n7323_i2,
  n7398_i2,
  n7459_i2,
  n7501_i2,
  n7518_i2,
  G563_i2,
  n7606_i2,
  G3358_i2,
  n7675_i2,
  G3410_i2,
  n7722_i2,
  n7747_i2,
  n7835_i2,
  G587_i2,
  G6046_i2,
  n7909_i2,
  G566_i2,
  G6070_i2,
  G3698_i2,
  n8086_i2,
  n8093_i2,
  G3752_i2,
  n8156_i2,
  n8199_i2,
  n2800_lo_buf_i2,
  G548_i2,
  G1715_i2,
  G569_i2,
  G1761_i2,
  G4043_i2,
  G4101_i2,
  G551_i2,
  G2034_i2,
  G4743_i2,
  G5271_i2,
  G5790_i2,
  G6122_i2,
  G2082_i2,
  n2812_lo_buf_i2,
  n2668_lo_buf_i2,
  n2680_lo_buf_i2,
  G572_i2,
  G6125_i2,
  G4395_i2,
  n2656_lo_buf_i2,
  G554_i2,
  G4452_i2,
  G2358_i2,
  n2644_lo_buf_i2,
  G2410_i2,
  n2632_lo_buf_i2,
  n2620_lo_buf_i2,
  G6131_i2,
  G4693_i2,
  G5209_i2,
  G5741_i2,
  G6082_i2,
  G6119_i2,
  n2608_lo_buf_i2,
  n2596_lo_buf_i2,
  n2584_lo_buf_i2,
  n2572_lo_buf_i2,
  n2704_lo_buf_i2,
  G557_i2,
  G5936_i2,
  G5442_i2,
  G4926_i2,
  G6134_i2,
  G3929_i2,
  G4425_i2,
  G4947_i2,
  n2764_lo_buf_i2,
  G2689_i2,
  n2560_lo_buf_i2,
  n2824_lo_buf_i2,
  G575_i2,
  G2740_i2,
  G4749_i2,
  n2548_lo_buf_i2,
  n2536_lo_buf_i2,
  n2524_lo_buf_i2,
  G875_i2,
  G1064_i2,
  G1253_i2,
  G6140_i2,
  G5151_i2,
  G5686_i2,
  G6061_i2,
  G4803_i2,
  G5332_i2,
  G5844_i2,
  G6114_i2,
  G4806_i2,
  G3881_i2,
  G4370_i2,
  G4896_i2,
  G5001_i2,
  G3121_i2,
  n2512_lo_buf_i2,
  G4085_i2,
  G4605_i2,
  G5118_i2,
  G4997_i2,
  n2500_lo_buf_i2,
  n2716_lo_buf_i2,
  G560_i2,
  G1895_i2,
  G3064_i2,
  G3269_i2,
  G3569_i2,
  G3022_i2,
  G1196_i2,
  G1007_i2,
  G818_i2,
  G674_i2,
  G5041_i2,
  G5562_i2,
  G6005_i2,
  G5214_i2,
  G5746_i2,
  G6087_i2,
  G6086_i2,
  G5745_i2,
  G5213_i2,
  G5893_i2,
  G5391_i2,
  G4864_i2,
  G6143_i2,
  G6008_i2,
  G5565_i2,
  G5044_i2,
  G3813_i2,
  G4325_i2,
  G4834_i2,
  G4993_i2,
  G3989_i2,
  G4490_i2,
  G5011_i2,
  G5112_i2,
  n2776_lo_buf_i2,
  G3298_i2,
  G3073_i2,
  G3265_i2,
  G3624_i2,
  G1642_i2,
  G1980_i2,
  n2488_lo_buf_i2,
  G626_i2,
  G1139_i2,
  G950_i2,
  G707_i2,
  G545_i2,
  G4217_i2,
  G4716_i2,
  G5244_i2,
  G3136_i2,
  G3499_i2,
  G3885_i2,
  G5243_i2,
  G3886_i2,
  G4375_i2,
  G4901_i2,
  G5054_i2,
  G4374_i2,
  G4900_i2,
  G5053_i2,
  G5242_i2,
  G4034_i2,
  G4556_i2,
  G5064_i2,
  G5172_i2,
  G2030_i2,
  G3016_i2,
  G3520_i2,
  G3261_i2,
  G3620_i2,
  G4220_i2,
  G4719_i2,
  G5247_i2,
  G5109_i2,
  G1638_i2,
  G1976_i2,
  G3560_i2,
  G3205_i2,
  G3193_i2,
  G3367_i2,
  G3670_i2,
  G1400_i2,
  G1280_i2,
  G902_i2,
  G659_i2,
  G983_i2,
  G740_i2,
  G2917_i2,
  G3391_i2,
  G3494_i2,
  G1512_i2,
  G1854_i2,
  G2203_i2,
  G3493_i2,
  G3069_i2,
  G3574_i2,
  G3319_i2,
  G3667_i2,
  G3068_i2,
  G3573_i2,
  G3666_i2,
  G3318_i2,
  G3492_i2,
  G3241_i2,
  G3722_i2,
  G3422_i2,
  G1445_i2,
  G3257_i2,
  G3616_i2,
  G1634_i2,
  G1972_i2,
  G2256_i2,
  G3394_i2,
  G3557_i2,
  G3364_i2,
  G3719_i2,
  G2253_i2,
  G1583_i2,
  G1917_i2,
  G1727_i2,
  G2061_i2,
  G935_i2,
  G692_i2,
  G2136_i2,
  G1507_i2,
  G1849_i2,
  G2198_i2,
  G2197_i2,
  G1848_i2,
  G1689_i2,
  G2016_i2,
  G2314_i2,
  G2313_i2,
  G1688_i2,
  G2015_i2,
  G1847_i2,
  G2196_i2,
  G2118_i2,
  G1777_i2,
  G1630_i2,
  G1968_i2,
  G2309_i2,
  G2139_i2,
  G1580_i2,
  G2250_i2,
  G1914_i2,
  G1724_i2,
  G2058_i2,
  n2728_lo_buf_i2
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input n2491_lo;input n2575_lo;input n2587_lo;input n2599_lo;input n2611_lo;input n2623_lo;input n2635_lo;input n2647_lo;input n2659_lo;input n2671_lo;input n2683_lo;input n2734_lo;input n2746_lo;input n2758_lo;input n2770_lo;input n2782_lo;input n2785_lo;input n2794_lo;input n2797_lo;input n2806_lo;input n2809_lo;input n2818_lo;input n2821_lo;input n2830_lo;input n2833_lo;input n2836_lo;input n2839_lo;input n2842_lo;input n2845_lo;input n2848_lo;input n2851_lo;input n2854_lo;input n2857_lo;input n2860_lo;input n2863_lo;input n4871_o2;input n4893_o2;input n4938_o2;input n5056_o2;input n5100_o2;input n5122_o2;input n5254_o2;input n5276_o2;input n5316_o2;input n5434_o2;input n5473_o2;input n5494_o2;input n5620_o2;input n5643_o2;input n5682_o2;input n5798_o2;input n5839_o2;input n5867_o2;input n6052_o2;input n6087_o2;input n6153_o2;input n6408_o2;input n6454_o2;input n6509_o2;input n6775_o2;input n6818_o2;input n6892_o2;input n5779_o2;input n5780_o2;input n7156_o2;input n5792_o2;input n7205_o2;input n5842_o2;input n5863_o2;input n7263_o2;input n5881_o2;input n5930_o2;input n5959_o2;input n5981_o2;input n6042_o2;input n6075_o2;input n6103_o2;input n7610_o2;input n6169_o2;input n7665_o2;input n6205_o2;input n6239_o2;input n7788_o2;input n6309_o2;input n6461_o2;input n6476_o2;input n325_inv;input n6545_o2;input G578_o2;input G5106_o2;input n6713_o2;input G5164_o2;input n343_inv;input n6810_o2;input n6973_o2;input n352_inv;input n7053_o2;input G581_o2;input G5467_o2;input n7231_o2;input G5527_o2;input n370_inv;input n7304_o2;input n7530_o2;input n379_inv;input n7653_o2;input G584_o2;input G5820_o2;input n7148_o2;input n7149_o2;input n7224_o2;input n7916_o2;input G5868_o2;input n406_inv;input n7280_o2;input n7313_o2;input n8056_o2;input n7323_o2;input n7398_o2;input n7459_o2;input n7501_o2;input n7518_o2;input G563_o2;input n7606_o2;input n439_inv;input n7675_o2;input G3410_o2;input n7722_o2;input n7747_o2;input n7835_o2;input G587_o2;input G6046_o2;input n7909_o2;input G566_o2;input G6070_o2;input n472_inv;input n8086_o2;input n8093_o2;input G3752_o2;input n484_inv;input n8199_o2;input n2800_lo_buf_o2;input G548_o2;input n496_inv;input G569_o2;input G1761_o2;input n505_inv;input G4101_o2;input G551_o2;input n514_inv;input G4743_o2;input G5271_o2;input G5790_o2;input G6122_o2;input G2082_o2;input n2812_lo_buf_o2;input n2668_lo_buf_o2;input n2680_lo_buf_o2;input G572_o2;input G6125_o2;input n547_inv;input n2656_lo_buf_o2;input G554_o2;input G4452_o2;input n559_inv;input n2644_lo_buf_o2;input G2410_o2;input n2632_lo_buf_o2;input n2620_lo_buf_o2;input G6131_o2;input G4693_o2;input G5209_o2;input G5741_o2;input G6082_o2;input G6119_o2;input n2608_lo_buf_o2;input n2596_lo_buf_o2;input n2584_lo_buf_o2;input n2572_lo_buf_o2;input n2704_lo_buf_o2;input G557_o2;input G5936_o2;input G5442_o2;input G4926_o2;input G6134_o2;input G3929_o2;input G4425_o2;input G4947_o2;input n2764_lo_buf_o2;input n634_inv;input n2560_lo_buf_o2;input n2824_lo_buf_o2;input G575_o2;input G2740_o2;input n649_inv;input n2548_lo_buf_o2;input n2536_lo_buf_o2;input n2524_lo_buf_o2;input G875_o2;input G1064_o2;input G1253_o2;input G6140_o2;input G5151_o2;input G5686_o2;input G6061_o2;input G4803_o2;input G5332_o2;input G5844_o2;input G6114_o2;input G4806_o2;input G3881_o2;input G4370_o2;input G4896_o2;input G5001_o2;input G3121_o2;input n2512_lo_buf_o2;input G4085_o2;input G4605_o2;input G5118_o2;input G4997_o2;input n2500_lo_buf_o2;input n2716_lo_buf_o2;input G560_o2;input G1895_o2;input G3064_o2;input G3269_o2;input G3569_o2;input n748_inv;input G1196_o2;input G1007_o2;input G818_o2;input G674_o2;input G5041_o2;input G5562_o2;input G6005_o2;input G5214_o2;input G5746_o2;input G6087_o2;input G6086_o2;input G5745_o2;input G5213_o2;input G5893_o2;input G5391_o2;input G4864_o2;input G6143_o2;input G6008_o2;input G5565_o2;input G5044_o2;input G3813_o2;input G4325_o2;input G4834_o2;input G4993_o2;input G3989_o2;input G4490_o2;input G5011_o2;input G5112_o2;input n2776_lo_buf_o2;input G3298_o2;input G3073_o2;input G3265_o2;input G3624_o2;input G1642_o2;input G1980_o2;input n2488_lo_buf_o2;input G626_o2;input G1139_o2;input G950_o2;input G707_o2;input G545_o2;input G4217_o2;input G4716_o2;input G5244_o2;input G3136_o2;input G3499_o2;input G3885_o2;input G5243_o2;input G3886_o2;input G4375_o2;input G4901_o2;input G5054_o2;input G4374_o2;input G4900_o2;input G5053_o2;input G5242_o2;input G4034_o2;input G4556_o2;input G5064_o2;input G5172_o2;input G2030_o2;input G3016_o2;input G3520_o2;input G3261_o2;input G3620_o2;input G4220_o2;input G4719_o2;input G5247_o2;input G5109_o2;input G1638_o2;input G1976_o2;input G3560_o2;input G3205_o2;input G3193_o2;input G3367_o2;input G3670_o2;input n979_inv;input G1280_o2;input G902_o2;input G659_o2;input G983_o2;input G740_o2;input G2917_o2;input G3391_o2;input G3494_o2;input G1512_o2;input G1854_o2;input G2203_o2;input G3493_o2;input G3069_o2;input G3574_o2;input G3319_o2;input G3667_o2;input G3068_o2;input G3573_o2;input G3666_o2;input G3318_o2;input G3492_o2;input G3241_o2;input G3722_o2;input G3422_o2;input G1445_o2;input G3257_o2;input G3616_o2;input G1634_o2;input G1972_o2;input G2256_o2;input G3394_o2;input G3557_o2;input G3364_o2;input G3719_o2;input G2253_o2;input G1583_o2;input G1917_o2;input G1727_o2;input G2061_o2;input G935_o2;input G692_o2;input G2136_o2;input G1507_o2;input G1849_o2;input G2198_o2;input G2197_o2;input G1848_o2;input G1689_o2;input G2016_o2;input G2314_o2;input G2313_o2;input G1688_o2;input G2015_o2;input G1847_o2;input G2196_o2;input G2118_o2;input G1777_o2;input G1630_o2;input G1968_o2;input G2309_o2;input G2139_o2;input G1580_o2;input G2250_o2;input G1914_o2;input G1724_o2;input G2058_o2;input n2728_lo_buf_o2;
  output G6257;output G6258;output G6259;output G6260;output G6261;output G6262;output G6263;output G6264;output G6265;output G6266;output G6267;output G6268;output G6269;output G6270;output G6271;output G6272;output G6273;output G6274;output G6275;output G6276;output G6277;output G6278;output G6279;output G6280;output G6281;output G6282;output G6283;output G6284;output G6285;output G6286;output G6287;output G6288;output n2491_li;output n2575_li;output n2587_li;output n2599_li;output n2611_li;output n2623_li;output n2635_li;output n2647_li;output n2659_li;output n2671_li;output n2683_li;output n2734_li;output n2746_li;output n2758_li;output n2770_li;output n2782_li;output n2785_li;output n2794_li;output n2797_li;output n2806_li;output n2809_li;output n2818_li;output n2821_li;output n2830_li;output n2833_li;output n2836_li;output n2839_li;output n2842_li;output n2845_li;output n2848_li;output n2851_li;output n2854_li;output n2857_li;output n2860_li;output n2863_li;output n4871_i2;output n4893_i2;output n4938_i2;output n5056_i2;output n5100_i2;output n5122_i2;output n5254_i2;output n5276_i2;output n5316_i2;output n5434_i2;output n5473_i2;output n5494_i2;output n5620_i2;output n5643_i2;output n5682_i2;output n5798_i2;output n5839_i2;output n5867_i2;output n6052_i2;output n6087_i2;output n6153_i2;output n6408_i2;output n6454_i2;output n6509_i2;output n6775_i2;output n6818_i2;output n6892_i2;output n5779_i2;output n5780_i2;output n7156_i2;output n5792_i2;output n7205_i2;output n5842_i2;output n5863_i2;output n7263_i2;output n5881_i2;output n5930_i2;output n5959_i2;output n5981_i2;output n6042_i2;output n6075_i2;output n6103_i2;output n7610_i2;output n6169_i2;output n7665_i2;output n6205_i2;output n6239_i2;output n7788_i2;output n6309_i2;output n6461_i2;output n6476_i2;output n6521_i2;output n6545_i2;output G578_i2;output G5106_i2;output n6713_i2;output G5164_i2;output n6771_i2;output n6810_i2;output n6973_i2;output n6995_i2;output n7053_i2;output G581_i2;output G5467_i2;output n7231_i2;output G5527_i2;output n7277_i2;output n7304_i2;output n7530_i2;output n7595_i2;output n7653_i2;output G584_i2;output G5820_i2;output n7148_i2;output n7149_i2;output n7224_i2;output n7916_i2;output G5868_i2;output n7958_i2;output n7280_i2;output n7313_i2;output n8056_i2;output n7323_i2;output n7398_i2;output n7459_i2;output n7501_i2;output n7518_i2;output G563_i2;output n7606_i2;output G3358_i2;output n7675_i2;output G3410_i2;output n7722_i2;output n7747_i2;output n7835_i2;output G587_i2;output G6046_i2;output n7909_i2;output G566_i2;output G6070_i2;output G3698_i2;output n8086_i2;output n8093_i2;output G3752_i2;output n8156_i2;output n8199_i2;output n2800_lo_buf_i2;output G548_i2;output G1715_i2;output G569_i2;output G1761_i2;output G4043_i2;output G4101_i2;output G551_i2;output G2034_i2;output G4743_i2;output G5271_i2;output G5790_i2;output G6122_i2;output G2082_i2;output n2812_lo_buf_i2;output n2668_lo_buf_i2;output n2680_lo_buf_i2;output G572_i2;output G6125_i2;output G4395_i2;output n2656_lo_buf_i2;output G554_i2;output G4452_i2;output G2358_i2;output n2644_lo_buf_i2;output G2410_i2;output n2632_lo_buf_i2;output n2620_lo_buf_i2;output G6131_i2;output G4693_i2;output G5209_i2;output G5741_i2;output G6082_i2;output G6119_i2;output n2608_lo_buf_i2;output n2596_lo_buf_i2;output n2584_lo_buf_i2;output n2572_lo_buf_i2;output n2704_lo_buf_i2;output G557_i2;output G5936_i2;output G5442_i2;output G4926_i2;output G6134_i2;output G3929_i2;output G4425_i2;output G4947_i2;output n2764_lo_buf_i2;output G2689_i2;output n2560_lo_buf_i2;output n2824_lo_buf_i2;output G575_i2;output G2740_i2;output G4749_i2;output n2548_lo_buf_i2;output n2536_lo_buf_i2;output n2524_lo_buf_i2;output G875_i2;output G1064_i2;output G1253_i2;output G6140_i2;output G5151_i2;output G5686_i2;output G6061_i2;output G4803_i2;output G5332_i2;output G5844_i2;output G6114_i2;output G4806_i2;output G3881_i2;output G4370_i2;output G4896_i2;output G5001_i2;output G3121_i2;output n2512_lo_buf_i2;output G4085_i2;output G4605_i2;output G5118_i2;output G4997_i2;output n2500_lo_buf_i2;output n2716_lo_buf_i2;output G560_i2;output G1895_i2;output G3064_i2;output G3269_i2;output G3569_i2;output G3022_i2;output G1196_i2;output G1007_i2;output G818_i2;output G674_i2;output G5041_i2;output G5562_i2;output G6005_i2;output G5214_i2;output G5746_i2;output G6087_i2;output G6086_i2;output G5745_i2;output G5213_i2;output G5893_i2;output G5391_i2;output G4864_i2;output G6143_i2;output G6008_i2;output G5565_i2;output G5044_i2;output G3813_i2;output G4325_i2;output G4834_i2;output G4993_i2;output G3989_i2;output G4490_i2;output G5011_i2;output G5112_i2;output n2776_lo_buf_i2;output G3298_i2;output G3073_i2;output G3265_i2;output G3624_i2;output G1642_i2;output G1980_i2;output n2488_lo_buf_i2;output G626_i2;output G1139_i2;output G950_i2;output G707_i2;output G545_i2;output G4217_i2;output G4716_i2;output G5244_i2;output G3136_i2;output G3499_i2;output G3885_i2;output G5243_i2;output G3886_i2;output G4375_i2;output G4901_i2;output G5054_i2;output G4374_i2;output G4900_i2;output G5053_i2;output G5242_i2;output G4034_i2;output G4556_i2;output G5064_i2;output G5172_i2;output G2030_i2;output G3016_i2;output G3520_i2;output G3261_i2;output G3620_i2;output G4220_i2;output G4719_i2;output G5247_i2;output G5109_i2;output G1638_i2;output G1976_i2;output G3560_i2;output G3205_i2;output G3193_i2;output G3367_i2;output G3670_i2;output G1400_i2;output G1280_i2;output G902_i2;output G659_i2;output G983_i2;output G740_i2;output G2917_i2;output G3391_i2;output G3494_i2;output G1512_i2;output G1854_i2;output G2203_i2;output G3493_i2;output G3069_i2;output G3574_i2;output G3319_i2;output G3667_i2;output G3068_i2;output G3573_i2;output G3666_i2;output G3318_i2;output G3492_i2;output G3241_i2;output G3722_i2;output G3422_i2;output G1445_i2;output G3257_i2;output G3616_i2;output G1634_i2;output G1972_i2;output G2256_i2;output G3394_i2;output G3557_i2;output G3364_i2;output G3719_i2;output G2253_i2;output G1583_i2;output G1917_i2;output G1727_i2;output G2061_i2;output G935_i2;output G692_i2;output G2136_i2;output G1507_i2;output G1849_i2;output G2198_i2;output G2197_i2;output G1848_i2;output G1689_i2;output G2016_i2;output G2314_i2;output G2313_i2;output G1688_i2;output G2015_i2;output G1847_i2;output G2196_i2;output G2118_i2;output G1777_i2;output G1630_i2;output G1968_i2;output G2309_i2;output G2139_i2;output G1580_i2;output G2250_i2;output G1914_i2;output G1724_i2;output G2058_i2;output n2728_lo_buf_i2;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire n2491_lo_p;
  wire n2491_lo_n;
  wire n2575_lo_p;
  wire n2575_lo_n;
  wire n2587_lo_p;
  wire n2587_lo_n;
  wire n2599_lo_p;
  wire n2599_lo_n;
  wire n2611_lo_p;
  wire n2611_lo_n;
  wire n2623_lo_p;
  wire n2623_lo_n;
  wire n2635_lo_p;
  wire n2635_lo_n;
  wire n2647_lo_p;
  wire n2647_lo_n;
  wire n2659_lo_p;
  wire n2659_lo_n;
  wire n2671_lo_p;
  wire n2671_lo_n;
  wire n2683_lo_p;
  wire n2683_lo_n;
  wire n2734_lo_p;
  wire n2734_lo_n;
  wire n2746_lo_p;
  wire n2746_lo_n;
  wire n2758_lo_p;
  wire n2758_lo_n;
  wire n2770_lo_p;
  wire n2770_lo_n;
  wire n2782_lo_p;
  wire n2782_lo_n;
  wire n2785_lo_p;
  wire n2785_lo_n;
  wire n2794_lo_p;
  wire n2794_lo_n;
  wire n2797_lo_p;
  wire n2797_lo_n;
  wire n2806_lo_p;
  wire n2806_lo_n;
  wire n2809_lo_p;
  wire n2809_lo_n;
  wire n2818_lo_p;
  wire n2818_lo_n;
  wire n2821_lo_p;
  wire n2821_lo_n;
  wire n2830_lo_p;
  wire n2830_lo_n;
  wire n2833_lo_p;
  wire n2833_lo_n;
  wire n2836_lo_p;
  wire n2836_lo_n;
  wire n2839_lo_p;
  wire n2839_lo_n;
  wire n2842_lo_p;
  wire n2842_lo_n;
  wire n2845_lo_p;
  wire n2845_lo_n;
  wire n2848_lo_p;
  wire n2848_lo_n;
  wire n2851_lo_p;
  wire n2851_lo_n;
  wire n2854_lo_p;
  wire n2854_lo_n;
  wire n2857_lo_p;
  wire n2857_lo_n;
  wire n2860_lo_p;
  wire n2860_lo_n;
  wire n2863_lo_p;
  wire n2863_lo_n;
  wire n4871_o2_p;
  wire n4871_o2_n;
  wire n4893_o2_p;
  wire n4893_o2_n;
  wire n4938_o2_p;
  wire n4938_o2_n;
  wire n5056_o2_p;
  wire n5056_o2_n;
  wire n5100_o2_p;
  wire n5100_o2_n;
  wire n5122_o2_p;
  wire n5122_o2_n;
  wire n5254_o2_p;
  wire n5254_o2_n;
  wire n5276_o2_p;
  wire n5276_o2_n;
  wire n5316_o2_p;
  wire n5316_o2_n;
  wire n5434_o2_p;
  wire n5434_o2_n;
  wire n5473_o2_p;
  wire n5473_o2_n;
  wire n5494_o2_p;
  wire n5494_o2_n;
  wire n5620_o2_p;
  wire n5620_o2_n;
  wire n5643_o2_p;
  wire n5643_o2_n;
  wire n5682_o2_p;
  wire n5682_o2_n;
  wire n5798_o2_p;
  wire n5798_o2_n;
  wire n5839_o2_p;
  wire n5839_o2_n;
  wire n5867_o2_p;
  wire n5867_o2_n;
  wire n6052_o2_p;
  wire n6052_o2_n;
  wire n6087_o2_p;
  wire n6087_o2_n;
  wire n6153_o2_p;
  wire n6153_o2_n;
  wire n6408_o2_p;
  wire n6408_o2_n;
  wire n6454_o2_p;
  wire n6454_o2_n;
  wire n6509_o2_p;
  wire n6509_o2_n;
  wire n6775_o2_p;
  wire n6775_o2_n;
  wire n6818_o2_p;
  wire n6818_o2_n;
  wire n6892_o2_p;
  wire n6892_o2_n;
  wire n5779_o2_p;
  wire n5779_o2_n;
  wire n5780_o2_p;
  wire n5780_o2_n;
  wire n7156_o2_p;
  wire n7156_o2_n;
  wire n5792_o2_p;
  wire n5792_o2_n;
  wire n7205_o2_p;
  wire n7205_o2_n;
  wire n5842_o2_p;
  wire n5842_o2_n;
  wire n5863_o2_p;
  wire n5863_o2_n;
  wire n7263_o2_p;
  wire n7263_o2_n;
  wire n5881_o2_p;
  wire n5881_o2_n;
  wire n5930_o2_p;
  wire n5930_o2_n;
  wire n5959_o2_p;
  wire n5959_o2_n;
  wire n5981_o2_p;
  wire n5981_o2_n;
  wire n6042_o2_p;
  wire n6042_o2_n;
  wire n6075_o2_p;
  wire n6075_o2_n;
  wire n6103_o2_p;
  wire n6103_o2_n;
  wire n7610_o2_p;
  wire n7610_o2_n;
  wire n6169_o2_p;
  wire n6169_o2_n;
  wire n7665_o2_p;
  wire n7665_o2_n;
  wire n6205_o2_p;
  wire n6205_o2_n;
  wire n6239_o2_p;
  wire n6239_o2_n;
  wire n7788_o2_p;
  wire n7788_o2_n;
  wire n6309_o2_p;
  wire n6309_o2_n;
  wire n6461_o2_p;
  wire n6461_o2_n;
  wire n6476_o2_p;
  wire n6476_o2_n;
  wire n325_inv_p;
  wire n325_inv_n;
  wire n6545_o2_p;
  wire n6545_o2_n;
  wire G578_o2_p;
  wire G578_o2_n;
  wire G5106_o2_p;
  wire G5106_o2_n;
  wire n6713_o2_p;
  wire n6713_o2_n;
  wire G5164_o2_p;
  wire G5164_o2_n;
  wire n343_inv_p;
  wire n343_inv_n;
  wire n6810_o2_p;
  wire n6810_o2_n;
  wire n6973_o2_p;
  wire n6973_o2_n;
  wire n352_inv_p;
  wire n352_inv_n;
  wire n7053_o2_p;
  wire n7053_o2_n;
  wire G581_o2_p;
  wire G581_o2_n;
  wire G5467_o2_p;
  wire G5467_o2_n;
  wire n7231_o2_p;
  wire n7231_o2_n;
  wire G5527_o2_p;
  wire G5527_o2_n;
  wire n370_inv_p;
  wire n370_inv_n;
  wire n7304_o2_p;
  wire n7304_o2_n;
  wire n7530_o2_p;
  wire n7530_o2_n;
  wire n379_inv_p;
  wire n379_inv_n;
  wire n7653_o2_p;
  wire n7653_o2_n;
  wire G584_o2_p;
  wire G584_o2_n;
  wire G5820_o2_p;
  wire G5820_o2_n;
  wire n7148_o2_p;
  wire n7148_o2_n;
  wire n7149_o2_p;
  wire n7149_o2_n;
  wire n7224_o2_p;
  wire n7224_o2_n;
  wire n7916_o2_p;
  wire n7916_o2_n;
  wire G5868_o2_p;
  wire G5868_o2_n;
  wire n406_inv_p;
  wire n406_inv_n;
  wire n7280_o2_p;
  wire n7280_o2_n;
  wire n7313_o2_p;
  wire n7313_o2_n;
  wire n8056_o2_p;
  wire n8056_o2_n;
  wire n7323_o2_p;
  wire n7323_o2_n;
  wire n7398_o2_p;
  wire n7398_o2_n;
  wire n7459_o2_p;
  wire n7459_o2_n;
  wire n7501_o2_p;
  wire n7501_o2_n;
  wire n7518_o2_p;
  wire n7518_o2_n;
  wire G563_o2_p;
  wire G563_o2_n;
  wire n7606_o2_p;
  wire n7606_o2_n;
  wire n439_inv_p;
  wire n439_inv_n;
  wire n7675_o2_p;
  wire n7675_o2_n;
  wire G3410_o2_p;
  wire G3410_o2_n;
  wire n7722_o2_p;
  wire n7722_o2_n;
  wire n7747_o2_p;
  wire n7747_o2_n;
  wire n7835_o2_p;
  wire n7835_o2_n;
  wire G587_o2_p;
  wire G587_o2_n;
  wire G6046_o2_p;
  wire G6046_o2_n;
  wire n7909_o2_p;
  wire n7909_o2_n;
  wire G566_o2_p;
  wire G566_o2_n;
  wire G6070_o2_p;
  wire G6070_o2_n;
  wire n472_inv_p;
  wire n472_inv_n;
  wire n8086_o2_p;
  wire n8086_o2_n;
  wire n8093_o2_p;
  wire n8093_o2_n;
  wire G3752_o2_p;
  wire G3752_o2_n;
  wire n484_inv_p;
  wire n484_inv_n;
  wire n8199_o2_p;
  wire n8199_o2_n;
  wire n2800_lo_buf_o2_p;
  wire n2800_lo_buf_o2_n;
  wire G548_o2_p;
  wire G548_o2_n;
  wire n496_inv_p;
  wire n496_inv_n;
  wire G569_o2_p;
  wire G569_o2_n;
  wire G1761_o2_p;
  wire G1761_o2_n;
  wire n505_inv_p;
  wire n505_inv_n;
  wire G4101_o2_p;
  wire G4101_o2_n;
  wire G551_o2_p;
  wire G551_o2_n;
  wire n514_inv_p;
  wire n514_inv_n;
  wire G4743_o2_p;
  wire G4743_o2_n;
  wire G5271_o2_p;
  wire G5271_o2_n;
  wire G5790_o2_p;
  wire G5790_o2_n;
  wire G6122_o2_p;
  wire G6122_o2_n;
  wire G2082_o2_p;
  wire G2082_o2_n;
  wire n2812_lo_buf_o2_p;
  wire n2812_lo_buf_o2_n;
  wire n2668_lo_buf_o2_p;
  wire n2668_lo_buf_o2_n;
  wire n2680_lo_buf_o2_p;
  wire n2680_lo_buf_o2_n;
  wire G572_o2_p;
  wire G572_o2_n;
  wire G6125_o2_p;
  wire G6125_o2_n;
  wire n547_inv_p;
  wire n547_inv_n;
  wire n2656_lo_buf_o2_p;
  wire n2656_lo_buf_o2_n;
  wire G554_o2_p;
  wire G554_o2_n;
  wire G4452_o2_p;
  wire G4452_o2_n;
  wire n559_inv_p;
  wire n559_inv_n;
  wire n2644_lo_buf_o2_p;
  wire n2644_lo_buf_o2_n;
  wire G2410_o2_p;
  wire G2410_o2_n;
  wire n2632_lo_buf_o2_p;
  wire n2632_lo_buf_o2_n;
  wire n2620_lo_buf_o2_p;
  wire n2620_lo_buf_o2_n;
  wire G6131_o2_p;
  wire G6131_o2_n;
  wire G4693_o2_p;
  wire G4693_o2_n;
  wire G5209_o2_p;
  wire G5209_o2_n;
  wire G5741_o2_p;
  wire G5741_o2_n;
  wire G6082_o2_p;
  wire G6082_o2_n;
  wire G6119_o2_p;
  wire G6119_o2_n;
  wire n2608_lo_buf_o2_p;
  wire n2608_lo_buf_o2_n;
  wire n2596_lo_buf_o2_p;
  wire n2596_lo_buf_o2_n;
  wire n2584_lo_buf_o2_p;
  wire n2584_lo_buf_o2_n;
  wire n2572_lo_buf_o2_p;
  wire n2572_lo_buf_o2_n;
  wire n2704_lo_buf_o2_p;
  wire n2704_lo_buf_o2_n;
  wire G557_o2_p;
  wire G557_o2_n;
  wire G5936_o2_p;
  wire G5936_o2_n;
  wire G5442_o2_p;
  wire G5442_o2_n;
  wire G4926_o2_p;
  wire G4926_o2_n;
  wire G6134_o2_p;
  wire G6134_o2_n;
  wire G3929_o2_p;
  wire G3929_o2_n;
  wire G4425_o2_p;
  wire G4425_o2_n;
  wire G4947_o2_p;
  wire G4947_o2_n;
  wire n2764_lo_buf_o2_p;
  wire n2764_lo_buf_o2_n;
  wire n634_inv_p;
  wire n634_inv_n;
  wire n2560_lo_buf_o2_p;
  wire n2560_lo_buf_o2_n;
  wire n2824_lo_buf_o2_p;
  wire n2824_lo_buf_o2_n;
  wire G575_o2_p;
  wire G575_o2_n;
  wire G2740_o2_p;
  wire G2740_o2_n;
  wire n649_inv_p;
  wire n649_inv_n;
  wire n2548_lo_buf_o2_p;
  wire n2548_lo_buf_o2_n;
  wire n2536_lo_buf_o2_p;
  wire n2536_lo_buf_o2_n;
  wire n2524_lo_buf_o2_p;
  wire n2524_lo_buf_o2_n;
  wire G875_o2_p;
  wire G875_o2_n;
  wire G1064_o2_p;
  wire G1064_o2_n;
  wire G1253_o2_p;
  wire G1253_o2_n;
  wire G6140_o2_p;
  wire G6140_o2_n;
  wire G5151_o2_p;
  wire G5151_o2_n;
  wire G5686_o2_p;
  wire G5686_o2_n;
  wire G6061_o2_p;
  wire G6061_o2_n;
  wire G4803_o2_p;
  wire G4803_o2_n;
  wire G5332_o2_p;
  wire G5332_o2_n;
  wire G5844_o2_p;
  wire G5844_o2_n;
  wire G6114_o2_p;
  wire G6114_o2_n;
  wire G4806_o2_p;
  wire G4806_o2_n;
  wire G3881_o2_p;
  wire G3881_o2_n;
  wire G4370_o2_p;
  wire G4370_o2_n;
  wire G4896_o2_p;
  wire G4896_o2_n;
  wire G5001_o2_p;
  wire G5001_o2_n;
  wire G3121_o2_p;
  wire G3121_o2_n;
  wire n2512_lo_buf_o2_p;
  wire n2512_lo_buf_o2_n;
  wire G4085_o2_p;
  wire G4085_o2_n;
  wire G4605_o2_p;
  wire G4605_o2_n;
  wire G5118_o2_p;
  wire G5118_o2_n;
  wire G4997_o2_p;
  wire G4997_o2_n;
  wire n2500_lo_buf_o2_p;
  wire n2500_lo_buf_o2_n;
  wire n2716_lo_buf_o2_p;
  wire n2716_lo_buf_o2_n;
  wire G560_o2_p;
  wire G560_o2_n;
  wire G1895_o2_p;
  wire G1895_o2_n;
  wire G3064_o2_p;
  wire G3064_o2_n;
  wire G3269_o2_p;
  wire G3269_o2_n;
  wire G3569_o2_p;
  wire G3569_o2_n;
  wire n748_inv_p;
  wire n748_inv_n;
  wire G1196_o2_p;
  wire G1196_o2_n;
  wire G1007_o2_p;
  wire G1007_o2_n;
  wire G818_o2_p;
  wire G818_o2_n;
  wire G674_o2_p;
  wire G674_o2_n;
  wire G5041_o2_p;
  wire G5041_o2_n;
  wire G5562_o2_p;
  wire G5562_o2_n;
  wire G6005_o2_p;
  wire G6005_o2_n;
  wire G5214_o2_p;
  wire G5214_o2_n;
  wire G5746_o2_p;
  wire G5746_o2_n;
  wire G6087_o2_p;
  wire G6087_o2_n;
  wire G6086_o2_p;
  wire G6086_o2_n;
  wire G5745_o2_p;
  wire G5745_o2_n;
  wire G5213_o2_p;
  wire G5213_o2_n;
  wire G5893_o2_p;
  wire G5893_o2_n;
  wire G5391_o2_p;
  wire G5391_o2_n;
  wire G4864_o2_p;
  wire G4864_o2_n;
  wire G6143_o2_p;
  wire G6143_o2_n;
  wire G6008_o2_p;
  wire G6008_o2_n;
  wire G5565_o2_p;
  wire G5565_o2_n;
  wire G5044_o2_p;
  wire G5044_o2_n;
  wire G3813_o2_p;
  wire G3813_o2_n;
  wire G4325_o2_p;
  wire G4325_o2_n;
  wire G4834_o2_p;
  wire G4834_o2_n;
  wire G4993_o2_p;
  wire G4993_o2_n;
  wire G3989_o2_p;
  wire G3989_o2_n;
  wire G4490_o2_p;
  wire G4490_o2_n;
  wire G5011_o2_p;
  wire G5011_o2_n;
  wire G5112_o2_p;
  wire G5112_o2_n;
  wire n2776_lo_buf_o2_p;
  wire n2776_lo_buf_o2_n;
  wire G3298_o2_p;
  wire G3298_o2_n;
  wire G3073_o2_p;
  wire G3073_o2_n;
  wire G3265_o2_p;
  wire G3265_o2_n;
  wire G3624_o2_p;
  wire G3624_o2_n;
  wire G1642_o2_p;
  wire G1642_o2_n;
  wire G1980_o2_p;
  wire G1980_o2_n;
  wire n2488_lo_buf_o2_p;
  wire n2488_lo_buf_o2_n;
  wire G626_o2_p;
  wire G626_o2_n;
  wire G1139_o2_p;
  wire G1139_o2_n;
  wire G950_o2_p;
  wire G950_o2_n;
  wire G707_o2_p;
  wire G707_o2_n;
  wire G545_o2_p;
  wire G545_o2_n;
  wire G4217_o2_p;
  wire G4217_o2_n;
  wire G4716_o2_p;
  wire G4716_o2_n;
  wire G5244_o2_p;
  wire G5244_o2_n;
  wire G3136_o2_p;
  wire G3136_o2_n;
  wire G3499_o2_p;
  wire G3499_o2_n;
  wire G3885_o2_p;
  wire G3885_o2_n;
  wire G5243_o2_p;
  wire G5243_o2_n;
  wire G3886_o2_p;
  wire G3886_o2_n;
  wire G4375_o2_p;
  wire G4375_o2_n;
  wire G4901_o2_p;
  wire G4901_o2_n;
  wire G5054_o2_p;
  wire G5054_o2_n;
  wire G4374_o2_p;
  wire G4374_o2_n;
  wire G4900_o2_p;
  wire G4900_o2_n;
  wire G5053_o2_p;
  wire G5053_o2_n;
  wire G5242_o2_p;
  wire G5242_o2_n;
  wire G4034_o2_p;
  wire G4034_o2_n;
  wire G4556_o2_p;
  wire G4556_o2_n;
  wire G5064_o2_p;
  wire G5064_o2_n;
  wire G5172_o2_p;
  wire G5172_o2_n;
  wire G2030_o2_p;
  wire G2030_o2_n;
  wire G3016_o2_p;
  wire G3016_o2_n;
  wire G3520_o2_p;
  wire G3520_o2_n;
  wire G3261_o2_p;
  wire G3261_o2_n;
  wire G3620_o2_p;
  wire G3620_o2_n;
  wire G4220_o2_p;
  wire G4220_o2_n;
  wire G4719_o2_p;
  wire G4719_o2_n;
  wire G5247_o2_p;
  wire G5247_o2_n;
  wire G5109_o2_p;
  wire G5109_o2_n;
  wire G1638_o2_p;
  wire G1638_o2_n;
  wire G1976_o2_p;
  wire G1976_o2_n;
  wire G3560_o2_p;
  wire G3560_o2_n;
  wire G3205_o2_p;
  wire G3205_o2_n;
  wire G3193_o2_p;
  wire G3193_o2_n;
  wire G3367_o2_p;
  wire G3367_o2_n;
  wire G3670_o2_p;
  wire G3670_o2_n;
  wire n979_inv_p;
  wire n979_inv_n;
  wire G1280_o2_p;
  wire G1280_o2_n;
  wire G902_o2_p;
  wire G902_o2_n;
  wire G659_o2_p;
  wire G659_o2_n;
  wire G983_o2_p;
  wire G983_o2_n;
  wire G740_o2_p;
  wire G740_o2_n;
  wire G2917_o2_p;
  wire G2917_o2_n;
  wire G3391_o2_p;
  wire G3391_o2_n;
  wire G3494_o2_p;
  wire G3494_o2_n;
  wire G1512_o2_p;
  wire G1512_o2_n;
  wire G1854_o2_p;
  wire G1854_o2_n;
  wire G2203_o2_p;
  wire G2203_o2_n;
  wire G3493_o2_p;
  wire G3493_o2_n;
  wire G3069_o2_p;
  wire G3069_o2_n;
  wire G3574_o2_p;
  wire G3574_o2_n;
  wire G3319_o2_p;
  wire G3319_o2_n;
  wire G3667_o2_p;
  wire G3667_o2_n;
  wire G3068_o2_p;
  wire G3068_o2_n;
  wire G3573_o2_p;
  wire G3573_o2_n;
  wire G3666_o2_p;
  wire G3666_o2_n;
  wire G3318_o2_p;
  wire G3318_o2_n;
  wire G3492_o2_p;
  wire G3492_o2_n;
  wire G3241_o2_p;
  wire G3241_o2_n;
  wire G3722_o2_p;
  wire G3722_o2_n;
  wire G3422_o2_p;
  wire G3422_o2_n;
  wire G1445_o2_p;
  wire G1445_o2_n;
  wire G3257_o2_p;
  wire G3257_o2_n;
  wire G3616_o2_p;
  wire G3616_o2_n;
  wire G1634_o2_p;
  wire G1634_o2_n;
  wire G1972_o2_p;
  wire G1972_o2_n;
  wire G2256_o2_p;
  wire G2256_o2_n;
  wire G3394_o2_p;
  wire G3394_o2_n;
  wire G3557_o2_p;
  wire G3557_o2_n;
  wire G3364_o2_p;
  wire G3364_o2_n;
  wire G3719_o2_p;
  wire G3719_o2_n;
  wire G2253_o2_p;
  wire G2253_o2_n;
  wire G1583_o2_p;
  wire G1583_o2_n;
  wire G1917_o2_p;
  wire G1917_o2_n;
  wire G1727_o2_p;
  wire G1727_o2_n;
  wire G2061_o2_p;
  wire G2061_o2_n;
  wire G935_o2_p;
  wire G935_o2_n;
  wire G692_o2_p;
  wire G692_o2_n;
  wire G2136_o2_p;
  wire G2136_o2_n;
  wire G1507_o2_p;
  wire G1507_o2_n;
  wire G1849_o2_p;
  wire G1849_o2_n;
  wire G2198_o2_p;
  wire G2198_o2_n;
  wire G2197_o2_p;
  wire G2197_o2_n;
  wire G1848_o2_p;
  wire G1848_o2_n;
  wire G1689_o2_p;
  wire G1689_o2_n;
  wire G2016_o2_p;
  wire G2016_o2_n;
  wire G2314_o2_p;
  wire G2314_o2_n;
  wire G2313_o2_p;
  wire G2313_o2_n;
  wire G1688_o2_p;
  wire G1688_o2_n;
  wire G2015_o2_p;
  wire G2015_o2_n;
  wire G1847_o2_p;
  wire G1847_o2_n;
  wire G2196_o2_p;
  wire G2196_o2_n;
  wire G2118_o2_p;
  wire G2118_o2_n;
  wire G1777_o2_p;
  wire G1777_o2_n;
  wire G1630_o2_p;
  wire G1630_o2_n;
  wire G1968_o2_p;
  wire G1968_o2_n;
  wire G2309_o2_p;
  wire G2309_o2_n;
  wire G2139_o2_p;
  wire G2139_o2_n;
  wire G1580_o2_p;
  wire G1580_o2_n;
  wire G2250_o2_p;
  wire G2250_o2_n;
  wire G1914_o2_p;
  wire G1914_o2_n;
  wire G1724_o2_p;
  wire G1724_o2_n;
  wire G2058_o2_p;
  wire G2058_o2_n;
  wire n2728_lo_buf_o2_p;
  wire n2728_lo_buf_o2_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire g686_p;
  wire g686_n;
  wire g687_p;
  wire g687_n;
  wire g688_p;
  wire g688_n;
  wire g689_p;
  wire g689_n;
  wire g690_p;
  wire g690_n;
  wire g691_p;
  wire g691_n;
  wire g692_p;
  wire g692_n;
  wire g693_p;
  wire g693_n;
  wire g694_p;
  wire g694_n;
  wire g695_p;
  wire g695_n;
  wire g696_p;
  wire g696_n;
  wire g697_p;
  wire g697_n;
  wire g698_p;
  wire g698_n;
  wire g699_p;
  wire g699_n;
  wire g700_p;
  wire g700_n;
  wire g701_p;
  wire g701_n;
  wire g702_p;
  wire g702_n;
  wire g703_p;
  wire g703_n;
  wire g704_p;
  wire g704_n;
  wire g705_p;
  wire g705_n;
  wire g706_p;
  wire g706_n;
  wire g707_p;
  wire g707_n;
  wire g708_p;
  wire g708_n;
  wire g709_p;
  wire g709_n;
  wire g710_p;
  wire g710_n;
  wire g711_p;
  wire g711_n;
  wire g712_p;
  wire g712_n;
  wire g713_p;
  wire g713_n;
  wire g714_p;
  wire g714_n;
  wire g715_p;
  wire g715_n;
  wire g716_p;
  wire g716_n;
  wire g717_p;
  wire g717_n;
  wire g718_p;
  wire g718_n;
  wire g719_p;
  wire g719_n;
  wire g720_p;
  wire g720_n;
  wire g721_p;
  wire g721_n;
  wire g722_p;
  wire g722_n;
  wire g723_p;
  wire g723_n;
  wire g724_p;
  wire g724_n;
  wire g725_p;
  wire g725_n;
  wire g726_p;
  wire g726_n;
  wire g727_p;
  wire g727_n;
  wire g728_p;
  wire g728_n;
  wire g729_p;
  wire g729_n;
  wire g730_p;
  wire g730_n;
  wire g731_p;
  wire g731_n;
  wire g732_p;
  wire g732_n;
  wire g733_p;
  wire g733_n;
  wire g734_p;
  wire g734_n;
  wire g735_p;
  wire g735_n;
  wire g736_p;
  wire g736_n;
  wire g737_p;
  wire g737_n;
  wire g738_p;
  wire g738_n;
  wire g739_p;
  wire g739_n;
  wire g740_p;
  wire g740_n;
  wire g741_p;
  wire g741_n;
  wire g742_p;
  wire g742_n;
  wire g743_p;
  wire g743_n;
  wire g744_p;
  wire g744_n;
  wire g745_p;
  wire g745_n;
  wire g746_p;
  wire g746_n;
  wire g747_p;
  wire g747_n;
  wire g748_p;
  wire g748_n;
  wire g749_p;
  wire g749_n;
  wire g750_p;
  wire g750_n;
  wire g751_p;
  wire g751_n;
  wire g752_p;
  wire g752_n;
  wire g753_p;
  wire g753_n;
  wire g754_p;
  wire g754_n;
  wire g755_p;
  wire g755_n;
  wire g756_p;
  wire g756_n;
  wire g757_p;
  wire g757_n;
  wire g758_p;
  wire g758_n;
  wire g759_p;
  wire g759_n;
  wire g760_p;
  wire g760_n;
  wire g761_p;
  wire g761_n;
  wire g762_p;
  wire g762_n;
  wire g763_p;
  wire g763_n;
  wire g764_p;
  wire g764_n;
  wire g765_p;
  wire g765_n;
  wire g766_p;
  wire g766_n;
  wire g767_p;
  wire g767_n;
  wire g768_p;
  wire g768_n;
  wire g769_p;
  wire g769_n;
  wire g770_p;
  wire g770_n;
  wire g771_p;
  wire g771_n;
  wire g772_p;
  wire g772_n;
  wire g773_p;
  wire g773_n;
  wire g774_p;
  wire g774_n;
  wire g775_p;
  wire g775_n;
  wire g776_p;
  wire g776_n;
  wire g777_p;
  wire g777_n;
  wire g778_p;
  wire g778_n;
  wire g779_p;
  wire g779_n;
  wire g780_p;
  wire g780_n;
  wire g781_p;
  wire g781_n;
  wire g782_p;
  wire g782_n;
  wire g783_p;
  wire g783_n;
  wire g784_p;
  wire g784_n;
  wire g785_p;
  wire g785_n;
  wire g786_p;
  wire g786_n;
  wire g787_p;
  wire g787_n;
  wire g788_p;
  wire g788_n;
  wire g789_p;
  wire g789_n;
  wire g790_p;
  wire g790_n;
  wire g791_p;
  wire g791_n;
  wire g792_p;
  wire g792_n;
  wire g793_p;
  wire g793_n;
  wire g794_p;
  wire g794_n;
  wire g795_p;
  wire g795_n;
  wire g796_p;
  wire g796_n;
  wire g797_p;
  wire g797_n;
  wire g798_p;
  wire g798_n;
  wire g799_p;
  wire g799_n;
  wire g800_p;
  wire g800_n;
  wire g801_p;
  wire g801_n;
  wire g802_p;
  wire g802_n;
  wire g803_p;
  wire g803_n;
  wire g804_p;
  wire g804_n;
  wire g805_p;
  wire g805_n;
  wire g806_p;
  wire g806_n;
  wire g807_p;
  wire g807_n;
  wire g808_p;
  wire g808_n;
  wire g809_p;
  wire g809_n;
  wire g810_p;
  wire g810_n;
  wire g811_p;
  wire g811_n;
  wire g812_p;
  wire g812_n;
  wire g813_p;
  wire g813_n;
  wire g814_p;
  wire g814_n;
  wire g815_p;
  wire g815_n;
  wire g816_p;
  wire g816_n;
  wire g817_p;
  wire g817_n;
  wire g818_p;
  wire g818_n;
  wire g819_p;
  wire g819_n;
  wire g820_p;
  wire g820_n;
  wire g821_p;
  wire g821_n;
  wire g822_p;
  wire g822_n;
  wire g823_p;
  wire g823_n;
  wire g824_p;
  wire g824_n;
  wire g825_p;
  wire g825_n;
  wire g826_p;
  wire g826_n;
  wire g827_p;
  wire g827_n;
  wire g828_p;
  wire g828_n;
  wire g829_p;
  wire g829_n;
  wire g830_p;
  wire g830_n;
  wire g831_p;
  wire g831_n;
  wire g832_p;
  wire g832_n;
  wire g833_p;
  wire g833_n;
  wire g834_p;
  wire g834_n;
  wire g835_p;
  wire g835_n;
  wire g836_p;
  wire g836_n;
  wire g837_p;
  wire g837_n;
  wire g838_p;
  wire g838_n;
  wire g839_p;
  wire g839_n;
  wire g840_p;
  wire g840_n;
  wire g841_p;
  wire g841_n;
  wire g842_p;
  wire g842_n;
  wire g843_p;
  wire g843_n;
  wire g844_p;
  wire g844_n;
  wire g845_p;
  wire g845_n;
  wire g846_p;
  wire g846_n;
  wire g847_p;
  wire g847_n;
  wire g848_p;
  wire g848_n;
  wire g849_p;
  wire g849_n;
  wire g850_p;
  wire g850_n;
  wire g851_p;
  wire g851_n;
  wire g852_p;
  wire g852_n;
  wire g853_p;
  wire g853_n;
  wire g854_p;
  wire g854_n;
  wire g855_p;
  wire g855_n;
  wire g856_p;
  wire g856_n;
  wire g857_p;
  wire g857_n;
  wire g858_p;
  wire g858_n;
  wire g859_p;
  wire g859_n;
  wire g860_p;
  wire g860_n;
  wire g861_p;
  wire g861_n;
  wire g862_p;
  wire g862_n;
  wire g863_p;
  wire g863_n;
  wire g864_p;
  wire g864_n;
  wire g865_p;
  wire g865_n;
  wire g866_p;
  wire g866_n;
  wire g867_p;
  wire g867_n;
  wire g868_p;
  wire g868_n;
  wire g869_p;
  wire g869_n;
  wire g870_p;
  wire g870_n;
  wire g871_p;
  wire g871_n;
  wire g872_p;
  wire g872_n;
  wire g873_p;
  wire g873_n;
  wire g874_p;
  wire g874_n;
  wire g875_p;
  wire g875_n;
  wire g876_p;
  wire g876_n;
  wire g877_p;
  wire g877_n;
  wire g878_p;
  wire g878_n;
  wire g879_p;
  wire g879_n;
  wire g880_p;
  wire g880_n;
  wire g881_p;
  wire g881_n;
  wire g882_p;
  wire g882_n;
  wire g883_p;
  wire g883_n;
  wire g884_p;
  wire g884_n;
  wire g885_p;
  wire g885_n;
  wire g886_p;
  wire g886_n;
  wire g887_p;
  wire g887_n;
  wire g888_p;
  wire g888_n;
  wire g889_p;
  wire g889_n;
  wire g890_p;
  wire g890_n;
  wire g891_p;
  wire g891_n;
  wire g892_p;
  wire g892_n;
  wire g893_p;
  wire g893_n;
  wire g894_p;
  wire g894_n;
  wire g895_p;
  wire g895_n;
  wire g896_p;
  wire g896_n;
  wire g897_p;
  wire g897_n;
  wire g898_p;
  wire g898_n;
  wire g899_p;
  wire g899_n;
  wire g900_p;
  wire g900_n;
  wire g901_p;
  wire g901_n;
  wire g902_p;
  wire g902_n;
  wire g903_p;
  wire g903_n;
  wire g904_p;
  wire g904_n;
  wire g905_p;
  wire g905_n;
  wire g906_p;
  wire g906_n;
  wire g907_p;
  wire g907_n;
  wire g908_p;
  wire g908_n;
  wire g909_p;
  wire g909_n;
  wire g910_p;
  wire g910_n;
  wire g911_p;
  wire g911_n;
  wire g912_p;
  wire g912_n;
  wire g913_p;
  wire g913_n;
  wire g914_p;
  wire g914_n;
  wire g915_p;
  wire g915_n;
  wire g916_p;
  wire g916_n;
  wire g917_p;
  wire g917_n;
  wire g918_p;
  wire g918_n;
  wire g919_p;
  wire g919_n;
  wire g920_p;
  wire g920_n;
  wire g921_p;
  wire g921_n;
  wire g922_p;
  wire g922_n;
  wire g923_p;
  wire g923_n;
  wire g924_p;
  wire g924_n;
  wire g925_p;
  wire g925_n;
  wire g926_p;
  wire g926_n;
  wire g927_p;
  wire g927_n;
  wire g928_p;
  wire g928_n;
  wire g929_p;
  wire g929_n;
  wire g930_p;
  wire g930_n;
  wire g931_p;
  wire g931_n;
  wire g932_p;
  wire g932_n;
  wire g933_p;
  wire g933_n;
  wire g934_p;
  wire g934_n;
  wire g935_p;
  wire g935_n;
  wire g936_p;
  wire g936_n;
  wire g937_p;
  wire g937_n;
  wire g938_p;
  wire g938_n;
  wire g939_p;
  wire g939_n;
  wire g940_p;
  wire g940_n;
  wire g941_p;
  wire g941_n;
  wire g942_p;
  wire g942_n;
  wire g943_p;
  wire g943_n;
  wire g944_p;
  wire g944_n;
  wire g945_p;
  wire g945_n;
  wire g946_p;
  wire g946_n;
  wire g947_p;
  wire g947_n;
  wire g948_p;
  wire g948_n;
  wire g949_p;
  wire g949_n;
  wire g950_p;
  wire g950_n;
  wire g951_p;
  wire g951_n;
  wire g952_p;
  wire g952_n;
  wire g953_p;
  wire g953_n;
  wire g954_p;
  wire g954_n;
  wire g955_p;
  wire g955_n;
  wire g956_p;
  wire g956_n;
  wire g957_p;
  wire g957_n;
  wire g958_p;
  wire g958_n;
  wire g959_p;
  wire g959_n;
  wire g960_p;
  wire g960_n;
  wire g961_p;
  wire g961_n;
  wire g962_p;
  wire g962_n;
  wire g963_p;
  wire g963_n;
  wire g964_p;
  wire g964_n;
  wire g965_p;
  wire g965_n;
  wire g966_p;
  wire g966_n;
  wire g967_p;
  wire g967_n;
  wire g968_p;
  wire g968_n;
  wire g969_p;
  wire g969_n;
  wire g970_p;
  wire g970_n;
  wire g971_p;
  wire g971_n;
  wire g972_p;
  wire g972_n;
  wire g973_p;
  wire g973_n;
  wire g974_p;
  wire g974_n;
  wire g975_p;
  wire g975_n;
  wire g976_p;
  wire g976_n;
  wire g977_p;
  wire g977_n;
  wire g978_p;
  wire g978_n;
  wire g979_p;
  wire g979_n;
  wire g980_p;
  wire g980_n;
  wire g981_p;
  wire g981_n;
  wire g982_p;
  wire g982_n;
  wire g983_p;
  wire g983_n;
  wire g984_p;
  wire g984_n;
  wire g985_p;
  wire g985_n;
  wire g986_p;
  wire g986_n;
  wire g987_p;
  wire g987_n;
  wire g988_p;
  wire g988_n;
  wire g989_p;
  wire g989_n;
  wire g990_p;
  wire g990_n;
  wire g991_p;
  wire g991_n;
  wire g992_p;
  wire g992_n;
  wire g993_p;
  wire g993_n;
  wire g994_p;
  wire g994_n;
  wire g995_p;
  wire g995_n;
  wire g996_p;
  wire g996_n;
  wire g997_p;
  wire g997_n;
  wire g998_p;
  wire g998_n;
  wire g999_p;
  wire g999_n;
  wire g1000_p;
  wire g1000_n;
  wire g1001_p;
  wire g1001_n;
  wire g1002_p;
  wire g1002_n;
  wire g1003_p;
  wire g1003_n;
  wire g1004_p;
  wire g1004_n;
  wire g1005_p;
  wire g1005_n;
  wire g1006_p;
  wire g1006_n;
  wire g1007_p;
  wire g1007_n;
  wire g1008_p;
  wire g1008_n;
  wire g1009_p;
  wire g1009_n;
  wire g1010_p;
  wire g1010_n;
  wire g1011_p;
  wire g1011_n;
  wire g1012_p;
  wire g1012_n;
  wire g1013_p;
  wire g1013_n;
  wire g1014_p;
  wire g1014_n;
  wire g1015_p;
  wire g1015_n;
  wire g1016_p;
  wire g1016_n;
  wire g1017_p;
  wire g1017_n;
  wire g1018_p;
  wire g1018_n;
  wire g1019_p;
  wire g1019_n;
  wire g1020_p;
  wire g1020_n;
  wire g1021_p;
  wire g1021_n;
  wire g1022_p;
  wire g1022_n;
  wire g1023_p;
  wire g1023_n;
  wire g1024_p;
  wire g1024_n;
  wire g1025_p;
  wire g1025_n;
  wire g1026_p;
  wire g1026_n;
  wire g1027_p;
  wire g1027_n;
  wire g1028_p;
  wire g1028_n;
  wire g1029_p;
  wire g1029_n;
  wire g1030_p;
  wire g1030_n;
  wire g1031_p;
  wire g1031_n;
  wire g1032_p;
  wire g1032_n;
  wire g1033_p;
  wire g1033_n;
  wire g1034_p;
  wire g1034_n;
  wire g1035_p;
  wire g1035_n;
  wire g1036_p;
  wire g1036_n;
  wire g1037_p;
  wire g1037_n;
  wire g1038_p;
  wire g1038_n;
  wire g1039_p;
  wire g1039_n;
  wire g1040_p;
  wire g1040_n;
  wire g1041_p;
  wire g1041_n;
  wire g1042_p;
  wire g1042_n;
  wire g1043_p;
  wire g1043_n;
  wire g1044_p;
  wire g1044_n;
  wire g1045_p;
  wire g1045_n;
  wire g1046_p;
  wire g1046_n;
  wire g1047_p;
  wire g1047_n;
  wire g1048_p;
  wire g1048_n;
  wire g1049_p;
  wire g1049_n;
  wire g1050_p;
  wire g1050_n;
  wire g1051_p;
  wire g1051_n;
  wire g1052_p;
  wire g1052_n;
  wire g1053_p;
  wire g1053_n;
  wire g1054_p;
  wire g1054_n;
  wire g1055_p;
  wire g1055_n;
  wire g1056_p;
  wire g1056_n;
  wire g1057_p;
  wire g1057_n;
  wire g1058_p;
  wire g1058_n;
  wire g1059_p;
  wire g1059_n;
  wire g1060_p;
  wire g1060_n;
  wire g1061_p;
  wire g1061_n;
  wire g1062_p;
  wire g1062_n;
  wire g1063_p;
  wire g1063_n;
  wire g1064_p;
  wire g1064_n;
  wire g1065_p;
  wire g1065_n;
  wire g1066_p;
  wire g1066_n;
  wire g1067_p;
  wire g1067_n;
  wire g1068_p;
  wire g1068_n;
  wire g1069_p;
  wire g1069_n;
  wire g1070_p;
  wire g1070_n;
  wire g1071_p;
  wire g1071_n;
  wire g1072_p;
  wire g1072_n;
  wire g1073_p;
  wire g1073_n;
  wire g1074_p;
  wire g1074_n;
  wire g1075_p;
  wire g1075_n;
  wire g1076_p;
  wire g1076_n;
  wire g1077_p;
  wire g1077_n;
  wire g1078_p;
  wire g1078_n;
  wire g1079_p;
  wire g1079_n;
  wire g1080_p;
  wire g1080_n;
  wire g1081_p;
  wire g1081_n;
  wire g1082_p;
  wire g1082_n;
  wire g1083_p;
  wire g1083_n;
  wire g1084_p;
  wire g1084_n;
  wire g1085_p;
  wire g1085_n;
  wire g1086_p;
  wire g1086_n;
  wire g1087_p;
  wire g1087_n;
  wire g1088_p;
  wire g1088_n;
  wire g1089_p;
  wire g1089_n;
  wire g1090_p;
  wire g1090_n;
  wire g1091_p;
  wire g1091_n;
  wire g1092_p;
  wire g1092_n;
  wire g1093_p;
  wire g1093_n;
  wire g1094_p;
  wire g1094_n;
  wire g1095_p;
  wire g1095_n;
  wire g1096_p;
  wire g1096_n;
  wire g1097_p;
  wire g1097_n;
  wire g1098_p;
  wire g1098_n;
  wire g1099_p;
  wire g1099_n;
  wire g1100_p;
  wire g1100_n;
  wire g1101_p;
  wire g1101_n;
  wire g1102_p;
  wire g1102_n;
  wire g1103_p;
  wire g1103_n;
  wire g1104_p;
  wire g1104_n;
  wire g1105_p;
  wire g1105_n;
  wire g1106_p;
  wire g1106_n;
  wire g1107_p;
  wire g1107_n;
  wire g1108_p;
  wire g1108_n;
  wire g1109_p;
  wire g1109_n;
  wire g1110_p;
  wire g1110_n;
  wire g1111_p;
  wire g1111_n;
  wire g1112_p;
  wire g1112_n;
  wire g1113_p;
  wire g1113_n;
  wire g1114_p;
  wire g1114_n;
  wire g1115_p;
  wire g1115_n;
  wire g1116_p;
  wire g1116_n;
  wire g1117_p;
  wire g1117_n;
  wire g1118_p;
  wire g1118_n;
  wire g1119_p;
  wire g1119_n;
  wire g1120_p;
  wire g1120_n;
  wire g1121_p;
  wire g1121_n;
  wire g1122_p;
  wire g1122_n;
  wire g1123_p;
  wire g1123_n;
  wire g1124_p;
  wire g1124_n;
  wire g1125_p;
  wire g1125_n;
  wire g1126_p;
  wire g1126_n;
  wire g1127_p;
  wire g1127_n;
  wire g1128_p;
  wire g1128_n;
  wire g1129_p;
  wire g1129_n;
  wire g1130_p;
  wire g1130_n;
  wire g1131_p;
  wire g1131_n;
  wire g1132_p;
  wire g1132_n;
  wire g1133_p;
  wire g1133_n;
  wire g1134_p;
  wire g1134_n;
  wire g1135_p;
  wire g1135_n;
  wire g1136_p;
  wire g1136_n;
  wire g1137_p;
  wire g1137_n;
  wire g1138_p;
  wire g1138_n;
  wire g1139_p;
  wire g1139_n;
  wire g1140_p;
  wire g1140_n;
  wire g1141_p;
  wire g1141_n;
  wire g1142_p;
  wire g1142_n;
  wire g1143_p;
  wire g1143_n;
  wire g1144_p;
  wire g1144_n;
  wire g1145_p;
  wire g1145_n;
  wire g1146_p;
  wire g1146_n;
  wire g1147_p;
  wire g1147_n;
  wire g1148_p;
  wire g1148_n;
  wire g1149_p;
  wire g1149_n;
  wire g1150_p;
  wire g1150_n;
  wire g1151_p;
  wire g1151_n;
  wire g1152_p;
  wire g1152_n;
  wire g1153_p;
  wire g1153_n;
  wire g1154_p;
  wire g1154_n;
  wire g1155_p;
  wire g1155_n;
  wire g1156_p;
  wire g1156_n;
  wire g1157_p;
  wire g1157_n;
  wire g1158_p;
  wire g1158_n;
  wire g1159_p;
  wire g1159_n;
  wire g1160_p;
  wire g1160_n;
  wire g1161_p;
  wire g1161_n;
  wire g1162_p;
  wire g1162_n;
  wire g1163_p;
  wire g1163_n;
  wire g1164_p;
  wire g1164_n;
  wire g1165_p;
  wire g1165_n;
  wire g1166_p;
  wire g1166_n;
  wire g1167_p;
  wire g1167_n;
  wire g1168_p;
  wire g1168_n;
  wire g1169_p;
  wire g1169_n;
  wire g1170_p;
  wire g1170_n;
  wire g1171_p;
  wire g1171_n;
  wire g1172_p;
  wire g1172_n;
  wire g1173_p;
  wire g1173_n;
  wire g1174_p;
  wire g1174_n;
  wire g1175_p;
  wire g1175_n;
  wire g1176_p;
  wire g1176_n;
  wire g1177_p;
  wire g1177_n;
  wire g1178_p;
  wire g1178_n;
  wire g1179_p;
  wire g1179_n;
  wire g1180_p;
  wire g1180_n;
  wire g1181_p;
  wire g1181_n;
  wire g1182_p;
  wire g1182_n;
  wire g1183_p;
  wire g1183_n;
  wire g1184_p;
  wire g1184_n;
  wire g1185_p;
  wire g1185_n;
  wire g1186_p;
  wire g1186_n;
  wire g1187_p;
  wire g1187_n;
  wire g1188_p;
  wire g1188_n;
  wire g1189_p;
  wire g1189_n;
  wire g1190_p;
  wire g1190_n;
  wire g1191_p;
  wire g1191_n;
  wire g1192_p;
  wire g1192_n;
  wire g1193_p;
  wire g1193_n;
  wire g1194_p;
  wire g1194_n;
  wire g1195_p;
  wire g1195_n;
  wire g1196_p;
  wire g1196_n;
  wire g1197_p;
  wire g1197_n;
  wire g1198_p;
  wire g1198_n;
  wire g1199_p;
  wire g1199_n;
  wire g1200_p;
  wire g1200_n;
  wire g1201_p;
  wire g1201_n;
  wire g1202_p;
  wire g1202_n;
  wire g1203_p;
  wire g1203_n;
  wire g1204_p;
  wire g1204_n;
  wire g1205_p;
  wire g1205_n;
  wire g1206_p;
  wire g1206_n;
  wire g1207_p;
  wire g1207_n;
  wire g1208_p;
  wire g1208_n;
  wire g1209_p;
  wire g1209_n;
  wire g1210_p;
  wire g1210_n;
  wire g1211_p;
  wire g1211_n;
  wire g1212_p;
  wire g1212_n;
  wire g1213_p;
  wire g1213_n;
  wire g1214_p;
  wire g1214_n;
  wire g1215_p;
  wire g1215_n;
  wire g1216_p;
  wire g1216_n;
  wire g1217_p;
  wire g1217_n;
  wire g1218_p;
  wire g1218_n;
  wire g1219_p;
  wire g1219_n;
  wire g1220_p;
  wire g1220_n;
  wire g1221_p;
  wire g1221_n;
  wire g1222_p;
  wire g1222_n;
  wire g1223_p;
  wire g1223_n;
  wire g1224_p;
  wire g1224_n;
  wire g1225_p;
  wire g1225_n;
  wire g1226_p;
  wire g1226_n;
  wire g1227_p;
  wire g1227_n;
  wire g1228_p;
  wire g1228_n;
  wire g1229_p;
  wire g1229_n;
  wire g1230_p;
  wire g1230_n;
  wire g1231_p;
  wire g1231_n;
  wire g1232_p;
  wire g1232_n;
  wire g1233_p;
  wire g1233_n;
  wire g1234_p;
  wire g1234_n;
  wire g1235_p;
  wire g1235_n;
  wire g1236_p;
  wire g1236_n;
  wire g1237_p;
  wire g1237_n;
  wire g1238_p;
  wire g1238_n;
  wire g1239_p;
  wire g1239_n;
  wire g1240_p;
  wire g1240_n;
  wire g1241_p;
  wire g1241_n;
  wire g1242_p;
  wire g1242_n;
  wire g1243_p;
  wire g1243_n;
  wire g1244_p;
  wire g1244_n;
  wire g1245_p;
  wire g1245_n;
  wire g1246_p;
  wire g1246_n;
  wire g1247_p;
  wire g1247_n;
  wire g1248_p;
  wire g1248_n;
  wire g1249_p;
  wire g1249_n;
  wire g1250_p;
  wire g1250_n;
  wire g1251_p;
  wire g1251_n;
  wire g1252_p;
  wire g1252_n;
  wire g1253_p;
  wire g1253_n;
  wire g1254_p;
  wire g1254_n;
  wire g1255_p;
  wire g1255_n;
  wire g1256_p;
  wire g1256_n;
  wire g1257_p;
  wire g1257_n;
  wire g1258_p;
  wire g1258_n;
  wire g1259_p;
  wire g1259_n;
  wire g1260_p;
  wire g1260_n;
  wire g1261_p;
  wire g1261_n;
  wire g1262_p;
  wire g1262_n;
  wire g1263_p;
  wire g1263_n;
  wire g1264_p;
  wire g1264_n;
  wire g1265_p;
  wire g1265_n;
  wire g1266_p;
  wire g1266_n;
  wire g1267_p;
  wire g1267_n;
  wire g1268_p;
  wire g1268_n;
  wire g1269_p;
  wire g1269_n;
  wire g1270_p;
  wire g1270_n;
  wire g1271_p;
  wire g1271_n;
  wire g1272_p;
  wire g1272_n;
  wire g1273_p;
  wire g1273_n;
  wire g1274_p;
  wire g1274_n;
  wire g1275_p;
  wire g1275_n;
  wire g1276_p;
  wire g1276_n;
  wire g1277_p;
  wire g1277_n;
  wire g1278_p;
  wire g1278_n;
  wire g1279_p;
  wire g1279_n;
  wire g1280_p;
  wire g1280_n;
  wire g1281_p;
  wire g1281_n;
  wire g1282_p;
  wire g1282_n;
  wire g1283_p;
  wire g1283_n;
  wire g1284_p;
  wire g1284_n;
  wire g1285_p;
  wire g1285_n;
  wire g1286_p;
  wire g1286_n;
  wire g1287_p;
  wire g1287_n;
  wire g1288_p;
  wire g1288_n;
  wire g1289_p;
  wire g1289_n;
  wire g1290_p;
  wire g1290_n;
  wire g1291_p;
  wire g1291_n;
  wire g1292_p;
  wire g1292_n;
  wire g1293_p;
  wire g1293_n;
  wire g1294_p;
  wire g1294_n;
  wire g1295_p;
  wire g1295_n;
  wire g1296_p;
  wire g1296_n;
  wire g1297_p;
  wire g1297_n;
  wire g1298_p;
  wire g1298_n;
  wire g1299_p;
  wire g1299_n;
  wire g1300_p;
  wire g1300_n;
  wire g1301_p;
  wire g1301_n;
  wire g1302_p;
  wire g1302_n;
  wire g1303_p;
  wire g1303_n;
  wire g1304_p;
  wire g1304_n;
  wire g1305_p;
  wire g1305_n;
  wire g1306_p;
  wire g1306_n;
  wire g1307_p;
  wire g1307_n;
  wire g1308_p;
  wire g1308_n;
  wire g1309_p;
  wire g1309_n;
  wire g1310_p;
  wire g1310_n;
  wire g1311_p;
  wire g1311_n;
  wire g1312_p;
  wire g1312_n;
  wire g1313_p;
  wire g1313_n;
  wire g1314_p;
  wire g1314_n;
  wire g1315_p;
  wire g1315_n;
  wire g1316_p;
  wire g1316_n;
  wire g1317_p;
  wire g1317_n;
  wire g1318_p;
  wire g1318_n;
  wire g1319_p;
  wire g1319_n;
  wire g1320_p;
  wire g1320_n;
  wire g1321_p;
  wire g1321_n;
  wire g1322_p;
  wire g1322_n;
  wire g1323_p;
  wire g1323_n;
  wire g1324_p;
  wire g1324_n;
  wire g1325_p;
  wire g1325_n;
  wire g1326_p;
  wire g1326_n;
  wire g1327_p;
  wire g1327_n;
  wire g1328_p;
  wire g1328_n;
  wire g1329_p;
  wire g1329_n;
  wire g1330_p;
  wire g1330_n;
  wire g1331_p;
  wire g1331_n;
  wire g1332_p;
  wire g1332_n;
  wire g1333_p;
  wire g1333_n;
  wire g1334_p;
  wire g1334_n;
  wire g1335_p;
  wire g1335_n;
  wire g1336_p;
  wire g1336_n;
  wire g1337_p;
  wire g1337_n;
  wire g1338_p;
  wire g1338_n;
  wire g1339_p;
  wire g1339_n;
  wire g1340_p;
  wire g1340_n;
  wire g1341_p;
  wire g1341_n;
  wire g1342_p;
  wire g1342_n;
  wire g1343_p;
  wire g1343_n;
  wire g1344_p;
  wire g1344_n;
  wire g1345_p;
  wire g1345_n;
  wire g1346_p;
  wire g1346_n;
  wire g1347_p;
  wire g1347_n;
  wire g1348_p;
  wire g1348_n;
  wire g1349_p;
  wire g1349_n;
  wire g1350_p;
  wire g1350_n;
  wire g1351_p;
  wire g1351_n;
  wire g1352_p;
  wire g1352_n;
  wire g1353_p;
  wire g1353_n;
  wire g1354_p;
  wire g1354_n;
  wire g1355_p;
  wire g1355_n;
  wire g1356_p;
  wire g1356_n;
  wire g1357_p;
  wire g1357_n;
  wire g1358_p;
  wire g1358_n;
  wire g1359_p;
  wire g1359_n;
  wire g1360_p;
  wire g1360_n;
  wire g1361_p;
  wire g1361_n;
  wire g1362_p;
  wire g1362_n;
  wire g1363_p;
  wire g1363_n;
  wire g1364_p;
  wire g1364_n;
  wire g1365_p;
  wire g1365_n;
  wire g1366_p;
  wire g1366_n;
  wire g1367_p;
  wire g1367_n;
  wire g1368_p;
  wire g1368_n;
  wire g1369_p;
  wire g1369_n;
  wire g1370_p;
  wire g1370_n;
  wire g1371_p;
  wire g1371_n;
  wire g1372_p;
  wire g1372_n;
  wire g1373_p;
  wire g1373_n;
  wire g1374_p;
  wire g1374_n;
  wire g1375_p;
  wire g1375_n;
  wire g1376_p;
  wire g1376_n;
  wire g1377_p;
  wire g1377_n;
  wire g1378_p;
  wire g1378_n;
  wire g1379_p;
  wire g1379_n;
  wire g1380_p;
  wire g1380_n;
  wire g1381_p;
  wire g1381_n;
  wire g1382_p;
  wire g1382_n;
  wire g1383_p;
  wire g1383_n;
  wire g1384_p;
  wire g1384_n;
  wire g1385_p;
  wire g1385_n;
  wire g1386_p;
  wire g1386_n;
  wire g1387_p;
  wire g1387_n;
  wire g1388_p;
  wire g1388_n;
  wire g1389_p;
  wire g1389_n;
  wire g1390_p;
  wire g1390_n;
  wire g1391_p;
  wire g1391_n;
  wire g1392_p;
  wire g1392_n;
  wire g1393_p;
  wire g1393_n;
  wire g1394_p;
  wire g1394_n;
  wire g1395_p;
  wire g1395_n;
  wire g1396_p;
  wire g1396_n;
  wire g1397_p;
  wire g1397_n;
  wire g1398_p;
  wire g1398_n;
  wire g1399_p;
  wire g1399_n;
  wire g1400_p;
  wire g1400_n;
  wire g1401_p;
  wire g1401_n;
  wire g1402_p;
  wire g1402_n;
  wire g1403_p;
  wire g1403_n;
  wire g1404_p;
  wire g1404_n;
  wire g1405_p;
  wire g1405_n;
  wire g1406_p;
  wire g1406_n;
  wire g1407_p;
  wire g1407_n;
  wire g1408_p;
  wire g1408_n;
  wire g1409_p;
  wire g1409_n;
  wire g1410_p;
  wire g1410_n;
  wire g1411_p;
  wire g1411_n;
  wire g1412_p;
  wire g1412_n;
  wire g1413_p;
  wire g1413_n;
  wire g1414_p;
  wire g1414_n;
  wire g1415_p;
  wire g1415_n;
  wire g1416_p;
  wire g1416_n;
  wire g1417_p;
  wire g1417_n;
  wire g1418_p;
  wire g1418_n;
  wire g1419_p;
  wire g1419_n;
  wire g1420_p;
  wire g1420_n;
  wire g1421_p;
  wire g1421_n;
  wire g1422_p;
  wire g1422_n;
  wire g1423_p;
  wire g1423_n;
  wire g1424_p;
  wire g1424_n;
  wire g1425_p;
  wire g1425_n;
  wire g1426_p;
  wire g1426_n;
  wire g1427_p;
  wire g1427_n;
  wire g1428_p;
  wire g1428_n;
  wire g1429_p;
  wire g1429_n;
  wire g1430_p;
  wire g1430_n;
  wire g1431_p;
  wire g1431_n;
  wire g1432_p;
  wire g1432_n;
  wire g1433_p;
  wire g1433_n;
  wire g1434_p;
  wire g1434_n;
  wire g1435_p;
  wire g1435_n;
  wire g1436_p;
  wire g1436_n;
  wire g1437_p;
  wire g1437_n;
  wire g1438_p;
  wire g1438_n;
  wire g1439_p;
  wire g1439_n;
  wire g1440_p;
  wire g1440_n;
  wire g1441_p;
  wire g1441_n;
  wire g1442_p;
  wire g1442_n;
  wire g1443_p;
  wire g1443_n;
  wire g1444_p;
  wire g1444_n;
  wire g1445_p;
  wire g1445_n;
  wire g1446_p;
  wire g1446_n;
  wire g1447_p;
  wire g1447_n;
  wire g1448_p;
  wire g1448_n;
  wire g1449_p;
  wire g1449_n;
  wire g1450_p;
  wire g1450_n;
  wire g1451_p;
  wire g1451_n;
  wire g1452_p;
  wire g1452_n;
  wire g1453_p;
  wire g1453_n;
  wire g1454_p;
  wire g1454_n;
  wire g1455_p;
  wire g1455_n;
  wire g1456_p;
  wire g1456_n;
  wire g1457_p;
  wire g1457_n;
  wire g1458_p;
  wire g1458_n;
  wire g1459_p;
  wire g1459_n;
  wire g1460_p;
  wire g1460_n;
  wire g1461_p;
  wire g1461_n;
  wire g1462_p;
  wire g1462_n;
  wire g1463_p;
  wire g1463_n;
  wire g1464_p;
  wire g1464_n;
  wire g1465_p;
  wire g1465_n;
  wire g1466_p;
  wire g1466_n;
  wire g1467_p;
  wire g1467_n;
  wire g1468_p;
  wire g1468_n;
  wire g1469_p;
  wire g1469_n;
  wire g1470_p;
  wire g1470_n;
  wire g1471_p;
  wire g1471_n;
  wire g1472_p;
  wire g1472_n;
  wire g1473_p;
  wire g1473_n;
  wire g1474_p;
  wire g1474_n;
  wire g1475_p;
  wire g1475_n;
  wire g1476_p;
  wire g1476_n;
  wire g1477_p;
  wire g1477_n;
  wire g1478_p;
  wire g1478_n;
  wire g1479_p;
  wire g1479_n;
  wire g1480_p;
  wire g1480_n;
  wire g1481_p;
  wire g1481_n;
  wire g1482_p;
  wire g1482_n;
  wire g1483_p;
  wire g1483_n;
  wire g1484_p;
  wire g1484_n;
  wire g1485_p;
  wire g1485_n;
  wire g1486_p;
  wire g1486_n;
  wire g1487_p;
  wire g1487_n;
  wire g1488_p;
  wire g1488_n;
  wire g1489_p;
  wire g1489_n;
  wire g1490_p;
  wire g1490_n;
  wire g1491_p;
  wire g1491_n;
  wire g1492_p;
  wire g1492_n;
  wire g1493_p;
  wire g1493_n;
  wire g1494_p;
  wire g1494_n;
  wire g1495_p;
  wire g1495_n;
  wire g1496_p;
  wire g1496_n;
  wire g1497_p;
  wire g1497_n;
  wire g1498_p;
  wire g1498_n;
  wire g1499_p;
  wire g1499_n;
  wire g1500_p;
  wire g1500_n;
  wire g1501_p;
  wire g1501_n;
  wire g1502_p;
  wire g1502_n;
  wire g1503_p;
  wire g1503_n;
  wire g1504_p;
  wire g1504_n;
  wire g1505_p;
  wire g1505_n;
  wire g1506_p;
  wire g1506_n;
  wire g1507_p;
  wire g1507_n;
  wire g1508_p;
  wire g1508_n;
  wire g1509_p;
  wire g1509_n;
  wire g1510_p;
  wire g1510_n;
  wire g1511_p;
  wire g1511_n;
  wire g1512_p;
  wire g1512_n;
  wire g1513_p;
  wire g1513_n;
  wire g1514_p;
  wire g1514_n;
  wire g1515_p;
  wire g1515_n;
  wire g1516_p;
  wire g1516_n;
  wire g1517_p;
  wire g1517_n;
  wire g1518_p;
  wire g1518_n;
  wire g1519_p;
  wire g1519_n;
  wire g1520_p;
  wire g1520_n;
  wire g1521_p;
  wire g1521_n;
  wire g1522_p;
  wire g1522_n;
  wire g1523_p;
  wire g1523_n;
  wire g1524_p;
  wire g1524_n;
  wire g1525_p;
  wire g1525_n;
  wire g1526_p;
  wire g1526_n;
  wire g1527_p;
  wire g1527_n;
  wire g1528_p;
  wire g1528_n;
  wire g1529_p;
  wire g1529_n;
  wire g1530_p;
  wire g1530_n;
  wire g1531_p;
  wire g1531_n;
  wire g1532_p;
  wire g1532_n;
  wire g1533_p;
  wire g1533_n;
  wire g1534_p;
  wire g1534_n;
  wire g1535_p;
  wire g1535_n;
  wire g1536_p;
  wire g1536_n;
  wire g1537_p;
  wire g1537_n;
  wire g1538_p;
  wire g1538_n;
  wire g1539_p;
  wire g1539_n;
  wire g1540_p;
  wire g1540_n;
  wire g1541_p;
  wire g1541_n;
  wire g1542_p;
  wire g1542_n;
  wire g1543_p;
  wire g1543_n;
  wire g1544_p;
  wire g1544_n;
  wire g1545_p;
  wire g1545_n;
  wire g1546_p;
  wire g1546_n;
  wire g1547_p;
  wire g1547_n;
  wire g1548_p;
  wire g1548_n;
  wire g1549_p;
  wire g1549_n;
  wire g1550_p;
  wire g1550_n;
  wire g1551_p;
  wire g1551_n;
  wire g1552_p;
  wire g1552_n;
  wire g1553_p;
  wire g1553_n;
  wire g1554_p;
  wire g1554_n;
  wire g1555_p;
  wire g1555_n;
  wire g1556_p;
  wire g1556_n;
  wire g1557_p;
  wire g1557_n;
  wire g1558_p;
  wire g1558_n;
  wire g1559_p;
  wire g1559_n;
  wire g1560_p;
  wire g1560_n;
  wire g1561_p;
  wire g1561_n;
  wire g1562_p;
  wire g1562_n;
  wire g1563_p;
  wire g1563_n;
  wire g1564_p;
  wire g1564_n;
  wire g1565_p;
  wire g1565_n;
  wire g1566_p;
  wire g1566_n;
  wire g1567_p;
  wire g1567_n;
  wire g1568_p;
  wire g1568_n;
  wire g1569_p;
  wire g1569_n;
  wire g1570_p;
  wire g1570_n;
  wire g1571_p;
  wire g1571_n;
  wire g1572_p;
  wire g1572_n;
  wire g1573_p;
  wire g1573_n;
  wire g1574_p;
  wire g1574_n;
  wire g1575_p;
  wire g1575_n;
  wire g1576_p;
  wire g1576_n;
  wire g1577_p;
  wire g1577_n;
  wire g1578_p;
  wire g1578_n;
  wire g1579_p;
  wire g1579_n;
  wire g1580_p;
  wire g1580_n;
  wire g1581_p;
  wire g1581_n;
  wire g1582_p;
  wire g1582_n;
  wire g1583_p;
  wire g1583_n;
  wire g1584_p;
  wire g1584_n;
  wire g1585_p;
  wire g1585_n;
  wire g1586_p;
  wire g1586_n;
  wire g1587_p;
  wire g1587_n;
  wire g1588_p;
  wire g1588_n;
  wire g1589_p;
  wire g1589_n;
  wire g1590_p;
  wire g1590_n;
  wire g1591_p;
  wire g1591_n;
  wire g1592_p;
  wire g1592_n;
  wire g1593_p;
  wire g1593_n;
  wire g1594_p;
  wire g1594_n;
  wire g1595_p;
  wire g1595_n;
  wire g1596_p;
  wire g1596_n;
  wire g1597_p;
  wire g1597_n;
  wire g1598_p;
  wire g1598_n;
  wire g1599_p;
  wire g1599_n;
  wire g1600_p;
  wire g1600_n;
  wire g1601_p;
  wire g1601_n;
  wire g1602_p;
  wire g1602_n;
  wire g1603_p;
  wire g1603_n;
  wire g1604_p;
  wire g1604_n;
  wire g1605_p;
  wire g1605_n;
  wire g1606_p;
  wire g1606_n;
  wire g1607_p;
  wire g1607_n;
  wire g1608_p;
  wire g1608_n;
  wire g1609_p;
  wire g1609_n;
  wire g1610_p;
  wire g1610_n;
  wire g1611_p;
  wire g1611_n;
  wire g1612_p;
  wire g1612_n;
  wire g1613_p;
  wire g1613_n;
  wire g1614_p;
  wire g1614_n;
  wire g1615_p;
  wire g1615_n;
  wire g1616_p;
  wire g1616_n;
  wire g1617_p;
  wire g1617_n;
  wire g1618_p;
  wire g1618_n;
  wire g1619_p;
  wire g1619_n;
  wire g1620_p;
  wire g1620_n;
  wire g1621_p;
  wire g1621_n;
  wire g1622_p;
  wire g1622_n;
  wire g1623_p;
  wire g1623_n;
  wire g1624_p;
  wire g1624_n;
  wire g1625_p;
  wire g1625_n;
  wire g1626_p;
  wire g1626_n;
  wire g1627_p;
  wire g1627_n;
  wire g1628_p;
  wire g1628_n;
  wire g1629_p;
  wire g1629_n;
  wire g1630_p;
  wire g1630_n;
  wire g1631_p;
  wire g1631_n;
  wire g1632_p;
  wire g1632_n;
  wire g1633_p;
  wire g1633_n;
  wire g1634_p;
  wire g1634_n;
  wire g1635_p;
  wire g1635_n;
  wire g1636_p;
  wire g1636_n;
  wire g1637_p;
  wire g1637_n;
  wire g1638_p;
  wire g1638_n;
  wire g1639_p;
  wire g1639_n;
  wire g1640_p;
  wire g1640_n;
  wire g1641_p;
  wire g1641_n;
  wire g1642_p;
  wire g1642_n;
  wire g1643_p;
  wire g1643_n;
  wire g1644_p;
  wire g1644_n;
  wire g1645_p;
  wire g1645_n;
  wire g1646_p;
  wire g1646_n;
  wire g1647_p;
  wire g1647_n;
  wire g1648_p;
  wire g1648_n;
  wire g1649_p;
  wire g1649_n;
  wire g1650_p;
  wire g1650_n;
  wire g1651_p;
  wire g1651_n;
  wire g1652_p;
  wire g1652_n;
  wire g1653_p;
  wire g1653_n;
  wire g1654_p;
  wire g1654_n;
  wire g1655_p;
  wire g1655_n;
  wire g1656_p;
  wire g1656_n;
  wire g1657_p;
  wire g1657_n;
  wire g1658_p;
  wire g1658_n;
  wire g1659_p;
  wire g1659_n;
  wire g1660_p;
  wire g1660_n;
  wire g1661_p;
  wire g1661_n;
  wire g1662_p;
  wire g1662_n;
  wire g1663_p;
  wire g1663_n;
  wire g1664_p;
  wire g1664_n;
  wire g1665_p;
  wire g1665_n;
  wire g1666_p;
  wire g1666_n;
  wire g1667_p;
  wire g1667_n;
  wire g1668_p;
  wire g1668_n;
  wire g1669_p;
  wire g1669_n;
  wire g1670_p;
  wire g1670_n;
  wire g1671_p;
  wire g1671_n;
  wire g1672_p;
  wire g1672_n;
  wire g1673_p;
  wire g1673_n;
  wire g1674_p;
  wire g1674_n;
  wire g1675_p;
  wire g1675_n;
  wire g1676_p;
  wire g1676_n;
  wire g1677_p;
  wire g1677_n;
  wire g1678_p;
  wire g1678_n;
  wire g1679_p;
  wire g1679_n;
  wire g1680_p;
  wire g1680_n;
  wire g1681_p;
  wire g1681_n;
  wire g1682_p;
  wire g1682_n;
  wire g1683_p;
  wire g1683_n;
  wire g1684_p;
  wire g1684_n;
  wire g1685_p;
  wire g1685_n;
  wire g1686_p;
  wire g1686_n;
  wire g1687_p;
  wire g1687_n;
  wire g1688_p;
  wire g1688_n;
  wire g1689_p;
  wire g1689_n;
  wire g1690_p;
  wire g1690_n;
  wire g1691_p;
  wire g1691_n;
  wire g1692_p;
  wire g1692_n;
  wire g1693_p;
  wire g1693_n;
  wire g1694_p;
  wire g1694_n;
  wire g1695_p;
  wire g1695_n;
  wire g1696_p;
  wire g1696_n;
  wire g1697_p;
  wire g1697_n;
  wire g1698_p;
  wire g1698_n;
  wire g1699_p;
  wire g1699_n;
  wire g1700_p;
  wire g1700_n;
  wire g1701_p;
  wire g1701_n;
  wire g1702_p;
  wire g1702_n;
  wire g1703_p;
  wire g1703_n;
  wire g1704_p;
  wire g1704_n;
  wire g1705_p;
  wire g1705_n;
  wire g1706_p;
  wire g1706_n;
  wire g1707_p;
  wire g1707_n;
  wire g1708_p;
  wire g1708_n;
  wire g1709_p;
  wire g1709_n;
  wire g1710_p;
  wire g1710_n;
  wire g1711_p;
  wire g1711_n;
  wire g1712_p;
  wire g1712_n;
  wire g1713_p;
  wire g1713_n;
  wire g1714_p;
  wire g1714_n;
  wire g1715_p;
  wire g1715_n;
  wire g1716_p;
  wire g1716_n;
  wire g1717_p;
  wire g1717_n;
  wire g1718_p;
  wire g1718_n;
  wire g1719_p;
  wire g1719_n;
  wire g1720_p;
  wire g1720_n;
  wire g1721_p;
  wire g1721_n;
  wire g1722_p;
  wire g1722_n;
  wire g1723_p;
  wire g1723_n;
  wire g1724_p;
  wire g1724_n;
  wire g1725_p;
  wire g1725_n;
  wire g1726_p;
  wire g1726_n;
  wire g1727_p;
  wire g1727_n;
  wire g1728_p;
  wire g1728_n;
  wire g1729_p;
  wire g1729_n;
  wire g1730_p;
  wire g1730_n;
  wire g1731_p;
  wire g1731_n;
  wire g1732_p;
  wire g1732_n;
  wire g1733_p;
  wire g1733_n;
  wire g1734_p;
  wire g1734_n;
  wire g1735_p;
  wire g1735_n;
  wire g1736_p;
  wire g1736_n;
  wire g1737_p;
  wire g1737_n;
  wire g1738_p;
  wire g1738_n;
  wire g1739_p;
  wire g1739_n;
  wire g1740_p;
  wire g1740_n;
  wire g1741_p;
  wire g1741_n;
  wire g1742_p;
  wire g1742_n;
  wire g1743_p;
  wire g1743_n;
  wire g1744_p;
  wire g1744_n;
  wire g1745_p;
  wire g1745_n;
  wire g1746_p;
  wire g1746_n;
  wire g1747_p;
  wire g1747_n;
  wire g1748_p;
  wire g1748_n;
  wire g1749_p;
  wire g1749_n;
  wire g1750_p;
  wire g1750_n;
  wire g1751_p;
  wire g1751_n;
  wire g1752_p;
  wire g1752_n;
  wire g1753_p;
  wire g1753_n;
  wire g1754_p;
  wire g1754_n;
  wire g1755_p;
  wire g1755_n;
  wire g1756_p;
  wire g1756_n;
  wire g1757_p;
  wire g1757_n;
  wire g1758_p;
  wire g1758_n;
  wire g1759_p;
  wire g1759_n;
  wire g1760_p;
  wire g1760_n;
  wire g1761_p;
  wire g1761_n;
  wire g1762_p;
  wire g1762_n;
  wire g1763_p;
  wire g1763_n;
  wire g1764_p;
  wire g1764_n;
  wire g1765_p;
  wire g1765_n;
  wire g1766_p;
  wire g1766_n;
  wire g1767_p;
  wire g1767_n;
  wire g1768_p;
  wire g1768_n;
  wire g1769_p;
  wire g1769_n;
  wire g1770_p;
  wire g1770_n;
  wire g1771_p;
  wire g1771_n;
  wire g1772_p;
  wire g1772_n;
  wire g1773_p;
  wire g1773_n;
  wire g1774_p;
  wire g1774_n;
  wire g1775_p;
  wire g1775_n;
  wire g1776_p;
  wire g1776_n;
  wire g1777_p;
  wire g1777_n;
  wire g1778_p;
  wire g1778_n;
  wire g1779_p;
  wire g1779_n;
  wire g1780_p;
  wire g1780_n;
  wire g1781_p;
  wire g1781_n;
  wire g1782_p;
  wire g1782_n;
  wire g1783_p;
  wire g1783_n;
  wire g1784_p;
  wire g1784_n;
  wire g1785_p;
  wire g1785_n;
  wire g1786_p;
  wire g1786_n;
  wire g1787_p;
  wire g1787_n;
  wire g1788_p;
  wire g1788_n;
  wire g1789_p;
  wire g1789_n;
  wire g1790_p;
  wire g1790_n;
  wire g1791_p;
  wire g1791_n;
  wire g1792_p;
  wire g1792_n;
  wire g1793_p;
  wire g1793_n;
  wire g1794_p;
  wire g1794_n;
  wire g1795_p;
  wire g1795_n;
  wire g1796_p;
  wire g1796_n;
  wire g1797_p;
  wire g1797_n;
  wire g1798_p;
  wire g1798_n;
  wire g1799_p;
  wire g1799_n;
  wire g1800_p;
  wire g1800_n;
  wire g1801_p;
  wire g1801_n;
  wire g1802_p;
  wire g1802_n;
  wire g1803_p;
  wire g1803_n;
  wire g1804_p;
  wire g1804_n;
  wire g1805_p;
  wire g1805_n;
  wire g1806_p;
  wire g1806_n;
  wire g1807_p;
  wire g1807_n;
  wire g1808_p;
  wire g1808_n;
  wire g1809_p;
  wire g1809_n;
  wire g1810_p;
  wire g1810_n;
  wire g1811_p;
  wire g1811_n;
  wire g1812_p;
  wire g1812_n;
  wire g1813_p;
  wire g1813_n;
  wire g1814_p;
  wire g1814_n;
  wire g1815_p;
  wire g1815_n;
  wire g1816_p;
  wire g1816_n;
  wire g1817_p;
  wire g1817_n;
  wire g1818_p;
  wire g1818_n;
  wire g1819_p;
  wire g1819_n;
  wire g1820_p;
  wire g1820_n;
  wire g1821_p;
  wire g1821_n;
  wire g1822_p;
  wire g1822_n;
  wire g1823_p;
  wire g1823_n;
  wire g1824_p;
  wire g1824_n;
  wire g1825_p;
  wire g1825_n;
  wire g1826_p;
  wire g1826_n;
  wire g1827_p;
  wire g1827_n;
  wire g1828_p;
  wire g1828_n;
  wire g1829_p;
  wire g1829_n;
  wire g1830_p;
  wire g1830_n;
  wire g1831_p;
  wire g1831_n;
  wire g1832_p;
  wire g1832_n;
  wire g1833_p;
  wire g1833_n;
  wire g1834_p;
  wire g1834_n;
  wire g1835_p;
  wire g1835_n;
  wire g1836_p;
  wire g1836_n;
  wire g1837_p;
  wire g1837_n;
  wire g1838_p;
  wire g1838_n;
  wire g1839_p;
  wire g1839_n;
  wire g1840_p;
  wire g1840_n;
  wire g1841_p;
  wire g1841_n;
  wire g1842_p;
  wire g1842_n;
  wire g1843_p;
  wire g1843_n;
  wire g1844_p;
  wire g1844_n;
  wire g1845_p;
  wire g1845_n;
  wire g1846_p;
  wire g1846_n;
  wire g1847_p;
  wire g1847_n;
  wire g1848_p;
  wire g1848_n;
  wire g1849_p;
  wire g1849_n;
  wire g1850_p;
  wire g1850_n;
  wire g1851_p;
  wire g1851_n;
  wire g1852_p;
  wire g1852_n;
  wire g1853_p;
  wire g1853_n;
  wire g1854_p;
  wire g1854_n;
  wire g1855_p;
  wire g1855_n;
  wire g1856_p;
  wire g1856_n;
  wire g1857_p;
  wire g1857_n;
  wire g1858_p;
  wire g1858_n;
  wire g1859_p;
  wire g1859_n;
  wire g1860_p;
  wire g1860_n;
  wire g1861_p;
  wire g1861_n;
  wire g1862_p;
  wire g1862_n;
  wire g1863_p;
  wire g1863_n;
  wire g1864_p;
  wire g1864_n;
  wire g1865_p;
  wire g1865_n;
  wire g1866_p;
  wire g1866_n;
  wire g1867_p;
  wire g1867_n;
  wire g1868_p;
  wire g1868_n;
  wire g1869_p;
  wire g1869_n;
  wire g1870_p;
  wire g1870_n;
  wire g1871_p;
  wire g1871_n;
  wire g1872_p;
  wire g1872_n;
  wire g1873_p;
  wire g1873_n;
  wire g1874_p;
  wire g1874_n;
  wire g1875_p;
  wire g1875_n;
  wire g1876_p;
  wire g1876_n;
  wire g1877_p;
  wire g1877_n;
  wire g1878_p;
  wire g1878_n;
  wire g1879_p;
  wire g1879_n;
  wire g1880_p;
  wire g1880_n;
  wire g1881_p;
  wire g1881_n;
  wire g1882_p;
  wire g1882_n;
  wire g1883_p;
  wire g1883_n;
  wire g1884_p;
  wire g1884_n;
  wire g1885_p;
  wire g1885_n;
  wire g1886_p;
  wire g1886_n;
  wire g1887_p;
  wire g1887_n;
  wire g1888_p;
  wire g1888_n;
  wire g1889_p;
  wire g1889_n;
  wire g1890_p;
  wire g1890_n;
  wire g1891_p;
  wire g1891_n;
  wire g1892_p;
  wire g1892_n;
  wire g1893_p;
  wire g1893_n;
  wire g1894_p;
  wire g1894_n;
  wire g1895_p;
  wire g1895_n;
  wire g1896_p;
  wire g1896_n;
  wire g1897_p;
  wire g1897_n;
  wire g1898_p;
  wire g1898_n;
  wire g1899_p;
  wire g1899_n;
  wire g1900_p;
  wire g1900_n;
  wire g1901_p;
  wire g1901_n;
  wire g1902_p;
  wire g1902_n;
  wire g1903_p;
  wire g1903_n;
  wire g1904_p;
  wire g1904_n;
  wire g1905_p;
  wire g1905_n;
  wire g1906_p;
  wire g1906_n;
  wire g1907_p;
  wire g1907_n;
  wire g1908_p;
  wire g1908_n;
  wire g1909_p;
  wire g1909_n;
  wire g1910_p;
  wire g1910_n;
  wire g1911_p;
  wire g1911_n;
  wire g1912_p;
  wire g1912_n;
  wire g1913_p;
  wire g1913_n;
  wire g1914_p;
  wire g1914_n;
  wire g1915_p;
  wire g1915_n;
  wire g1916_p;
  wire g1916_n;
  wire g1917_p;
  wire g1917_n;
  wire g1918_p;
  wire g1918_n;
  wire g1919_p;
  wire g1919_n;
  wire g1920_p;
  wire g1920_n;
  wire g1921_p;
  wire g1921_n;
  wire g1922_p;
  wire g1922_n;
  wire g1923_p;
  wire g1923_n;
  wire g1924_p;
  wire g1924_n;
  wire g1925_p;
  wire g1925_n;
  wire g1926_p;
  wire g1926_n;
  wire g1927_p;
  wire g1927_n;
  wire g1928_p;
  wire g1928_n;
  wire g1929_p;
  wire g1929_n;
  wire g1930_p;
  wire g1930_n;
  wire g1931_p;
  wire g1931_n;
  wire g1932_p;
  wire g1932_n;
  wire g1933_p;
  wire g1933_n;
  wire g1934_p;
  wire g1934_n;
  wire g1935_p;
  wire g1935_n;
  wire g1936_p;
  wire g1936_n;
  wire g1937_p;
  wire g1937_n;
  wire g1938_p;
  wire g1938_n;
  wire g1939_p;
  wire g1939_n;
  wire g1940_p;
  wire g1940_n;
  wire g1941_p;
  wire g1941_n;
  wire g1942_p;
  wire g1942_n;
  wire g1943_p;
  wire g1943_n;
  wire g1944_p;
  wire g1944_n;
  wire g1945_p;
  wire g1945_n;
  wire g1946_p;
  wire g1946_n;
  wire g1947_p;
  wire g1947_n;
  wire g1948_p;
  wire g1948_n;
  wire g1949_p;
  wire g1949_n;
  wire g1950_p;
  wire g1950_n;
  wire g1951_p;
  wire g1951_n;
  wire g1952_p;
  wire g1952_n;
  wire g1953_p;
  wire g1953_n;
  wire g1954_p;
  wire g1954_n;
  wire g1955_p;
  wire g1955_n;
  wire g1956_p;
  wire g1956_n;
  wire g1957_p;
  wire g1957_n;
  wire g1958_p;
  wire g1958_n;
  wire g1959_p;
  wire g1959_n;
  wire g1960_p;
  wire g1960_n;
  wire g1961_p;
  wire g1961_n;
  wire g1962_p;
  wire g1962_n;
  wire g1963_p;
  wire g1963_n;
  wire g1964_p;
  wire g1964_n;
  wire g1965_p;
  wire g1965_n;
  wire g1966_p;
  wire g1966_n;
  wire g1967_p;
  wire g1967_n;
  wire g1968_p;
  wire g1968_n;
  wire g1969_p;
  wire g1969_n;
  wire g1970_p;
  wire g1970_n;
  wire g1971_p;
  wire g1971_n;
  wire g1972_p;
  wire g1972_n;
  wire g1973_p;
  wire g1973_n;
  wire g1974_p;
  wire g1974_n;
  wire g1975_p;
  wire g1975_n;
  wire g1976_p;
  wire g1976_n;
  wire g1977_p;
  wire g1977_n;
  wire g1978_p;
  wire g1978_n;
  wire g1979_p;
  wire g1979_n;
  wire g1980_p;
  wire g1980_n;
  wire g1981_p;
  wire g1981_n;
  wire g1982_p;
  wire g1982_n;
  wire g1983_p;
  wire g1983_n;
  wire g1984_p;
  wire g1984_n;
  wire g1985_p;
  wire g1985_n;
  wire g1986_p;
  wire g1986_n;
  wire g1987_p;
  wire g1987_n;
  wire g1988_p;
  wire g1988_n;
  wire g1989_p;
  wire g1989_n;
  wire g1990_p;
  wire g1990_n;
  wire g1991_p;
  wire g1991_n;
  wire g1992_p;
  wire g1992_n;
  wire g1993_p;
  wire g1993_n;
  wire g1994_p;
  wire g1994_n;
  wire g1995_p;
  wire g1995_n;
  wire g1996_p;
  wire g1996_n;
  wire g1997_p;
  wire g1997_n;
  wire g1998_p;
  wire g1998_n;
  wire g1999_p;
  wire g1999_n;
  wire g2000_p;
  wire g2000_n;
  wire g2001_p;
  wire g2001_n;
  wire g2002_p;
  wire g2002_n;
  wire g2003_p;
  wire g2003_n;
  wire g2004_p;
  wire g2004_n;
  wire g2005_p;
  wire g2005_n;
  wire g2006_p;
  wire g2006_n;
  wire g2007_p;
  wire g2007_n;
  wire g2008_p;
  wire g2008_n;
  wire g2009_p;
  wire g2009_n;
  wire g2010_p;
  wire g2010_n;
  wire g2011_p;
  wire g2011_n;
  wire g2012_p;
  wire g2012_n;
  wire g2013_p;
  wire g2013_n;
  wire g2014_p;
  wire g2014_n;
  wire g2015_p;
  wire g2015_n;
  wire g2016_p;
  wire g2016_n;
  wire g2017_p;
  wire g2017_n;
  wire g2018_p;
  wire g2018_n;
  wire g2019_p;
  wire g2019_n;
  wire g2020_p;
  wire g2020_n;
  wire g2021_p;
  wire g2021_n;
  wire g2022_p;
  wire g2022_n;
  wire g2023_p;
  wire g2023_n;
  wire g2024_p;
  wire g2024_n;
  wire g2025_p;
  wire g2025_n;
  wire g2026_p;
  wire g2026_n;
  wire g2027_p;
  wire g2027_n;
  wire g2028_p;
  wire g2028_n;
  wire g2029_p;
  wire g2029_n;
  wire g2030_p;
  wire g2030_n;
  wire g2031_p;
  wire g2031_n;
  wire g2032_p;
  wire g2032_n;
  wire g2033_p;
  wire g2033_n;
  wire g2034_p;
  wire g2034_n;
  wire g2035_p;
  wire g2035_n;
  wire g2036_p;
  wire g2036_n;
  wire g2037_p;
  wire g2037_n;
  wire g2038_p;
  wire g2038_n;
  wire g2039_p;
  wire g2039_n;
  wire g2040_p;
  wire g2040_n;
  wire g2041_p;
  wire g2041_n;
  wire g2042_p;
  wire g2042_n;
  wire g2043_p;
  wire g2043_n;
  wire g2044_p;
  wire g2044_n;
  wire g2045_p;
  wire g2045_n;
  wire g2046_p;
  wire g2046_n;
  wire g2047_p;
  wire g2047_n;
  wire g2048_p;
  wire g2048_n;
  wire g2049_p;
  wire g2049_n;
  wire g2050_p;
  wire g2050_n;
  wire g2051_p;
  wire g2051_n;
  wire g2052_p;
  wire g2052_n;
  wire g2053_p;
  wire g2053_n;
  wire g2054_p;
  wire g2054_n;
  wire g2055_p;
  wire g2055_n;
  wire g2056_p;
  wire g2056_n;
  wire g2057_p;
  wire g2057_n;
  wire g2058_p;
  wire g2058_n;
  wire g2059_p;
  wire g2059_n;
  wire g2060_p;
  wire g2060_n;
  wire g2061_p;
  wire g2061_n;
  wire g2062_p;
  wire g2062_n;
  wire g2063_p;
  wire g2063_n;
  wire g2064_p;
  wire g2064_n;
  wire g2065_p;
  wire g2065_n;
  wire g2066_p;
  wire g2066_n;
  wire g2067_p;
  wire g2067_n;
  wire g2068_p;
  wire g2068_n;
  wire g2069_p;
  wire g2069_n;
  wire g2070_p;
  wire g2070_n;
  wire g2071_p;
  wire g2071_n;
  wire g2072_p;
  wire g2072_n;
  wire g2073_p;
  wire g2073_n;
  wire g2074_p;
  wire g2074_n;
  wire g2075_p;
  wire g2075_n;
  wire g2076_p;
  wire g2076_n;
  wire g2077_p;
  wire g2077_n;
  wire g2078_p;
  wire g2078_n;
  wire g2079_p;
  wire g2079_n;
  wire g2080_p;
  wire g2080_n;
  wire g2081_p;
  wire g2081_n;
  wire g2082_p;
  wire g2082_n;
  wire g2083_p;
  wire g2083_n;
  wire g2084_p;
  wire g2084_n;
  wire g2085_p;
  wire g2085_n;
  wire g2086_p;
  wire g2086_n;
  wire g2087_p;
  wire g2087_n;
  wire g2088_p;
  wire g2088_n;
  wire g2089_p;
  wire g2089_n;
  wire g2090_p;
  wire g2090_n;
  wire g2091_p;
  wire g2091_n;
  wire g2092_p;
  wire g2092_n;
  wire g2093_p;
  wire g2093_n;
  wire g2094_p;
  wire g2094_n;
  wire g2095_p;
  wire g2095_n;
  wire g2096_p;
  wire g2096_n;
  wire g2097_p;
  wire g2097_n;
  wire g2098_p;
  wire g2098_n;
  wire g2099_p;
  wire g2099_n;
  wire g2100_p;
  wire g2100_n;
  wire g2101_p;
  wire g2101_n;
  wire g2102_p;
  wire g2102_n;
  wire g2103_p;
  wire g2103_n;
  wire g2104_p;
  wire g2104_n;
  wire g2105_p;
  wire g2105_n;
  wire g2106_p;
  wire g2106_n;
  wire g2107_p;
  wire g2107_n;
  wire g2108_p;
  wire g2108_n;
  wire g2109_p;
  wire g2109_n;
  wire g2110_p;
  wire g2110_n;
  wire g2111_p;
  wire g2111_n;
  wire g2112_p;
  wire g2112_n;
  wire g2113_p;
  wire g2113_n;
  wire g2114_p;
  wire g2114_n;
  wire g2115_p;
  wire g2115_n;
  wire g2116_p;
  wire g2116_n;
  wire g2117_p;
  wire g2117_n;
  wire g2118_p;
  wire g2118_n;
  wire g2119_p;
  wire g2119_n;
  wire g2120_p;
  wire g2120_n;
  wire g2121_p;
  wire g2121_n;
  wire g2122_p;
  wire g2122_n;
  wire g2123_p;
  wire g2123_n;
  wire g2124_p;
  wire g2124_n;
  wire g2125_p;
  wire g2125_n;
  wire g2126_p;
  wire g2126_n;
  wire g2127_p;
  wire g2127_n;
  wire g2128_p;
  wire g2128_n;
  wire g2129_p;
  wire g2129_n;
  wire g2130_p;
  wire g2130_n;
  wire g2131_p;
  wire g2131_n;
  wire g2132_p;
  wire g2132_n;
  wire g2133_p;
  wire g2133_n;
  wire g2134_p;
  wire g2134_n;
  wire g2135_p;
  wire g2135_n;
  wire g2136_p;
  wire g2136_n;
  wire g2137_p;
  wire g2137_n;
  wire g2138_p;
  wire g2138_n;
  wire g2139_p;
  wire g2139_n;
  wire g2140_p;
  wire g2140_n;
  wire g2141_p;
  wire g2141_n;
  wire g2142_p;
  wire g2142_n;
  wire g2143_p;
  wire g2143_n;
  wire g2144_p;
  wire g2144_n;
  wire g2145_p;
  wire g2145_n;
  wire g2146_p;
  wire g2146_n;
  wire g2147_p;
  wire g2147_n;
  wire g2148_p;
  wire g2148_n;
  wire g2149_p;
  wire g2149_n;
  wire g2150_p;
  wire g2150_n;
  wire g2151_p;
  wire g2151_n;
  wire g2152_p;
  wire g2152_n;
  wire g2153_p;
  wire g2153_n;
  wire g2154_p;
  wire g2154_n;
  wire g2155_p;
  wire g2155_n;
  wire g2156_p;
  wire g2156_n;
  wire g2157_p;
  wire g2157_n;
  wire g2158_p;
  wire g2158_n;
  wire g2159_p;
  wire g2159_n;
  wire g2160_p;
  wire g2160_n;
  wire g2161_p;
  wire g2161_n;
  wire g2162_p;
  wire g2162_n;
  wire g2163_p;
  wire g2163_n;
  wire g2164_p;
  wire g2164_n;
  wire g2165_p;
  wire g2165_n;
  wire g2166_p;
  wire g2166_n;
  wire g2167_p;
  wire g2167_n;
  wire g2168_p;
  wire g2168_n;
  wire g2169_p;
  wire g2169_n;
  wire g2170_p;
  wire g2170_n;
  wire g2171_p;
  wire g2171_n;
  wire g2172_p;
  wire g2172_n;
  wire g2173_p;
  wire g2173_n;
  wire g2174_p;
  wire g2174_n;
  wire g2175_p;
  wire g2175_n;
  wire g2176_p;
  wire g2176_n;
  wire g2177_p;
  wire g2177_n;
  wire g2178_p;
  wire g2178_n;
  wire g2179_p;
  wire g2179_n;
  wire g2180_p;
  wire g2180_n;
  wire g2181_p;
  wire g2181_n;
  wire g2182_p;
  wire g2182_n;
  wire g2183_p;
  wire g2183_n;
  wire g2184_p;
  wire g2184_n;
  wire g2185_p;
  wire g2185_n;
  wire g2186_p;
  wire g2186_n;
  wire g2187_p;
  wire g2187_n;
  wire g2188_p;
  wire g2188_n;
  wire g2189_p;
  wire g2189_n;
  wire g2190_p;
  wire g2190_n;
  wire g2191_p;
  wire g2191_n;
  wire g2192_p;
  wire g2192_n;
  wire g2193_p;
  wire g2193_n;
  wire g2194_p;
  wire g2194_n;
  wire g2195_p;
  wire g2195_n;
  wire g2196_p;
  wire g2196_n;
  wire g2197_p;
  wire g2197_n;
  wire g2198_p;
  wire g2198_n;
  wire g2199_p;
  wire g2199_n;
  wire g2200_p;
  wire g2200_n;
  wire g2201_p;
  wire g2201_n;
  wire g2202_p;
  wire g2202_n;
  wire g2203_p;
  wire g2203_n;
  wire g2204_p;
  wire g2204_n;
  wire g2205_p;
  wire g2205_n;
  wire g2206_p;
  wire g2206_n;
  wire g2207_p;
  wire g2207_n;
  wire g2208_p;
  wire g2208_n;
  wire g2209_p;
  wire g2209_n;
  wire g2210_p;
  wire g2210_n;
  wire g2211_p;
  wire g2211_n;
  wire g2212_p;
  wire g2212_n;
  wire g2213_p;
  wire g2213_n;
  wire g2214_p;
  wire g2214_n;
  wire g2215_p;
  wire g2215_n;
  wire g2216_p;
  wire g2216_n;
  wire g2217_p;
  wire g2217_n;
  wire g2218_p;
  wire g2218_n;
  wire g2219_p;
  wire g2219_n;
  wire g2220_p;
  wire g2220_n;
  wire g2221_p;
  wire g2221_n;
  wire g2222_p;
  wire g2222_n;
  wire g2223_p;
  wire g2223_n;
  wire g2224_p;
  wire g2224_n;
  wire g2225_p;
  wire g2225_n;
  wire g2226_p;
  wire g2226_n;
  wire g2227_p;
  wire g2227_n;
  wire g2228_p;
  wire g2228_n;
  wire g2229_p;
  wire g2229_n;
  wire g2230_p;
  wire g2230_n;
  wire g2231_p;
  wire g2231_n;
  wire g2232_p;
  wire g2232_n;
  wire g2233_p;
  wire g2233_n;
  wire g2234_p;
  wire g2234_n;
  wire g2235_p;
  wire g2235_n;
  wire g2236_p;
  wire g2236_n;
  wire g2237_p;
  wire g2237_n;
  wire g2238_p;
  wire g2238_n;
  wire g2239_p;
  wire g2239_n;
  wire g2240_p;
  wire g2240_n;
  wire g2241_p;
  wire g2241_n;
  wire g2242_p;
  wire g2242_n;
  wire g2243_p;
  wire g2243_n;
  wire g2244_p;
  wire g2244_n;
  wire g2245_p;
  wire g2245_n;
  wire g2246_p;
  wire g2246_n;
  wire g2247_p;
  wire g2247_n;
  wire g2248_p;
  wire g2248_n;
  wire g2249_p;
  wire g2249_n;
  wire g2250_p;
  wire g2250_n;
  wire g2251_p;
  wire g2251_n;
  wire g2252_p;
  wire g2252_n;
  wire g2253_p;
  wire g2253_n;
  wire g2254_p;
  wire g2254_n;
  wire g2255_p;
  wire g2255_n;
  wire g2256_p;
  wire g2256_n;
  wire g2257_p;
  wire g2257_n;
  wire g2258_p;
  wire g2258_n;
  wire g2259_p;
  wire g2259_n;
  wire g2260_p;
  wire g2260_n;
  wire g2261_p;
  wire g2261_n;
  wire g2262_p;
  wire g2262_n;
  wire g2263_p;
  wire g2263_n;
  wire g2264_p;
  wire g2264_n;
  wire g2265_p;
  wire g2265_n;
  wire g2266_p;
  wire g2266_n;
  wire g2267_p;
  wire g2267_n;
  wire g2268_p;
  wire g2268_n;
  wire g2269_p;
  wire g2269_n;
  wire g2270_p;
  wire g2270_n;
  wire g2271_p;
  wire g2271_n;
  wire g2272_p;
  wire g2272_n;
  wire g2273_p;
  wire g2273_n;
  wire g2274_p;
  wire g2274_n;
  wire g2275_p;
  wire g2275_n;
  wire g2276_p;
  wire g2276_n;
  wire g2277_p;
  wire g2277_n;
  wire g2278_p;
  wire g2278_n;
  wire g2279_p;
  wire g2279_n;
  wire g2280_p;
  wire g2280_n;
  wire g2281_p;
  wire g2281_n;
  wire g2282_p;
  wire g2282_n;
  wire g2283_p;
  wire g2283_n;
  wire g2284_p;
  wire g2284_n;
  wire g2285_p;
  wire g2285_n;
  wire g2286_p;
  wire g2286_n;
  wire g2287_p;
  wire g2287_n;
  wire g2288_p;
  wire g2288_n;
  wire g2289_p;
  wire g2289_n;
  wire g2290_p;
  wire g2290_n;
  wire g2291_p;
  wire g2291_n;
  wire g2292_p;
  wire g2292_n;
  wire g2293_p;
  wire g2293_n;
  wire g2294_p;
  wire g2294_n;
  wire g2295_p;
  wire g2295_n;
  wire g2296_p;
  wire g2296_n;
  wire g2297_p;
  wire g2297_n;
  wire g2298_p;
  wire g2298_n;
  wire g2299_p;
  wire g2299_n;
  wire g2300_p;
  wire g2300_n;
  wire g2301_p;
  wire g2301_n;
  wire g2302_p;
  wire g2302_n;
  wire g2303_p;
  wire g2303_n;
  wire g2304_p;
  wire g2304_n;
  wire g2305_p;
  wire g2305_n;
  wire g2306_p;
  wire g2306_n;
  wire g2307_p;
  wire g2307_n;
  wire g2308_p;
  wire g2308_n;
  wire g2309_p;
  wire g2309_n;
  wire g2310_p;
  wire g2310_n;
  wire g2311_p;
  wire g2311_n;
  wire g2312_p;
  wire g2312_n;
  wire g2313_p;
  wire g2313_n;
  wire g2314_p;
  wire g2314_n;
  wire g2315_p;
  wire g2315_n;
  wire g2316_p;
  wire g2316_n;
  wire g2317_p;
  wire g2317_n;
  wire g2318_p;
  wire g2318_n;
  wire g2319_p;
  wire g2319_n;
  wire g2320_p;
  wire g2320_n;
  wire g2321_p;
  wire g2321_n;
  wire g2322_p;
  wire g2322_n;
  wire g2323_p;
  wire g2323_n;
  wire g2324_p;
  wire g2324_n;
  wire g2325_p;
  wire g2325_n;
  wire g2326_p;
  wire g2326_n;
  wire g2327_p;
  wire g2327_n;
  wire g2328_p;
  wire g2328_n;
  wire g2329_p;
  wire g2329_n;
  wire g2330_p;
  wire g2330_n;
  wire g2331_p;
  wire g2331_n;
  wire g2332_p;
  wire g2332_n;
  wire g2333_p;
  wire g2333_n;
  wire g2334_p;
  wire g2334_n;
  wire g2335_p;
  wire g2335_n;
  wire g2336_p;
  wire g2336_n;
  wire g2337_p;
  wire g2337_n;
  wire g2338_p;
  wire g2338_n;
  wire g2339_p;
  wire g2339_n;
  wire g2340_p;
  wire g2340_n;
  wire g2341_p;
  wire g2341_n;
  wire g2342_p;
  wire g2342_n;
  wire g2343_p;
  wire g2343_n;
  wire g2344_p;
  wire g2344_n;
  wire g2345_p;
  wire g2345_n;
  wire g2346_p;
  wire g2346_n;
  wire g2347_p;
  wire g2347_n;
  wire g2348_p;
  wire g2348_n;
  wire g2349_p;
  wire g2349_n;
  wire g2350_p;
  wire g2350_n;
  wire g2351_p;
  wire g2351_n;
  wire g2352_p;
  wire g2352_n;
  wire g2353_p;
  wire g2353_n;
  wire g2354_p;
  wire g2354_n;
  wire g2355_p;
  wire g2355_n;
  wire g2356_p;
  wire g2356_n;
  wire g2357_p;
  wire g2357_n;
  wire g2358_p;
  wire g2358_n;
  wire g2359_p;
  wire g2359_n;
  wire g2360_p;
  wire g2360_n;
  wire g2361_p;
  wire g2361_n;
  wire g2362_p;
  wire g2362_n;
  wire g2363_p;
  wire g2363_n;
  wire g2364_p;
  wire g2364_n;
  wire g2365_p;
  wire g2365_n;
  wire g2366_p;
  wire g2366_n;
  wire g2367_p;
  wire g2367_n;
  wire g2368_p;
  wire g2368_n;
  wire g2369_p;
  wire g2369_n;
  wire g2370_p;
  wire g2370_n;
  wire g2371_p;
  wire g2371_n;
  wire g2372_p;
  wire g2372_n;
  wire g2373_p;
  wire g2373_n;
  wire g2374_p;
  wire g2374_n;
  wire g2375_p;
  wire g2375_n;
  wire g2376_p;
  wire g2376_n;
  wire g2377_p;
  wire g2377_n;
  wire g2378_p;
  wire g2378_n;
  wire g2379_p;
  wire g2379_n;
  wire g2380_p;
  wire g2380_n;
  wire g2381_p;
  wire g2381_n;
  wire g2382_p;
  wire g2382_n;
  wire g2383_p;
  wire g2383_n;
  wire g2384_p;
  wire g2384_n;
  wire g2385_p;
  wire g2385_n;
  wire g2386_p;
  wire g2386_n;
  wire g2387_p;
  wire g2387_n;
  wire g2388_p;
  wire g2388_n;
  wire g2389_p;
  wire g2389_n;
  wire g2390_p;
  wire g2390_n;
  wire g2391_p;
  wire g2391_n;
  wire g2392_p;
  wire g2392_n;
  wire g2393_p;
  wire g2393_n;
  wire g2394_p;
  wire g2394_n;
  wire g2395_p;
  wire g2395_n;
  wire g2396_p;
  wire g2396_n;
  wire g2397_p;
  wire g2397_n;
  wire g2398_p;
  wire g2398_n;
  wire g2399_p;
  wire g2399_n;
  wire g2400_p;
  wire g2400_n;
  wire g2401_p;
  wire g2401_n;
  wire g2402_p;
  wire g2402_n;
  wire g2403_p;
  wire g2403_n;
  wire g2404_p;
  wire g2404_n;
  wire g2405_p;
  wire g2405_n;
  wire g2406_p;
  wire g2406_n;
  wire g2407_p;
  wire g2407_n;
  wire g2408_p;
  wire g2408_n;
  wire g2409_p;
  wire g2409_n;
  wire g2410_p;
  wire g2410_n;
  wire g2411_p;
  wire g2411_n;
  wire g2412_p;
  wire g2412_n;
  wire g2413_p;
  wire g2413_n;
  wire g2414_p;
  wire g2414_n;
  wire g2415_p;
  wire g2415_n;
  wire g2416_p;
  wire g2416_n;
  wire g2417_p;
  wire g2417_n;
  wire g2418_p;
  wire g2418_n;
  wire g2419_p;
  wire g2419_n;
  wire g2420_p;
  wire g2420_n;
  wire g2421_p;
  wire g2421_n;
  wire g2422_p;
  wire g2422_n;
  wire g2423_p;
  wire g2423_n;
  wire g2424_p;
  wire g2424_n;
  wire g2425_p;
  wire g2425_n;
  wire g2426_p;
  wire g2426_n;
  wire g2427_p;
  wire g2427_n;
  wire g2428_p;
  wire g2428_n;
  wire g2429_p;
  wire g2429_n;
  wire g2430_p;
  wire g2430_n;
  wire g2431_p;
  wire g2431_n;
  wire g2432_p;
  wire g2432_n;
  wire g2433_p;
  wire g2433_n;
  wire g2434_p;
  wire g2434_n;
  wire g2435_p;
  wire g2435_n;
  wire g2436_p;
  wire g2436_n;
  wire g2437_p;
  wire g2437_n;
  wire g2438_p;
  wire g2438_n;
  wire g2439_p;
  wire g2439_n;
  wire g2440_p;
  wire g2440_n;
  wire g2441_p;
  wire g2441_n;
  wire g2442_p;
  wire g2442_n;
  wire g2443_p;
  wire g2443_n;
  wire g2444_p;
  wire g2444_n;
  wire g2445_p;
  wire g2445_n;
  wire g2446_p;
  wire g2446_n;
  wire g2447_p;
  wire g2447_n;
  wire g2448_p;
  wire g2448_n;
  wire g2449_p;
  wire g2449_n;
  wire g2450_p;
  wire g2450_n;
  wire g2451_p;
  wire g2451_n;
  wire g2452_p;
  wire g2452_n;
  wire g2453_p;
  wire g2453_n;
  wire g2454_p;
  wire g2454_n;
  wire g2455_p;
  wire g2455_n;
  wire g2456_p;
  wire g2456_n;
  wire g2457_p;
  wire g2457_n;
  wire g2458_p;
  wire g2458_n;
  wire g2459_p;
  wire g2459_n;
  wire g2460_p;
  wire g2460_n;
  wire g2461_p;
  wire g2461_n;
  wire g2462_p;
  wire g2462_n;
  wire g2463_p;
  wire g2463_n;
  wire g2464_p;
  wire g2464_n;
  wire g2465_p;
  wire g2465_n;
  wire g2466_p;
  wire g2466_n;
  wire g2467_p;
  wire g2467_n;
  wire g2468_p;
  wire g2468_n;
  wire g2469_p;
  wire g2469_n;
  wire g2470_p;
  wire g2470_n;
  wire g2471_p;
  wire g2471_n;
  wire g2472_p;
  wire g2472_n;
  wire g2473_p;
  wire g2473_n;
  wire g2474_p;
  wire g2474_n;
  wire g2475_p;
  wire g2475_n;
  wire g2476_p;
  wire g2476_n;
  wire g2477_p;
  wire g2477_n;
  wire g2478_p;
  wire g2478_n;
  wire g2479_p;
  wire g2479_n;
  wire g2480_p;
  wire g2480_n;
  wire g2481_p;
  wire g2481_n;
  wire g2482_p;
  wire g2482_n;
  wire g2483_p;
  wire g2483_n;
  wire g2484_p;
  wire g2484_n;
  wire g2485_p;
  wire g2485_n;
  wire g2486_p;
  wire g2486_n;
  wire g2487_p;
  wire g2487_n;
  wire g2488_p;
  wire g2488_n;
  wire g2489_p;
  wire g2489_n;
  wire g2490_p;
  wire g2490_n;
  wire g2491_p;
  wire g2491_n;
  wire g2492_p;
  wire g2492_n;
  wire g2493_p;
  wire g2493_n;
  wire g2494_p;
  wire g2494_n;
  wire g2495_p;
  wire g2495_n;
  wire g2496_p;
  wire g2496_n;
  wire g2497_p;
  wire g2497_n;
  wire g2498_p;
  wire g2498_n;
  wire g2499_p;
  wire g2499_n;
  wire g2500_p;
  wire g2500_n;
  wire g2501_p;
  wire g2501_n;
  wire g2502_p;
  wire g2502_n;
  wire g2503_p;
  wire g2503_n;
  wire g2504_p;
  wire g2504_n;
  wire g2505_p;
  wire g2505_n;
  wire g2506_p;
  wire g2506_n;
  wire g2507_p;
  wire g2507_n;
  wire g2508_p;
  wire g2508_n;
  wire g2509_p;
  wire g2509_n;
  wire g2510_p;
  wire g2510_n;
  wire g2511_p;
  wire g2511_n;
  wire g2512_p;
  wire g2512_n;
  wire g2513_p;
  wire g2513_n;
  wire g2514_p;
  wire g2514_n;
  wire g2515_p;
  wire g2515_n;
  wire g2516_p;
  wire g2516_n;
  wire g2517_p;
  wire g2517_n;
  wire g2518_p;
  wire g2518_n;
  wire g2519_p;
  wire g2519_n;
  wire g2520_p;
  wire g2520_n;
  wire g2521_p;
  wire g2521_n;
  wire g2522_p;
  wire g2522_n;
  wire g2523_p;
  wire g2523_n;
  wire g2524_p;
  wire g2524_n;
  wire g2525_p;
  wire g2525_n;
  wire g2526_p;
  wire g2526_n;
  wire g2527_p;
  wire g2527_n;
  wire g2528_p;
  wire g2528_n;
  wire g2529_p;
  wire g2529_n;
  wire g2530_p;
  wire g2530_n;
  wire g2531_p;
  wire g2531_n;
  wire g2532_p;
  wire g2532_n;
  wire g2533_p;
  wire g2533_n;
  wire g2534_p;
  wire g2534_n;
  wire g2535_p;
  wire g2535_n;
  wire g2536_p;
  wire g2536_n;
  wire g2537_p;
  wire g2537_n;
  wire g2538_p;
  wire g2538_n;
  wire g2539_p;
  wire g2539_n;
  wire g2540_p;
  wire g2540_n;
  wire g2541_p;
  wire g2541_n;
  wire g2542_p;
  wire g2542_n;
  wire g2543_p;
  wire g2543_n;
  wire g2544_p;
  wire g2544_n;
  wire g2545_p;
  wire g2545_n;
  wire g2546_p;
  wire g2546_n;
  wire g2547_p;
  wire g2547_n;
  wire g2548_p;
  wire g2548_n;
  wire g2549_p;
  wire g2549_n;
  wire g2550_p;
  wire g2550_n;
  wire g2551_p;
  wire g2551_n;
  wire g2552_p;
  wire g2552_n;
  wire g2553_p;
  wire g2553_n;
  wire g2554_p;
  wire g2554_n;
  wire g2555_p;
  wire g2555_n;
  wire g2556_p;
  wire g2556_n;
  wire g2557_p;
  wire g2557_n;
  wire g2558_p;
  wire g2558_n;
  wire g2559_p;
  wire g2559_n;
  wire g2560_p;
  wire g2560_n;
  wire g2561_p;
  wire g2561_n;
  wire g2562_p;
  wire g2562_n;
  wire g2563_p;
  wire g2563_n;
  wire g2564_p;
  wire g2564_n;
  wire g2565_p;
  wire g2565_n;
  wire g2566_p;
  wire g2566_n;
  wire g2567_p;
  wire g2567_n;
  wire g2568_p;
  wire g2568_n;
  wire g2569_p;
  wire g2569_n;
  wire g2570_p;
  wire g2570_n;
  wire g2571_p;
  wire g2571_n;
  wire g2572_p;
  wire g2572_n;
  wire g2573_p;
  wire g2573_n;
  wire g2574_p;
  wire g2574_n;
  wire g2575_p;
  wire g2575_n;
  wire g2576_p;
  wire g2576_n;
  wire g2577_p;
  wire g2577_n;
  wire g2578_p;
  wire g2578_n;
  wire g2579_p;
  wire g2579_n;
  wire g2580_p;
  wire g2580_n;
  wire g2581_p;
  wire g2581_n;
  wire g2582_p;
  wire g2582_n;
  wire g2583_p;
  wire g2583_n;
  wire g2584_p;
  wire g2584_n;
  wire g2585_p;
  wire g2585_n;
  wire g2586_p;
  wire g2586_n;
  wire g2587_p;
  wire g2587_n;
  wire g2588_p;
  wire g2588_n;
  wire g2589_p;
  wire g2589_n;
  wire g2590_p;
  wire g2590_n;
  wire g2591_p;
  wire g2591_n;
  wire g2592_p;
  wire g2592_n;
  wire g2593_p;
  wire g2593_n;
  wire g2594_p;
  wire g2594_n;
  wire g2595_p;
  wire g2595_n;
  wire g2596_p;
  wire g2596_n;
  wire g2597_p;
  wire g2597_n;
  wire g2598_p;
  wire g2598_n;
  wire g2599_p;
  wire g2599_n;
  wire g2600_p;
  wire g2600_n;
  wire g2601_p;
  wire g2601_n;
  wire g2602_p;
  wire g2602_n;
  wire g2603_p;
  wire g2603_n;
  wire g2604_p;
  wire g2604_n;
  wire g2605_p;
  wire g2605_n;
  wire g2606_p;
  wire g2606_n;
  wire g2607_p;
  wire g2607_n;
  wire g2608_p;
  wire g2608_n;
  wire g2609_p;
  wire g2609_n;
  wire g2610_p;
  wire g2610_n;
  wire g2611_p;
  wire g2611_n;
  wire g2612_p;
  wire g2612_n;
  wire g2613_p;
  wire g2613_n;
  wire g2614_p;
  wire g2614_n;
  wire g2615_p;
  wire g2615_n;
  wire g2616_p;
  wire g2616_n;
  wire g2617_p;
  wire g2617_n;
  wire g2618_p;
  wire g2618_n;
  wire g2619_p;
  wire g2619_n;
  wire g2620_p;
  wire g2620_n;
  wire g2621_p;
  wire g2621_n;
  wire g2622_p;
  wire g2622_n;
  wire g2623_p;
  wire g2623_n;
  wire g2624_p;
  wire g2624_n;
  wire g2625_p;
  wire g2625_n;
  wire g2626_p;
  wire g2626_n;
  wire g2627_p;
  wire g2627_n;
  wire g2628_p;
  wire g2628_n;
  wire g2629_p;
  wire g2629_n;
  wire g2630_p;
  wire g2630_n;
  wire g2631_p;
  wire g2631_n;
  wire g2632_p;
  wire g2632_n;
  wire g2633_p;
  wire g2633_n;
  wire g2634_p;
  wire g2634_n;
  wire g2635_p;
  wire g2635_n;
  wire g2636_p;
  wire g2636_n;
  wire g2637_p;
  wire g2637_n;
  wire g2638_p;
  wire g2638_n;
  wire g2639_p;
  wire g2639_n;
  wire g2640_p;
  wire g2640_n;
  wire g2641_p;
  wire g2641_n;
  wire g2642_p;
  wire g2642_n;
  wire g2643_p;
  wire g2643_n;
  wire g2644_p;
  wire g2644_n;
  wire g2645_p;
  wire g2645_n;
  wire g2646_p;
  wire g2646_n;
  wire g2647_p;
  wire g2647_n;
  wire g2648_p;
  wire g2648_n;
  wire g2649_p;
  wire g2649_n;
  wire g2650_p;
  wire g2650_n;
  wire g2651_p;
  wire g2651_n;
  wire g2652_p;
  wire g2652_n;
  wire g2653_p;
  wire g2653_n;
  wire g2654_p;
  wire g2654_n;
  wire g2655_p;
  wire g2655_n;
  wire g2656_p;
  wire g2656_n;
  wire g2657_p;
  wire g2657_n;
  wire g2658_p;
  wire g2658_n;
  wire g2659_p;
  wire g2659_n;
  wire g2660_p;
  wire g2660_n;
  wire g2661_p;
  wire g2661_n;
  wire g2662_p;
  wire g2662_n;
  wire g2663_p;
  wire g2663_n;
  wire g2664_p;
  wire g2664_n;
  wire g2665_p;
  wire g2665_n;
  wire g2666_p;
  wire g2666_n;
  wire g2667_p;
  wire g2667_n;
  wire g2668_p;
  wire g2668_n;
  wire g2669_p;
  wire g2669_n;
  wire g2670_p;
  wire g2670_n;
  wire g2671_p;
  wire g2671_n;
  wire g2672_p;
  wire g2672_n;
  wire g2673_p;
  wire g2673_n;
  wire g2674_p;
  wire g2674_n;
  wire g2675_p;
  wire g2675_n;
  wire g2676_p;
  wire g2676_n;
  wire g2677_p;
  wire g2677_n;
  wire g2678_p;
  wire g2678_n;
  wire g2679_p;
  wire g2679_n;
  wire g2680_p;
  wire g2680_n;
  wire g2681_p;
  wire g2681_n;
  wire g2682_p;
  wire g2682_n;
  wire g2683_p;
  wire g2683_n;
  wire g2684_p;
  wire g2684_n;
  wire g2685_p;
  wire g2685_n;
  wire g2686_p;
  wire g2686_n;
  wire g2687_p;
  wire g2687_n;
  wire g2688_p;
  wire g2688_n;
  wire g2689_p;
  wire g2689_n;
  wire g2690_p;
  wire g2690_n;
  wire g2691_p;
  wire g2691_n;
  wire g2692_p;
  wire g2692_n;
  wire g2693_p;
  wire g2693_n;
  wire g2694_p;
  wire g2694_n;
  wire g2695_p;
  wire g2695_n;
  wire g2696_p;
  wire g2696_n;
  wire g2697_p;
  wire g2697_n;
  wire g2698_p;
  wire g2698_n;
  wire g2699_p;
  wire g2699_n;
  wire g2700_p;
  wire g2700_n;
  wire g2701_p;
  wire g2701_n;
  wire g2702_p;
  wire g2702_n;
  wire g2703_p;
  wire g2703_n;
  wire g2704_p;
  wire g2704_n;
  wire g2705_p;
  wire g2705_n;
  wire g2706_p;
  wire g2706_n;
  wire g2707_p;
  wire g2707_n;
  wire g2708_p;
  wire g2708_n;
  wire g2709_p;
  wire g2709_n;
  wire g2710_p;
  wire g2710_n;
  wire g2711_p;
  wire g2711_n;
  wire g2712_p;
  wire g2712_n;
  wire g2713_p;
  wire g2713_n;
  wire g2714_p;
  wire g2714_n;
  wire g2715_p;
  wire g2715_n;
  wire g2716_p;
  wire g2716_n;
  wire g2717_p;
  wire g2717_n;
  wire g2718_p;
  wire g2718_n;
  wire g2719_p;
  wire g2719_n;
  wire g2720_p;
  wire g2720_n;
  wire g2721_p;
  wire g2721_n;
  wire g2722_p;
  wire g2722_n;
  wire g2723_p;
  wire g2723_n;
  wire g2724_p;
  wire g2724_n;
  wire g2725_p;
  wire g2725_n;
  wire g2726_p;
  wire g2726_n;
  wire g2727_p;
  wire g2727_n;
  wire g2728_p;
  wire g2728_n;
  wire g2729_p;
  wire g2729_n;
  wire g2730_p;
  wire g2730_n;
  wire g2731_p;
  wire g2731_n;
  wire g2732_p;
  wire g2732_n;
  wire g2733_p;
  wire g2733_n;
  wire g2734_p;
  wire g2734_n;
  wire g2735_p;
  wire g2735_n;
  wire g2736_p;
  wire g2736_n;
  wire g2737_p;
  wire g2737_n;
  wire g2738_p;
  wire g2738_n;
  wire g2739_p;
  wire g2739_n;
  wire g2740_p;
  wire g2740_n;
  wire g2741_p;
  wire g2741_n;
  wire g2742_p;
  wire g2742_n;
  wire g2743_p;
  wire g2743_n;
  wire g2744_p;
  wire g2744_n;
  wire n4938_o2_p_spl_;
  wire n5122_o2_p_spl_;
  wire n5316_o2_p_spl_;
  wire n5494_o2_p_spl_;
  wire n5682_o2_p_spl_;
  wire n5867_o2_p_spl_;
  wire n6153_o2_p_spl_;
  wire n6509_o2_p_spl_;
  wire n6892_o2_p_spl_;
  wire n7263_o2_p_spl_;
  wire n7788_o2_p_spl_;
  wire G5164_o2_p_spl_;
  wire G5527_o2_p_spl_;
  wire G5868_o2_p_spl_;
  wire G6070_o2_p_spl_;
  wire G6125_o2_p_spl_;
  wire G6134_o2_p_spl_;
  wire G6143_o2_p_spl_;
  wire G6143_o2_p_spl_0;
  wire g460_p_spl_;
  wire g459_p_spl_;
  wire g461_p_spl_;
  wire g461_p_spl_0;
  wire G6008_o2_n_spl_;
  wire G6005_o2_n_spl_;
  wire G6008_o2_p_spl_;
  wire G6005_o2_p_spl_;
  wire g465_n_spl_;
  wire g465_n_spl_0;
  wire g465_p_spl_;
  wire g465_p_spl_0;
  wire g469_p_spl_;
  wire g468_p_spl_;
  wire g470_p_spl_;
  wire g470_p_spl_0;
  wire G5893_o2_n_spl_;
  wire G5893_o2_n_spl_0;
  wire G5893_o2_p_spl_;
  wire G5893_o2_p_spl_0;
  wire g477_n_spl_;
  wire g476_n_spl_;
  wire g477_p_spl_;
  wire g476_p_spl_;
  wire g478_n_spl_;
  wire g478_n_spl_0;
  wire g478_p_spl_;
  wire g478_p_spl_0;
  wire g482_p_spl_;
  wire g481_p_spl_;
  wire g483_p_spl_;
  wire g483_p_spl_0;
  wire n2863_lo_p_spl_;
  wire n2863_lo_p_spl_0;
  wire n2863_lo_p_spl_00;
  wire n2863_lo_p_spl_000;
  wire n2863_lo_p_spl_01;
  wire n2863_lo_p_spl_1;
  wire n2863_lo_p_spl_10;
  wire n2863_lo_p_spl_11;
  wire n2863_lo_n_spl_;
  wire n2863_lo_n_spl_0;
  wire n2863_lo_n_spl_00;
  wire n2863_lo_n_spl_000;
  wire n2863_lo_n_spl_01;
  wire n2863_lo_n_spl_1;
  wire n2863_lo_n_spl_10;
  wire n2863_lo_n_spl_11;
  wire g488_n_spl_;
  wire g487_n_spl_;
  wire g488_p_spl_;
  wire g487_p_spl_;
  wire g489_n_spl_;
  wire g489_n_spl_0;
  wire g489_p_spl_;
  wire g489_p_spl_0;
  wire g493_n_spl_;
  wire g492_n_spl_;
  wire g493_p_spl_;
  wire g492_p_spl_;
  wire g494_n_spl_;
  wire g494_n_spl_0;
  wire g494_p_spl_;
  wire g494_p_spl_0;
  wire g498_p_spl_;
  wire g497_p_spl_;
  wire g499_p_spl_;
  wire g499_p_spl_0;
  wire G5565_o2_n_spl_;
  wire G5562_o2_n_spl_;
  wire G5565_o2_p_spl_;
  wire G5562_o2_p_spl_;
  wire g503_n_spl_;
  wire g503_n_spl_0;
  wire g503_p_spl_;
  wire g503_p_spl_0;
  wire g507_n_spl_;
  wire g506_n_spl_;
  wire g507_p_spl_;
  wire g506_p_spl_;
  wire g508_n_spl_;
  wire g508_n_spl_0;
  wire g508_p_spl_;
  wire g508_p_spl_0;
  wire g512_n_spl_;
  wire g511_n_spl_;
  wire g512_p_spl_;
  wire g511_p_spl_;
  wire g513_n_spl_;
  wire g513_n_spl_0;
  wire g513_p_spl_;
  wire g513_p_spl_0;
  wire g517_p_spl_;
  wire g516_p_spl_;
  wire g518_p_spl_;
  wire g518_p_spl_0;
  wire G5391_o2_n_spl_;
  wire G5391_o2_n_spl_0;
  wire G5391_o2_p_spl_;
  wire G5391_o2_p_spl_0;
  wire g525_n_spl_;
  wire g524_n_spl_;
  wire g525_p_spl_;
  wire g524_p_spl_;
  wire g526_n_spl_;
  wire g526_n_spl_0;
  wire g526_p_spl_;
  wire g526_p_spl_0;
  wire g530_n_spl_;
  wire g529_n_spl_;
  wire g530_p_spl_;
  wire g529_p_spl_;
  wire g531_n_spl_;
  wire g531_n_spl_0;
  wire g531_p_spl_;
  wire g531_p_spl_0;
  wire g535_n_spl_;
  wire g534_n_spl_;
  wire g535_p_spl_;
  wire g534_p_spl_;
  wire g536_n_spl_;
  wire g536_n_spl_0;
  wire g536_p_spl_;
  wire g536_p_spl_0;
  wire g540_p_spl_;
  wire g539_p_spl_;
  wire g541_p_spl_;
  wire g541_p_spl_0;
  wire n2851_lo_p_spl_;
  wire n2851_lo_p_spl_0;
  wire n2851_lo_p_spl_00;
  wire n2851_lo_p_spl_1;
  wire n2623_lo_p_spl_;
  wire n2851_lo_n_spl_;
  wire n2851_lo_n_spl_0;
  wire n2851_lo_n_spl_00;
  wire n2851_lo_n_spl_1;
  wire n2623_lo_n_spl_;
  wire g546_n_spl_;
  wire g545_n_spl_;
  wire g546_p_spl_;
  wire g545_p_spl_;
  wire g547_n_spl_;
  wire g547_n_spl_0;
  wire g547_p_spl_;
  wire g547_p_spl_0;
  wire g551_n_spl_;
  wire g550_n_spl_;
  wire g551_p_spl_;
  wire g550_p_spl_;
  wire g552_n_spl_;
  wire g552_n_spl_0;
  wire g552_p_spl_;
  wire g552_p_spl_0;
  wire g556_n_spl_;
  wire g555_n_spl_;
  wire g556_p_spl_;
  wire g555_p_spl_;
  wire g557_n_spl_;
  wire g557_n_spl_0;
  wire g557_p_spl_;
  wire g557_p_spl_0;
  wire g561_n_spl_;
  wire g560_n_spl_;
  wire g561_p_spl_;
  wire g560_p_spl_;
  wire g562_n_spl_;
  wire g562_n_spl_0;
  wire g562_p_spl_;
  wire g562_p_spl_0;
  wire g566_p_spl_;
  wire g565_p_spl_;
  wire g567_p_spl_;
  wire g567_p_spl_0;
  wire G5044_o2_n_spl_;
  wire G5041_o2_n_spl_;
  wire G5044_o2_p_spl_;
  wire G5041_o2_p_spl_;
  wire g571_n_spl_;
  wire g571_n_spl_0;
  wire g571_p_spl_;
  wire g571_p_spl_0;
  wire n2635_lo_p_spl_;
  wire n2635_lo_n_spl_;
  wire g575_n_spl_;
  wire g574_n_spl_;
  wire g575_p_spl_;
  wire g574_p_spl_;
  wire g576_n_spl_;
  wire g576_n_spl_0;
  wire g576_p_spl_;
  wire g576_p_spl_0;
  wire g580_n_spl_;
  wire g579_n_spl_;
  wire g580_p_spl_;
  wire g579_p_spl_;
  wire g581_n_spl_;
  wire g581_n_spl_0;
  wire g581_p_spl_;
  wire g581_p_spl_0;
  wire g585_n_spl_;
  wire g584_n_spl_;
  wire g585_p_spl_;
  wire g584_p_spl_;
  wire g586_n_spl_;
  wire g586_n_spl_0;
  wire g586_p_spl_;
  wire g586_p_spl_0;
  wire g590_n_spl_;
  wire g589_n_spl_;
  wire g590_p_spl_;
  wire g589_p_spl_;
  wire g591_n_spl_;
  wire g591_n_spl_0;
  wire g591_p_spl_;
  wire g591_p_spl_0;
  wire g595_p_spl_;
  wire g594_p_spl_;
  wire g596_p_spl_;
  wire g596_p_spl_0;
  wire G4864_o2_n_spl_;
  wire G4864_o2_n_spl_0;
  wire G4864_o2_p_spl_;
  wire G4864_o2_p_spl_0;
  wire g603_n_spl_;
  wire g602_n_spl_;
  wire g603_p_spl_;
  wire g602_p_spl_;
  wire g604_n_spl_;
  wire g604_n_spl_0;
  wire g604_p_spl_;
  wire g604_p_spl_0;
  wire n2647_lo_p_spl_;
  wire n2647_lo_n_spl_;
  wire g608_n_spl_;
  wire g607_n_spl_;
  wire g608_p_spl_;
  wire g607_p_spl_;
  wire g609_n_spl_;
  wire g609_n_spl_0;
  wire g609_p_spl_;
  wire g609_p_spl_0;
  wire g613_n_spl_;
  wire g612_n_spl_;
  wire g613_p_spl_;
  wire g612_p_spl_;
  wire g614_n_spl_;
  wire g614_n_spl_0;
  wire g614_p_spl_;
  wire g614_p_spl_0;
  wire g618_n_spl_;
  wire g617_n_spl_;
  wire g618_p_spl_;
  wire g617_p_spl_;
  wire g619_n_spl_;
  wire g619_n_spl_0;
  wire g619_p_spl_;
  wire g619_p_spl_0;
  wire g623_n_spl_;
  wire g622_n_spl_;
  wire g623_p_spl_;
  wire g622_p_spl_;
  wire g624_n_spl_;
  wire g624_n_spl_0;
  wire g624_p_spl_;
  wire g624_p_spl_0;
  wire g628_p_spl_;
  wire g627_p_spl_;
  wire g629_p_spl_;
  wire g629_p_spl_0;
  wire n2671_lo_p_spl_;
  wire n2671_lo_p_spl_0;
  wire n2671_lo_n_spl_;
  wire n2671_lo_n_spl_0;
  wire g634_n_spl_;
  wire g633_n_spl_;
  wire g634_p_spl_;
  wire g633_p_spl_;
  wire g635_n_spl_;
  wire g635_n_spl_0;
  wire g635_p_spl_;
  wire g635_p_spl_0;
  wire n2659_lo_p_spl_;
  wire n2659_lo_n_spl_;
  wire g639_n_spl_;
  wire g638_n_spl_;
  wire g639_p_spl_;
  wire g638_p_spl_;
  wire g640_n_spl_;
  wire g640_n_spl_0;
  wire g640_p_spl_;
  wire g640_p_spl_0;
  wire g644_n_spl_;
  wire g643_n_spl_;
  wire g644_p_spl_;
  wire g643_p_spl_;
  wire g645_n_spl_;
  wire g645_n_spl_0;
  wire g645_p_spl_;
  wire g645_p_spl_0;
  wire g649_n_spl_;
  wire g648_n_spl_;
  wire g649_p_spl_;
  wire g648_p_spl_;
  wire g650_n_spl_;
  wire g650_n_spl_0;
  wire g650_p_spl_;
  wire g650_p_spl_0;
  wire g654_n_spl_;
  wire g653_n_spl_;
  wire g654_p_spl_;
  wire g653_p_spl_;
  wire g655_n_spl_;
  wire g655_n_spl_0;
  wire g655_p_spl_;
  wire g655_p_spl_0;
  wire g659_p_spl_;
  wire g658_p_spl_;
  wire g660_p_spl_;
  wire g660_p_spl_0;
  wire g665_n_spl_;
  wire g664_n_spl_;
  wire g665_p_spl_;
  wire g664_p_spl_;
  wire g666_n_spl_;
  wire g666_n_spl_0;
  wire g666_p_spl_;
  wire g666_p_spl_0;
  wire g670_n_spl_;
  wire g669_n_spl_;
  wire g670_p_spl_;
  wire g669_p_spl_;
  wire g671_n_spl_;
  wire g671_n_spl_0;
  wire g671_p_spl_;
  wire g671_p_spl_0;
  wire g675_n_spl_;
  wire g674_n_spl_;
  wire g675_p_spl_;
  wire g674_p_spl_;
  wire g676_n_spl_;
  wire g676_n_spl_0;
  wire g676_p_spl_;
  wire g676_p_spl_0;
  wire g680_p_spl_;
  wire g679_p_spl_;
  wire g681_p_spl_;
  wire g681_p_spl_0;
  wire g686_n_spl_;
  wire g685_n_spl_;
  wire g686_p_spl_;
  wire g685_p_spl_;
  wire g687_n_spl_;
  wire g687_n_spl_0;
  wire g687_p_spl_;
  wire g692_n_spl_;
  wire g692_n_spl_0;
  wire n2824_lo_buf_o2_p_spl_;
  wire n2824_lo_buf_o2_p_spl_0;
  wire n2824_lo_buf_o2_p_spl_00;
  wire n2824_lo_buf_o2_p_spl_000;
  wire n2824_lo_buf_o2_p_spl_001;
  wire n2824_lo_buf_o2_p_spl_01;
  wire n2824_lo_buf_o2_p_spl_010;
  wire n2824_lo_buf_o2_p_spl_1;
  wire n2824_lo_buf_o2_p_spl_10;
  wire n2824_lo_buf_o2_p_spl_11;
  wire n6461_o2_p_spl_;
  wire n6461_o2_p_spl_0;
  wire n6461_o2_p_spl_00;
  wire n6461_o2_p_spl_1;
  wire n2824_lo_buf_o2_n_spl_;
  wire n2824_lo_buf_o2_n_spl_0;
  wire n2824_lo_buf_o2_n_spl_00;
  wire n2824_lo_buf_o2_n_spl_000;
  wire n2824_lo_buf_o2_n_spl_001;
  wire n2824_lo_buf_o2_n_spl_01;
  wire n2824_lo_buf_o2_n_spl_010;
  wire n2824_lo_buf_o2_n_spl_1;
  wire n2824_lo_buf_o2_n_spl_10;
  wire n2824_lo_buf_o2_n_spl_11;
  wire n6461_o2_n_spl_;
  wire n6461_o2_n_spl_0;
  wire n6461_o2_n_spl_1;
  wire g698_n_spl_;
  wire g697_p_spl_;
  wire n2836_lo_p_spl_;
  wire n2836_lo_p_spl_0;
  wire n2836_lo_p_spl_00;
  wire n2836_lo_p_spl_000;
  wire n2836_lo_p_spl_001;
  wire n2836_lo_p_spl_01;
  wire n2836_lo_p_spl_010;
  wire n2836_lo_p_spl_011;
  wire n2836_lo_p_spl_1;
  wire n2836_lo_p_spl_10;
  wire n2836_lo_p_spl_100;
  wire n2836_lo_p_spl_101;
  wire n2836_lo_p_spl_11;
  wire n2836_lo_p_spl_110;
  wire n2836_lo_n_spl_;
  wire n2836_lo_n_spl_0;
  wire n2836_lo_n_spl_00;
  wire n2836_lo_n_spl_000;
  wire n2836_lo_n_spl_001;
  wire n2836_lo_n_spl_01;
  wire n2836_lo_n_spl_010;
  wire n2836_lo_n_spl_011;
  wire n2836_lo_n_spl_1;
  wire n2836_lo_n_spl_10;
  wire n2836_lo_n_spl_100;
  wire n2836_lo_n_spl_101;
  wire n2836_lo_n_spl_11;
  wire n2836_lo_n_spl_110;
  wire G5109_o2_p_spl_;
  wire G626_o2_n_spl_;
  wire G5109_o2_n_spl_;
  wire G626_o2_p_spl_;
  wire g701_n_spl_;
  wire g701_n_spl_0;
  wire g701_p_spl_;
  wire g701_p_spl_0;
  wire g699_p_spl_;
  wire g705_n_spl_;
  wire g704_n_spl_;
  wire g705_p_spl_;
  wire g704_p_spl_;
  wire g706_n_spl_;
  wire g706_n_spl_0;
  wire g706_p_spl_;
  wire g706_p_spl_0;
  wire g709_n_spl_;
  wire g700_p_spl_;
  wire n2848_lo_p_spl_;
  wire n2848_lo_p_spl_0;
  wire n2848_lo_p_spl_00;
  wire n2848_lo_p_spl_000;
  wire n2848_lo_p_spl_001;
  wire n2848_lo_p_spl_01;
  wire n2848_lo_p_spl_010;
  wire n2848_lo_p_spl_1;
  wire n2848_lo_p_spl_10;
  wire n2848_lo_p_spl_11;
  wire n2848_lo_n_spl_;
  wire n2848_lo_n_spl_0;
  wire n2848_lo_n_spl_00;
  wire n2848_lo_n_spl_000;
  wire n2848_lo_n_spl_001;
  wire n2848_lo_n_spl_01;
  wire n2848_lo_n_spl_010;
  wire n2848_lo_n_spl_1;
  wire n2848_lo_n_spl_10;
  wire n2848_lo_n_spl_11;
  wire G5172_o2_n_spl_;
  wire G5172_o2_n_spl_0;
  wire G5172_o2_p_spl_;
  wire G5172_o2_p_spl_0;
  wire g715_n_spl_;
  wire g714_n_spl_;
  wire g715_p_spl_;
  wire g714_p_spl_;
  wire g716_n_spl_;
  wire g716_n_spl_0;
  wire g716_p_spl_;
  wire g716_p_spl_0;
  wire n6309_o2_p_spl_;
  wire n6309_o2_p_spl_0;
  wire n6309_o2_n_spl_;
  wire n6309_o2_n_spl_0;
  wire g720_n_spl_;
  wire g719_n_spl_;
  wire g720_p_spl_;
  wire g719_p_spl_;
  wire g721_n_spl_;
  wire g721_n_spl_0;
  wire g721_p_spl_;
  wire g721_p_spl_0;
  wire g710_p_spl_;
  wire g725_n_spl_;
  wire g724_n_spl_;
  wire g725_p_spl_;
  wire g724_p_spl_;
  wire g726_n_spl_;
  wire g726_n_spl_0;
  wire g726_p_spl_;
  wire g726_p_spl_0;
  wire g729_n_spl_;
  wire g711_p_spl_;
  wire n2764_lo_buf_o2_p_spl_;
  wire n2764_lo_buf_o2_p_spl_0;
  wire n2764_lo_buf_o2_p_spl_00;
  wire n2764_lo_buf_o2_p_spl_1;
  wire n8086_o2_p_spl_;
  wire n8086_o2_p_spl_0;
  wire n8086_o2_p_spl_00;
  wire n8086_o2_p_spl_01;
  wire n8086_o2_p_spl_1;
  wire n2764_lo_buf_o2_n_spl_;
  wire n2764_lo_buf_o2_n_spl_0;
  wire n2764_lo_buf_o2_n_spl_00;
  wire n2764_lo_buf_o2_n_spl_1;
  wire n8086_o2_n_spl_;
  wire n8086_o2_n_spl_0;
  wire n8086_o2_n_spl_00;
  wire n8086_o2_n_spl_1;
  wire G3257_o2_p_spl_;
  wire G3257_o2_p_spl_0;
  wire G3257_o2_n_spl_;
  wire G3257_o2_n_spl_0;
  wire g734_n_spl_;
  wire g731_p_spl_;
  wire n2860_lo_p_spl_;
  wire n2860_lo_p_spl_0;
  wire n2860_lo_p_spl_00;
  wire n2860_lo_p_spl_01;
  wire n2860_lo_p_spl_1;
  wire n2860_lo_p_spl_10;
  wire n2860_lo_n_spl_;
  wire n2860_lo_n_spl_0;
  wire n2860_lo_n_spl_00;
  wire n2860_lo_n_spl_01;
  wire n2860_lo_n_spl_1;
  wire n2860_lo_n_spl_10;
  wire g738_n_spl_;
  wire g737_n_spl_;
  wire g738_p_spl_;
  wire g737_p_spl_;
  wire g739_n_spl_;
  wire g739_n_spl_0;
  wire g739_p_spl_;
  wire g739_p_spl_0;
  wire n6239_o2_p_spl_;
  wire n6239_o2_p_spl_0;
  wire n6239_o2_n_spl_;
  wire n6239_o2_n_spl_0;
  wire g743_n_spl_;
  wire g742_n_spl_;
  wire g743_p_spl_;
  wire g742_p_spl_;
  wire g744_n_spl_;
  wire g744_n_spl_0;
  wire g744_p_spl_;
  wire g744_p_spl_0;
  wire g748_n_spl_;
  wire g747_n_spl_;
  wire g748_p_spl_;
  wire g747_p_spl_;
  wire g749_n_spl_;
  wire g749_n_spl_0;
  wire g749_p_spl_;
  wire g749_p_spl_0;
  wire g753_n_spl_;
  wire g752_n_spl_;
  wire g753_p_spl_;
  wire g752_p_spl_;
  wire g754_n_spl_;
  wire g754_n_spl_0;
  wire g754_p_spl_;
  wire g754_p_spl_0;
  wire g730_p_spl_;
  wire g758_n_spl_;
  wire g757_n_spl_;
  wire g758_p_spl_;
  wire g757_p_spl_;
  wire g759_n_spl_;
  wire g759_n_spl_0;
  wire g759_p_spl_;
  wire g759_p_spl_0;
  wire n2776_lo_buf_o2_p_spl_;
  wire n2776_lo_buf_o2_p_spl_0;
  wire n2776_lo_buf_o2_p_spl_00;
  wire n2776_lo_buf_o2_p_spl_000;
  wire n2776_lo_buf_o2_p_spl_001;
  wire n2776_lo_buf_o2_p_spl_01;
  wire n2776_lo_buf_o2_p_spl_010;
  wire n2776_lo_buf_o2_p_spl_011;
  wire n2776_lo_buf_o2_p_spl_1;
  wire n2776_lo_buf_o2_p_spl_10;
  wire n2776_lo_buf_o2_p_spl_100;
  wire n2776_lo_buf_o2_p_spl_101;
  wire n2776_lo_buf_o2_p_spl_11;
  wire n2776_lo_buf_o2_n_spl_;
  wire n2776_lo_buf_o2_n_spl_0;
  wire n2776_lo_buf_o2_n_spl_00;
  wire n2776_lo_buf_o2_n_spl_000;
  wire n2776_lo_buf_o2_n_spl_001;
  wire n2776_lo_buf_o2_n_spl_01;
  wire n2776_lo_buf_o2_n_spl_010;
  wire n2776_lo_buf_o2_n_spl_011;
  wire n2776_lo_buf_o2_n_spl_1;
  wire n2776_lo_buf_o2_n_spl_10;
  wire n2776_lo_buf_o2_n_spl_100;
  wire n2776_lo_buf_o2_n_spl_101;
  wire n2776_lo_buf_o2_n_spl_11;
  wire g762_n_spl_;
  wire g736_p_spl_;
  wire n7909_o2_p_spl_;
  wire n7909_o2_p_spl_0;
  wire n7909_o2_p_spl_00;
  wire n7909_o2_p_spl_01;
  wire n7909_o2_p_spl_1;
  wire n7909_o2_p_spl_10;
  wire n7909_o2_n_spl_;
  wire n7909_o2_n_spl_0;
  wire n7909_o2_n_spl_00;
  wire n7909_o2_n_spl_1;
  wire g766_n_spl_;
  wire g765_n_spl_;
  wire g766_p_spl_;
  wire g765_p_spl_;
  wire g767_n_spl_;
  wire g767_n_spl_0;
  wire g767_p_spl_;
  wire g767_p_spl_0;
  wire g735_p_spl_;
  wire g771_n_spl_;
  wire g770_n_spl_;
  wire g771_p_spl_;
  wire g770_p_spl_;
  wire g772_n_spl_;
  wire g772_n_spl_0;
  wire g772_p_spl_;
  wire g772_p_spl_0;
  wire g775_n_spl_;
  wire g763_p_spl_;
  wire n2488_lo_buf_o2_p_spl_;
  wire n2488_lo_buf_o2_p_spl_0;
  wire n2488_lo_buf_o2_p_spl_00;
  wire n2488_lo_buf_o2_p_spl_1;
  wire n2704_lo_buf_o2_p_spl_;
  wire n2704_lo_buf_o2_p_spl_0;
  wire n2488_lo_buf_o2_n_spl_;
  wire n2488_lo_buf_o2_n_spl_0;
  wire n2488_lo_buf_o2_n_spl_00;
  wire n2488_lo_buf_o2_n_spl_1;
  wire n2704_lo_buf_o2_n_spl_;
  wire n2704_lo_buf_o2_n_spl_0;
  wire G1580_o2_n_spl_;
  wire G1507_o2_n_spl_;
  wire G1580_o2_p_spl_;
  wire G1507_o2_p_spl_;
  wire g778_n_spl_;
  wire g778_n_spl_0;
  wire g778_p_spl_;
  wire g778_p_spl_0;
  wire n2785_lo_p_spl_;
  wire n2785_lo_p_spl_0;
  wire n2785_lo_p_spl_00;
  wire n2785_lo_p_spl_000;
  wire n2785_lo_p_spl_001;
  wire n2785_lo_p_spl_01;
  wire n2785_lo_p_spl_010;
  wire n2785_lo_p_spl_011;
  wire n2785_lo_p_spl_1;
  wire n2785_lo_p_spl_10;
  wire n2785_lo_p_spl_100;
  wire n2785_lo_p_spl_101;
  wire n2785_lo_p_spl_11;
  wire n2785_lo_p_spl_110;
  wire n2785_lo_p_spl_111;
  wire n2785_lo_n_spl_;
  wire n2785_lo_n_spl_0;
  wire n2785_lo_n_spl_00;
  wire n2785_lo_n_spl_000;
  wire n2785_lo_n_spl_001;
  wire n2785_lo_n_spl_01;
  wire n2785_lo_n_spl_010;
  wire n2785_lo_n_spl_011;
  wire n2785_lo_n_spl_1;
  wire n2785_lo_n_spl_10;
  wire n2785_lo_n_spl_100;
  wire n2785_lo_n_spl_101;
  wire n2785_lo_n_spl_11;
  wire n2785_lo_n_spl_110;
  wire n2785_lo_n_spl_111;
  wire g781_n_spl_;
  wire g777_p_spl_;
  wire G3364_o2_p_spl_;
  wire G659_o2_n_spl_;
  wire G3364_o2_n_spl_;
  wire G659_o2_p_spl_;
  wire g784_n_spl_;
  wire g784_n_spl_0;
  wire g784_p_spl_;
  wire g784_p_spl_0;
  wire g788_n_spl_;
  wire g787_n_spl_;
  wire g788_p_spl_;
  wire g787_p_spl_;
  wire g789_n_spl_;
  wire g789_n_spl_0;
  wire g789_p_spl_;
  wire g789_p_spl_0;
  wire g793_n_spl_;
  wire g792_n_spl_;
  wire g793_p_spl_;
  wire g792_p_spl_;
  wire g794_n_spl_;
  wire g794_n_spl_0;
  wire g794_p_spl_;
  wire g794_p_spl_0;
  wire g776_p_spl_;
  wire g798_n_spl_;
  wire g797_n_spl_;
  wire g798_p_spl_;
  wire g797_p_spl_;
  wire g799_n_spl_;
  wire g799_n_spl_0;
  wire g799_p_spl_;
  wire g799_p_spl_0;
  wire g802_n_spl_;
  wire g782_p_spl_;
  wire n2716_lo_buf_o2_p_spl_;
  wire n2716_lo_buf_o2_p_spl_0;
  wire n2716_lo_buf_o2_p_spl_00;
  wire n2716_lo_buf_o2_p_spl_000;
  wire n2716_lo_buf_o2_p_spl_01;
  wire n2716_lo_buf_o2_p_spl_1;
  wire n2716_lo_buf_o2_p_spl_10;
  wire n2716_lo_buf_o2_p_spl_11;
  wire n2716_lo_buf_o2_n_spl_;
  wire n2716_lo_buf_o2_n_spl_0;
  wire n2716_lo_buf_o2_n_spl_00;
  wire n2716_lo_buf_o2_n_spl_000;
  wire n2716_lo_buf_o2_n_spl_01;
  wire n2716_lo_buf_o2_n_spl_1;
  wire n2716_lo_buf_o2_n_spl_10;
  wire n2716_lo_buf_o2_n_spl_11;
  wire G1630_o2_p_spl_;
  wire G1630_o2_p_spl_0;
  wire G1630_o2_n_spl_;
  wire G1630_o2_n_spl_0;
  wire n2500_lo_buf_o2_p_spl_;
  wire n2500_lo_buf_o2_p_spl_0;
  wire n2500_lo_buf_o2_p_spl_00;
  wire n2500_lo_buf_o2_p_spl_01;
  wire n2500_lo_buf_o2_p_spl_1;
  wire n2500_lo_buf_o2_n_spl_;
  wire n2500_lo_buf_o2_n_spl_0;
  wire n2500_lo_buf_o2_n_spl_00;
  wire n2500_lo_buf_o2_n_spl_1;
  wire g808_n_spl_;
  wire g807_n_spl_;
  wire g808_p_spl_;
  wire g807_p_spl_;
  wire g809_n_spl_;
  wire g809_n_spl_0;
  wire g809_p_spl_;
  wire g809_p_spl_0;
  wire g783_p_spl_;
  wire g813_n_spl_;
  wire g812_n_spl_;
  wire g813_p_spl_;
  wire g812_p_spl_;
  wire g814_n_spl_;
  wire g814_n_spl_0;
  wire g814_p_spl_;
  wire g814_p_spl_0;
  wire n2812_lo_buf_o2_p_spl_;
  wire n2812_lo_buf_o2_p_spl_0;
  wire n2812_lo_buf_o2_p_spl_00;
  wire n2812_lo_buf_o2_p_spl_01;
  wire n2812_lo_buf_o2_p_spl_1;
  wire n5779_o2_p_spl_;
  wire n5779_o2_p_spl_0;
  wire n5779_o2_p_spl_1;
  wire n2812_lo_buf_o2_n_spl_;
  wire n2812_lo_buf_o2_n_spl_0;
  wire n2812_lo_buf_o2_n_spl_00;
  wire n2812_lo_buf_o2_n_spl_01;
  wire n2812_lo_buf_o2_n_spl_1;
  wire n5779_o2_n_spl_;
  wire n5779_o2_n_spl_0;
  wire n2800_lo_buf_o2_p_spl_;
  wire n2800_lo_buf_o2_n_spl_;
  wire n5792_o2_p_spl_;
  wire n5792_o2_p_spl_0;
  wire n5792_o2_p_spl_1;
  wire n5792_o2_n_spl_;
  wire n5792_o2_n_spl_0;
  wire n5792_o2_n_spl_1;
  wire g821_n_spl_;
  wire g820_n_spl_;
  wire g821_p_spl_;
  wire g820_p_spl_;
  wire g822_n_spl_;
  wire g822_n_spl_0;
  wire g822_p_spl_;
  wire g822_p_spl_0;
  wire g823_n_spl_;
  wire g819_n_spl_;
  wire g823_p_spl_;
  wire g819_p_spl_;
  wire g824_n_spl_;
  wire g824_n_spl_0;
  wire g824_p_spl_;
  wire g824_p_spl_0;
  wire g828_n_spl_;
  wire g827_n_spl_;
  wire g828_p_spl_;
  wire g827_p_spl_;
  wire g829_n_spl_;
  wire g829_n_spl_0;
  wire g829_p_spl_;
  wire g829_p_spl_0;
  wire g830_n_spl_;
  wire g818_n_spl_;
  wire g830_p_spl_;
  wire g818_p_spl_;
  wire g831_n_spl_;
  wire g831_n_spl_0;
  wire g831_p_spl_;
  wire g831_p_spl_0;
  wire g835_n_spl_;
  wire g834_n_spl_;
  wire g835_p_spl_;
  wire g834_p_spl_;
  wire g836_n_spl_;
  wire g836_n_spl_0;
  wire g836_p_spl_;
  wire g836_p_spl_0;
  wire G4034_o2_n_spl_;
  wire G4034_o2_n_spl_0;
  wire G4034_o2_p_spl_;
  wire G4034_o2_p_spl_0;
  wire g846_n_spl_;
  wire g845_n_spl_;
  wire g846_p_spl_;
  wire g845_p_spl_;
  wire g847_n_spl_;
  wire g847_n_spl_0;
  wire g847_p_spl_;
  wire g847_p_spl_0;
  wire n5842_o2_p_spl_;
  wire n5842_o2_p_spl_0;
  wire n5842_o2_p_spl_1;
  wire n5842_o2_n_spl_;
  wire n5842_o2_n_spl_0;
  wire g851_n_spl_;
  wire g850_n_spl_;
  wire g851_p_spl_;
  wire g850_p_spl_;
  wire g852_n_spl_;
  wire g852_n_spl_0;
  wire g852_p_spl_;
  wire g852_p_spl_0;
  wire g853_n_spl_;
  wire g842_n_spl_;
  wire g853_p_spl_;
  wire g842_p_spl_;
  wire g854_n_spl_;
  wire g854_n_spl_0;
  wire g854_p_spl_;
  wire g854_p_spl_0;
  wire g858_n_spl_;
  wire g857_n_spl_;
  wire g858_p_spl_;
  wire g857_p_spl_;
  wire g859_n_spl_;
  wire g859_n_spl_0;
  wire g859_p_spl_;
  wire g859_p_spl_0;
  wire g860_n_spl_;
  wire g839_n_spl_;
  wire g860_p_spl_;
  wire g839_p_spl_;
  wire g865_n_spl_;
  wire g864_n_spl_;
  wire g865_p_spl_;
  wire g864_p_spl_;
  wire g866_n_spl_;
  wire g866_n_spl_0;
  wire g866_p_spl_;
  wire g866_p_spl_0;
  wire n5863_o2_p_spl_;
  wire n5863_o2_p_spl_0;
  wire n5863_o2_p_spl_1;
  wire n5863_o2_n_spl_;
  wire n5863_o2_n_spl_0;
  wire g870_n_spl_;
  wire g869_n_spl_;
  wire g870_p_spl_;
  wire g869_p_spl_;
  wire g871_n_spl_;
  wire g871_n_spl_0;
  wire g871_p_spl_;
  wire g871_p_spl_0;
  wire G4220_o2_n_spl_;
  wire G4217_o2_n_spl_;
  wire G4220_o2_p_spl_;
  wire G4217_o2_p_spl_;
  wire g875_n_spl_;
  wire g875_n_spl_0;
  wire g875_p_spl_;
  wire g875_p_spl_0;
  wire n5881_o2_p_spl_;
  wire n5881_o2_p_spl_0;
  wire n5881_o2_p_spl_1;
  wire n5881_o2_n_spl_;
  wire n5881_o2_n_spl_0;
  wire g879_n_spl_;
  wire g878_n_spl_;
  wire g879_p_spl_;
  wire g878_p_spl_;
  wire g880_n_spl_;
  wire g880_n_spl_0;
  wire g880_p_spl_;
  wire g880_p_spl_0;
  wire g881_n_spl_;
  wire g874_n_spl_;
  wire g881_p_spl_;
  wire g874_p_spl_;
  wire g882_n_spl_;
  wire g882_n_spl_0;
  wire g882_p_spl_;
  wire g882_p_spl_0;
  wire g886_n_spl_;
  wire g885_n_spl_;
  wire g886_p_spl_;
  wire g885_p_spl_;
  wire g887_n_spl_;
  wire g887_n_spl_0;
  wire g887_p_spl_;
  wire g887_p_spl_0;
  wire n5930_o2_p_spl_;
  wire n5930_o2_p_spl_0;
  wire n5930_o2_p_spl_1;
  wire n5930_o2_n_spl_;
  wire n5930_o2_n_spl_0;
  wire n5930_o2_n_spl_1;
  wire g895_n_spl_;
  wire g894_n_spl_;
  wire g895_p_spl_;
  wire g894_p_spl_;
  wire g896_n_spl_;
  wire g896_n_spl_0;
  wire g896_p_spl_;
  wire g896_p_spl_0;
  wire g897_n_spl_;
  wire g893_n_spl_;
  wire g897_p_spl_;
  wire g893_p_spl_;
  wire g898_n_spl_;
  wire g898_n_spl_0;
  wire g898_p_spl_;
  wire g898_p_spl_0;
  wire g902_n_spl_;
  wire g901_n_spl_;
  wire g902_p_spl_;
  wire g901_p_spl_;
  wire g903_n_spl_;
  wire g903_n_spl_0;
  wire g903_p_spl_;
  wire g903_p_spl_0;
  wire g904_n_spl_;
  wire g890_n_spl_;
  wire g904_p_spl_;
  wire g890_p_spl_;
  wire g905_n_spl_;
  wire g905_n_spl_0;
  wire g905_p_spl_;
  wire g905_p_spl_0;
  wire g909_n_spl_;
  wire g908_n_spl_;
  wire g909_p_spl_;
  wire g908_p_spl_;
  wire g910_n_spl_;
  wire g910_n_spl_0;
  wire g910_p_spl_;
  wire g910_p_spl_0;
  wire G4556_o2_n_spl_;
  wire G4556_o2_n_spl_0;
  wire G4556_o2_p_spl_;
  wire G4556_o2_p_spl_0;
  wire g920_n_spl_;
  wire g919_n_spl_;
  wire g920_p_spl_;
  wire g919_p_spl_;
  wire g921_n_spl_;
  wire g921_n_spl_0;
  wire g921_p_spl_;
  wire g921_p_spl_0;
  wire n5959_o2_p_spl_;
  wire n5959_o2_p_spl_0;
  wire n5959_o2_p_spl_1;
  wire n5959_o2_n_spl_;
  wire n5959_o2_n_spl_0;
  wire g925_n_spl_;
  wire g924_n_spl_;
  wire g925_p_spl_;
  wire g924_p_spl_;
  wire g926_n_spl_;
  wire g926_n_spl_0;
  wire g926_p_spl_;
  wire g926_p_spl_0;
  wire g927_n_spl_;
  wire g916_n_spl_;
  wire g927_p_spl_;
  wire g916_p_spl_;
  wire g928_n_spl_;
  wire g928_n_spl_0;
  wire g928_p_spl_;
  wire g928_p_spl_0;
  wire g932_n_spl_;
  wire g931_n_spl_;
  wire g932_p_spl_;
  wire g931_p_spl_;
  wire g933_n_spl_;
  wire g933_n_spl_0;
  wire g933_p_spl_;
  wire g933_p_spl_0;
  wire g934_n_spl_;
  wire g913_n_spl_;
  wire g934_p_spl_;
  wire g913_p_spl_;
  wire g939_n_spl_;
  wire g938_n_spl_;
  wire g939_p_spl_;
  wire g938_p_spl_;
  wire g940_n_spl_;
  wire g940_n_spl_0;
  wire g940_p_spl_;
  wire g940_p_spl_0;
  wire n5981_o2_p_spl_;
  wire n5981_o2_p_spl_0;
  wire n5981_o2_p_spl_1;
  wire n5981_o2_n_spl_;
  wire n5981_o2_n_spl_0;
  wire g944_n_spl_;
  wire g943_n_spl_;
  wire g944_p_spl_;
  wire g943_p_spl_;
  wire g945_n_spl_;
  wire g945_n_spl_0;
  wire g945_p_spl_;
  wire g945_p_spl_0;
  wire G4719_o2_n_spl_;
  wire G4716_o2_n_spl_;
  wire G4719_o2_p_spl_;
  wire G4716_o2_p_spl_;
  wire g949_n_spl_;
  wire g949_n_spl_0;
  wire g949_p_spl_;
  wire g949_p_spl_0;
  wire n6042_o2_p_spl_;
  wire n6042_o2_p_spl_0;
  wire n6042_o2_p_spl_1;
  wire n6042_o2_n_spl_;
  wire n6042_o2_n_spl_0;
  wire g953_n_spl_;
  wire g952_n_spl_;
  wire g953_p_spl_;
  wire g952_p_spl_;
  wire g954_n_spl_;
  wire g954_n_spl_0;
  wire g954_p_spl_;
  wire g954_p_spl_0;
  wire g955_n_spl_;
  wire g948_n_spl_;
  wire g955_p_spl_;
  wire g948_p_spl_;
  wire g956_n_spl_;
  wire g956_n_spl_0;
  wire g956_p_spl_;
  wire g956_p_spl_0;
  wire g960_n_spl_;
  wire g959_n_spl_;
  wire g960_p_spl_;
  wire g959_p_spl_;
  wire g961_n_spl_;
  wire g961_n_spl_0;
  wire g961_p_spl_;
  wire g961_p_spl_0;
  wire n6075_o2_p_spl_;
  wire n6075_o2_p_spl_0;
  wire n6075_o2_n_spl_;
  wire n6075_o2_n_spl_0;
  wire n6075_o2_n_spl_1;
  wire g969_n_spl_;
  wire g968_n_spl_;
  wire g969_p_spl_;
  wire g968_p_spl_;
  wire g970_n_spl_;
  wire g970_n_spl_0;
  wire g970_p_spl_;
  wire g970_p_spl_0;
  wire g971_n_spl_;
  wire g967_n_spl_;
  wire g971_p_spl_;
  wire g967_p_spl_;
  wire g972_n_spl_;
  wire g972_n_spl_0;
  wire g972_p_spl_;
  wire g972_p_spl_0;
  wire g976_n_spl_;
  wire g975_n_spl_;
  wire g976_p_spl_;
  wire g975_p_spl_;
  wire g977_n_spl_;
  wire g977_n_spl_0;
  wire g977_p_spl_;
  wire g977_p_spl_0;
  wire g978_n_spl_;
  wire g964_n_spl_;
  wire g978_p_spl_;
  wire g964_p_spl_;
  wire g979_n_spl_;
  wire g979_n_spl_0;
  wire g979_p_spl_;
  wire g979_p_spl_0;
  wire g983_n_spl_;
  wire g982_n_spl_;
  wire g983_p_spl_;
  wire g982_p_spl_;
  wire g984_n_spl_;
  wire g984_n_spl_0;
  wire g984_p_spl_;
  wire g984_p_spl_0;
  wire G5064_o2_n_spl_;
  wire G5064_o2_n_spl_0;
  wire G5064_o2_p_spl_;
  wire G5064_o2_p_spl_0;
  wire g994_n_spl_;
  wire g993_n_spl_;
  wire g994_p_spl_;
  wire g993_p_spl_;
  wire g995_n_spl_;
  wire g995_n_spl_0;
  wire g995_p_spl_;
  wire g995_p_spl_0;
  wire n6103_o2_p_spl_;
  wire n6103_o2_p_spl_0;
  wire n6103_o2_n_spl_;
  wire n6103_o2_n_spl_0;
  wire g999_n_spl_;
  wire g998_n_spl_;
  wire g999_p_spl_;
  wire g998_p_spl_;
  wire g1000_n_spl_;
  wire g1000_n_spl_0;
  wire g1000_p_spl_;
  wire g1000_p_spl_0;
  wire g1001_n_spl_;
  wire g990_n_spl_;
  wire g1001_p_spl_;
  wire g990_p_spl_;
  wire g1002_n_spl_;
  wire g1002_n_spl_0;
  wire g1002_p_spl_;
  wire g1002_p_spl_0;
  wire g1006_n_spl_;
  wire g1005_n_spl_;
  wire g1006_p_spl_;
  wire g1005_p_spl_;
  wire g1007_n_spl_;
  wire g1007_n_spl_0;
  wire g1007_p_spl_;
  wire g1007_p_spl_0;
  wire g1008_n_spl_;
  wire g987_n_spl_;
  wire g1008_p_spl_;
  wire g987_p_spl_;
  wire G5247_o2_n_spl_;
  wire G5244_o2_n_spl_;
  wire G5247_o2_p_spl_;
  wire G5244_o2_p_spl_;
  wire g1010_n_spl_;
  wire g1010_n_spl_0;
  wire g1010_p_spl_;
  wire g1010_p_spl_0;
  wire n6205_o2_p_spl_;
  wire n6205_o2_p_spl_0;
  wire n6205_o2_n_spl_;
  wire n6205_o2_n_spl_0;
  wire g1014_n_spl_;
  wire g1013_n_spl_;
  wire g1014_p_spl_;
  wire g1013_p_spl_;
  wire g1015_n_spl_;
  wire g1015_n_spl_0;
  wire g1015_p_spl_;
  wire g1015_p_spl_0;
  wire g1019_n_spl_;
  wire g1018_n_spl_;
  wire g1019_p_spl_;
  wire g1018_p_spl_;
  wire g1020_n_spl_;
  wire g1020_n_spl_0;
  wire g1020_p_spl_;
  wire g1020_p_spl_0;
  wire g1024_n_spl_;
  wire g1023_n_spl_;
  wire g1024_p_spl_;
  wire g1023_p_spl_;
  wire g1025_n_spl_;
  wire g1025_n_spl_0;
  wire g1025_p_spl_;
  wire g1025_p_spl_0;
  wire g1029_n_spl_;
  wire g1028_n_spl_;
  wire g1029_p_spl_;
  wire g1028_p_spl_;
  wire g1030_n_spl_;
  wire g1030_n_spl_0;
  wire g1030_p_spl_;
  wire g1030_p_spl_0;
  wire g1034_n_spl_;
  wire g1033_n_spl_;
  wire g1034_p_spl_;
  wire g1033_p_spl_;
  wire g1035_n_spl_;
  wire g1035_n_spl_0;
  wire g1035_p_spl_;
  wire g1035_p_spl_0;
  wire g764_p_spl_;
  wire g1039_n_spl_;
  wire g1038_n_spl_;
  wire g1040_n_spl_;
  wire g817_n_spl_;
  wire g804_p_spl_;
  wire n2797_lo_p_spl_;
  wire n2797_lo_p_spl_0;
  wire n2797_lo_p_spl_00;
  wire n2797_lo_p_spl_000;
  wire n2797_lo_p_spl_001;
  wire n2797_lo_p_spl_01;
  wire n2797_lo_p_spl_010;
  wire n2797_lo_p_spl_011;
  wire n2797_lo_p_spl_1;
  wire n2797_lo_p_spl_10;
  wire n2797_lo_p_spl_100;
  wire n2797_lo_p_spl_101;
  wire n2797_lo_p_spl_11;
  wire n2797_lo_n_spl_;
  wire n2797_lo_n_spl_0;
  wire n2797_lo_n_spl_00;
  wire n2797_lo_n_spl_000;
  wire n2797_lo_n_spl_001;
  wire n2797_lo_n_spl_01;
  wire n2797_lo_n_spl_010;
  wire n2797_lo_n_spl_011;
  wire n2797_lo_n_spl_1;
  wire n2797_lo_n_spl_10;
  wire n2797_lo_n_spl_100;
  wire n2797_lo_n_spl_101;
  wire n2797_lo_n_spl_11;
  wire G3422_o2_n_spl_;
  wire G3422_o2_n_spl_0;
  wire G3422_o2_p_spl_;
  wire G3422_o2_p_spl_0;
  wire g1049_n_spl_;
  wire g1048_n_spl_;
  wire g1049_p_spl_;
  wire g1048_p_spl_;
  wire g1050_n_spl_;
  wire g1050_n_spl_0;
  wire g1050_p_spl_;
  wire g1050_p_spl_0;
  wire n7835_o2_p_spl_;
  wire n7835_o2_p_spl_0;
  wire n7835_o2_p_spl_00;
  wire n7835_o2_p_spl_1;
  wire n7835_o2_n_spl_;
  wire n7835_o2_n_spl_0;
  wire n7835_o2_n_spl_00;
  wire n7835_o2_n_spl_1;
  wire g1054_n_spl_;
  wire g1053_n_spl_;
  wire g1054_p_spl_;
  wire g1053_p_spl_;
  wire g1055_n_spl_;
  wire g1055_n_spl_0;
  wire g1055_p_spl_;
  wire g1055_p_spl_0;
  wire g1059_n_spl_;
  wire g1058_n_spl_;
  wire g1059_p_spl_;
  wire g1058_p_spl_;
  wire g1060_n_spl_;
  wire g1060_n_spl_0;
  wire g1060_p_spl_;
  wire g1060_p_spl_0;
  wire g1064_n_spl_;
  wire g1063_n_spl_;
  wire g1064_p_spl_;
  wire g1063_p_spl_;
  wire g1065_n_spl_;
  wire g1065_n_spl_0;
  wire g1065_p_spl_;
  wire g1065_p_spl_0;
  wire g803_p_spl_;
  wire g1069_n_spl_;
  wire g1068_n_spl_;
  wire g1069_p_spl_;
  wire g1068_p_spl_;
  wire g1070_n_spl_;
  wire g1070_n_spl_0;
  wire g1070_p_spl_;
  wire g1070_p_spl_0;
  wire n2728_lo_buf_o2_p_spl_;
  wire n2728_lo_buf_o2_p_spl_0;
  wire n2728_lo_buf_o2_p_spl_00;
  wire n2728_lo_buf_o2_p_spl_000;
  wire n2728_lo_buf_o2_p_spl_001;
  wire n2728_lo_buf_o2_p_spl_01;
  wire n2728_lo_buf_o2_p_spl_010;
  wire n2728_lo_buf_o2_p_spl_011;
  wire n2728_lo_buf_o2_p_spl_1;
  wire n2728_lo_buf_o2_p_spl_10;
  wire n2728_lo_buf_o2_p_spl_100;
  wire n2728_lo_buf_o2_p_spl_101;
  wire n2728_lo_buf_o2_p_spl_11;
  wire n2728_lo_buf_o2_p_spl_110;
  wire n2728_lo_buf_o2_p_spl_111;
  wire n2728_lo_buf_o2_n_spl_;
  wire n2728_lo_buf_o2_n_spl_0;
  wire n2728_lo_buf_o2_n_spl_00;
  wire n2728_lo_buf_o2_n_spl_000;
  wire n2728_lo_buf_o2_n_spl_001;
  wire n2728_lo_buf_o2_n_spl_01;
  wire n2728_lo_buf_o2_n_spl_010;
  wire n2728_lo_buf_o2_n_spl_011;
  wire n2728_lo_buf_o2_n_spl_1;
  wire n2728_lo_buf_o2_n_spl_10;
  wire n2728_lo_buf_o2_n_spl_100;
  wire n2728_lo_buf_o2_n_spl_101;
  wire n2728_lo_buf_o2_n_spl_11;
  wire n2728_lo_buf_o2_n_spl_110;
  wire n2728_lo_buf_o2_n_spl_111;
  wire g1073_n_spl_;
  wire g1045_p_spl_;
  wire n2512_lo_buf_o2_p_spl_;
  wire n2512_lo_buf_o2_p_spl_0;
  wire n2512_lo_buf_o2_p_spl_00;
  wire n2512_lo_buf_o2_p_spl_01;
  wire n2512_lo_buf_o2_p_spl_1;
  wire n2512_lo_buf_o2_p_spl_10;
  wire n2512_lo_buf_o2_n_spl_;
  wire n2512_lo_buf_o2_n_spl_0;
  wire n2512_lo_buf_o2_n_spl_00;
  wire n2512_lo_buf_o2_n_spl_1;
  wire g1077_n_spl_;
  wire g1076_n_spl_;
  wire g1077_p_spl_;
  wire g1076_p_spl_;
  wire g1078_n_spl_;
  wire g1078_n_spl_0;
  wire g1078_p_spl_;
  wire g1078_p_spl_0;
  wire g1082_n_spl_;
  wire g1081_n_spl_;
  wire g1082_p_spl_;
  wire g1081_p_spl_;
  wire g1083_n_spl_;
  wire g1083_n_spl_0;
  wire g1083_p_spl_;
  wire g1083_p_spl_0;
  wire g1087_n_spl_;
  wire g1086_n_spl_;
  wire g1087_p_spl_;
  wire g1086_p_spl_;
  wire g1088_n_spl_;
  wire g1088_n_spl_0;
  wire g1088_p_spl_;
  wire g1088_p_spl_0;
  wire g1044_p_spl_;
  wire g1092_n_spl_;
  wire g1091_n_spl_;
  wire g1092_p_spl_;
  wire g1091_p_spl_;
  wire g1093_n_spl_;
  wire g1093_n_spl_0;
  wire g1093_p_spl_;
  wire g1093_p_spl_0;
  wire g1096_n_spl_;
  wire g1074_p_spl_;
  wire g1043_n_spl_;
  wire g1043_n_spl_0;
  wire g1105_n_spl_;
  wire g1104_n_spl_;
  wire g1105_p_spl_;
  wire g1104_p_spl_;
  wire g1106_n_spl_;
  wire g1106_n_spl_0;
  wire g1106_p_spl_;
  wire g1106_p_spl_0;
  wire g1110_n_spl_;
  wire g1109_n_spl_;
  wire g1110_p_spl_;
  wire g1109_p_spl_;
  wire g1111_n_spl_;
  wire g1111_n_spl_0;
  wire g1111_p_spl_;
  wire g1111_p_spl_0;
  wire g1115_n_spl_;
  wire g1114_n_spl_;
  wire g1115_p_spl_;
  wire g1114_p_spl_;
  wire g1116_n_spl_;
  wire g1116_n_spl_0;
  wire g1116_p_spl_;
  wire g1116_p_spl_0;
  wire g1120_n_spl_;
  wire g1119_n_spl_;
  wire g1120_p_spl_;
  wire g1119_p_spl_;
  wire g1121_n_spl_;
  wire g1121_n_spl_0;
  wire g1121_p_spl_;
  wire g1121_p_spl_0;
  wire g1130_n_spl_;
  wire g1129_n_spl_;
  wire g1130_p_spl_;
  wire g1129_p_spl_;
  wire g1131_n_spl_;
  wire g1131_n_spl_0;
  wire g1131_p_spl_;
  wire g1131_p_spl_0;
  wire g1135_n_spl_;
  wire g1134_n_spl_;
  wire g1135_p_spl_;
  wire g1134_p_spl_;
  wire g1136_n_spl_;
  wire g1136_n_spl_0;
  wire g1136_p_spl_;
  wire g1136_p_spl_0;
  wire g1140_n_spl_;
  wire g1139_n_spl_;
  wire g1140_p_spl_;
  wire g1139_p_spl_;
  wire g1141_n_spl_;
  wire g1141_n_spl_0;
  wire g1141_p_spl_;
  wire g1141_p_spl_0;
  wire g1145_n_spl_;
  wire g1144_n_spl_;
  wire g1145_p_spl_;
  wire g1144_p_spl_;
  wire g1146_n_spl_;
  wire g1146_n_spl_0;
  wire g1146_p_spl_;
  wire g1146_p_spl_0;
  wire g1158_n_spl_;
  wire g1157_n_spl_;
  wire g1158_p_spl_;
  wire g1157_p_spl_;
  wire g1159_n_spl_;
  wire g1159_n_spl_0;
  wire g1159_p_spl_;
  wire g1159_p_spl_0;
  wire n6169_o2_p_spl_;
  wire n6169_o2_p_spl_0;
  wire n6169_o2_n_spl_;
  wire n6169_o2_n_spl_0;
  wire g1163_n_spl_;
  wire g1162_n_spl_;
  wire g1163_p_spl_;
  wire g1162_p_spl_;
  wire g1164_n_spl_;
  wire g1164_n_spl_0;
  wire g1164_p_spl_;
  wire g1164_p_spl_0;
  wire g1165_n_spl_;
  wire g1154_n_spl_;
  wire g1165_p_spl_;
  wire g1154_p_spl_;
  wire g1166_n_spl_;
  wire g1166_n_spl_0;
  wire g1166_p_spl_;
  wire g1166_p_spl_0;
  wire g1170_n_spl_;
  wire g1169_n_spl_;
  wire g1170_p_spl_;
  wire g1169_p_spl_;
  wire g1171_n_spl_;
  wire g1171_n_spl_0;
  wire g1171_p_spl_;
  wire g1171_p_spl_0;
  wire g1178_n_spl_;
  wire g1177_n_spl_;
  wire g1178_p_spl_;
  wire g1177_p_spl_;
  wire g1179_n_spl_;
  wire g1179_n_spl_0;
  wire g1179_p_spl_;
  wire g1179_p_spl_0;
  wire g1183_n_spl_;
  wire g1182_n_spl_;
  wire g1183_p_spl_;
  wire g1182_p_spl_;
  wire g1184_n_spl_;
  wire g1184_n_spl_0;
  wire g1184_p_spl_;
  wire g1184_p_spl_0;
  wire g1185_n_spl_;
  wire g1174_n_spl_;
  wire g1185_p_spl_;
  wire g1174_p_spl_;
  wire g1186_n_spl_;
  wire g1186_n_spl_0;
  wire g1186_p_spl_;
  wire g1186_p_spl_0;
  wire g1190_n_spl_;
  wire g1189_n_spl_;
  wire g1190_p_spl_;
  wire g1189_p_spl_;
  wire g1191_n_spl_;
  wire g1191_n_spl_0;
  wire g1191_p_spl_;
  wire g1191_p_spl_0;
  wire g1198_n_spl_;
  wire g1197_n_spl_;
  wire g1198_p_spl_;
  wire g1197_p_spl_;
  wire g1199_n_spl_;
  wire g1199_n_spl_0;
  wire g1199_p_spl_;
  wire g1199_p_spl_0;
  wire g1203_n_spl_;
  wire g1202_n_spl_;
  wire g1203_p_spl_;
  wire g1202_p_spl_;
  wire g1204_n_spl_;
  wire g1204_n_spl_0;
  wire g1204_p_spl_;
  wire g1204_p_spl_0;
  wire g1210_n_spl_;
  wire g1209_n_spl_;
  wire g1211_n_spl_;
  wire n2734_lo_p_spl_;
  wire n2734_lo_p_spl_0;
  wire n2734_lo_p_spl_00;
  wire n2734_lo_p_spl_000;
  wire n2734_lo_p_spl_001;
  wire n2734_lo_p_spl_01;
  wire n2734_lo_p_spl_010;
  wire n2734_lo_p_spl_011;
  wire n2734_lo_p_spl_1;
  wire n2734_lo_p_spl_10;
  wire n2734_lo_p_spl_100;
  wire n2734_lo_p_spl_101;
  wire n2734_lo_p_spl_11;
  wire n2734_lo_p_spl_110;
  wire n2734_lo_p_spl_111;
  wire n2734_lo_n_spl_;
  wire n2734_lo_n_spl_0;
  wire n2734_lo_n_spl_00;
  wire n2734_lo_n_spl_000;
  wire n2734_lo_n_spl_001;
  wire n2734_lo_n_spl_01;
  wire n2734_lo_n_spl_010;
  wire n2734_lo_n_spl_011;
  wire n2734_lo_n_spl_1;
  wire n2734_lo_n_spl_10;
  wire n2734_lo_n_spl_100;
  wire n2734_lo_n_spl_101;
  wire n2734_lo_n_spl_11;
  wire n2734_lo_n_spl_110;
  wire n2734_lo_n_spl_111;
  wire g1009_n_spl_;
  wire g1009_n_spl_0;
  wire g1009_p_spl_;
  wire g935_n_spl_;
  wire g935_n_spl_0;
  wire g935_p_spl_;
  wire g861_n_spl_;
  wire g861_n_spl_0;
  wire g861_p_spl_;
  wire g1214_n_spl_;
  wire g1098_n_spl_;
  wire n7148_o2_p_spl_;
  wire n7148_o2_p_spl_0;
  wire n7148_o2_p_spl_1;
  wire n7148_o2_n_spl_;
  wire n7148_o2_n_spl_0;
  wire G2917_o2_n_spl_;
  wire G1280_o2_n_spl_;
  wire G2917_o2_p_spl_;
  wire G1280_o2_p_spl_;
  wire g1233_n_spl_;
  wire g1233_n_spl_0;
  wire g1233_p_spl_;
  wire g1233_p_spl_0;
  wire n7224_o2_p_spl_;
  wire n7224_o2_p_spl_0;
  wire n7224_o2_p_spl_1;
  wire n7224_o2_n_spl_;
  wire n7224_o2_n_spl_0;
  wire g1237_n_spl_;
  wire g1236_n_spl_;
  wire g1237_p_spl_;
  wire g1236_p_spl_;
  wire g1238_n_spl_;
  wire g1238_n_spl_0;
  wire g1238_p_spl_;
  wire g1238_p_spl_0;
  wire g1239_n_spl_;
  wire g1232_n_spl_;
  wire g1239_p_spl_;
  wire g1232_p_spl_;
  wire g1240_n_spl_;
  wire g1240_n_spl_0;
  wire g1240_p_spl_;
  wire g1240_p_spl_0;
  wire g1244_n_spl_;
  wire g1243_n_spl_;
  wire g1244_p_spl_;
  wire g1243_p_spl_;
  wire g1245_n_spl_;
  wire g1245_n_spl_0;
  wire g1245_p_spl_;
  wire g1245_p_spl_0;
  wire n7280_o2_p_spl_;
  wire n7280_o2_p_spl_0;
  wire n7280_o2_p_spl_1;
  wire n7280_o2_n_spl_;
  wire n7280_o2_n_spl_0;
  wire n7280_o2_n_spl_1;
  wire g1253_n_spl_;
  wire g1252_n_spl_;
  wire g1253_p_spl_;
  wire g1252_p_spl_;
  wire g1254_n_spl_;
  wire g1254_n_spl_0;
  wire g1254_p_spl_;
  wire g1254_p_spl_0;
  wire g1255_n_spl_;
  wire g1251_n_spl_;
  wire g1255_p_spl_;
  wire g1251_p_spl_;
  wire g1256_n_spl_;
  wire g1256_n_spl_0;
  wire g1256_p_spl_;
  wire g1256_p_spl_0;
  wire g1260_n_spl_;
  wire g1259_n_spl_;
  wire g1260_p_spl_;
  wire g1259_p_spl_;
  wire g1261_n_spl_;
  wire g1261_n_spl_0;
  wire g1261_p_spl_;
  wire g1261_p_spl_0;
  wire g1262_n_spl_;
  wire g1248_n_spl_;
  wire g1262_p_spl_;
  wire g1248_p_spl_;
  wire g1263_n_spl_;
  wire g1263_n_spl_0;
  wire g1263_p_spl_;
  wire g1263_p_spl_0;
  wire g1267_n_spl_;
  wire g1266_n_spl_;
  wire g1267_p_spl_;
  wire g1266_p_spl_;
  wire g1268_n_spl_;
  wire g1268_n_spl_0;
  wire g1268_p_spl_;
  wire g1268_p_spl_0;
  wire G3241_o2_n_spl_;
  wire G3241_o2_n_spl_0;
  wire G3241_o2_p_spl_;
  wire G3241_o2_p_spl_0;
  wire g1278_n_spl_;
  wire g1277_n_spl_;
  wire g1278_p_spl_;
  wire g1277_p_spl_;
  wire g1279_n_spl_;
  wire g1279_n_spl_0;
  wire g1279_p_spl_;
  wire g1279_p_spl_0;
  wire n7313_o2_p_spl_;
  wire n7313_o2_p_spl_0;
  wire n7313_o2_p_spl_1;
  wire n7313_o2_n_spl_;
  wire n7313_o2_n_spl_0;
  wire g1283_n_spl_;
  wire g1282_n_spl_;
  wire g1283_p_spl_;
  wire g1282_p_spl_;
  wire g1284_n_spl_;
  wire g1284_n_spl_0;
  wire g1284_p_spl_;
  wire g1284_p_spl_0;
  wire g1285_n_spl_;
  wire g1274_n_spl_;
  wire g1285_p_spl_;
  wire g1274_p_spl_;
  wire g1286_n_spl_;
  wire g1286_n_spl_0;
  wire g1286_p_spl_;
  wire g1286_p_spl_0;
  wire g1290_n_spl_;
  wire g1289_n_spl_;
  wire g1290_p_spl_;
  wire g1289_p_spl_;
  wire g1291_n_spl_;
  wire g1291_n_spl_0;
  wire g1291_p_spl_;
  wire g1291_p_spl_0;
  wire g1292_n_spl_;
  wire g1271_n_spl_;
  wire g1292_p_spl_;
  wire g1271_p_spl_;
  wire g1297_n_spl_;
  wire g1296_n_spl_;
  wire g1297_p_spl_;
  wire g1296_p_spl_;
  wire g1298_n_spl_;
  wire g1298_n_spl_0;
  wire g1298_p_spl_;
  wire g1298_p_spl_0;
  wire n7323_o2_p_spl_;
  wire n7323_o2_p_spl_0;
  wire n7323_o2_p_spl_1;
  wire n7323_o2_n_spl_;
  wire n7323_o2_n_spl_0;
  wire g1302_n_spl_;
  wire g1301_n_spl_;
  wire g1302_p_spl_;
  wire g1301_p_spl_;
  wire g1303_n_spl_;
  wire g1303_n_spl_0;
  wire g1303_p_spl_;
  wire g1303_p_spl_0;
  wire G3394_o2_n_spl_;
  wire G3391_o2_n_spl_;
  wire G3394_o2_p_spl_;
  wire G3391_o2_p_spl_;
  wire g1307_n_spl_;
  wire g1307_n_spl_0;
  wire g1307_p_spl_;
  wire g1307_p_spl_0;
  wire n7398_o2_p_spl_;
  wire n7398_o2_p_spl_0;
  wire n7398_o2_p_spl_1;
  wire n7398_o2_n_spl_;
  wire n7398_o2_n_spl_0;
  wire g1311_n_spl_;
  wire g1310_n_spl_;
  wire g1311_p_spl_;
  wire g1310_p_spl_;
  wire g1312_n_spl_;
  wire g1312_n_spl_0;
  wire g1312_p_spl_;
  wire g1312_p_spl_0;
  wire g1313_n_spl_;
  wire g1306_n_spl_;
  wire g1313_p_spl_;
  wire g1306_p_spl_;
  wire g1314_n_spl_;
  wire g1314_n_spl_0;
  wire g1314_p_spl_;
  wire g1314_p_spl_0;
  wire g1318_n_spl_;
  wire g1317_n_spl_;
  wire g1318_p_spl_;
  wire g1317_p_spl_;
  wire g1319_n_spl_;
  wire g1319_n_spl_0;
  wire g1319_p_spl_;
  wire g1319_p_spl_0;
  wire n7459_o2_p_spl_;
  wire n7459_o2_p_spl_0;
  wire n7459_o2_p_spl_1;
  wire n7459_o2_n_spl_;
  wire n7459_o2_n_spl_0;
  wire n7459_o2_n_spl_1;
  wire g1327_n_spl_;
  wire g1326_n_spl_;
  wire g1327_p_spl_;
  wire g1326_p_spl_;
  wire g1328_n_spl_;
  wire g1328_n_spl_0;
  wire g1328_p_spl_;
  wire g1328_p_spl_0;
  wire g1329_n_spl_;
  wire g1325_n_spl_;
  wire g1329_p_spl_;
  wire g1325_p_spl_;
  wire g1330_n_spl_;
  wire g1330_n_spl_0;
  wire g1330_p_spl_;
  wire g1330_p_spl_0;
  wire g1334_n_spl_;
  wire g1333_n_spl_;
  wire g1334_p_spl_;
  wire g1333_p_spl_;
  wire g1335_n_spl_;
  wire g1335_n_spl_0;
  wire g1335_p_spl_;
  wire g1335_p_spl_0;
  wire g1336_n_spl_;
  wire g1322_n_spl_;
  wire g1336_p_spl_;
  wire g1322_p_spl_;
  wire g1337_n_spl_;
  wire g1337_n_spl_0;
  wire g1337_p_spl_;
  wire g1337_p_spl_0;
  wire g1341_n_spl_;
  wire g1340_n_spl_;
  wire g1341_p_spl_;
  wire g1340_p_spl_;
  wire g1342_n_spl_;
  wire g1342_n_spl_0;
  wire g1342_p_spl_;
  wire g1342_p_spl_0;
  wire G3722_o2_n_spl_;
  wire G3722_o2_n_spl_0;
  wire G3722_o2_p_spl_;
  wire G3722_o2_p_spl_0;
  wire g1352_n_spl_;
  wire g1351_n_spl_;
  wire g1352_p_spl_;
  wire g1351_p_spl_;
  wire g1353_n_spl_;
  wire g1353_n_spl_0;
  wire g1353_p_spl_;
  wire g1353_p_spl_0;
  wire n7501_o2_p_spl_;
  wire n7501_o2_p_spl_0;
  wire n7501_o2_p_spl_1;
  wire n7501_o2_n_spl_;
  wire n7501_o2_n_spl_0;
  wire g1357_n_spl_;
  wire g1356_n_spl_;
  wire g1357_p_spl_;
  wire g1356_p_spl_;
  wire g1358_n_spl_;
  wire g1358_n_spl_0;
  wire g1358_p_spl_;
  wire g1358_p_spl_0;
  wire g1359_n_spl_;
  wire g1348_n_spl_;
  wire g1359_p_spl_;
  wire g1348_p_spl_;
  wire g1360_n_spl_;
  wire g1360_n_spl_0;
  wire g1360_p_spl_;
  wire g1360_p_spl_0;
  wire g1364_n_spl_;
  wire g1363_n_spl_;
  wire g1364_p_spl_;
  wire g1363_p_spl_;
  wire g1365_n_spl_;
  wire g1365_n_spl_0;
  wire g1365_p_spl_;
  wire g1365_p_spl_0;
  wire g1366_n_spl_;
  wire g1345_n_spl_;
  wire g1366_p_spl_;
  wire g1345_p_spl_;
  wire G3719_o2_p_spl_;
  wire G902_o2_n_spl_;
  wire G3719_o2_n_spl_;
  wire G902_o2_p_spl_;
  wire g1371_n_spl_;
  wire g1371_n_spl_0;
  wire g1371_p_spl_;
  wire g1371_p_spl_0;
  wire g1372_n_spl_;
  wire g1370_n_spl_;
  wire g1372_p_spl_;
  wire g1370_p_spl_;
  wire g1373_n_spl_;
  wire g1373_n_spl_0;
  wire g1373_p_spl_;
  wire g1373_p_spl_0;
  wire n7518_o2_p_spl_;
  wire n7518_o2_p_spl_0;
  wire n7518_o2_p_spl_1;
  wire n7518_o2_n_spl_;
  wire n7518_o2_n_spl_0;
  wire g1377_n_spl_;
  wire g1376_n_spl_;
  wire g1377_p_spl_;
  wire g1376_p_spl_;
  wire g1378_n_spl_;
  wire g1378_n_spl_0;
  wire g1378_p_spl_;
  wire g1378_p_spl_0;
  wire n7606_o2_p_spl_;
  wire n7606_o2_p_spl_0;
  wire n7606_o2_p_spl_00;
  wire n7606_o2_p_spl_1;
  wire n7606_o2_n_spl_;
  wire n7606_o2_n_spl_0;
  wire n7606_o2_n_spl_1;
  wire g1386_n_spl_;
  wire g1385_n_spl_;
  wire g1386_p_spl_;
  wire g1385_p_spl_;
  wire g1387_n_spl_;
  wire g1387_n_spl_0;
  wire g1387_p_spl_;
  wire g1387_p_spl_0;
  wire g1388_n_spl_;
  wire g1384_n_spl_;
  wire g1388_p_spl_;
  wire g1384_p_spl_;
  wire g1389_n_spl_;
  wire g1389_n_spl_0;
  wire g1389_p_spl_;
  wire g1389_p_spl_0;
  wire g1393_n_spl_;
  wire g1392_n_spl_;
  wire g1393_p_spl_;
  wire g1392_p_spl_;
  wire g1394_n_spl_;
  wire g1394_n_spl_0;
  wire g1394_p_spl_;
  wire g1394_p_spl_0;
  wire g1395_n_spl_;
  wire g1381_n_spl_;
  wire g1395_p_spl_;
  wire g1381_p_spl_;
  wire g1396_n_spl_;
  wire g1396_n_spl_0;
  wire g1396_p_spl_;
  wire g1396_p_spl_0;
  wire g1400_n_spl_;
  wire g1399_n_spl_;
  wire g1400_p_spl_;
  wire g1399_p_spl_;
  wire g1401_n_spl_;
  wire g1401_n_spl_0;
  wire g1401_p_spl_;
  wire g1401_p_spl_0;
  wire G3616_o2_p_spl_;
  wire G3616_o2_p_spl_0;
  wire G3616_o2_n_spl_;
  wire G3616_o2_n_spl_0;
  wire n7675_o2_p_spl_;
  wire n7675_o2_p_spl_0;
  wire n7675_o2_p_spl_00;
  wire n7675_o2_p_spl_1;
  wire n7675_o2_n_spl_;
  wire n7675_o2_n_spl_0;
  wire n7675_o2_n_spl_00;
  wire n7675_o2_n_spl_1;
  wire g1414_n_spl_;
  wire g1413_n_spl_;
  wire g1414_p_spl_;
  wire g1413_p_spl_;
  wire g1415_n_spl_;
  wire g1415_n_spl_0;
  wire g1415_p_spl_;
  wire g1415_p_spl_0;
  wire g1416_n_spl_;
  wire g1410_n_spl_;
  wire g1416_p_spl_;
  wire g1410_p_spl_;
  wire g1417_n_spl_;
  wire g1417_n_spl_0;
  wire g1417_p_spl_;
  wire g1417_p_spl_0;
  wire g1421_n_spl_;
  wire g1420_n_spl_;
  wire g1421_p_spl_;
  wire g1420_p_spl_;
  wire g1422_n_spl_;
  wire g1422_n_spl_0;
  wire g1422_p_spl_;
  wire g1422_p_spl_0;
  wire g1423_n_spl_;
  wire g1407_n_spl_;
  wire g1423_p_spl_;
  wire g1407_p_spl_;
  wire g1424_n_spl_;
  wire g1424_n_spl_0;
  wire g1424_p_spl_;
  wire g1424_p_spl_0;
  wire g1428_n_spl_;
  wire g1427_n_spl_;
  wire g1428_p_spl_;
  wire g1427_p_spl_;
  wire g1429_n_spl_;
  wire g1429_n_spl_0;
  wire g1429_p_spl_;
  wire g1429_p_spl_0;
  wire g1430_n_spl_;
  wire g1404_n_spl_;
  wire g1430_p_spl_;
  wire g1404_p_spl_;
  wire g1431_n_spl_;
  wire g1431_n_spl_0;
  wire g1431_p_spl_;
  wire g1431_p_spl_0;
  wire n2809_lo_p_spl_;
  wire n2809_lo_p_spl_0;
  wire n2809_lo_p_spl_00;
  wire n2809_lo_p_spl_000;
  wire n2809_lo_p_spl_001;
  wire n2809_lo_p_spl_01;
  wire n2809_lo_p_spl_1;
  wire n2809_lo_p_spl_10;
  wire n2809_lo_p_spl_11;
  wire n2809_lo_n_spl_;
  wire n2809_lo_n_spl_0;
  wire n2809_lo_n_spl_00;
  wire n2809_lo_n_spl_000;
  wire n2809_lo_n_spl_001;
  wire n2809_lo_n_spl_01;
  wire n2809_lo_n_spl_1;
  wire n2809_lo_n_spl_10;
  wire n2809_lo_n_spl_11;
  wire g1435_n_spl_;
  wire g1434_n_spl_;
  wire g1435_p_spl_;
  wire g1434_p_spl_;
  wire g1436_n_spl_;
  wire g1436_n_spl_0;
  wire g1436_p_spl_;
  wire g1436_p_spl_0;
  wire G3557_o2_n_spl_;
  wire G3494_o2_n_spl_;
  wire G3557_o2_p_spl_;
  wire G3494_o2_p_spl_;
  wire g1449_n_spl_;
  wire g1449_n_spl_0;
  wire g1449_p_spl_;
  wire g1449_p_spl_0;
  wire n7722_o2_p_spl_;
  wire n7722_o2_p_spl_0;
  wire n7722_o2_p_spl_00;
  wire n7722_o2_p_spl_01;
  wire n7722_o2_p_spl_1;
  wire n7722_o2_n_spl_;
  wire n7722_o2_n_spl_0;
  wire n7722_o2_n_spl_00;
  wire n7722_o2_n_spl_1;
  wire g1453_n_spl_;
  wire g1452_n_spl_;
  wire g1453_p_spl_;
  wire g1452_p_spl_;
  wire g1454_n_spl_;
  wire g1454_n_spl_0;
  wire g1454_p_spl_;
  wire g1454_p_spl_0;
  wire g1455_n_spl_;
  wire g1448_n_spl_;
  wire g1455_p_spl_;
  wire g1448_p_spl_;
  wire g1456_n_spl_;
  wire g1456_n_spl_0;
  wire g1456_p_spl_;
  wire g1456_p_spl_0;
  wire g1460_n_spl_;
  wire g1459_n_spl_;
  wire g1460_p_spl_;
  wire g1459_p_spl_;
  wire g1461_n_spl_;
  wire g1461_n_spl_0;
  wire g1461_p_spl_;
  wire g1461_p_spl_0;
  wire g1462_n_spl_;
  wire g1445_n_spl_;
  wire g1462_p_spl_;
  wire g1445_p_spl_;
  wire g1463_n_spl_;
  wire g1463_n_spl_0;
  wire g1463_p_spl_;
  wire g1463_p_spl_0;
  wire g1467_n_spl_;
  wire g1466_n_spl_;
  wire g1467_p_spl_;
  wire g1466_p_spl_;
  wire g1468_n_spl_;
  wire g1468_n_spl_0;
  wire g1468_p_spl_;
  wire g1468_p_spl_0;
  wire g1469_n_spl_;
  wire g1442_n_spl_;
  wire g1469_p_spl_;
  wire g1442_p_spl_;
  wire g1470_n_spl_;
  wire g1470_n_spl_0;
  wire g1470_p_spl_;
  wire g1470_p_spl_0;
  wire g1474_n_spl_;
  wire g1473_n_spl_;
  wire g1474_p_spl_;
  wire g1473_p_spl_;
  wire g1475_n_spl_;
  wire g1475_n_spl_0;
  wire g1475_p_spl_;
  wire g1475_p_spl_0;
  wire g1476_n_spl_;
  wire g1439_n_spl_;
  wire g1476_p_spl_;
  wire g1439_p_spl_;
  wire G1724_o2_p_spl_;
  wire G692_o2_n_spl_;
  wire G1724_o2_n_spl_;
  wire G692_o2_p_spl_;
  wire g1478_n_spl_;
  wire g1478_n_spl_0;
  wire g1478_p_spl_;
  wire g1478_p_spl_0;
  wire g1482_n_spl_;
  wire g1481_n_spl_;
  wire g1482_p_spl_;
  wire g1481_p_spl_;
  wire g1483_n_spl_;
  wire g1483_n_spl_0;
  wire g1483_p_spl_;
  wire g1483_p_spl_0;
  wire g1487_n_spl_;
  wire g1486_n_spl_;
  wire g1487_p_spl_;
  wire g1486_p_spl_;
  wire g1488_n_spl_;
  wire g1488_n_spl_0;
  wire g1488_p_spl_;
  wire g1488_p_spl_0;
  wire g1492_n_spl_;
  wire g1491_n_spl_;
  wire g1492_p_spl_;
  wire g1491_p_spl_;
  wire g1493_n_spl_;
  wire g1493_n_spl_0;
  wire g1493_p_spl_;
  wire g1493_p_spl_0;
  wire g1497_n_spl_;
  wire g1496_n_spl_;
  wire g1497_p_spl_;
  wire g1496_p_spl_;
  wire g1498_n_spl_;
  wire g1498_n_spl_0;
  wire g1498_p_spl_;
  wire g1498_p_spl_0;
  wire g1097_p_spl_;
  wire g1502_n_spl_;
  wire g1501_n_spl_;
  wire g1502_p_spl_;
  wire g1501_p_spl_;
  wire g1503_n_spl_;
  wire g1503_n_spl_0;
  wire g1503_p_spl_;
  wire g1503_p_spl_0;
  wire g1506_n_spl_;
  wire g1215_p_spl_;
  wire g1510_n_spl_;
  wire g1509_n_spl_;
  wire g1510_p_spl_;
  wire g1509_p_spl_;
  wire g1511_n_spl_;
  wire g1511_n_spl_0;
  wire g1511_p_spl_;
  wire g1511_p_spl_0;
  wire n7747_o2_p_spl_;
  wire n7747_o2_p_spl_0;
  wire n7747_o2_p_spl_00;
  wire n7747_o2_p_spl_01;
  wire n7747_o2_p_spl_1;
  wire n7747_o2_n_spl_;
  wire n7747_o2_n_spl_0;
  wire n7747_o2_n_spl_00;
  wire n7747_o2_n_spl_1;
  wire g1515_n_spl_;
  wire g1514_n_spl_;
  wire g1515_p_spl_;
  wire g1514_p_spl_;
  wire g1516_n_spl_;
  wire g1516_n_spl_0;
  wire g1516_p_spl_;
  wire g1516_p_spl_0;
  wire g1520_n_spl_;
  wire g1519_n_spl_;
  wire g1520_p_spl_;
  wire g1519_p_spl_;
  wire g1521_n_spl_;
  wire g1521_n_spl_0;
  wire g1521_p_spl_;
  wire g1521_p_spl_0;
  wire g1525_n_spl_;
  wire g1524_n_spl_;
  wire g1525_p_spl_;
  wire g1524_p_spl_;
  wire g1526_n_spl_;
  wire g1526_n_spl_0;
  wire g1526_p_spl_;
  wire g1526_p_spl_0;
  wire g1530_n_spl_;
  wire g1529_n_spl_;
  wire g1530_p_spl_;
  wire g1529_p_spl_;
  wire g1531_n_spl_;
  wire g1531_n_spl_0;
  wire g1531_p_spl_;
  wire g1531_p_spl_0;
  wire g1535_n_spl_;
  wire g1534_n_spl_;
  wire g1535_p_spl_;
  wire g1534_p_spl_;
  wire g1536_n_spl_;
  wire g1536_n_spl_0;
  wire g1536_p_spl_;
  wire g1536_p_spl_0;
  wire g1075_p_spl_;
  wire g1540_n_spl_;
  wire g1539_n_spl_;
  wire g1540_p_spl_;
  wire g1539_p_spl_;
  wire g1541_n_spl_;
  wire g1541_n_spl_0;
  wire g1541_p_spl_;
  wire g1541_p_spl_0;
  wire g1231_p_spl_;
  wire g1552_n_spl_;
  wire g1551_n_spl_;
  wire g1552_p_spl_;
  wire g1551_p_spl_;
  wire g1553_n_spl_;
  wire g1553_n_spl_0;
  wire g1553_p_spl_;
  wire g1557_n_spl_;
  wire g1556_n_spl_;
  wire g1557_p_spl_;
  wire g1556_p_spl_;
  wire g1558_n_spl_;
  wire g1558_n_spl_0;
  wire g1558_p_spl_;
  wire g1567_n_spl_;
  wire g1566_n_spl_;
  wire g1567_p_spl_;
  wire g1566_p_spl_;
  wire g1568_n_spl_;
  wire g1568_n_spl_0;
  wire g1568_p_spl_;
  wire g1572_n_spl_;
  wire g1571_n_spl_;
  wire g1572_p_spl_;
  wire g1571_p_spl_;
  wire g1573_n_spl_;
  wire g1573_n_spl_0;
  wire g1573_p_spl_;
  wire g1582_n_spl_;
  wire g1581_n_spl_;
  wire g1582_p_spl_;
  wire g1581_p_spl_;
  wire g1583_n_spl_;
  wire g1583_n_spl_0;
  wire g1583_p_spl_;
  wire g1587_n_spl_;
  wire g1586_n_spl_;
  wire g1587_p_spl_;
  wire g1586_p_spl_;
  wire g1588_n_spl_;
  wire g1588_n_spl_0;
  wire g1588_p_spl_;
  wire g1101_n_spl_;
  wire g1101_n_spl_0;
  wire g1126_n_spl_;
  wire g1126_n_spl_0;
  wire g1151_n_spl_;
  wire g1151_n_spl_0;
  wire g1206_n_spl_;
  wire g1206_n_spl_0;
  wire g1544_n_spl_;
  wire g1507_p_spl_;
  wire g1608_n_spl_;
  wire g1607_n_spl_;
  wire g1608_p_spl_;
  wire g1607_p_spl_;
  wire g1609_n_spl_;
  wire g1609_n_spl_0;
  wire g1609_p_spl_;
  wire g1609_p_spl_0;
  wire g1613_n_spl_;
  wire g1612_n_spl_;
  wire g1613_p_spl_;
  wire g1612_p_spl_;
  wire g1614_n_spl_;
  wire g1614_n_spl_0;
  wire g1614_p_spl_;
  wire g1614_p_spl_0;
  wire g1623_n_spl_;
  wire g1622_n_spl_;
  wire g1623_p_spl_;
  wire g1622_p_spl_;
  wire g1624_n_spl_;
  wire g1624_n_spl_0;
  wire g1624_p_spl_;
  wire g1624_p_spl_0;
  wire g1628_n_spl_;
  wire g1627_n_spl_;
  wire g1628_p_spl_;
  wire g1627_p_spl_;
  wire g1629_n_spl_;
  wire g1629_n_spl_0;
  wire g1629_p_spl_;
  wire g1629_p_spl_0;
  wire g1633_n_spl_;
  wire g1632_n_spl_;
  wire g1633_p_spl_;
  wire g1632_p_spl_;
  wire g1634_n_spl_;
  wire g1634_n_spl_0;
  wire g1634_p_spl_;
  wire g1634_p_spl_0;
  wire g1638_n_spl_;
  wire g1637_n_spl_;
  wire g1638_p_spl_;
  wire g1637_p_spl_;
  wire g1639_n_spl_;
  wire g1639_n_spl_0;
  wire g1639_p_spl_;
  wire g1639_p_spl_0;
  wire g1648_n_spl_;
  wire g1647_n_spl_;
  wire g1648_p_spl_;
  wire g1647_p_spl_;
  wire g1649_n_spl_;
  wire g1649_n_spl_0;
  wire g1649_p_spl_;
  wire g1649_p_spl_0;
  wire g1653_n_spl_;
  wire g1652_n_spl_;
  wire g1653_p_spl_;
  wire g1652_p_spl_;
  wire g1654_n_spl_;
  wire g1654_n_spl_0;
  wire g1654_p_spl_;
  wire g1654_p_spl_0;
  wire g1658_n_spl_;
  wire g1657_n_spl_;
  wire g1658_p_spl_;
  wire g1657_p_spl_;
  wire g1659_n_spl_;
  wire g1659_n_spl_0;
  wire g1659_p_spl_;
  wire g1659_p_spl_0;
  wire g1663_n_spl_;
  wire g1662_n_spl_;
  wire g1663_p_spl_;
  wire g1662_p_spl_;
  wire g1664_n_spl_;
  wire g1664_n_spl_0;
  wire g1664_p_spl_;
  wire g1664_p_spl_0;
  wire g1679_n_spl_;
  wire g1678_n_spl_;
  wire g1679_p_spl_;
  wire g1678_p_spl_;
  wire g1680_n_spl_;
  wire g1680_n_spl_0;
  wire g1680_p_spl_;
  wire g1680_p_spl_0;
  wire g1684_n_spl_;
  wire g1683_n_spl_;
  wire g1684_p_spl_;
  wire g1683_p_spl_;
  wire g1685_n_spl_;
  wire g1685_n_spl_0;
  wire g1685_p_spl_;
  wire g1685_p_spl_0;
  wire g1686_n_spl_;
  wire g1675_n_spl_;
  wire g1686_p_spl_;
  wire g1675_p_spl_;
  wire g1687_n_spl_;
  wire g1687_n_spl_0;
  wire g1687_p_spl_;
  wire g1687_p_spl_0;
  wire g1691_n_spl_;
  wire g1690_n_spl_;
  wire g1691_p_spl_;
  wire g1690_p_spl_;
  wire g1692_n_spl_;
  wire g1692_n_spl_0;
  wire g1692_p_spl_;
  wire g1692_p_spl_0;
  wire g1693_n_spl_;
  wire g1672_n_spl_;
  wire g1693_p_spl_;
  wire g1672_p_spl_;
  wire g1694_n_spl_;
  wire g1694_n_spl_0;
  wire g1694_p_spl_;
  wire g1694_p_spl_0;
  wire g1698_n_spl_;
  wire g1697_n_spl_;
  wire g1698_p_spl_;
  wire g1697_p_spl_;
  wire g1699_n_spl_;
  wire g1699_n_spl_0;
  wire g1699_p_spl_;
  wire g1699_p_spl_0;
  wire g1709_n_spl_;
  wire g1708_n_spl_;
  wire g1709_p_spl_;
  wire g1708_p_spl_;
  wire g1710_n_spl_;
  wire g1710_n_spl_0;
  wire g1710_p_spl_;
  wire g1710_p_spl_0;
  wire g1714_n_spl_;
  wire g1713_n_spl_;
  wire g1714_p_spl_;
  wire g1713_p_spl_;
  wire g1715_n_spl_;
  wire g1715_n_spl_0;
  wire g1715_p_spl_;
  wire g1715_p_spl_0;
  wire g1716_n_spl_;
  wire g1705_n_spl_;
  wire g1716_p_spl_;
  wire g1705_p_spl_;
  wire g1717_n_spl_;
  wire g1717_n_spl_0;
  wire g1717_p_spl_;
  wire g1717_p_spl_0;
  wire g1721_n_spl_;
  wire g1720_n_spl_;
  wire g1721_p_spl_;
  wire g1720_p_spl_;
  wire g1722_n_spl_;
  wire g1722_n_spl_0;
  wire g1722_p_spl_;
  wire g1722_p_spl_0;
  wire n2668_lo_buf_o2_p_spl_;
  wire n2668_lo_buf_o2_p_spl_0;
  wire n2668_lo_buf_o2_p_spl_00;
  wire n2668_lo_buf_o2_p_spl_1;
  wire n2668_lo_buf_o2_n_spl_;
  wire n2668_lo_buf_o2_n_spl_0;
  wire g1726_n_spl_;
  wire g1725_n_spl_;
  wire g1726_p_spl_;
  wire g1725_p_spl_;
  wire g1727_n_spl_;
  wire g1727_n_spl_0;
  wire g1727_p_spl_;
  wire g1727_p_spl_0;
  wire n2656_lo_buf_o2_p_spl_;
  wire n2656_lo_buf_o2_p_spl_0;
  wire n2656_lo_buf_o2_p_spl_1;
  wire n2656_lo_buf_o2_n_spl_;
  wire n2656_lo_buf_o2_n_spl_0;
  wire g1731_n_spl_;
  wire g1730_n_spl_;
  wire g1731_p_spl_;
  wire g1730_p_spl_;
  wire g1732_n_spl_;
  wire g1732_n_spl_0;
  wire g1732_p_spl_;
  wire g1732_p_spl_0;
  wire G2139_o2_n_spl_;
  wire G2136_o2_n_spl_;
  wire G2139_o2_p_spl_;
  wire G2136_o2_p_spl_;
  wire g1736_n_spl_;
  wire g1736_n_spl_0;
  wire g1736_p_spl_;
  wire g1736_p_spl_0;
  wire n2644_lo_buf_o2_p_spl_;
  wire n2644_lo_buf_o2_p_spl_0;
  wire n2644_lo_buf_o2_p_spl_1;
  wire n2644_lo_buf_o2_n_spl_;
  wire n2644_lo_buf_o2_n_spl_0;
  wire g1740_n_spl_;
  wire g1739_n_spl_;
  wire g1740_p_spl_;
  wire g1739_p_spl_;
  wire g1741_n_spl_;
  wire g1741_n_spl_0;
  wire g1741_p_spl_;
  wire g1741_p_spl_0;
  wire g1742_n_spl_;
  wire g1735_n_spl_;
  wire g1742_p_spl_;
  wire g1735_p_spl_;
  wire g1743_n_spl_;
  wire g1743_n_spl_0;
  wire g1743_p_spl_;
  wire g1743_p_spl_0;
  wire g1747_n_spl_;
  wire g1746_n_spl_;
  wire g1747_p_spl_;
  wire g1746_p_spl_;
  wire g1748_n_spl_;
  wire g1748_n_spl_0;
  wire g1748_p_spl_;
  wire g1748_p_spl_0;
  wire n2632_lo_buf_o2_p_spl_;
  wire n2632_lo_buf_o2_p_spl_0;
  wire n2632_lo_buf_o2_p_spl_1;
  wire n2632_lo_buf_o2_n_spl_;
  wire n2632_lo_buf_o2_n_spl_0;
  wire n2632_lo_buf_o2_n_spl_1;
  wire g1756_n_spl_;
  wire g1755_n_spl_;
  wire g1756_p_spl_;
  wire g1755_p_spl_;
  wire g1757_n_spl_;
  wire g1757_n_spl_0;
  wire g1757_p_spl_;
  wire g1757_p_spl_0;
  wire g1758_n_spl_;
  wire g1754_n_spl_;
  wire g1758_p_spl_;
  wire g1754_p_spl_;
  wire g1759_n_spl_;
  wire g1759_n_spl_0;
  wire g1759_p_spl_;
  wire g1759_p_spl_0;
  wire g1763_n_spl_;
  wire g1762_n_spl_;
  wire g1763_p_spl_;
  wire g1762_p_spl_;
  wire g1764_n_spl_;
  wire g1764_n_spl_0;
  wire g1764_p_spl_;
  wire g1764_p_spl_0;
  wire g1765_n_spl_;
  wire g1751_n_spl_;
  wire g1765_p_spl_;
  wire g1751_p_spl_;
  wire g1766_n_spl_;
  wire g1766_n_spl_0;
  wire g1766_p_spl_;
  wire g1766_p_spl_0;
  wire n2746_lo_p_spl_;
  wire n2746_lo_p_spl_0;
  wire n2746_lo_p_spl_00;
  wire n2746_lo_p_spl_000;
  wire n2746_lo_p_spl_001;
  wire n2746_lo_p_spl_01;
  wire n2746_lo_p_spl_010;
  wire n2746_lo_p_spl_011;
  wire n2746_lo_p_spl_1;
  wire n2746_lo_p_spl_10;
  wire n2746_lo_p_spl_100;
  wire n2746_lo_p_spl_101;
  wire n2746_lo_p_spl_11;
  wire n2746_lo_p_spl_110;
  wire n2746_lo_n_spl_;
  wire n2746_lo_n_spl_0;
  wire n2746_lo_n_spl_00;
  wire n2746_lo_n_spl_000;
  wire n2746_lo_n_spl_001;
  wire n2746_lo_n_spl_01;
  wire n2746_lo_n_spl_010;
  wire n2746_lo_n_spl_011;
  wire n2746_lo_n_spl_1;
  wire n2746_lo_n_spl_10;
  wire n2746_lo_n_spl_100;
  wire n2746_lo_n_spl_101;
  wire n2746_lo_n_spl_11;
  wire n2746_lo_n_spl_110;
  wire g1770_n_spl_;
  wire g1769_n_spl_;
  wire g1770_p_spl_;
  wire g1769_p_spl_;
  wire g1771_n_spl_;
  wire g1771_n_spl_0;
  wire g1771_p_spl_;
  wire g1771_p_spl_0;
  wire G2309_o2_p_spl_;
  wire G2309_o2_p_spl_0;
  wire G2309_o2_n_spl_;
  wire G2309_o2_n_spl_0;
  wire n2620_lo_buf_o2_p_spl_;
  wire n2620_lo_buf_o2_p_spl_0;
  wire n2620_lo_buf_o2_p_spl_00;
  wire n2620_lo_buf_o2_p_spl_1;
  wire n2620_lo_buf_o2_n_spl_;
  wire n2620_lo_buf_o2_n_spl_0;
  wire n2620_lo_buf_o2_n_spl_1;
  wire g1784_n_spl_;
  wire g1783_n_spl_;
  wire g1784_p_spl_;
  wire g1783_p_spl_;
  wire g1785_n_spl_;
  wire g1785_n_spl_0;
  wire g1785_p_spl_;
  wire g1785_p_spl_0;
  wire g1786_n_spl_;
  wire g1780_n_spl_;
  wire g1786_p_spl_;
  wire g1780_p_spl_;
  wire g1787_n_spl_;
  wire g1787_n_spl_0;
  wire g1787_p_spl_;
  wire g1787_p_spl_0;
  wire g1791_n_spl_;
  wire g1790_n_spl_;
  wire g1791_p_spl_;
  wire g1790_p_spl_;
  wire g1792_n_spl_;
  wire g1792_n_spl_0;
  wire g1792_p_spl_;
  wire g1792_p_spl_0;
  wire g1793_n_spl_;
  wire g1777_n_spl_;
  wire g1793_p_spl_;
  wire g1777_p_spl_;
  wire g1794_n_spl_;
  wire g1794_n_spl_0;
  wire g1794_p_spl_;
  wire g1794_p_spl_0;
  wire g1798_n_spl_;
  wire g1797_n_spl_;
  wire g1798_p_spl_;
  wire g1797_p_spl_;
  wire g1799_n_spl_;
  wire g1799_n_spl_0;
  wire g1799_p_spl_;
  wire g1799_p_spl_0;
  wire g1800_n_spl_;
  wire g1774_n_spl_;
  wire g1800_p_spl_;
  wire g1774_p_spl_;
  wire g1293_n_spl_;
  wire g1293_n_spl_0;
  wire g1293_p_spl_;
  wire g1367_n_spl_;
  wire g1367_n_spl_0;
  wire g1367_p_spl_;
  wire g1477_n_spl_;
  wire g1477_n_spl_0;
  wire g1477_p_spl_;
  wire n2821_lo_p_spl_;
  wire n2821_lo_p_spl_0;
  wire n2821_lo_p_spl_1;
  wire n2821_lo_n_spl_;
  wire n2821_lo_n_spl_0;
  wire n2821_lo_n_spl_1;
  wire g1823_n_spl_;
  wire g1822_n_spl_;
  wire g1823_p_spl_;
  wire g1822_p_spl_;
  wire g1824_n_spl_;
  wire g1824_n_spl_0;
  wire g1824_p_spl_;
  wire g1824_p_spl_0;
  wire g1828_n_spl_;
  wire g1827_n_spl_;
  wire g1828_p_spl_;
  wire g1827_p_spl_;
  wire g1829_n_spl_;
  wire g1829_n_spl_0;
  wire g1829_p_spl_;
  wire g1829_p_spl_0;
  wire G19_p_spl_;
  wire G19_p_spl_0;
  wire G19_p_spl_00;
  wire G19_p_spl_000;
  wire G19_p_spl_001;
  wire G19_p_spl_01;
  wire G19_p_spl_010;
  wire G19_p_spl_011;
  wire G19_p_spl_1;
  wire G19_p_spl_10;
  wire G19_p_spl_100;
  wire G19_p_spl_11;
  wire G16_p_spl_;
  wire G16_p_spl_0;
  wire G16_p_spl_1;
  wire G19_n_spl_;
  wire G19_n_spl_0;
  wire G19_n_spl_00;
  wire G19_n_spl_000;
  wire G19_n_spl_001;
  wire G19_n_spl_01;
  wire G19_n_spl_010;
  wire G19_n_spl_011;
  wire G19_n_spl_1;
  wire G19_n_spl_10;
  wire G19_n_spl_11;
  wire G16_n_spl_;
  wire G16_n_spl_0;
  wire G18_p_spl_;
  wire G18_p_spl_0;
  wire G18_p_spl_00;
  wire G18_p_spl_000;
  wire G18_p_spl_001;
  wire G18_p_spl_01;
  wire G18_p_spl_010;
  wire G18_p_spl_011;
  wire G18_p_spl_1;
  wire G18_p_spl_10;
  wire G18_p_spl_100;
  wire G18_p_spl_101;
  wire G18_p_spl_11;
  wire G18_p_spl_110;
  wire G18_n_spl_;
  wire G18_n_spl_0;
  wire G18_n_spl_00;
  wire G18_n_spl_000;
  wire G18_n_spl_001;
  wire G18_n_spl_01;
  wire G18_n_spl_010;
  wire G18_n_spl_011;
  wire G18_n_spl_1;
  wire G18_n_spl_10;
  wire G18_n_spl_100;
  wire G18_n_spl_101;
  wire G18_n_spl_11;
  wire G18_n_spl_110;
  wire G18_n_spl_111;
  wire G17_p_spl_;
  wire G17_p_spl_0;
  wire G17_p_spl_00;
  wire G17_p_spl_000;
  wire G17_p_spl_001;
  wire G17_p_spl_01;
  wire G17_p_spl_010;
  wire G17_p_spl_011;
  wire G17_p_spl_1;
  wire G17_p_spl_10;
  wire G17_p_spl_100;
  wire G17_p_spl_101;
  wire G17_p_spl_11;
  wire G17_p_spl_110;
  wire G17_p_spl_111;
  wire G17_n_spl_;
  wire G17_n_spl_0;
  wire G17_n_spl_00;
  wire G17_n_spl_000;
  wire G17_n_spl_001;
  wire G17_n_spl_01;
  wire G17_n_spl_010;
  wire G17_n_spl_011;
  wire G17_n_spl_1;
  wire G17_n_spl_10;
  wire G17_n_spl_100;
  wire G17_n_spl_101;
  wire G17_n_spl_11;
  wire G17_n_spl_110;
  wire G15_p_spl_;
  wire G15_p_spl_0;
  wire G15_p_spl_00;
  wire G15_p_spl_1;
  wire G15_n_spl_;
  wire G15_n_spl_0;
  wire G15_n_spl_1;
  wire g1836_n_spl_;
  wire g1835_p_spl_;
  wire g1836_p_spl_;
  wire g1835_n_spl_;
  wire g1837_n_spl_;
  wire g1837_p_spl_;
  wire g1838_n_spl_;
  wire g1838_n_spl_0;
  wire g1834_n_spl_;
  wire g1838_p_spl_;
  wire g1838_p_spl_0;
  wire g1834_p_spl_;
  wire g1839_n_spl_;
  wire g1839_n_spl_0;
  wire g1839_p_spl_;
  wire g1839_p_spl_0;
  wire g1843_n_spl_;
  wire g1842_n_spl_;
  wire g1843_p_spl_;
  wire g1842_p_spl_;
  wire g1844_n_spl_;
  wire g1844_n_spl_0;
  wire g1844_p_spl_;
  wire g1844_p_spl_0;
  wire g1845_n_spl_;
  wire g1833_n_spl_;
  wire g1845_p_spl_;
  wire g1833_p_spl_;
  wire g1848_n_spl_;
  wire g1847_n_spl_;
  wire g1848_p_spl_;
  wire g1847_p_spl_;
  wire g1849_n_spl_;
  wire g1849_n_spl_0;
  wire g1849_p_spl_;
  wire g1849_p_spl_0;
  wire g1853_n_spl_;
  wire g1852_n_spl_;
  wire g1853_p_spl_;
  wire g1852_p_spl_;
  wire g1854_n_spl_;
  wire g1854_n_spl_0;
  wire g1854_p_spl_;
  wire g1854_p_spl_0;
  wire g1858_n_spl_;
  wire g1857_n_spl_;
  wire g1858_p_spl_;
  wire g1857_p_spl_;
  wire g1859_n_spl_;
  wire g1859_n_spl_0;
  wire g1859_p_spl_;
  wire g1859_p_spl_0;
  wire g1863_n_spl_;
  wire g1862_n_spl_;
  wire g1863_p_spl_;
  wire g1862_p_spl_;
  wire g1864_n_spl_;
  wire g1864_n_spl_0;
  wire g1864_p_spl_;
  wire g1864_p_spl_0;
  wire n2572_lo_buf_o2_p_spl_;
  wire n2572_lo_buf_o2_p_spl_0;
  wire n2572_lo_buf_o2_p_spl_00;
  wire n2572_lo_buf_o2_p_spl_01;
  wire n2572_lo_buf_o2_p_spl_1;
  wire n2572_lo_buf_o2_p_spl_10;
  wire n2572_lo_buf_o2_n_spl_;
  wire n2572_lo_buf_o2_n_spl_0;
  wire n2572_lo_buf_o2_n_spl_00;
  wire n2572_lo_buf_o2_n_spl_1;
  wire g1871_n_spl_;
  wire g1870_n_spl_;
  wire g1871_p_spl_;
  wire g1870_p_spl_;
  wire g1872_n_spl_;
  wire g1872_n_spl_0;
  wire g1872_p_spl_;
  wire g1872_p_spl_0;
  wire G1968_o2_p_spl_;
  wire G1968_o2_p_spl_0;
  wire G1968_o2_n_spl_;
  wire G1968_o2_n_spl_0;
  wire n2560_lo_buf_o2_p_spl_;
  wire n2560_lo_buf_o2_p_spl_0;
  wire n2560_lo_buf_o2_p_spl_00;
  wire n2560_lo_buf_o2_p_spl_01;
  wire n2560_lo_buf_o2_p_spl_1;
  wire n2560_lo_buf_o2_n_spl_;
  wire n2560_lo_buf_o2_n_spl_0;
  wire n2560_lo_buf_o2_n_spl_00;
  wire n2560_lo_buf_o2_n_spl_1;
  wire g1879_n_spl_;
  wire g1878_n_spl_;
  wire g1879_p_spl_;
  wire g1878_p_spl_;
  wire g1880_n_spl_;
  wire g1880_n_spl_0;
  wire g1880_p_spl_;
  wire g1880_p_spl_0;
  wire g1881_n_spl_;
  wire g1875_n_spl_;
  wire g1881_p_spl_;
  wire g1875_p_spl_;
  wire g1882_n_spl_;
  wire g1882_n_spl_0;
  wire g1882_p_spl_;
  wire g1882_p_spl_0;
  wire g1886_n_spl_;
  wire g1885_n_spl_;
  wire g1886_p_spl_;
  wire g1885_p_spl_;
  wire g1887_n_spl_;
  wire g1887_n_spl_0;
  wire g1887_p_spl_;
  wire g1887_p_spl_0;
  wire G1914_o2_n_spl_;
  wire G1849_o2_n_spl_;
  wire G1914_o2_p_spl_;
  wire G1849_o2_p_spl_;
  wire g1894_n_spl_;
  wire g1894_n_spl_0;
  wire g1894_p_spl_;
  wire g1894_p_spl_0;
  wire n2548_lo_buf_o2_p_spl_;
  wire n2548_lo_buf_o2_p_spl_0;
  wire n2548_lo_buf_o2_p_spl_00;
  wire n2548_lo_buf_o2_p_spl_01;
  wire n2548_lo_buf_o2_p_spl_1;
  wire n2548_lo_buf_o2_n_spl_;
  wire n2548_lo_buf_o2_n_spl_0;
  wire n2548_lo_buf_o2_n_spl_00;
  wire n2548_lo_buf_o2_n_spl_1;
  wire g1898_n_spl_;
  wire g1897_n_spl_;
  wire g1898_p_spl_;
  wire g1897_p_spl_;
  wire g1899_n_spl_;
  wire g1899_n_spl_0;
  wire g1899_p_spl_;
  wire g1899_p_spl_0;
  wire g1900_n_spl_;
  wire g1893_n_spl_;
  wire g1900_p_spl_;
  wire g1893_p_spl_;
  wire g1901_n_spl_;
  wire g1901_n_spl_0;
  wire g1901_p_spl_;
  wire g1901_p_spl_0;
  wire g1905_n_spl_;
  wire g1904_n_spl_;
  wire g1905_p_spl_;
  wire g1904_p_spl_;
  wire g1906_n_spl_;
  wire g1906_n_spl_0;
  wire g1906_p_spl_;
  wire g1906_p_spl_0;
  wire g1907_n_spl_;
  wire g1890_n_spl_;
  wire g1907_p_spl_;
  wire g1890_p_spl_;
  wire g1908_n_spl_;
  wire g1908_n_spl_0;
  wire g1908_p_spl_;
  wire g1908_p_spl_0;
  wire g1912_n_spl_;
  wire g1911_n_spl_;
  wire g1912_p_spl_;
  wire g1911_p_spl_;
  wire g1913_n_spl_;
  wire g1913_n_spl_0;
  wire g1913_p_spl_;
  wire g1913_p_spl_0;
  wire G1777_o2_n_spl_;
  wire G1777_o2_n_spl_0;
  wire G1777_o2_p_spl_;
  wire G1777_o2_p_spl_0;
  wire g1924_n_spl_;
  wire g1923_n_spl_;
  wire g1924_p_spl_;
  wire g1923_p_spl_;
  wire g1925_n_spl_;
  wire g1925_n_spl_0;
  wire g1925_p_spl_;
  wire g1925_p_spl_0;
  wire n2536_lo_buf_o2_p_spl_;
  wire n2536_lo_buf_o2_p_spl_0;
  wire n2536_lo_buf_o2_p_spl_00;
  wire n2536_lo_buf_o2_p_spl_01;
  wire n2536_lo_buf_o2_p_spl_1;
  wire n2536_lo_buf_o2_n_spl_;
  wire n2536_lo_buf_o2_n_spl_0;
  wire n2536_lo_buf_o2_n_spl_00;
  wire n2536_lo_buf_o2_n_spl_1;
  wire g1929_n_spl_;
  wire g1928_n_spl_;
  wire g1929_p_spl_;
  wire g1928_p_spl_;
  wire g1930_n_spl_;
  wire g1930_n_spl_0;
  wire g1930_p_spl_;
  wire g1930_p_spl_0;
  wire g1931_n_spl_;
  wire g1922_n_spl_;
  wire g1931_p_spl_;
  wire g1922_p_spl_;
  wire g1932_n_spl_;
  wire g1932_n_spl_0;
  wire g1932_p_spl_;
  wire g1932_p_spl_0;
  wire g1936_n_spl_;
  wire g1935_n_spl_;
  wire g1936_p_spl_;
  wire g1935_p_spl_;
  wire g1937_n_spl_;
  wire g1937_n_spl_0;
  wire g1937_p_spl_;
  wire g1937_p_spl_0;
  wire g1938_n_spl_;
  wire g1919_n_spl_;
  wire g1938_p_spl_;
  wire g1919_p_spl_;
  wire g1939_n_spl_;
  wire g1939_n_spl_0;
  wire g1939_p_spl_;
  wire g1939_p_spl_0;
  wire g1943_n_spl_;
  wire g1942_n_spl_;
  wire g1943_p_spl_;
  wire g1942_p_spl_;
  wire g1944_n_spl_;
  wire g1944_n_spl_0;
  wire g1944_p_spl_;
  wire g1944_p_spl_0;
  wire g1945_n_spl_;
  wire g1916_n_spl_;
  wire g1945_p_spl_;
  wire g1916_p_spl_;
  wire g1946_n_spl_;
  wire g1946_n_spl_0;
  wire g1946_p_spl_;
  wire g1946_p_spl_0;
  wire g1950_n_spl_;
  wire g1949_n_spl_;
  wire g1950_p_spl_;
  wire g1949_p_spl_;
  wire g1951_n_spl_;
  wire g1951_n_spl_0;
  wire g1951_p_spl_;
  wire g1951_p_spl_0;
  wire g1967_n_spl_;
  wire g1966_n_spl_;
  wire g1967_p_spl_;
  wire g1966_p_spl_;
  wire g1968_n_spl_;
  wire g1968_n_spl_0;
  wire g1968_p_spl_;
  wire g1968_p_spl_0;
  wire n2524_lo_buf_o2_p_spl_;
  wire n2524_lo_buf_o2_p_spl_0;
  wire n2524_lo_buf_o2_p_spl_00;
  wire n2524_lo_buf_o2_p_spl_1;
  wire n2524_lo_buf_o2_n_spl_;
  wire n2524_lo_buf_o2_n_spl_0;
  wire n2524_lo_buf_o2_n_spl_00;
  wire n2524_lo_buf_o2_n_spl_1;
  wire g1972_n_spl_;
  wire g1971_n_spl_;
  wire g1972_p_spl_;
  wire g1971_p_spl_;
  wire g1973_n_spl_;
  wire g1973_n_spl_0;
  wire g1973_p_spl_;
  wire g1973_p_spl_0;
  wire g1974_n_spl_;
  wire g1963_n_spl_;
  wire g1974_p_spl_;
  wire g1963_p_spl_;
  wire g1975_n_spl_;
  wire g1975_n_spl_0;
  wire g1975_p_spl_;
  wire g1975_p_spl_0;
  wire g1979_n_spl_;
  wire g1978_n_spl_;
  wire g1979_p_spl_;
  wire g1978_p_spl_;
  wire g1980_n_spl_;
  wire g1980_n_spl_0;
  wire g1980_p_spl_;
  wire g1980_p_spl_0;
  wire g1981_n_spl_;
  wire g1960_n_spl_;
  wire g1981_p_spl_;
  wire g1960_p_spl_;
  wire g1982_n_spl_;
  wire g1982_n_spl_0;
  wire g1982_p_spl_;
  wire g1982_p_spl_0;
  wire g1986_n_spl_;
  wire g1985_n_spl_;
  wire g1986_p_spl_;
  wire g1985_p_spl_;
  wire g1987_n_spl_;
  wire g1987_n_spl_0;
  wire g1987_p_spl_;
  wire g1987_p_spl_0;
  wire g1988_n_spl_;
  wire g1957_n_spl_;
  wire g1988_p_spl_;
  wire g1957_p_spl_;
  wire g1989_n_spl_;
  wire g1989_n_spl_0;
  wire g1989_p_spl_;
  wire g1989_p_spl_0;
  wire g1993_n_spl_;
  wire g1992_n_spl_;
  wire g1993_p_spl_;
  wire g1992_p_spl_;
  wire g1994_n_spl_;
  wire g1994_n_spl_0;
  wire g1994_p_spl_;
  wire g1994_p_spl_0;
  wire G2250_o2_n_spl_;
  wire G2198_o2_n_spl_;
  wire G2250_o2_p_spl_;
  wire G2198_o2_p_spl_;
  wire g2003_n_spl_;
  wire g2003_n_spl_0;
  wire g2003_p_spl_;
  wire g2003_p_spl_0;
  wire n2608_lo_buf_o2_p_spl_;
  wire n2608_lo_buf_o2_p_spl_0;
  wire n2608_lo_buf_o2_p_spl_00;
  wire n2608_lo_buf_o2_p_spl_1;
  wire n2608_lo_buf_o2_n_spl_;
  wire n2608_lo_buf_o2_n_spl_0;
  wire n2608_lo_buf_o2_n_spl_1;
  wire g2007_n_spl_;
  wire g2006_n_spl_;
  wire g2007_p_spl_;
  wire g2006_p_spl_;
  wire g2008_n_spl_;
  wire g2008_n_spl_0;
  wire g2008_p_spl_;
  wire g2008_p_spl_0;
  wire g2009_n_spl_;
  wire g2002_n_spl_;
  wire g2009_p_spl_;
  wire g2002_p_spl_;
  wire g2010_n_spl_;
  wire g2010_n_spl_0;
  wire g2010_p_spl_;
  wire g2010_p_spl_0;
  wire g2014_n_spl_;
  wire g2013_n_spl_;
  wire g2014_p_spl_;
  wire g2013_p_spl_;
  wire g2015_n_spl_;
  wire g2015_n_spl_0;
  wire g2015_p_spl_;
  wire g2015_p_spl_0;
  wire g2016_n_spl_;
  wire g1999_n_spl_;
  wire g2016_p_spl_;
  wire g1999_p_spl_;
  wire g2017_n_spl_;
  wire g2017_n_spl_0;
  wire g2017_p_spl_;
  wire g2017_p_spl_0;
  wire g2021_n_spl_;
  wire g2020_n_spl_;
  wire g2021_p_spl_;
  wire g2020_p_spl_;
  wire g2022_n_spl_;
  wire g2022_n_spl_0;
  wire g2022_p_spl_;
  wire g2022_p_spl_0;
  wire G2118_o2_n_spl_;
  wire G2118_o2_n_spl_0;
  wire G2118_o2_p_spl_;
  wire G2118_o2_p_spl_0;
  wire g2033_n_spl_;
  wire g2032_n_spl_;
  wire g2033_p_spl_;
  wire g2032_p_spl_;
  wire g2034_n_spl_;
  wire g2034_n_spl_0;
  wire g2034_p_spl_;
  wire g2034_p_spl_0;
  wire n2596_lo_buf_o2_p_spl_;
  wire n2596_lo_buf_o2_p_spl_0;
  wire n2596_lo_buf_o2_p_spl_00;
  wire n2596_lo_buf_o2_p_spl_1;
  wire n2596_lo_buf_o2_n_spl_;
  wire n2596_lo_buf_o2_n_spl_0;
  wire n2596_lo_buf_o2_n_spl_1;
  wire g2038_n_spl_;
  wire g2037_n_spl_;
  wire g2038_p_spl_;
  wire g2037_p_spl_;
  wire g2039_n_spl_;
  wire g2039_n_spl_0;
  wire g2039_p_spl_;
  wire g2039_p_spl_0;
  wire g2040_n_spl_;
  wire g2031_n_spl_;
  wire g2040_p_spl_;
  wire g2031_p_spl_;
  wire g2041_n_spl_;
  wire g2041_n_spl_0;
  wire g2041_p_spl_;
  wire g2041_p_spl_0;
  wire g2045_n_spl_;
  wire g2044_n_spl_;
  wire g2045_p_spl_;
  wire g2044_p_spl_;
  wire g2046_n_spl_;
  wire g2046_n_spl_0;
  wire g2046_p_spl_;
  wire g2046_p_spl_0;
  wire g2047_n_spl_;
  wire g2028_n_spl_;
  wire g2047_p_spl_;
  wire g2028_p_spl_;
  wire g2048_n_spl_;
  wire g2048_n_spl_0;
  wire g2048_p_spl_;
  wire g2048_p_spl_0;
  wire g2052_n_spl_;
  wire g2051_n_spl_;
  wire g2052_p_spl_;
  wire g2051_p_spl_;
  wire g2053_n_spl_;
  wire g2053_n_spl_0;
  wire g2053_p_spl_;
  wire g2053_p_spl_0;
  wire g2054_n_spl_;
  wire g2025_n_spl_;
  wire g2054_p_spl_;
  wire g2025_p_spl_;
  wire g2055_n_spl_;
  wire g2055_n_spl_0;
  wire g2055_p_spl_;
  wire g2055_p_spl_0;
  wire n2758_lo_p_spl_;
  wire n2758_lo_p_spl_0;
  wire n2758_lo_p_spl_00;
  wire n2758_lo_p_spl_000;
  wire n2758_lo_p_spl_001;
  wire n2758_lo_p_spl_01;
  wire n2758_lo_p_spl_1;
  wire n2758_lo_p_spl_10;
  wire n2758_lo_p_spl_11;
  wire n2758_lo_n_spl_;
  wire n2758_lo_n_spl_0;
  wire n2758_lo_n_spl_00;
  wire n2758_lo_n_spl_000;
  wire n2758_lo_n_spl_001;
  wire n2758_lo_n_spl_01;
  wire n2758_lo_n_spl_1;
  wire n2758_lo_n_spl_10;
  wire n2758_lo_n_spl_11;
  wire g2059_n_spl_;
  wire g2058_n_spl_;
  wire g2059_p_spl_;
  wire g2058_p_spl_;
  wire g2060_n_spl_;
  wire g2060_n_spl_0;
  wire g2060_p_spl_;
  wire g2060_p_spl_0;
  wire G2058_o2_p_spl_;
  wire G935_o2_n_spl_;
  wire G2058_o2_n_spl_;
  wire G935_o2_p_spl_;
  wire g2076_n_spl_;
  wire g2076_n_spl_0;
  wire g2076_p_spl_;
  wire g2076_p_spl_0;
  wire g2077_n_spl_;
  wire g2075_n_spl_;
  wire g2077_p_spl_;
  wire g2075_p_spl_;
  wire g2078_n_spl_;
  wire g2078_n_spl_0;
  wire g2078_p_spl_;
  wire g2078_p_spl_0;
  wire n2584_lo_buf_o2_p_spl_;
  wire n2584_lo_buf_o2_p_spl_0;
  wire n2584_lo_buf_o2_p_spl_00;
  wire n2584_lo_buf_o2_p_spl_1;
  wire n2584_lo_buf_o2_n_spl_;
  wire n2584_lo_buf_o2_n_spl_0;
  wire n2584_lo_buf_o2_n_spl_00;
  wire n2584_lo_buf_o2_n_spl_1;
  wire g2082_n_spl_;
  wire g2081_n_spl_;
  wire g2082_p_spl_;
  wire g2081_p_spl_;
  wire g2083_n_spl_;
  wire g2083_n_spl_0;
  wire g2083_p_spl_;
  wire g2083_p_spl_0;
  wire g2084_n_spl_;
  wire g2072_n_spl_;
  wire g2084_p_spl_;
  wire g2072_p_spl_;
  wire g2085_n_spl_;
  wire g2085_n_spl_0;
  wire g2085_p_spl_;
  wire g2085_p_spl_0;
  wire g2089_n_spl_;
  wire g2088_n_spl_;
  wire g2089_p_spl_;
  wire g2088_p_spl_;
  wire g2090_n_spl_;
  wire g2090_n_spl_0;
  wire g2090_p_spl_;
  wire g2090_p_spl_0;
  wire g2091_n_spl_;
  wire g2069_n_spl_;
  wire g2091_p_spl_;
  wire g2069_p_spl_;
  wire g2092_n_spl_;
  wire g2092_n_spl_0;
  wire g2092_p_spl_;
  wire g2092_p_spl_0;
  wire g2096_n_spl_;
  wire g2095_n_spl_;
  wire g2096_p_spl_;
  wire g2095_p_spl_;
  wire g2097_n_spl_;
  wire g2097_n_spl_0;
  wire g2097_p_spl_;
  wire g2097_p_spl_0;
  wire g2098_n_spl_;
  wire g2066_n_spl_;
  wire g2098_p_spl_;
  wire g2066_p_spl_;
  wire g2099_n_spl_;
  wire g2099_n_spl_0;
  wire g2099_p_spl_;
  wire g2099_p_spl_0;
  wire g2103_n_spl_;
  wire g2102_n_spl_;
  wire g2103_p_spl_;
  wire g2102_p_spl_;
  wire g2104_n_spl_;
  wire g2104_n_spl_0;
  wire g2104_p_spl_;
  wire g2104_p_spl_0;
  wire g2110_n_spl_;
  wire g2109_n_spl_;
  wire g2110_p_spl_;
  wire g2109_p_spl_;
  wire g2111_n_spl_;
  wire g2111_n_spl_0;
  wire g2111_p_spl_;
  wire g2111_p_spl_0;
  wire g2115_n_spl_;
  wire g2114_n_spl_;
  wire g2115_p_spl_;
  wire g2114_p_spl_;
  wire g2116_n_spl_;
  wire g2116_n_spl_0;
  wire g2116_p_spl_;
  wire g2116_p_spl_0;
  wire g2120_n_spl_;
  wire g2119_n_spl_;
  wire g2120_p_spl_;
  wire g2119_p_spl_;
  wire g2121_n_spl_;
  wire g2121_n_spl_0;
  wire g2121_p_spl_;
  wire g2121_p_spl_0;
  wire g2125_n_spl_;
  wire g2124_n_spl_;
  wire g2125_p_spl_;
  wire g2124_p_spl_;
  wire g2126_n_spl_;
  wire g2126_n_spl_0;
  wire g2126_p_spl_;
  wire g2126_p_spl_0;
  wire g1508_p_spl_;
  wire g2130_n_spl_;
  wire g2129_n_spl_;
  wire g2131_n_spl_;
  wire g1563_n_spl_;
  wire g1563_n_spl_0;
  wire g1578_n_spl_;
  wire g1578_n_spl_0;
  wire g1593_n_spl_;
  wire g1593_n_spl_0;
  wire g1602_n_spl_;
  wire g1545_n_spl_;
  wire g1599_n_spl_;
  wire g1546_n_spl_;
  wire g1596_n_spl_;
  wire g1547_n_spl_;
  wire g1605_n_spl_;
  wire g1548_n_spl_;
  wire g1220_n_spl_;
  wire g1220_n_spl_0;
  wire g1225_n_spl_;
  wire g1225_n_spl_0;
  wire g1230_n_spl_;
  wire g1230_n_spl_0;
  wire g2167_n_spl_;
  wire g2166_n_spl_;
  wire g2167_p_spl_;
  wire g2166_p_spl_;
  wire g2168_n_spl_;
  wire g2168_n_spl_0;
  wire g2168_p_spl_;
  wire g2172_n_spl_;
  wire g2171_n_spl_;
  wire g2172_p_spl_;
  wire g2171_p_spl_;
  wire g2173_n_spl_;
  wire g2173_n_spl_0;
  wire g2173_p_spl_;
  wire g2182_n_spl_;
  wire g2181_n_spl_;
  wire g2182_p_spl_;
  wire g2181_p_spl_;
  wire g2183_n_spl_;
  wire g2183_n_spl_0;
  wire g2183_p_spl_;
  wire g2187_n_spl_;
  wire g2186_n_spl_;
  wire g2187_p_spl_;
  wire g2186_p_spl_;
  wire g2188_n_spl_;
  wire g2188_n_spl_0;
  wire g2188_p_spl_;
  wire g1606_p_spl_;
  wire g1619_n_spl_;
  wire g1619_n_spl_0;
  wire g1644_n_spl_;
  wire g1644_n_spl_0;
  wire g1669_n_spl_;
  wire g1669_n_spl_0;
  wire g1724_n_spl_;
  wire g1724_n_spl_0;
  wire g1801_n_spl_;
  wire g1801_n_spl_0;
  wire g1801_p_spl_;
  wire g2134_n_spl_;
  wire g1832_n_spl_;
  wire g2226_n_spl_;
  wire g2225_n_spl_;
  wire g2226_p_spl_;
  wire g2225_p_spl_;
  wire g2227_n_spl_;
  wire g2227_n_spl_0;
  wire g2227_p_spl_;
  wire g2227_p_spl_0;
  wire g2231_n_spl_;
  wire g2230_n_spl_;
  wire g2231_p_spl_;
  wire g2230_p_spl_;
  wire g2232_n_spl_;
  wire g2232_n_spl_0;
  wire g2232_p_spl_;
  wire g2232_p_spl_0;
  wire g2233_n_spl_;
  wire g2222_n_spl_;
  wire g2233_p_spl_;
  wire g2222_p_spl_;
  wire g2234_n_spl_;
  wire g2234_n_spl_0;
  wire g2234_p_spl_;
  wire g2234_p_spl_0;
  wire g2238_n_spl_;
  wire g2237_n_spl_;
  wire g2238_p_spl_;
  wire g2237_p_spl_;
  wire g2239_n_spl_;
  wire g2239_n_spl_0;
  wire g2239_p_spl_;
  wire g2239_p_spl_0;
  wire g2257_n_spl_;
  wire g2256_n_spl_;
  wire g2257_p_spl_;
  wire g2256_p_spl_;
  wire g2258_n_spl_;
  wire g2258_n_spl_0;
  wire g2258_p_spl_;
  wire g2258_p_spl_0;
  wire g2262_n_spl_;
  wire g2261_n_spl_;
  wire g2262_p_spl_;
  wire g2261_p_spl_;
  wire g2263_n_spl_;
  wire g2263_n_spl_0;
  wire g2263_p_spl_;
  wire g2263_p_spl_0;
  wire g2264_n_spl_;
  wire g2253_n_spl_;
  wire g2264_p_spl_;
  wire g2253_p_spl_;
  wire g2265_n_spl_;
  wire g2265_n_spl_0;
  wire g2265_p_spl_;
  wire g2265_p_spl_0;
  wire g2269_n_spl_;
  wire g2268_n_spl_;
  wire g2269_p_spl_;
  wire g2268_p_spl_;
  wire g2270_n_spl_;
  wire g2270_n_spl_0;
  wire g2270_p_spl_;
  wire g2270_p_spl_0;
  wire g2271_n_spl_;
  wire g2250_n_spl_;
  wire g2271_p_spl_;
  wire g2250_p_spl_;
  wire g2272_n_spl_;
  wire g2272_n_spl_0;
  wire g2272_p_spl_;
  wire g2272_p_spl_0;
  wire g2276_n_spl_;
  wire g2275_n_spl_;
  wire g2276_p_spl_;
  wire g2275_p_spl_;
  wire g2277_n_spl_;
  wire g2277_n_spl_0;
  wire g2277_p_spl_;
  wire g2277_p_spl_0;
  wire g2278_n_spl_;
  wire g2247_n_spl_;
  wire g2278_p_spl_;
  wire g2247_p_spl_;
  wire g2279_n_spl_;
  wire g2279_n_spl_0;
  wire g2279_p_spl_;
  wire g2279_p_spl_0;
  wire g2283_n_spl_;
  wire g2282_n_spl_;
  wire g2283_p_spl_;
  wire g2282_p_spl_;
  wire g2284_n_spl_;
  wire g2284_n_spl_0;
  wire g2284_p_spl_;
  wire g2284_p_spl_0;
  wire G7_p_spl_;
  wire G7_p_spl_0;
  wire G7_p_spl_1;
  wire G7_n_spl_;
  wire G7_n_spl_0;
  wire G6_p_spl_;
  wire G6_p_spl_0;
  wire G6_p_spl_1;
  wire G6_n_spl_;
  wire G6_n_spl_0;
  wire g2288_n_spl_;
  wire g2287_p_spl_;
  wire g2288_p_spl_;
  wire g2287_n_spl_;
  wire g2289_n_spl_;
  wire g2289_p_spl_;
  wire g2290_n_spl_;
  wire g2290_n_spl_0;
  wire g2290_p_spl_;
  wire g2290_p_spl_0;
  wire G5_p_spl_;
  wire G5_p_spl_0;
  wire G5_n_spl_;
  wire G5_n_spl_0;
  wire g2294_n_spl_;
  wire g2293_p_spl_;
  wire g2294_p_spl_;
  wire g2293_n_spl_;
  wire g2295_n_spl_;
  wire g2295_p_spl_;
  wire g2296_p_spl_;
  wire G13_p_spl_;
  wire G13_p_spl_0;
  wire G13_p_spl_00;
  wire G13_p_spl_1;
  wire G13_n_spl_;
  wire G13_n_spl_0;
  wire G13_n_spl_1;
  wire G12_p_spl_;
  wire G12_p_spl_0;
  wire G12_p_spl_00;
  wire G12_p_spl_1;
  wire G12_n_spl_;
  wire G12_n_spl_0;
  wire G12_n_spl_1;
  wire g2299_n_spl_;
  wire g2298_p_spl_;
  wire g2299_p_spl_;
  wire g2298_n_spl_;
  wire g2300_n_spl_;
  wire g2300_p_spl_;
  wire g2301_n_spl_;
  wire g2301_n_spl_0;
  wire g2301_p_spl_;
  wire g2301_p_spl_0;
  wire G11_p_spl_;
  wire G11_p_spl_0;
  wire G11_p_spl_00;
  wire G11_p_spl_1;
  wire G11_n_spl_;
  wire G11_n_spl_0;
  wire G11_n_spl_1;
  wire g2305_n_spl_;
  wire g2304_p_spl_;
  wire g2305_p_spl_;
  wire g2304_n_spl_;
  wire g2306_n_spl_;
  wire g2306_p_spl_;
  wire g2307_n_spl_;
  wire g2307_n_spl_0;
  wire g2303_n_spl_;
  wire g2307_p_spl_;
  wire g2307_p_spl_0;
  wire g2303_p_spl_;
  wire g2308_n_spl_;
  wire g2308_n_spl_0;
  wire g2308_p_spl_;
  wire g2308_p_spl_0;
  wire g2312_n_spl_;
  wire g2311_n_spl_;
  wire g2312_p_spl_;
  wire g2311_p_spl_;
  wire g2313_n_spl_;
  wire g2313_n_spl_0;
  wire g2313_p_spl_;
  wire g2313_p_spl_0;
  wire G10_p_spl_;
  wire G10_p_spl_0;
  wire G10_p_spl_1;
  wire G10_n_spl_;
  wire G10_n_spl_0;
  wire G10_n_spl_1;
  wire g2320_n_spl_;
  wire g2319_p_spl_;
  wire g2320_p_spl_;
  wire g2319_n_spl_;
  wire g2321_n_spl_;
  wire g2321_p_spl_;
  wire g2322_n_spl_;
  wire g2322_n_spl_0;
  wire g2318_n_spl_;
  wire g2322_p_spl_;
  wire g2322_p_spl_0;
  wire g2318_p_spl_;
  wire g2323_n_spl_;
  wire g2323_n_spl_0;
  wire g2323_p_spl_;
  wire g2323_p_spl_0;
  wire g2327_n_spl_;
  wire g2326_n_spl_;
  wire g2327_p_spl_;
  wire g2326_p_spl_;
  wire g2328_n_spl_;
  wire g2328_n_spl_0;
  wire g2328_p_spl_;
  wire g2328_p_spl_0;
  wire g2341_n_spl_;
  wire g2340_n_spl_;
  wire g2341_p_spl_;
  wire g2340_p_spl_;
  wire g2342_n_spl_;
  wire g2342_n_spl_0;
  wire g2342_p_spl_;
  wire g2347_n_spl_;
  wire g2347_n_spl_0;
  wire g2216_p_spl_;
  wire g2356_n_spl_;
  wire g2355_n_spl_;
  wire g2356_p_spl_;
  wire g2355_p_spl_;
  wire g2357_n_spl_;
  wire g2357_n_spl_0;
  wire g2357_p_spl_;
  wire g2357_p_spl_0;
  wire g2361_n_spl_;
  wire g2360_n_spl_;
  wire g2361_p_spl_;
  wire g2360_p_spl_;
  wire g2362_n_spl_;
  wire g2362_n_spl_0;
  wire g2362_p_spl_;
  wire g2362_p_spl_0;
  wire g2363_n_spl_;
  wire g2352_n_spl_;
  wire g2363_p_spl_;
  wire g2352_p_spl_;
  wire g2364_n_spl_;
  wire g2364_n_spl_0;
  wire g2364_p_spl_;
  wire g2364_p_spl_0;
  wire g2368_n_spl_;
  wire g2367_n_spl_;
  wire g2368_p_spl_;
  wire g2367_p_spl_;
  wire g2369_n_spl_;
  wire g2369_n_spl_0;
  wire g2369_p_spl_;
  wire g2369_p_spl_0;
  wire g2376_n_spl_;
  wire g2375_n_spl_;
  wire g2376_p_spl_;
  wire g2375_p_spl_;
  wire g2377_n_spl_;
  wire g2377_n_spl_0;
  wire g2377_p_spl_;
  wire g2377_p_spl_0;
  wire g2381_n_spl_;
  wire g2380_n_spl_;
  wire g2381_p_spl_;
  wire g2380_p_spl_;
  wire g2382_n_spl_;
  wire g2382_n_spl_0;
  wire g2382_p_spl_;
  wire g2382_p_spl_0;
  wire g2383_n_spl_;
  wire g2372_n_spl_;
  wire g2383_p_spl_;
  wire g2372_p_spl_;
  wire g2384_n_spl_;
  wire g2384_n_spl_0;
  wire g2384_p_spl_;
  wire g2389_n_spl_;
  wire g2389_n_spl_0;
  wire g2163_n_spl_;
  wire g2163_n_spl_0;
  wire g2178_n_spl_;
  wire g2178_n_spl_0;
  wire g2193_n_spl_;
  wire g2193_n_spl_0;
  wire g2198_n_spl_;
  wire g2198_n_spl_0;
  wire g2201_n_spl_;
  wire g2135_n_spl_;
  wire g2204_n_spl_;
  wire g2136_n_spl_;
  wire g2207_n_spl_;
  wire g2137_n_spl_;
  wire g2210_n_spl_;
  wire g2138_n_spl_;
  wire g1846_n_spl_;
  wire g1846_n_spl_0;
  wire g1846_p_spl_;
  wire G20_p_spl_;
  wire G20_p_spl_0;
  wire G20_p_spl_00;
  wire G20_p_spl_01;
  wire G20_p_spl_1;
  wire G20_p_spl_10;
  wire G20_n_spl_;
  wire G20_n_spl_0;
  wire G20_n_spl_00;
  wire G20_n_spl_01;
  wire G20_n_spl_1;
  wire g2411_n_spl_;
  wire g2410_n_spl_;
  wire g2411_p_spl_;
  wire g2410_p_spl_;
  wire g2412_n_spl_;
  wire g2412_n_spl_0;
  wire g2412_p_spl_;
  wire g2416_n_spl_;
  wire g2415_n_spl_;
  wire g2416_p_spl_;
  wire g2415_p_spl_;
  wire g2417_n_spl_;
  wire g2417_n_spl_0;
  wire g2417_p_spl_;
  wire g2426_n_spl_;
  wire g2425_n_spl_;
  wire g2426_p_spl_;
  wire g2425_p_spl_;
  wire g2427_n_spl_;
  wire g2427_n_spl_0;
  wire g2427_p_spl_;
  wire g2431_n_spl_;
  wire g2430_n_spl_;
  wire g2431_p_spl_;
  wire g2430_p_spl_;
  wire g2432_n_spl_;
  wire g2432_n_spl_0;
  wire g2432_p_spl_;
  wire g2444_n_spl_;
  wire g2443_n_spl_;
  wire g2444_p_spl_;
  wire g2443_p_spl_;
  wire g2445_n_spl_;
  wire g2445_n_spl_0;
  wire g2445_p_spl_;
  wire g2445_p_spl_0;
  wire g2449_n_spl_;
  wire g2448_n_spl_;
  wire g2450_n_spl_;
  wire g2450_n_spl_0;
  wire g2459_n_spl_;
  wire g2458_n_spl_;
  wire g2459_p_spl_;
  wire g2458_p_spl_;
  wire g2460_n_spl_;
  wire g2460_n_spl_0;
  wire g2460_p_spl_;
  wire g2460_p_spl_0;
  wire g2464_p_spl_;
  wire g2463_p_spl_;
  wire g2465_p_spl_;
  wire g2465_p_spl_0;
  wire g1806_n_spl_;
  wire g1806_n_spl_0;
  wire g1811_n_spl_;
  wire g1811_n_spl_0;
  wire g1816_n_spl_;
  wire g1816_n_spl_0;
  wire g1831_n_spl_;
  wire g1831_n_spl_0;
  wire g2296_n_spl_;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_1;
  wire G4_n_spl_;
  wire g2483_n_spl_;
  wire g2482_p_spl_;
  wire g2483_p_spl_;
  wire g2482_n_spl_;
  wire g2484_n_spl_;
  wire g2484_p_spl_;
  wire g2485_p_spl_;
  wire G9_p_spl_;
  wire G9_p_spl_0;
  wire G9_p_spl_00;
  wire G9_p_spl_1;
  wire G9_n_spl_;
  wire G9_n_spl_0;
  wire g2493_n_spl_;
  wire g2492_p_spl_;
  wire g2493_p_spl_;
  wire g2492_n_spl_;
  wire g2494_n_spl_;
  wire g2494_p_spl_;
  wire g2495_n_spl_;
  wire g2495_n_spl_0;
  wire g2491_n_spl_;
  wire g2495_p_spl_;
  wire g2495_p_spl_0;
  wire g2491_p_spl_;
  wire g2496_n_spl_;
  wire g2496_n_spl_0;
  wire g2496_p_spl_;
  wire g2496_p_spl_0;
  wire g2500_n_spl_;
  wire g2499_n_spl_;
  wire g2500_p_spl_;
  wire g2499_p_spl_;
  wire g2501_n_spl_;
  wire g2501_n_spl_0;
  wire g2501_p_spl_;
  wire g2501_p_spl_0;
  wire g1869_n_spl_;
  wire g1869_n_spl_0;
  wire g1996_n_spl_;
  wire g1996_n_spl_0;
  wire g2106_n_spl_;
  wire g2106_n_spl_0;
  wire G2_p_spl_;
  wire G2_p_spl_0;
  wire G2_n_spl_;
  wire n2770_lo_p_spl_;
  wire g2530_n_spl_;
  wire g2529_n_spl_;
  wire g2530_p_spl_;
  wire g2529_p_spl_;
  wire g2531_n_spl_;
  wire g2531_n_spl_0;
  wire g2531_p_spl_;
  wire g2536_n_spl_;
  wire g2536_n_spl_0;
  wire G3_p_spl_;
  wire G3_p_spl_0;
  wire G3_n_spl_;
  wire g2540_p_spl_;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire G8_p_spl_1;
  wire G8_n_spl_;
  wire G8_n_spl_0;
  wire g2543_n_spl_;
  wire g2542_p_spl_;
  wire g2543_p_spl_;
  wire g2542_n_spl_;
  wire g2544_n_spl_;
  wire g2544_p_spl_;
  wire g2545_n_spl_;
  wire g2545_n_spl_0;
  wire g2545_p_spl_;
  wire g2545_p_spl_0;
  wire g2549_n_spl_;
  wire g2548_p_spl_;
  wire g2549_p_spl_;
  wire g2548_n_spl_;
  wire g2550_n_spl_;
  wire g2550_p_spl_;
  wire g2551_n_spl_;
  wire g2551_n_spl_0;
  wire g2547_n_spl_;
  wire g2551_p_spl_;
  wire g2551_p_spl_0;
  wire g2547_p_spl_;
  wire g2552_n_spl_;
  wire g2552_n_spl_0;
  wire g2552_p_spl_;
  wire g2557_n_spl_;
  wire g2557_n_spl_0;
  wire G14_p_spl_;
  wire G14_p_spl_0;
  wire G14_p_spl_00;
  wire G14_p_spl_1;
  wire G14_n_spl_;
  wire G14_n_spl_0;
  wire G14_n_spl_1;
  wire g2560_n_spl_;
  wire g2559_p_spl_;
  wire g2560_p_spl_;
  wire g2559_n_spl_;
  wire g2561_n_spl_;
  wire g2561_p_spl_;
  wire g2562_n_spl_;
  wire g2562_n_spl_0;
  wire g2562_p_spl_;
  wire g2562_p_spl_0;
  wire g2566_n_spl_;
  wire g2565_p_spl_;
  wire g2566_p_spl_;
  wire g2565_n_spl_;
  wire g2567_n_spl_;
  wire g2567_p_spl_;
  wire g2568_n_spl_;
  wire g2568_n_spl_0;
  wire g2564_n_spl_;
  wire g2568_p_spl_;
  wire g2568_p_spl_0;
  wire g2564_p_spl_;
  wire g2569_n_spl_;
  wire g2569_n_spl_0;
  wire g2569_p_spl_;
  wire g2569_p_spl_0;
  wire g2573_n_spl_;
  wire g2572_n_spl_;
  wire g2573_p_spl_;
  wire g2572_p_spl_;
  wire g2574_n_spl_;
  wire g2574_n_spl_0;
  wire g2574_p_spl_;
  wire g2574_p_spl_0;
  wire g2579_n_spl_;
  wire g2579_p_spl_;
  wire g2580_n_spl_;
  wire g2580_n_spl_0;
  wire g2580_p_spl_;
  wire g2580_p_spl_0;
  wire g2584_n_spl_;
  wire g2583_n_spl_;
  wire g2584_p_spl_;
  wire g2583_p_spl_;
  wire g2585_n_spl_;
  wire g2585_n_spl_0;
  wire g2585_p_spl_;
  wire g2585_p_spl_0;
  wire g2586_n_spl_;
  wire g2577_n_spl_;
  wire g2586_p_spl_;
  wire g2577_p_spl_;
  wire g2587_n_spl_;
  wire g2587_n_spl_0;
  wire g2587_p_spl_;
  wire g2592_n_spl_;
  wire g2592_n_spl_0;
  wire g2422_n_spl_;
  wire g2422_n_spl_0;
  wire g2437_n_spl_;
  wire g2437_n_spl_0;
  wire g2452_n_spl_;
  wire g2452_n_spl_0;
  wire g2467_n_spl_;
  wire g2467_n_spl_0;
  wire g2512_n_spl_;
  wire g2332_n_spl_;
  wire g2518_n_spl_;
  wire g2333_n_spl_;
  wire g2515_n_spl_;
  wire g2334_n_spl_;
  wire g2519_p_spl_;
  wire g2335_n_spl_;
  wire g2509_n_spl_;
  wire g2349_n_spl_;
  wire g2506_p_spl_;
  wire g2390_p_spl_;
  wire g2485_n_spl_;
  wire g2613_n_spl_;
  wire g2612_p_spl_;
  wire g2612_n_spl_;
  wire g2614_n_spl_;
  wire g2615_p_spl_;
  wire g2621_n_spl_;
  wire g2621_p_spl_;
  wire g2622_n_spl_;
  wire g2622_n_spl_0;
  wire g2622_p_spl_;
  wire g2622_p_spl_0;
  wire g2626_p_spl_;
  wire g2625_p_spl_;
  wire g2627_p_spl_;
  wire g2627_p_spl_0;
  wire g2634_n_spl_;
  wire g2634_p_spl_;
  wire g2635_n_spl_;
  wire g2635_n_spl_0;
  wire g2635_p_spl_;
  wire g2635_p_spl_0;
  wire g2639_n_spl_;
  wire g2638_n_spl_;
  wire g2639_p_spl_;
  wire g2638_p_spl_;
  wire g2640_n_spl_;
  wire g2640_n_spl_0;
  wire g2640_p_spl_;
  wire g2640_p_spl_0;
  wire g2641_n_spl_;
  wire g2632_n_spl_;
  wire g2641_p_spl_;
  wire g2632_p_spl_;
  wire g2642_n_spl_;
  wire g2642_n_spl_0;
  wire g2642_p_spl_;
  wire g2646_n_spl_;
  wire g2645_n_spl_;
  wire g2646_p_spl_;
  wire g2645_p_spl_;
  wire g2647_n_spl_;
  wire g2647_n_spl_0;
  wire g2647_p_spl_;
  wire g2654_n_spl_;
  wire g2653_n_spl_;
  wire g2654_p_spl_;
  wire g2653_p_spl_;
  wire g2655_n_spl_;
  wire g2655_n_spl_0;
  wire g2655_p_spl_;
  wire g2655_p_spl_0;
  wire g2659_p_spl_;
  wire g2658_p_spl_;
  wire g2660_p_spl_;
  wire g2660_p_spl_0;
  wire g2215_n_spl_;
  wire g2215_n_spl_0;
  wire g2241_n_spl_;
  wire g2241_n_spl_0;
  wire g2286_n_spl_;
  wire g2286_n_spl_0;
  wire g2297_n_spl_;
  wire g2297_n_spl_0;
  wire g2330_n_spl_;
  wire g2330_n_spl_0;
  wire g2607_p_spl_;
  wire g2694_n_spl_;
  wire g2694_p_spl_;
  wire g2695_n_spl_;
  wire g2695_n_spl_0;
  wire g2695_p_spl_;
  wire g2700_n_spl_;
  wire g2700_n_spl_0;
  wire g2705_n_spl_;
  wire g2704_n_spl_;
  wire g2705_p_spl_;
  wire g2704_p_spl_;
  wire g2706_n_spl_;
  wire g2706_n_spl_0;
  wire g2706_p_spl_;
  wire g2711_n_spl_;
  wire g2711_n_spl_0;
  wire g2616_n_spl_;
  wire g2616_n_spl_0;
  wire g2629_n_spl_;
  wire g2629_n_spl_0;
  wire g2662_n_spl_;
  wire g2662_n_spl_0;
  wire g2688_n_spl_;
  wire g2523_n_spl_;
  wire g2685_n_spl_;
  wire g2524_n_spl_;
  wire g2679_n_spl_;
  wire g2541_n_spl_;
  wire g2541_n_spl_0;
  wire g2682_p_spl_;
  wire g2558_p_spl_;
  wire g2677_p_spl_;
  wire g2593_p_spl_;
  wire g2409_n_spl_;
  wire g2409_n_spl_0;
  wire g2486_n_spl_;
  wire g2486_n_spl_0;
  wire g2503_n_spl_;
  wire g2503_n_spl_0;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    n2491_lo_p,
    n2491_lo
  );


  not

  (
    n2491_lo_n,
    n2491_lo
  );


  buf

  (
    n2575_lo_p,
    n2575_lo
  );


  not

  (
    n2575_lo_n,
    n2575_lo
  );


  buf

  (
    n2587_lo_p,
    n2587_lo
  );


  not

  (
    n2587_lo_n,
    n2587_lo
  );


  buf

  (
    n2599_lo_p,
    n2599_lo
  );


  not

  (
    n2599_lo_n,
    n2599_lo
  );


  buf

  (
    n2611_lo_p,
    n2611_lo
  );


  not

  (
    n2611_lo_n,
    n2611_lo
  );


  buf

  (
    n2623_lo_p,
    n2623_lo
  );


  not

  (
    n2623_lo_n,
    n2623_lo
  );


  buf

  (
    n2635_lo_p,
    n2635_lo
  );


  not

  (
    n2635_lo_n,
    n2635_lo
  );


  buf

  (
    n2647_lo_p,
    n2647_lo
  );


  not

  (
    n2647_lo_n,
    n2647_lo
  );


  buf

  (
    n2659_lo_p,
    n2659_lo
  );


  not

  (
    n2659_lo_n,
    n2659_lo
  );


  buf

  (
    n2671_lo_p,
    n2671_lo
  );


  not

  (
    n2671_lo_n,
    n2671_lo
  );


  buf

  (
    n2683_lo_p,
    n2683_lo
  );


  not

  (
    n2683_lo_n,
    n2683_lo
  );


  buf

  (
    n2734_lo_p,
    n2734_lo
  );


  not

  (
    n2734_lo_n,
    n2734_lo
  );


  buf

  (
    n2746_lo_p,
    n2746_lo
  );


  not

  (
    n2746_lo_n,
    n2746_lo
  );


  buf

  (
    n2758_lo_p,
    n2758_lo
  );


  not

  (
    n2758_lo_n,
    n2758_lo
  );


  buf

  (
    n2770_lo_p,
    n2770_lo
  );


  not

  (
    n2770_lo_n,
    n2770_lo
  );


  buf

  (
    n2782_lo_p,
    n2782_lo
  );


  not

  (
    n2782_lo_n,
    n2782_lo
  );


  buf

  (
    n2785_lo_p,
    n2785_lo
  );


  not

  (
    n2785_lo_n,
    n2785_lo
  );


  buf

  (
    n2794_lo_p,
    n2794_lo
  );


  not

  (
    n2794_lo_n,
    n2794_lo
  );


  buf

  (
    n2797_lo_p,
    n2797_lo
  );


  not

  (
    n2797_lo_n,
    n2797_lo
  );


  buf

  (
    n2806_lo_p,
    n2806_lo
  );


  not

  (
    n2806_lo_n,
    n2806_lo
  );


  buf

  (
    n2809_lo_p,
    n2809_lo
  );


  not

  (
    n2809_lo_n,
    n2809_lo
  );


  buf

  (
    n2818_lo_p,
    n2818_lo
  );


  not

  (
    n2818_lo_n,
    n2818_lo
  );


  buf

  (
    n2821_lo_p,
    n2821_lo
  );


  not

  (
    n2821_lo_n,
    n2821_lo
  );


  buf

  (
    n2830_lo_p,
    n2830_lo
  );


  not

  (
    n2830_lo_n,
    n2830_lo
  );


  buf

  (
    n2833_lo_p,
    n2833_lo
  );


  not

  (
    n2833_lo_n,
    n2833_lo
  );


  buf

  (
    n2836_lo_p,
    n2836_lo
  );


  not

  (
    n2836_lo_n,
    n2836_lo
  );


  buf

  (
    n2839_lo_p,
    n2839_lo
  );


  not

  (
    n2839_lo_n,
    n2839_lo
  );


  buf

  (
    n2842_lo_p,
    n2842_lo
  );


  not

  (
    n2842_lo_n,
    n2842_lo
  );


  buf

  (
    n2845_lo_p,
    n2845_lo
  );


  not

  (
    n2845_lo_n,
    n2845_lo
  );


  buf

  (
    n2848_lo_p,
    n2848_lo
  );


  not

  (
    n2848_lo_n,
    n2848_lo
  );


  buf

  (
    n2851_lo_p,
    n2851_lo
  );


  not

  (
    n2851_lo_n,
    n2851_lo
  );


  buf

  (
    n2854_lo_p,
    n2854_lo
  );


  not

  (
    n2854_lo_n,
    n2854_lo
  );


  buf

  (
    n2857_lo_p,
    n2857_lo
  );


  not

  (
    n2857_lo_n,
    n2857_lo
  );


  buf

  (
    n2860_lo_p,
    n2860_lo
  );


  not

  (
    n2860_lo_n,
    n2860_lo
  );


  buf

  (
    n2863_lo_p,
    n2863_lo
  );


  not

  (
    n2863_lo_n,
    n2863_lo
  );


  buf

  (
    n4871_o2_p,
    n4871_o2
  );


  not

  (
    n4871_o2_n,
    n4871_o2
  );


  buf

  (
    n4893_o2_p,
    n4893_o2
  );


  not

  (
    n4893_o2_n,
    n4893_o2
  );


  buf

  (
    n4938_o2_p,
    n4938_o2
  );


  not

  (
    n4938_o2_n,
    n4938_o2
  );


  buf

  (
    n5056_o2_p,
    n5056_o2
  );


  not

  (
    n5056_o2_n,
    n5056_o2
  );


  buf

  (
    n5100_o2_p,
    n5100_o2
  );


  not

  (
    n5100_o2_n,
    n5100_o2
  );


  buf

  (
    n5122_o2_p,
    n5122_o2
  );


  not

  (
    n5122_o2_n,
    n5122_o2
  );


  buf

  (
    n5254_o2_p,
    n5254_o2
  );


  not

  (
    n5254_o2_n,
    n5254_o2
  );


  buf

  (
    n5276_o2_p,
    n5276_o2
  );


  not

  (
    n5276_o2_n,
    n5276_o2
  );


  buf

  (
    n5316_o2_p,
    n5316_o2
  );


  not

  (
    n5316_o2_n,
    n5316_o2
  );


  buf

  (
    n5434_o2_p,
    n5434_o2
  );


  not

  (
    n5434_o2_n,
    n5434_o2
  );


  buf

  (
    n5473_o2_p,
    n5473_o2
  );


  not

  (
    n5473_o2_n,
    n5473_o2
  );


  buf

  (
    n5494_o2_p,
    n5494_o2
  );


  not

  (
    n5494_o2_n,
    n5494_o2
  );


  buf

  (
    n5620_o2_p,
    n5620_o2
  );


  not

  (
    n5620_o2_n,
    n5620_o2
  );


  buf

  (
    n5643_o2_p,
    n5643_o2
  );


  not

  (
    n5643_o2_n,
    n5643_o2
  );


  buf

  (
    n5682_o2_p,
    n5682_o2
  );


  not

  (
    n5682_o2_n,
    n5682_o2
  );


  buf

  (
    n5798_o2_p,
    n5798_o2
  );


  not

  (
    n5798_o2_n,
    n5798_o2
  );


  buf

  (
    n5839_o2_p,
    n5839_o2
  );


  not

  (
    n5839_o2_n,
    n5839_o2
  );


  buf

  (
    n5867_o2_p,
    n5867_o2
  );


  not

  (
    n5867_o2_n,
    n5867_o2
  );


  buf

  (
    n6052_o2_p,
    n6052_o2
  );


  not

  (
    n6052_o2_n,
    n6052_o2
  );


  buf

  (
    n6087_o2_p,
    n6087_o2
  );


  not

  (
    n6087_o2_n,
    n6087_o2
  );


  buf

  (
    n6153_o2_p,
    n6153_o2
  );


  not

  (
    n6153_o2_n,
    n6153_o2
  );


  buf

  (
    n6408_o2_p,
    n6408_o2
  );


  not

  (
    n6408_o2_n,
    n6408_o2
  );


  buf

  (
    n6454_o2_p,
    n6454_o2
  );


  not

  (
    n6454_o2_n,
    n6454_o2
  );


  buf

  (
    n6509_o2_p,
    n6509_o2
  );


  not

  (
    n6509_o2_n,
    n6509_o2
  );


  buf

  (
    n6775_o2_p,
    n6775_o2
  );


  not

  (
    n6775_o2_n,
    n6775_o2
  );


  buf

  (
    n6818_o2_p,
    n6818_o2
  );


  not

  (
    n6818_o2_n,
    n6818_o2
  );


  buf

  (
    n6892_o2_p,
    n6892_o2
  );


  not

  (
    n6892_o2_n,
    n6892_o2
  );


  buf

  (
    n5779_o2_p,
    n5779_o2
  );


  not

  (
    n5779_o2_n,
    n5779_o2
  );


  buf

  (
    n5780_o2_p,
    n5780_o2
  );


  not

  (
    n5780_o2_n,
    n5780_o2
  );


  buf

  (
    n7156_o2_p,
    n7156_o2
  );


  not

  (
    n7156_o2_n,
    n7156_o2
  );


  buf

  (
    n5792_o2_p,
    n5792_o2
  );


  not

  (
    n5792_o2_n,
    n5792_o2
  );


  buf

  (
    n7205_o2_p,
    n7205_o2
  );


  not

  (
    n7205_o2_n,
    n7205_o2
  );


  buf

  (
    n5842_o2_p,
    n5842_o2
  );


  not

  (
    n5842_o2_n,
    n5842_o2
  );


  buf

  (
    n5863_o2_p,
    n5863_o2
  );


  not

  (
    n5863_o2_n,
    n5863_o2
  );


  buf

  (
    n7263_o2_p,
    n7263_o2
  );


  not

  (
    n7263_o2_n,
    n7263_o2
  );


  buf

  (
    n5881_o2_p,
    n5881_o2
  );


  not

  (
    n5881_o2_n,
    n5881_o2
  );


  buf

  (
    n5930_o2_p,
    n5930_o2
  );


  not

  (
    n5930_o2_n,
    n5930_o2
  );


  buf

  (
    n5959_o2_p,
    n5959_o2
  );


  not

  (
    n5959_o2_n,
    n5959_o2
  );


  buf

  (
    n5981_o2_p,
    n5981_o2
  );


  not

  (
    n5981_o2_n,
    n5981_o2
  );


  buf

  (
    n6042_o2_p,
    n6042_o2
  );


  not

  (
    n6042_o2_n,
    n6042_o2
  );


  buf

  (
    n6075_o2_p,
    n6075_o2
  );


  not

  (
    n6075_o2_n,
    n6075_o2
  );


  buf

  (
    n6103_o2_p,
    n6103_o2
  );


  not

  (
    n6103_o2_n,
    n6103_o2
  );


  buf

  (
    n7610_o2_p,
    n7610_o2
  );


  not

  (
    n7610_o2_n,
    n7610_o2
  );


  buf

  (
    n6169_o2_p,
    n6169_o2
  );


  not

  (
    n6169_o2_n,
    n6169_o2
  );


  buf

  (
    n7665_o2_p,
    n7665_o2
  );


  not

  (
    n7665_o2_n,
    n7665_o2
  );


  buf

  (
    n6205_o2_p,
    n6205_o2
  );


  not

  (
    n6205_o2_n,
    n6205_o2
  );


  buf

  (
    n6239_o2_p,
    n6239_o2
  );


  not

  (
    n6239_o2_n,
    n6239_o2
  );


  buf

  (
    n7788_o2_p,
    n7788_o2
  );


  not

  (
    n7788_o2_n,
    n7788_o2
  );


  buf

  (
    n6309_o2_p,
    n6309_o2
  );


  not

  (
    n6309_o2_n,
    n6309_o2
  );


  buf

  (
    n6461_o2_p,
    n6461_o2
  );


  not

  (
    n6461_o2_n,
    n6461_o2
  );


  buf

  (
    n6476_o2_p,
    n6476_o2
  );


  not

  (
    n6476_o2_n,
    n6476_o2
  );


  buf

  (
    n325_inv_p,
    n325_inv
  );


  not

  (
    n325_inv_n,
    n325_inv
  );


  buf

  (
    n6545_o2_p,
    n6545_o2
  );


  not

  (
    n6545_o2_n,
    n6545_o2
  );


  buf

  (
    G578_o2_p,
    G578_o2
  );


  not

  (
    G578_o2_n,
    G578_o2
  );


  buf

  (
    G5106_o2_p,
    G5106_o2
  );


  not

  (
    G5106_o2_n,
    G5106_o2
  );


  buf

  (
    n6713_o2_p,
    n6713_o2
  );


  not

  (
    n6713_o2_n,
    n6713_o2
  );


  buf

  (
    G5164_o2_p,
    G5164_o2
  );


  not

  (
    G5164_o2_n,
    G5164_o2
  );


  buf

  (
    n343_inv_p,
    n343_inv
  );


  not

  (
    n343_inv_n,
    n343_inv
  );


  buf

  (
    n6810_o2_p,
    n6810_o2
  );


  not

  (
    n6810_o2_n,
    n6810_o2
  );


  buf

  (
    n6973_o2_p,
    n6973_o2
  );


  not

  (
    n6973_o2_n,
    n6973_o2
  );


  buf

  (
    n352_inv_p,
    n352_inv
  );


  not

  (
    n352_inv_n,
    n352_inv
  );


  buf

  (
    n7053_o2_p,
    n7053_o2
  );


  not

  (
    n7053_o2_n,
    n7053_o2
  );


  buf

  (
    G581_o2_p,
    G581_o2
  );


  not

  (
    G581_o2_n,
    G581_o2
  );


  buf

  (
    G5467_o2_p,
    G5467_o2
  );


  not

  (
    G5467_o2_n,
    G5467_o2
  );


  buf

  (
    n7231_o2_p,
    n7231_o2
  );


  not

  (
    n7231_o2_n,
    n7231_o2
  );


  buf

  (
    G5527_o2_p,
    G5527_o2
  );


  not

  (
    G5527_o2_n,
    G5527_o2
  );


  buf

  (
    n370_inv_p,
    n370_inv
  );


  not

  (
    n370_inv_n,
    n370_inv
  );


  buf

  (
    n7304_o2_p,
    n7304_o2
  );


  not

  (
    n7304_o2_n,
    n7304_o2
  );


  buf

  (
    n7530_o2_p,
    n7530_o2
  );


  not

  (
    n7530_o2_n,
    n7530_o2
  );


  buf

  (
    n379_inv_p,
    n379_inv
  );


  not

  (
    n379_inv_n,
    n379_inv
  );


  buf

  (
    n7653_o2_p,
    n7653_o2
  );


  not

  (
    n7653_o2_n,
    n7653_o2
  );


  buf

  (
    G584_o2_p,
    G584_o2
  );


  not

  (
    G584_o2_n,
    G584_o2
  );


  buf

  (
    G5820_o2_p,
    G5820_o2
  );


  not

  (
    G5820_o2_n,
    G5820_o2
  );


  buf

  (
    n7148_o2_p,
    n7148_o2
  );


  not

  (
    n7148_o2_n,
    n7148_o2
  );


  buf

  (
    n7149_o2_p,
    n7149_o2
  );


  not

  (
    n7149_o2_n,
    n7149_o2
  );


  buf

  (
    n7224_o2_p,
    n7224_o2
  );


  not

  (
    n7224_o2_n,
    n7224_o2
  );


  buf

  (
    n7916_o2_p,
    n7916_o2
  );


  not

  (
    n7916_o2_n,
    n7916_o2
  );


  buf

  (
    G5868_o2_p,
    G5868_o2
  );


  not

  (
    G5868_o2_n,
    G5868_o2
  );


  buf

  (
    n406_inv_p,
    n406_inv
  );


  not

  (
    n406_inv_n,
    n406_inv
  );


  buf

  (
    n7280_o2_p,
    n7280_o2
  );


  not

  (
    n7280_o2_n,
    n7280_o2
  );


  buf

  (
    n7313_o2_p,
    n7313_o2
  );


  not

  (
    n7313_o2_n,
    n7313_o2
  );


  buf

  (
    n8056_o2_p,
    n8056_o2
  );


  not

  (
    n8056_o2_n,
    n8056_o2
  );


  buf

  (
    n7323_o2_p,
    n7323_o2
  );


  not

  (
    n7323_o2_n,
    n7323_o2
  );


  buf

  (
    n7398_o2_p,
    n7398_o2
  );


  not

  (
    n7398_o2_n,
    n7398_o2
  );


  buf

  (
    n7459_o2_p,
    n7459_o2
  );


  not

  (
    n7459_o2_n,
    n7459_o2
  );


  buf

  (
    n7501_o2_p,
    n7501_o2
  );


  not

  (
    n7501_o2_n,
    n7501_o2
  );


  buf

  (
    n7518_o2_p,
    n7518_o2
  );


  not

  (
    n7518_o2_n,
    n7518_o2
  );


  buf

  (
    G563_o2_p,
    G563_o2
  );


  not

  (
    G563_o2_n,
    G563_o2
  );


  buf

  (
    n7606_o2_p,
    n7606_o2
  );


  not

  (
    n7606_o2_n,
    n7606_o2
  );


  buf

  (
    n439_inv_p,
    n439_inv
  );


  not

  (
    n439_inv_n,
    n439_inv
  );


  buf

  (
    n7675_o2_p,
    n7675_o2
  );


  not

  (
    n7675_o2_n,
    n7675_o2
  );


  buf

  (
    G3410_o2_p,
    G3410_o2
  );


  not

  (
    G3410_o2_n,
    G3410_o2
  );


  buf

  (
    n7722_o2_p,
    n7722_o2
  );


  not

  (
    n7722_o2_n,
    n7722_o2
  );


  buf

  (
    n7747_o2_p,
    n7747_o2
  );


  not

  (
    n7747_o2_n,
    n7747_o2
  );


  buf

  (
    n7835_o2_p,
    n7835_o2
  );


  not

  (
    n7835_o2_n,
    n7835_o2
  );


  buf

  (
    G587_o2_p,
    G587_o2
  );


  not

  (
    G587_o2_n,
    G587_o2
  );


  buf

  (
    G6046_o2_p,
    G6046_o2
  );


  not

  (
    G6046_o2_n,
    G6046_o2
  );


  buf

  (
    n7909_o2_p,
    n7909_o2
  );


  not

  (
    n7909_o2_n,
    n7909_o2
  );


  buf

  (
    G566_o2_p,
    G566_o2
  );


  not

  (
    G566_o2_n,
    G566_o2
  );


  buf

  (
    G6070_o2_p,
    G6070_o2
  );


  not

  (
    G6070_o2_n,
    G6070_o2
  );


  buf

  (
    n472_inv_p,
    n472_inv
  );


  not

  (
    n472_inv_n,
    n472_inv
  );


  buf

  (
    n8086_o2_p,
    n8086_o2
  );


  not

  (
    n8086_o2_n,
    n8086_o2
  );


  buf

  (
    n8093_o2_p,
    n8093_o2
  );


  not

  (
    n8093_o2_n,
    n8093_o2
  );


  buf

  (
    G3752_o2_p,
    G3752_o2
  );


  not

  (
    G3752_o2_n,
    G3752_o2
  );


  buf

  (
    n484_inv_p,
    n484_inv
  );


  not

  (
    n484_inv_n,
    n484_inv
  );


  buf

  (
    n8199_o2_p,
    n8199_o2
  );


  not

  (
    n8199_o2_n,
    n8199_o2
  );


  buf

  (
    n2800_lo_buf_o2_p,
    n2800_lo_buf_o2
  );


  not

  (
    n2800_lo_buf_o2_n,
    n2800_lo_buf_o2
  );


  buf

  (
    G548_o2_p,
    G548_o2
  );


  not

  (
    G548_o2_n,
    G548_o2
  );


  buf

  (
    n496_inv_p,
    n496_inv
  );


  not

  (
    n496_inv_n,
    n496_inv
  );


  buf

  (
    G569_o2_p,
    G569_o2
  );


  not

  (
    G569_o2_n,
    G569_o2
  );


  buf

  (
    G1761_o2_p,
    G1761_o2
  );


  not

  (
    G1761_o2_n,
    G1761_o2
  );


  buf

  (
    n505_inv_p,
    n505_inv
  );


  not

  (
    n505_inv_n,
    n505_inv
  );


  buf

  (
    G4101_o2_p,
    G4101_o2
  );


  not

  (
    G4101_o2_n,
    G4101_o2
  );


  buf

  (
    G551_o2_p,
    G551_o2
  );


  not

  (
    G551_o2_n,
    G551_o2
  );


  buf

  (
    n514_inv_p,
    n514_inv
  );


  not

  (
    n514_inv_n,
    n514_inv
  );


  buf

  (
    G4743_o2_p,
    G4743_o2
  );


  not

  (
    G4743_o2_n,
    G4743_o2
  );


  buf

  (
    G5271_o2_p,
    G5271_o2
  );


  not

  (
    G5271_o2_n,
    G5271_o2
  );


  buf

  (
    G5790_o2_p,
    G5790_o2
  );


  not

  (
    G5790_o2_n,
    G5790_o2
  );


  buf

  (
    G6122_o2_p,
    G6122_o2
  );


  not

  (
    G6122_o2_n,
    G6122_o2
  );


  buf

  (
    G2082_o2_p,
    G2082_o2
  );


  not

  (
    G2082_o2_n,
    G2082_o2
  );


  buf

  (
    n2812_lo_buf_o2_p,
    n2812_lo_buf_o2
  );


  not

  (
    n2812_lo_buf_o2_n,
    n2812_lo_buf_o2
  );


  buf

  (
    n2668_lo_buf_o2_p,
    n2668_lo_buf_o2
  );


  not

  (
    n2668_lo_buf_o2_n,
    n2668_lo_buf_o2
  );


  buf

  (
    n2680_lo_buf_o2_p,
    n2680_lo_buf_o2
  );


  not

  (
    n2680_lo_buf_o2_n,
    n2680_lo_buf_o2
  );


  buf

  (
    G572_o2_p,
    G572_o2
  );


  not

  (
    G572_o2_n,
    G572_o2
  );


  buf

  (
    G6125_o2_p,
    G6125_o2
  );


  not

  (
    G6125_o2_n,
    G6125_o2
  );


  buf

  (
    n547_inv_p,
    n547_inv
  );


  not

  (
    n547_inv_n,
    n547_inv
  );


  buf

  (
    n2656_lo_buf_o2_p,
    n2656_lo_buf_o2
  );


  not

  (
    n2656_lo_buf_o2_n,
    n2656_lo_buf_o2
  );


  buf

  (
    G554_o2_p,
    G554_o2
  );


  not

  (
    G554_o2_n,
    G554_o2
  );


  buf

  (
    G4452_o2_p,
    G4452_o2
  );


  not

  (
    G4452_o2_n,
    G4452_o2
  );


  buf

  (
    n559_inv_p,
    n559_inv
  );


  not

  (
    n559_inv_n,
    n559_inv
  );


  buf

  (
    n2644_lo_buf_o2_p,
    n2644_lo_buf_o2
  );


  not

  (
    n2644_lo_buf_o2_n,
    n2644_lo_buf_o2
  );


  buf

  (
    G2410_o2_p,
    G2410_o2
  );


  not

  (
    G2410_o2_n,
    G2410_o2
  );


  buf

  (
    n2632_lo_buf_o2_p,
    n2632_lo_buf_o2
  );


  not

  (
    n2632_lo_buf_o2_n,
    n2632_lo_buf_o2
  );


  buf

  (
    n2620_lo_buf_o2_p,
    n2620_lo_buf_o2
  );


  not

  (
    n2620_lo_buf_o2_n,
    n2620_lo_buf_o2
  );


  buf

  (
    G6131_o2_p,
    G6131_o2
  );


  not

  (
    G6131_o2_n,
    G6131_o2
  );


  buf

  (
    G4693_o2_p,
    G4693_o2
  );


  not

  (
    G4693_o2_n,
    G4693_o2
  );


  buf

  (
    G5209_o2_p,
    G5209_o2
  );


  not

  (
    G5209_o2_n,
    G5209_o2
  );


  buf

  (
    G5741_o2_p,
    G5741_o2
  );


  not

  (
    G5741_o2_n,
    G5741_o2
  );


  buf

  (
    G6082_o2_p,
    G6082_o2
  );


  not

  (
    G6082_o2_n,
    G6082_o2
  );


  buf

  (
    G6119_o2_p,
    G6119_o2
  );


  not

  (
    G6119_o2_n,
    G6119_o2
  );


  buf

  (
    n2608_lo_buf_o2_p,
    n2608_lo_buf_o2
  );


  not

  (
    n2608_lo_buf_o2_n,
    n2608_lo_buf_o2
  );


  buf

  (
    n2596_lo_buf_o2_p,
    n2596_lo_buf_o2
  );


  not

  (
    n2596_lo_buf_o2_n,
    n2596_lo_buf_o2
  );


  buf

  (
    n2584_lo_buf_o2_p,
    n2584_lo_buf_o2
  );


  not

  (
    n2584_lo_buf_o2_n,
    n2584_lo_buf_o2
  );


  buf

  (
    n2572_lo_buf_o2_p,
    n2572_lo_buf_o2
  );


  not

  (
    n2572_lo_buf_o2_n,
    n2572_lo_buf_o2
  );


  buf

  (
    n2704_lo_buf_o2_p,
    n2704_lo_buf_o2
  );


  not

  (
    n2704_lo_buf_o2_n,
    n2704_lo_buf_o2
  );


  buf

  (
    G557_o2_p,
    G557_o2
  );


  not

  (
    G557_o2_n,
    G557_o2
  );


  buf

  (
    G5936_o2_p,
    G5936_o2
  );


  not

  (
    G5936_o2_n,
    G5936_o2
  );


  buf

  (
    G5442_o2_p,
    G5442_o2
  );


  not

  (
    G5442_o2_n,
    G5442_o2
  );


  buf

  (
    G4926_o2_p,
    G4926_o2
  );


  not

  (
    G4926_o2_n,
    G4926_o2
  );


  buf

  (
    G6134_o2_p,
    G6134_o2
  );


  not

  (
    G6134_o2_n,
    G6134_o2
  );


  buf

  (
    G3929_o2_p,
    G3929_o2
  );


  not

  (
    G3929_o2_n,
    G3929_o2
  );


  buf

  (
    G4425_o2_p,
    G4425_o2
  );


  not

  (
    G4425_o2_n,
    G4425_o2
  );


  buf

  (
    G4947_o2_p,
    G4947_o2
  );


  not

  (
    G4947_o2_n,
    G4947_o2
  );


  buf

  (
    n2764_lo_buf_o2_p,
    n2764_lo_buf_o2
  );


  not

  (
    n2764_lo_buf_o2_n,
    n2764_lo_buf_o2
  );


  buf

  (
    n634_inv_p,
    n634_inv
  );


  not

  (
    n634_inv_n,
    n634_inv
  );


  buf

  (
    n2560_lo_buf_o2_p,
    n2560_lo_buf_o2
  );


  not

  (
    n2560_lo_buf_o2_n,
    n2560_lo_buf_o2
  );


  buf

  (
    n2824_lo_buf_o2_p,
    n2824_lo_buf_o2
  );


  not

  (
    n2824_lo_buf_o2_n,
    n2824_lo_buf_o2
  );


  buf

  (
    G575_o2_p,
    G575_o2
  );


  not

  (
    G575_o2_n,
    G575_o2
  );


  buf

  (
    G2740_o2_p,
    G2740_o2
  );


  not

  (
    G2740_o2_n,
    G2740_o2
  );


  buf

  (
    n649_inv_p,
    n649_inv
  );


  not

  (
    n649_inv_n,
    n649_inv
  );


  buf

  (
    n2548_lo_buf_o2_p,
    n2548_lo_buf_o2
  );


  not

  (
    n2548_lo_buf_o2_n,
    n2548_lo_buf_o2
  );


  buf

  (
    n2536_lo_buf_o2_p,
    n2536_lo_buf_o2
  );


  not

  (
    n2536_lo_buf_o2_n,
    n2536_lo_buf_o2
  );


  buf

  (
    n2524_lo_buf_o2_p,
    n2524_lo_buf_o2
  );


  not

  (
    n2524_lo_buf_o2_n,
    n2524_lo_buf_o2
  );


  buf

  (
    G875_o2_p,
    G875_o2
  );


  not

  (
    G875_o2_n,
    G875_o2
  );


  buf

  (
    G1064_o2_p,
    G1064_o2
  );


  not

  (
    G1064_o2_n,
    G1064_o2
  );


  buf

  (
    G1253_o2_p,
    G1253_o2
  );


  not

  (
    G1253_o2_n,
    G1253_o2
  );


  buf

  (
    G6140_o2_p,
    G6140_o2
  );


  not

  (
    G6140_o2_n,
    G6140_o2
  );


  buf

  (
    G5151_o2_p,
    G5151_o2
  );


  not

  (
    G5151_o2_n,
    G5151_o2
  );


  buf

  (
    G5686_o2_p,
    G5686_o2
  );


  not

  (
    G5686_o2_n,
    G5686_o2
  );


  buf

  (
    G6061_o2_p,
    G6061_o2
  );


  not

  (
    G6061_o2_n,
    G6061_o2
  );


  buf

  (
    G4803_o2_p,
    G4803_o2
  );


  not

  (
    G4803_o2_n,
    G4803_o2
  );


  buf

  (
    G5332_o2_p,
    G5332_o2
  );


  not

  (
    G5332_o2_n,
    G5332_o2
  );


  buf

  (
    G5844_o2_p,
    G5844_o2
  );


  not

  (
    G5844_o2_n,
    G5844_o2
  );


  buf

  (
    G6114_o2_p,
    G6114_o2
  );


  not

  (
    G6114_o2_n,
    G6114_o2
  );


  buf

  (
    G4806_o2_p,
    G4806_o2
  );


  not

  (
    G4806_o2_n,
    G4806_o2
  );


  buf

  (
    G3881_o2_p,
    G3881_o2
  );


  not

  (
    G3881_o2_n,
    G3881_o2
  );


  buf

  (
    G4370_o2_p,
    G4370_o2
  );


  not

  (
    G4370_o2_n,
    G4370_o2
  );


  buf

  (
    G4896_o2_p,
    G4896_o2
  );


  not

  (
    G4896_o2_n,
    G4896_o2
  );


  buf

  (
    G5001_o2_p,
    G5001_o2
  );


  not

  (
    G5001_o2_n,
    G5001_o2
  );


  buf

  (
    G3121_o2_p,
    G3121_o2
  );


  not

  (
    G3121_o2_n,
    G3121_o2
  );


  buf

  (
    n2512_lo_buf_o2_p,
    n2512_lo_buf_o2
  );


  not

  (
    n2512_lo_buf_o2_n,
    n2512_lo_buf_o2
  );


  buf

  (
    G4085_o2_p,
    G4085_o2
  );


  not

  (
    G4085_o2_n,
    G4085_o2
  );


  buf

  (
    G4605_o2_p,
    G4605_o2
  );


  not

  (
    G4605_o2_n,
    G4605_o2
  );


  buf

  (
    G5118_o2_p,
    G5118_o2
  );


  not

  (
    G5118_o2_n,
    G5118_o2
  );


  buf

  (
    G4997_o2_p,
    G4997_o2
  );


  not

  (
    G4997_o2_n,
    G4997_o2
  );


  buf

  (
    n2500_lo_buf_o2_p,
    n2500_lo_buf_o2
  );


  not

  (
    n2500_lo_buf_o2_n,
    n2500_lo_buf_o2
  );


  buf

  (
    n2716_lo_buf_o2_p,
    n2716_lo_buf_o2
  );


  not

  (
    n2716_lo_buf_o2_n,
    n2716_lo_buf_o2
  );


  buf

  (
    G560_o2_p,
    G560_o2
  );


  not

  (
    G560_o2_n,
    G560_o2
  );


  buf

  (
    G1895_o2_p,
    G1895_o2
  );


  not

  (
    G1895_o2_n,
    G1895_o2
  );


  buf

  (
    G3064_o2_p,
    G3064_o2
  );


  not

  (
    G3064_o2_n,
    G3064_o2
  );


  buf

  (
    G3269_o2_p,
    G3269_o2
  );


  not

  (
    G3269_o2_n,
    G3269_o2
  );


  buf

  (
    G3569_o2_p,
    G3569_o2
  );


  not

  (
    G3569_o2_n,
    G3569_o2
  );


  buf

  (
    n748_inv_p,
    n748_inv
  );


  not

  (
    n748_inv_n,
    n748_inv
  );


  buf

  (
    G1196_o2_p,
    G1196_o2
  );


  not

  (
    G1196_o2_n,
    G1196_o2
  );


  buf

  (
    G1007_o2_p,
    G1007_o2
  );


  not

  (
    G1007_o2_n,
    G1007_o2
  );


  buf

  (
    G818_o2_p,
    G818_o2
  );


  not

  (
    G818_o2_n,
    G818_o2
  );


  buf

  (
    G674_o2_p,
    G674_o2
  );


  not

  (
    G674_o2_n,
    G674_o2
  );


  buf

  (
    G5041_o2_p,
    G5041_o2
  );


  not

  (
    G5041_o2_n,
    G5041_o2
  );


  buf

  (
    G5562_o2_p,
    G5562_o2
  );


  not

  (
    G5562_o2_n,
    G5562_o2
  );


  buf

  (
    G6005_o2_p,
    G6005_o2
  );


  not

  (
    G6005_o2_n,
    G6005_o2
  );


  buf

  (
    G5214_o2_p,
    G5214_o2
  );


  not

  (
    G5214_o2_n,
    G5214_o2
  );


  buf

  (
    G5746_o2_p,
    G5746_o2
  );


  not

  (
    G5746_o2_n,
    G5746_o2
  );


  buf

  (
    G6087_o2_p,
    G6087_o2
  );


  not

  (
    G6087_o2_n,
    G6087_o2
  );


  buf

  (
    G6086_o2_p,
    G6086_o2
  );


  not

  (
    G6086_o2_n,
    G6086_o2
  );


  buf

  (
    G5745_o2_p,
    G5745_o2
  );


  not

  (
    G5745_o2_n,
    G5745_o2
  );


  buf

  (
    G5213_o2_p,
    G5213_o2
  );


  not

  (
    G5213_o2_n,
    G5213_o2
  );


  buf

  (
    G5893_o2_p,
    G5893_o2
  );


  not

  (
    G5893_o2_n,
    G5893_o2
  );


  buf

  (
    G5391_o2_p,
    G5391_o2
  );


  not

  (
    G5391_o2_n,
    G5391_o2
  );


  buf

  (
    G4864_o2_p,
    G4864_o2
  );


  not

  (
    G4864_o2_n,
    G4864_o2
  );


  buf

  (
    G6143_o2_p,
    G6143_o2
  );


  not

  (
    G6143_o2_n,
    G6143_o2
  );


  buf

  (
    G6008_o2_p,
    G6008_o2
  );


  not

  (
    G6008_o2_n,
    G6008_o2
  );


  buf

  (
    G5565_o2_p,
    G5565_o2
  );


  not

  (
    G5565_o2_n,
    G5565_o2
  );


  buf

  (
    G5044_o2_p,
    G5044_o2
  );


  not

  (
    G5044_o2_n,
    G5044_o2
  );


  buf

  (
    G3813_o2_p,
    G3813_o2
  );


  not

  (
    G3813_o2_n,
    G3813_o2
  );


  buf

  (
    G4325_o2_p,
    G4325_o2
  );


  not

  (
    G4325_o2_n,
    G4325_o2
  );


  buf

  (
    G4834_o2_p,
    G4834_o2
  );


  not

  (
    G4834_o2_n,
    G4834_o2
  );


  buf

  (
    G4993_o2_p,
    G4993_o2
  );


  not

  (
    G4993_o2_n,
    G4993_o2
  );


  buf

  (
    G3989_o2_p,
    G3989_o2
  );


  not

  (
    G3989_o2_n,
    G3989_o2
  );


  buf

  (
    G4490_o2_p,
    G4490_o2
  );


  not

  (
    G4490_o2_n,
    G4490_o2
  );


  buf

  (
    G5011_o2_p,
    G5011_o2
  );


  not

  (
    G5011_o2_n,
    G5011_o2
  );


  buf

  (
    G5112_o2_p,
    G5112_o2
  );


  not

  (
    G5112_o2_n,
    G5112_o2
  );


  buf

  (
    n2776_lo_buf_o2_p,
    n2776_lo_buf_o2
  );


  not

  (
    n2776_lo_buf_o2_n,
    n2776_lo_buf_o2
  );


  buf

  (
    G3298_o2_p,
    G3298_o2
  );


  not

  (
    G3298_o2_n,
    G3298_o2
  );


  buf

  (
    G3073_o2_p,
    G3073_o2
  );


  not

  (
    G3073_o2_n,
    G3073_o2
  );


  buf

  (
    G3265_o2_p,
    G3265_o2
  );


  not

  (
    G3265_o2_n,
    G3265_o2
  );


  buf

  (
    G3624_o2_p,
    G3624_o2
  );


  not

  (
    G3624_o2_n,
    G3624_o2
  );


  buf

  (
    G1642_o2_p,
    G1642_o2
  );


  not

  (
    G1642_o2_n,
    G1642_o2
  );


  buf

  (
    G1980_o2_p,
    G1980_o2
  );


  not

  (
    G1980_o2_n,
    G1980_o2
  );


  buf

  (
    n2488_lo_buf_o2_p,
    n2488_lo_buf_o2
  );


  not

  (
    n2488_lo_buf_o2_n,
    n2488_lo_buf_o2
  );


  buf

  (
    G626_o2_p,
    G626_o2
  );


  not

  (
    G626_o2_n,
    G626_o2
  );


  buf

  (
    G1139_o2_p,
    G1139_o2
  );


  not

  (
    G1139_o2_n,
    G1139_o2
  );


  buf

  (
    G950_o2_p,
    G950_o2
  );


  not

  (
    G950_o2_n,
    G950_o2
  );


  buf

  (
    G707_o2_p,
    G707_o2
  );


  not

  (
    G707_o2_n,
    G707_o2
  );


  buf

  (
    G545_o2_p,
    G545_o2
  );


  not

  (
    G545_o2_n,
    G545_o2
  );


  buf

  (
    G4217_o2_p,
    G4217_o2
  );


  not

  (
    G4217_o2_n,
    G4217_o2
  );


  buf

  (
    G4716_o2_p,
    G4716_o2
  );


  not

  (
    G4716_o2_n,
    G4716_o2
  );


  buf

  (
    G5244_o2_p,
    G5244_o2
  );


  not

  (
    G5244_o2_n,
    G5244_o2
  );


  buf

  (
    G3136_o2_p,
    G3136_o2
  );


  not

  (
    G3136_o2_n,
    G3136_o2
  );


  buf

  (
    G3499_o2_p,
    G3499_o2
  );


  not

  (
    G3499_o2_n,
    G3499_o2
  );


  buf

  (
    G3885_o2_p,
    G3885_o2
  );


  not

  (
    G3885_o2_n,
    G3885_o2
  );


  buf

  (
    G5243_o2_p,
    G5243_o2
  );


  not

  (
    G5243_o2_n,
    G5243_o2
  );


  buf

  (
    G3886_o2_p,
    G3886_o2
  );


  not

  (
    G3886_o2_n,
    G3886_o2
  );


  buf

  (
    G4375_o2_p,
    G4375_o2
  );


  not

  (
    G4375_o2_n,
    G4375_o2
  );


  buf

  (
    G4901_o2_p,
    G4901_o2
  );


  not

  (
    G4901_o2_n,
    G4901_o2
  );


  buf

  (
    G5054_o2_p,
    G5054_o2
  );


  not

  (
    G5054_o2_n,
    G5054_o2
  );


  buf

  (
    G4374_o2_p,
    G4374_o2
  );


  not

  (
    G4374_o2_n,
    G4374_o2
  );


  buf

  (
    G4900_o2_p,
    G4900_o2
  );


  not

  (
    G4900_o2_n,
    G4900_o2
  );


  buf

  (
    G5053_o2_p,
    G5053_o2
  );


  not

  (
    G5053_o2_n,
    G5053_o2
  );


  buf

  (
    G5242_o2_p,
    G5242_o2
  );


  not

  (
    G5242_o2_n,
    G5242_o2
  );


  buf

  (
    G4034_o2_p,
    G4034_o2
  );


  not

  (
    G4034_o2_n,
    G4034_o2
  );


  buf

  (
    G4556_o2_p,
    G4556_o2
  );


  not

  (
    G4556_o2_n,
    G4556_o2
  );


  buf

  (
    G5064_o2_p,
    G5064_o2
  );


  not

  (
    G5064_o2_n,
    G5064_o2
  );


  buf

  (
    G5172_o2_p,
    G5172_o2
  );


  not

  (
    G5172_o2_n,
    G5172_o2
  );


  buf

  (
    G2030_o2_p,
    G2030_o2
  );


  not

  (
    G2030_o2_n,
    G2030_o2
  );


  buf

  (
    G3016_o2_p,
    G3016_o2
  );


  not

  (
    G3016_o2_n,
    G3016_o2
  );


  buf

  (
    G3520_o2_p,
    G3520_o2
  );


  not

  (
    G3520_o2_n,
    G3520_o2
  );


  buf

  (
    G3261_o2_p,
    G3261_o2
  );


  not

  (
    G3261_o2_n,
    G3261_o2
  );


  buf

  (
    G3620_o2_p,
    G3620_o2
  );


  not

  (
    G3620_o2_n,
    G3620_o2
  );


  buf

  (
    G4220_o2_p,
    G4220_o2
  );


  not

  (
    G4220_o2_n,
    G4220_o2
  );


  buf

  (
    G4719_o2_p,
    G4719_o2
  );


  not

  (
    G4719_o2_n,
    G4719_o2
  );


  buf

  (
    G5247_o2_p,
    G5247_o2
  );


  not

  (
    G5247_o2_n,
    G5247_o2
  );


  buf

  (
    G5109_o2_p,
    G5109_o2
  );


  not

  (
    G5109_o2_n,
    G5109_o2
  );


  buf

  (
    G1638_o2_p,
    G1638_o2
  );


  not

  (
    G1638_o2_n,
    G1638_o2
  );


  buf

  (
    G1976_o2_p,
    G1976_o2
  );


  not

  (
    G1976_o2_n,
    G1976_o2
  );


  buf

  (
    G3560_o2_p,
    G3560_o2
  );


  not

  (
    G3560_o2_n,
    G3560_o2
  );


  buf

  (
    G3205_o2_p,
    G3205_o2
  );


  not

  (
    G3205_o2_n,
    G3205_o2
  );


  buf

  (
    G3193_o2_p,
    G3193_o2
  );


  not

  (
    G3193_o2_n,
    G3193_o2
  );


  buf

  (
    G3367_o2_p,
    G3367_o2
  );


  not

  (
    G3367_o2_n,
    G3367_o2
  );


  buf

  (
    G3670_o2_p,
    G3670_o2
  );


  not

  (
    G3670_o2_n,
    G3670_o2
  );


  buf

  (
    n979_inv_p,
    n979_inv
  );


  not

  (
    n979_inv_n,
    n979_inv
  );


  buf

  (
    G1280_o2_p,
    G1280_o2
  );


  not

  (
    G1280_o2_n,
    G1280_o2
  );


  buf

  (
    G902_o2_p,
    G902_o2
  );


  not

  (
    G902_o2_n,
    G902_o2
  );


  buf

  (
    G659_o2_p,
    G659_o2
  );


  not

  (
    G659_o2_n,
    G659_o2
  );


  buf

  (
    G983_o2_p,
    G983_o2
  );


  not

  (
    G983_o2_n,
    G983_o2
  );


  buf

  (
    G740_o2_p,
    G740_o2
  );


  not

  (
    G740_o2_n,
    G740_o2
  );


  buf

  (
    G2917_o2_p,
    G2917_o2
  );


  not

  (
    G2917_o2_n,
    G2917_o2
  );


  buf

  (
    G3391_o2_p,
    G3391_o2
  );


  not

  (
    G3391_o2_n,
    G3391_o2
  );


  buf

  (
    G3494_o2_p,
    G3494_o2
  );


  not

  (
    G3494_o2_n,
    G3494_o2
  );


  buf

  (
    G1512_o2_p,
    G1512_o2
  );


  not

  (
    G1512_o2_n,
    G1512_o2
  );


  buf

  (
    G1854_o2_p,
    G1854_o2
  );


  not

  (
    G1854_o2_n,
    G1854_o2
  );


  buf

  (
    G2203_o2_p,
    G2203_o2
  );


  not

  (
    G2203_o2_n,
    G2203_o2
  );


  buf

  (
    G3493_o2_p,
    G3493_o2
  );


  not

  (
    G3493_o2_n,
    G3493_o2
  );


  buf

  (
    G3069_o2_p,
    G3069_o2
  );


  not

  (
    G3069_o2_n,
    G3069_o2
  );


  buf

  (
    G3574_o2_p,
    G3574_o2
  );


  not

  (
    G3574_o2_n,
    G3574_o2
  );


  buf

  (
    G3319_o2_p,
    G3319_o2
  );


  not

  (
    G3319_o2_n,
    G3319_o2
  );


  buf

  (
    G3667_o2_p,
    G3667_o2
  );


  not

  (
    G3667_o2_n,
    G3667_o2
  );


  buf

  (
    G3068_o2_p,
    G3068_o2
  );


  not

  (
    G3068_o2_n,
    G3068_o2
  );


  buf

  (
    G3573_o2_p,
    G3573_o2
  );


  not

  (
    G3573_o2_n,
    G3573_o2
  );


  buf

  (
    G3666_o2_p,
    G3666_o2
  );


  not

  (
    G3666_o2_n,
    G3666_o2
  );


  buf

  (
    G3318_o2_p,
    G3318_o2
  );


  not

  (
    G3318_o2_n,
    G3318_o2
  );


  buf

  (
    G3492_o2_p,
    G3492_o2
  );


  not

  (
    G3492_o2_n,
    G3492_o2
  );


  buf

  (
    G3241_o2_p,
    G3241_o2
  );


  not

  (
    G3241_o2_n,
    G3241_o2
  );


  buf

  (
    G3722_o2_p,
    G3722_o2
  );


  not

  (
    G3722_o2_n,
    G3722_o2
  );


  buf

  (
    G3422_o2_p,
    G3422_o2
  );


  not

  (
    G3422_o2_n,
    G3422_o2
  );


  buf

  (
    G1445_o2_p,
    G1445_o2
  );


  not

  (
    G1445_o2_n,
    G1445_o2
  );


  buf

  (
    G3257_o2_p,
    G3257_o2
  );


  not

  (
    G3257_o2_n,
    G3257_o2
  );


  buf

  (
    G3616_o2_p,
    G3616_o2
  );


  not

  (
    G3616_o2_n,
    G3616_o2
  );


  buf

  (
    G1634_o2_p,
    G1634_o2
  );


  not

  (
    G1634_o2_n,
    G1634_o2
  );


  buf

  (
    G1972_o2_p,
    G1972_o2
  );


  not

  (
    G1972_o2_n,
    G1972_o2
  );


  buf

  (
    G2256_o2_p,
    G2256_o2
  );


  not

  (
    G2256_o2_n,
    G2256_o2
  );


  buf

  (
    G3394_o2_p,
    G3394_o2
  );


  not

  (
    G3394_o2_n,
    G3394_o2
  );


  buf

  (
    G3557_o2_p,
    G3557_o2
  );


  not

  (
    G3557_o2_n,
    G3557_o2
  );


  buf

  (
    G3364_o2_p,
    G3364_o2
  );


  not

  (
    G3364_o2_n,
    G3364_o2
  );


  buf

  (
    G3719_o2_p,
    G3719_o2
  );


  not

  (
    G3719_o2_n,
    G3719_o2
  );


  buf

  (
    G2253_o2_p,
    G2253_o2
  );


  not

  (
    G2253_o2_n,
    G2253_o2
  );


  buf

  (
    G1583_o2_p,
    G1583_o2
  );


  not

  (
    G1583_o2_n,
    G1583_o2
  );


  buf

  (
    G1917_o2_p,
    G1917_o2
  );


  not

  (
    G1917_o2_n,
    G1917_o2
  );


  buf

  (
    G1727_o2_p,
    G1727_o2
  );


  not

  (
    G1727_o2_n,
    G1727_o2
  );


  buf

  (
    G2061_o2_p,
    G2061_o2
  );


  not

  (
    G2061_o2_n,
    G2061_o2
  );


  buf

  (
    G935_o2_p,
    G935_o2
  );


  not

  (
    G935_o2_n,
    G935_o2
  );


  buf

  (
    G692_o2_p,
    G692_o2
  );


  not

  (
    G692_o2_n,
    G692_o2
  );


  buf

  (
    G2136_o2_p,
    G2136_o2
  );


  not

  (
    G2136_o2_n,
    G2136_o2
  );


  buf

  (
    G1507_o2_p,
    G1507_o2
  );


  not

  (
    G1507_o2_n,
    G1507_o2
  );


  buf

  (
    G1849_o2_p,
    G1849_o2
  );


  not

  (
    G1849_o2_n,
    G1849_o2
  );


  buf

  (
    G2198_o2_p,
    G2198_o2
  );


  not

  (
    G2198_o2_n,
    G2198_o2
  );


  buf

  (
    G2197_o2_p,
    G2197_o2
  );


  not

  (
    G2197_o2_n,
    G2197_o2
  );


  buf

  (
    G1848_o2_p,
    G1848_o2
  );


  not

  (
    G1848_o2_n,
    G1848_o2
  );


  buf

  (
    G1689_o2_p,
    G1689_o2
  );


  not

  (
    G1689_o2_n,
    G1689_o2
  );


  buf

  (
    G2016_o2_p,
    G2016_o2
  );


  not

  (
    G2016_o2_n,
    G2016_o2
  );


  buf

  (
    G2314_o2_p,
    G2314_o2
  );


  not

  (
    G2314_o2_n,
    G2314_o2
  );


  buf

  (
    G2313_o2_p,
    G2313_o2
  );


  not

  (
    G2313_o2_n,
    G2313_o2
  );


  buf

  (
    G1688_o2_p,
    G1688_o2
  );


  not

  (
    G1688_o2_n,
    G1688_o2
  );


  buf

  (
    G2015_o2_p,
    G2015_o2
  );


  not

  (
    G2015_o2_n,
    G2015_o2
  );


  buf

  (
    G1847_o2_p,
    G1847_o2
  );


  not

  (
    G1847_o2_n,
    G1847_o2
  );


  buf

  (
    G2196_o2_p,
    G2196_o2
  );


  not

  (
    G2196_o2_n,
    G2196_o2
  );


  buf

  (
    G2118_o2_p,
    G2118_o2
  );


  not

  (
    G2118_o2_n,
    G2118_o2
  );


  buf

  (
    G1777_o2_p,
    G1777_o2
  );


  not

  (
    G1777_o2_n,
    G1777_o2
  );


  buf

  (
    G1630_o2_p,
    G1630_o2
  );


  not

  (
    G1630_o2_n,
    G1630_o2
  );


  buf

  (
    G1968_o2_p,
    G1968_o2
  );


  not

  (
    G1968_o2_n,
    G1968_o2
  );


  buf

  (
    G2309_o2_p,
    G2309_o2
  );


  not

  (
    G2309_o2_n,
    G2309_o2
  );


  buf

  (
    G2139_o2_p,
    G2139_o2
  );


  not

  (
    G2139_o2_n,
    G2139_o2
  );


  buf

  (
    G1580_o2_p,
    G1580_o2
  );


  not

  (
    G1580_o2_n,
    G1580_o2
  );


  buf

  (
    G2250_o2_p,
    G2250_o2
  );


  not

  (
    G2250_o2_n,
    G2250_o2
  );


  buf

  (
    G1914_o2_p,
    G1914_o2
  );


  not

  (
    G1914_o2_n,
    G1914_o2
  );


  buf

  (
    G1724_o2_p,
    G1724_o2
  );


  not

  (
    G1724_o2_n,
    G1724_o2
  );


  buf

  (
    G2058_o2_p,
    G2058_o2
  );


  not

  (
    G2058_o2_n,
    G2058_o2
  );


  buf

  (
    n2728_lo_buf_o2_p,
    n2728_lo_buf_o2
  );


  not

  (
    n2728_lo_buf_o2_n,
    n2728_lo_buf_o2
  );


  and

  (
    g405_p,
    n2683_lo_p,
    n2491_lo_p
  );


  or

  (
    g406_n,
    n4938_o2_p_spl_,
    n4893_o2_n
  );


  or

  (
    g407_n,
    n4938_o2_p_spl_,
    n4871_o2_p
  );


  and

  (
    g408_p,
    g407_n,
    g406_n
  );


  or

  (
    g409_n,
    n5122_o2_p_spl_,
    n5100_o2_n
  );


  or

  (
    g410_n,
    n5122_o2_p_spl_,
    n5056_o2_p
  );


  and

  (
    g411_p,
    g410_n,
    g409_n
  );


  or

  (
    g412_n,
    n5316_o2_p_spl_,
    n5276_o2_n
  );


  or

  (
    g413_n,
    n5316_o2_p_spl_,
    n5254_o2_p
  );


  and

  (
    g414_p,
    g413_n,
    g412_n
  );


  or

  (
    g415_n,
    n5494_o2_p_spl_,
    n5473_o2_n
  );


  or

  (
    g416_n,
    n5494_o2_p_spl_,
    n5434_o2_p
  );


  and

  (
    g417_p,
    g416_n,
    g415_n
  );


  or

  (
    g418_n,
    n5682_o2_p_spl_,
    n5643_o2_n
  );


  or

  (
    g419_n,
    n5682_o2_p_spl_,
    n5620_o2_p
  );


  and

  (
    g420_p,
    g419_n,
    g418_n
  );


  or

  (
    g421_n,
    n5867_o2_p_spl_,
    n5839_o2_n
  );


  or

  (
    g422_n,
    n5867_o2_p_spl_,
    n5798_o2_p
  );


  and

  (
    g423_p,
    g422_n,
    g421_n
  );


  or

  (
    g424_n,
    n6153_o2_p_spl_,
    n6087_o2_n
  );


  or

  (
    g425_n,
    n6153_o2_p_spl_,
    n6052_o2_p
  );


  and

  (
    g426_p,
    g425_n,
    g424_n
  );


  or

  (
    g427_n,
    n6509_o2_p_spl_,
    n6454_o2_n
  );


  or

  (
    g428_n,
    n6509_o2_p_spl_,
    n6408_o2_p
  );


  and

  (
    g429_p,
    g428_n,
    g427_n
  );


  or

  (
    g430_n,
    n6892_o2_p_spl_,
    n6818_o2_n
  );


  or

  (
    g431_n,
    n6892_o2_p_spl_,
    n6775_o2_p
  );


  and

  (
    g432_p,
    g431_n,
    g430_n
  );


  or

  (
    g433_n,
    n7263_o2_p_spl_,
    n7205_o2_n
  );


  or

  (
    g434_n,
    n7263_o2_p_spl_,
    n7156_o2_p
  );


  and

  (
    g435_p,
    g434_n,
    g433_n
  );


  or

  (
    g436_n,
    n7788_o2_p_spl_,
    n7665_o2_n
  );


  or

  (
    g437_n,
    n7788_o2_p_spl_,
    n7610_o2_p
  );


  and

  (
    g438_p,
    g437_n,
    g436_n
  );


  or

  (
    g439_n,
    G5164_o2_p_spl_,
    G5106_o2_n
  );


  or

  (
    g440_n,
    G5164_o2_p_spl_,
    G578_o2_p
  );


  and

  (
    g441_p,
    g440_n,
    g439_n
  );


  or

  (
    g442_n,
    G5527_o2_p_spl_,
    G5467_o2_n
  );


  or

  (
    g443_n,
    G5527_o2_p_spl_,
    G581_o2_p
  );


  and

  (
    g444_p,
    g443_n,
    g442_n
  );


  or

  (
    g445_n,
    G5868_o2_p_spl_,
    G5820_o2_n
  );


  or

  (
    g446_n,
    G5868_o2_p_spl_,
    G584_o2_p
  );


  and

  (
    g447_p,
    g446_n,
    g445_n
  );


  or

  (
    g448_n,
    G6070_o2_p_spl_,
    G6046_o2_n
  );


  or

  (
    g449_n,
    G6070_o2_p_spl_,
    G587_o2_p
  );


  and

  (
    g450_p,
    g449_n,
    g448_n
  );


  or

  (
    g451_n,
    G6125_o2_p_spl_,
    G6122_o2_n
  );


  and

  (
    g452_p,
    g451_n,
    G6125_o2_p_spl_
  );


  or

  (
    g453_n,
    G6134_o2_p_spl_,
    G6119_o2_n
  );


  or

  (
    g454_n,
    G6134_o2_p_spl_,
    G6131_o2_p
  );


  and

  (
    g455_p,
    g454_n,
    g453_n
  );


  or

  (
    g456_n,
    G6143_o2_p_spl_0,
    G6114_o2_n
  );


  or

  (
    g457_n,
    G6143_o2_p_spl_0,
    G6140_o2_p
  );


  and

  (
    g458_p,
    g457_n,
    g456_n
  );


  and

  (
    g459_p,
    G6086_o2_n,
    G6087_o2_n
  );


  or

  (
    g459_n,
    G6086_o2_p,
    G6087_o2_p
  );


  and

  (
    g460_p,
    G6143_o2_n,
    G6082_o2_p
  );


  or

  (
    g460_n,
    G6143_o2_p_spl_,
    G6082_o2_n
  );


  and

  (
    g461_p,
    g460_n,
    g459_n
  );


  or

  (
    g461_n,
    g460_p_spl_,
    g459_p_spl_
  );


  or

  (
    g462_n,
    g461_p_spl_0,
    g459_p_spl_
  );


  or

  (
    g463_n,
    g461_p_spl_0,
    g460_p_spl_
  );


  and

  (
    g464_p,
    g463_n,
    g462_n
  );


  and

  (
    g465_p,
    G6008_o2_n_spl_,
    G6005_o2_n_spl_
  );


  or

  (
    g465_n,
    G6008_o2_p_spl_,
    G6005_o2_p_spl_
  );


  and

  (
    g466_p,
    g465_n_spl_0,
    G6008_o2_n_spl_
  );


  or

  (
    g466_n,
    g465_p_spl_0,
    G6008_o2_p_spl_
  );


  and

  (
    g467_p,
    g465_n_spl_0,
    G6005_o2_n_spl_
  );


  or

  (
    g467_n,
    g465_p_spl_0,
    G6005_o2_p_spl_
  );


  and

  (
    g468_p,
    g467_n,
    g466_n
  );


  or

  (
    g468_n,
    g467_p,
    g466_p
  );


  and

  (
    g469_p,
    g461_n,
    G6061_o2_p
  );


  or

  (
    g469_n,
    g461_p_spl_,
    G6061_o2_n
  );


  and

  (
    g470_p,
    g469_n,
    g468_n
  );


  or

  (
    g470_n,
    g469_p_spl_,
    g468_p_spl_
  );


  or

  (
    g471_n,
    g470_p_spl_0,
    g468_p_spl_
  );


  or

  (
    g472_n,
    g470_p_spl_0,
    g469_p_spl_
  );


  and

  (
    g473_p,
    g472_n,
    g471_n
  );


  and

  (
    g474_p,
    G5893_o2_n_spl_0,
    G5844_o2_p
  );


  or

  (
    g474_n,
    G5893_o2_p_spl_0,
    G5844_o2_n
  );


  and

  (
    g475_p,
    G5893_o2_n_spl_0,
    G875_o2_n
  );


  or

  (
    g475_n,
    G5893_o2_p_spl_0,
    G875_o2_p
  );


  and

  (
    g476_p,
    g475_n,
    g474_n
  );


  or

  (
    g476_n,
    g475_p,
    g474_p
  );


  and

  (
    g477_p,
    G5936_o2_n,
    G5790_o2_p
  );


  or

  (
    g477_n,
    G5936_o2_p,
    G5790_o2_n
  );


  and

  (
    g478_p,
    g477_n_spl_,
    g476_n_spl_
  );


  or

  (
    g478_n,
    g477_p_spl_,
    g476_p_spl_
  );


  and

  (
    g479_p,
    g478_n_spl_0,
    g476_n_spl_
  );


  or

  (
    g479_n,
    g478_p_spl_0,
    g476_p_spl_
  );


  and

  (
    g480_p,
    g478_n_spl_0,
    g477_n_spl_
  );


  or

  (
    g480_n,
    g478_p_spl_0,
    g477_p_spl_
  );


  and

  (
    g481_p,
    g480_n,
    g479_n
  );


  or

  (
    g481_n,
    g480_p,
    g479_p
  );


  and

  (
    g482_p,
    g470_n,
    g465_n_spl_
  );


  or

  (
    g482_n,
    g470_p_spl_,
    g465_p_spl_
  );


  and

  (
    g483_p,
    g482_n,
    g481_n
  );


  or

  (
    g483_n,
    g482_p_spl_,
    g481_p_spl_
  );


  or

  (
    g484_n,
    g483_p_spl_0,
    g481_p_spl_
  );


  or

  (
    g485_n,
    g483_p_spl_0,
    g482_p_spl_
  );


  and

  (
    g486_p,
    g485_n,
    g484_n
  );


  and

  (
    g487_p,
    G5745_o2_n,
    G5746_o2_n
  );


  or

  (
    g487_n,
    G5745_o2_p,
    G5746_o2_p
  );


  and

  (
    g488_p,
    n2863_lo_p_spl_000,
    n2575_lo_p
  );


  or

  (
    g488_n,
    n2863_lo_n_spl_000,
    n2575_lo_n
  );


  and

  (
    g489_p,
    g488_n_spl_,
    g487_n_spl_
  );


  or

  (
    g489_n,
    g488_p_spl_,
    g487_p_spl_
  );


  and

  (
    g490_p,
    g489_n_spl_0,
    g487_n_spl_
  );


  or

  (
    g490_n,
    g489_p_spl_0,
    g487_p_spl_
  );


  and

  (
    g491_p,
    g489_n_spl_0,
    g488_n_spl_
  );


  or

  (
    g491_n,
    g489_p_spl_0,
    g488_p_spl_
  );


  and

  (
    g492_p,
    g491_n,
    g490_n
  );


  or

  (
    g492_n,
    g491_p,
    g490_p
  );


  and

  (
    g493_p,
    G5893_o2_n_spl_,
    G5741_o2_p
  );


  or

  (
    g493_n,
    G5893_o2_p_spl_,
    G5741_o2_n
  );


  and

  (
    g494_p,
    g493_n_spl_,
    g492_n_spl_
  );


  or

  (
    g494_n,
    g493_p_spl_,
    g492_p_spl_
  );


  and

  (
    g495_p,
    g494_n_spl_0,
    g492_n_spl_
  );


  or

  (
    g495_n,
    g494_p_spl_0,
    g492_p_spl_
  );


  and

  (
    g496_p,
    g494_n_spl_0,
    g493_n_spl_
  );


  or

  (
    g496_n,
    g494_p_spl_0,
    g493_p_spl_
  );


  and

  (
    g497_p,
    g496_n,
    g495_n
  );


  or

  (
    g497_n,
    g496_p,
    g495_p
  );


  and

  (
    g498_p,
    g483_n,
    g478_n_spl_
  );


  or

  (
    g498_n,
    g483_p_spl_,
    g478_p_spl_
  );


  and

  (
    g499_p,
    g498_n,
    g497_n
  );


  or

  (
    g499_n,
    g498_p_spl_,
    g497_p_spl_
  );


  or

  (
    g500_n,
    g499_p_spl_0,
    g497_p_spl_
  );


  or

  (
    g501_n,
    g499_p_spl_0,
    g498_p_spl_
  );


  and

  (
    g502_p,
    g501_n,
    g500_n
  );


  and

  (
    g503_p,
    G5565_o2_n_spl_,
    G5562_o2_n_spl_
  );


  or

  (
    g503_n,
    G5565_o2_p_spl_,
    G5562_o2_p_spl_
  );


  and

  (
    g504_p,
    g503_n_spl_0,
    G5565_o2_n_spl_
  );


  or

  (
    g504_n,
    g503_p_spl_0,
    G5565_o2_p_spl_
  );


  and

  (
    g505_p,
    g503_n_spl_0,
    G5562_o2_n_spl_
  );


  or

  (
    g505_n,
    g503_p_spl_0,
    G5562_o2_p_spl_
  );


  and

  (
    g506_p,
    g505_n,
    g504_n
  );


  or

  (
    g506_n,
    g505_p,
    g504_p
  );


  and

  (
    g507_p,
    n2863_lo_p_spl_000,
    n2587_lo_p
  );


  or

  (
    g507_n,
    n2863_lo_n_spl_000,
    n2587_lo_n
  );


  and

  (
    g508_p,
    g507_n_spl_,
    g506_n_spl_
  );


  or

  (
    g508_n,
    g507_p_spl_,
    g506_p_spl_
  );


  and

  (
    g509_p,
    g508_n_spl_0,
    g506_n_spl_
  );


  or

  (
    g509_n,
    g508_p_spl_0,
    g506_p_spl_
  );


  and

  (
    g510_p,
    g508_n_spl_0,
    g507_n_spl_
  );


  or

  (
    g510_n,
    g508_p_spl_0,
    g507_p_spl_
  );


  and

  (
    g511_p,
    g510_n,
    g509_n
  );


  or

  (
    g511_n,
    g510_p,
    g509_p
  );


  and

  (
    g512_p,
    g489_n_spl_,
    G5686_o2_p
  );


  or

  (
    g512_n,
    g489_p_spl_,
    G5686_o2_n
  );


  and

  (
    g513_p,
    g512_n_spl_,
    g511_n_spl_
  );


  or

  (
    g513_n,
    g512_p_spl_,
    g511_p_spl_
  );


  and

  (
    g514_p,
    g513_n_spl_0,
    g511_n_spl_
  );


  or

  (
    g514_n,
    g513_p_spl_0,
    g511_p_spl_
  );


  and

  (
    g515_p,
    g513_n_spl_0,
    g512_n_spl_
  );


  or

  (
    g515_n,
    g513_p_spl_0,
    g512_p_spl_
  );


  and

  (
    g516_p,
    g515_n,
    g514_n
  );


  or

  (
    g516_n,
    g515_p,
    g514_p
  );


  and

  (
    g517_p,
    g499_n,
    g494_n_spl_
  );


  or

  (
    g517_n,
    g499_p_spl_,
    g494_p_spl_
  );


  and

  (
    g518_p,
    g517_n,
    g516_n
  );


  or

  (
    g518_n,
    g517_p_spl_,
    g516_p_spl_
  );


  or

  (
    g519_n,
    g518_p_spl_0,
    g516_p_spl_
  );


  or

  (
    g520_n,
    g518_p_spl_0,
    g517_p_spl_
  );


  and

  (
    g521_p,
    g520_n,
    g519_n
  );


  and

  (
    g522_p,
    G5391_o2_n_spl_0,
    G5332_o2_p
  );


  or

  (
    g522_n,
    G5391_o2_p_spl_0,
    G5332_o2_n
  );


  and

  (
    g523_p,
    G5391_o2_n_spl_0,
    G1064_o2_n
  );


  or

  (
    g523_n,
    G5391_o2_p_spl_0,
    G1064_o2_p
  );


  and

  (
    g524_p,
    g523_n,
    g522_n
  );


  or

  (
    g524_n,
    g523_p,
    g522_p
  );


  and

  (
    g525_p,
    G5442_o2_n,
    G5271_o2_p
  );


  or

  (
    g525_n,
    G5442_o2_p,
    G5271_o2_n
  );


  and

  (
    g526_p,
    g525_n_spl_,
    g524_n_spl_
  );


  or

  (
    g526_n,
    g525_p_spl_,
    g524_p_spl_
  );


  and

  (
    g527_p,
    g526_n_spl_0,
    g524_n_spl_
  );


  or

  (
    g527_n,
    g526_p_spl_0,
    g524_p_spl_
  );


  and

  (
    g528_p,
    g526_n_spl_0,
    g525_n_spl_
  );


  or

  (
    g528_n,
    g526_p_spl_0,
    g525_p_spl_
  );


  and

  (
    g529_p,
    g528_n,
    g527_n
  );


  or

  (
    g529_n,
    g528_p,
    g527_p
  );


  and

  (
    g530_p,
    n2863_lo_p_spl_00,
    n2599_lo_p
  );


  or

  (
    g530_n,
    n2863_lo_n_spl_00,
    n2599_lo_n
  );


  and

  (
    g531_p,
    g530_n_spl_,
    g529_n_spl_
  );


  or

  (
    g531_n,
    g530_p_spl_,
    g529_p_spl_
  );


  and

  (
    g532_p,
    g531_n_spl_0,
    g529_n_spl_
  );


  or

  (
    g532_n,
    g531_p_spl_0,
    g529_p_spl_
  );


  and

  (
    g533_p,
    g531_n_spl_0,
    g530_n_spl_
  );


  or

  (
    g533_n,
    g531_p_spl_0,
    g530_p_spl_
  );


  and

  (
    g534_p,
    g533_n,
    g532_n
  );


  or

  (
    g534_n,
    g533_p,
    g532_p
  );


  and

  (
    g535_p,
    g508_n_spl_,
    g503_n_spl_
  );


  or

  (
    g535_n,
    g508_p_spl_,
    g503_p_spl_
  );


  and

  (
    g536_p,
    g535_n_spl_,
    g534_n_spl_
  );


  or

  (
    g536_n,
    g535_p_spl_,
    g534_p_spl_
  );


  and

  (
    g537_p,
    g536_n_spl_0,
    g534_n_spl_
  );


  or

  (
    g537_n,
    g536_p_spl_0,
    g534_p_spl_
  );


  and

  (
    g538_p,
    g536_n_spl_0,
    g535_n_spl_
  );


  or

  (
    g538_n,
    g536_p_spl_0,
    g535_p_spl_
  );


  and

  (
    g539_p,
    g538_n,
    g537_n
  );


  or

  (
    g539_n,
    g538_p,
    g537_p
  );


  and

  (
    g540_p,
    g518_n,
    g513_n_spl_
  );


  or

  (
    g540_n,
    g518_p_spl_,
    g513_p_spl_
  );


  and

  (
    g541_p,
    g540_n,
    g539_n
  );


  or

  (
    g541_n,
    g540_p_spl_,
    g539_p_spl_
  );


  or

  (
    g542_n,
    g541_p_spl_0,
    g539_p_spl_
  );


  or

  (
    g543_n,
    g541_p_spl_0,
    g540_p_spl_
  );


  and

  (
    g544_p,
    g543_n,
    g542_n
  );


  and

  (
    g545_p,
    G5213_o2_n,
    G5214_o2_n
  );


  or

  (
    g545_n,
    G5213_o2_p,
    G5214_o2_p
  );


  and

  (
    g546_p,
    n2851_lo_p_spl_00,
    n2623_lo_p_spl_
  );


  or

  (
    g546_n,
    n2851_lo_n_spl_00,
    n2623_lo_n_spl_
  );


  and

  (
    g547_p,
    g546_n_spl_,
    g545_n_spl_
  );


  or

  (
    g547_n,
    g546_p_spl_,
    g545_p_spl_
  );


  and

  (
    g548_p,
    g547_n_spl_0,
    g545_n_spl_
  );


  or

  (
    g548_n,
    g547_p_spl_0,
    g545_p_spl_
  );


  and

  (
    g549_p,
    g547_n_spl_0,
    g546_n_spl_
  );


  or

  (
    g549_n,
    g547_p_spl_0,
    g546_p_spl_
  );


  and

  (
    g550_p,
    g549_n,
    g548_n
  );


  or

  (
    g550_n,
    g549_p,
    g548_p
  );


  and

  (
    g551_p,
    G5391_o2_n_spl_,
    G5209_o2_p
  );


  or

  (
    g551_n,
    G5391_o2_p_spl_,
    G5209_o2_n
  );


  and

  (
    g552_p,
    g551_n_spl_,
    g550_n_spl_
  );


  or

  (
    g552_n,
    g551_p_spl_,
    g550_p_spl_
  );


  and

  (
    g553_p,
    g552_n_spl_0,
    g550_n_spl_
  );


  or

  (
    g553_n,
    g552_p_spl_0,
    g550_p_spl_
  );


  and

  (
    g554_p,
    g552_n_spl_0,
    g551_n_spl_
  );


  or

  (
    g554_n,
    g552_p_spl_0,
    g551_p_spl_
  );


  and

  (
    g555_p,
    g554_n,
    g553_n
  );


  or

  (
    g555_n,
    g554_p,
    g553_p
  );


  and

  (
    g556_p,
    n2863_lo_p_spl_01,
    n2611_lo_p
  );


  or

  (
    g556_n,
    n2863_lo_n_spl_01,
    n2611_lo_n
  );


  and

  (
    g557_p,
    g556_n_spl_,
    g555_n_spl_
  );


  or

  (
    g557_n,
    g556_p_spl_,
    g555_p_spl_
  );


  and

  (
    g558_p,
    g557_n_spl_0,
    g555_n_spl_
  );


  or

  (
    g558_n,
    g557_p_spl_0,
    g555_p_spl_
  );


  and

  (
    g559_p,
    g557_n_spl_0,
    g556_n_spl_
  );


  or

  (
    g559_n,
    g557_p_spl_0,
    g556_p_spl_
  );


  and

  (
    g560_p,
    g559_n,
    g558_n
  );


  or

  (
    g560_n,
    g559_p,
    g558_p
  );


  and

  (
    g561_p,
    g531_n_spl_,
    g526_n_spl_
  );


  or

  (
    g561_n,
    g531_p_spl_,
    g526_p_spl_
  );


  and

  (
    g562_p,
    g561_n_spl_,
    g560_n_spl_
  );


  or

  (
    g562_n,
    g561_p_spl_,
    g560_p_spl_
  );


  and

  (
    g563_p,
    g562_n_spl_0,
    g560_n_spl_
  );


  or

  (
    g563_n,
    g562_p_spl_0,
    g560_p_spl_
  );


  and

  (
    g564_p,
    g562_n_spl_0,
    g561_n_spl_
  );


  or

  (
    g564_n,
    g562_p_spl_0,
    g561_p_spl_
  );


  and

  (
    g565_p,
    g564_n,
    g563_n
  );


  or

  (
    g565_n,
    g564_p,
    g563_p
  );


  and

  (
    g566_p,
    g541_n,
    g536_n_spl_
  );


  or

  (
    g566_n,
    g541_p_spl_,
    g536_p_spl_
  );


  and

  (
    g567_p,
    g566_n,
    g565_n
  );


  or

  (
    g567_n,
    g566_p_spl_,
    g565_p_spl_
  );


  or

  (
    g568_n,
    g567_p_spl_0,
    g565_p_spl_
  );


  or

  (
    g569_n,
    g567_p_spl_0,
    g566_p_spl_
  );


  and

  (
    g570_p,
    g569_n,
    g568_n
  );


  and

  (
    g571_p,
    G5044_o2_n_spl_,
    G5041_o2_n_spl_
  );


  or

  (
    g571_n,
    G5044_o2_p_spl_,
    G5041_o2_p_spl_
  );


  and

  (
    g572_p,
    g571_n_spl_0,
    G5044_o2_n_spl_
  );


  or

  (
    g572_n,
    g571_p_spl_0,
    G5044_o2_p_spl_
  );


  and

  (
    g573_p,
    g571_n_spl_0,
    G5041_o2_n_spl_
  );


  or

  (
    g573_n,
    g571_p_spl_0,
    G5041_o2_p_spl_
  );


  and

  (
    g574_p,
    g573_n,
    g572_n
  );


  or

  (
    g574_n,
    g573_p,
    g572_p
  );


  and

  (
    g575_p,
    n2851_lo_p_spl_00,
    n2635_lo_p_spl_
  );


  or

  (
    g575_n,
    n2851_lo_n_spl_00,
    n2635_lo_n_spl_
  );


  and

  (
    g576_p,
    g575_n_spl_,
    g574_n_spl_
  );


  or

  (
    g576_n,
    g575_p_spl_,
    g574_p_spl_
  );


  and

  (
    g577_p,
    g576_n_spl_0,
    g574_n_spl_
  );


  or

  (
    g577_n,
    g576_p_spl_0,
    g574_p_spl_
  );


  and

  (
    g578_p,
    g576_n_spl_0,
    g575_n_spl_
  );


  or

  (
    g578_n,
    g576_p_spl_0,
    g575_p_spl_
  );


  and

  (
    g579_p,
    g578_n,
    g577_n
  );


  or

  (
    g579_n,
    g578_p,
    g577_p
  );


  and

  (
    g580_p,
    g547_n_spl_,
    G5151_o2_p
  );


  or

  (
    g580_n,
    g547_p_spl_,
    G5151_o2_n
  );


  and

  (
    g581_p,
    g580_n_spl_,
    g579_n_spl_
  );


  or

  (
    g581_n,
    g580_p_spl_,
    g579_p_spl_
  );


  and

  (
    g582_p,
    g581_n_spl_0,
    g579_n_spl_
  );


  or

  (
    g582_n,
    g581_p_spl_0,
    g579_p_spl_
  );


  and

  (
    g583_p,
    g581_n_spl_0,
    g580_n_spl_
  );


  or

  (
    g583_n,
    g581_p_spl_0,
    g580_p_spl_
  );


  and

  (
    g584_p,
    g583_n,
    g582_n
  );


  or

  (
    g584_n,
    g583_p,
    g582_p
  );


  and

  (
    g585_p,
    n2863_lo_p_spl_01,
    n2623_lo_p_spl_
  );


  or

  (
    g585_n,
    n2863_lo_n_spl_01,
    n2623_lo_n_spl_
  );


  and

  (
    g586_p,
    g585_n_spl_,
    g584_n_spl_
  );


  or

  (
    g586_n,
    g585_p_spl_,
    g584_p_spl_
  );


  and

  (
    g587_p,
    g586_n_spl_0,
    g584_n_spl_
  );


  or

  (
    g587_n,
    g586_p_spl_0,
    g584_p_spl_
  );


  and

  (
    g588_p,
    g586_n_spl_0,
    g585_n_spl_
  );


  or

  (
    g588_n,
    g586_p_spl_0,
    g585_p_spl_
  );


  and

  (
    g589_p,
    g588_n,
    g587_n
  );


  or

  (
    g589_n,
    g588_p,
    g587_p
  );


  and

  (
    g590_p,
    g557_n_spl_,
    g552_n_spl_
  );


  or

  (
    g590_n,
    g557_p_spl_,
    g552_p_spl_
  );


  and

  (
    g591_p,
    g590_n_spl_,
    g589_n_spl_
  );


  or

  (
    g591_n,
    g590_p_spl_,
    g589_p_spl_
  );


  and

  (
    g592_p,
    g591_n_spl_0,
    g589_n_spl_
  );


  or

  (
    g592_n,
    g591_p_spl_0,
    g589_p_spl_
  );


  and

  (
    g593_p,
    g591_n_spl_0,
    g590_n_spl_
  );


  or

  (
    g593_n,
    g591_p_spl_0,
    g590_p_spl_
  );


  and

  (
    g594_p,
    g593_n,
    g592_n
  );


  or

  (
    g594_n,
    g593_p,
    g592_p
  );


  and

  (
    g595_p,
    g567_n,
    g562_n_spl_
  );


  or

  (
    g595_n,
    g567_p_spl_,
    g562_p_spl_
  );


  and

  (
    g596_p,
    g595_n,
    g594_n
  );


  or

  (
    g596_n,
    g595_p_spl_,
    g594_p_spl_
  );


  or

  (
    g597_n,
    g596_p_spl_0,
    g594_p_spl_
  );


  or

  (
    g598_n,
    g596_p_spl_0,
    g595_p_spl_
  );


  and

  (
    g599_p,
    g598_n,
    g597_n
  );


  and

  (
    g600_p,
    G4864_o2_n_spl_0,
    G4803_o2_p
  );


  or

  (
    g600_n,
    G4864_o2_p_spl_0,
    G4803_o2_n
  );


  and

  (
    g601_p,
    G4864_o2_n_spl_0,
    G1253_o2_n
  );


  or

  (
    g601_n,
    G4864_o2_p_spl_0,
    G1253_o2_p
  );


  and

  (
    g602_p,
    g601_n,
    g600_n
  );


  or

  (
    g602_n,
    g601_p,
    g600_p
  );


  and

  (
    g603_p,
    G4926_o2_n,
    G4743_o2_p
  );


  or

  (
    g603_n,
    G4926_o2_p,
    G4743_o2_n
  );


  and

  (
    g604_p,
    g603_n_spl_,
    g602_n_spl_
  );


  or

  (
    g604_n,
    g603_p_spl_,
    g602_p_spl_
  );


  and

  (
    g605_p,
    g604_n_spl_0,
    g602_n_spl_
  );


  or

  (
    g605_n,
    g604_p_spl_0,
    g602_p_spl_
  );


  and

  (
    g606_p,
    g604_n_spl_0,
    g603_n_spl_
  );


  or

  (
    g606_n,
    g604_p_spl_0,
    g603_p_spl_
  );


  and

  (
    g607_p,
    g606_n,
    g605_n
  );


  or

  (
    g607_n,
    g606_p,
    g605_p
  );


  and

  (
    g608_p,
    n2851_lo_p_spl_0,
    n2647_lo_p_spl_
  );


  or

  (
    g608_n,
    n2851_lo_n_spl_0,
    n2647_lo_n_spl_
  );


  and

  (
    g609_p,
    g608_n_spl_,
    g607_n_spl_
  );


  or

  (
    g609_n,
    g608_p_spl_,
    g607_p_spl_
  );


  and

  (
    g610_p,
    g609_n_spl_0,
    g607_n_spl_
  );


  or

  (
    g610_n,
    g609_p_spl_0,
    g607_p_spl_
  );


  and

  (
    g611_p,
    g609_n_spl_0,
    g608_n_spl_
  );


  or

  (
    g611_n,
    g609_p_spl_0,
    g608_p_spl_
  );


  and

  (
    g612_p,
    g611_n,
    g610_n
  );


  or

  (
    g612_n,
    g611_p,
    g610_p
  );


  and

  (
    g613_p,
    g576_n_spl_,
    g571_n_spl_
  );


  or

  (
    g613_n,
    g576_p_spl_,
    g571_p_spl_
  );


  and

  (
    g614_p,
    g613_n_spl_,
    g612_n_spl_
  );


  or

  (
    g614_n,
    g613_p_spl_,
    g612_p_spl_
  );


  and

  (
    g615_p,
    g614_n_spl_0,
    g612_n_spl_
  );


  or

  (
    g615_n,
    g614_p_spl_0,
    g612_p_spl_
  );


  and

  (
    g616_p,
    g614_n_spl_0,
    g613_n_spl_
  );


  or

  (
    g616_n,
    g614_p_spl_0,
    g613_p_spl_
  );


  and

  (
    g617_p,
    g616_n,
    g615_n
  );


  or

  (
    g617_n,
    g616_p,
    g615_p
  );


  and

  (
    g618_p,
    n2863_lo_p_spl_10,
    n2635_lo_p_spl_
  );


  or

  (
    g618_n,
    n2863_lo_n_spl_10,
    n2635_lo_n_spl_
  );


  and

  (
    g619_p,
    g618_n_spl_,
    g617_n_spl_
  );


  or

  (
    g619_n,
    g618_p_spl_,
    g617_p_spl_
  );


  and

  (
    g620_p,
    g619_n_spl_0,
    g617_n_spl_
  );


  or

  (
    g620_n,
    g619_p_spl_0,
    g617_p_spl_
  );


  and

  (
    g621_p,
    g619_n_spl_0,
    g618_n_spl_
  );


  or

  (
    g621_n,
    g619_p_spl_0,
    g618_p_spl_
  );


  and

  (
    g622_p,
    g621_n,
    g620_n
  );


  or

  (
    g622_n,
    g621_p,
    g620_p
  );


  and

  (
    g623_p,
    g586_n_spl_,
    g581_n_spl_
  );


  or

  (
    g623_n,
    g586_p_spl_,
    g581_p_spl_
  );


  and

  (
    g624_p,
    g623_n_spl_,
    g622_n_spl_
  );


  or

  (
    g624_n,
    g623_p_spl_,
    g622_p_spl_
  );


  and

  (
    g625_p,
    g624_n_spl_0,
    g622_n_spl_
  );


  or

  (
    g625_n,
    g624_p_spl_0,
    g622_p_spl_
  );


  and

  (
    g626_p,
    g624_n_spl_0,
    g623_n_spl_
  );


  or

  (
    g626_n,
    g624_p_spl_0,
    g623_p_spl_
  );


  and

  (
    g627_p,
    g626_n,
    g625_n
  );


  or

  (
    g627_n,
    g626_p,
    g625_p
  );


  and

  (
    g628_p,
    g596_n,
    g591_n_spl_
  );


  or

  (
    g628_n,
    g596_p_spl_,
    g591_p_spl_
  );


  and

  (
    g629_p,
    g628_n,
    g627_n
  );


  or

  (
    g629_n,
    g628_p_spl_,
    g627_p_spl_
  );


  or

  (
    g630_n,
    g629_p_spl_0,
    g627_p_spl_
  );


  or

  (
    g631_n,
    g629_p_spl_0,
    g628_p_spl_
  );


  and

  (
    g632_p,
    g631_n,
    g630_n
  );


  and

  (
    g633_p,
    n2839_lo_p,
    n2671_lo_p_spl_0
  );


  or

  (
    g633_n,
    n2839_lo_n,
    n2671_lo_n_spl_0
  );


  and

  (
    g634_p,
    G4864_o2_n_spl_,
    G4693_o2_p
  );


  or

  (
    g634_n,
    G4864_o2_p_spl_,
    G4693_o2_n
  );


  and

  (
    g635_p,
    g634_n_spl_,
    g633_n_spl_
  );


  or

  (
    g635_n,
    g634_p_spl_,
    g633_p_spl_
  );


  and

  (
    g636_p,
    g635_n_spl_0,
    g633_n_spl_
  );


  or

  (
    g636_n,
    g635_p_spl_0,
    g633_p_spl_
  );


  and

  (
    g637_p,
    g635_n_spl_0,
    g634_n_spl_
  );


  or

  (
    g637_n,
    g635_p_spl_0,
    g634_p_spl_
  );


  and

  (
    g638_p,
    g637_n,
    g636_n
  );


  or

  (
    g638_n,
    g637_p,
    g636_p
  );


  and

  (
    g639_p,
    n2851_lo_p_spl_1,
    n2659_lo_p_spl_
  );


  or

  (
    g639_n,
    n2851_lo_n_spl_1,
    n2659_lo_n_spl_
  );


  and

  (
    g640_p,
    g639_n_spl_,
    g638_n_spl_
  );


  or

  (
    g640_n,
    g639_p_spl_,
    g638_p_spl_
  );


  and

  (
    g641_p,
    g640_n_spl_0,
    g638_n_spl_
  );


  or

  (
    g641_n,
    g640_p_spl_0,
    g638_p_spl_
  );


  and

  (
    g642_p,
    g640_n_spl_0,
    g639_n_spl_
  );


  or

  (
    g642_n,
    g640_p_spl_0,
    g639_p_spl_
  );


  and

  (
    g643_p,
    g642_n,
    g641_n
  );


  or

  (
    g643_n,
    g642_p,
    g641_p
  );


  and

  (
    g644_p,
    g609_n_spl_,
    g604_n_spl_
  );


  or

  (
    g644_n,
    g609_p_spl_,
    g604_p_spl_
  );


  and

  (
    g645_p,
    g644_n_spl_,
    g643_n_spl_
  );


  or

  (
    g645_n,
    g644_p_spl_,
    g643_p_spl_
  );


  and

  (
    g646_p,
    g645_n_spl_0,
    g643_n_spl_
  );


  or

  (
    g646_n,
    g645_p_spl_0,
    g643_p_spl_
  );


  and

  (
    g647_p,
    g645_n_spl_0,
    g644_n_spl_
  );


  or

  (
    g647_n,
    g645_p_spl_0,
    g644_p_spl_
  );


  and

  (
    g648_p,
    g647_n,
    g646_n
  );


  or

  (
    g648_n,
    g647_p,
    g646_p
  );


  and

  (
    g649_p,
    n2863_lo_p_spl_10,
    n2647_lo_p_spl_
  );


  or

  (
    g649_n,
    n2863_lo_n_spl_10,
    n2647_lo_n_spl_
  );


  and

  (
    g650_p,
    g649_n_spl_,
    g648_n_spl_
  );


  or

  (
    g650_n,
    g649_p_spl_,
    g648_p_spl_
  );


  and

  (
    g651_p,
    g650_n_spl_0,
    g648_n_spl_
  );


  or

  (
    g651_n,
    g650_p_spl_0,
    g648_p_spl_
  );


  and

  (
    g652_p,
    g650_n_spl_0,
    g649_n_spl_
  );


  or

  (
    g652_n,
    g650_p_spl_0,
    g649_p_spl_
  );


  and

  (
    g653_p,
    g652_n,
    g651_n
  );


  or

  (
    g653_n,
    g652_p,
    g651_p
  );


  and

  (
    g654_p,
    g619_n_spl_,
    g614_n_spl_
  );


  or

  (
    g654_n,
    g619_p_spl_,
    g614_p_spl_
  );


  and

  (
    g655_p,
    g654_n_spl_,
    g653_n_spl_
  );


  or

  (
    g655_n,
    g654_p_spl_,
    g653_p_spl_
  );


  and

  (
    g656_p,
    g655_n_spl_0,
    g653_n_spl_
  );


  or

  (
    g656_n,
    g655_p_spl_0,
    g653_p_spl_
  );


  and

  (
    g657_p,
    g655_n_spl_0,
    g654_n_spl_
  );


  or

  (
    g657_n,
    g655_p_spl_0,
    g654_p_spl_
  );


  and

  (
    g658_p,
    g657_n,
    g656_n
  );


  or

  (
    g658_n,
    g657_p,
    g656_p
  );


  and

  (
    g659_p,
    g629_n,
    g624_n_spl_
  );


  or

  (
    g659_n,
    g629_p_spl_,
    g624_p_spl_
  );


  and

  (
    g660_p,
    g659_n,
    g658_n
  );


  or

  (
    g660_n,
    g659_p_spl_,
    g658_p_spl_
  );


  or

  (
    g661_n,
    g660_p_spl_0,
    g658_p_spl_
  );


  or

  (
    g662_n,
    g660_p_spl_0,
    g659_p_spl_
  );


  and

  (
    g663_p,
    g662_n,
    g661_n
  );


  and

  (
    g664_p,
    n2851_lo_p_spl_1,
    n2671_lo_p_spl_0
  );


  or

  (
    g664_n,
    n2851_lo_n_spl_1,
    n2671_lo_n_spl_0
  );


  and

  (
    g665_p,
    g640_n_spl_,
    g635_n_spl_
  );


  or

  (
    g665_n,
    g640_p_spl_,
    g635_p_spl_
  );


  and

  (
    g666_p,
    g665_n_spl_,
    g664_n_spl_
  );


  or

  (
    g666_n,
    g665_p_spl_,
    g664_p_spl_
  );


  and

  (
    g667_p,
    g666_n_spl_0,
    g664_n_spl_
  );


  or

  (
    g667_n,
    g666_p_spl_0,
    g664_p_spl_
  );


  and

  (
    g668_p,
    g666_n_spl_0,
    g665_n_spl_
  );


  or

  (
    g668_n,
    g666_p_spl_0,
    g665_p_spl_
  );


  and

  (
    g669_p,
    g668_n,
    g667_n
  );


  or

  (
    g669_n,
    g668_p,
    g667_p
  );


  and

  (
    g670_p,
    n2863_lo_p_spl_11,
    n2659_lo_p_spl_
  );


  or

  (
    g670_n,
    n2863_lo_n_spl_11,
    n2659_lo_n_spl_
  );


  and

  (
    g671_p,
    g670_n_spl_,
    g669_n_spl_
  );


  or

  (
    g671_n,
    g670_p_spl_,
    g669_p_spl_
  );


  and

  (
    g672_p,
    g671_n_spl_0,
    g669_n_spl_
  );


  or

  (
    g672_n,
    g671_p_spl_0,
    g669_p_spl_
  );


  and

  (
    g673_p,
    g671_n_spl_0,
    g670_n_spl_
  );


  or

  (
    g673_n,
    g671_p_spl_0,
    g670_p_spl_
  );


  and

  (
    g674_p,
    g673_n,
    g672_n
  );


  or

  (
    g674_n,
    g673_p,
    g672_p
  );


  and

  (
    g675_p,
    g650_n_spl_,
    g645_n_spl_
  );


  or

  (
    g675_n,
    g650_p_spl_,
    g645_p_spl_
  );


  and

  (
    g676_p,
    g675_n_spl_,
    g674_n_spl_
  );


  or

  (
    g676_n,
    g675_p_spl_,
    g674_p_spl_
  );


  and

  (
    g677_p,
    g676_n_spl_0,
    g674_n_spl_
  );


  or

  (
    g677_n,
    g676_p_spl_0,
    g674_p_spl_
  );


  and

  (
    g678_p,
    g676_n_spl_0,
    g675_n_spl_
  );


  or

  (
    g678_n,
    g676_p_spl_0,
    g675_p_spl_
  );


  and

  (
    g679_p,
    g678_n,
    g677_n
  );


  or

  (
    g679_n,
    g678_p,
    g677_p
  );


  and

  (
    g680_p,
    g660_n,
    g655_n_spl_
  );


  or

  (
    g680_n,
    g660_p_spl_,
    g655_p_spl_
  );


  and

  (
    g681_p,
    g680_n,
    g679_n
  );


  or

  (
    g681_n,
    g680_p_spl_,
    g679_p_spl_
  );


  or

  (
    g682_n,
    g681_p_spl_0,
    g679_p_spl_
  );


  or

  (
    g683_n,
    g681_p_spl_0,
    g680_p_spl_
  );


  and

  (
    g684_p,
    g683_n,
    g682_n
  );


  and

  (
    g685_p,
    n2863_lo_p_spl_11,
    n2671_lo_p_spl_
  );


  or

  (
    g685_n,
    n2863_lo_n_spl_11,
    n2671_lo_n_spl_
  );


  and

  (
    g686_p,
    g671_n_spl_,
    g666_n_spl_
  );


  or

  (
    g686_n,
    g671_p_spl_,
    g666_p_spl_
  );


  and

  (
    g687_p,
    g686_n_spl_,
    g685_n_spl_
  );


  or

  (
    g687_n,
    g686_p_spl_,
    g685_p_spl_
  );


  and

  (
    g688_p,
    g687_n_spl_0,
    g685_n_spl_
  );


  or

  (
    g688_n,
    g687_p_spl_,
    g685_p_spl_
  );


  and

  (
    g689_p,
    g687_n_spl_0,
    g686_n_spl_
  );


  or

  (
    g689_n,
    g687_p_spl_,
    g686_p_spl_
  );


  and

  (
    g690_p,
    g689_n,
    g688_n
  );


  or

  (
    g690_n,
    g689_p,
    g688_p
  );


  and

  (
    g691_p,
    g681_n,
    g676_n_spl_
  );


  or

  (
    g691_n,
    g681_p_spl_,
    g676_p_spl_
  );


  or

  (
    g692_n,
    g691_p,
    g690_p
  );


  and

  (
    g693_p,
    g692_n_spl_0,
    g687_n_spl_
  );


  and

  (
    g694_p,
    g692_n_spl_0,
    g690_n
  );


  and

  (
    g695_p,
    g692_n_spl_,
    g691_n
  );


  or

  (
    g696_n,
    g695_p,
    g694_p
  );


  and

  (
    g697_p,
    n2824_lo_buf_o2_p_spl_000,
    n6461_o2_p_spl_00
  );


  or

  (
    g697_n,
    n2824_lo_buf_o2_n_spl_000,
    n6461_o2_n_spl_0
  );


  and

  (
    g698_p,
    G5053_o2_n,
    G5054_o2_n
  );


  or

  (
    g698_n,
    G5053_o2_p,
    G5054_o2_p
  );


  and

  (
    g699_p,
    g698_n_spl_,
    g697_n
  );


  or

  (
    g699_n,
    g698_p,
    g697_p_spl_
  );


  and

  (
    g700_p,
    n6461_o2_p_spl_00,
    n2836_lo_p_spl_000
  );


  or

  (
    g700_n,
    n6461_o2_n_spl_0,
    n2836_lo_n_spl_000
  );


  and

  (
    g701_p,
    G5109_o2_p_spl_,
    G626_o2_n_spl_
  );


  or

  (
    g701_n,
    G5109_o2_n_spl_,
    G626_o2_p_spl_
  );


  and

  (
    g702_p,
    g701_n_spl_0,
    G5109_o2_p_spl_
  );


  or

  (
    g702_n,
    g701_p_spl_0,
    G5109_o2_n_spl_
  );


  and

  (
    g703_p,
    g701_n_spl_0,
    G626_o2_n_spl_
  );


  or

  (
    g703_n,
    g701_p_spl_0,
    G626_o2_p_spl_
  );


  and

  (
    g704_p,
    g703_n,
    g702_n
  );


  or

  (
    g704_n,
    g703_p,
    g702_p
  );


  and

  (
    g705_p,
    g699_n,
    G4993_o2_p
  );


  or

  (
    g705_n,
    g699_p_spl_,
    G4993_o2_n
  );


  and

  (
    g706_p,
    g705_n_spl_,
    g704_n_spl_
  );


  or

  (
    g706_n,
    g705_p_spl_,
    g704_p_spl_
  );


  and

  (
    g707_p,
    g706_n_spl_0,
    g704_n_spl_
  );


  or

  (
    g707_n,
    g706_p_spl_0,
    g704_p_spl_
  );


  and

  (
    g708_p,
    g706_n_spl_0,
    g705_n_spl_
  );


  or

  (
    g708_n,
    g706_p_spl_0,
    g705_p_spl_
  );


  and

  (
    g709_p,
    g708_n,
    g707_n
  );


  or

  (
    g709_n,
    g708_p,
    g707_p
  );


  and

  (
    g710_p,
    g709_n_spl_,
    g700_n
  );


  or

  (
    g710_n,
    g709_p,
    g700_p_spl_
  );


  and

  (
    g711_p,
    n6461_o2_p_spl_0,
    n2848_lo_p_spl_000
  );


  or

  (
    g711_n,
    n6461_o2_n_spl_1,
    n2848_lo_n_spl_000
  );


  and

  (
    g712_p,
    G5172_o2_n_spl_0,
    G5112_o2_p
  );


  or

  (
    g712_n,
    G5172_o2_p_spl_0,
    G5112_o2_n
  );


  and

  (
    g713_p,
    G5172_o2_n_spl_0,
    G674_o2_n
  );


  or

  (
    g713_n,
    G5172_o2_p_spl_0,
    G674_o2_p
  );


  and

  (
    g714_p,
    g713_n,
    g712_n
  );


  or

  (
    g714_n,
    g713_p,
    g712_p
  );


  and

  (
    g715_p,
    g701_n_spl_,
    G4997_o2_p
  );


  or

  (
    g715_n,
    g701_p_spl_,
    G4997_o2_n
  );


  and

  (
    g716_p,
    g715_n_spl_,
    g714_n_spl_
  );


  or

  (
    g716_n,
    g715_p_spl_,
    g714_p_spl_
  );


  and

  (
    g717_p,
    g716_n_spl_0,
    g714_n_spl_
  );


  or

  (
    g717_n,
    g716_p_spl_0,
    g714_p_spl_
  );


  and

  (
    g718_p,
    g716_n_spl_0,
    g715_n_spl_
  );


  or

  (
    g718_n,
    g716_p_spl_0,
    g715_p_spl_
  );


  and

  (
    g719_p,
    g718_n,
    g717_n
  );


  or

  (
    g719_n,
    g718_p,
    g717_p
  );


  and

  (
    g720_p,
    n6309_o2_p_spl_0,
    n2836_lo_p_spl_000
  );


  or

  (
    g720_n,
    n6309_o2_n_spl_0,
    n2836_lo_n_spl_000
  );


  and

  (
    g721_p,
    g720_n_spl_,
    g719_n_spl_
  );


  or

  (
    g721_n,
    g720_p_spl_,
    g719_p_spl_
  );


  and

  (
    g722_p,
    g721_n_spl_0,
    g719_n_spl_
  );


  or

  (
    g722_n,
    g721_p_spl_0,
    g719_p_spl_
  );


  and

  (
    g723_p,
    g721_n_spl_0,
    g720_n_spl_
  );


  or

  (
    g723_n,
    g721_p_spl_0,
    g720_p_spl_
  );


  and

  (
    g724_p,
    g723_n,
    g722_n
  );


  or

  (
    g724_n,
    g723_p,
    g722_p
  );


  and

  (
    g725_p,
    g710_n,
    g706_n_spl_
  );


  or

  (
    g725_n,
    g710_p_spl_,
    g706_p_spl_
  );


  and

  (
    g726_p,
    g725_n_spl_,
    g724_n_spl_
  );


  or

  (
    g726_n,
    g725_p_spl_,
    g724_p_spl_
  );


  and

  (
    g727_p,
    g726_n_spl_0,
    g724_n_spl_
  );


  or

  (
    g727_n,
    g726_p_spl_0,
    g724_p_spl_
  );


  and

  (
    g728_p,
    g726_n_spl_0,
    g725_n_spl_
  );


  or

  (
    g728_n,
    g726_p_spl_0,
    g725_p_spl_
  );


  and

  (
    g729_p,
    g728_n,
    g727_n
  );


  or

  (
    g729_n,
    g728_p,
    g727_p
  );


  and

  (
    g730_p,
    g729_n_spl_,
    g711_n
  );


  or

  (
    g730_n,
    g729_p,
    g711_p_spl_
  );


  and

  (
    g731_p,
    n2764_lo_buf_o2_p_spl_00,
    n8086_o2_p_spl_00
  );


  or

  (
    g731_n,
    n2764_lo_buf_o2_n_spl_00,
    n8086_o2_n_spl_00
  );


  and

  (
    g732_p,
    G3257_o2_p_spl_0,
    G3205_o2_n
  );


  or

  (
    g732_n,
    G3257_o2_n_spl_0,
    G3205_o2_p
  );


  and

  (
    g733_p,
    G3257_o2_p_spl_0,
    G3136_o2_n
  );


  or

  (
    g733_n,
    G3257_o2_n_spl_0,
    G3136_o2_p
  );


  and

  (
    g734_p,
    g733_n,
    g732_n
  );


  or

  (
    g734_n,
    g733_p,
    g732_p
  );


  and

  (
    g735_p,
    g734_n_spl_,
    g731_n
  );


  or

  (
    g735_n,
    g734_p,
    g731_p_spl_
  );


  and

  (
    g736_p,
    n6461_o2_p_spl_1,
    n2860_lo_p_spl_00
  );


  or

  (
    g736_n,
    n6461_o2_n_spl_1,
    n2860_lo_n_spl_00
  );


  and

  (
    g737_p,
    G5242_o2_n,
    G5243_o2_p
  );


  or

  (
    g737_n,
    G5242_o2_p,
    G5243_o2_n
  );


  and

  (
    g738_p,
    G5172_o2_n_spl_,
    G5001_o2_p
  );


  or

  (
    g738_n,
    G5172_o2_p_spl_,
    G5001_o2_n
  );


  and

  (
    g739_p,
    g738_n_spl_,
    g737_n_spl_
  );


  or

  (
    g739_n,
    g738_p_spl_,
    g737_p_spl_
  );


  and

  (
    g740_p,
    g739_n_spl_0,
    g737_n_spl_
  );


  or

  (
    g740_n,
    g739_p_spl_0,
    g737_p_spl_
  );


  and

  (
    g741_p,
    g739_n_spl_0,
    g738_n_spl_
  );


  or

  (
    g741_n,
    g739_p_spl_0,
    g738_p_spl_
  );


  and

  (
    g742_p,
    g741_n,
    g740_n
  );


  or

  (
    g742_n,
    g741_p,
    g740_p
  );


  and

  (
    g743_p,
    n6239_o2_p_spl_0,
    n2836_lo_p_spl_001
  );


  or

  (
    g743_n,
    n6239_o2_n_spl_0,
    n2836_lo_n_spl_001
  );


  and

  (
    g744_p,
    g743_n_spl_,
    g742_n_spl_
  );


  or

  (
    g744_n,
    g743_p_spl_,
    g742_p_spl_
  );


  and

  (
    g745_p,
    g744_n_spl_0,
    g742_n_spl_
  );


  or

  (
    g745_n,
    g744_p_spl_0,
    g742_p_spl_
  );


  and

  (
    g746_p,
    g744_n_spl_0,
    g743_n_spl_
  );


  or

  (
    g746_n,
    g744_p_spl_0,
    g743_p_spl_
  );


  and

  (
    g747_p,
    g746_n,
    g745_n
  );


  or

  (
    g747_n,
    g746_p,
    g745_p
  );


  and

  (
    g748_p,
    g721_n_spl_,
    g716_n_spl_
  );


  or

  (
    g748_n,
    g721_p_spl_,
    g716_p_spl_
  );


  and

  (
    g749_p,
    g748_n_spl_,
    g747_n_spl_
  );


  or

  (
    g749_n,
    g748_p_spl_,
    g747_p_spl_
  );


  and

  (
    g750_p,
    g749_n_spl_0,
    g747_n_spl_
  );


  or

  (
    g750_n,
    g749_p_spl_0,
    g747_p_spl_
  );


  and

  (
    g751_p,
    g749_n_spl_0,
    g748_n_spl_
  );


  or

  (
    g751_n,
    g749_p_spl_0,
    g748_p_spl_
  );


  and

  (
    g752_p,
    g751_n,
    g750_n
  );


  or

  (
    g752_n,
    g751_p,
    g750_p
  );


  and

  (
    g753_p,
    n6309_o2_p_spl_0,
    n2848_lo_p_spl_000
  );


  or

  (
    g753_n,
    n6309_o2_n_spl_0,
    n2848_lo_n_spl_000
  );


  and

  (
    g754_p,
    g753_n_spl_,
    g752_n_spl_
  );


  or

  (
    g754_n,
    g753_p_spl_,
    g752_p_spl_
  );


  and

  (
    g755_p,
    g754_n_spl_0,
    g752_n_spl_
  );


  or

  (
    g755_n,
    g754_p_spl_0,
    g752_p_spl_
  );


  and

  (
    g756_p,
    g754_n_spl_0,
    g753_n_spl_
  );


  or

  (
    g756_n,
    g754_p_spl_0,
    g753_p_spl_
  );


  and

  (
    g757_p,
    g756_n,
    g755_n
  );


  or

  (
    g757_n,
    g756_p,
    g755_p
  );


  and

  (
    g758_p,
    g730_n,
    g726_n_spl_
  );


  or

  (
    g758_n,
    g730_p_spl_,
    g726_p_spl_
  );


  and

  (
    g759_p,
    g758_n_spl_,
    g757_n_spl_
  );


  or

  (
    g759_n,
    g758_p_spl_,
    g757_p_spl_
  );


  and

  (
    g760_p,
    g759_n_spl_0,
    g757_n_spl_
  );


  or

  (
    g760_n,
    g759_p_spl_0,
    g757_p_spl_
  );


  and

  (
    g761_p,
    g759_n_spl_0,
    g758_n_spl_
  );


  or

  (
    g761_n,
    g759_p_spl_0,
    g758_p_spl_
  );


  and

  (
    g762_p,
    g761_n,
    g760_n
  );


  or

  (
    g762_n,
    g761_p,
    g760_p
  );


  and

  (
    g763_p,
    n2776_lo_buf_o2_p_spl_000,
    n8086_o2_p_spl_00
  );


  or

  (
    g763_n,
    n2776_lo_buf_o2_n_spl_000,
    n8086_o2_n_spl_00
  );


  and

  (
    g764_p,
    g762_n_spl_,
    g736_n
  );


  or

  (
    g764_n,
    g762_p,
    g736_p_spl_
  );


  and

  (
    g765_p,
    G3318_o2_n,
    G3319_o2_n
  );


  or

  (
    g765_n,
    G3318_o2_p,
    G3319_o2_p
  );


  and

  (
    g766_p,
    n2764_lo_buf_o2_p_spl_00,
    n7909_o2_p_spl_00
  );


  or

  (
    g766_n,
    n2764_lo_buf_o2_n_spl_00,
    n7909_o2_n_spl_00
  );


  and

  (
    g767_p,
    g766_n_spl_,
    g765_n_spl_
  );


  or

  (
    g767_n,
    g766_p_spl_,
    g765_p_spl_
  );


  and

  (
    g768_p,
    g767_n_spl_0,
    g765_n_spl_
  );


  or

  (
    g768_n,
    g767_p_spl_0,
    g765_p_spl_
  );


  and

  (
    g769_p,
    g767_n_spl_0,
    g766_n_spl_
  );


  or

  (
    g769_n,
    g767_p_spl_0,
    g766_p_spl_
  );


  and

  (
    g770_p,
    g769_n,
    g768_n
  );


  or

  (
    g770_n,
    g769_p,
    g768_p
  );


  and

  (
    g771_p,
    g735_n,
    G3257_o2_p_spl_
  );


  or

  (
    g771_n,
    g735_p_spl_,
    G3257_o2_n_spl_
  );


  and

  (
    g772_p,
    g771_n_spl_,
    g770_n_spl_
  );


  or

  (
    g772_n,
    g771_p_spl_,
    g770_p_spl_
  );


  and

  (
    g773_p,
    g772_n_spl_0,
    g770_n_spl_
  );


  or

  (
    g773_n,
    g772_p_spl_0,
    g770_p_spl_
  );


  and

  (
    g774_p,
    g772_n_spl_0,
    g771_n_spl_
  );


  or

  (
    g774_n,
    g772_p_spl_0,
    g771_p_spl_
  );


  and

  (
    g775_p,
    g774_n,
    g773_n
  );


  or

  (
    g775_n,
    g774_p,
    g773_p
  );


  and

  (
    g776_p,
    g775_n_spl_,
    g763_n
  );


  or

  (
    g776_n,
    g775_p,
    g763_p_spl_
  );


  and

  (
    g777_p,
    n2488_lo_buf_o2_p_spl_00,
    n2704_lo_buf_o2_p_spl_0
  );


  or

  (
    g777_n,
    n2488_lo_buf_o2_n_spl_00,
    n2704_lo_buf_o2_n_spl_0
  );


  and

  (
    g778_p,
    G1580_o2_n_spl_,
    G1507_o2_n_spl_
  );


  or

  (
    g778_n,
    G1580_o2_p_spl_,
    G1507_o2_p_spl_
  );


  and

  (
    g779_p,
    g778_n_spl_0,
    G1580_o2_n_spl_
  );


  or

  (
    g779_n,
    g778_p_spl_0,
    G1580_o2_p_spl_
  );


  and

  (
    g780_p,
    g778_n_spl_0,
    G1507_o2_n_spl_
  );


  or

  (
    g780_n,
    g778_p_spl_0,
    G1507_o2_p_spl_
  );


  and

  (
    g781_p,
    g780_n,
    g779_n
  );


  or

  (
    g781_n,
    g780_p,
    g779_p
  );


  and

  (
    g782_p,
    n8086_o2_p_spl_01,
    n2785_lo_p_spl_000
  );


  or

  (
    g782_n,
    n8086_o2_n_spl_0,
    n2785_lo_n_spl_000
  );


  and

  (
    g783_p,
    g781_n_spl_,
    g777_n
  );


  or

  (
    g783_n,
    g781_p,
    g777_p_spl_
  );


  and

  (
    g784_p,
    G3364_o2_p_spl_,
    G659_o2_n_spl_
  );


  or

  (
    g784_n,
    G3364_o2_n_spl_,
    G659_o2_p_spl_
  );


  and

  (
    g785_p,
    g784_n_spl_0,
    G3364_o2_p_spl_
  );


  or

  (
    g785_n,
    g784_p_spl_0,
    G3364_o2_n_spl_
  );


  and

  (
    g786_p,
    g784_n_spl_0,
    G659_o2_n_spl_
  );


  or

  (
    g786_n,
    g784_p_spl_0,
    G659_o2_p_spl_
  );


  and

  (
    g787_p,
    g786_n,
    g785_n
  );


  or

  (
    g787_n,
    g786_p,
    g785_p
  );


  and

  (
    g788_p,
    g767_n_spl_,
    G3261_o2_p
  );


  or

  (
    g788_n,
    g767_p_spl_,
    G3261_o2_n
  );


  and

  (
    g789_p,
    g788_n_spl_,
    g787_n_spl_
  );


  or

  (
    g789_n,
    g788_p_spl_,
    g787_p_spl_
  );


  and

  (
    g790_p,
    g789_n_spl_0,
    g787_n_spl_
  );


  or

  (
    g790_n,
    g789_p_spl_0,
    g787_p_spl_
  );


  and

  (
    g791_p,
    g789_n_spl_0,
    g788_n_spl_
  );


  or

  (
    g791_n,
    g789_p_spl_0,
    g788_p_spl_
  );


  and

  (
    g792_p,
    g791_n,
    g790_n
  );


  or

  (
    g792_n,
    g791_p,
    g790_p
  );


  and

  (
    g793_p,
    n2776_lo_buf_o2_p_spl_000,
    n7909_o2_p_spl_00
  );


  or

  (
    g793_n,
    n2776_lo_buf_o2_n_spl_000,
    n7909_o2_n_spl_00
  );


  and

  (
    g794_p,
    g793_n_spl_,
    g792_n_spl_
  );


  or

  (
    g794_n,
    g793_p_spl_,
    g792_p_spl_
  );


  and

  (
    g795_p,
    g794_n_spl_0,
    g792_n_spl_
  );


  or

  (
    g795_n,
    g794_p_spl_0,
    g792_p_spl_
  );


  and

  (
    g796_p,
    g794_n_spl_0,
    g793_n_spl_
  );


  or

  (
    g796_n,
    g794_p_spl_0,
    g793_p_spl_
  );


  and

  (
    g797_p,
    g796_n,
    g795_n
  );


  or

  (
    g797_n,
    g796_p,
    g795_p
  );


  and

  (
    g798_p,
    g776_n,
    g772_n_spl_
  );


  or

  (
    g798_n,
    g776_p_spl_,
    g772_p_spl_
  );


  and

  (
    g799_p,
    g798_n_spl_,
    g797_n_spl_
  );


  or

  (
    g799_n,
    g798_p_spl_,
    g797_p_spl_
  );


  and

  (
    g800_p,
    g799_n_spl_0,
    g797_n_spl_
  );


  or

  (
    g800_n,
    g799_p_spl_0,
    g797_p_spl_
  );


  and

  (
    g801_p,
    g799_n_spl_0,
    g798_n_spl_
  );


  or

  (
    g801_n,
    g799_p_spl_0,
    g798_p_spl_
  );


  and

  (
    g802_p,
    g801_n,
    g800_n
  );


  or

  (
    g802_n,
    g801_p,
    g800_p
  );


  and

  (
    g803_p,
    g802_n_spl_,
    g782_n
  );


  or

  (
    g803_n,
    g802_p,
    g782_p_spl_
  );


  and

  (
    g804_p,
    n2488_lo_buf_o2_p_spl_00,
    n2716_lo_buf_o2_p_spl_000
  );


  or

  (
    g804_n,
    n2488_lo_buf_o2_n_spl_00,
    n2716_lo_buf_o2_n_spl_000
  );


  and

  (
    g805_p,
    G1630_o2_p_spl_0,
    G1583_o2_n
  );


  or

  (
    g805_n,
    G1630_o2_n_spl_0,
    G1583_o2_p
  );


  and

  (
    g806_p,
    G1630_o2_p_spl_0,
    G1512_o2_n
  );


  or

  (
    g806_n,
    G1630_o2_n_spl_0,
    G1512_o2_p
  );


  and

  (
    g807_p,
    g806_n,
    g805_n
  );


  or

  (
    g807_n,
    g806_p,
    g805_p
  );


  and

  (
    g808_p,
    n2500_lo_buf_o2_p_spl_00,
    n2704_lo_buf_o2_p_spl_0
  );


  or

  (
    g808_n,
    n2500_lo_buf_o2_n_spl_00,
    n2704_lo_buf_o2_n_spl_0
  );


  and

  (
    g809_p,
    g808_n_spl_,
    g807_n_spl_
  );


  or

  (
    g809_n,
    g808_p_spl_,
    g807_p_spl_
  );


  and

  (
    g810_p,
    g809_n_spl_0,
    g807_n_spl_
  );


  or

  (
    g810_n,
    g809_p_spl_0,
    g807_p_spl_
  );


  and

  (
    g811_p,
    g809_n_spl_0,
    g808_n_spl_
  );


  or

  (
    g811_n,
    g809_p_spl_0,
    g808_p_spl_
  );


  and

  (
    g812_p,
    g811_n,
    g810_n
  );


  or

  (
    g812_n,
    g811_p,
    g810_p
  );


  and

  (
    g813_p,
    g783_n,
    g778_n_spl_
  );


  or

  (
    g813_n,
    g783_p_spl_,
    g778_p_spl_
  );


  and

  (
    g814_p,
    g813_n_spl_,
    g812_n_spl_
  );


  or

  (
    g814_n,
    g813_p_spl_,
    g812_p_spl_
  );


  and

  (
    g815_p,
    g814_n_spl_0,
    g812_n_spl_
  );


  or

  (
    g815_n,
    g814_p_spl_0,
    g812_p_spl_
  );


  and

  (
    g816_p,
    g814_n_spl_0,
    g813_n_spl_
  );


  or

  (
    g816_n,
    g814_p_spl_0,
    g813_p_spl_
  );


  and

  (
    g817_p,
    g816_n,
    g815_n
  );


  or

  (
    g817_n,
    g816_p,
    g815_p
  );


  and

  (
    g818_p,
    n2812_lo_buf_o2_p_spl_00,
    n5779_o2_p_spl_0
  );


  or

  (
    g818_n,
    n2812_lo_buf_o2_n_spl_00,
    n5779_o2_n_spl_0
  );


  and

  (
    g819_p,
    n2800_lo_buf_o2_p_spl_,
    n5779_o2_p_spl_0
  );


  or

  (
    g819_n,
    n2800_lo_buf_o2_n_spl_,
    n5779_o2_n_spl_0
  );


  and

  (
    g820_p,
    G3886_o2_n,
    G3885_o2_n
  );


  or

  (
    g820_n,
    G3886_o2_p,
    G3885_o2_p
  );


  and

  (
    g821_p,
    n2800_lo_buf_o2_p_spl_,
    n5792_o2_p_spl_0
  );


  or

  (
    g821_n,
    n2800_lo_buf_o2_n_spl_,
    n5792_o2_n_spl_0
  );


  and

  (
    g822_p,
    g821_n_spl_,
    g820_n_spl_
  );


  or

  (
    g822_n,
    g821_p_spl_,
    g820_p_spl_
  );


  and

  (
    g823_p,
    g822_n_spl_0,
    G3813_o2_p
  );


  or

  (
    g823_n,
    g822_p_spl_0,
    G3813_o2_n
  );


  and

  (
    g824_p,
    g823_n_spl_,
    g819_n_spl_
  );


  or

  (
    g824_n,
    g823_p_spl_,
    g819_p_spl_
  );


  and

  (
    g825_p,
    g824_n_spl_0,
    g819_n_spl_
  );


  or

  (
    g825_n,
    g824_p_spl_0,
    g819_p_spl_
  );


  and

  (
    g826_p,
    g824_n_spl_0,
    g823_n_spl_
  );


  or

  (
    g826_n,
    g824_p_spl_0,
    g823_p_spl_
  );


  and

  (
    g827_p,
    g826_n,
    g825_n
  );


  or

  (
    g827_n,
    g826_p,
    g825_p
  );


  and

  (
    g828_p,
    n2812_lo_buf_o2_p_spl_00,
    n5792_o2_p_spl_0
  );


  or

  (
    g828_n,
    n2812_lo_buf_o2_n_spl_00,
    n5792_o2_n_spl_0
  );


  and

  (
    g829_p,
    g828_n_spl_,
    g827_n_spl_
  );


  or

  (
    g829_n,
    g828_p_spl_,
    g827_p_spl_
  );


  and

  (
    g830_p,
    g829_n_spl_0,
    g824_n_spl_
  );


  or

  (
    g830_n,
    g829_p_spl_0,
    g824_p_spl_
  );


  and

  (
    g831_p,
    g830_n_spl_,
    g818_n_spl_
  );


  or

  (
    g831_n,
    g830_p_spl_,
    g818_p_spl_
  );


  and

  (
    g832_p,
    g831_n_spl_0,
    g818_n_spl_
  );


  or

  (
    g832_n,
    g831_p_spl_0,
    g818_p_spl_
  );


  and

  (
    g833_p,
    g831_n_spl_0,
    g830_n_spl_
  );


  or

  (
    g833_n,
    g831_p_spl_0,
    g830_p_spl_
  );


  and

  (
    g834_p,
    g833_n,
    g832_n
  );


  or

  (
    g834_n,
    g833_p,
    g832_p
  );


  and

  (
    g835_p,
    n2824_lo_buf_o2_p_spl_000,
    n5792_o2_p_spl_1
  );


  or

  (
    g835_n,
    n2824_lo_buf_o2_n_spl_000,
    n5792_o2_n_spl_1
  );


  and

  (
    g836_p,
    g835_n_spl_,
    g834_n_spl_
  );


  or

  (
    g836_n,
    g835_p_spl_,
    g834_p_spl_
  );


  and

  (
    g837_p,
    g836_n_spl_0,
    g834_n_spl_
  );


  or

  (
    g837_n,
    g836_p_spl_0,
    g834_p_spl_
  );


  and

  (
    g838_p,
    g836_n_spl_0,
    g835_n_spl_
  );


  or

  (
    g838_n,
    g836_p_spl_0,
    g835_p_spl_
  );


  and

  (
    g839_p,
    g838_n,
    g837_n
  );


  or

  (
    g839_n,
    g838_p,
    g837_p
  );


  and

  (
    g840_p,
    g829_n_spl_0,
    g827_n_spl_
  );


  or

  (
    g840_n,
    g829_p_spl_0,
    g827_p_spl_
  );


  and

  (
    g841_p,
    g829_n_spl_,
    g828_n_spl_
  );


  or

  (
    g841_n,
    g829_p_spl_,
    g828_p_spl_
  );


  and

  (
    g842_p,
    g841_n,
    g840_n
  );


  or

  (
    g842_n,
    g841_p,
    g840_p
  );


  and

  (
    g843_p,
    g822_n_spl_0,
    g820_n_spl_
  );


  or

  (
    g843_n,
    g822_p_spl_0,
    g820_p_spl_
  );


  and

  (
    g844_p,
    g822_n_spl_,
    g821_n_spl_
  );


  or

  (
    g844_n,
    g822_p_spl_,
    g821_p_spl_
  );


  and

  (
    g845_p,
    g844_n,
    g843_n
  );


  or

  (
    g845_n,
    g844_p,
    g843_p
  );


  and

  (
    g846_p,
    G4034_o2_n_spl_0,
    G3881_o2_p
  );


  or

  (
    g846_n,
    G4034_o2_p_spl_0,
    G3881_o2_n
  );


  and

  (
    g847_p,
    g846_n_spl_,
    g845_n_spl_
  );


  or

  (
    g847_n,
    g846_p_spl_,
    g845_p_spl_
  );


  and

  (
    g848_p,
    g847_n_spl_0,
    g845_n_spl_
  );


  or

  (
    g848_n,
    g847_p_spl_0,
    g845_p_spl_
  );


  and

  (
    g849_p,
    g847_n_spl_0,
    g846_n_spl_
  );


  or

  (
    g849_n,
    g847_p_spl_0,
    g846_p_spl_
  );


  and

  (
    g850_p,
    g849_n,
    g848_n
  );


  or

  (
    g850_n,
    g849_p,
    g848_p
  );


  and

  (
    g851_p,
    n2812_lo_buf_o2_p_spl_01,
    n5842_o2_p_spl_0
  );


  or

  (
    g851_n,
    n2812_lo_buf_o2_n_spl_01,
    n5842_o2_n_spl_0
  );


  and

  (
    g852_p,
    g851_n_spl_,
    g850_n_spl_
  );


  or

  (
    g852_n,
    g851_p_spl_,
    g850_p_spl_
  );


  and

  (
    g853_p,
    g852_n_spl_0,
    g847_n_spl_
  );


  or

  (
    g853_n,
    g852_p_spl_0,
    g847_p_spl_
  );


  and

  (
    g854_p,
    g853_n_spl_,
    g842_n_spl_
  );


  or

  (
    g854_n,
    g853_p_spl_,
    g842_p_spl_
  );


  and

  (
    g855_p,
    g854_n_spl_0,
    g842_n_spl_
  );


  or

  (
    g855_n,
    g854_p_spl_0,
    g842_p_spl_
  );


  and

  (
    g856_p,
    g854_n_spl_0,
    g853_n_spl_
  );


  or

  (
    g856_n,
    g854_p_spl_0,
    g853_p_spl_
  );


  and

  (
    g857_p,
    g856_n,
    g855_n
  );


  or

  (
    g857_n,
    g856_p,
    g855_p
  );


  and

  (
    g858_p,
    n2824_lo_buf_o2_p_spl_001,
    n5842_o2_p_spl_0
  );


  or

  (
    g858_n,
    n2824_lo_buf_o2_n_spl_001,
    n5842_o2_n_spl_0
  );


  and

  (
    g859_p,
    g858_n_spl_,
    g857_n_spl_
  );


  or

  (
    g859_n,
    g858_p_spl_,
    g857_p_spl_
  );


  and

  (
    g860_p,
    g859_n_spl_0,
    g854_n_spl_
  );


  or

  (
    g860_n,
    g859_p_spl_0,
    g854_p_spl_
  );


  and

  (
    g861_p,
    g860_n_spl_,
    g839_n_spl_
  );


  or

  (
    g861_n,
    g860_p_spl_,
    g839_p_spl_
  );


  and

  (
    g862_p,
    G4034_o2_n_spl_0,
    G3989_o2_p
  );


  or

  (
    g862_n,
    G4034_o2_p_spl_0,
    G3989_o2_n
  );


  and

  (
    g863_p,
    G4034_o2_n_spl_,
    G1196_o2_n
  );


  or

  (
    g863_n,
    G4034_o2_p_spl_,
    G1196_o2_p
  );


  and

  (
    g864_p,
    g863_n,
    g862_n
  );


  or

  (
    g864_n,
    g863_p,
    g862_p
  );


  and

  (
    g865_p,
    G4085_o2_n,
    G3929_o2_p
  );


  or

  (
    g865_n,
    G4085_o2_p,
    G3929_o2_n
  );


  and

  (
    g866_p,
    g865_n_spl_,
    g864_n_spl_
  );


  or

  (
    g866_n,
    g865_p_spl_,
    g864_p_spl_
  );


  and

  (
    g867_p,
    g866_n_spl_0,
    g864_n_spl_
  );


  or

  (
    g867_n,
    g866_p_spl_0,
    g864_p_spl_
  );


  and

  (
    g868_p,
    g866_n_spl_0,
    g865_n_spl_
  );


  or

  (
    g868_n,
    g866_p_spl_0,
    g865_p_spl_
  );


  and

  (
    g869_p,
    g868_n,
    g867_n
  );


  or

  (
    g869_n,
    g868_p,
    g867_p
  );


  and

  (
    g870_p,
    n2812_lo_buf_o2_p_spl_01,
    n5863_o2_p_spl_0
  );


  or

  (
    g870_n,
    n2812_lo_buf_o2_n_spl_01,
    n5863_o2_n_spl_0
  );


  and

  (
    g871_p,
    g870_n_spl_,
    g869_n_spl_
  );


  or

  (
    g871_n,
    g870_p_spl_,
    g869_p_spl_
  );


  and

  (
    g872_p,
    g871_n_spl_0,
    g869_n_spl_
  );


  or

  (
    g872_n,
    g871_p_spl_0,
    g869_p_spl_
  );


  and

  (
    g873_p,
    g871_n_spl_0,
    g870_n_spl_
  );


  or

  (
    g873_n,
    g871_p_spl_0,
    g870_p_spl_
  );


  and

  (
    g874_p,
    g873_n,
    g872_n
  );


  or

  (
    g874_n,
    g873_p,
    g872_p
  );


  and

  (
    g875_p,
    G4220_o2_n_spl_,
    G4217_o2_n_spl_
  );


  or

  (
    g875_n,
    G4220_o2_p_spl_,
    G4217_o2_p_spl_
  );


  and

  (
    g876_p,
    g875_n_spl_0,
    G4220_o2_n_spl_
  );


  or

  (
    g876_n,
    g875_p_spl_0,
    G4220_o2_p_spl_
  );


  and

  (
    g877_p,
    g875_n_spl_0,
    G4217_o2_n_spl_
  );


  or

  (
    g877_n,
    g875_p_spl_0,
    G4217_o2_p_spl_
  );


  and

  (
    g878_p,
    g877_n,
    g876_n
  );


  or

  (
    g878_n,
    g877_p,
    g876_p
  );


  and

  (
    g879_p,
    n2812_lo_buf_o2_p_spl_1,
    n5881_o2_p_spl_0
  );


  or

  (
    g879_n,
    n2812_lo_buf_o2_n_spl_1,
    n5881_o2_n_spl_0
  );


  and

  (
    g880_p,
    g879_n_spl_,
    g878_n_spl_
  );


  or

  (
    g880_n,
    g879_p_spl_,
    g878_p_spl_
  );


  and

  (
    g881_p,
    g880_n_spl_0,
    g875_n_spl_
  );


  or

  (
    g881_n,
    g880_p_spl_0,
    g875_p_spl_
  );


  and

  (
    g882_p,
    g881_n_spl_,
    g874_n_spl_
  );


  or

  (
    g882_n,
    g881_p_spl_,
    g874_p_spl_
  );


  and

  (
    g883_p,
    g882_n_spl_0,
    g874_n_spl_
  );


  or

  (
    g883_n,
    g882_p_spl_0,
    g874_p_spl_
  );


  and

  (
    g884_p,
    g882_n_spl_0,
    g881_n_spl_
  );


  or

  (
    g884_n,
    g882_p_spl_0,
    g881_p_spl_
  );


  and

  (
    g885_p,
    g884_n,
    g883_n
  );


  or

  (
    g885_n,
    g884_p,
    g883_p
  );


  and

  (
    g886_p,
    n2824_lo_buf_o2_p_spl_001,
    n5881_o2_p_spl_0
  );


  or

  (
    g886_n,
    n2824_lo_buf_o2_n_spl_001,
    n5881_o2_n_spl_0
  );


  and

  (
    g887_p,
    g886_n_spl_,
    g885_n_spl_
  );


  or

  (
    g887_n,
    g886_p_spl_,
    g885_p_spl_
  );


  and

  (
    g888_p,
    g887_n_spl_0,
    g885_n_spl_
  );


  or

  (
    g888_n,
    g887_p_spl_0,
    g885_p_spl_
  );


  and

  (
    g889_p,
    g887_n_spl_0,
    g886_n_spl_
  );


  or

  (
    g889_n,
    g887_p_spl_0,
    g886_p_spl_
  );


  and

  (
    g890_p,
    g889_n,
    g888_n
  );


  or

  (
    g890_n,
    g889_p,
    g888_p
  );


  and

  (
    g891_p,
    g880_n_spl_0,
    g878_n_spl_
  );


  or

  (
    g891_n,
    g880_p_spl_0,
    g878_p_spl_
  );


  and

  (
    g892_p,
    g880_n_spl_,
    g879_n_spl_
  );


  or

  (
    g892_n,
    g880_p_spl_,
    g879_p_spl_
  );


  and

  (
    g893_p,
    g892_n,
    g891_n
  );


  or

  (
    g893_n,
    g892_p,
    g891_p
  );


  and

  (
    g894_p,
    G4374_o2_n,
    G4375_o2_n
  );


  or

  (
    g894_n,
    G4374_o2_p,
    G4375_o2_p
  );


  and

  (
    g895_p,
    n2812_lo_buf_o2_p_spl_1,
    n5930_o2_p_spl_0
  );


  or

  (
    g895_n,
    n2812_lo_buf_o2_n_spl_1,
    n5930_o2_n_spl_0
  );


  and

  (
    g896_p,
    g895_n_spl_,
    g894_n_spl_
  );


  or

  (
    g896_n,
    g895_p_spl_,
    g894_p_spl_
  );


  and

  (
    g897_p,
    g896_n_spl_0,
    G4325_o2_p
  );


  or

  (
    g897_n,
    g896_p_spl_0,
    G4325_o2_n
  );


  and

  (
    g898_p,
    g897_n_spl_,
    g893_n_spl_
  );


  or

  (
    g898_n,
    g897_p_spl_,
    g893_p_spl_
  );


  and

  (
    g899_p,
    g898_n_spl_0,
    g893_n_spl_
  );


  or

  (
    g899_n,
    g898_p_spl_0,
    g893_p_spl_
  );


  and

  (
    g900_p,
    g898_n_spl_0,
    g897_n_spl_
  );


  or

  (
    g900_n,
    g898_p_spl_0,
    g897_p_spl_
  );


  and

  (
    g901_p,
    g900_n,
    g899_n
  );


  or

  (
    g901_n,
    g900_p,
    g899_p
  );


  and

  (
    g902_p,
    n2824_lo_buf_o2_p_spl_010,
    n5930_o2_p_spl_0
  );


  or

  (
    g902_n,
    n2824_lo_buf_o2_n_spl_010,
    n5930_o2_n_spl_0
  );


  and

  (
    g903_p,
    g902_n_spl_,
    g901_n_spl_
  );


  or

  (
    g903_n,
    g902_p_spl_,
    g901_p_spl_
  );


  and

  (
    g904_p,
    g903_n_spl_0,
    g898_n_spl_
  );


  or

  (
    g904_n,
    g903_p_spl_0,
    g898_p_spl_
  );


  and

  (
    g905_p,
    g904_n_spl_,
    g890_n_spl_
  );


  or

  (
    g905_n,
    g904_p_spl_,
    g890_p_spl_
  );


  and

  (
    g906_p,
    g905_n_spl_0,
    g890_n_spl_
  );


  or

  (
    g906_n,
    g905_p_spl_0,
    g890_p_spl_
  );


  and

  (
    g907_p,
    g905_n_spl_0,
    g904_n_spl_
  );


  or

  (
    g907_n,
    g905_p_spl_0,
    g904_p_spl_
  );


  and

  (
    g908_p,
    g907_n,
    g906_n
  );


  or

  (
    g908_n,
    g907_p,
    g906_p
  );


  and

  (
    g909_p,
    n5930_o2_p_spl_1,
    n2836_lo_p_spl_001
  );


  or

  (
    g909_n,
    n5930_o2_n_spl_1,
    n2836_lo_n_spl_001
  );


  and

  (
    g910_p,
    g909_n_spl_,
    g908_n_spl_
  );


  or

  (
    g910_n,
    g909_p_spl_,
    g908_p_spl_
  );


  and

  (
    g911_p,
    g910_n_spl_0,
    g908_n_spl_
  );


  or

  (
    g911_n,
    g910_p_spl_0,
    g908_p_spl_
  );


  and

  (
    g912_p,
    g910_n_spl_0,
    g909_n_spl_
  );


  or

  (
    g912_n,
    g910_p_spl_0,
    g909_p_spl_
  );


  and

  (
    g913_p,
    g912_n,
    g911_n
  );


  or

  (
    g913_n,
    g912_p,
    g911_p
  );


  and

  (
    g914_p,
    g903_n_spl_0,
    g901_n_spl_
  );


  or

  (
    g914_n,
    g903_p_spl_0,
    g901_p_spl_
  );


  and

  (
    g915_p,
    g903_n_spl_,
    g902_n_spl_
  );


  or

  (
    g915_n,
    g903_p_spl_,
    g902_p_spl_
  );


  and

  (
    g916_p,
    g915_n,
    g914_n
  );


  or

  (
    g916_n,
    g915_p,
    g914_p
  );


  and

  (
    g917_p,
    g896_n_spl_0,
    g894_n_spl_
  );


  or

  (
    g917_n,
    g896_p_spl_0,
    g894_p_spl_
  );


  and

  (
    g918_p,
    g896_n_spl_,
    g895_n_spl_
  );


  or

  (
    g918_n,
    g896_p_spl_,
    g895_p_spl_
  );


  and

  (
    g919_p,
    g918_n,
    g917_n
  );


  or

  (
    g919_n,
    g918_p,
    g917_p
  );


  and

  (
    g920_p,
    G4556_o2_n_spl_0,
    G4370_o2_p
  );


  or

  (
    g920_n,
    G4556_o2_p_spl_0,
    G4370_o2_n
  );


  and

  (
    g921_p,
    g920_n_spl_,
    g919_n_spl_
  );


  or

  (
    g921_n,
    g920_p_spl_,
    g919_p_spl_
  );


  and

  (
    g922_p,
    g921_n_spl_0,
    g919_n_spl_
  );


  or

  (
    g922_n,
    g921_p_spl_0,
    g919_p_spl_
  );


  and

  (
    g923_p,
    g921_n_spl_0,
    g920_n_spl_
  );


  or

  (
    g923_n,
    g921_p_spl_0,
    g920_p_spl_
  );


  and

  (
    g924_p,
    g923_n,
    g922_n
  );


  or

  (
    g924_n,
    g923_p,
    g922_p
  );


  and

  (
    g925_p,
    n2824_lo_buf_o2_p_spl_010,
    n5959_o2_p_spl_0
  );


  or

  (
    g925_n,
    n2824_lo_buf_o2_n_spl_010,
    n5959_o2_n_spl_0
  );


  and

  (
    g926_p,
    g925_n_spl_,
    g924_n_spl_
  );


  or

  (
    g926_n,
    g925_p_spl_,
    g924_p_spl_
  );


  and

  (
    g927_p,
    g926_n_spl_0,
    g921_n_spl_
  );


  or

  (
    g927_n,
    g926_p_spl_0,
    g921_p_spl_
  );


  and

  (
    g928_p,
    g927_n_spl_,
    g916_n_spl_
  );


  or

  (
    g928_n,
    g927_p_spl_,
    g916_p_spl_
  );


  and

  (
    g929_p,
    g928_n_spl_0,
    g916_n_spl_
  );


  or

  (
    g929_n,
    g928_p_spl_0,
    g916_p_spl_
  );


  and

  (
    g930_p,
    g928_n_spl_0,
    g927_n_spl_
  );


  or

  (
    g930_n,
    g928_p_spl_0,
    g927_p_spl_
  );


  and

  (
    g931_p,
    g930_n,
    g929_n
  );


  or

  (
    g931_n,
    g930_p,
    g929_p
  );


  and

  (
    g932_p,
    n5959_o2_p_spl_0,
    n2836_lo_p_spl_010
  );


  or

  (
    g932_n,
    n5959_o2_n_spl_0,
    n2836_lo_n_spl_010
  );


  and

  (
    g933_p,
    g932_n_spl_,
    g931_n_spl_
  );


  or

  (
    g933_n,
    g932_p_spl_,
    g931_p_spl_
  );


  and

  (
    g934_p,
    g933_n_spl_0,
    g928_n_spl_
  );


  or

  (
    g934_n,
    g933_p_spl_0,
    g928_p_spl_
  );


  and

  (
    g935_p,
    g934_n_spl_,
    g913_n_spl_
  );


  or

  (
    g935_n,
    g934_p_spl_,
    g913_p_spl_
  );


  and

  (
    g936_p,
    G4556_o2_n_spl_0,
    G4490_o2_p
  );


  or

  (
    g936_n,
    G4556_o2_p_spl_0,
    G4490_o2_n
  );


  and

  (
    g937_p,
    G4556_o2_n_spl_,
    G1007_o2_n
  );


  or

  (
    g937_n,
    G4556_o2_p_spl_,
    G1007_o2_p
  );


  and

  (
    g938_p,
    g937_n,
    g936_n
  );


  or

  (
    g938_n,
    g937_p,
    g936_p
  );


  and

  (
    g939_p,
    G4605_o2_n,
    G4425_o2_p
  );


  or

  (
    g939_n,
    G4605_o2_p,
    G4425_o2_n
  );


  and

  (
    g940_p,
    g939_n_spl_,
    g938_n_spl_
  );


  or

  (
    g940_n,
    g939_p_spl_,
    g938_p_spl_
  );


  and

  (
    g941_p,
    g940_n_spl_0,
    g938_n_spl_
  );


  or

  (
    g941_n,
    g940_p_spl_0,
    g938_p_spl_
  );


  and

  (
    g942_p,
    g940_n_spl_0,
    g939_n_spl_
  );


  or

  (
    g942_n,
    g940_p_spl_0,
    g939_p_spl_
  );


  and

  (
    g943_p,
    g942_n,
    g941_n
  );


  or

  (
    g943_n,
    g942_p,
    g941_p
  );


  and

  (
    g944_p,
    n2824_lo_buf_o2_p_spl_01,
    n5981_o2_p_spl_0
  );


  or

  (
    g944_n,
    n2824_lo_buf_o2_n_spl_01,
    n5981_o2_n_spl_0
  );


  and

  (
    g945_p,
    g944_n_spl_,
    g943_n_spl_
  );


  or

  (
    g945_n,
    g944_p_spl_,
    g943_p_spl_
  );


  and

  (
    g946_p,
    g945_n_spl_0,
    g943_n_spl_
  );


  or

  (
    g946_n,
    g945_p_spl_0,
    g943_p_spl_
  );


  and

  (
    g947_p,
    g945_n_spl_0,
    g944_n_spl_
  );


  or

  (
    g947_n,
    g945_p_spl_0,
    g944_p_spl_
  );


  and

  (
    g948_p,
    g947_n,
    g946_n
  );


  or

  (
    g948_n,
    g947_p,
    g946_p
  );


  and

  (
    g949_p,
    G4719_o2_n_spl_,
    G4716_o2_n_spl_
  );


  or

  (
    g949_n,
    G4719_o2_p_spl_,
    G4716_o2_p_spl_
  );


  and

  (
    g950_p,
    g949_n_spl_0,
    G4719_o2_n_spl_
  );


  or

  (
    g950_n,
    g949_p_spl_0,
    G4719_o2_p_spl_
  );


  and

  (
    g951_p,
    g949_n_spl_0,
    G4716_o2_n_spl_
  );


  or

  (
    g951_n,
    g949_p_spl_0,
    G4716_o2_p_spl_
  );


  and

  (
    g952_p,
    g951_n,
    g950_n
  );


  or

  (
    g952_n,
    g951_p,
    g950_p
  );


  and

  (
    g953_p,
    n2824_lo_buf_o2_p_spl_10,
    n6042_o2_p_spl_0
  );


  or

  (
    g953_n,
    n2824_lo_buf_o2_n_spl_10,
    n6042_o2_n_spl_0
  );


  and

  (
    g954_p,
    g953_n_spl_,
    g952_n_spl_
  );


  or

  (
    g954_n,
    g953_p_spl_,
    g952_p_spl_
  );


  and

  (
    g955_p,
    g954_n_spl_0,
    g949_n_spl_
  );


  or

  (
    g955_n,
    g954_p_spl_0,
    g949_p_spl_
  );


  and

  (
    g956_p,
    g955_n_spl_,
    g948_n_spl_
  );


  or

  (
    g956_n,
    g955_p_spl_,
    g948_p_spl_
  );


  and

  (
    g957_p,
    g956_n_spl_0,
    g948_n_spl_
  );


  or

  (
    g957_n,
    g956_p_spl_0,
    g948_p_spl_
  );


  and

  (
    g958_p,
    g956_n_spl_0,
    g955_n_spl_
  );


  or

  (
    g958_n,
    g956_p_spl_0,
    g955_p_spl_
  );


  and

  (
    g959_p,
    g958_n,
    g957_n
  );


  or

  (
    g959_n,
    g958_p,
    g957_p
  );


  and

  (
    g960_p,
    n6042_o2_p_spl_0,
    n2836_lo_p_spl_010
  );


  or

  (
    g960_n,
    n6042_o2_n_spl_0,
    n2836_lo_n_spl_010
  );


  and

  (
    g961_p,
    g960_n_spl_,
    g959_n_spl_
  );


  or

  (
    g961_n,
    g960_p_spl_,
    g959_p_spl_
  );


  and

  (
    g962_p,
    g961_n_spl_0,
    g959_n_spl_
  );


  or

  (
    g962_n,
    g961_p_spl_0,
    g959_p_spl_
  );


  and

  (
    g963_p,
    g961_n_spl_0,
    g960_n_spl_
  );


  or

  (
    g963_n,
    g961_p_spl_0,
    g960_p_spl_
  );


  and

  (
    g964_p,
    g963_n,
    g962_n
  );


  or

  (
    g964_n,
    g963_p,
    g962_p
  );


  and

  (
    g965_p,
    g954_n_spl_0,
    g952_n_spl_
  );


  or

  (
    g965_n,
    g954_p_spl_0,
    g952_p_spl_
  );


  and

  (
    g966_p,
    g954_n_spl_,
    g953_n_spl_
  );


  or

  (
    g966_n,
    g954_p_spl_,
    g953_p_spl_
  );


  and

  (
    g967_p,
    g966_n,
    g965_n
  );


  or

  (
    g967_n,
    g966_p,
    g965_p
  );


  and

  (
    g968_p,
    G4900_o2_n,
    G4901_o2_n
  );


  or

  (
    g968_n,
    G4900_o2_p,
    G4901_o2_p
  );


  and

  (
    g969_p,
    n2824_lo_buf_o2_p_spl_10,
    n6075_o2_p_spl_0
  );


  or

  (
    g969_n,
    n2824_lo_buf_o2_n_spl_10,
    n6075_o2_n_spl_0
  );


  and

  (
    g970_p,
    g969_n_spl_,
    g968_n_spl_
  );


  or

  (
    g970_n,
    g969_p_spl_,
    g968_p_spl_
  );


  and

  (
    g971_p,
    g970_n_spl_0,
    G4834_o2_p
  );


  or

  (
    g971_n,
    g970_p_spl_0,
    G4834_o2_n
  );


  and

  (
    g972_p,
    g971_n_spl_,
    g967_n_spl_
  );


  or

  (
    g972_n,
    g971_p_spl_,
    g967_p_spl_
  );


  and

  (
    g973_p,
    g972_n_spl_0,
    g967_n_spl_
  );


  or

  (
    g973_n,
    g972_p_spl_0,
    g967_p_spl_
  );


  and

  (
    g974_p,
    g972_n_spl_0,
    g971_n_spl_
  );


  or

  (
    g974_n,
    g972_p_spl_0,
    g971_p_spl_
  );


  and

  (
    g975_p,
    g974_n,
    g973_n
  );


  or

  (
    g975_n,
    g974_p,
    g973_p
  );


  and

  (
    g976_p,
    n6075_o2_p_spl_0,
    n2836_lo_p_spl_011
  );


  or

  (
    g976_n,
    n6075_o2_n_spl_0,
    n2836_lo_n_spl_011
  );


  and

  (
    g977_p,
    g976_n_spl_,
    g975_n_spl_
  );


  or

  (
    g977_n,
    g976_p_spl_,
    g975_p_spl_
  );


  and

  (
    g978_p,
    g977_n_spl_0,
    g972_n_spl_
  );


  or

  (
    g978_n,
    g977_p_spl_0,
    g972_p_spl_
  );


  and

  (
    g979_p,
    g978_n_spl_,
    g964_n_spl_
  );


  or

  (
    g979_n,
    g978_p_spl_,
    g964_p_spl_
  );


  and

  (
    g980_p,
    g979_n_spl_0,
    g964_n_spl_
  );


  or

  (
    g980_n,
    g979_p_spl_0,
    g964_p_spl_
  );


  and

  (
    g981_p,
    g979_n_spl_0,
    g978_n_spl_
  );


  or

  (
    g981_n,
    g979_p_spl_0,
    g978_p_spl_
  );


  and

  (
    g982_p,
    g981_n,
    g980_n
  );


  or

  (
    g982_n,
    g981_p,
    g980_p
  );


  and

  (
    g983_p,
    n6075_o2_p_spl_,
    n2848_lo_p_spl_001
  );


  or

  (
    g983_n,
    n6075_o2_n_spl_1,
    n2848_lo_n_spl_001
  );


  and

  (
    g984_p,
    g983_n_spl_,
    g982_n_spl_
  );


  or

  (
    g984_n,
    g983_p_spl_,
    g982_p_spl_
  );


  and

  (
    g985_p,
    g984_n_spl_0,
    g982_n_spl_
  );


  or

  (
    g985_n,
    g984_p_spl_0,
    g982_p_spl_
  );


  and

  (
    g986_p,
    g984_n_spl_0,
    g983_n_spl_
  );


  or

  (
    g986_n,
    g984_p_spl_0,
    g983_p_spl_
  );


  and

  (
    g987_p,
    g986_n,
    g985_n
  );


  or

  (
    g987_n,
    g986_p,
    g985_p
  );


  and

  (
    g988_p,
    g977_n_spl_0,
    g975_n_spl_
  );


  or

  (
    g988_n,
    g977_p_spl_0,
    g975_p_spl_
  );


  and

  (
    g989_p,
    g977_n_spl_,
    g976_n_spl_
  );


  or

  (
    g989_n,
    g977_p_spl_,
    g976_p_spl_
  );


  and

  (
    g990_p,
    g989_n,
    g988_n
  );


  or

  (
    g990_n,
    g989_p,
    g988_p
  );


  and

  (
    g991_p,
    g970_n_spl_0,
    g968_n_spl_
  );


  or

  (
    g991_n,
    g970_p_spl_0,
    g968_p_spl_
  );


  and

  (
    g992_p,
    g970_n_spl_,
    g969_n_spl_
  );


  or

  (
    g992_n,
    g970_p_spl_,
    g969_p_spl_
  );


  and

  (
    g993_p,
    g992_n,
    g991_n
  );


  or

  (
    g993_n,
    g992_p,
    g991_p
  );


  and

  (
    g994_p,
    G5064_o2_n_spl_0,
    G4896_o2_p
  );


  or

  (
    g994_n,
    G5064_o2_p_spl_0,
    G4896_o2_n
  );


  and

  (
    g995_p,
    g994_n_spl_,
    g993_n_spl_
  );


  or

  (
    g995_n,
    g994_p_spl_,
    g993_p_spl_
  );


  and

  (
    g996_p,
    g995_n_spl_0,
    g993_n_spl_
  );


  or

  (
    g996_n,
    g995_p_spl_0,
    g993_p_spl_
  );


  and

  (
    g997_p,
    g995_n_spl_0,
    g994_n_spl_
  );


  or

  (
    g997_n,
    g995_p_spl_0,
    g994_p_spl_
  );


  and

  (
    g998_p,
    g997_n,
    g996_n
  );


  or

  (
    g998_n,
    g997_p,
    g996_p
  );


  and

  (
    g999_p,
    n6103_o2_p_spl_0,
    n2836_lo_p_spl_011
  );


  or

  (
    g999_n,
    n6103_o2_n_spl_0,
    n2836_lo_n_spl_011
  );


  and

  (
    g1000_p,
    g999_n_spl_,
    g998_n_spl_
  );


  or

  (
    g1000_n,
    g999_p_spl_,
    g998_p_spl_
  );


  and

  (
    g1001_p,
    g1000_n_spl_0,
    g995_n_spl_
  );


  or

  (
    g1001_n,
    g1000_p_spl_0,
    g995_p_spl_
  );


  and

  (
    g1002_p,
    g1001_n_spl_,
    g990_n_spl_
  );


  or

  (
    g1002_n,
    g1001_p_spl_,
    g990_p_spl_
  );


  and

  (
    g1003_p,
    g1002_n_spl_0,
    g990_n_spl_
  );


  or

  (
    g1003_n,
    g1002_p_spl_0,
    g990_p_spl_
  );


  and

  (
    g1004_p,
    g1002_n_spl_0,
    g1001_n_spl_
  );


  or

  (
    g1004_n,
    g1002_p_spl_0,
    g1001_p_spl_
  );


  and

  (
    g1005_p,
    g1004_n,
    g1003_n
  );


  or

  (
    g1005_n,
    g1004_p,
    g1003_p
  );


  and

  (
    g1006_p,
    n6103_o2_p_spl_0,
    n2848_lo_p_spl_001
  );


  or

  (
    g1006_n,
    n6103_o2_n_spl_0,
    n2848_lo_n_spl_001
  );


  and

  (
    g1007_p,
    g1006_n_spl_,
    g1005_n_spl_
  );


  or

  (
    g1007_n,
    g1006_p_spl_,
    g1005_p_spl_
  );


  and

  (
    g1008_p,
    g1007_n_spl_0,
    g1002_n_spl_
  );


  or

  (
    g1008_n,
    g1007_p_spl_0,
    g1002_p_spl_
  );


  and

  (
    g1009_p,
    g1008_n_spl_,
    g987_n_spl_
  );


  or

  (
    g1009_n,
    g1008_p_spl_,
    g987_p_spl_
  );


  and

  (
    g1010_p,
    G5247_o2_n_spl_,
    G5244_o2_n_spl_
  );


  or

  (
    g1010_n,
    G5247_o2_p_spl_,
    G5244_o2_p_spl_
  );


  and

  (
    g1011_p,
    g1010_n_spl_0,
    G5247_o2_n_spl_
  );


  or

  (
    g1011_n,
    g1010_p_spl_0,
    G5247_o2_p_spl_
  );


  and

  (
    g1012_p,
    g1010_n_spl_0,
    G5244_o2_n_spl_
  );


  or

  (
    g1012_n,
    g1010_p_spl_0,
    G5244_o2_p_spl_
  );


  and

  (
    g1013_p,
    g1012_n,
    g1011_n
  );


  or

  (
    g1013_n,
    g1012_p,
    g1011_p
  );


  and

  (
    g1014_p,
    n6205_o2_p_spl_0,
    n2836_lo_p_spl_100
  );


  or

  (
    g1014_n,
    n6205_o2_n_spl_0,
    n2836_lo_n_spl_100
  );


  and

  (
    g1015_p,
    g1014_n_spl_,
    g1013_n_spl_
  );


  or

  (
    g1015_n,
    g1014_p_spl_,
    g1013_p_spl_
  );


  and

  (
    g1016_p,
    g1015_n_spl_0,
    g1013_n_spl_
  );


  or

  (
    g1016_n,
    g1015_p_spl_0,
    g1013_p_spl_
  );


  and

  (
    g1017_p,
    g1015_n_spl_0,
    g1014_n_spl_
  );


  or

  (
    g1017_n,
    g1015_p_spl_0,
    g1014_p_spl_
  );


  and

  (
    g1018_p,
    g1017_n,
    g1016_n
  );


  or

  (
    g1018_n,
    g1017_p,
    g1016_p
  );


  and

  (
    g1019_p,
    g744_n_spl_,
    g739_n_spl_
  );


  or

  (
    g1019_n,
    g744_p_spl_,
    g739_p_spl_
  );


  and

  (
    g1020_p,
    g1019_n_spl_,
    g1018_n_spl_
  );


  or

  (
    g1020_n,
    g1019_p_spl_,
    g1018_p_spl_
  );


  and

  (
    g1021_p,
    g1020_n_spl_0,
    g1018_n_spl_
  );


  or

  (
    g1021_n,
    g1020_p_spl_0,
    g1018_p_spl_
  );


  and

  (
    g1022_p,
    g1020_n_spl_0,
    g1019_n_spl_
  );


  or

  (
    g1022_n,
    g1020_p_spl_0,
    g1019_p_spl_
  );


  and

  (
    g1023_p,
    g1022_n,
    g1021_n
  );


  or

  (
    g1023_n,
    g1022_p,
    g1021_p
  );


  and

  (
    g1024_p,
    n6239_o2_p_spl_0,
    n2848_lo_p_spl_010
  );


  or

  (
    g1024_n,
    n6239_o2_n_spl_0,
    n2848_lo_n_spl_010
  );


  and

  (
    g1025_p,
    g1024_n_spl_,
    g1023_n_spl_
  );


  or

  (
    g1025_n,
    g1024_p_spl_,
    g1023_p_spl_
  );


  and

  (
    g1026_p,
    g1025_n_spl_0,
    g1023_n_spl_
  );


  or

  (
    g1026_n,
    g1025_p_spl_0,
    g1023_p_spl_
  );


  and

  (
    g1027_p,
    g1025_n_spl_0,
    g1024_n_spl_
  );


  or

  (
    g1027_n,
    g1025_p_spl_0,
    g1024_p_spl_
  );


  and

  (
    g1028_p,
    g1027_n,
    g1026_n
  );


  or

  (
    g1028_n,
    g1027_p,
    g1026_p
  );


  and

  (
    g1029_p,
    g754_n_spl_,
    g749_n_spl_
  );


  or

  (
    g1029_n,
    g754_p_spl_,
    g749_p_spl_
  );


  and

  (
    g1030_p,
    g1029_n_spl_,
    g1028_n_spl_
  );


  or

  (
    g1030_n,
    g1029_p_spl_,
    g1028_p_spl_
  );


  and

  (
    g1031_p,
    g1030_n_spl_0,
    g1028_n_spl_
  );


  or

  (
    g1031_n,
    g1030_p_spl_0,
    g1028_p_spl_
  );


  and

  (
    g1032_p,
    g1030_n_spl_0,
    g1029_n_spl_
  );


  or

  (
    g1032_n,
    g1030_p_spl_0,
    g1029_p_spl_
  );


  and

  (
    g1033_p,
    g1032_n,
    g1031_n
  );


  or

  (
    g1033_n,
    g1032_p,
    g1031_p
  );


  and

  (
    g1034_p,
    n6309_o2_p_spl_,
    n2860_lo_p_spl_00
  );


  or

  (
    g1034_n,
    n6309_o2_n_spl_,
    n2860_lo_n_spl_00
  );


  and

  (
    g1035_p,
    g1034_n_spl_,
    g1033_n_spl_
  );


  or

  (
    g1035_n,
    g1034_p_spl_,
    g1033_p_spl_
  );


  and

  (
    g1036_p,
    g1035_n_spl_0,
    g1033_n_spl_
  );


  or

  (
    g1036_n,
    g1035_p_spl_0,
    g1033_p_spl_
  );


  and

  (
    g1037_p,
    g1035_n_spl_0,
    g1034_n_spl_
  );


  or

  (
    g1037_n,
    g1035_p_spl_0,
    g1034_p_spl_
  );


  and

  (
    g1038_p,
    g1037_n,
    g1036_n
  );


  or

  (
    g1038_n,
    g1037_p,
    g1036_p
  );


  and

  (
    g1039_p,
    g764_n,
    g759_n_spl_
  );


  or

  (
    g1039_n,
    g764_p_spl_,
    g759_p_spl_
  );


  and

  (
    g1040_p,
    g1039_n_spl_,
    g1038_n_spl_
  );


  or

  (
    g1040_n,
    g1039_p,
    g1038_p
  );


  and

  (
    g1041_p,
    g1040_n_spl_,
    g1038_n_spl_
  );


  and

  (
    g1042_p,
    g1040_n_spl_,
    g1039_n_spl_
  );


  or

  (
    g1043_n,
    g1042_p,
    g1041_p
  );


  and

  (
    g1044_p,
    g817_n_spl_,
    g804_n
  );


  or

  (
    g1044_n,
    g817_p,
    g804_p_spl_
  );


  and

  (
    g1045_p,
    n8086_o2_p_spl_01,
    n2797_lo_p_spl_000
  );


  or

  (
    g1045_n,
    n8086_o2_n_spl_1,
    n2797_lo_n_spl_000
  );


  and

  (
    g1046_p,
    G3422_o2_n_spl_0,
    G3367_o2_p
  );


  or

  (
    g1046_n,
    G3422_o2_p_spl_0,
    G3367_o2_n
  );


  and

  (
    g1047_p,
    G3422_o2_n_spl_0,
    G707_o2_n
  );


  or

  (
    g1047_n,
    G3422_o2_p_spl_0,
    G707_o2_p
  );


  and

  (
    g1048_p,
    g1047_n,
    g1046_n
  );


  or

  (
    g1048_n,
    g1047_p,
    g1046_p
  );


  and

  (
    g1049_p,
    g784_n_spl_,
    G3265_o2_p
  );


  or

  (
    g1049_n,
    g784_p_spl_,
    G3265_o2_n
  );


  and

  (
    g1050_p,
    g1049_n_spl_,
    g1048_n_spl_
  );


  or

  (
    g1050_n,
    g1049_p_spl_,
    g1048_p_spl_
  );


  and

  (
    g1051_p,
    g1050_n_spl_0,
    g1048_n_spl_
  );


  or

  (
    g1051_n,
    g1050_p_spl_0,
    g1048_p_spl_
  );


  and

  (
    g1052_p,
    g1050_n_spl_0,
    g1049_n_spl_
  );


  or

  (
    g1052_n,
    g1050_p_spl_0,
    g1049_p_spl_
  );


  and

  (
    g1053_p,
    g1052_n,
    g1051_n
  );


  or

  (
    g1053_n,
    g1052_p,
    g1051_p
  );


  and

  (
    g1054_p,
    n2776_lo_buf_o2_p_spl_001,
    n7835_o2_p_spl_00
  );


  or

  (
    g1054_n,
    n2776_lo_buf_o2_n_spl_001,
    n7835_o2_n_spl_00
  );


  and

  (
    g1055_p,
    g1054_n_spl_,
    g1053_n_spl_
  );


  or

  (
    g1055_n,
    g1054_p_spl_,
    g1053_p_spl_
  );


  and

  (
    g1056_p,
    g1055_n_spl_0,
    g1053_n_spl_
  );


  or

  (
    g1056_n,
    g1055_p_spl_0,
    g1053_p_spl_
  );


  and

  (
    g1057_p,
    g1055_n_spl_0,
    g1054_n_spl_
  );


  or

  (
    g1057_n,
    g1055_p_spl_0,
    g1054_p_spl_
  );


  and

  (
    g1058_p,
    g1057_n,
    g1056_n
  );


  or

  (
    g1058_n,
    g1057_p,
    g1056_p
  );


  and

  (
    g1059_p,
    g794_n_spl_,
    g789_n_spl_
  );


  or

  (
    g1059_n,
    g794_p_spl_,
    g789_p_spl_
  );


  and

  (
    g1060_p,
    g1059_n_spl_,
    g1058_n_spl_
  );


  or

  (
    g1060_n,
    g1059_p_spl_,
    g1058_p_spl_
  );


  and

  (
    g1061_p,
    g1060_n_spl_0,
    g1058_n_spl_
  );


  or

  (
    g1061_n,
    g1060_p_spl_0,
    g1058_p_spl_
  );


  and

  (
    g1062_p,
    g1060_n_spl_0,
    g1059_n_spl_
  );


  or

  (
    g1062_n,
    g1060_p_spl_0,
    g1059_p_spl_
  );


  and

  (
    g1063_p,
    g1062_n,
    g1061_n
  );


  or

  (
    g1063_n,
    g1062_p,
    g1061_p
  );


  and

  (
    g1064_p,
    n7909_o2_p_spl_01,
    n2785_lo_p_spl_000
  );


  or

  (
    g1064_n,
    n7909_o2_n_spl_0,
    n2785_lo_n_spl_000
  );


  and

  (
    g1065_p,
    g1064_n_spl_,
    g1063_n_spl_
  );


  or

  (
    g1065_n,
    g1064_p_spl_,
    g1063_p_spl_
  );


  and

  (
    g1066_p,
    g1065_n_spl_0,
    g1063_n_spl_
  );


  or

  (
    g1066_n,
    g1065_p_spl_0,
    g1063_p_spl_
  );


  and

  (
    g1067_p,
    g1065_n_spl_0,
    g1064_n_spl_
  );


  or

  (
    g1067_n,
    g1065_p_spl_0,
    g1064_p_spl_
  );


  and

  (
    g1068_p,
    g1067_n,
    g1066_n
  );


  or

  (
    g1068_n,
    g1067_p,
    g1066_p
  );


  and

  (
    g1069_p,
    g803_n,
    g799_n_spl_
  );


  or

  (
    g1069_n,
    g803_p_spl_,
    g799_p_spl_
  );


  and

  (
    g1070_p,
    g1069_n_spl_,
    g1068_n_spl_
  );


  or

  (
    g1070_n,
    g1069_p_spl_,
    g1068_p_spl_
  );


  and

  (
    g1071_p,
    g1070_n_spl_0,
    g1068_n_spl_
  );


  or

  (
    g1071_n,
    g1070_p_spl_0,
    g1068_p_spl_
  );


  and

  (
    g1072_p,
    g1070_n_spl_0,
    g1069_n_spl_
  );


  or

  (
    g1072_n,
    g1070_p_spl_0,
    g1069_p_spl_
  );


  and

  (
    g1073_p,
    g1072_n,
    g1071_n
  );


  or

  (
    g1073_n,
    g1072_p,
    g1071_p
  );


  and

  (
    g1074_p,
    n2728_lo_buf_o2_p_spl_000,
    n2488_lo_buf_o2_p_spl_0
  );


  or

  (
    g1074_n,
    n2728_lo_buf_o2_n_spl_000,
    n2488_lo_buf_o2_n_spl_0
  );


  and

  (
    g1075_p,
    g1073_n_spl_,
    g1045_n
  );


  or

  (
    g1075_n,
    g1073_p,
    g1045_p_spl_
  );


  and

  (
    g1076_p,
    G1688_o2_n,
    G1689_o2_n
  );


  or

  (
    g1076_n,
    G1688_o2_p,
    G1689_o2_p
  );


  and

  (
    g1077_p,
    n2512_lo_buf_o2_p_spl_00,
    n2704_lo_buf_o2_p_spl_
  );


  or

  (
    g1077_n,
    n2512_lo_buf_o2_n_spl_00,
    n2704_lo_buf_o2_n_spl_
  );


  and

  (
    g1078_p,
    g1077_n_spl_,
    g1076_n_spl_
  );


  or

  (
    g1078_n,
    g1077_p_spl_,
    g1076_p_spl_
  );


  and

  (
    g1079_p,
    g1078_n_spl_0,
    g1076_n_spl_
  );


  or

  (
    g1079_n,
    g1078_p_spl_0,
    g1076_p_spl_
  );


  and

  (
    g1080_p,
    g1078_n_spl_0,
    g1077_n_spl_
  );


  or

  (
    g1080_n,
    g1078_p_spl_0,
    g1077_p_spl_
  );


  and

  (
    g1081_p,
    g1080_n,
    g1079_n
  );


  or

  (
    g1081_n,
    g1080_p,
    g1079_p
  );


  and

  (
    g1082_p,
    g809_n_spl_,
    G1630_o2_p_spl_
  );


  or

  (
    g1082_n,
    g809_p_spl_,
    G1630_o2_n_spl_
  );


  and

  (
    g1083_p,
    g1082_n_spl_,
    g1081_n_spl_
  );


  or

  (
    g1083_n,
    g1082_p_spl_,
    g1081_p_spl_
  );


  and

  (
    g1084_p,
    g1083_n_spl_0,
    g1081_n_spl_
  );


  or

  (
    g1084_n,
    g1083_p_spl_0,
    g1081_p_spl_
  );


  and

  (
    g1085_p,
    g1083_n_spl_0,
    g1082_n_spl_
  );


  or

  (
    g1085_n,
    g1083_p_spl_0,
    g1082_p_spl_
  );


  and

  (
    g1086_p,
    g1085_n,
    g1084_n
  );


  or

  (
    g1086_n,
    g1085_p,
    g1084_p
  );


  and

  (
    g1087_p,
    n2716_lo_buf_o2_p_spl_000,
    n2500_lo_buf_o2_p_spl_00
  );


  or

  (
    g1087_n,
    n2716_lo_buf_o2_n_spl_000,
    n2500_lo_buf_o2_n_spl_00
  );


  and

  (
    g1088_p,
    g1087_n_spl_,
    g1086_n_spl_
  );


  or

  (
    g1088_n,
    g1087_p_spl_,
    g1086_p_spl_
  );


  and

  (
    g1089_p,
    g1088_n_spl_0,
    g1086_n_spl_
  );


  or

  (
    g1089_n,
    g1088_p_spl_0,
    g1086_p_spl_
  );


  and

  (
    g1090_p,
    g1088_n_spl_0,
    g1087_n_spl_
  );


  or

  (
    g1090_n,
    g1088_p_spl_0,
    g1087_p_spl_
  );


  and

  (
    g1091_p,
    g1090_n,
    g1089_n
  );


  or

  (
    g1091_n,
    g1090_p,
    g1089_p
  );


  and

  (
    g1092_p,
    g1044_n,
    g814_n_spl_
  );


  or

  (
    g1092_n,
    g1044_p_spl_,
    g814_p_spl_
  );


  and

  (
    g1093_p,
    g1092_n_spl_,
    g1091_n_spl_
  );


  or

  (
    g1093_n,
    g1092_p_spl_,
    g1091_p_spl_
  );


  and

  (
    g1094_p,
    g1093_n_spl_0,
    g1091_n_spl_
  );


  or

  (
    g1094_n,
    g1093_p_spl_0,
    g1091_p_spl_
  );


  and

  (
    g1095_p,
    g1093_n_spl_0,
    g1092_n_spl_
  );


  or

  (
    g1095_n,
    g1093_p_spl_0,
    g1092_p_spl_
  );


  and

  (
    g1096_p,
    g1095_n,
    g1094_n
  );


  or

  (
    g1096_n,
    g1095_p,
    g1094_p
  );


  and

  (
    g1097_p,
    g1096_n_spl_,
    g1074_n
  );


  or

  (
    g1097_n,
    g1096_p,
    g1074_p_spl_
  );


  or

  (
    g1098_n,
    g1043_n_spl_0,
    g1040_p
  );


  and

  (
    g1099_p,
    n2824_lo_buf_o2_p_spl_11,
    n5779_o2_p_spl_1
  );


  or

  (
    g1099_n,
    n2824_lo_buf_o2_n_spl_11,
    n5779_o2_n_spl_
  );


  and

  (
    g1100_p,
    g836_n_spl_,
    g831_n_spl_
  );


  or

  (
    g1100_n,
    g836_p_spl_,
    g831_p_spl_
  );


  or

  (
    g1101_n,
    g1100_p,
    g1099_p
  );


  and

  (
    g1102_p,
    g852_n_spl_0,
    g850_n_spl_
  );


  or

  (
    g1102_n,
    g852_p_spl_0,
    g850_p_spl_
  );


  and

  (
    g1103_p,
    g852_n_spl_,
    g851_n_spl_
  );


  or

  (
    g1103_n,
    g852_p_spl_,
    g851_p_spl_
  );


  and

  (
    g1104_p,
    g1103_n,
    g1102_n
  );


  or

  (
    g1104_n,
    g1103_p,
    g1102_p
  );


  and

  (
    g1105_p,
    g871_n_spl_,
    g866_n_spl_
  );


  or

  (
    g1105_n,
    g871_p_spl_,
    g866_p_spl_
  );


  and

  (
    g1106_p,
    g1105_n_spl_,
    g1104_n_spl_
  );


  or

  (
    g1106_n,
    g1105_p_spl_,
    g1104_p_spl_
  );


  and

  (
    g1107_p,
    g1106_n_spl_0,
    g1104_n_spl_
  );


  or

  (
    g1107_n,
    g1106_p_spl_0,
    g1104_p_spl_
  );


  and

  (
    g1108_p,
    g1106_n_spl_0,
    g1105_n_spl_
  );


  or

  (
    g1108_n,
    g1106_p_spl_0,
    g1105_p_spl_
  );


  and

  (
    g1109_p,
    g1108_n,
    g1107_n
  );


  or

  (
    g1109_n,
    g1108_p,
    g1107_p
  );


  and

  (
    g1110_p,
    n2824_lo_buf_o2_p_spl_11,
    n5863_o2_p_spl_0
  );


  or

  (
    g1110_n,
    n2824_lo_buf_o2_n_spl_11,
    n5863_o2_n_spl_0
  );


  and

  (
    g1111_p,
    g1110_n_spl_,
    g1109_n_spl_
  );


  or

  (
    g1111_n,
    g1110_p_spl_,
    g1109_p_spl_
  );


  and

  (
    g1112_p,
    g1111_n_spl_0,
    g1109_n_spl_
  );


  or

  (
    g1112_n,
    g1111_p_spl_0,
    g1109_p_spl_
  );


  and

  (
    g1113_p,
    g1111_n_spl_0,
    g1110_n_spl_
  );


  or

  (
    g1113_n,
    g1111_p_spl_0,
    g1110_p_spl_
  );


  and

  (
    g1114_p,
    g1113_n,
    g1112_n
  );


  or

  (
    g1114_n,
    g1113_p,
    g1112_p
  );


  and

  (
    g1115_p,
    g887_n_spl_,
    g882_n_spl_
  );


  or

  (
    g1115_n,
    g887_p_spl_,
    g882_p_spl_
  );


  and

  (
    g1116_p,
    g1115_n_spl_,
    g1114_n_spl_
  );


  or

  (
    g1116_n,
    g1115_p_spl_,
    g1114_p_spl_
  );


  and

  (
    g1117_p,
    g1116_n_spl_0,
    g1114_n_spl_
  );


  or

  (
    g1117_n,
    g1116_p_spl_0,
    g1114_p_spl_
  );


  and

  (
    g1118_p,
    g1116_n_spl_0,
    g1115_n_spl_
  );


  or

  (
    g1118_n,
    g1116_p_spl_0,
    g1115_p_spl_
  );


  and

  (
    g1119_p,
    g1118_n,
    g1117_n
  );


  or

  (
    g1119_n,
    g1118_p,
    g1117_p
  );


  and

  (
    g1120_p,
    n5881_o2_p_spl_1,
    n2836_lo_p_spl_100
  );


  or

  (
    g1120_n,
    n5881_o2_n_spl_,
    n2836_lo_n_spl_100
  );


  and

  (
    g1121_p,
    g1120_n_spl_,
    g1119_n_spl_
  );


  or

  (
    g1121_n,
    g1120_p_spl_,
    g1119_p_spl_
  );


  and

  (
    g1122_p,
    g1121_n_spl_0,
    g1119_n_spl_
  );


  or

  (
    g1122_n,
    g1121_p_spl_0,
    g1119_p_spl_
  );


  and

  (
    g1123_p,
    g1121_n_spl_0,
    g1120_n_spl_
  );


  or

  (
    g1123_n,
    g1121_p_spl_0,
    g1120_p_spl_
  );


  and

  (
    g1124_p,
    g1123_n,
    g1122_n
  );


  or

  (
    g1124_n,
    g1123_p,
    g1122_p
  );


  and

  (
    g1125_p,
    g910_n_spl_,
    g905_n_spl_
  );


  or

  (
    g1125_n,
    g910_p_spl_,
    g905_p_spl_
  );


  or

  (
    g1126_n,
    g1125_p,
    g1124_p
  );


  and

  (
    g1127_p,
    g926_n_spl_0,
    g924_n_spl_
  );


  or

  (
    g1127_n,
    g926_p_spl_0,
    g924_p_spl_
  );


  and

  (
    g1128_p,
    g926_n_spl_,
    g925_n_spl_
  );


  or

  (
    g1128_n,
    g926_p_spl_,
    g925_p_spl_
  );


  and

  (
    g1129_p,
    g1128_n,
    g1127_n
  );


  or

  (
    g1129_n,
    g1128_p,
    g1127_p
  );


  and

  (
    g1130_p,
    g945_n_spl_,
    g940_n_spl_
  );


  or

  (
    g1130_n,
    g945_p_spl_,
    g940_p_spl_
  );


  and

  (
    g1131_p,
    g1130_n_spl_,
    g1129_n_spl_
  );


  or

  (
    g1131_n,
    g1130_p_spl_,
    g1129_p_spl_
  );


  and

  (
    g1132_p,
    g1131_n_spl_0,
    g1129_n_spl_
  );


  or

  (
    g1132_n,
    g1131_p_spl_0,
    g1129_p_spl_
  );


  and

  (
    g1133_p,
    g1131_n_spl_0,
    g1130_n_spl_
  );


  or

  (
    g1133_n,
    g1131_p_spl_0,
    g1130_p_spl_
  );


  and

  (
    g1134_p,
    g1133_n,
    g1132_n
  );


  or

  (
    g1134_n,
    g1133_p,
    g1132_p
  );


  and

  (
    g1135_p,
    n5981_o2_p_spl_0,
    n2836_lo_p_spl_101
  );


  or

  (
    g1135_n,
    n5981_o2_n_spl_0,
    n2836_lo_n_spl_101
  );


  and

  (
    g1136_p,
    g1135_n_spl_,
    g1134_n_spl_
  );


  or

  (
    g1136_n,
    g1135_p_spl_,
    g1134_p_spl_
  );


  and

  (
    g1137_p,
    g1136_n_spl_0,
    g1134_n_spl_
  );


  or

  (
    g1137_n,
    g1136_p_spl_0,
    g1134_p_spl_
  );


  and

  (
    g1138_p,
    g1136_n_spl_0,
    g1135_n_spl_
  );


  or

  (
    g1138_n,
    g1136_p_spl_0,
    g1135_p_spl_
  );


  and

  (
    g1139_p,
    g1138_n,
    g1137_n
  );


  or

  (
    g1139_n,
    g1138_p,
    g1137_p
  );


  and

  (
    g1140_p,
    g961_n_spl_,
    g956_n_spl_
  );


  or

  (
    g1140_n,
    g961_p_spl_,
    g956_p_spl_
  );


  and

  (
    g1141_p,
    g1140_n_spl_,
    g1139_n_spl_
  );


  or

  (
    g1141_n,
    g1140_p_spl_,
    g1139_p_spl_
  );


  and

  (
    g1142_p,
    g1141_n_spl_0,
    g1139_n_spl_
  );


  or

  (
    g1142_n,
    g1141_p_spl_0,
    g1139_p_spl_
  );


  and

  (
    g1143_p,
    g1141_n_spl_0,
    g1140_n_spl_
  );


  or

  (
    g1143_n,
    g1141_p_spl_0,
    g1140_p_spl_
  );


  and

  (
    g1144_p,
    g1143_n,
    g1142_n
  );


  or

  (
    g1144_n,
    g1143_p,
    g1142_p
  );


  and

  (
    g1145_p,
    n6042_o2_p_spl_1,
    n2848_lo_p_spl_010
  );


  or

  (
    g1145_n,
    n6042_o2_n_spl_,
    n2848_lo_n_spl_010
  );


  and

  (
    g1146_p,
    g1145_n_spl_,
    g1144_n_spl_
  );


  or

  (
    g1146_n,
    g1145_p_spl_,
    g1144_p_spl_
  );


  and

  (
    g1147_p,
    g1146_n_spl_0,
    g1144_n_spl_
  );


  or

  (
    g1147_n,
    g1146_p_spl_0,
    g1144_p_spl_
  );


  and

  (
    g1148_p,
    g1146_n_spl_0,
    g1145_n_spl_
  );


  or

  (
    g1148_n,
    g1146_p_spl_0,
    g1145_p_spl_
  );


  and

  (
    g1149_p,
    g1148_n,
    g1147_n
  );


  or

  (
    g1149_n,
    g1148_p,
    g1147_p
  );


  and

  (
    g1150_p,
    g984_n_spl_,
    g979_n_spl_
  );


  or

  (
    g1150_n,
    g984_p_spl_,
    g979_p_spl_
  );


  or

  (
    g1151_n,
    g1150_p,
    g1149_p
  );


  and

  (
    g1152_p,
    g1000_n_spl_0,
    g998_n_spl_
  );


  or

  (
    g1152_n,
    g1000_p_spl_0,
    g998_p_spl_
  );


  and

  (
    g1153_p,
    g1000_n_spl_,
    g999_n_spl_
  );


  or

  (
    g1153_n,
    g1000_p_spl_,
    g999_p_spl_
  );


  and

  (
    g1154_p,
    g1153_n,
    g1152_n
  );


  or

  (
    g1154_n,
    g1153_p,
    g1152_p
  );


  and

  (
    g1155_p,
    G5064_o2_n_spl_0,
    G5011_o2_p
  );


  or

  (
    g1155_n,
    G5064_o2_p_spl_0,
    G5011_o2_n
  );


  and

  (
    g1156_p,
    G5064_o2_n_spl_,
    G818_o2_n
  );


  or

  (
    g1156_n,
    G5064_o2_p_spl_,
    G818_o2_p
  );


  and

  (
    g1157_p,
    g1156_n,
    g1155_n
  );


  or

  (
    g1157_n,
    g1156_p,
    g1155_p
  );


  and

  (
    g1158_p,
    G5118_o2_n,
    G4947_o2_p
  );


  or

  (
    g1158_n,
    G5118_o2_p,
    G4947_o2_n
  );


  and

  (
    g1159_p,
    g1158_n_spl_,
    g1157_n_spl_
  );


  or

  (
    g1159_n,
    g1158_p_spl_,
    g1157_p_spl_
  );


  and

  (
    g1160_p,
    g1159_n_spl_0,
    g1157_n_spl_
  );


  or

  (
    g1160_n,
    g1159_p_spl_0,
    g1157_p_spl_
  );


  and

  (
    g1161_p,
    g1159_n_spl_0,
    g1158_n_spl_
  );


  or

  (
    g1161_n,
    g1159_p_spl_0,
    g1158_p_spl_
  );


  and

  (
    g1162_p,
    g1161_n,
    g1160_n
  );


  or

  (
    g1162_n,
    g1161_p,
    g1160_p
  );


  and

  (
    g1163_p,
    n6169_o2_p_spl_0,
    n2836_lo_p_spl_101
  );


  or

  (
    g1163_n,
    n6169_o2_n_spl_0,
    n2836_lo_n_spl_101
  );


  and

  (
    g1164_p,
    g1163_n_spl_,
    g1162_n_spl_
  );


  or

  (
    g1164_n,
    g1163_p_spl_,
    g1162_p_spl_
  );


  and

  (
    g1165_p,
    g1164_n_spl_0,
    g1159_n_spl_
  );


  or

  (
    g1165_n,
    g1164_p_spl_0,
    g1159_p_spl_
  );


  and

  (
    g1166_p,
    g1165_n_spl_,
    g1154_n_spl_
  );


  or

  (
    g1166_n,
    g1165_p_spl_,
    g1154_p_spl_
  );


  and

  (
    g1167_p,
    g1166_n_spl_0,
    g1154_n_spl_
  );


  or

  (
    g1167_n,
    g1166_p_spl_0,
    g1154_p_spl_
  );


  and

  (
    g1168_p,
    g1166_n_spl_0,
    g1165_n_spl_
  );


  or

  (
    g1168_n,
    g1166_p_spl_0,
    g1165_p_spl_
  );


  and

  (
    g1169_p,
    g1168_n,
    g1167_n
  );


  or

  (
    g1169_n,
    g1168_p,
    g1167_p
  );


  and

  (
    g1170_p,
    n6169_o2_p_spl_0,
    n2848_lo_p_spl_01
  );


  or

  (
    g1170_n,
    n6169_o2_n_spl_0,
    n2848_lo_n_spl_01
  );


  and

  (
    g1171_p,
    g1170_n_spl_,
    g1169_n_spl_
  );


  or

  (
    g1171_n,
    g1170_p_spl_,
    g1169_p_spl_
  );


  and

  (
    g1172_p,
    g1171_n_spl_0,
    g1169_n_spl_
  );


  or

  (
    g1172_n,
    g1171_p_spl_0,
    g1169_p_spl_
  );


  and

  (
    g1173_p,
    g1171_n_spl_0,
    g1170_n_spl_
  );


  or

  (
    g1173_n,
    g1171_p_spl_0,
    g1170_p_spl_
  );


  and

  (
    g1174_p,
    g1173_n,
    g1172_n
  );


  or

  (
    g1174_n,
    g1173_p,
    g1172_p
  );


  and

  (
    g1175_p,
    g1164_n_spl_0,
    g1162_n_spl_
  );


  or

  (
    g1175_n,
    g1164_p_spl_0,
    g1162_p_spl_
  );


  and

  (
    g1176_p,
    g1164_n_spl_,
    g1163_n_spl_
  );


  or

  (
    g1176_n,
    g1164_p_spl_,
    g1163_p_spl_
  );


  and

  (
    g1177_p,
    g1176_n,
    g1175_n
  );


  or

  (
    g1177_n,
    g1176_p,
    g1175_p
  );


  and

  (
    g1178_p,
    g1015_n_spl_,
    g1010_n_spl_
  );


  or

  (
    g1178_n,
    g1015_p_spl_,
    g1010_p_spl_
  );


  and

  (
    g1179_p,
    g1178_n_spl_,
    g1177_n_spl_
  );


  or

  (
    g1179_n,
    g1178_p_spl_,
    g1177_p_spl_
  );


  and

  (
    g1180_p,
    g1179_n_spl_0,
    g1177_n_spl_
  );


  or

  (
    g1180_n,
    g1179_p_spl_0,
    g1177_p_spl_
  );


  and

  (
    g1181_p,
    g1179_n_spl_0,
    g1178_n_spl_
  );


  or

  (
    g1181_n,
    g1179_p_spl_0,
    g1178_p_spl_
  );


  and

  (
    g1182_p,
    g1181_n,
    g1180_n
  );


  or

  (
    g1182_n,
    g1181_p,
    g1180_p
  );


  and

  (
    g1183_p,
    n6205_o2_p_spl_0,
    n2848_lo_p_spl_10
  );


  or

  (
    g1183_n,
    n6205_o2_n_spl_0,
    n2848_lo_n_spl_10
  );


  and

  (
    g1184_p,
    g1183_n_spl_,
    g1182_n_spl_
  );


  or

  (
    g1184_n,
    g1183_p_spl_,
    g1182_p_spl_
  );


  and

  (
    g1185_p,
    g1184_n_spl_0,
    g1179_n_spl_
  );


  or

  (
    g1185_n,
    g1184_p_spl_0,
    g1179_p_spl_
  );


  and

  (
    g1186_p,
    g1185_n_spl_,
    g1174_n_spl_
  );


  or

  (
    g1186_n,
    g1185_p_spl_,
    g1174_p_spl_
  );


  and

  (
    g1187_p,
    g1186_n_spl_0,
    g1174_n_spl_
  );


  or

  (
    g1187_n,
    g1186_p_spl_0,
    g1174_p_spl_
  );


  and

  (
    g1188_p,
    g1186_n_spl_0,
    g1185_n_spl_
  );


  or

  (
    g1188_n,
    g1186_p_spl_0,
    g1185_p_spl_
  );


  and

  (
    g1189_p,
    g1188_n,
    g1187_n
  );


  or

  (
    g1189_n,
    g1188_p,
    g1187_p
  );


  and

  (
    g1190_p,
    n6205_o2_p_spl_,
    n2860_lo_p_spl_01
  );


  or

  (
    g1190_n,
    n6205_o2_n_spl_,
    n2860_lo_n_spl_01
  );


  and

  (
    g1191_p,
    g1190_n_spl_,
    g1189_n_spl_
  );


  or

  (
    g1191_n,
    g1190_p_spl_,
    g1189_p_spl_
  );


  and

  (
    g1192_p,
    g1191_n_spl_0,
    g1189_n_spl_
  );


  or

  (
    g1192_n,
    g1191_p_spl_0,
    g1189_p_spl_
  );


  and

  (
    g1193_p,
    g1191_n_spl_0,
    g1190_n_spl_
  );


  or

  (
    g1193_n,
    g1191_p_spl_0,
    g1190_p_spl_
  );


  and

  (
    g1194_p,
    g1193_n,
    g1192_n
  );


  or

  (
    g1194_n,
    g1193_p,
    g1192_p
  );


  and

  (
    g1195_p,
    g1184_n_spl_0,
    g1182_n_spl_
  );


  or

  (
    g1195_n,
    g1184_p_spl_0,
    g1182_p_spl_
  );


  and

  (
    g1196_p,
    g1184_n_spl_,
    g1183_n_spl_
  );


  or

  (
    g1196_n,
    g1184_p_spl_,
    g1183_p_spl_
  );


  and

  (
    g1197_p,
    g1196_n,
    g1195_n
  );


  or

  (
    g1197_n,
    g1196_p,
    g1195_p
  );


  and

  (
    g1198_p,
    g1025_n_spl_,
    g1020_n_spl_
  );


  or

  (
    g1198_n,
    g1025_p_spl_,
    g1020_p_spl_
  );


  and

  (
    g1199_p,
    g1198_n_spl_,
    g1197_n_spl_
  );


  or

  (
    g1199_n,
    g1198_p_spl_,
    g1197_p_spl_
  );


  and

  (
    g1200_p,
    g1199_n_spl_0,
    g1197_n_spl_
  );


  or

  (
    g1200_n,
    g1199_p_spl_0,
    g1197_p_spl_
  );


  and

  (
    g1201_p,
    g1199_n_spl_0,
    g1198_n_spl_
  );


  or

  (
    g1201_n,
    g1199_p_spl_0,
    g1198_p_spl_
  );


  and

  (
    g1202_p,
    g1201_n,
    g1200_n
  );


  or

  (
    g1202_n,
    g1201_p,
    g1200_p
  );


  and

  (
    g1203_p,
    n6239_o2_p_spl_,
    n2860_lo_p_spl_01
  );


  or

  (
    g1203_n,
    n6239_o2_n_spl_,
    n2860_lo_n_spl_01
  );


  and

  (
    g1204_p,
    g1203_n_spl_,
    g1202_n_spl_
  );


  or

  (
    g1204_n,
    g1203_p_spl_,
    g1202_p_spl_
  );


  and

  (
    g1205_p,
    g1204_n_spl_0,
    g1199_n_spl_
  );


  or

  (
    g1205_n,
    g1204_p_spl_0,
    g1199_p_spl_
  );


  or

  (
    g1206_n,
    g1205_p,
    g1194_p
  );


  and

  (
    g1207_p,
    g1204_n_spl_0,
    g1202_n_spl_
  );


  or

  (
    g1207_n,
    g1204_p_spl_0,
    g1202_p_spl_
  );


  and

  (
    g1208_p,
    g1204_n_spl_,
    g1203_n_spl_
  );


  or

  (
    g1208_n,
    g1204_p_spl_,
    g1203_p_spl_
  );


  and

  (
    g1209_p,
    g1208_n,
    g1207_n
  );


  or

  (
    g1209_n,
    g1208_p,
    g1207_p
  );


  and

  (
    g1210_p,
    g1035_n_spl_,
    g1030_n_spl_
  );


  or

  (
    g1210_n,
    g1035_p_spl_,
    g1030_p_spl_
  );


  and

  (
    g1211_p,
    g1210_n_spl_,
    g1209_n_spl_
  );


  or

  (
    g1211_n,
    g1210_p,
    g1209_p
  );


  and

  (
    g1212_p,
    g1211_n_spl_,
    g1209_n_spl_
  );


  and

  (
    g1213_p,
    g1211_n_spl_,
    g1210_n_spl_
  );


  or

  (
    g1214_n,
    g1213_p,
    g1212_p
  );


  and

  (
    g1215_p,
    n2488_lo_buf_o2_p_spl_1,
    n2734_lo_p_spl_000
  );


  or

  (
    g1215_n,
    n2488_lo_buf_o2_n_spl_1,
    n2734_lo_n_spl_000
  );


  and

  (
    g1216_p,
    g1009_n_spl_0,
    g987_n_spl_
  );


  or

  (
    g1216_n,
    g1009_p_spl_,
    g987_p_spl_
  );


  and

  (
    g1217_p,
    g1009_n_spl_0,
    g1008_n_spl_
  );


  or

  (
    g1217_n,
    g1009_p_spl_,
    g1008_p_spl_
  );


  and

  (
    g1218_p,
    g1217_n,
    g1216_n
  );


  or

  (
    g1218_n,
    g1217_p,
    g1216_p
  );


  and

  (
    g1219_p,
    n6103_o2_p_spl_,
    n2860_lo_p_spl_10
  );


  or

  (
    g1219_n,
    n6103_o2_n_spl_,
    n2860_lo_n_spl_10
  );


  or

  (
    g1220_n,
    g1219_p,
    g1218_p
  );


  and

  (
    g1221_p,
    g935_n_spl_0,
    g913_n_spl_
  );


  or

  (
    g1221_n,
    g935_p_spl_,
    g913_p_spl_
  );


  and

  (
    g1222_p,
    g935_n_spl_0,
    g934_n_spl_
  );


  or

  (
    g1222_n,
    g935_p_spl_,
    g934_p_spl_
  );


  and

  (
    g1223_p,
    g1222_n,
    g1221_n
  );


  or

  (
    g1223_n,
    g1222_p,
    g1221_p
  );


  and

  (
    g1224_p,
    n5959_o2_p_spl_1,
    n2848_lo_p_spl_10
  );


  or

  (
    g1224_n,
    n5959_o2_n_spl_,
    n2848_lo_n_spl_10
  );


  or

  (
    g1225_n,
    g1224_p,
    g1223_p
  );


  and

  (
    g1226_p,
    g861_n_spl_0,
    g839_n_spl_
  );


  or

  (
    g1226_n,
    g861_p_spl_,
    g839_p_spl_
  );


  and

  (
    g1227_p,
    g861_n_spl_0,
    g860_n_spl_
  );


  or

  (
    g1227_n,
    g861_p_spl_,
    g860_p_spl_
  );


  and

  (
    g1228_p,
    g1227_n,
    g1226_n
  );


  or

  (
    g1228_n,
    g1227_p,
    g1226_p
  );


  and

  (
    g1229_p,
    n5842_o2_p_spl_1,
    n2836_lo_p_spl_110
  );


  or

  (
    g1229_n,
    n5842_o2_n_spl_,
    n2836_lo_n_spl_110
  );


  or

  (
    g1230_n,
    g1229_p,
    g1228_p
  );


  and

  (
    g1231_p,
    g1214_n_spl_,
    g1098_n_spl_
  );


  and

  (
    g1232_p,
    n2764_lo_buf_o2_p_spl_0,
    n7148_o2_p_spl_0
  );


  or

  (
    g1232_n,
    n2764_lo_buf_o2_n_spl_0,
    n7148_o2_n_spl_0
  );


  and

  (
    g1233_p,
    G2917_o2_n_spl_,
    G1280_o2_n_spl_
  );


  or

  (
    g1233_n,
    G2917_o2_p_spl_,
    G1280_o2_p_spl_
  );


  and

  (
    g1234_p,
    g1233_n_spl_0,
    G1280_o2_n_spl_
  );


  or

  (
    g1234_n,
    g1233_p_spl_0,
    G1280_o2_p_spl_
  );


  and

  (
    g1235_p,
    g1233_n_spl_0,
    G2917_o2_n_spl_
  );


  or

  (
    g1235_n,
    g1233_p_spl_0,
    G2917_o2_p_spl_
  );


  and

  (
    g1236_p,
    g1235_n,
    g1234_n
  );


  or

  (
    g1236_n,
    g1235_p,
    g1234_p
  );


  and

  (
    g1237_p,
    n2764_lo_buf_o2_p_spl_1,
    n7224_o2_p_spl_0
  );


  or

  (
    g1237_n,
    n2764_lo_buf_o2_n_spl_1,
    n7224_o2_n_spl_0
  );


  and

  (
    g1238_p,
    g1237_n_spl_,
    g1236_n_spl_
  );


  or

  (
    g1238_n,
    g1237_p_spl_,
    g1236_p_spl_
  );


  and

  (
    g1239_p,
    g1238_n_spl_0,
    g1233_n_spl_
  );


  or

  (
    g1239_n,
    g1238_p_spl_0,
    g1233_p_spl_
  );


  and

  (
    g1240_p,
    g1239_n_spl_,
    g1232_n_spl_
  );


  or

  (
    g1240_n,
    g1239_p_spl_,
    g1232_p_spl_
  );


  and

  (
    g1241_p,
    g1240_n_spl_0,
    g1232_n_spl_
  );


  or

  (
    g1241_n,
    g1240_p_spl_0,
    g1232_p_spl_
  );


  and

  (
    g1242_p,
    g1240_n_spl_0,
    g1239_n_spl_
  );


  or

  (
    g1242_n,
    g1240_p_spl_0,
    g1239_p_spl_
  );


  and

  (
    g1243_p,
    g1242_n,
    g1241_n
  );


  or

  (
    g1243_n,
    g1242_p,
    g1241_p
  );


  and

  (
    g1244_p,
    n2776_lo_buf_o2_p_spl_001,
    n7224_o2_p_spl_0
  );


  or

  (
    g1244_n,
    n2776_lo_buf_o2_n_spl_001,
    n7224_o2_n_spl_0
  );


  and

  (
    g1245_p,
    g1244_n_spl_,
    g1243_n_spl_
  );


  or

  (
    g1245_n,
    g1244_p_spl_,
    g1243_p_spl_
  );


  and

  (
    g1246_p,
    g1245_n_spl_0,
    g1243_n_spl_
  );


  or

  (
    g1246_n,
    g1245_p_spl_0,
    g1243_p_spl_
  );


  and

  (
    g1247_p,
    g1245_n_spl_0,
    g1244_n_spl_
  );


  or

  (
    g1247_n,
    g1245_p_spl_0,
    g1244_p_spl_
  );


  and

  (
    g1248_p,
    g1247_n,
    g1246_n
  );


  or

  (
    g1248_n,
    g1247_p,
    g1246_p
  );


  and

  (
    g1249_p,
    g1238_n_spl_0,
    g1236_n_spl_
  );


  or

  (
    g1249_n,
    g1238_p_spl_0,
    g1236_p_spl_
  );


  and

  (
    g1250_p,
    g1238_n_spl_,
    g1237_n_spl_
  );


  or

  (
    g1250_n,
    g1238_p_spl_,
    g1237_p_spl_
  );


  and

  (
    g1251_p,
    g1250_n,
    g1249_n
  );


  or

  (
    g1251_n,
    g1250_p,
    g1249_p
  );


  and

  (
    g1252_p,
    G3068_o2_n,
    G3069_o2_n
  );


  or

  (
    g1252_n,
    G3068_o2_p,
    G3069_o2_p
  );


  and

  (
    g1253_p,
    n2764_lo_buf_o2_p_spl_1,
    n7280_o2_p_spl_0
  );


  or

  (
    g1253_n,
    n2764_lo_buf_o2_n_spl_1,
    n7280_o2_n_spl_0
  );


  and

  (
    g1254_p,
    g1253_n_spl_,
    g1252_n_spl_
  );


  or

  (
    g1254_n,
    g1253_p_spl_,
    g1252_p_spl_
  );


  and

  (
    g1255_p,
    g1254_n_spl_0,
    G3016_o2_p
  );


  or

  (
    g1255_n,
    g1254_p_spl_0,
    G3016_o2_n
  );


  and

  (
    g1256_p,
    g1255_n_spl_,
    g1251_n_spl_
  );


  or

  (
    g1256_n,
    g1255_p_spl_,
    g1251_p_spl_
  );


  and

  (
    g1257_p,
    g1256_n_spl_0,
    g1251_n_spl_
  );


  or

  (
    g1257_n,
    g1256_p_spl_0,
    g1251_p_spl_
  );


  and

  (
    g1258_p,
    g1256_n_spl_0,
    g1255_n_spl_
  );


  or

  (
    g1258_n,
    g1256_p_spl_0,
    g1255_p_spl_
  );


  and

  (
    g1259_p,
    g1258_n,
    g1257_n
  );


  or

  (
    g1259_n,
    g1258_p,
    g1257_p
  );


  and

  (
    g1260_p,
    n2776_lo_buf_o2_p_spl_010,
    n7280_o2_p_spl_0
  );


  or

  (
    g1260_n,
    n2776_lo_buf_o2_n_spl_010,
    n7280_o2_n_spl_0
  );


  and

  (
    g1261_p,
    g1260_n_spl_,
    g1259_n_spl_
  );


  or

  (
    g1261_n,
    g1260_p_spl_,
    g1259_p_spl_
  );


  and

  (
    g1262_p,
    g1261_n_spl_0,
    g1256_n_spl_
  );


  or

  (
    g1262_n,
    g1261_p_spl_0,
    g1256_p_spl_
  );


  and

  (
    g1263_p,
    g1262_n_spl_,
    g1248_n_spl_
  );


  or

  (
    g1263_n,
    g1262_p_spl_,
    g1248_p_spl_
  );


  and

  (
    g1264_p,
    g1263_n_spl_0,
    g1248_n_spl_
  );


  or

  (
    g1264_n,
    g1263_p_spl_0,
    g1248_p_spl_
  );


  and

  (
    g1265_p,
    g1263_n_spl_0,
    g1262_n_spl_
  );


  or

  (
    g1265_n,
    g1263_p_spl_0,
    g1262_p_spl_
  );


  and

  (
    g1266_p,
    g1265_n,
    g1264_n
  );


  or

  (
    g1266_n,
    g1265_p,
    g1264_p
  );


  and

  (
    g1267_p,
    n7280_o2_p_spl_1,
    n2785_lo_p_spl_001
  );


  or

  (
    g1267_n,
    n7280_o2_n_spl_1,
    n2785_lo_n_spl_001
  );


  and

  (
    g1268_p,
    g1267_n_spl_,
    g1266_n_spl_
  );


  or

  (
    g1268_n,
    g1267_p_spl_,
    g1266_p_spl_
  );


  and

  (
    g1269_p,
    g1268_n_spl_0,
    g1266_n_spl_
  );


  or

  (
    g1269_n,
    g1268_p_spl_0,
    g1266_p_spl_
  );


  and

  (
    g1270_p,
    g1268_n_spl_0,
    g1267_n_spl_
  );


  or

  (
    g1270_n,
    g1268_p_spl_0,
    g1267_p_spl_
  );


  and

  (
    g1271_p,
    g1270_n,
    g1269_n
  );


  or

  (
    g1271_n,
    g1270_p,
    g1269_p
  );


  and

  (
    g1272_p,
    g1261_n_spl_0,
    g1259_n_spl_
  );


  or

  (
    g1272_n,
    g1261_p_spl_0,
    g1259_p_spl_
  );


  and

  (
    g1273_p,
    g1261_n_spl_,
    g1260_n_spl_
  );


  or

  (
    g1273_n,
    g1261_p_spl_,
    g1260_p_spl_
  );


  and

  (
    g1274_p,
    g1273_n,
    g1272_n
  );


  or

  (
    g1274_n,
    g1273_p,
    g1272_p
  );


  and

  (
    g1275_p,
    g1254_n_spl_0,
    g1252_n_spl_
  );


  or

  (
    g1275_n,
    g1254_p_spl_0,
    g1252_p_spl_
  );


  and

  (
    g1276_p,
    g1254_n_spl_,
    g1253_n_spl_
  );


  or

  (
    g1276_n,
    g1254_p_spl_,
    g1253_p_spl_
  );


  and

  (
    g1277_p,
    g1276_n,
    g1275_n
  );


  or

  (
    g1277_n,
    g1276_p,
    g1275_p
  );


  and

  (
    g1278_p,
    G3241_o2_n_spl_0,
    G3064_o2_p
  );


  or

  (
    g1278_n,
    G3241_o2_p_spl_0,
    G3064_o2_n
  );


  and

  (
    g1279_p,
    g1278_n_spl_,
    g1277_n_spl_
  );


  or

  (
    g1279_n,
    g1278_p_spl_,
    g1277_p_spl_
  );


  and

  (
    g1280_p,
    g1279_n_spl_0,
    g1277_n_spl_
  );


  or

  (
    g1280_n,
    g1279_p_spl_0,
    g1277_p_spl_
  );


  and

  (
    g1281_p,
    g1279_n_spl_0,
    g1278_n_spl_
  );


  or

  (
    g1281_n,
    g1279_p_spl_0,
    g1278_p_spl_
  );


  and

  (
    g1282_p,
    g1281_n,
    g1280_n
  );


  or

  (
    g1282_n,
    g1281_p,
    g1280_p
  );


  and

  (
    g1283_p,
    n2776_lo_buf_o2_p_spl_010,
    n7313_o2_p_spl_0
  );


  or

  (
    g1283_n,
    n2776_lo_buf_o2_n_spl_010,
    n7313_o2_n_spl_0
  );


  and

  (
    g1284_p,
    g1283_n_spl_,
    g1282_n_spl_
  );


  or

  (
    g1284_n,
    g1283_p_spl_,
    g1282_p_spl_
  );


  and

  (
    g1285_p,
    g1284_n_spl_0,
    g1279_n_spl_
  );


  or

  (
    g1285_n,
    g1284_p_spl_0,
    g1279_p_spl_
  );


  and

  (
    g1286_p,
    g1285_n_spl_,
    g1274_n_spl_
  );


  or

  (
    g1286_n,
    g1285_p_spl_,
    g1274_p_spl_
  );


  and

  (
    g1287_p,
    g1286_n_spl_0,
    g1274_n_spl_
  );


  or

  (
    g1287_n,
    g1286_p_spl_0,
    g1274_p_spl_
  );


  and

  (
    g1288_p,
    g1286_n_spl_0,
    g1285_n_spl_
  );


  or

  (
    g1288_n,
    g1286_p_spl_0,
    g1285_p_spl_
  );


  and

  (
    g1289_p,
    g1288_n,
    g1287_n
  );


  or

  (
    g1289_n,
    g1288_p,
    g1287_p
  );


  and

  (
    g1290_p,
    n7313_o2_p_spl_0,
    n2785_lo_p_spl_001
  );


  or

  (
    g1290_n,
    n7313_o2_n_spl_0,
    n2785_lo_n_spl_001
  );


  and

  (
    g1291_p,
    g1290_n_spl_,
    g1289_n_spl_
  );


  or

  (
    g1291_n,
    g1290_p_spl_,
    g1289_p_spl_
  );


  and

  (
    g1292_p,
    g1291_n_spl_0,
    g1286_n_spl_
  );


  or

  (
    g1292_n,
    g1291_p_spl_0,
    g1286_p_spl_
  );


  and

  (
    g1293_p,
    g1292_n_spl_,
    g1271_n_spl_
  );


  or

  (
    g1293_n,
    g1292_p_spl_,
    g1271_p_spl_
  );


  and

  (
    g1294_p,
    G3241_o2_n_spl_0,
    G3193_o2_p
  );


  or

  (
    g1294_n,
    G3241_o2_p_spl_0,
    G3193_o2_n
  );


  and

  (
    g1295_p,
    G3241_o2_n_spl_,
    G1139_o2_n
  );


  or

  (
    g1295_n,
    G3241_o2_p_spl_,
    G1139_o2_p
  );


  and

  (
    g1296_p,
    g1295_n,
    g1294_n
  );


  or

  (
    g1296_n,
    g1295_p,
    g1294_p
  );


  and

  (
    g1297_p,
    G3298_o2_n,
    G3121_o2_p
  );


  or

  (
    g1297_n,
    G3298_o2_p,
    G3121_o2_n
  );


  and

  (
    g1298_p,
    g1297_n_spl_,
    g1296_n_spl_
  );


  or

  (
    g1298_n,
    g1297_p_spl_,
    g1296_p_spl_
  );


  and

  (
    g1299_p,
    g1298_n_spl_0,
    g1296_n_spl_
  );


  or

  (
    g1299_n,
    g1298_p_spl_0,
    g1296_p_spl_
  );


  and

  (
    g1300_p,
    g1298_n_spl_0,
    g1297_n_spl_
  );


  or

  (
    g1300_n,
    g1298_p_spl_0,
    g1297_p_spl_
  );


  and

  (
    g1301_p,
    g1300_n,
    g1299_n
  );


  or

  (
    g1301_n,
    g1300_p,
    g1299_p
  );


  and

  (
    g1302_p,
    n2776_lo_buf_o2_p_spl_011,
    n7323_o2_p_spl_0
  );


  or

  (
    g1302_n,
    n2776_lo_buf_o2_n_spl_011,
    n7323_o2_n_spl_0
  );


  and

  (
    g1303_p,
    g1302_n_spl_,
    g1301_n_spl_
  );


  or

  (
    g1303_n,
    g1302_p_spl_,
    g1301_p_spl_
  );


  and

  (
    g1304_p,
    g1303_n_spl_0,
    g1301_n_spl_
  );


  or

  (
    g1304_n,
    g1303_p_spl_0,
    g1301_p_spl_
  );


  and

  (
    g1305_p,
    g1303_n_spl_0,
    g1302_n_spl_
  );


  or

  (
    g1305_n,
    g1303_p_spl_0,
    g1302_p_spl_
  );


  and

  (
    g1306_p,
    g1305_n,
    g1304_n
  );


  or

  (
    g1306_n,
    g1305_p,
    g1304_p
  );


  and

  (
    g1307_p,
    G3394_o2_n_spl_,
    G3391_o2_n_spl_
  );


  or

  (
    g1307_n,
    G3394_o2_p_spl_,
    G3391_o2_p_spl_
  );


  and

  (
    g1308_p,
    g1307_n_spl_0,
    G3394_o2_n_spl_
  );


  or

  (
    g1308_n,
    g1307_p_spl_0,
    G3394_o2_p_spl_
  );


  and

  (
    g1309_p,
    g1307_n_spl_0,
    G3391_o2_n_spl_
  );


  or

  (
    g1309_n,
    g1307_p_spl_0,
    G3391_o2_p_spl_
  );


  and

  (
    g1310_p,
    g1309_n,
    g1308_n
  );


  or

  (
    g1310_n,
    g1309_p,
    g1308_p
  );


  and

  (
    g1311_p,
    n2776_lo_buf_o2_p_spl_011,
    n7398_o2_p_spl_0
  );


  or

  (
    g1311_n,
    n2776_lo_buf_o2_n_spl_011,
    n7398_o2_n_spl_0
  );


  and

  (
    g1312_p,
    g1311_n_spl_,
    g1310_n_spl_
  );


  or

  (
    g1312_n,
    g1311_p_spl_,
    g1310_p_spl_
  );


  and

  (
    g1313_p,
    g1312_n_spl_0,
    g1307_n_spl_
  );


  or

  (
    g1313_n,
    g1312_p_spl_0,
    g1307_p_spl_
  );


  and

  (
    g1314_p,
    g1313_n_spl_,
    g1306_n_spl_
  );


  or

  (
    g1314_n,
    g1313_p_spl_,
    g1306_p_spl_
  );


  and

  (
    g1315_p,
    g1314_n_spl_0,
    g1306_n_spl_
  );


  or

  (
    g1315_n,
    g1314_p_spl_0,
    g1306_p_spl_
  );


  and

  (
    g1316_p,
    g1314_n_spl_0,
    g1313_n_spl_
  );


  or

  (
    g1316_n,
    g1314_p_spl_0,
    g1313_p_spl_
  );


  and

  (
    g1317_p,
    g1316_n,
    g1315_n
  );


  or

  (
    g1317_n,
    g1316_p,
    g1315_p
  );


  and

  (
    g1318_p,
    n7398_o2_p_spl_0,
    n2785_lo_p_spl_010
  );


  or

  (
    g1318_n,
    n7398_o2_n_spl_0,
    n2785_lo_n_spl_010
  );


  and

  (
    g1319_p,
    g1318_n_spl_,
    g1317_n_spl_
  );


  or

  (
    g1319_n,
    g1318_p_spl_,
    g1317_p_spl_
  );


  and

  (
    g1320_p,
    g1319_n_spl_0,
    g1317_n_spl_
  );


  or

  (
    g1320_n,
    g1319_p_spl_0,
    g1317_p_spl_
  );


  and

  (
    g1321_p,
    g1319_n_spl_0,
    g1318_n_spl_
  );


  or

  (
    g1321_n,
    g1319_p_spl_0,
    g1318_p_spl_
  );


  and

  (
    g1322_p,
    g1321_n,
    g1320_n
  );


  or

  (
    g1322_n,
    g1321_p,
    g1320_p
  );


  and

  (
    g1323_p,
    g1312_n_spl_0,
    g1310_n_spl_
  );


  or

  (
    g1323_n,
    g1312_p_spl_0,
    g1310_p_spl_
  );


  and

  (
    g1324_p,
    g1312_n_spl_,
    g1311_n_spl_
  );


  or

  (
    g1324_n,
    g1312_p_spl_,
    g1311_p_spl_
  );


  and

  (
    g1325_p,
    g1324_n,
    g1323_n
  );


  or

  (
    g1325_n,
    g1324_p,
    g1323_p
  );


  and

  (
    g1326_p,
    G3573_o2_n,
    G3574_o2_n
  );


  or

  (
    g1326_n,
    G3573_o2_p,
    G3574_o2_p
  );


  and

  (
    g1327_p,
    n2776_lo_buf_o2_p_spl_100,
    n7459_o2_p_spl_0
  );


  or

  (
    g1327_n,
    n2776_lo_buf_o2_n_spl_100,
    n7459_o2_n_spl_0
  );


  and

  (
    g1328_p,
    g1327_n_spl_,
    g1326_n_spl_
  );


  or

  (
    g1328_n,
    g1327_p_spl_,
    g1326_p_spl_
  );


  and

  (
    g1329_p,
    g1328_n_spl_0,
    G3520_o2_p
  );


  or

  (
    g1329_n,
    g1328_p_spl_0,
    G3520_o2_n
  );


  and

  (
    g1330_p,
    g1329_n_spl_,
    g1325_n_spl_
  );


  or

  (
    g1330_n,
    g1329_p_spl_,
    g1325_p_spl_
  );


  and

  (
    g1331_p,
    g1330_n_spl_0,
    g1325_n_spl_
  );


  or

  (
    g1331_n,
    g1330_p_spl_0,
    g1325_p_spl_
  );


  and

  (
    g1332_p,
    g1330_n_spl_0,
    g1329_n_spl_
  );


  or

  (
    g1332_n,
    g1330_p_spl_0,
    g1329_p_spl_
  );


  and

  (
    g1333_p,
    g1332_n,
    g1331_n
  );


  or

  (
    g1333_n,
    g1332_p,
    g1331_p
  );


  and

  (
    g1334_p,
    n7459_o2_p_spl_0,
    n2785_lo_p_spl_010
  );


  or

  (
    g1334_n,
    n7459_o2_n_spl_0,
    n2785_lo_n_spl_010
  );


  and

  (
    g1335_p,
    g1334_n_spl_,
    g1333_n_spl_
  );


  or

  (
    g1335_n,
    g1334_p_spl_,
    g1333_p_spl_
  );


  and

  (
    g1336_p,
    g1335_n_spl_0,
    g1330_n_spl_
  );


  or

  (
    g1336_n,
    g1335_p_spl_0,
    g1330_p_spl_
  );


  and

  (
    g1337_p,
    g1336_n_spl_,
    g1322_n_spl_
  );


  or

  (
    g1337_n,
    g1336_p_spl_,
    g1322_p_spl_
  );


  and

  (
    g1338_p,
    g1337_n_spl_0,
    g1322_n_spl_
  );


  or

  (
    g1338_n,
    g1337_p_spl_0,
    g1322_p_spl_
  );


  and

  (
    g1339_p,
    g1337_n_spl_0,
    g1336_n_spl_
  );


  or

  (
    g1339_n,
    g1337_p_spl_0,
    g1336_p_spl_
  );


  and

  (
    g1340_p,
    g1339_n,
    g1338_n
  );


  or

  (
    g1340_n,
    g1339_p,
    g1338_p
  );


  and

  (
    g1341_p,
    n7459_o2_p_spl_1,
    n2797_lo_p_spl_000
  );


  or

  (
    g1341_n,
    n7459_o2_n_spl_1,
    n2797_lo_n_spl_000
  );


  and

  (
    g1342_p,
    g1341_n_spl_,
    g1340_n_spl_
  );


  or

  (
    g1342_n,
    g1341_p_spl_,
    g1340_p_spl_
  );


  and

  (
    g1343_p,
    g1342_n_spl_0,
    g1340_n_spl_
  );


  or

  (
    g1343_n,
    g1342_p_spl_0,
    g1340_p_spl_
  );


  and

  (
    g1344_p,
    g1342_n_spl_0,
    g1341_n_spl_
  );


  or

  (
    g1344_n,
    g1342_p_spl_0,
    g1341_p_spl_
  );


  and

  (
    g1345_p,
    g1344_n,
    g1343_n
  );


  or

  (
    g1345_n,
    g1344_p,
    g1343_p
  );


  and

  (
    g1346_p,
    g1335_n_spl_0,
    g1333_n_spl_
  );


  or

  (
    g1346_n,
    g1335_p_spl_0,
    g1333_p_spl_
  );


  and

  (
    g1347_p,
    g1335_n_spl_,
    g1334_n_spl_
  );


  or

  (
    g1347_n,
    g1335_p_spl_,
    g1334_p_spl_
  );


  and

  (
    g1348_p,
    g1347_n,
    g1346_n
  );


  or

  (
    g1348_n,
    g1347_p,
    g1346_p
  );


  and

  (
    g1349_p,
    g1328_n_spl_0,
    g1326_n_spl_
  );


  or

  (
    g1349_n,
    g1328_p_spl_0,
    g1326_p_spl_
  );


  and

  (
    g1350_p,
    g1328_n_spl_,
    g1327_n_spl_
  );


  or

  (
    g1350_n,
    g1328_p_spl_,
    g1327_p_spl_
  );


  and

  (
    g1351_p,
    g1350_n,
    g1349_n
  );


  or

  (
    g1351_n,
    g1350_p,
    g1349_p
  );


  and

  (
    g1352_p,
    G3722_o2_n_spl_0,
    G3569_o2_p
  );


  or

  (
    g1352_n,
    G3722_o2_p_spl_0,
    G3569_o2_n
  );


  and

  (
    g1353_p,
    g1352_n_spl_,
    g1351_n_spl_
  );


  or

  (
    g1353_n,
    g1352_p_spl_,
    g1351_p_spl_
  );


  and

  (
    g1354_p,
    g1353_n_spl_0,
    g1351_n_spl_
  );


  or

  (
    g1354_n,
    g1353_p_spl_0,
    g1351_p_spl_
  );


  and

  (
    g1355_p,
    g1353_n_spl_0,
    g1352_n_spl_
  );


  or

  (
    g1355_n,
    g1353_p_spl_0,
    g1352_p_spl_
  );


  and

  (
    g1356_p,
    g1355_n,
    g1354_n
  );


  or

  (
    g1356_n,
    g1355_p,
    g1354_p
  );


  and

  (
    g1357_p,
    n7501_o2_p_spl_0,
    n2785_lo_p_spl_011
  );


  or

  (
    g1357_n,
    n7501_o2_n_spl_0,
    n2785_lo_n_spl_011
  );


  and

  (
    g1358_p,
    g1357_n_spl_,
    g1356_n_spl_
  );


  or

  (
    g1358_n,
    g1357_p_spl_,
    g1356_p_spl_
  );


  and

  (
    g1359_p,
    g1358_n_spl_0,
    g1353_n_spl_
  );


  or

  (
    g1359_n,
    g1358_p_spl_0,
    g1353_p_spl_
  );


  and

  (
    g1360_p,
    g1359_n_spl_,
    g1348_n_spl_
  );


  or

  (
    g1360_n,
    g1359_p_spl_,
    g1348_p_spl_
  );


  and

  (
    g1361_p,
    g1360_n_spl_0,
    g1348_n_spl_
  );


  or

  (
    g1361_n,
    g1360_p_spl_0,
    g1348_p_spl_
  );


  and

  (
    g1362_p,
    g1360_n_spl_0,
    g1359_n_spl_
  );


  or

  (
    g1362_n,
    g1360_p_spl_0,
    g1359_p_spl_
  );


  and

  (
    g1363_p,
    g1362_n,
    g1361_n
  );


  or

  (
    g1363_n,
    g1362_p,
    g1361_p
  );


  and

  (
    g1364_p,
    n7501_o2_p_spl_0,
    n2797_lo_p_spl_001
  );


  or

  (
    g1364_n,
    n7501_o2_n_spl_0,
    n2797_lo_n_spl_001
  );


  and

  (
    g1365_p,
    g1364_n_spl_,
    g1363_n_spl_
  );


  or

  (
    g1365_n,
    g1364_p_spl_,
    g1363_p_spl_
  );


  and

  (
    g1366_p,
    g1365_n_spl_0,
    g1360_n_spl_
  );


  or

  (
    g1366_n,
    g1365_p_spl_0,
    g1360_p_spl_
  );


  and

  (
    g1367_p,
    g1366_n_spl_,
    g1345_n_spl_
  );


  or

  (
    g1367_n,
    g1366_p_spl_,
    g1345_p_spl_
  );


  and

  (
    g1368_p,
    G3722_o2_n_spl_0,
    G3670_o2_p
  );


  or

  (
    g1368_n,
    G3722_o2_p_spl_0,
    G3670_o2_n
  );


  and

  (
    g1369_p,
    G3722_o2_n_spl_,
    G950_o2_n
  );


  or

  (
    g1369_n,
    G3722_o2_p_spl_,
    G950_o2_p
  );


  and

  (
    g1370_p,
    g1369_n,
    g1368_n
  );


  or

  (
    g1370_n,
    g1369_p,
    g1368_p
  );


  and

  (
    g1371_p,
    G3719_o2_p_spl_,
    G902_o2_n_spl_
  );


  or

  (
    g1371_n,
    G3719_o2_n_spl_,
    G902_o2_p_spl_
  );


  and

  (
    g1372_p,
    g1371_n_spl_0,
    G3624_o2_p
  );


  or

  (
    g1372_n,
    g1371_p_spl_0,
    G3624_o2_n
  );


  and

  (
    g1373_p,
    g1372_n_spl_,
    g1370_n_spl_
  );


  or

  (
    g1373_n,
    g1372_p_spl_,
    g1370_p_spl_
  );


  and

  (
    g1374_p,
    g1373_n_spl_0,
    g1370_n_spl_
  );


  or

  (
    g1374_n,
    g1373_p_spl_0,
    g1370_p_spl_
  );


  and

  (
    g1375_p,
    g1373_n_spl_0,
    g1372_n_spl_
  );


  or

  (
    g1375_n,
    g1373_p_spl_0,
    g1372_p_spl_
  );


  and

  (
    g1376_p,
    g1375_n,
    g1374_n
  );


  or

  (
    g1376_n,
    g1375_p,
    g1374_p
  );


  and

  (
    g1377_p,
    n7518_o2_p_spl_0,
    n2785_lo_p_spl_011
  );


  or

  (
    g1377_n,
    n7518_o2_n_spl_0,
    n2785_lo_n_spl_011
  );


  and

  (
    g1378_p,
    g1377_n_spl_,
    g1376_n_spl_
  );


  or

  (
    g1378_n,
    g1377_p_spl_,
    g1376_p_spl_
  );


  and

  (
    g1379_p,
    g1378_n_spl_0,
    g1376_n_spl_
  );


  or

  (
    g1379_n,
    g1378_p_spl_0,
    g1376_p_spl_
  );


  and

  (
    g1380_p,
    g1378_n_spl_0,
    g1377_n_spl_
  );


  or

  (
    g1380_n,
    g1378_p_spl_0,
    g1377_p_spl_
  );


  and

  (
    g1381_p,
    g1380_n,
    g1379_n
  );


  or

  (
    g1381_n,
    g1380_p,
    g1379_p
  );


  and

  (
    g1382_p,
    g1371_n_spl_0,
    G3719_o2_p_spl_
  );


  or

  (
    g1382_n,
    g1371_p_spl_0,
    G3719_o2_n_spl_
  );


  and

  (
    g1383_p,
    g1371_n_spl_,
    G902_o2_n_spl_
  );


  or

  (
    g1383_n,
    g1371_p_spl_,
    G902_o2_p_spl_
  );


  and

  (
    g1384_p,
    g1383_n,
    g1382_n
  );


  or

  (
    g1384_n,
    g1383_p,
    g1382_p
  );


  and

  (
    g1385_p,
    G3666_o2_n,
    G3667_o2_n
  );


  or

  (
    g1385_n,
    G3666_o2_p,
    G3667_o2_p
  );


  and

  (
    g1386_p,
    n2776_lo_buf_o2_p_spl_100,
    n7606_o2_p_spl_00
  );


  or

  (
    g1386_n,
    n2776_lo_buf_o2_n_spl_100,
    n7606_o2_n_spl_0
  );


  and

  (
    g1387_p,
    g1386_n_spl_,
    g1385_n_spl_
  );


  or

  (
    g1387_n,
    g1386_p_spl_,
    g1385_p_spl_
  );


  and

  (
    g1388_p,
    g1387_n_spl_0,
    G3620_o2_p
  );


  or

  (
    g1388_n,
    g1387_p_spl_0,
    G3620_o2_n
  );


  and

  (
    g1389_p,
    g1388_n_spl_,
    g1384_n_spl_
  );


  or

  (
    g1389_n,
    g1388_p_spl_,
    g1384_p_spl_
  );


  and

  (
    g1390_p,
    g1389_n_spl_0,
    g1384_n_spl_
  );


  or

  (
    g1390_n,
    g1389_p_spl_0,
    g1384_p_spl_
  );


  and

  (
    g1391_p,
    g1389_n_spl_0,
    g1388_n_spl_
  );


  or

  (
    g1391_n,
    g1389_p_spl_0,
    g1388_p_spl_
  );


  and

  (
    g1392_p,
    g1391_n,
    g1390_n
  );


  or

  (
    g1392_n,
    g1391_p,
    g1390_p
  );


  and

  (
    g1393_p,
    n7606_o2_p_spl_00,
    n2785_lo_p_spl_100
  );


  or

  (
    g1393_n,
    n7606_o2_n_spl_0,
    n2785_lo_n_spl_100
  );


  and

  (
    g1394_p,
    g1393_n_spl_,
    g1392_n_spl_
  );


  or

  (
    g1394_n,
    g1393_p_spl_,
    g1392_p_spl_
  );


  and

  (
    g1395_p,
    g1394_n_spl_0,
    g1389_n_spl_
  );


  or

  (
    g1395_n,
    g1394_p_spl_0,
    g1389_p_spl_
  );


  and

  (
    g1396_p,
    g1395_n_spl_,
    g1381_n_spl_
  );


  or

  (
    g1396_n,
    g1395_p_spl_,
    g1381_p_spl_
  );


  and

  (
    g1397_p,
    g1396_n_spl_0,
    g1381_n_spl_
  );


  or

  (
    g1397_n,
    g1396_p_spl_0,
    g1381_p_spl_
  );


  and

  (
    g1398_p,
    g1396_n_spl_0,
    g1395_n_spl_
  );


  or

  (
    g1398_n,
    g1396_p_spl_0,
    g1395_p_spl_
  );


  and

  (
    g1399_p,
    g1398_n,
    g1397_n
  );


  or

  (
    g1399_n,
    g1398_p,
    g1397_p
  );


  and

  (
    g1400_p,
    n7606_o2_p_spl_0,
    n2797_lo_p_spl_001
  );


  or

  (
    g1400_n,
    n7606_o2_n_spl_1,
    n2797_lo_n_spl_001
  );


  and

  (
    g1401_p,
    g1400_n_spl_,
    g1399_n_spl_
  );


  or

  (
    g1401_n,
    g1400_p_spl_,
    g1399_p_spl_
  );


  and

  (
    g1402_p,
    g1401_n_spl_0,
    g1399_n_spl_
  );


  or

  (
    g1402_n,
    g1401_p_spl_0,
    g1399_p_spl_
  );


  and

  (
    g1403_p,
    g1401_n_spl_0,
    g1400_n_spl_
  );


  or

  (
    g1403_n,
    g1401_p_spl_0,
    g1400_p_spl_
  );


  and

  (
    g1404_p,
    g1403_n,
    g1402_n
  );


  or

  (
    g1404_n,
    g1403_p,
    g1402_p
  );


  and

  (
    g1405_p,
    g1394_n_spl_0,
    g1392_n_spl_
  );


  or

  (
    g1405_n,
    g1394_p_spl_0,
    g1392_p_spl_
  );


  and

  (
    g1406_p,
    g1394_n_spl_,
    g1393_n_spl_
  );


  or

  (
    g1406_n,
    g1394_p_spl_,
    g1393_p_spl_
  );


  and

  (
    g1407_p,
    g1406_n,
    g1405_n
  );


  or

  (
    g1407_n,
    g1406_p,
    g1405_p
  );


  and

  (
    g1408_p,
    g1387_n_spl_0,
    g1385_n_spl_
  );


  or

  (
    g1408_n,
    g1387_p_spl_0,
    g1385_p_spl_
  );


  and

  (
    g1409_p,
    g1387_n_spl_,
    g1386_n_spl_
  );


  or

  (
    g1409_n,
    g1387_p_spl_,
    g1386_p_spl_
  );


  and

  (
    g1410_p,
    g1409_n,
    g1408_n
  );


  or

  (
    g1410_n,
    g1409_p,
    g1408_p
  );


  and

  (
    g1411_p,
    G3616_o2_p_spl_0,
    G3560_o2_n
  );


  or

  (
    g1411_n,
    G3616_o2_n_spl_0,
    G3560_o2_p
  );


  and

  (
    g1412_p,
    G3616_o2_p_spl_0,
    G3499_o2_n
  );


  or

  (
    g1412_n,
    G3616_o2_n_spl_0,
    G3499_o2_p
  );


  and

  (
    g1413_p,
    g1412_n,
    g1411_n
  );


  or

  (
    g1413_n,
    g1412_p,
    g1411_p
  );


  and

  (
    g1414_p,
    n2776_lo_buf_o2_p_spl_101,
    n7675_o2_p_spl_00
  );


  or

  (
    g1414_n,
    n2776_lo_buf_o2_n_spl_101,
    n7675_o2_n_spl_00
  );


  and

  (
    g1415_p,
    g1414_n_spl_,
    g1413_n_spl_
  );


  or

  (
    g1415_n,
    g1414_p_spl_,
    g1413_p_spl_
  );


  and

  (
    g1416_p,
    g1415_n_spl_0,
    G3616_o2_p_spl_
  );


  or

  (
    g1416_n,
    g1415_p_spl_0,
    G3616_o2_n_spl_
  );


  and

  (
    g1417_p,
    g1416_n_spl_,
    g1410_n_spl_
  );


  or

  (
    g1417_n,
    g1416_p_spl_,
    g1410_p_spl_
  );


  and

  (
    g1418_p,
    g1417_n_spl_0,
    g1410_n_spl_
  );


  or

  (
    g1418_n,
    g1417_p_spl_0,
    g1410_p_spl_
  );


  and

  (
    g1419_p,
    g1417_n_spl_0,
    g1416_n_spl_
  );


  or

  (
    g1419_n,
    g1417_p_spl_0,
    g1416_p_spl_
  );


  and

  (
    g1420_p,
    g1419_n,
    g1418_n
  );


  or

  (
    g1420_n,
    g1419_p,
    g1418_p
  );


  and

  (
    g1421_p,
    n7675_o2_p_spl_00,
    n2785_lo_p_spl_100
  );


  or

  (
    g1421_n,
    n7675_o2_n_spl_00,
    n2785_lo_n_spl_100
  );


  and

  (
    g1422_p,
    g1421_n_spl_,
    g1420_n_spl_
  );


  or

  (
    g1422_n,
    g1421_p_spl_,
    g1420_p_spl_
  );


  and

  (
    g1423_p,
    g1422_n_spl_0,
    g1417_n_spl_
  );


  or

  (
    g1423_n,
    g1422_p_spl_0,
    g1417_p_spl_
  );


  and

  (
    g1424_p,
    g1423_n_spl_,
    g1407_n_spl_
  );


  or

  (
    g1424_n,
    g1423_p_spl_,
    g1407_p_spl_
  );


  and

  (
    g1425_p,
    g1424_n_spl_0,
    g1407_n_spl_
  );


  or

  (
    g1425_n,
    g1424_p_spl_0,
    g1407_p_spl_
  );


  and

  (
    g1426_p,
    g1424_n_spl_0,
    g1423_n_spl_
  );


  or

  (
    g1426_n,
    g1424_p_spl_0,
    g1423_p_spl_
  );


  and

  (
    g1427_p,
    g1426_n,
    g1425_n
  );


  or

  (
    g1427_n,
    g1426_p,
    g1425_p
  );


  and

  (
    g1428_p,
    n7675_o2_p_spl_0,
    n2797_lo_p_spl_010
  );


  or

  (
    g1428_n,
    n7675_o2_n_spl_0,
    n2797_lo_n_spl_010
  );


  and

  (
    g1429_p,
    g1428_n_spl_,
    g1427_n_spl_
  );


  or

  (
    g1429_n,
    g1428_p_spl_,
    g1427_p_spl_
  );


  and

  (
    g1430_p,
    g1429_n_spl_0,
    g1424_n_spl_
  );


  or

  (
    g1430_n,
    g1429_p_spl_0,
    g1424_p_spl_
  );


  and

  (
    g1431_p,
    g1430_n_spl_,
    g1404_n_spl_
  );


  or

  (
    g1431_n,
    g1430_p_spl_,
    g1404_p_spl_
  );


  and

  (
    g1432_p,
    g1431_n_spl_0,
    g1404_n_spl_
  );


  or

  (
    g1432_n,
    g1431_p_spl_0,
    g1404_p_spl_
  );


  and

  (
    g1433_p,
    g1431_n_spl_0,
    g1430_n_spl_
  );


  or

  (
    g1433_n,
    g1431_p_spl_0,
    g1430_p_spl_
  );


  and

  (
    g1434_p,
    g1433_n,
    g1432_n
  );


  or

  (
    g1434_n,
    g1433_p,
    g1432_p
  );


  and

  (
    g1435_p,
    n7675_o2_p_spl_1,
    n2809_lo_p_spl_000
  );


  or

  (
    g1435_n,
    n7675_o2_n_spl_1,
    n2809_lo_n_spl_000
  );


  and

  (
    g1436_p,
    g1435_n_spl_,
    g1434_n_spl_
  );


  or

  (
    g1436_n,
    g1435_p_spl_,
    g1434_p_spl_
  );


  and

  (
    g1437_p,
    g1436_n_spl_0,
    g1434_n_spl_
  );


  or

  (
    g1437_n,
    g1436_p_spl_0,
    g1434_p_spl_
  );


  and

  (
    g1438_p,
    g1436_n_spl_0,
    g1435_n_spl_
  );


  or

  (
    g1438_n,
    g1436_p_spl_0,
    g1435_p_spl_
  );


  and

  (
    g1439_p,
    g1438_n,
    g1437_n
  );


  or

  (
    g1439_n,
    g1438_p,
    g1437_p
  );


  and

  (
    g1440_p,
    g1429_n_spl_0,
    g1427_n_spl_
  );


  or

  (
    g1440_n,
    g1429_p_spl_0,
    g1427_p_spl_
  );


  and

  (
    g1441_p,
    g1429_n_spl_,
    g1428_n_spl_
  );


  or

  (
    g1441_n,
    g1429_p_spl_,
    g1428_p_spl_
  );


  and

  (
    g1442_p,
    g1441_n,
    g1440_n
  );


  or

  (
    g1442_n,
    g1441_p,
    g1440_p
  );


  and

  (
    g1443_p,
    g1422_n_spl_0,
    g1420_n_spl_
  );


  or

  (
    g1443_n,
    g1422_p_spl_0,
    g1420_p_spl_
  );


  and

  (
    g1444_p,
    g1422_n_spl_,
    g1421_n_spl_
  );


  or

  (
    g1444_n,
    g1422_p_spl_,
    g1421_p_spl_
  );


  and

  (
    g1445_p,
    g1444_n,
    g1443_n
  );


  or

  (
    g1445_n,
    g1444_p,
    g1443_p
  );


  and

  (
    g1446_p,
    g1415_n_spl_0,
    g1413_n_spl_
  );


  or

  (
    g1446_n,
    g1415_p_spl_0,
    g1413_p_spl_
  );


  and

  (
    g1447_p,
    g1415_n_spl_,
    g1414_n_spl_
  );


  or

  (
    g1447_n,
    g1415_p_spl_,
    g1414_p_spl_
  );


  and

  (
    g1448_p,
    g1447_n,
    g1446_n
  );


  or

  (
    g1448_n,
    g1447_p,
    g1446_p
  );


  and

  (
    g1449_p,
    G3557_o2_n_spl_,
    G3494_o2_n_spl_
  );


  or

  (
    g1449_n,
    G3557_o2_p_spl_,
    G3494_o2_p_spl_
  );


  and

  (
    g1450_p,
    g1449_n_spl_0,
    G3557_o2_n_spl_
  );


  or

  (
    g1450_n,
    g1449_p_spl_0,
    G3557_o2_p_spl_
  );


  and

  (
    g1451_p,
    g1449_n_spl_0,
    G3494_o2_n_spl_
  );


  or

  (
    g1451_n,
    g1449_p_spl_0,
    G3494_o2_p_spl_
  );


  and

  (
    g1452_p,
    g1451_n,
    g1450_n
  );


  or

  (
    g1452_n,
    g1451_p,
    g1450_p
  );


  and

  (
    g1453_p,
    n2776_lo_buf_o2_p_spl_101,
    n7722_o2_p_spl_00
  );


  or

  (
    g1453_n,
    n2776_lo_buf_o2_n_spl_101,
    n7722_o2_n_spl_00
  );


  and

  (
    g1454_p,
    g1453_n_spl_,
    g1452_n_spl_
  );


  or

  (
    g1454_n,
    g1453_p_spl_,
    g1452_p_spl_
  );


  and

  (
    g1455_p,
    g1454_n_spl_0,
    g1449_n_spl_
  );


  or

  (
    g1455_n,
    g1454_p_spl_0,
    g1449_p_spl_
  );


  and

  (
    g1456_p,
    g1455_n_spl_,
    g1448_n_spl_
  );


  or

  (
    g1456_n,
    g1455_p_spl_,
    g1448_p_spl_
  );


  and

  (
    g1457_p,
    g1456_n_spl_0,
    g1448_n_spl_
  );


  or

  (
    g1457_n,
    g1456_p_spl_0,
    g1448_p_spl_
  );


  and

  (
    g1458_p,
    g1456_n_spl_0,
    g1455_n_spl_
  );


  or

  (
    g1458_n,
    g1456_p_spl_0,
    g1455_p_spl_
  );


  and

  (
    g1459_p,
    g1458_n,
    g1457_n
  );


  or

  (
    g1459_n,
    g1458_p,
    g1457_p
  );


  and

  (
    g1460_p,
    n7722_o2_p_spl_00,
    n2785_lo_p_spl_101
  );


  or

  (
    g1460_n,
    n7722_o2_n_spl_00,
    n2785_lo_n_spl_101
  );


  and

  (
    g1461_p,
    g1460_n_spl_,
    g1459_n_spl_
  );


  or

  (
    g1461_n,
    g1460_p_spl_,
    g1459_p_spl_
  );


  and

  (
    g1462_p,
    g1461_n_spl_0,
    g1456_n_spl_
  );


  or

  (
    g1462_n,
    g1461_p_spl_0,
    g1456_p_spl_
  );


  and

  (
    g1463_p,
    g1462_n_spl_,
    g1445_n_spl_
  );


  or

  (
    g1463_n,
    g1462_p_spl_,
    g1445_p_spl_
  );


  and

  (
    g1464_p,
    g1463_n_spl_0,
    g1445_n_spl_
  );


  or

  (
    g1464_n,
    g1463_p_spl_0,
    g1445_p_spl_
  );


  and

  (
    g1465_p,
    g1463_n_spl_0,
    g1462_n_spl_
  );


  or

  (
    g1465_n,
    g1463_p_spl_0,
    g1462_p_spl_
  );


  and

  (
    g1466_p,
    g1465_n,
    g1464_n
  );


  or

  (
    g1466_n,
    g1465_p,
    g1464_p
  );


  and

  (
    g1467_p,
    n7722_o2_p_spl_01,
    n2797_lo_p_spl_010
  );


  or

  (
    g1467_n,
    n7722_o2_n_spl_0,
    n2797_lo_n_spl_010
  );


  and

  (
    g1468_p,
    g1467_n_spl_,
    g1466_n_spl_
  );


  or

  (
    g1468_n,
    g1467_p_spl_,
    g1466_p_spl_
  );


  and

  (
    g1469_p,
    g1468_n_spl_0,
    g1463_n_spl_
  );


  or

  (
    g1469_n,
    g1468_p_spl_0,
    g1463_p_spl_
  );


  and

  (
    g1470_p,
    g1469_n_spl_,
    g1442_n_spl_
  );


  or

  (
    g1470_n,
    g1469_p_spl_,
    g1442_p_spl_
  );


  and

  (
    g1471_p,
    g1470_n_spl_0,
    g1442_n_spl_
  );


  or

  (
    g1471_n,
    g1470_p_spl_0,
    g1442_p_spl_
  );


  and

  (
    g1472_p,
    g1470_n_spl_0,
    g1469_n_spl_
  );


  or

  (
    g1472_n,
    g1470_p_spl_0,
    g1469_p_spl_
  );


  and

  (
    g1473_p,
    g1472_n,
    g1471_n
  );


  or

  (
    g1473_n,
    g1472_p,
    g1471_p
  );


  and

  (
    g1474_p,
    n7722_o2_p_spl_01,
    n2809_lo_p_spl_000
  );


  or

  (
    g1474_n,
    n7722_o2_n_spl_1,
    n2809_lo_n_spl_000
  );


  and

  (
    g1475_p,
    g1474_n_spl_,
    g1473_n_spl_
  );


  or

  (
    g1475_n,
    g1474_p_spl_,
    g1473_p_spl_
  );


  and

  (
    g1476_p,
    g1475_n_spl_0,
    g1470_n_spl_
  );


  or

  (
    g1476_n,
    g1475_p_spl_0,
    g1470_p_spl_
  );


  and

  (
    g1477_p,
    g1476_n_spl_,
    g1439_n_spl_
  );


  or

  (
    g1477_n,
    g1476_p_spl_,
    g1439_p_spl_
  );


  and

  (
    g1478_p,
    G1724_o2_p_spl_,
    G692_o2_n_spl_
  );


  or

  (
    g1478_n,
    G1724_o2_n_spl_,
    G692_o2_p_spl_
  );


  and

  (
    g1479_p,
    g1478_n_spl_0,
    G1724_o2_p_spl_
  );


  or

  (
    g1479_n,
    g1478_p_spl_0,
    G1724_o2_n_spl_
  );


  and

  (
    g1480_p,
    g1478_n_spl_0,
    G692_o2_n_spl_
  );


  or

  (
    g1480_n,
    g1478_p_spl_0,
    G692_o2_p_spl_
  );


  and

  (
    g1481_p,
    g1480_n,
    g1479_n
  );


  or

  (
    g1481_n,
    g1480_p,
    g1479_p
  );


  and

  (
    g1482_p,
    g1078_n_spl_,
    G1634_o2_p
  );


  or

  (
    g1482_n,
    g1078_p_spl_,
    G1634_o2_n
  );


  and

  (
    g1483_p,
    g1482_n_spl_,
    g1481_n_spl_
  );


  or

  (
    g1483_n,
    g1482_p_spl_,
    g1481_p_spl_
  );


  and

  (
    g1484_p,
    g1483_n_spl_0,
    g1481_n_spl_
  );


  or

  (
    g1484_n,
    g1483_p_spl_0,
    g1481_p_spl_
  );


  and

  (
    g1485_p,
    g1483_n_spl_0,
    g1482_n_spl_
  );


  or

  (
    g1485_n,
    g1483_p_spl_0,
    g1482_p_spl_
  );


  and

  (
    g1486_p,
    g1485_n,
    g1484_n
  );


  or

  (
    g1486_n,
    g1485_p,
    g1484_p
  );


  and

  (
    g1487_p,
    n2716_lo_buf_o2_p_spl_00,
    n2512_lo_buf_o2_p_spl_00
  );


  or

  (
    g1487_n,
    n2716_lo_buf_o2_n_spl_00,
    n2512_lo_buf_o2_n_spl_00
  );


  and

  (
    g1488_p,
    g1487_n_spl_,
    g1486_n_spl_
  );


  or

  (
    g1488_n,
    g1487_p_spl_,
    g1486_p_spl_
  );


  and

  (
    g1489_p,
    g1488_n_spl_0,
    g1486_n_spl_
  );


  or

  (
    g1489_n,
    g1488_p_spl_0,
    g1486_p_spl_
  );


  and

  (
    g1490_p,
    g1488_n_spl_0,
    g1487_n_spl_
  );


  or

  (
    g1490_n,
    g1488_p_spl_0,
    g1487_p_spl_
  );


  and

  (
    g1491_p,
    g1490_n,
    g1489_n
  );


  or

  (
    g1491_n,
    g1490_p,
    g1489_p
  );


  and

  (
    g1492_p,
    g1088_n_spl_,
    g1083_n_spl_
  );


  or

  (
    g1492_n,
    g1088_p_spl_,
    g1083_p_spl_
  );


  and

  (
    g1493_p,
    g1492_n_spl_,
    g1491_n_spl_
  );


  or

  (
    g1493_n,
    g1492_p_spl_,
    g1491_p_spl_
  );


  and

  (
    g1494_p,
    g1493_n_spl_0,
    g1491_n_spl_
  );


  or

  (
    g1494_n,
    g1493_p_spl_0,
    g1491_p_spl_
  );


  and

  (
    g1495_p,
    g1493_n_spl_0,
    g1492_n_spl_
  );


  or

  (
    g1495_n,
    g1493_p_spl_0,
    g1492_p_spl_
  );


  and

  (
    g1496_p,
    g1495_n,
    g1494_n
  );


  or

  (
    g1496_n,
    g1495_p,
    g1494_p
  );


  and

  (
    g1497_p,
    n2728_lo_buf_o2_p_spl_000,
    n2500_lo_buf_o2_p_spl_01
  );


  or

  (
    g1497_n,
    n2728_lo_buf_o2_n_spl_000,
    n2500_lo_buf_o2_n_spl_0
  );


  and

  (
    g1498_p,
    g1497_n_spl_,
    g1496_n_spl_
  );


  or

  (
    g1498_n,
    g1497_p_spl_,
    g1496_p_spl_
  );


  and

  (
    g1499_p,
    g1498_n_spl_0,
    g1496_n_spl_
  );


  or

  (
    g1499_n,
    g1498_p_spl_0,
    g1496_p_spl_
  );


  and

  (
    g1500_p,
    g1498_n_spl_0,
    g1497_n_spl_
  );


  or

  (
    g1500_n,
    g1498_p_spl_0,
    g1497_p_spl_
  );


  and

  (
    g1501_p,
    g1500_n,
    g1499_n
  );


  or

  (
    g1501_n,
    g1500_p,
    g1499_p
  );


  and

  (
    g1502_p,
    g1097_n,
    g1093_n_spl_
  );


  or

  (
    g1502_n,
    g1097_p_spl_,
    g1093_p_spl_
  );


  and

  (
    g1503_p,
    g1502_n_spl_,
    g1501_n_spl_
  );


  or

  (
    g1503_n,
    g1502_p_spl_,
    g1501_p_spl_
  );


  and

  (
    g1504_p,
    g1503_n_spl_0,
    g1501_n_spl_
  );


  or

  (
    g1504_n,
    g1503_p_spl_0,
    g1501_p_spl_
  );


  and

  (
    g1505_p,
    g1503_n_spl_0,
    g1502_n_spl_
  );


  or

  (
    g1505_n,
    g1503_p_spl_0,
    g1502_p_spl_
  );


  and

  (
    g1506_p,
    g1505_n,
    g1504_n
  );


  or

  (
    g1506_n,
    g1505_p,
    g1504_p
  );


  and

  (
    g1507_p,
    n8086_o2_p_spl_1,
    n2809_lo_p_spl_001
  );


  or

  (
    g1507_n,
    n8086_o2_n_spl_1,
    n2809_lo_n_spl_001
  );


  and

  (
    g1508_p,
    g1506_n_spl_,
    g1215_n
  );


  or

  (
    g1508_n,
    g1506_p,
    g1215_p_spl_
  );


  and

  (
    g1509_p,
    G3492_o2_n,
    G3493_o2_p
  );


  or

  (
    g1509_n,
    G3492_o2_p,
    G3493_o2_n
  );


  and

  (
    g1510_p,
    G3422_o2_n_spl_,
    G3269_o2_p
  );


  or

  (
    g1510_n,
    G3422_o2_p_spl_,
    G3269_o2_n
  );


  and

  (
    g1511_p,
    g1510_n_spl_,
    g1509_n_spl_
  );


  or

  (
    g1511_n,
    g1510_p_spl_,
    g1509_p_spl_
  );


  and

  (
    g1512_p,
    g1511_n_spl_0,
    g1509_n_spl_
  );


  or

  (
    g1512_n,
    g1511_p_spl_0,
    g1509_p_spl_
  );


  and

  (
    g1513_p,
    g1511_n_spl_0,
    g1510_n_spl_
  );


  or

  (
    g1513_n,
    g1511_p_spl_0,
    g1510_p_spl_
  );


  and

  (
    g1514_p,
    g1513_n,
    g1512_n
  );


  or

  (
    g1514_n,
    g1513_p,
    g1512_p
  );


  and

  (
    g1515_p,
    n2776_lo_buf_o2_p_spl_11,
    n7747_o2_p_spl_00
  );


  or

  (
    g1515_n,
    n2776_lo_buf_o2_n_spl_11,
    n7747_o2_n_spl_00
  );


  and

  (
    g1516_p,
    g1515_n_spl_,
    g1514_n_spl_
  );


  or

  (
    g1516_n,
    g1515_p_spl_,
    g1514_p_spl_
  );


  and

  (
    g1517_p,
    g1516_n_spl_0,
    g1514_n_spl_
  );


  or

  (
    g1517_n,
    g1516_p_spl_0,
    g1514_p_spl_
  );


  and

  (
    g1518_p,
    g1516_n_spl_0,
    g1515_n_spl_
  );


  or

  (
    g1518_n,
    g1516_p_spl_0,
    g1515_p_spl_
  );


  and

  (
    g1519_p,
    g1518_n,
    g1517_n
  );


  or

  (
    g1519_n,
    g1518_p,
    g1517_p
  );


  and

  (
    g1520_p,
    g1055_n_spl_,
    g1050_n_spl_
  );


  or

  (
    g1520_n,
    g1055_p_spl_,
    g1050_p_spl_
  );


  and

  (
    g1521_p,
    g1520_n_spl_,
    g1519_n_spl_
  );


  or

  (
    g1521_n,
    g1520_p_spl_,
    g1519_p_spl_
  );


  and

  (
    g1522_p,
    g1521_n_spl_0,
    g1519_n_spl_
  );


  or

  (
    g1522_n,
    g1521_p_spl_0,
    g1519_p_spl_
  );


  and

  (
    g1523_p,
    g1521_n_spl_0,
    g1520_n_spl_
  );


  or

  (
    g1523_n,
    g1521_p_spl_0,
    g1520_p_spl_
  );


  and

  (
    g1524_p,
    g1523_n,
    g1522_n
  );


  or

  (
    g1524_n,
    g1523_p,
    g1522_p
  );


  and

  (
    g1525_p,
    n7835_o2_p_spl_00,
    n2785_lo_p_spl_101
  );


  or

  (
    g1525_n,
    n7835_o2_n_spl_00,
    n2785_lo_n_spl_101
  );


  and

  (
    g1526_p,
    g1525_n_spl_,
    g1524_n_spl_
  );


  or

  (
    g1526_n,
    g1525_p_spl_,
    g1524_p_spl_
  );


  and

  (
    g1527_p,
    g1526_n_spl_0,
    g1524_n_spl_
  );


  or

  (
    g1527_n,
    g1526_p_spl_0,
    g1524_p_spl_
  );


  and

  (
    g1528_p,
    g1526_n_spl_0,
    g1525_n_spl_
  );


  or

  (
    g1528_n,
    g1526_p_spl_0,
    g1525_p_spl_
  );


  and

  (
    g1529_p,
    g1528_n,
    g1527_n
  );


  or

  (
    g1529_n,
    g1528_p,
    g1527_p
  );


  and

  (
    g1530_p,
    g1065_n_spl_,
    g1060_n_spl_
  );


  or

  (
    g1530_n,
    g1065_p_spl_,
    g1060_p_spl_
  );


  and

  (
    g1531_p,
    g1530_n_spl_,
    g1529_n_spl_
  );


  or

  (
    g1531_n,
    g1530_p_spl_,
    g1529_p_spl_
  );


  and

  (
    g1532_p,
    g1531_n_spl_0,
    g1529_n_spl_
  );


  or

  (
    g1532_n,
    g1531_p_spl_0,
    g1529_p_spl_
  );


  and

  (
    g1533_p,
    g1531_n_spl_0,
    g1530_n_spl_
  );


  or

  (
    g1533_n,
    g1531_p_spl_0,
    g1530_p_spl_
  );


  and

  (
    g1534_p,
    g1533_n,
    g1532_n
  );


  or

  (
    g1534_n,
    g1533_p,
    g1532_p
  );


  and

  (
    g1535_p,
    n7909_o2_p_spl_01,
    n2797_lo_p_spl_011
  );


  or

  (
    g1535_n,
    n7909_o2_n_spl_1,
    n2797_lo_n_spl_011
  );


  and

  (
    g1536_p,
    g1535_n_spl_,
    g1534_n_spl_
  );


  or

  (
    g1536_n,
    g1535_p_spl_,
    g1534_p_spl_
  );


  and

  (
    g1537_p,
    g1536_n_spl_0,
    g1534_n_spl_
  );


  or

  (
    g1537_n,
    g1536_p_spl_0,
    g1534_p_spl_
  );


  and

  (
    g1538_p,
    g1536_n_spl_0,
    g1535_n_spl_
  );


  or

  (
    g1538_n,
    g1536_p_spl_0,
    g1535_p_spl_
  );


  and

  (
    g1539_p,
    g1538_n,
    g1537_n
  );


  or

  (
    g1539_n,
    g1538_p,
    g1537_p
  );


  and

  (
    g1540_p,
    g1075_n,
    g1070_n_spl_
  );


  or

  (
    g1540_n,
    g1075_p_spl_,
    g1070_p_spl_
  );


  and

  (
    g1541_p,
    g1540_n_spl_,
    g1539_n_spl_
  );


  or

  (
    g1541_n,
    g1540_p_spl_,
    g1539_p_spl_
  );


  and

  (
    g1542_p,
    g1541_n_spl_0,
    g1539_n_spl_
  );


  or

  (
    g1542_n,
    g1541_p_spl_0,
    g1539_p_spl_
  );


  and

  (
    g1543_p,
    g1541_n_spl_0,
    g1540_n_spl_
  );


  or

  (
    g1543_n,
    g1541_p_spl_0,
    g1540_p_spl_
  );


  and

  (
    g1544_p,
    g1543_n,
    g1542_n
  );


  or

  (
    g1544_n,
    g1543_p,
    g1542_p
  );


  or

  (
    g1545_n,
    n6075_o2_n_spl_1,
    n2860_lo_n_spl_10
  );


  or

  (
    g1546_n,
    n5930_o2_n_spl_1,
    n2848_lo_n_spl_11
  );


  or

  (
    g1547_n,
    n5792_o2_n_spl_1,
    n2836_lo_n_spl_110
  );


  or

  (
    g1548_n,
    g1231_p_spl_,
    g1211_p
  );


  and

  (
    g1549_p,
    g859_n_spl_0,
    g857_n_spl_
  );


  or

  (
    g1549_n,
    g859_p_spl_0,
    g857_p_spl_
  );


  and

  (
    g1550_p,
    g859_n_spl_,
    g858_n_spl_
  );


  or

  (
    g1550_n,
    g859_p_spl_,
    g858_p_spl_
  );


  and

  (
    g1551_p,
    g1550_n,
    g1549_n
  );


  or

  (
    g1551_n,
    g1550_p,
    g1549_p
  );


  and

  (
    g1552_p,
    g1111_n_spl_,
    g1106_n_spl_
  );


  or

  (
    g1552_n,
    g1111_p_spl_,
    g1106_p_spl_
  );


  and

  (
    g1553_p,
    g1552_n_spl_,
    g1551_n_spl_
  );


  or

  (
    g1553_n,
    g1552_p_spl_,
    g1551_p_spl_
  );


  and

  (
    g1554_p,
    g1553_n_spl_0,
    g1551_n_spl_
  );


  or

  (
    g1554_n,
    g1553_p_spl_,
    g1551_p_spl_
  );


  and

  (
    g1555_p,
    g1553_n_spl_0,
    g1552_n_spl_
  );


  or

  (
    g1555_n,
    g1553_p_spl_,
    g1552_p_spl_
  );


  and

  (
    g1556_p,
    g1555_n,
    g1554_n
  );


  or

  (
    g1556_n,
    g1555_p,
    g1554_p
  );


  and

  (
    g1557_p,
    n5863_o2_p_spl_1,
    n2836_lo_p_spl_110
  );


  or

  (
    g1557_n,
    n5863_o2_n_spl_,
    n2836_lo_n_spl_11
  );


  and

  (
    g1558_p,
    g1557_n_spl_,
    g1556_n_spl_
  );


  or

  (
    g1558_n,
    g1557_p_spl_,
    g1556_p_spl_
  );


  and

  (
    g1559_p,
    g1558_n_spl_0,
    g1556_n_spl_
  );


  or

  (
    g1559_n,
    g1558_p_spl_,
    g1556_p_spl_
  );


  and

  (
    g1560_p,
    g1558_n_spl_0,
    g1557_n_spl_
  );


  or

  (
    g1560_n,
    g1558_p_spl_,
    g1557_p_spl_
  );


  and

  (
    g1561_p,
    g1560_n,
    g1559_n
  );


  or

  (
    g1561_n,
    g1560_p,
    g1559_p
  );


  and

  (
    g1562_p,
    g1121_n_spl_,
    g1116_n_spl_
  );


  or

  (
    g1562_n,
    g1121_p_spl_,
    g1116_p_spl_
  );


  or

  (
    g1563_n,
    g1562_p,
    g1561_p
  );


  and

  (
    g1564_p,
    g933_n_spl_0,
    g931_n_spl_
  );


  or

  (
    g1564_n,
    g933_p_spl_0,
    g931_p_spl_
  );


  and

  (
    g1565_p,
    g933_n_spl_,
    g932_n_spl_
  );


  or

  (
    g1565_n,
    g933_p_spl_,
    g932_p_spl_
  );


  and

  (
    g1566_p,
    g1565_n,
    g1564_n
  );


  or

  (
    g1566_n,
    g1565_p,
    g1564_p
  );


  and

  (
    g1567_p,
    g1136_n_spl_,
    g1131_n_spl_
  );


  or

  (
    g1567_n,
    g1136_p_spl_,
    g1131_p_spl_
  );


  and

  (
    g1568_p,
    g1567_n_spl_,
    g1566_n_spl_
  );


  or

  (
    g1568_n,
    g1567_p_spl_,
    g1566_p_spl_
  );


  and

  (
    g1569_p,
    g1568_n_spl_0,
    g1566_n_spl_
  );


  or

  (
    g1569_n,
    g1568_p_spl_,
    g1566_p_spl_
  );


  and

  (
    g1570_p,
    g1568_n_spl_0,
    g1567_n_spl_
  );


  or

  (
    g1570_n,
    g1568_p_spl_,
    g1567_p_spl_
  );


  and

  (
    g1571_p,
    g1570_n,
    g1569_n
  );


  or

  (
    g1571_n,
    g1570_p,
    g1569_p
  );


  and

  (
    g1572_p,
    n5981_o2_p_spl_1,
    n2848_lo_p_spl_11
  );


  or

  (
    g1572_n,
    n5981_o2_n_spl_,
    n2848_lo_n_spl_11
  );


  and

  (
    g1573_p,
    g1572_n_spl_,
    g1571_n_spl_
  );


  or

  (
    g1573_n,
    g1572_p_spl_,
    g1571_p_spl_
  );


  and

  (
    g1574_p,
    g1573_n_spl_0,
    g1571_n_spl_
  );


  or

  (
    g1574_n,
    g1573_p_spl_,
    g1571_p_spl_
  );


  and

  (
    g1575_p,
    g1573_n_spl_0,
    g1572_n_spl_
  );


  or

  (
    g1575_n,
    g1573_p_spl_,
    g1572_p_spl_
  );


  and

  (
    g1576_p,
    g1575_n,
    g1574_n
  );


  or

  (
    g1576_n,
    g1575_p,
    g1574_p
  );


  and

  (
    g1577_p,
    g1146_n_spl_,
    g1141_n_spl_
  );


  or

  (
    g1577_n,
    g1146_p_spl_,
    g1141_p_spl_
  );


  or

  (
    g1578_n,
    g1577_p,
    g1576_p
  );


  and

  (
    g1579_p,
    g1007_n_spl_0,
    g1005_n_spl_
  );


  or

  (
    g1579_n,
    g1007_p_spl_0,
    g1005_p_spl_
  );


  and

  (
    g1580_p,
    g1007_n_spl_,
    g1006_n_spl_
  );


  or

  (
    g1580_n,
    g1007_p_spl_,
    g1006_p_spl_
  );


  and

  (
    g1581_p,
    g1580_n,
    g1579_n
  );


  or

  (
    g1581_n,
    g1580_p,
    g1579_p
  );


  and

  (
    g1582_p,
    g1171_n_spl_,
    g1166_n_spl_
  );


  or

  (
    g1582_n,
    g1171_p_spl_,
    g1166_p_spl_
  );


  and

  (
    g1583_p,
    g1582_n_spl_,
    g1581_n_spl_
  );


  or

  (
    g1583_n,
    g1582_p_spl_,
    g1581_p_spl_
  );


  and

  (
    g1584_p,
    g1583_n_spl_0,
    g1581_n_spl_
  );


  or

  (
    g1584_n,
    g1583_p_spl_,
    g1581_p_spl_
  );


  and

  (
    g1585_p,
    g1583_n_spl_0,
    g1582_n_spl_
  );


  or

  (
    g1585_n,
    g1583_p_spl_,
    g1582_p_spl_
  );


  and

  (
    g1586_p,
    g1585_n,
    g1584_n
  );


  or

  (
    g1586_n,
    g1585_p,
    g1584_p
  );


  and

  (
    g1587_p,
    n6169_o2_p_spl_,
    n2860_lo_p_spl_10
  );


  or

  (
    g1587_n,
    n6169_o2_n_spl_,
    n2860_lo_n_spl_1
  );


  and

  (
    g1588_p,
    g1587_n_spl_,
    g1586_n_spl_
  );


  or

  (
    g1588_n,
    g1587_p_spl_,
    g1586_p_spl_
  );


  and

  (
    g1589_p,
    g1588_n_spl_0,
    g1586_n_spl_
  );


  or

  (
    g1589_n,
    g1588_p_spl_,
    g1586_p_spl_
  );


  and

  (
    g1590_p,
    g1588_n_spl_0,
    g1587_n_spl_
  );


  or

  (
    g1590_n,
    g1588_p_spl_,
    g1587_p_spl_
  );


  and

  (
    g1591_p,
    g1590_n,
    g1589_n
  );


  or

  (
    g1591_n,
    g1590_p,
    g1589_p
  );


  and

  (
    g1592_p,
    g1191_n_spl_,
    g1186_n_spl_
  );


  or

  (
    g1592_n,
    g1191_p_spl_,
    g1186_p_spl_
  );


  or

  (
    g1593_n,
    g1592_p,
    g1591_p
  );


  and

  (
    g1594_p,
    g1101_n_spl_0,
    g1099_n
  );


  and

  (
    g1595_p,
    g1101_n_spl_0,
    g1100_n
  );


  or

  (
    g1596_n,
    g1595_p,
    g1594_p
  );


  and

  (
    g1597_p,
    g1126_n_spl_0,
    g1124_n
  );


  and

  (
    g1598_p,
    g1126_n_spl_0,
    g1125_n
  );


  or

  (
    g1599_n,
    g1598_p,
    g1597_p
  );


  and

  (
    g1600_p,
    g1151_n_spl_0,
    g1149_n
  );


  and

  (
    g1601_p,
    g1151_n_spl_0,
    g1150_n
  );


  or

  (
    g1602_n,
    g1601_p,
    g1600_p
  );


  and

  (
    g1603_p,
    g1206_n_spl_0,
    g1194_n
  );


  and

  (
    g1604_p,
    g1206_n_spl_0,
    g1205_n
  );


  or

  (
    g1605_n,
    g1604_p,
    g1603_p
  );


  and

  (
    g1606_p,
    g1544_n_spl_,
    g1507_n
  );


  or

  (
    g1606_n,
    g1544_p,
    g1507_p_spl_
  );


  and

  (
    g1607_p,
    n2776_lo_buf_o2_p_spl_11,
    n7148_o2_p_spl_0
  );


  or

  (
    g1607_n,
    n2776_lo_buf_o2_n_spl_11,
    n7148_o2_n_spl_0
  );


  and

  (
    g1608_p,
    g1245_n_spl_,
    g1240_n_spl_
  );


  or

  (
    g1608_n,
    g1245_p_spl_,
    g1240_p_spl_
  );


  and

  (
    g1609_p,
    g1608_n_spl_,
    g1607_n_spl_
  );


  or

  (
    g1609_n,
    g1608_p_spl_,
    g1607_p_spl_
  );


  and

  (
    g1610_p,
    g1609_n_spl_0,
    g1607_n_spl_
  );


  or

  (
    g1610_n,
    g1609_p_spl_0,
    g1607_p_spl_
  );


  and

  (
    g1611_p,
    g1609_n_spl_0,
    g1608_n_spl_
  );


  or

  (
    g1611_n,
    g1609_p_spl_0,
    g1608_p_spl_
  );


  and

  (
    g1612_p,
    g1611_n,
    g1610_n
  );


  or

  (
    g1612_n,
    g1611_p,
    g1610_p
  );


  and

  (
    g1613_p,
    n7224_o2_p_spl_1,
    n2785_lo_p_spl_110
  );


  or

  (
    g1613_n,
    n7224_o2_n_spl_,
    n2785_lo_n_spl_110
  );


  and

  (
    g1614_p,
    g1613_n_spl_,
    g1612_n_spl_
  );


  or

  (
    g1614_n,
    g1613_p_spl_,
    g1612_p_spl_
  );


  and

  (
    g1615_p,
    g1614_n_spl_0,
    g1612_n_spl_
  );


  or

  (
    g1615_n,
    g1614_p_spl_0,
    g1612_p_spl_
  );


  and

  (
    g1616_p,
    g1614_n_spl_0,
    g1613_n_spl_
  );


  or

  (
    g1616_n,
    g1614_p_spl_0,
    g1613_p_spl_
  );


  and

  (
    g1617_p,
    g1616_n,
    g1615_n
  );


  or

  (
    g1617_n,
    g1616_p,
    g1615_p
  );


  and

  (
    g1618_p,
    g1268_n_spl_,
    g1263_n_spl_
  );


  or

  (
    g1618_n,
    g1268_p_spl_,
    g1263_p_spl_
  );


  or

  (
    g1619_n,
    g1618_p,
    g1617_p
  );


  and

  (
    g1620_p,
    g1284_n_spl_0,
    g1282_n_spl_
  );


  or

  (
    g1620_n,
    g1284_p_spl_0,
    g1282_p_spl_
  );


  and

  (
    g1621_p,
    g1284_n_spl_,
    g1283_n_spl_
  );


  or

  (
    g1621_n,
    g1284_p_spl_,
    g1283_p_spl_
  );


  and

  (
    g1622_p,
    g1621_n,
    g1620_n
  );


  or

  (
    g1622_n,
    g1621_p,
    g1620_p
  );


  and

  (
    g1623_p,
    g1303_n_spl_,
    g1298_n_spl_
  );


  or

  (
    g1623_n,
    g1303_p_spl_,
    g1298_p_spl_
  );


  and

  (
    g1624_p,
    g1623_n_spl_,
    g1622_n_spl_
  );


  or

  (
    g1624_n,
    g1623_p_spl_,
    g1622_p_spl_
  );


  and

  (
    g1625_p,
    g1624_n_spl_0,
    g1622_n_spl_
  );


  or

  (
    g1625_n,
    g1624_p_spl_0,
    g1622_p_spl_
  );


  and

  (
    g1626_p,
    g1624_n_spl_0,
    g1623_n_spl_
  );


  or

  (
    g1626_n,
    g1624_p_spl_0,
    g1623_p_spl_
  );


  and

  (
    g1627_p,
    g1626_n,
    g1625_n
  );


  or

  (
    g1627_n,
    g1626_p,
    g1625_p
  );


  and

  (
    g1628_p,
    n7323_o2_p_spl_0,
    n2785_lo_p_spl_110
  );


  or

  (
    g1628_n,
    n7323_o2_n_spl_0,
    n2785_lo_n_spl_110
  );


  and

  (
    g1629_p,
    g1628_n_spl_,
    g1627_n_spl_
  );


  or

  (
    g1629_n,
    g1628_p_spl_,
    g1627_p_spl_
  );


  and

  (
    g1630_p,
    g1629_n_spl_0,
    g1627_n_spl_
  );


  or

  (
    g1630_n,
    g1629_p_spl_0,
    g1627_p_spl_
  );


  and

  (
    g1631_p,
    g1629_n_spl_0,
    g1628_n_spl_
  );


  or

  (
    g1631_n,
    g1629_p_spl_0,
    g1628_p_spl_
  );


  and

  (
    g1632_p,
    g1631_n,
    g1630_n
  );


  or

  (
    g1632_n,
    g1631_p,
    g1630_p
  );


  and

  (
    g1633_p,
    g1319_n_spl_,
    g1314_n_spl_
  );


  or

  (
    g1633_n,
    g1319_p_spl_,
    g1314_p_spl_
  );


  and

  (
    g1634_p,
    g1633_n_spl_,
    g1632_n_spl_
  );


  or

  (
    g1634_n,
    g1633_p_spl_,
    g1632_p_spl_
  );


  and

  (
    g1635_p,
    g1634_n_spl_0,
    g1632_n_spl_
  );


  or

  (
    g1635_n,
    g1634_p_spl_0,
    g1632_p_spl_
  );


  and

  (
    g1636_p,
    g1634_n_spl_0,
    g1633_n_spl_
  );


  or

  (
    g1636_n,
    g1634_p_spl_0,
    g1633_p_spl_
  );


  and

  (
    g1637_p,
    g1636_n,
    g1635_n
  );


  or

  (
    g1637_n,
    g1636_p,
    g1635_p
  );


  and

  (
    g1638_p,
    n7398_o2_p_spl_1,
    n2797_lo_p_spl_011
  );


  or

  (
    g1638_n,
    n7398_o2_n_spl_,
    n2797_lo_n_spl_011
  );


  and

  (
    g1639_p,
    g1638_n_spl_,
    g1637_n_spl_
  );


  or

  (
    g1639_n,
    g1638_p_spl_,
    g1637_p_spl_
  );


  and

  (
    g1640_p,
    g1639_n_spl_0,
    g1637_n_spl_
  );


  or

  (
    g1640_n,
    g1639_p_spl_0,
    g1637_p_spl_
  );


  and

  (
    g1641_p,
    g1639_n_spl_0,
    g1638_n_spl_
  );


  or

  (
    g1641_n,
    g1639_p_spl_0,
    g1638_p_spl_
  );


  and

  (
    g1642_p,
    g1641_n,
    g1640_n
  );


  or

  (
    g1642_n,
    g1641_p,
    g1640_p
  );


  and

  (
    g1643_p,
    g1342_n_spl_,
    g1337_n_spl_
  );


  or

  (
    g1643_n,
    g1342_p_spl_,
    g1337_p_spl_
  );


  or

  (
    g1644_n,
    g1643_p,
    g1642_p
  );


  and

  (
    g1645_p,
    g1358_n_spl_0,
    g1356_n_spl_
  );


  or

  (
    g1645_n,
    g1358_p_spl_0,
    g1356_p_spl_
  );


  and

  (
    g1646_p,
    g1358_n_spl_,
    g1357_n_spl_
  );


  or

  (
    g1646_n,
    g1358_p_spl_,
    g1357_p_spl_
  );


  and

  (
    g1647_p,
    g1646_n,
    g1645_n
  );


  or

  (
    g1647_n,
    g1646_p,
    g1645_p
  );


  and

  (
    g1648_p,
    g1378_n_spl_,
    g1373_n_spl_
  );


  or

  (
    g1648_n,
    g1378_p_spl_,
    g1373_p_spl_
  );


  and

  (
    g1649_p,
    g1648_n_spl_,
    g1647_n_spl_
  );


  or

  (
    g1649_n,
    g1648_p_spl_,
    g1647_p_spl_
  );


  and

  (
    g1650_p,
    g1649_n_spl_0,
    g1647_n_spl_
  );


  or

  (
    g1650_n,
    g1649_p_spl_0,
    g1647_p_spl_
  );


  and

  (
    g1651_p,
    g1649_n_spl_0,
    g1648_n_spl_
  );


  or

  (
    g1651_n,
    g1649_p_spl_0,
    g1648_p_spl_
  );


  and

  (
    g1652_p,
    g1651_n,
    g1650_n
  );


  or

  (
    g1652_n,
    g1651_p,
    g1650_p
  );


  and

  (
    g1653_p,
    n7518_o2_p_spl_0,
    n2797_lo_p_spl_100
  );


  or

  (
    g1653_n,
    n7518_o2_n_spl_0,
    n2797_lo_n_spl_100
  );


  and

  (
    g1654_p,
    g1653_n_spl_,
    g1652_n_spl_
  );


  or

  (
    g1654_n,
    g1653_p_spl_,
    g1652_p_spl_
  );


  and

  (
    g1655_p,
    g1654_n_spl_0,
    g1652_n_spl_
  );


  or

  (
    g1655_n,
    g1654_p_spl_0,
    g1652_p_spl_
  );


  and

  (
    g1656_p,
    g1654_n_spl_0,
    g1653_n_spl_
  );


  or

  (
    g1656_n,
    g1654_p_spl_0,
    g1653_p_spl_
  );


  and

  (
    g1657_p,
    g1656_n,
    g1655_n
  );


  or

  (
    g1657_n,
    g1656_p,
    g1655_p
  );


  and

  (
    g1658_p,
    g1401_n_spl_,
    g1396_n_spl_
  );


  or

  (
    g1658_n,
    g1401_p_spl_,
    g1396_p_spl_
  );


  and

  (
    g1659_p,
    g1658_n_spl_,
    g1657_n_spl_
  );


  or

  (
    g1659_n,
    g1658_p_spl_,
    g1657_p_spl_
  );


  and

  (
    g1660_p,
    g1659_n_spl_0,
    g1657_n_spl_
  );


  or

  (
    g1660_n,
    g1659_p_spl_0,
    g1657_p_spl_
  );


  and

  (
    g1661_p,
    g1659_n_spl_0,
    g1658_n_spl_
  );


  or

  (
    g1661_n,
    g1659_p_spl_0,
    g1658_p_spl_
  );


  and

  (
    g1662_p,
    g1661_n,
    g1660_n
  );


  or

  (
    g1662_n,
    g1661_p,
    g1660_p
  );


  and

  (
    g1663_p,
    n7606_o2_p_spl_1,
    n2809_lo_p_spl_001
  );


  or

  (
    g1663_n,
    n7606_o2_n_spl_1,
    n2809_lo_n_spl_001
  );


  and

  (
    g1664_p,
    g1663_n_spl_,
    g1662_n_spl_
  );


  or

  (
    g1664_n,
    g1663_p_spl_,
    g1662_p_spl_
  );


  and

  (
    g1665_p,
    g1664_n_spl_0,
    g1662_n_spl_
  );


  or

  (
    g1665_n,
    g1664_p_spl_0,
    g1662_p_spl_
  );


  and

  (
    g1666_p,
    g1664_n_spl_0,
    g1663_n_spl_
  );


  or

  (
    g1666_n,
    g1664_p_spl_0,
    g1663_p_spl_
  );


  and

  (
    g1667_p,
    g1666_n,
    g1665_n
  );


  or

  (
    g1667_n,
    g1666_p,
    g1665_p
  );


  and

  (
    g1668_p,
    g1436_n_spl_,
    g1431_n_spl_
  );


  or

  (
    g1668_n,
    g1436_p_spl_,
    g1431_p_spl_
  );


  or

  (
    g1669_n,
    g1668_p,
    g1667_p
  );


  and

  (
    g1670_p,
    g1468_n_spl_0,
    g1466_n_spl_
  );


  or

  (
    g1670_n,
    g1468_p_spl_0,
    g1466_p_spl_
  );


  and

  (
    g1671_p,
    g1468_n_spl_,
    g1467_n_spl_
  );


  or

  (
    g1671_n,
    g1468_p_spl_,
    g1467_p_spl_
  );


  and

  (
    g1672_p,
    g1671_n,
    g1670_n
  );


  or

  (
    g1672_n,
    g1671_p,
    g1670_p
  );


  and

  (
    g1673_p,
    g1461_n_spl_0,
    g1459_n_spl_
  );


  or

  (
    g1673_n,
    g1461_p_spl_0,
    g1459_p_spl_
  );


  and

  (
    g1674_p,
    g1461_n_spl_,
    g1460_n_spl_
  );


  or

  (
    g1674_n,
    g1461_p_spl_,
    g1460_p_spl_
  );


  and

  (
    g1675_p,
    g1674_n,
    g1673_n
  );


  or

  (
    g1675_n,
    g1674_p,
    g1673_p
  );


  and

  (
    g1676_p,
    g1454_n_spl_0,
    g1452_n_spl_
  );


  or

  (
    g1676_n,
    g1454_p_spl_0,
    g1452_p_spl_
  );


  and

  (
    g1677_p,
    g1454_n_spl_,
    g1453_n_spl_
  );


  or

  (
    g1677_n,
    g1454_p_spl_,
    g1453_p_spl_
  );


  and

  (
    g1678_p,
    g1677_n,
    g1676_n
  );


  or

  (
    g1678_n,
    g1677_p,
    g1676_p
  );


  and

  (
    g1679_p,
    g1516_n_spl_,
    g1511_n_spl_
  );


  or

  (
    g1679_n,
    g1516_p_spl_,
    g1511_p_spl_
  );


  and

  (
    g1680_p,
    g1679_n_spl_,
    g1678_n_spl_
  );


  or

  (
    g1680_n,
    g1679_p_spl_,
    g1678_p_spl_
  );


  and

  (
    g1681_p,
    g1680_n_spl_0,
    g1678_n_spl_
  );


  or

  (
    g1681_n,
    g1680_p_spl_0,
    g1678_p_spl_
  );


  and

  (
    g1682_p,
    g1680_n_spl_0,
    g1679_n_spl_
  );


  or

  (
    g1682_n,
    g1680_p_spl_0,
    g1679_p_spl_
  );


  and

  (
    g1683_p,
    g1682_n,
    g1681_n
  );


  or

  (
    g1683_n,
    g1682_p,
    g1681_p
  );


  and

  (
    g1684_p,
    n7747_o2_p_spl_00,
    n2785_lo_p_spl_111
  );


  or

  (
    g1684_n,
    n7747_o2_n_spl_00,
    n2785_lo_n_spl_111
  );


  and

  (
    g1685_p,
    g1684_n_spl_,
    g1683_n_spl_
  );


  or

  (
    g1685_n,
    g1684_p_spl_,
    g1683_p_spl_
  );


  and

  (
    g1686_p,
    g1685_n_spl_0,
    g1680_n_spl_
  );


  or

  (
    g1686_n,
    g1685_p_spl_0,
    g1680_p_spl_
  );


  and

  (
    g1687_p,
    g1686_n_spl_,
    g1675_n_spl_
  );


  or

  (
    g1687_n,
    g1686_p_spl_,
    g1675_p_spl_
  );


  and

  (
    g1688_p,
    g1687_n_spl_0,
    g1675_n_spl_
  );


  or

  (
    g1688_n,
    g1687_p_spl_0,
    g1675_p_spl_
  );


  and

  (
    g1689_p,
    g1687_n_spl_0,
    g1686_n_spl_
  );


  or

  (
    g1689_n,
    g1687_p_spl_0,
    g1686_p_spl_
  );


  and

  (
    g1690_p,
    g1689_n,
    g1688_n
  );


  or

  (
    g1690_n,
    g1689_p,
    g1688_p
  );


  and

  (
    g1691_p,
    n7747_o2_p_spl_01,
    n2797_lo_p_spl_100
  );


  or

  (
    g1691_n,
    n7747_o2_n_spl_0,
    n2797_lo_n_spl_100
  );


  and

  (
    g1692_p,
    g1691_n_spl_,
    g1690_n_spl_
  );


  or

  (
    g1692_n,
    g1691_p_spl_,
    g1690_p_spl_
  );


  and

  (
    g1693_p,
    g1692_n_spl_0,
    g1687_n_spl_
  );


  or

  (
    g1693_n,
    g1692_p_spl_0,
    g1687_p_spl_
  );


  and

  (
    g1694_p,
    g1693_n_spl_,
    g1672_n_spl_
  );


  or

  (
    g1694_n,
    g1693_p_spl_,
    g1672_p_spl_
  );


  and

  (
    g1695_p,
    g1694_n_spl_0,
    g1672_n_spl_
  );


  or

  (
    g1695_n,
    g1694_p_spl_0,
    g1672_p_spl_
  );


  and

  (
    g1696_p,
    g1694_n_spl_0,
    g1693_n_spl_
  );


  or

  (
    g1696_n,
    g1694_p_spl_0,
    g1693_p_spl_
  );


  and

  (
    g1697_p,
    g1696_n,
    g1695_n
  );


  or

  (
    g1697_n,
    g1696_p,
    g1695_p
  );


  and

  (
    g1698_p,
    n7747_o2_p_spl_01,
    n2809_lo_p_spl_01
  );


  or

  (
    g1698_n,
    n7747_o2_n_spl_1,
    n2809_lo_n_spl_01
  );


  and

  (
    g1699_p,
    g1698_n_spl_,
    g1697_n_spl_
  );


  or

  (
    g1699_n,
    g1698_p_spl_,
    g1697_p_spl_
  );


  and

  (
    g1700_p,
    g1699_n_spl_0,
    g1697_n_spl_
  );


  or

  (
    g1700_n,
    g1699_p_spl_0,
    g1697_p_spl_
  );


  and

  (
    g1701_p,
    g1699_n_spl_0,
    g1698_n_spl_
  );


  or

  (
    g1701_n,
    g1699_p_spl_0,
    g1698_p_spl_
  );


  and

  (
    g1702_p,
    g1701_n,
    g1700_n
  );


  or

  (
    g1702_n,
    g1701_p,
    g1700_p
  );


  and

  (
    g1703_p,
    g1692_n_spl_0,
    g1690_n_spl_
  );


  or

  (
    g1703_n,
    g1692_p_spl_0,
    g1690_p_spl_
  );


  and

  (
    g1704_p,
    g1692_n_spl_,
    g1691_n_spl_
  );


  or

  (
    g1704_n,
    g1692_p_spl_,
    g1691_p_spl_
  );


  and

  (
    g1705_p,
    g1704_n,
    g1703_n
  );


  or

  (
    g1705_n,
    g1704_p,
    g1703_p
  );


  and

  (
    g1706_p,
    g1685_n_spl_0,
    g1683_n_spl_
  );


  or

  (
    g1706_n,
    g1685_p_spl_0,
    g1683_p_spl_
  );


  and

  (
    g1707_p,
    g1685_n_spl_,
    g1684_n_spl_
  );


  or

  (
    g1707_n,
    g1685_p_spl_,
    g1684_p_spl_
  );


  and

  (
    g1708_p,
    g1707_n,
    g1706_n
  );


  or

  (
    g1708_n,
    g1707_p,
    g1706_p
  );


  and

  (
    g1709_p,
    g1526_n_spl_,
    g1521_n_spl_
  );


  or

  (
    g1709_n,
    g1526_p_spl_,
    g1521_p_spl_
  );


  and

  (
    g1710_p,
    g1709_n_spl_,
    g1708_n_spl_
  );


  or

  (
    g1710_n,
    g1709_p_spl_,
    g1708_p_spl_
  );


  and

  (
    g1711_p,
    g1710_n_spl_0,
    g1708_n_spl_
  );


  or

  (
    g1711_n,
    g1710_p_spl_0,
    g1708_p_spl_
  );


  and

  (
    g1712_p,
    g1710_n_spl_0,
    g1709_n_spl_
  );


  or

  (
    g1712_n,
    g1710_p_spl_0,
    g1709_p_spl_
  );


  and

  (
    g1713_p,
    g1712_n,
    g1711_n
  );


  or

  (
    g1713_n,
    g1712_p,
    g1711_p
  );


  and

  (
    g1714_p,
    n7835_o2_p_spl_0,
    n2797_lo_p_spl_101
  );


  or

  (
    g1714_n,
    n7835_o2_n_spl_0,
    n2797_lo_n_spl_101
  );


  and

  (
    g1715_p,
    g1714_n_spl_,
    g1713_n_spl_
  );


  or

  (
    g1715_n,
    g1714_p_spl_,
    g1713_p_spl_
  );


  and

  (
    g1716_p,
    g1715_n_spl_0,
    g1710_n_spl_
  );


  or

  (
    g1716_n,
    g1715_p_spl_0,
    g1710_p_spl_
  );


  and

  (
    g1717_p,
    g1716_n_spl_,
    g1705_n_spl_
  );


  or

  (
    g1717_n,
    g1716_p_spl_,
    g1705_p_spl_
  );


  and

  (
    g1718_p,
    g1717_n_spl_0,
    g1705_n_spl_
  );


  or

  (
    g1718_n,
    g1717_p_spl_0,
    g1705_p_spl_
  );


  and

  (
    g1719_p,
    g1717_n_spl_0,
    g1716_n_spl_
  );


  or

  (
    g1719_n,
    g1717_p_spl_0,
    g1716_p_spl_
  );


  and

  (
    g1720_p,
    g1719_n,
    g1718_n
  );


  or

  (
    g1720_n,
    g1719_p,
    g1718_p
  );


  and

  (
    g1721_p,
    n7835_o2_p_spl_1,
    n2809_lo_p_spl_01
  );


  or

  (
    g1721_n,
    n7835_o2_n_spl_1,
    n2809_lo_n_spl_01
  );


  and

  (
    g1722_p,
    g1721_n_spl_,
    g1720_n_spl_
  );


  or

  (
    g1722_n,
    g1721_p_spl_,
    g1720_p_spl_
  );


  and

  (
    g1723_p,
    g1722_n_spl_0,
    g1717_n_spl_
  );


  or

  (
    g1723_n,
    g1722_p_spl_0,
    g1717_p_spl_
  );


  or

  (
    g1724_n,
    g1723_p,
    g1702_p
  );


  and

  (
    g1725_p,
    n2716_lo_buf_o2_p_spl_01,
    n2668_lo_buf_o2_p_spl_00
  );


  or

  (
    g1725_n,
    n2716_lo_buf_o2_n_spl_01,
    n2668_lo_buf_o2_n_spl_0
  );


  and

  (
    g1726_p,
    G2030_o2_n,
    G1895_o2_p
  );


  or

  (
    g1726_n,
    G2030_o2_p,
    G1895_o2_n
  );


  and

  (
    g1727_p,
    g1726_n_spl_,
    g1725_n_spl_
  );


  or

  (
    g1727_n,
    g1726_p_spl_,
    g1725_p_spl_
  );


  and

  (
    g1728_p,
    g1727_n_spl_0,
    g1725_n_spl_
  );


  or

  (
    g1728_n,
    g1727_p_spl_0,
    g1725_p_spl_
  );


  and

  (
    g1729_p,
    g1727_n_spl_0,
    g1726_n_spl_
  );


  or

  (
    g1729_n,
    g1727_p_spl_0,
    g1726_p_spl_
  );


  and

  (
    g1730_p,
    g1729_n,
    g1728_n
  );


  or

  (
    g1730_n,
    g1729_p,
    g1728_p
  );


  and

  (
    g1731_p,
    n2728_lo_buf_o2_p_spl_001,
    n2656_lo_buf_o2_p_spl_0
  );


  or

  (
    g1731_n,
    n2728_lo_buf_o2_n_spl_001,
    n2656_lo_buf_o2_n_spl_0
  );


  and

  (
    g1732_p,
    g1731_n_spl_,
    g1730_n_spl_
  );


  or

  (
    g1732_n,
    g1731_p_spl_,
    g1730_p_spl_
  );


  and

  (
    g1733_p,
    g1732_n_spl_0,
    g1730_n_spl_
  );


  or

  (
    g1733_n,
    g1732_p_spl_0,
    g1730_p_spl_
  );


  and

  (
    g1734_p,
    g1732_n_spl_0,
    g1731_n_spl_
  );


  or

  (
    g1734_n,
    g1732_p_spl_0,
    g1731_p_spl_
  );


  and

  (
    g1735_p,
    g1734_n,
    g1733_n
  );


  or

  (
    g1735_n,
    g1734_p,
    g1733_p
  );


  and

  (
    g1736_p,
    G2139_o2_n_spl_,
    G2136_o2_n_spl_
  );


  or

  (
    g1736_n,
    G2139_o2_p_spl_,
    G2136_o2_p_spl_
  );


  and

  (
    g1737_p,
    g1736_n_spl_0,
    G2139_o2_n_spl_
  );


  or

  (
    g1737_n,
    g1736_p_spl_0,
    G2139_o2_p_spl_
  );


  and

  (
    g1738_p,
    g1736_n_spl_0,
    G2136_o2_n_spl_
  );


  or

  (
    g1738_n,
    g1736_p_spl_0,
    G2136_o2_p_spl_
  );


  and

  (
    g1739_p,
    g1738_n,
    g1737_n
  );


  or

  (
    g1739_n,
    g1738_p,
    g1737_p
  );


  and

  (
    g1740_p,
    n2728_lo_buf_o2_p_spl_001,
    n2644_lo_buf_o2_p_spl_0
  );


  or

  (
    g1740_n,
    n2728_lo_buf_o2_n_spl_001,
    n2644_lo_buf_o2_n_spl_0
  );


  and

  (
    g1741_p,
    g1740_n_spl_,
    g1739_n_spl_
  );


  or

  (
    g1741_n,
    g1740_p_spl_,
    g1739_p_spl_
  );


  and

  (
    g1742_p,
    g1741_n_spl_0,
    g1736_n_spl_
  );


  or

  (
    g1742_n,
    g1741_p_spl_0,
    g1736_p_spl_
  );


  and

  (
    g1743_p,
    g1742_n_spl_,
    g1735_n_spl_
  );


  or

  (
    g1743_n,
    g1742_p_spl_,
    g1735_p_spl_
  );


  and

  (
    g1744_p,
    g1743_n_spl_0,
    g1735_n_spl_
  );


  or

  (
    g1744_n,
    g1743_p_spl_0,
    g1735_p_spl_
  );


  and

  (
    g1745_p,
    g1743_n_spl_0,
    g1742_n_spl_
  );


  or

  (
    g1745_n,
    g1743_p_spl_0,
    g1742_p_spl_
  );


  and

  (
    g1746_p,
    g1745_n,
    g1744_n
  );


  or

  (
    g1746_n,
    g1745_p,
    g1744_p
  );


  and

  (
    g1747_p,
    n2644_lo_buf_o2_p_spl_0,
    n2734_lo_p_spl_000
  );


  or

  (
    g1747_n,
    n2644_lo_buf_o2_n_spl_0,
    n2734_lo_n_spl_000
  );


  and

  (
    g1748_p,
    g1747_n_spl_,
    g1746_n_spl_
  );


  or

  (
    g1748_n,
    g1747_p_spl_,
    g1746_p_spl_
  );


  and

  (
    g1749_p,
    g1748_n_spl_0,
    g1746_n_spl_
  );


  or

  (
    g1749_n,
    g1748_p_spl_0,
    g1746_p_spl_
  );


  and

  (
    g1750_p,
    g1748_n_spl_0,
    g1747_n_spl_
  );


  or

  (
    g1750_n,
    g1748_p_spl_0,
    g1747_p_spl_
  );


  and

  (
    g1751_p,
    g1750_n,
    g1749_n
  );


  or

  (
    g1751_n,
    g1750_p,
    g1749_p
  );


  and

  (
    g1752_p,
    g1741_n_spl_0,
    g1739_n_spl_
  );


  or

  (
    g1752_n,
    g1741_p_spl_0,
    g1739_p_spl_
  );


  and

  (
    g1753_p,
    g1741_n_spl_,
    g1740_n_spl_
  );


  or

  (
    g1753_n,
    g1741_p_spl_,
    g1740_p_spl_
  );


  and

  (
    g1754_p,
    g1753_n,
    g1752_n
  );


  or

  (
    g1754_n,
    g1753_p,
    g1752_p
  );


  and

  (
    g1755_p,
    G2313_o2_n,
    G2314_o2_n
  );


  or

  (
    g1755_n,
    G2313_o2_p,
    G2314_o2_p
  );


  and

  (
    g1756_p,
    n2728_lo_buf_o2_p_spl_010,
    n2632_lo_buf_o2_p_spl_0
  );


  or

  (
    g1756_n,
    n2728_lo_buf_o2_n_spl_010,
    n2632_lo_buf_o2_n_spl_0
  );


  and

  (
    g1757_p,
    g1756_n_spl_,
    g1755_n_spl_
  );


  or

  (
    g1757_n,
    g1756_p_spl_,
    g1755_p_spl_
  );


  and

  (
    g1758_p,
    g1757_n_spl_0,
    G2256_o2_p
  );


  or

  (
    g1758_n,
    g1757_p_spl_0,
    G2256_o2_n
  );


  and

  (
    g1759_p,
    g1758_n_spl_,
    g1754_n_spl_
  );


  or

  (
    g1759_n,
    g1758_p_spl_,
    g1754_p_spl_
  );


  and

  (
    g1760_p,
    g1759_n_spl_0,
    g1754_n_spl_
  );


  or

  (
    g1760_n,
    g1759_p_spl_0,
    g1754_p_spl_
  );


  and

  (
    g1761_p,
    g1759_n_spl_0,
    g1758_n_spl_
  );


  or

  (
    g1761_n,
    g1759_p_spl_0,
    g1758_p_spl_
  );


  and

  (
    g1762_p,
    g1761_n,
    g1760_n
  );


  or

  (
    g1762_n,
    g1761_p,
    g1760_p
  );


  and

  (
    g1763_p,
    n2632_lo_buf_o2_p_spl_0,
    n2734_lo_p_spl_001
  );


  or

  (
    g1763_n,
    n2632_lo_buf_o2_n_spl_0,
    n2734_lo_n_spl_001
  );


  and

  (
    g1764_p,
    g1763_n_spl_,
    g1762_n_spl_
  );


  or

  (
    g1764_n,
    g1763_p_spl_,
    g1762_p_spl_
  );


  and

  (
    g1765_p,
    g1764_n_spl_0,
    g1759_n_spl_
  );


  or

  (
    g1765_n,
    g1764_p_spl_0,
    g1759_p_spl_
  );


  and

  (
    g1766_p,
    g1765_n_spl_,
    g1751_n_spl_
  );


  or

  (
    g1766_n,
    g1765_p_spl_,
    g1751_p_spl_
  );


  and

  (
    g1767_p,
    g1766_n_spl_0,
    g1751_n_spl_
  );


  or

  (
    g1767_n,
    g1766_p_spl_0,
    g1751_p_spl_
  );


  and

  (
    g1768_p,
    g1766_n_spl_0,
    g1765_n_spl_
  );


  or

  (
    g1768_n,
    g1766_p_spl_0,
    g1765_p_spl_
  );


  and

  (
    g1769_p,
    g1768_n,
    g1767_n
  );


  or

  (
    g1769_n,
    g1768_p,
    g1767_p
  );


  and

  (
    g1770_p,
    n2632_lo_buf_o2_p_spl_1,
    n2746_lo_p_spl_000
  );


  or

  (
    g1770_n,
    n2632_lo_buf_o2_n_spl_1,
    n2746_lo_n_spl_000
  );


  and

  (
    g1771_p,
    g1770_n_spl_,
    g1769_n_spl_
  );


  or

  (
    g1771_n,
    g1770_p_spl_,
    g1769_p_spl_
  );


  and

  (
    g1772_p,
    g1771_n_spl_0,
    g1769_n_spl_
  );


  or

  (
    g1772_n,
    g1771_p_spl_0,
    g1769_p_spl_
  );


  and

  (
    g1773_p,
    g1771_n_spl_0,
    g1770_n_spl_
  );


  or

  (
    g1773_n,
    g1771_p_spl_0,
    g1770_p_spl_
  );


  and

  (
    g1774_p,
    g1773_n,
    g1772_n
  );


  or

  (
    g1774_n,
    g1773_p,
    g1772_p
  );


  and

  (
    g1775_p,
    g1764_n_spl_0,
    g1762_n_spl_
  );


  or

  (
    g1775_n,
    g1764_p_spl_0,
    g1762_p_spl_
  );


  and

  (
    g1776_p,
    g1764_n_spl_,
    g1763_n_spl_
  );


  or

  (
    g1776_n,
    g1764_p_spl_,
    g1763_p_spl_
  );


  and

  (
    g1777_p,
    g1776_n,
    g1775_n
  );


  or

  (
    g1777_n,
    g1776_p,
    g1775_p
  );


  and

  (
    g1778_p,
    g1757_n_spl_0,
    g1755_n_spl_
  );


  or

  (
    g1778_n,
    g1757_p_spl_0,
    g1755_p_spl_
  );


  and

  (
    g1779_p,
    g1757_n_spl_,
    g1756_n_spl_
  );


  or

  (
    g1779_n,
    g1757_p_spl_,
    g1756_p_spl_
  );


  and

  (
    g1780_p,
    g1779_n,
    g1778_n
  );


  or

  (
    g1780_n,
    g1779_p,
    g1778_p
  );


  and

  (
    g1781_p,
    G2309_o2_p_spl_0,
    G2253_o2_n
  );


  or

  (
    g1781_n,
    G2309_o2_n_spl_0,
    G2253_o2_p
  );


  and

  (
    g1782_p,
    G2309_o2_p_spl_0,
    G2203_o2_n
  );


  or

  (
    g1782_n,
    G2309_o2_n_spl_0,
    G2203_o2_p
  );


  and

  (
    g1783_p,
    g1782_n,
    g1781_n
  );


  or

  (
    g1783_n,
    g1782_p,
    g1781_p
  );


  and

  (
    g1784_p,
    n2728_lo_buf_o2_p_spl_010,
    n2620_lo_buf_o2_p_spl_00
  );


  or

  (
    g1784_n,
    n2728_lo_buf_o2_n_spl_010,
    n2620_lo_buf_o2_n_spl_0
  );


  and

  (
    g1785_p,
    g1784_n_spl_,
    g1783_n_spl_
  );


  or

  (
    g1785_n,
    g1784_p_spl_,
    g1783_p_spl_
  );


  and

  (
    g1786_p,
    g1785_n_spl_0,
    G2309_o2_p_spl_
  );


  or

  (
    g1786_n,
    g1785_p_spl_0,
    G2309_o2_n_spl_
  );


  and

  (
    g1787_p,
    g1786_n_spl_,
    g1780_n_spl_
  );


  or

  (
    g1787_n,
    g1786_p_spl_,
    g1780_p_spl_
  );


  and

  (
    g1788_p,
    g1787_n_spl_0,
    g1780_n_spl_
  );


  or

  (
    g1788_n,
    g1787_p_spl_0,
    g1780_p_spl_
  );


  and

  (
    g1789_p,
    g1787_n_spl_0,
    g1786_n_spl_
  );


  or

  (
    g1789_n,
    g1787_p_spl_0,
    g1786_p_spl_
  );


  and

  (
    g1790_p,
    g1789_n,
    g1788_n
  );


  or

  (
    g1790_n,
    g1789_p,
    g1788_p
  );


  and

  (
    g1791_p,
    n2620_lo_buf_o2_p_spl_00,
    n2734_lo_p_spl_001
  );


  or

  (
    g1791_n,
    n2620_lo_buf_o2_n_spl_0,
    n2734_lo_n_spl_001
  );


  and

  (
    g1792_p,
    g1791_n_spl_,
    g1790_n_spl_
  );


  or

  (
    g1792_n,
    g1791_p_spl_,
    g1790_p_spl_
  );


  and

  (
    g1793_p,
    g1792_n_spl_0,
    g1787_n_spl_
  );


  or

  (
    g1793_n,
    g1792_p_spl_0,
    g1787_p_spl_
  );


  and

  (
    g1794_p,
    g1793_n_spl_,
    g1777_n_spl_
  );


  or

  (
    g1794_n,
    g1793_p_spl_,
    g1777_p_spl_
  );


  and

  (
    g1795_p,
    g1794_n_spl_0,
    g1777_n_spl_
  );


  or

  (
    g1795_n,
    g1794_p_spl_0,
    g1777_p_spl_
  );


  and

  (
    g1796_p,
    g1794_n_spl_0,
    g1793_n_spl_
  );


  or

  (
    g1796_n,
    g1794_p_spl_0,
    g1793_p_spl_
  );


  and

  (
    g1797_p,
    g1796_n,
    g1795_n
  );


  or

  (
    g1797_n,
    g1796_p,
    g1795_p
  );


  and

  (
    g1798_p,
    n2620_lo_buf_o2_p_spl_0,
    n2746_lo_p_spl_000
  );


  or

  (
    g1798_n,
    n2620_lo_buf_o2_n_spl_1,
    n2746_lo_n_spl_000
  );


  and

  (
    g1799_p,
    g1798_n_spl_,
    g1797_n_spl_
  );


  or

  (
    g1799_n,
    g1798_p_spl_,
    g1797_p_spl_
  );


  and

  (
    g1800_p,
    g1799_n_spl_0,
    g1794_n_spl_
  );


  or

  (
    g1800_n,
    g1799_p_spl_0,
    g1794_p_spl_
  );


  and

  (
    g1801_p,
    g1800_n_spl_,
    g1774_n_spl_
  );


  or

  (
    g1801_n,
    g1800_p_spl_,
    g1774_p_spl_
  );


  and

  (
    g1802_p,
    g1293_n_spl_0,
    g1271_n_spl_
  );


  or

  (
    g1802_n,
    g1293_p_spl_,
    g1271_p_spl_
  );


  and

  (
    g1803_p,
    g1293_n_spl_0,
    g1292_n_spl_
  );


  or

  (
    g1803_n,
    g1293_p_spl_,
    g1292_p_spl_
  );


  and

  (
    g1804_p,
    g1803_n,
    g1802_n
  );


  or

  (
    g1804_n,
    g1803_p,
    g1802_p
  );


  and

  (
    g1805_p,
    n7313_o2_p_spl_1,
    n2797_lo_p_spl_101
  );


  or

  (
    g1805_n,
    n7313_o2_n_spl_,
    n2797_lo_n_spl_101
  );


  or

  (
    g1806_n,
    g1805_p,
    g1804_p
  );


  and

  (
    g1807_p,
    g1367_n_spl_0,
    g1345_n_spl_
  );


  or

  (
    g1807_n,
    g1367_p_spl_,
    g1345_p_spl_
  );


  and

  (
    g1808_p,
    g1367_n_spl_0,
    g1366_n_spl_
  );


  or

  (
    g1808_n,
    g1367_p_spl_,
    g1366_p_spl_
  );


  and

  (
    g1809_p,
    g1808_n,
    g1807_n
  );


  or

  (
    g1809_n,
    g1808_p,
    g1807_p
  );


  and

  (
    g1810_p,
    n7501_o2_p_spl_1,
    n2809_lo_p_spl_10
  );


  or

  (
    g1810_n,
    n7501_o2_n_spl_,
    n2809_lo_n_spl_10
  );


  or

  (
    g1811_n,
    g1810_p,
    g1809_p
  );


  and

  (
    g1812_p,
    g1477_n_spl_0,
    g1439_n_spl_
  );


  or

  (
    g1812_n,
    g1477_p_spl_,
    g1439_p_spl_
  );


  and

  (
    g1813_p,
    g1477_n_spl_0,
    g1476_n_spl_
  );


  or

  (
    g1813_n,
    g1477_p_spl_,
    g1476_p_spl_
  );


  and

  (
    g1814_p,
    g1813_n,
    g1812_n
  );


  or

  (
    g1814_n,
    g1813_p,
    g1812_p
  );


  and

  (
    g1815_p,
    n7722_o2_p_spl_1,
    n2821_lo_p_spl_0
  );


  or

  (
    g1815_n,
    n7722_o2_n_spl_1,
    n2821_lo_n_spl_0
  );


  or

  (
    g1816_n,
    g1815_p,
    g1814_p
  );


  and

  (
    g1817_p,
    g1722_n_spl_0,
    g1720_n_spl_
  );


  or

  (
    g1817_n,
    g1722_p_spl_0,
    g1720_p_spl_
  );


  and

  (
    g1818_p,
    g1722_n_spl_,
    g1721_n_spl_
  );


  or

  (
    g1818_n,
    g1722_p_spl_,
    g1721_p_spl_
  );


  and

  (
    g1819_p,
    g1818_n,
    g1817_n
  );


  or

  (
    g1819_n,
    g1818_p,
    g1817_p
  );


  and

  (
    g1820_p,
    g1715_n_spl_0,
    g1713_n_spl_
  );


  or

  (
    g1820_n,
    g1715_p_spl_0,
    g1713_p_spl_
  );


  and

  (
    g1821_p,
    g1715_n_spl_,
    g1714_n_spl_
  );


  or

  (
    g1821_n,
    g1715_p_spl_,
    g1714_p_spl_
  );


  and

  (
    g1822_p,
    g1821_n,
    g1820_n
  );


  or

  (
    g1822_n,
    g1821_p,
    g1820_p
  );


  and

  (
    g1823_p,
    g1536_n_spl_,
    g1531_n_spl_
  );


  or

  (
    g1823_n,
    g1536_p_spl_,
    g1531_p_spl_
  );


  and

  (
    g1824_p,
    g1823_n_spl_,
    g1822_n_spl_
  );


  or

  (
    g1824_n,
    g1823_p_spl_,
    g1822_p_spl_
  );


  and

  (
    g1825_p,
    g1824_n_spl_0,
    g1822_n_spl_
  );


  or

  (
    g1825_n,
    g1824_p_spl_0,
    g1822_p_spl_
  );


  and

  (
    g1826_p,
    g1824_n_spl_0,
    g1823_n_spl_
  );


  or

  (
    g1826_n,
    g1824_p_spl_0,
    g1823_p_spl_
  );


  and

  (
    g1827_p,
    g1826_n,
    g1825_n
  );


  or

  (
    g1827_n,
    g1826_p,
    g1825_p
  );


  and

  (
    g1828_p,
    n7909_o2_p_spl_10,
    n2809_lo_p_spl_10
  );


  or

  (
    g1828_n,
    n7909_o2_n_spl_1,
    n2809_lo_n_spl_10
  );


  and

  (
    g1829_p,
    g1828_n_spl_,
    g1827_n_spl_
  );


  or

  (
    g1829_n,
    g1828_p_spl_,
    g1827_p_spl_
  );


  and

  (
    g1830_p,
    g1829_n_spl_0,
    g1824_n_spl_
  );


  or

  (
    g1830_n,
    g1829_p_spl_0,
    g1824_p_spl_
  );


  or

  (
    g1831_n,
    g1830_p,
    g1819_p
  );


  or

  (
    g1832_n,
    n2488_lo_buf_o2_n_spl_1,
    n2746_lo_n_spl_001
  );


  and

  (
    g1833_p,
    G19_p_spl_000,
    G16_p_spl_0
  );


  or

  (
    g1833_n,
    G19_n_spl_000,
    G16_n_spl_0
  );


  and

  (
    g1834_p,
    G18_p_spl_000,
    G16_p_spl_0
  );


  or

  (
    g1834_n,
    G18_n_spl_000,
    G16_n_spl_0
  );


  and

  (
    g1835_p,
    G17_p_spl_000,
    G16_p_spl_1
  );


  or

  (
    g1835_n,
    G17_n_spl_000,
    G16_n_spl_
  );


  and

  (
    g1836_p,
    G18_p_spl_000,
    G15_p_spl_00
  );


  or

  (
    g1836_n,
    G18_n_spl_000,
    G15_n_spl_0
  );


  and

  (
    g1837_p,
    g1836_n_spl_,
    g1835_p_spl_
  );


  or

  (
    g1837_n,
    g1836_p_spl_,
    g1835_n_spl_
  );


  and

  (
    g1838_p,
    g1837_n_spl_,
    g1835_p_spl_
  );


  or

  (
    g1838_n,
    g1837_p_spl_,
    g1835_n_spl_
  );


  and

  (
    g1839_p,
    g1838_n_spl_0,
    g1834_n_spl_
  );


  or

  (
    g1839_n,
    g1838_p_spl_0,
    g1834_p_spl_
  );


  and

  (
    g1840_p,
    g1839_n_spl_0,
    g1834_n_spl_
  );


  or

  (
    g1840_n,
    g1839_p_spl_0,
    g1834_p_spl_
  );


  and

  (
    g1841_p,
    g1839_n_spl_0,
    g1838_n_spl_0
  );


  or

  (
    g1841_n,
    g1839_p_spl_0,
    g1838_p_spl_0
  );


  and

  (
    g1842_p,
    g1841_n,
    g1840_n
  );


  or

  (
    g1842_n,
    g1841_p,
    g1840_p
  );


  and

  (
    g1843_p,
    G19_p_spl_000,
    G15_p_spl_00
  );


  or

  (
    g1843_n,
    G19_n_spl_000,
    G15_n_spl_0
  );


  and

  (
    g1844_p,
    g1843_n_spl_,
    g1842_n_spl_
  );


  or

  (
    g1844_n,
    g1843_p_spl_,
    g1842_p_spl_
  );


  and

  (
    g1845_p,
    g1844_n_spl_0,
    g1839_n_spl_
  );


  or

  (
    g1845_n,
    g1844_p_spl_0,
    g1839_p_spl_
  );


  and

  (
    g1846_p,
    g1845_n_spl_,
    g1833_n_spl_
  );


  or

  (
    g1846_n,
    g1845_p_spl_,
    g1833_p_spl_
  );


  and

  (
    g1847_p,
    n2728_lo_buf_o2_p_spl_011,
    n2668_lo_buf_o2_p_spl_00
  );


  or

  (
    g1847_n,
    n2728_lo_buf_o2_n_spl_011,
    n2668_lo_buf_o2_n_spl_0
  );


  and

  (
    g1848_p,
    g1732_n_spl_,
    g1727_n_spl_
  );


  or

  (
    g1848_n,
    g1732_p_spl_,
    g1727_p_spl_
  );


  and

  (
    g1849_p,
    g1848_n_spl_,
    g1847_n_spl_
  );


  or

  (
    g1849_n,
    g1848_p_spl_,
    g1847_p_spl_
  );


  and

  (
    g1850_p,
    g1849_n_spl_0,
    g1847_n_spl_
  );


  or

  (
    g1850_n,
    g1849_p_spl_0,
    g1847_p_spl_
  );


  and

  (
    g1851_p,
    g1849_n_spl_0,
    g1848_n_spl_
  );


  or

  (
    g1851_n,
    g1849_p_spl_0,
    g1848_p_spl_
  );


  and

  (
    g1852_p,
    g1851_n,
    g1850_n
  );


  or

  (
    g1852_n,
    g1851_p,
    g1850_p
  );


  and

  (
    g1853_p,
    n2656_lo_buf_o2_p_spl_0,
    n2734_lo_p_spl_010
  );


  or

  (
    g1853_n,
    n2656_lo_buf_o2_n_spl_0,
    n2734_lo_n_spl_010
  );


  and

  (
    g1854_p,
    g1853_n_spl_,
    g1852_n_spl_
  );


  or

  (
    g1854_n,
    g1853_p_spl_,
    g1852_p_spl_
  );


  and

  (
    g1855_p,
    g1854_n_spl_0,
    g1852_n_spl_
  );


  or

  (
    g1855_n,
    g1854_p_spl_0,
    g1852_p_spl_
  );


  and

  (
    g1856_p,
    g1854_n_spl_0,
    g1853_n_spl_
  );


  or

  (
    g1856_n,
    g1854_p_spl_0,
    g1853_p_spl_
  );


  and

  (
    g1857_p,
    g1856_n,
    g1855_n
  );


  or

  (
    g1857_n,
    g1856_p,
    g1855_p
  );


  and

  (
    g1858_p,
    g1748_n_spl_,
    g1743_n_spl_
  );


  or

  (
    g1858_n,
    g1748_p_spl_,
    g1743_p_spl_
  );


  and

  (
    g1859_p,
    g1858_n_spl_,
    g1857_n_spl_
  );


  or

  (
    g1859_n,
    g1858_p_spl_,
    g1857_p_spl_
  );


  and

  (
    g1860_p,
    g1859_n_spl_0,
    g1857_n_spl_
  );


  or

  (
    g1860_n,
    g1859_p_spl_0,
    g1857_p_spl_
  );


  and

  (
    g1861_p,
    g1859_n_spl_0,
    g1858_n_spl_
  );


  or

  (
    g1861_n,
    g1859_p_spl_0,
    g1858_p_spl_
  );


  and

  (
    g1862_p,
    g1861_n,
    g1860_n
  );


  or

  (
    g1862_n,
    g1861_p,
    g1860_p
  );


  and

  (
    g1863_p,
    n2644_lo_buf_o2_p_spl_1,
    n2746_lo_p_spl_001
  );


  or

  (
    g1863_n,
    n2644_lo_buf_o2_n_spl_,
    n2746_lo_n_spl_001
  );


  and

  (
    g1864_p,
    g1863_n_spl_,
    g1862_n_spl_
  );


  or

  (
    g1864_n,
    g1863_p_spl_,
    g1862_p_spl_
  );


  and

  (
    g1865_p,
    g1864_n_spl_0,
    g1862_n_spl_
  );


  or

  (
    g1865_n,
    g1864_p_spl_0,
    g1862_p_spl_
  );


  and

  (
    g1866_p,
    g1864_n_spl_0,
    g1863_n_spl_
  );


  or

  (
    g1866_n,
    g1864_p_spl_0,
    g1863_p_spl_
  );


  and

  (
    g1867_p,
    g1866_n,
    g1865_n
  );


  or

  (
    g1867_n,
    g1866_p,
    g1865_p
  );


  and

  (
    g1868_p,
    g1771_n_spl_,
    g1766_n_spl_
  );


  or

  (
    g1868_n,
    g1771_p_spl_,
    g1766_p_spl_
  );


  or

  (
    g1869_n,
    g1868_p,
    g1867_p
  );


  and

  (
    g1870_p,
    G2015_o2_n,
    G2016_o2_n
  );


  or

  (
    g1870_n,
    G2015_o2_p,
    G2016_o2_p
  );


  and

  (
    g1871_p,
    n2716_lo_buf_o2_p_spl_01,
    n2572_lo_buf_o2_p_spl_00
  );


  or

  (
    g1871_n,
    n2716_lo_buf_o2_n_spl_01,
    n2572_lo_buf_o2_n_spl_00
  );


  and

  (
    g1872_p,
    g1871_n_spl_,
    g1870_n_spl_
  );


  or

  (
    g1872_n,
    g1871_p_spl_,
    g1870_p_spl_
  );


  and

  (
    g1873_p,
    g1872_n_spl_0,
    g1870_n_spl_
  );


  or

  (
    g1873_n,
    g1872_p_spl_0,
    g1870_p_spl_
  );


  and

  (
    g1874_p,
    g1872_n_spl_0,
    g1871_n_spl_
  );


  or

  (
    g1874_n,
    g1872_p_spl_0,
    g1871_p_spl_
  );


  and

  (
    g1875_p,
    g1874_n,
    g1873_n
  );


  or

  (
    g1875_n,
    g1874_p,
    g1873_p
  );


  and

  (
    g1876_p,
    G1968_o2_p_spl_0,
    G1917_o2_n
  );


  or

  (
    g1876_n,
    G1968_o2_n_spl_0,
    G1917_o2_p
  );


  and

  (
    g1877_p,
    G1968_o2_p_spl_0,
    G1854_o2_n
  );


  or

  (
    g1877_n,
    G1968_o2_n_spl_0,
    G1854_o2_p
  );


  and

  (
    g1878_p,
    g1877_n,
    g1876_n
  );


  or

  (
    g1878_n,
    g1877_p,
    g1876_p
  );


  and

  (
    g1879_p,
    n2716_lo_buf_o2_p_spl_10,
    n2560_lo_buf_o2_p_spl_00
  );


  or

  (
    g1879_n,
    n2716_lo_buf_o2_n_spl_10,
    n2560_lo_buf_o2_n_spl_00
  );


  and

  (
    g1880_p,
    g1879_n_spl_,
    g1878_n_spl_
  );


  or

  (
    g1880_n,
    g1879_p_spl_,
    g1878_p_spl_
  );


  and

  (
    g1881_p,
    g1880_n_spl_0,
    G1968_o2_p_spl_
  );


  or

  (
    g1881_n,
    g1880_p_spl_0,
    G1968_o2_n_spl_
  );


  and

  (
    g1882_p,
    g1881_n_spl_,
    g1875_n_spl_
  );


  or

  (
    g1882_n,
    g1881_p_spl_,
    g1875_p_spl_
  );


  and

  (
    g1883_p,
    g1882_n_spl_0,
    g1875_n_spl_
  );


  or

  (
    g1883_n,
    g1882_p_spl_0,
    g1875_p_spl_
  );


  and

  (
    g1884_p,
    g1882_n_spl_0,
    g1881_n_spl_
  );


  or

  (
    g1884_n,
    g1882_p_spl_0,
    g1881_p_spl_
  );


  and

  (
    g1885_p,
    g1884_n,
    g1883_n
  );


  or

  (
    g1885_n,
    g1884_p,
    g1883_p
  );


  and

  (
    g1886_p,
    n2728_lo_buf_o2_p_spl_011,
    n2560_lo_buf_o2_p_spl_00
  );


  or

  (
    g1886_n,
    n2728_lo_buf_o2_n_spl_011,
    n2560_lo_buf_o2_n_spl_00
  );


  and

  (
    g1887_p,
    g1886_n_spl_,
    g1885_n_spl_
  );


  or

  (
    g1887_n,
    g1886_p_spl_,
    g1885_p_spl_
  );


  and

  (
    g1888_p,
    g1887_n_spl_0,
    g1885_n_spl_
  );


  or

  (
    g1888_n,
    g1887_p_spl_0,
    g1885_p_spl_
  );


  and

  (
    g1889_p,
    g1887_n_spl_0,
    g1886_n_spl_
  );


  or

  (
    g1889_n,
    g1887_p_spl_0,
    g1886_p_spl_
  );


  and

  (
    g1890_p,
    g1889_n,
    g1888_n
  );


  or

  (
    g1890_n,
    g1889_p,
    g1888_p
  );


  and

  (
    g1891_p,
    g1880_n_spl_0,
    g1878_n_spl_
  );


  or

  (
    g1891_n,
    g1880_p_spl_0,
    g1878_p_spl_
  );


  and

  (
    g1892_p,
    g1880_n_spl_,
    g1879_n_spl_
  );


  or

  (
    g1892_n,
    g1880_p_spl_,
    g1879_p_spl_
  );


  and

  (
    g1893_p,
    g1892_n,
    g1891_n
  );


  or

  (
    g1893_n,
    g1892_p,
    g1891_p
  );


  and

  (
    g1894_p,
    G1914_o2_n_spl_,
    G1849_o2_n_spl_
  );


  or

  (
    g1894_n,
    G1914_o2_p_spl_,
    G1849_o2_p_spl_
  );


  and

  (
    g1895_p,
    g1894_n_spl_0,
    G1914_o2_n_spl_
  );


  or

  (
    g1895_n,
    g1894_p_spl_0,
    G1914_o2_p_spl_
  );


  and

  (
    g1896_p,
    g1894_n_spl_0,
    G1849_o2_n_spl_
  );


  or

  (
    g1896_n,
    g1894_p_spl_0,
    G1849_o2_p_spl_
  );


  and

  (
    g1897_p,
    g1896_n,
    g1895_n
  );


  or

  (
    g1897_n,
    g1896_p,
    g1895_p
  );


  and

  (
    g1898_p,
    n2716_lo_buf_o2_p_spl_10,
    n2548_lo_buf_o2_p_spl_00
  );


  or

  (
    g1898_n,
    n2716_lo_buf_o2_n_spl_10,
    n2548_lo_buf_o2_n_spl_00
  );


  and

  (
    g1899_p,
    g1898_n_spl_,
    g1897_n_spl_
  );


  or

  (
    g1899_n,
    g1898_p_spl_,
    g1897_p_spl_
  );


  and

  (
    g1900_p,
    g1899_n_spl_0,
    g1894_n_spl_
  );


  or

  (
    g1900_n,
    g1899_p_spl_0,
    g1894_p_spl_
  );


  and

  (
    g1901_p,
    g1900_n_spl_,
    g1893_n_spl_
  );


  or

  (
    g1901_n,
    g1900_p_spl_,
    g1893_p_spl_
  );


  and

  (
    g1902_p,
    g1901_n_spl_0,
    g1893_n_spl_
  );


  or

  (
    g1902_n,
    g1901_p_spl_0,
    g1893_p_spl_
  );


  and

  (
    g1903_p,
    g1901_n_spl_0,
    g1900_n_spl_
  );


  or

  (
    g1903_n,
    g1901_p_spl_0,
    g1900_p_spl_
  );


  and

  (
    g1904_p,
    g1903_n,
    g1902_n
  );


  or

  (
    g1904_n,
    g1903_p,
    g1902_p
  );


  and

  (
    g1905_p,
    n2728_lo_buf_o2_p_spl_100,
    n2548_lo_buf_o2_p_spl_00
  );


  or

  (
    g1905_n,
    n2728_lo_buf_o2_n_spl_100,
    n2548_lo_buf_o2_n_spl_00
  );


  and

  (
    g1906_p,
    g1905_n_spl_,
    g1904_n_spl_
  );


  or

  (
    g1906_n,
    g1905_p_spl_,
    g1904_p_spl_
  );


  and

  (
    g1907_p,
    g1906_n_spl_0,
    g1901_n_spl_
  );


  or

  (
    g1907_n,
    g1906_p_spl_0,
    g1901_p_spl_
  );


  and

  (
    g1908_p,
    g1907_n_spl_,
    g1890_n_spl_
  );


  or

  (
    g1908_n,
    g1907_p_spl_,
    g1890_p_spl_
  );


  and

  (
    g1909_p,
    g1908_n_spl_0,
    g1890_n_spl_
  );


  or

  (
    g1909_n,
    g1908_p_spl_0,
    g1890_p_spl_
  );


  and

  (
    g1910_p,
    g1908_n_spl_0,
    g1907_n_spl_
  );


  or

  (
    g1910_n,
    g1908_p_spl_0,
    g1907_p_spl_
  );


  and

  (
    g1911_p,
    g1910_n,
    g1909_n
  );


  or

  (
    g1911_n,
    g1910_p,
    g1909_p
  );


  and

  (
    g1912_p,
    n2548_lo_buf_o2_p_spl_01,
    n2734_lo_p_spl_010
  );


  or

  (
    g1912_n,
    n2548_lo_buf_o2_n_spl_0,
    n2734_lo_n_spl_010
  );


  and

  (
    g1913_p,
    g1912_n_spl_,
    g1911_n_spl_
  );


  or

  (
    g1913_n,
    g1912_p_spl_,
    g1911_p_spl_
  );


  and

  (
    g1914_p,
    g1913_n_spl_0,
    g1911_n_spl_
  );


  or

  (
    g1914_n,
    g1913_p_spl_0,
    g1911_p_spl_
  );


  and

  (
    g1915_p,
    g1913_n_spl_0,
    g1912_n_spl_
  );


  or

  (
    g1915_n,
    g1913_p_spl_0,
    g1912_p_spl_
  );


  and

  (
    g1916_p,
    g1915_n,
    g1914_n
  );


  or

  (
    g1916_n,
    g1915_p,
    g1914_p
  );


  and

  (
    g1917_p,
    g1906_n_spl_0,
    g1904_n_spl_
  );


  or

  (
    g1917_n,
    g1906_p_spl_0,
    g1904_p_spl_
  );


  and

  (
    g1918_p,
    g1906_n_spl_,
    g1905_n_spl_
  );


  or

  (
    g1918_n,
    g1906_p_spl_,
    g1905_p_spl_
  );


  and

  (
    g1919_p,
    g1918_n,
    g1917_n
  );


  or

  (
    g1919_n,
    g1918_p,
    g1917_p
  );


  and

  (
    g1920_p,
    g1899_n_spl_0,
    g1897_n_spl_
  );


  or

  (
    g1920_n,
    g1899_p_spl_0,
    g1897_p_spl_
  );


  and

  (
    g1921_p,
    g1899_n_spl_,
    g1898_n_spl_
  );


  or

  (
    g1921_n,
    g1899_p_spl_,
    g1898_p_spl_
  );


  and

  (
    g1922_p,
    g1921_n,
    g1920_n
  );


  or

  (
    g1922_n,
    g1921_p,
    g1920_p
  );


  and

  (
    g1923_p,
    G1847_o2_n,
    G1848_o2_p
  );


  or

  (
    g1923_n,
    G1847_o2_p,
    G1848_o2_n
  );


  and

  (
    g1924_p,
    G1777_o2_n_spl_0,
    G1642_o2_p
  );


  or

  (
    g1924_n,
    G1777_o2_p_spl_0,
    G1642_o2_n
  );


  and

  (
    g1925_p,
    g1924_n_spl_,
    g1923_n_spl_
  );


  or

  (
    g1925_n,
    g1924_p_spl_,
    g1923_p_spl_
  );


  and

  (
    g1926_p,
    g1925_n_spl_0,
    g1923_n_spl_
  );


  or

  (
    g1926_n,
    g1925_p_spl_0,
    g1923_p_spl_
  );


  and

  (
    g1927_p,
    g1925_n_spl_0,
    g1924_n_spl_
  );


  or

  (
    g1927_n,
    g1925_p_spl_0,
    g1924_p_spl_
  );


  and

  (
    g1928_p,
    g1927_n,
    g1926_n
  );


  or

  (
    g1928_n,
    g1927_p,
    g1926_p
  );


  and

  (
    g1929_p,
    n2716_lo_buf_o2_p_spl_11,
    n2536_lo_buf_o2_p_spl_00
  );


  or

  (
    g1929_n,
    n2716_lo_buf_o2_n_spl_11,
    n2536_lo_buf_o2_n_spl_00
  );


  and

  (
    g1930_p,
    g1929_n_spl_,
    g1928_n_spl_
  );


  or

  (
    g1930_n,
    g1929_p_spl_,
    g1928_p_spl_
  );


  and

  (
    g1931_p,
    g1930_n_spl_0,
    g1925_n_spl_
  );


  or

  (
    g1931_n,
    g1930_p_spl_0,
    g1925_p_spl_
  );


  and

  (
    g1932_p,
    g1931_n_spl_,
    g1922_n_spl_
  );


  or

  (
    g1932_n,
    g1931_p_spl_,
    g1922_p_spl_
  );


  and

  (
    g1933_p,
    g1932_n_spl_0,
    g1922_n_spl_
  );


  or

  (
    g1933_n,
    g1932_p_spl_0,
    g1922_p_spl_
  );


  and

  (
    g1934_p,
    g1932_n_spl_0,
    g1931_n_spl_
  );


  or

  (
    g1934_n,
    g1932_p_spl_0,
    g1931_p_spl_
  );


  and

  (
    g1935_p,
    g1934_n,
    g1933_n
  );


  or

  (
    g1935_n,
    g1934_p,
    g1933_p
  );


  and

  (
    g1936_p,
    n2728_lo_buf_o2_p_spl_100,
    n2536_lo_buf_o2_p_spl_00
  );


  or

  (
    g1936_n,
    n2728_lo_buf_o2_n_spl_100,
    n2536_lo_buf_o2_n_spl_00
  );


  and

  (
    g1937_p,
    g1936_n_spl_,
    g1935_n_spl_
  );


  or

  (
    g1937_n,
    g1936_p_spl_,
    g1935_p_spl_
  );


  and

  (
    g1938_p,
    g1937_n_spl_0,
    g1932_n_spl_
  );


  or

  (
    g1938_n,
    g1937_p_spl_0,
    g1932_p_spl_
  );


  and

  (
    g1939_p,
    g1938_n_spl_,
    g1919_n_spl_
  );


  or

  (
    g1939_n,
    g1938_p_spl_,
    g1919_p_spl_
  );


  and

  (
    g1940_p,
    g1939_n_spl_0,
    g1919_n_spl_
  );


  or

  (
    g1940_n,
    g1939_p_spl_0,
    g1919_p_spl_
  );


  and

  (
    g1941_p,
    g1939_n_spl_0,
    g1938_n_spl_
  );


  or

  (
    g1941_n,
    g1939_p_spl_0,
    g1938_p_spl_
  );


  and

  (
    g1942_p,
    g1941_n,
    g1940_n
  );


  or

  (
    g1942_n,
    g1941_p,
    g1940_p
  );


  and

  (
    g1943_p,
    n2536_lo_buf_o2_p_spl_01,
    n2734_lo_p_spl_011
  );


  or

  (
    g1943_n,
    n2536_lo_buf_o2_n_spl_0,
    n2734_lo_n_spl_011
  );


  and

  (
    g1944_p,
    g1943_n_spl_,
    g1942_n_spl_
  );


  or

  (
    g1944_n,
    g1943_p_spl_,
    g1942_p_spl_
  );


  and

  (
    g1945_p,
    g1944_n_spl_0,
    g1939_n_spl_
  );


  or

  (
    g1945_n,
    g1944_p_spl_0,
    g1939_p_spl_
  );


  and

  (
    g1946_p,
    g1945_n_spl_,
    g1916_n_spl_
  );


  or

  (
    g1946_n,
    g1945_p_spl_,
    g1916_p_spl_
  );


  and

  (
    g1947_p,
    g1946_n_spl_0,
    g1916_n_spl_
  );


  or

  (
    g1947_n,
    g1946_p_spl_0,
    g1916_p_spl_
  );


  and

  (
    g1948_p,
    g1946_n_spl_0,
    g1945_n_spl_
  );


  or

  (
    g1948_n,
    g1946_p_spl_0,
    g1945_p_spl_
  );


  and

  (
    g1949_p,
    g1948_n,
    g1947_n
  );


  or

  (
    g1949_n,
    g1948_p,
    g1947_p
  );


  and

  (
    g1950_p,
    n2536_lo_buf_o2_p_spl_01,
    n2746_lo_p_spl_001
  );


  or

  (
    g1950_n,
    n2536_lo_buf_o2_n_spl_1,
    n2746_lo_n_spl_010
  );


  and

  (
    g1951_p,
    g1950_n_spl_,
    g1949_n_spl_
  );


  or

  (
    g1951_n,
    g1950_p_spl_,
    g1949_p_spl_
  );


  and

  (
    g1952_p,
    g1951_n_spl_0,
    g1949_n_spl_
  );


  or

  (
    g1952_n,
    g1951_p_spl_0,
    g1949_p_spl_
  );


  and

  (
    g1953_p,
    g1951_n_spl_0,
    g1950_n_spl_
  );


  or

  (
    g1953_n,
    g1951_p_spl_0,
    g1950_p_spl_
  );


  and

  (
    g1954_p,
    g1953_n,
    g1952_n
  );


  or

  (
    g1954_n,
    g1953_p,
    g1952_p
  );


  and

  (
    g1955_p,
    g1944_n_spl_0,
    g1942_n_spl_
  );


  or

  (
    g1955_n,
    g1944_p_spl_0,
    g1942_p_spl_
  );


  and

  (
    g1956_p,
    g1944_n_spl_,
    g1943_n_spl_
  );


  or

  (
    g1956_n,
    g1944_p_spl_,
    g1943_p_spl_
  );


  and

  (
    g1957_p,
    g1956_n,
    g1955_n
  );


  or

  (
    g1957_n,
    g1956_p,
    g1955_p
  );


  and

  (
    g1958_p,
    g1937_n_spl_0,
    g1935_n_spl_
  );


  or

  (
    g1958_n,
    g1937_p_spl_0,
    g1935_p_spl_
  );


  and

  (
    g1959_p,
    g1937_n_spl_,
    g1936_n_spl_
  );


  or

  (
    g1959_n,
    g1937_p_spl_,
    g1936_p_spl_
  );


  and

  (
    g1960_p,
    g1959_n,
    g1958_n
  );


  or

  (
    g1960_n,
    g1959_p,
    g1958_p
  );


  and

  (
    g1961_p,
    g1930_n_spl_0,
    g1928_n_spl_
  );


  or

  (
    g1961_n,
    g1930_p_spl_0,
    g1928_p_spl_
  );


  and

  (
    g1962_p,
    g1930_n_spl_,
    g1929_n_spl_
  );


  or

  (
    g1962_n,
    g1930_p_spl_,
    g1929_p_spl_
  );


  and

  (
    g1963_p,
    g1962_n,
    g1961_n
  );


  or

  (
    g1963_n,
    g1962_p,
    g1961_p
  );


  and

  (
    g1964_p,
    G1777_o2_n_spl_0,
    G1727_o2_p
  );


  or

  (
    g1964_n,
    G1777_o2_p_spl_0,
    G1727_o2_n
  );


  and

  (
    g1965_p,
    G1777_o2_n_spl_,
    G740_o2_n
  );


  or

  (
    g1965_n,
    G1777_o2_p_spl_,
    G740_o2_p
  );


  and

  (
    g1966_p,
    g1965_n,
    g1964_n
  );


  or

  (
    g1966_n,
    g1965_p,
    g1964_p
  );


  and

  (
    g1967_p,
    g1478_n_spl_,
    G1638_o2_p
  );


  or

  (
    g1967_n,
    g1478_p_spl_,
    G1638_o2_n
  );


  and

  (
    g1968_p,
    g1967_n_spl_,
    g1966_n_spl_
  );


  or

  (
    g1968_n,
    g1967_p_spl_,
    g1966_p_spl_
  );


  and

  (
    g1969_p,
    g1968_n_spl_0,
    g1966_n_spl_
  );


  or

  (
    g1969_n,
    g1968_p_spl_0,
    g1966_p_spl_
  );


  and

  (
    g1970_p,
    g1968_n_spl_0,
    g1967_n_spl_
  );


  or

  (
    g1970_n,
    g1968_p_spl_0,
    g1967_p_spl_
  );


  and

  (
    g1971_p,
    g1970_n,
    g1969_n
  );


  or

  (
    g1971_n,
    g1970_p,
    g1969_p
  );


  and

  (
    g1972_p,
    n2716_lo_buf_o2_p_spl_11,
    n2524_lo_buf_o2_p_spl_00
  );


  or

  (
    g1972_n,
    n2716_lo_buf_o2_n_spl_11,
    n2524_lo_buf_o2_n_spl_00
  );


  and

  (
    g1973_p,
    g1972_n_spl_,
    g1971_n_spl_
  );


  or

  (
    g1973_n,
    g1972_p_spl_,
    g1971_p_spl_
  );


  and

  (
    g1974_p,
    g1973_n_spl_0,
    g1968_n_spl_
  );


  or

  (
    g1974_n,
    g1973_p_spl_0,
    g1968_p_spl_
  );


  and

  (
    g1975_p,
    g1974_n_spl_,
    g1963_n_spl_
  );


  or

  (
    g1975_n,
    g1974_p_spl_,
    g1963_p_spl_
  );


  and

  (
    g1976_p,
    g1975_n_spl_0,
    g1963_n_spl_
  );


  or

  (
    g1976_n,
    g1975_p_spl_0,
    g1963_p_spl_
  );


  and

  (
    g1977_p,
    g1975_n_spl_0,
    g1974_n_spl_
  );


  or

  (
    g1977_n,
    g1975_p_spl_0,
    g1974_p_spl_
  );


  and

  (
    g1978_p,
    g1977_n,
    g1976_n
  );


  or

  (
    g1978_n,
    g1977_p,
    g1976_p
  );


  and

  (
    g1979_p,
    n2728_lo_buf_o2_p_spl_101,
    n2524_lo_buf_o2_p_spl_00
  );


  or

  (
    g1979_n,
    n2728_lo_buf_o2_n_spl_101,
    n2524_lo_buf_o2_n_spl_00
  );


  and

  (
    g1980_p,
    g1979_n_spl_,
    g1978_n_spl_
  );


  or

  (
    g1980_n,
    g1979_p_spl_,
    g1978_p_spl_
  );


  and

  (
    g1981_p,
    g1980_n_spl_0,
    g1975_n_spl_
  );


  or

  (
    g1981_n,
    g1980_p_spl_0,
    g1975_p_spl_
  );


  and

  (
    g1982_p,
    g1981_n_spl_,
    g1960_n_spl_
  );


  or

  (
    g1982_n,
    g1981_p_spl_,
    g1960_p_spl_
  );


  and

  (
    g1983_p,
    g1982_n_spl_0,
    g1960_n_spl_
  );


  or

  (
    g1983_n,
    g1982_p_spl_0,
    g1960_p_spl_
  );


  and

  (
    g1984_p,
    g1982_n_spl_0,
    g1981_n_spl_
  );


  or

  (
    g1984_n,
    g1982_p_spl_0,
    g1981_p_spl_
  );


  and

  (
    g1985_p,
    g1984_n,
    g1983_n
  );


  or

  (
    g1985_n,
    g1984_p,
    g1983_p
  );


  and

  (
    g1986_p,
    n2524_lo_buf_o2_p_spl_0,
    n2734_lo_p_spl_011
  );


  or

  (
    g1986_n,
    n2524_lo_buf_o2_n_spl_0,
    n2734_lo_n_spl_011
  );


  and

  (
    g1987_p,
    g1986_n_spl_,
    g1985_n_spl_
  );


  or

  (
    g1987_n,
    g1986_p_spl_,
    g1985_p_spl_
  );


  and

  (
    g1988_p,
    g1987_n_spl_0,
    g1982_n_spl_
  );


  or

  (
    g1988_n,
    g1987_p_spl_0,
    g1982_p_spl_
  );


  and

  (
    g1989_p,
    g1988_n_spl_,
    g1957_n_spl_
  );


  or

  (
    g1989_n,
    g1988_p_spl_,
    g1957_p_spl_
  );


  and

  (
    g1990_p,
    g1989_n_spl_0,
    g1957_n_spl_
  );


  or

  (
    g1990_n,
    g1989_p_spl_0,
    g1957_p_spl_
  );


  and

  (
    g1991_p,
    g1989_n_spl_0,
    g1988_n_spl_
  );


  or

  (
    g1991_n,
    g1989_p_spl_0,
    g1988_p_spl_
  );


  and

  (
    g1992_p,
    g1991_n,
    g1990_n
  );


  or

  (
    g1992_n,
    g1991_p,
    g1990_p
  );


  and

  (
    g1993_p,
    n2524_lo_buf_o2_p_spl_1,
    n2746_lo_p_spl_010
  );


  or

  (
    g1993_n,
    n2524_lo_buf_o2_n_spl_1,
    n2746_lo_n_spl_010
  );


  and

  (
    g1994_p,
    g1993_n_spl_,
    g1992_n_spl_
  );


  or

  (
    g1994_n,
    g1993_p_spl_,
    g1992_p_spl_
  );


  and

  (
    g1995_p,
    g1994_n_spl_0,
    g1989_n_spl_
  );


  or

  (
    g1995_n,
    g1994_p_spl_0,
    g1989_p_spl_
  );


  or

  (
    g1996_n,
    g1995_p,
    g1954_p
  );


  and

  (
    g1997_p,
    g1792_n_spl_0,
    g1790_n_spl_
  );


  or

  (
    g1997_n,
    g1792_p_spl_0,
    g1790_p_spl_
  );


  and

  (
    g1998_p,
    g1792_n_spl_,
    g1791_n_spl_
  );


  or

  (
    g1998_n,
    g1792_p_spl_,
    g1791_p_spl_
  );


  and

  (
    g1999_p,
    g1998_n,
    g1997_n
  );


  or

  (
    g1999_n,
    g1998_p,
    g1997_p
  );


  and

  (
    g2000_p,
    g1785_n_spl_0,
    g1783_n_spl_
  );


  or

  (
    g2000_n,
    g1785_p_spl_0,
    g1783_p_spl_
  );


  and

  (
    g2001_p,
    g1785_n_spl_,
    g1784_n_spl_
  );


  or

  (
    g2001_n,
    g1785_p_spl_,
    g1784_p_spl_
  );


  and

  (
    g2002_p,
    g2001_n,
    g2000_n
  );


  or

  (
    g2002_n,
    g2001_p,
    g2000_p
  );


  and

  (
    g2003_p,
    G2250_o2_n_spl_,
    G2198_o2_n_spl_
  );


  or

  (
    g2003_n,
    G2250_o2_p_spl_,
    G2198_o2_p_spl_
  );


  and

  (
    g2004_p,
    g2003_n_spl_0,
    G2250_o2_n_spl_
  );


  or

  (
    g2004_n,
    g2003_p_spl_0,
    G2250_o2_p_spl_
  );


  and

  (
    g2005_p,
    g2003_n_spl_0,
    G2198_o2_n_spl_
  );


  or

  (
    g2005_n,
    g2003_p_spl_0,
    G2198_o2_p_spl_
  );


  and

  (
    g2006_p,
    g2005_n,
    g2004_n
  );


  or

  (
    g2006_n,
    g2005_p,
    g2004_p
  );


  and

  (
    g2007_p,
    n2728_lo_buf_o2_p_spl_101,
    n2608_lo_buf_o2_p_spl_00
  );


  or

  (
    g2007_n,
    n2728_lo_buf_o2_n_spl_101,
    n2608_lo_buf_o2_n_spl_0
  );


  and

  (
    g2008_p,
    g2007_n_spl_,
    g2006_n_spl_
  );


  or

  (
    g2008_n,
    g2007_p_spl_,
    g2006_p_spl_
  );


  and

  (
    g2009_p,
    g2008_n_spl_0,
    g2003_n_spl_
  );


  or

  (
    g2009_n,
    g2008_p_spl_0,
    g2003_p_spl_
  );


  and

  (
    g2010_p,
    g2009_n_spl_,
    g2002_n_spl_
  );


  or

  (
    g2010_n,
    g2009_p_spl_,
    g2002_p_spl_
  );


  and

  (
    g2011_p,
    g2010_n_spl_0,
    g2002_n_spl_
  );


  or

  (
    g2011_n,
    g2010_p_spl_0,
    g2002_p_spl_
  );


  and

  (
    g2012_p,
    g2010_n_spl_0,
    g2009_n_spl_
  );


  or

  (
    g2012_n,
    g2010_p_spl_0,
    g2009_p_spl_
  );


  and

  (
    g2013_p,
    g2012_n,
    g2011_n
  );


  or

  (
    g2013_n,
    g2012_p,
    g2011_p
  );


  and

  (
    g2014_p,
    n2608_lo_buf_o2_p_spl_00,
    n2734_lo_p_spl_100
  );


  or

  (
    g2014_n,
    n2608_lo_buf_o2_n_spl_0,
    n2734_lo_n_spl_100
  );


  and

  (
    g2015_p,
    g2014_n_spl_,
    g2013_n_spl_
  );


  or

  (
    g2015_n,
    g2014_p_spl_,
    g2013_p_spl_
  );


  and

  (
    g2016_p,
    g2015_n_spl_0,
    g2010_n_spl_
  );


  or

  (
    g2016_n,
    g2015_p_spl_0,
    g2010_p_spl_
  );


  and

  (
    g2017_p,
    g2016_n_spl_,
    g1999_n_spl_
  );


  or

  (
    g2017_n,
    g2016_p_spl_,
    g1999_p_spl_
  );


  and

  (
    g2018_p,
    g2017_n_spl_0,
    g1999_n_spl_
  );


  or

  (
    g2018_n,
    g2017_p_spl_0,
    g1999_p_spl_
  );


  and

  (
    g2019_p,
    g2017_n_spl_0,
    g2016_n_spl_
  );


  or

  (
    g2019_n,
    g2017_p_spl_0,
    g2016_p_spl_
  );


  and

  (
    g2020_p,
    g2019_n,
    g2018_n
  );


  or

  (
    g2020_n,
    g2019_p,
    g2018_p
  );


  and

  (
    g2021_p,
    n2608_lo_buf_o2_p_spl_0,
    n2746_lo_p_spl_010
  );


  or

  (
    g2021_n,
    n2608_lo_buf_o2_n_spl_1,
    n2746_lo_n_spl_011
  );


  and

  (
    g2022_p,
    g2021_n_spl_,
    g2020_n_spl_
  );


  or

  (
    g2022_n,
    g2021_p_spl_,
    g2020_p_spl_
  );


  and

  (
    g2023_p,
    g2022_n_spl_0,
    g2020_n_spl_
  );


  or

  (
    g2023_n,
    g2022_p_spl_0,
    g2020_p_spl_
  );


  and

  (
    g2024_p,
    g2022_n_spl_0,
    g2021_n_spl_
  );


  or

  (
    g2024_n,
    g2022_p_spl_0,
    g2021_p_spl_
  );


  and

  (
    g2025_p,
    g2024_n,
    g2023_n
  );


  or

  (
    g2025_n,
    g2024_p,
    g2023_p
  );


  and

  (
    g2026_p,
    g2015_n_spl_0,
    g2013_n_spl_
  );


  or

  (
    g2026_n,
    g2015_p_spl_0,
    g2013_p_spl_
  );


  and

  (
    g2027_p,
    g2015_n_spl_,
    g2014_n_spl_
  );


  or

  (
    g2027_n,
    g2015_p_spl_,
    g2014_p_spl_
  );


  and

  (
    g2028_p,
    g2027_n,
    g2026_n
  );


  or

  (
    g2028_n,
    g2027_p,
    g2026_p
  );


  and

  (
    g2029_p,
    g2008_n_spl_0,
    g2006_n_spl_
  );


  or

  (
    g2029_n,
    g2008_p_spl_0,
    g2006_p_spl_
  );


  and

  (
    g2030_p,
    g2008_n_spl_,
    g2007_n_spl_
  );


  or

  (
    g2030_n,
    g2008_p_spl_,
    g2007_p_spl_
  );


  and

  (
    g2031_p,
    g2030_n,
    g2029_n
  );


  or

  (
    g2031_n,
    g2030_p,
    g2029_p
  );


  and

  (
    g2032_p,
    G2196_o2_n,
    G2197_o2_p
  );


  or

  (
    g2032_n,
    G2196_o2_p,
    G2197_o2_n
  );


  and

  (
    g2033_p,
    G2118_o2_n_spl_0,
    G1980_o2_p
  );


  or

  (
    g2033_n,
    G2118_o2_p_spl_0,
    G1980_o2_n
  );


  and

  (
    g2034_p,
    g2033_n_spl_,
    g2032_n_spl_
  );


  or

  (
    g2034_n,
    g2033_p_spl_,
    g2032_p_spl_
  );


  and

  (
    g2035_p,
    g2034_n_spl_0,
    g2032_n_spl_
  );


  or

  (
    g2035_n,
    g2034_p_spl_0,
    g2032_p_spl_
  );


  and

  (
    g2036_p,
    g2034_n_spl_0,
    g2033_n_spl_
  );


  or

  (
    g2036_n,
    g2034_p_spl_0,
    g2033_p_spl_
  );


  and

  (
    g2037_p,
    g2036_n,
    g2035_n
  );


  or

  (
    g2037_n,
    g2036_p,
    g2035_p
  );


  and

  (
    g2038_p,
    n2728_lo_buf_o2_p_spl_110,
    n2596_lo_buf_o2_p_spl_00
  );


  or

  (
    g2038_n,
    n2728_lo_buf_o2_n_spl_110,
    n2596_lo_buf_o2_n_spl_0
  );


  and

  (
    g2039_p,
    g2038_n_spl_,
    g2037_n_spl_
  );


  or

  (
    g2039_n,
    g2038_p_spl_,
    g2037_p_spl_
  );


  and

  (
    g2040_p,
    g2039_n_spl_0,
    g2034_n_spl_
  );


  or

  (
    g2040_n,
    g2039_p_spl_0,
    g2034_p_spl_
  );


  and

  (
    g2041_p,
    g2040_n_spl_,
    g2031_n_spl_
  );


  or

  (
    g2041_n,
    g2040_p_spl_,
    g2031_p_spl_
  );


  and

  (
    g2042_p,
    g2041_n_spl_0,
    g2031_n_spl_
  );


  or

  (
    g2042_n,
    g2041_p_spl_0,
    g2031_p_spl_
  );


  and

  (
    g2043_p,
    g2041_n_spl_0,
    g2040_n_spl_
  );


  or

  (
    g2043_n,
    g2041_p_spl_0,
    g2040_p_spl_
  );


  and

  (
    g2044_p,
    g2043_n,
    g2042_n
  );


  or

  (
    g2044_n,
    g2043_p,
    g2042_p
  );


  and

  (
    g2045_p,
    n2596_lo_buf_o2_p_spl_00,
    n2734_lo_p_spl_100
  );


  or

  (
    g2045_n,
    n2596_lo_buf_o2_n_spl_0,
    n2734_lo_n_spl_100
  );


  and

  (
    g2046_p,
    g2045_n_spl_,
    g2044_n_spl_
  );


  or

  (
    g2046_n,
    g2045_p_spl_,
    g2044_p_spl_
  );


  and

  (
    g2047_p,
    g2046_n_spl_0,
    g2041_n_spl_
  );


  or

  (
    g2047_n,
    g2046_p_spl_0,
    g2041_p_spl_
  );


  and

  (
    g2048_p,
    g2047_n_spl_,
    g2028_n_spl_
  );


  or

  (
    g2048_n,
    g2047_p_spl_,
    g2028_p_spl_
  );


  and

  (
    g2049_p,
    g2048_n_spl_0,
    g2028_n_spl_
  );


  or

  (
    g2049_n,
    g2048_p_spl_0,
    g2028_p_spl_
  );


  and

  (
    g2050_p,
    g2048_n_spl_0,
    g2047_n_spl_
  );


  or

  (
    g2050_n,
    g2048_p_spl_0,
    g2047_p_spl_
  );


  and

  (
    g2051_p,
    g2050_n,
    g2049_n
  );


  or

  (
    g2051_n,
    g2050_p,
    g2049_p
  );


  and

  (
    g2052_p,
    n2596_lo_buf_o2_p_spl_0,
    n2746_lo_p_spl_011
  );


  or

  (
    g2052_n,
    n2596_lo_buf_o2_n_spl_1,
    n2746_lo_n_spl_011
  );


  and

  (
    g2053_p,
    g2052_n_spl_,
    g2051_n_spl_
  );


  or

  (
    g2053_n,
    g2052_p_spl_,
    g2051_p_spl_
  );


  and

  (
    g2054_p,
    g2053_n_spl_0,
    g2048_n_spl_
  );


  or

  (
    g2054_n,
    g2053_p_spl_0,
    g2048_p_spl_
  );


  and

  (
    g2055_p,
    g2054_n_spl_,
    g2025_n_spl_
  );


  or

  (
    g2055_n,
    g2054_p_spl_,
    g2025_p_spl_
  );


  and

  (
    g2056_p,
    g2055_n_spl_0,
    g2025_n_spl_
  );


  or

  (
    g2056_n,
    g2055_p_spl_0,
    g2025_p_spl_
  );


  and

  (
    g2057_p,
    g2055_n_spl_0,
    g2054_n_spl_
  );


  or

  (
    g2057_n,
    g2055_p_spl_0,
    g2054_p_spl_
  );


  and

  (
    g2058_p,
    g2057_n,
    g2056_n
  );


  or

  (
    g2058_n,
    g2057_p,
    g2056_p
  );


  and

  (
    g2059_p,
    n2596_lo_buf_o2_p_spl_1,
    n2758_lo_p_spl_000
  );


  or

  (
    g2059_n,
    n2596_lo_buf_o2_n_spl_1,
    n2758_lo_n_spl_000
  );


  and

  (
    g2060_p,
    g2059_n_spl_,
    g2058_n_spl_
  );


  or

  (
    g2060_n,
    g2059_p_spl_,
    g2058_p_spl_
  );


  and

  (
    g2061_p,
    g2060_n_spl_0,
    g2058_n_spl_
  );


  or

  (
    g2061_n,
    g2060_p_spl_0,
    g2058_p_spl_
  );


  and

  (
    g2062_p,
    g2060_n_spl_0,
    g2059_n_spl_
  );


  or

  (
    g2062_n,
    g2060_p_spl_0,
    g2059_p_spl_
  );


  and

  (
    g2063_p,
    g2062_n,
    g2061_n
  );


  or

  (
    g2063_n,
    g2062_p,
    g2061_p
  );


  and

  (
    g2064_p,
    g2053_n_spl_0,
    g2051_n_spl_
  );


  or

  (
    g2064_n,
    g2053_p_spl_0,
    g2051_p_spl_
  );


  and

  (
    g2065_p,
    g2053_n_spl_,
    g2052_n_spl_
  );


  or

  (
    g2065_n,
    g2053_p_spl_,
    g2052_p_spl_
  );


  and

  (
    g2066_p,
    g2065_n,
    g2064_n
  );


  or

  (
    g2066_n,
    g2065_p,
    g2064_p
  );


  and

  (
    g2067_p,
    g2046_n_spl_0,
    g2044_n_spl_
  );


  or

  (
    g2067_n,
    g2046_p_spl_0,
    g2044_p_spl_
  );


  and

  (
    g2068_p,
    g2046_n_spl_,
    g2045_n_spl_
  );


  or

  (
    g2068_n,
    g2046_p_spl_,
    g2045_p_spl_
  );


  and

  (
    g2069_p,
    g2068_n,
    g2067_n
  );


  or

  (
    g2069_n,
    g2068_p,
    g2067_p
  );


  and

  (
    g2070_p,
    g2039_n_spl_0,
    g2037_n_spl_
  );


  or

  (
    g2070_n,
    g2039_p_spl_0,
    g2037_p_spl_
  );


  and

  (
    g2071_p,
    g2039_n_spl_,
    g2038_n_spl_
  );


  or

  (
    g2071_n,
    g2039_p_spl_,
    g2038_p_spl_
  );


  and

  (
    g2072_p,
    g2071_n,
    g2070_n
  );


  or

  (
    g2072_n,
    g2071_p,
    g2070_p
  );


  and

  (
    g2073_p,
    G2118_o2_n_spl_0,
    G2061_o2_p
  );


  or

  (
    g2073_n,
    G2118_o2_p_spl_0,
    G2061_o2_n
  );


  and

  (
    g2074_p,
    G2118_o2_n_spl_,
    G983_o2_n
  );


  or

  (
    g2074_n,
    G2118_o2_p_spl_,
    G983_o2_p
  );


  and

  (
    g2075_p,
    g2074_n,
    g2073_n
  );


  or

  (
    g2075_n,
    g2074_p,
    g2073_p
  );


  and

  (
    g2076_p,
    G2058_o2_p_spl_,
    G935_o2_n_spl_
  );


  or

  (
    g2076_n,
    G2058_o2_n_spl_,
    G935_o2_p_spl_
  );


  and

  (
    g2077_p,
    g2076_n_spl_0,
    G1976_o2_p
  );


  or

  (
    g2077_n,
    g2076_p_spl_0,
    G1976_o2_n
  );


  and

  (
    g2078_p,
    g2077_n_spl_,
    g2075_n_spl_
  );


  or

  (
    g2078_n,
    g2077_p_spl_,
    g2075_p_spl_
  );


  and

  (
    g2079_p,
    g2078_n_spl_0,
    g2075_n_spl_
  );


  or

  (
    g2079_n,
    g2078_p_spl_0,
    g2075_p_spl_
  );


  and

  (
    g2080_p,
    g2078_n_spl_0,
    g2077_n_spl_
  );


  or

  (
    g2080_n,
    g2078_p_spl_0,
    g2077_p_spl_
  );


  and

  (
    g2081_p,
    g2080_n,
    g2079_n
  );


  or

  (
    g2081_n,
    g2080_p,
    g2079_p
  );


  and

  (
    g2082_p,
    n2728_lo_buf_o2_p_spl_110,
    n2584_lo_buf_o2_p_spl_00
  );


  or

  (
    g2082_n,
    n2728_lo_buf_o2_n_spl_110,
    n2584_lo_buf_o2_n_spl_00
  );


  and

  (
    g2083_p,
    g2082_n_spl_,
    g2081_n_spl_
  );


  or

  (
    g2083_n,
    g2082_p_spl_,
    g2081_p_spl_
  );


  and

  (
    g2084_p,
    g2083_n_spl_0,
    g2078_n_spl_
  );


  or

  (
    g2084_n,
    g2083_p_spl_0,
    g2078_p_spl_
  );


  and

  (
    g2085_p,
    g2084_n_spl_,
    g2072_n_spl_
  );


  or

  (
    g2085_n,
    g2084_p_spl_,
    g2072_p_spl_
  );


  and

  (
    g2086_p,
    g2085_n_spl_0,
    g2072_n_spl_
  );


  or

  (
    g2086_n,
    g2085_p_spl_0,
    g2072_p_spl_
  );


  and

  (
    g2087_p,
    g2085_n_spl_0,
    g2084_n_spl_
  );


  or

  (
    g2087_n,
    g2085_p_spl_0,
    g2084_p_spl_
  );


  and

  (
    g2088_p,
    g2087_n,
    g2086_n
  );


  or

  (
    g2088_n,
    g2087_p,
    g2086_p
  );


  and

  (
    g2089_p,
    n2584_lo_buf_o2_p_spl_00,
    n2734_lo_p_spl_101
  );


  or

  (
    g2089_n,
    n2584_lo_buf_o2_n_spl_00,
    n2734_lo_n_spl_101
  );


  and

  (
    g2090_p,
    g2089_n_spl_,
    g2088_n_spl_
  );


  or

  (
    g2090_n,
    g2089_p_spl_,
    g2088_p_spl_
  );


  and

  (
    g2091_p,
    g2090_n_spl_0,
    g2085_n_spl_
  );


  or

  (
    g2091_n,
    g2090_p_spl_0,
    g2085_p_spl_
  );


  and

  (
    g2092_p,
    g2091_n_spl_,
    g2069_n_spl_
  );


  or

  (
    g2092_n,
    g2091_p_spl_,
    g2069_p_spl_
  );


  and

  (
    g2093_p,
    g2092_n_spl_0,
    g2069_n_spl_
  );


  or

  (
    g2093_n,
    g2092_p_spl_0,
    g2069_p_spl_
  );


  and

  (
    g2094_p,
    g2092_n_spl_0,
    g2091_n_spl_
  );


  or

  (
    g2094_n,
    g2092_p_spl_0,
    g2091_p_spl_
  );


  and

  (
    g2095_p,
    g2094_n,
    g2093_n
  );


  or

  (
    g2095_n,
    g2094_p,
    g2093_p
  );


  and

  (
    g2096_p,
    n2584_lo_buf_o2_p_spl_0,
    n2746_lo_p_spl_011
  );


  or

  (
    g2096_n,
    n2584_lo_buf_o2_n_spl_0,
    n2746_lo_n_spl_100
  );


  and

  (
    g2097_p,
    g2096_n_spl_,
    g2095_n_spl_
  );


  or

  (
    g2097_n,
    g2096_p_spl_,
    g2095_p_spl_
  );


  and

  (
    g2098_p,
    g2097_n_spl_0,
    g2092_n_spl_
  );


  or

  (
    g2098_n,
    g2097_p_spl_0,
    g2092_p_spl_
  );


  and

  (
    g2099_p,
    g2098_n_spl_,
    g2066_n_spl_
  );


  or

  (
    g2099_n,
    g2098_p_spl_,
    g2066_p_spl_
  );


  and

  (
    g2100_p,
    g2099_n_spl_0,
    g2066_n_spl_
  );


  or

  (
    g2100_n,
    g2099_p_spl_0,
    g2066_p_spl_
  );


  and

  (
    g2101_p,
    g2099_n_spl_0,
    g2098_n_spl_
  );


  or

  (
    g2101_n,
    g2099_p_spl_0,
    g2098_p_spl_
  );


  and

  (
    g2102_p,
    g2101_n,
    g2100_n
  );


  or

  (
    g2102_n,
    g2101_p,
    g2100_p
  );


  and

  (
    g2103_p,
    n2584_lo_buf_o2_p_spl_1,
    n2758_lo_p_spl_000
  );


  or

  (
    g2103_n,
    n2584_lo_buf_o2_n_spl_1,
    n2758_lo_n_spl_000
  );


  and

  (
    g2104_p,
    g2103_n_spl_,
    g2102_n_spl_
  );


  or

  (
    g2104_n,
    g2103_p_spl_,
    g2102_p_spl_
  );


  and

  (
    g2105_p,
    g2104_n_spl_0,
    g2099_n_spl_
  );


  or

  (
    g2105_n,
    g2104_p_spl_0,
    g2099_p_spl_
  );


  or

  (
    g2106_n,
    g2105_p,
    g2063_p
  );


  and

  (
    g2107_p,
    g1973_n_spl_0,
    g1971_n_spl_
  );


  or

  (
    g2107_n,
    g1973_p_spl_0,
    g1971_p_spl_
  );


  and

  (
    g2108_p,
    g1973_n_spl_,
    g1972_n_spl_
  );


  or

  (
    g2108_n,
    g1973_p_spl_,
    g1972_p_spl_
  );


  and

  (
    g2109_p,
    g2108_n,
    g2107_n
  );


  or

  (
    g2109_n,
    g2108_p,
    g2107_p
  );


  and

  (
    g2110_p,
    g1488_n_spl_,
    g1483_n_spl_
  );


  or

  (
    g2110_n,
    g1488_p_spl_,
    g1483_p_spl_
  );


  and

  (
    g2111_p,
    g2110_n_spl_,
    g2109_n_spl_
  );


  or

  (
    g2111_n,
    g2110_p_spl_,
    g2109_p_spl_
  );


  and

  (
    g2112_p,
    g2111_n_spl_0,
    g2109_n_spl_
  );


  or

  (
    g2112_n,
    g2111_p_spl_0,
    g2109_p_spl_
  );


  and

  (
    g2113_p,
    g2111_n_spl_0,
    g2110_n_spl_
  );


  or

  (
    g2113_n,
    g2111_p_spl_0,
    g2110_p_spl_
  );


  and

  (
    g2114_p,
    g2113_n,
    g2112_n
  );


  or

  (
    g2114_n,
    g2113_p,
    g2112_p
  );


  and

  (
    g2115_p,
    n2728_lo_buf_o2_p_spl_111,
    n2512_lo_buf_o2_p_spl_01
  );


  or

  (
    g2115_n,
    n2728_lo_buf_o2_n_spl_111,
    n2512_lo_buf_o2_n_spl_0
  );


  and

  (
    g2116_p,
    g2115_n_spl_,
    g2114_n_spl_
  );


  or

  (
    g2116_n,
    g2115_p_spl_,
    g2114_p_spl_
  );


  and

  (
    g2117_p,
    g2116_n_spl_0,
    g2114_n_spl_
  );


  or

  (
    g2117_n,
    g2116_p_spl_0,
    g2114_p_spl_
  );


  and

  (
    g2118_p,
    g2116_n_spl_0,
    g2115_n_spl_
  );


  or

  (
    g2118_n,
    g2116_p_spl_0,
    g2115_p_spl_
  );


  and

  (
    g2119_p,
    g2118_n,
    g2117_n
  );


  or

  (
    g2119_n,
    g2118_p,
    g2117_p
  );


  and

  (
    g2120_p,
    g1498_n_spl_,
    g1493_n_spl_
  );


  or

  (
    g2120_n,
    g1498_p_spl_,
    g1493_p_spl_
  );


  and

  (
    g2121_p,
    g2120_n_spl_,
    g2119_n_spl_
  );


  or

  (
    g2121_n,
    g2120_p_spl_,
    g2119_p_spl_
  );


  and

  (
    g2122_p,
    g2121_n_spl_0,
    g2119_n_spl_
  );


  or

  (
    g2122_n,
    g2121_p_spl_0,
    g2119_p_spl_
  );


  and

  (
    g2123_p,
    g2121_n_spl_0,
    g2120_n_spl_
  );


  or

  (
    g2123_n,
    g2121_p_spl_0,
    g2120_p_spl_
  );


  and

  (
    g2124_p,
    g2123_n,
    g2122_n
  );


  or

  (
    g2124_n,
    g2123_p,
    g2122_p
  );


  and

  (
    g2125_p,
    n2500_lo_buf_o2_p_spl_01,
    n2734_lo_p_spl_101
  );


  or

  (
    g2125_n,
    n2500_lo_buf_o2_n_spl_1,
    n2734_lo_n_spl_101
  );


  and

  (
    g2126_p,
    g2125_n_spl_,
    g2124_n_spl_
  );


  or

  (
    g2126_n,
    g2125_p_spl_,
    g2124_p_spl_
  );


  and

  (
    g2127_p,
    g2126_n_spl_0,
    g2124_n_spl_
  );


  or

  (
    g2127_n,
    g2126_p_spl_0,
    g2124_p_spl_
  );


  and

  (
    g2128_p,
    g2126_n_spl_0,
    g2125_n_spl_
  );


  or

  (
    g2128_n,
    g2126_p_spl_0,
    g2125_p_spl_
  );


  and

  (
    g2129_p,
    g2128_n,
    g2127_n
  );


  or

  (
    g2129_n,
    g2128_p,
    g2127_p
  );


  and

  (
    g2130_p,
    g1508_n,
    g1503_n_spl_
  );


  or

  (
    g2130_n,
    g1508_p_spl_,
    g1503_p_spl_
  );


  and

  (
    g2131_p,
    g2130_n_spl_,
    g2129_n_spl_
  );


  or

  (
    g2131_n,
    g2130_p,
    g2129_p
  );


  and

  (
    g2132_p,
    g2131_n_spl_,
    g2129_n_spl_
  );


  and

  (
    g2133_p,
    g2131_n_spl_,
    g2130_n_spl_
  );


  or

  (
    g2134_n,
    g2133_p,
    g2132_p
  );


  or

  (
    g2135_n,
    n7280_o2_n_spl_1,
    n2797_lo_n_spl_11
  );


  or

  (
    g2136_n,
    n7459_o2_n_spl_1,
    n2809_lo_n_spl_11
  );


  or

  (
    g2137_n,
    n7675_o2_n_spl_1,
    n2821_lo_n_spl_0
  );


  or

  (
    g2138_n,
    n7835_o2_n_spl_1,
    n2821_lo_n_spl_1
  );


  and

  (
    g2139_p,
    g1558_n_spl_,
    g1553_n_spl_
  );


  and

  (
    g2140_p,
    g1573_n_spl_,
    g1568_n_spl_
  );


  and

  (
    g2141_p,
    g1588_n_spl_,
    g1583_n_spl_
  );


  and

  (
    g2142_p,
    g1563_n_spl_0,
    g1562_n
  );


  and

  (
    g2143_p,
    g1578_n_spl_0,
    g1577_n
  );


  and

  (
    g2144_p,
    g1593_n_spl_0,
    g1592_n
  );


  and

  (
    g2145_p,
    g1593_n_spl_0,
    g1591_n
  );


  and

  (
    g2146_p,
    g1578_n_spl_0,
    g1576_n
  );


  and

  (
    g2147_p,
    g1563_n_spl_0,
    g1561_n
  );


  and

  (
    g2148_p,
    g1602_n_spl_,
    g1545_n_spl_
  );


  and

  (
    g2149_p,
    g1599_n_spl_,
    g1546_n_spl_
  );


  and

  (
    g2150_p,
    g1596_n_spl_,
    g1547_n_spl_
  );


  and

  (
    g2151_p,
    g1605_n_spl_,
    g1548_n_spl_
  );


  and

  (
    g2152_p,
    g1220_n_spl_0,
    g1218_n
  );


  and

  (
    g2153_p,
    g1220_n_spl_0,
    g1219_n
  );


  or

  (
    g2154_n,
    g2153_p,
    g2152_p
  );


  and

  (
    g2155_p,
    g1225_n_spl_0,
    g1223_n
  );


  and

  (
    g2156_p,
    g1225_n_spl_0,
    g1224_n
  );


  or

  (
    g2157_n,
    g2156_p,
    g2155_p
  );


  and

  (
    g2158_p,
    g1230_n_spl_0,
    g1228_n
  );


  and

  (
    g2159_p,
    g1230_n_spl_0,
    g1229_n
  );


  or

  (
    g2160_n,
    g2159_p,
    g2158_p
  );


  and

  (
    g2161_p,
    n7148_o2_p_spl_1,
    n2785_lo_p_spl_111
  );


  or

  (
    g2161_n,
    n7148_o2_n_spl_,
    n2785_lo_n_spl_111
  );


  and

  (
    g2162_p,
    g1614_n_spl_,
    g1609_n_spl_
  );


  or

  (
    g2162_n,
    g1614_p_spl_,
    g1609_p_spl_
  );


  or

  (
    g2163_n,
    g2162_p,
    g2161_p
  );


  and

  (
    g2164_p,
    g1291_n_spl_0,
    g1289_n_spl_
  );


  or

  (
    g2164_n,
    g1291_p_spl_0,
    g1289_p_spl_
  );


  and

  (
    g2165_p,
    g1291_n_spl_,
    g1290_n_spl_
  );


  or

  (
    g2165_n,
    g1291_p_spl_,
    g1290_p_spl_
  );


  and

  (
    g2166_p,
    g2165_n,
    g2164_n
  );


  or

  (
    g2166_n,
    g2165_p,
    g2164_p
  );


  and

  (
    g2167_p,
    g1629_n_spl_,
    g1624_n_spl_
  );


  or

  (
    g2167_n,
    g1629_p_spl_,
    g1624_p_spl_
  );


  and

  (
    g2168_p,
    g2167_n_spl_,
    g2166_n_spl_
  );


  or

  (
    g2168_n,
    g2167_p_spl_,
    g2166_p_spl_
  );


  and

  (
    g2169_p,
    g2168_n_spl_0,
    g2166_n_spl_
  );


  or

  (
    g2169_n,
    g2168_p_spl_,
    g2166_p_spl_
  );


  and

  (
    g2170_p,
    g2168_n_spl_0,
    g2167_n_spl_
  );


  or

  (
    g2170_n,
    g2168_p_spl_,
    g2167_p_spl_
  );


  and

  (
    g2171_p,
    g2170_n,
    g2169_n
  );


  or

  (
    g2171_n,
    g2170_p,
    g2169_p
  );


  and

  (
    g2172_p,
    n7323_o2_p_spl_1,
    n2797_lo_p_spl_11
  );


  or

  (
    g2172_n,
    n7323_o2_n_spl_,
    n2797_lo_n_spl_11
  );


  and

  (
    g2173_p,
    g2172_n_spl_,
    g2171_n_spl_
  );


  or

  (
    g2173_n,
    g2172_p_spl_,
    g2171_p_spl_
  );


  and

  (
    g2174_p,
    g2173_n_spl_0,
    g2171_n_spl_
  );


  or

  (
    g2174_n,
    g2173_p_spl_,
    g2171_p_spl_
  );


  and

  (
    g2175_p,
    g2173_n_spl_0,
    g2172_n_spl_
  );


  or

  (
    g2175_n,
    g2173_p_spl_,
    g2172_p_spl_
  );


  and

  (
    g2176_p,
    g2175_n,
    g2174_n
  );


  or

  (
    g2176_n,
    g2175_p,
    g2174_p
  );


  and

  (
    g2177_p,
    g1639_n_spl_,
    g1634_n_spl_
  );


  or

  (
    g2177_n,
    g1639_p_spl_,
    g1634_p_spl_
  );


  or

  (
    g2178_n,
    g2177_p,
    g2176_p
  );


  and

  (
    g2179_p,
    g1365_n_spl_0,
    g1363_n_spl_
  );


  or

  (
    g2179_n,
    g1365_p_spl_0,
    g1363_p_spl_
  );


  and

  (
    g2180_p,
    g1365_n_spl_,
    g1364_n_spl_
  );


  or

  (
    g2180_n,
    g1365_p_spl_,
    g1364_p_spl_
  );


  and

  (
    g2181_p,
    g2180_n,
    g2179_n
  );


  or

  (
    g2181_n,
    g2180_p,
    g2179_p
  );


  and

  (
    g2182_p,
    g1654_n_spl_,
    g1649_n_spl_
  );


  or

  (
    g2182_n,
    g1654_p_spl_,
    g1649_p_spl_
  );


  and

  (
    g2183_p,
    g2182_n_spl_,
    g2181_n_spl_
  );


  or

  (
    g2183_n,
    g2182_p_spl_,
    g2181_p_spl_
  );


  and

  (
    g2184_p,
    g2183_n_spl_0,
    g2181_n_spl_
  );


  or

  (
    g2184_n,
    g2183_p_spl_,
    g2181_p_spl_
  );


  and

  (
    g2185_p,
    g2183_n_spl_0,
    g2182_n_spl_
  );


  or

  (
    g2185_n,
    g2183_p_spl_,
    g2182_p_spl_
  );


  and

  (
    g2186_p,
    g2185_n,
    g2184_n
  );


  or

  (
    g2186_n,
    g2185_p,
    g2184_p
  );


  and

  (
    g2187_p,
    n7518_o2_p_spl_1,
    n2809_lo_p_spl_11
  );


  or

  (
    g2187_n,
    n7518_o2_n_spl_,
    n2809_lo_n_spl_11
  );


  and

  (
    g2188_p,
    g2187_n_spl_,
    g2186_n_spl_
  );


  or

  (
    g2188_n,
    g2187_p_spl_,
    g2186_p_spl_
  );


  and

  (
    g2189_p,
    g2188_n_spl_0,
    g2186_n_spl_
  );


  or

  (
    g2189_n,
    g2188_p_spl_,
    g2186_p_spl_
  );


  and

  (
    g2190_p,
    g2188_n_spl_0,
    g2187_n_spl_
  );


  or

  (
    g2190_n,
    g2188_p_spl_,
    g2187_p_spl_
  );


  and

  (
    g2191_p,
    g2190_n,
    g2189_n
  );


  or

  (
    g2191_n,
    g2190_p,
    g2189_p
  );


  and

  (
    g2192_p,
    g1664_n_spl_,
    g1659_n_spl_
  );


  or

  (
    g2192_n,
    g1664_p_spl_,
    g1659_p_spl_
  );


  or

  (
    g2193_n,
    g2192_p,
    g2191_p
  );


  and

  (
    g2194_p,
    g1829_n_spl_0,
    g1827_n_spl_
  );


  or

  (
    g2194_n,
    g1829_p_spl_0,
    g1827_p_spl_
  );


  and

  (
    g2195_p,
    g1829_n_spl_,
    g1828_n_spl_
  );


  or

  (
    g2195_n,
    g1829_p_spl_,
    g1828_p_spl_
  );


  and

  (
    g2196_p,
    g2195_n,
    g2194_n
  );


  or

  (
    g2196_n,
    g2195_p,
    g2194_p
  );


  and

  (
    g2197_p,
    g1606_n,
    g1541_n_spl_
  );


  or

  (
    g2197_n,
    g1606_p_spl_,
    g1541_p_spl_
  );


  or

  (
    g2198_n,
    g2197_p,
    g2196_p
  );


  and

  (
    g2199_p,
    g1619_n_spl_0,
    g1617_n
  );


  and

  (
    g2200_p,
    g1619_n_spl_0,
    g1618_n
  );


  or

  (
    g2201_n,
    g2200_p,
    g2199_p
  );


  and

  (
    g2202_p,
    g1644_n_spl_0,
    g1642_n
  );


  and

  (
    g2203_p,
    g1644_n_spl_0,
    g1643_n
  );


  or

  (
    g2204_n,
    g2203_p,
    g2202_p
  );


  and

  (
    g2205_p,
    g1669_n_spl_0,
    g1667_n
  );


  and

  (
    g2206_p,
    g1669_n_spl_0,
    g1668_n
  );


  or

  (
    g2207_n,
    g2206_p,
    g2205_p
  );


  and

  (
    g2208_p,
    g1724_n_spl_0,
    g1702_n
  );


  and

  (
    g2209_p,
    g1724_n_spl_0,
    g1723_n
  );


  or

  (
    g2210_n,
    g2209_p,
    g2208_p
  );


  and

  (
    g2211_p,
    g1801_n_spl_0,
    g1774_n_spl_
  );


  or

  (
    g2211_n,
    g1801_p_spl_,
    g1774_p_spl_
  );


  and

  (
    g2212_p,
    g1801_n_spl_0,
    g1800_n_spl_
  );


  or

  (
    g2212_n,
    g1801_p_spl_,
    g1800_p_spl_
  );


  and

  (
    g2213_p,
    g2212_n,
    g2211_n
  );


  or

  (
    g2213_n,
    g2212_p,
    g2211_p
  );


  and

  (
    g2214_p,
    n2620_lo_buf_o2_p_spl_1,
    n2758_lo_p_spl_001
  );


  or

  (
    g2214_n,
    n2620_lo_buf_o2_n_spl_1,
    n2758_lo_n_spl_001
  );


  or

  (
    g2215_n,
    g2214_p,
    g2213_p
  );


  and

  (
    g2216_p,
    g2134_n_spl_,
    g1832_n_spl_
  );


  and

  (
    g2217_p,
    g1994_n_spl_0,
    g1992_n_spl_
  );


  or

  (
    g2217_n,
    g1994_p_spl_0,
    g1992_p_spl_
  );


  and

  (
    g2218_p,
    g1994_n_spl_,
    g1993_n_spl_
  );


  or

  (
    g2218_n,
    g1994_p_spl_,
    g1993_p_spl_
  );


  and

  (
    g2219_p,
    g2218_n,
    g2217_n
  );


  or

  (
    g2219_n,
    g2218_p,
    g2217_p
  );


  and

  (
    g2220_p,
    g1987_n_spl_0,
    g1985_n_spl_
  );


  or

  (
    g2220_n,
    g1987_p_spl_0,
    g1985_p_spl_
  );


  and

  (
    g2221_p,
    g1987_n_spl_,
    g1986_n_spl_
  );


  or

  (
    g2221_n,
    g1987_p_spl_,
    g1986_p_spl_
  );


  and

  (
    g2222_p,
    g2221_n,
    g2220_n
  );


  or

  (
    g2222_n,
    g2221_p,
    g2220_p
  );


  and

  (
    g2223_p,
    g1980_n_spl_0,
    g1978_n_spl_
  );


  or

  (
    g2223_n,
    g1980_p_spl_0,
    g1978_p_spl_
  );


  and

  (
    g2224_p,
    g1980_n_spl_,
    g1979_n_spl_
  );


  or

  (
    g2224_n,
    g1980_p_spl_,
    g1979_p_spl_
  );


  and

  (
    g2225_p,
    g2224_n,
    g2223_n
  );


  or

  (
    g2225_n,
    g2224_p,
    g2223_p
  );


  and

  (
    g2226_p,
    g2116_n_spl_,
    g2111_n_spl_
  );


  or

  (
    g2226_n,
    g2116_p_spl_,
    g2111_p_spl_
  );


  and

  (
    g2227_p,
    g2226_n_spl_,
    g2225_n_spl_
  );


  or

  (
    g2227_n,
    g2226_p_spl_,
    g2225_p_spl_
  );


  and

  (
    g2228_p,
    g2227_n_spl_0,
    g2225_n_spl_
  );


  or

  (
    g2228_n,
    g2227_p_spl_0,
    g2225_p_spl_
  );


  and

  (
    g2229_p,
    g2227_n_spl_0,
    g2226_n_spl_
  );


  or

  (
    g2229_n,
    g2227_p_spl_0,
    g2226_p_spl_
  );


  and

  (
    g2230_p,
    g2229_n,
    g2228_n
  );


  or

  (
    g2230_n,
    g2229_p,
    g2228_p
  );


  and

  (
    g2231_p,
    n2512_lo_buf_o2_p_spl_01,
    n2734_lo_p_spl_110
  );


  or

  (
    g2231_n,
    n2512_lo_buf_o2_n_spl_1,
    n2734_lo_n_spl_110
  );


  and

  (
    g2232_p,
    g2231_n_spl_,
    g2230_n_spl_
  );


  or

  (
    g2232_n,
    g2231_p_spl_,
    g2230_p_spl_
  );


  and

  (
    g2233_p,
    g2232_n_spl_0,
    g2227_n_spl_
  );


  or

  (
    g2233_n,
    g2232_p_spl_0,
    g2227_p_spl_
  );


  and

  (
    g2234_p,
    g2233_n_spl_,
    g2222_n_spl_
  );


  or

  (
    g2234_n,
    g2233_p_spl_,
    g2222_p_spl_
  );


  and

  (
    g2235_p,
    g2234_n_spl_0,
    g2222_n_spl_
  );


  or

  (
    g2235_n,
    g2234_p_spl_0,
    g2222_p_spl_
  );


  and

  (
    g2236_p,
    g2234_n_spl_0,
    g2233_n_spl_
  );


  or

  (
    g2236_n,
    g2234_p_spl_0,
    g2233_p_spl_
  );


  and

  (
    g2237_p,
    g2236_n,
    g2235_n
  );


  or

  (
    g2237_n,
    g2236_p,
    g2235_p
  );


  and

  (
    g2238_p,
    n2512_lo_buf_o2_p_spl_10,
    n2746_lo_p_spl_100
  );


  or

  (
    g2238_n,
    n2512_lo_buf_o2_n_spl_1,
    n2746_lo_n_spl_100
  );


  and

  (
    g2239_p,
    g2238_n_spl_,
    g2237_n_spl_
  );


  or

  (
    g2239_n,
    g2238_p_spl_,
    g2237_p_spl_
  );


  and

  (
    g2240_p,
    g2239_n_spl_0,
    g2234_n_spl_
  );


  or

  (
    g2240_n,
    g2239_p_spl_0,
    g2234_p_spl_
  );


  or

  (
    g2241_n,
    g2240_p,
    g2219_p
  );


  and

  (
    g2242_p,
    g2104_n_spl_0,
    g2102_n_spl_
  );


  or

  (
    g2242_n,
    g2104_p_spl_0,
    g2102_p_spl_
  );


  and

  (
    g2243_p,
    g2104_n_spl_,
    g2103_n_spl_
  );


  or

  (
    g2243_n,
    g2104_p_spl_,
    g2103_p_spl_
  );


  and

  (
    g2244_p,
    g2243_n,
    g2242_n
  );


  or

  (
    g2244_n,
    g2243_p,
    g2242_p
  );


  and

  (
    g2245_p,
    g2097_n_spl_0,
    g2095_n_spl_
  );


  or

  (
    g2245_n,
    g2097_p_spl_0,
    g2095_p_spl_
  );


  and

  (
    g2246_p,
    g2097_n_spl_,
    g2096_n_spl_
  );


  or

  (
    g2246_n,
    g2097_p_spl_,
    g2096_p_spl_
  );


  and

  (
    g2247_p,
    g2246_n,
    g2245_n
  );


  or

  (
    g2247_n,
    g2246_p,
    g2245_p
  );


  and

  (
    g2248_p,
    g2090_n_spl_0,
    g2088_n_spl_
  );


  or

  (
    g2248_n,
    g2090_p_spl_0,
    g2088_p_spl_
  );


  and

  (
    g2249_p,
    g2090_n_spl_,
    g2089_n_spl_
  );


  or

  (
    g2249_n,
    g2090_p_spl_,
    g2089_p_spl_
  );


  and

  (
    g2250_p,
    g2249_n,
    g2248_n
  );


  or

  (
    g2250_n,
    g2249_p,
    g2248_p
  );


  and

  (
    g2251_p,
    g2083_n_spl_0,
    g2081_n_spl_
  );


  or

  (
    g2251_n,
    g2083_p_spl_0,
    g2081_p_spl_
  );


  and

  (
    g2252_p,
    g2083_n_spl_,
    g2082_n_spl_
  );


  or

  (
    g2252_n,
    g2083_p_spl_,
    g2082_p_spl_
  );


  and

  (
    g2253_p,
    g2252_n,
    g2251_n
  );


  or

  (
    g2253_n,
    g2252_p,
    g2251_p
  );


  and

  (
    g2254_p,
    g2076_n_spl_0,
    G2058_o2_p_spl_
  );


  or

  (
    g2254_n,
    g2076_p_spl_0,
    G2058_o2_n_spl_
  );


  and

  (
    g2255_p,
    g2076_n_spl_,
    G935_o2_n_spl_
  );


  or

  (
    g2255_n,
    g2076_p_spl_,
    G935_o2_p_spl_
  );


  and

  (
    g2256_p,
    g2255_n,
    g2254_n
  );


  or

  (
    g2256_n,
    g2255_p,
    g2254_p
  );


  and

  (
    g2257_p,
    g1872_n_spl_,
    G1972_o2_p
  );


  or

  (
    g2257_n,
    g1872_p_spl_,
    G1972_o2_n
  );


  and

  (
    g2258_p,
    g2257_n_spl_,
    g2256_n_spl_
  );


  or

  (
    g2258_n,
    g2257_p_spl_,
    g2256_p_spl_
  );


  and

  (
    g2259_p,
    g2258_n_spl_0,
    g2256_n_spl_
  );


  or

  (
    g2259_n,
    g2258_p_spl_0,
    g2256_p_spl_
  );


  and

  (
    g2260_p,
    g2258_n_spl_0,
    g2257_n_spl_
  );


  or

  (
    g2260_n,
    g2258_p_spl_0,
    g2257_p_spl_
  );


  and

  (
    g2261_p,
    g2260_n,
    g2259_n
  );


  or

  (
    g2261_n,
    g2260_p,
    g2259_p
  );


  and

  (
    g2262_p,
    n2728_lo_buf_o2_p_spl_111,
    n2572_lo_buf_o2_p_spl_00
  );


  or

  (
    g2262_n,
    n2728_lo_buf_o2_n_spl_111,
    n2572_lo_buf_o2_n_spl_00
  );


  and

  (
    g2263_p,
    g2262_n_spl_,
    g2261_n_spl_
  );


  or

  (
    g2263_n,
    g2262_p_spl_,
    g2261_p_spl_
  );


  and

  (
    g2264_p,
    g2263_n_spl_0,
    g2258_n_spl_
  );


  or

  (
    g2264_n,
    g2263_p_spl_0,
    g2258_p_spl_
  );


  and

  (
    g2265_p,
    g2264_n_spl_,
    g2253_n_spl_
  );


  or

  (
    g2265_n,
    g2264_p_spl_,
    g2253_p_spl_
  );


  and

  (
    g2266_p,
    g2265_n_spl_0,
    g2253_n_spl_
  );


  or

  (
    g2266_n,
    g2265_p_spl_0,
    g2253_p_spl_
  );


  and

  (
    g2267_p,
    g2265_n_spl_0,
    g2264_n_spl_
  );


  or

  (
    g2267_n,
    g2265_p_spl_0,
    g2264_p_spl_
  );


  and

  (
    g2268_p,
    g2267_n,
    g2266_n
  );


  or

  (
    g2268_n,
    g2267_p,
    g2266_p
  );


  and

  (
    g2269_p,
    n2572_lo_buf_o2_p_spl_01,
    n2734_lo_p_spl_110
  );


  or

  (
    g2269_n,
    n2572_lo_buf_o2_n_spl_0,
    n2734_lo_n_spl_110
  );


  and

  (
    g2270_p,
    g2269_n_spl_,
    g2268_n_spl_
  );


  or

  (
    g2270_n,
    g2269_p_spl_,
    g2268_p_spl_
  );


  and

  (
    g2271_p,
    g2270_n_spl_0,
    g2265_n_spl_
  );


  or

  (
    g2271_n,
    g2270_p_spl_0,
    g2265_p_spl_
  );


  and

  (
    g2272_p,
    g2271_n_spl_,
    g2250_n_spl_
  );


  or

  (
    g2272_n,
    g2271_p_spl_,
    g2250_p_spl_
  );


  and

  (
    g2273_p,
    g2272_n_spl_0,
    g2250_n_spl_
  );


  or

  (
    g2273_n,
    g2272_p_spl_0,
    g2250_p_spl_
  );


  and

  (
    g2274_p,
    g2272_n_spl_0,
    g2271_n_spl_
  );


  or

  (
    g2274_n,
    g2272_p_spl_0,
    g2271_p_spl_
  );


  and

  (
    g2275_p,
    g2274_n,
    g2273_n
  );


  or

  (
    g2275_n,
    g2274_p,
    g2273_p
  );


  and

  (
    g2276_p,
    n2572_lo_buf_o2_p_spl_01,
    n2746_lo_p_spl_100
  );


  or

  (
    g2276_n,
    n2572_lo_buf_o2_n_spl_1,
    n2746_lo_n_spl_101
  );


  and

  (
    g2277_p,
    g2276_n_spl_,
    g2275_n_spl_
  );


  or

  (
    g2277_n,
    g2276_p_spl_,
    g2275_p_spl_
  );


  and

  (
    g2278_p,
    g2277_n_spl_0,
    g2272_n_spl_
  );


  or

  (
    g2278_n,
    g2277_p_spl_0,
    g2272_p_spl_
  );


  and

  (
    g2279_p,
    g2278_n_spl_,
    g2247_n_spl_
  );


  or

  (
    g2279_n,
    g2278_p_spl_,
    g2247_p_spl_
  );


  and

  (
    g2280_p,
    g2279_n_spl_0,
    g2247_n_spl_
  );


  or

  (
    g2280_n,
    g2279_p_spl_0,
    g2247_p_spl_
  );


  and

  (
    g2281_p,
    g2279_n_spl_0,
    g2278_n_spl_
  );


  or

  (
    g2281_n,
    g2279_p_spl_0,
    g2278_p_spl_
  );


  and

  (
    g2282_p,
    g2281_n,
    g2280_n
  );


  or

  (
    g2282_n,
    g2281_p,
    g2280_p
  );


  and

  (
    g2283_p,
    n2572_lo_buf_o2_p_spl_10,
    n2758_lo_p_spl_001
  );


  or

  (
    g2283_n,
    n2572_lo_buf_o2_n_spl_1,
    n2758_lo_n_spl_001
  );


  and

  (
    g2284_p,
    g2283_n_spl_,
    g2282_n_spl_
  );


  or

  (
    g2284_n,
    g2283_p_spl_,
    g2282_p_spl_
  );


  and

  (
    g2285_p,
    g2284_n_spl_0,
    g2279_n_spl_
  );


  or

  (
    g2285_n,
    g2284_p_spl_0,
    g2279_p_spl_
  );


  or

  (
    g2286_n,
    g2285_p,
    g2244_p
  );


  and

  (
    g2287_p,
    G17_p_spl_000,
    G7_p_spl_0
  );


  or

  (
    g2287_n,
    G17_n_spl_000,
    G7_n_spl_0
  );


  and

  (
    g2288_p,
    G18_p_spl_001,
    G6_p_spl_0
  );


  or

  (
    g2288_n,
    G18_n_spl_001,
    G6_n_spl_0
  );


  and

  (
    g2289_p,
    g2288_n_spl_,
    g2287_p_spl_
  );


  or

  (
    g2289_n,
    g2288_p_spl_,
    g2287_n_spl_
  );


  and

  (
    g2290_p,
    g2289_n_spl_,
    g2287_p_spl_
  );


  or

  (
    g2290_n,
    g2289_p_spl_,
    g2287_n_spl_
  );


  and

  (
    g2291_p,
    g2289_n_spl_,
    g2288_n_spl_
  );


  or

  (
    g2291_n,
    g2289_p_spl_,
    g2288_p_spl_
  );


  and

  (
    g2292_p,
    g2291_n,
    g2290_n_spl_0
  );


  or

  (
    g2292_n,
    g2291_p,
    g2290_p_spl_0
  );


  and

  (
    g2293_p,
    G17_p_spl_001,
    G6_p_spl_0
  );


  or

  (
    g2293_n,
    G17_n_spl_001,
    G6_n_spl_0
  );


  and

  (
    g2294_p,
    G18_p_spl_001,
    G5_p_spl_0
  );


  or

  (
    g2294_n,
    G18_n_spl_001,
    G5_n_spl_0
  );


  and

  (
    g2295_p,
    g2294_n_spl_,
    g2293_p_spl_
  );


  or

  (
    g2295_n,
    g2294_p_spl_,
    g2293_n_spl_
  );


  and

  (
    g2296_p,
    g2295_n_spl_,
    g2293_p_spl_
  );


  or

  (
    g2296_n,
    g2295_p_spl_,
    g2293_n_spl_
  );


  or

  (
    g2297_n,
    g2296_p_spl_,
    g2292_p
  );


  and

  (
    g2298_p,
    G17_p_spl_001,
    G13_p_spl_00
  );


  or

  (
    g2298_n,
    G17_n_spl_001,
    G13_n_spl_0
  );


  and

  (
    g2299_p,
    G18_p_spl_010,
    G12_p_spl_00
  );


  or

  (
    g2299_n,
    G18_n_spl_010,
    G12_n_spl_0
  );


  and

  (
    g2300_p,
    g2299_n_spl_,
    g2298_p_spl_
  );


  or

  (
    g2300_n,
    g2299_p_spl_,
    g2298_n_spl_
  );


  and

  (
    g2301_p,
    g2300_n_spl_,
    g2298_p_spl_
  );


  or

  (
    g2301_n,
    g2300_p_spl_,
    g2298_n_spl_
  );


  and

  (
    g2302_p,
    g2300_n_spl_,
    g2299_n_spl_
  );


  or

  (
    g2302_n,
    g2300_p_spl_,
    g2299_p_spl_
  );


  and

  (
    g2303_p,
    g2302_n,
    g2301_n_spl_0
  );


  or

  (
    g2303_n,
    g2302_p,
    g2301_p_spl_0
  );


  and

  (
    g2304_p,
    G17_p_spl_010,
    G12_p_spl_00
  );


  or

  (
    g2304_n,
    G17_n_spl_010,
    G12_n_spl_0
  );


  and

  (
    g2305_p,
    G18_p_spl_010,
    G11_p_spl_00
  );


  or

  (
    g2305_n,
    G18_n_spl_010,
    G11_n_spl_0
  );


  and

  (
    g2306_p,
    g2305_n_spl_,
    g2304_p_spl_
  );


  or

  (
    g2306_n,
    g2305_p_spl_,
    g2304_n_spl_
  );


  and

  (
    g2307_p,
    g2306_n_spl_,
    g2304_p_spl_
  );


  or

  (
    g2307_n,
    g2306_p_spl_,
    g2304_n_spl_
  );


  and

  (
    g2308_p,
    g2307_n_spl_0,
    g2303_n_spl_
  );


  or

  (
    g2308_n,
    g2307_p_spl_0,
    g2303_p_spl_
  );


  and

  (
    g2309_p,
    g2308_n_spl_0,
    g2303_n_spl_
  );


  or

  (
    g2309_n,
    g2308_p_spl_0,
    g2303_p_spl_
  );


  and

  (
    g2310_p,
    g2308_n_spl_0,
    g2307_n_spl_0
  );


  or

  (
    g2310_n,
    g2308_p_spl_0,
    g2307_p_spl_0
  );


  and

  (
    g2311_p,
    g2310_n,
    g2309_n
  );


  or

  (
    g2311_n,
    g2310_p,
    g2309_p
  );


  and

  (
    g2312_p,
    G19_p_spl_001,
    G11_p_spl_00
  );


  or

  (
    g2312_n,
    G19_n_spl_001,
    G11_n_spl_0
  );


  and

  (
    g2313_p,
    g2312_n_spl_,
    g2311_n_spl_
  );


  or

  (
    g2313_n,
    g2312_p_spl_,
    g2311_p_spl_
  );


  and

  (
    g2314_p,
    g2313_n_spl_0,
    g2311_n_spl_
  );


  or

  (
    g2314_n,
    g2313_p_spl_0,
    g2311_p_spl_
  );


  and

  (
    g2315_p,
    g2313_n_spl_0,
    g2312_n_spl_
  );


  or

  (
    g2315_n,
    g2313_p_spl_0,
    g2312_p_spl_
  );


  and

  (
    g2316_p,
    g2315_n,
    g2314_n
  );


  or

  (
    g2316_n,
    g2315_p,
    g2314_p
  );


  and

  (
    g2317_p,
    g2306_n_spl_,
    g2305_n_spl_
  );


  or

  (
    g2317_n,
    g2306_p_spl_,
    g2305_p_spl_
  );


  and

  (
    g2318_p,
    g2317_n,
    g2307_n_spl_
  );


  or

  (
    g2318_n,
    g2317_p,
    g2307_p_spl_
  );


  and

  (
    g2319_p,
    G17_p_spl_010,
    G11_p_spl_0
  );


  or

  (
    g2319_n,
    G17_n_spl_010,
    G11_n_spl_1
  );


  and

  (
    g2320_p,
    G18_p_spl_011,
    G10_p_spl_0
  );


  or

  (
    g2320_n,
    G18_n_spl_011,
    G10_n_spl_0
  );


  and

  (
    g2321_p,
    g2320_n_spl_,
    g2319_p_spl_
  );


  or

  (
    g2321_n,
    g2320_p_spl_,
    g2319_n_spl_
  );


  and

  (
    g2322_p,
    g2321_n_spl_,
    g2319_p_spl_
  );


  or

  (
    g2322_n,
    g2321_p_spl_,
    g2319_n_spl_
  );


  and

  (
    g2323_p,
    g2322_n_spl_0,
    g2318_n_spl_
  );


  or

  (
    g2323_n,
    g2322_p_spl_0,
    g2318_p_spl_
  );


  and

  (
    g2324_p,
    g2323_n_spl_0,
    g2318_n_spl_
  );


  or

  (
    g2324_n,
    g2323_p_spl_0,
    g2318_p_spl_
  );


  and

  (
    g2325_p,
    g2323_n_spl_0,
    g2322_n_spl_0
  );


  or

  (
    g2325_n,
    g2323_p_spl_0,
    g2322_p_spl_0
  );


  and

  (
    g2326_p,
    g2325_n,
    g2324_n
  );


  or

  (
    g2326_n,
    g2325_p,
    g2324_p
  );


  and

  (
    g2327_p,
    G19_p_spl_001,
    G10_p_spl_0
  );


  or

  (
    g2327_n,
    G19_n_spl_001,
    G10_n_spl_0
  );


  and

  (
    g2328_p,
    g2327_n_spl_,
    g2326_n_spl_
  );


  or

  (
    g2328_n,
    g2327_p_spl_,
    g2326_p_spl_
  );


  and

  (
    g2329_p,
    g2328_n_spl_0,
    g2323_n_spl_
  );


  or

  (
    g2329_n,
    g2328_p_spl_0,
    g2323_p_spl_
  );


  or

  (
    g2330_n,
    g2329_p,
    g2316_p
  );


  and

  (
    g2331_p,
    n7909_o2_p_spl_10,
    n2821_lo_p_spl_0
  );


  or

  (
    g2332_n,
    n2632_lo_buf_o2_n_spl_1,
    n2758_lo_n_spl_01
  );


  or

  (
    g2333_n,
    n2584_lo_buf_o2_n_spl_1,
    n2770_lo_n
  );


  or

  (
    g2334_n,
    n2524_lo_buf_o2_n_spl_1,
    n2758_lo_n_spl_01
  );


  or

  (
    g2335_n,
    G18_n_spl_011,
    G1_n
  );


  and

  (
    g2336_p,
    g2173_n_spl_,
    g2168_n_spl_
  );


  and

  (
    g2337_p,
    g2188_n_spl_,
    g2183_n_spl_
  );


  and

  (
    g2338_p,
    g1475_n_spl_0,
    g1473_n_spl_
  );


  or

  (
    g2338_n,
    g1475_p_spl_0,
    g1473_p_spl_
  );


  and

  (
    g2339_p,
    g1475_n_spl_,
    g1474_n_spl_
  );


  or

  (
    g2339_n,
    g1475_p_spl_,
    g1474_p_spl_
  );


  and

  (
    g2340_p,
    g2339_n,
    g2338_n
  );


  or

  (
    g2340_n,
    g2339_p,
    g2338_p
  );


  and

  (
    g2341_p,
    g1699_n_spl_,
    g1694_n_spl_
  );


  or

  (
    g2341_n,
    g1699_p_spl_,
    g1694_p_spl_
  );


  and

  (
    g2342_p,
    g2341_n_spl_,
    g2340_n_spl_
  );


  or

  (
    g2342_n,
    g2341_p_spl_,
    g2340_p_spl_
  );


  and

  (
    g2343_p,
    g2342_n_spl_0,
    g2340_n_spl_
  );


  or

  (
    g2343_n,
    g2342_p_spl_,
    g2340_p_spl_
  );


  and

  (
    g2344_p,
    g2342_n_spl_0,
    g2341_n_spl_
  );


  or

  (
    g2344_n,
    g2342_p_spl_,
    g2341_p_spl_
  );


  and

  (
    g2345_p,
    g2344_n,
    g2343_n
  );


  or

  (
    g2345_n,
    g2344_p,
    g2343_p
  );


  and

  (
    g2346_p,
    n7747_o2_p_spl_1,
    n2821_lo_p_spl_1
  );


  or

  (
    g2346_n,
    n7747_o2_n_spl_1,
    n2821_lo_n_spl_1
  );


  or

  (
    g2347_n,
    g2346_p,
    g2345_p
  );


  and

  (
    g2348_p,
    g2347_n_spl_0,
    g2342_n_spl_
  );


  or

  (
    g2349_n,
    g2216_p_spl_,
    g2131_p
  );


  and

  (
    g2350_p,
    g2270_n_spl_0,
    g2268_n_spl_
  );


  or

  (
    g2350_n,
    g2270_p_spl_0,
    g2268_p_spl_
  );


  and

  (
    g2351_p,
    g2270_n_spl_,
    g2269_n_spl_
  );


  or

  (
    g2351_n,
    g2270_p_spl_,
    g2269_p_spl_
  );


  and

  (
    g2352_p,
    g2351_n,
    g2350_n
  );


  or

  (
    g2352_n,
    g2351_p,
    g2350_p
  );


  and

  (
    g2353_p,
    g2263_n_spl_0,
    g2261_n_spl_
  );


  or

  (
    g2353_n,
    g2263_p_spl_0,
    g2261_p_spl_
  );


  and

  (
    g2354_p,
    g2263_n_spl_,
    g2262_n_spl_
  );


  or

  (
    g2354_n,
    g2263_p_spl_,
    g2262_p_spl_
  );


  and

  (
    g2355_p,
    g2354_n,
    g2353_n
  );


  or

  (
    g2355_n,
    g2354_p,
    g2353_p
  );


  and

  (
    g2356_p,
    g1887_n_spl_,
    g1882_n_spl_
  );


  or

  (
    g2356_n,
    g1887_p_spl_,
    g1882_p_spl_
  );


  and

  (
    g2357_p,
    g2356_n_spl_,
    g2355_n_spl_
  );


  or

  (
    g2357_n,
    g2356_p_spl_,
    g2355_p_spl_
  );


  and

  (
    g2358_p,
    g2357_n_spl_0,
    g2355_n_spl_
  );


  or

  (
    g2358_n,
    g2357_p_spl_0,
    g2355_p_spl_
  );


  and

  (
    g2359_p,
    g2357_n_spl_0,
    g2356_n_spl_
  );


  or

  (
    g2359_n,
    g2357_p_spl_0,
    g2356_p_spl_
  );


  and

  (
    g2360_p,
    g2359_n,
    g2358_n
  );


  or

  (
    g2360_n,
    g2359_p,
    g2358_p
  );


  and

  (
    g2361_p,
    n2560_lo_buf_o2_p_spl_01,
    n2734_lo_p_spl_111
  );


  or

  (
    g2361_n,
    n2560_lo_buf_o2_n_spl_0,
    n2734_lo_n_spl_111
  );


  and

  (
    g2362_p,
    g2361_n_spl_,
    g2360_n_spl_
  );


  or

  (
    g2362_n,
    g2361_p_spl_,
    g2360_p_spl_
  );


  and

  (
    g2363_p,
    g2362_n_spl_0,
    g2357_n_spl_
  );


  or

  (
    g2363_n,
    g2362_p_spl_0,
    g2357_p_spl_
  );


  and

  (
    g2364_p,
    g2363_n_spl_,
    g2352_n_spl_
  );


  or

  (
    g2364_n,
    g2363_p_spl_,
    g2352_p_spl_
  );


  and

  (
    g2365_p,
    g2364_n_spl_0,
    g2352_n_spl_
  );


  or

  (
    g2365_n,
    g2364_p_spl_0,
    g2352_p_spl_
  );


  and

  (
    g2366_p,
    g2364_n_spl_0,
    g2363_n_spl_
  );


  or

  (
    g2366_n,
    g2364_p_spl_0,
    g2363_p_spl_
  );


  and

  (
    g2367_p,
    g2366_n,
    g2365_n
  );


  or

  (
    g2367_n,
    g2366_p,
    g2365_p
  );


  and

  (
    g2368_p,
    n2560_lo_buf_o2_p_spl_01,
    n2746_lo_p_spl_101
  );


  or

  (
    g2368_n,
    n2560_lo_buf_o2_n_spl_1,
    n2746_lo_n_spl_101
  );


  and

  (
    g2369_p,
    g2368_n_spl_,
    g2367_n_spl_
  );


  or

  (
    g2369_n,
    g2368_p_spl_,
    g2367_p_spl_
  );


  and

  (
    g2370_p,
    g2369_n_spl_0,
    g2367_n_spl_
  );


  or

  (
    g2370_n,
    g2369_p_spl_0,
    g2367_p_spl_
  );


  and

  (
    g2371_p,
    g2369_n_spl_0,
    g2368_n_spl_
  );


  or

  (
    g2371_n,
    g2369_p_spl_0,
    g2368_p_spl_
  );


  and

  (
    g2372_p,
    g2371_n,
    g2370_n
  );


  or

  (
    g2372_n,
    g2371_p,
    g2370_p
  );


  and

  (
    g2373_p,
    g2362_n_spl_0,
    g2360_n_spl_
  );


  or

  (
    g2373_n,
    g2362_p_spl_0,
    g2360_p_spl_
  );


  and

  (
    g2374_p,
    g2362_n_spl_,
    g2361_n_spl_
  );


  or

  (
    g2374_n,
    g2362_p_spl_,
    g2361_p_spl_
  );


  and

  (
    g2375_p,
    g2374_n,
    g2373_n
  );


  or

  (
    g2375_n,
    g2374_p,
    g2373_p
  );


  and

  (
    g2376_p,
    g1913_n_spl_,
    g1908_n_spl_
  );


  or

  (
    g2376_n,
    g1913_p_spl_,
    g1908_p_spl_
  );


  and

  (
    g2377_p,
    g2376_n_spl_,
    g2375_n_spl_
  );


  or

  (
    g2377_n,
    g2376_p_spl_,
    g2375_p_spl_
  );


  and

  (
    g2378_p,
    g2377_n_spl_0,
    g2375_n_spl_
  );


  or

  (
    g2378_n,
    g2377_p_spl_0,
    g2375_p_spl_
  );


  and

  (
    g2379_p,
    g2377_n_spl_0,
    g2376_n_spl_
  );


  or

  (
    g2379_n,
    g2377_p_spl_0,
    g2376_p_spl_
  );


  and

  (
    g2380_p,
    g2379_n,
    g2378_n
  );


  or

  (
    g2380_n,
    g2379_p,
    g2378_p
  );


  and

  (
    g2381_p,
    n2548_lo_buf_o2_p_spl_01,
    n2746_lo_p_spl_101
  );


  or

  (
    g2381_n,
    n2548_lo_buf_o2_n_spl_1,
    n2746_lo_n_spl_110
  );


  and

  (
    g2382_p,
    g2381_n_spl_,
    g2380_n_spl_
  );


  or

  (
    g2382_n,
    g2381_p_spl_,
    g2380_p_spl_
  );


  and

  (
    g2383_p,
    g2382_n_spl_0,
    g2377_n_spl_
  );


  or

  (
    g2383_n,
    g2382_p_spl_0,
    g2377_p_spl_
  );


  and

  (
    g2384_p,
    g2383_n_spl_,
    g2372_n_spl_
  );


  or

  (
    g2384_n,
    g2383_p_spl_,
    g2372_p_spl_
  );


  and

  (
    g2385_p,
    g2384_n_spl_0,
    g2372_n_spl_
  );


  or

  (
    g2385_n,
    g2384_p_spl_,
    g2372_p_spl_
  );


  and

  (
    g2386_p,
    g2384_n_spl_0,
    g2383_n_spl_
  );


  or

  (
    g2386_n,
    g2384_p_spl_,
    g2383_p_spl_
  );


  and

  (
    g2387_p,
    g2386_n,
    g2385_n
  );


  or

  (
    g2387_n,
    g2386_p,
    g2385_p
  );


  and

  (
    g2388_p,
    n2548_lo_buf_o2_p_spl_1,
    n2758_lo_p_spl_01
  );


  or

  (
    g2388_n,
    n2548_lo_buf_o2_n_spl_1,
    n2758_lo_n_spl_10
  );


  or

  (
    g2389_n,
    g2388_p,
    g2387_p
  );


  and

  (
    g2390_p,
    g2389_n_spl_0,
    g2384_n_spl_
  );


  and

  (
    g2391_p,
    g2163_n_spl_0,
    g2161_n
  );


  and

  (
    g2392_p,
    g2347_n_spl_0,
    g2346_n
  );


  and

  (
    g2393_p,
    g2163_n_spl_0,
    g2162_n
  );


  and

  (
    g2394_p,
    g2178_n_spl_0,
    g2177_n
  );


  and

  (
    g2395_p,
    g2193_n_spl_0,
    g2192_n
  );


  and

  (
    g2396_p,
    g2198_n_spl_0,
    g2197_n
  );


  and

  (
    g2397_p,
    g2178_n_spl_0,
    g2176_n
  );


  and

  (
    g2398_p,
    g2193_n_spl_0,
    g2191_n
  );


  and

  (
    g2399_p,
    g2198_n_spl_0,
    g2196_n
  );


  and

  (
    g2400_p,
    g2347_n_spl_,
    g2345_n
  );


  and

  (
    g2401_p,
    g2201_n_spl_,
    g2135_n_spl_
  );


  and

  (
    g2402_p,
    g2204_n_spl_,
    g2136_n_spl_
  );


  and

  (
    g2403_p,
    g2207_n_spl_,
    g2137_n_spl_
  );


  and

  (
    g2404_p,
    g2210_n_spl_,
    g2138_n_spl_
  );


  and

  (
    g2405_p,
    g1846_n_spl_0,
    g1833_n_spl_
  );


  or

  (
    g2405_n,
    g1846_p_spl_,
    g1833_p_spl_
  );


  and

  (
    g2406_p,
    g1846_n_spl_0,
    g1845_n_spl_
  );


  or

  (
    g2406_n,
    g1846_p_spl_,
    g1845_p_spl_
  );


  and

  (
    g2407_p,
    g2406_n,
    g2405_n
  );


  or

  (
    g2407_n,
    g2406_p,
    g2405_p
  );


  and

  (
    g2408_p,
    G20_p_spl_00,
    G15_p_spl_0
  );


  or

  (
    g2408_n,
    G20_n_spl_00,
    G15_n_spl_1
  );


  or

  (
    g2409_n,
    g2408_p,
    g2407_p
  );


  and

  (
    g2410_p,
    n2668_lo_buf_o2_p_spl_0,
    n2734_lo_p_spl_111
  );


  or

  (
    g2410_n,
    n2668_lo_buf_o2_n_spl_,
    n2734_lo_n_spl_111
  );


  and

  (
    g2411_p,
    g1854_n_spl_,
    g1849_n_spl_
  );


  or

  (
    g2411_n,
    g1854_p_spl_,
    g1849_p_spl_
  );


  and

  (
    g2412_p,
    g2411_n_spl_,
    g2410_n_spl_
  );


  or

  (
    g2412_n,
    g2411_p_spl_,
    g2410_p_spl_
  );


  and

  (
    g2413_p,
    g2412_n_spl_0,
    g2410_n_spl_
  );


  or

  (
    g2413_n,
    g2412_p_spl_,
    g2410_p_spl_
  );


  and

  (
    g2414_p,
    g2412_n_spl_0,
    g2411_n_spl_
  );


  or

  (
    g2414_n,
    g2412_p_spl_,
    g2411_p_spl_
  );


  and

  (
    g2415_p,
    g2414_n,
    g2413_n
  );


  or

  (
    g2415_n,
    g2414_p,
    g2413_p
  );


  and

  (
    g2416_p,
    n2656_lo_buf_o2_p_spl_1,
    n2746_lo_p_spl_110
  );


  or

  (
    g2416_n,
    n2656_lo_buf_o2_n_spl_,
    n2746_lo_n_spl_110
  );


  and

  (
    g2417_p,
    g2416_n_spl_,
    g2415_n_spl_
  );


  or

  (
    g2417_n,
    g2416_p_spl_,
    g2415_p_spl_
  );


  and

  (
    g2418_p,
    g2417_n_spl_0,
    g2415_n_spl_
  );


  or

  (
    g2418_n,
    g2417_p_spl_,
    g2415_p_spl_
  );


  and

  (
    g2419_p,
    g2417_n_spl_0,
    g2416_n_spl_
  );


  or

  (
    g2419_n,
    g2417_p_spl_,
    g2416_p_spl_
  );


  and

  (
    g2420_p,
    g2419_n,
    g2418_n
  );


  or

  (
    g2420_n,
    g2419_p,
    g2418_p
  );


  and

  (
    g2421_p,
    g1864_n_spl_,
    g1859_n_spl_
  );


  or

  (
    g2421_n,
    g1864_p_spl_,
    g1859_p_spl_
  );


  or

  (
    g2422_n,
    g2421_p,
    g2420_p
  );


  and

  (
    g2423_p,
    g1799_n_spl_0,
    g1797_n_spl_
  );


  or

  (
    g2423_n,
    g1799_p_spl_0,
    g1797_p_spl_
  );


  and

  (
    g2424_p,
    g1799_n_spl_,
    g1798_n_spl_
  );


  or

  (
    g2424_n,
    g1799_p_spl_,
    g1798_p_spl_
  );


  and

  (
    g2425_p,
    g2424_n,
    g2423_n
  );


  or

  (
    g2425_n,
    g2424_p,
    g2423_p
  );


  and

  (
    g2426_p,
    g2022_n_spl_,
    g2017_n_spl_
  );


  or

  (
    g2426_n,
    g2022_p_spl_,
    g2017_p_spl_
  );


  and

  (
    g2427_p,
    g2426_n_spl_,
    g2425_n_spl_
  );


  or

  (
    g2427_n,
    g2426_p_spl_,
    g2425_p_spl_
  );


  and

  (
    g2428_p,
    g2427_n_spl_0,
    g2425_n_spl_
  );


  or

  (
    g2428_n,
    g2427_p_spl_,
    g2425_p_spl_
  );


  and

  (
    g2429_p,
    g2427_n_spl_0,
    g2426_n_spl_
  );


  or

  (
    g2429_n,
    g2427_p_spl_,
    g2426_p_spl_
  );


  and

  (
    g2430_p,
    g2429_n,
    g2428_n
  );


  or

  (
    g2430_n,
    g2429_p,
    g2428_p
  );


  and

  (
    g2431_p,
    n2608_lo_buf_o2_p_spl_1,
    n2758_lo_p_spl_01
  );


  or

  (
    g2431_n,
    n2608_lo_buf_o2_n_spl_1,
    n2758_lo_n_spl_10
  );


  and

  (
    g2432_p,
    g2431_n_spl_,
    g2430_n_spl_
  );


  or

  (
    g2432_n,
    g2431_p_spl_,
    g2430_p_spl_
  );


  and

  (
    g2433_p,
    g2432_n_spl_0,
    g2430_n_spl_
  );


  or

  (
    g2433_n,
    g2432_p_spl_,
    g2430_p_spl_
  );


  and

  (
    g2434_p,
    g2432_n_spl_0,
    g2431_n_spl_
  );


  or

  (
    g2434_n,
    g2432_p_spl_,
    g2431_p_spl_
  );


  and

  (
    g2435_p,
    g2434_n,
    g2433_n
  );


  or

  (
    g2435_n,
    g2434_p,
    g2433_p
  );


  and

  (
    g2436_p,
    g2060_n_spl_,
    g2055_n_spl_
  );


  or

  (
    g2436_n,
    g2060_p_spl_,
    g2055_p_spl_
  );


  or

  (
    g2437_n,
    g2436_p,
    g2435_p
  );


  and

  (
    g2438_p,
    g2239_n_spl_0,
    g2237_n_spl_
  );


  or

  (
    g2438_n,
    g2239_p_spl_0,
    g2237_p_spl_
  );


  and

  (
    g2439_p,
    g2239_n_spl_,
    g2238_n_spl_
  );


  or

  (
    g2439_n,
    g2239_p_spl_,
    g2238_p_spl_
  );


  and

  (
    g2440_p,
    g2439_n,
    g2438_n
  );


  or

  (
    g2440_n,
    g2439_p,
    g2438_p
  );


  and

  (
    g2441_p,
    g2232_n_spl_0,
    g2230_n_spl_
  );


  or

  (
    g2441_n,
    g2232_p_spl_0,
    g2230_p_spl_
  );


  and

  (
    g2442_p,
    g2232_n_spl_,
    g2231_n_spl_
  );


  or

  (
    g2442_n,
    g2232_p_spl_,
    g2231_p_spl_
  );


  and

  (
    g2443_p,
    g2442_n,
    g2441_n
  );


  or

  (
    g2443_n,
    g2442_p,
    g2441_p
  );


  and

  (
    g2444_p,
    g2126_n_spl_,
    g2121_n_spl_
  );


  or

  (
    g2444_n,
    g2126_p_spl_,
    g2121_p_spl_
  );


  and

  (
    g2445_p,
    g2444_n_spl_,
    g2443_n_spl_
  );


  or

  (
    g2445_n,
    g2444_p_spl_,
    g2443_p_spl_
  );


  and

  (
    g2446_p,
    g2445_n_spl_0,
    g2443_n_spl_
  );


  or

  (
    g2446_n,
    g2445_p_spl_0,
    g2443_p_spl_
  );


  and

  (
    g2447_p,
    g2445_n_spl_0,
    g2444_n_spl_
  );


  or

  (
    g2447_n,
    g2445_p_spl_0,
    g2444_p_spl_
  );


  and

  (
    g2448_p,
    g2447_n,
    g2446_n
  );


  or

  (
    g2448_n,
    g2447_p,
    g2446_p
  );


  and

  (
    g2449_p,
    n2500_lo_buf_o2_p_spl_1,
    n2746_lo_p_spl_110
  );


  or

  (
    g2449_n,
    n2500_lo_buf_o2_n_spl_1,
    n2746_lo_n_spl_11
  );


  and

  (
    g2450_p,
    g2449_n_spl_,
    g2448_n_spl_
  );


  or

  (
    g2450_n,
    g2449_p,
    g2448_p
  );


  and

  (
    g2451_p,
    g2450_n_spl_0,
    g2445_n_spl_
  );


  or

  (
    g2451_n,
    g2450_p,
    g2445_p_spl_
  );


  or

  (
    g2452_n,
    g2451_p,
    g2440_p
  );


  and

  (
    g2453_p,
    g2284_n_spl_0,
    g2282_n_spl_
  );


  or

  (
    g2453_n,
    g2284_p_spl_0,
    g2282_p_spl_
  );


  and

  (
    g2454_p,
    g2284_n_spl_,
    g2283_n_spl_
  );


  or

  (
    g2454_n,
    g2284_p_spl_,
    g2283_p_spl_
  );


  and

  (
    g2455_p,
    g2454_n,
    g2453_n
  );


  or

  (
    g2455_n,
    g2454_p,
    g2453_p
  );


  and

  (
    g2456_p,
    g2277_n_spl_0,
    g2275_n_spl_
  );


  or

  (
    g2456_n,
    g2277_p_spl_0,
    g2275_p_spl_
  );


  and

  (
    g2457_p,
    g2277_n_spl_,
    g2276_n_spl_
  );


  or

  (
    g2457_n,
    g2277_p_spl_,
    g2276_p_spl_
  );


  and

  (
    g2458_p,
    g2457_n,
    g2456_n
  );


  or

  (
    g2458_n,
    g2457_p,
    g2456_p
  );


  and

  (
    g2459_p,
    g2369_n_spl_,
    g2364_n_spl_
  );


  or

  (
    g2459_n,
    g2369_p_spl_,
    g2364_p_spl_
  );


  and

  (
    g2460_p,
    g2459_n_spl_,
    g2458_n_spl_
  );


  or

  (
    g2460_n,
    g2459_p_spl_,
    g2458_p_spl_
  );


  and

  (
    g2461_p,
    g2460_n_spl_0,
    g2458_n_spl_
  );


  or

  (
    g2461_n,
    g2460_p_spl_0,
    g2458_p_spl_
  );


  and

  (
    g2462_p,
    g2460_n_spl_0,
    g2459_n_spl_
  );


  or

  (
    g2462_n,
    g2460_p_spl_0,
    g2459_p_spl_
  );


  and

  (
    g2463_p,
    g2462_n,
    g2461_n
  );


  or

  (
    g2463_n,
    g2462_p,
    g2461_p
  );


  and

  (
    g2464_p,
    n2560_lo_buf_o2_p_spl_1,
    n2758_lo_p_spl_10
  );


  or

  (
    g2464_n,
    n2560_lo_buf_o2_n_spl_1,
    n2758_lo_n_spl_11
  );


  and

  (
    g2465_p,
    g2464_n,
    g2463_n
  );


  or

  (
    g2465_n,
    g2464_p_spl_,
    g2463_p_spl_
  );


  and

  (
    g2466_p,
    g2465_n,
    g2460_n_spl_
  );


  or

  (
    g2466_n,
    g2465_p_spl_0,
    g2460_p_spl_
  );


  or

  (
    g2467_n,
    g2466_p,
    g2455_p
  );


  and

  (
    g2468_p,
    g1806_n_spl_0,
    g1804_n
  );


  and

  (
    g2469_p,
    g1806_n_spl_0,
    g1805_n
  );


  or

  (
    g2470_n,
    g2469_p,
    g2468_p
  );


  and

  (
    g2471_p,
    g1811_n_spl_0,
    g1809_n
  );


  and

  (
    g2472_p,
    g1811_n_spl_0,
    g1810_n
  );


  or

  (
    g2473_n,
    g2472_p,
    g2471_p
  );


  and

  (
    g2474_p,
    g1816_n_spl_0,
    g1814_n
  );


  and

  (
    g2475_p,
    g1816_n_spl_0,
    g1815_n
  );


  or

  (
    g2476_n,
    g2475_p,
    g2474_p
  );


  and

  (
    g2477_p,
    g1831_n_spl_0,
    g1819_n
  );


  and

  (
    g2478_p,
    g1831_n_spl_0,
    g1830_n
  );


  or

  (
    g2479_n,
    g2478_p,
    g2477_p
  );


  and

  (
    g2480_p,
    g2295_n_spl_,
    g2294_n_spl_
  );


  or

  (
    g2480_n,
    g2295_p_spl_,
    g2294_p_spl_
  );


  and

  (
    g2481_p,
    g2480_n,
    g2296_n_spl_
  );


  or

  (
    g2481_n,
    g2480_p,
    g2296_p_spl_
  );


  and

  (
    g2482_p,
    G17_p_spl_011,
    G5_p_spl_0
  );


  or

  (
    g2482_n,
    G17_n_spl_011,
    G5_n_spl_0
  );


  and

  (
    g2483_p,
    G18_p_spl_011,
    G4_p_spl_0
  );


  or

  (
    g2483_n,
    G18_n_spl_100,
    G4_n_spl_
  );


  and

  (
    g2484_p,
    g2483_n_spl_,
    g2482_p_spl_
  );


  or

  (
    g2484_n,
    g2483_p_spl_,
    g2482_n_spl_
  );


  and

  (
    g2485_p,
    g2484_n_spl_,
    g2482_p_spl_
  );


  or

  (
    g2485_n,
    g2484_p_spl_,
    g2482_n_spl_
  );


  or

  (
    g2486_n,
    g2485_p_spl_,
    g2481_p
  );


  and

  (
    g2487_p,
    g2328_n_spl_0,
    g2326_n_spl_
  );


  or

  (
    g2487_n,
    g2328_p_spl_0,
    g2326_p_spl_
  );


  and

  (
    g2488_p,
    g2328_n_spl_,
    g2327_n_spl_
  );


  or

  (
    g2488_n,
    g2328_p_spl_,
    g2327_p_spl_
  );


  and

  (
    g2489_p,
    g2488_n,
    g2487_n
  );


  or

  (
    g2489_n,
    g2488_p,
    g2487_p
  );


  and

  (
    g2490_p,
    g2321_n_spl_,
    g2320_n_spl_
  );


  or

  (
    g2490_n,
    g2321_p_spl_,
    g2320_p_spl_
  );


  and

  (
    g2491_p,
    g2490_n,
    g2322_n_spl_
  );


  or

  (
    g2491_n,
    g2490_p,
    g2322_p_spl_
  );


  and

  (
    g2492_p,
    G17_p_spl_011,
    G10_p_spl_1
  );


  or

  (
    g2492_n,
    G17_n_spl_011,
    G10_n_spl_1
  );


  and

  (
    g2493_p,
    G18_p_spl_100,
    G9_p_spl_00
  );


  or

  (
    g2493_n,
    G18_n_spl_100,
    G9_n_spl_0
  );


  and

  (
    g2494_p,
    g2493_n_spl_,
    g2492_p_spl_
  );


  or

  (
    g2494_n,
    g2493_p_spl_,
    g2492_n_spl_
  );


  and

  (
    g2495_p,
    g2494_n_spl_,
    g2492_p_spl_
  );


  or

  (
    g2495_n,
    g2494_p_spl_,
    g2492_n_spl_
  );


  and

  (
    g2496_p,
    g2495_n_spl_0,
    g2491_n_spl_
  );


  or

  (
    g2496_n,
    g2495_p_spl_0,
    g2491_p_spl_
  );


  and

  (
    g2497_p,
    g2496_n_spl_0,
    g2491_n_spl_
  );


  or

  (
    g2497_n,
    g2496_p_spl_0,
    g2491_p_spl_
  );


  and

  (
    g2498_p,
    g2496_n_spl_0,
    g2495_n_spl_0
  );


  or

  (
    g2498_n,
    g2496_p_spl_0,
    g2495_p_spl_0
  );


  and

  (
    g2499_p,
    g2498_n,
    g2497_n
  );


  or

  (
    g2499_n,
    g2498_p,
    g2497_p
  );


  and

  (
    g2500_p,
    G19_p_spl_010,
    G9_p_spl_00
  );


  or

  (
    g2500_n,
    G19_n_spl_010,
    G9_n_spl_0
  );


  and

  (
    g2501_p,
    g2500_n_spl_,
    g2499_n_spl_
  );


  or

  (
    g2501_n,
    g2500_p_spl_,
    g2499_p_spl_
  );


  and

  (
    g2502_p,
    g2501_n_spl_0,
    g2496_n_spl_
  );


  or

  (
    g2502_n,
    g2501_p_spl_0,
    g2496_p_spl_
  );


  or

  (
    g2503_n,
    g2502_p,
    g2489_p
  );


  or

  (
    g2504_n,
    g2465_p_spl_0,
    g2463_p_spl_
  );


  or

  (
    g2505_n,
    g2465_p_spl_,
    g2464_p_spl_
  );


  and

  (
    g2506_p,
    g2505_n,
    g2504_n
  );


  and

  (
    g2507_p,
    g2450_n_spl_0,
    g2448_n_spl_
  );


  and

  (
    g2508_p,
    g2450_n_spl_,
    g2449_n_spl_
  );


  or

  (
    g2509_n,
    g2508_p,
    g2507_p
  );


  and

  (
    g2510_p,
    g1869_n_spl_0,
    g1867_n
  );


  and

  (
    g2511_p,
    g1869_n_spl_0,
    g1868_n
  );


  or

  (
    g2512_n,
    g2511_p,
    g2510_p
  );


  and

  (
    g2513_p,
    g1996_n_spl_0,
    g1954_n
  );


  and

  (
    g2514_p,
    g1996_n_spl_0,
    g1995_n
  );


  or

  (
    g2515_n,
    g2514_p,
    g2513_p
  );


  and

  (
    g2516_p,
    g2106_n_spl_0,
    g2063_n
  );


  and

  (
    g2517_p,
    g2106_n_spl_0,
    g2105_n
  );


  or

  (
    g2518_n,
    g2517_p,
    g2516_p
  );


  and

  (
    g2519_p,
    G17_p_spl_100,
    G2_p_spl_0
  );


  or

  (
    g2519_n,
    G17_n_spl_100,
    G2_n_spl_
  );


  and

  (
    g2520_p,
    n2668_lo_buf_o2_p_spl_1,
    n2746_lo_p_spl_11
  );


  and

  (
    g2521_p,
    n2572_lo_buf_o2_p_spl_10,
    n2770_lo_p_spl_
  );


  and

  (
    g2522_p,
    n2512_lo_buf_o2_p_spl_10,
    n2758_lo_p_spl_10
  );


  or

  (
    g2523_n,
    G20_n_spl_00,
    G10_n_spl_1
  );


  or

  (
    g2524_n,
    G19_n_spl_010,
    G5_n_spl_
  );


  and

  (
    g2525_p,
    g2417_n_spl_,
    g2412_n_spl_
  );


  and

  (
    g2526_p,
    g2432_n_spl_,
    g2427_n_spl_
  );


  and

  (
    g2527_p,
    g2382_n_spl_0,
    g2380_n_spl_
  );


  or

  (
    g2527_n,
    g2382_p_spl_0,
    g2380_p_spl_
  );


  and

  (
    g2528_p,
    g2382_n_spl_,
    g2381_n_spl_
  );


  or

  (
    g2528_n,
    g2382_p_spl_,
    g2381_p_spl_
  );


  and

  (
    g2529_p,
    g2528_n,
    g2527_n
  );


  or

  (
    g2529_n,
    g2528_p,
    g2527_p
  );


  and

  (
    g2530_p,
    g1951_n_spl_,
    g1946_n_spl_
  );


  or

  (
    g2530_n,
    g1951_p_spl_,
    g1946_p_spl_
  );


  and

  (
    g2531_p,
    g2530_n_spl_,
    g2529_n_spl_
  );


  or

  (
    g2531_n,
    g2530_p_spl_,
    g2529_p_spl_
  );


  and

  (
    g2532_p,
    g2531_n_spl_0,
    g2529_n_spl_
  );


  or

  (
    g2532_n,
    g2531_p_spl_,
    g2529_p_spl_
  );


  and

  (
    g2533_p,
    g2531_n_spl_0,
    g2530_n_spl_
  );


  or

  (
    g2533_n,
    g2531_p_spl_,
    g2530_p_spl_
  );


  and

  (
    g2534_p,
    g2533_n,
    g2532_n
  );


  or

  (
    g2534_n,
    g2533_p,
    g2532_p
  );


  and

  (
    g2535_p,
    n2536_lo_buf_o2_p_spl_1,
    n2758_lo_p_spl_11
  );


  or

  (
    g2535_n,
    n2536_lo_buf_o2_n_spl_1,
    n2758_lo_n_spl_11
  );


  or

  (
    g2536_n,
    g2535_p,
    g2534_p
  );


  and

  (
    g2537_p,
    g2536_n_spl_0,
    g2531_n_spl_
  );


  and

  (
    g2538_p,
    G17_p_spl_100,
    G3_p_spl_0
  );


  or

  (
    g2538_n,
    G17_n_spl_100,
    G3_n_spl_
  );


  and

  (
    g2539_p,
    G18_p_spl_100,
    G2_p_spl_0
  );


  or

  (
    g2539_n,
    G18_n_spl_101,
    G2_n_spl_
  );


  and

  (
    g2540_p,
    g2539_n,
    g2538_p
  );


  or

  (
    g2541_n,
    g2540_p_spl_,
    g2538_n
  );


  and

  (
    g2542_p,
    G17_p_spl_101,
    G9_p_spl_0
  );


  or

  (
    g2542_n,
    G17_n_spl_101,
    G9_n_spl_
  );


  and

  (
    g2543_p,
    G18_p_spl_101,
    G8_p_spl_0
  );


  or

  (
    g2543_n,
    G18_n_spl_101,
    G8_n_spl_0
  );


  and

  (
    g2544_p,
    g2543_n_spl_,
    g2542_p_spl_
  );


  or

  (
    g2544_n,
    g2543_p_spl_,
    g2542_n_spl_
  );


  and

  (
    g2545_p,
    g2544_n_spl_,
    g2542_p_spl_
  );


  or

  (
    g2545_n,
    g2544_p_spl_,
    g2542_n_spl_
  );


  and

  (
    g2546_p,
    g2544_n_spl_,
    g2543_n_spl_
  );


  or

  (
    g2546_n,
    g2544_p_spl_,
    g2543_p_spl_
  );


  and

  (
    g2547_p,
    g2546_n,
    g2545_n_spl_0
  );


  or

  (
    g2547_n,
    g2546_p,
    g2545_p_spl_0
  );


  and

  (
    g2548_p,
    G17_p_spl_101,
    G8_p_spl_0
  );


  or

  (
    g2548_n,
    G17_n_spl_101,
    G8_n_spl_0
  );


  and

  (
    g2549_p,
    G18_p_spl_101,
    G7_p_spl_0
  );


  or

  (
    g2549_n,
    G18_n_spl_110,
    G7_n_spl_0
  );


  and

  (
    g2550_p,
    g2549_n_spl_,
    g2548_p_spl_
  );


  or

  (
    g2550_n,
    g2549_p_spl_,
    g2548_n_spl_
  );


  and

  (
    g2551_p,
    g2550_n_spl_,
    g2548_p_spl_
  );


  or

  (
    g2551_n,
    g2550_p_spl_,
    g2548_n_spl_
  );


  and

  (
    g2552_p,
    g2551_n_spl_0,
    g2547_n_spl_
  );


  or

  (
    g2552_n,
    g2551_p_spl_0,
    g2547_p_spl_
  );


  and

  (
    g2553_p,
    g2552_n_spl_0,
    g2547_n_spl_
  );


  or

  (
    g2553_n,
    g2552_p_spl_,
    g2547_p_spl_
  );


  and

  (
    g2554_p,
    g2552_n_spl_0,
    g2551_n_spl_0
  );


  or

  (
    g2554_n,
    g2552_p_spl_,
    g2551_p_spl_0
  );


  and

  (
    g2555_p,
    g2554_n,
    g2553_n
  );


  or

  (
    g2555_n,
    g2554_p,
    g2553_p
  );


  and

  (
    g2556_p,
    G19_p_spl_010,
    G7_p_spl_1
  );


  or

  (
    g2556_n,
    G19_n_spl_011,
    G7_n_spl_
  );


  or

  (
    g2557_n,
    g2556_p,
    g2555_p
  );


  and

  (
    g2558_p,
    g2557_n_spl_0,
    g2552_n_spl_
  );


  and

  (
    g2559_p,
    G17_p_spl_110,
    G15_p_spl_1
  );


  or

  (
    g2559_n,
    G17_n_spl_110,
    G15_n_spl_1
  );


  and

  (
    g2560_p,
    G18_p_spl_110,
    G14_p_spl_00
  );


  or

  (
    g2560_n,
    G18_n_spl_110,
    G14_n_spl_0
  );


  and

  (
    g2561_p,
    g2560_n_spl_,
    g2559_p_spl_
  );


  or

  (
    g2561_n,
    g2560_p_spl_,
    g2559_n_spl_
  );


  and

  (
    g2562_p,
    g2561_n_spl_,
    g2559_p_spl_
  );


  or

  (
    g2562_n,
    g2561_p_spl_,
    g2559_n_spl_
  );


  and

  (
    g2563_p,
    g2561_n_spl_,
    g2560_n_spl_
  );


  or

  (
    g2563_n,
    g2561_p_spl_,
    g2560_p_spl_
  );


  and

  (
    g2564_p,
    g2563_n,
    g2562_n_spl_0
  );


  or

  (
    g2564_n,
    g2563_p,
    g2562_p_spl_0
  );


  and

  (
    g2565_p,
    G17_p_spl_110,
    G14_p_spl_00
  );


  or

  (
    g2565_n,
    G17_n_spl_110,
    G14_n_spl_0
  );


  and

  (
    g2566_p,
    G18_p_spl_110,
    G13_p_spl_00
  );


  or

  (
    g2566_n,
    G18_n_spl_111,
    G13_n_spl_0
  );


  and

  (
    g2567_p,
    g2566_n_spl_,
    g2565_p_spl_
  );


  or

  (
    g2567_n,
    g2566_p_spl_,
    g2565_n_spl_
  );


  and

  (
    g2568_p,
    g2567_n_spl_,
    g2565_p_spl_
  );


  or

  (
    g2568_n,
    g2567_p_spl_,
    g2565_n_spl_
  );


  and

  (
    g2569_p,
    g2568_n_spl_0,
    g2564_n_spl_
  );


  or

  (
    g2569_n,
    g2568_p_spl_0,
    g2564_p_spl_
  );


  and

  (
    g2570_p,
    g2569_n_spl_0,
    g2564_n_spl_
  );


  or

  (
    g2570_n,
    g2569_p_spl_0,
    g2564_p_spl_
  );


  and

  (
    g2571_p,
    g2569_n_spl_0,
    g2568_n_spl_0
  );


  or

  (
    g2571_n,
    g2569_p_spl_0,
    g2568_p_spl_0
  );


  and

  (
    g2572_p,
    g2571_n,
    g2570_n
  );


  or

  (
    g2572_n,
    g2571_p,
    g2570_p
  );


  and

  (
    g2573_p,
    G19_p_spl_011,
    G13_p_spl_0
  );


  or

  (
    g2573_n,
    G19_n_spl_011,
    G13_n_spl_1
  );


  and

  (
    g2574_p,
    g2573_n_spl_,
    g2572_n_spl_
  );


  or

  (
    g2574_n,
    g2573_p_spl_,
    g2572_p_spl_
  );


  and

  (
    g2575_p,
    g2574_n_spl_0,
    g2572_n_spl_
  );


  or

  (
    g2575_n,
    g2574_p_spl_0,
    g2572_p_spl_
  );


  and

  (
    g2576_p,
    g2574_n_spl_0,
    g2573_n_spl_
  );


  or

  (
    g2576_n,
    g2574_p_spl_0,
    g2573_p_spl_
  );


  and

  (
    g2577_p,
    g2576_n,
    g2575_n
  );


  or

  (
    g2577_n,
    g2576_p,
    g2575_p
  );


  and

  (
    g2578_p,
    g2567_n_spl_,
    g2566_n_spl_
  );


  or

  (
    g2578_n,
    g2567_p_spl_,
    g2566_p_spl_
  );


  and

  (
    g2579_p,
    g2578_n,
    g2568_n_spl_
  );


  or

  (
    g2579_n,
    g2578_p,
    g2568_p_spl_
  );


  and

  (
    g2580_p,
    g2579_n_spl_,
    g2301_n_spl_0
  );


  or

  (
    g2580_n,
    g2579_p_spl_,
    g2301_p_spl_0
  );


  and

  (
    g2581_p,
    g2580_n_spl_0,
    g2579_n_spl_
  );


  or

  (
    g2581_n,
    g2580_p_spl_0,
    g2579_p_spl_
  );


  and

  (
    g2582_p,
    g2580_n_spl_0,
    g2301_n_spl_
  );


  or

  (
    g2582_n,
    g2580_p_spl_0,
    g2301_p_spl_
  );


  and

  (
    g2583_p,
    g2582_n,
    g2581_n
  );


  or

  (
    g2583_n,
    g2582_p,
    g2581_p
  );


  and

  (
    g2584_p,
    G19_p_spl_011,
    G12_p_spl_0
  );


  or

  (
    g2584_n,
    G19_n_spl_10,
    G12_n_spl_1
  );


  and

  (
    g2585_p,
    g2584_n_spl_,
    g2583_n_spl_
  );


  or

  (
    g2585_n,
    g2584_p_spl_,
    g2583_p_spl_
  );


  and

  (
    g2586_p,
    g2585_n_spl_0,
    g2580_n_spl_
  );


  or

  (
    g2586_n,
    g2585_p_spl_0,
    g2580_p_spl_
  );


  and

  (
    g2587_p,
    g2586_n_spl_,
    g2577_n_spl_
  );


  or

  (
    g2587_n,
    g2586_p_spl_,
    g2577_p_spl_
  );


  and

  (
    g2588_p,
    g2587_n_spl_0,
    g2577_n_spl_
  );


  or

  (
    g2588_n,
    g2587_p_spl_,
    g2577_p_spl_
  );


  and

  (
    g2589_p,
    g2587_n_spl_0,
    g2586_n_spl_
  );


  or

  (
    g2589_n,
    g2587_p_spl_,
    g2586_p_spl_
  );


  and

  (
    g2590_p,
    g2589_n,
    g2588_n
  );


  or

  (
    g2590_n,
    g2589_p,
    g2588_p
  );


  and

  (
    g2591_p,
    G20_p_spl_00,
    G12_p_spl_1
  );


  or

  (
    g2591_n,
    G20_n_spl_01,
    G12_n_spl_1
  );


  or

  (
    g2592_n,
    g2591_p,
    g2590_p
  );


  and

  (
    g2593_p,
    g2592_n_spl_0,
    g2587_n_spl_
  );


  and

  (
    g2594_p,
    g2536_n_spl_0,
    g2535_n
  );


  and

  (
    g2595_p,
    g2422_n_spl_0,
    g2421_n
  );


  and

  (
    g2596_p,
    g2437_n_spl_0,
    g2436_n
  );


  and

  (
    g2597_p,
    g2452_n_spl_0,
    g2451_n
  );


  and

  (
    g2598_p,
    g2467_n_spl_0,
    g2466_n
  );


  and

  (
    g2599_p,
    g2422_n_spl_0,
    g2420_n
  );


  and

  (
    g2600_p,
    g2437_n_spl_0,
    g2435_n
  );


  and

  (
    g2601_p,
    g2467_n_spl_0,
    g2455_n
  );


  and

  (
    g2602_p,
    g2452_n_spl_0,
    g2440_n
  );


  and

  (
    g2603_p,
    g2536_n_spl_,
    g2534_n
  );


  and

  (
    g2604_p,
    g2512_n_spl_,
    g2332_n_spl_
  );


  and

  (
    g2605_p,
    g2518_n_spl_,
    g2333_n_spl_
  );


  and

  (
    g2606_p,
    g2515_n_spl_,
    g2334_n_spl_
  );


  and

  (
    g2607_p,
    g2519_p_spl_,
    g2335_n_spl_
  );


  and

  (
    g2608_p,
    g2509_n_spl_,
    g2349_n_spl_
  );


  or

  (
    g2609_n,
    g2506_p_spl_,
    g2390_p_spl_
  );


  and

  (
    g2610_p,
    g2484_n_spl_,
    g2483_n_spl_
  );


  or

  (
    g2610_n,
    g2484_p_spl_,
    g2483_p_spl_
  );


  and

  (
    g2611_p,
    g2610_n,
    g2485_n_spl_
  );


  or

  (
    g2611_n,
    g2610_p,
    g2485_p_spl_
  );


  and

  (
    g2612_p,
    G17_p_spl_111,
    G4_p_spl_0
  );


  or

  (
    g2612_n,
    G17_n_spl_11,
    G4_n_spl_
  );


  and

  (
    g2613_p,
    G18_p_spl_11,
    G3_p_spl_0
  );


  or

  (
    g2613_n,
    G18_n_spl_111,
    G3_n_spl_
  );


  and

  (
    g2614_p,
    g2613_n_spl_,
    g2612_p_spl_
  );


  or

  (
    g2614_n,
    g2613_p,
    g2612_n_spl_
  );


  and

  (
    g2615_p,
    g2614_n_spl_,
    g2612_p_spl_
  );


  or

  (
    g2615_n,
    g2614_p,
    g2612_n_spl_
  );


  or

  (
    g2616_n,
    g2615_p_spl_,
    g2611_p
  );


  and

  (
    g2617_p,
    g2501_n_spl_0,
    g2499_n_spl_
  );


  or

  (
    g2617_n,
    g2501_p_spl_0,
    g2499_p_spl_
  );


  and

  (
    g2618_p,
    g2501_n_spl_,
    g2500_n_spl_
  );


  or

  (
    g2618_n,
    g2501_p_spl_,
    g2500_p_spl_
  );


  and

  (
    g2619_p,
    g2618_n,
    g2617_n
  );


  or

  (
    g2619_n,
    g2618_p,
    g2617_p
  );


  and

  (
    g2620_p,
    g2494_n_spl_,
    g2493_n_spl_
  );


  or

  (
    g2620_n,
    g2494_p_spl_,
    g2493_p_spl_
  );


  and

  (
    g2621_p,
    g2620_n,
    g2495_n_spl_
  );


  or

  (
    g2621_n,
    g2620_p,
    g2495_p_spl_
  );


  and

  (
    g2622_p,
    g2621_n_spl_,
    g2545_n_spl_0
  );


  or

  (
    g2622_n,
    g2621_p_spl_,
    g2545_p_spl_0
  );


  and

  (
    g2623_p,
    g2622_n_spl_0,
    g2621_n_spl_
  );


  or

  (
    g2623_n,
    g2622_p_spl_0,
    g2621_p_spl_
  );


  and

  (
    g2624_p,
    g2622_n_spl_0,
    g2545_n_spl_
  );


  or

  (
    g2624_n,
    g2622_p_spl_0,
    g2545_p_spl_
  );


  and

  (
    g2625_p,
    g2624_n,
    g2623_n
  );


  or

  (
    g2625_n,
    g2624_p,
    g2623_p
  );


  and

  (
    g2626_p,
    G19_p_spl_100,
    G8_p_spl_1
  );


  or

  (
    g2626_n,
    G19_n_spl_10,
    G8_n_spl_
  );


  and

  (
    g2627_p,
    g2626_n,
    g2625_n
  );


  or

  (
    g2627_n,
    g2626_p_spl_,
    g2625_p_spl_
  );


  and

  (
    g2628_p,
    g2627_n,
    g2622_n_spl_
  );


  or

  (
    g2628_n,
    g2627_p_spl_0,
    g2622_p_spl_
  );


  or

  (
    g2629_n,
    g2628_p,
    g2619_p
  );


  and

  (
    g2630_p,
    g1844_n_spl_0,
    g1842_n_spl_
  );


  or

  (
    g2630_n,
    g1844_p_spl_0,
    g1842_p_spl_
  );


  and

  (
    g2631_p,
    g1844_n_spl_,
    g1843_n_spl_
  );


  or

  (
    g2631_n,
    g1844_p_spl_,
    g1843_p_spl_
  );


  and

  (
    g2632_p,
    g2631_n,
    g2630_n
  );


  or

  (
    g2632_n,
    g2631_p,
    g2630_p
  );


  and

  (
    g2633_p,
    g1837_n_spl_,
    g1836_n_spl_
  );


  or

  (
    g2633_n,
    g1837_p_spl_,
    g1836_p_spl_
  );


  and

  (
    g2634_p,
    g2633_n,
    g1838_n_spl_
  );


  or

  (
    g2634_n,
    g2633_p,
    g1838_p_spl_
  );


  and

  (
    g2635_p,
    g2634_n_spl_,
    g2562_n_spl_0
  );


  or

  (
    g2635_n,
    g2634_p_spl_,
    g2562_p_spl_0
  );


  and

  (
    g2636_p,
    g2635_n_spl_0,
    g2634_n_spl_
  );


  or

  (
    g2636_n,
    g2635_p_spl_0,
    g2634_p_spl_
  );


  and

  (
    g2637_p,
    g2635_n_spl_0,
    g2562_n_spl_
  );


  or

  (
    g2637_n,
    g2635_p_spl_0,
    g2562_p_spl_
  );


  and

  (
    g2638_p,
    g2637_n,
    g2636_n
  );


  or

  (
    g2638_n,
    g2637_p,
    g2636_p
  );


  and

  (
    g2639_p,
    G19_p_spl_100,
    G14_p_spl_0
  );


  or

  (
    g2639_n,
    G19_n_spl_11,
    G14_n_spl_1
  );


  and

  (
    g2640_p,
    g2639_n_spl_,
    g2638_n_spl_
  );


  or

  (
    g2640_n,
    g2639_p_spl_,
    g2638_p_spl_
  );


  and

  (
    g2641_p,
    g2640_n_spl_0,
    g2635_n_spl_
  );


  or

  (
    g2641_n,
    g2640_p_spl_0,
    g2635_p_spl_
  );


  and

  (
    g2642_p,
    g2641_n_spl_,
    g2632_n_spl_
  );


  or

  (
    g2642_n,
    g2641_p_spl_,
    g2632_p_spl_
  );


  and

  (
    g2643_p,
    g2642_n_spl_0,
    g2632_n_spl_
  );


  or

  (
    g2643_n,
    g2642_p_spl_,
    g2632_p_spl_
  );


  and

  (
    g2644_p,
    g2642_n_spl_0,
    g2641_n_spl_
  );


  or

  (
    g2644_n,
    g2642_p_spl_,
    g2641_p_spl_
  );


  and

  (
    g2645_p,
    g2644_n,
    g2643_n
  );


  or

  (
    g2645_n,
    g2644_p,
    g2643_p
  );


  and

  (
    g2646_p,
    G20_p_spl_01,
    G14_p_spl_1
  );


  or

  (
    g2646_n,
    G20_n_spl_01,
    G14_n_spl_1
  );


  and

  (
    g2647_p,
    g2646_n_spl_,
    g2645_n_spl_
  );


  or

  (
    g2647_n,
    g2646_p_spl_,
    g2645_p_spl_
  );


  and

  (
    g2648_p,
    g2647_n_spl_0,
    g2645_n_spl_
  );


  or

  (
    g2648_n,
    g2647_p_spl_,
    g2645_p_spl_
  );


  and

  (
    g2649_p,
    g2647_n_spl_0,
    g2646_n_spl_
  );


  or

  (
    g2649_n,
    g2647_p_spl_,
    g2646_p_spl_
  );


  and

  (
    g2650_p,
    g2649_n,
    g2648_n
  );


  or

  (
    g2650_n,
    g2649_p,
    g2648_p
  );


  and

  (
    g2651_p,
    g2640_n_spl_0,
    g2638_n_spl_
  );


  or

  (
    g2651_n,
    g2640_p_spl_0,
    g2638_p_spl_
  );


  and

  (
    g2652_p,
    g2640_n_spl_,
    g2639_n_spl_
  );


  or

  (
    g2652_n,
    g2640_p_spl_,
    g2639_p_spl_
  );


  and

  (
    g2653_p,
    g2652_n,
    g2651_n
  );


  or

  (
    g2653_n,
    g2652_p,
    g2651_p
  );


  and

  (
    g2654_p,
    g2574_n_spl_,
    g2569_n_spl_
  );


  or

  (
    g2654_n,
    g2574_p_spl_,
    g2569_p_spl_
  );


  and

  (
    g2655_p,
    g2654_n_spl_,
    g2653_n_spl_
  );


  or

  (
    g2655_n,
    g2654_p_spl_,
    g2653_p_spl_
  );


  and

  (
    g2656_p,
    g2655_n_spl_0,
    g2653_n_spl_
  );


  or

  (
    g2656_n,
    g2655_p_spl_0,
    g2653_p_spl_
  );


  and

  (
    g2657_p,
    g2655_n_spl_0,
    g2654_n_spl_
  );


  or

  (
    g2657_n,
    g2655_p_spl_0,
    g2654_p_spl_
  );


  and

  (
    g2658_p,
    g2657_n,
    g2656_n
  );


  or

  (
    g2658_n,
    g2657_p,
    g2656_p
  );


  and

  (
    g2659_p,
    G20_p_spl_01,
    G13_p_spl_1
  );


  or

  (
    g2659_n,
    G20_n_spl_1,
    G13_n_spl_1
  );


  and

  (
    g2660_p,
    g2659_n,
    g2658_n
  );


  or

  (
    g2660_n,
    g2659_p_spl_,
    g2658_p_spl_
  );


  and

  (
    g2661_p,
    g2660_n,
    g2655_n_spl_
  );


  or

  (
    g2661_n,
    g2660_p_spl_0,
    g2655_p_spl_
  );


  or

  (
    g2662_n,
    g2661_p,
    g2650_p
  );


  and

  (
    g2663_p,
    g2215_n_spl_0,
    g2213_n
  );


  and

  (
    g2664_p,
    g2215_n_spl_0,
    g2214_n
  );


  or

  (
    g2665_n,
    g2664_p,
    g2663_p
  );


  and

  (
    g2666_p,
    g2389_n_spl_0,
    g2387_n
  );


  and

  (
    g2667_p,
    g2389_n_spl_,
    g2388_n
  );


  or

  (
    g2668_n,
    g2667_p,
    g2666_p
  );


  and

  (
    g2669_p,
    g2241_n_spl_0,
    g2219_n
  );


  and

  (
    g2670_p,
    g2241_n_spl_0,
    g2240_n
  );


  or

  (
    g2671_n,
    g2670_p,
    g2669_p
  );


  and

  (
    g2672_p,
    g2286_n_spl_0,
    g2244_n
  );


  and

  (
    g2673_p,
    g2286_n_spl_0,
    g2285_n
  );


  or

  (
    g2674_n,
    g2673_p,
    g2672_p
  );


  or

  (
    g2675_n,
    g2660_p_spl_0,
    g2658_p_spl_
  );


  or

  (
    g2676_n,
    g2660_p_spl_,
    g2659_p_spl_
  );


  and

  (
    g2677_p,
    g2676_n,
    g2675_n
  );


  and

  (
    g2678_p,
    g2614_n_spl_,
    g2613_n_spl_
  );


  or

  (
    g2679_n,
    g2678_p,
    g2615_p_spl_
  );


  or

  (
    g2680_n,
    g2627_p_spl_0,
    g2625_p_spl_
  );


  or

  (
    g2681_n,
    g2627_p_spl_,
    g2626_p_spl_
  );


  and

  (
    g2682_p,
    g2681_n,
    g2680_n
  );


  and

  (
    g2683_p,
    g2297_n_spl_0,
    g2292_n
  );


  and

  (
    g2684_p,
    g2297_n_spl_0,
    g2296_n_spl_
  );


  or

  (
    g2685_n,
    g2684_p,
    g2683_p
  );


  and

  (
    g2686_p,
    g2330_n_spl_0,
    g2316_n
  );


  and

  (
    g2687_p,
    g2330_n_spl_0,
    g2329_n
  );


  or

  (
    g2688_n,
    g2687_p,
    g2686_p
  );


  and

  (
    g2689_p,
    G20_p_spl_10,
    G9_p_spl_1
  );


  and

  (
    g2690_p,
    G19_p_spl_10,
    G4_p_spl_1
  );


  and

  (
    g2691_p,
    g2647_n_spl_,
    g2642_n_spl_
  );


  or

  (
    g2692_n,
    g2607_p_spl_,
    g2519_n
  );


  and

  (
    g2693_p,
    g2550_n_spl_,
    g2549_n_spl_
  );


  or

  (
    g2693_n,
    g2550_p_spl_,
    g2549_p_spl_
  );


  and

  (
    g2694_p,
    g2693_n,
    g2551_n_spl_
  );


  or

  (
    g2694_n,
    g2693_p,
    g2551_p_spl_
  );


  and

  (
    g2695_p,
    g2694_n_spl_,
    g2290_n_spl_0
  );


  or

  (
    g2695_n,
    g2694_p_spl_,
    g2290_p_spl_0
  );


  and

  (
    g2696_p,
    g2695_n_spl_0,
    g2694_n_spl_
  );


  or

  (
    g2696_n,
    g2695_p_spl_,
    g2694_p_spl_
  );


  and

  (
    g2697_p,
    g2695_n_spl_0,
    g2290_n_spl_
  );


  or

  (
    g2697_n,
    g2695_p_spl_,
    g2290_p_spl_
  );


  and

  (
    g2698_p,
    g2697_n,
    g2696_n
  );


  or

  (
    g2698_n,
    g2697_p,
    g2696_p
  );


  and

  (
    g2699_p,
    G19_p_spl_11,
    G6_p_spl_1
  );


  or

  (
    g2699_n,
    G19_n_spl_11,
    G6_n_spl_
  );


  or

  (
    g2700_n,
    g2699_p,
    g2698_p
  );


  and

  (
    g2701_p,
    g2700_n_spl_0,
    g2695_n_spl_
  );


  and

  (
    g2702_p,
    g2585_n_spl_0,
    g2583_n_spl_
  );


  or

  (
    g2702_n,
    g2585_p_spl_0,
    g2583_p_spl_
  );


  and

  (
    g2703_p,
    g2585_n_spl_,
    g2584_n_spl_
  );


  or

  (
    g2703_n,
    g2585_p_spl_,
    g2584_p_spl_
  );


  and

  (
    g2704_p,
    g2703_n,
    g2702_n
  );


  or

  (
    g2704_n,
    g2703_p,
    g2702_p
  );


  and

  (
    g2705_p,
    g2313_n_spl_,
    g2308_n_spl_
  );


  or

  (
    g2705_n,
    g2313_p_spl_,
    g2308_p_spl_
  );


  and

  (
    g2706_p,
    g2705_n_spl_,
    g2704_n_spl_
  );


  or

  (
    g2706_n,
    g2705_p_spl_,
    g2704_p_spl_
  );


  and

  (
    g2707_p,
    g2706_n_spl_0,
    g2704_n_spl_
  );


  or

  (
    g2707_n,
    g2706_p_spl_,
    g2704_p_spl_
  );


  and

  (
    g2708_p,
    g2706_n_spl_0,
    g2705_n_spl_
  );


  or

  (
    g2708_n,
    g2706_p_spl_,
    g2705_p_spl_
  );


  and

  (
    g2709_p,
    g2708_n,
    g2707_n
  );


  or

  (
    g2709_n,
    g2708_p,
    g2707_p
  );


  and

  (
    g2710_p,
    G20_p_spl_10,
    G11_p_spl_1
  );


  or

  (
    g2710_n,
    G20_n_spl_1,
    G11_n_spl_1
  );


  or

  (
    g2711_n,
    g2710_p,
    g2709_p
  );


  and

  (
    g2712_p,
    g2711_n_spl_0,
    g2706_n_spl_
  );


  and

  (
    g2713_p,
    g2711_n_spl_0,
    g2710_n
  );


  and

  (
    g2714_p,
    g2700_n_spl_0,
    g2699_n
  );


  and

  (
    g2715_p,
    g2616_n_spl_0,
    g2615_n
  );


  and

  (
    g2716_p,
    g2629_n_spl_0,
    g2628_n
  );


  and

  (
    g2717_p,
    g2662_n_spl_0,
    g2661_n
  );


  and

  (
    g2718_p,
    g2662_n_spl_0,
    g2650_n
  );


  and

  (
    g2719_p,
    g2616_n_spl_0,
    g2611_n
  );


  and

  (
    g2720_p,
    g2629_n_spl_0,
    g2619_n
  );


  and

  (
    g2721_p,
    g2700_n_spl_,
    g2698_n
  );


  and

  (
    g2722_p,
    g2711_n_spl_,
    g2709_n
  );


  and

  (
    g2723_p,
    g2688_n_spl_,
    g2523_n_spl_
  );


  and

  (
    g2724_p,
    g2685_n_spl_,
    g2524_n_spl_
  );


  and

  (
    g2725_p,
    g2679_n_spl_,
    g2541_n_spl_0
  );


  or

  (
    g2726_n,
    g2682_p_spl_,
    g2558_p_spl_
  );


  or

  (
    g2727_n,
    g2677_p_spl_,
    g2593_p_spl_
  );


  and

  (
    g2728_p,
    g2409_n_spl_0,
    g2407_n
  );


  and

  (
    g2729_p,
    g2409_n_spl_0,
    g2408_n
  );


  or

  (
    g2730_n,
    g2729_p,
    g2728_p
  );


  or

  (
    g2731_n,
    g2540_p_spl_,
    g2539_p
  );


  and

  (
    g2732_p,
    g2731_n,
    g2541_n_spl_0
  );


  and

  (
    g2733_p,
    g2592_n_spl_0,
    g2590_n
  );


  and

  (
    g2734_p,
    g2592_n_spl_,
    g2591_n
  );


  or

  (
    g2735_n,
    g2734_p,
    g2733_p
  );


  and

  (
    g2736_p,
    g2557_n_spl_0,
    g2555_n
  );


  and

  (
    g2737_p,
    g2557_n_spl_,
    g2556_n
  );


  or

  (
    g2738_n,
    g2737_p,
    g2736_p
  );


  and

  (
    g2739_p,
    g2486_n_spl_0,
    g2481_n
  );


  and

  (
    g2740_p,
    g2486_n_spl_0,
    g2485_n_spl_
  );


  or

  (
    g2741_n,
    g2740_p,
    g2739_p
  );


  and

  (
    g2742_p,
    g2503_n_spl_0,
    g2489_n
  );


  and

  (
    g2743_p,
    g2503_n_spl_0,
    g2502_n
  );


  or

  (
    g2744_n,
    g2743_p,
    g2742_p
  );


  buf

  (
    G6257,
    g405_p
  );


  buf

  (
    G6258,
    g408_p
  );


  buf

  (
    G6259,
    g411_p
  );


  buf

  (
    G6260,
    g414_p
  );


  buf

  (
    G6261,
    g417_p
  );


  buf

  (
    G6262,
    g420_p
  );


  buf

  (
    G6263,
    g423_p
  );


  buf

  (
    G6264,
    g426_p
  );


  buf

  (
    G6265,
    g429_p
  );


  buf

  (
    G6266,
    g432_p
  );


  buf

  (
    G6267,
    g435_p
  );


  buf

  (
    G6268,
    g438_p
  );


  buf

  (
    G6269,
    g441_p
  );


  buf

  (
    G6270,
    g444_p
  );


  buf

  (
    G6271,
    g447_p
  );


  buf

  (
    G6272,
    g450_p
  );


  buf

  (
    G6273,
    g452_p
  );


  buf

  (
    G6274,
    g455_p
  );


  buf

  (
    G6275,
    g458_p
  );


  buf

  (
    G6276,
    g464_p
  );


  buf

  (
    G6277,
    g473_p
  );


  buf

  (
    G6278,
    g486_p
  );


  buf

  (
    G6279,
    g502_p
  );


  buf

  (
    G6280,
    g521_p
  );


  buf

  (
    G6281,
    g544_p
  );


  buf

  (
    G6282,
    g570_p
  );


  buf

  (
    G6283,
    g599_p
  );


  buf

  (
    G6284,
    g632_p
  );


  buf

  (
    G6285,
    g663_p
  );


  buf

  (
    G6286,
    g684_p
  );


  buf

  (
    G6287,
    g693_p
  );


  not

  (
    G6288,
    g696_n
  );


  buf

  (
    n2491_li,
    n6461_o2_p_spl_1
  );


  buf

  (
    n2575_li,
    n6042_o2_p_spl_1
  );


  buf

  (
    n2587_li,
    n5981_o2_p_spl_1
  );


  buf

  (
    n2599_li,
    n5959_o2_p_spl_1
  );


  buf

  (
    n2611_li,
    n5930_o2_p_spl_1
  );


  buf

  (
    n2623_li,
    n5881_o2_p_spl_1
  );


  buf

  (
    n2635_li,
    n5863_o2_p_spl_1
  );


  buf

  (
    n2647_li,
    n5842_o2_p_spl_1
  );


  buf

  (
    n2659_li,
    n5792_o2_p_spl_1
  );


  buf

  (
    n2671_li,
    n5779_o2_p_spl_1
  );


  buf

  (
    n2683_li,
    n5780_o2_p
  );


  buf

  (
    n2734_li,
    G22_p
  );


  buf

  (
    n2746_li,
    G23_p
  );


  buf

  (
    n2758_li,
    G24_p
  );


  buf

  (
    n2770_li,
    G25_p
  );


  buf

  (
    n2782_li,
    G26_p
  );


  buf

  (
    n2785_li,
    n2782_lo_p
  );


  buf

  (
    n2794_li,
    G27_p
  );


  buf

  (
    n2797_li,
    n2794_lo_p
  );


  buf

  (
    n2806_li,
    G28_p
  );


  buf

  (
    n2809_li,
    n2806_lo_p
  );


  buf

  (
    n2818_li,
    G29_p
  );


  buf

  (
    n2821_li,
    n2818_lo_p
  );


  buf

  (
    n2830_li,
    G30_p
  );


  buf

  (
    n2833_li,
    n2830_lo_p
  );


  buf

  (
    n2836_li,
    n2833_lo_p
  );


  buf

  (
    n2839_li,
    n2836_lo_p_spl_11
  );


  buf

  (
    n2842_li,
    G31_p
  );


  buf

  (
    n2845_li,
    n2842_lo_p
  );


  buf

  (
    n2848_li,
    n2845_lo_p
  );


  buf

  (
    n2851_li,
    n2848_lo_p_spl_11
  );


  buf

  (
    n2854_li,
    G32_p
  );


  buf

  (
    n2857_li,
    n2854_lo_p
  );


  buf

  (
    n2860_li,
    n2857_lo_p
  );


  buf

  (
    n2863_li,
    n2860_lo_p_spl_1
  );


  buf

  (
    n4871_i2,
    n6476_o2_p
  );


  buf

  (
    n4893_i2,
    n325_inv_p
  );


  buf

  (
    n4938_i2,
    n6545_o2_p
  );


  buf

  (
    n5056_i2,
    n6713_o2_p
  );


  buf

  (
    n5100_i2,
    n343_inv_p
  );


  buf

  (
    n5122_i2,
    n6810_o2_p
  );


  buf

  (
    n5254_i2,
    n6973_o2_p
  );


  buf

  (
    n5276_i2,
    n352_inv_p
  );


  buf

  (
    n5316_i2,
    n7053_o2_p
  );


  buf

  (
    n5434_i2,
    n7231_o2_p
  );


  buf

  (
    n5473_i2,
    n370_inv_p
  );


  buf

  (
    n5494_i2,
    n7304_o2_p
  );


  buf

  (
    n5620_i2,
    n7530_o2_p
  );


  buf

  (
    n5643_i2,
    n379_inv_p
  );


  buf

  (
    n5682_i2,
    n7653_o2_p
  );


  buf

  (
    n5798_i2,
    n7916_o2_p
  );


  buf

  (
    n5839_i2,
    n406_inv_p
  );


  buf

  (
    n5867_i2,
    n8056_o2_p
  );


  buf

  (
    n6052_i2,
    G563_o2_p
  );


  buf

  (
    n6087_i2,
    n439_inv_p
  );


  buf

  (
    n6153_i2,
    G3410_o2_p
  );


  buf

  (
    n6408_i2,
    G566_o2_p
  );


  buf

  (
    n6454_i2,
    n472_inv_p
  );


  buf

  (
    n6509_i2,
    G3752_o2_p
  );


  buf

  (
    n6775_i2,
    G569_o2_p
  );


  buf

  (
    n6818_i2,
    n505_inv_p
  );


  buf

  (
    n6892_i2,
    G4101_o2_p
  );


  buf

  (
    n5779_i2,
    n7148_o2_p_spl_1
  );


  buf

  (
    n5780_i2,
    n7149_o2_p
  );


  buf

  (
    n7156_i2,
    G572_o2_p
  );


  buf

  (
    n5792_i2,
    n7224_o2_p_spl_1
  );


  buf

  (
    n7205_i2,
    n547_inv_p
  );


  buf

  (
    n5842_i2,
    n7280_o2_p_spl_1
  );


  buf

  (
    n5863_i2,
    n7313_o2_p_spl_1
  );


  buf

  (
    n7263_i2,
    G4452_o2_p
  );


  buf

  (
    n5881_i2,
    n7323_o2_p_spl_1
  );


  buf

  (
    n5930_i2,
    n7398_o2_p_spl_1
  );


  buf

  (
    n5959_i2,
    n7459_o2_p_spl_1
  );


  buf

  (
    n5981_i2,
    n7501_o2_p_spl_1
  );


  buf

  (
    n6042_i2,
    n7518_o2_p_spl_1
  );


  buf

  (
    n6075_i2,
    n7606_o2_p_spl_1
  );


  buf

  (
    n6103_i2,
    n7675_o2_p_spl_1
  );


  buf

  (
    n7610_i2,
    G575_o2_p
  );


  buf

  (
    n6169_i2,
    n7722_o2_p_spl_1
  );


  buf

  (
    n7665_i2,
    n649_inv_p
  );


  buf

  (
    n6205_i2,
    n7747_o2_p_spl_1
  );


  buf

  (
    n6239_i2,
    n7835_o2_p_spl_1
  );


  buf

  (
    n7788_i2,
    G4806_o2_p
  );


  buf

  (
    n6309_i2,
    n7909_o2_p_spl_1
  );


  buf

  (
    n6461_i2,
    n8086_o2_p_spl_1
  );


  buf

  (
    n6476_i2,
    n8093_o2_p
  );


  buf

  (
    n6521_i2,
    n484_inv_p
  );


  buf

  (
    n6545_i2,
    n8199_o2_p
  );


  buf

  (
    G578_i2,
    g697_p_spl_
  );


  buf

  (
    G5106_i2,
    g698_n_spl_
  );


  buf

  (
    n6713_i2,
    G548_o2_p
  );


  buf

  (
    G5164_i2,
    g699_p_spl_
  );


  buf

  (
    n6771_i2,
    n496_inv_p
  );


  buf

  (
    n6810_i2,
    G1761_o2_p
  );


  buf

  (
    n6973_i2,
    G551_o2_p
  );


  buf

  (
    n6995_i2,
    n514_inv_p
  );


  buf

  (
    n7053_i2,
    G2082_o2_p
  );


  buf

  (
    G581_i2,
    g700_p_spl_
  );


  buf

  (
    G5467_i2,
    g709_n_spl_
  );


  buf

  (
    n7231_i2,
    G554_o2_p
  );


  buf

  (
    G5527_i2,
    g710_p_spl_
  );


  buf

  (
    n7277_i2,
    n559_inv_p
  );


  buf

  (
    n7304_i2,
    G2410_o2_p
  );


  buf

  (
    n7530_i2,
    G557_o2_p
  );


  buf

  (
    n7595_i2,
    n634_inv_p
  );


  buf

  (
    n7653_i2,
    G2740_o2_p
  );


  buf

  (
    G584_i2,
    g711_p_spl_
  );


  buf

  (
    G5820_i2,
    g729_n_spl_
  );


  buf

  (
    n7148_i2,
    n2668_lo_buf_o2_p_spl_1
  );


  buf

  (
    n7149_i2,
    n2680_lo_buf_o2_p
  );


  buf

  (
    n7224_i2,
    n2656_lo_buf_o2_p_spl_1
  );


  buf

  (
    n7916_i2,
    G560_o2_p
  );


  buf

  (
    G5868_i2,
    g730_p_spl_
  );


  buf

  (
    n7958_i2,
    n748_inv_p
  );


  buf

  (
    n7280_i2,
    n2644_lo_buf_o2_p_spl_1
  );


  buf

  (
    n7313_i2,
    n2632_lo_buf_o2_p_spl_1
  );


  buf

  (
    n8056_i2,
    G3073_o2_p
  );


  buf

  (
    n7323_i2,
    n2620_lo_buf_o2_p_spl_1
  );


  buf

  (
    n7398_i2,
    n2608_lo_buf_o2_p_spl_1
  );


  buf

  (
    n7459_i2,
    n2596_lo_buf_o2_p_spl_1
  );


  buf

  (
    n7501_i2,
    n2584_lo_buf_o2_p_spl_1
  );


  buf

  (
    n7518_i2,
    n2572_lo_buf_o2_p_spl_1
  );


  buf

  (
    G563_i2,
    g731_p_spl_
  );


  buf

  (
    n7606_i2,
    n2560_lo_buf_o2_p_spl_1
  );


  buf

  (
    G3358_i2,
    g734_n_spl_
  );


  buf

  (
    n7675_i2,
    n2548_lo_buf_o2_p_spl_1
  );


  buf

  (
    G3410_i2,
    g735_p_spl_
  );


  buf

  (
    n7722_i2,
    n2536_lo_buf_o2_p_spl_1
  );


  buf

  (
    n7747_i2,
    n2524_lo_buf_o2_p_spl_1
  );


  buf

  (
    n7835_i2,
    n2512_lo_buf_o2_p_spl_1
  );


  buf

  (
    G587_i2,
    g736_p_spl_
  );


  buf

  (
    G6046_i2,
    g762_n_spl_
  );


  buf

  (
    n7909_i2,
    n2500_lo_buf_o2_p_spl_1
  );


  buf

  (
    G566_i2,
    g763_p_spl_
  );


  buf

  (
    G6070_i2,
    g764_p_spl_
  );


  buf

  (
    G3698_i2,
    g775_n_spl_
  );


  buf

  (
    n8086_i2,
    n2488_lo_buf_o2_p_spl_1
  );


  buf

  (
    n8093_i2,
    G545_o2_p
  );


  buf

  (
    G3752_i2,
    g776_p_spl_
  );


  buf

  (
    n8156_i2,
    n979_inv_p
  );


  buf

  (
    n8199_i2,
    G1445_o2_p
  );


  buf

  (
    n2800_lo_buf_i2,
    n2797_lo_p_spl_11
  );


  buf

  (
    G548_i2,
    g777_p_spl_
  );


  buf

  (
    G1715_i2,
    g781_n_spl_
  );


  buf

  (
    G569_i2,
    g782_p_spl_
  );


  buf

  (
    G1761_i2,
    g783_p_spl_
  );


  buf

  (
    G4043_i2,
    g802_n_spl_
  );


  buf

  (
    G4101_i2,
    g803_p_spl_
  );


  buf

  (
    G551_i2,
    g804_p_spl_
  );


  buf

  (
    G2034_i2,
    g817_n_spl_
  );


  buf

  (
    G4743_i2,
    g861_n_spl_
  );


  buf

  (
    G5271_i2,
    g935_n_spl_
  );


  buf

  (
    G5790_i2,
    g1009_n_spl_
  );


  buf

  (
    G6122_i2,
    g1043_n_spl_0
  );


  buf

  (
    G2082_i2,
    g1044_p_spl_
  );


  buf

  (
    n2812_lo_buf_i2,
    n2809_lo_p_spl_11
  );


  buf

  (
    n2668_lo_buf_i2,
    G16_p_spl_1
  );


  buf

  (
    n2680_lo_buf_i2,
    G17_p_spl_111
  );


  buf

  (
    G572_i2,
    g1045_p_spl_
  );


  buf

  (
    G6125_i2,
    g1043_n_spl_
  );


  buf

  (
    G4395_i2,
    g1073_n_spl_
  );


  buf

  (
    n2656_lo_buf_i2,
    G15_p_spl_1
  );


  buf

  (
    G554_i2,
    g1074_p_spl_
  );


  buf

  (
    G4452_i2,
    g1075_p_spl_
  );


  buf

  (
    G2358_i2,
    g1096_n_spl_
  );


  buf

  (
    n2644_lo_buf_i2,
    G14_p_spl_1
  );


  buf

  (
    G2410_i2,
    g1097_p_spl_
  );


  buf

  (
    n2632_lo_buf_i2,
    G13_p_spl_1
  );


  buf

  (
    n2620_lo_buf_i2,
    G12_p_spl_1
  );


  not

  (
    G6131_i2,
    g1098_n_spl_
  );


  buf

  (
    G4693_i2,
    g1101_n_spl_
  );


  buf

  (
    G5209_i2,
    g1126_n_spl_
  );


  buf

  (
    G5741_i2,
    g1151_n_spl_
  );


  buf

  (
    G6082_i2,
    g1206_n_spl_
  );


  buf

  (
    G6119_i2,
    g1214_n_spl_
  );


  buf

  (
    n2608_lo_buf_i2,
    G11_p_spl_1
  );


  buf

  (
    n2596_lo_buf_i2,
    G10_p_spl_1
  );


  buf

  (
    n2584_lo_buf_i2,
    G9_p_spl_1
  );


  buf

  (
    n2572_lo_buf_i2,
    G8_p_spl_1
  );


  buf

  (
    n2704_lo_buf_i2,
    G19_p_spl_11
  );


  buf

  (
    G557_i2,
    g1215_p_spl_
  );


  not

  (
    G5936_i2,
    g1220_n_spl_
  );


  not

  (
    G5442_i2,
    g1225_n_spl_
  );


  not

  (
    G4926_i2,
    g1230_n_spl_
  );


  buf

  (
    G6134_i2,
    g1231_p_spl_
  );


  buf

  (
    G3929_i2,
    g1293_n_spl_
  );


  buf

  (
    G4425_i2,
    g1367_n_spl_
  );


  buf

  (
    G4947_i2,
    g1477_n_spl_
  );


  buf

  (
    n2764_lo_buf_i2,
    n2758_lo_p_spl_11
  );


  buf

  (
    G2689_i2,
    g1506_n_spl_
  );


  buf

  (
    n2560_lo_buf_i2,
    G7_p_spl_1
  );


  buf

  (
    n2824_lo_buf_i2,
    n2821_lo_p_spl_1
  );


  buf

  (
    G575_i2,
    g1507_p_spl_
  );


  buf

  (
    G2740_i2,
    g1508_p_spl_
  );


  buf

  (
    G4749_i2,
    g1544_n_spl_
  );


  buf

  (
    n2548_lo_buf_i2,
    G6_p_spl_1
  );


  buf

  (
    n2536_lo_buf_i2,
    G5_p_spl_
  );


  buf

  (
    n2524_lo_buf_i2,
    G4_p_spl_1
  );


  not

  (
    G875_i2,
    g1545_n_spl_
  );


  not

  (
    G1064_i2,
    g1546_n_spl_
  );


  not

  (
    G1253_i2,
    g1547_n_spl_
  );


  not

  (
    G6140_i2,
    g1548_n_spl_
  );


  buf

  (
    G5151_i2,
    g1563_n_spl_
  );


  buf

  (
    G5686_i2,
    g1578_n_spl_
  );


  buf

  (
    G6061_i2,
    g1593_n_spl_
  );


  buf

  (
    G4803_i2,
    g1596_n_spl_
  );


  buf

  (
    G5332_i2,
    g1599_n_spl_
  );


  buf

  (
    G5844_i2,
    g1602_n_spl_
  );


  buf

  (
    G6114_i2,
    g1605_n_spl_
  );


  buf

  (
    G4806_i2,
    g1606_p_spl_
  );


  buf

  (
    G3881_i2,
    g1619_n_spl_
  );


  buf

  (
    G4370_i2,
    g1644_n_spl_
  );


  buf

  (
    G4896_i2,
    g1669_n_spl_
  );


  buf

  (
    G5001_i2,
    g1724_n_spl_
  );


  buf

  (
    G3121_i2,
    g1801_n_spl_
  );


  buf

  (
    n2512_lo_buf_i2,
    G3_p_spl_
  );


  not

  (
    G4085_i2,
    g1806_n_spl_
  );


  not

  (
    G4605_i2,
    g1811_n_spl_
  );


  not

  (
    G5118_i2,
    g1816_n_spl_
  );


  buf

  (
    G4997_i2,
    g1831_n_spl_
  );


  buf

  (
    n2500_lo_buf_i2,
    G2_p_spl_
  );


  buf

  (
    n2716_lo_buf_i2,
    G20_p_spl_1
  );


  not

  (
    G560_i2,
    g1832_n_spl_
  );


  buf

  (
    G1895_i2,
    g1846_n_spl_
  );


  buf

  (
    G3064_i2,
    g1869_n_spl_
  );


  buf

  (
    G3269_i2,
    g1996_n_spl_
  );


  buf

  (
    G3569_i2,
    g2106_n_spl_
  );


  buf

  (
    G3022_i2,
    g2134_n_spl_
  );


  not

  (
    G1196_i2,
    g2135_n_spl_
  );


  not

  (
    G1007_i2,
    g2136_n_spl_
  );


  not

  (
    G818_i2,
    g2137_n_spl_
  );


  not

  (
    G674_i2,
    g2138_n_spl_
  );


  buf

  (
    G5041_i2,
    g2139_p
  );


  buf

  (
    G5562_i2,
    g2140_p
  );


  buf

  (
    G6005_i2,
    g2141_p
  );


  buf

  (
    G5214_i2,
    g2142_p
  );


  buf

  (
    G5746_i2,
    g2143_p
  );


  buf

  (
    G6087_i2,
    g2144_p
  );


  buf

  (
    G6086_i2,
    g2145_p
  );


  buf

  (
    G5745_i2,
    g2146_p
  );


  buf

  (
    G5213_i2,
    g2147_p
  );


  buf

  (
    G5893_i2,
    g2148_p
  );


  buf

  (
    G5391_i2,
    g2149_p
  );


  buf

  (
    G4864_i2,
    g2150_p
  );


  buf

  (
    G6143_i2,
    g2151_p
  );


  not

  (
    G6008_i2,
    g2154_n
  );


  not

  (
    G5565_i2,
    g2157_n
  );


  not

  (
    G5044_i2,
    g2160_n
  );


  buf

  (
    G3813_i2,
    g2163_n_spl_
  );


  buf

  (
    G4325_i2,
    g2178_n_spl_
  );


  buf

  (
    G4834_i2,
    g2193_n_spl_
  );


  buf

  (
    G4993_i2,
    g2198_n_spl_
  );


  buf

  (
    G3989_i2,
    g2201_n_spl_
  );


  buf

  (
    G4490_i2,
    g2204_n_spl_
  );


  buf

  (
    G5011_i2,
    g2207_n_spl_
  );


  buf

  (
    G5112_i2,
    g2210_n_spl_
  );


  buf

  (
    n2776_lo_buf_i2,
    n2770_lo_p_spl_
  );


  not

  (
    G3298_i2,
    g2215_n_spl_
  );


  buf

  (
    G3073_i2,
    g2216_p_spl_
  );


  buf

  (
    G3265_i2,
    g2241_n_spl_
  );


  buf

  (
    G3624_i2,
    g2286_n_spl_
  );


  buf

  (
    G1642_i2,
    g2297_n_spl_
  );


  buf

  (
    G1980_i2,
    g2330_n_spl_
  );


  buf

  (
    n2488_lo_buf_i2,
    G1_p
  );


  buf

  (
    G626_i2,
    g2331_p
  );


  not

  (
    G1139_i2,
    g2332_n_spl_
  );


  not

  (
    G950_i2,
    g2333_n_spl_
  );


  not

  (
    G707_i2,
    g2334_n_spl_
  );


  not

  (
    G545_i2,
    g2335_n_spl_
  );


  buf

  (
    G4217_i2,
    g2336_p
  );


  buf

  (
    G4716_i2,
    g2337_p
  );


  buf

  (
    G5244_i2,
    g2348_p
  );


  not

  (
    G3136_i2,
    g2349_n_spl_
  );


  buf

  (
    G3499_i2,
    g2390_p_spl_
  );


  buf

  (
    G3885_i2,
    g2391_p
  );


  not

  (
    G5243_i2,
    g2392_p
  );


  buf

  (
    G3886_i2,
    g2393_p
  );


  buf

  (
    G4375_i2,
    g2394_p
  );


  buf

  (
    G4901_i2,
    g2395_p
  );


  buf

  (
    G5054_i2,
    g2396_p
  );


  buf

  (
    G4374_i2,
    g2397_p
  );


  buf

  (
    G4900_i2,
    g2398_p
  );


  buf

  (
    G5053_i2,
    g2399_p
  );


  buf

  (
    G5242_i2,
    g2400_p
  );


  buf

  (
    G4034_i2,
    g2401_p
  );


  buf

  (
    G4556_i2,
    g2402_p
  );


  buf

  (
    G5064_i2,
    g2403_p
  );


  buf

  (
    G5172_i2,
    g2404_p
  );


  not

  (
    G2030_i2,
    g2409_n_spl_
  );


  buf

  (
    G3016_i2,
    g2422_n_spl_
  );


  buf

  (
    G3520_i2,
    g2437_n_spl_
  );


  buf

  (
    G3261_i2,
    g2452_n_spl_
  );


  buf

  (
    G3620_i2,
    g2467_n_spl_
  );


  not

  (
    G4220_i2,
    g2470_n
  );


  not

  (
    G4719_i2,
    g2473_n
  );


  not

  (
    G5247_i2,
    g2476_n
  );


  buf

  (
    G5109_i2,
    g2479_n
  );


  buf

  (
    G1638_i2,
    g2486_n_spl_
  );


  buf

  (
    G1976_i2,
    g2503_n_spl_
  );


  buf

  (
    G3560_i2,
    g2506_p_spl_
  );


  not

  (
    G3205_i2,
    g2509_n_spl_
  );


  buf

  (
    G3193_i2,
    g2512_n_spl_
  );


  buf

  (
    G3367_i2,
    g2515_n_spl_
  );


  buf

  (
    G3670_i2,
    g2518_n_spl_
  );


  buf

  (
    G1400_i2,
    g2519_p_spl_
  );


  buf

  (
    G1280_i2,
    g2520_p
  );


  buf

  (
    G902_i2,
    g2521_p
  );


  buf

  (
    G659_i2,
    g2522_p
  );


  not

  (
    G983_i2,
    g2523_n_spl_
  );


  not

  (
    G740_i2,
    g2524_n_spl_
  );


  buf

  (
    G2917_i2,
    g2525_p
  );


  buf

  (
    G3391_i2,
    g2526_p
  );


  buf

  (
    G3494_i2,
    g2537_p
  );


  not

  (
    G1512_i2,
    g2541_n_spl_
  );


  buf

  (
    G1854_i2,
    g2558_p_spl_
  );


  buf

  (
    G2203_i2,
    g2593_p_spl_
  );


  not

  (
    G3493_i2,
    g2594_p
  );


  buf

  (
    G3069_i2,
    g2595_p
  );


  buf

  (
    G3574_i2,
    g2596_p
  );


  buf

  (
    G3319_i2,
    g2597_p
  );


  buf

  (
    G3667_i2,
    g2598_p
  );


  buf

  (
    G3068_i2,
    g2599_p
  );


  buf

  (
    G3573_i2,
    g2600_p
  );


  buf

  (
    G3666_i2,
    g2601_p
  );


  buf

  (
    G3318_i2,
    g2602_p
  );


  buf

  (
    G3492_i2,
    g2603_p
  );


  buf

  (
    G3241_i2,
    g2604_p
  );


  buf

  (
    G3722_i2,
    g2605_p
  );


  buf

  (
    G3422_i2,
    g2606_p
  );


  buf

  (
    G1445_i2,
    g2607_p_spl_
  );


  not

  (
    G3257_i2,
    g2608_p
  );


  buf

  (
    G3616_i2,
    g2609_n
  );


  buf

  (
    G1634_i2,
    g2616_n_spl_
  );


  buf

  (
    G1972_i2,
    g2629_n_spl_
  );


  buf

  (
    G2256_i2,
    g2662_n_spl_
  );


  not

  (
    G3394_i2,
    g2665_n
  );


  not

  (
    G3557_i2,
    g2668_n
  );


  buf

  (
    G3364_i2,
    g2671_n
  );


  buf

  (
    G3719_i2,
    g2674_n
  );


  buf

  (
    G2253_i2,
    g2677_p_spl_
  );


  not

  (
    G1583_i2,
    g2679_n_spl_
  );


  buf

  (
    G1917_i2,
    g2682_p_spl_
  );


  buf

  (
    G1727_i2,
    g2685_n_spl_
  );


  buf

  (
    G2061_i2,
    g2688_n_spl_
  );


  buf

  (
    G935_i2,
    g2689_p
  );


  buf

  (
    G692_i2,
    g2690_p
  );


  buf

  (
    G2136_i2,
    g2691_p
  );


  not

  (
    G1507_i2,
    g2692_n
  );


  buf

  (
    G1849_i2,
    g2701_p
  );


  buf

  (
    G2198_i2,
    g2712_p
  );


  not

  (
    G2197_i2,
    g2713_p
  );


  not

  (
    G1848_i2,
    g2714_p
  );


  buf

  (
    G1689_i2,
    g2715_p
  );


  buf

  (
    G2016_i2,
    g2716_p
  );


  buf

  (
    G2314_i2,
    g2717_p
  );


  buf

  (
    G2313_i2,
    g2718_p
  );


  buf

  (
    G1688_i2,
    g2719_p
  );


  buf

  (
    G2015_i2,
    g2720_p
  );


  buf

  (
    G1847_i2,
    g2721_p
  );


  buf

  (
    G2196_i2,
    g2722_p
  );


  buf

  (
    G2118_i2,
    g2723_p
  );


  buf

  (
    G1777_i2,
    g2724_p
  );


  not

  (
    G1630_i2,
    g2725_p
  );


  buf

  (
    G1968_i2,
    g2726_n
  );


  buf

  (
    G2309_i2,
    g2727_n
  );


  not

  (
    G2139_i2,
    g2730_n
  );


  buf

  (
    G1580_i2,
    g2732_p
  );


  not

  (
    G2250_i2,
    g2735_n
  );


  not

  (
    G1914_i2,
    g2738_n
  );


  buf

  (
    G1724_i2,
    g2741_n
  );


  buf

  (
    G2058_i2,
    g2744_n
  );


  buf

  (
    n2728_lo_buf_i2,
    G21_p
  );


  buf

  (
    n4938_o2_p_spl_,
    n4938_o2_p
  );


  buf

  (
    n5122_o2_p_spl_,
    n5122_o2_p
  );


  buf

  (
    n5316_o2_p_spl_,
    n5316_o2_p
  );


  buf

  (
    n5494_o2_p_spl_,
    n5494_o2_p
  );


  buf

  (
    n5682_o2_p_spl_,
    n5682_o2_p
  );


  buf

  (
    n5867_o2_p_spl_,
    n5867_o2_p
  );


  buf

  (
    n6153_o2_p_spl_,
    n6153_o2_p
  );


  buf

  (
    n6509_o2_p_spl_,
    n6509_o2_p
  );


  buf

  (
    n6892_o2_p_spl_,
    n6892_o2_p
  );


  buf

  (
    n7263_o2_p_spl_,
    n7263_o2_p
  );


  buf

  (
    n7788_o2_p_spl_,
    n7788_o2_p
  );


  buf

  (
    G5164_o2_p_spl_,
    G5164_o2_p
  );


  buf

  (
    G5527_o2_p_spl_,
    G5527_o2_p
  );


  buf

  (
    G5868_o2_p_spl_,
    G5868_o2_p
  );


  buf

  (
    G6070_o2_p_spl_,
    G6070_o2_p
  );


  buf

  (
    G6125_o2_p_spl_,
    G6125_o2_p
  );


  buf

  (
    G6134_o2_p_spl_,
    G6134_o2_p
  );


  buf

  (
    G6143_o2_p_spl_,
    G6143_o2_p
  );


  buf

  (
    G6143_o2_p_spl_0,
    G6143_o2_p_spl_
  );


  buf

  (
    g460_p_spl_,
    g460_p
  );


  buf

  (
    g459_p_spl_,
    g459_p
  );


  buf

  (
    g461_p_spl_,
    g461_p
  );


  buf

  (
    g461_p_spl_0,
    g461_p_spl_
  );


  buf

  (
    G6008_o2_n_spl_,
    G6008_o2_n
  );


  buf

  (
    G6005_o2_n_spl_,
    G6005_o2_n
  );


  buf

  (
    G6008_o2_p_spl_,
    G6008_o2_p
  );


  buf

  (
    G6005_o2_p_spl_,
    G6005_o2_p
  );


  buf

  (
    g465_n_spl_,
    g465_n
  );


  buf

  (
    g465_n_spl_0,
    g465_n_spl_
  );


  buf

  (
    g465_p_spl_,
    g465_p
  );


  buf

  (
    g465_p_spl_0,
    g465_p_spl_
  );


  buf

  (
    g469_p_spl_,
    g469_p
  );


  buf

  (
    g468_p_spl_,
    g468_p
  );


  buf

  (
    g470_p_spl_,
    g470_p
  );


  buf

  (
    g470_p_spl_0,
    g470_p_spl_
  );


  buf

  (
    G5893_o2_n_spl_,
    G5893_o2_n
  );


  buf

  (
    G5893_o2_n_spl_0,
    G5893_o2_n_spl_
  );


  buf

  (
    G5893_o2_p_spl_,
    G5893_o2_p
  );


  buf

  (
    G5893_o2_p_spl_0,
    G5893_o2_p_spl_
  );


  buf

  (
    g477_n_spl_,
    g477_n
  );


  buf

  (
    g476_n_spl_,
    g476_n
  );


  buf

  (
    g477_p_spl_,
    g477_p
  );


  buf

  (
    g476_p_spl_,
    g476_p
  );


  buf

  (
    g478_n_spl_,
    g478_n
  );


  buf

  (
    g478_n_spl_0,
    g478_n_spl_
  );


  buf

  (
    g478_p_spl_,
    g478_p
  );


  buf

  (
    g478_p_spl_0,
    g478_p_spl_
  );


  buf

  (
    g482_p_spl_,
    g482_p
  );


  buf

  (
    g481_p_spl_,
    g481_p
  );


  buf

  (
    g483_p_spl_,
    g483_p
  );


  buf

  (
    g483_p_spl_0,
    g483_p_spl_
  );


  buf

  (
    n2863_lo_p_spl_,
    n2863_lo_p
  );


  buf

  (
    n2863_lo_p_spl_0,
    n2863_lo_p_spl_
  );


  buf

  (
    n2863_lo_p_spl_00,
    n2863_lo_p_spl_0
  );


  buf

  (
    n2863_lo_p_spl_000,
    n2863_lo_p_spl_00
  );


  buf

  (
    n2863_lo_p_spl_01,
    n2863_lo_p_spl_0
  );


  buf

  (
    n2863_lo_p_spl_1,
    n2863_lo_p_spl_
  );


  buf

  (
    n2863_lo_p_spl_10,
    n2863_lo_p_spl_1
  );


  buf

  (
    n2863_lo_p_spl_11,
    n2863_lo_p_spl_1
  );


  buf

  (
    n2863_lo_n_spl_,
    n2863_lo_n
  );


  buf

  (
    n2863_lo_n_spl_0,
    n2863_lo_n_spl_
  );


  buf

  (
    n2863_lo_n_spl_00,
    n2863_lo_n_spl_0
  );


  buf

  (
    n2863_lo_n_spl_000,
    n2863_lo_n_spl_00
  );


  buf

  (
    n2863_lo_n_spl_01,
    n2863_lo_n_spl_0
  );


  buf

  (
    n2863_lo_n_spl_1,
    n2863_lo_n_spl_
  );


  buf

  (
    n2863_lo_n_spl_10,
    n2863_lo_n_spl_1
  );


  buf

  (
    n2863_lo_n_spl_11,
    n2863_lo_n_spl_1
  );


  buf

  (
    g488_n_spl_,
    g488_n
  );


  buf

  (
    g487_n_spl_,
    g487_n
  );


  buf

  (
    g488_p_spl_,
    g488_p
  );


  buf

  (
    g487_p_spl_,
    g487_p
  );


  buf

  (
    g489_n_spl_,
    g489_n
  );


  buf

  (
    g489_n_spl_0,
    g489_n_spl_
  );


  buf

  (
    g489_p_spl_,
    g489_p
  );


  buf

  (
    g489_p_spl_0,
    g489_p_spl_
  );


  buf

  (
    g493_n_spl_,
    g493_n
  );


  buf

  (
    g492_n_spl_,
    g492_n
  );


  buf

  (
    g493_p_spl_,
    g493_p
  );


  buf

  (
    g492_p_spl_,
    g492_p
  );


  buf

  (
    g494_n_spl_,
    g494_n
  );


  buf

  (
    g494_n_spl_0,
    g494_n_spl_
  );


  buf

  (
    g494_p_spl_,
    g494_p
  );


  buf

  (
    g494_p_spl_0,
    g494_p_spl_
  );


  buf

  (
    g498_p_spl_,
    g498_p
  );


  buf

  (
    g497_p_spl_,
    g497_p
  );


  buf

  (
    g499_p_spl_,
    g499_p
  );


  buf

  (
    g499_p_spl_0,
    g499_p_spl_
  );


  buf

  (
    G5565_o2_n_spl_,
    G5565_o2_n
  );


  buf

  (
    G5562_o2_n_spl_,
    G5562_o2_n
  );


  buf

  (
    G5565_o2_p_spl_,
    G5565_o2_p
  );


  buf

  (
    G5562_o2_p_spl_,
    G5562_o2_p
  );


  buf

  (
    g503_n_spl_,
    g503_n
  );


  buf

  (
    g503_n_spl_0,
    g503_n_spl_
  );


  buf

  (
    g503_p_spl_,
    g503_p
  );


  buf

  (
    g503_p_spl_0,
    g503_p_spl_
  );


  buf

  (
    g507_n_spl_,
    g507_n
  );


  buf

  (
    g506_n_spl_,
    g506_n
  );


  buf

  (
    g507_p_spl_,
    g507_p
  );


  buf

  (
    g506_p_spl_,
    g506_p
  );


  buf

  (
    g508_n_spl_,
    g508_n
  );


  buf

  (
    g508_n_spl_0,
    g508_n_spl_
  );


  buf

  (
    g508_p_spl_,
    g508_p
  );


  buf

  (
    g508_p_spl_0,
    g508_p_spl_
  );


  buf

  (
    g512_n_spl_,
    g512_n
  );


  buf

  (
    g511_n_spl_,
    g511_n
  );


  buf

  (
    g512_p_spl_,
    g512_p
  );


  buf

  (
    g511_p_spl_,
    g511_p
  );


  buf

  (
    g513_n_spl_,
    g513_n
  );


  buf

  (
    g513_n_spl_0,
    g513_n_spl_
  );


  buf

  (
    g513_p_spl_,
    g513_p
  );


  buf

  (
    g513_p_spl_0,
    g513_p_spl_
  );


  buf

  (
    g517_p_spl_,
    g517_p
  );


  buf

  (
    g516_p_spl_,
    g516_p
  );


  buf

  (
    g518_p_spl_,
    g518_p
  );


  buf

  (
    g518_p_spl_0,
    g518_p_spl_
  );


  buf

  (
    G5391_o2_n_spl_,
    G5391_o2_n
  );


  buf

  (
    G5391_o2_n_spl_0,
    G5391_o2_n_spl_
  );


  buf

  (
    G5391_o2_p_spl_,
    G5391_o2_p
  );


  buf

  (
    G5391_o2_p_spl_0,
    G5391_o2_p_spl_
  );


  buf

  (
    g525_n_spl_,
    g525_n
  );


  buf

  (
    g524_n_spl_,
    g524_n
  );


  buf

  (
    g525_p_spl_,
    g525_p
  );


  buf

  (
    g524_p_spl_,
    g524_p
  );


  buf

  (
    g526_n_spl_,
    g526_n
  );


  buf

  (
    g526_n_spl_0,
    g526_n_spl_
  );


  buf

  (
    g526_p_spl_,
    g526_p
  );


  buf

  (
    g526_p_spl_0,
    g526_p_spl_
  );


  buf

  (
    g530_n_spl_,
    g530_n
  );


  buf

  (
    g529_n_spl_,
    g529_n
  );


  buf

  (
    g530_p_spl_,
    g530_p
  );


  buf

  (
    g529_p_spl_,
    g529_p
  );


  buf

  (
    g531_n_spl_,
    g531_n
  );


  buf

  (
    g531_n_spl_0,
    g531_n_spl_
  );


  buf

  (
    g531_p_spl_,
    g531_p
  );


  buf

  (
    g531_p_spl_0,
    g531_p_spl_
  );


  buf

  (
    g535_n_spl_,
    g535_n
  );


  buf

  (
    g534_n_spl_,
    g534_n
  );


  buf

  (
    g535_p_spl_,
    g535_p
  );


  buf

  (
    g534_p_spl_,
    g534_p
  );


  buf

  (
    g536_n_spl_,
    g536_n
  );


  buf

  (
    g536_n_spl_0,
    g536_n_spl_
  );


  buf

  (
    g536_p_spl_,
    g536_p
  );


  buf

  (
    g536_p_spl_0,
    g536_p_spl_
  );


  buf

  (
    g540_p_spl_,
    g540_p
  );


  buf

  (
    g539_p_spl_,
    g539_p
  );


  buf

  (
    g541_p_spl_,
    g541_p
  );


  buf

  (
    g541_p_spl_0,
    g541_p_spl_
  );


  buf

  (
    n2851_lo_p_spl_,
    n2851_lo_p
  );


  buf

  (
    n2851_lo_p_spl_0,
    n2851_lo_p_spl_
  );


  buf

  (
    n2851_lo_p_spl_00,
    n2851_lo_p_spl_0
  );


  buf

  (
    n2851_lo_p_spl_1,
    n2851_lo_p_spl_
  );


  buf

  (
    n2623_lo_p_spl_,
    n2623_lo_p
  );


  buf

  (
    n2851_lo_n_spl_,
    n2851_lo_n
  );


  buf

  (
    n2851_lo_n_spl_0,
    n2851_lo_n_spl_
  );


  buf

  (
    n2851_lo_n_spl_00,
    n2851_lo_n_spl_0
  );


  buf

  (
    n2851_lo_n_spl_1,
    n2851_lo_n_spl_
  );


  buf

  (
    n2623_lo_n_spl_,
    n2623_lo_n
  );


  buf

  (
    g546_n_spl_,
    g546_n
  );


  buf

  (
    g545_n_spl_,
    g545_n
  );


  buf

  (
    g546_p_spl_,
    g546_p
  );


  buf

  (
    g545_p_spl_,
    g545_p
  );


  buf

  (
    g547_n_spl_,
    g547_n
  );


  buf

  (
    g547_n_spl_0,
    g547_n_spl_
  );


  buf

  (
    g547_p_spl_,
    g547_p
  );


  buf

  (
    g547_p_spl_0,
    g547_p_spl_
  );


  buf

  (
    g551_n_spl_,
    g551_n
  );


  buf

  (
    g550_n_spl_,
    g550_n
  );


  buf

  (
    g551_p_spl_,
    g551_p
  );


  buf

  (
    g550_p_spl_,
    g550_p
  );


  buf

  (
    g552_n_spl_,
    g552_n
  );


  buf

  (
    g552_n_spl_0,
    g552_n_spl_
  );


  buf

  (
    g552_p_spl_,
    g552_p
  );


  buf

  (
    g552_p_spl_0,
    g552_p_spl_
  );


  buf

  (
    g556_n_spl_,
    g556_n
  );


  buf

  (
    g555_n_spl_,
    g555_n
  );


  buf

  (
    g556_p_spl_,
    g556_p
  );


  buf

  (
    g555_p_spl_,
    g555_p
  );


  buf

  (
    g557_n_spl_,
    g557_n
  );


  buf

  (
    g557_n_spl_0,
    g557_n_spl_
  );


  buf

  (
    g557_p_spl_,
    g557_p
  );


  buf

  (
    g557_p_spl_0,
    g557_p_spl_
  );


  buf

  (
    g561_n_spl_,
    g561_n
  );


  buf

  (
    g560_n_spl_,
    g560_n
  );


  buf

  (
    g561_p_spl_,
    g561_p
  );


  buf

  (
    g560_p_spl_,
    g560_p
  );


  buf

  (
    g562_n_spl_,
    g562_n
  );


  buf

  (
    g562_n_spl_0,
    g562_n_spl_
  );


  buf

  (
    g562_p_spl_,
    g562_p
  );


  buf

  (
    g562_p_spl_0,
    g562_p_spl_
  );


  buf

  (
    g566_p_spl_,
    g566_p
  );


  buf

  (
    g565_p_spl_,
    g565_p
  );


  buf

  (
    g567_p_spl_,
    g567_p
  );


  buf

  (
    g567_p_spl_0,
    g567_p_spl_
  );


  buf

  (
    G5044_o2_n_spl_,
    G5044_o2_n
  );


  buf

  (
    G5041_o2_n_spl_,
    G5041_o2_n
  );


  buf

  (
    G5044_o2_p_spl_,
    G5044_o2_p
  );


  buf

  (
    G5041_o2_p_spl_,
    G5041_o2_p
  );


  buf

  (
    g571_n_spl_,
    g571_n
  );


  buf

  (
    g571_n_spl_0,
    g571_n_spl_
  );


  buf

  (
    g571_p_spl_,
    g571_p
  );


  buf

  (
    g571_p_spl_0,
    g571_p_spl_
  );


  buf

  (
    n2635_lo_p_spl_,
    n2635_lo_p
  );


  buf

  (
    n2635_lo_n_spl_,
    n2635_lo_n
  );


  buf

  (
    g575_n_spl_,
    g575_n
  );


  buf

  (
    g574_n_spl_,
    g574_n
  );


  buf

  (
    g575_p_spl_,
    g575_p
  );


  buf

  (
    g574_p_spl_,
    g574_p
  );


  buf

  (
    g576_n_spl_,
    g576_n
  );


  buf

  (
    g576_n_spl_0,
    g576_n_spl_
  );


  buf

  (
    g576_p_spl_,
    g576_p
  );


  buf

  (
    g576_p_spl_0,
    g576_p_spl_
  );


  buf

  (
    g580_n_spl_,
    g580_n
  );


  buf

  (
    g579_n_spl_,
    g579_n
  );


  buf

  (
    g580_p_spl_,
    g580_p
  );


  buf

  (
    g579_p_spl_,
    g579_p
  );


  buf

  (
    g581_n_spl_,
    g581_n
  );


  buf

  (
    g581_n_spl_0,
    g581_n_spl_
  );


  buf

  (
    g581_p_spl_,
    g581_p
  );


  buf

  (
    g581_p_spl_0,
    g581_p_spl_
  );


  buf

  (
    g585_n_spl_,
    g585_n
  );


  buf

  (
    g584_n_spl_,
    g584_n
  );


  buf

  (
    g585_p_spl_,
    g585_p
  );


  buf

  (
    g584_p_spl_,
    g584_p
  );


  buf

  (
    g586_n_spl_,
    g586_n
  );


  buf

  (
    g586_n_spl_0,
    g586_n_spl_
  );


  buf

  (
    g586_p_spl_,
    g586_p
  );


  buf

  (
    g586_p_spl_0,
    g586_p_spl_
  );


  buf

  (
    g590_n_spl_,
    g590_n
  );


  buf

  (
    g589_n_spl_,
    g589_n
  );


  buf

  (
    g590_p_spl_,
    g590_p
  );


  buf

  (
    g589_p_spl_,
    g589_p
  );


  buf

  (
    g591_n_spl_,
    g591_n
  );


  buf

  (
    g591_n_spl_0,
    g591_n_spl_
  );


  buf

  (
    g591_p_spl_,
    g591_p
  );


  buf

  (
    g591_p_spl_0,
    g591_p_spl_
  );


  buf

  (
    g595_p_spl_,
    g595_p
  );


  buf

  (
    g594_p_spl_,
    g594_p
  );


  buf

  (
    g596_p_spl_,
    g596_p
  );


  buf

  (
    g596_p_spl_0,
    g596_p_spl_
  );


  buf

  (
    G4864_o2_n_spl_,
    G4864_o2_n
  );


  buf

  (
    G4864_o2_n_spl_0,
    G4864_o2_n_spl_
  );


  buf

  (
    G4864_o2_p_spl_,
    G4864_o2_p
  );


  buf

  (
    G4864_o2_p_spl_0,
    G4864_o2_p_spl_
  );


  buf

  (
    g603_n_spl_,
    g603_n
  );


  buf

  (
    g602_n_spl_,
    g602_n
  );


  buf

  (
    g603_p_spl_,
    g603_p
  );


  buf

  (
    g602_p_spl_,
    g602_p
  );


  buf

  (
    g604_n_spl_,
    g604_n
  );


  buf

  (
    g604_n_spl_0,
    g604_n_spl_
  );


  buf

  (
    g604_p_spl_,
    g604_p
  );


  buf

  (
    g604_p_spl_0,
    g604_p_spl_
  );


  buf

  (
    n2647_lo_p_spl_,
    n2647_lo_p
  );


  buf

  (
    n2647_lo_n_spl_,
    n2647_lo_n
  );


  buf

  (
    g608_n_spl_,
    g608_n
  );


  buf

  (
    g607_n_spl_,
    g607_n
  );


  buf

  (
    g608_p_spl_,
    g608_p
  );


  buf

  (
    g607_p_spl_,
    g607_p
  );


  buf

  (
    g609_n_spl_,
    g609_n
  );


  buf

  (
    g609_n_spl_0,
    g609_n_spl_
  );


  buf

  (
    g609_p_spl_,
    g609_p
  );


  buf

  (
    g609_p_spl_0,
    g609_p_spl_
  );


  buf

  (
    g613_n_spl_,
    g613_n
  );


  buf

  (
    g612_n_spl_,
    g612_n
  );


  buf

  (
    g613_p_spl_,
    g613_p
  );


  buf

  (
    g612_p_spl_,
    g612_p
  );


  buf

  (
    g614_n_spl_,
    g614_n
  );


  buf

  (
    g614_n_spl_0,
    g614_n_spl_
  );


  buf

  (
    g614_p_spl_,
    g614_p
  );


  buf

  (
    g614_p_spl_0,
    g614_p_spl_
  );


  buf

  (
    g618_n_spl_,
    g618_n
  );


  buf

  (
    g617_n_spl_,
    g617_n
  );


  buf

  (
    g618_p_spl_,
    g618_p
  );


  buf

  (
    g617_p_spl_,
    g617_p
  );


  buf

  (
    g619_n_spl_,
    g619_n
  );


  buf

  (
    g619_n_spl_0,
    g619_n_spl_
  );


  buf

  (
    g619_p_spl_,
    g619_p
  );


  buf

  (
    g619_p_spl_0,
    g619_p_spl_
  );


  buf

  (
    g623_n_spl_,
    g623_n
  );


  buf

  (
    g622_n_spl_,
    g622_n
  );


  buf

  (
    g623_p_spl_,
    g623_p
  );


  buf

  (
    g622_p_spl_,
    g622_p
  );


  buf

  (
    g624_n_spl_,
    g624_n
  );


  buf

  (
    g624_n_spl_0,
    g624_n_spl_
  );


  buf

  (
    g624_p_spl_,
    g624_p
  );


  buf

  (
    g624_p_spl_0,
    g624_p_spl_
  );


  buf

  (
    g628_p_spl_,
    g628_p
  );


  buf

  (
    g627_p_spl_,
    g627_p
  );


  buf

  (
    g629_p_spl_,
    g629_p
  );


  buf

  (
    g629_p_spl_0,
    g629_p_spl_
  );


  buf

  (
    n2671_lo_p_spl_,
    n2671_lo_p
  );


  buf

  (
    n2671_lo_p_spl_0,
    n2671_lo_p_spl_
  );


  buf

  (
    n2671_lo_n_spl_,
    n2671_lo_n
  );


  buf

  (
    n2671_lo_n_spl_0,
    n2671_lo_n_spl_
  );


  buf

  (
    g634_n_spl_,
    g634_n
  );


  buf

  (
    g633_n_spl_,
    g633_n
  );


  buf

  (
    g634_p_spl_,
    g634_p
  );


  buf

  (
    g633_p_spl_,
    g633_p
  );


  buf

  (
    g635_n_spl_,
    g635_n
  );


  buf

  (
    g635_n_spl_0,
    g635_n_spl_
  );


  buf

  (
    g635_p_spl_,
    g635_p
  );


  buf

  (
    g635_p_spl_0,
    g635_p_spl_
  );


  buf

  (
    n2659_lo_p_spl_,
    n2659_lo_p
  );


  buf

  (
    n2659_lo_n_spl_,
    n2659_lo_n
  );


  buf

  (
    g639_n_spl_,
    g639_n
  );


  buf

  (
    g638_n_spl_,
    g638_n
  );


  buf

  (
    g639_p_spl_,
    g639_p
  );


  buf

  (
    g638_p_spl_,
    g638_p
  );


  buf

  (
    g640_n_spl_,
    g640_n
  );


  buf

  (
    g640_n_spl_0,
    g640_n_spl_
  );


  buf

  (
    g640_p_spl_,
    g640_p
  );


  buf

  (
    g640_p_spl_0,
    g640_p_spl_
  );


  buf

  (
    g644_n_spl_,
    g644_n
  );


  buf

  (
    g643_n_spl_,
    g643_n
  );


  buf

  (
    g644_p_spl_,
    g644_p
  );


  buf

  (
    g643_p_spl_,
    g643_p
  );


  buf

  (
    g645_n_spl_,
    g645_n
  );


  buf

  (
    g645_n_spl_0,
    g645_n_spl_
  );


  buf

  (
    g645_p_spl_,
    g645_p
  );


  buf

  (
    g645_p_spl_0,
    g645_p_spl_
  );


  buf

  (
    g649_n_spl_,
    g649_n
  );


  buf

  (
    g648_n_spl_,
    g648_n
  );


  buf

  (
    g649_p_spl_,
    g649_p
  );


  buf

  (
    g648_p_spl_,
    g648_p
  );


  buf

  (
    g650_n_spl_,
    g650_n
  );


  buf

  (
    g650_n_spl_0,
    g650_n_spl_
  );


  buf

  (
    g650_p_spl_,
    g650_p
  );


  buf

  (
    g650_p_spl_0,
    g650_p_spl_
  );


  buf

  (
    g654_n_spl_,
    g654_n
  );


  buf

  (
    g653_n_spl_,
    g653_n
  );


  buf

  (
    g654_p_spl_,
    g654_p
  );


  buf

  (
    g653_p_spl_,
    g653_p
  );


  buf

  (
    g655_n_spl_,
    g655_n
  );


  buf

  (
    g655_n_spl_0,
    g655_n_spl_
  );


  buf

  (
    g655_p_spl_,
    g655_p
  );


  buf

  (
    g655_p_spl_0,
    g655_p_spl_
  );


  buf

  (
    g659_p_spl_,
    g659_p
  );


  buf

  (
    g658_p_spl_,
    g658_p
  );


  buf

  (
    g660_p_spl_,
    g660_p
  );


  buf

  (
    g660_p_spl_0,
    g660_p_spl_
  );


  buf

  (
    g665_n_spl_,
    g665_n
  );


  buf

  (
    g664_n_spl_,
    g664_n
  );


  buf

  (
    g665_p_spl_,
    g665_p
  );


  buf

  (
    g664_p_spl_,
    g664_p
  );


  buf

  (
    g666_n_spl_,
    g666_n
  );


  buf

  (
    g666_n_spl_0,
    g666_n_spl_
  );


  buf

  (
    g666_p_spl_,
    g666_p
  );


  buf

  (
    g666_p_spl_0,
    g666_p_spl_
  );


  buf

  (
    g670_n_spl_,
    g670_n
  );


  buf

  (
    g669_n_spl_,
    g669_n
  );


  buf

  (
    g670_p_spl_,
    g670_p
  );


  buf

  (
    g669_p_spl_,
    g669_p
  );


  buf

  (
    g671_n_spl_,
    g671_n
  );


  buf

  (
    g671_n_spl_0,
    g671_n_spl_
  );


  buf

  (
    g671_p_spl_,
    g671_p
  );


  buf

  (
    g671_p_spl_0,
    g671_p_spl_
  );


  buf

  (
    g675_n_spl_,
    g675_n
  );


  buf

  (
    g674_n_spl_,
    g674_n
  );


  buf

  (
    g675_p_spl_,
    g675_p
  );


  buf

  (
    g674_p_spl_,
    g674_p
  );


  buf

  (
    g676_n_spl_,
    g676_n
  );


  buf

  (
    g676_n_spl_0,
    g676_n_spl_
  );


  buf

  (
    g676_p_spl_,
    g676_p
  );


  buf

  (
    g676_p_spl_0,
    g676_p_spl_
  );


  buf

  (
    g680_p_spl_,
    g680_p
  );


  buf

  (
    g679_p_spl_,
    g679_p
  );


  buf

  (
    g681_p_spl_,
    g681_p
  );


  buf

  (
    g681_p_spl_0,
    g681_p_spl_
  );


  buf

  (
    g686_n_spl_,
    g686_n
  );


  buf

  (
    g685_n_spl_,
    g685_n
  );


  buf

  (
    g686_p_spl_,
    g686_p
  );


  buf

  (
    g685_p_spl_,
    g685_p
  );


  buf

  (
    g687_n_spl_,
    g687_n
  );


  buf

  (
    g687_n_spl_0,
    g687_n_spl_
  );


  buf

  (
    g687_p_spl_,
    g687_p
  );


  buf

  (
    g692_n_spl_,
    g692_n
  );


  buf

  (
    g692_n_spl_0,
    g692_n_spl_
  );


  buf

  (
    n2824_lo_buf_o2_p_spl_,
    n2824_lo_buf_o2_p
  );


  buf

  (
    n2824_lo_buf_o2_p_spl_0,
    n2824_lo_buf_o2_p_spl_
  );


  buf

  (
    n2824_lo_buf_o2_p_spl_00,
    n2824_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2824_lo_buf_o2_p_spl_000,
    n2824_lo_buf_o2_p_spl_00
  );


  buf

  (
    n2824_lo_buf_o2_p_spl_001,
    n2824_lo_buf_o2_p_spl_00
  );


  buf

  (
    n2824_lo_buf_o2_p_spl_01,
    n2824_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2824_lo_buf_o2_p_spl_010,
    n2824_lo_buf_o2_p_spl_01
  );


  buf

  (
    n2824_lo_buf_o2_p_spl_1,
    n2824_lo_buf_o2_p_spl_
  );


  buf

  (
    n2824_lo_buf_o2_p_spl_10,
    n2824_lo_buf_o2_p_spl_1
  );


  buf

  (
    n2824_lo_buf_o2_p_spl_11,
    n2824_lo_buf_o2_p_spl_1
  );


  buf

  (
    n6461_o2_p_spl_,
    n6461_o2_p
  );


  buf

  (
    n6461_o2_p_spl_0,
    n6461_o2_p_spl_
  );


  buf

  (
    n6461_o2_p_spl_00,
    n6461_o2_p_spl_0
  );


  buf

  (
    n6461_o2_p_spl_1,
    n6461_o2_p_spl_
  );


  buf

  (
    n2824_lo_buf_o2_n_spl_,
    n2824_lo_buf_o2_n
  );


  buf

  (
    n2824_lo_buf_o2_n_spl_0,
    n2824_lo_buf_o2_n_spl_
  );


  buf

  (
    n2824_lo_buf_o2_n_spl_00,
    n2824_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2824_lo_buf_o2_n_spl_000,
    n2824_lo_buf_o2_n_spl_00
  );


  buf

  (
    n2824_lo_buf_o2_n_spl_001,
    n2824_lo_buf_o2_n_spl_00
  );


  buf

  (
    n2824_lo_buf_o2_n_spl_01,
    n2824_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2824_lo_buf_o2_n_spl_010,
    n2824_lo_buf_o2_n_spl_01
  );


  buf

  (
    n2824_lo_buf_o2_n_spl_1,
    n2824_lo_buf_o2_n_spl_
  );


  buf

  (
    n2824_lo_buf_o2_n_spl_10,
    n2824_lo_buf_o2_n_spl_1
  );


  buf

  (
    n2824_lo_buf_o2_n_spl_11,
    n2824_lo_buf_o2_n_spl_1
  );


  buf

  (
    n6461_o2_n_spl_,
    n6461_o2_n
  );


  buf

  (
    n6461_o2_n_spl_0,
    n6461_o2_n_spl_
  );


  buf

  (
    n6461_o2_n_spl_1,
    n6461_o2_n_spl_
  );


  buf

  (
    g698_n_spl_,
    g698_n
  );


  buf

  (
    g697_p_spl_,
    g697_p
  );


  buf

  (
    n2836_lo_p_spl_,
    n2836_lo_p
  );


  buf

  (
    n2836_lo_p_spl_0,
    n2836_lo_p_spl_
  );


  buf

  (
    n2836_lo_p_spl_00,
    n2836_lo_p_spl_0
  );


  buf

  (
    n2836_lo_p_spl_000,
    n2836_lo_p_spl_00
  );


  buf

  (
    n2836_lo_p_spl_001,
    n2836_lo_p_spl_00
  );


  buf

  (
    n2836_lo_p_spl_01,
    n2836_lo_p_spl_0
  );


  buf

  (
    n2836_lo_p_spl_010,
    n2836_lo_p_spl_01
  );


  buf

  (
    n2836_lo_p_spl_011,
    n2836_lo_p_spl_01
  );


  buf

  (
    n2836_lo_p_spl_1,
    n2836_lo_p_spl_
  );


  buf

  (
    n2836_lo_p_spl_10,
    n2836_lo_p_spl_1
  );


  buf

  (
    n2836_lo_p_spl_100,
    n2836_lo_p_spl_10
  );


  buf

  (
    n2836_lo_p_spl_101,
    n2836_lo_p_spl_10
  );


  buf

  (
    n2836_lo_p_spl_11,
    n2836_lo_p_spl_1
  );


  buf

  (
    n2836_lo_p_spl_110,
    n2836_lo_p_spl_11
  );


  buf

  (
    n2836_lo_n_spl_,
    n2836_lo_n
  );


  buf

  (
    n2836_lo_n_spl_0,
    n2836_lo_n_spl_
  );


  buf

  (
    n2836_lo_n_spl_00,
    n2836_lo_n_spl_0
  );


  buf

  (
    n2836_lo_n_spl_000,
    n2836_lo_n_spl_00
  );


  buf

  (
    n2836_lo_n_spl_001,
    n2836_lo_n_spl_00
  );


  buf

  (
    n2836_lo_n_spl_01,
    n2836_lo_n_spl_0
  );


  buf

  (
    n2836_lo_n_spl_010,
    n2836_lo_n_spl_01
  );


  buf

  (
    n2836_lo_n_spl_011,
    n2836_lo_n_spl_01
  );


  buf

  (
    n2836_lo_n_spl_1,
    n2836_lo_n_spl_
  );


  buf

  (
    n2836_lo_n_spl_10,
    n2836_lo_n_spl_1
  );


  buf

  (
    n2836_lo_n_spl_100,
    n2836_lo_n_spl_10
  );


  buf

  (
    n2836_lo_n_spl_101,
    n2836_lo_n_spl_10
  );


  buf

  (
    n2836_lo_n_spl_11,
    n2836_lo_n_spl_1
  );


  buf

  (
    n2836_lo_n_spl_110,
    n2836_lo_n_spl_11
  );


  buf

  (
    G5109_o2_p_spl_,
    G5109_o2_p
  );


  buf

  (
    G626_o2_n_spl_,
    G626_o2_n
  );


  buf

  (
    G5109_o2_n_spl_,
    G5109_o2_n
  );


  buf

  (
    G626_o2_p_spl_,
    G626_o2_p
  );


  buf

  (
    g701_n_spl_,
    g701_n
  );


  buf

  (
    g701_n_spl_0,
    g701_n_spl_
  );


  buf

  (
    g701_p_spl_,
    g701_p
  );


  buf

  (
    g701_p_spl_0,
    g701_p_spl_
  );


  buf

  (
    g699_p_spl_,
    g699_p
  );


  buf

  (
    g705_n_spl_,
    g705_n
  );


  buf

  (
    g704_n_spl_,
    g704_n
  );


  buf

  (
    g705_p_spl_,
    g705_p
  );


  buf

  (
    g704_p_spl_,
    g704_p
  );


  buf

  (
    g706_n_spl_,
    g706_n
  );


  buf

  (
    g706_n_spl_0,
    g706_n_spl_
  );


  buf

  (
    g706_p_spl_,
    g706_p
  );


  buf

  (
    g706_p_spl_0,
    g706_p_spl_
  );


  buf

  (
    g709_n_spl_,
    g709_n
  );


  buf

  (
    g700_p_spl_,
    g700_p
  );


  buf

  (
    n2848_lo_p_spl_,
    n2848_lo_p
  );


  buf

  (
    n2848_lo_p_spl_0,
    n2848_lo_p_spl_
  );


  buf

  (
    n2848_lo_p_spl_00,
    n2848_lo_p_spl_0
  );


  buf

  (
    n2848_lo_p_spl_000,
    n2848_lo_p_spl_00
  );


  buf

  (
    n2848_lo_p_spl_001,
    n2848_lo_p_spl_00
  );


  buf

  (
    n2848_lo_p_spl_01,
    n2848_lo_p_spl_0
  );


  buf

  (
    n2848_lo_p_spl_010,
    n2848_lo_p_spl_01
  );


  buf

  (
    n2848_lo_p_spl_1,
    n2848_lo_p_spl_
  );


  buf

  (
    n2848_lo_p_spl_10,
    n2848_lo_p_spl_1
  );


  buf

  (
    n2848_lo_p_spl_11,
    n2848_lo_p_spl_1
  );


  buf

  (
    n2848_lo_n_spl_,
    n2848_lo_n
  );


  buf

  (
    n2848_lo_n_spl_0,
    n2848_lo_n_spl_
  );


  buf

  (
    n2848_lo_n_spl_00,
    n2848_lo_n_spl_0
  );


  buf

  (
    n2848_lo_n_spl_000,
    n2848_lo_n_spl_00
  );


  buf

  (
    n2848_lo_n_spl_001,
    n2848_lo_n_spl_00
  );


  buf

  (
    n2848_lo_n_spl_01,
    n2848_lo_n_spl_0
  );


  buf

  (
    n2848_lo_n_spl_010,
    n2848_lo_n_spl_01
  );


  buf

  (
    n2848_lo_n_spl_1,
    n2848_lo_n_spl_
  );


  buf

  (
    n2848_lo_n_spl_10,
    n2848_lo_n_spl_1
  );


  buf

  (
    n2848_lo_n_spl_11,
    n2848_lo_n_spl_1
  );


  buf

  (
    G5172_o2_n_spl_,
    G5172_o2_n
  );


  buf

  (
    G5172_o2_n_spl_0,
    G5172_o2_n_spl_
  );


  buf

  (
    G5172_o2_p_spl_,
    G5172_o2_p
  );


  buf

  (
    G5172_o2_p_spl_0,
    G5172_o2_p_spl_
  );


  buf

  (
    g715_n_spl_,
    g715_n
  );


  buf

  (
    g714_n_spl_,
    g714_n
  );


  buf

  (
    g715_p_spl_,
    g715_p
  );


  buf

  (
    g714_p_spl_,
    g714_p
  );


  buf

  (
    g716_n_spl_,
    g716_n
  );


  buf

  (
    g716_n_spl_0,
    g716_n_spl_
  );


  buf

  (
    g716_p_spl_,
    g716_p
  );


  buf

  (
    g716_p_spl_0,
    g716_p_spl_
  );


  buf

  (
    n6309_o2_p_spl_,
    n6309_o2_p
  );


  buf

  (
    n6309_o2_p_spl_0,
    n6309_o2_p_spl_
  );


  buf

  (
    n6309_o2_n_spl_,
    n6309_o2_n
  );


  buf

  (
    n6309_o2_n_spl_0,
    n6309_o2_n_spl_
  );


  buf

  (
    g720_n_spl_,
    g720_n
  );


  buf

  (
    g719_n_spl_,
    g719_n
  );


  buf

  (
    g720_p_spl_,
    g720_p
  );


  buf

  (
    g719_p_spl_,
    g719_p
  );


  buf

  (
    g721_n_spl_,
    g721_n
  );


  buf

  (
    g721_n_spl_0,
    g721_n_spl_
  );


  buf

  (
    g721_p_spl_,
    g721_p
  );


  buf

  (
    g721_p_spl_0,
    g721_p_spl_
  );


  buf

  (
    g710_p_spl_,
    g710_p
  );


  buf

  (
    g725_n_spl_,
    g725_n
  );


  buf

  (
    g724_n_spl_,
    g724_n
  );


  buf

  (
    g725_p_spl_,
    g725_p
  );


  buf

  (
    g724_p_spl_,
    g724_p
  );


  buf

  (
    g726_n_spl_,
    g726_n
  );


  buf

  (
    g726_n_spl_0,
    g726_n_spl_
  );


  buf

  (
    g726_p_spl_,
    g726_p
  );


  buf

  (
    g726_p_spl_0,
    g726_p_spl_
  );


  buf

  (
    g729_n_spl_,
    g729_n
  );


  buf

  (
    g711_p_spl_,
    g711_p
  );


  buf

  (
    n2764_lo_buf_o2_p_spl_,
    n2764_lo_buf_o2_p
  );


  buf

  (
    n2764_lo_buf_o2_p_spl_0,
    n2764_lo_buf_o2_p_spl_
  );


  buf

  (
    n2764_lo_buf_o2_p_spl_00,
    n2764_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2764_lo_buf_o2_p_spl_1,
    n2764_lo_buf_o2_p_spl_
  );


  buf

  (
    n8086_o2_p_spl_,
    n8086_o2_p
  );


  buf

  (
    n8086_o2_p_spl_0,
    n8086_o2_p_spl_
  );


  buf

  (
    n8086_o2_p_spl_00,
    n8086_o2_p_spl_0
  );


  buf

  (
    n8086_o2_p_spl_01,
    n8086_o2_p_spl_0
  );


  buf

  (
    n8086_o2_p_spl_1,
    n8086_o2_p_spl_
  );


  buf

  (
    n2764_lo_buf_o2_n_spl_,
    n2764_lo_buf_o2_n
  );


  buf

  (
    n2764_lo_buf_o2_n_spl_0,
    n2764_lo_buf_o2_n_spl_
  );


  buf

  (
    n2764_lo_buf_o2_n_spl_00,
    n2764_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2764_lo_buf_o2_n_spl_1,
    n2764_lo_buf_o2_n_spl_
  );


  buf

  (
    n8086_o2_n_spl_,
    n8086_o2_n
  );


  buf

  (
    n8086_o2_n_spl_0,
    n8086_o2_n_spl_
  );


  buf

  (
    n8086_o2_n_spl_00,
    n8086_o2_n_spl_0
  );


  buf

  (
    n8086_o2_n_spl_1,
    n8086_o2_n_spl_
  );


  buf

  (
    G3257_o2_p_spl_,
    G3257_o2_p
  );


  buf

  (
    G3257_o2_p_spl_0,
    G3257_o2_p_spl_
  );


  buf

  (
    G3257_o2_n_spl_,
    G3257_o2_n
  );


  buf

  (
    G3257_o2_n_spl_0,
    G3257_o2_n_spl_
  );


  buf

  (
    g734_n_spl_,
    g734_n
  );


  buf

  (
    g731_p_spl_,
    g731_p
  );


  buf

  (
    n2860_lo_p_spl_,
    n2860_lo_p
  );


  buf

  (
    n2860_lo_p_spl_0,
    n2860_lo_p_spl_
  );


  buf

  (
    n2860_lo_p_spl_00,
    n2860_lo_p_spl_0
  );


  buf

  (
    n2860_lo_p_spl_01,
    n2860_lo_p_spl_0
  );


  buf

  (
    n2860_lo_p_spl_1,
    n2860_lo_p_spl_
  );


  buf

  (
    n2860_lo_p_spl_10,
    n2860_lo_p_spl_1
  );


  buf

  (
    n2860_lo_n_spl_,
    n2860_lo_n
  );


  buf

  (
    n2860_lo_n_spl_0,
    n2860_lo_n_spl_
  );


  buf

  (
    n2860_lo_n_spl_00,
    n2860_lo_n_spl_0
  );


  buf

  (
    n2860_lo_n_spl_01,
    n2860_lo_n_spl_0
  );


  buf

  (
    n2860_lo_n_spl_1,
    n2860_lo_n_spl_
  );


  buf

  (
    n2860_lo_n_spl_10,
    n2860_lo_n_spl_1
  );


  buf

  (
    g738_n_spl_,
    g738_n
  );


  buf

  (
    g737_n_spl_,
    g737_n
  );


  buf

  (
    g738_p_spl_,
    g738_p
  );


  buf

  (
    g737_p_spl_,
    g737_p
  );


  buf

  (
    g739_n_spl_,
    g739_n
  );


  buf

  (
    g739_n_spl_0,
    g739_n_spl_
  );


  buf

  (
    g739_p_spl_,
    g739_p
  );


  buf

  (
    g739_p_spl_0,
    g739_p_spl_
  );


  buf

  (
    n6239_o2_p_spl_,
    n6239_o2_p
  );


  buf

  (
    n6239_o2_p_spl_0,
    n6239_o2_p_spl_
  );


  buf

  (
    n6239_o2_n_spl_,
    n6239_o2_n
  );


  buf

  (
    n6239_o2_n_spl_0,
    n6239_o2_n_spl_
  );


  buf

  (
    g743_n_spl_,
    g743_n
  );


  buf

  (
    g742_n_spl_,
    g742_n
  );


  buf

  (
    g743_p_spl_,
    g743_p
  );


  buf

  (
    g742_p_spl_,
    g742_p
  );


  buf

  (
    g744_n_spl_,
    g744_n
  );


  buf

  (
    g744_n_spl_0,
    g744_n_spl_
  );


  buf

  (
    g744_p_spl_,
    g744_p
  );


  buf

  (
    g744_p_spl_0,
    g744_p_spl_
  );


  buf

  (
    g748_n_spl_,
    g748_n
  );


  buf

  (
    g747_n_spl_,
    g747_n
  );


  buf

  (
    g748_p_spl_,
    g748_p
  );


  buf

  (
    g747_p_spl_,
    g747_p
  );


  buf

  (
    g749_n_spl_,
    g749_n
  );


  buf

  (
    g749_n_spl_0,
    g749_n_spl_
  );


  buf

  (
    g749_p_spl_,
    g749_p
  );


  buf

  (
    g749_p_spl_0,
    g749_p_spl_
  );


  buf

  (
    g753_n_spl_,
    g753_n
  );


  buf

  (
    g752_n_spl_,
    g752_n
  );


  buf

  (
    g753_p_spl_,
    g753_p
  );


  buf

  (
    g752_p_spl_,
    g752_p
  );


  buf

  (
    g754_n_spl_,
    g754_n
  );


  buf

  (
    g754_n_spl_0,
    g754_n_spl_
  );


  buf

  (
    g754_p_spl_,
    g754_p
  );


  buf

  (
    g754_p_spl_0,
    g754_p_spl_
  );


  buf

  (
    g730_p_spl_,
    g730_p
  );


  buf

  (
    g758_n_spl_,
    g758_n
  );


  buf

  (
    g757_n_spl_,
    g757_n
  );


  buf

  (
    g758_p_spl_,
    g758_p
  );


  buf

  (
    g757_p_spl_,
    g757_p
  );


  buf

  (
    g759_n_spl_,
    g759_n
  );


  buf

  (
    g759_n_spl_0,
    g759_n_spl_
  );


  buf

  (
    g759_p_spl_,
    g759_p
  );


  buf

  (
    g759_p_spl_0,
    g759_p_spl_
  );


  buf

  (
    n2776_lo_buf_o2_p_spl_,
    n2776_lo_buf_o2_p
  );


  buf

  (
    n2776_lo_buf_o2_p_spl_0,
    n2776_lo_buf_o2_p_spl_
  );


  buf

  (
    n2776_lo_buf_o2_p_spl_00,
    n2776_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2776_lo_buf_o2_p_spl_000,
    n2776_lo_buf_o2_p_spl_00
  );


  buf

  (
    n2776_lo_buf_o2_p_spl_001,
    n2776_lo_buf_o2_p_spl_00
  );


  buf

  (
    n2776_lo_buf_o2_p_spl_01,
    n2776_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2776_lo_buf_o2_p_spl_010,
    n2776_lo_buf_o2_p_spl_01
  );


  buf

  (
    n2776_lo_buf_o2_p_spl_011,
    n2776_lo_buf_o2_p_spl_01
  );


  buf

  (
    n2776_lo_buf_o2_p_spl_1,
    n2776_lo_buf_o2_p_spl_
  );


  buf

  (
    n2776_lo_buf_o2_p_spl_10,
    n2776_lo_buf_o2_p_spl_1
  );


  buf

  (
    n2776_lo_buf_o2_p_spl_100,
    n2776_lo_buf_o2_p_spl_10
  );


  buf

  (
    n2776_lo_buf_o2_p_spl_101,
    n2776_lo_buf_o2_p_spl_10
  );


  buf

  (
    n2776_lo_buf_o2_p_spl_11,
    n2776_lo_buf_o2_p_spl_1
  );


  buf

  (
    n2776_lo_buf_o2_n_spl_,
    n2776_lo_buf_o2_n
  );


  buf

  (
    n2776_lo_buf_o2_n_spl_0,
    n2776_lo_buf_o2_n_spl_
  );


  buf

  (
    n2776_lo_buf_o2_n_spl_00,
    n2776_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2776_lo_buf_o2_n_spl_000,
    n2776_lo_buf_o2_n_spl_00
  );


  buf

  (
    n2776_lo_buf_o2_n_spl_001,
    n2776_lo_buf_o2_n_spl_00
  );


  buf

  (
    n2776_lo_buf_o2_n_spl_01,
    n2776_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2776_lo_buf_o2_n_spl_010,
    n2776_lo_buf_o2_n_spl_01
  );


  buf

  (
    n2776_lo_buf_o2_n_spl_011,
    n2776_lo_buf_o2_n_spl_01
  );


  buf

  (
    n2776_lo_buf_o2_n_spl_1,
    n2776_lo_buf_o2_n_spl_
  );


  buf

  (
    n2776_lo_buf_o2_n_spl_10,
    n2776_lo_buf_o2_n_spl_1
  );


  buf

  (
    n2776_lo_buf_o2_n_spl_100,
    n2776_lo_buf_o2_n_spl_10
  );


  buf

  (
    n2776_lo_buf_o2_n_spl_101,
    n2776_lo_buf_o2_n_spl_10
  );


  buf

  (
    n2776_lo_buf_o2_n_spl_11,
    n2776_lo_buf_o2_n_spl_1
  );


  buf

  (
    g762_n_spl_,
    g762_n
  );


  buf

  (
    g736_p_spl_,
    g736_p
  );


  buf

  (
    n7909_o2_p_spl_,
    n7909_o2_p
  );


  buf

  (
    n7909_o2_p_spl_0,
    n7909_o2_p_spl_
  );


  buf

  (
    n7909_o2_p_spl_00,
    n7909_o2_p_spl_0
  );


  buf

  (
    n7909_o2_p_spl_01,
    n7909_o2_p_spl_0
  );


  buf

  (
    n7909_o2_p_spl_1,
    n7909_o2_p_spl_
  );


  buf

  (
    n7909_o2_p_spl_10,
    n7909_o2_p_spl_1
  );


  buf

  (
    n7909_o2_n_spl_,
    n7909_o2_n
  );


  buf

  (
    n7909_o2_n_spl_0,
    n7909_o2_n_spl_
  );


  buf

  (
    n7909_o2_n_spl_00,
    n7909_o2_n_spl_0
  );


  buf

  (
    n7909_o2_n_spl_1,
    n7909_o2_n_spl_
  );


  buf

  (
    g766_n_spl_,
    g766_n
  );


  buf

  (
    g765_n_spl_,
    g765_n
  );


  buf

  (
    g766_p_spl_,
    g766_p
  );


  buf

  (
    g765_p_spl_,
    g765_p
  );


  buf

  (
    g767_n_spl_,
    g767_n
  );


  buf

  (
    g767_n_spl_0,
    g767_n_spl_
  );


  buf

  (
    g767_p_spl_,
    g767_p
  );


  buf

  (
    g767_p_spl_0,
    g767_p_spl_
  );


  buf

  (
    g735_p_spl_,
    g735_p
  );


  buf

  (
    g771_n_spl_,
    g771_n
  );


  buf

  (
    g770_n_spl_,
    g770_n
  );


  buf

  (
    g771_p_spl_,
    g771_p
  );


  buf

  (
    g770_p_spl_,
    g770_p
  );


  buf

  (
    g772_n_spl_,
    g772_n
  );


  buf

  (
    g772_n_spl_0,
    g772_n_spl_
  );


  buf

  (
    g772_p_spl_,
    g772_p
  );


  buf

  (
    g772_p_spl_0,
    g772_p_spl_
  );


  buf

  (
    g775_n_spl_,
    g775_n
  );


  buf

  (
    g763_p_spl_,
    g763_p
  );


  buf

  (
    n2488_lo_buf_o2_p_spl_,
    n2488_lo_buf_o2_p
  );


  buf

  (
    n2488_lo_buf_o2_p_spl_0,
    n2488_lo_buf_o2_p_spl_
  );


  buf

  (
    n2488_lo_buf_o2_p_spl_00,
    n2488_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2488_lo_buf_o2_p_spl_1,
    n2488_lo_buf_o2_p_spl_
  );


  buf

  (
    n2704_lo_buf_o2_p_spl_,
    n2704_lo_buf_o2_p
  );


  buf

  (
    n2704_lo_buf_o2_p_spl_0,
    n2704_lo_buf_o2_p_spl_
  );


  buf

  (
    n2488_lo_buf_o2_n_spl_,
    n2488_lo_buf_o2_n
  );


  buf

  (
    n2488_lo_buf_o2_n_spl_0,
    n2488_lo_buf_o2_n_spl_
  );


  buf

  (
    n2488_lo_buf_o2_n_spl_00,
    n2488_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2488_lo_buf_o2_n_spl_1,
    n2488_lo_buf_o2_n_spl_
  );


  buf

  (
    n2704_lo_buf_o2_n_spl_,
    n2704_lo_buf_o2_n
  );


  buf

  (
    n2704_lo_buf_o2_n_spl_0,
    n2704_lo_buf_o2_n_spl_
  );


  buf

  (
    G1580_o2_n_spl_,
    G1580_o2_n
  );


  buf

  (
    G1507_o2_n_spl_,
    G1507_o2_n
  );


  buf

  (
    G1580_o2_p_spl_,
    G1580_o2_p
  );


  buf

  (
    G1507_o2_p_spl_,
    G1507_o2_p
  );


  buf

  (
    g778_n_spl_,
    g778_n
  );


  buf

  (
    g778_n_spl_0,
    g778_n_spl_
  );


  buf

  (
    g778_p_spl_,
    g778_p
  );


  buf

  (
    g778_p_spl_0,
    g778_p_spl_
  );


  buf

  (
    n2785_lo_p_spl_,
    n2785_lo_p
  );


  buf

  (
    n2785_lo_p_spl_0,
    n2785_lo_p_spl_
  );


  buf

  (
    n2785_lo_p_spl_00,
    n2785_lo_p_spl_0
  );


  buf

  (
    n2785_lo_p_spl_000,
    n2785_lo_p_spl_00
  );


  buf

  (
    n2785_lo_p_spl_001,
    n2785_lo_p_spl_00
  );


  buf

  (
    n2785_lo_p_spl_01,
    n2785_lo_p_spl_0
  );


  buf

  (
    n2785_lo_p_spl_010,
    n2785_lo_p_spl_01
  );


  buf

  (
    n2785_lo_p_spl_011,
    n2785_lo_p_spl_01
  );


  buf

  (
    n2785_lo_p_spl_1,
    n2785_lo_p_spl_
  );


  buf

  (
    n2785_lo_p_spl_10,
    n2785_lo_p_spl_1
  );


  buf

  (
    n2785_lo_p_spl_100,
    n2785_lo_p_spl_10
  );


  buf

  (
    n2785_lo_p_spl_101,
    n2785_lo_p_spl_10
  );


  buf

  (
    n2785_lo_p_spl_11,
    n2785_lo_p_spl_1
  );


  buf

  (
    n2785_lo_p_spl_110,
    n2785_lo_p_spl_11
  );


  buf

  (
    n2785_lo_p_spl_111,
    n2785_lo_p_spl_11
  );


  buf

  (
    n2785_lo_n_spl_,
    n2785_lo_n
  );


  buf

  (
    n2785_lo_n_spl_0,
    n2785_lo_n_spl_
  );


  buf

  (
    n2785_lo_n_spl_00,
    n2785_lo_n_spl_0
  );


  buf

  (
    n2785_lo_n_spl_000,
    n2785_lo_n_spl_00
  );


  buf

  (
    n2785_lo_n_spl_001,
    n2785_lo_n_spl_00
  );


  buf

  (
    n2785_lo_n_spl_01,
    n2785_lo_n_spl_0
  );


  buf

  (
    n2785_lo_n_spl_010,
    n2785_lo_n_spl_01
  );


  buf

  (
    n2785_lo_n_spl_011,
    n2785_lo_n_spl_01
  );


  buf

  (
    n2785_lo_n_spl_1,
    n2785_lo_n_spl_
  );


  buf

  (
    n2785_lo_n_spl_10,
    n2785_lo_n_spl_1
  );


  buf

  (
    n2785_lo_n_spl_100,
    n2785_lo_n_spl_10
  );


  buf

  (
    n2785_lo_n_spl_101,
    n2785_lo_n_spl_10
  );


  buf

  (
    n2785_lo_n_spl_11,
    n2785_lo_n_spl_1
  );


  buf

  (
    n2785_lo_n_spl_110,
    n2785_lo_n_spl_11
  );


  buf

  (
    n2785_lo_n_spl_111,
    n2785_lo_n_spl_11
  );


  buf

  (
    g781_n_spl_,
    g781_n
  );


  buf

  (
    g777_p_spl_,
    g777_p
  );


  buf

  (
    G3364_o2_p_spl_,
    G3364_o2_p
  );


  buf

  (
    G659_o2_n_spl_,
    G659_o2_n
  );


  buf

  (
    G3364_o2_n_spl_,
    G3364_o2_n
  );


  buf

  (
    G659_o2_p_spl_,
    G659_o2_p
  );


  buf

  (
    g784_n_spl_,
    g784_n
  );


  buf

  (
    g784_n_spl_0,
    g784_n_spl_
  );


  buf

  (
    g784_p_spl_,
    g784_p
  );


  buf

  (
    g784_p_spl_0,
    g784_p_spl_
  );


  buf

  (
    g788_n_spl_,
    g788_n
  );


  buf

  (
    g787_n_spl_,
    g787_n
  );


  buf

  (
    g788_p_spl_,
    g788_p
  );


  buf

  (
    g787_p_spl_,
    g787_p
  );


  buf

  (
    g789_n_spl_,
    g789_n
  );


  buf

  (
    g789_n_spl_0,
    g789_n_spl_
  );


  buf

  (
    g789_p_spl_,
    g789_p
  );


  buf

  (
    g789_p_spl_0,
    g789_p_spl_
  );


  buf

  (
    g793_n_spl_,
    g793_n
  );


  buf

  (
    g792_n_spl_,
    g792_n
  );


  buf

  (
    g793_p_spl_,
    g793_p
  );


  buf

  (
    g792_p_spl_,
    g792_p
  );


  buf

  (
    g794_n_spl_,
    g794_n
  );


  buf

  (
    g794_n_spl_0,
    g794_n_spl_
  );


  buf

  (
    g794_p_spl_,
    g794_p
  );


  buf

  (
    g794_p_spl_0,
    g794_p_spl_
  );


  buf

  (
    g776_p_spl_,
    g776_p
  );


  buf

  (
    g798_n_spl_,
    g798_n
  );


  buf

  (
    g797_n_spl_,
    g797_n
  );


  buf

  (
    g798_p_spl_,
    g798_p
  );


  buf

  (
    g797_p_spl_,
    g797_p
  );


  buf

  (
    g799_n_spl_,
    g799_n
  );


  buf

  (
    g799_n_spl_0,
    g799_n_spl_
  );


  buf

  (
    g799_p_spl_,
    g799_p
  );


  buf

  (
    g799_p_spl_0,
    g799_p_spl_
  );


  buf

  (
    g802_n_spl_,
    g802_n
  );


  buf

  (
    g782_p_spl_,
    g782_p
  );


  buf

  (
    n2716_lo_buf_o2_p_spl_,
    n2716_lo_buf_o2_p
  );


  buf

  (
    n2716_lo_buf_o2_p_spl_0,
    n2716_lo_buf_o2_p_spl_
  );


  buf

  (
    n2716_lo_buf_o2_p_spl_00,
    n2716_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2716_lo_buf_o2_p_spl_000,
    n2716_lo_buf_o2_p_spl_00
  );


  buf

  (
    n2716_lo_buf_o2_p_spl_01,
    n2716_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2716_lo_buf_o2_p_spl_1,
    n2716_lo_buf_o2_p_spl_
  );


  buf

  (
    n2716_lo_buf_o2_p_spl_10,
    n2716_lo_buf_o2_p_spl_1
  );


  buf

  (
    n2716_lo_buf_o2_p_spl_11,
    n2716_lo_buf_o2_p_spl_1
  );


  buf

  (
    n2716_lo_buf_o2_n_spl_,
    n2716_lo_buf_o2_n
  );


  buf

  (
    n2716_lo_buf_o2_n_spl_0,
    n2716_lo_buf_o2_n_spl_
  );


  buf

  (
    n2716_lo_buf_o2_n_spl_00,
    n2716_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2716_lo_buf_o2_n_spl_000,
    n2716_lo_buf_o2_n_spl_00
  );


  buf

  (
    n2716_lo_buf_o2_n_spl_01,
    n2716_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2716_lo_buf_o2_n_spl_1,
    n2716_lo_buf_o2_n_spl_
  );


  buf

  (
    n2716_lo_buf_o2_n_spl_10,
    n2716_lo_buf_o2_n_spl_1
  );


  buf

  (
    n2716_lo_buf_o2_n_spl_11,
    n2716_lo_buf_o2_n_spl_1
  );


  buf

  (
    G1630_o2_p_spl_,
    G1630_o2_p
  );


  buf

  (
    G1630_o2_p_spl_0,
    G1630_o2_p_spl_
  );


  buf

  (
    G1630_o2_n_spl_,
    G1630_o2_n
  );


  buf

  (
    G1630_o2_n_spl_0,
    G1630_o2_n_spl_
  );


  buf

  (
    n2500_lo_buf_o2_p_spl_,
    n2500_lo_buf_o2_p
  );


  buf

  (
    n2500_lo_buf_o2_p_spl_0,
    n2500_lo_buf_o2_p_spl_
  );


  buf

  (
    n2500_lo_buf_o2_p_spl_00,
    n2500_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2500_lo_buf_o2_p_spl_01,
    n2500_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2500_lo_buf_o2_p_spl_1,
    n2500_lo_buf_o2_p_spl_
  );


  buf

  (
    n2500_lo_buf_o2_n_spl_,
    n2500_lo_buf_o2_n
  );


  buf

  (
    n2500_lo_buf_o2_n_spl_0,
    n2500_lo_buf_o2_n_spl_
  );


  buf

  (
    n2500_lo_buf_o2_n_spl_00,
    n2500_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2500_lo_buf_o2_n_spl_1,
    n2500_lo_buf_o2_n_spl_
  );


  buf

  (
    g808_n_spl_,
    g808_n
  );


  buf

  (
    g807_n_spl_,
    g807_n
  );


  buf

  (
    g808_p_spl_,
    g808_p
  );


  buf

  (
    g807_p_spl_,
    g807_p
  );


  buf

  (
    g809_n_spl_,
    g809_n
  );


  buf

  (
    g809_n_spl_0,
    g809_n_spl_
  );


  buf

  (
    g809_p_spl_,
    g809_p
  );


  buf

  (
    g809_p_spl_0,
    g809_p_spl_
  );


  buf

  (
    g783_p_spl_,
    g783_p
  );


  buf

  (
    g813_n_spl_,
    g813_n
  );


  buf

  (
    g812_n_spl_,
    g812_n
  );


  buf

  (
    g813_p_spl_,
    g813_p
  );


  buf

  (
    g812_p_spl_,
    g812_p
  );


  buf

  (
    g814_n_spl_,
    g814_n
  );


  buf

  (
    g814_n_spl_0,
    g814_n_spl_
  );


  buf

  (
    g814_p_spl_,
    g814_p
  );


  buf

  (
    g814_p_spl_0,
    g814_p_spl_
  );


  buf

  (
    n2812_lo_buf_o2_p_spl_,
    n2812_lo_buf_o2_p
  );


  buf

  (
    n2812_lo_buf_o2_p_spl_0,
    n2812_lo_buf_o2_p_spl_
  );


  buf

  (
    n2812_lo_buf_o2_p_spl_00,
    n2812_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2812_lo_buf_o2_p_spl_01,
    n2812_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2812_lo_buf_o2_p_spl_1,
    n2812_lo_buf_o2_p_spl_
  );


  buf

  (
    n5779_o2_p_spl_,
    n5779_o2_p
  );


  buf

  (
    n5779_o2_p_spl_0,
    n5779_o2_p_spl_
  );


  buf

  (
    n5779_o2_p_spl_1,
    n5779_o2_p_spl_
  );


  buf

  (
    n2812_lo_buf_o2_n_spl_,
    n2812_lo_buf_o2_n
  );


  buf

  (
    n2812_lo_buf_o2_n_spl_0,
    n2812_lo_buf_o2_n_spl_
  );


  buf

  (
    n2812_lo_buf_o2_n_spl_00,
    n2812_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2812_lo_buf_o2_n_spl_01,
    n2812_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2812_lo_buf_o2_n_spl_1,
    n2812_lo_buf_o2_n_spl_
  );


  buf

  (
    n5779_o2_n_spl_,
    n5779_o2_n
  );


  buf

  (
    n5779_o2_n_spl_0,
    n5779_o2_n_spl_
  );


  buf

  (
    n2800_lo_buf_o2_p_spl_,
    n2800_lo_buf_o2_p
  );


  buf

  (
    n2800_lo_buf_o2_n_spl_,
    n2800_lo_buf_o2_n
  );


  buf

  (
    n5792_o2_p_spl_,
    n5792_o2_p
  );


  buf

  (
    n5792_o2_p_spl_0,
    n5792_o2_p_spl_
  );


  buf

  (
    n5792_o2_p_spl_1,
    n5792_o2_p_spl_
  );


  buf

  (
    n5792_o2_n_spl_,
    n5792_o2_n
  );


  buf

  (
    n5792_o2_n_spl_0,
    n5792_o2_n_spl_
  );


  buf

  (
    n5792_o2_n_spl_1,
    n5792_o2_n_spl_
  );


  buf

  (
    g821_n_spl_,
    g821_n
  );


  buf

  (
    g820_n_spl_,
    g820_n
  );


  buf

  (
    g821_p_spl_,
    g821_p
  );


  buf

  (
    g820_p_spl_,
    g820_p
  );


  buf

  (
    g822_n_spl_,
    g822_n
  );


  buf

  (
    g822_n_spl_0,
    g822_n_spl_
  );


  buf

  (
    g822_p_spl_,
    g822_p
  );


  buf

  (
    g822_p_spl_0,
    g822_p_spl_
  );


  buf

  (
    g823_n_spl_,
    g823_n
  );


  buf

  (
    g819_n_spl_,
    g819_n
  );


  buf

  (
    g823_p_spl_,
    g823_p
  );


  buf

  (
    g819_p_spl_,
    g819_p
  );


  buf

  (
    g824_n_spl_,
    g824_n
  );


  buf

  (
    g824_n_spl_0,
    g824_n_spl_
  );


  buf

  (
    g824_p_spl_,
    g824_p
  );


  buf

  (
    g824_p_spl_0,
    g824_p_spl_
  );


  buf

  (
    g828_n_spl_,
    g828_n
  );


  buf

  (
    g827_n_spl_,
    g827_n
  );


  buf

  (
    g828_p_spl_,
    g828_p
  );


  buf

  (
    g827_p_spl_,
    g827_p
  );


  buf

  (
    g829_n_spl_,
    g829_n
  );


  buf

  (
    g829_n_spl_0,
    g829_n_spl_
  );


  buf

  (
    g829_p_spl_,
    g829_p
  );


  buf

  (
    g829_p_spl_0,
    g829_p_spl_
  );


  buf

  (
    g830_n_spl_,
    g830_n
  );


  buf

  (
    g818_n_spl_,
    g818_n
  );


  buf

  (
    g830_p_spl_,
    g830_p
  );


  buf

  (
    g818_p_spl_,
    g818_p
  );


  buf

  (
    g831_n_spl_,
    g831_n
  );


  buf

  (
    g831_n_spl_0,
    g831_n_spl_
  );


  buf

  (
    g831_p_spl_,
    g831_p
  );


  buf

  (
    g831_p_spl_0,
    g831_p_spl_
  );


  buf

  (
    g835_n_spl_,
    g835_n
  );


  buf

  (
    g834_n_spl_,
    g834_n
  );


  buf

  (
    g835_p_spl_,
    g835_p
  );


  buf

  (
    g834_p_spl_,
    g834_p
  );


  buf

  (
    g836_n_spl_,
    g836_n
  );


  buf

  (
    g836_n_spl_0,
    g836_n_spl_
  );


  buf

  (
    g836_p_spl_,
    g836_p
  );


  buf

  (
    g836_p_spl_0,
    g836_p_spl_
  );


  buf

  (
    G4034_o2_n_spl_,
    G4034_o2_n
  );


  buf

  (
    G4034_o2_n_spl_0,
    G4034_o2_n_spl_
  );


  buf

  (
    G4034_o2_p_spl_,
    G4034_o2_p
  );


  buf

  (
    G4034_o2_p_spl_0,
    G4034_o2_p_spl_
  );


  buf

  (
    g846_n_spl_,
    g846_n
  );


  buf

  (
    g845_n_spl_,
    g845_n
  );


  buf

  (
    g846_p_spl_,
    g846_p
  );


  buf

  (
    g845_p_spl_,
    g845_p
  );


  buf

  (
    g847_n_spl_,
    g847_n
  );


  buf

  (
    g847_n_spl_0,
    g847_n_spl_
  );


  buf

  (
    g847_p_spl_,
    g847_p
  );


  buf

  (
    g847_p_spl_0,
    g847_p_spl_
  );


  buf

  (
    n5842_o2_p_spl_,
    n5842_o2_p
  );


  buf

  (
    n5842_o2_p_spl_0,
    n5842_o2_p_spl_
  );


  buf

  (
    n5842_o2_p_spl_1,
    n5842_o2_p_spl_
  );


  buf

  (
    n5842_o2_n_spl_,
    n5842_o2_n
  );


  buf

  (
    n5842_o2_n_spl_0,
    n5842_o2_n_spl_
  );


  buf

  (
    g851_n_spl_,
    g851_n
  );


  buf

  (
    g850_n_spl_,
    g850_n
  );


  buf

  (
    g851_p_spl_,
    g851_p
  );


  buf

  (
    g850_p_spl_,
    g850_p
  );


  buf

  (
    g852_n_spl_,
    g852_n
  );


  buf

  (
    g852_n_spl_0,
    g852_n_spl_
  );


  buf

  (
    g852_p_spl_,
    g852_p
  );


  buf

  (
    g852_p_spl_0,
    g852_p_spl_
  );


  buf

  (
    g853_n_spl_,
    g853_n
  );


  buf

  (
    g842_n_spl_,
    g842_n
  );


  buf

  (
    g853_p_spl_,
    g853_p
  );


  buf

  (
    g842_p_spl_,
    g842_p
  );


  buf

  (
    g854_n_spl_,
    g854_n
  );


  buf

  (
    g854_n_spl_0,
    g854_n_spl_
  );


  buf

  (
    g854_p_spl_,
    g854_p
  );


  buf

  (
    g854_p_spl_0,
    g854_p_spl_
  );


  buf

  (
    g858_n_spl_,
    g858_n
  );


  buf

  (
    g857_n_spl_,
    g857_n
  );


  buf

  (
    g858_p_spl_,
    g858_p
  );


  buf

  (
    g857_p_spl_,
    g857_p
  );


  buf

  (
    g859_n_spl_,
    g859_n
  );


  buf

  (
    g859_n_spl_0,
    g859_n_spl_
  );


  buf

  (
    g859_p_spl_,
    g859_p
  );


  buf

  (
    g859_p_spl_0,
    g859_p_spl_
  );


  buf

  (
    g860_n_spl_,
    g860_n
  );


  buf

  (
    g839_n_spl_,
    g839_n
  );


  buf

  (
    g860_p_spl_,
    g860_p
  );


  buf

  (
    g839_p_spl_,
    g839_p
  );


  buf

  (
    g865_n_spl_,
    g865_n
  );


  buf

  (
    g864_n_spl_,
    g864_n
  );


  buf

  (
    g865_p_spl_,
    g865_p
  );


  buf

  (
    g864_p_spl_,
    g864_p
  );


  buf

  (
    g866_n_spl_,
    g866_n
  );


  buf

  (
    g866_n_spl_0,
    g866_n_spl_
  );


  buf

  (
    g866_p_spl_,
    g866_p
  );


  buf

  (
    g866_p_spl_0,
    g866_p_spl_
  );


  buf

  (
    n5863_o2_p_spl_,
    n5863_o2_p
  );


  buf

  (
    n5863_o2_p_spl_0,
    n5863_o2_p_spl_
  );


  buf

  (
    n5863_o2_p_spl_1,
    n5863_o2_p_spl_
  );


  buf

  (
    n5863_o2_n_spl_,
    n5863_o2_n
  );


  buf

  (
    n5863_o2_n_spl_0,
    n5863_o2_n_spl_
  );


  buf

  (
    g870_n_spl_,
    g870_n
  );


  buf

  (
    g869_n_spl_,
    g869_n
  );


  buf

  (
    g870_p_spl_,
    g870_p
  );


  buf

  (
    g869_p_spl_,
    g869_p
  );


  buf

  (
    g871_n_spl_,
    g871_n
  );


  buf

  (
    g871_n_spl_0,
    g871_n_spl_
  );


  buf

  (
    g871_p_spl_,
    g871_p
  );


  buf

  (
    g871_p_spl_0,
    g871_p_spl_
  );


  buf

  (
    G4220_o2_n_spl_,
    G4220_o2_n
  );


  buf

  (
    G4217_o2_n_spl_,
    G4217_o2_n
  );


  buf

  (
    G4220_o2_p_spl_,
    G4220_o2_p
  );


  buf

  (
    G4217_o2_p_spl_,
    G4217_o2_p
  );


  buf

  (
    g875_n_spl_,
    g875_n
  );


  buf

  (
    g875_n_spl_0,
    g875_n_spl_
  );


  buf

  (
    g875_p_spl_,
    g875_p
  );


  buf

  (
    g875_p_spl_0,
    g875_p_spl_
  );


  buf

  (
    n5881_o2_p_spl_,
    n5881_o2_p
  );


  buf

  (
    n5881_o2_p_spl_0,
    n5881_o2_p_spl_
  );


  buf

  (
    n5881_o2_p_spl_1,
    n5881_o2_p_spl_
  );


  buf

  (
    n5881_o2_n_spl_,
    n5881_o2_n
  );


  buf

  (
    n5881_o2_n_spl_0,
    n5881_o2_n_spl_
  );


  buf

  (
    g879_n_spl_,
    g879_n
  );


  buf

  (
    g878_n_spl_,
    g878_n
  );


  buf

  (
    g879_p_spl_,
    g879_p
  );


  buf

  (
    g878_p_spl_,
    g878_p
  );


  buf

  (
    g880_n_spl_,
    g880_n
  );


  buf

  (
    g880_n_spl_0,
    g880_n_spl_
  );


  buf

  (
    g880_p_spl_,
    g880_p
  );


  buf

  (
    g880_p_spl_0,
    g880_p_spl_
  );


  buf

  (
    g881_n_spl_,
    g881_n
  );


  buf

  (
    g874_n_spl_,
    g874_n
  );


  buf

  (
    g881_p_spl_,
    g881_p
  );


  buf

  (
    g874_p_spl_,
    g874_p
  );


  buf

  (
    g882_n_spl_,
    g882_n
  );


  buf

  (
    g882_n_spl_0,
    g882_n_spl_
  );


  buf

  (
    g882_p_spl_,
    g882_p
  );


  buf

  (
    g882_p_spl_0,
    g882_p_spl_
  );


  buf

  (
    g886_n_spl_,
    g886_n
  );


  buf

  (
    g885_n_spl_,
    g885_n
  );


  buf

  (
    g886_p_spl_,
    g886_p
  );


  buf

  (
    g885_p_spl_,
    g885_p
  );


  buf

  (
    g887_n_spl_,
    g887_n
  );


  buf

  (
    g887_n_spl_0,
    g887_n_spl_
  );


  buf

  (
    g887_p_spl_,
    g887_p
  );


  buf

  (
    g887_p_spl_0,
    g887_p_spl_
  );


  buf

  (
    n5930_o2_p_spl_,
    n5930_o2_p
  );


  buf

  (
    n5930_o2_p_spl_0,
    n5930_o2_p_spl_
  );


  buf

  (
    n5930_o2_p_spl_1,
    n5930_o2_p_spl_
  );


  buf

  (
    n5930_o2_n_spl_,
    n5930_o2_n
  );


  buf

  (
    n5930_o2_n_spl_0,
    n5930_o2_n_spl_
  );


  buf

  (
    n5930_o2_n_spl_1,
    n5930_o2_n_spl_
  );


  buf

  (
    g895_n_spl_,
    g895_n
  );


  buf

  (
    g894_n_spl_,
    g894_n
  );


  buf

  (
    g895_p_spl_,
    g895_p
  );


  buf

  (
    g894_p_spl_,
    g894_p
  );


  buf

  (
    g896_n_spl_,
    g896_n
  );


  buf

  (
    g896_n_spl_0,
    g896_n_spl_
  );


  buf

  (
    g896_p_spl_,
    g896_p
  );


  buf

  (
    g896_p_spl_0,
    g896_p_spl_
  );


  buf

  (
    g897_n_spl_,
    g897_n
  );


  buf

  (
    g893_n_spl_,
    g893_n
  );


  buf

  (
    g897_p_spl_,
    g897_p
  );


  buf

  (
    g893_p_spl_,
    g893_p
  );


  buf

  (
    g898_n_spl_,
    g898_n
  );


  buf

  (
    g898_n_spl_0,
    g898_n_spl_
  );


  buf

  (
    g898_p_spl_,
    g898_p
  );


  buf

  (
    g898_p_spl_0,
    g898_p_spl_
  );


  buf

  (
    g902_n_spl_,
    g902_n
  );


  buf

  (
    g901_n_spl_,
    g901_n
  );


  buf

  (
    g902_p_spl_,
    g902_p
  );


  buf

  (
    g901_p_spl_,
    g901_p
  );


  buf

  (
    g903_n_spl_,
    g903_n
  );


  buf

  (
    g903_n_spl_0,
    g903_n_spl_
  );


  buf

  (
    g903_p_spl_,
    g903_p
  );


  buf

  (
    g903_p_spl_0,
    g903_p_spl_
  );


  buf

  (
    g904_n_spl_,
    g904_n
  );


  buf

  (
    g890_n_spl_,
    g890_n
  );


  buf

  (
    g904_p_spl_,
    g904_p
  );


  buf

  (
    g890_p_spl_,
    g890_p
  );


  buf

  (
    g905_n_spl_,
    g905_n
  );


  buf

  (
    g905_n_spl_0,
    g905_n_spl_
  );


  buf

  (
    g905_p_spl_,
    g905_p
  );


  buf

  (
    g905_p_spl_0,
    g905_p_spl_
  );


  buf

  (
    g909_n_spl_,
    g909_n
  );


  buf

  (
    g908_n_spl_,
    g908_n
  );


  buf

  (
    g909_p_spl_,
    g909_p
  );


  buf

  (
    g908_p_spl_,
    g908_p
  );


  buf

  (
    g910_n_spl_,
    g910_n
  );


  buf

  (
    g910_n_spl_0,
    g910_n_spl_
  );


  buf

  (
    g910_p_spl_,
    g910_p
  );


  buf

  (
    g910_p_spl_0,
    g910_p_spl_
  );


  buf

  (
    G4556_o2_n_spl_,
    G4556_o2_n
  );


  buf

  (
    G4556_o2_n_spl_0,
    G4556_o2_n_spl_
  );


  buf

  (
    G4556_o2_p_spl_,
    G4556_o2_p
  );


  buf

  (
    G4556_o2_p_spl_0,
    G4556_o2_p_spl_
  );


  buf

  (
    g920_n_spl_,
    g920_n
  );


  buf

  (
    g919_n_spl_,
    g919_n
  );


  buf

  (
    g920_p_spl_,
    g920_p
  );


  buf

  (
    g919_p_spl_,
    g919_p
  );


  buf

  (
    g921_n_spl_,
    g921_n
  );


  buf

  (
    g921_n_spl_0,
    g921_n_spl_
  );


  buf

  (
    g921_p_spl_,
    g921_p
  );


  buf

  (
    g921_p_spl_0,
    g921_p_spl_
  );


  buf

  (
    n5959_o2_p_spl_,
    n5959_o2_p
  );


  buf

  (
    n5959_o2_p_spl_0,
    n5959_o2_p_spl_
  );


  buf

  (
    n5959_o2_p_spl_1,
    n5959_o2_p_spl_
  );


  buf

  (
    n5959_o2_n_spl_,
    n5959_o2_n
  );


  buf

  (
    n5959_o2_n_spl_0,
    n5959_o2_n_spl_
  );


  buf

  (
    g925_n_spl_,
    g925_n
  );


  buf

  (
    g924_n_spl_,
    g924_n
  );


  buf

  (
    g925_p_spl_,
    g925_p
  );


  buf

  (
    g924_p_spl_,
    g924_p
  );


  buf

  (
    g926_n_spl_,
    g926_n
  );


  buf

  (
    g926_n_spl_0,
    g926_n_spl_
  );


  buf

  (
    g926_p_spl_,
    g926_p
  );


  buf

  (
    g926_p_spl_0,
    g926_p_spl_
  );


  buf

  (
    g927_n_spl_,
    g927_n
  );


  buf

  (
    g916_n_spl_,
    g916_n
  );


  buf

  (
    g927_p_spl_,
    g927_p
  );


  buf

  (
    g916_p_spl_,
    g916_p
  );


  buf

  (
    g928_n_spl_,
    g928_n
  );


  buf

  (
    g928_n_spl_0,
    g928_n_spl_
  );


  buf

  (
    g928_p_spl_,
    g928_p
  );


  buf

  (
    g928_p_spl_0,
    g928_p_spl_
  );


  buf

  (
    g932_n_spl_,
    g932_n
  );


  buf

  (
    g931_n_spl_,
    g931_n
  );


  buf

  (
    g932_p_spl_,
    g932_p
  );


  buf

  (
    g931_p_spl_,
    g931_p
  );


  buf

  (
    g933_n_spl_,
    g933_n
  );


  buf

  (
    g933_n_spl_0,
    g933_n_spl_
  );


  buf

  (
    g933_p_spl_,
    g933_p
  );


  buf

  (
    g933_p_spl_0,
    g933_p_spl_
  );


  buf

  (
    g934_n_spl_,
    g934_n
  );


  buf

  (
    g913_n_spl_,
    g913_n
  );


  buf

  (
    g934_p_spl_,
    g934_p
  );


  buf

  (
    g913_p_spl_,
    g913_p
  );


  buf

  (
    g939_n_spl_,
    g939_n
  );


  buf

  (
    g938_n_spl_,
    g938_n
  );


  buf

  (
    g939_p_spl_,
    g939_p
  );


  buf

  (
    g938_p_spl_,
    g938_p
  );


  buf

  (
    g940_n_spl_,
    g940_n
  );


  buf

  (
    g940_n_spl_0,
    g940_n_spl_
  );


  buf

  (
    g940_p_spl_,
    g940_p
  );


  buf

  (
    g940_p_spl_0,
    g940_p_spl_
  );


  buf

  (
    n5981_o2_p_spl_,
    n5981_o2_p
  );


  buf

  (
    n5981_o2_p_spl_0,
    n5981_o2_p_spl_
  );


  buf

  (
    n5981_o2_p_spl_1,
    n5981_o2_p_spl_
  );


  buf

  (
    n5981_o2_n_spl_,
    n5981_o2_n
  );


  buf

  (
    n5981_o2_n_spl_0,
    n5981_o2_n_spl_
  );


  buf

  (
    g944_n_spl_,
    g944_n
  );


  buf

  (
    g943_n_spl_,
    g943_n
  );


  buf

  (
    g944_p_spl_,
    g944_p
  );


  buf

  (
    g943_p_spl_,
    g943_p
  );


  buf

  (
    g945_n_spl_,
    g945_n
  );


  buf

  (
    g945_n_spl_0,
    g945_n_spl_
  );


  buf

  (
    g945_p_spl_,
    g945_p
  );


  buf

  (
    g945_p_spl_0,
    g945_p_spl_
  );


  buf

  (
    G4719_o2_n_spl_,
    G4719_o2_n
  );


  buf

  (
    G4716_o2_n_spl_,
    G4716_o2_n
  );


  buf

  (
    G4719_o2_p_spl_,
    G4719_o2_p
  );


  buf

  (
    G4716_o2_p_spl_,
    G4716_o2_p
  );


  buf

  (
    g949_n_spl_,
    g949_n
  );


  buf

  (
    g949_n_spl_0,
    g949_n_spl_
  );


  buf

  (
    g949_p_spl_,
    g949_p
  );


  buf

  (
    g949_p_spl_0,
    g949_p_spl_
  );


  buf

  (
    n6042_o2_p_spl_,
    n6042_o2_p
  );


  buf

  (
    n6042_o2_p_spl_0,
    n6042_o2_p_spl_
  );


  buf

  (
    n6042_o2_p_spl_1,
    n6042_o2_p_spl_
  );


  buf

  (
    n6042_o2_n_spl_,
    n6042_o2_n
  );


  buf

  (
    n6042_o2_n_spl_0,
    n6042_o2_n_spl_
  );


  buf

  (
    g953_n_spl_,
    g953_n
  );


  buf

  (
    g952_n_spl_,
    g952_n
  );


  buf

  (
    g953_p_spl_,
    g953_p
  );


  buf

  (
    g952_p_spl_,
    g952_p
  );


  buf

  (
    g954_n_spl_,
    g954_n
  );


  buf

  (
    g954_n_spl_0,
    g954_n_spl_
  );


  buf

  (
    g954_p_spl_,
    g954_p
  );


  buf

  (
    g954_p_spl_0,
    g954_p_spl_
  );


  buf

  (
    g955_n_spl_,
    g955_n
  );


  buf

  (
    g948_n_spl_,
    g948_n
  );


  buf

  (
    g955_p_spl_,
    g955_p
  );


  buf

  (
    g948_p_spl_,
    g948_p
  );


  buf

  (
    g956_n_spl_,
    g956_n
  );


  buf

  (
    g956_n_spl_0,
    g956_n_spl_
  );


  buf

  (
    g956_p_spl_,
    g956_p
  );


  buf

  (
    g956_p_spl_0,
    g956_p_spl_
  );


  buf

  (
    g960_n_spl_,
    g960_n
  );


  buf

  (
    g959_n_spl_,
    g959_n
  );


  buf

  (
    g960_p_spl_,
    g960_p
  );


  buf

  (
    g959_p_spl_,
    g959_p
  );


  buf

  (
    g961_n_spl_,
    g961_n
  );


  buf

  (
    g961_n_spl_0,
    g961_n_spl_
  );


  buf

  (
    g961_p_spl_,
    g961_p
  );


  buf

  (
    g961_p_spl_0,
    g961_p_spl_
  );


  buf

  (
    n6075_o2_p_spl_,
    n6075_o2_p
  );


  buf

  (
    n6075_o2_p_spl_0,
    n6075_o2_p_spl_
  );


  buf

  (
    n6075_o2_n_spl_,
    n6075_o2_n
  );


  buf

  (
    n6075_o2_n_spl_0,
    n6075_o2_n_spl_
  );


  buf

  (
    n6075_o2_n_spl_1,
    n6075_o2_n_spl_
  );


  buf

  (
    g969_n_spl_,
    g969_n
  );


  buf

  (
    g968_n_spl_,
    g968_n
  );


  buf

  (
    g969_p_spl_,
    g969_p
  );


  buf

  (
    g968_p_spl_,
    g968_p
  );


  buf

  (
    g970_n_spl_,
    g970_n
  );


  buf

  (
    g970_n_spl_0,
    g970_n_spl_
  );


  buf

  (
    g970_p_spl_,
    g970_p
  );


  buf

  (
    g970_p_spl_0,
    g970_p_spl_
  );


  buf

  (
    g971_n_spl_,
    g971_n
  );


  buf

  (
    g967_n_spl_,
    g967_n
  );


  buf

  (
    g971_p_spl_,
    g971_p
  );


  buf

  (
    g967_p_spl_,
    g967_p
  );


  buf

  (
    g972_n_spl_,
    g972_n
  );


  buf

  (
    g972_n_spl_0,
    g972_n_spl_
  );


  buf

  (
    g972_p_spl_,
    g972_p
  );


  buf

  (
    g972_p_spl_0,
    g972_p_spl_
  );


  buf

  (
    g976_n_spl_,
    g976_n
  );


  buf

  (
    g975_n_spl_,
    g975_n
  );


  buf

  (
    g976_p_spl_,
    g976_p
  );


  buf

  (
    g975_p_spl_,
    g975_p
  );


  buf

  (
    g977_n_spl_,
    g977_n
  );


  buf

  (
    g977_n_spl_0,
    g977_n_spl_
  );


  buf

  (
    g977_p_spl_,
    g977_p
  );


  buf

  (
    g977_p_spl_0,
    g977_p_spl_
  );


  buf

  (
    g978_n_spl_,
    g978_n
  );


  buf

  (
    g964_n_spl_,
    g964_n
  );


  buf

  (
    g978_p_spl_,
    g978_p
  );


  buf

  (
    g964_p_spl_,
    g964_p
  );


  buf

  (
    g979_n_spl_,
    g979_n
  );


  buf

  (
    g979_n_spl_0,
    g979_n_spl_
  );


  buf

  (
    g979_p_spl_,
    g979_p
  );


  buf

  (
    g979_p_spl_0,
    g979_p_spl_
  );


  buf

  (
    g983_n_spl_,
    g983_n
  );


  buf

  (
    g982_n_spl_,
    g982_n
  );


  buf

  (
    g983_p_spl_,
    g983_p
  );


  buf

  (
    g982_p_spl_,
    g982_p
  );


  buf

  (
    g984_n_spl_,
    g984_n
  );


  buf

  (
    g984_n_spl_0,
    g984_n_spl_
  );


  buf

  (
    g984_p_spl_,
    g984_p
  );


  buf

  (
    g984_p_spl_0,
    g984_p_spl_
  );


  buf

  (
    G5064_o2_n_spl_,
    G5064_o2_n
  );


  buf

  (
    G5064_o2_n_spl_0,
    G5064_o2_n_spl_
  );


  buf

  (
    G5064_o2_p_spl_,
    G5064_o2_p
  );


  buf

  (
    G5064_o2_p_spl_0,
    G5064_o2_p_spl_
  );


  buf

  (
    g994_n_spl_,
    g994_n
  );


  buf

  (
    g993_n_spl_,
    g993_n
  );


  buf

  (
    g994_p_spl_,
    g994_p
  );


  buf

  (
    g993_p_spl_,
    g993_p
  );


  buf

  (
    g995_n_spl_,
    g995_n
  );


  buf

  (
    g995_n_spl_0,
    g995_n_spl_
  );


  buf

  (
    g995_p_spl_,
    g995_p
  );


  buf

  (
    g995_p_spl_0,
    g995_p_spl_
  );


  buf

  (
    n6103_o2_p_spl_,
    n6103_o2_p
  );


  buf

  (
    n6103_o2_p_spl_0,
    n6103_o2_p_spl_
  );


  buf

  (
    n6103_o2_n_spl_,
    n6103_o2_n
  );


  buf

  (
    n6103_o2_n_spl_0,
    n6103_o2_n_spl_
  );


  buf

  (
    g999_n_spl_,
    g999_n
  );


  buf

  (
    g998_n_spl_,
    g998_n
  );


  buf

  (
    g999_p_spl_,
    g999_p
  );


  buf

  (
    g998_p_spl_,
    g998_p
  );


  buf

  (
    g1000_n_spl_,
    g1000_n
  );


  buf

  (
    g1000_n_spl_0,
    g1000_n_spl_
  );


  buf

  (
    g1000_p_spl_,
    g1000_p
  );


  buf

  (
    g1000_p_spl_0,
    g1000_p_spl_
  );


  buf

  (
    g1001_n_spl_,
    g1001_n
  );


  buf

  (
    g990_n_spl_,
    g990_n
  );


  buf

  (
    g1001_p_spl_,
    g1001_p
  );


  buf

  (
    g990_p_spl_,
    g990_p
  );


  buf

  (
    g1002_n_spl_,
    g1002_n
  );


  buf

  (
    g1002_n_spl_0,
    g1002_n_spl_
  );


  buf

  (
    g1002_p_spl_,
    g1002_p
  );


  buf

  (
    g1002_p_spl_0,
    g1002_p_spl_
  );


  buf

  (
    g1006_n_spl_,
    g1006_n
  );


  buf

  (
    g1005_n_spl_,
    g1005_n
  );


  buf

  (
    g1006_p_spl_,
    g1006_p
  );


  buf

  (
    g1005_p_spl_,
    g1005_p
  );


  buf

  (
    g1007_n_spl_,
    g1007_n
  );


  buf

  (
    g1007_n_spl_0,
    g1007_n_spl_
  );


  buf

  (
    g1007_p_spl_,
    g1007_p
  );


  buf

  (
    g1007_p_spl_0,
    g1007_p_spl_
  );


  buf

  (
    g1008_n_spl_,
    g1008_n
  );


  buf

  (
    g987_n_spl_,
    g987_n
  );


  buf

  (
    g1008_p_spl_,
    g1008_p
  );


  buf

  (
    g987_p_spl_,
    g987_p
  );


  buf

  (
    G5247_o2_n_spl_,
    G5247_o2_n
  );


  buf

  (
    G5244_o2_n_spl_,
    G5244_o2_n
  );


  buf

  (
    G5247_o2_p_spl_,
    G5247_o2_p
  );


  buf

  (
    G5244_o2_p_spl_,
    G5244_o2_p
  );


  buf

  (
    g1010_n_spl_,
    g1010_n
  );


  buf

  (
    g1010_n_spl_0,
    g1010_n_spl_
  );


  buf

  (
    g1010_p_spl_,
    g1010_p
  );


  buf

  (
    g1010_p_spl_0,
    g1010_p_spl_
  );


  buf

  (
    n6205_o2_p_spl_,
    n6205_o2_p
  );


  buf

  (
    n6205_o2_p_spl_0,
    n6205_o2_p_spl_
  );


  buf

  (
    n6205_o2_n_spl_,
    n6205_o2_n
  );


  buf

  (
    n6205_o2_n_spl_0,
    n6205_o2_n_spl_
  );


  buf

  (
    g1014_n_spl_,
    g1014_n
  );


  buf

  (
    g1013_n_spl_,
    g1013_n
  );


  buf

  (
    g1014_p_spl_,
    g1014_p
  );


  buf

  (
    g1013_p_spl_,
    g1013_p
  );


  buf

  (
    g1015_n_spl_,
    g1015_n
  );


  buf

  (
    g1015_n_spl_0,
    g1015_n_spl_
  );


  buf

  (
    g1015_p_spl_,
    g1015_p
  );


  buf

  (
    g1015_p_spl_0,
    g1015_p_spl_
  );


  buf

  (
    g1019_n_spl_,
    g1019_n
  );


  buf

  (
    g1018_n_spl_,
    g1018_n
  );


  buf

  (
    g1019_p_spl_,
    g1019_p
  );


  buf

  (
    g1018_p_spl_,
    g1018_p
  );


  buf

  (
    g1020_n_spl_,
    g1020_n
  );


  buf

  (
    g1020_n_spl_0,
    g1020_n_spl_
  );


  buf

  (
    g1020_p_spl_,
    g1020_p
  );


  buf

  (
    g1020_p_spl_0,
    g1020_p_spl_
  );


  buf

  (
    g1024_n_spl_,
    g1024_n
  );


  buf

  (
    g1023_n_spl_,
    g1023_n
  );


  buf

  (
    g1024_p_spl_,
    g1024_p
  );


  buf

  (
    g1023_p_spl_,
    g1023_p
  );


  buf

  (
    g1025_n_spl_,
    g1025_n
  );


  buf

  (
    g1025_n_spl_0,
    g1025_n_spl_
  );


  buf

  (
    g1025_p_spl_,
    g1025_p
  );


  buf

  (
    g1025_p_spl_0,
    g1025_p_spl_
  );


  buf

  (
    g1029_n_spl_,
    g1029_n
  );


  buf

  (
    g1028_n_spl_,
    g1028_n
  );


  buf

  (
    g1029_p_spl_,
    g1029_p
  );


  buf

  (
    g1028_p_spl_,
    g1028_p
  );


  buf

  (
    g1030_n_spl_,
    g1030_n
  );


  buf

  (
    g1030_n_spl_0,
    g1030_n_spl_
  );


  buf

  (
    g1030_p_spl_,
    g1030_p
  );


  buf

  (
    g1030_p_spl_0,
    g1030_p_spl_
  );


  buf

  (
    g1034_n_spl_,
    g1034_n
  );


  buf

  (
    g1033_n_spl_,
    g1033_n
  );


  buf

  (
    g1034_p_spl_,
    g1034_p
  );


  buf

  (
    g1033_p_spl_,
    g1033_p
  );


  buf

  (
    g1035_n_spl_,
    g1035_n
  );


  buf

  (
    g1035_n_spl_0,
    g1035_n_spl_
  );


  buf

  (
    g1035_p_spl_,
    g1035_p
  );


  buf

  (
    g1035_p_spl_0,
    g1035_p_spl_
  );


  buf

  (
    g764_p_spl_,
    g764_p
  );


  buf

  (
    g1039_n_spl_,
    g1039_n
  );


  buf

  (
    g1038_n_spl_,
    g1038_n
  );


  buf

  (
    g1040_n_spl_,
    g1040_n
  );


  buf

  (
    g817_n_spl_,
    g817_n
  );


  buf

  (
    g804_p_spl_,
    g804_p
  );


  buf

  (
    n2797_lo_p_spl_,
    n2797_lo_p
  );


  buf

  (
    n2797_lo_p_spl_0,
    n2797_lo_p_spl_
  );


  buf

  (
    n2797_lo_p_spl_00,
    n2797_lo_p_spl_0
  );


  buf

  (
    n2797_lo_p_spl_000,
    n2797_lo_p_spl_00
  );


  buf

  (
    n2797_lo_p_spl_001,
    n2797_lo_p_spl_00
  );


  buf

  (
    n2797_lo_p_spl_01,
    n2797_lo_p_spl_0
  );


  buf

  (
    n2797_lo_p_spl_010,
    n2797_lo_p_spl_01
  );


  buf

  (
    n2797_lo_p_spl_011,
    n2797_lo_p_spl_01
  );


  buf

  (
    n2797_lo_p_spl_1,
    n2797_lo_p_spl_
  );


  buf

  (
    n2797_lo_p_spl_10,
    n2797_lo_p_spl_1
  );


  buf

  (
    n2797_lo_p_spl_100,
    n2797_lo_p_spl_10
  );


  buf

  (
    n2797_lo_p_spl_101,
    n2797_lo_p_spl_10
  );


  buf

  (
    n2797_lo_p_spl_11,
    n2797_lo_p_spl_1
  );


  buf

  (
    n2797_lo_n_spl_,
    n2797_lo_n
  );


  buf

  (
    n2797_lo_n_spl_0,
    n2797_lo_n_spl_
  );


  buf

  (
    n2797_lo_n_spl_00,
    n2797_lo_n_spl_0
  );


  buf

  (
    n2797_lo_n_spl_000,
    n2797_lo_n_spl_00
  );


  buf

  (
    n2797_lo_n_spl_001,
    n2797_lo_n_spl_00
  );


  buf

  (
    n2797_lo_n_spl_01,
    n2797_lo_n_spl_0
  );


  buf

  (
    n2797_lo_n_spl_010,
    n2797_lo_n_spl_01
  );


  buf

  (
    n2797_lo_n_spl_011,
    n2797_lo_n_spl_01
  );


  buf

  (
    n2797_lo_n_spl_1,
    n2797_lo_n_spl_
  );


  buf

  (
    n2797_lo_n_spl_10,
    n2797_lo_n_spl_1
  );


  buf

  (
    n2797_lo_n_spl_100,
    n2797_lo_n_spl_10
  );


  buf

  (
    n2797_lo_n_spl_101,
    n2797_lo_n_spl_10
  );


  buf

  (
    n2797_lo_n_spl_11,
    n2797_lo_n_spl_1
  );


  buf

  (
    G3422_o2_n_spl_,
    G3422_o2_n
  );


  buf

  (
    G3422_o2_n_spl_0,
    G3422_o2_n_spl_
  );


  buf

  (
    G3422_o2_p_spl_,
    G3422_o2_p
  );


  buf

  (
    G3422_o2_p_spl_0,
    G3422_o2_p_spl_
  );


  buf

  (
    g1049_n_spl_,
    g1049_n
  );


  buf

  (
    g1048_n_spl_,
    g1048_n
  );


  buf

  (
    g1049_p_spl_,
    g1049_p
  );


  buf

  (
    g1048_p_spl_,
    g1048_p
  );


  buf

  (
    g1050_n_spl_,
    g1050_n
  );


  buf

  (
    g1050_n_spl_0,
    g1050_n_spl_
  );


  buf

  (
    g1050_p_spl_,
    g1050_p
  );


  buf

  (
    g1050_p_spl_0,
    g1050_p_spl_
  );


  buf

  (
    n7835_o2_p_spl_,
    n7835_o2_p
  );


  buf

  (
    n7835_o2_p_spl_0,
    n7835_o2_p_spl_
  );


  buf

  (
    n7835_o2_p_spl_00,
    n7835_o2_p_spl_0
  );


  buf

  (
    n7835_o2_p_spl_1,
    n7835_o2_p_spl_
  );


  buf

  (
    n7835_o2_n_spl_,
    n7835_o2_n
  );


  buf

  (
    n7835_o2_n_spl_0,
    n7835_o2_n_spl_
  );


  buf

  (
    n7835_o2_n_spl_00,
    n7835_o2_n_spl_0
  );


  buf

  (
    n7835_o2_n_spl_1,
    n7835_o2_n_spl_
  );


  buf

  (
    g1054_n_spl_,
    g1054_n
  );


  buf

  (
    g1053_n_spl_,
    g1053_n
  );


  buf

  (
    g1054_p_spl_,
    g1054_p
  );


  buf

  (
    g1053_p_spl_,
    g1053_p
  );


  buf

  (
    g1055_n_spl_,
    g1055_n
  );


  buf

  (
    g1055_n_spl_0,
    g1055_n_spl_
  );


  buf

  (
    g1055_p_spl_,
    g1055_p
  );


  buf

  (
    g1055_p_spl_0,
    g1055_p_spl_
  );


  buf

  (
    g1059_n_spl_,
    g1059_n
  );


  buf

  (
    g1058_n_spl_,
    g1058_n
  );


  buf

  (
    g1059_p_spl_,
    g1059_p
  );


  buf

  (
    g1058_p_spl_,
    g1058_p
  );


  buf

  (
    g1060_n_spl_,
    g1060_n
  );


  buf

  (
    g1060_n_spl_0,
    g1060_n_spl_
  );


  buf

  (
    g1060_p_spl_,
    g1060_p
  );


  buf

  (
    g1060_p_spl_0,
    g1060_p_spl_
  );


  buf

  (
    g1064_n_spl_,
    g1064_n
  );


  buf

  (
    g1063_n_spl_,
    g1063_n
  );


  buf

  (
    g1064_p_spl_,
    g1064_p
  );


  buf

  (
    g1063_p_spl_,
    g1063_p
  );


  buf

  (
    g1065_n_spl_,
    g1065_n
  );


  buf

  (
    g1065_n_spl_0,
    g1065_n_spl_
  );


  buf

  (
    g1065_p_spl_,
    g1065_p
  );


  buf

  (
    g1065_p_spl_0,
    g1065_p_spl_
  );


  buf

  (
    g803_p_spl_,
    g803_p
  );


  buf

  (
    g1069_n_spl_,
    g1069_n
  );


  buf

  (
    g1068_n_spl_,
    g1068_n
  );


  buf

  (
    g1069_p_spl_,
    g1069_p
  );


  buf

  (
    g1068_p_spl_,
    g1068_p
  );


  buf

  (
    g1070_n_spl_,
    g1070_n
  );


  buf

  (
    g1070_n_spl_0,
    g1070_n_spl_
  );


  buf

  (
    g1070_p_spl_,
    g1070_p
  );


  buf

  (
    g1070_p_spl_0,
    g1070_p_spl_
  );


  buf

  (
    n2728_lo_buf_o2_p_spl_,
    n2728_lo_buf_o2_p
  );


  buf

  (
    n2728_lo_buf_o2_p_spl_0,
    n2728_lo_buf_o2_p_spl_
  );


  buf

  (
    n2728_lo_buf_o2_p_spl_00,
    n2728_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2728_lo_buf_o2_p_spl_000,
    n2728_lo_buf_o2_p_spl_00
  );


  buf

  (
    n2728_lo_buf_o2_p_spl_001,
    n2728_lo_buf_o2_p_spl_00
  );


  buf

  (
    n2728_lo_buf_o2_p_spl_01,
    n2728_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2728_lo_buf_o2_p_spl_010,
    n2728_lo_buf_o2_p_spl_01
  );


  buf

  (
    n2728_lo_buf_o2_p_spl_011,
    n2728_lo_buf_o2_p_spl_01
  );


  buf

  (
    n2728_lo_buf_o2_p_spl_1,
    n2728_lo_buf_o2_p_spl_
  );


  buf

  (
    n2728_lo_buf_o2_p_spl_10,
    n2728_lo_buf_o2_p_spl_1
  );


  buf

  (
    n2728_lo_buf_o2_p_spl_100,
    n2728_lo_buf_o2_p_spl_10
  );


  buf

  (
    n2728_lo_buf_o2_p_spl_101,
    n2728_lo_buf_o2_p_spl_10
  );


  buf

  (
    n2728_lo_buf_o2_p_spl_11,
    n2728_lo_buf_o2_p_spl_1
  );


  buf

  (
    n2728_lo_buf_o2_p_spl_110,
    n2728_lo_buf_o2_p_spl_11
  );


  buf

  (
    n2728_lo_buf_o2_p_spl_111,
    n2728_lo_buf_o2_p_spl_11
  );


  buf

  (
    n2728_lo_buf_o2_n_spl_,
    n2728_lo_buf_o2_n
  );


  buf

  (
    n2728_lo_buf_o2_n_spl_0,
    n2728_lo_buf_o2_n_spl_
  );


  buf

  (
    n2728_lo_buf_o2_n_spl_00,
    n2728_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2728_lo_buf_o2_n_spl_000,
    n2728_lo_buf_o2_n_spl_00
  );


  buf

  (
    n2728_lo_buf_o2_n_spl_001,
    n2728_lo_buf_o2_n_spl_00
  );


  buf

  (
    n2728_lo_buf_o2_n_spl_01,
    n2728_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2728_lo_buf_o2_n_spl_010,
    n2728_lo_buf_o2_n_spl_01
  );


  buf

  (
    n2728_lo_buf_o2_n_spl_011,
    n2728_lo_buf_o2_n_spl_01
  );


  buf

  (
    n2728_lo_buf_o2_n_spl_1,
    n2728_lo_buf_o2_n_spl_
  );


  buf

  (
    n2728_lo_buf_o2_n_spl_10,
    n2728_lo_buf_o2_n_spl_1
  );


  buf

  (
    n2728_lo_buf_o2_n_spl_100,
    n2728_lo_buf_o2_n_spl_10
  );


  buf

  (
    n2728_lo_buf_o2_n_spl_101,
    n2728_lo_buf_o2_n_spl_10
  );


  buf

  (
    n2728_lo_buf_o2_n_spl_11,
    n2728_lo_buf_o2_n_spl_1
  );


  buf

  (
    n2728_lo_buf_o2_n_spl_110,
    n2728_lo_buf_o2_n_spl_11
  );


  buf

  (
    n2728_lo_buf_o2_n_spl_111,
    n2728_lo_buf_o2_n_spl_11
  );


  buf

  (
    g1073_n_spl_,
    g1073_n
  );


  buf

  (
    g1045_p_spl_,
    g1045_p
  );


  buf

  (
    n2512_lo_buf_o2_p_spl_,
    n2512_lo_buf_o2_p
  );


  buf

  (
    n2512_lo_buf_o2_p_spl_0,
    n2512_lo_buf_o2_p_spl_
  );


  buf

  (
    n2512_lo_buf_o2_p_spl_00,
    n2512_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2512_lo_buf_o2_p_spl_01,
    n2512_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2512_lo_buf_o2_p_spl_1,
    n2512_lo_buf_o2_p_spl_
  );


  buf

  (
    n2512_lo_buf_o2_p_spl_10,
    n2512_lo_buf_o2_p_spl_1
  );


  buf

  (
    n2512_lo_buf_o2_n_spl_,
    n2512_lo_buf_o2_n
  );


  buf

  (
    n2512_lo_buf_o2_n_spl_0,
    n2512_lo_buf_o2_n_spl_
  );


  buf

  (
    n2512_lo_buf_o2_n_spl_00,
    n2512_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2512_lo_buf_o2_n_spl_1,
    n2512_lo_buf_o2_n_spl_
  );


  buf

  (
    g1077_n_spl_,
    g1077_n
  );


  buf

  (
    g1076_n_spl_,
    g1076_n
  );


  buf

  (
    g1077_p_spl_,
    g1077_p
  );


  buf

  (
    g1076_p_spl_,
    g1076_p
  );


  buf

  (
    g1078_n_spl_,
    g1078_n
  );


  buf

  (
    g1078_n_spl_0,
    g1078_n_spl_
  );


  buf

  (
    g1078_p_spl_,
    g1078_p
  );


  buf

  (
    g1078_p_spl_0,
    g1078_p_spl_
  );


  buf

  (
    g1082_n_spl_,
    g1082_n
  );


  buf

  (
    g1081_n_spl_,
    g1081_n
  );


  buf

  (
    g1082_p_spl_,
    g1082_p
  );


  buf

  (
    g1081_p_spl_,
    g1081_p
  );


  buf

  (
    g1083_n_spl_,
    g1083_n
  );


  buf

  (
    g1083_n_spl_0,
    g1083_n_spl_
  );


  buf

  (
    g1083_p_spl_,
    g1083_p
  );


  buf

  (
    g1083_p_spl_0,
    g1083_p_spl_
  );


  buf

  (
    g1087_n_spl_,
    g1087_n
  );


  buf

  (
    g1086_n_spl_,
    g1086_n
  );


  buf

  (
    g1087_p_spl_,
    g1087_p
  );


  buf

  (
    g1086_p_spl_,
    g1086_p
  );


  buf

  (
    g1088_n_spl_,
    g1088_n
  );


  buf

  (
    g1088_n_spl_0,
    g1088_n_spl_
  );


  buf

  (
    g1088_p_spl_,
    g1088_p
  );


  buf

  (
    g1088_p_spl_0,
    g1088_p_spl_
  );


  buf

  (
    g1044_p_spl_,
    g1044_p
  );


  buf

  (
    g1092_n_spl_,
    g1092_n
  );


  buf

  (
    g1091_n_spl_,
    g1091_n
  );


  buf

  (
    g1092_p_spl_,
    g1092_p
  );


  buf

  (
    g1091_p_spl_,
    g1091_p
  );


  buf

  (
    g1093_n_spl_,
    g1093_n
  );


  buf

  (
    g1093_n_spl_0,
    g1093_n_spl_
  );


  buf

  (
    g1093_p_spl_,
    g1093_p
  );


  buf

  (
    g1093_p_spl_0,
    g1093_p_spl_
  );


  buf

  (
    g1096_n_spl_,
    g1096_n
  );


  buf

  (
    g1074_p_spl_,
    g1074_p
  );


  buf

  (
    g1043_n_spl_,
    g1043_n
  );


  buf

  (
    g1043_n_spl_0,
    g1043_n_spl_
  );


  buf

  (
    g1105_n_spl_,
    g1105_n
  );


  buf

  (
    g1104_n_spl_,
    g1104_n
  );


  buf

  (
    g1105_p_spl_,
    g1105_p
  );


  buf

  (
    g1104_p_spl_,
    g1104_p
  );


  buf

  (
    g1106_n_spl_,
    g1106_n
  );


  buf

  (
    g1106_n_spl_0,
    g1106_n_spl_
  );


  buf

  (
    g1106_p_spl_,
    g1106_p
  );


  buf

  (
    g1106_p_spl_0,
    g1106_p_spl_
  );


  buf

  (
    g1110_n_spl_,
    g1110_n
  );


  buf

  (
    g1109_n_spl_,
    g1109_n
  );


  buf

  (
    g1110_p_spl_,
    g1110_p
  );


  buf

  (
    g1109_p_spl_,
    g1109_p
  );


  buf

  (
    g1111_n_spl_,
    g1111_n
  );


  buf

  (
    g1111_n_spl_0,
    g1111_n_spl_
  );


  buf

  (
    g1111_p_spl_,
    g1111_p
  );


  buf

  (
    g1111_p_spl_0,
    g1111_p_spl_
  );


  buf

  (
    g1115_n_spl_,
    g1115_n
  );


  buf

  (
    g1114_n_spl_,
    g1114_n
  );


  buf

  (
    g1115_p_spl_,
    g1115_p
  );


  buf

  (
    g1114_p_spl_,
    g1114_p
  );


  buf

  (
    g1116_n_spl_,
    g1116_n
  );


  buf

  (
    g1116_n_spl_0,
    g1116_n_spl_
  );


  buf

  (
    g1116_p_spl_,
    g1116_p
  );


  buf

  (
    g1116_p_spl_0,
    g1116_p_spl_
  );


  buf

  (
    g1120_n_spl_,
    g1120_n
  );


  buf

  (
    g1119_n_spl_,
    g1119_n
  );


  buf

  (
    g1120_p_spl_,
    g1120_p
  );


  buf

  (
    g1119_p_spl_,
    g1119_p
  );


  buf

  (
    g1121_n_spl_,
    g1121_n
  );


  buf

  (
    g1121_n_spl_0,
    g1121_n_spl_
  );


  buf

  (
    g1121_p_spl_,
    g1121_p
  );


  buf

  (
    g1121_p_spl_0,
    g1121_p_spl_
  );


  buf

  (
    g1130_n_spl_,
    g1130_n
  );


  buf

  (
    g1129_n_spl_,
    g1129_n
  );


  buf

  (
    g1130_p_spl_,
    g1130_p
  );


  buf

  (
    g1129_p_spl_,
    g1129_p
  );


  buf

  (
    g1131_n_spl_,
    g1131_n
  );


  buf

  (
    g1131_n_spl_0,
    g1131_n_spl_
  );


  buf

  (
    g1131_p_spl_,
    g1131_p
  );


  buf

  (
    g1131_p_spl_0,
    g1131_p_spl_
  );


  buf

  (
    g1135_n_spl_,
    g1135_n
  );


  buf

  (
    g1134_n_spl_,
    g1134_n
  );


  buf

  (
    g1135_p_spl_,
    g1135_p
  );


  buf

  (
    g1134_p_spl_,
    g1134_p
  );


  buf

  (
    g1136_n_spl_,
    g1136_n
  );


  buf

  (
    g1136_n_spl_0,
    g1136_n_spl_
  );


  buf

  (
    g1136_p_spl_,
    g1136_p
  );


  buf

  (
    g1136_p_spl_0,
    g1136_p_spl_
  );


  buf

  (
    g1140_n_spl_,
    g1140_n
  );


  buf

  (
    g1139_n_spl_,
    g1139_n
  );


  buf

  (
    g1140_p_spl_,
    g1140_p
  );


  buf

  (
    g1139_p_spl_,
    g1139_p
  );


  buf

  (
    g1141_n_spl_,
    g1141_n
  );


  buf

  (
    g1141_n_spl_0,
    g1141_n_spl_
  );


  buf

  (
    g1141_p_spl_,
    g1141_p
  );


  buf

  (
    g1141_p_spl_0,
    g1141_p_spl_
  );


  buf

  (
    g1145_n_spl_,
    g1145_n
  );


  buf

  (
    g1144_n_spl_,
    g1144_n
  );


  buf

  (
    g1145_p_spl_,
    g1145_p
  );


  buf

  (
    g1144_p_spl_,
    g1144_p
  );


  buf

  (
    g1146_n_spl_,
    g1146_n
  );


  buf

  (
    g1146_n_spl_0,
    g1146_n_spl_
  );


  buf

  (
    g1146_p_spl_,
    g1146_p
  );


  buf

  (
    g1146_p_spl_0,
    g1146_p_spl_
  );


  buf

  (
    g1158_n_spl_,
    g1158_n
  );


  buf

  (
    g1157_n_spl_,
    g1157_n
  );


  buf

  (
    g1158_p_spl_,
    g1158_p
  );


  buf

  (
    g1157_p_spl_,
    g1157_p
  );


  buf

  (
    g1159_n_spl_,
    g1159_n
  );


  buf

  (
    g1159_n_spl_0,
    g1159_n_spl_
  );


  buf

  (
    g1159_p_spl_,
    g1159_p
  );


  buf

  (
    g1159_p_spl_0,
    g1159_p_spl_
  );


  buf

  (
    n6169_o2_p_spl_,
    n6169_o2_p
  );


  buf

  (
    n6169_o2_p_spl_0,
    n6169_o2_p_spl_
  );


  buf

  (
    n6169_o2_n_spl_,
    n6169_o2_n
  );


  buf

  (
    n6169_o2_n_spl_0,
    n6169_o2_n_spl_
  );


  buf

  (
    g1163_n_spl_,
    g1163_n
  );


  buf

  (
    g1162_n_spl_,
    g1162_n
  );


  buf

  (
    g1163_p_spl_,
    g1163_p
  );


  buf

  (
    g1162_p_spl_,
    g1162_p
  );


  buf

  (
    g1164_n_spl_,
    g1164_n
  );


  buf

  (
    g1164_n_spl_0,
    g1164_n_spl_
  );


  buf

  (
    g1164_p_spl_,
    g1164_p
  );


  buf

  (
    g1164_p_spl_0,
    g1164_p_spl_
  );


  buf

  (
    g1165_n_spl_,
    g1165_n
  );


  buf

  (
    g1154_n_spl_,
    g1154_n
  );


  buf

  (
    g1165_p_spl_,
    g1165_p
  );


  buf

  (
    g1154_p_spl_,
    g1154_p
  );


  buf

  (
    g1166_n_spl_,
    g1166_n
  );


  buf

  (
    g1166_n_spl_0,
    g1166_n_spl_
  );


  buf

  (
    g1166_p_spl_,
    g1166_p
  );


  buf

  (
    g1166_p_spl_0,
    g1166_p_spl_
  );


  buf

  (
    g1170_n_spl_,
    g1170_n
  );


  buf

  (
    g1169_n_spl_,
    g1169_n
  );


  buf

  (
    g1170_p_spl_,
    g1170_p
  );


  buf

  (
    g1169_p_spl_,
    g1169_p
  );


  buf

  (
    g1171_n_spl_,
    g1171_n
  );


  buf

  (
    g1171_n_spl_0,
    g1171_n_spl_
  );


  buf

  (
    g1171_p_spl_,
    g1171_p
  );


  buf

  (
    g1171_p_spl_0,
    g1171_p_spl_
  );


  buf

  (
    g1178_n_spl_,
    g1178_n
  );


  buf

  (
    g1177_n_spl_,
    g1177_n
  );


  buf

  (
    g1178_p_spl_,
    g1178_p
  );


  buf

  (
    g1177_p_spl_,
    g1177_p
  );


  buf

  (
    g1179_n_spl_,
    g1179_n
  );


  buf

  (
    g1179_n_spl_0,
    g1179_n_spl_
  );


  buf

  (
    g1179_p_spl_,
    g1179_p
  );


  buf

  (
    g1179_p_spl_0,
    g1179_p_spl_
  );


  buf

  (
    g1183_n_spl_,
    g1183_n
  );


  buf

  (
    g1182_n_spl_,
    g1182_n
  );


  buf

  (
    g1183_p_spl_,
    g1183_p
  );


  buf

  (
    g1182_p_spl_,
    g1182_p
  );


  buf

  (
    g1184_n_spl_,
    g1184_n
  );


  buf

  (
    g1184_n_spl_0,
    g1184_n_spl_
  );


  buf

  (
    g1184_p_spl_,
    g1184_p
  );


  buf

  (
    g1184_p_spl_0,
    g1184_p_spl_
  );


  buf

  (
    g1185_n_spl_,
    g1185_n
  );


  buf

  (
    g1174_n_spl_,
    g1174_n
  );


  buf

  (
    g1185_p_spl_,
    g1185_p
  );


  buf

  (
    g1174_p_spl_,
    g1174_p
  );


  buf

  (
    g1186_n_spl_,
    g1186_n
  );


  buf

  (
    g1186_n_spl_0,
    g1186_n_spl_
  );


  buf

  (
    g1186_p_spl_,
    g1186_p
  );


  buf

  (
    g1186_p_spl_0,
    g1186_p_spl_
  );


  buf

  (
    g1190_n_spl_,
    g1190_n
  );


  buf

  (
    g1189_n_spl_,
    g1189_n
  );


  buf

  (
    g1190_p_spl_,
    g1190_p
  );


  buf

  (
    g1189_p_spl_,
    g1189_p
  );


  buf

  (
    g1191_n_spl_,
    g1191_n
  );


  buf

  (
    g1191_n_spl_0,
    g1191_n_spl_
  );


  buf

  (
    g1191_p_spl_,
    g1191_p
  );


  buf

  (
    g1191_p_spl_0,
    g1191_p_spl_
  );


  buf

  (
    g1198_n_spl_,
    g1198_n
  );


  buf

  (
    g1197_n_spl_,
    g1197_n
  );


  buf

  (
    g1198_p_spl_,
    g1198_p
  );


  buf

  (
    g1197_p_spl_,
    g1197_p
  );


  buf

  (
    g1199_n_spl_,
    g1199_n
  );


  buf

  (
    g1199_n_spl_0,
    g1199_n_spl_
  );


  buf

  (
    g1199_p_spl_,
    g1199_p
  );


  buf

  (
    g1199_p_spl_0,
    g1199_p_spl_
  );


  buf

  (
    g1203_n_spl_,
    g1203_n
  );


  buf

  (
    g1202_n_spl_,
    g1202_n
  );


  buf

  (
    g1203_p_spl_,
    g1203_p
  );


  buf

  (
    g1202_p_spl_,
    g1202_p
  );


  buf

  (
    g1204_n_spl_,
    g1204_n
  );


  buf

  (
    g1204_n_spl_0,
    g1204_n_spl_
  );


  buf

  (
    g1204_p_spl_,
    g1204_p
  );


  buf

  (
    g1204_p_spl_0,
    g1204_p_spl_
  );


  buf

  (
    g1210_n_spl_,
    g1210_n
  );


  buf

  (
    g1209_n_spl_,
    g1209_n
  );


  buf

  (
    g1211_n_spl_,
    g1211_n
  );


  buf

  (
    n2734_lo_p_spl_,
    n2734_lo_p
  );


  buf

  (
    n2734_lo_p_spl_0,
    n2734_lo_p_spl_
  );


  buf

  (
    n2734_lo_p_spl_00,
    n2734_lo_p_spl_0
  );


  buf

  (
    n2734_lo_p_spl_000,
    n2734_lo_p_spl_00
  );


  buf

  (
    n2734_lo_p_spl_001,
    n2734_lo_p_spl_00
  );


  buf

  (
    n2734_lo_p_spl_01,
    n2734_lo_p_spl_0
  );


  buf

  (
    n2734_lo_p_spl_010,
    n2734_lo_p_spl_01
  );


  buf

  (
    n2734_lo_p_spl_011,
    n2734_lo_p_spl_01
  );


  buf

  (
    n2734_lo_p_spl_1,
    n2734_lo_p_spl_
  );


  buf

  (
    n2734_lo_p_spl_10,
    n2734_lo_p_spl_1
  );


  buf

  (
    n2734_lo_p_spl_100,
    n2734_lo_p_spl_10
  );


  buf

  (
    n2734_lo_p_spl_101,
    n2734_lo_p_spl_10
  );


  buf

  (
    n2734_lo_p_spl_11,
    n2734_lo_p_spl_1
  );


  buf

  (
    n2734_lo_p_spl_110,
    n2734_lo_p_spl_11
  );


  buf

  (
    n2734_lo_p_spl_111,
    n2734_lo_p_spl_11
  );


  buf

  (
    n2734_lo_n_spl_,
    n2734_lo_n
  );


  buf

  (
    n2734_lo_n_spl_0,
    n2734_lo_n_spl_
  );


  buf

  (
    n2734_lo_n_spl_00,
    n2734_lo_n_spl_0
  );


  buf

  (
    n2734_lo_n_spl_000,
    n2734_lo_n_spl_00
  );


  buf

  (
    n2734_lo_n_spl_001,
    n2734_lo_n_spl_00
  );


  buf

  (
    n2734_lo_n_spl_01,
    n2734_lo_n_spl_0
  );


  buf

  (
    n2734_lo_n_spl_010,
    n2734_lo_n_spl_01
  );


  buf

  (
    n2734_lo_n_spl_011,
    n2734_lo_n_spl_01
  );


  buf

  (
    n2734_lo_n_spl_1,
    n2734_lo_n_spl_
  );


  buf

  (
    n2734_lo_n_spl_10,
    n2734_lo_n_spl_1
  );


  buf

  (
    n2734_lo_n_spl_100,
    n2734_lo_n_spl_10
  );


  buf

  (
    n2734_lo_n_spl_101,
    n2734_lo_n_spl_10
  );


  buf

  (
    n2734_lo_n_spl_11,
    n2734_lo_n_spl_1
  );


  buf

  (
    n2734_lo_n_spl_110,
    n2734_lo_n_spl_11
  );


  buf

  (
    n2734_lo_n_spl_111,
    n2734_lo_n_spl_11
  );


  buf

  (
    g1009_n_spl_,
    g1009_n
  );


  buf

  (
    g1009_n_spl_0,
    g1009_n_spl_
  );


  buf

  (
    g1009_p_spl_,
    g1009_p
  );


  buf

  (
    g935_n_spl_,
    g935_n
  );


  buf

  (
    g935_n_spl_0,
    g935_n_spl_
  );


  buf

  (
    g935_p_spl_,
    g935_p
  );


  buf

  (
    g861_n_spl_,
    g861_n
  );


  buf

  (
    g861_n_spl_0,
    g861_n_spl_
  );


  buf

  (
    g861_p_spl_,
    g861_p
  );


  buf

  (
    g1214_n_spl_,
    g1214_n
  );


  buf

  (
    g1098_n_spl_,
    g1098_n
  );


  buf

  (
    n7148_o2_p_spl_,
    n7148_o2_p
  );


  buf

  (
    n7148_o2_p_spl_0,
    n7148_o2_p_spl_
  );


  buf

  (
    n7148_o2_p_spl_1,
    n7148_o2_p_spl_
  );


  buf

  (
    n7148_o2_n_spl_,
    n7148_o2_n
  );


  buf

  (
    n7148_o2_n_spl_0,
    n7148_o2_n_spl_
  );


  buf

  (
    G2917_o2_n_spl_,
    G2917_o2_n
  );


  buf

  (
    G1280_o2_n_spl_,
    G1280_o2_n
  );


  buf

  (
    G2917_o2_p_spl_,
    G2917_o2_p
  );


  buf

  (
    G1280_o2_p_spl_,
    G1280_o2_p
  );


  buf

  (
    g1233_n_spl_,
    g1233_n
  );


  buf

  (
    g1233_n_spl_0,
    g1233_n_spl_
  );


  buf

  (
    g1233_p_spl_,
    g1233_p
  );


  buf

  (
    g1233_p_spl_0,
    g1233_p_spl_
  );


  buf

  (
    n7224_o2_p_spl_,
    n7224_o2_p
  );


  buf

  (
    n7224_o2_p_spl_0,
    n7224_o2_p_spl_
  );


  buf

  (
    n7224_o2_p_spl_1,
    n7224_o2_p_spl_
  );


  buf

  (
    n7224_o2_n_spl_,
    n7224_o2_n
  );


  buf

  (
    n7224_o2_n_spl_0,
    n7224_o2_n_spl_
  );


  buf

  (
    g1237_n_spl_,
    g1237_n
  );


  buf

  (
    g1236_n_spl_,
    g1236_n
  );


  buf

  (
    g1237_p_spl_,
    g1237_p
  );


  buf

  (
    g1236_p_spl_,
    g1236_p
  );


  buf

  (
    g1238_n_spl_,
    g1238_n
  );


  buf

  (
    g1238_n_spl_0,
    g1238_n_spl_
  );


  buf

  (
    g1238_p_spl_,
    g1238_p
  );


  buf

  (
    g1238_p_spl_0,
    g1238_p_spl_
  );


  buf

  (
    g1239_n_spl_,
    g1239_n
  );


  buf

  (
    g1232_n_spl_,
    g1232_n
  );


  buf

  (
    g1239_p_spl_,
    g1239_p
  );


  buf

  (
    g1232_p_spl_,
    g1232_p
  );


  buf

  (
    g1240_n_spl_,
    g1240_n
  );


  buf

  (
    g1240_n_spl_0,
    g1240_n_spl_
  );


  buf

  (
    g1240_p_spl_,
    g1240_p
  );


  buf

  (
    g1240_p_spl_0,
    g1240_p_spl_
  );


  buf

  (
    g1244_n_spl_,
    g1244_n
  );


  buf

  (
    g1243_n_spl_,
    g1243_n
  );


  buf

  (
    g1244_p_spl_,
    g1244_p
  );


  buf

  (
    g1243_p_spl_,
    g1243_p
  );


  buf

  (
    g1245_n_spl_,
    g1245_n
  );


  buf

  (
    g1245_n_spl_0,
    g1245_n_spl_
  );


  buf

  (
    g1245_p_spl_,
    g1245_p
  );


  buf

  (
    g1245_p_spl_0,
    g1245_p_spl_
  );


  buf

  (
    n7280_o2_p_spl_,
    n7280_o2_p
  );


  buf

  (
    n7280_o2_p_spl_0,
    n7280_o2_p_spl_
  );


  buf

  (
    n7280_o2_p_spl_1,
    n7280_o2_p_spl_
  );


  buf

  (
    n7280_o2_n_spl_,
    n7280_o2_n
  );


  buf

  (
    n7280_o2_n_spl_0,
    n7280_o2_n_spl_
  );


  buf

  (
    n7280_o2_n_spl_1,
    n7280_o2_n_spl_
  );


  buf

  (
    g1253_n_spl_,
    g1253_n
  );


  buf

  (
    g1252_n_spl_,
    g1252_n
  );


  buf

  (
    g1253_p_spl_,
    g1253_p
  );


  buf

  (
    g1252_p_spl_,
    g1252_p
  );


  buf

  (
    g1254_n_spl_,
    g1254_n
  );


  buf

  (
    g1254_n_spl_0,
    g1254_n_spl_
  );


  buf

  (
    g1254_p_spl_,
    g1254_p
  );


  buf

  (
    g1254_p_spl_0,
    g1254_p_spl_
  );


  buf

  (
    g1255_n_spl_,
    g1255_n
  );


  buf

  (
    g1251_n_spl_,
    g1251_n
  );


  buf

  (
    g1255_p_spl_,
    g1255_p
  );


  buf

  (
    g1251_p_spl_,
    g1251_p
  );


  buf

  (
    g1256_n_spl_,
    g1256_n
  );


  buf

  (
    g1256_n_spl_0,
    g1256_n_spl_
  );


  buf

  (
    g1256_p_spl_,
    g1256_p
  );


  buf

  (
    g1256_p_spl_0,
    g1256_p_spl_
  );


  buf

  (
    g1260_n_spl_,
    g1260_n
  );


  buf

  (
    g1259_n_spl_,
    g1259_n
  );


  buf

  (
    g1260_p_spl_,
    g1260_p
  );


  buf

  (
    g1259_p_spl_,
    g1259_p
  );


  buf

  (
    g1261_n_spl_,
    g1261_n
  );


  buf

  (
    g1261_n_spl_0,
    g1261_n_spl_
  );


  buf

  (
    g1261_p_spl_,
    g1261_p
  );


  buf

  (
    g1261_p_spl_0,
    g1261_p_spl_
  );


  buf

  (
    g1262_n_spl_,
    g1262_n
  );


  buf

  (
    g1248_n_spl_,
    g1248_n
  );


  buf

  (
    g1262_p_spl_,
    g1262_p
  );


  buf

  (
    g1248_p_spl_,
    g1248_p
  );


  buf

  (
    g1263_n_spl_,
    g1263_n
  );


  buf

  (
    g1263_n_spl_0,
    g1263_n_spl_
  );


  buf

  (
    g1263_p_spl_,
    g1263_p
  );


  buf

  (
    g1263_p_spl_0,
    g1263_p_spl_
  );


  buf

  (
    g1267_n_spl_,
    g1267_n
  );


  buf

  (
    g1266_n_spl_,
    g1266_n
  );


  buf

  (
    g1267_p_spl_,
    g1267_p
  );


  buf

  (
    g1266_p_spl_,
    g1266_p
  );


  buf

  (
    g1268_n_spl_,
    g1268_n
  );


  buf

  (
    g1268_n_spl_0,
    g1268_n_spl_
  );


  buf

  (
    g1268_p_spl_,
    g1268_p
  );


  buf

  (
    g1268_p_spl_0,
    g1268_p_spl_
  );


  buf

  (
    G3241_o2_n_spl_,
    G3241_o2_n
  );


  buf

  (
    G3241_o2_n_spl_0,
    G3241_o2_n_spl_
  );


  buf

  (
    G3241_o2_p_spl_,
    G3241_o2_p
  );


  buf

  (
    G3241_o2_p_spl_0,
    G3241_o2_p_spl_
  );


  buf

  (
    g1278_n_spl_,
    g1278_n
  );


  buf

  (
    g1277_n_spl_,
    g1277_n
  );


  buf

  (
    g1278_p_spl_,
    g1278_p
  );


  buf

  (
    g1277_p_spl_,
    g1277_p
  );


  buf

  (
    g1279_n_spl_,
    g1279_n
  );


  buf

  (
    g1279_n_spl_0,
    g1279_n_spl_
  );


  buf

  (
    g1279_p_spl_,
    g1279_p
  );


  buf

  (
    g1279_p_spl_0,
    g1279_p_spl_
  );


  buf

  (
    n7313_o2_p_spl_,
    n7313_o2_p
  );


  buf

  (
    n7313_o2_p_spl_0,
    n7313_o2_p_spl_
  );


  buf

  (
    n7313_o2_p_spl_1,
    n7313_o2_p_spl_
  );


  buf

  (
    n7313_o2_n_spl_,
    n7313_o2_n
  );


  buf

  (
    n7313_o2_n_spl_0,
    n7313_o2_n_spl_
  );


  buf

  (
    g1283_n_spl_,
    g1283_n
  );


  buf

  (
    g1282_n_spl_,
    g1282_n
  );


  buf

  (
    g1283_p_spl_,
    g1283_p
  );


  buf

  (
    g1282_p_spl_,
    g1282_p
  );


  buf

  (
    g1284_n_spl_,
    g1284_n
  );


  buf

  (
    g1284_n_spl_0,
    g1284_n_spl_
  );


  buf

  (
    g1284_p_spl_,
    g1284_p
  );


  buf

  (
    g1284_p_spl_0,
    g1284_p_spl_
  );


  buf

  (
    g1285_n_spl_,
    g1285_n
  );


  buf

  (
    g1274_n_spl_,
    g1274_n
  );


  buf

  (
    g1285_p_spl_,
    g1285_p
  );


  buf

  (
    g1274_p_spl_,
    g1274_p
  );


  buf

  (
    g1286_n_spl_,
    g1286_n
  );


  buf

  (
    g1286_n_spl_0,
    g1286_n_spl_
  );


  buf

  (
    g1286_p_spl_,
    g1286_p
  );


  buf

  (
    g1286_p_spl_0,
    g1286_p_spl_
  );


  buf

  (
    g1290_n_spl_,
    g1290_n
  );


  buf

  (
    g1289_n_spl_,
    g1289_n
  );


  buf

  (
    g1290_p_spl_,
    g1290_p
  );


  buf

  (
    g1289_p_spl_,
    g1289_p
  );


  buf

  (
    g1291_n_spl_,
    g1291_n
  );


  buf

  (
    g1291_n_spl_0,
    g1291_n_spl_
  );


  buf

  (
    g1291_p_spl_,
    g1291_p
  );


  buf

  (
    g1291_p_spl_0,
    g1291_p_spl_
  );


  buf

  (
    g1292_n_spl_,
    g1292_n
  );


  buf

  (
    g1271_n_spl_,
    g1271_n
  );


  buf

  (
    g1292_p_spl_,
    g1292_p
  );


  buf

  (
    g1271_p_spl_,
    g1271_p
  );


  buf

  (
    g1297_n_spl_,
    g1297_n
  );


  buf

  (
    g1296_n_spl_,
    g1296_n
  );


  buf

  (
    g1297_p_spl_,
    g1297_p
  );


  buf

  (
    g1296_p_spl_,
    g1296_p
  );


  buf

  (
    g1298_n_spl_,
    g1298_n
  );


  buf

  (
    g1298_n_spl_0,
    g1298_n_spl_
  );


  buf

  (
    g1298_p_spl_,
    g1298_p
  );


  buf

  (
    g1298_p_spl_0,
    g1298_p_spl_
  );


  buf

  (
    n7323_o2_p_spl_,
    n7323_o2_p
  );


  buf

  (
    n7323_o2_p_spl_0,
    n7323_o2_p_spl_
  );


  buf

  (
    n7323_o2_p_spl_1,
    n7323_o2_p_spl_
  );


  buf

  (
    n7323_o2_n_spl_,
    n7323_o2_n
  );


  buf

  (
    n7323_o2_n_spl_0,
    n7323_o2_n_spl_
  );


  buf

  (
    g1302_n_spl_,
    g1302_n
  );


  buf

  (
    g1301_n_spl_,
    g1301_n
  );


  buf

  (
    g1302_p_spl_,
    g1302_p
  );


  buf

  (
    g1301_p_spl_,
    g1301_p
  );


  buf

  (
    g1303_n_spl_,
    g1303_n
  );


  buf

  (
    g1303_n_spl_0,
    g1303_n_spl_
  );


  buf

  (
    g1303_p_spl_,
    g1303_p
  );


  buf

  (
    g1303_p_spl_0,
    g1303_p_spl_
  );


  buf

  (
    G3394_o2_n_spl_,
    G3394_o2_n
  );


  buf

  (
    G3391_o2_n_spl_,
    G3391_o2_n
  );


  buf

  (
    G3394_o2_p_spl_,
    G3394_o2_p
  );


  buf

  (
    G3391_o2_p_spl_,
    G3391_o2_p
  );


  buf

  (
    g1307_n_spl_,
    g1307_n
  );


  buf

  (
    g1307_n_spl_0,
    g1307_n_spl_
  );


  buf

  (
    g1307_p_spl_,
    g1307_p
  );


  buf

  (
    g1307_p_spl_0,
    g1307_p_spl_
  );


  buf

  (
    n7398_o2_p_spl_,
    n7398_o2_p
  );


  buf

  (
    n7398_o2_p_spl_0,
    n7398_o2_p_spl_
  );


  buf

  (
    n7398_o2_p_spl_1,
    n7398_o2_p_spl_
  );


  buf

  (
    n7398_o2_n_spl_,
    n7398_o2_n
  );


  buf

  (
    n7398_o2_n_spl_0,
    n7398_o2_n_spl_
  );


  buf

  (
    g1311_n_spl_,
    g1311_n
  );


  buf

  (
    g1310_n_spl_,
    g1310_n
  );


  buf

  (
    g1311_p_spl_,
    g1311_p
  );


  buf

  (
    g1310_p_spl_,
    g1310_p
  );


  buf

  (
    g1312_n_spl_,
    g1312_n
  );


  buf

  (
    g1312_n_spl_0,
    g1312_n_spl_
  );


  buf

  (
    g1312_p_spl_,
    g1312_p
  );


  buf

  (
    g1312_p_spl_0,
    g1312_p_spl_
  );


  buf

  (
    g1313_n_spl_,
    g1313_n
  );


  buf

  (
    g1306_n_spl_,
    g1306_n
  );


  buf

  (
    g1313_p_spl_,
    g1313_p
  );


  buf

  (
    g1306_p_spl_,
    g1306_p
  );


  buf

  (
    g1314_n_spl_,
    g1314_n
  );


  buf

  (
    g1314_n_spl_0,
    g1314_n_spl_
  );


  buf

  (
    g1314_p_spl_,
    g1314_p
  );


  buf

  (
    g1314_p_spl_0,
    g1314_p_spl_
  );


  buf

  (
    g1318_n_spl_,
    g1318_n
  );


  buf

  (
    g1317_n_spl_,
    g1317_n
  );


  buf

  (
    g1318_p_spl_,
    g1318_p
  );


  buf

  (
    g1317_p_spl_,
    g1317_p
  );


  buf

  (
    g1319_n_spl_,
    g1319_n
  );


  buf

  (
    g1319_n_spl_0,
    g1319_n_spl_
  );


  buf

  (
    g1319_p_spl_,
    g1319_p
  );


  buf

  (
    g1319_p_spl_0,
    g1319_p_spl_
  );


  buf

  (
    n7459_o2_p_spl_,
    n7459_o2_p
  );


  buf

  (
    n7459_o2_p_spl_0,
    n7459_o2_p_spl_
  );


  buf

  (
    n7459_o2_p_spl_1,
    n7459_o2_p_spl_
  );


  buf

  (
    n7459_o2_n_spl_,
    n7459_o2_n
  );


  buf

  (
    n7459_o2_n_spl_0,
    n7459_o2_n_spl_
  );


  buf

  (
    n7459_o2_n_spl_1,
    n7459_o2_n_spl_
  );


  buf

  (
    g1327_n_spl_,
    g1327_n
  );


  buf

  (
    g1326_n_spl_,
    g1326_n
  );


  buf

  (
    g1327_p_spl_,
    g1327_p
  );


  buf

  (
    g1326_p_spl_,
    g1326_p
  );


  buf

  (
    g1328_n_spl_,
    g1328_n
  );


  buf

  (
    g1328_n_spl_0,
    g1328_n_spl_
  );


  buf

  (
    g1328_p_spl_,
    g1328_p
  );


  buf

  (
    g1328_p_spl_0,
    g1328_p_spl_
  );


  buf

  (
    g1329_n_spl_,
    g1329_n
  );


  buf

  (
    g1325_n_spl_,
    g1325_n
  );


  buf

  (
    g1329_p_spl_,
    g1329_p
  );


  buf

  (
    g1325_p_spl_,
    g1325_p
  );


  buf

  (
    g1330_n_spl_,
    g1330_n
  );


  buf

  (
    g1330_n_spl_0,
    g1330_n_spl_
  );


  buf

  (
    g1330_p_spl_,
    g1330_p
  );


  buf

  (
    g1330_p_spl_0,
    g1330_p_spl_
  );


  buf

  (
    g1334_n_spl_,
    g1334_n
  );


  buf

  (
    g1333_n_spl_,
    g1333_n
  );


  buf

  (
    g1334_p_spl_,
    g1334_p
  );


  buf

  (
    g1333_p_spl_,
    g1333_p
  );


  buf

  (
    g1335_n_spl_,
    g1335_n
  );


  buf

  (
    g1335_n_spl_0,
    g1335_n_spl_
  );


  buf

  (
    g1335_p_spl_,
    g1335_p
  );


  buf

  (
    g1335_p_spl_0,
    g1335_p_spl_
  );


  buf

  (
    g1336_n_spl_,
    g1336_n
  );


  buf

  (
    g1322_n_spl_,
    g1322_n
  );


  buf

  (
    g1336_p_spl_,
    g1336_p
  );


  buf

  (
    g1322_p_spl_,
    g1322_p
  );


  buf

  (
    g1337_n_spl_,
    g1337_n
  );


  buf

  (
    g1337_n_spl_0,
    g1337_n_spl_
  );


  buf

  (
    g1337_p_spl_,
    g1337_p
  );


  buf

  (
    g1337_p_spl_0,
    g1337_p_spl_
  );


  buf

  (
    g1341_n_spl_,
    g1341_n
  );


  buf

  (
    g1340_n_spl_,
    g1340_n
  );


  buf

  (
    g1341_p_spl_,
    g1341_p
  );


  buf

  (
    g1340_p_spl_,
    g1340_p
  );


  buf

  (
    g1342_n_spl_,
    g1342_n
  );


  buf

  (
    g1342_n_spl_0,
    g1342_n_spl_
  );


  buf

  (
    g1342_p_spl_,
    g1342_p
  );


  buf

  (
    g1342_p_spl_0,
    g1342_p_spl_
  );


  buf

  (
    G3722_o2_n_spl_,
    G3722_o2_n
  );


  buf

  (
    G3722_o2_n_spl_0,
    G3722_o2_n_spl_
  );


  buf

  (
    G3722_o2_p_spl_,
    G3722_o2_p
  );


  buf

  (
    G3722_o2_p_spl_0,
    G3722_o2_p_spl_
  );


  buf

  (
    g1352_n_spl_,
    g1352_n
  );


  buf

  (
    g1351_n_spl_,
    g1351_n
  );


  buf

  (
    g1352_p_spl_,
    g1352_p
  );


  buf

  (
    g1351_p_spl_,
    g1351_p
  );


  buf

  (
    g1353_n_spl_,
    g1353_n
  );


  buf

  (
    g1353_n_spl_0,
    g1353_n_spl_
  );


  buf

  (
    g1353_p_spl_,
    g1353_p
  );


  buf

  (
    g1353_p_spl_0,
    g1353_p_spl_
  );


  buf

  (
    n7501_o2_p_spl_,
    n7501_o2_p
  );


  buf

  (
    n7501_o2_p_spl_0,
    n7501_o2_p_spl_
  );


  buf

  (
    n7501_o2_p_spl_1,
    n7501_o2_p_spl_
  );


  buf

  (
    n7501_o2_n_spl_,
    n7501_o2_n
  );


  buf

  (
    n7501_o2_n_spl_0,
    n7501_o2_n_spl_
  );


  buf

  (
    g1357_n_spl_,
    g1357_n
  );


  buf

  (
    g1356_n_spl_,
    g1356_n
  );


  buf

  (
    g1357_p_spl_,
    g1357_p
  );


  buf

  (
    g1356_p_spl_,
    g1356_p
  );


  buf

  (
    g1358_n_spl_,
    g1358_n
  );


  buf

  (
    g1358_n_spl_0,
    g1358_n_spl_
  );


  buf

  (
    g1358_p_spl_,
    g1358_p
  );


  buf

  (
    g1358_p_spl_0,
    g1358_p_spl_
  );


  buf

  (
    g1359_n_spl_,
    g1359_n
  );


  buf

  (
    g1348_n_spl_,
    g1348_n
  );


  buf

  (
    g1359_p_spl_,
    g1359_p
  );


  buf

  (
    g1348_p_spl_,
    g1348_p
  );


  buf

  (
    g1360_n_spl_,
    g1360_n
  );


  buf

  (
    g1360_n_spl_0,
    g1360_n_spl_
  );


  buf

  (
    g1360_p_spl_,
    g1360_p
  );


  buf

  (
    g1360_p_spl_0,
    g1360_p_spl_
  );


  buf

  (
    g1364_n_spl_,
    g1364_n
  );


  buf

  (
    g1363_n_spl_,
    g1363_n
  );


  buf

  (
    g1364_p_spl_,
    g1364_p
  );


  buf

  (
    g1363_p_spl_,
    g1363_p
  );


  buf

  (
    g1365_n_spl_,
    g1365_n
  );


  buf

  (
    g1365_n_spl_0,
    g1365_n_spl_
  );


  buf

  (
    g1365_p_spl_,
    g1365_p
  );


  buf

  (
    g1365_p_spl_0,
    g1365_p_spl_
  );


  buf

  (
    g1366_n_spl_,
    g1366_n
  );


  buf

  (
    g1345_n_spl_,
    g1345_n
  );


  buf

  (
    g1366_p_spl_,
    g1366_p
  );


  buf

  (
    g1345_p_spl_,
    g1345_p
  );


  buf

  (
    G3719_o2_p_spl_,
    G3719_o2_p
  );


  buf

  (
    G902_o2_n_spl_,
    G902_o2_n
  );


  buf

  (
    G3719_o2_n_spl_,
    G3719_o2_n
  );


  buf

  (
    G902_o2_p_spl_,
    G902_o2_p
  );


  buf

  (
    g1371_n_spl_,
    g1371_n
  );


  buf

  (
    g1371_n_spl_0,
    g1371_n_spl_
  );


  buf

  (
    g1371_p_spl_,
    g1371_p
  );


  buf

  (
    g1371_p_spl_0,
    g1371_p_spl_
  );


  buf

  (
    g1372_n_spl_,
    g1372_n
  );


  buf

  (
    g1370_n_spl_,
    g1370_n
  );


  buf

  (
    g1372_p_spl_,
    g1372_p
  );


  buf

  (
    g1370_p_spl_,
    g1370_p
  );


  buf

  (
    g1373_n_spl_,
    g1373_n
  );


  buf

  (
    g1373_n_spl_0,
    g1373_n_spl_
  );


  buf

  (
    g1373_p_spl_,
    g1373_p
  );


  buf

  (
    g1373_p_spl_0,
    g1373_p_spl_
  );


  buf

  (
    n7518_o2_p_spl_,
    n7518_o2_p
  );


  buf

  (
    n7518_o2_p_spl_0,
    n7518_o2_p_spl_
  );


  buf

  (
    n7518_o2_p_spl_1,
    n7518_o2_p_spl_
  );


  buf

  (
    n7518_o2_n_spl_,
    n7518_o2_n
  );


  buf

  (
    n7518_o2_n_spl_0,
    n7518_o2_n_spl_
  );


  buf

  (
    g1377_n_spl_,
    g1377_n
  );


  buf

  (
    g1376_n_spl_,
    g1376_n
  );


  buf

  (
    g1377_p_spl_,
    g1377_p
  );


  buf

  (
    g1376_p_spl_,
    g1376_p
  );


  buf

  (
    g1378_n_spl_,
    g1378_n
  );


  buf

  (
    g1378_n_spl_0,
    g1378_n_spl_
  );


  buf

  (
    g1378_p_spl_,
    g1378_p
  );


  buf

  (
    g1378_p_spl_0,
    g1378_p_spl_
  );


  buf

  (
    n7606_o2_p_spl_,
    n7606_o2_p
  );


  buf

  (
    n7606_o2_p_spl_0,
    n7606_o2_p_spl_
  );


  buf

  (
    n7606_o2_p_spl_00,
    n7606_o2_p_spl_0
  );


  buf

  (
    n7606_o2_p_spl_1,
    n7606_o2_p_spl_
  );


  buf

  (
    n7606_o2_n_spl_,
    n7606_o2_n
  );


  buf

  (
    n7606_o2_n_spl_0,
    n7606_o2_n_spl_
  );


  buf

  (
    n7606_o2_n_spl_1,
    n7606_o2_n_spl_
  );


  buf

  (
    g1386_n_spl_,
    g1386_n
  );


  buf

  (
    g1385_n_spl_,
    g1385_n
  );


  buf

  (
    g1386_p_spl_,
    g1386_p
  );


  buf

  (
    g1385_p_spl_,
    g1385_p
  );


  buf

  (
    g1387_n_spl_,
    g1387_n
  );


  buf

  (
    g1387_n_spl_0,
    g1387_n_spl_
  );


  buf

  (
    g1387_p_spl_,
    g1387_p
  );


  buf

  (
    g1387_p_spl_0,
    g1387_p_spl_
  );


  buf

  (
    g1388_n_spl_,
    g1388_n
  );


  buf

  (
    g1384_n_spl_,
    g1384_n
  );


  buf

  (
    g1388_p_spl_,
    g1388_p
  );


  buf

  (
    g1384_p_spl_,
    g1384_p
  );


  buf

  (
    g1389_n_spl_,
    g1389_n
  );


  buf

  (
    g1389_n_spl_0,
    g1389_n_spl_
  );


  buf

  (
    g1389_p_spl_,
    g1389_p
  );


  buf

  (
    g1389_p_spl_0,
    g1389_p_spl_
  );


  buf

  (
    g1393_n_spl_,
    g1393_n
  );


  buf

  (
    g1392_n_spl_,
    g1392_n
  );


  buf

  (
    g1393_p_spl_,
    g1393_p
  );


  buf

  (
    g1392_p_spl_,
    g1392_p
  );


  buf

  (
    g1394_n_spl_,
    g1394_n
  );


  buf

  (
    g1394_n_spl_0,
    g1394_n_spl_
  );


  buf

  (
    g1394_p_spl_,
    g1394_p
  );


  buf

  (
    g1394_p_spl_0,
    g1394_p_spl_
  );


  buf

  (
    g1395_n_spl_,
    g1395_n
  );


  buf

  (
    g1381_n_spl_,
    g1381_n
  );


  buf

  (
    g1395_p_spl_,
    g1395_p
  );


  buf

  (
    g1381_p_spl_,
    g1381_p
  );


  buf

  (
    g1396_n_spl_,
    g1396_n
  );


  buf

  (
    g1396_n_spl_0,
    g1396_n_spl_
  );


  buf

  (
    g1396_p_spl_,
    g1396_p
  );


  buf

  (
    g1396_p_spl_0,
    g1396_p_spl_
  );


  buf

  (
    g1400_n_spl_,
    g1400_n
  );


  buf

  (
    g1399_n_spl_,
    g1399_n
  );


  buf

  (
    g1400_p_spl_,
    g1400_p
  );


  buf

  (
    g1399_p_spl_,
    g1399_p
  );


  buf

  (
    g1401_n_spl_,
    g1401_n
  );


  buf

  (
    g1401_n_spl_0,
    g1401_n_spl_
  );


  buf

  (
    g1401_p_spl_,
    g1401_p
  );


  buf

  (
    g1401_p_spl_0,
    g1401_p_spl_
  );


  buf

  (
    G3616_o2_p_spl_,
    G3616_o2_p
  );


  buf

  (
    G3616_o2_p_spl_0,
    G3616_o2_p_spl_
  );


  buf

  (
    G3616_o2_n_spl_,
    G3616_o2_n
  );


  buf

  (
    G3616_o2_n_spl_0,
    G3616_o2_n_spl_
  );


  buf

  (
    n7675_o2_p_spl_,
    n7675_o2_p
  );


  buf

  (
    n7675_o2_p_spl_0,
    n7675_o2_p_spl_
  );


  buf

  (
    n7675_o2_p_spl_00,
    n7675_o2_p_spl_0
  );


  buf

  (
    n7675_o2_p_spl_1,
    n7675_o2_p_spl_
  );


  buf

  (
    n7675_o2_n_spl_,
    n7675_o2_n
  );


  buf

  (
    n7675_o2_n_spl_0,
    n7675_o2_n_spl_
  );


  buf

  (
    n7675_o2_n_spl_00,
    n7675_o2_n_spl_0
  );


  buf

  (
    n7675_o2_n_spl_1,
    n7675_o2_n_spl_
  );


  buf

  (
    g1414_n_spl_,
    g1414_n
  );


  buf

  (
    g1413_n_spl_,
    g1413_n
  );


  buf

  (
    g1414_p_spl_,
    g1414_p
  );


  buf

  (
    g1413_p_spl_,
    g1413_p
  );


  buf

  (
    g1415_n_spl_,
    g1415_n
  );


  buf

  (
    g1415_n_spl_0,
    g1415_n_spl_
  );


  buf

  (
    g1415_p_spl_,
    g1415_p
  );


  buf

  (
    g1415_p_spl_0,
    g1415_p_spl_
  );


  buf

  (
    g1416_n_spl_,
    g1416_n
  );


  buf

  (
    g1410_n_spl_,
    g1410_n
  );


  buf

  (
    g1416_p_spl_,
    g1416_p
  );


  buf

  (
    g1410_p_spl_,
    g1410_p
  );


  buf

  (
    g1417_n_spl_,
    g1417_n
  );


  buf

  (
    g1417_n_spl_0,
    g1417_n_spl_
  );


  buf

  (
    g1417_p_spl_,
    g1417_p
  );


  buf

  (
    g1417_p_spl_0,
    g1417_p_spl_
  );


  buf

  (
    g1421_n_spl_,
    g1421_n
  );


  buf

  (
    g1420_n_spl_,
    g1420_n
  );


  buf

  (
    g1421_p_spl_,
    g1421_p
  );


  buf

  (
    g1420_p_spl_,
    g1420_p
  );


  buf

  (
    g1422_n_spl_,
    g1422_n
  );


  buf

  (
    g1422_n_spl_0,
    g1422_n_spl_
  );


  buf

  (
    g1422_p_spl_,
    g1422_p
  );


  buf

  (
    g1422_p_spl_0,
    g1422_p_spl_
  );


  buf

  (
    g1423_n_spl_,
    g1423_n
  );


  buf

  (
    g1407_n_spl_,
    g1407_n
  );


  buf

  (
    g1423_p_spl_,
    g1423_p
  );


  buf

  (
    g1407_p_spl_,
    g1407_p
  );


  buf

  (
    g1424_n_spl_,
    g1424_n
  );


  buf

  (
    g1424_n_spl_0,
    g1424_n_spl_
  );


  buf

  (
    g1424_p_spl_,
    g1424_p
  );


  buf

  (
    g1424_p_spl_0,
    g1424_p_spl_
  );


  buf

  (
    g1428_n_spl_,
    g1428_n
  );


  buf

  (
    g1427_n_spl_,
    g1427_n
  );


  buf

  (
    g1428_p_spl_,
    g1428_p
  );


  buf

  (
    g1427_p_spl_,
    g1427_p
  );


  buf

  (
    g1429_n_spl_,
    g1429_n
  );


  buf

  (
    g1429_n_spl_0,
    g1429_n_spl_
  );


  buf

  (
    g1429_p_spl_,
    g1429_p
  );


  buf

  (
    g1429_p_spl_0,
    g1429_p_spl_
  );


  buf

  (
    g1430_n_spl_,
    g1430_n
  );


  buf

  (
    g1404_n_spl_,
    g1404_n
  );


  buf

  (
    g1430_p_spl_,
    g1430_p
  );


  buf

  (
    g1404_p_spl_,
    g1404_p
  );


  buf

  (
    g1431_n_spl_,
    g1431_n
  );


  buf

  (
    g1431_n_spl_0,
    g1431_n_spl_
  );


  buf

  (
    g1431_p_spl_,
    g1431_p
  );


  buf

  (
    g1431_p_spl_0,
    g1431_p_spl_
  );


  buf

  (
    n2809_lo_p_spl_,
    n2809_lo_p
  );


  buf

  (
    n2809_lo_p_spl_0,
    n2809_lo_p_spl_
  );


  buf

  (
    n2809_lo_p_spl_00,
    n2809_lo_p_spl_0
  );


  buf

  (
    n2809_lo_p_spl_000,
    n2809_lo_p_spl_00
  );


  buf

  (
    n2809_lo_p_spl_001,
    n2809_lo_p_spl_00
  );


  buf

  (
    n2809_lo_p_spl_01,
    n2809_lo_p_spl_0
  );


  buf

  (
    n2809_lo_p_spl_1,
    n2809_lo_p_spl_
  );


  buf

  (
    n2809_lo_p_spl_10,
    n2809_lo_p_spl_1
  );


  buf

  (
    n2809_lo_p_spl_11,
    n2809_lo_p_spl_1
  );


  buf

  (
    n2809_lo_n_spl_,
    n2809_lo_n
  );


  buf

  (
    n2809_lo_n_spl_0,
    n2809_lo_n_spl_
  );


  buf

  (
    n2809_lo_n_spl_00,
    n2809_lo_n_spl_0
  );


  buf

  (
    n2809_lo_n_spl_000,
    n2809_lo_n_spl_00
  );


  buf

  (
    n2809_lo_n_spl_001,
    n2809_lo_n_spl_00
  );


  buf

  (
    n2809_lo_n_spl_01,
    n2809_lo_n_spl_0
  );


  buf

  (
    n2809_lo_n_spl_1,
    n2809_lo_n_spl_
  );


  buf

  (
    n2809_lo_n_spl_10,
    n2809_lo_n_spl_1
  );


  buf

  (
    n2809_lo_n_spl_11,
    n2809_lo_n_spl_1
  );


  buf

  (
    g1435_n_spl_,
    g1435_n
  );


  buf

  (
    g1434_n_spl_,
    g1434_n
  );


  buf

  (
    g1435_p_spl_,
    g1435_p
  );


  buf

  (
    g1434_p_spl_,
    g1434_p
  );


  buf

  (
    g1436_n_spl_,
    g1436_n
  );


  buf

  (
    g1436_n_spl_0,
    g1436_n_spl_
  );


  buf

  (
    g1436_p_spl_,
    g1436_p
  );


  buf

  (
    g1436_p_spl_0,
    g1436_p_spl_
  );


  buf

  (
    G3557_o2_n_spl_,
    G3557_o2_n
  );


  buf

  (
    G3494_o2_n_spl_,
    G3494_o2_n
  );


  buf

  (
    G3557_o2_p_spl_,
    G3557_o2_p
  );


  buf

  (
    G3494_o2_p_spl_,
    G3494_o2_p
  );


  buf

  (
    g1449_n_spl_,
    g1449_n
  );


  buf

  (
    g1449_n_spl_0,
    g1449_n_spl_
  );


  buf

  (
    g1449_p_spl_,
    g1449_p
  );


  buf

  (
    g1449_p_spl_0,
    g1449_p_spl_
  );


  buf

  (
    n7722_o2_p_spl_,
    n7722_o2_p
  );


  buf

  (
    n7722_o2_p_spl_0,
    n7722_o2_p_spl_
  );


  buf

  (
    n7722_o2_p_spl_00,
    n7722_o2_p_spl_0
  );


  buf

  (
    n7722_o2_p_spl_01,
    n7722_o2_p_spl_0
  );


  buf

  (
    n7722_o2_p_spl_1,
    n7722_o2_p_spl_
  );


  buf

  (
    n7722_o2_n_spl_,
    n7722_o2_n
  );


  buf

  (
    n7722_o2_n_spl_0,
    n7722_o2_n_spl_
  );


  buf

  (
    n7722_o2_n_spl_00,
    n7722_o2_n_spl_0
  );


  buf

  (
    n7722_o2_n_spl_1,
    n7722_o2_n_spl_
  );


  buf

  (
    g1453_n_spl_,
    g1453_n
  );


  buf

  (
    g1452_n_spl_,
    g1452_n
  );


  buf

  (
    g1453_p_spl_,
    g1453_p
  );


  buf

  (
    g1452_p_spl_,
    g1452_p
  );


  buf

  (
    g1454_n_spl_,
    g1454_n
  );


  buf

  (
    g1454_n_spl_0,
    g1454_n_spl_
  );


  buf

  (
    g1454_p_spl_,
    g1454_p
  );


  buf

  (
    g1454_p_spl_0,
    g1454_p_spl_
  );


  buf

  (
    g1455_n_spl_,
    g1455_n
  );


  buf

  (
    g1448_n_spl_,
    g1448_n
  );


  buf

  (
    g1455_p_spl_,
    g1455_p
  );


  buf

  (
    g1448_p_spl_,
    g1448_p
  );


  buf

  (
    g1456_n_spl_,
    g1456_n
  );


  buf

  (
    g1456_n_spl_0,
    g1456_n_spl_
  );


  buf

  (
    g1456_p_spl_,
    g1456_p
  );


  buf

  (
    g1456_p_spl_0,
    g1456_p_spl_
  );


  buf

  (
    g1460_n_spl_,
    g1460_n
  );


  buf

  (
    g1459_n_spl_,
    g1459_n
  );


  buf

  (
    g1460_p_spl_,
    g1460_p
  );


  buf

  (
    g1459_p_spl_,
    g1459_p
  );


  buf

  (
    g1461_n_spl_,
    g1461_n
  );


  buf

  (
    g1461_n_spl_0,
    g1461_n_spl_
  );


  buf

  (
    g1461_p_spl_,
    g1461_p
  );


  buf

  (
    g1461_p_spl_0,
    g1461_p_spl_
  );


  buf

  (
    g1462_n_spl_,
    g1462_n
  );


  buf

  (
    g1445_n_spl_,
    g1445_n
  );


  buf

  (
    g1462_p_spl_,
    g1462_p
  );


  buf

  (
    g1445_p_spl_,
    g1445_p
  );


  buf

  (
    g1463_n_spl_,
    g1463_n
  );


  buf

  (
    g1463_n_spl_0,
    g1463_n_spl_
  );


  buf

  (
    g1463_p_spl_,
    g1463_p
  );


  buf

  (
    g1463_p_spl_0,
    g1463_p_spl_
  );


  buf

  (
    g1467_n_spl_,
    g1467_n
  );


  buf

  (
    g1466_n_spl_,
    g1466_n
  );


  buf

  (
    g1467_p_spl_,
    g1467_p
  );


  buf

  (
    g1466_p_spl_,
    g1466_p
  );


  buf

  (
    g1468_n_spl_,
    g1468_n
  );


  buf

  (
    g1468_n_spl_0,
    g1468_n_spl_
  );


  buf

  (
    g1468_p_spl_,
    g1468_p
  );


  buf

  (
    g1468_p_spl_0,
    g1468_p_spl_
  );


  buf

  (
    g1469_n_spl_,
    g1469_n
  );


  buf

  (
    g1442_n_spl_,
    g1442_n
  );


  buf

  (
    g1469_p_spl_,
    g1469_p
  );


  buf

  (
    g1442_p_spl_,
    g1442_p
  );


  buf

  (
    g1470_n_spl_,
    g1470_n
  );


  buf

  (
    g1470_n_spl_0,
    g1470_n_spl_
  );


  buf

  (
    g1470_p_spl_,
    g1470_p
  );


  buf

  (
    g1470_p_spl_0,
    g1470_p_spl_
  );


  buf

  (
    g1474_n_spl_,
    g1474_n
  );


  buf

  (
    g1473_n_spl_,
    g1473_n
  );


  buf

  (
    g1474_p_spl_,
    g1474_p
  );


  buf

  (
    g1473_p_spl_,
    g1473_p
  );


  buf

  (
    g1475_n_spl_,
    g1475_n
  );


  buf

  (
    g1475_n_spl_0,
    g1475_n_spl_
  );


  buf

  (
    g1475_p_spl_,
    g1475_p
  );


  buf

  (
    g1475_p_spl_0,
    g1475_p_spl_
  );


  buf

  (
    g1476_n_spl_,
    g1476_n
  );


  buf

  (
    g1439_n_spl_,
    g1439_n
  );


  buf

  (
    g1476_p_spl_,
    g1476_p
  );


  buf

  (
    g1439_p_spl_,
    g1439_p
  );


  buf

  (
    G1724_o2_p_spl_,
    G1724_o2_p
  );


  buf

  (
    G692_o2_n_spl_,
    G692_o2_n
  );


  buf

  (
    G1724_o2_n_spl_,
    G1724_o2_n
  );


  buf

  (
    G692_o2_p_spl_,
    G692_o2_p
  );


  buf

  (
    g1478_n_spl_,
    g1478_n
  );


  buf

  (
    g1478_n_spl_0,
    g1478_n_spl_
  );


  buf

  (
    g1478_p_spl_,
    g1478_p
  );


  buf

  (
    g1478_p_spl_0,
    g1478_p_spl_
  );


  buf

  (
    g1482_n_spl_,
    g1482_n
  );


  buf

  (
    g1481_n_spl_,
    g1481_n
  );


  buf

  (
    g1482_p_spl_,
    g1482_p
  );


  buf

  (
    g1481_p_spl_,
    g1481_p
  );


  buf

  (
    g1483_n_spl_,
    g1483_n
  );


  buf

  (
    g1483_n_spl_0,
    g1483_n_spl_
  );


  buf

  (
    g1483_p_spl_,
    g1483_p
  );


  buf

  (
    g1483_p_spl_0,
    g1483_p_spl_
  );


  buf

  (
    g1487_n_spl_,
    g1487_n
  );


  buf

  (
    g1486_n_spl_,
    g1486_n
  );


  buf

  (
    g1487_p_spl_,
    g1487_p
  );


  buf

  (
    g1486_p_spl_,
    g1486_p
  );


  buf

  (
    g1488_n_spl_,
    g1488_n
  );


  buf

  (
    g1488_n_spl_0,
    g1488_n_spl_
  );


  buf

  (
    g1488_p_spl_,
    g1488_p
  );


  buf

  (
    g1488_p_spl_0,
    g1488_p_spl_
  );


  buf

  (
    g1492_n_spl_,
    g1492_n
  );


  buf

  (
    g1491_n_spl_,
    g1491_n
  );


  buf

  (
    g1492_p_spl_,
    g1492_p
  );


  buf

  (
    g1491_p_spl_,
    g1491_p
  );


  buf

  (
    g1493_n_spl_,
    g1493_n
  );


  buf

  (
    g1493_n_spl_0,
    g1493_n_spl_
  );


  buf

  (
    g1493_p_spl_,
    g1493_p
  );


  buf

  (
    g1493_p_spl_0,
    g1493_p_spl_
  );


  buf

  (
    g1497_n_spl_,
    g1497_n
  );


  buf

  (
    g1496_n_spl_,
    g1496_n
  );


  buf

  (
    g1497_p_spl_,
    g1497_p
  );


  buf

  (
    g1496_p_spl_,
    g1496_p
  );


  buf

  (
    g1498_n_spl_,
    g1498_n
  );


  buf

  (
    g1498_n_spl_0,
    g1498_n_spl_
  );


  buf

  (
    g1498_p_spl_,
    g1498_p
  );


  buf

  (
    g1498_p_spl_0,
    g1498_p_spl_
  );


  buf

  (
    g1097_p_spl_,
    g1097_p
  );


  buf

  (
    g1502_n_spl_,
    g1502_n
  );


  buf

  (
    g1501_n_spl_,
    g1501_n
  );


  buf

  (
    g1502_p_spl_,
    g1502_p
  );


  buf

  (
    g1501_p_spl_,
    g1501_p
  );


  buf

  (
    g1503_n_spl_,
    g1503_n
  );


  buf

  (
    g1503_n_spl_0,
    g1503_n_spl_
  );


  buf

  (
    g1503_p_spl_,
    g1503_p
  );


  buf

  (
    g1503_p_spl_0,
    g1503_p_spl_
  );


  buf

  (
    g1506_n_spl_,
    g1506_n
  );


  buf

  (
    g1215_p_spl_,
    g1215_p
  );


  buf

  (
    g1510_n_spl_,
    g1510_n
  );


  buf

  (
    g1509_n_spl_,
    g1509_n
  );


  buf

  (
    g1510_p_spl_,
    g1510_p
  );


  buf

  (
    g1509_p_spl_,
    g1509_p
  );


  buf

  (
    g1511_n_spl_,
    g1511_n
  );


  buf

  (
    g1511_n_spl_0,
    g1511_n_spl_
  );


  buf

  (
    g1511_p_spl_,
    g1511_p
  );


  buf

  (
    g1511_p_spl_0,
    g1511_p_spl_
  );


  buf

  (
    n7747_o2_p_spl_,
    n7747_o2_p
  );


  buf

  (
    n7747_o2_p_spl_0,
    n7747_o2_p_spl_
  );


  buf

  (
    n7747_o2_p_spl_00,
    n7747_o2_p_spl_0
  );


  buf

  (
    n7747_o2_p_spl_01,
    n7747_o2_p_spl_0
  );


  buf

  (
    n7747_o2_p_spl_1,
    n7747_o2_p_spl_
  );


  buf

  (
    n7747_o2_n_spl_,
    n7747_o2_n
  );


  buf

  (
    n7747_o2_n_spl_0,
    n7747_o2_n_spl_
  );


  buf

  (
    n7747_o2_n_spl_00,
    n7747_o2_n_spl_0
  );


  buf

  (
    n7747_o2_n_spl_1,
    n7747_o2_n_spl_
  );


  buf

  (
    g1515_n_spl_,
    g1515_n
  );


  buf

  (
    g1514_n_spl_,
    g1514_n
  );


  buf

  (
    g1515_p_spl_,
    g1515_p
  );


  buf

  (
    g1514_p_spl_,
    g1514_p
  );


  buf

  (
    g1516_n_spl_,
    g1516_n
  );


  buf

  (
    g1516_n_spl_0,
    g1516_n_spl_
  );


  buf

  (
    g1516_p_spl_,
    g1516_p
  );


  buf

  (
    g1516_p_spl_0,
    g1516_p_spl_
  );


  buf

  (
    g1520_n_spl_,
    g1520_n
  );


  buf

  (
    g1519_n_spl_,
    g1519_n
  );


  buf

  (
    g1520_p_spl_,
    g1520_p
  );


  buf

  (
    g1519_p_spl_,
    g1519_p
  );


  buf

  (
    g1521_n_spl_,
    g1521_n
  );


  buf

  (
    g1521_n_spl_0,
    g1521_n_spl_
  );


  buf

  (
    g1521_p_spl_,
    g1521_p
  );


  buf

  (
    g1521_p_spl_0,
    g1521_p_spl_
  );


  buf

  (
    g1525_n_spl_,
    g1525_n
  );


  buf

  (
    g1524_n_spl_,
    g1524_n
  );


  buf

  (
    g1525_p_spl_,
    g1525_p
  );


  buf

  (
    g1524_p_spl_,
    g1524_p
  );


  buf

  (
    g1526_n_spl_,
    g1526_n
  );


  buf

  (
    g1526_n_spl_0,
    g1526_n_spl_
  );


  buf

  (
    g1526_p_spl_,
    g1526_p
  );


  buf

  (
    g1526_p_spl_0,
    g1526_p_spl_
  );


  buf

  (
    g1530_n_spl_,
    g1530_n
  );


  buf

  (
    g1529_n_spl_,
    g1529_n
  );


  buf

  (
    g1530_p_spl_,
    g1530_p
  );


  buf

  (
    g1529_p_spl_,
    g1529_p
  );


  buf

  (
    g1531_n_spl_,
    g1531_n
  );


  buf

  (
    g1531_n_spl_0,
    g1531_n_spl_
  );


  buf

  (
    g1531_p_spl_,
    g1531_p
  );


  buf

  (
    g1531_p_spl_0,
    g1531_p_spl_
  );


  buf

  (
    g1535_n_spl_,
    g1535_n
  );


  buf

  (
    g1534_n_spl_,
    g1534_n
  );


  buf

  (
    g1535_p_spl_,
    g1535_p
  );


  buf

  (
    g1534_p_spl_,
    g1534_p
  );


  buf

  (
    g1536_n_spl_,
    g1536_n
  );


  buf

  (
    g1536_n_spl_0,
    g1536_n_spl_
  );


  buf

  (
    g1536_p_spl_,
    g1536_p
  );


  buf

  (
    g1536_p_spl_0,
    g1536_p_spl_
  );


  buf

  (
    g1075_p_spl_,
    g1075_p
  );


  buf

  (
    g1540_n_spl_,
    g1540_n
  );


  buf

  (
    g1539_n_spl_,
    g1539_n
  );


  buf

  (
    g1540_p_spl_,
    g1540_p
  );


  buf

  (
    g1539_p_spl_,
    g1539_p
  );


  buf

  (
    g1541_n_spl_,
    g1541_n
  );


  buf

  (
    g1541_n_spl_0,
    g1541_n_spl_
  );


  buf

  (
    g1541_p_spl_,
    g1541_p
  );


  buf

  (
    g1541_p_spl_0,
    g1541_p_spl_
  );


  buf

  (
    g1231_p_spl_,
    g1231_p
  );


  buf

  (
    g1552_n_spl_,
    g1552_n
  );


  buf

  (
    g1551_n_spl_,
    g1551_n
  );


  buf

  (
    g1552_p_spl_,
    g1552_p
  );


  buf

  (
    g1551_p_spl_,
    g1551_p
  );


  buf

  (
    g1553_n_spl_,
    g1553_n
  );


  buf

  (
    g1553_n_spl_0,
    g1553_n_spl_
  );


  buf

  (
    g1553_p_spl_,
    g1553_p
  );


  buf

  (
    g1557_n_spl_,
    g1557_n
  );


  buf

  (
    g1556_n_spl_,
    g1556_n
  );


  buf

  (
    g1557_p_spl_,
    g1557_p
  );


  buf

  (
    g1556_p_spl_,
    g1556_p
  );


  buf

  (
    g1558_n_spl_,
    g1558_n
  );


  buf

  (
    g1558_n_spl_0,
    g1558_n_spl_
  );


  buf

  (
    g1558_p_spl_,
    g1558_p
  );


  buf

  (
    g1567_n_spl_,
    g1567_n
  );


  buf

  (
    g1566_n_spl_,
    g1566_n
  );


  buf

  (
    g1567_p_spl_,
    g1567_p
  );


  buf

  (
    g1566_p_spl_,
    g1566_p
  );


  buf

  (
    g1568_n_spl_,
    g1568_n
  );


  buf

  (
    g1568_n_spl_0,
    g1568_n_spl_
  );


  buf

  (
    g1568_p_spl_,
    g1568_p
  );


  buf

  (
    g1572_n_spl_,
    g1572_n
  );


  buf

  (
    g1571_n_spl_,
    g1571_n
  );


  buf

  (
    g1572_p_spl_,
    g1572_p
  );


  buf

  (
    g1571_p_spl_,
    g1571_p
  );


  buf

  (
    g1573_n_spl_,
    g1573_n
  );


  buf

  (
    g1573_n_spl_0,
    g1573_n_spl_
  );


  buf

  (
    g1573_p_spl_,
    g1573_p
  );


  buf

  (
    g1582_n_spl_,
    g1582_n
  );


  buf

  (
    g1581_n_spl_,
    g1581_n
  );


  buf

  (
    g1582_p_spl_,
    g1582_p
  );


  buf

  (
    g1581_p_spl_,
    g1581_p
  );


  buf

  (
    g1583_n_spl_,
    g1583_n
  );


  buf

  (
    g1583_n_spl_0,
    g1583_n_spl_
  );


  buf

  (
    g1583_p_spl_,
    g1583_p
  );


  buf

  (
    g1587_n_spl_,
    g1587_n
  );


  buf

  (
    g1586_n_spl_,
    g1586_n
  );


  buf

  (
    g1587_p_spl_,
    g1587_p
  );


  buf

  (
    g1586_p_spl_,
    g1586_p
  );


  buf

  (
    g1588_n_spl_,
    g1588_n
  );


  buf

  (
    g1588_n_spl_0,
    g1588_n_spl_
  );


  buf

  (
    g1588_p_spl_,
    g1588_p
  );


  buf

  (
    g1101_n_spl_,
    g1101_n
  );


  buf

  (
    g1101_n_spl_0,
    g1101_n_spl_
  );


  buf

  (
    g1126_n_spl_,
    g1126_n
  );


  buf

  (
    g1126_n_spl_0,
    g1126_n_spl_
  );


  buf

  (
    g1151_n_spl_,
    g1151_n
  );


  buf

  (
    g1151_n_spl_0,
    g1151_n_spl_
  );


  buf

  (
    g1206_n_spl_,
    g1206_n
  );


  buf

  (
    g1206_n_spl_0,
    g1206_n_spl_
  );


  buf

  (
    g1544_n_spl_,
    g1544_n
  );


  buf

  (
    g1507_p_spl_,
    g1507_p
  );


  buf

  (
    g1608_n_spl_,
    g1608_n
  );


  buf

  (
    g1607_n_spl_,
    g1607_n
  );


  buf

  (
    g1608_p_spl_,
    g1608_p
  );


  buf

  (
    g1607_p_spl_,
    g1607_p
  );


  buf

  (
    g1609_n_spl_,
    g1609_n
  );


  buf

  (
    g1609_n_spl_0,
    g1609_n_spl_
  );


  buf

  (
    g1609_p_spl_,
    g1609_p
  );


  buf

  (
    g1609_p_spl_0,
    g1609_p_spl_
  );


  buf

  (
    g1613_n_spl_,
    g1613_n
  );


  buf

  (
    g1612_n_spl_,
    g1612_n
  );


  buf

  (
    g1613_p_spl_,
    g1613_p
  );


  buf

  (
    g1612_p_spl_,
    g1612_p
  );


  buf

  (
    g1614_n_spl_,
    g1614_n
  );


  buf

  (
    g1614_n_spl_0,
    g1614_n_spl_
  );


  buf

  (
    g1614_p_spl_,
    g1614_p
  );


  buf

  (
    g1614_p_spl_0,
    g1614_p_spl_
  );


  buf

  (
    g1623_n_spl_,
    g1623_n
  );


  buf

  (
    g1622_n_spl_,
    g1622_n
  );


  buf

  (
    g1623_p_spl_,
    g1623_p
  );


  buf

  (
    g1622_p_spl_,
    g1622_p
  );


  buf

  (
    g1624_n_spl_,
    g1624_n
  );


  buf

  (
    g1624_n_spl_0,
    g1624_n_spl_
  );


  buf

  (
    g1624_p_spl_,
    g1624_p
  );


  buf

  (
    g1624_p_spl_0,
    g1624_p_spl_
  );


  buf

  (
    g1628_n_spl_,
    g1628_n
  );


  buf

  (
    g1627_n_spl_,
    g1627_n
  );


  buf

  (
    g1628_p_spl_,
    g1628_p
  );


  buf

  (
    g1627_p_spl_,
    g1627_p
  );


  buf

  (
    g1629_n_spl_,
    g1629_n
  );


  buf

  (
    g1629_n_spl_0,
    g1629_n_spl_
  );


  buf

  (
    g1629_p_spl_,
    g1629_p
  );


  buf

  (
    g1629_p_spl_0,
    g1629_p_spl_
  );


  buf

  (
    g1633_n_spl_,
    g1633_n
  );


  buf

  (
    g1632_n_spl_,
    g1632_n
  );


  buf

  (
    g1633_p_spl_,
    g1633_p
  );


  buf

  (
    g1632_p_spl_,
    g1632_p
  );


  buf

  (
    g1634_n_spl_,
    g1634_n
  );


  buf

  (
    g1634_n_spl_0,
    g1634_n_spl_
  );


  buf

  (
    g1634_p_spl_,
    g1634_p
  );


  buf

  (
    g1634_p_spl_0,
    g1634_p_spl_
  );


  buf

  (
    g1638_n_spl_,
    g1638_n
  );


  buf

  (
    g1637_n_spl_,
    g1637_n
  );


  buf

  (
    g1638_p_spl_,
    g1638_p
  );


  buf

  (
    g1637_p_spl_,
    g1637_p
  );


  buf

  (
    g1639_n_spl_,
    g1639_n
  );


  buf

  (
    g1639_n_spl_0,
    g1639_n_spl_
  );


  buf

  (
    g1639_p_spl_,
    g1639_p
  );


  buf

  (
    g1639_p_spl_0,
    g1639_p_spl_
  );


  buf

  (
    g1648_n_spl_,
    g1648_n
  );


  buf

  (
    g1647_n_spl_,
    g1647_n
  );


  buf

  (
    g1648_p_spl_,
    g1648_p
  );


  buf

  (
    g1647_p_spl_,
    g1647_p
  );


  buf

  (
    g1649_n_spl_,
    g1649_n
  );


  buf

  (
    g1649_n_spl_0,
    g1649_n_spl_
  );


  buf

  (
    g1649_p_spl_,
    g1649_p
  );


  buf

  (
    g1649_p_spl_0,
    g1649_p_spl_
  );


  buf

  (
    g1653_n_spl_,
    g1653_n
  );


  buf

  (
    g1652_n_spl_,
    g1652_n
  );


  buf

  (
    g1653_p_spl_,
    g1653_p
  );


  buf

  (
    g1652_p_spl_,
    g1652_p
  );


  buf

  (
    g1654_n_spl_,
    g1654_n
  );


  buf

  (
    g1654_n_spl_0,
    g1654_n_spl_
  );


  buf

  (
    g1654_p_spl_,
    g1654_p
  );


  buf

  (
    g1654_p_spl_0,
    g1654_p_spl_
  );


  buf

  (
    g1658_n_spl_,
    g1658_n
  );


  buf

  (
    g1657_n_spl_,
    g1657_n
  );


  buf

  (
    g1658_p_spl_,
    g1658_p
  );


  buf

  (
    g1657_p_spl_,
    g1657_p
  );


  buf

  (
    g1659_n_spl_,
    g1659_n
  );


  buf

  (
    g1659_n_spl_0,
    g1659_n_spl_
  );


  buf

  (
    g1659_p_spl_,
    g1659_p
  );


  buf

  (
    g1659_p_spl_0,
    g1659_p_spl_
  );


  buf

  (
    g1663_n_spl_,
    g1663_n
  );


  buf

  (
    g1662_n_spl_,
    g1662_n
  );


  buf

  (
    g1663_p_spl_,
    g1663_p
  );


  buf

  (
    g1662_p_spl_,
    g1662_p
  );


  buf

  (
    g1664_n_spl_,
    g1664_n
  );


  buf

  (
    g1664_n_spl_0,
    g1664_n_spl_
  );


  buf

  (
    g1664_p_spl_,
    g1664_p
  );


  buf

  (
    g1664_p_spl_0,
    g1664_p_spl_
  );


  buf

  (
    g1679_n_spl_,
    g1679_n
  );


  buf

  (
    g1678_n_spl_,
    g1678_n
  );


  buf

  (
    g1679_p_spl_,
    g1679_p
  );


  buf

  (
    g1678_p_spl_,
    g1678_p
  );


  buf

  (
    g1680_n_spl_,
    g1680_n
  );


  buf

  (
    g1680_n_spl_0,
    g1680_n_spl_
  );


  buf

  (
    g1680_p_spl_,
    g1680_p
  );


  buf

  (
    g1680_p_spl_0,
    g1680_p_spl_
  );


  buf

  (
    g1684_n_spl_,
    g1684_n
  );


  buf

  (
    g1683_n_spl_,
    g1683_n
  );


  buf

  (
    g1684_p_spl_,
    g1684_p
  );


  buf

  (
    g1683_p_spl_,
    g1683_p
  );


  buf

  (
    g1685_n_spl_,
    g1685_n
  );


  buf

  (
    g1685_n_spl_0,
    g1685_n_spl_
  );


  buf

  (
    g1685_p_spl_,
    g1685_p
  );


  buf

  (
    g1685_p_spl_0,
    g1685_p_spl_
  );


  buf

  (
    g1686_n_spl_,
    g1686_n
  );


  buf

  (
    g1675_n_spl_,
    g1675_n
  );


  buf

  (
    g1686_p_spl_,
    g1686_p
  );


  buf

  (
    g1675_p_spl_,
    g1675_p
  );


  buf

  (
    g1687_n_spl_,
    g1687_n
  );


  buf

  (
    g1687_n_spl_0,
    g1687_n_spl_
  );


  buf

  (
    g1687_p_spl_,
    g1687_p
  );


  buf

  (
    g1687_p_spl_0,
    g1687_p_spl_
  );


  buf

  (
    g1691_n_spl_,
    g1691_n
  );


  buf

  (
    g1690_n_spl_,
    g1690_n
  );


  buf

  (
    g1691_p_spl_,
    g1691_p
  );


  buf

  (
    g1690_p_spl_,
    g1690_p
  );


  buf

  (
    g1692_n_spl_,
    g1692_n
  );


  buf

  (
    g1692_n_spl_0,
    g1692_n_spl_
  );


  buf

  (
    g1692_p_spl_,
    g1692_p
  );


  buf

  (
    g1692_p_spl_0,
    g1692_p_spl_
  );


  buf

  (
    g1693_n_spl_,
    g1693_n
  );


  buf

  (
    g1672_n_spl_,
    g1672_n
  );


  buf

  (
    g1693_p_spl_,
    g1693_p
  );


  buf

  (
    g1672_p_spl_,
    g1672_p
  );


  buf

  (
    g1694_n_spl_,
    g1694_n
  );


  buf

  (
    g1694_n_spl_0,
    g1694_n_spl_
  );


  buf

  (
    g1694_p_spl_,
    g1694_p
  );


  buf

  (
    g1694_p_spl_0,
    g1694_p_spl_
  );


  buf

  (
    g1698_n_spl_,
    g1698_n
  );


  buf

  (
    g1697_n_spl_,
    g1697_n
  );


  buf

  (
    g1698_p_spl_,
    g1698_p
  );


  buf

  (
    g1697_p_spl_,
    g1697_p
  );


  buf

  (
    g1699_n_spl_,
    g1699_n
  );


  buf

  (
    g1699_n_spl_0,
    g1699_n_spl_
  );


  buf

  (
    g1699_p_spl_,
    g1699_p
  );


  buf

  (
    g1699_p_spl_0,
    g1699_p_spl_
  );


  buf

  (
    g1709_n_spl_,
    g1709_n
  );


  buf

  (
    g1708_n_spl_,
    g1708_n
  );


  buf

  (
    g1709_p_spl_,
    g1709_p
  );


  buf

  (
    g1708_p_spl_,
    g1708_p
  );


  buf

  (
    g1710_n_spl_,
    g1710_n
  );


  buf

  (
    g1710_n_spl_0,
    g1710_n_spl_
  );


  buf

  (
    g1710_p_spl_,
    g1710_p
  );


  buf

  (
    g1710_p_spl_0,
    g1710_p_spl_
  );


  buf

  (
    g1714_n_spl_,
    g1714_n
  );


  buf

  (
    g1713_n_spl_,
    g1713_n
  );


  buf

  (
    g1714_p_spl_,
    g1714_p
  );


  buf

  (
    g1713_p_spl_,
    g1713_p
  );


  buf

  (
    g1715_n_spl_,
    g1715_n
  );


  buf

  (
    g1715_n_spl_0,
    g1715_n_spl_
  );


  buf

  (
    g1715_p_spl_,
    g1715_p
  );


  buf

  (
    g1715_p_spl_0,
    g1715_p_spl_
  );


  buf

  (
    g1716_n_spl_,
    g1716_n
  );


  buf

  (
    g1705_n_spl_,
    g1705_n
  );


  buf

  (
    g1716_p_spl_,
    g1716_p
  );


  buf

  (
    g1705_p_spl_,
    g1705_p
  );


  buf

  (
    g1717_n_spl_,
    g1717_n
  );


  buf

  (
    g1717_n_spl_0,
    g1717_n_spl_
  );


  buf

  (
    g1717_p_spl_,
    g1717_p
  );


  buf

  (
    g1717_p_spl_0,
    g1717_p_spl_
  );


  buf

  (
    g1721_n_spl_,
    g1721_n
  );


  buf

  (
    g1720_n_spl_,
    g1720_n
  );


  buf

  (
    g1721_p_spl_,
    g1721_p
  );


  buf

  (
    g1720_p_spl_,
    g1720_p
  );


  buf

  (
    g1722_n_spl_,
    g1722_n
  );


  buf

  (
    g1722_n_spl_0,
    g1722_n_spl_
  );


  buf

  (
    g1722_p_spl_,
    g1722_p
  );


  buf

  (
    g1722_p_spl_0,
    g1722_p_spl_
  );


  buf

  (
    n2668_lo_buf_o2_p_spl_,
    n2668_lo_buf_o2_p
  );


  buf

  (
    n2668_lo_buf_o2_p_spl_0,
    n2668_lo_buf_o2_p_spl_
  );


  buf

  (
    n2668_lo_buf_o2_p_spl_00,
    n2668_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2668_lo_buf_o2_p_spl_1,
    n2668_lo_buf_o2_p_spl_
  );


  buf

  (
    n2668_lo_buf_o2_n_spl_,
    n2668_lo_buf_o2_n
  );


  buf

  (
    n2668_lo_buf_o2_n_spl_0,
    n2668_lo_buf_o2_n_spl_
  );


  buf

  (
    g1726_n_spl_,
    g1726_n
  );


  buf

  (
    g1725_n_spl_,
    g1725_n
  );


  buf

  (
    g1726_p_spl_,
    g1726_p
  );


  buf

  (
    g1725_p_spl_,
    g1725_p
  );


  buf

  (
    g1727_n_spl_,
    g1727_n
  );


  buf

  (
    g1727_n_spl_0,
    g1727_n_spl_
  );


  buf

  (
    g1727_p_spl_,
    g1727_p
  );


  buf

  (
    g1727_p_spl_0,
    g1727_p_spl_
  );


  buf

  (
    n2656_lo_buf_o2_p_spl_,
    n2656_lo_buf_o2_p
  );


  buf

  (
    n2656_lo_buf_o2_p_spl_0,
    n2656_lo_buf_o2_p_spl_
  );


  buf

  (
    n2656_lo_buf_o2_p_spl_1,
    n2656_lo_buf_o2_p_spl_
  );


  buf

  (
    n2656_lo_buf_o2_n_spl_,
    n2656_lo_buf_o2_n
  );


  buf

  (
    n2656_lo_buf_o2_n_spl_0,
    n2656_lo_buf_o2_n_spl_
  );


  buf

  (
    g1731_n_spl_,
    g1731_n
  );


  buf

  (
    g1730_n_spl_,
    g1730_n
  );


  buf

  (
    g1731_p_spl_,
    g1731_p
  );


  buf

  (
    g1730_p_spl_,
    g1730_p
  );


  buf

  (
    g1732_n_spl_,
    g1732_n
  );


  buf

  (
    g1732_n_spl_0,
    g1732_n_spl_
  );


  buf

  (
    g1732_p_spl_,
    g1732_p
  );


  buf

  (
    g1732_p_spl_0,
    g1732_p_spl_
  );


  buf

  (
    G2139_o2_n_spl_,
    G2139_o2_n
  );


  buf

  (
    G2136_o2_n_spl_,
    G2136_o2_n
  );


  buf

  (
    G2139_o2_p_spl_,
    G2139_o2_p
  );


  buf

  (
    G2136_o2_p_spl_,
    G2136_o2_p
  );


  buf

  (
    g1736_n_spl_,
    g1736_n
  );


  buf

  (
    g1736_n_spl_0,
    g1736_n_spl_
  );


  buf

  (
    g1736_p_spl_,
    g1736_p
  );


  buf

  (
    g1736_p_spl_0,
    g1736_p_spl_
  );


  buf

  (
    n2644_lo_buf_o2_p_spl_,
    n2644_lo_buf_o2_p
  );


  buf

  (
    n2644_lo_buf_o2_p_spl_0,
    n2644_lo_buf_o2_p_spl_
  );


  buf

  (
    n2644_lo_buf_o2_p_spl_1,
    n2644_lo_buf_o2_p_spl_
  );


  buf

  (
    n2644_lo_buf_o2_n_spl_,
    n2644_lo_buf_o2_n
  );


  buf

  (
    n2644_lo_buf_o2_n_spl_0,
    n2644_lo_buf_o2_n_spl_
  );


  buf

  (
    g1740_n_spl_,
    g1740_n
  );


  buf

  (
    g1739_n_spl_,
    g1739_n
  );


  buf

  (
    g1740_p_spl_,
    g1740_p
  );


  buf

  (
    g1739_p_spl_,
    g1739_p
  );


  buf

  (
    g1741_n_spl_,
    g1741_n
  );


  buf

  (
    g1741_n_spl_0,
    g1741_n_spl_
  );


  buf

  (
    g1741_p_spl_,
    g1741_p
  );


  buf

  (
    g1741_p_spl_0,
    g1741_p_spl_
  );


  buf

  (
    g1742_n_spl_,
    g1742_n
  );


  buf

  (
    g1735_n_spl_,
    g1735_n
  );


  buf

  (
    g1742_p_spl_,
    g1742_p
  );


  buf

  (
    g1735_p_spl_,
    g1735_p
  );


  buf

  (
    g1743_n_spl_,
    g1743_n
  );


  buf

  (
    g1743_n_spl_0,
    g1743_n_spl_
  );


  buf

  (
    g1743_p_spl_,
    g1743_p
  );


  buf

  (
    g1743_p_spl_0,
    g1743_p_spl_
  );


  buf

  (
    g1747_n_spl_,
    g1747_n
  );


  buf

  (
    g1746_n_spl_,
    g1746_n
  );


  buf

  (
    g1747_p_spl_,
    g1747_p
  );


  buf

  (
    g1746_p_spl_,
    g1746_p
  );


  buf

  (
    g1748_n_spl_,
    g1748_n
  );


  buf

  (
    g1748_n_spl_0,
    g1748_n_spl_
  );


  buf

  (
    g1748_p_spl_,
    g1748_p
  );


  buf

  (
    g1748_p_spl_0,
    g1748_p_spl_
  );


  buf

  (
    n2632_lo_buf_o2_p_spl_,
    n2632_lo_buf_o2_p
  );


  buf

  (
    n2632_lo_buf_o2_p_spl_0,
    n2632_lo_buf_o2_p_spl_
  );


  buf

  (
    n2632_lo_buf_o2_p_spl_1,
    n2632_lo_buf_o2_p_spl_
  );


  buf

  (
    n2632_lo_buf_o2_n_spl_,
    n2632_lo_buf_o2_n
  );


  buf

  (
    n2632_lo_buf_o2_n_spl_0,
    n2632_lo_buf_o2_n_spl_
  );


  buf

  (
    n2632_lo_buf_o2_n_spl_1,
    n2632_lo_buf_o2_n_spl_
  );


  buf

  (
    g1756_n_spl_,
    g1756_n
  );


  buf

  (
    g1755_n_spl_,
    g1755_n
  );


  buf

  (
    g1756_p_spl_,
    g1756_p
  );


  buf

  (
    g1755_p_spl_,
    g1755_p
  );


  buf

  (
    g1757_n_spl_,
    g1757_n
  );


  buf

  (
    g1757_n_spl_0,
    g1757_n_spl_
  );


  buf

  (
    g1757_p_spl_,
    g1757_p
  );


  buf

  (
    g1757_p_spl_0,
    g1757_p_spl_
  );


  buf

  (
    g1758_n_spl_,
    g1758_n
  );


  buf

  (
    g1754_n_spl_,
    g1754_n
  );


  buf

  (
    g1758_p_spl_,
    g1758_p
  );


  buf

  (
    g1754_p_spl_,
    g1754_p
  );


  buf

  (
    g1759_n_spl_,
    g1759_n
  );


  buf

  (
    g1759_n_spl_0,
    g1759_n_spl_
  );


  buf

  (
    g1759_p_spl_,
    g1759_p
  );


  buf

  (
    g1759_p_spl_0,
    g1759_p_spl_
  );


  buf

  (
    g1763_n_spl_,
    g1763_n
  );


  buf

  (
    g1762_n_spl_,
    g1762_n
  );


  buf

  (
    g1763_p_spl_,
    g1763_p
  );


  buf

  (
    g1762_p_spl_,
    g1762_p
  );


  buf

  (
    g1764_n_spl_,
    g1764_n
  );


  buf

  (
    g1764_n_spl_0,
    g1764_n_spl_
  );


  buf

  (
    g1764_p_spl_,
    g1764_p
  );


  buf

  (
    g1764_p_spl_0,
    g1764_p_spl_
  );


  buf

  (
    g1765_n_spl_,
    g1765_n
  );


  buf

  (
    g1751_n_spl_,
    g1751_n
  );


  buf

  (
    g1765_p_spl_,
    g1765_p
  );


  buf

  (
    g1751_p_spl_,
    g1751_p
  );


  buf

  (
    g1766_n_spl_,
    g1766_n
  );


  buf

  (
    g1766_n_spl_0,
    g1766_n_spl_
  );


  buf

  (
    g1766_p_spl_,
    g1766_p
  );


  buf

  (
    g1766_p_spl_0,
    g1766_p_spl_
  );


  buf

  (
    n2746_lo_p_spl_,
    n2746_lo_p
  );


  buf

  (
    n2746_lo_p_spl_0,
    n2746_lo_p_spl_
  );


  buf

  (
    n2746_lo_p_spl_00,
    n2746_lo_p_spl_0
  );


  buf

  (
    n2746_lo_p_spl_000,
    n2746_lo_p_spl_00
  );


  buf

  (
    n2746_lo_p_spl_001,
    n2746_lo_p_spl_00
  );


  buf

  (
    n2746_lo_p_spl_01,
    n2746_lo_p_spl_0
  );


  buf

  (
    n2746_lo_p_spl_010,
    n2746_lo_p_spl_01
  );


  buf

  (
    n2746_lo_p_spl_011,
    n2746_lo_p_spl_01
  );


  buf

  (
    n2746_lo_p_spl_1,
    n2746_lo_p_spl_
  );


  buf

  (
    n2746_lo_p_spl_10,
    n2746_lo_p_spl_1
  );


  buf

  (
    n2746_lo_p_spl_100,
    n2746_lo_p_spl_10
  );


  buf

  (
    n2746_lo_p_spl_101,
    n2746_lo_p_spl_10
  );


  buf

  (
    n2746_lo_p_spl_11,
    n2746_lo_p_spl_1
  );


  buf

  (
    n2746_lo_p_spl_110,
    n2746_lo_p_spl_11
  );


  buf

  (
    n2746_lo_n_spl_,
    n2746_lo_n
  );


  buf

  (
    n2746_lo_n_spl_0,
    n2746_lo_n_spl_
  );


  buf

  (
    n2746_lo_n_spl_00,
    n2746_lo_n_spl_0
  );


  buf

  (
    n2746_lo_n_spl_000,
    n2746_lo_n_spl_00
  );


  buf

  (
    n2746_lo_n_spl_001,
    n2746_lo_n_spl_00
  );


  buf

  (
    n2746_lo_n_spl_01,
    n2746_lo_n_spl_0
  );


  buf

  (
    n2746_lo_n_spl_010,
    n2746_lo_n_spl_01
  );


  buf

  (
    n2746_lo_n_spl_011,
    n2746_lo_n_spl_01
  );


  buf

  (
    n2746_lo_n_spl_1,
    n2746_lo_n_spl_
  );


  buf

  (
    n2746_lo_n_spl_10,
    n2746_lo_n_spl_1
  );


  buf

  (
    n2746_lo_n_spl_100,
    n2746_lo_n_spl_10
  );


  buf

  (
    n2746_lo_n_spl_101,
    n2746_lo_n_spl_10
  );


  buf

  (
    n2746_lo_n_spl_11,
    n2746_lo_n_spl_1
  );


  buf

  (
    n2746_lo_n_spl_110,
    n2746_lo_n_spl_11
  );


  buf

  (
    g1770_n_spl_,
    g1770_n
  );


  buf

  (
    g1769_n_spl_,
    g1769_n
  );


  buf

  (
    g1770_p_spl_,
    g1770_p
  );


  buf

  (
    g1769_p_spl_,
    g1769_p
  );


  buf

  (
    g1771_n_spl_,
    g1771_n
  );


  buf

  (
    g1771_n_spl_0,
    g1771_n_spl_
  );


  buf

  (
    g1771_p_spl_,
    g1771_p
  );


  buf

  (
    g1771_p_spl_0,
    g1771_p_spl_
  );


  buf

  (
    G2309_o2_p_spl_,
    G2309_o2_p
  );


  buf

  (
    G2309_o2_p_spl_0,
    G2309_o2_p_spl_
  );


  buf

  (
    G2309_o2_n_spl_,
    G2309_o2_n
  );


  buf

  (
    G2309_o2_n_spl_0,
    G2309_o2_n_spl_
  );


  buf

  (
    n2620_lo_buf_o2_p_spl_,
    n2620_lo_buf_o2_p
  );


  buf

  (
    n2620_lo_buf_o2_p_spl_0,
    n2620_lo_buf_o2_p_spl_
  );


  buf

  (
    n2620_lo_buf_o2_p_spl_00,
    n2620_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2620_lo_buf_o2_p_spl_1,
    n2620_lo_buf_o2_p_spl_
  );


  buf

  (
    n2620_lo_buf_o2_n_spl_,
    n2620_lo_buf_o2_n
  );


  buf

  (
    n2620_lo_buf_o2_n_spl_0,
    n2620_lo_buf_o2_n_spl_
  );


  buf

  (
    n2620_lo_buf_o2_n_spl_1,
    n2620_lo_buf_o2_n_spl_
  );


  buf

  (
    g1784_n_spl_,
    g1784_n
  );


  buf

  (
    g1783_n_spl_,
    g1783_n
  );


  buf

  (
    g1784_p_spl_,
    g1784_p
  );


  buf

  (
    g1783_p_spl_,
    g1783_p
  );


  buf

  (
    g1785_n_spl_,
    g1785_n
  );


  buf

  (
    g1785_n_spl_0,
    g1785_n_spl_
  );


  buf

  (
    g1785_p_spl_,
    g1785_p
  );


  buf

  (
    g1785_p_spl_0,
    g1785_p_spl_
  );


  buf

  (
    g1786_n_spl_,
    g1786_n
  );


  buf

  (
    g1780_n_spl_,
    g1780_n
  );


  buf

  (
    g1786_p_spl_,
    g1786_p
  );


  buf

  (
    g1780_p_spl_,
    g1780_p
  );


  buf

  (
    g1787_n_spl_,
    g1787_n
  );


  buf

  (
    g1787_n_spl_0,
    g1787_n_spl_
  );


  buf

  (
    g1787_p_spl_,
    g1787_p
  );


  buf

  (
    g1787_p_spl_0,
    g1787_p_spl_
  );


  buf

  (
    g1791_n_spl_,
    g1791_n
  );


  buf

  (
    g1790_n_spl_,
    g1790_n
  );


  buf

  (
    g1791_p_spl_,
    g1791_p
  );


  buf

  (
    g1790_p_spl_,
    g1790_p
  );


  buf

  (
    g1792_n_spl_,
    g1792_n
  );


  buf

  (
    g1792_n_spl_0,
    g1792_n_spl_
  );


  buf

  (
    g1792_p_spl_,
    g1792_p
  );


  buf

  (
    g1792_p_spl_0,
    g1792_p_spl_
  );


  buf

  (
    g1793_n_spl_,
    g1793_n
  );


  buf

  (
    g1777_n_spl_,
    g1777_n
  );


  buf

  (
    g1793_p_spl_,
    g1793_p
  );


  buf

  (
    g1777_p_spl_,
    g1777_p
  );


  buf

  (
    g1794_n_spl_,
    g1794_n
  );


  buf

  (
    g1794_n_spl_0,
    g1794_n_spl_
  );


  buf

  (
    g1794_p_spl_,
    g1794_p
  );


  buf

  (
    g1794_p_spl_0,
    g1794_p_spl_
  );


  buf

  (
    g1798_n_spl_,
    g1798_n
  );


  buf

  (
    g1797_n_spl_,
    g1797_n
  );


  buf

  (
    g1798_p_spl_,
    g1798_p
  );


  buf

  (
    g1797_p_spl_,
    g1797_p
  );


  buf

  (
    g1799_n_spl_,
    g1799_n
  );


  buf

  (
    g1799_n_spl_0,
    g1799_n_spl_
  );


  buf

  (
    g1799_p_spl_,
    g1799_p
  );


  buf

  (
    g1799_p_spl_0,
    g1799_p_spl_
  );


  buf

  (
    g1800_n_spl_,
    g1800_n
  );


  buf

  (
    g1774_n_spl_,
    g1774_n
  );


  buf

  (
    g1800_p_spl_,
    g1800_p
  );


  buf

  (
    g1774_p_spl_,
    g1774_p
  );


  buf

  (
    g1293_n_spl_,
    g1293_n
  );


  buf

  (
    g1293_n_spl_0,
    g1293_n_spl_
  );


  buf

  (
    g1293_p_spl_,
    g1293_p
  );


  buf

  (
    g1367_n_spl_,
    g1367_n
  );


  buf

  (
    g1367_n_spl_0,
    g1367_n_spl_
  );


  buf

  (
    g1367_p_spl_,
    g1367_p
  );


  buf

  (
    g1477_n_spl_,
    g1477_n
  );


  buf

  (
    g1477_n_spl_0,
    g1477_n_spl_
  );


  buf

  (
    g1477_p_spl_,
    g1477_p
  );


  buf

  (
    n2821_lo_p_spl_,
    n2821_lo_p
  );


  buf

  (
    n2821_lo_p_spl_0,
    n2821_lo_p_spl_
  );


  buf

  (
    n2821_lo_p_spl_1,
    n2821_lo_p_spl_
  );


  buf

  (
    n2821_lo_n_spl_,
    n2821_lo_n
  );


  buf

  (
    n2821_lo_n_spl_0,
    n2821_lo_n_spl_
  );


  buf

  (
    n2821_lo_n_spl_1,
    n2821_lo_n_spl_
  );


  buf

  (
    g1823_n_spl_,
    g1823_n
  );


  buf

  (
    g1822_n_spl_,
    g1822_n
  );


  buf

  (
    g1823_p_spl_,
    g1823_p
  );


  buf

  (
    g1822_p_spl_,
    g1822_p
  );


  buf

  (
    g1824_n_spl_,
    g1824_n
  );


  buf

  (
    g1824_n_spl_0,
    g1824_n_spl_
  );


  buf

  (
    g1824_p_spl_,
    g1824_p
  );


  buf

  (
    g1824_p_spl_0,
    g1824_p_spl_
  );


  buf

  (
    g1828_n_spl_,
    g1828_n
  );


  buf

  (
    g1827_n_spl_,
    g1827_n
  );


  buf

  (
    g1828_p_spl_,
    g1828_p
  );


  buf

  (
    g1827_p_spl_,
    g1827_p
  );


  buf

  (
    g1829_n_spl_,
    g1829_n
  );


  buf

  (
    g1829_n_spl_0,
    g1829_n_spl_
  );


  buf

  (
    g1829_p_spl_,
    g1829_p
  );


  buf

  (
    g1829_p_spl_0,
    g1829_p_spl_
  );


  buf

  (
    G19_p_spl_,
    G19_p
  );


  buf

  (
    G19_p_spl_0,
    G19_p_spl_
  );


  buf

  (
    G19_p_spl_00,
    G19_p_spl_0
  );


  buf

  (
    G19_p_spl_000,
    G19_p_spl_00
  );


  buf

  (
    G19_p_spl_001,
    G19_p_spl_00
  );


  buf

  (
    G19_p_spl_01,
    G19_p_spl_0
  );


  buf

  (
    G19_p_spl_010,
    G19_p_spl_01
  );


  buf

  (
    G19_p_spl_011,
    G19_p_spl_01
  );


  buf

  (
    G19_p_spl_1,
    G19_p_spl_
  );


  buf

  (
    G19_p_spl_10,
    G19_p_spl_1
  );


  buf

  (
    G19_p_spl_100,
    G19_p_spl_10
  );


  buf

  (
    G19_p_spl_11,
    G19_p_spl_1
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    G16_p_spl_0,
    G16_p_spl_
  );


  buf

  (
    G16_p_spl_1,
    G16_p_spl_
  );


  buf

  (
    G19_n_spl_,
    G19_n
  );


  buf

  (
    G19_n_spl_0,
    G19_n_spl_
  );


  buf

  (
    G19_n_spl_00,
    G19_n_spl_0
  );


  buf

  (
    G19_n_spl_000,
    G19_n_spl_00
  );


  buf

  (
    G19_n_spl_001,
    G19_n_spl_00
  );


  buf

  (
    G19_n_spl_01,
    G19_n_spl_0
  );


  buf

  (
    G19_n_spl_010,
    G19_n_spl_01
  );


  buf

  (
    G19_n_spl_011,
    G19_n_spl_01
  );


  buf

  (
    G19_n_spl_1,
    G19_n_spl_
  );


  buf

  (
    G19_n_spl_10,
    G19_n_spl_1
  );


  buf

  (
    G19_n_spl_11,
    G19_n_spl_1
  );


  buf

  (
    G16_n_spl_,
    G16_n
  );


  buf

  (
    G16_n_spl_0,
    G16_n_spl_
  );


  buf

  (
    G18_p_spl_,
    G18_p
  );


  buf

  (
    G18_p_spl_0,
    G18_p_spl_
  );


  buf

  (
    G18_p_spl_00,
    G18_p_spl_0
  );


  buf

  (
    G18_p_spl_000,
    G18_p_spl_00
  );


  buf

  (
    G18_p_spl_001,
    G18_p_spl_00
  );


  buf

  (
    G18_p_spl_01,
    G18_p_spl_0
  );


  buf

  (
    G18_p_spl_010,
    G18_p_spl_01
  );


  buf

  (
    G18_p_spl_011,
    G18_p_spl_01
  );


  buf

  (
    G18_p_spl_1,
    G18_p_spl_
  );


  buf

  (
    G18_p_spl_10,
    G18_p_spl_1
  );


  buf

  (
    G18_p_spl_100,
    G18_p_spl_10
  );


  buf

  (
    G18_p_spl_101,
    G18_p_spl_10
  );


  buf

  (
    G18_p_spl_11,
    G18_p_spl_1
  );


  buf

  (
    G18_p_spl_110,
    G18_p_spl_11
  );


  buf

  (
    G18_n_spl_,
    G18_n
  );


  buf

  (
    G18_n_spl_0,
    G18_n_spl_
  );


  buf

  (
    G18_n_spl_00,
    G18_n_spl_0
  );


  buf

  (
    G18_n_spl_000,
    G18_n_spl_00
  );


  buf

  (
    G18_n_spl_001,
    G18_n_spl_00
  );


  buf

  (
    G18_n_spl_01,
    G18_n_spl_0
  );


  buf

  (
    G18_n_spl_010,
    G18_n_spl_01
  );


  buf

  (
    G18_n_spl_011,
    G18_n_spl_01
  );


  buf

  (
    G18_n_spl_1,
    G18_n_spl_
  );


  buf

  (
    G18_n_spl_10,
    G18_n_spl_1
  );


  buf

  (
    G18_n_spl_100,
    G18_n_spl_10
  );


  buf

  (
    G18_n_spl_101,
    G18_n_spl_10
  );


  buf

  (
    G18_n_spl_11,
    G18_n_spl_1
  );


  buf

  (
    G18_n_spl_110,
    G18_n_spl_11
  );


  buf

  (
    G18_n_spl_111,
    G18_n_spl_11
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


  buf

  (
    G17_p_spl_0,
    G17_p_spl_
  );


  buf

  (
    G17_p_spl_00,
    G17_p_spl_0
  );


  buf

  (
    G17_p_spl_000,
    G17_p_spl_00
  );


  buf

  (
    G17_p_spl_001,
    G17_p_spl_00
  );


  buf

  (
    G17_p_spl_01,
    G17_p_spl_0
  );


  buf

  (
    G17_p_spl_010,
    G17_p_spl_01
  );


  buf

  (
    G17_p_spl_011,
    G17_p_spl_01
  );


  buf

  (
    G17_p_spl_1,
    G17_p_spl_
  );


  buf

  (
    G17_p_spl_10,
    G17_p_spl_1
  );


  buf

  (
    G17_p_spl_100,
    G17_p_spl_10
  );


  buf

  (
    G17_p_spl_101,
    G17_p_spl_10
  );


  buf

  (
    G17_p_spl_11,
    G17_p_spl_1
  );


  buf

  (
    G17_p_spl_110,
    G17_p_spl_11
  );


  buf

  (
    G17_p_spl_111,
    G17_p_spl_11
  );


  buf

  (
    G17_n_spl_,
    G17_n
  );


  buf

  (
    G17_n_spl_0,
    G17_n_spl_
  );


  buf

  (
    G17_n_spl_00,
    G17_n_spl_0
  );


  buf

  (
    G17_n_spl_000,
    G17_n_spl_00
  );


  buf

  (
    G17_n_spl_001,
    G17_n_spl_00
  );


  buf

  (
    G17_n_spl_01,
    G17_n_spl_0
  );


  buf

  (
    G17_n_spl_010,
    G17_n_spl_01
  );


  buf

  (
    G17_n_spl_011,
    G17_n_spl_01
  );


  buf

  (
    G17_n_spl_1,
    G17_n_spl_
  );


  buf

  (
    G17_n_spl_10,
    G17_n_spl_1
  );


  buf

  (
    G17_n_spl_100,
    G17_n_spl_10
  );


  buf

  (
    G17_n_spl_101,
    G17_n_spl_10
  );


  buf

  (
    G17_n_spl_11,
    G17_n_spl_1
  );


  buf

  (
    G17_n_spl_110,
    G17_n_spl_11
  );


  buf

  (
    G15_p_spl_,
    G15_p
  );


  buf

  (
    G15_p_spl_0,
    G15_p_spl_
  );


  buf

  (
    G15_p_spl_00,
    G15_p_spl_0
  );


  buf

  (
    G15_p_spl_1,
    G15_p_spl_
  );


  buf

  (
    G15_n_spl_,
    G15_n
  );


  buf

  (
    G15_n_spl_0,
    G15_n_spl_
  );


  buf

  (
    G15_n_spl_1,
    G15_n_spl_
  );


  buf

  (
    g1836_n_spl_,
    g1836_n
  );


  buf

  (
    g1835_p_spl_,
    g1835_p
  );


  buf

  (
    g1836_p_spl_,
    g1836_p
  );


  buf

  (
    g1835_n_spl_,
    g1835_n
  );


  buf

  (
    g1837_n_spl_,
    g1837_n
  );


  buf

  (
    g1837_p_spl_,
    g1837_p
  );


  buf

  (
    g1838_n_spl_,
    g1838_n
  );


  buf

  (
    g1838_n_spl_0,
    g1838_n_spl_
  );


  buf

  (
    g1834_n_spl_,
    g1834_n
  );


  buf

  (
    g1838_p_spl_,
    g1838_p
  );


  buf

  (
    g1838_p_spl_0,
    g1838_p_spl_
  );


  buf

  (
    g1834_p_spl_,
    g1834_p
  );


  buf

  (
    g1839_n_spl_,
    g1839_n
  );


  buf

  (
    g1839_n_spl_0,
    g1839_n_spl_
  );


  buf

  (
    g1839_p_spl_,
    g1839_p
  );


  buf

  (
    g1839_p_spl_0,
    g1839_p_spl_
  );


  buf

  (
    g1843_n_spl_,
    g1843_n
  );


  buf

  (
    g1842_n_spl_,
    g1842_n
  );


  buf

  (
    g1843_p_spl_,
    g1843_p
  );


  buf

  (
    g1842_p_spl_,
    g1842_p
  );


  buf

  (
    g1844_n_spl_,
    g1844_n
  );


  buf

  (
    g1844_n_spl_0,
    g1844_n_spl_
  );


  buf

  (
    g1844_p_spl_,
    g1844_p
  );


  buf

  (
    g1844_p_spl_0,
    g1844_p_spl_
  );


  buf

  (
    g1845_n_spl_,
    g1845_n
  );


  buf

  (
    g1833_n_spl_,
    g1833_n
  );


  buf

  (
    g1845_p_spl_,
    g1845_p
  );


  buf

  (
    g1833_p_spl_,
    g1833_p
  );


  buf

  (
    g1848_n_spl_,
    g1848_n
  );


  buf

  (
    g1847_n_spl_,
    g1847_n
  );


  buf

  (
    g1848_p_spl_,
    g1848_p
  );


  buf

  (
    g1847_p_spl_,
    g1847_p
  );


  buf

  (
    g1849_n_spl_,
    g1849_n
  );


  buf

  (
    g1849_n_spl_0,
    g1849_n_spl_
  );


  buf

  (
    g1849_p_spl_,
    g1849_p
  );


  buf

  (
    g1849_p_spl_0,
    g1849_p_spl_
  );


  buf

  (
    g1853_n_spl_,
    g1853_n
  );


  buf

  (
    g1852_n_spl_,
    g1852_n
  );


  buf

  (
    g1853_p_spl_,
    g1853_p
  );


  buf

  (
    g1852_p_spl_,
    g1852_p
  );


  buf

  (
    g1854_n_spl_,
    g1854_n
  );


  buf

  (
    g1854_n_spl_0,
    g1854_n_spl_
  );


  buf

  (
    g1854_p_spl_,
    g1854_p
  );


  buf

  (
    g1854_p_spl_0,
    g1854_p_spl_
  );


  buf

  (
    g1858_n_spl_,
    g1858_n
  );


  buf

  (
    g1857_n_spl_,
    g1857_n
  );


  buf

  (
    g1858_p_spl_,
    g1858_p
  );


  buf

  (
    g1857_p_spl_,
    g1857_p
  );


  buf

  (
    g1859_n_spl_,
    g1859_n
  );


  buf

  (
    g1859_n_spl_0,
    g1859_n_spl_
  );


  buf

  (
    g1859_p_spl_,
    g1859_p
  );


  buf

  (
    g1859_p_spl_0,
    g1859_p_spl_
  );


  buf

  (
    g1863_n_spl_,
    g1863_n
  );


  buf

  (
    g1862_n_spl_,
    g1862_n
  );


  buf

  (
    g1863_p_spl_,
    g1863_p
  );


  buf

  (
    g1862_p_spl_,
    g1862_p
  );


  buf

  (
    g1864_n_spl_,
    g1864_n
  );


  buf

  (
    g1864_n_spl_0,
    g1864_n_spl_
  );


  buf

  (
    g1864_p_spl_,
    g1864_p
  );


  buf

  (
    g1864_p_spl_0,
    g1864_p_spl_
  );


  buf

  (
    n2572_lo_buf_o2_p_spl_,
    n2572_lo_buf_o2_p
  );


  buf

  (
    n2572_lo_buf_o2_p_spl_0,
    n2572_lo_buf_o2_p_spl_
  );


  buf

  (
    n2572_lo_buf_o2_p_spl_00,
    n2572_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2572_lo_buf_o2_p_spl_01,
    n2572_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2572_lo_buf_o2_p_spl_1,
    n2572_lo_buf_o2_p_spl_
  );


  buf

  (
    n2572_lo_buf_o2_p_spl_10,
    n2572_lo_buf_o2_p_spl_1
  );


  buf

  (
    n2572_lo_buf_o2_n_spl_,
    n2572_lo_buf_o2_n
  );


  buf

  (
    n2572_lo_buf_o2_n_spl_0,
    n2572_lo_buf_o2_n_spl_
  );


  buf

  (
    n2572_lo_buf_o2_n_spl_00,
    n2572_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2572_lo_buf_o2_n_spl_1,
    n2572_lo_buf_o2_n_spl_
  );


  buf

  (
    g1871_n_spl_,
    g1871_n
  );


  buf

  (
    g1870_n_spl_,
    g1870_n
  );


  buf

  (
    g1871_p_spl_,
    g1871_p
  );


  buf

  (
    g1870_p_spl_,
    g1870_p
  );


  buf

  (
    g1872_n_spl_,
    g1872_n
  );


  buf

  (
    g1872_n_spl_0,
    g1872_n_spl_
  );


  buf

  (
    g1872_p_spl_,
    g1872_p
  );


  buf

  (
    g1872_p_spl_0,
    g1872_p_spl_
  );


  buf

  (
    G1968_o2_p_spl_,
    G1968_o2_p
  );


  buf

  (
    G1968_o2_p_spl_0,
    G1968_o2_p_spl_
  );


  buf

  (
    G1968_o2_n_spl_,
    G1968_o2_n
  );


  buf

  (
    G1968_o2_n_spl_0,
    G1968_o2_n_spl_
  );


  buf

  (
    n2560_lo_buf_o2_p_spl_,
    n2560_lo_buf_o2_p
  );


  buf

  (
    n2560_lo_buf_o2_p_spl_0,
    n2560_lo_buf_o2_p_spl_
  );


  buf

  (
    n2560_lo_buf_o2_p_spl_00,
    n2560_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2560_lo_buf_o2_p_spl_01,
    n2560_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2560_lo_buf_o2_p_spl_1,
    n2560_lo_buf_o2_p_spl_
  );


  buf

  (
    n2560_lo_buf_o2_n_spl_,
    n2560_lo_buf_o2_n
  );


  buf

  (
    n2560_lo_buf_o2_n_spl_0,
    n2560_lo_buf_o2_n_spl_
  );


  buf

  (
    n2560_lo_buf_o2_n_spl_00,
    n2560_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2560_lo_buf_o2_n_spl_1,
    n2560_lo_buf_o2_n_spl_
  );


  buf

  (
    g1879_n_spl_,
    g1879_n
  );


  buf

  (
    g1878_n_spl_,
    g1878_n
  );


  buf

  (
    g1879_p_spl_,
    g1879_p
  );


  buf

  (
    g1878_p_spl_,
    g1878_p
  );


  buf

  (
    g1880_n_spl_,
    g1880_n
  );


  buf

  (
    g1880_n_spl_0,
    g1880_n_spl_
  );


  buf

  (
    g1880_p_spl_,
    g1880_p
  );


  buf

  (
    g1880_p_spl_0,
    g1880_p_spl_
  );


  buf

  (
    g1881_n_spl_,
    g1881_n
  );


  buf

  (
    g1875_n_spl_,
    g1875_n
  );


  buf

  (
    g1881_p_spl_,
    g1881_p
  );


  buf

  (
    g1875_p_spl_,
    g1875_p
  );


  buf

  (
    g1882_n_spl_,
    g1882_n
  );


  buf

  (
    g1882_n_spl_0,
    g1882_n_spl_
  );


  buf

  (
    g1882_p_spl_,
    g1882_p
  );


  buf

  (
    g1882_p_spl_0,
    g1882_p_spl_
  );


  buf

  (
    g1886_n_spl_,
    g1886_n
  );


  buf

  (
    g1885_n_spl_,
    g1885_n
  );


  buf

  (
    g1886_p_spl_,
    g1886_p
  );


  buf

  (
    g1885_p_spl_,
    g1885_p
  );


  buf

  (
    g1887_n_spl_,
    g1887_n
  );


  buf

  (
    g1887_n_spl_0,
    g1887_n_spl_
  );


  buf

  (
    g1887_p_spl_,
    g1887_p
  );


  buf

  (
    g1887_p_spl_0,
    g1887_p_spl_
  );


  buf

  (
    G1914_o2_n_spl_,
    G1914_o2_n
  );


  buf

  (
    G1849_o2_n_spl_,
    G1849_o2_n
  );


  buf

  (
    G1914_o2_p_spl_,
    G1914_o2_p
  );


  buf

  (
    G1849_o2_p_spl_,
    G1849_o2_p
  );


  buf

  (
    g1894_n_spl_,
    g1894_n
  );


  buf

  (
    g1894_n_spl_0,
    g1894_n_spl_
  );


  buf

  (
    g1894_p_spl_,
    g1894_p
  );


  buf

  (
    g1894_p_spl_0,
    g1894_p_spl_
  );


  buf

  (
    n2548_lo_buf_o2_p_spl_,
    n2548_lo_buf_o2_p
  );


  buf

  (
    n2548_lo_buf_o2_p_spl_0,
    n2548_lo_buf_o2_p_spl_
  );


  buf

  (
    n2548_lo_buf_o2_p_spl_00,
    n2548_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2548_lo_buf_o2_p_spl_01,
    n2548_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2548_lo_buf_o2_p_spl_1,
    n2548_lo_buf_o2_p_spl_
  );


  buf

  (
    n2548_lo_buf_o2_n_spl_,
    n2548_lo_buf_o2_n
  );


  buf

  (
    n2548_lo_buf_o2_n_spl_0,
    n2548_lo_buf_o2_n_spl_
  );


  buf

  (
    n2548_lo_buf_o2_n_spl_00,
    n2548_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2548_lo_buf_o2_n_spl_1,
    n2548_lo_buf_o2_n_spl_
  );


  buf

  (
    g1898_n_spl_,
    g1898_n
  );


  buf

  (
    g1897_n_spl_,
    g1897_n
  );


  buf

  (
    g1898_p_spl_,
    g1898_p
  );


  buf

  (
    g1897_p_spl_,
    g1897_p
  );


  buf

  (
    g1899_n_spl_,
    g1899_n
  );


  buf

  (
    g1899_n_spl_0,
    g1899_n_spl_
  );


  buf

  (
    g1899_p_spl_,
    g1899_p
  );


  buf

  (
    g1899_p_spl_0,
    g1899_p_spl_
  );


  buf

  (
    g1900_n_spl_,
    g1900_n
  );


  buf

  (
    g1893_n_spl_,
    g1893_n
  );


  buf

  (
    g1900_p_spl_,
    g1900_p
  );


  buf

  (
    g1893_p_spl_,
    g1893_p
  );


  buf

  (
    g1901_n_spl_,
    g1901_n
  );


  buf

  (
    g1901_n_spl_0,
    g1901_n_spl_
  );


  buf

  (
    g1901_p_spl_,
    g1901_p
  );


  buf

  (
    g1901_p_spl_0,
    g1901_p_spl_
  );


  buf

  (
    g1905_n_spl_,
    g1905_n
  );


  buf

  (
    g1904_n_spl_,
    g1904_n
  );


  buf

  (
    g1905_p_spl_,
    g1905_p
  );


  buf

  (
    g1904_p_spl_,
    g1904_p
  );


  buf

  (
    g1906_n_spl_,
    g1906_n
  );


  buf

  (
    g1906_n_spl_0,
    g1906_n_spl_
  );


  buf

  (
    g1906_p_spl_,
    g1906_p
  );


  buf

  (
    g1906_p_spl_0,
    g1906_p_spl_
  );


  buf

  (
    g1907_n_spl_,
    g1907_n
  );


  buf

  (
    g1890_n_spl_,
    g1890_n
  );


  buf

  (
    g1907_p_spl_,
    g1907_p
  );


  buf

  (
    g1890_p_spl_,
    g1890_p
  );


  buf

  (
    g1908_n_spl_,
    g1908_n
  );


  buf

  (
    g1908_n_spl_0,
    g1908_n_spl_
  );


  buf

  (
    g1908_p_spl_,
    g1908_p
  );


  buf

  (
    g1908_p_spl_0,
    g1908_p_spl_
  );


  buf

  (
    g1912_n_spl_,
    g1912_n
  );


  buf

  (
    g1911_n_spl_,
    g1911_n
  );


  buf

  (
    g1912_p_spl_,
    g1912_p
  );


  buf

  (
    g1911_p_spl_,
    g1911_p
  );


  buf

  (
    g1913_n_spl_,
    g1913_n
  );


  buf

  (
    g1913_n_spl_0,
    g1913_n_spl_
  );


  buf

  (
    g1913_p_spl_,
    g1913_p
  );


  buf

  (
    g1913_p_spl_0,
    g1913_p_spl_
  );


  buf

  (
    G1777_o2_n_spl_,
    G1777_o2_n
  );


  buf

  (
    G1777_o2_n_spl_0,
    G1777_o2_n_spl_
  );


  buf

  (
    G1777_o2_p_spl_,
    G1777_o2_p
  );


  buf

  (
    G1777_o2_p_spl_0,
    G1777_o2_p_spl_
  );


  buf

  (
    g1924_n_spl_,
    g1924_n
  );


  buf

  (
    g1923_n_spl_,
    g1923_n
  );


  buf

  (
    g1924_p_spl_,
    g1924_p
  );


  buf

  (
    g1923_p_spl_,
    g1923_p
  );


  buf

  (
    g1925_n_spl_,
    g1925_n
  );


  buf

  (
    g1925_n_spl_0,
    g1925_n_spl_
  );


  buf

  (
    g1925_p_spl_,
    g1925_p
  );


  buf

  (
    g1925_p_spl_0,
    g1925_p_spl_
  );


  buf

  (
    n2536_lo_buf_o2_p_spl_,
    n2536_lo_buf_o2_p
  );


  buf

  (
    n2536_lo_buf_o2_p_spl_0,
    n2536_lo_buf_o2_p_spl_
  );


  buf

  (
    n2536_lo_buf_o2_p_spl_00,
    n2536_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2536_lo_buf_o2_p_spl_01,
    n2536_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2536_lo_buf_o2_p_spl_1,
    n2536_lo_buf_o2_p_spl_
  );


  buf

  (
    n2536_lo_buf_o2_n_spl_,
    n2536_lo_buf_o2_n
  );


  buf

  (
    n2536_lo_buf_o2_n_spl_0,
    n2536_lo_buf_o2_n_spl_
  );


  buf

  (
    n2536_lo_buf_o2_n_spl_00,
    n2536_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2536_lo_buf_o2_n_spl_1,
    n2536_lo_buf_o2_n_spl_
  );


  buf

  (
    g1929_n_spl_,
    g1929_n
  );


  buf

  (
    g1928_n_spl_,
    g1928_n
  );


  buf

  (
    g1929_p_spl_,
    g1929_p
  );


  buf

  (
    g1928_p_spl_,
    g1928_p
  );


  buf

  (
    g1930_n_spl_,
    g1930_n
  );


  buf

  (
    g1930_n_spl_0,
    g1930_n_spl_
  );


  buf

  (
    g1930_p_spl_,
    g1930_p
  );


  buf

  (
    g1930_p_spl_0,
    g1930_p_spl_
  );


  buf

  (
    g1931_n_spl_,
    g1931_n
  );


  buf

  (
    g1922_n_spl_,
    g1922_n
  );


  buf

  (
    g1931_p_spl_,
    g1931_p
  );


  buf

  (
    g1922_p_spl_,
    g1922_p
  );


  buf

  (
    g1932_n_spl_,
    g1932_n
  );


  buf

  (
    g1932_n_spl_0,
    g1932_n_spl_
  );


  buf

  (
    g1932_p_spl_,
    g1932_p
  );


  buf

  (
    g1932_p_spl_0,
    g1932_p_spl_
  );


  buf

  (
    g1936_n_spl_,
    g1936_n
  );


  buf

  (
    g1935_n_spl_,
    g1935_n
  );


  buf

  (
    g1936_p_spl_,
    g1936_p
  );


  buf

  (
    g1935_p_spl_,
    g1935_p
  );


  buf

  (
    g1937_n_spl_,
    g1937_n
  );


  buf

  (
    g1937_n_spl_0,
    g1937_n_spl_
  );


  buf

  (
    g1937_p_spl_,
    g1937_p
  );


  buf

  (
    g1937_p_spl_0,
    g1937_p_spl_
  );


  buf

  (
    g1938_n_spl_,
    g1938_n
  );


  buf

  (
    g1919_n_spl_,
    g1919_n
  );


  buf

  (
    g1938_p_spl_,
    g1938_p
  );


  buf

  (
    g1919_p_spl_,
    g1919_p
  );


  buf

  (
    g1939_n_spl_,
    g1939_n
  );


  buf

  (
    g1939_n_spl_0,
    g1939_n_spl_
  );


  buf

  (
    g1939_p_spl_,
    g1939_p
  );


  buf

  (
    g1939_p_spl_0,
    g1939_p_spl_
  );


  buf

  (
    g1943_n_spl_,
    g1943_n
  );


  buf

  (
    g1942_n_spl_,
    g1942_n
  );


  buf

  (
    g1943_p_spl_,
    g1943_p
  );


  buf

  (
    g1942_p_spl_,
    g1942_p
  );


  buf

  (
    g1944_n_spl_,
    g1944_n
  );


  buf

  (
    g1944_n_spl_0,
    g1944_n_spl_
  );


  buf

  (
    g1944_p_spl_,
    g1944_p
  );


  buf

  (
    g1944_p_spl_0,
    g1944_p_spl_
  );


  buf

  (
    g1945_n_spl_,
    g1945_n
  );


  buf

  (
    g1916_n_spl_,
    g1916_n
  );


  buf

  (
    g1945_p_spl_,
    g1945_p
  );


  buf

  (
    g1916_p_spl_,
    g1916_p
  );


  buf

  (
    g1946_n_spl_,
    g1946_n
  );


  buf

  (
    g1946_n_spl_0,
    g1946_n_spl_
  );


  buf

  (
    g1946_p_spl_,
    g1946_p
  );


  buf

  (
    g1946_p_spl_0,
    g1946_p_spl_
  );


  buf

  (
    g1950_n_spl_,
    g1950_n
  );


  buf

  (
    g1949_n_spl_,
    g1949_n
  );


  buf

  (
    g1950_p_spl_,
    g1950_p
  );


  buf

  (
    g1949_p_spl_,
    g1949_p
  );


  buf

  (
    g1951_n_spl_,
    g1951_n
  );


  buf

  (
    g1951_n_spl_0,
    g1951_n_spl_
  );


  buf

  (
    g1951_p_spl_,
    g1951_p
  );


  buf

  (
    g1951_p_spl_0,
    g1951_p_spl_
  );


  buf

  (
    g1967_n_spl_,
    g1967_n
  );


  buf

  (
    g1966_n_spl_,
    g1966_n
  );


  buf

  (
    g1967_p_spl_,
    g1967_p
  );


  buf

  (
    g1966_p_spl_,
    g1966_p
  );


  buf

  (
    g1968_n_spl_,
    g1968_n
  );


  buf

  (
    g1968_n_spl_0,
    g1968_n_spl_
  );


  buf

  (
    g1968_p_spl_,
    g1968_p
  );


  buf

  (
    g1968_p_spl_0,
    g1968_p_spl_
  );


  buf

  (
    n2524_lo_buf_o2_p_spl_,
    n2524_lo_buf_o2_p
  );


  buf

  (
    n2524_lo_buf_o2_p_spl_0,
    n2524_lo_buf_o2_p_spl_
  );


  buf

  (
    n2524_lo_buf_o2_p_spl_00,
    n2524_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2524_lo_buf_o2_p_spl_1,
    n2524_lo_buf_o2_p_spl_
  );


  buf

  (
    n2524_lo_buf_o2_n_spl_,
    n2524_lo_buf_o2_n
  );


  buf

  (
    n2524_lo_buf_o2_n_spl_0,
    n2524_lo_buf_o2_n_spl_
  );


  buf

  (
    n2524_lo_buf_o2_n_spl_00,
    n2524_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2524_lo_buf_o2_n_spl_1,
    n2524_lo_buf_o2_n_spl_
  );


  buf

  (
    g1972_n_spl_,
    g1972_n
  );


  buf

  (
    g1971_n_spl_,
    g1971_n
  );


  buf

  (
    g1972_p_spl_,
    g1972_p
  );


  buf

  (
    g1971_p_spl_,
    g1971_p
  );


  buf

  (
    g1973_n_spl_,
    g1973_n
  );


  buf

  (
    g1973_n_spl_0,
    g1973_n_spl_
  );


  buf

  (
    g1973_p_spl_,
    g1973_p
  );


  buf

  (
    g1973_p_spl_0,
    g1973_p_spl_
  );


  buf

  (
    g1974_n_spl_,
    g1974_n
  );


  buf

  (
    g1963_n_spl_,
    g1963_n
  );


  buf

  (
    g1974_p_spl_,
    g1974_p
  );


  buf

  (
    g1963_p_spl_,
    g1963_p
  );


  buf

  (
    g1975_n_spl_,
    g1975_n
  );


  buf

  (
    g1975_n_spl_0,
    g1975_n_spl_
  );


  buf

  (
    g1975_p_spl_,
    g1975_p
  );


  buf

  (
    g1975_p_spl_0,
    g1975_p_spl_
  );


  buf

  (
    g1979_n_spl_,
    g1979_n
  );


  buf

  (
    g1978_n_spl_,
    g1978_n
  );


  buf

  (
    g1979_p_spl_,
    g1979_p
  );


  buf

  (
    g1978_p_spl_,
    g1978_p
  );


  buf

  (
    g1980_n_spl_,
    g1980_n
  );


  buf

  (
    g1980_n_spl_0,
    g1980_n_spl_
  );


  buf

  (
    g1980_p_spl_,
    g1980_p
  );


  buf

  (
    g1980_p_spl_0,
    g1980_p_spl_
  );


  buf

  (
    g1981_n_spl_,
    g1981_n
  );


  buf

  (
    g1960_n_spl_,
    g1960_n
  );


  buf

  (
    g1981_p_spl_,
    g1981_p
  );


  buf

  (
    g1960_p_spl_,
    g1960_p
  );


  buf

  (
    g1982_n_spl_,
    g1982_n
  );


  buf

  (
    g1982_n_spl_0,
    g1982_n_spl_
  );


  buf

  (
    g1982_p_spl_,
    g1982_p
  );


  buf

  (
    g1982_p_spl_0,
    g1982_p_spl_
  );


  buf

  (
    g1986_n_spl_,
    g1986_n
  );


  buf

  (
    g1985_n_spl_,
    g1985_n
  );


  buf

  (
    g1986_p_spl_,
    g1986_p
  );


  buf

  (
    g1985_p_spl_,
    g1985_p
  );


  buf

  (
    g1987_n_spl_,
    g1987_n
  );


  buf

  (
    g1987_n_spl_0,
    g1987_n_spl_
  );


  buf

  (
    g1987_p_spl_,
    g1987_p
  );


  buf

  (
    g1987_p_spl_0,
    g1987_p_spl_
  );


  buf

  (
    g1988_n_spl_,
    g1988_n
  );


  buf

  (
    g1957_n_spl_,
    g1957_n
  );


  buf

  (
    g1988_p_spl_,
    g1988_p
  );


  buf

  (
    g1957_p_spl_,
    g1957_p
  );


  buf

  (
    g1989_n_spl_,
    g1989_n
  );


  buf

  (
    g1989_n_spl_0,
    g1989_n_spl_
  );


  buf

  (
    g1989_p_spl_,
    g1989_p
  );


  buf

  (
    g1989_p_spl_0,
    g1989_p_spl_
  );


  buf

  (
    g1993_n_spl_,
    g1993_n
  );


  buf

  (
    g1992_n_spl_,
    g1992_n
  );


  buf

  (
    g1993_p_spl_,
    g1993_p
  );


  buf

  (
    g1992_p_spl_,
    g1992_p
  );


  buf

  (
    g1994_n_spl_,
    g1994_n
  );


  buf

  (
    g1994_n_spl_0,
    g1994_n_spl_
  );


  buf

  (
    g1994_p_spl_,
    g1994_p
  );


  buf

  (
    g1994_p_spl_0,
    g1994_p_spl_
  );


  buf

  (
    G2250_o2_n_spl_,
    G2250_o2_n
  );


  buf

  (
    G2198_o2_n_spl_,
    G2198_o2_n
  );


  buf

  (
    G2250_o2_p_spl_,
    G2250_o2_p
  );


  buf

  (
    G2198_o2_p_spl_,
    G2198_o2_p
  );


  buf

  (
    g2003_n_spl_,
    g2003_n
  );


  buf

  (
    g2003_n_spl_0,
    g2003_n_spl_
  );


  buf

  (
    g2003_p_spl_,
    g2003_p
  );


  buf

  (
    g2003_p_spl_0,
    g2003_p_spl_
  );


  buf

  (
    n2608_lo_buf_o2_p_spl_,
    n2608_lo_buf_o2_p
  );


  buf

  (
    n2608_lo_buf_o2_p_spl_0,
    n2608_lo_buf_o2_p_spl_
  );


  buf

  (
    n2608_lo_buf_o2_p_spl_00,
    n2608_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2608_lo_buf_o2_p_spl_1,
    n2608_lo_buf_o2_p_spl_
  );


  buf

  (
    n2608_lo_buf_o2_n_spl_,
    n2608_lo_buf_o2_n
  );


  buf

  (
    n2608_lo_buf_o2_n_spl_0,
    n2608_lo_buf_o2_n_spl_
  );


  buf

  (
    n2608_lo_buf_o2_n_spl_1,
    n2608_lo_buf_o2_n_spl_
  );


  buf

  (
    g2007_n_spl_,
    g2007_n
  );


  buf

  (
    g2006_n_spl_,
    g2006_n
  );


  buf

  (
    g2007_p_spl_,
    g2007_p
  );


  buf

  (
    g2006_p_spl_,
    g2006_p
  );


  buf

  (
    g2008_n_spl_,
    g2008_n
  );


  buf

  (
    g2008_n_spl_0,
    g2008_n_spl_
  );


  buf

  (
    g2008_p_spl_,
    g2008_p
  );


  buf

  (
    g2008_p_spl_0,
    g2008_p_spl_
  );


  buf

  (
    g2009_n_spl_,
    g2009_n
  );


  buf

  (
    g2002_n_spl_,
    g2002_n
  );


  buf

  (
    g2009_p_spl_,
    g2009_p
  );


  buf

  (
    g2002_p_spl_,
    g2002_p
  );


  buf

  (
    g2010_n_spl_,
    g2010_n
  );


  buf

  (
    g2010_n_spl_0,
    g2010_n_spl_
  );


  buf

  (
    g2010_p_spl_,
    g2010_p
  );


  buf

  (
    g2010_p_spl_0,
    g2010_p_spl_
  );


  buf

  (
    g2014_n_spl_,
    g2014_n
  );


  buf

  (
    g2013_n_spl_,
    g2013_n
  );


  buf

  (
    g2014_p_spl_,
    g2014_p
  );


  buf

  (
    g2013_p_spl_,
    g2013_p
  );


  buf

  (
    g2015_n_spl_,
    g2015_n
  );


  buf

  (
    g2015_n_spl_0,
    g2015_n_spl_
  );


  buf

  (
    g2015_p_spl_,
    g2015_p
  );


  buf

  (
    g2015_p_spl_0,
    g2015_p_spl_
  );


  buf

  (
    g2016_n_spl_,
    g2016_n
  );


  buf

  (
    g1999_n_spl_,
    g1999_n
  );


  buf

  (
    g2016_p_spl_,
    g2016_p
  );


  buf

  (
    g1999_p_spl_,
    g1999_p
  );


  buf

  (
    g2017_n_spl_,
    g2017_n
  );


  buf

  (
    g2017_n_spl_0,
    g2017_n_spl_
  );


  buf

  (
    g2017_p_spl_,
    g2017_p
  );


  buf

  (
    g2017_p_spl_0,
    g2017_p_spl_
  );


  buf

  (
    g2021_n_spl_,
    g2021_n
  );


  buf

  (
    g2020_n_spl_,
    g2020_n
  );


  buf

  (
    g2021_p_spl_,
    g2021_p
  );


  buf

  (
    g2020_p_spl_,
    g2020_p
  );


  buf

  (
    g2022_n_spl_,
    g2022_n
  );


  buf

  (
    g2022_n_spl_0,
    g2022_n_spl_
  );


  buf

  (
    g2022_p_spl_,
    g2022_p
  );


  buf

  (
    g2022_p_spl_0,
    g2022_p_spl_
  );


  buf

  (
    G2118_o2_n_spl_,
    G2118_o2_n
  );


  buf

  (
    G2118_o2_n_spl_0,
    G2118_o2_n_spl_
  );


  buf

  (
    G2118_o2_p_spl_,
    G2118_o2_p
  );


  buf

  (
    G2118_o2_p_spl_0,
    G2118_o2_p_spl_
  );


  buf

  (
    g2033_n_spl_,
    g2033_n
  );


  buf

  (
    g2032_n_spl_,
    g2032_n
  );


  buf

  (
    g2033_p_spl_,
    g2033_p
  );


  buf

  (
    g2032_p_spl_,
    g2032_p
  );


  buf

  (
    g2034_n_spl_,
    g2034_n
  );


  buf

  (
    g2034_n_spl_0,
    g2034_n_spl_
  );


  buf

  (
    g2034_p_spl_,
    g2034_p
  );


  buf

  (
    g2034_p_spl_0,
    g2034_p_spl_
  );


  buf

  (
    n2596_lo_buf_o2_p_spl_,
    n2596_lo_buf_o2_p
  );


  buf

  (
    n2596_lo_buf_o2_p_spl_0,
    n2596_lo_buf_o2_p_spl_
  );


  buf

  (
    n2596_lo_buf_o2_p_spl_00,
    n2596_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2596_lo_buf_o2_p_spl_1,
    n2596_lo_buf_o2_p_spl_
  );


  buf

  (
    n2596_lo_buf_o2_n_spl_,
    n2596_lo_buf_o2_n
  );


  buf

  (
    n2596_lo_buf_o2_n_spl_0,
    n2596_lo_buf_o2_n_spl_
  );


  buf

  (
    n2596_lo_buf_o2_n_spl_1,
    n2596_lo_buf_o2_n_spl_
  );


  buf

  (
    g2038_n_spl_,
    g2038_n
  );


  buf

  (
    g2037_n_spl_,
    g2037_n
  );


  buf

  (
    g2038_p_spl_,
    g2038_p
  );


  buf

  (
    g2037_p_spl_,
    g2037_p
  );


  buf

  (
    g2039_n_spl_,
    g2039_n
  );


  buf

  (
    g2039_n_spl_0,
    g2039_n_spl_
  );


  buf

  (
    g2039_p_spl_,
    g2039_p
  );


  buf

  (
    g2039_p_spl_0,
    g2039_p_spl_
  );


  buf

  (
    g2040_n_spl_,
    g2040_n
  );


  buf

  (
    g2031_n_spl_,
    g2031_n
  );


  buf

  (
    g2040_p_spl_,
    g2040_p
  );


  buf

  (
    g2031_p_spl_,
    g2031_p
  );


  buf

  (
    g2041_n_spl_,
    g2041_n
  );


  buf

  (
    g2041_n_spl_0,
    g2041_n_spl_
  );


  buf

  (
    g2041_p_spl_,
    g2041_p
  );


  buf

  (
    g2041_p_spl_0,
    g2041_p_spl_
  );


  buf

  (
    g2045_n_spl_,
    g2045_n
  );


  buf

  (
    g2044_n_spl_,
    g2044_n
  );


  buf

  (
    g2045_p_spl_,
    g2045_p
  );


  buf

  (
    g2044_p_spl_,
    g2044_p
  );


  buf

  (
    g2046_n_spl_,
    g2046_n
  );


  buf

  (
    g2046_n_spl_0,
    g2046_n_spl_
  );


  buf

  (
    g2046_p_spl_,
    g2046_p
  );


  buf

  (
    g2046_p_spl_0,
    g2046_p_spl_
  );


  buf

  (
    g2047_n_spl_,
    g2047_n
  );


  buf

  (
    g2028_n_spl_,
    g2028_n
  );


  buf

  (
    g2047_p_spl_,
    g2047_p
  );


  buf

  (
    g2028_p_spl_,
    g2028_p
  );


  buf

  (
    g2048_n_spl_,
    g2048_n
  );


  buf

  (
    g2048_n_spl_0,
    g2048_n_spl_
  );


  buf

  (
    g2048_p_spl_,
    g2048_p
  );


  buf

  (
    g2048_p_spl_0,
    g2048_p_spl_
  );


  buf

  (
    g2052_n_spl_,
    g2052_n
  );


  buf

  (
    g2051_n_spl_,
    g2051_n
  );


  buf

  (
    g2052_p_spl_,
    g2052_p
  );


  buf

  (
    g2051_p_spl_,
    g2051_p
  );


  buf

  (
    g2053_n_spl_,
    g2053_n
  );


  buf

  (
    g2053_n_spl_0,
    g2053_n_spl_
  );


  buf

  (
    g2053_p_spl_,
    g2053_p
  );


  buf

  (
    g2053_p_spl_0,
    g2053_p_spl_
  );


  buf

  (
    g2054_n_spl_,
    g2054_n
  );


  buf

  (
    g2025_n_spl_,
    g2025_n
  );


  buf

  (
    g2054_p_spl_,
    g2054_p
  );


  buf

  (
    g2025_p_spl_,
    g2025_p
  );


  buf

  (
    g2055_n_spl_,
    g2055_n
  );


  buf

  (
    g2055_n_spl_0,
    g2055_n_spl_
  );


  buf

  (
    g2055_p_spl_,
    g2055_p
  );


  buf

  (
    g2055_p_spl_0,
    g2055_p_spl_
  );


  buf

  (
    n2758_lo_p_spl_,
    n2758_lo_p
  );


  buf

  (
    n2758_lo_p_spl_0,
    n2758_lo_p_spl_
  );


  buf

  (
    n2758_lo_p_spl_00,
    n2758_lo_p_spl_0
  );


  buf

  (
    n2758_lo_p_spl_000,
    n2758_lo_p_spl_00
  );


  buf

  (
    n2758_lo_p_spl_001,
    n2758_lo_p_spl_00
  );


  buf

  (
    n2758_lo_p_spl_01,
    n2758_lo_p_spl_0
  );


  buf

  (
    n2758_lo_p_spl_1,
    n2758_lo_p_spl_
  );


  buf

  (
    n2758_lo_p_spl_10,
    n2758_lo_p_spl_1
  );


  buf

  (
    n2758_lo_p_spl_11,
    n2758_lo_p_spl_1
  );


  buf

  (
    n2758_lo_n_spl_,
    n2758_lo_n
  );


  buf

  (
    n2758_lo_n_spl_0,
    n2758_lo_n_spl_
  );


  buf

  (
    n2758_lo_n_spl_00,
    n2758_lo_n_spl_0
  );


  buf

  (
    n2758_lo_n_spl_000,
    n2758_lo_n_spl_00
  );


  buf

  (
    n2758_lo_n_spl_001,
    n2758_lo_n_spl_00
  );


  buf

  (
    n2758_lo_n_spl_01,
    n2758_lo_n_spl_0
  );


  buf

  (
    n2758_lo_n_spl_1,
    n2758_lo_n_spl_
  );


  buf

  (
    n2758_lo_n_spl_10,
    n2758_lo_n_spl_1
  );


  buf

  (
    n2758_lo_n_spl_11,
    n2758_lo_n_spl_1
  );


  buf

  (
    g2059_n_spl_,
    g2059_n
  );


  buf

  (
    g2058_n_spl_,
    g2058_n
  );


  buf

  (
    g2059_p_spl_,
    g2059_p
  );


  buf

  (
    g2058_p_spl_,
    g2058_p
  );


  buf

  (
    g2060_n_spl_,
    g2060_n
  );


  buf

  (
    g2060_n_spl_0,
    g2060_n_spl_
  );


  buf

  (
    g2060_p_spl_,
    g2060_p
  );


  buf

  (
    g2060_p_spl_0,
    g2060_p_spl_
  );


  buf

  (
    G2058_o2_p_spl_,
    G2058_o2_p
  );


  buf

  (
    G935_o2_n_spl_,
    G935_o2_n
  );


  buf

  (
    G2058_o2_n_spl_,
    G2058_o2_n
  );


  buf

  (
    G935_o2_p_spl_,
    G935_o2_p
  );


  buf

  (
    g2076_n_spl_,
    g2076_n
  );


  buf

  (
    g2076_n_spl_0,
    g2076_n_spl_
  );


  buf

  (
    g2076_p_spl_,
    g2076_p
  );


  buf

  (
    g2076_p_spl_0,
    g2076_p_spl_
  );


  buf

  (
    g2077_n_spl_,
    g2077_n
  );


  buf

  (
    g2075_n_spl_,
    g2075_n
  );


  buf

  (
    g2077_p_spl_,
    g2077_p
  );


  buf

  (
    g2075_p_spl_,
    g2075_p
  );


  buf

  (
    g2078_n_spl_,
    g2078_n
  );


  buf

  (
    g2078_n_spl_0,
    g2078_n_spl_
  );


  buf

  (
    g2078_p_spl_,
    g2078_p
  );


  buf

  (
    g2078_p_spl_0,
    g2078_p_spl_
  );


  buf

  (
    n2584_lo_buf_o2_p_spl_,
    n2584_lo_buf_o2_p
  );


  buf

  (
    n2584_lo_buf_o2_p_spl_0,
    n2584_lo_buf_o2_p_spl_
  );


  buf

  (
    n2584_lo_buf_o2_p_spl_00,
    n2584_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2584_lo_buf_o2_p_spl_1,
    n2584_lo_buf_o2_p_spl_
  );


  buf

  (
    n2584_lo_buf_o2_n_spl_,
    n2584_lo_buf_o2_n
  );


  buf

  (
    n2584_lo_buf_o2_n_spl_0,
    n2584_lo_buf_o2_n_spl_
  );


  buf

  (
    n2584_lo_buf_o2_n_spl_00,
    n2584_lo_buf_o2_n_spl_0
  );


  buf

  (
    n2584_lo_buf_o2_n_spl_1,
    n2584_lo_buf_o2_n_spl_
  );


  buf

  (
    g2082_n_spl_,
    g2082_n
  );


  buf

  (
    g2081_n_spl_,
    g2081_n
  );


  buf

  (
    g2082_p_spl_,
    g2082_p
  );


  buf

  (
    g2081_p_spl_,
    g2081_p
  );


  buf

  (
    g2083_n_spl_,
    g2083_n
  );


  buf

  (
    g2083_n_spl_0,
    g2083_n_spl_
  );


  buf

  (
    g2083_p_spl_,
    g2083_p
  );


  buf

  (
    g2083_p_spl_0,
    g2083_p_spl_
  );


  buf

  (
    g2084_n_spl_,
    g2084_n
  );


  buf

  (
    g2072_n_spl_,
    g2072_n
  );


  buf

  (
    g2084_p_spl_,
    g2084_p
  );


  buf

  (
    g2072_p_spl_,
    g2072_p
  );


  buf

  (
    g2085_n_spl_,
    g2085_n
  );


  buf

  (
    g2085_n_spl_0,
    g2085_n_spl_
  );


  buf

  (
    g2085_p_spl_,
    g2085_p
  );


  buf

  (
    g2085_p_spl_0,
    g2085_p_spl_
  );


  buf

  (
    g2089_n_spl_,
    g2089_n
  );


  buf

  (
    g2088_n_spl_,
    g2088_n
  );


  buf

  (
    g2089_p_spl_,
    g2089_p
  );


  buf

  (
    g2088_p_spl_,
    g2088_p
  );


  buf

  (
    g2090_n_spl_,
    g2090_n
  );


  buf

  (
    g2090_n_spl_0,
    g2090_n_spl_
  );


  buf

  (
    g2090_p_spl_,
    g2090_p
  );


  buf

  (
    g2090_p_spl_0,
    g2090_p_spl_
  );


  buf

  (
    g2091_n_spl_,
    g2091_n
  );


  buf

  (
    g2069_n_spl_,
    g2069_n
  );


  buf

  (
    g2091_p_spl_,
    g2091_p
  );


  buf

  (
    g2069_p_spl_,
    g2069_p
  );


  buf

  (
    g2092_n_spl_,
    g2092_n
  );


  buf

  (
    g2092_n_spl_0,
    g2092_n_spl_
  );


  buf

  (
    g2092_p_spl_,
    g2092_p
  );


  buf

  (
    g2092_p_spl_0,
    g2092_p_spl_
  );


  buf

  (
    g2096_n_spl_,
    g2096_n
  );


  buf

  (
    g2095_n_spl_,
    g2095_n
  );


  buf

  (
    g2096_p_spl_,
    g2096_p
  );


  buf

  (
    g2095_p_spl_,
    g2095_p
  );


  buf

  (
    g2097_n_spl_,
    g2097_n
  );


  buf

  (
    g2097_n_spl_0,
    g2097_n_spl_
  );


  buf

  (
    g2097_p_spl_,
    g2097_p
  );


  buf

  (
    g2097_p_spl_0,
    g2097_p_spl_
  );


  buf

  (
    g2098_n_spl_,
    g2098_n
  );


  buf

  (
    g2066_n_spl_,
    g2066_n
  );


  buf

  (
    g2098_p_spl_,
    g2098_p
  );


  buf

  (
    g2066_p_spl_,
    g2066_p
  );


  buf

  (
    g2099_n_spl_,
    g2099_n
  );


  buf

  (
    g2099_n_spl_0,
    g2099_n_spl_
  );


  buf

  (
    g2099_p_spl_,
    g2099_p
  );


  buf

  (
    g2099_p_spl_0,
    g2099_p_spl_
  );


  buf

  (
    g2103_n_spl_,
    g2103_n
  );


  buf

  (
    g2102_n_spl_,
    g2102_n
  );


  buf

  (
    g2103_p_spl_,
    g2103_p
  );


  buf

  (
    g2102_p_spl_,
    g2102_p
  );


  buf

  (
    g2104_n_spl_,
    g2104_n
  );


  buf

  (
    g2104_n_spl_0,
    g2104_n_spl_
  );


  buf

  (
    g2104_p_spl_,
    g2104_p
  );


  buf

  (
    g2104_p_spl_0,
    g2104_p_spl_
  );


  buf

  (
    g2110_n_spl_,
    g2110_n
  );


  buf

  (
    g2109_n_spl_,
    g2109_n
  );


  buf

  (
    g2110_p_spl_,
    g2110_p
  );


  buf

  (
    g2109_p_spl_,
    g2109_p
  );


  buf

  (
    g2111_n_spl_,
    g2111_n
  );


  buf

  (
    g2111_n_spl_0,
    g2111_n_spl_
  );


  buf

  (
    g2111_p_spl_,
    g2111_p
  );


  buf

  (
    g2111_p_spl_0,
    g2111_p_spl_
  );


  buf

  (
    g2115_n_spl_,
    g2115_n
  );


  buf

  (
    g2114_n_spl_,
    g2114_n
  );


  buf

  (
    g2115_p_spl_,
    g2115_p
  );


  buf

  (
    g2114_p_spl_,
    g2114_p
  );


  buf

  (
    g2116_n_spl_,
    g2116_n
  );


  buf

  (
    g2116_n_spl_0,
    g2116_n_spl_
  );


  buf

  (
    g2116_p_spl_,
    g2116_p
  );


  buf

  (
    g2116_p_spl_0,
    g2116_p_spl_
  );


  buf

  (
    g2120_n_spl_,
    g2120_n
  );


  buf

  (
    g2119_n_spl_,
    g2119_n
  );


  buf

  (
    g2120_p_spl_,
    g2120_p
  );


  buf

  (
    g2119_p_spl_,
    g2119_p
  );


  buf

  (
    g2121_n_spl_,
    g2121_n
  );


  buf

  (
    g2121_n_spl_0,
    g2121_n_spl_
  );


  buf

  (
    g2121_p_spl_,
    g2121_p
  );


  buf

  (
    g2121_p_spl_0,
    g2121_p_spl_
  );


  buf

  (
    g2125_n_spl_,
    g2125_n
  );


  buf

  (
    g2124_n_spl_,
    g2124_n
  );


  buf

  (
    g2125_p_spl_,
    g2125_p
  );


  buf

  (
    g2124_p_spl_,
    g2124_p
  );


  buf

  (
    g2126_n_spl_,
    g2126_n
  );


  buf

  (
    g2126_n_spl_0,
    g2126_n_spl_
  );


  buf

  (
    g2126_p_spl_,
    g2126_p
  );


  buf

  (
    g2126_p_spl_0,
    g2126_p_spl_
  );


  buf

  (
    g1508_p_spl_,
    g1508_p
  );


  buf

  (
    g2130_n_spl_,
    g2130_n
  );


  buf

  (
    g2129_n_spl_,
    g2129_n
  );


  buf

  (
    g2131_n_spl_,
    g2131_n
  );


  buf

  (
    g1563_n_spl_,
    g1563_n
  );


  buf

  (
    g1563_n_spl_0,
    g1563_n_spl_
  );


  buf

  (
    g1578_n_spl_,
    g1578_n
  );


  buf

  (
    g1578_n_spl_0,
    g1578_n_spl_
  );


  buf

  (
    g1593_n_spl_,
    g1593_n
  );


  buf

  (
    g1593_n_spl_0,
    g1593_n_spl_
  );


  buf

  (
    g1602_n_spl_,
    g1602_n
  );


  buf

  (
    g1545_n_spl_,
    g1545_n
  );


  buf

  (
    g1599_n_spl_,
    g1599_n
  );


  buf

  (
    g1546_n_spl_,
    g1546_n
  );


  buf

  (
    g1596_n_spl_,
    g1596_n
  );


  buf

  (
    g1547_n_spl_,
    g1547_n
  );


  buf

  (
    g1605_n_spl_,
    g1605_n
  );


  buf

  (
    g1548_n_spl_,
    g1548_n
  );


  buf

  (
    g1220_n_spl_,
    g1220_n
  );


  buf

  (
    g1220_n_spl_0,
    g1220_n_spl_
  );


  buf

  (
    g1225_n_spl_,
    g1225_n
  );


  buf

  (
    g1225_n_spl_0,
    g1225_n_spl_
  );


  buf

  (
    g1230_n_spl_,
    g1230_n
  );


  buf

  (
    g1230_n_spl_0,
    g1230_n_spl_
  );


  buf

  (
    g2167_n_spl_,
    g2167_n
  );


  buf

  (
    g2166_n_spl_,
    g2166_n
  );


  buf

  (
    g2167_p_spl_,
    g2167_p
  );


  buf

  (
    g2166_p_spl_,
    g2166_p
  );


  buf

  (
    g2168_n_spl_,
    g2168_n
  );


  buf

  (
    g2168_n_spl_0,
    g2168_n_spl_
  );


  buf

  (
    g2168_p_spl_,
    g2168_p
  );


  buf

  (
    g2172_n_spl_,
    g2172_n
  );


  buf

  (
    g2171_n_spl_,
    g2171_n
  );


  buf

  (
    g2172_p_spl_,
    g2172_p
  );


  buf

  (
    g2171_p_spl_,
    g2171_p
  );


  buf

  (
    g2173_n_spl_,
    g2173_n
  );


  buf

  (
    g2173_n_spl_0,
    g2173_n_spl_
  );


  buf

  (
    g2173_p_spl_,
    g2173_p
  );


  buf

  (
    g2182_n_spl_,
    g2182_n
  );


  buf

  (
    g2181_n_spl_,
    g2181_n
  );


  buf

  (
    g2182_p_spl_,
    g2182_p
  );


  buf

  (
    g2181_p_spl_,
    g2181_p
  );


  buf

  (
    g2183_n_spl_,
    g2183_n
  );


  buf

  (
    g2183_n_spl_0,
    g2183_n_spl_
  );


  buf

  (
    g2183_p_spl_,
    g2183_p
  );


  buf

  (
    g2187_n_spl_,
    g2187_n
  );


  buf

  (
    g2186_n_spl_,
    g2186_n
  );


  buf

  (
    g2187_p_spl_,
    g2187_p
  );


  buf

  (
    g2186_p_spl_,
    g2186_p
  );


  buf

  (
    g2188_n_spl_,
    g2188_n
  );


  buf

  (
    g2188_n_spl_0,
    g2188_n_spl_
  );


  buf

  (
    g2188_p_spl_,
    g2188_p
  );


  buf

  (
    g1606_p_spl_,
    g1606_p
  );


  buf

  (
    g1619_n_spl_,
    g1619_n
  );


  buf

  (
    g1619_n_spl_0,
    g1619_n_spl_
  );


  buf

  (
    g1644_n_spl_,
    g1644_n
  );


  buf

  (
    g1644_n_spl_0,
    g1644_n_spl_
  );


  buf

  (
    g1669_n_spl_,
    g1669_n
  );


  buf

  (
    g1669_n_spl_0,
    g1669_n_spl_
  );


  buf

  (
    g1724_n_spl_,
    g1724_n
  );


  buf

  (
    g1724_n_spl_0,
    g1724_n_spl_
  );


  buf

  (
    g1801_n_spl_,
    g1801_n
  );


  buf

  (
    g1801_n_spl_0,
    g1801_n_spl_
  );


  buf

  (
    g1801_p_spl_,
    g1801_p
  );


  buf

  (
    g2134_n_spl_,
    g2134_n
  );


  buf

  (
    g1832_n_spl_,
    g1832_n
  );


  buf

  (
    g2226_n_spl_,
    g2226_n
  );


  buf

  (
    g2225_n_spl_,
    g2225_n
  );


  buf

  (
    g2226_p_spl_,
    g2226_p
  );


  buf

  (
    g2225_p_spl_,
    g2225_p
  );


  buf

  (
    g2227_n_spl_,
    g2227_n
  );


  buf

  (
    g2227_n_spl_0,
    g2227_n_spl_
  );


  buf

  (
    g2227_p_spl_,
    g2227_p
  );


  buf

  (
    g2227_p_spl_0,
    g2227_p_spl_
  );


  buf

  (
    g2231_n_spl_,
    g2231_n
  );


  buf

  (
    g2230_n_spl_,
    g2230_n
  );


  buf

  (
    g2231_p_spl_,
    g2231_p
  );


  buf

  (
    g2230_p_spl_,
    g2230_p
  );


  buf

  (
    g2232_n_spl_,
    g2232_n
  );


  buf

  (
    g2232_n_spl_0,
    g2232_n_spl_
  );


  buf

  (
    g2232_p_spl_,
    g2232_p
  );


  buf

  (
    g2232_p_spl_0,
    g2232_p_spl_
  );


  buf

  (
    g2233_n_spl_,
    g2233_n
  );


  buf

  (
    g2222_n_spl_,
    g2222_n
  );


  buf

  (
    g2233_p_spl_,
    g2233_p
  );


  buf

  (
    g2222_p_spl_,
    g2222_p
  );


  buf

  (
    g2234_n_spl_,
    g2234_n
  );


  buf

  (
    g2234_n_spl_0,
    g2234_n_spl_
  );


  buf

  (
    g2234_p_spl_,
    g2234_p
  );


  buf

  (
    g2234_p_spl_0,
    g2234_p_spl_
  );


  buf

  (
    g2238_n_spl_,
    g2238_n
  );


  buf

  (
    g2237_n_spl_,
    g2237_n
  );


  buf

  (
    g2238_p_spl_,
    g2238_p
  );


  buf

  (
    g2237_p_spl_,
    g2237_p
  );


  buf

  (
    g2239_n_spl_,
    g2239_n
  );


  buf

  (
    g2239_n_spl_0,
    g2239_n_spl_
  );


  buf

  (
    g2239_p_spl_,
    g2239_p
  );


  buf

  (
    g2239_p_spl_0,
    g2239_p_spl_
  );


  buf

  (
    g2257_n_spl_,
    g2257_n
  );


  buf

  (
    g2256_n_spl_,
    g2256_n
  );


  buf

  (
    g2257_p_spl_,
    g2257_p
  );


  buf

  (
    g2256_p_spl_,
    g2256_p
  );


  buf

  (
    g2258_n_spl_,
    g2258_n
  );


  buf

  (
    g2258_n_spl_0,
    g2258_n_spl_
  );


  buf

  (
    g2258_p_spl_,
    g2258_p
  );


  buf

  (
    g2258_p_spl_0,
    g2258_p_spl_
  );


  buf

  (
    g2262_n_spl_,
    g2262_n
  );


  buf

  (
    g2261_n_spl_,
    g2261_n
  );


  buf

  (
    g2262_p_spl_,
    g2262_p
  );


  buf

  (
    g2261_p_spl_,
    g2261_p
  );


  buf

  (
    g2263_n_spl_,
    g2263_n
  );


  buf

  (
    g2263_n_spl_0,
    g2263_n_spl_
  );


  buf

  (
    g2263_p_spl_,
    g2263_p
  );


  buf

  (
    g2263_p_spl_0,
    g2263_p_spl_
  );


  buf

  (
    g2264_n_spl_,
    g2264_n
  );


  buf

  (
    g2253_n_spl_,
    g2253_n
  );


  buf

  (
    g2264_p_spl_,
    g2264_p
  );


  buf

  (
    g2253_p_spl_,
    g2253_p
  );


  buf

  (
    g2265_n_spl_,
    g2265_n
  );


  buf

  (
    g2265_n_spl_0,
    g2265_n_spl_
  );


  buf

  (
    g2265_p_spl_,
    g2265_p
  );


  buf

  (
    g2265_p_spl_0,
    g2265_p_spl_
  );


  buf

  (
    g2269_n_spl_,
    g2269_n
  );


  buf

  (
    g2268_n_spl_,
    g2268_n
  );


  buf

  (
    g2269_p_spl_,
    g2269_p
  );


  buf

  (
    g2268_p_spl_,
    g2268_p
  );


  buf

  (
    g2270_n_spl_,
    g2270_n
  );


  buf

  (
    g2270_n_spl_0,
    g2270_n_spl_
  );


  buf

  (
    g2270_p_spl_,
    g2270_p
  );


  buf

  (
    g2270_p_spl_0,
    g2270_p_spl_
  );


  buf

  (
    g2271_n_spl_,
    g2271_n
  );


  buf

  (
    g2250_n_spl_,
    g2250_n
  );


  buf

  (
    g2271_p_spl_,
    g2271_p
  );


  buf

  (
    g2250_p_spl_,
    g2250_p
  );


  buf

  (
    g2272_n_spl_,
    g2272_n
  );


  buf

  (
    g2272_n_spl_0,
    g2272_n_spl_
  );


  buf

  (
    g2272_p_spl_,
    g2272_p
  );


  buf

  (
    g2272_p_spl_0,
    g2272_p_spl_
  );


  buf

  (
    g2276_n_spl_,
    g2276_n
  );


  buf

  (
    g2275_n_spl_,
    g2275_n
  );


  buf

  (
    g2276_p_spl_,
    g2276_p
  );


  buf

  (
    g2275_p_spl_,
    g2275_p
  );


  buf

  (
    g2277_n_spl_,
    g2277_n
  );


  buf

  (
    g2277_n_spl_0,
    g2277_n_spl_
  );


  buf

  (
    g2277_p_spl_,
    g2277_p
  );


  buf

  (
    g2277_p_spl_0,
    g2277_p_spl_
  );


  buf

  (
    g2278_n_spl_,
    g2278_n
  );


  buf

  (
    g2247_n_spl_,
    g2247_n
  );


  buf

  (
    g2278_p_spl_,
    g2278_p
  );


  buf

  (
    g2247_p_spl_,
    g2247_p
  );


  buf

  (
    g2279_n_spl_,
    g2279_n
  );


  buf

  (
    g2279_n_spl_0,
    g2279_n_spl_
  );


  buf

  (
    g2279_p_spl_,
    g2279_p
  );


  buf

  (
    g2279_p_spl_0,
    g2279_p_spl_
  );


  buf

  (
    g2283_n_spl_,
    g2283_n
  );


  buf

  (
    g2282_n_spl_,
    g2282_n
  );


  buf

  (
    g2283_p_spl_,
    g2283_p
  );


  buf

  (
    g2282_p_spl_,
    g2282_p
  );


  buf

  (
    g2284_n_spl_,
    g2284_n
  );


  buf

  (
    g2284_n_spl_0,
    g2284_n_spl_
  );


  buf

  (
    g2284_p_spl_,
    g2284_p
  );


  buf

  (
    g2284_p_spl_0,
    g2284_p_spl_
  );


  buf

  (
    G7_p_spl_,
    G7_p
  );


  buf

  (
    G7_p_spl_0,
    G7_p_spl_
  );


  buf

  (
    G7_p_spl_1,
    G7_p_spl_
  );


  buf

  (
    G7_n_spl_,
    G7_n
  );


  buf

  (
    G7_n_spl_0,
    G7_n_spl_
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G6_p_spl_0,
    G6_p_spl_
  );


  buf

  (
    G6_p_spl_1,
    G6_p_spl_
  );


  buf

  (
    G6_n_spl_,
    G6_n
  );


  buf

  (
    G6_n_spl_0,
    G6_n_spl_
  );


  buf

  (
    g2288_n_spl_,
    g2288_n
  );


  buf

  (
    g2287_p_spl_,
    g2287_p
  );


  buf

  (
    g2288_p_spl_,
    g2288_p
  );


  buf

  (
    g2287_n_spl_,
    g2287_n
  );


  buf

  (
    g2289_n_spl_,
    g2289_n
  );


  buf

  (
    g2289_p_spl_,
    g2289_p
  );


  buf

  (
    g2290_n_spl_,
    g2290_n
  );


  buf

  (
    g2290_n_spl_0,
    g2290_n_spl_
  );


  buf

  (
    g2290_p_spl_,
    g2290_p
  );


  buf

  (
    g2290_p_spl_0,
    g2290_p_spl_
  );


  buf

  (
    G5_p_spl_,
    G5_p
  );


  buf

  (
    G5_p_spl_0,
    G5_p_spl_
  );


  buf

  (
    G5_n_spl_,
    G5_n
  );


  buf

  (
    G5_n_spl_0,
    G5_n_spl_
  );


  buf

  (
    g2294_n_spl_,
    g2294_n
  );


  buf

  (
    g2293_p_spl_,
    g2293_p
  );


  buf

  (
    g2294_p_spl_,
    g2294_p
  );


  buf

  (
    g2293_n_spl_,
    g2293_n
  );


  buf

  (
    g2295_n_spl_,
    g2295_n
  );


  buf

  (
    g2295_p_spl_,
    g2295_p
  );


  buf

  (
    g2296_p_spl_,
    g2296_p
  );


  buf

  (
    G13_p_spl_,
    G13_p
  );


  buf

  (
    G13_p_spl_0,
    G13_p_spl_
  );


  buf

  (
    G13_p_spl_00,
    G13_p_spl_0
  );


  buf

  (
    G13_p_spl_1,
    G13_p_spl_
  );


  buf

  (
    G13_n_spl_,
    G13_n
  );


  buf

  (
    G13_n_spl_0,
    G13_n_spl_
  );


  buf

  (
    G13_n_spl_1,
    G13_n_spl_
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G12_p_spl_0,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_00,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_1,
    G12_p_spl_
  );


  buf

  (
    G12_n_spl_,
    G12_n
  );


  buf

  (
    G12_n_spl_0,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_1,
    G12_n_spl_
  );


  buf

  (
    g2299_n_spl_,
    g2299_n
  );


  buf

  (
    g2298_p_spl_,
    g2298_p
  );


  buf

  (
    g2299_p_spl_,
    g2299_p
  );


  buf

  (
    g2298_n_spl_,
    g2298_n
  );


  buf

  (
    g2300_n_spl_,
    g2300_n
  );


  buf

  (
    g2300_p_spl_,
    g2300_p
  );


  buf

  (
    g2301_n_spl_,
    g2301_n
  );


  buf

  (
    g2301_n_spl_0,
    g2301_n_spl_
  );


  buf

  (
    g2301_p_spl_,
    g2301_p
  );


  buf

  (
    g2301_p_spl_0,
    g2301_p_spl_
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    G11_p_spl_0,
    G11_p_spl_
  );


  buf

  (
    G11_p_spl_00,
    G11_p_spl_0
  );


  buf

  (
    G11_p_spl_1,
    G11_p_spl_
  );


  buf

  (
    G11_n_spl_,
    G11_n
  );


  buf

  (
    G11_n_spl_0,
    G11_n_spl_
  );


  buf

  (
    G11_n_spl_1,
    G11_n_spl_
  );


  buf

  (
    g2305_n_spl_,
    g2305_n
  );


  buf

  (
    g2304_p_spl_,
    g2304_p
  );


  buf

  (
    g2305_p_spl_,
    g2305_p
  );


  buf

  (
    g2304_n_spl_,
    g2304_n
  );


  buf

  (
    g2306_n_spl_,
    g2306_n
  );


  buf

  (
    g2306_p_spl_,
    g2306_p
  );


  buf

  (
    g2307_n_spl_,
    g2307_n
  );


  buf

  (
    g2307_n_spl_0,
    g2307_n_spl_
  );


  buf

  (
    g2303_n_spl_,
    g2303_n
  );


  buf

  (
    g2307_p_spl_,
    g2307_p
  );


  buf

  (
    g2307_p_spl_0,
    g2307_p_spl_
  );


  buf

  (
    g2303_p_spl_,
    g2303_p
  );


  buf

  (
    g2308_n_spl_,
    g2308_n
  );


  buf

  (
    g2308_n_spl_0,
    g2308_n_spl_
  );


  buf

  (
    g2308_p_spl_,
    g2308_p
  );


  buf

  (
    g2308_p_spl_0,
    g2308_p_spl_
  );


  buf

  (
    g2312_n_spl_,
    g2312_n
  );


  buf

  (
    g2311_n_spl_,
    g2311_n
  );


  buf

  (
    g2312_p_spl_,
    g2312_p
  );


  buf

  (
    g2311_p_spl_,
    g2311_p
  );


  buf

  (
    g2313_n_spl_,
    g2313_n
  );


  buf

  (
    g2313_n_spl_0,
    g2313_n_spl_
  );


  buf

  (
    g2313_p_spl_,
    g2313_p
  );


  buf

  (
    g2313_p_spl_0,
    g2313_p_spl_
  );


  buf

  (
    G10_p_spl_,
    G10_p
  );


  buf

  (
    G10_p_spl_0,
    G10_p_spl_
  );


  buf

  (
    G10_p_spl_1,
    G10_p_spl_
  );


  buf

  (
    G10_n_spl_,
    G10_n
  );


  buf

  (
    G10_n_spl_0,
    G10_n_spl_
  );


  buf

  (
    G10_n_spl_1,
    G10_n_spl_
  );


  buf

  (
    g2320_n_spl_,
    g2320_n
  );


  buf

  (
    g2319_p_spl_,
    g2319_p
  );


  buf

  (
    g2320_p_spl_,
    g2320_p
  );


  buf

  (
    g2319_n_spl_,
    g2319_n
  );


  buf

  (
    g2321_n_spl_,
    g2321_n
  );


  buf

  (
    g2321_p_spl_,
    g2321_p
  );


  buf

  (
    g2322_n_spl_,
    g2322_n
  );


  buf

  (
    g2322_n_spl_0,
    g2322_n_spl_
  );


  buf

  (
    g2318_n_spl_,
    g2318_n
  );


  buf

  (
    g2322_p_spl_,
    g2322_p
  );


  buf

  (
    g2322_p_spl_0,
    g2322_p_spl_
  );


  buf

  (
    g2318_p_spl_,
    g2318_p
  );


  buf

  (
    g2323_n_spl_,
    g2323_n
  );


  buf

  (
    g2323_n_spl_0,
    g2323_n_spl_
  );


  buf

  (
    g2323_p_spl_,
    g2323_p
  );


  buf

  (
    g2323_p_spl_0,
    g2323_p_spl_
  );


  buf

  (
    g2327_n_spl_,
    g2327_n
  );


  buf

  (
    g2326_n_spl_,
    g2326_n
  );


  buf

  (
    g2327_p_spl_,
    g2327_p
  );


  buf

  (
    g2326_p_spl_,
    g2326_p
  );


  buf

  (
    g2328_n_spl_,
    g2328_n
  );


  buf

  (
    g2328_n_spl_0,
    g2328_n_spl_
  );


  buf

  (
    g2328_p_spl_,
    g2328_p
  );


  buf

  (
    g2328_p_spl_0,
    g2328_p_spl_
  );


  buf

  (
    g2341_n_spl_,
    g2341_n
  );


  buf

  (
    g2340_n_spl_,
    g2340_n
  );


  buf

  (
    g2341_p_spl_,
    g2341_p
  );


  buf

  (
    g2340_p_spl_,
    g2340_p
  );


  buf

  (
    g2342_n_spl_,
    g2342_n
  );


  buf

  (
    g2342_n_spl_0,
    g2342_n_spl_
  );


  buf

  (
    g2342_p_spl_,
    g2342_p
  );


  buf

  (
    g2347_n_spl_,
    g2347_n
  );


  buf

  (
    g2347_n_spl_0,
    g2347_n_spl_
  );


  buf

  (
    g2216_p_spl_,
    g2216_p
  );


  buf

  (
    g2356_n_spl_,
    g2356_n
  );


  buf

  (
    g2355_n_spl_,
    g2355_n
  );


  buf

  (
    g2356_p_spl_,
    g2356_p
  );


  buf

  (
    g2355_p_spl_,
    g2355_p
  );


  buf

  (
    g2357_n_spl_,
    g2357_n
  );


  buf

  (
    g2357_n_spl_0,
    g2357_n_spl_
  );


  buf

  (
    g2357_p_spl_,
    g2357_p
  );


  buf

  (
    g2357_p_spl_0,
    g2357_p_spl_
  );


  buf

  (
    g2361_n_spl_,
    g2361_n
  );


  buf

  (
    g2360_n_spl_,
    g2360_n
  );


  buf

  (
    g2361_p_spl_,
    g2361_p
  );


  buf

  (
    g2360_p_spl_,
    g2360_p
  );


  buf

  (
    g2362_n_spl_,
    g2362_n
  );


  buf

  (
    g2362_n_spl_0,
    g2362_n_spl_
  );


  buf

  (
    g2362_p_spl_,
    g2362_p
  );


  buf

  (
    g2362_p_spl_0,
    g2362_p_spl_
  );


  buf

  (
    g2363_n_spl_,
    g2363_n
  );


  buf

  (
    g2352_n_spl_,
    g2352_n
  );


  buf

  (
    g2363_p_spl_,
    g2363_p
  );


  buf

  (
    g2352_p_spl_,
    g2352_p
  );


  buf

  (
    g2364_n_spl_,
    g2364_n
  );


  buf

  (
    g2364_n_spl_0,
    g2364_n_spl_
  );


  buf

  (
    g2364_p_spl_,
    g2364_p
  );


  buf

  (
    g2364_p_spl_0,
    g2364_p_spl_
  );


  buf

  (
    g2368_n_spl_,
    g2368_n
  );


  buf

  (
    g2367_n_spl_,
    g2367_n
  );


  buf

  (
    g2368_p_spl_,
    g2368_p
  );


  buf

  (
    g2367_p_spl_,
    g2367_p
  );


  buf

  (
    g2369_n_spl_,
    g2369_n
  );


  buf

  (
    g2369_n_spl_0,
    g2369_n_spl_
  );


  buf

  (
    g2369_p_spl_,
    g2369_p
  );


  buf

  (
    g2369_p_spl_0,
    g2369_p_spl_
  );


  buf

  (
    g2376_n_spl_,
    g2376_n
  );


  buf

  (
    g2375_n_spl_,
    g2375_n
  );


  buf

  (
    g2376_p_spl_,
    g2376_p
  );


  buf

  (
    g2375_p_spl_,
    g2375_p
  );


  buf

  (
    g2377_n_spl_,
    g2377_n
  );


  buf

  (
    g2377_n_spl_0,
    g2377_n_spl_
  );


  buf

  (
    g2377_p_spl_,
    g2377_p
  );


  buf

  (
    g2377_p_spl_0,
    g2377_p_spl_
  );


  buf

  (
    g2381_n_spl_,
    g2381_n
  );


  buf

  (
    g2380_n_spl_,
    g2380_n
  );


  buf

  (
    g2381_p_spl_,
    g2381_p
  );


  buf

  (
    g2380_p_spl_,
    g2380_p
  );


  buf

  (
    g2382_n_spl_,
    g2382_n
  );


  buf

  (
    g2382_n_spl_0,
    g2382_n_spl_
  );


  buf

  (
    g2382_p_spl_,
    g2382_p
  );


  buf

  (
    g2382_p_spl_0,
    g2382_p_spl_
  );


  buf

  (
    g2383_n_spl_,
    g2383_n
  );


  buf

  (
    g2372_n_spl_,
    g2372_n
  );


  buf

  (
    g2383_p_spl_,
    g2383_p
  );


  buf

  (
    g2372_p_spl_,
    g2372_p
  );


  buf

  (
    g2384_n_spl_,
    g2384_n
  );


  buf

  (
    g2384_n_spl_0,
    g2384_n_spl_
  );


  buf

  (
    g2384_p_spl_,
    g2384_p
  );


  buf

  (
    g2389_n_spl_,
    g2389_n
  );


  buf

  (
    g2389_n_spl_0,
    g2389_n_spl_
  );


  buf

  (
    g2163_n_spl_,
    g2163_n
  );


  buf

  (
    g2163_n_spl_0,
    g2163_n_spl_
  );


  buf

  (
    g2178_n_spl_,
    g2178_n
  );


  buf

  (
    g2178_n_spl_0,
    g2178_n_spl_
  );


  buf

  (
    g2193_n_spl_,
    g2193_n
  );


  buf

  (
    g2193_n_spl_0,
    g2193_n_spl_
  );


  buf

  (
    g2198_n_spl_,
    g2198_n
  );


  buf

  (
    g2198_n_spl_0,
    g2198_n_spl_
  );


  buf

  (
    g2201_n_spl_,
    g2201_n
  );


  buf

  (
    g2135_n_spl_,
    g2135_n
  );


  buf

  (
    g2204_n_spl_,
    g2204_n
  );


  buf

  (
    g2136_n_spl_,
    g2136_n
  );


  buf

  (
    g2207_n_spl_,
    g2207_n
  );


  buf

  (
    g2137_n_spl_,
    g2137_n
  );


  buf

  (
    g2210_n_spl_,
    g2210_n
  );


  buf

  (
    g2138_n_spl_,
    g2138_n
  );


  buf

  (
    g1846_n_spl_,
    g1846_n
  );


  buf

  (
    g1846_n_spl_0,
    g1846_n_spl_
  );


  buf

  (
    g1846_p_spl_,
    g1846_p
  );


  buf

  (
    G20_p_spl_,
    G20_p
  );


  buf

  (
    G20_p_spl_0,
    G20_p_spl_
  );


  buf

  (
    G20_p_spl_00,
    G20_p_spl_0
  );


  buf

  (
    G20_p_spl_01,
    G20_p_spl_0
  );


  buf

  (
    G20_p_spl_1,
    G20_p_spl_
  );


  buf

  (
    G20_p_spl_10,
    G20_p_spl_1
  );


  buf

  (
    G20_n_spl_,
    G20_n
  );


  buf

  (
    G20_n_spl_0,
    G20_n_spl_
  );


  buf

  (
    G20_n_spl_00,
    G20_n_spl_0
  );


  buf

  (
    G20_n_spl_01,
    G20_n_spl_0
  );


  buf

  (
    G20_n_spl_1,
    G20_n_spl_
  );


  buf

  (
    g2411_n_spl_,
    g2411_n
  );


  buf

  (
    g2410_n_spl_,
    g2410_n
  );


  buf

  (
    g2411_p_spl_,
    g2411_p
  );


  buf

  (
    g2410_p_spl_,
    g2410_p
  );


  buf

  (
    g2412_n_spl_,
    g2412_n
  );


  buf

  (
    g2412_n_spl_0,
    g2412_n_spl_
  );


  buf

  (
    g2412_p_spl_,
    g2412_p
  );


  buf

  (
    g2416_n_spl_,
    g2416_n
  );


  buf

  (
    g2415_n_spl_,
    g2415_n
  );


  buf

  (
    g2416_p_spl_,
    g2416_p
  );


  buf

  (
    g2415_p_spl_,
    g2415_p
  );


  buf

  (
    g2417_n_spl_,
    g2417_n
  );


  buf

  (
    g2417_n_spl_0,
    g2417_n_spl_
  );


  buf

  (
    g2417_p_spl_,
    g2417_p
  );


  buf

  (
    g2426_n_spl_,
    g2426_n
  );


  buf

  (
    g2425_n_spl_,
    g2425_n
  );


  buf

  (
    g2426_p_spl_,
    g2426_p
  );


  buf

  (
    g2425_p_spl_,
    g2425_p
  );


  buf

  (
    g2427_n_spl_,
    g2427_n
  );


  buf

  (
    g2427_n_spl_0,
    g2427_n_spl_
  );


  buf

  (
    g2427_p_spl_,
    g2427_p
  );


  buf

  (
    g2431_n_spl_,
    g2431_n
  );


  buf

  (
    g2430_n_spl_,
    g2430_n
  );


  buf

  (
    g2431_p_spl_,
    g2431_p
  );


  buf

  (
    g2430_p_spl_,
    g2430_p
  );


  buf

  (
    g2432_n_spl_,
    g2432_n
  );


  buf

  (
    g2432_n_spl_0,
    g2432_n_spl_
  );


  buf

  (
    g2432_p_spl_,
    g2432_p
  );


  buf

  (
    g2444_n_spl_,
    g2444_n
  );


  buf

  (
    g2443_n_spl_,
    g2443_n
  );


  buf

  (
    g2444_p_spl_,
    g2444_p
  );


  buf

  (
    g2443_p_spl_,
    g2443_p
  );


  buf

  (
    g2445_n_spl_,
    g2445_n
  );


  buf

  (
    g2445_n_spl_0,
    g2445_n_spl_
  );


  buf

  (
    g2445_p_spl_,
    g2445_p
  );


  buf

  (
    g2445_p_spl_0,
    g2445_p_spl_
  );


  buf

  (
    g2449_n_spl_,
    g2449_n
  );


  buf

  (
    g2448_n_spl_,
    g2448_n
  );


  buf

  (
    g2450_n_spl_,
    g2450_n
  );


  buf

  (
    g2450_n_spl_0,
    g2450_n_spl_
  );


  buf

  (
    g2459_n_spl_,
    g2459_n
  );


  buf

  (
    g2458_n_spl_,
    g2458_n
  );


  buf

  (
    g2459_p_spl_,
    g2459_p
  );


  buf

  (
    g2458_p_spl_,
    g2458_p
  );


  buf

  (
    g2460_n_spl_,
    g2460_n
  );


  buf

  (
    g2460_n_spl_0,
    g2460_n_spl_
  );


  buf

  (
    g2460_p_spl_,
    g2460_p
  );


  buf

  (
    g2460_p_spl_0,
    g2460_p_spl_
  );


  buf

  (
    g2464_p_spl_,
    g2464_p
  );


  buf

  (
    g2463_p_spl_,
    g2463_p
  );


  buf

  (
    g2465_p_spl_,
    g2465_p
  );


  buf

  (
    g2465_p_spl_0,
    g2465_p_spl_
  );


  buf

  (
    g1806_n_spl_,
    g1806_n
  );


  buf

  (
    g1806_n_spl_0,
    g1806_n_spl_
  );


  buf

  (
    g1811_n_spl_,
    g1811_n
  );


  buf

  (
    g1811_n_spl_0,
    g1811_n_spl_
  );


  buf

  (
    g1816_n_spl_,
    g1816_n
  );


  buf

  (
    g1816_n_spl_0,
    g1816_n_spl_
  );


  buf

  (
    g1831_n_spl_,
    g1831_n
  );


  buf

  (
    g1831_n_spl_0,
    g1831_n_spl_
  );


  buf

  (
    g2296_n_spl_,
    g2296_n
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    g2483_n_spl_,
    g2483_n
  );


  buf

  (
    g2482_p_spl_,
    g2482_p
  );


  buf

  (
    g2483_p_spl_,
    g2483_p
  );


  buf

  (
    g2482_n_spl_,
    g2482_n
  );


  buf

  (
    g2484_n_spl_,
    g2484_n
  );


  buf

  (
    g2484_p_spl_,
    g2484_p
  );


  buf

  (
    g2485_p_spl_,
    g2485_p
  );


  buf

  (
    G9_p_spl_,
    G9_p
  );


  buf

  (
    G9_p_spl_0,
    G9_p_spl_
  );


  buf

  (
    G9_p_spl_00,
    G9_p_spl_0
  );


  buf

  (
    G9_p_spl_1,
    G9_p_spl_
  );


  buf

  (
    G9_n_spl_,
    G9_n
  );


  buf

  (
    G9_n_spl_0,
    G9_n_spl_
  );


  buf

  (
    g2493_n_spl_,
    g2493_n
  );


  buf

  (
    g2492_p_spl_,
    g2492_p
  );


  buf

  (
    g2493_p_spl_,
    g2493_p
  );


  buf

  (
    g2492_n_spl_,
    g2492_n
  );


  buf

  (
    g2494_n_spl_,
    g2494_n
  );


  buf

  (
    g2494_p_spl_,
    g2494_p
  );


  buf

  (
    g2495_n_spl_,
    g2495_n
  );


  buf

  (
    g2495_n_spl_0,
    g2495_n_spl_
  );


  buf

  (
    g2491_n_spl_,
    g2491_n
  );


  buf

  (
    g2495_p_spl_,
    g2495_p
  );


  buf

  (
    g2495_p_spl_0,
    g2495_p_spl_
  );


  buf

  (
    g2491_p_spl_,
    g2491_p
  );


  buf

  (
    g2496_n_spl_,
    g2496_n
  );


  buf

  (
    g2496_n_spl_0,
    g2496_n_spl_
  );


  buf

  (
    g2496_p_spl_,
    g2496_p
  );


  buf

  (
    g2496_p_spl_0,
    g2496_p_spl_
  );


  buf

  (
    g2500_n_spl_,
    g2500_n
  );


  buf

  (
    g2499_n_spl_,
    g2499_n
  );


  buf

  (
    g2500_p_spl_,
    g2500_p
  );


  buf

  (
    g2499_p_spl_,
    g2499_p
  );


  buf

  (
    g2501_n_spl_,
    g2501_n
  );


  buf

  (
    g2501_n_spl_0,
    g2501_n_spl_
  );


  buf

  (
    g2501_p_spl_,
    g2501_p
  );


  buf

  (
    g2501_p_spl_0,
    g2501_p_spl_
  );


  buf

  (
    g1869_n_spl_,
    g1869_n
  );


  buf

  (
    g1869_n_spl_0,
    g1869_n_spl_
  );


  buf

  (
    g1996_n_spl_,
    g1996_n
  );


  buf

  (
    g1996_n_spl_0,
    g1996_n_spl_
  );


  buf

  (
    g2106_n_spl_,
    g2106_n
  );


  buf

  (
    g2106_n_spl_0,
    g2106_n_spl_
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G2_p_spl_0,
    G2_p_spl_
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    n2770_lo_p_spl_,
    n2770_lo_p
  );


  buf

  (
    g2530_n_spl_,
    g2530_n
  );


  buf

  (
    g2529_n_spl_,
    g2529_n
  );


  buf

  (
    g2530_p_spl_,
    g2530_p
  );


  buf

  (
    g2529_p_spl_,
    g2529_p
  );


  buf

  (
    g2531_n_spl_,
    g2531_n
  );


  buf

  (
    g2531_n_spl_0,
    g2531_n_spl_
  );


  buf

  (
    g2531_p_spl_,
    g2531_p
  );


  buf

  (
    g2536_n_spl_,
    g2536_n
  );


  buf

  (
    g2536_n_spl_0,
    g2536_n_spl_
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G3_p_spl_0,
    G3_p_spl_
  );


  buf

  (
    G3_n_spl_,
    G3_n
  );


  buf

  (
    g2540_p_spl_,
    g2540_p
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_1,
    G8_p_spl_
  );


  buf

  (
    G8_n_spl_,
    G8_n
  );


  buf

  (
    G8_n_spl_0,
    G8_n_spl_
  );


  buf

  (
    g2543_n_spl_,
    g2543_n
  );


  buf

  (
    g2542_p_spl_,
    g2542_p
  );


  buf

  (
    g2543_p_spl_,
    g2543_p
  );


  buf

  (
    g2542_n_spl_,
    g2542_n
  );


  buf

  (
    g2544_n_spl_,
    g2544_n
  );


  buf

  (
    g2544_p_spl_,
    g2544_p
  );


  buf

  (
    g2545_n_spl_,
    g2545_n
  );


  buf

  (
    g2545_n_spl_0,
    g2545_n_spl_
  );


  buf

  (
    g2545_p_spl_,
    g2545_p
  );


  buf

  (
    g2545_p_spl_0,
    g2545_p_spl_
  );


  buf

  (
    g2549_n_spl_,
    g2549_n
  );


  buf

  (
    g2548_p_spl_,
    g2548_p
  );


  buf

  (
    g2549_p_spl_,
    g2549_p
  );


  buf

  (
    g2548_n_spl_,
    g2548_n
  );


  buf

  (
    g2550_n_spl_,
    g2550_n
  );


  buf

  (
    g2550_p_spl_,
    g2550_p
  );


  buf

  (
    g2551_n_spl_,
    g2551_n
  );


  buf

  (
    g2551_n_spl_0,
    g2551_n_spl_
  );


  buf

  (
    g2547_n_spl_,
    g2547_n
  );


  buf

  (
    g2551_p_spl_,
    g2551_p
  );


  buf

  (
    g2551_p_spl_0,
    g2551_p_spl_
  );


  buf

  (
    g2547_p_spl_,
    g2547_p
  );


  buf

  (
    g2552_n_spl_,
    g2552_n
  );


  buf

  (
    g2552_n_spl_0,
    g2552_n_spl_
  );


  buf

  (
    g2552_p_spl_,
    g2552_p
  );


  buf

  (
    g2557_n_spl_,
    g2557_n
  );


  buf

  (
    g2557_n_spl_0,
    g2557_n_spl_
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G14_p_spl_0,
    G14_p_spl_
  );


  buf

  (
    G14_p_spl_00,
    G14_p_spl_0
  );


  buf

  (
    G14_p_spl_1,
    G14_p_spl_
  );


  buf

  (
    G14_n_spl_,
    G14_n
  );


  buf

  (
    G14_n_spl_0,
    G14_n_spl_
  );


  buf

  (
    G14_n_spl_1,
    G14_n_spl_
  );


  buf

  (
    g2560_n_spl_,
    g2560_n
  );


  buf

  (
    g2559_p_spl_,
    g2559_p
  );


  buf

  (
    g2560_p_spl_,
    g2560_p
  );


  buf

  (
    g2559_n_spl_,
    g2559_n
  );


  buf

  (
    g2561_n_spl_,
    g2561_n
  );


  buf

  (
    g2561_p_spl_,
    g2561_p
  );


  buf

  (
    g2562_n_spl_,
    g2562_n
  );


  buf

  (
    g2562_n_spl_0,
    g2562_n_spl_
  );


  buf

  (
    g2562_p_spl_,
    g2562_p
  );


  buf

  (
    g2562_p_spl_0,
    g2562_p_spl_
  );


  buf

  (
    g2566_n_spl_,
    g2566_n
  );


  buf

  (
    g2565_p_spl_,
    g2565_p
  );


  buf

  (
    g2566_p_spl_,
    g2566_p
  );


  buf

  (
    g2565_n_spl_,
    g2565_n
  );


  buf

  (
    g2567_n_spl_,
    g2567_n
  );


  buf

  (
    g2567_p_spl_,
    g2567_p
  );


  buf

  (
    g2568_n_spl_,
    g2568_n
  );


  buf

  (
    g2568_n_spl_0,
    g2568_n_spl_
  );


  buf

  (
    g2564_n_spl_,
    g2564_n
  );


  buf

  (
    g2568_p_spl_,
    g2568_p
  );


  buf

  (
    g2568_p_spl_0,
    g2568_p_spl_
  );


  buf

  (
    g2564_p_spl_,
    g2564_p
  );


  buf

  (
    g2569_n_spl_,
    g2569_n
  );


  buf

  (
    g2569_n_spl_0,
    g2569_n_spl_
  );


  buf

  (
    g2569_p_spl_,
    g2569_p
  );


  buf

  (
    g2569_p_spl_0,
    g2569_p_spl_
  );


  buf

  (
    g2573_n_spl_,
    g2573_n
  );


  buf

  (
    g2572_n_spl_,
    g2572_n
  );


  buf

  (
    g2573_p_spl_,
    g2573_p
  );


  buf

  (
    g2572_p_spl_,
    g2572_p
  );


  buf

  (
    g2574_n_spl_,
    g2574_n
  );


  buf

  (
    g2574_n_spl_0,
    g2574_n_spl_
  );


  buf

  (
    g2574_p_spl_,
    g2574_p
  );


  buf

  (
    g2574_p_spl_0,
    g2574_p_spl_
  );


  buf

  (
    g2579_n_spl_,
    g2579_n
  );


  buf

  (
    g2579_p_spl_,
    g2579_p
  );


  buf

  (
    g2580_n_spl_,
    g2580_n
  );


  buf

  (
    g2580_n_spl_0,
    g2580_n_spl_
  );


  buf

  (
    g2580_p_spl_,
    g2580_p
  );


  buf

  (
    g2580_p_spl_0,
    g2580_p_spl_
  );


  buf

  (
    g2584_n_spl_,
    g2584_n
  );


  buf

  (
    g2583_n_spl_,
    g2583_n
  );


  buf

  (
    g2584_p_spl_,
    g2584_p
  );


  buf

  (
    g2583_p_spl_,
    g2583_p
  );


  buf

  (
    g2585_n_spl_,
    g2585_n
  );


  buf

  (
    g2585_n_spl_0,
    g2585_n_spl_
  );


  buf

  (
    g2585_p_spl_,
    g2585_p
  );


  buf

  (
    g2585_p_spl_0,
    g2585_p_spl_
  );


  buf

  (
    g2586_n_spl_,
    g2586_n
  );


  buf

  (
    g2577_n_spl_,
    g2577_n
  );


  buf

  (
    g2586_p_spl_,
    g2586_p
  );


  buf

  (
    g2577_p_spl_,
    g2577_p
  );


  buf

  (
    g2587_n_spl_,
    g2587_n
  );


  buf

  (
    g2587_n_spl_0,
    g2587_n_spl_
  );


  buf

  (
    g2587_p_spl_,
    g2587_p
  );


  buf

  (
    g2592_n_spl_,
    g2592_n
  );


  buf

  (
    g2592_n_spl_0,
    g2592_n_spl_
  );


  buf

  (
    g2422_n_spl_,
    g2422_n
  );


  buf

  (
    g2422_n_spl_0,
    g2422_n_spl_
  );


  buf

  (
    g2437_n_spl_,
    g2437_n
  );


  buf

  (
    g2437_n_spl_0,
    g2437_n_spl_
  );


  buf

  (
    g2452_n_spl_,
    g2452_n
  );


  buf

  (
    g2452_n_spl_0,
    g2452_n_spl_
  );


  buf

  (
    g2467_n_spl_,
    g2467_n
  );


  buf

  (
    g2467_n_spl_0,
    g2467_n_spl_
  );


  buf

  (
    g2512_n_spl_,
    g2512_n
  );


  buf

  (
    g2332_n_spl_,
    g2332_n
  );


  buf

  (
    g2518_n_spl_,
    g2518_n
  );


  buf

  (
    g2333_n_spl_,
    g2333_n
  );


  buf

  (
    g2515_n_spl_,
    g2515_n
  );


  buf

  (
    g2334_n_spl_,
    g2334_n
  );


  buf

  (
    g2519_p_spl_,
    g2519_p
  );


  buf

  (
    g2335_n_spl_,
    g2335_n
  );


  buf

  (
    g2509_n_spl_,
    g2509_n
  );


  buf

  (
    g2349_n_spl_,
    g2349_n
  );


  buf

  (
    g2506_p_spl_,
    g2506_p
  );


  buf

  (
    g2390_p_spl_,
    g2390_p
  );


  buf

  (
    g2485_n_spl_,
    g2485_n
  );


  buf

  (
    g2613_n_spl_,
    g2613_n
  );


  buf

  (
    g2612_p_spl_,
    g2612_p
  );


  buf

  (
    g2612_n_spl_,
    g2612_n
  );


  buf

  (
    g2614_n_spl_,
    g2614_n
  );


  buf

  (
    g2615_p_spl_,
    g2615_p
  );


  buf

  (
    g2621_n_spl_,
    g2621_n
  );


  buf

  (
    g2621_p_spl_,
    g2621_p
  );


  buf

  (
    g2622_n_spl_,
    g2622_n
  );


  buf

  (
    g2622_n_spl_0,
    g2622_n_spl_
  );


  buf

  (
    g2622_p_spl_,
    g2622_p
  );


  buf

  (
    g2622_p_spl_0,
    g2622_p_spl_
  );


  buf

  (
    g2626_p_spl_,
    g2626_p
  );


  buf

  (
    g2625_p_spl_,
    g2625_p
  );


  buf

  (
    g2627_p_spl_,
    g2627_p
  );


  buf

  (
    g2627_p_spl_0,
    g2627_p_spl_
  );


  buf

  (
    g2634_n_spl_,
    g2634_n
  );


  buf

  (
    g2634_p_spl_,
    g2634_p
  );


  buf

  (
    g2635_n_spl_,
    g2635_n
  );


  buf

  (
    g2635_n_spl_0,
    g2635_n_spl_
  );


  buf

  (
    g2635_p_spl_,
    g2635_p
  );


  buf

  (
    g2635_p_spl_0,
    g2635_p_spl_
  );


  buf

  (
    g2639_n_spl_,
    g2639_n
  );


  buf

  (
    g2638_n_spl_,
    g2638_n
  );


  buf

  (
    g2639_p_spl_,
    g2639_p
  );


  buf

  (
    g2638_p_spl_,
    g2638_p
  );


  buf

  (
    g2640_n_spl_,
    g2640_n
  );


  buf

  (
    g2640_n_spl_0,
    g2640_n_spl_
  );


  buf

  (
    g2640_p_spl_,
    g2640_p
  );


  buf

  (
    g2640_p_spl_0,
    g2640_p_spl_
  );


  buf

  (
    g2641_n_spl_,
    g2641_n
  );


  buf

  (
    g2632_n_spl_,
    g2632_n
  );


  buf

  (
    g2641_p_spl_,
    g2641_p
  );


  buf

  (
    g2632_p_spl_,
    g2632_p
  );


  buf

  (
    g2642_n_spl_,
    g2642_n
  );


  buf

  (
    g2642_n_spl_0,
    g2642_n_spl_
  );


  buf

  (
    g2642_p_spl_,
    g2642_p
  );


  buf

  (
    g2646_n_spl_,
    g2646_n
  );


  buf

  (
    g2645_n_spl_,
    g2645_n
  );


  buf

  (
    g2646_p_spl_,
    g2646_p
  );


  buf

  (
    g2645_p_spl_,
    g2645_p
  );


  buf

  (
    g2647_n_spl_,
    g2647_n
  );


  buf

  (
    g2647_n_spl_0,
    g2647_n_spl_
  );


  buf

  (
    g2647_p_spl_,
    g2647_p
  );


  buf

  (
    g2654_n_spl_,
    g2654_n
  );


  buf

  (
    g2653_n_spl_,
    g2653_n
  );


  buf

  (
    g2654_p_spl_,
    g2654_p
  );


  buf

  (
    g2653_p_spl_,
    g2653_p
  );


  buf

  (
    g2655_n_spl_,
    g2655_n
  );


  buf

  (
    g2655_n_spl_0,
    g2655_n_spl_
  );


  buf

  (
    g2655_p_spl_,
    g2655_p
  );


  buf

  (
    g2655_p_spl_0,
    g2655_p_spl_
  );


  buf

  (
    g2659_p_spl_,
    g2659_p
  );


  buf

  (
    g2658_p_spl_,
    g2658_p
  );


  buf

  (
    g2660_p_spl_,
    g2660_p
  );


  buf

  (
    g2660_p_spl_0,
    g2660_p_spl_
  );


  buf

  (
    g2215_n_spl_,
    g2215_n
  );


  buf

  (
    g2215_n_spl_0,
    g2215_n_spl_
  );


  buf

  (
    g2241_n_spl_,
    g2241_n
  );


  buf

  (
    g2241_n_spl_0,
    g2241_n_spl_
  );


  buf

  (
    g2286_n_spl_,
    g2286_n
  );


  buf

  (
    g2286_n_spl_0,
    g2286_n_spl_
  );


  buf

  (
    g2297_n_spl_,
    g2297_n
  );


  buf

  (
    g2297_n_spl_0,
    g2297_n_spl_
  );


  buf

  (
    g2330_n_spl_,
    g2330_n
  );


  buf

  (
    g2330_n_spl_0,
    g2330_n_spl_
  );


  buf

  (
    g2607_p_spl_,
    g2607_p
  );


  buf

  (
    g2694_n_spl_,
    g2694_n
  );


  buf

  (
    g2694_p_spl_,
    g2694_p
  );


  buf

  (
    g2695_n_spl_,
    g2695_n
  );


  buf

  (
    g2695_n_spl_0,
    g2695_n_spl_
  );


  buf

  (
    g2695_p_spl_,
    g2695_p
  );


  buf

  (
    g2700_n_spl_,
    g2700_n
  );


  buf

  (
    g2700_n_spl_0,
    g2700_n_spl_
  );


  buf

  (
    g2705_n_spl_,
    g2705_n
  );


  buf

  (
    g2704_n_spl_,
    g2704_n
  );


  buf

  (
    g2705_p_spl_,
    g2705_p
  );


  buf

  (
    g2704_p_spl_,
    g2704_p
  );


  buf

  (
    g2706_n_spl_,
    g2706_n
  );


  buf

  (
    g2706_n_spl_0,
    g2706_n_spl_
  );


  buf

  (
    g2706_p_spl_,
    g2706_p
  );


  buf

  (
    g2711_n_spl_,
    g2711_n
  );


  buf

  (
    g2711_n_spl_0,
    g2711_n_spl_
  );


  buf

  (
    g2616_n_spl_,
    g2616_n
  );


  buf

  (
    g2616_n_spl_0,
    g2616_n_spl_
  );


  buf

  (
    g2629_n_spl_,
    g2629_n
  );


  buf

  (
    g2629_n_spl_0,
    g2629_n_spl_
  );


  buf

  (
    g2662_n_spl_,
    g2662_n
  );


  buf

  (
    g2662_n_spl_0,
    g2662_n_spl_
  );


  buf

  (
    g2688_n_spl_,
    g2688_n
  );


  buf

  (
    g2523_n_spl_,
    g2523_n
  );


  buf

  (
    g2685_n_spl_,
    g2685_n
  );


  buf

  (
    g2524_n_spl_,
    g2524_n
  );


  buf

  (
    g2679_n_spl_,
    g2679_n
  );


  buf

  (
    g2541_n_spl_,
    g2541_n
  );


  buf

  (
    g2541_n_spl_0,
    g2541_n_spl_
  );


  buf

  (
    g2682_p_spl_,
    g2682_p
  );


  buf

  (
    g2558_p_spl_,
    g2558_p
  );


  buf

  (
    g2677_p_spl_,
    g2677_p
  );


  buf

  (
    g2593_p_spl_,
    g2593_p
  );


  buf

  (
    g2409_n_spl_,
    g2409_n
  );


  buf

  (
    g2409_n_spl_0,
    g2409_n_spl_
  );


  buf

  (
    g2486_n_spl_,
    g2486_n
  );


  buf

  (
    g2486_n_spl_0,
    g2486_n_spl_
  );


  buf

  (
    g2503_n_spl_,
    g2503_n
  );


  buf

  (
    g2503_n_spl_0,
    g2503_n_spl_
  );


endmodule
