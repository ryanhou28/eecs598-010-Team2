
module mymod
(
  G1_p,
  G1_n,
  G2_p,
  G2_n,
  G3_p,
  G3_n,
  G4_p,
  G4_n,
  G5_p,
  G5_n,
  G6_p,
  G6_n,
  G7_p,
  G7_n,
  G8_p,
  G8_n,
  G9_p,
  G9_n,
  G10_p,
  G10_n,
  G11_p,
  G11_n,
  G12_p,
  G12_n,
  G13_p,
  G13_n,
  G14_p,
  G14_n,
  G15_p,
  G15_n,
  G16_p,
  G16_n,
  G17_p,
  G17_n,
  G18_p,
  G18_n,
  G19_p,
  G19_n,
  G20_p,
  G20_n,
  G21_p,
  G21_n,
  G22_p,
  G22_n,
  G23_p,
  G23_n,
  G24_p,
  G24_n,
  G25_p,
  G25_n,
  G26_p,
  G26_n,
  G27_p,
  G27_n,
  G28_p,
  G28_n,
  G29_p,
  G29_n,
  G30_p,
  G30_n,
  G31_p,
  G31_n,
  G32_p,
  G32_n,
  G33_p,
  G33_n,
  G34_p,
  G34_n,
  G35_p,
  G35_n,
  G36_p,
  G36_n,
  G37_p,
  G37_n,
  G38_p,
  G38_n,
  G39_p,
  G39_n,
  G40_p,
  G40_n,
  G41_p,
  G41_n,
  G468_n,
  G469_n,
  G470_n,
  G471_n,
  G472_n,
  G473_n,
  G474_n,
  G475_n,
  G476_n,
  G477_n,
  G478_n,
  G479_n,
  G480_n,
  G481_n,
  G482_n,
  G483_n,
  G484_n,
  G485_n,
  G486_n,
  G487_n,
  G488_n,
  G489_n,
  G490_n,
  G491_n,
  G492_n,
  G493_n,
  G494_n,
  G495_n,
  G496_n,
  G497_n,
  G498_n,
  G499_n
);

  input G1_p;input G1_n;input G2_p;input G2_n;input G3_p;input G3_n;input G4_p;input G4_n;input G5_p;input G5_n;input G6_p;input G6_n;input G7_p;input G7_n;input G8_p;input G8_n;input G9_p;input G9_n;input G10_p;input G10_n;input G11_p;input G11_n;input G12_p;input G12_n;input G13_p;input G13_n;input G14_p;input G14_n;input G15_p;input G15_n;input G16_p;input G16_n;input G17_p;input G17_n;input G18_p;input G18_n;input G19_p;input G19_n;input G20_p;input G20_n;input G21_p;input G21_n;input G22_p;input G22_n;input G23_p;input G23_n;input G24_p;input G24_n;input G25_p;input G25_n;input G26_p;input G26_n;input G27_p;input G27_n;input G28_p;input G28_n;input G29_p;input G29_n;input G30_p;input G30_n;input G31_p;input G31_n;input G32_p;input G32_n;input G33_p;input G33_n;input G34_p;input G34_n;input G35_p;input G35_n;input G36_p;input G36_n;input G37_p;input G37_n;input G38_p;input G38_n;input G39_p;input G39_n;input G40_p;input G40_n;input G41_p;input G41_n;
  output G468_n;output G469_n;output G470_n;output G471_n;output G472_n;output G473_n;output G474_n;output G475_n;output G476_n;output G477_n;output G478_n;output G479_n;output G480_n;output G481_n;output G482_n;output G483_n;output G484_n;output G485_n;output G486_n;output G487_n;output G488_n;output G489_n;output G490_n;output G491_n;output G492_n;output G493_n;output G494_n;output G495_n;output G496_n;output G497_n;output G498_n;output G499_n;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire g42_p;
  wire g42_n;
  wire g43_p;
  wire g43_n;
  wire g44_p;
  wire g44_n;
  wire g45_p;
  wire g45_n;
  wire g46_p;
  wire g46_n;
  wire g47_p;
  wire g47_n;
  wire g48_p;
  wire g48_n;
  wire g49_p;
  wire g49_n;
  wire g50_p;
  wire g50_n;
  wire g51_p;
  wire g51_n;
  wire g52_p;
  wire g52_n;
  wire g53_p;
  wire g53_n;
  wire g54_p;
  wire g54_n;
  wire g55_p;
  wire g55_n;
  wire g56_p;
  wire g56_n;
  wire g57_p;
  wire g57_n;
  wire g58_p;
  wire g58_n;
  wire g59_p;
  wire g59_n;
  wire g60_p;
  wire g60_n;
  wire g61_p;
  wire g61_n;
  wire g62_p;
  wire g62_n;
  wire g63_p;
  wire g63_n;
  wire g64_p;
  wire g64_n;
  wire g65_p;
  wire g65_n;
  wire g66_p;
  wire g66_n;
  wire g67_p;
  wire g67_n;
  wire g68_p;
  wire g68_n;
  wire g69_p;
  wire g69_n;
  wire g70_p;
  wire g70_n;
  wire g71_p;
  wire g71_n;
  wire g72_p;
  wire g72_n;
  wire g73_p;
  wire g73_n;
  wire g74_p;
  wire g74_n;
  wire g75_p;
  wire g75_n;
  wire g76_p;
  wire g76_n;
  wire g77_p;
  wire g77_n;
  wire g78_p;
  wire g78_n;
  wire g79_p;
  wire g79_n;
  wire g80_p;
  wire g80_n;
  wire g81_p;
  wire g81_n;
  wire g82_p;
  wire g82_n;
  wire g83_p;
  wire g83_n;
  wire g84_p;
  wire g84_n;
  wire g85_p;
  wire g85_n;
  wire g86_p;
  wire g86_n;
  wire g87_p;
  wire g87_n;
  wire g88_p;
  wire g88_n;
  wire g89_p;
  wire g89_n;
  wire g90_p;
  wire g90_n;
  wire g91_p;
  wire g91_n;
  wire g92_p;
  wire g92_n;
  wire g93_p;
  wire g93_n;
  wire g94_p;
  wire g94_n;
  wire g95_p;
  wire g95_n;
  wire g96_p;
  wire g96_n;
  wire g97_p;
  wire g97_n;
  wire g98_p;
  wire g98_n;
  wire g99_p;
  wire g99_n;
  wire g100_p;
  wire g100_n;
  wire g101_p;
  wire g101_n;
  wire g102_p;
  wire g102_n;
  wire g103_p;
  wire g103_n;
  wire g104_p;
  wire g104_n;
  wire g105_p;
  wire g105_n;
  wire g106_p;
  wire g106_n;
  wire g107_p;
  wire g107_n;
  wire g108_p;
  wire g108_n;
  wire g109_p;
  wire g109_n;
  wire g110_p;
  wire g110_n;
  wire g111_p;
  wire g111_n;
  wire g112_p;
  wire g112_n;
  wire g113_p;
  wire g113_n;
  wire g114_p;
  wire g114_n;
  wire g115_p;
  wire g115_n;
  wire g116_p;
  wire g116_n;
  wire g117_p;
  wire g117_n;
  wire g118_p;
  wire g118_n;
  wire g119_p;
  wire g119_n;
  wire g120_p;
  wire g120_n;
  wire g121_p;
  wire g121_n;
  wire g122_p;
  wire g122_n;
  wire g123_p;
  wire g123_n;
  wire g124_p;
  wire g124_n;
  wire g125_p;
  wire g125_n;
  wire g126_p;
  wire g126_n;
  wire g127_p;
  wire g127_n;
  wire g128_p;
  wire g128_n;
  wire g129_p;
  wire g129_n;
  wire g130_p;
  wire g130_n;
  wire g131_p;
  wire g131_n;
  wire g132_p;
  wire g132_n;
  wire g133_p;
  wire g133_n;
  wire g134_p;
  wire g134_n;
  wire g135_p;
  wire g135_n;
  wire g136_p;
  wire g136_n;
  wire g137_p;
  wire g137_n;
  wire g138_p;
  wire g138_n;
  wire g139_p;
  wire g139_n;
  wire g140_p;
  wire g140_n;
  wire g141_p;
  wire g141_n;
  wire g142_p;
  wire g142_n;
  wire g143_p;
  wire g143_n;
  wire g144_p;
  wire g144_n;
  wire g145_p;
  wire g145_n;
  wire g146_p;
  wire g146_n;
  wire g147_p;
  wire g147_n;
  wire g148_p;
  wire g148_n;
  wire g149_p;
  wire g149_n;
  wire g150_p;
  wire g150_n;
  wire g151_p;
  wire g151_n;
  wire g152_p;
  wire g152_n;
  wire g153_p;
  wire g153_n;
  wire g154_p;
  wire g154_n;
  wire g155_p;
  wire g155_n;
  wire g156_p;
  wire g156_n;
  wire g157_p;
  wire g157_n;
  wire g158_p;
  wire g158_n;
  wire g159_p;
  wire g159_n;
  wire g160_p;
  wire g160_n;
  wire g161_p;
  wire g161_n;
  wire g162_p;
  wire g162_n;
  wire g163_p;
  wire g163_n;
  wire g164_p;
  wire g164_n;
  wire g165_p;
  wire g165_n;
  wire g166_p;
  wire g166_n;
  wire g167_p;
  wire g167_n;
  wire g168_p;
  wire g168_n;
  wire g169_p;
  wire g169_n;
  wire g170_p;
  wire g170_n;
  wire g171_p;
  wire g171_n;
  wire g172_p;
  wire g172_n;
  wire g173_p;
  wire g173_n;
  wire g174_p;
  wire g174_n;
  wire g175_p;
  wire g175_n;
  wire g176_p;
  wire g176_n;
  wire g177_p;
  wire g177_n;
  wire g178_p;
  wire g178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire G1_n_spl_;
  wire G1_n_spl_0;
  wire G1_n_spl_00;
  wire G1_n_spl_1;
  wire G5_n_spl_;
  wire G5_n_spl_0;
  wire G5_n_spl_00;
  wire G5_n_spl_1;
  wire G1_p_spl_;
  wire G1_p_spl_0;
  wire G1_p_spl_00;
  wire G1_p_spl_1;
  wire G5_p_spl_;
  wire G5_p_spl_0;
  wire G5_p_spl_00;
  wire G5_p_spl_1;
  wire G9_n_spl_;
  wire G9_n_spl_0;
  wire G9_n_spl_00;
  wire G9_n_spl_1;
  wire G13_n_spl_;
  wire G13_n_spl_0;
  wire G13_n_spl_00;
  wire G13_n_spl_1;
  wire G9_p_spl_;
  wire G9_p_spl_0;
  wire G9_p_spl_00;
  wire G9_p_spl_1;
  wire G13_p_spl_;
  wire G13_p_spl_0;
  wire G13_p_spl_00;
  wire G13_p_spl_1;
  wire g44_n_spl_;
  wire g47_p_spl_;
  wire g44_p_spl_;
  wire g47_n_spl_;
  wire G41_p_spl_;
  wire G41_p_spl_0;
  wire G41_p_spl_00;
  wire G41_p_spl_01;
  wire G41_p_spl_1;
  wire G41_p_spl_10;
  wire G41_p_spl_11;
  wire G41_n_spl_;
  wire G41_n_spl_0;
  wire G41_n_spl_00;
  wire G41_n_spl_01;
  wire G41_n_spl_1;
  wire G41_n_spl_10;
  wire G41_n_spl_11;
  wire G17_n_spl_;
  wire G17_n_spl_0;
  wire G17_n_spl_00;
  wire G17_n_spl_1;
  wire G18_n_spl_;
  wire G18_n_spl_0;
  wire G18_n_spl_00;
  wire G18_n_spl_1;
  wire G17_p_spl_;
  wire G17_p_spl_0;
  wire G17_p_spl_00;
  wire G17_p_spl_1;
  wire G18_p_spl_;
  wire G18_p_spl_0;
  wire G18_p_spl_00;
  wire G18_p_spl_1;
  wire G19_n_spl_;
  wire G19_n_spl_0;
  wire G19_n_spl_00;
  wire G19_n_spl_1;
  wire G20_n_spl_;
  wire G20_n_spl_0;
  wire G20_n_spl_00;
  wire G20_n_spl_1;
  wire G19_p_spl_;
  wire G19_p_spl_0;
  wire G19_p_spl_00;
  wire G19_p_spl_1;
  wire G20_p_spl_;
  wire G20_p_spl_0;
  wire G20_p_spl_00;
  wire G20_p_spl_1;
  wire g54_n_spl_;
  wire g57_p_spl_;
  wire g54_p_spl_;
  wire g57_n_spl_;
  wire G21_n_spl_;
  wire G21_n_spl_0;
  wire G21_n_spl_00;
  wire G21_n_spl_1;
  wire G22_n_spl_;
  wire G22_n_spl_0;
  wire G22_n_spl_00;
  wire G22_n_spl_1;
  wire G21_p_spl_;
  wire G21_p_spl_0;
  wire G21_p_spl_00;
  wire G21_p_spl_1;
  wire G22_p_spl_;
  wire G22_p_spl_0;
  wire G22_p_spl_00;
  wire G22_p_spl_1;
  wire G23_n_spl_;
  wire G23_n_spl_0;
  wire G23_n_spl_00;
  wire G23_n_spl_1;
  wire G24_n_spl_;
  wire G24_n_spl_0;
  wire G24_n_spl_00;
  wire G24_n_spl_1;
  wire G23_p_spl_;
  wire G23_p_spl_0;
  wire G23_p_spl_00;
  wire G23_p_spl_1;
  wire G24_p_spl_;
  wire G24_p_spl_0;
  wire G24_p_spl_00;
  wire G24_p_spl_1;
  wire g63_n_spl_;
  wire g66_p_spl_;
  wire g63_p_spl_;
  wire g66_n_spl_;
  wire g60_n_spl_;
  wire g60_n_spl_0;
  wire g60_n_spl_1;
  wire g69_n_spl_;
  wire g69_n_spl_0;
  wire g69_n_spl_1;
  wire g60_p_spl_;
  wire g60_p_spl_0;
  wire g60_p_spl_1;
  wire g69_p_spl_;
  wire g69_p_spl_0;
  wire g69_p_spl_1;
  wire g51_n_spl_;
  wire g72_p_spl_;
  wire g51_p_spl_;
  wire g72_n_spl_;
  wire g50_p_spl_;
  wire g75_n_spl_;
  wire g50_n_spl_;
  wire g75_p_spl_;
  wire G25_n_spl_;
  wire G25_n_spl_0;
  wire G25_n_spl_00;
  wire G25_n_spl_1;
  wire G29_n_spl_;
  wire G29_n_spl_0;
  wire G29_n_spl_00;
  wire G29_n_spl_1;
  wire G25_p_spl_;
  wire G25_p_spl_0;
  wire G25_p_spl_00;
  wire G25_p_spl_1;
  wire G29_p_spl_;
  wire G29_p_spl_0;
  wire G29_p_spl_00;
  wire G29_p_spl_1;
  wire g81_n_spl_;
  wire g84_p_spl_;
  wire g81_p_spl_;
  wire g84_n_spl_;
  wire G6_n_spl_;
  wire G6_n_spl_0;
  wire G6_n_spl_00;
  wire G6_n_spl_1;
  wire G6_p_spl_;
  wire G6_p_spl_0;
  wire G6_p_spl_00;
  wire G6_p_spl_1;
  wire G7_n_spl_;
  wire G7_n_spl_0;
  wire G7_n_spl_00;
  wire G7_n_spl_1;
  wire G8_n_spl_;
  wire G8_n_spl_0;
  wire G8_n_spl_00;
  wire G8_n_spl_1;
  wire G7_p_spl_;
  wire G7_p_spl_0;
  wire G7_p_spl_00;
  wire G7_p_spl_1;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire G8_p_spl_00;
  wire G8_p_spl_1;
  wire g91_n_spl_;
  wire g94_p_spl_;
  wire g91_p_spl_;
  wire g94_n_spl_;
  wire G2_n_spl_;
  wire G2_n_spl_0;
  wire G2_n_spl_00;
  wire G2_n_spl_1;
  wire G2_p_spl_;
  wire G2_p_spl_0;
  wire G2_p_spl_00;
  wire G2_p_spl_1;
  wire G3_n_spl_;
  wire G3_n_spl_0;
  wire G3_n_spl_00;
  wire G3_n_spl_1;
  wire G4_n_spl_;
  wire G4_n_spl_0;
  wire G4_n_spl_00;
  wire G4_n_spl_1;
  wire G3_p_spl_;
  wire G3_p_spl_0;
  wire G3_p_spl_00;
  wire G3_p_spl_1;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_00;
  wire G4_p_spl_1;
  wire g100_n_spl_;
  wire g103_p_spl_;
  wire g100_p_spl_;
  wire g103_n_spl_;
  wire g97_n_spl_;
  wire g97_n_spl_0;
  wire g97_n_spl_1;
  wire g106_n_spl_;
  wire g106_n_spl_0;
  wire g106_n_spl_1;
  wire g97_p_spl_;
  wire g97_p_spl_0;
  wire g97_p_spl_1;
  wire g106_p_spl_;
  wire g106_p_spl_0;
  wire g106_p_spl_1;
  wire g88_n_spl_;
  wire g109_p_spl_;
  wire g88_p_spl_;
  wire g109_n_spl_;
  wire g87_p_spl_;
  wire g112_n_spl_;
  wire g87_n_spl_;
  wire g112_p_spl_;
  wire G26_n_spl_;
  wire G26_n_spl_0;
  wire G26_n_spl_00;
  wire G26_n_spl_1;
  wire G30_n_spl_;
  wire G30_n_spl_0;
  wire G30_n_spl_00;
  wire G30_n_spl_1;
  wire G26_p_spl_;
  wire G26_p_spl_0;
  wire G26_p_spl_00;
  wire G26_p_spl_1;
  wire G30_p_spl_;
  wire G30_p_spl_0;
  wire G30_p_spl_00;
  wire G30_p_spl_1;
  wire g118_n_spl_;
  wire g121_p_spl_;
  wire g118_p_spl_;
  wire g121_n_spl_;
  wire G14_n_spl_;
  wire G14_n_spl_0;
  wire G14_n_spl_00;
  wire G14_n_spl_1;
  wire G14_p_spl_;
  wire G14_p_spl_0;
  wire G14_p_spl_00;
  wire G14_p_spl_1;
  wire G15_n_spl_;
  wire G15_n_spl_0;
  wire G15_n_spl_00;
  wire G15_n_spl_1;
  wire G16_n_spl_;
  wire G16_n_spl_0;
  wire G16_n_spl_00;
  wire G16_n_spl_1;
  wire G15_p_spl_;
  wire G15_p_spl_0;
  wire G15_p_spl_00;
  wire G15_p_spl_1;
  wire G16_p_spl_;
  wire G16_p_spl_0;
  wire G16_p_spl_00;
  wire G16_p_spl_1;
  wire g128_n_spl_;
  wire g131_p_spl_;
  wire g128_p_spl_;
  wire g131_n_spl_;
  wire G10_n_spl_;
  wire G10_n_spl_0;
  wire G10_n_spl_00;
  wire G10_n_spl_1;
  wire G10_p_spl_;
  wire G10_p_spl_0;
  wire G10_p_spl_00;
  wire G10_p_spl_1;
  wire G11_n_spl_;
  wire G11_n_spl_0;
  wire G11_n_spl_00;
  wire G11_n_spl_1;
  wire G12_n_spl_;
  wire G12_n_spl_0;
  wire G12_n_spl_00;
  wire G12_n_spl_1;
  wire G11_p_spl_;
  wire G11_p_spl_0;
  wire G11_p_spl_00;
  wire G11_p_spl_1;
  wire G12_p_spl_;
  wire G12_p_spl_0;
  wire G12_p_spl_00;
  wire G12_p_spl_1;
  wire g137_n_spl_;
  wire g140_p_spl_;
  wire g137_p_spl_;
  wire g140_n_spl_;
  wire g134_n_spl_;
  wire g134_n_spl_0;
  wire g134_n_spl_1;
  wire g143_n_spl_;
  wire g143_n_spl_0;
  wire g143_n_spl_1;
  wire g134_p_spl_;
  wire g134_p_spl_0;
  wire g134_p_spl_1;
  wire g143_p_spl_;
  wire g143_p_spl_0;
  wire g143_p_spl_1;
  wire g125_n_spl_;
  wire g146_p_spl_;
  wire g125_p_spl_;
  wire g146_n_spl_;
  wire g124_p_spl_;
  wire g149_n_spl_;
  wire g124_n_spl_;
  wire g149_p_spl_;
  wire g115_n_spl_;
  wire g115_n_spl_0;
  wire g115_n_spl_00;
  wire g115_n_spl_01;
  wire g115_n_spl_1;
  wire g115_n_spl_10;
  wire g152_p_spl_;
  wire g152_p_spl_0;
  wire g152_p_spl_00;
  wire g152_p_spl_01;
  wire g152_p_spl_1;
  wire g152_p_spl_10;
  wire g115_p_spl_;
  wire g115_p_spl_0;
  wire g115_p_spl_00;
  wire g115_p_spl_01;
  wire g115_p_spl_1;
  wire g115_p_spl_10;
  wire g152_n_spl_;
  wire g152_n_spl_0;
  wire g152_n_spl_00;
  wire g152_n_spl_01;
  wire g152_n_spl_1;
  wire g152_n_spl_10;
  wire G28_n_spl_;
  wire G28_n_spl_0;
  wire G28_n_spl_00;
  wire G28_n_spl_1;
  wire G32_n_spl_;
  wire G32_n_spl_0;
  wire G32_n_spl_00;
  wire G32_n_spl_1;
  wire G28_p_spl_;
  wire G28_p_spl_0;
  wire G28_p_spl_00;
  wire G28_p_spl_1;
  wire G32_p_spl_;
  wire G32_p_spl_0;
  wire G32_p_spl_00;
  wire G32_p_spl_1;
  wire g156_n_spl_;
  wire g159_p_spl_;
  wire g156_p_spl_;
  wire g159_n_spl_;
  wire g163_n_spl_;
  wire g166_p_spl_;
  wire g163_p_spl_;
  wire g166_n_spl_;
  wire g162_p_spl_;
  wire g169_n_spl_;
  wire g162_n_spl_;
  wire g169_p_spl_;
  wire G27_n_spl_;
  wire G27_n_spl_0;
  wire G27_n_spl_00;
  wire G27_n_spl_1;
  wire G31_n_spl_;
  wire G31_n_spl_0;
  wire G31_n_spl_00;
  wire G31_n_spl_1;
  wire G27_p_spl_;
  wire G27_p_spl_0;
  wire G27_p_spl_00;
  wire G27_p_spl_1;
  wire G31_p_spl_;
  wire G31_p_spl_0;
  wire G31_p_spl_00;
  wire G31_p_spl_1;
  wire g175_n_spl_;
  wire g178_p_spl_;
  wire g175_p_spl_;
  wire g178_n_spl_;
  wire g182_n_spl_;
  wire g185_p_spl_;
  wire g182_p_spl_;
  wire g185_n_spl_;
  wire g181_p_spl_;
  wire g188_n_spl_;
  wire g181_n_spl_;
  wire g188_p_spl_;
  wire g172_p_spl_;
  wire g172_p_spl_0;
  wire g172_p_spl_00;
  wire g172_p_spl_01;
  wire g172_p_spl_1;
  wire g172_p_spl_10;
  wire g172_p_spl_11;
  wire g191_n_spl_;
  wire g191_n_spl_0;
  wire g191_n_spl_00;
  wire g191_n_spl_01;
  wire g191_n_spl_1;
  wire g191_n_spl_10;
  wire g191_n_spl_11;
  wire g172_n_spl_;
  wire g172_n_spl_0;
  wire g172_n_spl_00;
  wire g172_n_spl_01;
  wire g172_n_spl_1;
  wire g172_n_spl_10;
  wire g172_n_spl_11;
  wire g191_p_spl_;
  wire g191_p_spl_0;
  wire g191_p_spl_00;
  wire g191_p_spl_01;
  wire g191_p_spl_1;
  wire g191_p_spl_10;
  wire g191_p_spl_11;
  wire g195_n_spl_;
  wire g198_p_spl_;
  wire g195_p_spl_;
  wire g198_n_spl_;
  wire g205_n_spl_;
  wire g208_p_spl_;
  wire g205_p_spl_;
  wire g208_n_spl_;
  wire g211_n_spl_;
  wire g211_n_spl_0;
  wire g211_n_spl_1;
  wire g211_p_spl_;
  wire g211_p_spl_0;
  wire g211_p_spl_1;
  wire g202_n_spl_;
  wire g214_p_spl_;
  wire g202_p_spl_;
  wire g214_n_spl_;
  wire g201_p_spl_;
  wire g217_n_spl_;
  wire g201_n_spl_;
  wire g217_p_spl_;
  wire g223_n_spl_;
  wire g226_p_spl_;
  wire g223_p_spl_;
  wire g226_n_spl_;
  wire g233_n_spl_;
  wire g236_p_spl_;
  wire g233_p_spl_;
  wire g236_n_spl_;
  wire g239_n_spl_;
  wire g239_n_spl_0;
  wire g239_n_spl_1;
  wire g239_p_spl_;
  wire g239_p_spl_0;
  wire g239_p_spl_1;
  wire g230_n_spl_;
  wire g242_p_spl_;
  wire g230_p_spl_;
  wire g242_n_spl_;
  wire g229_p_spl_;
  wire g245_n_spl_;
  wire g229_n_spl_;
  wire g245_p_spl_;
  wire g251_n_spl_;
  wire g254_p_spl_;
  wire g251_p_spl_;
  wire g254_n_spl_;
  wire g258_n_spl_;
  wire g261_p_spl_;
  wire g258_p_spl_;
  wire g261_n_spl_;
  wire g257_p_spl_;
  wire g264_n_spl_;
  wire g257_n_spl_;
  wire g264_p_spl_;
  wire g78_n_spl_;
  wire g78_n_spl_0;
  wire g78_n_spl_00;
  wire g78_n_spl_01;
  wire g78_n_spl_1;
  wire g78_n_spl_10;
  wire g267_p_spl_;
  wire g267_p_spl_0;
  wire g267_p_spl_00;
  wire g267_p_spl_01;
  wire g267_p_spl_1;
  wire g267_p_spl_10;
  wire g78_p_spl_;
  wire g78_p_spl_0;
  wire g78_p_spl_00;
  wire g78_p_spl_01;
  wire g78_p_spl_1;
  wire g78_p_spl_10;
  wire g267_n_spl_;
  wire g267_n_spl_0;
  wire g267_n_spl_00;
  wire g267_n_spl_01;
  wire g267_n_spl_1;
  wire g267_n_spl_10;
  wire g248_p_spl_;
  wire g248_p_spl_0;
  wire g248_p_spl_00;
  wire g248_p_spl_01;
  wire g248_p_spl_1;
  wire g248_p_spl_10;
  wire g248_p_spl_11;
  wire g268_p_spl_;
  wire g248_n_spl_;
  wire g248_n_spl_0;
  wire g248_n_spl_00;
  wire g248_n_spl_01;
  wire g248_n_spl_1;
  wire g248_n_spl_10;
  wire g248_n_spl_11;
  wire g268_n_spl_;
  wire g270_p_spl_;
  wire g270_n_spl_;
  wire g269_n_spl_;
  wire g271_n_spl_;
  wire g269_p_spl_;
  wire g271_p_spl_;
  wire g220_p_spl_;
  wire g220_p_spl_0;
  wire g220_p_spl_00;
  wire g220_p_spl_01;
  wire g220_p_spl_1;
  wire g220_p_spl_10;
  wire g220_p_spl_11;
  wire g220_n_spl_;
  wire g220_n_spl_0;
  wire g220_n_spl_00;
  wire g220_n_spl_01;
  wire g220_n_spl_1;
  wire g220_n_spl_10;
  wire g220_n_spl_11;
  wire g274_n_spl_;
  wire g274_n_spl_0;
  wire g274_p_spl_;
  wire g274_p_spl_0;
  wire g192_p_spl_;
  wire g279_n_spl_;
  wire g192_n_spl_;
  wire g279_p_spl_;
  wire g153_p_spl_;
  wire g280_p_spl_;
  wire g153_n_spl_;
  wire g280_n_spl_;
  wire g281_p_spl_;
  wire g281_p_spl_0;
  wire g281_p_spl_1;
  wire g281_n_spl_;
  wire g281_n_spl_0;
  wire g281_n_spl_1;
  wire g298_p_spl_;
  wire g299_p_spl_;
  wire g298_n_spl_;
  wire g299_n_spl_;
  wire g300_p_spl_;
  wire g300_p_spl_0;
  wire g300_p_spl_1;
  wire g300_n_spl_;
  wire g300_n_spl_0;
  wire g300_n_spl_1;
  wire g317_p_spl_;
  wire g317_n_spl_;
  wire g318_p_spl_;
  wire g318_p_spl_0;
  wire g318_p_spl_1;
  wire g318_n_spl_;
  wire g318_n_spl_0;
  wire g318_n_spl_1;
  wire g335_p_spl_;
  wire g335_n_spl_;
  wire g336_p_spl_;
  wire g336_p_spl_0;
  wire g336_p_spl_1;
  wire g336_n_spl_;
  wire g336_n_spl_0;
  wire g336_n_spl_1;
  wire g359_n_spl_;
  wire g359_n_spl_0;
  wire g359_p_spl_;
  wire g359_p_spl_0;
  wire g361_p_spl_;
  wire g361_p_spl_0;
  wire g361_p_spl_1;
  wire g361_n_spl_;
  wire g361_n_spl_0;
  wire g361_n_spl_1;
  wire g378_p_spl_;
  wire g378_n_spl_;
  wire g379_p_spl_;
  wire g379_p_spl_0;
  wire g379_p_spl_1;
  wire g379_n_spl_;
  wire g379_n_spl_0;
  wire g379_n_spl_1;
  wire g397_p_spl_;
  wire g397_p_spl_0;
  wire g397_p_spl_1;
  wire g397_n_spl_;
  wire g397_n_spl_0;
  wire g397_n_spl_1;
  wire g414_p_spl_;
  wire g414_p_spl_0;
  wire g414_p_spl_1;
  wire g414_n_spl_;
  wire g414_n_spl_0;
  wire g414_n_spl_1;

  LA
  g_g42_p
  (
    .dout(g42_p),
    .din1(G1_n_spl_00),
    .din2(G5_n_spl_00)
  );


  FA
  g_g42_n
  (
    .dout(g42_n),
    .din1(G1_p_spl_00),
    .din2(G5_p_spl_00)
  );


  LA
  g_g43_p
  (
    .dout(g43_p),
    .din1(G1_p_spl_00),
    .din2(G5_p_spl_00)
  );


  FA
  g_g43_n
  (
    .dout(g43_n),
    .din1(G1_n_spl_00),
    .din2(G5_n_spl_00)
  );


  LA
  g_g44_p
  (
    .dout(g44_p),
    .din1(g42_n),
    .din2(g43_n)
  );


  FA
  g_g44_n
  (
    .dout(g44_n),
    .din1(g42_p),
    .din2(g43_p)
  );


  LA
  g_g45_p
  (
    .dout(g45_p),
    .din1(G9_n_spl_00),
    .din2(G13_n_spl_00)
  );


  FA
  g_g45_n
  (
    .dout(g45_n),
    .din1(G9_p_spl_00),
    .din2(G13_p_spl_00)
  );


  LA
  g_g46_p
  (
    .dout(g46_p),
    .din1(G9_p_spl_00),
    .din2(G13_p_spl_00)
  );


  FA
  g_g46_n
  (
    .dout(g46_n),
    .din1(G9_n_spl_00),
    .din2(G13_n_spl_00)
  );


  LA
  g_g47_p
  (
    .dout(g47_p),
    .din1(g45_n),
    .din2(g46_n)
  );


  FA
  g_g47_n
  (
    .dout(g47_n),
    .din1(g45_p),
    .din2(g46_p)
  );


  LA
  g_g48_p
  (
    .dout(g48_p),
    .din1(g44_n_spl_),
    .din2(g47_p_spl_)
  );


  FA
  g_g48_n
  (
    .dout(g48_n),
    .din1(g44_p_spl_),
    .din2(g47_n_spl_)
  );


  LA
  g_g49_p
  (
    .dout(g49_p),
    .din1(g44_p_spl_),
    .din2(g47_n_spl_)
  );


  FA
  g_g49_n
  (
    .dout(g49_n),
    .din1(g44_n_spl_),
    .din2(g47_p_spl_)
  );


  LA
  g_g50_p
  (
    .dout(g50_p),
    .din1(g48_n),
    .din2(g49_n)
  );


  FA
  g_g50_n
  (
    .dout(g50_n),
    .din1(g48_p),
    .din2(g49_p)
  );


  LA
  g_g51_p
  (
    .dout(g51_p),
    .din1(G33_p),
    .din2(G41_p_spl_00)
  );


  FA
  g_g51_n
  (
    .dout(g51_n),
    .din1(G33_n),
    .din2(G41_n_spl_00)
  );


  LA
  g_g52_p
  (
    .dout(g52_p),
    .din1(G17_n_spl_00),
    .din2(G18_n_spl_00)
  );


  FA
  g_g52_n
  (
    .dout(g52_n),
    .din1(G17_p_spl_00),
    .din2(G18_p_spl_00)
  );


  LA
  g_g53_p
  (
    .dout(g53_p),
    .din1(G17_p_spl_00),
    .din2(G18_p_spl_00)
  );


  FA
  g_g53_n
  (
    .dout(g53_n),
    .din1(G17_n_spl_00),
    .din2(G18_n_spl_00)
  );


  LA
  g_g54_p
  (
    .dout(g54_p),
    .din1(g52_n),
    .din2(g53_n)
  );


  FA
  g_g54_n
  (
    .dout(g54_n),
    .din1(g52_p),
    .din2(g53_p)
  );


  LA
  g_g55_p
  (
    .dout(g55_p),
    .din1(G19_n_spl_00),
    .din2(G20_n_spl_00)
  );


  FA
  g_g55_n
  (
    .dout(g55_n),
    .din1(G19_p_spl_00),
    .din2(G20_p_spl_00)
  );


  LA
  g_g56_p
  (
    .dout(g56_p),
    .din1(G19_p_spl_00),
    .din2(G20_p_spl_00)
  );


  FA
  g_g56_n
  (
    .dout(g56_n),
    .din1(G19_n_spl_00),
    .din2(G20_n_spl_00)
  );


  LA
  g_g57_p
  (
    .dout(g57_p),
    .din1(g55_n),
    .din2(g56_n)
  );


  FA
  g_g57_n
  (
    .dout(g57_n),
    .din1(g55_p),
    .din2(g56_p)
  );


  LA
  g_g58_p
  (
    .dout(g58_p),
    .din1(g54_n_spl_),
    .din2(g57_p_spl_)
  );


  FA
  g_g58_n
  (
    .dout(g58_n),
    .din1(g54_p_spl_),
    .din2(g57_n_spl_)
  );


  LA
  g_g59_p
  (
    .dout(g59_p),
    .din1(g54_p_spl_),
    .din2(g57_n_spl_)
  );


  FA
  g_g59_n
  (
    .dout(g59_n),
    .din1(g54_n_spl_),
    .din2(g57_p_spl_)
  );


  LA
  g_g60_p
  (
    .dout(g60_p),
    .din1(g58_n),
    .din2(g59_n)
  );


  FA
  g_g60_n
  (
    .dout(g60_n),
    .din1(g58_p),
    .din2(g59_p)
  );


  LA
  g_g61_p
  (
    .dout(g61_p),
    .din1(G21_n_spl_00),
    .din2(G22_n_spl_00)
  );


  FA
  g_g61_n
  (
    .dout(g61_n),
    .din1(G21_p_spl_00),
    .din2(G22_p_spl_00)
  );


  LA
  g_g62_p
  (
    .dout(g62_p),
    .din1(G21_p_spl_00),
    .din2(G22_p_spl_00)
  );


  FA
  g_g62_n
  (
    .dout(g62_n),
    .din1(G21_n_spl_00),
    .din2(G22_n_spl_00)
  );


  LA
  g_g63_p
  (
    .dout(g63_p),
    .din1(g61_n),
    .din2(g62_n)
  );


  FA
  g_g63_n
  (
    .dout(g63_n),
    .din1(g61_p),
    .din2(g62_p)
  );


  LA
  g_g64_p
  (
    .dout(g64_p),
    .din1(G23_n_spl_00),
    .din2(G24_n_spl_00)
  );


  FA
  g_g64_n
  (
    .dout(g64_n),
    .din1(G23_p_spl_00),
    .din2(G24_p_spl_00)
  );


  LA
  g_g65_p
  (
    .dout(g65_p),
    .din1(G23_p_spl_00),
    .din2(G24_p_spl_00)
  );


  FA
  g_g65_n
  (
    .dout(g65_n),
    .din1(G23_n_spl_00),
    .din2(G24_n_spl_00)
  );


  LA
  g_g66_p
  (
    .dout(g66_p),
    .din1(g64_n),
    .din2(g65_n)
  );


  FA
  g_g66_n
  (
    .dout(g66_n),
    .din1(g64_p),
    .din2(g65_p)
  );


  LA
  g_g67_p
  (
    .dout(g67_p),
    .din1(g63_n_spl_),
    .din2(g66_p_spl_)
  );


  FA
  g_g67_n
  (
    .dout(g67_n),
    .din1(g63_p_spl_),
    .din2(g66_n_spl_)
  );


  LA
  g_g68_p
  (
    .dout(g68_p),
    .din1(g63_p_spl_),
    .din2(g66_n_spl_)
  );


  FA
  g_g68_n
  (
    .dout(g68_n),
    .din1(g63_n_spl_),
    .din2(g66_p_spl_)
  );


  LA
  g_g69_p
  (
    .dout(g69_p),
    .din1(g67_n),
    .din2(g68_n)
  );


  FA
  g_g69_n
  (
    .dout(g69_n),
    .din1(g67_p),
    .din2(g68_p)
  );


  LA
  g_g70_p
  (
    .dout(g70_p),
    .din1(g60_n_spl_0),
    .din2(g69_n_spl_0)
  );


  FA
  g_g70_n
  (
    .dout(g70_n),
    .din1(g60_p_spl_0),
    .din2(g69_p_spl_0)
  );


  LA
  g_g71_p
  (
    .dout(g71_p),
    .din1(g60_p_spl_0),
    .din2(g69_p_spl_0)
  );


  FA
  g_g71_n
  (
    .dout(g71_n),
    .din1(g60_n_spl_0),
    .din2(g69_n_spl_0)
  );


  LA
  g_g72_p
  (
    .dout(g72_p),
    .din1(g70_n),
    .din2(g71_n)
  );


  FA
  g_g72_n
  (
    .dout(g72_n),
    .din1(g70_p),
    .din2(g71_p)
  );


  LA
  g_g73_p
  (
    .dout(g73_p),
    .din1(g51_n_spl_),
    .din2(g72_p_spl_)
  );


  FA
  g_g73_n
  (
    .dout(g73_n),
    .din1(g51_p_spl_),
    .din2(g72_n_spl_)
  );


  LA
  g_g74_p
  (
    .dout(g74_p),
    .din1(g51_p_spl_),
    .din2(g72_n_spl_)
  );


  FA
  g_g74_n
  (
    .dout(g74_n),
    .din1(g51_n_spl_),
    .din2(g72_p_spl_)
  );


  LA
  g_g75_p
  (
    .dout(g75_p),
    .din1(g73_n),
    .din2(g74_n)
  );


  FA
  g_g75_n
  (
    .dout(g75_n),
    .din1(g73_p),
    .din2(g74_p)
  );


  LA
  g_g76_p
  (
    .dout(g76_p),
    .din1(g50_p_spl_),
    .din2(g75_n_spl_)
  );


  FA
  g_g76_n
  (
    .dout(g76_n),
    .din1(g50_n_spl_),
    .din2(g75_p_spl_)
  );


  LA
  g_g77_p
  (
    .dout(g77_p),
    .din1(g50_n_spl_),
    .din2(g75_p_spl_)
  );


  FA
  g_g77_n
  (
    .dout(g77_n),
    .din1(g50_p_spl_),
    .din2(g75_n_spl_)
  );


  LA
  g_g78_p
  (
    .dout(g78_p),
    .din1(g76_n),
    .din2(g77_n)
  );


  FA
  g_g78_n
  (
    .dout(g78_n),
    .din1(g76_p),
    .din2(g77_p)
  );


  LA
  g_g79_p
  (
    .dout(g79_p),
    .din1(G17_n_spl_0),
    .din2(G21_n_spl_0)
  );


  FA
  g_g79_n
  (
    .dout(g79_n),
    .din1(G17_p_spl_0),
    .din2(G21_p_spl_0)
  );


  LA
  g_g80_p
  (
    .dout(g80_p),
    .din1(G17_p_spl_1),
    .din2(G21_p_spl_1)
  );


  FA
  g_g80_n
  (
    .dout(g80_n),
    .din1(G17_n_spl_1),
    .din2(G21_n_spl_1)
  );


  LA
  g_g81_p
  (
    .dout(g81_p),
    .din1(g79_n),
    .din2(g80_n)
  );


  FA
  g_g81_n
  (
    .dout(g81_n),
    .din1(g79_p),
    .din2(g80_p)
  );


  LA
  g_g82_p
  (
    .dout(g82_p),
    .din1(G25_n_spl_00),
    .din2(G29_n_spl_00)
  );


  FA
  g_g82_n
  (
    .dout(g82_n),
    .din1(G25_p_spl_00),
    .din2(G29_p_spl_00)
  );


  LA
  g_g83_p
  (
    .dout(g83_p),
    .din1(G25_p_spl_00),
    .din2(G29_p_spl_00)
  );


  FA
  g_g83_n
  (
    .dout(g83_n),
    .din1(G25_n_spl_00),
    .din2(G29_n_spl_00)
  );


  LA
  g_g84_p
  (
    .dout(g84_p),
    .din1(g82_n),
    .din2(g83_n)
  );


  FA
  g_g84_n
  (
    .dout(g84_n),
    .din1(g82_p),
    .din2(g83_p)
  );


  LA
  g_g85_p
  (
    .dout(g85_p),
    .din1(g81_n_spl_),
    .din2(g84_p_spl_)
  );


  FA
  g_g85_n
  (
    .dout(g85_n),
    .din1(g81_p_spl_),
    .din2(g84_n_spl_)
  );


  LA
  g_g86_p
  (
    .dout(g86_p),
    .din1(g81_p_spl_),
    .din2(g84_n_spl_)
  );


  FA
  g_g86_n
  (
    .dout(g86_n),
    .din1(g81_n_spl_),
    .din2(g84_p_spl_)
  );


  LA
  g_g87_p
  (
    .dout(g87_p),
    .din1(g85_n),
    .din2(g86_n)
  );


  FA
  g_g87_n
  (
    .dout(g87_n),
    .din1(g85_p),
    .din2(g86_p)
  );


  LA
  g_g88_p
  (
    .dout(g88_p),
    .din1(G37_p),
    .din2(G41_p_spl_00)
  );


  FA
  g_g88_n
  (
    .dout(g88_n),
    .din1(G37_n),
    .din2(G41_n_spl_00)
  );


  LA
  g_g89_p
  (
    .dout(g89_p),
    .din1(G5_n_spl_0),
    .din2(G6_n_spl_00)
  );


  FA
  g_g89_n
  (
    .dout(g89_n),
    .din1(G5_p_spl_0),
    .din2(G6_p_spl_00)
  );


  LA
  g_g90_p
  (
    .dout(g90_p),
    .din1(G5_p_spl_1),
    .din2(G6_p_spl_00)
  );


  FA
  g_g90_n
  (
    .dout(g90_n),
    .din1(G5_n_spl_1),
    .din2(G6_n_spl_00)
  );


  LA
  g_g91_p
  (
    .dout(g91_p),
    .din1(g89_n),
    .din2(g90_n)
  );


  FA
  g_g91_n
  (
    .dout(g91_n),
    .din1(g89_p),
    .din2(g90_p)
  );


  LA
  g_g92_p
  (
    .dout(g92_p),
    .din1(G7_n_spl_00),
    .din2(G8_n_spl_00)
  );


  FA
  g_g92_n
  (
    .dout(g92_n),
    .din1(G7_p_spl_00),
    .din2(G8_p_spl_00)
  );


  LA
  g_g93_p
  (
    .dout(g93_p),
    .din1(G7_p_spl_00),
    .din2(G8_p_spl_00)
  );


  FA
  g_g93_n
  (
    .dout(g93_n),
    .din1(G7_n_spl_00),
    .din2(G8_n_spl_00)
  );


  LA
  g_g94_p
  (
    .dout(g94_p),
    .din1(g92_n),
    .din2(g93_n)
  );


  FA
  g_g94_n
  (
    .dout(g94_n),
    .din1(g92_p),
    .din2(g93_p)
  );


  LA
  g_g95_p
  (
    .dout(g95_p),
    .din1(g91_n_spl_),
    .din2(g94_p_spl_)
  );


  FA
  g_g95_n
  (
    .dout(g95_n),
    .din1(g91_p_spl_),
    .din2(g94_n_spl_)
  );


  LA
  g_g96_p
  (
    .dout(g96_p),
    .din1(g91_p_spl_),
    .din2(g94_n_spl_)
  );


  FA
  g_g96_n
  (
    .dout(g96_n),
    .din1(g91_n_spl_),
    .din2(g94_p_spl_)
  );


  LA
  g_g97_p
  (
    .dout(g97_p),
    .din1(g95_n),
    .din2(g96_n)
  );


  FA
  g_g97_n
  (
    .dout(g97_n),
    .din1(g95_p),
    .din2(g96_p)
  );


  LA
  g_g98_p
  (
    .dout(g98_p),
    .din1(G1_n_spl_0),
    .din2(G2_n_spl_00)
  );


  FA
  g_g98_n
  (
    .dout(g98_n),
    .din1(G1_p_spl_0),
    .din2(G2_p_spl_00)
  );


  LA
  g_g99_p
  (
    .dout(g99_p),
    .din1(G1_p_spl_1),
    .din2(G2_p_spl_00)
  );


  FA
  g_g99_n
  (
    .dout(g99_n),
    .din1(G1_n_spl_1),
    .din2(G2_n_spl_00)
  );


  LA
  g_g100_p
  (
    .dout(g100_p),
    .din1(g98_n),
    .din2(g99_n)
  );


  FA
  g_g100_n
  (
    .dout(g100_n),
    .din1(g98_p),
    .din2(g99_p)
  );


  LA
  g_g101_p
  (
    .dout(g101_p),
    .din1(G3_n_spl_00),
    .din2(G4_n_spl_00)
  );


  FA
  g_g101_n
  (
    .dout(g101_n),
    .din1(G3_p_spl_00),
    .din2(G4_p_spl_00)
  );


  LA
  g_g102_p
  (
    .dout(g102_p),
    .din1(G3_p_spl_00),
    .din2(G4_p_spl_00)
  );


  FA
  g_g102_n
  (
    .dout(g102_n),
    .din1(G3_n_spl_00),
    .din2(G4_n_spl_00)
  );


  LA
  g_g103_p
  (
    .dout(g103_p),
    .din1(g101_n),
    .din2(g102_n)
  );


  FA
  g_g103_n
  (
    .dout(g103_n),
    .din1(g101_p),
    .din2(g102_p)
  );


  LA
  g_g104_p
  (
    .dout(g104_p),
    .din1(g100_n_spl_),
    .din2(g103_p_spl_)
  );


  FA
  g_g104_n
  (
    .dout(g104_n),
    .din1(g100_p_spl_),
    .din2(g103_n_spl_)
  );


  LA
  g_g105_p
  (
    .dout(g105_p),
    .din1(g100_p_spl_),
    .din2(g103_n_spl_)
  );


  FA
  g_g105_n
  (
    .dout(g105_n),
    .din1(g100_n_spl_),
    .din2(g103_p_spl_)
  );


  LA
  g_g106_p
  (
    .dout(g106_p),
    .din1(g104_n),
    .din2(g105_n)
  );


  FA
  g_g106_n
  (
    .dout(g106_n),
    .din1(g104_p),
    .din2(g105_p)
  );


  LA
  g_g107_p
  (
    .dout(g107_p),
    .din1(g97_n_spl_0),
    .din2(g106_n_spl_0)
  );


  FA
  g_g107_n
  (
    .dout(g107_n),
    .din1(g97_p_spl_0),
    .din2(g106_p_spl_0)
  );


  LA
  g_g108_p
  (
    .dout(g108_p),
    .din1(g97_p_spl_0),
    .din2(g106_p_spl_0)
  );


  FA
  g_g108_n
  (
    .dout(g108_n),
    .din1(g97_n_spl_0),
    .din2(g106_n_spl_0)
  );


  LA
  g_g109_p
  (
    .dout(g109_p),
    .din1(g107_n),
    .din2(g108_n)
  );


  FA
  g_g109_n
  (
    .dout(g109_n),
    .din1(g107_p),
    .din2(g108_p)
  );


  LA
  g_g110_p
  (
    .dout(g110_p),
    .din1(g88_n_spl_),
    .din2(g109_p_spl_)
  );


  FA
  g_g110_n
  (
    .dout(g110_n),
    .din1(g88_p_spl_),
    .din2(g109_n_spl_)
  );


  LA
  g_g111_p
  (
    .dout(g111_p),
    .din1(g88_p_spl_),
    .din2(g109_n_spl_)
  );


  FA
  g_g111_n
  (
    .dout(g111_n),
    .din1(g88_n_spl_),
    .din2(g109_p_spl_)
  );


  LA
  g_g112_p
  (
    .dout(g112_p),
    .din1(g110_n),
    .din2(g111_n)
  );


  FA
  g_g112_n
  (
    .dout(g112_n),
    .din1(g110_p),
    .din2(g111_p)
  );


  LA
  g_g113_p
  (
    .dout(g113_p),
    .din1(g87_p_spl_),
    .din2(g112_n_spl_)
  );


  FA
  g_g113_n
  (
    .dout(g113_n),
    .din1(g87_n_spl_),
    .din2(g112_p_spl_)
  );


  LA
  g_g114_p
  (
    .dout(g114_p),
    .din1(g87_n_spl_),
    .din2(g112_p_spl_)
  );


  FA
  g_g114_n
  (
    .dout(g114_n),
    .din1(g87_p_spl_),
    .din2(g112_n_spl_)
  );


  LA
  g_g115_p
  (
    .dout(g115_p),
    .din1(g113_n),
    .din2(g114_n)
  );


  FA
  g_g115_n
  (
    .dout(g115_n),
    .din1(g113_p),
    .din2(g114_p)
  );


  LA
  g_g116_p
  (
    .dout(g116_p),
    .din1(G18_n_spl_0),
    .din2(G22_n_spl_0)
  );


  FA
  g_g116_n
  (
    .dout(g116_n),
    .din1(G18_p_spl_0),
    .din2(G22_p_spl_0)
  );


  LA
  g_g117_p
  (
    .dout(g117_p),
    .din1(G18_p_spl_1),
    .din2(G22_p_spl_1)
  );


  FA
  g_g117_n
  (
    .dout(g117_n),
    .din1(G18_n_spl_1),
    .din2(G22_n_spl_1)
  );


  LA
  g_g118_p
  (
    .dout(g118_p),
    .din1(g116_n),
    .din2(g117_n)
  );


  FA
  g_g118_n
  (
    .dout(g118_n),
    .din1(g116_p),
    .din2(g117_p)
  );


  LA
  g_g119_p
  (
    .dout(g119_p),
    .din1(G26_n_spl_00),
    .din2(G30_n_spl_00)
  );


  FA
  g_g119_n
  (
    .dout(g119_n),
    .din1(G26_p_spl_00),
    .din2(G30_p_spl_00)
  );


  LA
  g_g120_p
  (
    .dout(g120_p),
    .din1(G26_p_spl_00),
    .din2(G30_p_spl_00)
  );


  FA
  g_g120_n
  (
    .dout(g120_n),
    .din1(G26_n_spl_00),
    .din2(G30_n_spl_00)
  );


  LA
  g_g121_p
  (
    .dout(g121_p),
    .din1(g119_n),
    .din2(g120_n)
  );


  FA
  g_g121_n
  (
    .dout(g121_n),
    .din1(g119_p),
    .din2(g120_p)
  );


  LA
  g_g122_p
  (
    .dout(g122_p),
    .din1(g118_n_spl_),
    .din2(g121_p_spl_)
  );


  FA
  g_g122_n
  (
    .dout(g122_n),
    .din1(g118_p_spl_),
    .din2(g121_n_spl_)
  );


  LA
  g_g123_p
  (
    .dout(g123_p),
    .din1(g118_p_spl_),
    .din2(g121_n_spl_)
  );


  FA
  g_g123_n
  (
    .dout(g123_n),
    .din1(g118_n_spl_),
    .din2(g121_p_spl_)
  );


  LA
  g_g124_p
  (
    .dout(g124_p),
    .din1(g122_n),
    .din2(g123_n)
  );


  FA
  g_g124_n
  (
    .dout(g124_n),
    .din1(g122_p),
    .din2(g123_p)
  );


  LA
  g_g125_p
  (
    .dout(g125_p),
    .din1(G38_p),
    .din2(G41_p_spl_01)
  );


  FA
  g_g125_n
  (
    .dout(g125_n),
    .din1(G38_n),
    .din2(G41_n_spl_01)
  );


  LA
  g_g126_p
  (
    .dout(g126_p),
    .din1(G13_n_spl_0),
    .din2(G14_n_spl_00)
  );


  FA
  g_g126_n
  (
    .dout(g126_n),
    .din1(G13_p_spl_0),
    .din2(G14_p_spl_00)
  );


  LA
  g_g127_p
  (
    .dout(g127_p),
    .din1(G13_p_spl_1),
    .din2(G14_p_spl_00)
  );


  FA
  g_g127_n
  (
    .dout(g127_n),
    .din1(G13_n_spl_1),
    .din2(G14_n_spl_00)
  );


  LA
  g_g128_p
  (
    .dout(g128_p),
    .din1(g126_n),
    .din2(g127_n)
  );


  FA
  g_g128_n
  (
    .dout(g128_n),
    .din1(g126_p),
    .din2(g127_p)
  );


  LA
  g_g129_p
  (
    .dout(g129_p),
    .din1(G15_n_spl_00),
    .din2(G16_n_spl_00)
  );


  FA
  g_g129_n
  (
    .dout(g129_n),
    .din1(G15_p_spl_00),
    .din2(G16_p_spl_00)
  );


  LA
  g_g130_p
  (
    .dout(g130_p),
    .din1(G15_p_spl_00),
    .din2(G16_p_spl_00)
  );


  FA
  g_g130_n
  (
    .dout(g130_n),
    .din1(G15_n_spl_00),
    .din2(G16_n_spl_00)
  );


  LA
  g_g131_p
  (
    .dout(g131_p),
    .din1(g129_n),
    .din2(g130_n)
  );


  FA
  g_g131_n
  (
    .dout(g131_n),
    .din1(g129_p),
    .din2(g130_p)
  );


  LA
  g_g132_p
  (
    .dout(g132_p),
    .din1(g128_n_spl_),
    .din2(g131_p_spl_)
  );


  FA
  g_g132_n
  (
    .dout(g132_n),
    .din1(g128_p_spl_),
    .din2(g131_n_spl_)
  );


  LA
  g_g133_p
  (
    .dout(g133_p),
    .din1(g128_p_spl_),
    .din2(g131_n_spl_)
  );


  FA
  g_g133_n
  (
    .dout(g133_n),
    .din1(g128_n_spl_),
    .din2(g131_p_spl_)
  );


  LA
  g_g134_p
  (
    .dout(g134_p),
    .din1(g132_n),
    .din2(g133_n)
  );


  FA
  g_g134_n
  (
    .dout(g134_n),
    .din1(g132_p),
    .din2(g133_p)
  );


  LA
  g_g135_p
  (
    .dout(g135_p),
    .din1(G9_n_spl_0),
    .din2(G10_n_spl_00)
  );


  FA
  g_g135_n
  (
    .dout(g135_n),
    .din1(G9_p_spl_0),
    .din2(G10_p_spl_00)
  );


  LA
  g_g136_p
  (
    .dout(g136_p),
    .din1(G9_p_spl_1),
    .din2(G10_p_spl_00)
  );


  FA
  g_g136_n
  (
    .dout(g136_n),
    .din1(G9_n_spl_1),
    .din2(G10_n_spl_00)
  );


  LA
  g_g137_p
  (
    .dout(g137_p),
    .din1(g135_n),
    .din2(g136_n)
  );


  FA
  g_g137_n
  (
    .dout(g137_n),
    .din1(g135_p),
    .din2(g136_p)
  );


  LA
  g_g138_p
  (
    .dout(g138_p),
    .din1(G11_n_spl_00),
    .din2(G12_n_spl_00)
  );


  FA
  g_g138_n
  (
    .dout(g138_n),
    .din1(G11_p_spl_00),
    .din2(G12_p_spl_00)
  );


  LA
  g_g139_p
  (
    .dout(g139_p),
    .din1(G11_p_spl_00),
    .din2(G12_p_spl_00)
  );


  FA
  g_g139_n
  (
    .dout(g139_n),
    .din1(G11_n_spl_00),
    .din2(G12_n_spl_00)
  );


  LA
  g_g140_p
  (
    .dout(g140_p),
    .din1(g138_n),
    .din2(g139_n)
  );


  FA
  g_g140_n
  (
    .dout(g140_n),
    .din1(g138_p),
    .din2(g139_p)
  );


  LA
  g_g141_p
  (
    .dout(g141_p),
    .din1(g137_n_spl_),
    .din2(g140_p_spl_)
  );


  FA
  g_g141_n
  (
    .dout(g141_n),
    .din1(g137_p_spl_),
    .din2(g140_n_spl_)
  );


  LA
  g_g142_p
  (
    .dout(g142_p),
    .din1(g137_p_spl_),
    .din2(g140_n_spl_)
  );


  FA
  g_g142_n
  (
    .dout(g142_n),
    .din1(g137_n_spl_),
    .din2(g140_p_spl_)
  );


  LA
  g_g143_p
  (
    .dout(g143_p),
    .din1(g141_n),
    .din2(g142_n)
  );


  FA
  g_g143_n
  (
    .dout(g143_n),
    .din1(g141_p),
    .din2(g142_p)
  );


  LA
  g_g144_p
  (
    .dout(g144_p),
    .din1(g134_n_spl_0),
    .din2(g143_n_spl_0)
  );


  FA
  g_g144_n
  (
    .dout(g144_n),
    .din1(g134_p_spl_0),
    .din2(g143_p_spl_0)
  );


  LA
  g_g145_p
  (
    .dout(g145_p),
    .din1(g134_p_spl_0),
    .din2(g143_p_spl_0)
  );


  FA
  g_g145_n
  (
    .dout(g145_n),
    .din1(g134_n_spl_0),
    .din2(g143_n_spl_0)
  );


  LA
  g_g146_p
  (
    .dout(g146_p),
    .din1(g144_n),
    .din2(g145_n)
  );


  FA
  g_g146_n
  (
    .dout(g146_n),
    .din1(g144_p),
    .din2(g145_p)
  );


  LA
  g_g147_p
  (
    .dout(g147_p),
    .din1(g125_n_spl_),
    .din2(g146_p_spl_)
  );


  FA
  g_g147_n
  (
    .dout(g147_n),
    .din1(g125_p_spl_),
    .din2(g146_n_spl_)
  );


  LA
  g_g148_p
  (
    .dout(g148_p),
    .din1(g125_p_spl_),
    .din2(g146_n_spl_)
  );


  FA
  g_g148_n
  (
    .dout(g148_n),
    .din1(g125_n_spl_),
    .din2(g146_p_spl_)
  );


  LA
  g_g149_p
  (
    .dout(g149_p),
    .din1(g147_n),
    .din2(g148_n)
  );


  FA
  g_g149_n
  (
    .dout(g149_n),
    .din1(g147_p),
    .din2(g148_p)
  );


  LA
  g_g150_p
  (
    .dout(g150_p),
    .din1(g124_p_spl_),
    .din2(g149_n_spl_)
  );


  FA
  g_g150_n
  (
    .dout(g150_n),
    .din1(g124_n_spl_),
    .din2(g149_p_spl_)
  );


  LA
  g_g151_p
  (
    .dout(g151_p),
    .din1(g124_n_spl_),
    .din2(g149_p_spl_)
  );


  FA
  g_g151_n
  (
    .dout(g151_n),
    .din1(g124_p_spl_),
    .din2(g149_n_spl_)
  );


  LA
  g_g152_p
  (
    .dout(g152_p),
    .din1(g150_n),
    .din2(g151_n)
  );


  FA
  g_g152_n
  (
    .dout(g152_n),
    .din1(g150_p),
    .din2(g151_p)
  );


  LA
  g_g153_p
  (
    .dout(g153_p),
    .din1(g115_n_spl_00),
    .din2(g152_p_spl_00)
  );


  FA
  g_g153_n
  (
    .dout(g153_n),
    .din1(g115_p_spl_00),
    .din2(g152_n_spl_00)
  );


  LA
  g_g154_p
  (
    .dout(g154_p),
    .din1(G20_n_spl_0),
    .din2(G24_n_spl_0)
  );


  FA
  g_g154_n
  (
    .dout(g154_n),
    .din1(G20_p_spl_0),
    .din2(G24_p_spl_0)
  );


  LA
  g_g155_p
  (
    .dout(g155_p),
    .din1(G20_p_spl_1),
    .din2(G24_p_spl_1)
  );


  FA
  g_g155_n
  (
    .dout(g155_n),
    .din1(G20_n_spl_1),
    .din2(G24_n_spl_1)
  );


  LA
  g_g156_p
  (
    .dout(g156_p),
    .din1(g154_n),
    .din2(g155_n)
  );


  FA
  g_g156_n
  (
    .dout(g156_n),
    .din1(g154_p),
    .din2(g155_p)
  );


  LA
  g_g157_p
  (
    .dout(g157_p),
    .din1(G28_n_spl_00),
    .din2(G32_n_spl_00)
  );


  FA
  g_g157_n
  (
    .dout(g157_n),
    .din1(G28_p_spl_00),
    .din2(G32_p_spl_00)
  );


  LA
  g_g158_p
  (
    .dout(g158_p),
    .din1(G28_p_spl_00),
    .din2(G32_p_spl_00)
  );


  FA
  g_g158_n
  (
    .dout(g158_n),
    .din1(G28_n_spl_00),
    .din2(G32_n_spl_00)
  );


  LA
  g_g159_p
  (
    .dout(g159_p),
    .din1(g157_n),
    .din2(g158_n)
  );


  FA
  g_g159_n
  (
    .dout(g159_n),
    .din1(g157_p),
    .din2(g158_p)
  );


  LA
  g_g160_p
  (
    .dout(g160_p),
    .din1(g156_n_spl_),
    .din2(g159_p_spl_)
  );


  FA
  g_g160_n
  (
    .dout(g160_n),
    .din1(g156_p_spl_),
    .din2(g159_n_spl_)
  );


  LA
  g_g161_p
  (
    .dout(g161_p),
    .din1(g156_p_spl_),
    .din2(g159_n_spl_)
  );


  FA
  g_g161_n
  (
    .dout(g161_n),
    .din1(g156_n_spl_),
    .din2(g159_p_spl_)
  );


  LA
  g_g162_p
  (
    .dout(g162_p),
    .din1(g160_n),
    .din2(g161_n)
  );


  FA
  g_g162_n
  (
    .dout(g162_n),
    .din1(g160_p),
    .din2(g161_p)
  );


  LA
  g_g163_p
  (
    .dout(g163_p),
    .din1(G40_p),
    .din2(G41_p_spl_01)
  );


  FA
  g_g163_n
  (
    .dout(g163_n),
    .din1(G40_n),
    .din2(G41_n_spl_01)
  );


  LA
  g_g164_p
  (
    .dout(g164_p),
    .din1(g97_n_spl_1),
    .din2(g134_n_spl_1)
  );


  FA
  g_g164_n
  (
    .dout(g164_n),
    .din1(g97_p_spl_1),
    .din2(g134_p_spl_1)
  );


  LA
  g_g165_p
  (
    .dout(g165_p),
    .din1(g97_p_spl_1),
    .din2(g134_p_spl_1)
  );


  FA
  g_g165_n
  (
    .dout(g165_n),
    .din1(g97_n_spl_1),
    .din2(g134_n_spl_1)
  );


  LA
  g_g166_p
  (
    .dout(g166_p),
    .din1(g164_n),
    .din2(g165_n)
  );


  FA
  g_g166_n
  (
    .dout(g166_n),
    .din1(g164_p),
    .din2(g165_p)
  );


  LA
  g_g167_p
  (
    .dout(g167_p),
    .din1(g163_n_spl_),
    .din2(g166_p_spl_)
  );


  FA
  g_g167_n
  (
    .dout(g167_n),
    .din1(g163_p_spl_),
    .din2(g166_n_spl_)
  );


  LA
  g_g168_p
  (
    .dout(g168_p),
    .din1(g163_p_spl_),
    .din2(g166_n_spl_)
  );


  FA
  g_g168_n
  (
    .dout(g168_n),
    .din1(g163_n_spl_),
    .din2(g166_p_spl_)
  );


  LA
  g_g169_p
  (
    .dout(g169_p),
    .din1(g167_n),
    .din2(g168_n)
  );


  FA
  g_g169_n
  (
    .dout(g169_n),
    .din1(g167_p),
    .din2(g168_p)
  );


  LA
  g_g170_p
  (
    .dout(g170_p),
    .din1(g162_p_spl_),
    .din2(g169_n_spl_)
  );


  FA
  g_g170_n
  (
    .dout(g170_n),
    .din1(g162_n_spl_),
    .din2(g169_p_spl_)
  );


  LA
  g_g171_p
  (
    .dout(g171_p),
    .din1(g162_n_spl_),
    .din2(g169_p_spl_)
  );


  FA
  g_g171_n
  (
    .dout(g171_n),
    .din1(g162_p_spl_),
    .din2(g169_n_spl_)
  );


  LA
  g_g172_p
  (
    .dout(g172_p),
    .din1(g170_n),
    .din2(g171_n)
  );


  FA
  g_g172_n
  (
    .dout(g172_n),
    .din1(g170_p),
    .din2(g171_p)
  );


  LA
  g_g173_p
  (
    .dout(g173_p),
    .din1(G19_n_spl_0),
    .din2(G23_n_spl_0)
  );


  FA
  g_g173_n
  (
    .dout(g173_n),
    .din1(G19_p_spl_0),
    .din2(G23_p_spl_0)
  );


  LA
  g_g174_p
  (
    .dout(g174_p),
    .din1(G19_p_spl_1),
    .din2(G23_p_spl_1)
  );


  FA
  g_g174_n
  (
    .dout(g174_n),
    .din1(G19_n_spl_1),
    .din2(G23_n_spl_1)
  );


  LA
  g_g175_p
  (
    .dout(g175_p),
    .din1(g173_n),
    .din2(g174_n)
  );


  FA
  g_g175_n
  (
    .dout(g175_n),
    .din1(g173_p),
    .din2(g174_p)
  );


  LA
  g_g176_p
  (
    .dout(g176_p),
    .din1(G27_n_spl_00),
    .din2(G31_n_spl_00)
  );


  FA
  g_g176_n
  (
    .dout(g176_n),
    .din1(G27_p_spl_00),
    .din2(G31_p_spl_00)
  );


  LA
  g_g177_p
  (
    .dout(g177_p),
    .din1(G27_p_spl_00),
    .din2(G31_p_spl_00)
  );


  FA
  g_g177_n
  (
    .dout(g177_n),
    .din1(G27_n_spl_00),
    .din2(G31_n_spl_00)
  );


  LA
  g_g178_p
  (
    .dout(g178_p),
    .din1(g176_n),
    .din2(g177_n)
  );


  FA
  g_g178_n
  (
    .dout(g178_n),
    .din1(g176_p),
    .din2(g177_p)
  );


  LA
  g_g179_p
  (
    .dout(g179_p),
    .din1(g175_n_spl_),
    .din2(g178_p_spl_)
  );


  FA
  g_g179_n
  (
    .dout(g179_n),
    .din1(g175_p_spl_),
    .din2(g178_n_spl_)
  );


  LA
  g_g180_p
  (
    .dout(g180_p),
    .din1(g175_p_spl_),
    .din2(g178_n_spl_)
  );


  FA
  g_g180_n
  (
    .dout(g180_n),
    .din1(g175_n_spl_),
    .din2(g178_p_spl_)
  );


  LA
  g_g181_p
  (
    .dout(g181_p),
    .din1(g179_n),
    .din2(g180_n)
  );


  FA
  g_g181_n
  (
    .dout(g181_n),
    .din1(g179_p),
    .din2(g180_p)
  );


  LA
  g_g182_p
  (
    .dout(g182_p),
    .din1(G39_p),
    .din2(G41_p_spl_10)
  );


  FA
  g_g182_n
  (
    .dout(g182_n),
    .din1(G39_n),
    .din2(G41_n_spl_10)
  );


  LA
  g_g183_p
  (
    .dout(g183_p),
    .din1(g106_n_spl_1),
    .din2(g143_n_spl_1)
  );


  FA
  g_g183_n
  (
    .dout(g183_n),
    .din1(g106_p_spl_1),
    .din2(g143_p_spl_1)
  );


  LA
  g_g184_p
  (
    .dout(g184_p),
    .din1(g106_p_spl_1),
    .din2(g143_p_spl_1)
  );


  FA
  g_g184_n
  (
    .dout(g184_n),
    .din1(g106_n_spl_1),
    .din2(g143_n_spl_1)
  );


  LA
  g_g185_p
  (
    .dout(g185_p),
    .din1(g183_n),
    .din2(g184_n)
  );


  FA
  g_g185_n
  (
    .dout(g185_n),
    .din1(g183_p),
    .din2(g184_p)
  );


  LA
  g_g186_p
  (
    .dout(g186_p),
    .din1(g182_n_spl_),
    .din2(g185_p_spl_)
  );


  FA
  g_g186_n
  (
    .dout(g186_n),
    .din1(g182_p_spl_),
    .din2(g185_n_spl_)
  );


  LA
  g_g187_p
  (
    .dout(g187_p),
    .din1(g182_p_spl_),
    .din2(g185_n_spl_)
  );


  FA
  g_g187_n
  (
    .dout(g187_n),
    .din1(g182_n_spl_),
    .din2(g185_p_spl_)
  );


  LA
  g_g188_p
  (
    .dout(g188_p),
    .din1(g186_n),
    .din2(g187_n)
  );


  FA
  g_g188_n
  (
    .dout(g188_n),
    .din1(g186_p),
    .din2(g187_p)
  );


  LA
  g_g189_p
  (
    .dout(g189_p),
    .din1(g181_p_spl_),
    .din2(g188_n_spl_)
  );


  FA
  g_g189_n
  (
    .dout(g189_n),
    .din1(g181_n_spl_),
    .din2(g188_p_spl_)
  );


  LA
  g_g190_p
  (
    .dout(g190_p),
    .din1(g181_n_spl_),
    .din2(g188_p_spl_)
  );


  FA
  g_g190_n
  (
    .dout(g190_n),
    .din1(g181_p_spl_),
    .din2(g188_n_spl_)
  );


  LA
  g_g191_p
  (
    .dout(g191_p),
    .din1(g189_n),
    .din2(g190_n)
  );


  FA
  g_g191_n
  (
    .dout(g191_n),
    .din1(g189_p),
    .din2(g190_p)
  );


  LA
  g_g192_p
  (
    .dout(g192_p),
    .din1(g172_p_spl_00),
    .din2(g191_n_spl_00)
  );


  FA
  g_g192_n
  (
    .dout(g192_n),
    .din1(g172_n_spl_00),
    .din2(g191_p_spl_00)
  );


  LA
  g_g193_p
  (
    .dout(g193_p),
    .din1(G4_n_spl_0),
    .din2(G8_n_spl_0)
  );


  FA
  g_g193_n
  (
    .dout(g193_n),
    .din1(G4_p_spl_0),
    .din2(G8_p_spl_0)
  );


  LA
  g_g194_p
  (
    .dout(g194_p),
    .din1(G4_p_spl_1),
    .din2(G8_p_spl_1)
  );


  FA
  g_g194_n
  (
    .dout(g194_n),
    .din1(G4_n_spl_1),
    .din2(G8_n_spl_1)
  );


  LA
  g_g195_p
  (
    .dout(g195_p),
    .din1(g193_n),
    .din2(g194_n)
  );


  FA
  g_g195_n
  (
    .dout(g195_n),
    .din1(g193_p),
    .din2(g194_p)
  );


  LA
  g_g196_p
  (
    .dout(g196_p),
    .din1(G12_n_spl_0),
    .din2(G16_n_spl_0)
  );


  FA
  g_g196_n
  (
    .dout(g196_n),
    .din1(G12_p_spl_0),
    .din2(G16_p_spl_0)
  );


  LA
  g_g197_p
  (
    .dout(g197_p),
    .din1(G12_p_spl_1),
    .din2(G16_p_spl_1)
  );


  FA
  g_g197_n
  (
    .dout(g197_n),
    .din1(G12_n_spl_1),
    .din2(G16_n_spl_1)
  );


  LA
  g_g198_p
  (
    .dout(g198_p),
    .din1(g196_n),
    .din2(g197_n)
  );


  FA
  g_g198_n
  (
    .dout(g198_n),
    .din1(g196_p),
    .din2(g197_p)
  );


  LA
  g_g199_p
  (
    .dout(g199_p),
    .din1(g195_n_spl_),
    .din2(g198_p_spl_)
  );


  FA
  g_g199_n
  (
    .dout(g199_n),
    .din1(g195_p_spl_),
    .din2(g198_n_spl_)
  );


  LA
  g_g200_p
  (
    .dout(g200_p),
    .din1(g195_p_spl_),
    .din2(g198_n_spl_)
  );


  FA
  g_g200_n
  (
    .dout(g200_n),
    .din1(g195_n_spl_),
    .din2(g198_p_spl_)
  );


  LA
  g_g201_p
  (
    .dout(g201_p),
    .din1(g199_n),
    .din2(g200_n)
  );


  FA
  g_g201_n
  (
    .dout(g201_n),
    .din1(g199_p),
    .din2(g200_p)
  );


  LA
  g_g202_p
  (
    .dout(g202_p),
    .din1(G36_p),
    .din2(G41_p_spl_10)
  );


  FA
  g_g202_n
  (
    .dout(g202_n),
    .din1(G36_n),
    .din2(G41_n_spl_10)
  );


  LA
  g_g203_p
  (
    .dout(g203_p),
    .din1(G29_n_spl_0),
    .din2(G30_n_spl_0)
  );


  FA
  g_g203_n
  (
    .dout(g203_n),
    .din1(G29_p_spl_0),
    .din2(G30_p_spl_0)
  );


  LA
  g_g204_p
  (
    .dout(g204_p),
    .din1(G29_p_spl_1),
    .din2(G30_p_spl_1)
  );


  FA
  g_g204_n
  (
    .dout(g204_n),
    .din1(G29_n_spl_1),
    .din2(G30_n_spl_1)
  );


  LA
  g_g205_p
  (
    .dout(g205_p),
    .din1(g203_n),
    .din2(g204_n)
  );


  FA
  g_g205_n
  (
    .dout(g205_n),
    .din1(g203_p),
    .din2(g204_p)
  );


  LA
  g_g206_p
  (
    .dout(g206_p),
    .din1(G31_n_spl_0),
    .din2(G32_n_spl_0)
  );


  FA
  g_g206_n
  (
    .dout(g206_n),
    .din1(G31_p_spl_0),
    .din2(G32_p_spl_0)
  );


  LA
  g_g207_p
  (
    .dout(g207_p),
    .din1(G31_p_spl_1),
    .din2(G32_p_spl_1)
  );


  FA
  g_g207_n
  (
    .dout(g207_n),
    .din1(G31_n_spl_1),
    .din2(G32_n_spl_1)
  );


  LA
  g_g208_p
  (
    .dout(g208_p),
    .din1(g206_n),
    .din2(g207_n)
  );


  FA
  g_g208_n
  (
    .dout(g208_n),
    .din1(g206_p),
    .din2(g207_p)
  );


  LA
  g_g209_p
  (
    .dout(g209_p),
    .din1(g205_n_spl_),
    .din2(g208_p_spl_)
  );


  FA
  g_g209_n
  (
    .dout(g209_n),
    .din1(g205_p_spl_),
    .din2(g208_n_spl_)
  );


  LA
  g_g210_p
  (
    .dout(g210_p),
    .din1(g205_p_spl_),
    .din2(g208_n_spl_)
  );


  FA
  g_g210_n
  (
    .dout(g210_n),
    .din1(g205_n_spl_),
    .din2(g208_p_spl_)
  );


  LA
  g_g211_p
  (
    .dout(g211_p),
    .din1(g209_n),
    .din2(g210_n)
  );


  FA
  g_g211_n
  (
    .dout(g211_n),
    .din1(g209_p),
    .din2(g210_p)
  );


  LA
  g_g212_p
  (
    .dout(g212_p),
    .din1(g69_n_spl_1),
    .din2(g211_n_spl_0)
  );


  FA
  g_g212_n
  (
    .dout(g212_n),
    .din1(g69_p_spl_1),
    .din2(g211_p_spl_0)
  );


  LA
  g_g213_p
  (
    .dout(g213_p),
    .din1(g69_p_spl_1),
    .din2(g211_p_spl_0)
  );


  FA
  g_g213_n
  (
    .dout(g213_n),
    .din1(g69_n_spl_1),
    .din2(g211_n_spl_0)
  );


  LA
  g_g214_p
  (
    .dout(g214_p),
    .din1(g212_n),
    .din2(g213_n)
  );


  FA
  g_g214_n
  (
    .dout(g214_n),
    .din1(g212_p),
    .din2(g213_p)
  );


  LA
  g_g215_p
  (
    .dout(g215_p),
    .din1(g202_n_spl_),
    .din2(g214_p_spl_)
  );


  FA
  g_g215_n
  (
    .dout(g215_n),
    .din1(g202_p_spl_),
    .din2(g214_n_spl_)
  );


  LA
  g_g216_p
  (
    .dout(g216_p),
    .din1(g202_p_spl_),
    .din2(g214_n_spl_)
  );


  FA
  g_g216_n
  (
    .dout(g216_n),
    .din1(g202_n_spl_),
    .din2(g214_p_spl_)
  );


  LA
  g_g217_p
  (
    .dout(g217_p),
    .din1(g215_n),
    .din2(g216_n)
  );


  FA
  g_g217_n
  (
    .dout(g217_n),
    .din1(g215_p),
    .din2(g216_p)
  );


  LA
  g_g218_p
  (
    .dout(g218_p),
    .din1(g201_p_spl_),
    .din2(g217_n_spl_)
  );


  FA
  g_g218_n
  (
    .dout(g218_n),
    .din1(g201_n_spl_),
    .din2(g217_p_spl_)
  );


  LA
  g_g219_p
  (
    .dout(g219_p),
    .din1(g201_n_spl_),
    .din2(g217_p_spl_)
  );


  FA
  g_g219_n
  (
    .dout(g219_n),
    .din1(g201_p_spl_),
    .din2(g217_n_spl_)
  );


  LA
  g_g220_p
  (
    .dout(g220_p),
    .din1(g218_n),
    .din2(g219_n)
  );


  FA
  g_g220_n
  (
    .dout(g220_n),
    .din1(g218_p),
    .din2(g219_p)
  );


  LA
  g_g221_p
  (
    .dout(g221_p),
    .din1(G3_n_spl_0),
    .din2(G7_n_spl_0)
  );


  FA
  g_g221_n
  (
    .dout(g221_n),
    .din1(G3_p_spl_0),
    .din2(G7_p_spl_0)
  );


  LA
  g_g222_p
  (
    .dout(g222_p),
    .din1(G3_p_spl_1),
    .din2(G7_p_spl_1)
  );


  FA
  g_g222_n
  (
    .dout(g222_n),
    .din1(G3_n_spl_1),
    .din2(G7_n_spl_1)
  );


  LA
  g_g223_p
  (
    .dout(g223_p),
    .din1(g221_n),
    .din2(g222_n)
  );


  FA
  g_g223_n
  (
    .dout(g223_n),
    .din1(g221_p),
    .din2(g222_p)
  );


  LA
  g_g224_p
  (
    .dout(g224_p),
    .din1(G11_n_spl_0),
    .din2(G15_n_spl_0)
  );


  FA
  g_g224_n
  (
    .dout(g224_n),
    .din1(G11_p_spl_0),
    .din2(G15_p_spl_0)
  );


  LA
  g_g225_p
  (
    .dout(g225_p),
    .din1(G11_p_spl_1),
    .din2(G15_p_spl_1)
  );


  FA
  g_g225_n
  (
    .dout(g225_n),
    .din1(G11_n_spl_1),
    .din2(G15_n_spl_1)
  );


  LA
  g_g226_p
  (
    .dout(g226_p),
    .din1(g224_n),
    .din2(g225_n)
  );


  FA
  g_g226_n
  (
    .dout(g226_n),
    .din1(g224_p),
    .din2(g225_p)
  );


  LA
  g_g227_p
  (
    .dout(g227_p),
    .din1(g223_n_spl_),
    .din2(g226_p_spl_)
  );


  FA
  g_g227_n
  (
    .dout(g227_n),
    .din1(g223_p_spl_),
    .din2(g226_n_spl_)
  );


  LA
  g_g228_p
  (
    .dout(g228_p),
    .din1(g223_p_spl_),
    .din2(g226_n_spl_)
  );


  FA
  g_g228_n
  (
    .dout(g228_n),
    .din1(g223_n_spl_),
    .din2(g226_p_spl_)
  );


  LA
  g_g229_p
  (
    .dout(g229_p),
    .din1(g227_n),
    .din2(g228_n)
  );


  FA
  g_g229_n
  (
    .dout(g229_n),
    .din1(g227_p),
    .din2(g228_p)
  );


  LA
  g_g230_p
  (
    .dout(g230_p),
    .din1(G35_p),
    .din2(G41_p_spl_11)
  );


  FA
  g_g230_n
  (
    .dout(g230_n),
    .din1(G35_n),
    .din2(G41_n_spl_11)
  );


  LA
  g_g231_p
  (
    .dout(g231_p),
    .din1(G25_n_spl_0),
    .din2(G26_n_spl_0)
  );


  FA
  g_g231_n
  (
    .dout(g231_n),
    .din1(G25_p_spl_0),
    .din2(G26_p_spl_0)
  );


  LA
  g_g232_p
  (
    .dout(g232_p),
    .din1(G25_p_spl_1),
    .din2(G26_p_spl_1)
  );


  FA
  g_g232_n
  (
    .dout(g232_n),
    .din1(G25_n_spl_1),
    .din2(G26_n_spl_1)
  );


  LA
  g_g233_p
  (
    .dout(g233_p),
    .din1(g231_n),
    .din2(g232_n)
  );


  FA
  g_g233_n
  (
    .dout(g233_n),
    .din1(g231_p),
    .din2(g232_p)
  );


  LA
  g_g234_p
  (
    .dout(g234_p),
    .din1(G27_n_spl_0),
    .din2(G28_n_spl_0)
  );


  FA
  g_g234_n
  (
    .dout(g234_n),
    .din1(G27_p_spl_0),
    .din2(G28_p_spl_0)
  );


  LA
  g_g235_p
  (
    .dout(g235_p),
    .din1(G27_p_spl_1),
    .din2(G28_p_spl_1)
  );


  FA
  g_g235_n
  (
    .dout(g235_n),
    .din1(G27_n_spl_1),
    .din2(G28_n_spl_1)
  );


  LA
  g_g236_p
  (
    .dout(g236_p),
    .din1(g234_n),
    .din2(g235_n)
  );


  FA
  g_g236_n
  (
    .dout(g236_n),
    .din1(g234_p),
    .din2(g235_p)
  );


  LA
  g_g237_p
  (
    .dout(g237_p),
    .din1(g233_n_spl_),
    .din2(g236_p_spl_)
  );


  FA
  g_g237_n
  (
    .dout(g237_n),
    .din1(g233_p_spl_),
    .din2(g236_n_spl_)
  );


  LA
  g_g238_p
  (
    .dout(g238_p),
    .din1(g233_p_spl_),
    .din2(g236_n_spl_)
  );


  FA
  g_g238_n
  (
    .dout(g238_n),
    .din1(g233_n_spl_),
    .din2(g236_p_spl_)
  );


  LA
  g_g239_p
  (
    .dout(g239_p),
    .din1(g237_n),
    .din2(g238_n)
  );


  FA
  g_g239_n
  (
    .dout(g239_n),
    .din1(g237_p),
    .din2(g238_p)
  );


  LA
  g_g240_p
  (
    .dout(g240_p),
    .din1(g60_n_spl_1),
    .din2(g239_n_spl_0)
  );


  FA
  g_g240_n
  (
    .dout(g240_n),
    .din1(g60_p_spl_1),
    .din2(g239_p_spl_0)
  );


  LA
  g_g241_p
  (
    .dout(g241_p),
    .din1(g60_p_spl_1),
    .din2(g239_p_spl_0)
  );


  FA
  g_g241_n
  (
    .dout(g241_n),
    .din1(g60_n_spl_1),
    .din2(g239_n_spl_0)
  );


  LA
  g_g242_p
  (
    .dout(g242_p),
    .din1(g240_n),
    .din2(g241_n)
  );


  FA
  g_g242_n
  (
    .dout(g242_n),
    .din1(g240_p),
    .din2(g241_p)
  );


  LA
  g_g243_p
  (
    .dout(g243_p),
    .din1(g230_n_spl_),
    .din2(g242_p_spl_)
  );


  FA
  g_g243_n
  (
    .dout(g243_n),
    .din1(g230_p_spl_),
    .din2(g242_n_spl_)
  );


  LA
  g_g244_p
  (
    .dout(g244_p),
    .din1(g230_p_spl_),
    .din2(g242_n_spl_)
  );


  FA
  g_g244_n
  (
    .dout(g244_n),
    .din1(g230_n_spl_),
    .din2(g242_p_spl_)
  );


  LA
  g_g245_p
  (
    .dout(g245_p),
    .din1(g243_n),
    .din2(g244_n)
  );


  FA
  g_g245_n
  (
    .dout(g245_n),
    .din1(g243_p),
    .din2(g244_p)
  );


  LA
  g_g246_p
  (
    .dout(g246_p),
    .din1(g229_p_spl_),
    .din2(g245_n_spl_)
  );


  FA
  g_g246_n
  (
    .dout(g246_n),
    .din1(g229_n_spl_),
    .din2(g245_p_spl_)
  );


  LA
  g_g247_p
  (
    .dout(g247_p),
    .din1(g229_n_spl_),
    .din2(g245_p_spl_)
  );


  FA
  g_g247_n
  (
    .dout(g247_n),
    .din1(g229_p_spl_),
    .din2(g245_n_spl_)
  );


  LA
  g_g248_p
  (
    .dout(g248_p),
    .din1(g246_n),
    .din2(g247_n)
  );


  FA
  g_g248_n
  (
    .dout(g248_n),
    .din1(g246_p),
    .din2(g247_p)
  );


  LA
  g_g249_p
  (
    .dout(g249_p),
    .din1(G2_n_spl_0),
    .din2(G6_n_spl_0)
  );


  FA
  g_g249_n
  (
    .dout(g249_n),
    .din1(G2_p_spl_0),
    .din2(G6_p_spl_0)
  );


  LA
  g_g250_p
  (
    .dout(g250_p),
    .din1(G2_p_spl_1),
    .din2(G6_p_spl_1)
  );


  FA
  g_g250_n
  (
    .dout(g250_n),
    .din1(G2_n_spl_1),
    .din2(G6_n_spl_1)
  );


  LA
  g_g251_p
  (
    .dout(g251_p),
    .din1(g249_n),
    .din2(g250_n)
  );


  FA
  g_g251_n
  (
    .dout(g251_n),
    .din1(g249_p),
    .din2(g250_p)
  );


  LA
  g_g252_p
  (
    .dout(g252_p),
    .din1(G10_n_spl_0),
    .din2(G14_n_spl_0)
  );


  FA
  g_g252_n
  (
    .dout(g252_n),
    .din1(G10_p_spl_0),
    .din2(G14_p_spl_0)
  );


  LA
  g_g253_p
  (
    .dout(g253_p),
    .din1(G10_p_spl_1),
    .din2(G14_p_spl_1)
  );


  FA
  g_g253_n
  (
    .dout(g253_n),
    .din1(G10_n_spl_1),
    .din2(G14_n_spl_1)
  );


  LA
  g_g254_p
  (
    .dout(g254_p),
    .din1(g252_n),
    .din2(g253_n)
  );


  FA
  g_g254_n
  (
    .dout(g254_n),
    .din1(g252_p),
    .din2(g253_p)
  );


  LA
  g_g255_p
  (
    .dout(g255_p),
    .din1(g251_n_spl_),
    .din2(g254_p_spl_)
  );


  FA
  g_g255_n
  (
    .dout(g255_n),
    .din1(g251_p_spl_),
    .din2(g254_n_spl_)
  );


  LA
  g_g256_p
  (
    .dout(g256_p),
    .din1(g251_p_spl_),
    .din2(g254_n_spl_)
  );


  FA
  g_g256_n
  (
    .dout(g256_n),
    .din1(g251_n_spl_),
    .din2(g254_p_spl_)
  );


  LA
  g_g257_p
  (
    .dout(g257_p),
    .din1(g255_n),
    .din2(g256_n)
  );


  FA
  g_g257_n
  (
    .dout(g257_n),
    .din1(g255_p),
    .din2(g256_p)
  );


  LA
  g_g258_p
  (
    .dout(g258_p),
    .din1(G34_p),
    .din2(G41_p_spl_11)
  );


  FA
  g_g258_n
  (
    .dout(g258_n),
    .din1(G34_n),
    .din2(G41_n_spl_11)
  );


  LA
  g_g259_p
  (
    .dout(g259_p),
    .din1(g211_n_spl_1),
    .din2(g239_n_spl_1)
  );


  FA
  g_g259_n
  (
    .dout(g259_n),
    .din1(g211_p_spl_1),
    .din2(g239_p_spl_1)
  );


  LA
  g_g260_p
  (
    .dout(g260_p),
    .din1(g211_p_spl_1),
    .din2(g239_p_spl_1)
  );


  FA
  g_g260_n
  (
    .dout(g260_n),
    .din1(g211_n_spl_1),
    .din2(g239_n_spl_1)
  );


  LA
  g_g261_p
  (
    .dout(g261_p),
    .din1(g259_n),
    .din2(g260_n)
  );


  FA
  g_g261_n
  (
    .dout(g261_n),
    .din1(g259_p),
    .din2(g260_p)
  );


  LA
  g_g262_p
  (
    .dout(g262_p),
    .din1(g258_n_spl_),
    .din2(g261_p_spl_)
  );


  FA
  g_g262_n
  (
    .dout(g262_n),
    .din1(g258_p_spl_),
    .din2(g261_n_spl_)
  );


  LA
  g_g263_p
  (
    .dout(g263_p),
    .din1(g258_p_spl_),
    .din2(g261_n_spl_)
  );


  FA
  g_g263_n
  (
    .dout(g263_n),
    .din1(g258_n_spl_),
    .din2(g261_p_spl_)
  );


  LA
  g_g264_p
  (
    .dout(g264_p),
    .din1(g262_n),
    .din2(g263_n)
  );


  FA
  g_g264_n
  (
    .dout(g264_n),
    .din1(g262_p),
    .din2(g263_p)
  );


  LA
  g_g265_p
  (
    .dout(g265_p),
    .din1(g257_p_spl_),
    .din2(g264_n_spl_)
  );


  FA
  g_g265_n
  (
    .dout(g265_n),
    .din1(g257_n_spl_),
    .din2(g264_p_spl_)
  );


  LA
  g_g266_p
  (
    .dout(g266_p),
    .din1(g257_n_spl_),
    .din2(g264_p_spl_)
  );


  FA
  g_g266_n
  (
    .dout(g266_n),
    .din1(g257_p_spl_),
    .din2(g264_n_spl_)
  );


  LA
  g_g267_p
  (
    .dout(g267_p),
    .din1(g265_n),
    .din2(g266_n)
  );


  FA
  g_g267_n
  (
    .dout(g267_n),
    .din1(g265_p),
    .din2(g266_p)
  );


  LA
  g_g268_p
  (
    .dout(g268_p),
    .din1(g78_n_spl_00),
    .din2(g267_p_spl_00)
  );


  FA
  g_g268_n
  (
    .dout(g268_n),
    .din1(g78_p_spl_00),
    .din2(g267_n_spl_00)
  );


  LA
  g_g269_p
  (
    .dout(g269_p),
    .din1(g248_p_spl_00),
    .din2(g268_p_spl_)
  );


  FA
  g_g269_n
  (
    .dout(g269_n),
    .din1(g248_n_spl_00),
    .din2(g268_n_spl_)
  );


  LA
  g_g270_p
  (
    .dout(g270_p),
    .din1(g78_p_spl_00),
    .din2(g267_n_spl_00)
  );


  FA
  g_g270_n
  (
    .dout(g270_n),
    .din1(g78_n_spl_00),
    .din2(g267_p_spl_00)
  );


  LA
  g_g271_p
  (
    .dout(g271_p),
    .din1(g248_p_spl_00),
    .din2(g270_p_spl_)
  );


  FA
  g_g271_n
  (
    .dout(g271_n),
    .din1(g248_n_spl_00),
    .din2(g270_n_spl_)
  );


  LA
  g_g272_p
  (
    .dout(g272_p),
    .din1(g269_n_spl_),
    .din2(g271_n_spl_)
  );


  FA
  g_g272_n
  (
    .dout(g272_n),
    .din1(g269_p_spl_),
    .din2(g271_p_spl_)
  );


  LA
  g_g273_p
  (
    .dout(g273_p),
    .din1(g220_p_spl_00),
    .din2(g272_n)
  );


  FA
  g_g273_n
  (
    .dout(g273_n),
    .din1(g220_n_spl_00),
    .din2(g272_p)
  );


  LA
  g_g274_p
  (
    .dout(g274_p),
    .din1(g220_p_spl_00),
    .din2(g248_n_spl_01)
  );


  FA
  g_g274_n
  (
    .dout(g274_n),
    .din1(g220_n_spl_00),
    .din2(g248_p_spl_01)
  );


  LA
  g_g275_p
  (
    .dout(g275_p),
    .din1(g220_n_spl_01),
    .din2(g248_p_spl_01)
  );


  FA
  g_g275_n
  (
    .dout(g275_n),
    .din1(g220_p_spl_01),
    .din2(g248_n_spl_01)
  );


  LA
  g_g276_p
  (
    .dout(g276_p),
    .din1(g274_n_spl_0),
    .din2(g275_n)
  );


  FA
  g_g276_n
  (
    .dout(g276_n),
    .din1(g274_p_spl_0),
    .din2(g275_p)
  );


  LA
  g_g277_p
  (
    .dout(g277_p),
    .din1(g267_p_spl_01),
    .din2(g276_n)
  );


  FA
  g_g277_n
  (
    .dout(g277_n),
    .din1(g267_n_spl_01),
    .din2(g276_p)
  );


  LA
  g_g278_p
  (
    .dout(g278_p),
    .din1(g78_p_spl_01),
    .din2(g277_p)
  );


  FA
  g_g278_n
  (
    .dout(g278_n),
    .din1(g78_n_spl_01),
    .din2(g277_n)
  );


  LA
  g_g279_p
  (
    .dout(g279_p),
    .din1(g273_n),
    .din2(g278_n)
  );


  FA
  g_g279_n
  (
    .dout(g279_n),
    .din1(g273_p),
    .din2(g278_p)
  );


  LA
  g_g280_p
  (
    .dout(g280_p),
    .din1(g192_p_spl_),
    .din2(g279_n_spl_)
  );


  FA
  g_g280_n
  (
    .dout(g280_n),
    .din1(g192_n_spl_),
    .din2(g279_p_spl_)
  );


  LA
  g_g281_p
  (
    .dout(g281_p),
    .din1(g153_p_spl_),
    .din2(g280_p_spl_)
  );


  FA
  g_g281_n
  (
    .dout(g281_n),
    .din1(g153_n_spl_),
    .din2(g280_n_spl_)
  );


  LA
  g_g282_p
  (
    .dout(g282_p),
    .din1(g78_n_spl_01),
    .din2(g281_p_spl_0)
  );


  FA
  g_g282_n
  (
    .dout(g282_n),
    .din1(g78_p_spl_01),
    .din2(g281_n_spl_0)
  );


  FA
  g_g283_n
  (
    .dout(g283_n),
    .din1(G1_p_spl_1),
    .din2(g282_n)
  );


  FA
  g_g284_n
  (
    .dout(g284_n),
    .din1(G1_n_spl_1),
    .din2(g282_p)
  );


  LA
  g_g285_p
  (
    .dout(g285_p),
    .din1(g283_n),
    .din2(g284_n)
  );


  LA
  g_g286_p
  (
    .dout(g286_p),
    .din1(g267_n_spl_01),
    .din2(g281_p_spl_0)
  );


  FA
  g_g286_n
  (
    .dout(g286_n),
    .din1(g267_p_spl_01),
    .din2(g281_n_spl_0)
  );


  FA
  g_g287_n
  (
    .dout(g287_n),
    .din1(G2_p_spl_1),
    .din2(g286_n)
  );


  FA
  g_g288_n
  (
    .dout(g288_n),
    .din1(G2_n_spl_1),
    .din2(g286_p)
  );


  LA
  g_g289_p
  (
    .dout(g289_p),
    .din1(g287_n),
    .din2(g288_n)
  );


  LA
  g_g290_p
  (
    .dout(g290_p),
    .din1(g248_n_spl_10),
    .din2(g281_p_spl_1)
  );


  FA
  g_g290_n
  (
    .dout(g290_n),
    .din1(g248_p_spl_10),
    .din2(g281_n_spl_1)
  );


  FA
  g_g291_n
  (
    .dout(g291_n),
    .din1(G3_p_spl_1),
    .din2(g290_n)
  );


  FA
  g_g292_n
  (
    .dout(g292_n),
    .din1(G3_n_spl_1),
    .din2(g290_p)
  );


  LA
  g_g293_p
  (
    .dout(g293_p),
    .din1(g291_n),
    .din2(g292_n)
  );


  LA
  g_g294_p
  (
    .dout(g294_p),
    .din1(g220_n_spl_01),
    .din2(g281_p_spl_1)
  );


  FA
  g_g294_n
  (
    .dout(g294_n),
    .din1(g220_p_spl_01),
    .din2(g281_n_spl_1)
  );


  FA
  g_g295_n
  (
    .dout(g295_n),
    .din1(G4_p_spl_1),
    .din2(g294_n)
  );


  FA
  g_g296_n
  (
    .dout(g296_n),
    .din1(G4_n_spl_1),
    .din2(g294_p)
  );


  LA
  g_g297_p
  (
    .dout(g297_p),
    .din1(g295_n),
    .din2(g296_n)
  );


  LA
  g_g298_p
  (
    .dout(g298_p),
    .din1(g153_p_spl_),
    .din2(g191_p_spl_00)
  );


  FA
  g_g298_n
  (
    .dout(g298_n),
    .din1(g153_n_spl_),
    .din2(g191_n_spl_00)
  );


  LA
  g_g299_p
  (
    .dout(g299_p),
    .din1(g172_n_spl_00),
    .din2(g279_n_spl_)
  );


  FA
  g_g299_n
  (
    .dout(g299_n),
    .din1(g172_p_spl_00),
    .din2(g279_p_spl_)
  );


  LA
  g_g300_p
  (
    .dout(g300_p),
    .din1(g298_p_spl_),
    .din2(g299_p_spl_)
  );


  FA
  g_g300_n
  (
    .dout(g300_n),
    .din1(g298_n_spl_),
    .din2(g299_n_spl_)
  );


  LA
  g_g301_p
  (
    .dout(g301_p),
    .din1(g78_n_spl_10),
    .din2(g300_p_spl_0)
  );


  FA
  g_g301_n
  (
    .dout(g301_n),
    .din1(g78_p_spl_10),
    .din2(g300_n_spl_0)
  );


  FA
  g_g302_n
  (
    .dout(g302_n),
    .din1(G5_p_spl_1),
    .din2(g301_n)
  );


  FA
  g_g303_n
  (
    .dout(g303_n),
    .din1(G5_n_spl_1),
    .din2(g301_p)
  );


  LA
  g_g304_p
  (
    .dout(g304_p),
    .din1(g302_n),
    .din2(g303_n)
  );


  LA
  g_g305_p
  (
    .dout(g305_p),
    .din1(g267_n_spl_10),
    .din2(g300_p_spl_0)
  );


  FA
  g_g305_n
  (
    .dout(g305_n),
    .din1(g267_p_spl_10),
    .din2(g300_n_spl_0)
  );


  FA
  g_g306_n
  (
    .dout(g306_n),
    .din1(G6_p_spl_1),
    .din2(g305_n)
  );


  FA
  g_g307_n
  (
    .dout(g307_n),
    .din1(G6_n_spl_1),
    .din2(g305_p)
  );


  LA
  g_g308_p
  (
    .dout(g308_p),
    .din1(g306_n),
    .din2(g307_n)
  );


  LA
  g_g309_p
  (
    .dout(g309_p),
    .din1(g248_n_spl_10),
    .din2(g300_p_spl_1)
  );


  FA
  g_g309_n
  (
    .dout(g309_n),
    .din1(g248_p_spl_10),
    .din2(g300_n_spl_1)
  );


  FA
  g_g310_n
  (
    .dout(g310_n),
    .din1(G7_p_spl_1),
    .din2(g309_n)
  );


  FA
  g_g311_n
  (
    .dout(g311_n),
    .din1(G7_n_spl_1),
    .din2(g309_p)
  );


  LA
  g_g312_p
  (
    .dout(g312_p),
    .din1(g310_n),
    .din2(g311_n)
  );


  LA
  g_g313_p
  (
    .dout(g313_p),
    .din1(g220_n_spl_10),
    .din2(g300_p_spl_1)
  );


  FA
  g_g313_n
  (
    .dout(g313_n),
    .din1(g220_p_spl_10),
    .din2(g300_n_spl_1)
  );


  FA
  g_g314_n
  (
    .dout(g314_n),
    .din1(G8_p_spl_1),
    .din2(g313_n)
  );


  FA
  g_g315_n
  (
    .dout(g315_n),
    .din1(G8_n_spl_1),
    .din2(g313_p)
  );


  LA
  g_g316_p
  (
    .dout(g316_p),
    .din1(g314_n),
    .din2(g315_n)
  );


  LA
  g_g317_p
  (
    .dout(g317_p),
    .din1(g115_p_spl_00),
    .din2(g152_n_spl_00)
  );


  FA
  g_g317_n
  (
    .dout(g317_n),
    .din1(g115_n_spl_00),
    .din2(g152_p_spl_00)
  );


  LA
  g_g318_p
  (
    .dout(g318_p),
    .din1(g280_p_spl_),
    .din2(g317_p_spl_)
  );


  FA
  g_g318_n
  (
    .dout(g318_n),
    .din1(g280_n_spl_),
    .din2(g317_n_spl_)
  );


  LA
  g_g319_p
  (
    .dout(g319_p),
    .din1(g78_n_spl_10),
    .din2(g318_p_spl_0)
  );


  FA
  g_g319_n
  (
    .dout(g319_n),
    .din1(g78_p_spl_10),
    .din2(g318_n_spl_0)
  );


  FA
  g_g320_n
  (
    .dout(g320_n),
    .din1(G9_p_spl_1),
    .din2(g319_n)
  );


  FA
  g_g321_n
  (
    .dout(g321_n),
    .din1(G9_n_spl_1),
    .din2(g319_p)
  );


  LA
  g_g322_p
  (
    .dout(g322_p),
    .din1(g320_n),
    .din2(g321_n)
  );


  LA
  g_g323_p
  (
    .dout(g323_p),
    .din1(g267_n_spl_10),
    .din2(g318_p_spl_0)
  );


  FA
  g_g323_n
  (
    .dout(g323_n),
    .din1(g267_p_spl_10),
    .din2(g318_n_spl_0)
  );


  FA
  g_g324_n
  (
    .dout(g324_n),
    .din1(G10_p_spl_1),
    .din2(g323_n)
  );


  FA
  g_g325_n
  (
    .dout(g325_n),
    .din1(G10_n_spl_1),
    .din2(g323_p)
  );


  LA
  g_g326_p
  (
    .dout(g326_p),
    .din1(g324_n),
    .din2(g325_n)
  );


  LA
  g_g327_p
  (
    .dout(g327_p),
    .din1(g248_n_spl_11),
    .din2(g318_p_spl_1)
  );


  FA
  g_g327_n
  (
    .dout(g327_n),
    .din1(g248_p_spl_11),
    .din2(g318_n_spl_1)
  );


  FA
  g_g328_n
  (
    .dout(g328_n),
    .din1(G11_p_spl_1),
    .din2(g327_n)
  );


  FA
  g_g329_n
  (
    .dout(g329_n),
    .din1(G11_n_spl_1),
    .din2(g327_p)
  );


  LA
  g_g330_p
  (
    .dout(g330_p),
    .din1(g328_n),
    .din2(g329_n)
  );


  LA
  g_g331_p
  (
    .dout(g331_p),
    .din1(g220_n_spl_10),
    .din2(g318_p_spl_1)
  );


  FA
  g_g331_n
  (
    .dout(g331_n),
    .din1(g220_p_spl_10),
    .din2(g318_n_spl_1)
  );


  FA
  g_g332_n
  (
    .dout(g332_n),
    .din1(G12_p_spl_1),
    .din2(g331_n)
  );


  FA
  g_g333_n
  (
    .dout(g333_n),
    .din1(G12_n_spl_1),
    .din2(g331_p)
  );


  LA
  g_g334_p
  (
    .dout(g334_p),
    .din1(g332_n),
    .din2(g333_n)
  );


  LA
  g_g335_p
  (
    .dout(g335_p),
    .din1(g191_p_spl_01),
    .din2(g317_p_spl_)
  );


  FA
  g_g335_n
  (
    .dout(g335_n),
    .din1(g191_n_spl_01),
    .din2(g317_n_spl_)
  );


  LA
  g_g336_p
  (
    .dout(g336_p),
    .din1(g299_p_spl_),
    .din2(g335_p_spl_)
  );


  FA
  g_g336_n
  (
    .dout(g336_n),
    .din1(g299_n_spl_),
    .din2(g335_n_spl_)
  );


  LA
  g_g337_p
  (
    .dout(g337_p),
    .din1(g78_n_spl_1),
    .din2(g336_p_spl_0)
  );


  FA
  g_g337_n
  (
    .dout(g337_n),
    .din1(g78_p_spl_1),
    .din2(g336_n_spl_0)
  );


  FA
  g_g338_n
  (
    .dout(g338_n),
    .din1(G13_p_spl_1),
    .din2(g337_n)
  );


  FA
  g_g339_n
  (
    .dout(g339_n),
    .din1(G13_n_spl_1),
    .din2(g337_p)
  );


  LA
  g_g340_p
  (
    .dout(g340_p),
    .din1(g338_n),
    .din2(g339_n)
  );


  LA
  g_g341_p
  (
    .dout(g341_p),
    .din1(g267_n_spl_1),
    .din2(g336_p_spl_0)
  );


  FA
  g_g341_n
  (
    .dout(g341_n),
    .din1(g267_p_spl_1),
    .din2(g336_n_spl_0)
  );


  FA
  g_g342_n
  (
    .dout(g342_n),
    .din1(G14_p_spl_1),
    .din2(g341_n)
  );


  FA
  g_g343_n
  (
    .dout(g343_n),
    .din1(G14_n_spl_1),
    .din2(g341_p)
  );


  LA
  g_g344_p
  (
    .dout(g344_p),
    .din1(g342_n),
    .din2(g343_n)
  );


  LA
  g_g345_p
  (
    .dout(g345_p),
    .din1(g248_n_spl_11),
    .din2(g336_p_spl_1)
  );


  FA
  g_g345_n
  (
    .dout(g345_n),
    .din1(g248_p_spl_11),
    .din2(g336_n_spl_1)
  );


  FA
  g_g346_n
  (
    .dout(g346_n),
    .din1(G15_p_spl_1),
    .din2(g345_n)
  );


  FA
  g_g347_n
  (
    .dout(g347_n),
    .din1(G15_n_spl_1),
    .din2(g345_p)
  );


  LA
  g_g348_p
  (
    .dout(g348_p),
    .din1(g346_n),
    .din2(g347_n)
  );


  LA
  g_g349_p
  (
    .dout(g349_p),
    .din1(g220_n_spl_11),
    .din2(g336_p_spl_1)
  );


  FA
  g_g349_n
  (
    .dout(g349_n),
    .din1(g220_p_spl_11),
    .din2(g336_n_spl_1)
  );


  FA
  g_g350_n
  (
    .dout(g350_n),
    .din1(G16_p_spl_1),
    .din2(g349_n)
  );


  FA
  g_g351_n
  (
    .dout(g351_n),
    .din1(G16_n_spl_1),
    .din2(g349_p)
  );


  LA
  g_g352_p
  (
    .dout(g352_p),
    .din1(g350_n),
    .din2(g351_n)
  );


  LA
  g_g353_p
  (
    .dout(g353_p),
    .din1(g298_n_spl_),
    .din2(g335_n_spl_)
  );


  FA
  g_g353_n
  (
    .dout(g353_n),
    .din1(g298_p_spl_),
    .din2(g335_p_spl_)
  );


  LA
  g_g354_p
  (
    .dout(g354_p),
    .din1(g172_p_spl_01),
    .din2(g353_n)
  );


  FA
  g_g354_n
  (
    .dout(g354_n),
    .din1(g172_n_spl_01),
    .din2(g353_p)
  );


  LA
  g_g355_p
  (
    .dout(g355_p),
    .din1(g172_n_spl_01),
    .din2(g191_p_spl_01)
  );


  FA
  g_g355_n
  (
    .dout(g355_n),
    .din1(g172_p_spl_01),
    .din2(g191_n_spl_01)
  );


  LA
  g_g356_p
  (
    .dout(g356_p),
    .din1(g192_n_spl_),
    .din2(g355_n)
  );


  FA
  g_g356_n
  (
    .dout(g356_n),
    .din1(g192_p_spl_),
    .din2(g355_p)
  );


  LA
  g_g357_p
  (
    .dout(g357_p),
    .din1(g152_p_spl_01),
    .din2(g356_n)
  );


  FA
  g_g357_n
  (
    .dout(g357_n),
    .din1(g152_n_spl_01),
    .din2(g356_p)
  );


  LA
  g_g358_p
  (
    .dout(g358_p),
    .din1(g115_p_spl_01),
    .din2(g357_p)
  );


  FA
  g_g358_n
  (
    .dout(g358_n),
    .din1(g115_n_spl_01),
    .din2(g357_n)
  );


  LA
  g_g359_p
  (
    .dout(g359_p),
    .din1(g354_n),
    .din2(g358_n)
  );


  FA
  g_g359_n
  (
    .dout(g359_n),
    .din1(g354_p),
    .din2(g358_p)
  );


  LA
  g_g360_p
  (
    .dout(g360_p),
    .din1(g268_p_spl_),
    .din2(g359_n_spl_0)
  );


  FA
  g_g360_n
  (
    .dout(g360_n),
    .din1(g268_n_spl_),
    .din2(g359_p_spl_0)
  );


  LA
  g_g361_p
  (
    .dout(g361_p),
    .din1(g274_p_spl_0),
    .din2(g360_p)
  );


  FA
  g_g361_n
  (
    .dout(g361_n),
    .din1(g274_n_spl_0),
    .din2(g360_n)
  );


  LA
  g_g362_p
  (
    .dout(g362_p),
    .din1(g115_n_spl_01),
    .din2(g361_p_spl_0)
  );


  FA
  g_g362_n
  (
    .dout(g362_n),
    .din1(g115_p_spl_01),
    .din2(g361_n_spl_0)
  );


  FA
  g_g363_n
  (
    .dout(g363_n),
    .din1(G17_p_spl_1),
    .din2(g362_n)
  );


  FA
  g_g364_n
  (
    .dout(g364_n),
    .din1(G17_n_spl_1),
    .din2(g362_p)
  );


  LA
  g_g365_p
  (
    .dout(g365_p),
    .din1(g363_n),
    .din2(g364_n)
  );


  LA
  g_g366_p
  (
    .dout(g366_p),
    .din1(g152_n_spl_01),
    .din2(g361_p_spl_0)
  );


  FA
  g_g366_n
  (
    .dout(g366_n),
    .din1(g152_p_spl_01),
    .din2(g361_n_spl_0)
  );


  FA
  g_g367_n
  (
    .dout(g367_n),
    .din1(G18_p_spl_1),
    .din2(g366_n)
  );


  FA
  g_g368_n
  (
    .dout(g368_n),
    .din1(G18_n_spl_1),
    .din2(g366_p)
  );


  LA
  g_g369_p
  (
    .dout(g369_p),
    .din1(g367_n),
    .din2(g368_n)
  );


  LA
  g_g370_p
  (
    .dout(g370_p),
    .din1(g191_n_spl_10),
    .din2(g361_p_spl_1)
  );


  FA
  g_g370_n
  (
    .dout(g370_n),
    .din1(g191_p_spl_10),
    .din2(g361_n_spl_1)
  );


  FA
  g_g371_n
  (
    .dout(g371_n),
    .din1(G19_p_spl_1),
    .din2(g370_n)
  );


  FA
  g_g372_n
  (
    .dout(g372_n),
    .din1(G19_n_spl_1),
    .din2(g370_p)
  );


  LA
  g_g373_p
  (
    .dout(g373_p),
    .din1(g371_n),
    .din2(g372_n)
  );


  LA
  g_g374_p
  (
    .dout(g374_p),
    .din1(g172_n_spl_10),
    .din2(g361_p_spl_1)
  );


  FA
  g_g374_n
  (
    .dout(g374_n),
    .din1(g172_p_spl_10),
    .din2(g361_n_spl_1)
  );


  FA
  g_g375_n
  (
    .dout(g375_n),
    .din1(G20_p_spl_1),
    .din2(g374_n)
  );


  FA
  g_g376_n
  (
    .dout(g376_n),
    .din1(G20_n_spl_1),
    .din2(g374_p)
  );


  LA
  g_g377_p
  (
    .dout(g377_p),
    .din1(g375_n),
    .din2(g376_n)
  );


  LA
  g_g378_p
  (
    .dout(g378_p),
    .din1(g220_n_spl_11),
    .din2(g359_n_spl_0)
  );


  FA
  g_g378_n
  (
    .dout(g378_n),
    .din1(g220_p_spl_11),
    .din2(g359_p_spl_0)
  );


  LA
  g_g379_p
  (
    .dout(g379_p),
    .din1(g269_p_spl_),
    .din2(g378_p_spl_)
  );


  FA
  g_g379_n
  (
    .dout(g379_n),
    .din1(g269_n_spl_),
    .din2(g378_n_spl_)
  );


  LA
  g_g380_p
  (
    .dout(g380_p),
    .din1(g115_n_spl_10),
    .din2(g379_p_spl_0)
  );


  FA
  g_g380_n
  (
    .dout(g380_n),
    .din1(g115_p_spl_10),
    .din2(g379_n_spl_0)
  );


  FA
  g_g381_n
  (
    .dout(g381_n),
    .din1(G21_p_spl_1),
    .din2(g380_n)
  );


  FA
  g_g382_n
  (
    .dout(g382_n),
    .din1(G21_n_spl_1),
    .din2(g380_p)
  );


  LA
  g_g383_p
  (
    .dout(g383_p),
    .din1(g381_n),
    .din2(g382_n)
  );


  LA
  g_g384_p
  (
    .dout(g384_p),
    .din1(g152_n_spl_10),
    .din2(g379_p_spl_0)
  );


  FA
  g_g384_n
  (
    .dout(g384_n),
    .din1(g152_p_spl_10),
    .din2(g379_n_spl_0)
  );


  FA
  g_g385_n
  (
    .dout(g385_n),
    .din1(G22_p_spl_1),
    .din2(g384_n)
  );


  FA
  g_g386_n
  (
    .dout(g386_n),
    .din1(G22_n_spl_1),
    .din2(g384_p)
  );


  LA
  g_g387_p
  (
    .dout(g387_p),
    .din1(g385_n),
    .din2(g386_n)
  );


  LA
  g_g388_p
  (
    .dout(g388_p),
    .din1(g191_n_spl_10),
    .din2(g379_p_spl_1)
  );


  FA
  g_g388_n
  (
    .dout(g388_n),
    .din1(g191_p_spl_10),
    .din2(g379_n_spl_1)
  );


  FA
  g_g389_n
  (
    .dout(g389_n),
    .din1(G23_p_spl_1),
    .din2(g388_n)
  );


  FA
  g_g390_n
  (
    .dout(g390_n),
    .din1(G23_n_spl_1),
    .din2(g388_p)
  );


  LA
  g_g391_p
  (
    .dout(g391_p),
    .din1(g389_n),
    .din2(g390_n)
  );


  LA
  g_g392_p
  (
    .dout(g392_p),
    .din1(g172_n_spl_10),
    .din2(g379_p_spl_1)
  );


  FA
  g_g392_n
  (
    .dout(g392_n),
    .din1(g172_p_spl_10),
    .din2(g379_n_spl_1)
  );


  FA
  g_g393_n
  (
    .dout(g393_n),
    .din1(G24_p_spl_1),
    .din2(g392_n)
  );


  FA
  g_g394_n
  (
    .dout(g394_n),
    .din1(G24_n_spl_1),
    .din2(g392_p)
  );


  LA
  g_g395_p
  (
    .dout(g395_p),
    .din1(g393_n),
    .din2(g394_n)
  );


  LA
  g_g396_p
  (
    .dout(g396_p),
    .din1(g270_p_spl_),
    .din2(g359_n_spl_)
  );


  FA
  g_g396_n
  (
    .dout(g396_n),
    .din1(g270_n_spl_),
    .din2(g359_p_spl_)
  );


  LA
  g_g397_p
  (
    .dout(g397_p),
    .din1(g274_p_spl_),
    .din2(g396_p)
  );


  FA
  g_g397_n
  (
    .dout(g397_n),
    .din1(g274_n_spl_),
    .din2(g396_n)
  );


  LA
  g_g398_p
  (
    .dout(g398_p),
    .din1(g115_n_spl_10),
    .din2(g397_p_spl_0)
  );


  FA
  g_g398_n
  (
    .dout(g398_n),
    .din1(g115_p_spl_10),
    .din2(g397_n_spl_0)
  );


  FA
  g_g399_n
  (
    .dout(g399_n),
    .din1(G25_p_spl_1),
    .din2(g398_n)
  );


  FA
  g_g400_n
  (
    .dout(g400_n),
    .din1(G25_n_spl_1),
    .din2(g398_p)
  );


  LA
  g_g401_p
  (
    .dout(g401_p),
    .din1(g399_n),
    .din2(g400_n)
  );


  LA
  g_g402_p
  (
    .dout(g402_p),
    .din1(g152_n_spl_10),
    .din2(g397_p_spl_0)
  );


  FA
  g_g402_n
  (
    .dout(g402_n),
    .din1(g152_p_spl_10),
    .din2(g397_n_spl_0)
  );


  FA
  g_g403_n
  (
    .dout(g403_n),
    .din1(G26_p_spl_1),
    .din2(g402_n)
  );


  FA
  g_g404_n
  (
    .dout(g404_n),
    .din1(G26_n_spl_1),
    .din2(g402_p)
  );


  LA
  g_g405_p
  (
    .dout(g405_p),
    .din1(g403_n),
    .din2(g404_n)
  );


  LA
  g_g406_p
  (
    .dout(g406_p),
    .din1(g191_n_spl_11),
    .din2(g397_p_spl_1)
  );


  FA
  g_g406_n
  (
    .dout(g406_n),
    .din1(g191_p_spl_11),
    .din2(g397_n_spl_1)
  );


  FA
  g_g407_n
  (
    .dout(g407_n),
    .din1(G27_p_spl_1),
    .din2(g406_n)
  );


  FA
  g_g408_n
  (
    .dout(g408_n),
    .din1(G27_n_spl_1),
    .din2(g406_p)
  );


  LA
  g_g409_p
  (
    .dout(g409_p),
    .din1(g407_n),
    .din2(g408_n)
  );


  LA
  g_g410_p
  (
    .dout(g410_p),
    .din1(g172_n_spl_11),
    .din2(g397_p_spl_1)
  );


  FA
  g_g410_n
  (
    .dout(g410_n),
    .din1(g172_p_spl_11),
    .din2(g397_n_spl_1)
  );


  FA
  g_g411_n
  (
    .dout(g411_n),
    .din1(G28_p_spl_1),
    .din2(g410_n)
  );


  FA
  g_g412_n
  (
    .dout(g412_n),
    .din1(G28_n_spl_1),
    .din2(g410_p)
  );


  LA
  g_g413_p
  (
    .dout(g413_p),
    .din1(g411_n),
    .din2(g412_n)
  );


  LA
  g_g414_p
  (
    .dout(g414_p),
    .din1(g271_p_spl_),
    .din2(g378_p_spl_)
  );


  FA
  g_g414_n
  (
    .dout(g414_n),
    .din1(g271_n_spl_),
    .din2(g378_n_spl_)
  );


  LA
  g_g415_p
  (
    .dout(g415_p),
    .din1(g115_n_spl_1),
    .din2(g414_p_spl_0)
  );


  FA
  g_g415_n
  (
    .dout(g415_n),
    .din1(g115_p_spl_1),
    .din2(g414_n_spl_0)
  );


  FA
  g_g416_n
  (
    .dout(g416_n),
    .din1(G29_p_spl_1),
    .din2(g415_n)
  );


  FA
  g_g417_n
  (
    .dout(g417_n),
    .din1(G29_n_spl_1),
    .din2(g415_p)
  );


  LA
  g_g418_p
  (
    .dout(g418_p),
    .din1(g416_n),
    .din2(g417_n)
  );


  LA
  g_g419_p
  (
    .dout(g419_p),
    .din1(g152_n_spl_1),
    .din2(g414_p_spl_0)
  );


  FA
  g_g419_n
  (
    .dout(g419_n),
    .din1(g152_p_spl_1),
    .din2(g414_n_spl_0)
  );


  FA
  g_g420_n
  (
    .dout(g420_n),
    .din1(G30_p_spl_1),
    .din2(g419_n)
  );


  FA
  g_g421_n
  (
    .dout(g421_n),
    .din1(G30_n_spl_1),
    .din2(g419_p)
  );


  LA
  g_g422_p
  (
    .dout(g422_p),
    .din1(g420_n),
    .din2(g421_n)
  );


  LA
  g_g423_p
  (
    .dout(g423_p),
    .din1(g191_n_spl_11),
    .din2(g414_p_spl_1)
  );


  FA
  g_g423_n
  (
    .dout(g423_n),
    .din1(g191_p_spl_11),
    .din2(g414_n_spl_1)
  );


  FA
  g_g424_n
  (
    .dout(g424_n),
    .din1(G31_p_spl_1),
    .din2(g423_n)
  );


  FA
  g_g425_n
  (
    .dout(g425_n),
    .din1(G31_n_spl_1),
    .din2(g423_p)
  );


  LA
  g_g426_p
  (
    .dout(g426_p),
    .din1(g424_n),
    .din2(g425_n)
  );


  LA
  g_g427_p
  (
    .dout(g427_p),
    .din1(g172_n_spl_11),
    .din2(g414_p_spl_1)
  );


  FA
  g_g427_n
  (
    .dout(g427_n),
    .din1(g172_p_spl_11),
    .din2(g414_n_spl_1)
  );


  FA
  g_g428_n
  (
    .dout(g428_n),
    .din1(G32_p_spl_1),
    .din2(g427_n)
  );


  FA
  g_g429_n
  (
    .dout(g429_n),
    .din1(G32_n_spl_1),
    .din2(g427_p)
  );


  LA
  g_g430_p
  (
    .dout(g430_p),
    .din1(g428_n),
    .din2(g429_n)
  );


  buf

  (
    G468_n,
    g285_p
  );


  buf

  (
    G469_n,
    g289_p
  );


  buf

  (
    G470_n,
    g293_p
  );


  buf

  (
    G471_n,
    g297_p
  );


  buf

  (
    G472_n,
    g304_p
  );


  buf

  (
    G473_n,
    g308_p
  );


  buf

  (
    G474_n,
    g312_p
  );


  buf

  (
    G475_n,
    g316_p
  );


  buf

  (
    G476_n,
    g322_p
  );


  buf

  (
    G477_n,
    g326_p
  );


  buf

  (
    G478_n,
    g330_p
  );


  buf

  (
    G479_n,
    g334_p
  );


  buf

  (
    G480_n,
    g340_p
  );


  buf

  (
    G481_n,
    g344_p
  );


  buf

  (
    G482_n,
    g348_p
  );


  buf

  (
    G483_n,
    g352_p
  );


  buf

  (
    G484_n,
    g365_p
  );


  buf

  (
    G485_n,
    g369_p
  );


  buf

  (
    G486_n,
    g373_p
  );


  buf

  (
    G487_n,
    g377_p
  );


  buf

  (
    G488_n,
    g383_p
  );


  buf

  (
    G489_n,
    g387_p
  );


  buf

  (
    G490_n,
    g391_p
  );


  buf

  (
    G491_n,
    g395_p
  );


  buf

  (
    G492_n,
    g401_p
  );


  buf

  (
    G493_n,
    g405_p
  );


  buf

  (
    G494_n,
    g409_p
  );


  buf

  (
    G495_n,
    g413_p
  );


  buf

  (
    G496_n,
    g418_p
  );


  buf

  (
    G497_n,
    g422_p
  );


  buf

  (
    G498_n,
    g426_p
  );


  buf

  (
    G499_n,
    g430_p
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G1_n_spl_0,
    G1_n_spl_
  );


  buf

  (
    G1_n_spl_00,
    G1_n_spl_0
  );


  buf

  (
    G1_n_spl_1,
    G1_n_spl_
  );


  buf

  (
    G5_n_spl_,
    G5_n
  );


  buf

  (
    G5_n_spl_0,
    G5_n_spl_
  );


  buf

  (
    G5_n_spl_00,
    G5_n_spl_0
  );


  buf

  (
    G5_n_spl_1,
    G5_n_spl_
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G1_p_spl_0,
    G1_p_spl_
  );


  buf

  (
    G1_p_spl_00,
    G1_p_spl_0
  );


  buf

  (
    G1_p_spl_1,
    G1_p_spl_
  );


  buf

  (
    G5_p_spl_,
    G5_p
  );


  buf

  (
    G5_p_spl_0,
    G5_p_spl_
  );


  buf

  (
    G5_p_spl_00,
    G5_p_spl_0
  );


  buf

  (
    G5_p_spl_1,
    G5_p_spl_
  );


  buf

  (
    G9_n_spl_,
    G9_n
  );


  buf

  (
    G9_n_spl_0,
    G9_n_spl_
  );


  buf

  (
    G9_n_spl_00,
    G9_n_spl_0
  );


  buf

  (
    G9_n_spl_1,
    G9_n_spl_
  );


  buf

  (
    G13_n_spl_,
    G13_n
  );


  buf

  (
    G13_n_spl_0,
    G13_n_spl_
  );


  buf

  (
    G13_n_spl_00,
    G13_n_spl_0
  );


  buf

  (
    G13_n_spl_1,
    G13_n_spl_
  );


  buf

  (
    G9_p_spl_,
    G9_p
  );


  buf

  (
    G9_p_spl_0,
    G9_p_spl_
  );


  buf

  (
    G9_p_spl_00,
    G9_p_spl_0
  );


  buf

  (
    G9_p_spl_1,
    G9_p_spl_
  );


  buf

  (
    G13_p_spl_,
    G13_p
  );


  buf

  (
    G13_p_spl_0,
    G13_p_spl_
  );


  buf

  (
    G13_p_spl_00,
    G13_p_spl_0
  );


  buf

  (
    G13_p_spl_1,
    G13_p_spl_
  );


  buf

  (
    g44_n_spl_,
    g44_n
  );


  buf

  (
    g47_p_spl_,
    g47_p
  );


  buf

  (
    g44_p_spl_,
    g44_p
  );


  buf

  (
    g47_n_spl_,
    g47_n
  );


  buf

  (
    G41_p_spl_,
    G41_p
  );


  buf

  (
    G41_p_spl_0,
    G41_p_spl_
  );


  buf

  (
    G41_p_spl_00,
    G41_p_spl_0
  );


  buf

  (
    G41_p_spl_01,
    G41_p_spl_0
  );


  buf

  (
    G41_p_spl_1,
    G41_p_spl_
  );


  buf

  (
    G41_p_spl_10,
    G41_p_spl_1
  );


  buf

  (
    G41_p_spl_11,
    G41_p_spl_1
  );


  buf

  (
    G41_n_spl_,
    G41_n
  );


  buf

  (
    G41_n_spl_0,
    G41_n_spl_
  );


  buf

  (
    G41_n_spl_00,
    G41_n_spl_0
  );


  buf

  (
    G41_n_spl_01,
    G41_n_spl_0
  );


  buf

  (
    G41_n_spl_1,
    G41_n_spl_
  );


  buf

  (
    G41_n_spl_10,
    G41_n_spl_1
  );


  buf

  (
    G41_n_spl_11,
    G41_n_spl_1
  );


  buf

  (
    G17_n_spl_,
    G17_n
  );


  buf

  (
    G17_n_spl_0,
    G17_n_spl_
  );


  buf

  (
    G17_n_spl_00,
    G17_n_spl_0
  );


  buf

  (
    G17_n_spl_1,
    G17_n_spl_
  );


  buf

  (
    G18_n_spl_,
    G18_n
  );


  buf

  (
    G18_n_spl_0,
    G18_n_spl_
  );


  buf

  (
    G18_n_spl_00,
    G18_n_spl_0
  );


  buf

  (
    G18_n_spl_1,
    G18_n_spl_
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


  buf

  (
    G17_p_spl_0,
    G17_p_spl_
  );


  buf

  (
    G17_p_spl_00,
    G17_p_spl_0
  );


  buf

  (
    G17_p_spl_1,
    G17_p_spl_
  );


  buf

  (
    G18_p_spl_,
    G18_p
  );


  buf

  (
    G18_p_spl_0,
    G18_p_spl_
  );


  buf

  (
    G18_p_spl_00,
    G18_p_spl_0
  );


  buf

  (
    G18_p_spl_1,
    G18_p_spl_
  );


  buf

  (
    G19_n_spl_,
    G19_n
  );


  buf

  (
    G19_n_spl_0,
    G19_n_spl_
  );


  buf

  (
    G19_n_spl_00,
    G19_n_spl_0
  );


  buf

  (
    G19_n_spl_1,
    G19_n_spl_
  );


  buf

  (
    G20_n_spl_,
    G20_n
  );


  buf

  (
    G20_n_spl_0,
    G20_n_spl_
  );


  buf

  (
    G20_n_spl_00,
    G20_n_spl_0
  );


  buf

  (
    G20_n_spl_1,
    G20_n_spl_
  );


  buf

  (
    G19_p_spl_,
    G19_p
  );


  buf

  (
    G19_p_spl_0,
    G19_p_spl_
  );


  buf

  (
    G19_p_spl_00,
    G19_p_spl_0
  );


  buf

  (
    G19_p_spl_1,
    G19_p_spl_
  );


  buf

  (
    G20_p_spl_,
    G20_p
  );


  buf

  (
    G20_p_spl_0,
    G20_p_spl_
  );


  buf

  (
    G20_p_spl_00,
    G20_p_spl_0
  );


  buf

  (
    G20_p_spl_1,
    G20_p_spl_
  );


  buf

  (
    g54_n_spl_,
    g54_n
  );


  buf

  (
    g57_p_spl_,
    g57_p
  );


  buf

  (
    g54_p_spl_,
    g54_p
  );


  buf

  (
    g57_n_spl_,
    g57_n
  );


  buf

  (
    G21_n_spl_,
    G21_n
  );


  buf

  (
    G21_n_spl_0,
    G21_n_spl_
  );


  buf

  (
    G21_n_spl_00,
    G21_n_spl_0
  );


  buf

  (
    G21_n_spl_1,
    G21_n_spl_
  );


  buf

  (
    G22_n_spl_,
    G22_n
  );


  buf

  (
    G22_n_spl_0,
    G22_n_spl_
  );


  buf

  (
    G22_n_spl_00,
    G22_n_spl_0
  );


  buf

  (
    G22_n_spl_1,
    G22_n_spl_
  );


  buf

  (
    G21_p_spl_,
    G21_p
  );


  buf

  (
    G21_p_spl_0,
    G21_p_spl_
  );


  buf

  (
    G21_p_spl_00,
    G21_p_spl_0
  );


  buf

  (
    G21_p_spl_1,
    G21_p_spl_
  );


  buf

  (
    G22_p_spl_,
    G22_p
  );


  buf

  (
    G22_p_spl_0,
    G22_p_spl_
  );


  buf

  (
    G22_p_spl_00,
    G22_p_spl_0
  );


  buf

  (
    G22_p_spl_1,
    G22_p_spl_
  );


  buf

  (
    G23_n_spl_,
    G23_n
  );


  buf

  (
    G23_n_spl_0,
    G23_n_spl_
  );


  buf

  (
    G23_n_spl_00,
    G23_n_spl_0
  );


  buf

  (
    G23_n_spl_1,
    G23_n_spl_
  );


  buf

  (
    G24_n_spl_,
    G24_n
  );


  buf

  (
    G24_n_spl_0,
    G24_n_spl_
  );


  buf

  (
    G24_n_spl_00,
    G24_n_spl_0
  );


  buf

  (
    G24_n_spl_1,
    G24_n_spl_
  );


  buf

  (
    G23_p_spl_,
    G23_p
  );


  buf

  (
    G23_p_spl_0,
    G23_p_spl_
  );


  buf

  (
    G23_p_spl_00,
    G23_p_spl_0
  );


  buf

  (
    G23_p_spl_1,
    G23_p_spl_
  );


  buf

  (
    G24_p_spl_,
    G24_p
  );


  buf

  (
    G24_p_spl_0,
    G24_p_spl_
  );


  buf

  (
    G24_p_spl_00,
    G24_p_spl_0
  );


  buf

  (
    G24_p_spl_1,
    G24_p_spl_
  );


  buf

  (
    g63_n_spl_,
    g63_n
  );


  buf

  (
    g66_p_spl_,
    g66_p
  );


  buf

  (
    g63_p_spl_,
    g63_p
  );


  buf

  (
    g66_n_spl_,
    g66_n
  );


  buf

  (
    g60_n_spl_,
    g60_n
  );


  buf

  (
    g60_n_spl_0,
    g60_n_spl_
  );


  buf

  (
    g60_n_spl_1,
    g60_n_spl_
  );


  buf

  (
    g69_n_spl_,
    g69_n
  );


  buf

  (
    g69_n_spl_0,
    g69_n_spl_
  );


  buf

  (
    g69_n_spl_1,
    g69_n_spl_
  );


  buf

  (
    g60_p_spl_,
    g60_p
  );


  buf

  (
    g60_p_spl_0,
    g60_p_spl_
  );


  buf

  (
    g60_p_spl_1,
    g60_p_spl_
  );


  buf

  (
    g69_p_spl_,
    g69_p
  );


  buf

  (
    g69_p_spl_0,
    g69_p_spl_
  );


  buf

  (
    g69_p_spl_1,
    g69_p_spl_
  );


  buf

  (
    g51_n_spl_,
    g51_n
  );


  buf

  (
    g72_p_spl_,
    g72_p
  );


  buf

  (
    g51_p_spl_,
    g51_p
  );


  buf

  (
    g72_n_spl_,
    g72_n
  );


  buf

  (
    g50_p_spl_,
    g50_p
  );


  buf

  (
    g75_n_spl_,
    g75_n
  );


  buf

  (
    g50_n_spl_,
    g50_n
  );


  buf

  (
    g75_p_spl_,
    g75_p
  );


  buf

  (
    G25_n_spl_,
    G25_n
  );


  buf

  (
    G25_n_spl_0,
    G25_n_spl_
  );


  buf

  (
    G25_n_spl_00,
    G25_n_spl_0
  );


  buf

  (
    G25_n_spl_1,
    G25_n_spl_
  );


  buf

  (
    G29_n_spl_,
    G29_n
  );


  buf

  (
    G29_n_spl_0,
    G29_n_spl_
  );


  buf

  (
    G29_n_spl_00,
    G29_n_spl_0
  );


  buf

  (
    G29_n_spl_1,
    G29_n_spl_
  );


  buf

  (
    G25_p_spl_,
    G25_p
  );


  buf

  (
    G25_p_spl_0,
    G25_p_spl_
  );


  buf

  (
    G25_p_spl_00,
    G25_p_spl_0
  );


  buf

  (
    G25_p_spl_1,
    G25_p_spl_
  );


  buf

  (
    G29_p_spl_,
    G29_p
  );


  buf

  (
    G29_p_spl_0,
    G29_p_spl_
  );


  buf

  (
    G29_p_spl_00,
    G29_p_spl_0
  );


  buf

  (
    G29_p_spl_1,
    G29_p_spl_
  );


  buf

  (
    g81_n_spl_,
    g81_n
  );


  buf

  (
    g84_p_spl_,
    g84_p
  );


  buf

  (
    g81_p_spl_,
    g81_p
  );


  buf

  (
    g84_n_spl_,
    g84_n
  );


  buf

  (
    G6_n_spl_,
    G6_n
  );


  buf

  (
    G6_n_spl_0,
    G6_n_spl_
  );


  buf

  (
    G6_n_spl_00,
    G6_n_spl_0
  );


  buf

  (
    G6_n_spl_1,
    G6_n_spl_
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G6_p_spl_0,
    G6_p_spl_
  );


  buf

  (
    G6_p_spl_00,
    G6_p_spl_0
  );


  buf

  (
    G6_p_spl_1,
    G6_p_spl_
  );


  buf

  (
    G7_n_spl_,
    G7_n
  );


  buf

  (
    G7_n_spl_0,
    G7_n_spl_
  );


  buf

  (
    G7_n_spl_00,
    G7_n_spl_0
  );


  buf

  (
    G7_n_spl_1,
    G7_n_spl_
  );


  buf

  (
    G8_n_spl_,
    G8_n
  );


  buf

  (
    G8_n_spl_0,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_00,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_1,
    G8_n_spl_
  );


  buf

  (
    G7_p_spl_,
    G7_p
  );


  buf

  (
    G7_p_spl_0,
    G7_p_spl_
  );


  buf

  (
    G7_p_spl_00,
    G7_p_spl_0
  );


  buf

  (
    G7_p_spl_1,
    G7_p_spl_
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_00,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_1,
    G8_p_spl_
  );


  buf

  (
    g91_n_spl_,
    g91_n
  );


  buf

  (
    g94_p_spl_,
    g94_p
  );


  buf

  (
    g91_p_spl_,
    g91_p
  );


  buf

  (
    g94_n_spl_,
    g94_n
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G2_n_spl_0,
    G2_n_spl_
  );


  buf

  (
    G2_n_spl_00,
    G2_n_spl_0
  );


  buf

  (
    G2_n_spl_1,
    G2_n_spl_
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G2_p_spl_0,
    G2_p_spl_
  );


  buf

  (
    G2_p_spl_00,
    G2_p_spl_0
  );


  buf

  (
    G2_p_spl_1,
    G2_p_spl_
  );


  buf

  (
    G3_n_spl_,
    G3_n
  );


  buf

  (
    G3_n_spl_0,
    G3_n_spl_
  );


  buf

  (
    G3_n_spl_00,
    G3_n_spl_0
  );


  buf

  (
    G3_n_spl_1,
    G3_n_spl_
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    G4_n_spl_0,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_00,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_1,
    G4_n_spl_
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G3_p_spl_0,
    G3_p_spl_
  );


  buf

  (
    G3_p_spl_00,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_1,
    G3_p_spl_
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_00,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    g100_n_spl_,
    g100_n
  );


  buf

  (
    g103_p_spl_,
    g103_p
  );


  buf

  (
    g100_p_spl_,
    g100_p
  );


  buf

  (
    g103_n_spl_,
    g103_n
  );


  buf

  (
    g97_n_spl_,
    g97_n
  );


  buf

  (
    g97_n_spl_0,
    g97_n_spl_
  );


  buf

  (
    g97_n_spl_1,
    g97_n_spl_
  );


  buf

  (
    g106_n_spl_,
    g106_n
  );


  buf

  (
    g106_n_spl_0,
    g106_n_spl_
  );


  buf

  (
    g106_n_spl_1,
    g106_n_spl_
  );


  buf

  (
    g97_p_spl_,
    g97_p
  );


  buf

  (
    g97_p_spl_0,
    g97_p_spl_
  );


  buf

  (
    g97_p_spl_1,
    g97_p_spl_
  );


  buf

  (
    g106_p_spl_,
    g106_p
  );


  buf

  (
    g106_p_spl_0,
    g106_p_spl_
  );


  buf

  (
    g106_p_spl_1,
    g106_p_spl_
  );


  buf

  (
    g88_n_spl_,
    g88_n
  );


  buf

  (
    g109_p_spl_,
    g109_p
  );


  buf

  (
    g88_p_spl_,
    g88_p
  );


  buf

  (
    g109_n_spl_,
    g109_n
  );


  buf

  (
    g87_p_spl_,
    g87_p
  );


  buf

  (
    g112_n_spl_,
    g112_n
  );


  buf

  (
    g87_n_spl_,
    g87_n
  );


  buf

  (
    g112_p_spl_,
    g112_p
  );


  buf

  (
    G26_n_spl_,
    G26_n
  );


  buf

  (
    G26_n_spl_0,
    G26_n_spl_
  );


  buf

  (
    G26_n_spl_00,
    G26_n_spl_0
  );


  buf

  (
    G26_n_spl_1,
    G26_n_spl_
  );


  buf

  (
    G30_n_spl_,
    G30_n
  );


  buf

  (
    G30_n_spl_0,
    G30_n_spl_
  );


  buf

  (
    G30_n_spl_00,
    G30_n_spl_0
  );


  buf

  (
    G30_n_spl_1,
    G30_n_spl_
  );


  buf

  (
    G26_p_spl_,
    G26_p
  );


  buf

  (
    G26_p_spl_0,
    G26_p_spl_
  );


  buf

  (
    G26_p_spl_00,
    G26_p_spl_0
  );


  buf

  (
    G26_p_spl_1,
    G26_p_spl_
  );


  buf

  (
    G30_p_spl_,
    G30_p
  );


  buf

  (
    G30_p_spl_0,
    G30_p_spl_
  );


  buf

  (
    G30_p_spl_00,
    G30_p_spl_0
  );


  buf

  (
    G30_p_spl_1,
    G30_p_spl_
  );


  buf

  (
    g118_n_spl_,
    g118_n
  );


  buf

  (
    g121_p_spl_,
    g121_p
  );


  buf

  (
    g118_p_spl_,
    g118_p
  );


  buf

  (
    g121_n_spl_,
    g121_n
  );


  buf

  (
    G14_n_spl_,
    G14_n
  );


  buf

  (
    G14_n_spl_0,
    G14_n_spl_
  );


  buf

  (
    G14_n_spl_00,
    G14_n_spl_0
  );


  buf

  (
    G14_n_spl_1,
    G14_n_spl_
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G14_p_spl_0,
    G14_p_spl_
  );


  buf

  (
    G14_p_spl_00,
    G14_p_spl_0
  );


  buf

  (
    G14_p_spl_1,
    G14_p_spl_
  );


  buf

  (
    G15_n_spl_,
    G15_n
  );


  buf

  (
    G15_n_spl_0,
    G15_n_spl_
  );


  buf

  (
    G15_n_spl_00,
    G15_n_spl_0
  );


  buf

  (
    G15_n_spl_1,
    G15_n_spl_
  );


  buf

  (
    G16_n_spl_,
    G16_n
  );


  buf

  (
    G16_n_spl_0,
    G16_n_spl_
  );


  buf

  (
    G16_n_spl_00,
    G16_n_spl_0
  );


  buf

  (
    G16_n_spl_1,
    G16_n_spl_
  );


  buf

  (
    G15_p_spl_,
    G15_p
  );


  buf

  (
    G15_p_spl_0,
    G15_p_spl_
  );


  buf

  (
    G15_p_spl_00,
    G15_p_spl_0
  );


  buf

  (
    G15_p_spl_1,
    G15_p_spl_
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    G16_p_spl_0,
    G16_p_spl_
  );


  buf

  (
    G16_p_spl_00,
    G16_p_spl_0
  );


  buf

  (
    G16_p_spl_1,
    G16_p_spl_
  );


  buf

  (
    g128_n_spl_,
    g128_n
  );


  buf

  (
    g131_p_spl_,
    g131_p
  );


  buf

  (
    g128_p_spl_,
    g128_p
  );


  buf

  (
    g131_n_spl_,
    g131_n
  );


  buf

  (
    G10_n_spl_,
    G10_n
  );


  buf

  (
    G10_n_spl_0,
    G10_n_spl_
  );


  buf

  (
    G10_n_spl_00,
    G10_n_spl_0
  );


  buf

  (
    G10_n_spl_1,
    G10_n_spl_
  );


  buf

  (
    G10_p_spl_,
    G10_p
  );


  buf

  (
    G10_p_spl_0,
    G10_p_spl_
  );


  buf

  (
    G10_p_spl_00,
    G10_p_spl_0
  );


  buf

  (
    G10_p_spl_1,
    G10_p_spl_
  );


  buf

  (
    G11_n_spl_,
    G11_n
  );


  buf

  (
    G11_n_spl_0,
    G11_n_spl_
  );


  buf

  (
    G11_n_spl_00,
    G11_n_spl_0
  );


  buf

  (
    G11_n_spl_1,
    G11_n_spl_
  );


  buf

  (
    G12_n_spl_,
    G12_n
  );


  buf

  (
    G12_n_spl_0,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_00,
    G12_n_spl_0
  );


  buf

  (
    G12_n_spl_1,
    G12_n_spl_
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    G11_p_spl_0,
    G11_p_spl_
  );


  buf

  (
    G11_p_spl_00,
    G11_p_spl_0
  );


  buf

  (
    G11_p_spl_1,
    G11_p_spl_
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G12_p_spl_0,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_00,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_1,
    G12_p_spl_
  );


  buf

  (
    g137_n_spl_,
    g137_n
  );


  buf

  (
    g140_p_spl_,
    g140_p
  );


  buf

  (
    g137_p_spl_,
    g137_p
  );


  buf

  (
    g140_n_spl_,
    g140_n
  );


  buf

  (
    g134_n_spl_,
    g134_n
  );


  buf

  (
    g134_n_spl_0,
    g134_n_spl_
  );


  buf

  (
    g134_n_spl_1,
    g134_n_spl_
  );


  buf

  (
    g143_n_spl_,
    g143_n
  );


  buf

  (
    g143_n_spl_0,
    g143_n_spl_
  );


  buf

  (
    g143_n_spl_1,
    g143_n_spl_
  );


  buf

  (
    g134_p_spl_,
    g134_p
  );


  buf

  (
    g134_p_spl_0,
    g134_p_spl_
  );


  buf

  (
    g134_p_spl_1,
    g134_p_spl_
  );


  buf

  (
    g143_p_spl_,
    g143_p
  );


  buf

  (
    g143_p_spl_0,
    g143_p_spl_
  );


  buf

  (
    g143_p_spl_1,
    g143_p_spl_
  );


  buf

  (
    g125_n_spl_,
    g125_n
  );


  buf

  (
    g146_p_spl_,
    g146_p
  );


  buf

  (
    g125_p_spl_,
    g125_p
  );


  buf

  (
    g146_n_spl_,
    g146_n
  );


  buf

  (
    g124_p_spl_,
    g124_p
  );


  buf

  (
    g149_n_spl_,
    g149_n
  );


  buf

  (
    g124_n_spl_,
    g124_n
  );


  buf

  (
    g149_p_spl_,
    g149_p
  );


  buf

  (
    g115_n_spl_,
    g115_n
  );


  buf

  (
    g115_n_spl_0,
    g115_n_spl_
  );


  buf

  (
    g115_n_spl_00,
    g115_n_spl_0
  );


  buf

  (
    g115_n_spl_01,
    g115_n_spl_0
  );


  buf

  (
    g115_n_spl_1,
    g115_n_spl_
  );


  buf

  (
    g115_n_spl_10,
    g115_n_spl_1
  );


  buf

  (
    g152_p_spl_,
    g152_p
  );


  buf

  (
    g152_p_spl_0,
    g152_p_spl_
  );


  buf

  (
    g152_p_spl_00,
    g152_p_spl_0
  );


  buf

  (
    g152_p_spl_01,
    g152_p_spl_0
  );


  buf

  (
    g152_p_spl_1,
    g152_p_spl_
  );


  buf

  (
    g152_p_spl_10,
    g152_p_spl_1
  );


  buf

  (
    g115_p_spl_,
    g115_p
  );


  buf

  (
    g115_p_spl_0,
    g115_p_spl_
  );


  buf

  (
    g115_p_spl_00,
    g115_p_spl_0
  );


  buf

  (
    g115_p_spl_01,
    g115_p_spl_0
  );


  buf

  (
    g115_p_spl_1,
    g115_p_spl_
  );


  buf

  (
    g115_p_spl_10,
    g115_p_spl_1
  );


  buf

  (
    g152_n_spl_,
    g152_n
  );


  buf

  (
    g152_n_spl_0,
    g152_n_spl_
  );


  buf

  (
    g152_n_spl_00,
    g152_n_spl_0
  );


  buf

  (
    g152_n_spl_01,
    g152_n_spl_0
  );


  buf

  (
    g152_n_spl_1,
    g152_n_spl_
  );


  buf

  (
    g152_n_spl_10,
    g152_n_spl_1
  );


  buf

  (
    G28_n_spl_,
    G28_n
  );


  buf

  (
    G28_n_spl_0,
    G28_n_spl_
  );


  buf

  (
    G28_n_spl_00,
    G28_n_spl_0
  );


  buf

  (
    G28_n_spl_1,
    G28_n_spl_
  );


  buf

  (
    G32_n_spl_,
    G32_n
  );


  buf

  (
    G32_n_spl_0,
    G32_n_spl_
  );


  buf

  (
    G32_n_spl_00,
    G32_n_spl_0
  );


  buf

  (
    G32_n_spl_1,
    G32_n_spl_
  );


  buf

  (
    G28_p_spl_,
    G28_p
  );


  buf

  (
    G28_p_spl_0,
    G28_p_spl_
  );


  buf

  (
    G28_p_spl_00,
    G28_p_spl_0
  );


  buf

  (
    G28_p_spl_1,
    G28_p_spl_
  );


  buf

  (
    G32_p_spl_,
    G32_p
  );


  buf

  (
    G32_p_spl_0,
    G32_p_spl_
  );


  buf

  (
    G32_p_spl_00,
    G32_p_spl_0
  );


  buf

  (
    G32_p_spl_1,
    G32_p_spl_
  );


  buf

  (
    g156_n_spl_,
    g156_n
  );


  buf

  (
    g159_p_spl_,
    g159_p
  );


  buf

  (
    g156_p_spl_,
    g156_p
  );


  buf

  (
    g159_n_spl_,
    g159_n
  );


  buf

  (
    g163_n_spl_,
    g163_n
  );


  buf

  (
    g166_p_spl_,
    g166_p
  );


  buf

  (
    g163_p_spl_,
    g163_p
  );


  buf

  (
    g166_n_spl_,
    g166_n
  );


  buf

  (
    g162_p_spl_,
    g162_p
  );


  buf

  (
    g169_n_spl_,
    g169_n
  );


  buf

  (
    g162_n_spl_,
    g162_n
  );


  buf

  (
    g169_p_spl_,
    g169_p
  );


  buf

  (
    G27_n_spl_,
    G27_n
  );


  buf

  (
    G27_n_spl_0,
    G27_n_spl_
  );


  buf

  (
    G27_n_spl_00,
    G27_n_spl_0
  );


  buf

  (
    G27_n_spl_1,
    G27_n_spl_
  );


  buf

  (
    G31_n_spl_,
    G31_n
  );


  buf

  (
    G31_n_spl_0,
    G31_n_spl_
  );


  buf

  (
    G31_n_spl_00,
    G31_n_spl_0
  );


  buf

  (
    G31_n_spl_1,
    G31_n_spl_
  );


  buf

  (
    G27_p_spl_,
    G27_p
  );


  buf

  (
    G27_p_spl_0,
    G27_p_spl_
  );


  buf

  (
    G27_p_spl_00,
    G27_p_spl_0
  );


  buf

  (
    G27_p_spl_1,
    G27_p_spl_
  );


  buf

  (
    G31_p_spl_,
    G31_p
  );


  buf

  (
    G31_p_spl_0,
    G31_p_spl_
  );


  buf

  (
    G31_p_spl_00,
    G31_p_spl_0
  );


  buf

  (
    G31_p_spl_1,
    G31_p_spl_
  );


  buf

  (
    g175_n_spl_,
    g175_n
  );


  buf

  (
    g178_p_spl_,
    g178_p
  );


  buf

  (
    g175_p_spl_,
    g175_p
  );


  buf

  (
    g178_n_spl_,
    g178_n
  );


  buf

  (
    g182_n_spl_,
    g182_n
  );


  buf

  (
    g185_p_spl_,
    g185_p
  );


  buf

  (
    g182_p_spl_,
    g182_p
  );


  buf

  (
    g185_n_spl_,
    g185_n
  );


  buf

  (
    g181_p_spl_,
    g181_p
  );


  buf

  (
    g188_n_spl_,
    g188_n
  );


  buf

  (
    g181_n_spl_,
    g181_n
  );


  buf

  (
    g188_p_spl_,
    g188_p
  );


  buf

  (
    g172_p_spl_,
    g172_p
  );


  buf

  (
    g172_p_spl_0,
    g172_p_spl_
  );


  buf

  (
    g172_p_spl_00,
    g172_p_spl_0
  );


  buf

  (
    g172_p_spl_01,
    g172_p_spl_0
  );


  buf

  (
    g172_p_spl_1,
    g172_p_spl_
  );


  buf

  (
    g172_p_spl_10,
    g172_p_spl_1
  );


  buf

  (
    g172_p_spl_11,
    g172_p_spl_1
  );


  buf

  (
    g191_n_spl_,
    g191_n
  );


  buf

  (
    g191_n_spl_0,
    g191_n_spl_
  );


  buf

  (
    g191_n_spl_00,
    g191_n_spl_0
  );


  buf

  (
    g191_n_spl_01,
    g191_n_spl_0
  );


  buf

  (
    g191_n_spl_1,
    g191_n_spl_
  );


  buf

  (
    g191_n_spl_10,
    g191_n_spl_1
  );


  buf

  (
    g191_n_spl_11,
    g191_n_spl_1
  );


  buf

  (
    g172_n_spl_,
    g172_n
  );


  buf

  (
    g172_n_spl_0,
    g172_n_spl_
  );


  buf

  (
    g172_n_spl_00,
    g172_n_spl_0
  );


  buf

  (
    g172_n_spl_01,
    g172_n_spl_0
  );


  buf

  (
    g172_n_spl_1,
    g172_n_spl_
  );


  buf

  (
    g172_n_spl_10,
    g172_n_spl_1
  );


  buf

  (
    g172_n_spl_11,
    g172_n_spl_1
  );


  buf

  (
    g191_p_spl_,
    g191_p
  );


  buf

  (
    g191_p_spl_0,
    g191_p_spl_
  );


  buf

  (
    g191_p_spl_00,
    g191_p_spl_0
  );


  buf

  (
    g191_p_spl_01,
    g191_p_spl_0
  );


  buf

  (
    g191_p_spl_1,
    g191_p_spl_
  );


  buf

  (
    g191_p_spl_10,
    g191_p_spl_1
  );


  buf

  (
    g191_p_spl_11,
    g191_p_spl_1
  );


  buf

  (
    g195_n_spl_,
    g195_n
  );


  buf

  (
    g198_p_spl_,
    g198_p
  );


  buf

  (
    g195_p_spl_,
    g195_p
  );


  buf

  (
    g198_n_spl_,
    g198_n
  );


  buf

  (
    g205_n_spl_,
    g205_n
  );


  buf

  (
    g208_p_spl_,
    g208_p
  );


  buf

  (
    g205_p_spl_,
    g205_p
  );


  buf

  (
    g208_n_spl_,
    g208_n
  );


  buf

  (
    g211_n_spl_,
    g211_n
  );


  buf

  (
    g211_n_spl_0,
    g211_n_spl_
  );


  buf

  (
    g211_n_spl_1,
    g211_n_spl_
  );


  buf

  (
    g211_p_spl_,
    g211_p
  );


  buf

  (
    g211_p_spl_0,
    g211_p_spl_
  );


  buf

  (
    g211_p_spl_1,
    g211_p_spl_
  );


  buf

  (
    g202_n_spl_,
    g202_n
  );


  buf

  (
    g214_p_spl_,
    g214_p
  );


  buf

  (
    g202_p_spl_,
    g202_p
  );


  buf

  (
    g214_n_spl_,
    g214_n
  );


  buf

  (
    g201_p_spl_,
    g201_p
  );


  buf

  (
    g217_n_spl_,
    g217_n
  );


  buf

  (
    g201_n_spl_,
    g201_n
  );


  buf

  (
    g217_p_spl_,
    g217_p
  );


  buf

  (
    g223_n_spl_,
    g223_n
  );


  buf

  (
    g226_p_spl_,
    g226_p
  );


  buf

  (
    g223_p_spl_,
    g223_p
  );


  buf

  (
    g226_n_spl_,
    g226_n
  );


  buf

  (
    g233_n_spl_,
    g233_n
  );


  buf

  (
    g236_p_spl_,
    g236_p
  );


  buf

  (
    g233_p_spl_,
    g233_p
  );


  buf

  (
    g236_n_spl_,
    g236_n
  );


  buf

  (
    g239_n_spl_,
    g239_n
  );


  buf

  (
    g239_n_spl_0,
    g239_n_spl_
  );


  buf

  (
    g239_n_spl_1,
    g239_n_spl_
  );


  buf

  (
    g239_p_spl_,
    g239_p
  );


  buf

  (
    g239_p_spl_0,
    g239_p_spl_
  );


  buf

  (
    g239_p_spl_1,
    g239_p_spl_
  );


  buf

  (
    g230_n_spl_,
    g230_n
  );


  buf

  (
    g242_p_spl_,
    g242_p
  );


  buf

  (
    g230_p_spl_,
    g230_p
  );


  buf

  (
    g242_n_spl_,
    g242_n
  );


  buf

  (
    g229_p_spl_,
    g229_p
  );


  buf

  (
    g245_n_spl_,
    g245_n
  );


  buf

  (
    g229_n_spl_,
    g229_n
  );


  buf

  (
    g245_p_spl_,
    g245_p
  );


  buf

  (
    g251_n_spl_,
    g251_n
  );


  buf

  (
    g254_p_spl_,
    g254_p
  );


  buf

  (
    g251_p_spl_,
    g251_p
  );


  buf

  (
    g254_n_spl_,
    g254_n
  );


  buf

  (
    g258_n_spl_,
    g258_n
  );


  buf

  (
    g261_p_spl_,
    g261_p
  );


  buf

  (
    g258_p_spl_,
    g258_p
  );


  buf

  (
    g261_n_spl_,
    g261_n
  );


  buf

  (
    g257_p_spl_,
    g257_p
  );


  buf

  (
    g264_n_spl_,
    g264_n
  );


  buf

  (
    g257_n_spl_,
    g257_n
  );


  buf

  (
    g264_p_spl_,
    g264_p
  );


  buf

  (
    g78_n_spl_,
    g78_n
  );


  buf

  (
    g78_n_spl_0,
    g78_n_spl_
  );


  buf

  (
    g78_n_spl_00,
    g78_n_spl_0
  );


  buf

  (
    g78_n_spl_01,
    g78_n_spl_0
  );


  buf

  (
    g78_n_spl_1,
    g78_n_spl_
  );


  buf

  (
    g78_n_spl_10,
    g78_n_spl_1
  );


  buf

  (
    g267_p_spl_,
    g267_p
  );


  buf

  (
    g267_p_spl_0,
    g267_p_spl_
  );


  buf

  (
    g267_p_spl_00,
    g267_p_spl_0
  );


  buf

  (
    g267_p_spl_01,
    g267_p_spl_0
  );


  buf

  (
    g267_p_spl_1,
    g267_p_spl_
  );


  buf

  (
    g267_p_spl_10,
    g267_p_spl_1
  );


  buf

  (
    g78_p_spl_,
    g78_p
  );


  buf

  (
    g78_p_spl_0,
    g78_p_spl_
  );


  buf

  (
    g78_p_spl_00,
    g78_p_spl_0
  );


  buf

  (
    g78_p_spl_01,
    g78_p_spl_0
  );


  buf

  (
    g78_p_spl_1,
    g78_p_spl_
  );


  buf

  (
    g78_p_spl_10,
    g78_p_spl_1
  );


  buf

  (
    g267_n_spl_,
    g267_n
  );


  buf

  (
    g267_n_spl_0,
    g267_n_spl_
  );


  buf

  (
    g267_n_spl_00,
    g267_n_spl_0
  );


  buf

  (
    g267_n_spl_01,
    g267_n_spl_0
  );


  buf

  (
    g267_n_spl_1,
    g267_n_spl_
  );


  buf

  (
    g267_n_spl_10,
    g267_n_spl_1
  );


  buf

  (
    g248_p_spl_,
    g248_p
  );


  buf

  (
    g248_p_spl_0,
    g248_p_spl_
  );


  buf

  (
    g248_p_spl_00,
    g248_p_spl_0
  );


  buf

  (
    g248_p_spl_01,
    g248_p_spl_0
  );


  buf

  (
    g248_p_spl_1,
    g248_p_spl_
  );


  buf

  (
    g248_p_spl_10,
    g248_p_spl_1
  );


  buf

  (
    g248_p_spl_11,
    g248_p_spl_1
  );


  buf

  (
    g268_p_spl_,
    g268_p
  );


  buf

  (
    g248_n_spl_,
    g248_n
  );


  buf

  (
    g248_n_spl_0,
    g248_n_spl_
  );


  buf

  (
    g248_n_spl_00,
    g248_n_spl_0
  );


  buf

  (
    g248_n_spl_01,
    g248_n_spl_0
  );


  buf

  (
    g248_n_spl_1,
    g248_n_spl_
  );


  buf

  (
    g248_n_spl_10,
    g248_n_spl_1
  );


  buf

  (
    g248_n_spl_11,
    g248_n_spl_1
  );


  buf

  (
    g268_n_spl_,
    g268_n
  );


  buf

  (
    g270_p_spl_,
    g270_p
  );


  buf

  (
    g270_n_spl_,
    g270_n
  );


  buf

  (
    g269_n_spl_,
    g269_n
  );


  buf

  (
    g271_n_spl_,
    g271_n
  );


  buf

  (
    g269_p_spl_,
    g269_p
  );


  buf

  (
    g271_p_spl_,
    g271_p
  );


  buf

  (
    g220_p_spl_,
    g220_p
  );


  buf

  (
    g220_p_spl_0,
    g220_p_spl_
  );


  buf

  (
    g220_p_spl_00,
    g220_p_spl_0
  );


  buf

  (
    g220_p_spl_01,
    g220_p_spl_0
  );


  buf

  (
    g220_p_spl_1,
    g220_p_spl_
  );


  buf

  (
    g220_p_spl_10,
    g220_p_spl_1
  );


  buf

  (
    g220_p_spl_11,
    g220_p_spl_1
  );


  buf

  (
    g220_n_spl_,
    g220_n
  );


  buf

  (
    g220_n_spl_0,
    g220_n_spl_
  );


  buf

  (
    g220_n_spl_00,
    g220_n_spl_0
  );


  buf

  (
    g220_n_spl_01,
    g220_n_spl_0
  );


  buf

  (
    g220_n_spl_1,
    g220_n_spl_
  );


  buf

  (
    g220_n_spl_10,
    g220_n_spl_1
  );


  buf

  (
    g220_n_spl_11,
    g220_n_spl_1
  );


  buf

  (
    g274_n_spl_,
    g274_n
  );


  buf

  (
    g274_n_spl_0,
    g274_n_spl_
  );


  buf

  (
    g274_p_spl_,
    g274_p
  );


  buf

  (
    g274_p_spl_0,
    g274_p_spl_
  );


  buf

  (
    g192_p_spl_,
    g192_p
  );


  buf

  (
    g279_n_spl_,
    g279_n
  );


  buf

  (
    g192_n_spl_,
    g192_n
  );


  buf

  (
    g279_p_spl_,
    g279_p
  );


  buf

  (
    g153_p_spl_,
    g153_p
  );


  buf

  (
    g280_p_spl_,
    g280_p
  );


  buf

  (
    g153_n_spl_,
    g153_n
  );


  buf

  (
    g280_n_spl_,
    g280_n
  );


  buf

  (
    g281_p_spl_,
    g281_p
  );


  buf

  (
    g281_p_spl_0,
    g281_p_spl_
  );


  buf

  (
    g281_p_spl_1,
    g281_p_spl_
  );


  buf

  (
    g281_n_spl_,
    g281_n
  );


  buf

  (
    g281_n_spl_0,
    g281_n_spl_
  );


  buf

  (
    g281_n_spl_1,
    g281_n_spl_
  );


  buf

  (
    g298_p_spl_,
    g298_p
  );


  buf

  (
    g299_p_spl_,
    g299_p
  );


  buf

  (
    g298_n_spl_,
    g298_n
  );


  buf

  (
    g299_n_spl_,
    g299_n
  );


  buf

  (
    g300_p_spl_,
    g300_p
  );


  buf

  (
    g300_p_spl_0,
    g300_p_spl_
  );


  buf

  (
    g300_p_spl_1,
    g300_p_spl_
  );


  buf

  (
    g300_n_spl_,
    g300_n
  );


  buf

  (
    g300_n_spl_0,
    g300_n_spl_
  );


  buf

  (
    g300_n_spl_1,
    g300_n_spl_
  );


  buf

  (
    g317_p_spl_,
    g317_p
  );


  buf

  (
    g317_n_spl_,
    g317_n
  );


  buf

  (
    g318_p_spl_,
    g318_p
  );


  buf

  (
    g318_p_spl_0,
    g318_p_spl_
  );


  buf

  (
    g318_p_spl_1,
    g318_p_spl_
  );


  buf

  (
    g318_n_spl_,
    g318_n
  );


  buf

  (
    g318_n_spl_0,
    g318_n_spl_
  );


  buf

  (
    g318_n_spl_1,
    g318_n_spl_
  );


  buf

  (
    g335_p_spl_,
    g335_p
  );


  buf

  (
    g335_n_spl_,
    g335_n
  );


  buf

  (
    g336_p_spl_,
    g336_p
  );


  buf

  (
    g336_p_spl_0,
    g336_p_spl_
  );


  buf

  (
    g336_p_spl_1,
    g336_p_spl_
  );


  buf

  (
    g336_n_spl_,
    g336_n
  );


  buf

  (
    g336_n_spl_0,
    g336_n_spl_
  );


  buf

  (
    g336_n_spl_1,
    g336_n_spl_
  );


  buf

  (
    g359_n_spl_,
    g359_n
  );


  buf

  (
    g359_n_spl_0,
    g359_n_spl_
  );


  buf

  (
    g359_p_spl_,
    g359_p
  );


  buf

  (
    g359_p_spl_0,
    g359_p_spl_
  );


  buf

  (
    g361_p_spl_,
    g361_p
  );


  buf

  (
    g361_p_spl_0,
    g361_p_spl_
  );


  buf

  (
    g361_p_spl_1,
    g361_p_spl_
  );


  buf

  (
    g361_n_spl_,
    g361_n
  );


  buf

  (
    g361_n_spl_0,
    g361_n_spl_
  );


  buf

  (
    g361_n_spl_1,
    g361_n_spl_
  );


  buf

  (
    g378_p_spl_,
    g378_p
  );


  buf

  (
    g378_n_spl_,
    g378_n
  );


  buf

  (
    g379_p_spl_,
    g379_p
  );


  buf

  (
    g379_p_spl_0,
    g379_p_spl_
  );


  buf

  (
    g379_p_spl_1,
    g379_p_spl_
  );


  buf

  (
    g379_n_spl_,
    g379_n
  );


  buf

  (
    g379_n_spl_0,
    g379_n_spl_
  );


  buf

  (
    g379_n_spl_1,
    g379_n_spl_
  );


  buf

  (
    g397_p_spl_,
    g397_p
  );


  buf

  (
    g397_p_spl_0,
    g397_p_spl_
  );


  buf

  (
    g397_p_spl_1,
    g397_p_spl_
  );


  buf

  (
    g397_n_spl_,
    g397_n
  );


  buf

  (
    g397_n_spl_0,
    g397_n_spl_
  );


  buf

  (
    g397_n_spl_1,
    g397_n_spl_
  );


  buf

  (
    g414_p_spl_,
    g414_p
  );


  buf

  (
    g414_p_spl_0,
    g414_p_spl_
  );


  buf

  (
    g414_p_spl_1,
    g414_p_spl_
  );


  buf

  (
    g414_n_spl_,
    g414_n
  );


  buf

  (
    g414_n_spl_0,
    g414_n_spl_
  );


  buf

  (
    g414_n_spl_1,
    g414_n_spl_
  );


endmodule
