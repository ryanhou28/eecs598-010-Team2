// Benchmark "mymod" written by ABC on Sun Oct 29 19:31:47 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36,
    G426, G427, G428, G429, G430, G431, G432  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36;
  output G426, G427, G428, G429, G430, G431, G432;
  reg n205_lo, n214_lo, n217_lo, n226_lo, n229_lo, n232_lo, n238_lo,
    n241_lo, n250_lo, n253_lo, n256_lo, n262_lo, n265_lo, n274_lo, n277_lo,
    n280_lo, n286_lo, n289_lo, n298_lo, n301_lo, n304_lo, n310_lo, n313_lo,
    n322_lo, n325_lo, n328_lo, n334_lo, n337_lo, n346_lo, n349_lo, n352_lo,
    n358_lo, n361_lo, n370_lo, n373_lo, n376_lo, n382_lo, n385_lo, n394_lo,
    n397_lo, n400_lo, n406_lo, n409_lo, n418_lo, n421_lo, n424_lo, n430_lo,
    n433_lo, n442_lo, n445_lo, n448_lo, n454_lo, n457_lo, n466_lo, n469_lo,
    n472_lo, n478_lo, n481_lo, n490_lo, n493_lo, n496_lo, n502_lo, n505_lo,
    n514_lo, n517_lo, n520_lo, n526_lo, n529_lo, n538_lo, n541_lo, n544_lo,
    n550_lo, n553_lo, n562_lo, n565_lo, n568_lo, n574_lo, n577_lo, n586_lo,
    n589_lo, n592_lo, n598_lo, n601_lo, n610_lo, n613_lo, n616_lo, n622_lo,
    n625_lo, n628_lo, n634_lo, n316_inv, n319_inv, n997_o2, n998_o2,
    n999_o2, n1000_o2, n1001_o2, n1002_o2, n1003_o2, n1004_o2, n1005_o2,
    n1015_o2, n1016_o2, n1017_o2, n1018_o2, n1019_o2, n1020_o2, n1021_o2,
    n1022_o2, n1023_o2, n376_1_inv, n235_lo_buf_o2, n283_lo_buf_o2,
    n331_lo_buf_o2, n379_lo_buf_o2, n427_lo_buf_o2, n475_lo_buf_o2,
    n523_lo_buf_o2, n571_lo_buf_o2, n619_lo_buf_o2, n406_1_inv, G223_o2,
    G226_o2, G229_o2, G232_o2, G235_o2, G238_o2, G242_o2, G246_o2, G250_o2,
    n259_lo_buf_o2, n307_lo_buf_o2, n355_lo_buf_o2, n403_lo_buf_o2,
    n451_lo_buf_o2, n499_lo_buf_o2, n547_lo_buf_o2, n595_lo_buf_o2,
    n631_lo_buf_o2, G213_o2, G318_o2, G358_o2, G259_o2, G263_o2, G266_o2,
    G269_o2, G272_o2, G275_o2, G278_o2, G281_o2, G284_o2, n211_lo_buf_o2,
    n247_lo_buf_o2, n295_lo_buf_o2, n343_lo_buf_o2, n391_lo_buf_o2,
    n439_lo_buf_o2, n487_lo_buf_o2, n535_lo_buf_o2, n583_lo_buf_o2,
    G158_o2, G184_o2, G186_o2, G188_o2, G190_o2, G192_o2, G194_o2, G196_o2,
    G198_o2, n223_lo_buf_o2, n271_lo_buf_o2, n319_lo_buf_o2,
    n367_lo_buf_o2, n415_lo_buf_o2, n463_lo_buf_o2, n511_lo_buf_o2,
    n559_lo_buf_o2, n607_lo_buf_o2, n580_inv, G154_o2, G159_o2, G162_o2,
    G165_o2, G168_o2, G171_o2, G174_o2, G177_o2, G180_o2;
  wire new_new_n420__, new_new_n422__, new_new_n424__, new_new_n426__,
    new_new_n428__, new_new_n430__, new_new_n432__, new_new_n434__,
    new_new_n436__, new_new_n438__, new_new_n440__, new_new_n442__,
    new_new_n444__, new_new_n446__, new_new_n448__, new_new_n450__,
    new_new_n452__, new_new_n454__, new_new_n456__, new_new_n458__,
    new_new_n460__, new_new_n462__, new_new_n464__, new_new_n466__,
    new_new_n468__, new_new_n470__, new_new_n472__, new_new_n474__,
    new_new_n476__, new_new_n478__, new_new_n480__, new_new_n482__,
    new_new_n484__, new_new_n486__, new_new_n488__, new_new_n490__,
    new_new_n492__, new_new_n493__, new_new_n495__, new_new_n496__,
    new_new_n498__, new_new_n500__, new_new_n502__, new_new_n503__,
    new_new_n505__, new_new_n506__, new_new_n507__, new_new_n508__,
    new_new_n510__, new_new_n512__, new_new_n513__, new_new_n515__,
    new_new_n516__, new_new_n519__, new_new_n520__, new_new_n522__,
    new_new_n523__, new_new_n524__, new_new_n526__, new_new_n527__,
    new_new_n528__, new_new_n529__, new_new_n530__, new_new_n532__,
    new_new_n533__, new_new_n534__, new_new_n536__, new_new_n538__,
    new_new_n539__, new_new_n540__, new_new_n542__, new_new_n543__,
    new_new_n544__, new_new_n545__, new_new_n546__, new_new_n547__,
    new_new_n548__, new_new_n549__, new_new_n550__, new_new_n552__,
    new_new_n553__, new_new_n554__, new_new_n555__, new_new_n556__,
    new_new_n558__, new_new_n559__, new_new_n560__, new_new_n562__,
    new_new_n563__, new_new_n564__, new_new_n565__, new_new_n566__,
    new_new_n567__, new_new_n568__, new_new_n569__, new_new_n570__,
    new_new_n572__, new_new_n573__, new_new_n574__, new_new_n575__,
    new_new_n576__, new_new_n578__, new_new_n579__, new_new_n580__,
    new_new_n582__, new_new_n583__, new_new_n584__, new_new_n585__,
    new_new_n586__, new_new_n587__, new_new_n588__, new_new_n590__,
    new_new_n592__, new_new_n593__, new_new_n594__, new_new_n595__,
    new_new_n596__, new_new_n599__, new_new_n600__, new_new_n602__,
    new_new_n603__, new_new_n604__, new_new_n606__, new_new_n607__,
    new_new_n608__, new_new_n609__, new_new_n610__, new_new_n612__,
    new_new_n613__, new_new_n614__, new_new_n616__, new_new_n618__,
    new_new_n619__, new_new_n620__, new_new_n622__, new_new_n623__,
    new_new_n624__, new_new_n625__, new_new_n626__, new_new_n627__,
    new_new_n628__, new_new_n630__, new_new_n632__, new_new_n633__,
    new_new_n634__, new_new_n635__, new_new_n636__, new_new_n639__,
    new_new_n640__, new_new_n642__, new_new_n643__, new_new_n644__,
    new_new_n646__, new_new_n647__, new_new_n648__, new_new_n650__,
    new_new_n652__, new_new_n653__, new_new_n654__, new_new_n656__,
    new_new_n659__, new_new_n660__, new_new_n662__, new_new_n663__,
    new_new_n664__, new_new_n666__, new_new_n668__, new_new_n669__,
    new_new_n670__, new_new_n672__, new_new_n674__, new_new_n676__,
    new_new_n678__, new_new_n680__, new_new_n682__, new_new_n684__,
    new_new_n686__, new_new_n688__, new_new_n690__, new_new_n692__,
    new_new_n694__, new_new_n696__, new_new_n698__, new_new_n700__,
    new_new_n702__, new_new_n704__, new_new_n706__, new_new_n708__,
    new_new_n710__, new_new_n712__, new_new_n714__, new_new_n716__,
    new_new_n718__, new_new_n720__, new_new_n722__, new_new_n724__,
    new_new_n726__, new_new_n728__, new_new_n730__, new_new_n732__,
    new_new_n735__, new_new_n737__, new_new_n739__, new_new_n741__,
    new_new_n743__, new_new_n745__, new_new_n747__, new_new_n749__,
    new_new_n751__, new_new_n752__, new_new_n754__, new_new_n756__,
    new_new_n758__, new_new_n760__, new_new_n762__, new_new_n764__,
    new_new_n766__, new_new_n768__, new_new_n770__, new_new_n771__,
    new_new_n772__, new_new_n773__, new_new_n774__, new_new_n775__,
    new_new_n776__, new_new_n777__, new_new_n778__, new_new_n779__,
    new_new_n780__, new_new_n781__, new_new_n782__, new_new_n783__,
    new_new_n784__, new_new_n785__, new_new_n786__, new_new_n787__,
    new_new_n788__, new_new_n789__, new_new_n790__, new_new_n791__,
    new_new_n792__, new_new_n793__, new_new_n794__, new_new_n796__,
    new_new_n798__, new_new_n800__, new_new_n802__, new_new_n804__,
    new_new_n806__, new_new_n808__, new_new_n810__, new_new_n812__,
    new_new_n814__, new_new_n816__, new_new_n818__, new_new_n820__,
    new_new_n822__, new_new_n824__, new_new_n826__, new_new_n828__,
    new_new_n830__, new_new_n832__, new_new_n834__, new_new_n836__,
    new_new_n838__, new_new_n840__, new_new_n842__, new_new_n844__,
    new_new_n846__, new_new_n848__, new_new_n849__, new_new_n850__,
    new_new_n851__, new_new_n852__, new_new_n853__, new_new_n854__,
    new_new_n855__, new_new_n856__, new_new_n857__, new_new_n858__,
    new_new_n859__, new_new_n860__, new_new_n861__, new_new_n862__,
    new_new_n863__, new_new_n864__, new_new_n865__, new_new_n866__,
    new_new_n867__, new_new_n868__, new_new_n869__, new_new_n870__,
    new_new_n871__, new_new_n872__, new_new_n873__, new_new_n874__,
    new_new_n875__, new_new_n876__, new_new_n877__, new_new_n878__,
    new_new_n879__, new_new_n880__, new_new_n881__, new_new_n882__,
    new_new_n883__, new_new_n884__, new_new_n885__, new_new_n886__,
    new_new_n887__, new_new_n888__, new_new_n889__, new_new_n890__,
    new_new_n891__, new_new_n892__, new_new_n893__, new_new_n894__,
    new_new_n895__, new_new_n896__, new_new_n897__, new_new_n898__,
    new_new_n899__, new_new_n900__, new_new_n901__, new_new_n902__,
    new_new_n903__, new_new_n904__, new_new_n905__, new_new_n906__,
    new_new_n907__, new_new_n908__, new_new_n909__, new_new_n910__,
    new_new_n911__, new_new_n912__, new_new_n913__, new_new_n914__,
    new_new_n915__, new_new_n916__, new_new_n917__, new_new_n918__,
    new_new_n919__, new_new_n920__, new_new_n921__, new_new_n922__,
    new_new_n923__, new_new_n924__, new_new_n925__, new_new_n926__,
    new_new_n927__, new_new_n928__, new_new_n929__, new_new_n930__,
    new_new_n931__, new_new_n932__, new_new_n933__, new_new_n934__,
    new_new_n935__, new_new_n936__, new_new_n937__, new_new_n938__,
    new_new_n939__, new_new_n940__, new_new_n941__, new_new_n942__,
    new_new_n943__, new_new_n944__, new_new_n945__, new_new_n946__,
    new_new_n947__, new_new_n948__, new_new_n949__, new_new_n950__,
    new_new_n951__, new_new_n952__, new_new_n953__, new_new_n954__,
    new_new_n955__, new_new_n956__, new_new_n957__, new_new_n958__,
    new_new_n959__, new_new_n960__, new_new_n961__, new_new_n962__,
    new_new_n963__, new_new_n964__, new_new_n965__, new_new_n966__,
    new_new_n967__, new_new_n968__, new_new_n969__, new_new_n970__,
    new_new_n971__, new_new_n972__, new_new_n973__, new_new_n974__,
    new_new_n975__, new_new_n976__, new_new_n977__, new_new_n978__,
    new_new_n979__, new_new_n980__, new_new_n981__, new_new_n982__,
    new_new_n983__, new_new_n984__, new_new_n985__, new_new_n986__,
    new_new_n987__, new_new_n988__, new_new_n989__, new_new_n990__,
    new_new_n991__, new_new_n992__, new_new_n993__, new_new_n994__,
    new_new_n995__, new_new_n996__, new_new_n997__, new_new_n998__,
    new_new_n999__, new_new_n1000__, new_new_n1001__, new_new_n1002__,
    new_new_n1003__, new_new_n1004__, new_new_n1005__, new_new_n1006__,
    new_new_n1007__, new_new_n1008__, new_new_n1009__, new_new_n1010__,
    new_new_n1011__, new_new_n1012__, new_new_n1013__, new_new_n1014__,
    new_new_n1015__, new_new_n1016__, new_new_n1017__, new_new_n1018__,
    new_new_n1019__, new_new_n1020__, new_new_n1021__, new_new_n1022__,
    new_new_n1023__, new_new_n1024__, new_new_n1025__, new_new_n1026__,
    new_new_n1027__, new_new_n1028__, new_new_n1029__, new_new_n1030__,
    new_new_n1031__, new_new_n1032__, new_new_n1033__, new_new_n1034__,
    new_new_n1035__, new_new_n1036__, new_new_n1037__, new_new_n1038__,
    new_new_n1039__, new_new_n1040__, new_new_n1041__, new_new_n1042__,
    new_new_n1043__, new_new_n1044__, new_new_n1045__, new_new_n1046__,
    new_new_n1047__, new_new_n1048__, new_new_n1049__, new_new_n1050__,
    new_new_n1051__, new_new_n1052__, new_new_n1053__, new_new_n1054__,
    new_new_n1055__, new_new_n1056__, new_new_n1057__, new_new_n1058__,
    new_new_n1059__, new_new_n1060__, new_new_n1061__, new_new_n1062__,
    new_new_n1063__, new_new_n1064__, new_new_n1065__, new_new_n1066__,
    new_new_n1067__, new_new_n1068__, new_new_n1069__, new_new_n1070__,
    new_new_n1071__, new_new_n1072__, new_new_n1073__, new_new_n1074__,
    new_new_n1075__, new_new_n1076__, new_new_n1077__, new_new_n1078__,
    new_new_n1079__, new_new_n1080__, new_new_n1081__, new_new_n1082__,
    new_new_n1083__, new_new_n1084__, new_new_n1085__, new_new_n1086__,
    new_new_n1087__, new_new_n1088__, new_new_n1089__, new_new_n1090__,
    new_new_n1091__, new_new_n1092__, new_new_n1093__, new_new_n1094__,
    new_new_n1095__, new_new_n1096__, new_new_n1097__, new_new_n1098__,
    new_new_n1099__, new_new_n1100__, new_new_n1101__, new_new_n1102__,
    new_new_n1103__, new_new_n1104__, new_new_n1105__, new_new_n1106__,
    new_new_n1107__, new_new_n1108__, new_new_n1304__, new_new_n1305__,
    new_new_n1306__, new_new_n1307__, new_new_n1308__, new_new_n1309__,
    new_new_n1310__, new_new_n1311__, new_new_n1312__, new_new_n1313__,
    new_new_n1314__, new_new_n1315__, new_new_n1316__, new_new_n1317__,
    new_new_n1318__, new_new_n1319__, new_new_n1320__, new_new_n1321__,
    new_new_n1322__, new_new_n1323__, new_new_n1324__, new_new_n1325__,
    new_new_n1326__, new_new_n1327__, new_new_n1328__, new_new_n1329__,
    new_new_n1330__, new_new_n1331__, new_new_n1332__, new_new_n1333__,
    new_new_n1334__, new_new_n1335__, new_new_n1336__, new_new_n1337__,
    new_new_n1338__, new_new_n1339__, new_new_n1340__, new_new_n1341__,
    new_new_n1342__, new_new_n1343__, new_new_n1344__, new_new_n1345__,
    new_new_n1346__, new_new_n1347__, new_new_n1348__, new_new_n1349__,
    new_new_n1350__, new_new_n1351__, new_new_n1352__, new_new_n1353__,
    new_new_n1354__, new_new_n1355__, new_new_n1356__, new_new_n1357__,
    new_new_n1358__, new_new_n1359__, new_new_n1360__, new_new_n1361__,
    new_new_n1362__, new_new_n1363__, new_new_n1364__, new_new_n1365__,
    new_new_n1366__, new_new_n1367__, new_new_n1368__, new_new_n1369__,
    new_new_n1370__, new_new_n1371__, new_new_n1372__, new_new_n1373__,
    new_new_n1374__, new_new_n1375__, new_new_n1376__, new_new_n1377__,
    new_new_n1378__, new_new_n1379__, new_new_n1380__, new_new_n1381__,
    new_new_n1382__, new_new_n1383__, new_new_n1384__, new_new_n1385__,
    new_new_n1386__, new_new_n1387__, new_new_n1388__, new_new_n1389__,
    new_new_n1390__, new_new_n1391__, new_new_n1392__, new_new_n1393__,
    new_new_n1394__, new_new_n1395__, new_new_n1396__, new_new_n1397__,
    new_new_n1398__, new_new_n1399__, new_new_n1400__, new_new_n1401__,
    new_new_n1402__, new_new_n1403__, new_new_n1404__, new_new_n1405__,
    new_new_n1406__, new_new_n1407__, new_new_n1408__, new_new_n1409__,
    new_new_n1410__, new_new_n1411__, new_new_n1412__, new_new_n1413__,
    new_new_n1414__, new_new_n1415__, new_new_n1416__, new_new_n1417__,
    new_new_n1418__, new_new_n1419__, new_new_n1420__, new_new_n1421__,
    new_new_n1422__, new_new_n1423__, new_new_n1424__, new_new_n1425__,
    new_new_n1426__, new_new_n1427__, new_new_n1428__, new_new_n1429__,
    new_new_n1430__, new_new_n1431__, new_new_n1432__, new_new_n1433__,
    new_new_n1434__, new_new_n1435__, new_new_n1436__, new_new_n1437__,
    new_new_n1438__, new_new_n1439__, new_new_n1440__, new_new_n1441__,
    new_new_n1442__, new_new_n1443__, new_new_n1444__, new_new_n1445__,
    new_new_n1446__, new_new_n1447__, new_new_n1448__, new_new_n1449__,
    new_new_n1450__, n2012, n2015, n2018, n2021, n2024, n2027, n2030,
    n2033, n2036, n2039, n2042, n2045, n2048, n2051, n2054, n2057, n2060,
    n2063, n2066, n2069, n2072, n2075, n2078, n2081, n2084, n2087, n2090,
    n2093, n2096, n2099, n2102, n2105, n2108, n2111, n2114, n2117, n2120,
    n2123, n2126, n2129, n2132, n2135, n2138, n2141, n2144, n2147, n2150,
    n2153, n2156, n2159, n2162, n2165, n2168, n2171, n2174, n2177, n2180,
    n2183, n2186, n2189, n2192, n2195, n2198, n2201, n2204, n2207, n2210,
    n2213, n2216, n2219, n2222, n2225, n2228, n2231, n2234, n2237, n2240,
    n2243, n2246, n2249, n2252, n2255, n2258, n2261, n2264, n2267, n2270,
    n2273, n2276, n2279, n2282, n2285, n2288, n2291, n2294, n2297, n2300,
    n2303, n2306, n2309, n2312, n2315, n2318, n2321, n2324, n2327, n2330,
    n2333, n2336, n2339, n2342, n2345, n2348, n2351, n2354, n2357, n2360,
    n2363, n2366, n2369, n2372, n2375, n2378, n2381, n2384, n2387, n2390,
    n2393, n2396, n2399, n2402, n2405, n2408, n2411, n2414, n2417, n2420,
    n2423, n2426, n2429, n2432, n2435, n2438, n2441, n2444, n2447, n2450,
    n2453, n2456, n2459, n2462, n2465, n2468, n2471, n2474, n2477, n2480,
    n2483, n2486, n2489, n2492, n2495, n2498, n2501, n2504, n2507, n2510,
    n2513, n2516, n2519, n2522, n2525, n2528, n2531, n2534, n2537, n2540,
    n2543, n2546, n2549, n2552, n2555, n2558, n2561, n2564, n2567, n2570,
    n2573;
  buf1  g000(.din(G1), .dout(new_new_n420__));
  buf1  g001(.din(G2), .dout(new_new_n422__));
  buf1  g002(.din(G3), .dout(new_new_n424__));
  buf1  g003(.din(G4), .dout(new_new_n426__));
  buf1  g004(.din(G5), .dout(new_new_n428__));
  buf1  g005(.din(G6), .dout(new_new_n430__));
  buf1  g006(.din(G7), .dout(new_new_n432__));
  buf1  g007(.din(G8), .dout(new_new_n434__));
  buf1  g008(.din(G9), .dout(new_new_n436__));
  buf1  g009(.din(G10), .dout(new_new_n438__));
  buf1  g010(.din(G11), .dout(new_new_n440__));
  buf1  g011(.din(G12), .dout(new_new_n442__));
  buf1  g012(.din(G13), .dout(new_new_n444__));
  buf1  g013(.din(G14), .dout(new_new_n446__));
  buf1  g014(.din(G15), .dout(new_new_n448__));
  buf1  g015(.din(G16), .dout(new_new_n450__));
  buf1  g016(.din(G17), .dout(new_new_n452__));
  buf1  g017(.din(G18), .dout(new_new_n454__));
  buf1  g018(.din(G19), .dout(new_new_n456__));
  buf1  g019(.din(G20), .dout(new_new_n458__));
  buf1  g020(.din(G21), .dout(new_new_n460__));
  buf1  g021(.din(G22), .dout(new_new_n462__));
  buf1  g022(.din(G23), .dout(new_new_n464__));
  buf1  g023(.din(G24), .dout(new_new_n466__));
  buf1  g024(.din(G25), .dout(new_new_n468__));
  buf1  g025(.din(G26), .dout(new_new_n470__));
  buf1  g026(.din(G27), .dout(new_new_n472__));
  buf1  g027(.din(G28), .dout(new_new_n474__));
  buf1  g028(.din(G29), .dout(new_new_n476__));
  buf1  g029(.din(G30), .dout(new_new_n478__));
  buf1  g030(.din(G31), .dout(new_new_n480__));
  buf1  g031(.din(G32), .dout(new_new_n482__));
  buf1  g032(.din(G33), .dout(new_new_n484__));
  buf1  g033(.din(G34), .dout(new_new_n486__));
  buf1  g034(.din(G35), .dout(new_new_n488__));
  buf1  g035(.din(G36), .dout(new_new_n490__));
  buf1  g036(.din(n205_lo), .dout(new_new_n492__));
  not1  g037(.din(n205_lo), .dout(new_new_n493__));
  not1  g038(.din(n214_lo), .dout(new_new_n495__));
  buf1  g039(.din(n217_lo), .dout(new_new_n496__));
  buf1  g040(.din(n226_lo), .dout(new_new_n498__));
  buf1  g041(.din(n229_lo), .dout(new_new_n500__));
  buf1  g042(.din(n232_lo), .dout(new_new_n502__));
  not1  g043(.din(n232_lo), .dout(new_new_n503__));
  not1  g044(.din(n238_lo), .dout(new_new_n505__));
  buf1  g045(.din(n241_lo), .dout(new_new_n506__));
  not1  g046(.din(n241_lo), .dout(new_new_n507__));
  buf1  g047(.din(n250_lo), .dout(new_new_n508__));
  buf1  g048(.din(n253_lo), .dout(new_new_n510__));
  buf1  g049(.din(n256_lo), .dout(new_new_n512__));
  not1  g050(.din(n256_lo), .dout(new_new_n513__));
  not1  g051(.din(n262_lo), .dout(new_new_n515__));
  buf1  g052(.din(n265_lo), .dout(new_new_n516__));
  not1  g053(.din(n274_lo), .dout(new_new_n519__));
  buf1  g054(.din(n277_lo), .dout(new_new_n520__));
  buf1  g055(.din(n280_lo), .dout(new_new_n522__));
  not1  g056(.din(n280_lo), .dout(new_new_n523__));
  buf1  g057(.din(n286_lo), .dout(new_new_n524__));
  buf1  g058(.din(n289_lo), .dout(new_new_n526__));
  not1  g059(.din(n289_lo), .dout(new_new_n527__));
  buf1  g060(.din(n298_lo), .dout(new_new_n528__));
  not1  g061(.din(n298_lo), .dout(new_new_n529__));
  buf1  g062(.din(n301_lo), .dout(new_new_n530__));
  buf1  g063(.din(n304_lo), .dout(new_new_n532__));
  not1  g064(.din(n304_lo), .dout(new_new_n533__));
  buf1  g065(.din(n310_lo), .dout(new_new_n534__));
  buf1  g066(.din(n313_lo), .dout(new_new_n536__));
  buf1  g067(.din(n322_lo), .dout(new_new_n538__));
  not1  g068(.din(n322_lo), .dout(new_new_n539__));
  buf1  g069(.din(n325_lo), .dout(new_new_n540__));
  buf1  g070(.din(n328_lo), .dout(new_new_n542__));
  not1  g071(.din(n328_lo), .dout(new_new_n543__));
  buf1  g072(.din(n334_lo), .dout(new_new_n544__));
  not1  g073(.din(n334_lo), .dout(new_new_n545__));
  buf1  g074(.din(n337_lo), .dout(new_new_n546__));
  not1  g075(.din(n337_lo), .dout(new_new_n547__));
  buf1  g076(.din(n346_lo), .dout(new_new_n548__));
  not1  g077(.din(n346_lo), .dout(new_new_n549__));
  buf1  g078(.din(n349_lo), .dout(new_new_n550__));
  buf1  g079(.din(n352_lo), .dout(new_new_n552__));
  not1  g080(.din(n352_lo), .dout(new_new_n553__));
  buf1  g081(.din(n358_lo), .dout(new_new_n554__));
  not1  g082(.din(n358_lo), .dout(new_new_n555__));
  buf1  g083(.din(n361_lo), .dout(new_new_n556__));
  buf1  g084(.din(n370_lo), .dout(new_new_n558__));
  not1  g085(.din(n370_lo), .dout(new_new_n559__));
  buf1  g086(.din(n373_lo), .dout(new_new_n560__));
  buf1  g087(.din(n376_lo), .dout(new_new_n562__));
  not1  g088(.din(n376_lo), .dout(new_new_n563__));
  buf1  g089(.din(n382_lo), .dout(new_new_n564__));
  not1  g090(.din(n382_lo), .dout(new_new_n565__));
  buf1  g091(.din(n385_lo), .dout(new_new_n566__));
  not1  g092(.din(n385_lo), .dout(new_new_n567__));
  buf1  g093(.din(n394_lo), .dout(new_new_n568__));
  not1  g094(.din(n394_lo), .dout(new_new_n569__));
  buf1  g095(.din(n397_lo), .dout(new_new_n570__));
  buf1  g096(.din(n400_lo), .dout(new_new_n572__));
  not1  g097(.din(n400_lo), .dout(new_new_n573__));
  buf1  g098(.din(n406_lo), .dout(new_new_n574__));
  not1  g099(.din(n406_lo), .dout(new_new_n575__));
  buf1  g100(.din(n409_lo), .dout(new_new_n576__));
  buf1  g101(.din(n418_lo), .dout(new_new_n578__));
  not1  g102(.din(n418_lo), .dout(new_new_n579__));
  buf1  g103(.din(n421_lo), .dout(new_new_n580__));
  buf1  g104(.din(n424_lo), .dout(new_new_n582__));
  not1  g105(.din(n424_lo), .dout(new_new_n583__));
  buf1  g106(.din(n430_lo), .dout(new_new_n584__));
  not1  g107(.din(n430_lo), .dout(new_new_n585__));
  buf1  g108(.din(n433_lo), .dout(new_new_n586__));
  not1  g109(.din(n433_lo), .dout(new_new_n587__));
  buf1  g110(.din(n442_lo), .dout(new_new_n588__));
  buf1  g111(.din(n445_lo), .dout(new_new_n590__));
  buf1  g112(.din(n448_lo), .dout(new_new_n592__));
  not1  g113(.din(n448_lo), .dout(new_new_n593__));
  buf1  g114(.din(n454_lo), .dout(new_new_n594__));
  not1  g115(.din(n454_lo), .dout(new_new_n595__));
  buf1  g116(.din(n457_lo), .dout(new_new_n596__));
  not1  g117(.din(n466_lo), .dout(new_new_n599__));
  buf1  g118(.din(n469_lo), .dout(new_new_n600__));
  buf1  g119(.din(n472_lo), .dout(new_new_n602__));
  not1  g120(.din(n472_lo), .dout(new_new_n603__));
  buf1  g121(.din(n478_lo), .dout(new_new_n604__));
  buf1  g122(.din(n481_lo), .dout(new_new_n606__));
  not1  g123(.din(n481_lo), .dout(new_new_n607__));
  buf1  g124(.din(n490_lo), .dout(new_new_n608__));
  not1  g125(.din(n490_lo), .dout(new_new_n609__));
  buf1  g126(.din(n493_lo), .dout(new_new_n610__));
  buf1  g127(.din(n496_lo), .dout(new_new_n612__));
  not1  g128(.din(n496_lo), .dout(new_new_n613__));
  buf1  g129(.din(n502_lo), .dout(new_new_n614__));
  buf1  g130(.din(n505_lo), .dout(new_new_n616__));
  buf1  g131(.din(n514_lo), .dout(new_new_n618__));
  not1  g132(.din(n514_lo), .dout(new_new_n619__));
  buf1  g133(.din(n517_lo), .dout(new_new_n620__));
  buf1  g134(.din(n520_lo), .dout(new_new_n622__));
  not1  g135(.din(n520_lo), .dout(new_new_n623__));
  buf1  g136(.din(n526_lo), .dout(new_new_n624__));
  not1  g137(.din(n526_lo), .dout(new_new_n625__));
  buf1  g138(.din(n529_lo), .dout(new_new_n626__));
  not1  g139(.din(n529_lo), .dout(new_new_n627__));
  buf1  g140(.din(n538_lo), .dout(new_new_n628__));
  buf1  g141(.din(n541_lo), .dout(new_new_n630__));
  buf1  g142(.din(n544_lo), .dout(new_new_n632__));
  not1  g143(.din(n544_lo), .dout(new_new_n633__));
  buf1  g144(.din(n550_lo), .dout(new_new_n634__));
  not1  g145(.din(n550_lo), .dout(new_new_n635__));
  buf1  g146(.din(n553_lo), .dout(new_new_n636__));
  not1  g147(.din(n562_lo), .dout(new_new_n639__));
  buf1  g148(.din(n565_lo), .dout(new_new_n640__));
  buf1  g149(.din(n568_lo), .dout(new_new_n642__));
  not1  g150(.din(n568_lo), .dout(new_new_n643__));
  buf1  g151(.din(n574_lo), .dout(new_new_n644__));
  buf1  g152(.din(n577_lo), .dout(new_new_n646__));
  not1  g153(.din(n577_lo), .dout(new_new_n647__));
  buf1  g154(.din(n586_lo), .dout(new_new_n648__));
  buf1  g155(.din(n589_lo), .dout(new_new_n650__));
  buf1  g156(.din(n592_lo), .dout(new_new_n652__));
  not1  g157(.din(n592_lo), .dout(new_new_n653__));
  buf1  g158(.din(n598_lo), .dout(new_new_n654__));
  buf1  g159(.din(n601_lo), .dout(new_new_n656__));
  not1  g160(.din(n610_lo), .dout(new_new_n659__));
  buf1  g161(.din(n613_lo), .dout(new_new_n660__));
  buf1  g162(.din(n616_lo), .dout(new_new_n662__));
  not1  g163(.din(n616_lo), .dout(new_new_n663__));
  buf1  g164(.din(n622_lo), .dout(new_new_n664__));
  buf1  g165(.din(n625_lo), .dout(new_new_n666__));
  buf1  g166(.din(n628_lo), .dout(new_new_n668__));
  not1  g167(.din(n628_lo), .dout(new_new_n669__));
  buf1  g168(.din(n634_lo), .dout(new_new_n670__));
  buf1  g169(.din(n316_inv), .dout(new_new_n672__));
  buf1  g170(.din(n319_inv), .dout(new_new_n674__));
  buf1  g171(.din(n997_o2), .dout(new_new_n676__));
  buf1  g172(.din(n998_o2), .dout(new_new_n678__));
  buf1  g173(.din(n999_o2), .dout(new_new_n680__));
  buf1  g174(.din(n1000_o2), .dout(new_new_n682__));
  buf1  g175(.din(n1001_o2), .dout(new_new_n684__));
  buf1  g176(.din(n1002_o2), .dout(new_new_n686__));
  buf1  g177(.din(n1003_o2), .dout(new_new_n688__));
  buf1  g178(.din(n1004_o2), .dout(new_new_n690__));
  buf1  g179(.din(n1005_o2), .dout(new_new_n692__));
  buf1  g180(.din(n1015_o2), .dout(new_new_n694__));
  buf1  g181(.din(n1016_o2), .dout(new_new_n696__));
  buf1  g182(.din(n1017_o2), .dout(new_new_n698__));
  buf1  g183(.din(n1018_o2), .dout(new_new_n700__));
  buf1  g184(.din(n1019_o2), .dout(new_new_n702__));
  buf1  g185(.din(n1020_o2), .dout(new_new_n704__));
  buf1  g186(.din(n1021_o2), .dout(new_new_n706__));
  buf1  g187(.din(n1022_o2), .dout(new_new_n708__));
  buf1  g188(.din(n1023_o2), .dout(new_new_n710__));
  buf1  g189(.din(n376_1_inv), .dout(new_new_n712__));
  buf1  g190(.din(n235_lo_buf_o2), .dout(new_new_n714__));
  buf1  g191(.din(n283_lo_buf_o2), .dout(new_new_n716__));
  buf1  g192(.din(n331_lo_buf_o2), .dout(new_new_n718__));
  buf1  g193(.din(n379_lo_buf_o2), .dout(new_new_n720__));
  buf1  g194(.din(n427_lo_buf_o2), .dout(new_new_n722__));
  buf1  g195(.din(n475_lo_buf_o2), .dout(new_new_n724__));
  buf1  g196(.din(n523_lo_buf_o2), .dout(new_new_n726__));
  buf1  g197(.din(n571_lo_buf_o2), .dout(new_new_n728__));
  buf1  g198(.din(n619_lo_buf_o2), .dout(new_new_n730__));
  buf1  g199(.din(n406_1_inv), .dout(new_new_n732__));
  not1  g200(.din(G223_o2), .dout(new_new_n735__));
  not1  g201(.din(G226_o2), .dout(new_new_n737__));
  not1  g202(.din(G229_o2), .dout(new_new_n739__));
  not1  g203(.din(G232_o2), .dout(new_new_n741__));
  not1  g204(.din(G235_o2), .dout(new_new_n743__));
  not1  g205(.din(G238_o2), .dout(new_new_n745__));
  not1  g206(.din(G242_o2), .dout(new_new_n747__));
  not1  g207(.din(G246_o2), .dout(new_new_n749__));
  not1  g208(.din(G250_o2), .dout(new_new_n751__));
  buf1  g209(.din(n259_lo_buf_o2), .dout(new_new_n752__));
  buf1  g210(.din(n307_lo_buf_o2), .dout(new_new_n754__));
  buf1  g211(.din(n355_lo_buf_o2), .dout(new_new_n756__));
  buf1  g212(.din(n403_lo_buf_o2), .dout(new_new_n758__));
  buf1  g213(.din(n451_lo_buf_o2), .dout(new_new_n760__));
  buf1  g214(.din(n499_lo_buf_o2), .dout(new_new_n762__));
  buf1  g215(.din(n547_lo_buf_o2), .dout(new_new_n764__));
  buf1  g216(.din(n595_lo_buf_o2), .dout(new_new_n766__));
  buf1  g217(.din(n631_lo_buf_o2), .dout(new_new_n768__));
  buf1  g218(.din(G213_o2), .dout(new_new_n770__));
  not1  g219(.din(G213_o2), .dout(new_new_n771__));
  buf1  g220(.din(G318_o2), .dout(new_new_n772__));
  not1  g221(.din(G318_o2), .dout(new_new_n773__));
  buf1  g222(.din(G358_o2), .dout(new_new_n774__));
  not1  g223(.din(G358_o2), .dout(new_new_n775__));
  buf1  g224(.din(G259_o2), .dout(new_new_n776__));
  not1  g225(.din(G259_o2), .dout(new_new_n777__));
  buf1  g226(.din(G263_o2), .dout(new_new_n778__));
  not1  g227(.din(G263_o2), .dout(new_new_n779__));
  buf1  g228(.din(G266_o2), .dout(new_new_n780__));
  not1  g229(.din(G266_o2), .dout(new_new_n781__));
  buf1  g230(.din(G269_o2), .dout(new_new_n782__));
  not1  g231(.din(G269_o2), .dout(new_new_n783__));
  buf1  g232(.din(G272_o2), .dout(new_new_n784__));
  not1  g233(.din(G272_o2), .dout(new_new_n785__));
  buf1  g234(.din(G275_o2), .dout(new_new_n786__));
  not1  g235(.din(G275_o2), .dout(new_new_n787__));
  buf1  g236(.din(G278_o2), .dout(new_new_n788__));
  not1  g237(.din(G278_o2), .dout(new_new_n789__));
  buf1  g238(.din(G281_o2), .dout(new_new_n790__));
  not1  g239(.din(G281_o2), .dout(new_new_n791__));
  buf1  g240(.din(G284_o2), .dout(new_new_n792__));
  not1  g241(.din(G284_o2), .dout(new_new_n793__));
  buf1  g242(.din(n211_lo_buf_o2), .dout(new_new_n794__));
  buf1  g243(.din(n247_lo_buf_o2), .dout(new_new_n796__));
  buf1  g244(.din(n295_lo_buf_o2), .dout(new_new_n798__));
  buf1  g245(.din(n343_lo_buf_o2), .dout(new_new_n800__));
  buf1  g246(.din(n391_lo_buf_o2), .dout(new_new_n802__));
  buf1  g247(.din(n439_lo_buf_o2), .dout(new_new_n804__));
  buf1  g248(.din(n487_lo_buf_o2), .dout(new_new_n806__));
  buf1  g249(.din(n535_lo_buf_o2), .dout(new_new_n808__));
  buf1  g250(.din(n583_lo_buf_o2), .dout(new_new_n810__));
  buf1  g251(.din(G158_o2), .dout(new_new_n812__));
  buf1  g252(.din(G184_o2), .dout(new_new_n814__));
  buf1  g253(.din(G186_o2), .dout(new_new_n816__));
  buf1  g254(.din(G188_o2), .dout(new_new_n818__));
  buf1  g255(.din(G190_o2), .dout(new_new_n820__));
  buf1  g256(.din(G192_o2), .dout(new_new_n822__));
  buf1  g257(.din(G194_o2), .dout(new_new_n824__));
  buf1  g258(.din(G196_o2), .dout(new_new_n826__));
  buf1  g259(.din(G198_o2), .dout(new_new_n828__));
  buf1  g260(.din(n223_lo_buf_o2), .dout(new_new_n830__));
  buf1  g261(.din(n271_lo_buf_o2), .dout(new_new_n832__));
  buf1  g262(.din(n319_lo_buf_o2), .dout(new_new_n834__));
  buf1  g263(.din(n367_lo_buf_o2), .dout(new_new_n836__));
  buf1  g264(.din(n415_lo_buf_o2), .dout(new_new_n838__));
  buf1  g265(.din(n463_lo_buf_o2), .dout(new_new_n840__));
  buf1  g266(.din(n511_lo_buf_o2), .dout(new_new_n842__));
  buf1  g267(.din(n559_lo_buf_o2), .dout(new_new_n844__));
  buf1  g268(.din(n607_lo_buf_o2), .dout(new_new_n846__));
  buf1  g269(.din(n580_inv), .dout(new_new_n848__));
  not1  g270(.din(n580_inv), .dout(new_new_n849__));
  buf1  g271(.din(G154_o2), .dout(new_new_n850__));
  not1  g272(.din(G154_o2), .dout(new_new_n851__));
  buf1  g273(.din(G159_o2), .dout(new_new_n852__));
  not1  g274(.din(G159_o2), .dout(new_new_n853__));
  buf1  g275(.din(G162_o2), .dout(new_new_n854__));
  not1  g276(.din(G162_o2), .dout(new_new_n855__));
  buf1  g277(.din(G165_o2), .dout(new_new_n856__));
  not1  g278(.din(G165_o2), .dout(new_new_n857__));
  buf1  g279(.din(G168_o2), .dout(new_new_n858__));
  not1  g280(.din(G168_o2), .dout(new_new_n859__));
  buf1  g281(.din(G171_o2), .dout(new_new_n860__));
  not1  g282(.din(G171_o2), .dout(new_new_n861__));
  buf1  g283(.din(G174_o2), .dout(new_new_n862__));
  not1  g284(.din(G174_o2), .dout(new_new_n863__));
  buf1  g285(.din(G177_o2), .dout(new_new_n864__));
  not1  g286(.din(G177_o2), .dout(new_new_n865__));
  buf1  g287(.din(G180_o2), .dout(new_new_n866__));
  not1  g288(.din(G180_o2), .dout(new_new_n867__));
  or1   g289(.dina(new_new_n1306__), .dinb(new_new_n495__), .dout(new_new_n868__));
  or1   g290(.dina(new_new_n1310__), .dinb(new_new_n505__), .dout(new_new_n869__));
  or1   g291(.dina(new_new_n1314__), .dinb(new_new_n515__), .dout(new_new_n870__));
  and1  g292(.dina(new_new_n868__), .dinb(new_new_n498__), .dout(new_new_n871__));
  and1  g293(.dina(new_new_n871__), .dinb(new_new_n869__), .dout(new_new_n872__));
  and1  g294(.dina(new_new_n872__), .dinb(new_new_n870__), .dout(new_new_n873__));
  and1  g295(.dina(new_new_n1318__), .dinb(new_new_n508__), .dout(new_new_n874__));
  and1  g296(.dina(new_new_n1325__), .dinb(new_new_n524__), .dout(new_new_n875__));
  and1  g297(.dina(new_new_n1332__), .dinb(new_new_n534__), .dout(new_new_n876__));
  or1   g298(.dina(new_new_n875__), .dinb(new_new_n874__), .dout(new_new_n877__));
  or1   g299(.dina(new_new_n877__), .dinb(new_new_n876__), .dout(new_new_n878__));
  or1   g300(.dina(new_new_n878__), .dinb(new_new_n519__), .dout(new_new_n879__));
  and1  g301(.dina(new_new_n1318__), .dinb(new_new_n528__), .dout(new_new_n880__));
  or1   g302(.dina(new_new_n1306__), .dinb(new_new_n529__), .dout(new_new_n881__));
  and1  g303(.dina(new_new_n1325__), .dinb(new_new_n544__), .dout(new_new_n882__));
  or1   g304(.dina(new_new_n1310__), .dinb(new_new_n545__), .dout(new_new_n883__));
  and1  g305(.dina(new_new_n1332__), .dinb(new_new_n554__), .dout(new_new_n884__));
  or1   g306(.dina(new_new_n1314__), .dinb(new_new_n555__), .dout(new_new_n885__));
  and1  g307(.dina(new_new_n883__), .dinb(new_new_n881__), .dout(new_new_n886__));
  or1   g308(.dina(new_new_n882__), .dinb(new_new_n880__), .dout(new_new_n887__));
  and1  g309(.dina(new_new_n886__), .dinb(new_new_n885__), .dout(new_new_n888__));
  or1   g310(.dina(new_new_n887__), .dinb(new_new_n884__), .dout(new_new_n889__));
  and1  g311(.dina(new_new_n888__), .dinb(new_new_n538__), .dout(new_new_n890__));
  or1   g312(.dina(new_new_n889__), .dinb(new_new_n539__), .dout(new_new_n891__));
  and1  g313(.dina(new_new_n1319__), .dinb(new_new_n548__), .dout(new_new_n892__));
  or1   g314(.dina(new_new_n1305__), .dinb(new_new_n549__), .dout(new_new_n893__));
  and1  g315(.dina(new_new_n1326__), .dinb(new_new_n564__), .dout(new_new_n894__));
  or1   g316(.dina(new_new_n1309__), .dinb(new_new_n565__), .dout(new_new_n895__));
  and1  g317(.dina(new_new_n1333__), .dinb(new_new_n574__), .dout(new_new_n896__));
  or1   g318(.dina(new_new_n1313__), .dinb(new_new_n575__), .dout(new_new_n897__));
  and1  g319(.dina(new_new_n895__), .dinb(new_new_n893__), .dout(new_new_n898__));
  or1   g320(.dina(new_new_n894__), .dinb(new_new_n892__), .dout(new_new_n899__));
  and1  g321(.dina(new_new_n898__), .dinb(new_new_n897__), .dout(new_new_n900__));
  or1   g322(.dina(new_new_n899__), .dinb(new_new_n896__), .dout(new_new_n901__));
  and1  g323(.dina(new_new_n900__), .dinb(new_new_n558__), .dout(new_new_n902__));
  or1   g324(.dina(new_new_n901__), .dinb(new_new_n559__), .dout(new_new_n903__));
  and1  g325(.dina(new_new_n1319__), .dinb(new_new_n568__), .dout(new_new_n904__));
  or1   g326(.dina(new_new_n1307__), .dinb(new_new_n569__), .dout(new_new_n905__));
  and1  g327(.dina(new_new_n1326__), .dinb(new_new_n584__), .dout(new_new_n906__));
  or1   g328(.dina(new_new_n1311__), .dinb(new_new_n585__), .dout(new_new_n907__));
  and1  g329(.dina(new_new_n1333__), .dinb(new_new_n594__), .dout(new_new_n908__));
  or1   g330(.dina(new_new_n1315__), .dinb(new_new_n595__), .dout(new_new_n909__));
  and1  g331(.dina(new_new_n907__), .dinb(new_new_n905__), .dout(new_new_n910__));
  or1   g332(.dina(new_new_n906__), .dinb(new_new_n904__), .dout(new_new_n911__));
  and1  g333(.dina(new_new_n910__), .dinb(new_new_n909__), .dout(new_new_n912__));
  or1   g334(.dina(new_new_n911__), .dinb(new_new_n908__), .dout(new_new_n913__));
  and1  g335(.dina(new_new_n912__), .dinb(new_new_n578__), .dout(new_new_n914__));
  or1   g336(.dina(new_new_n913__), .dinb(new_new_n579__), .dout(new_new_n915__));
  and1  g337(.dina(new_new_n1321__), .dinb(new_new_n588__), .dout(new_new_n916__));
  and1  g338(.dina(new_new_n1328__), .dinb(new_new_n604__), .dout(new_new_n917__));
  and1  g339(.dina(new_new_n1335__), .dinb(new_new_n614__), .dout(new_new_n918__));
  or1   g340(.dina(new_new_n917__), .dinb(new_new_n916__), .dout(new_new_n919__));
  or1   g341(.dina(new_new_n919__), .dinb(new_new_n918__), .dout(new_new_n920__));
  or1   g342(.dina(new_new_n920__), .dinb(new_new_n599__), .dout(new_new_n921__));
  and1  g343(.dina(new_new_n1321__), .dinb(new_new_n608__), .dout(new_new_n922__));
  or1   g344(.dina(new_new_n1307__), .dinb(new_new_n609__), .dout(new_new_n923__));
  and1  g345(.dina(new_new_n1328__), .dinb(new_new_n624__), .dout(new_new_n924__));
  or1   g346(.dina(new_new_n1311__), .dinb(new_new_n625__), .dout(new_new_n925__));
  and1  g347(.dina(new_new_n1335__), .dinb(new_new_n634__), .dout(new_new_n926__));
  or1   g348(.dina(new_new_n1315__), .dinb(new_new_n635__), .dout(new_new_n927__));
  and1  g349(.dina(new_new_n925__), .dinb(new_new_n923__), .dout(new_new_n928__));
  or1   g350(.dina(new_new_n924__), .dinb(new_new_n922__), .dout(new_new_n929__));
  and1  g351(.dina(new_new_n928__), .dinb(new_new_n927__), .dout(new_new_n930__));
  or1   g352(.dina(new_new_n929__), .dinb(new_new_n926__), .dout(new_new_n931__));
  and1  g353(.dina(new_new_n930__), .dinb(new_new_n618__), .dout(new_new_n932__));
  or1   g354(.dina(new_new_n931__), .dinb(new_new_n619__), .dout(new_new_n933__));
  and1  g355(.dina(new_new_n1322__), .dinb(new_new_n628__), .dout(new_new_n934__));
  and1  g356(.dina(new_new_n1329__), .dinb(new_new_n644__), .dout(new_new_n935__));
  and1  g357(.dina(new_new_n1336__), .dinb(new_new_n654__), .dout(new_new_n936__));
  or1   g358(.dina(new_new_n935__), .dinb(new_new_n934__), .dout(new_new_n937__));
  or1   g359(.dina(new_new_n937__), .dinb(new_new_n936__), .dout(new_new_n938__));
  or1   g360(.dina(new_new_n938__), .dinb(new_new_n639__), .dout(new_new_n939__));
  and1  g361(.dina(new_new_n1322__), .dinb(new_new_n648__), .dout(new_new_n940__));
  and1  g362(.dina(new_new_n1329__), .dinb(new_new_n664__), .dout(new_new_n941__));
  and1  g363(.dina(new_new_n1336__), .dinb(new_new_n670__), .dout(new_new_n942__));
  or1   g364(.dina(new_new_n941__), .dinb(new_new_n940__), .dout(new_new_n943__));
  or1   g365(.dina(new_new_n943__), .dinb(new_new_n942__), .dout(new_new_n944__));
  or1   g366(.dina(new_new_n944__), .dinb(new_new_n659__), .dout(new_new_n945__));
  and1  g367(.dina(new_new_n891__), .dinb(new_new_n1337__), .dout(new_new_n946__));
  and1  g368(.dina(new_new_n1339__), .dinb(new_new_n1340__), .dout(new_new_n947__));
  and1  g369(.dina(new_new_n947__), .dinb(new_new_n1341__), .dout(new_new_n948__));
  and1  g370(.dina(new_new_n948__), .dinb(new_new_n1342__), .dout(new_new_n949__));
  and1  g371(.dina(new_new_n949__), .dinb(new_new_n1343__), .dout(new_new_n950__));
  and1  g372(.dina(new_new_n950__), .dinb(new_new_n1344__), .dout(new_new_n951__));
  and1  g373(.dina(new_new_n951__), .dinb(new_new_n945__), .dout(new_new_n952__));
  or1   g374(.dina(new_new_n952__), .dinb(new_new_n873__), .dout(new_new_n953__));
  or1   g375(.dina(new_new_n1340__), .dinb(new_new_n1345__), .dout(new_new_n954__));
  and1  g376(.dina(new_new_n1346__), .dinb(new_new_n1339__), .dout(new_new_n955__));
  and1  g377(.dina(new_new_n955__), .dinb(new_new_n1341__), .dout(new_new_n956__));
  or1   g378(.dina(new_new_n1347__), .dinb(new_new_n1345__), .dout(new_new_n957__));
  or1   g379(.dina(new_new_n1348__), .dinb(new_new_n1342__), .dout(new_new_n958__));
  or1   g380(.dina(new_new_n958__), .dinb(new_new_n1349__), .dout(new_new_n959__));
  or1   g381(.dina(new_new_n1349__), .dinb(new_new_n1347__), .dout(new_new_n960__));
  or1   g382(.dina(new_new_n960__), .dinb(new_new_n1343__), .dout(new_new_n961__));
  and1  g383(.dina(new_new_n1350__), .dinb(new_new_n1338__), .dout(new_new_n962__));
  and1  g384(.dina(new_new_n962__), .dinb(new_new_n961__), .dout(new_new_n963__));
  or1   g385(.dina(new_new_n1348__), .dinb(new_new_n932__), .dout(new_new_n964__));
  or1   g386(.dina(new_new_n964__), .dinb(new_new_n1344__), .dout(new_new_n965__));
  and1  g387(.dina(new_new_n1346__), .dinb(new_new_n1337__), .dout(new_new_n966__));
  and1  g388(.dina(new_new_n966__), .dinb(new_new_n1350__), .dout(new_new_n967__));
  and1  g389(.dina(new_new_n967__), .dinb(new_new_n965__), .dout(new_new_n968__));
  and1  g390(.dina(new_new_n1351__), .dinb(new_new_n1352__), .dout(new_new_n969__));
  or1   g391(.dina(new_new_n1353__), .dinb(new_new_n1354__), .dout(new_new_n970__));
  and1  g392(.dina(new_new_n969__), .dinb(new_new_n1355__), .dout(new_new_n971__));
  or1   g393(.dina(new_new_n970__), .dinb(new_new_n1356__), .dout(new_new_n972__));
  and1  g394(.dina(new_new_n971__), .dinb(new_new_n1357__), .dout(new_new_n973__));
  or1   g395(.dina(new_new_n972__), .dinb(new_new_n1358__), .dout(new_new_n974__));
  and1  g396(.dina(new_new_n973__), .dinb(new_new_n1359__), .dout(new_new_n975__));
  or1   g397(.dina(new_new_n974__), .dinb(new_new_n1360__), .dout(new_new_n976__));
  and1  g398(.dina(new_new_n975__), .dinb(new_new_n1361__), .dout(new_new_n977__));
  or1   g399(.dina(new_new_n976__), .dinb(new_new_n1362__), .dout(new_new_n978__));
  and1  g400(.dina(new_new_n977__), .dinb(new_new_n1363__), .dout(new_new_n979__));
  or1   g401(.dina(new_new_n978__), .dinb(new_new_n1364__), .dout(new_new_n980__));
  and1  g402(.dina(new_new_n979__), .dinb(new_new_n1365__), .dout(new_new_n981__));
  or1   g403(.dina(new_new_n980__), .dinb(new_new_n1366__), .dout(new_new_n982__));
  and1  g404(.dina(new_new_n981__), .dinb(new_new_n1367__), .dout(new_new_n983__));
  or1   g405(.dina(new_new_n982__), .dinb(new_new_n1368__), .dout(new_new_n984__));
  and1  g406(.dina(new_new_n1372__), .dinb(new_new_n777__), .dout(new_new_n985__));
  and1  g407(.dina(new_new_n1380__), .dinb(new_new_n776__), .dout(new_new_n986__));
  or1   g408(.dina(new_new_n986__), .dinb(new_new_n985__), .dout(new_new_n987__));
  and1  g409(.dina(new_new_n812__), .dinb(new_new_n735__), .dout(new_new_n988__));
  and1  g410(.dina(new_new_n988__), .dinb(new_new_n987__), .dout(new_new_n989__));
  and1  g411(.dina(new_new_n1372__), .dinb(new_new_n779__), .dout(new_new_n990__));
  and1  g412(.dina(new_new_n1380__), .dinb(new_new_n778__), .dout(new_new_n991__));
  or1   g413(.dina(new_new_n991__), .dinb(new_new_n990__), .dout(new_new_n992__));
  and1  g414(.dina(new_new_n814__), .dinb(new_new_n737__), .dout(new_new_n993__));
  and1  g415(.dina(new_new_n993__), .dinb(new_new_n992__), .dout(new_new_n994__));
  and1  g416(.dina(new_new_n1371__), .dinb(new_new_n781__), .dout(new_new_n995__));
  and1  g417(.dina(new_new_n1381__), .dinb(new_new_n780__), .dout(new_new_n996__));
  or1   g418(.dina(new_new_n996__), .dinb(new_new_n995__), .dout(new_new_n997__));
  and1  g419(.dina(new_new_n816__), .dinb(new_new_n739__), .dout(new_new_n998__));
  and1  g420(.dina(new_new_n998__), .dinb(new_new_n997__), .dout(new_new_n999__));
  and1  g421(.dina(new_new_n1373__), .dinb(new_new_n783__), .dout(new_new_n1000__));
  and1  g422(.dina(new_new_n1381__), .dinb(new_new_n782__), .dout(new_new_n1001__));
  or1   g423(.dina(new_new_n1001__), .dinb(new_new_n1000__), .dout(new_new_n1002__));
  and1  g424(.dina(new_new_n818__), .dinb(new_new_n741__), .dout(new_new_n1003__));
  and1  g425(.dina(new_new_n1003__), .dinb(new_new_n1002__), .dout(new_new_n1004__));
  and1  g426(.dina(new_new_n1373__), .dinb(new_new_n785__), .dout(new_new_n1005__));
  and1  g427(.dina(new_new_n1383__), .dinb(new_new_n784__), .dout(new_new_n1006__));
  or1   g428(.dina(new_new_n1006__), .dinb(new_new_n1005__), .dout(new_new_n1007__));
  and1  g429(.dina(new_new_n820__), .dinb(new_new_n743__), .dout(new_new_n1008__));
  and1  g430(.dina(new_new_n1008__), .dinb(new_new_n1007__), .dout(new_new_n1009__));
  and1  g431(.dina(new_new_n1375__), .dinb(new_new_n787__), .dout(new_new_n1010__));
  and1  g432(.dina(new_new_n1383__), .dinb(new_new_n786__), .dout(new_new_n1011__));
  or1   g433(.dina(new_new_n1011__), .dinb(new_new_n1010__), .dout(new_new_n1012__));
  and1  g434(.dina(new_new_n822__), .dinb(new_new_n745__), .dout(new_new_n1013__));
  and1  g435(.dina(new_new_n1013__), .dinb(new_new_n1012__), .dout(new_new_n1014__));
  and1  g436(.dina(new_new_n1375__), .dinb(new_new_n789__), .dout(new_new_n1015__));
  and1  g437(.dina(new_new_n1382__), .dinb(new_new_n788__), .dout(new_new_n1016__));
  or1   g438(.dina(new_new_n1016__), .dinb(new_new_n1015__), .dout(new_new_n1017__));
  and1  g439(.dina(new_new_n824__), .dinb(new_new_n747__), .dout(new_new_n1018__));
  and1  g440(.dina(new_new_n1018__), .dinb(new_new_n1017__), .dout(new_new_n1019__));
  and1  g441(.dina(new_new_n1376__), .dinb(new_new_n791__), .dout(new_new_n1020__));
  and1  g442(.dina(new_new_n1385__), .dinb(new_new_n790__), .dout(new_new_n1021__));
  or1   g443(.dina(new_new_n1021__), .dinb(new_new_n1020__), .dout(new_new_n1022__));
  and1  g444(.dina(new_new_n826__), .dinb(new_new_n749__), .dout(new_new_n1023__));
  and1  g445(.dina(new_new_n1023__), .dinb(new_new_n1022__), .dout(new_new_n1024__));
  and1  g446(.dina(new_new_n1376__), .dinb(new_new_n793__), .dout(new_new_n1025__));
  and1  g447(.dina(new_new_n1385__), .dinb(new_new_n792__), .dout(new_new_n1026__));
  or1   g448(.dina(new_new_n1026__), .dinb(new_new_n1025__), .dout(new_new_n1027__));
  and1  g449(.dina(new_new_n828__), .dinb(new_new_n751__), .dout(new_new_n1028__));
  and1  g450(.dina(new_new_n1028__), .dinb(new_new_n1027__), .dout(new_new_n1029__));
  or1   g451(.dina(new_new_n994__), .dinb(new_new_n989__), .dout(new_new_n1030__));
  or1   g452(.dina(new_new_n1030__), .dinb(new_new_n999__), .dout(new_new_n1031__));
  or1   g453(.dina(new_new_n1031__), .dinb(new_new_n1004__), .dout(new_new_n1032__));
  or1   g454(.dina(new_new_n1032__), .dinb(new_new_n1009__), .dout(new_new_n1033__));
  or1   g455(.dina(new_new_n1033__), .dinb(new_new_n1014__), .dout(new_new_n1034__));
  or1   g456(.dina(new_new_n1034__), .dinb(new_new_n1019__), .dout(new_new_n1035__));
  or1   g457(.dina(new_new_n1035__), .dinb(new_new_n1024__), .dout(new_new_n1036__));
  or1   g458(.dina(new_new_n1036__), .dinb(new_new_n1029__), .dout(new_new_n1037__));
  and1  g459(.dina(new_new_n1390__), .dinb(new_new_n1352__), .dout(new_new_n1038__));
  and1  g460(.dina(new_new_n1398__), .dinb(new_new_n1354__), .dout(new_new_n1039__));
  or1   g461(.dina(new_new_n1039__), .dinb(new_new_n1038__), .dout(new_new_n1040__));
  and1  g462(.dina(new_new_n1390__), .dinb(new_new_n1351__), .dout(new_new_n1041__));
  and1  g463(.dina(new_new_n1398__), .dinb(new_new_n1353__), .dout(new_new_n1042__));
  or1   g464(.dina(new_new_n1042__), .dinb(new_new_n1041__), .dout(new_new_n1043__));
  and1  g465(.dina(new_new_n1389__), .dinb(new_new_n1355__), .dout(new_new_n1044__));
  and1  g466(.dina(new_new_n1399__), .dinb(new_new_n1356__), .dout(new_new_n1045__));
  or1   g467(.dina(new_new_n1045__), .dinb(new_new_n1044__), .dout(new_new_n1046__));
  and1  g468(.dina(new_new_n1391__), .dinb(new_new_n1357__), .dout(new_new_n1047__));
  and1  g469(.dina(new_new_n1399__), .dinb(new_new_n1358__), .dout(new_new_n1048__));
  or1   g470(.dina(new_new_n1048__), .dinb(new_new_n1047__), .dout(new_new_n1049__));
  and1  g471(.dina(new_new_n1391__), .dinb(new_new_n1359__), .dout(new_new_n1050__));
  and1  g472(.dina(new_new_n1400__), .dinb(new_new_n1360__), .dout(new_new_n1051__));
  or1   g473(.dina(new_new_n1051__), .dinb(new_new_n1050__), .dout(new_new_n1052__));
  and1  g474(.dina(new_new_n1393__), .dinb(new_new_n1361__), .dout(new_new_n1053__));
  and1  g475(.dina(new_new_n1400__), .dinb(new_new_n1362__), .dout(new_new_n1054__));
  or1   g476(.dina(new_new_n1054__), .dinb(new_new_n1053__), .dout(new_new_n1055__));
  and1  g477(.dina(new_new_n1393__), .dinb(new_new_n1363__), .dout(new_new_n1056__));
  and1  g478(.dina(new_new_n1402__), .dinb(new_new_n1364__), .dout(new_new_n1057__));
  or1   g479(.dina(new_new_n1057__), .dinb(new_new_n1056__), .dout(new_new_n1058__));
  and1  g480(.dina(new_new_n1394__), .dinb(new_new_n1365__), .dout(new_new_n1059__));
  and1  g481(.dina(new_new_n1402__), .dinb(new_new_n1366__), .dout(new_new_n1060__));
  or1   g482(.dina(new_new_n1060__), .dinb(new_new_n1059__), .dout(new_new_n1061__));
  and1  g483(.dina(new_new_n1394__), .dinb(new_new_n1367__), .dout(new_new_n1062__));
  and1  g484(.dina(new_new_n1403__), .dinb(new_new_n1368__), .dout(new_new_n1063__));
  or1   g485(.dina(new_new_n1063__), .dinb(new_new_n1062__), .dout(new_new_n1064__));
  and1  g486(.dina(new_new_n1405__), .dinb(new_new_n503__), .dout(new_new_n1065__));
  and1  g487(.dina(new_new_n1065__), .dinb(new_new_n1406__), .dout(new_new_n1066__));
  and1  g488(.dina(new_new_n1408__), .dinb(new_new_n523__), .dout(new_new_n1067__));
  and1  g489(.dina(new_new_n1067__), .dinb(new_new_n1409__), .dout(new_new_n1068__));
  and1  g490(.dina(new_new_n1411__), .dinb(new_new_n543__), .dout(new_new_n1069__));
  and1  g491(.dina(new_new_n1069__), .dinb(new_new_n1412__), .dout(new_new_n1070__));
  and1  g492(.dina(new_new_n1414__), .dinb(new_new_n563__), .dout(new_new_n1071__));
  and1  g493(.dina(new_new_n1071__), .dinb(new_new_n1415__), .dout(new_new_n1072__));
  and1  g494(.dina(new_new_n1417__), .dinb(new_new_n583__), .dout(new_new_n1073__));
  and1  g495(.dina(new_new_n1073__), .dinb(new_new_n1418__), .dout(new_new_n1074__));
  and1  g496(.dina(new_new_n1420__), .dinb(new_new_n603__), .dout(new_new_n1075__));
  and1  g497(.dina(new_new_n1075__), .dinb(new_new_n1421__), .dout(new_new_n1076__));
  and1  g498(.dina(new_new_n1423__), .dinb(new_new_n623__), .dout(new_new_n1077__));
  and1  g499(.dina(new_new_n1077__), .dinb(new_new_n1424__), .dout(new_new_n1078__));
  and1  g500(.dina(new_new_n1426__), .dinb(new_new_n643__), .dout(new_new_n1079__));
  and1  g501(.dina(new_new_n1079__), .dinb(new_new_n1427__), .dout(new_new_n1080__));
  and1  g502(.dina(new_new_n1429__), .dinb(new_new_n663__), .dout(new_new_n1081__));
  and1  g503(.dina(new_new_n1081__), .dinb(new_new_n1430__), .dout(new_new_n1082__));
  and1  g504(.dina(new_new_n1405__), .dinb(new_new_n513__), .dout(new_new_n1083__));
  and1  g505(.dina(new_new_n1408__), .dinb(new_new_n533__), .dout(new_new_n1084__));
  and1  g506(.dina(new_new_n1411__), .dinb(new_new_n553__), .dout(new_new_n1085__));
  and1  g507(.dina(new_new_n1414__), .dinb(new_new_n573__), .dout(new_new_n1086__));
  and1  g508(.dina(new_new_n1417__), .dinb(new_new_n593__), .dout(new_new_n1087__));
  and1  g509(.dina(new_new_n1420__), .dinb(new_new_n613__), .dout(new_new_n1088__));
  and1  g510(.dina(new_new_n1423__), .dinb(new_new_n633__), .dout(new_new_n1089__));
  and1  g511(.dina(new_new_n1426__), .dinb(new_new_n653__), .dout(new_new_n1090__));
  and1  g512(.dina(new_new_n1429__), .dinb(new_new_n669__), .dout(new_new_n1091__));
  or1   g513(.dina(new_new_n1431__), .dinb(new_new_n1432__), .dout(new_new_n1092__));
  or1   g514(.dina(new_new_n1092__), .dinb(new_new_n1433__), .dout(new_new_n1093__));
  or1   g515(.dina(new_new_n1093__), .dinb(new_new_n1434__), .dout(new_new_n1094__));
  or1   g516(.dina(new_new_n1094__), .dinb(new_new_n1435__), .dout(new_new_n1095__));
  or1   g517(.dina(new_new_n1095__), .dinb(new_new_n1436__), .dout(new_new_n1096__));
  or1   g518(.dina(new_new_n1096__), .dinb(new_new_n1437__), .dout(new_new_n1097__));
  or1   g519(.dina(new_new_n1097__), .dinb(new_new_n1438__), .dout(new_new_n1098__));
  or1   g520(.dina(new_new_n1098__), .dinb(new_new_n1439__), .dout(new_new_n1099__));
  and1  g521(.dina(new_new_n1440__), .dinb(new_new_n493__), .dout(new_new_n1100__));
  and1  g522(.dina(new_new_n1441__), .dinb(new_new_n507__), .dout(new_new_n1101__));
  and1  g523(.dina(new_new_n1442__), .dinb(new_new_n527__), .dout(new_new_n1102__));
  and1  g524(.dina(new_new_n1443__), .dinb(new_new_n547__), .dout(new_new_n1103__));
  and1  g525(.dina(new_new_n1444__), .dinb(new_new_n567__), .dout(new_new_n1104__));
  and1  g526(.dina(new_new_n1445__), .dinb(new_new_n587__), .dout(new_new_n1105__));
  and1  g527(.dina(new_new_n1446__), .dinb(new_new_n607__), .dout(new_new_n1106__));
  and1  g528(.dina(new_new_n1447__), .dinb(new_new_n627__), .dout(new_new_n1107__));
  and1  g529(.dina(new_new_n1448__), .dinb(new_new_n647__), .dout(new_new_n1108__));
  buf1  g530(.din(new_new_n672__), .dout(G426));
  buf1  g531(.din(new_new_n674__), .dout(G427));
  buf1  g532(.din(new_new_n732__), .dout(G428));
  not1  g533(.din(new_new_n953__), .dout(G429));
  not1  g534(.din(new_new_n956__), .dout(G430));
  not1  g535(.din(new_new_n963__), .dout(G431));
  not1  g536(.din(new_new_n968__), .dout(G432));
  buf1  g537(.din(new_new_n420__), .dout(n2012));
  buf1  g538(.din(new_new_n676__), .dout(n2015));
  buf1  g539(.din(new_new_n422__), .dout(n2018));
  buf1  g540(.din(new_new_n694__), .dout(n2021));
  buf1  g541(.din(new_new_n424__), .dout(n2024));
  buf1  g542(.din(new_new_n500__), .dout(n2027));
  buf1  g543(.din(new_new_n714__), .dout(n2030));
  buf1  g544(.din(new_new_n426__), .dout(n2033));
  buf1  g545(.din(new_new_n678__), .dout(n2036));
  buf1  g546(.din(new_new_n428__), .dout(n2039));
  buf1  g547(.din(new_new_n510__), .dout(n2042));
  buf1  g548(.din(new_new_n752__), .dout(n2045));
  buf1  g549(.din(new_new_n430__), .dout(n2048));
  buf1  g550(.din(new_new_n696__), .dout(n2051));
  buf1  g551(.din(new_new_n432__), .dout(n2054));
  buf1  g552(.din(new_new_n520__), .dout(n2057));
  buf1  g553(.din(new_new_n716__), .dout(n2060));
  buf1  g554(.din(new_new_n434__), .dout(n2063));
  buf1  g555(.din(new_new_n680__), .dout(n2066));
  buf1  g556(.din(new_new_n436__), .dout(n2069));
  buf1  g557(.din(new_new_n530__), .dout(n2072));
  buf1  g558(.din(new_new_n754__), .dout(n2075));
  buf1  g559(.din(new_new_n438__), .dout(n2078));
  buf1  g560(.din(new_new_n698__), .dout(n2081));
  buf1  g561(.din(new_new_n440__), .dout(n2084));
  buf1  g562(.din(new_new_n540__), .dout(n2087));
  buf1  g563(.din(new_new_n718__), .dout(n2090));
  buf1  g564(.din(new_new_n442__), .dout(n2093));
  buf1  g565(.din(new_new_n682__), .dout(n2096));
  buf1  g566(.din(new_new_n444__), .dout(n2099));
  buf1  g567(.din(new_new_n550__), .dout(n2102));
  buf1  g568(.din(new_new_n756__), .dout(n2105));
  buf1  g569(.din(new_new_n446__), .dout(n2108));
  buf1  g570(.din(new_new_n700__), .dout(n2111));
  buf1  g571(.din(new_new_n448__), .dout(n2114));
  buf1  g572(.din(new_new_n560__), .dout(n2117));
  buf1  g573(.din(new_new_n720__), .dout(n2120));
  buf1  g574(.din(new_new_n450__), .dout(n2123));
  buf1  g575(.din(new_new_n684__), .dout(n2126));
  buf1  g576(.din(new_new_n452__), .dout(n2129));
  buf1  g577(.din(new_new_n570__), .dout(n2132));
  buf1  g578(.din(new_new_n758__), .dout(n2135));
  buf1  g579(.din(new_new_n454__), .dout(n2138));
  buf1  g580(.din(new_new_n702__), .dout(n2141));
  buf1  g581(.din(new_new_n456__), .dout(n2144));
  buf1  g582(.din(new_new_n580__), .dout(n2147));
  buf1  g583(.din(new_new_n722__), .dout(n2150));
  buf1  g584(.din(new_new_n458__), .dout(n2153));
  buf1  g585(.din(new_new_n686__), .dout(n2156));
  buf1  g586(.din(new_new_n460__), .dout(n2159));
  buf1  g587(.din(new_new_n590__), .dout(n2162));
  buf1  g588(.din(new_new_n760__), .dout(n2165));
  buf1  g589(.din(new_new_n462__), .dout(n2168));
  buf1  g590(.din(new_new_n704__), .dout(n2171));
  buf1  g591(.din(new_new_n464__), .dout(n2174));
  buf1  g592(.din(new_new_n600__), .dout(n2177));
  buf1  g593(.din(new_new_n724__), .dout(n2180));
  buf1  g594(.din(new_new_n466__), .dout(n2183));
  buf1  g595(.din(new_new_n688__), .dout(n2186));
  buf1  g596(.din(new_new_n468__), .dout(n2189));
  buf1  g597(.din(new_new_n610__), .dout(n2192));
  buf1  g598(.din(new_new_n762__), .dout(n2195));
  buf1  g599(.din(new_new_n470__), .dout(n2198));
  buf1  g600(.din(new_new_n706__), .dout(n2201));
  buf1  g601(.din(new_new_n472__), .dout(n2204));
  buf1  g602(.din(new_new_n620__), .dout(n2207));
  buf1  g603(.din(new_new_n726__), .dout(n2210));
  buf1  g604(.din(new_new_n474__), .dout(n2213));
  buf1  g605(.din(new_new_n690__), .dout(n2216));
  buf1  g606(.din(new_new_n476__), .dout(n2219));
  buf1  g607(.din(new_new_n630__), .dout(n2222));
  buf1  g608(.din(new_new_n764__), .dout(n2225));
  buf1  g609(.din(new_new_n478__), .dout(n2228));
  buf1  g610(.din(new_new_n708__), .dout(n2231));
  buf1  g611(.din(new_new_n480__), .dout(n2234));
  buf1  g612(.din(new_new_n640__), .dout(n2237));
  buf1  g613(.din(new_new_n728__), .dout(n2240));
  buf1  g614(.din(new_new_n482__), .dout(n2243));
  buf1  g615(.din(new_new_n692__), .dout(n2246));
  buf1  g616(.din(new_new_n484__), .dout(n2249));
  buf1  g617(.din(new_new_n650__), .dout(n2252));
  buf1  g618(.din(new_new_n766__), .dout(n2255));
  buf1  g619(.din(new_new_n486__), .dout(n2258));
  buf1  g620(.din(new_new_n710__), .dout(n2261));
  buf1  g621(.din(new_new_n488__), .dout(n2264));
  buf1  g622(.din(new_new_n660__), .dout(n2267));
  buf1  g623(.din(new_new_n730__), .dout(n2270));
  buf1  g624(.din(new_new_n490__), .dout(n2273));
  buf1  g625(.din(new_new_n666__), .dout(n2276));
  buf1  g626(.din(new_new_n768__), .dout(n2279));
  buf1  g627(.din(new_new_n1449__), .dout(n2282));
  buf1  g628(.din(new_new_n1386__), .dout(n2285));
  buf1  g629(.din(new_new_n794__), .dout(n2288));
  buf1  g630(.din(new_new_n796__), .dout(n2291));
  buf1  g631(.din(new_new_n798__), .dout(n2294));
  buf1  g632(.din(new_new_n800__), .dout(n2297));
  buf1  g633(.din(new_new_n802__), .dout(n2300));
  buf1  g634(.din(new_new_n804__), .dout(n2303));
  buf1  g635(.din(new_new_n806__), .dout(n2306));
  buf1  g636(.din(new_new_n808__), .dout(n2309));
  buf1  g637(.din(new_new_n810__), .dout(n2312));
  buf1  g638(.din(new_new_n1404__), .dout(n2315));
  buf1  g639(.din(new_new_n1407__), .dout(n2318));
  buf1  g640(.din(new_new_n1410__), .dout(n2321));
  buf1  g641(.din(new_new_n1413__), .dout(n2324));
  buf1  g642(.din(new_new_n1416__), .dout(n2327));
  buf1  g643(.din(new_new_n1419__), .dout(n2330));
  buf1  g644(.din(new_new_n1422__), .dout(n2333));
  buf1  g645(.din(new_new_n1425__), .dout(n2336));
  buf1  g646(.din(new_new_n1428__), .dout(n2339));
  buf1  g647(.din(new_new_n1403__), .dout(n2342));
  buf1  g648(.din(new_new_n502__), .dout(n2345));
  buf1  g649(.din(new_new_n522__), .dout(n2348));
  buf1  g650(.din(new_new_n542__), .dout(n2351));
  buf1  g651(.din(new_new_n562__), .dout(n2354));
  buf1  g652(.din(new_new_n582__), .dout(n2357));
  buf1  g653(.din(new_new_n602__), .dout(n2360));
  buf1  g654(.din(new_new_n622__), .dout(n2363));
  buf1  g655(.din(new_new_n642__), .dout(n2366));
  buf1  g656(.din(new_new_n662__), .dout(n2369));
  buf1  g657(.din(new_new_n1450__), .dout(n2372));
  not1  g658(.din(new_new_n1406__), .dout(n2375));
  not1  g659(.din(new_new_n1409__), .dout(n2378));
  not1  g660(.din(new_new_n1412__), .dout(n2381));
  not1  g661(.din(new_new_n1415__), .dout(n2384));
  not1  g662(.din(new_new_n1418__), .dout(n2387));
  not1  g663(.din(new_new_n1421__), .dout(n2390));
  not1  g664(.din(new_new_n1424__), .dout(n2393));
  not1  g665(.din(new_new_n1427__), .dout(n2396));
  not1  g666(.din(new_new_n1430__), .dout(n2399));
  buf1  g667(.din(new_new_n512__), .dout(n2402));
  buf1  g668(.din(new_new_n532__), .dout(n2405));
  buf1  g669(.din(new_new_n552__), .dout(n2408));
  buf1  g670(.din(new_new_n572__), .dout(n2411));
  buf1  g671(.din(new_new_n592__), .dout(n2414));
  buf1  g672(.din(new_new_n612__), .dout(n2417));
  buf1  g673(.din(new_new_n632__), .dout(n2420));
  buf1  g674(.din(new_new_n652__), .dout(n2423));
  buf1  g675(.din(new_new_n668__), .dout(n2426));
  buf1  g676(.din(n2282), .dout(n2429));
  buf1  g677(.din(n2285), .dout(n2432));
  buf1  g678(.din(n2372), .dout(n2435));
  buf1  g679(.din(new_new_n1432__), .dout(n2438));
  buf1  g680(.din(new_new_n1431__), .dout(n2441));
  buf1  g681(.din(new_new_n1433__), .dout(n2444));
  buf1  g682(.din(new_new_n1434__), .dout(n2447));
  buf1  g683(.din(new_new_n1435__), .dout(n2450));
  buf1  g684(.din(new_new_n1436__), .dout(n2453));
  buf1  g685(.din(new_new_n1437__), .dout(n2456));
  buf1  g686(.din(new_new_n1438__), .dout(n2459));
  buf1  g687(.din(new_new_n1439__), .dout(n2462));
  buf1  g688(.din(new_new_n492__), .dout(n2465));
  buf1  g689(.din(new_new_n506__), .dout(n2468));
  buf1  g690(.din(new_new_n526__), .dout(n2471));
  buf1  g691(.din(new_new_n546__), .dout(n2474));
  buf1  g692(.din(new_new_n566__), .dout(n2477));
  buf1  g693(.din(new_new_n586__), .dout(n2480));
  buf1  g694(.din(new_new_n606__), .dout(n2483));
  buf1  g695(.din(new_new_n626__), .dout(n2486));
  buf1  g696(.din(new_new_n646__), .dout(n2489));
  buf1  g697(.din(new_new_n1083__), .dout(n2492));
  buf1  g698(.din(new_new_n1084__), .dout(n2495));
  buf1  g699(.din(new_new_n1085__), .dout(n2498));
  buf1  g700(.din(new_new_n1086__), .dout(n2501));
  buf1  g701(.din(new_new_n1087__), .dout(n2504));
  buf1  g702(.din(new_new_n1088__), .dout(n2507));
  buf1  g703(.din(new_new_n1089__), .dout(n2510));
  buf1  g704(.din(new_new_n1090__), .dout(n2513));
  buf1  g705(.din(new_new_n1091__), .dout(n2516));
  buf1  g706(.din(new_new_n1440__), .dout(n2519));
  buf1  g707(.din(new_new_n1441__), .dout(n2522));
  buf1  g708(.din(new_new_n1442__), .dout(n2525));
  buf1  g709(.din(new_new_n1443__), .dout(n2528));
  buf1  g710(.din(new_new_n1444__), .dout(n2531));
  buf1  g711(.din(new_new_n1445__), .dout(n2534));
  buf1  g712(.din(new_new_n1446__), .dout(n2537));
  buf1  g713(.din(new_new_n1447__), .dout(n2540));
  buf1  g714(.din(new_new_n1448__), .dout(n2543));
  buf1  g715(.din(new_new_n1099__), .dout(n2546));
  buf1  g716(.din(new_new_n1100__), .dout(n2549));
  buf1  g717(.din(new_new_n1101__), .dout(n2552));
  buf1  g718(.din(new_new_n1102__), .dout(n2555));
  buf1  g719(.din(new_new_n1103__), .dout(n2558));
  buf1  g720(.din(new_new_n1104__), .dout(n2561));
  buf1  g721(.din(new_new_n1105__), .dout(n2564));
  buf1  g722(.din(new_new_n1106__), .dout(n2567));
  buf1  g723(.din(new_new_n1107__), .dout(n2570));
  buf1  g724(.din(new_new_n1108__), .dout(n2573));
  buf1  g725(.din(new_new_n771__), .dout(new_new_n1304__));
  buf1  g726(.din(new_new_n1304__), .dout(new_new_n1305__));
  buf1  g727(.din(new_new_n1305__), .dout(new_new_n1306__));
  buf1  g728(.din(new_new_n1304__), .dout(new_new_n1307__));
  buf1  g729(.din(new_new_n773__), .dout(new_new_n1308__));
  buf1  g730(.din(new_new_n1308__), .dout(new_new_n1309__));
  buf1  g731(.din(new_new_n1309__), .dout(new_new_n1310__));
  buf1  g732(.din(new_new_n1308__), .dout(new_new_n1311__));
  buf1  g733(.din(new_new_n775__), .dout(new_new_n1312__));
  buf1  g734(.din(new_new_n1312__), .dout(new_new_n1313__));
  buf1  g735(.din(new_new_n1313__), .dout(new_new_n1314__));
  buf1  g736(.din(new_new_n1312__), .dout(new_new_n1315__));
  buf1  g737(.din(new_new_n770__), .dout(new_new_n1316__));
  buf1  g738(.din(new_new_n1316__), .dout(new_new_n1317__));
  buf1  g739(.din(new_new_n1317__), .dout(new_new_n1318__));
  buf1  g740(.din(new_new_n1317__), .dout(new_new_n1319__));
  buf1  g741(.din(new_new_n1316__), .dout(new_new_n1320__));
  buf1  g742(.din(new_new_n1320__), .dout(new_new_n1321__));
  buf1  g743(.din(new_new_n1320__), .dout(new_new_n1322__));
  buf1  g744(.din(new_new_n772__), .dout(new_new_n1323__));
  buf1  g745(.din(new_new_n1323__), .dout(new_new_n1324__));
  buf1  g746(.din(new_new_n1324__), .dout(new_new_n1325__));
  buf1  g747(.din(new_new_n1324__), .dout(new_new_n1326__));
  buf1  g748(.din(new_new_n1323__), .dout(new_new_n1327__));
  buf1  g749(.din(new_new_n1327__), .dout(new_new_n1328__));
  buf1  g750(.din(new_new_n1327__), .dout(new_new_n1329__));
  buf1  g751(.din(new_new_n774__), .dout(new_new_n1330__));
  buf1  g752(.din(new_new_n1330__), .dout(new_new_n1331__));
  buf1  g753(.din(new_new_n1331__), .dout(new_new_n1332__));
  buf1  g754(.din(new_new_n1331__), .dout(new_new_n1333__));
  buf1  g755(.din(new_new_n1330__), .dout(new_new_n1334__));
  buf1  g756(.din(new_new_n1334__), .dout(new_new_n1335__));
  buf1  g757(.din(new_new_n1334__), .dout(new_new_n1336__));
  buf1  g758(.din(new_new_n879__), .dout(new_new_n1337__));
  buf1  g759(.din(new_new_n946__), .dout(new_new_n1338__));
  buf1  g760(.din(new_new_n1338__), .dout(new_new_n1339__));
  buf1  g761(.din(new_new_n903__), .dout(new_new_n1340__));
  buf1  g762(.din(new_new_n915__), .dout(new_new_n1341__));
  buf1  g763(.din(new_new_n921__), .dout(new_new_n1342__));
  buf1  g764(.din(new_new_n933__), .dout(new_new_n1343__));
  buf1  g765(.din(new_new_n939__), .dout(new_new_n1344__));
  buf1  g766(.din(new_new_n890__), .dout(new_new_n1345__));
  buf1  g767(.din(new_new_n954__), .dout(new_new_n1346__));
  buf1  g768(.din(new_new_n902__), .dout(new_new_n1347__));
  buf1  g769(.din(new_new_n957__), .dout(new_new_n1348__));
  buf1  g770(.din(new_new_n914__), .dout(new_new_n1349__));
  buf1  g771(.din(new_new_n959__), .dout(new_new_n1350__));
  buf1  g772(.din(new_new_n853__), .dout(new_new_n1351__));
  buf1  g773(.din(new_new_n851__), .dout(new_new_n1352__));
  buf1  g774(.din(new_new_n852__), .dout(new_new_n1353__));
  buf1  g775(.din(new_new_n850__), .dout(new_new_n1354__));
  buf1  g776(.din(new_new_n855__), .dout(new_new_n1355__));
  buf1  g777(.din(new_new_n854__), .dout(new_new_n1356__));
  buf1  g778(.din(new_new_n857__), .dout(new_new_n1357__));
  buf1  g779(.din(new_new_n856__), .dout(new_new_n1358__));
  buf1  g780(.din(new_new_n859__), .dout(new_new_n1359__));
  buf1  g781(.din(new_new_n858__), .dout(new_new_n1360__));
  buf1  g782(.din(new_new_n861__), .dout(new_new_n1361__));
  buf1  g783(.din(new_new_n860__), .dout(new_new_n1362__));
  buf1  g784(.din(new_new_n863__), .dout(new_new_n1363__));
  buf1  g785(.din(new_new_n862__), .dout(new_new_n1364__));
  buf1  g786(.din(new_new_n865__), .dout(new_new_n1365__));
  buf1  g787(.din(new_new_n864__), .dout(new_new_n1366__));
  buf1  g788(.din(new_new_n867__), .dout(new_new_n1367__));
  buf1  g789(.din(new_new_n866__), .dout(new_new_n1368__));
  buf1  g790(.din(new_new_n849__), .dout(new_new_n1369__));
  buf1  g791(.din(new_new_n1369__), .dout(new_new_n1370__));
  buf1  g792(.din(new_new_n1370__), .dout(new_new_n1371__));
  buf1  g793(.din(new_new_n1371__), .dout(new_new_n1372__));
  buf1  g794(.din(new_new_n1370__), .dout(new_new_n1373__));
  buf1  g795(.din(new_new_n1369__), .dout(new_new_n1374__));
  buf1  g796(.din(new_new_n1374__), .dout(new_new_n1375__));
  buf1  g797(.din(new_new_n1374__), .dout(new_new_n1376__));
  buf1  g798(.din(new_new_n848__), .dout(new_new_n1377__));
  buf1  g799(.din(new_new_n1377__), .dout(new_new_n1378__));
  buf1  g800(.din(new_new_n1378__), .dout(new_new_n1379__));
  buf1  g801(.din(new_new_n1379__), .dout(new_new_n1380__));
  buf1  g802(.din(new_new_n1379__), .dout(new_new_n1381__));
  buf1  g803(.din(new_new_n1378__), .dout(new_new_n1382__));
  buf1  g804(.din(new_new_n1382__), .dout(new_new_n1383__));
  buf1  g805(.din(new_new_n1377__), .dout(new_new_n1384__));
  buf1  g806(.din(new_new_n1384__), .dout(new_new_n1385__));
  buf1  g807(.din(new_new_n1384__), .dout(new_new_n1386__));
  buf1  g808(.din(new_new_n983__), .dout(new_new_n1387__));
  buf1  g809(.din(new_new_n1387__), .dout(new_new_n1388__));
  buf1  g810(.din(new_new_n1388__), .dout(new_new_n1389__));
  buf1  g811(.din(new_new_n1389__), .dout(new_new_n1390__));
  buf1  g812(.din(new_new_n1388__), .dout(new_new_n1391__));
  buf1  g813(.din(new_new_n1387__), .dout(new_new_n1392__));
  buf1  g814(.din(new_new_n1392__), .dout(new_new_n1393__));
  buf1  g815(.din(new_new_n1392__), .dout(new_new_n1394__));
  buf1  g816(.din(new_new_n984__), .dout(new_new_n1395__));
  buf1  g817(.din(new_new_n1395__), .dout(new_new_n1396__));
  buf1  g818(.din(new_new_n1396__), .dout(new_new_n1397__));
  buf1  g819(.din(new_new_n1397__), .dout(new_new_n1398__));
  buf1  g820(.din(new_new_n1397__), .dout(new_new_n1399__));
  buf1  g821(.din(new_new_n1396__), .dout(new_new_n1400__));
  buf1  g822(.din(new_new_n1395__), .dout(new_new_n1401__));
  buf1  g823(.din(new_new_n1401__), .dout(new_new_n1402__));
  buf1  g824(.din(new_new_n1401__), .dout(new_new_n1403__));
  buf1  g825(.din(new_new_n830__), .dout(new_new_n1404__));
  buf1  g826(.din(new_new_n1404__), .dout(new_new_n1405__));
  buf1  g827(.din(new_new_n1040__), .dout(new_new_n1406__));
  buf1  g828(.din(new_new_n832__), .dout(new_new_n1407__));
  buf1  g829(.din(new_new_n1407__), .dout(new_new_n1408__));
  buf1  g830(.din(new_new_n1043__), .dout(new_new_n1409__));
  buf1  g831(.din(new_new_n834__), .dout(new_new_n1410__));
  buf1  g832(.din(new_new_n1410__), .dout(new_new_n1411__));
  buf1  g833(.din(new_new_n1046__), .dout(new_new_n1412__));
  buf1  g834(.din(new_new_n836__), .dout(new_new_n1413__));
  buf1  g835(.din(new_new_n1413__), .dout(new_new_n1414__));
  buf1  g836(.din(new_new_n1049__), .dout(new_new_n1415__));
  buf1  g837(.din(new_new_n838__), .dout(new_new_n1416__));
  buf1  g838(.din(new_new_n1416__), .dout(new_new_n1417__));
  buf1  g839(.din(new_new_n1052__), .dout(new_new_n1418__));
  buf1  g840(.din(new_new_n840__), .dout(new_new_n1419__));
  buf1  g841(.din(new_new_n1419__), .dout(new_new_n1420__));
  buf1  g842(.din(new_new_n1055__), .dout(new_new_n1421__));
  buf1  g843(.din(new_new_n842__), .dout(new_new_n1422__));
  buf1  g844(.din(new_new_n1422__), .dout(new_new_n1423__));
  buf1  g845(.din(new_new_n1058__), .dout(new_new_n1424__));
  buf1  g846(.din(new_new_n844__), .dout(new_new_n1425__));
  buf1  g847(.din(new_new_n1425__), .dout(new_new_n1426__));
  buf1  g848(.din(new_new_n1061__), .dout(new_new_n1427__));
  buf1  g849(.din(new_new_n846__), .dout(new_new_n1428__));
  buf1  g850(.din(new_new_n1428__), .dout(new_new_n1429__));
  buf1  g851(.din(new_new_n1064__), .dout(new_new_n1430__));
  buf1  g852(.din(new_new_n1068__), .dout(new_new_n1431__));
  buf1  g853(.din(new_new_n1066__), .dout(new_new_n1432__));
  buf1  g854(.din(new_new_n1070__), .dout(new_new_n1433__));
  buf1  g855(.din(new_new_n1072__), .dout(new_new_n1434__));
  buf1  g856(.din(new_new_n1074__), .dout(new_new_n1435__));
  buf1  g857(.din(new_new_n1076__), .dout(new_new_n1436__));
  buf1  g858(.din(new_new_n1078__), .dout(new_new_n1437__));
  buf1  g859(.din(new_new_n1080__), .dout(new_new_n1438__));
  buf1  g860(.din(new_new_n1082__), .dout(new_new_n1439__));
  buf1  g861(.din(new_new_n496__), .dout(new_new_n1440__));
  buf1  g862(.din(new_new_n516__), .dout(new_new_n1441__));
  buf1  g863(.din(new_new_n536__), .dout(new_new_n1442__));
  buf1  g864(.din(new_new_n556__), .dout(new_new_n1443__));
  buf1  g865(.din(new_new_n576__), .dout(new_new_n1444__));
  buf1  g866(.din(new_new_n596__), .dout(new_new_n1445__));
  buf1  g867(.din(new_new_n616__), .dout(new_new_n1446__));
  buf1  g868(.din(new_new_n636__), .dout(new_new_n1447__));
  buf1  g869(.din(new_new_n656__), .dout(new_new_n1448__));
  buf1  g870(.din(new_new_n712__), .dout(new_new_n1449__));
  buf1  g871(.din(new_new_n1037__), .dout(new_new_n1450__));
  always @ (posedge clock) begin
    n205_lo <= n2012;
    n214_lo <= n2015;
    n217_lo <= n2018;
    n226_lo <= n2021;
    n229_lo <= n2024;
    n232_lo <= n2027;
    n238_lo <= n2030;
    n241_lo <= n2033;
    n250_lo <= n2036;
    n253_lo <= n2039;
    n256_lo <= n2042;
    n262_lo <= n2045;
    n265_lo <= n2048;
    n274_lo <= n2051;
    n277_lo <= n2054;
    n280_lo <= n2057;
    n286_lo <= n2060;
    n289_lo <= n2063;
    n298_lo <= n2066;
    n301_lo <= n2069;
    n304_lo <= n2072;
    n310_lo <= n2075;
    n313_lo <= n2078;
    n322_lo <= n2081;
    n325_lo <= n2084;
    n328_lo <= n2087;
    n334_lo <= n2090;
    n337_lo <= n2093;
    n346_lo <= n2096;
    n349_lo <= n2099;
    n352_lo <= n2102;
    n358_lo <= n2105;
    n361_lo <= n2108;
    n370_lo <= n2111;
    n373_lo <= n2114;
    n376_lo <= n2117;
    n382_lo <= n2120;
    n385_lo <= n2123;
    n394_lo <= n2126;
    n397_lo <= n2129;
    n400_lo <= n2132;
    n406_lo <= n2135;
    n409_lo <= n2138;
    n418_lo <= n2141;
    n421_lo <= n2144;
    n424_lo <= n2147;
    n430_lo <= n2150;
    n433_lo <= n2153;
    n442_lo <= n2156;
    n445_lo <= n2159;
    n448_lo <= n2162;
    n454_lo <= n2165;
    n457_lo <= n2168;
    n466_lo <= n2171;
    n469_lo <= n2174;
    n472_lo <= n2177;
    n478_lo <= n2180;
    n481_lo <= n2183;
    n490_lo <= n2186;
    n493_lo <= n2189;
    n496_lo <= n2192;
    n502_lo <= n2195;
    n505_lo <= n2198;
    n514_lo <= n2201;
    n517_lo <= n2204;
    n520_lo <= n2207;
    n526_lo <= n2210;
    n529_lo <= n2213;
    n538_lo <= n2216;
    n541_lo <= n2219;
    n544_lo <= n2222;
    n550_lo <= n2225;
    n553_lo <= n2228;
    n562_lo <= n2231;
    n565_lo <= n2234;
    n568_lo <= n2237;
    n574_lo <= n2240;
    n577_lo <= n2243;
    n586_lo <= n2246;
    n589_lo <= n2249;
    n592_lo <= n2252;
    n598_lo <= n2255;
    n601_lo <= n2258;
    n610_lo <= n2261;
    n613_lo <= n2264;
    n616_lo <= n2267;
    n622_lo <= n2270;
    n625_lo <= n2273;
    n628_lo <= n2276;
    n634_lo <= n2279;
    n316_inv <= n2282;
    n319_inv <= n2285;
    n997_o2 <= n2288;
    n998_o2 <= n2291;
    n999_o2 <= n2294;
    n1000_o2 <= n2297;
    n1001_o2 <= n2300;
    n1002_o2 <= n2303;
    n1003_o2 <= n2306;
    n1004_o2 <= n2309;
    n1005_o2 <= n2312;
    n1015_o2 <= n2315;
    n1016_o2 <= n2318;
    n1017_o2 <= n2321;
    n1018_o2 <= n2324;
    n1019_o2 <= n2327;
    n1020_o2 <= n2330;
    n1021_o2 <= n2333;
    n1022_o2 <= n2336;
    n1023_o2 <= n2339;
    n376_1_inv <= n2342;
    n235_lo_buf_o2 <= n2345;
    n283_lo_buf_o2 <= n2348;
    n331_lo_buf_o2 <= n2351;
    n379_lo_buf_o2 <= n2354;
    n427_lo_buf_o2 <= n2357;
    n475_lo_buf_o2 <= n2360;
    n523_lo_buf_o2 <= n2363;
    n571_lo_buf_o2 <= n2366;
    n619_lo_buf_o2 <= n2369;
    n406_1_inv <= n2372;
    G223_o2 <= n2375;
    G226_o2 <= n2378;
    G229_o2 <= n2381;
    G232_o2 <= n2384;
    G235_o2 <= n2387;
    G238_o2 <= n2390;
    G242_o2 <= n2393;
    G246_o2 <= n2396;
    G250_o2 <= n2399;
    n259_lo_buf_o2 <= n2402;
    n307_lo_buf_o2 <= n2405;
    n355_lo_buf_o2 <= n2408;
    n403_lo_buf_o2 <= n2411;
    n451_lo_buf_o2 <= n2414;
    n499_lo_buf_o2 <= n2417;
    n547_lo_buf_o2 <= n2420;
    n595_lo_buf_o2 <= n2423;
    n631_lo_buf_o2 <= n2426;
    G213_o2 <= n2429;
    G318_o2 <= n2432;
    G358_o2 <= n2435;
    G259_o2 <= n2438;
    G263_o2 <= n2441;
    G266_o2 <= n2444;
    G269_o2 <= n2447;
    G272_o2 <= n2450;
    G275_o2 <= n2453;
    G278_o2 <= n2456;
    G281_o2 <= n2459;
    G284_o2 <= n2462;
    n211_lo_buf_o2 <= n2465;
    n247_lo_buf_o2 <= n2468;
    n295_lo_buf_o2 <= n2471;
    n343_lo_buf_o2 <= n2474;
    n391_lo_buf_o2 <= n2477;
    n439_lo_buf_o2 <= n2480;
    n487_lo_buf_o2 <= n2483;
    n535_lo_buf_o2 <= n2486;
    n583_lo_buf_o2 <= n2489;
    G158_o2 <= n2492;
    G184_o2 <= n2495;
    G186_o2 <= n2498;
    G188_o2 <= n2501;
    G190_o2 <= n2504;
    G192_o2 <= n2507;
    G194_o2 <= n2510;
    G196_o2 <= n2513;
    G198_o2 <= n2516;
    n223_lo_buf_o2 <= n2519;
    n271_lo_buf_o2 <= n2522;
    n319_lo_buf_o2 <= n2525;
    n367_lo_buf_o2 <= n2528;
    n415_lo_buf_o2 <= n2531;
    n463_lo_buf_o2 <= n2534;
    n511_lo_buf_o2 <= n2537;
    n559_lo_buf_o2 <= n2540;
    n607_lo_buf_o2 <= n2543;
    n580_inv <= n2546;
    G154_o2 <= n2549;
    G159_o2 <= n2552;
    G162_o2 <= n2555;
    G165_o2 <= n2558;
    G168_o2 <= n2561;
    G171_o2 <= n2564;
    G174_o2 <= n2567;
    G177_o2 <= n2570;
    G180_o2 <= n2573;
  end
  initial begin
    n205_lo <= 1'b0;
    n214_lo <= 1'b0;
    n217_lo <= 1'b0;
    n226_lo <= 1'b0;
    n229_lo <= 1'b0;
    n232_lo <= 1'b0;
    n238_lo <= 1'b0;
    n241_lo <= 1'b0;
    n250_lo <= 1'b0;
    n253_lo <= 1'b0;
    n256_lo <= 1'b0;
    n262_lo <= 1'b0;
    n265_lo <= 1'b0;
    n274_lo <= 1'b0;
    n277_lo <= 1'b0;
    n280_lo <= 1'b0;
    n286_lo <= 1'b0;
    n289_lo <= 1'b0;
    n298_lo <= 1'b0;
    n301_lo <= 1'b0;
    n304_lo <= 1'b0;
    n310_lo <= 1'b0;
    n313_lo <= 1'b0;
    n322_lo <= 1'b0;
    n325_lo <= 1'b0;
    n328_lo <= 1'b0;
    n334_lo <= 1'b0;
    n337_lo <= 1'b0;
    n346_lo <= 1'b0;
    n349_lo <= 1'b0;
    n352_lo <= 1'b0;
    n358_lo <= 1'b0;
    n361_lo <= 1'b0;
    n370_lo <= 1'b0;
    n373_lo <= 1'b0;
    n376_lo <= 1'b0;
    n382_lo <= 1'b0;
    n385_lo <= 1'b0;
    n394_lo <= 1'b0;
    n397_lo <= 1'b0;
    n400_lo <= 1'b0;
    n406_lo <= 1'b0;
    n409_lo <= 1'b0;
    n418_lo <= 1'b0;
    n421_lo <= 1'b0;
    n424_lo <= 1'b0;
    n430_lo <= 1'b0;
    n433_lo <= 1'b0;
    n442_lo <= 1'b0;
    n445_lo <= 1'b0;
    n448_lo <= 1'b0;
    n454_lo <= 1'b0;
    n457_lo <= 1'b0;
    n466_lo <= 1'b0;
    n469_lo <= 1'b0;
    n472_lo <= 1'b0;
    n478_lo <= 1'b0;
    n481_lo <= 1'b0;
    n490_lo <= 1'b0;
    n493_lo <= 1'b0;
    n496_lo <= 1'b0;
    n502_lo <= 1'b0;
    n505_lo <= 1'b0;
    n514_lo <= 1'b0;
    n517_lo <= 1'b0;
    n520_lo <= 1'b0;
    n526_lo <= 1'b0;
    n529_lo <= 1'b0;
    n538_lo <= 1'b0;
    n541_lo <= 1'b0;
    n544_lo <= 1'b0;
    n550_lo <= 1'b0;
    n553_lo <= 1'b0;
    n562_lo <= 1'b0;
    n565_lo <= 1'b0;
    n568_lo <= 1'b0;
    n574_lo <= 1'b0;
    n577_lo <= 1'b0;
    n586_lo <= 1'b0;
    n589_lo <= 1'b0;
    n592_lo <= 1'b0;
    n598_lo <= 1'b0;
    n601_lo <= 1'b0;
    n610_lo <= 1'b0;
    n613_lo <= 1'b0;
    n616_lo <= 1'b0;
    n622_lo <= 1'b0;
    n625_lo <= 1'b0;
    n628_lo <= 1'b0;
    n634_lo <= 1'b0;
    n316_inv <= 1'b0;
    n319_inv <= 1'b0;
    n997_o2 <= 1'b0;
    n998_o2 <= 1'b0;
    n999_o2 <= 1'b0;
    n1000_o2 <= 1'b0;
    n1001_o2 <= 1'b0;
    n1002_o2 <= 1'b0;
    n1003_o2 <= 1'b0;
    n1004_o2 <= 1'b0;
    n1005_o2 <= 1'b0;
    n1015_o2 <= 1'b0;
    n1016_o2 <= 1'b0;
    n1017_o2 <= 1'b0;
    n1018_o2 <= 1'b0;
    n1019_o2 <= 1'b0;
    n1020_o2 <= 1'b0;
    n1021_o2 <= 1'b0;
    n1022_o2 <= 1'b0;
    n1023_o2 <= 1'b0;
    n376_1_inv <= 1'b0;
    n235_lo_buf_o2 <= 1'b0;
    n283_lo_buf_o2 <= 1'b0;
    n331_lo_buf_o2 <= 1'b0;
    n379_lo_buf_o2 <= 1'b0;
    n427_lo_buf_o2 <= 1'b0;
    n475_lo_buf_o2 <= 1'b0;
    n523_lo_buf_o2 <= 1'b0;
    n571_lo_buf_o2 <= 1'b0;
    n619_lo_buf_o2 <= 1'b0;
    n406_1_inv <= 1'b0;
    G223_o2 <= 1'b0;
    G226_o2 <= 1'b0;
    G229_o2 <= 1'b0;
    G232_o2 <= 1'b0;
    G235_o2 <= 1'b0;
    G238_o2 <= 1'b0;
    G242_o2 <= 1'b0;
    G246_o2 <= 1'b0;
    G250_o2 <= 1'b0;
    n259_lo_buf_o2 <= 1'b0;
    n307_lo_buf_o2 <= 1'b0;
    n355_lo_buf_o2 <= 1'b0;
    n403_lo_buf_o2 <= 1'b0;
    n451_lo_buf_o2 <= 1'b0;
    n499_lo_buf_o2 <= 1'b0;
    n547_lo_buf_o2 <= 1'b0;
    n595_lo_buf_o2 <= 1'b0;
    n631_lo_buf_o2 <= 1'b0;
    G213_o2 <= 1'b0;
    G318_o2 <= 1'b0;
    G358_o2 <= 1'b0;
    G259_o2 <= 1'b0;
    G263_o2 <= 1'b0;
    G266_o2 <= 1'b0;
    G269_o2 <= 1'b0;
    G272_o2 <= 1'b0;
    G275_o2 <= 1'b0;
    G278_o2 <= 1'b0;
    G281_o2 <= 1'b0;
    G284_o2 <= 1'b0;
    n211_lo_buf_o2 <= 1'b0;
    n247_lo_buf_o2 <= 1'b0;
    n295_lo_buf_o2 <= 1'b0;
    n343_lo_buf_o2 <= 1'b0;
    n391_lo_buf_o2 <= 1'b0;
    n439_lo_buf_o2 <= 1'b0;
    n487_lo_buf_o2 <= 1'b0;
    n535_lo_buf_o2 <= 1'b0;
    n583_lo_buf_o2 <= 1'b0;
    G158_o2 <= 1'b0;
    G184_o2 <= 1'b0;
    G186_o2 <= 1'b0;
    G188_o2 <= 1'b0;
    G190_o2 <= 1'b0;
    G192_o2 <= 1'b0;
    G194_o2 <= 1'b0;
    G196_o2 <= 1'b0;
    G198_o2 <= 1'b0;
    n223_lo_buf_o2 <= 1'b0;
    n271_lo_buf_o2 <= 1'b0;
    n319_lo_buf_o2 <= 1'b0;
    n367_lo_buf_o2 <= 1'b0;
    n415_lo_buf_o2 <= 1'b0;
    n463_lo_buf_o2 <= 1'b0;
    n511_lo_buf_o2 <= 1'b0;
    n559_lo_buf_o2 <= 1'b0;
    n607_lo_buf_o2 <= 1'b0;
    n580_inv <= 1'b0;
    G154_o2 <= 1'b0;
    G159_o2 <= 1'b0;
    G162_o2 <= 1'b0;
    G165_o2 <= 1'b0;
    G168_o2 <= 1'b0;
    G171_o2 <= 1'b0;
    G174_o2 <= 1'b0;
    G177_o2 <= 1'b0;
    G180_o2 <= 1'b0;
  end
endmodule


