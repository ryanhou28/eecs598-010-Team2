
module mymod
(
  G1_p,
  G1_n,
  G2_p,
  G2_n,
  G3_p,
  G3_n,
  G4_p,
  G4_n,
  G5_p,
  G5_n,
  G6_p,
  G6_n,
  G7_p,
  G7_n,
  G8_p,
  G8_n,
  G9_p,
  G9_n,
  G10_p,
  G10_n,
  G11_p,
  G11_n,
  G12_p,
  G12_n,
  G13_p,
  G13_n,
  G14_p,
  G14_n,
  G15_p,
  G15_n,
  G16_p,
  G16_n,
  G17_p,
  G17_n,
  G18_p,
  G18_n,
  G19_p,
  G19_n,
  G20_p,
  G20_n,
  G21_p,
  G21_n,
  G22_p,
  G22_n,
  G23_p,
  G23_n,
  G24_p,
  G24_n,
  G25_p,
  G25_n,
  G26_p,
  G26_n,
  G27_p,
  G27_n,
  G28_p,
  G28_n,
  G29_p,
  G29_n,
  G30_p,
  G30_n,
  G31_p,
  G31_n,
  G32_p,
  G32_n,
  G33_p,
  G33_n,
  G34_p,
  G34_n,
  G35_p,
  G35_n,
  G36_p,
  G36_n,
  G37_p,
  G37_n,
  G38_p,
  G38_n,
  G39_p,
  G39_n,
  G40_p,
  G40_n,
  G41_p,
  G41_n,
  G42_p,
  G42_n,
  G43_p,
  G43_n,
  G44_p,
  G44_n,
  G45_p,
  G45_n,
  G46_p,
  G46_n,
  G47_p,
  G47_n,
  G48_p,
  G48_n,
  G49_p,
  G49_n,
  G50_p,
  G50_n,
  G51_p,
  G51_n,
  G52_p,
  G52_n,
  G53_p,
  G53_n,
  G54_p,
  G54_n,
  G55_p,
  G55_n,
  G56_p,
  G56_n,
  G57_p,
  G57_n,
  G58_p,
  G58_n,
  G59_p,
  G59_n,
  G60_p,
  G60_n,
  G61_p,
  G61_n,
  G62_p,
  G62_n,
  G63_p,
  G63_n,
  G64_p,
  G64_n,
  G65_p,
  G65_n,
  G66_p,
  G66_n,
  G67_p,
  G67_n,
  G68_p,
  G68_n,
  G69_p,
  G69_n,
  G70_p,
  G70_n,
  G71_p,
  G71_n,
  G72_p,
  G72_n,
  G73_p,
  G73_n,
  G74_p,
  G74_n,
  G75_p,
  G75_n,
  G76_p,
  G76_n,
  G77_p,
  G77_n,
  G78_p,
  G78_n,
  G79_p,
  G79_n,
  G80_p,
  G80_n,
  G81_p,
  G81_n,
  G82_p,
  G82_n,
  G83_p,
  G83_n,
  G84_p,
  G84_n,
  G85_p,
  G85_n,
  G86_p,
  G86_n,
  G87_p,
  G87_n,
  G88_p,
  G88_n,
  G89_p,
  G89_n,
  G90_p,
  G90_n,
  G91_p,
  G91_n,
  G92_p,
  G92_n,
  G93_p,
  G93_n,
  G94_p,
  G94_n,
  G95_p,
  G95_n,
  G96_p,
  G96_n,
  G97_p,
  G97_n,
  G98_p,
  G98_n,
  G99_p,
  G99_n,
  G100_p,
  G100_n,
  G101_p,
  G101_n,
  G102_p,
  G102_n,
  G103_p,
  G103_n,
  G104_p,
  G104_n,
  G105_p,
  G105_n,
  G106_p,
  G106_n,
  G107_p,
  G107_n,
  G108_p,
  G108_n,
  G109_p,
  G109_n,
  G110_p,
  G110_n,
  G111_p,
  G111_n,
  G112_p,
  G112_n,
  G113_p,
  G113_n,
  G114_p,
  G114_n,
  G115_p,
  G115_n,
  G116_p,
  G116_n,
  G117_p,
  G117_n,
  G118_p,
  G118_n,
  G119_p,
  G119_n,
  G120_p,
  G120_n,
  G121_p,
  G121_n,
  G122_p,
  G122_n,
  G123_p,
  G123_n,
  G124_p,
  G124_n,
  G125_p,
  G125_n,
  G126_p,
  G126_n,
  G127_p,
  G127_n,
  G128_p,
  G128_n,
  G129_p,
  G129_n,
  G130_p,
  G130_n,
  G131_p,
  G131_n,
  G132_p,
  G132_n,
  G133_p,
  G133_n,
  G134_p,
  G134_n,
  G135_p,
  G135_n,
  G136_p,
  G136_n,
  G137_p,
  G137_n,
  G138_p,
  G138_n,
  G139_p,
  G139_n,
  G140_p,
  G140_n,
  G141_p,
  G141_n,
  G142_p,
  G142_n,
  G143_p,
  G143_n,
  G144_p,
  G144_n,
  G145_p,
  G145_n,
  G146_p,
  G146_n,
  G147_p,
  G147_n,
  G148_p,
  G148_n,
  G149_p,
  G149_n,
  G150_p,
  G150_n,
  G151_p,
  G151_n,
  G152_p,
  G152_n,
  G153_p,
  G153_n,
  G154_p,
  G154_n,
  G155_p,
  G155_n,
  G156_p,
  G156_n,
  G157_p,
  G157_n,
  G158_p,
  G158_n,
  G159_p,
  G159_n,
  G160_p,
  G160_n,
  G161_p,
  G161_n,
  G162_p,
  G162_n,
  G163_p,
  G163_n,
  G164_p,
  G164_n,
  G165_p,
  G165_n,
  G166_p,
  G166_n,
  G167_p,
  G167_n,
  G168_p,
  G168_n,
  G169_p,
  G169_n,
  G170_p,
  G170_n,
  G171_p,
  G171_n,
  G172_p,
  G172_n,
  G173_p,
  G173_n,
  G174_p,
  G174_n,
  G175_p,
  G175_n,
  G176_p,
  G176_n,
  G177_p,
  G177_n,
  G178_p,
  G178_n,
  G5193_p,
  G5194_p,
  G5195_p,
  G5196_p,
  G5197_p,
  G5198_p,
  G5199_n,
  G5200_p,
  G5201_p,
  G5202_p,
  G5203_p,
  G5204_p,
  G5205_p,
  G5206_p,
  G5207_p,
  G5208_p,
  G5209_p,
  G5210_p,
  G5211_p,
  G5212_p,
  G5213_p,
  G5214_p,
  G5215_p,
  G5216_p,
  G5217_p,
  G5218_p,
  G5219_p,
  G5220_p,
  G5221_p,
  G5222_p,
  G5223_p,
  G5224_p,
  G5225_p,
  G5226_p,
  G5227_p,
  G5228_p,
  G5229_p,
  G5230_p,
  G5231_p,
  G5232_p,
  G5233_p,
  G5234_p,
  G5235_p,
  G5236_p,
  G5237_p,
  G5238_n,
  G5239_p,
  G5240_p,
  G5241_n,
  G5242_n,
  G5243_n,
  G5244_n,
  G5245_p,
  G5246_n,
  G5247_p,
  G5248_n,
  G5249_p,
  G5250_n,
  G5251_p,
  G5252_p,
  G5253_n,
  G5254_n,
  G5255_n,
  G5256_p,
  G5257_n,
  G5258_n,
  G5259_n,
  G5260_p,
  G5261_n,
  G5262_n,
  G5263_n,
  G5264_n,
  G5265_p,
  G5266_p,
  G5267_p,
  G5268_p,
  G5269_p,
  G5270_n,
  G5271_p,
  G5272_p,
  G5273_p,
  G5274_n,
  G5275_p,
  G5276_n,
  G5277_p,
  G5278_p,
  G5279_p,
  G5280_n,
  G5281_p,
  G5282_p,
  G5283_p,
  G5284_p,
  G5285_n,
  G5286_n,
  G5287_n,
  G5288_n,
  G5289_n,
  G5290_n,
  G5291_n,
  G5292_n,
  G5293_n,
  G5294_p,
  G5295_p,
  G5296_p,
  G5297_p,
  G5298_p,
  G5299_p,
  G5300_p,
  G5301_p,
  G5302_p,
  G5303_p,
  G5304_p,
  G5305_p,
  G5306_p,
  G5307_p,
  G5308_p,
  G5309_p,
  G5310_p,
  G5311_p,
  G5312_n,
  G5313_n,
  G5314_p,
  G5315_p
);

  input G1_p;input G1_n;input G2_p;input G2_n;input G3_p;input G3_n;input G4_p;input G4_n;input G5_p;input G5_n;input G6_p;input G6_n;input G7_p;input G7_n;input G8_p;input G8_n;input G9_p;input G9_n;input G10_p;input G10_n;input G11_p;input G11_n;input G12_p;input G12_n;input G13_p;input G13_n;input G14_p;input G14_n;input G15_p;input G15_n;input G16_p;input G16_n;input G17_p;input G17_n;input G18_p;input G18_n;input G19_p;input G19_n;input G20_p;input G20_n;input G21_p;input G21_n;input G22_p;input G22_n;input G23_p;input G23_n;input G24_p;input G24_n;input G25_p;input G25_n;input G26_p;input G26_n;input G27_p;input G27_n;input G28_p;input G28_n;input G29_p;input G29_n;input G30_p;input G30_n;input G31_p;input G31_n;input G32_p;input G32_n;input G33_p;input G33_n;input G34_p;input G34_n;input G35_p;input G35_n;input G36_p;input G36_n;input G37_p;input G37_n;input G38_p;input G38_n;input G39_p;input G39_n;input G40_p;input G40_n;input G41_p;input G41_n;input G42_p;input G42_n;input G43_p;input G43_n;input G44_p;input G44_n;input G45_p;input G45_n;input G46_p;input G46_n;input G47_p;input G47_n;input G48_p;input G48_n;input G49_p;input G49_n;input G50_p;input G50_n;input G51_p;input G51_n;input G52_p;input G52_n;input G53_p;input G53_n;input G54_p;input G54_n;input G55_p;input G55_n;input G56_p;input G56_n;input G57_p;input G57_n;input G58_p;input G58_n;input G59_p;input G59_n;input G60_p;input G60_n;input G61_p;input G61_n;input G62_p;input G62_n;input G63_p;input G63_n;input G64_p;input G64_n;input G65_p;input G65_n;input G66_p;input G66_n;input G67_p;input G67_n;input G68_p;input G68_n;input G69_p;input G69_n;input G70_p;input G70_n;input G71_p;input G71_n;input G72_p;input G72_n;input G73_p;input G73_n;input G74_p;input G74_n;input G75_p;input G75_n;input G76_p;input G76_n;input G77_p;input G77_n;input G78_p;input G78_n;input G79_p;input G79_n;input G80_p;input G80_n;input G81_p;input G81_n;input G82_p;input G82_n;input G83_p;input G83_n;input G84_p;input G84_n;input G85_p;input G85_n;input G86_p;input G86_n;input G87_p;input G87_n;input G88_p;input G88_n;input G89_p;input G89_n;input G90_p;input G90_n;input G91_p;input G91_n;input G92_p;input G92_n;input G93_p;input G93_n;input G94_p;input G94_n;input G95_p;input G95_n;input G96_p;input G96_n;input G97_p;input G97_n;input G98_p;input G98_n;input G99_p;input G99_n;input G100_p;input G100_n;input G101_p;input G101_n;input G102_p;input G102_n;input G103_p;input G103_n;input G104_p;input G104_n;input G105_p;input G105_n;input G106_p;input G106_n;input G107_p;input G107_n;input G108_p;input G108_n;input G109_p;input G109_n;input G110_p;input G110_n;input G111_p;input G111_n;input G112_p;input G112_n;input G113_p;input G113_n;input G114_p;input G114_n;input G115_p;input G115_n;input G116_p;input G116_n;input G117_p;input G117_n;input G118_p;input G118_n;input G119_p;input G119_n;input G120_p;input G120_n;input G121_p;input G121_n;input G122_p;input G122_n;input G123_p;input G123_n;input G124_p;input G124_n;input G125_p;input G125_n;input G126_p;input G126_n;input G127_p;input G127_n;input G128_p;input G128_n;input G129_p;input G129_n;input G130_p;input G130_n;input G131_p;input G131_n;input G132_p;input G132_n;input G133_p;input G133_n;input G134_p;input G134_n;input G135_p;input G135_n;input G136_p;input G136_n;input G137_p;input G137_n;input G138_p;input G138_n;input G139_p;input G139_n;input G140_p;input G140_n;input G141_p;input G141_n;input G142_p;input G142_n;input G143_p;input G143_n;input G144_p;input G144_n;input G145_p;input G145_n;input G146_p;input G146_n;input G147_p;input G147_n;input G148_p;input G148_n;input G149_p;input G149_n;input G150_p;input G150_n;input G151_p;input G151_n;input G152_p;input G152_n;input G153_p;input G153_n;input G154_p;input G154_n;input G155_p;input G155_n;input G156_p;input G156_n;input G157_p;input G157_n;input G158_p;input G158_n;input G159_p;input G159_n;input G160_p;input G160_n;input G161_p;input G161_n;input G162_p;input G162_n;input G163_p;input G163_n;input G164_p;input G164_n;input G165_p;input G165_n;input G166_p;input G166_n;input G167_p;input G167_n;input G168_p;input G168_n;input G169_p;input G169_n;input G170_p;input G170_n;input G171_p;input G171_n;input G172_p;input G172_n;input G173_p;input G173_n;input G174_p;input G174_n;input G175_p;input G175_n;input G176_p;input G176_n;input G177_p;input G177_n;input G178_p;input G178_n;
  output G5193_p;output G5194_p;output G5195_p;output G5196_p;output G5197_p;output G5198_p;output G5199_n;output G5200_p;output G5201_p;output G5202_p;output G5203_p;output G5204_p;output G5205_p;output G5206_p;output G5207_p;output G5208_p;output G5209_p;output G5210_p;output G5211_p;output G5212_p;output G5213_p;output G5214_p;output G5215_p;output G5216_p;output G5217_p;output G5218_p;output G5219_p;output G5220_p;output G5221_p;output G5222_p;output G5223_p;output G5224_p;output G5225_p;output G5226_p;output G5227_p;output G5228_p;output G5229_p;output G5230_p;output G5231_p;output G5232_p;output G5233_p;output G5234_p;output G5235_p;output G5236_p;output G5237_p;output G5238_n;output G5239_p;output G5240_p;output G5241_n;output G5242_n;output G5243_n;output G5244_n;output G5245_p;output G5246_n;output G5247_p;output G5248_n;output G5249_p;output G5250_n;output G5251_p;output G5252_p;output G5253_n;output G5254_n;output G5255_n;output G5256_p;output G5257_n;output G5258_n;output G5259_n;output G5260_p;output G5261_n;output G5262_n;output G5263_n;output G5264_n;output G5265_p;output G5266_p;output G5267_p;output G5268_p;output G5269_p;output G5270_n;output G5271_p;output G5272_p;output G5273_p;output G5274_n;output G5275_p;output G5276_n;output G5277_p;output G5278_p;output G5279_p;output G5280_n;output G5281_p;output G5282_p;output G5283_p;output G5284_p;output G5285_n;output G5286_n;output G5287_n;output G5288_n;output G5289_n;output G5290_n;output G5291_n;output G5292_n;output G5293_n;output G5294_p;output G5295_p;output G5296_p;output G5297_p;output G5298_p;output G5299_p;output G5300_p;output G5301_p;output G5302_p;output G5303_p;output G5304_p;output G5305_p;output G5306_p;output G5307_p;output G5308_p;output G5309_p;output G5310_p;output G5311_p;output G5312_n;output G5313_n;output G5314_p;output G5315_p;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire G51_p;
  wire G51_n;
  wire G52_p;
  wire G52_n;
  wire G53_p;
  wire G53_n;
  wire G54_p;
  wire G54_n;
  wire G55_p;
  wire G55_n;
  wire G56_p;
  wire G56_n;
  wire G57_p;
  wire G57_n;
  wire G58_p;
  wire G58_n;
  wire G59_p;
  wire G59_n;
  wire G60_p;
  wire G60_n;
  wire G61_p;
  wire G61_n;
  wire G62_p;
  wire G62_n;
  wire G63_p;
  wire G63_n;
  wire G64_p;
  wire G64_n;
  wire G65_p;
  wire G65_n;
  wire G66_p;
  wire G66_n;
  wire G67_p;
  wire G67_n;
  wire G68_p;
  wire G68_n;
  wire G69_p;
  wire G69_n;
  wire G70_p;
  wire G70_n;
  wire G71_p;
  wire G71_n;
  wire G72_p;
  wire G72_n;
  wire G73_p;
  wire G73_n;
  wire G74_p;
  wire G74_n;
  wire G75_p;
  wire G75_n;
  wire G76_p;
  wire G76_n;
  wire G77_p;
  wire G77_n;
  wire G78_p;
  wire G78_n;
  wire G79_p;
  wire G79_n;
  wire G80_p;
  wire G80_n;
  wire G81_p;
  wire G81_n;
  wire G82_p;
  wire G82_n;
  wire G83_p;
  wire G83_n;
  wire G84_p;
  wire G84_n;
  wire G85_p;
  wire G85_n;
  wire G86_p;
  wire G86_n;
  wire G87_p;
  wire G87_n;
  wire G88_p;
  wire G88_n;
  wire G89_p;
  wire G89_n;
  wire G90_p;
  wire G90_n;
  wire G91_p;
  wire G91_n;
  wire G92_p;
  wire G92_n;
  wire G93_p;
  wire G93_n;
  wire G94_p;
  wire G94_n;
  wire G95_p;
  wire G95_n;
  wire G96_p;
  wire G96_n;
  wire G97_p;
  wire G97_n;
  wire G98_p;
  wire G98_n;
  wire G99_p;
  wire G99_n;
  wire G100_p;
  wire G100_n;
  wire G101_p;
  wire G101_n;
  wire G102_p;
  wire G102_n;
  wire G103_p;
  wire G103_n;
  wire G104_p;
  wire G104_n;
  wire G105_p;
  wire G105_n;
  wire G106_p;
  wire G106_n;
  wire G107_p;
  wire G107_n;
  wire G108_p;
  wire G108_n;
  wire G109_p;
  wire G109_n;
  wire G110_p;
  wire G110_n;
  wire G111_p;
  wire G111_n;
  wire G112_p;
  wire G112_n;
  wire G113_p;
  wire G113_n;
  wire G114_p;
  wire G114_n;
  wire G115_p;
  wire G115_n;
  wire G116_p;
  wire G116_n;
  wire G117_p;
  wire G117_n;
  wire G118_p;
  wire G118_n;
  wire G119_p;
  wire G119_n;
  wire G120_p;
  wire G120_n;
  wire G121_p;
  wire G121_n;
  wire G122_p;
  wire G122_n;
  wire G123_p;
  wire G123_n;
  wire G124_p;
  wire G124_n;
  wire G125_p;
  wire G125_n;
  wire G126_p;
  wire G126_n;
  wire G127_p;
  wire G127_n;
  wire G128_p;
  wire G128_n;
  wire G129_p;
  wire G129_n;
  wire G130_p;
  wire G130_n;
  wire G131_p;
  wire G131_n;
  wire G132_p;
  wire G132_n;
  wire G133_p;
  wire G133_n;
  wire G134_p;
  wire G134_n;
  wire G135_p;
  wire G135_n;
  wire G136_p;
  wire G136_n;
  wire G137_p;
  wire G137_n;
  wire G138_p;
  wire G138_n;
  wire G139_p;
  wire G139_n;
  wire G140_p;
  wire G140_n;
  wire G141_p;
  wire G141_n;
  wire G142_p;
  wire G142_n;
  wire G143_p;
  wire G143_n;
  wire G144_p;
  wire G144_n;
  wire G145_p;
  wire G145_n;
  wire G146_p;
  wire G146_n;
  wire G147_p;
  wire G147_n;
  wire G148_p;
  wire G148_n;
  wire G149_p;
  wire G149_n;
  wire G150_p;
  wire G150_n;
  wire G151_p;
  wire G151_n;
  wire G152_p;
  wire G152_n;
  wire G153_p;
  wire G153_n;
  wire G154_p;
  wire G154_n;
  wire G155_p;
  wire G155_n;
  wire G156_p;
  wire G156_n;
  wire G157_p;
  wire G157_n;
  wire G158_p;
  wire G158_n;
  wire G159_p;
  wire G159_n;
  wire G160_p;
  wire G160_n;
  wire G161_p;
  wire G161_n;
  wire G162_p;
  wire G162_n;
  wire G163_p;
  wire G163_n;
  wire G164_p;
  wire G164_n;
  wire G165_p;
  wire G165_n;
  wire G166_p;
  wire G166_n;
  wire G167_p;
  wire G167_n;
  wire G168_p;
  wire G168_n;
  wire G169_p;
  wire G169_n;
  wire G170_p;
  wire G170_n;
  wire G171_p;
  wire G171_n;
  wire G172_p;
  wire G172_n;
  wire G173_p;
  wire G173_n;
  wire G174_p;
  wire G174_n;
  wire G175_p;
  wire G175_n;
  wire G176_p;
  wire G176_n;
  wire G177_p;
  wire G177_n;
  wire G178_p;
  wire G178_n;
  wire ffc_0_p;
  wire ffc_0_n;
  wire ffc_1_p;
  wire ffc_1_n;
  wire ffc_2_p;
  wire ffc_2_n;
  wire ffc_3_p;
  wire ffc_3_n;
  wire ffc_4_p;
  wire ffc_4_n;
  wire ffc_5_p;
  wire ffc_5_n;
  wire ffc_6_p;
  wire ffc_6_n;
  wire ffc_7_p;
  wire ffc_7_n;
  wire ffc_8_p;
  wire ffc_8_n;
  wire ffc_9_p;
  wire ffc_9_n;
  wire ffc_10_p;
  wire ffc_10_n;
  wire ffc_11_p;
  wire ffc_11_n;
  wire ffc_12_p;
  wire ffc_12_n;
  wire ffc_13_p;
  wire ffc_13_n;
  wire ffc_14_p;
  wire ffc_14_n;
  wire ffc_15_p;
  wire ffc_15_n;
  wire ffc_16_p;
  wire ffc_16_n;
  wire ffc_17_p;
  wire ffc_17_n;
  wire ffc_18_p;
  wire ffc_18_n;
  wire ffc_19_p;
  wire ffc_19_n;
  wire ffc_20_p;
  wire ffc_20_n;
  wire ffc_21_p;
  wire ffc_21_n;
  wire ffc_22_p;
  wire ffc_22_n;
  wire ffc_23_p;
  wire ffc_23_n;
  wire ffc_24_p;
  wire ffc_24_n;
  wire ffc_25_p;
  wire ffc_25_n;
  wire ffc_26_p;
  wire ffc_26_n;
  wire ffc_27_p;
  wire ffc_27_n;
  wire ffc_28_p;
  wire ffc_28_n;
  wire ffc_29_p;
  wire ffc_29_n;
  wire ffc_30_p;
  wire ffc_30_n;
  wire ffc_31_p;
  wire ffc_31_n;
  wire ffc_32_p;
  wire ffc_32_n;
  wire ffc_33_p;
  wire ffc_33_n;
  wire ffc_34_p;
  wire ffc_34_n;
  wire ffc_35_p;
  wire ffc_35_n;
  wire ffc_36_p;
  wire ffc_36_n;
  wire ffc_37_p;
  wire ffc_37_n;
  wire ffc_38_p;
  wire ffc_38_n;
  wire ffc_39_p;
  wire ffc_39_n;
  wire ffc_40_p;
  wire ffc_40_n;
  wire ffc_41_p;
  wire ffc_41_n;
  wire ffc_42_p;
  wire ffc_42_n;
  wire ffc_43_p;
  wire ffc_43_n;
  wire ffc_44_p;
  wire ffc_44_n;
  wire ffc_45_p;
  wire ffc_45_n;
  wire ffc_46_p;
  wire ffc_46_n;
  wire ffc_47_p;
  wire ffc_47_n;
  wire ffc_48_p;
  wire ffc_48_n;
  wire ffc_49_p;
  wire ffc_49_n;
  wire ffc_50_p;
  wire ffc_50_n;
  wire ffc_51_p;
  wire ffc_51_n;
  wire ffc_52_p;
  wire ffc_52_n;
  wire ffc_53_p;
  wire ffc_53_n;
  wire ffc_54_p;
  wire ffc_54_n;
  wire ffc_55_p;
  wire ffc_55_n;
  wire ffc_56_p;
  wire ffc_56_n;
  wire ffc_57_p;
  wire ffc_57_n;
  wire ffc_58_p;
  wire ffc_58_n;
  wire ffc_59_p;
  wire ffc_59_n;
  wire ffc_60_p;
  wire ffc_60_n;
  wire ffc_61_p;
  wire ffc_61_n;
  wire ffc_62_p;
  wire ffc_62_n;
  wire ffc_63_p;
  wire ffc_63_n;
  wire ffc_64_p;
  wire ffc_64_n;
  wire ffc_65_p;
  wire ffc_65_n;
  wire ffc_66_p;
  wire ffc_66_n;
  wire ffc_67_p;
  wire ffc_67_n;
  wire ffc_68_p;
  wire ffc_68_n;
  wire ffc_69_p;
  wire ffc_69_n;
  wire ffc_70_p;
  wire ffc_70_n;
  wire ffc_71_p;
  wire ffc_71_n;
  wire ffc_72_p;
  wire ffc_72_n;
  wire ffc_73_p;
  wire ffc_73_n;
  wire ffc_74_p;
  wire ffc_74_n;
  wire ffc_75_p;
  wire ffc_75_n;
  wire ffc_76_p;
  wire ffc_76_n;
  wire ffc_77_p;
  wire ffc_77_n;
  wire ffc_78_p;
  wire ffc_78_n;
  wire ffc_79_p;
  wire ffc_79_n;
  wire ffc_80_p;
  wire ffc_80_n;
  wire ffc_81_p;
  wire ffc_81_n;
  wire ffc_82_p;
  wire ffc_82_n;
  wire ffc_83_p;
  wire ffc_83_n;
  wire ffc_84_p;
  wire ffc_84_n;
  wire ffc_85_p;
  wire ffc_85_n;
  wire ffc_86_p;
  wire ffc_86_n;
  wire ffc_87_p;
  wire ffc_87_n;
  wire ffc_88_p;
  wire ffc_88_n;
  wire ffc_89_p;
  wire ffc_89_n;
  wire ffc_90_p;
  wire ffc_90_n;
  wire ffc_91_p;
  wire ffc_91_n;
  wire ffc_92_p;
  wire ffc_92_n;
  wire ffc_93_p;
  wire ffc_93_n;
  wire ffc_94_p;
  wire ffc_94_n;
  wire ffc_95_p;
  wire ffc_95_n;
  wire ffc_96_p;
  wire ffc_96_n;
  wire ffc_97_p;
  wire ffc_97_n;
  wire ffc_98_p;
  wire ffc_98_n;
  wire ffc_99_p;
  wire ffc_99_n;
  wire ffc_100_p;
  wire ffc_100_n;
  wire ffc_101_p;
  wire ffc_101_n;
  wire ffc_102_p;
  wire ffc_102_n;
  wire ffc_103_p;
  wire ffc_103_n;
  wire ffc_104_p;
  wire ffc_104_n;
  wire ffc_105_p;
  wire ffc_105_n;
  wire ffc_106_p;
  wire ffc_106_n;
  wire ffc_107_p;
  wire ffc_107_n;
  wire ffc_108_p;
  wire ffc_108_n;
  wire ffc_109_p;
  wire ffc_109_n;
  wire ffc_110_p;
  wire ffc_110_n;
  wire ffc_111_p;
  wire ffc_111_n;
  wire ffc_112_p;
  wire ffc_112_n;
  wire ffc_113_p;
  wire ffc_113_n;
  wire ffc_114_p;
  wire ffc_114_n;
  wire ffc_115_p;
  wire ffc_115_n;
  wire ffc_116_p;
  wire ffc_116_n;
  wire ffc_117_p;
  wire ffc_117_n;
  wire ffc_118_p;
  wire ffc_118_n;
  wire ffc_119_p;
  wire ffc_119_n;
  wire ffc_120_p;
  wire ffc_120_n;
  wire ffc_121_p;
  wire ffc_121_n;
  wire ffc_122_p;
  wire ffc_122_n;
  wire ffc_123_p;
  wire ffc_123_n;
  wire ffc_124_p;
  wire ffc_124_n;
  wire ffc_125_p;
  wire ffc_125_n;
  wire ffc_126_p;
  wire ffc_126_n;
  wire ffc_127_p;
  wire ffc_127_n;
  wire ffc_128_p;
  wire ffc_128_n;
  wire ffc_129_p;
  wire ffc_129_n;
  wire ffc_130_p;
  wire ffc_130_n;
  wire ffc_131_p;
  wire ffc_131_n;
  wire ffc_132_p;
  wire ffc_132_n;
  wire ffc_133_p;
  wire ffc_133_n;
  wire ffc_134_p;
  wire ffc_134_n;
  wire ffc_135_p;
  wire ffc_135_n;
  wire ffc_136_p;
  wire ffc_136_n;
  wire ffc_137_p;
  wire ffc_137_n;
  wire ffc_138_p;
  wire ffc_138_n;
  wire ffc_139_p;
  wire ffc_139_n;
  wire ffc_140_p;
  wire ffc_140_n;
  wire ffc_141_p;
  wire ffc_141_n;
  wire ffc_142_p;
  wire ffc_142_n;
  wire ffc_143_p;
  wire ffc_143_n;
  wire ffc_144_p;
  wire ffc_144_n;
  wire ffc_145_p;
  wire ffc_145_n;
  wire ffc_146_p;
  wire ffc_146_n;
  wire ffc_147_p;
  wire ffc_147_n;
  wire ffc_148_p;
  wire ffc_148_n;
  wire ffc_149_p;
  wire ffc_149_n;
  wire ffc_150_p;
  wire ffc_150_n;
  wire ffc_151_p;
  wire ffc_151_n;
  wire ffc_152_p;
  wire ffc_152_n;
  wire ffc_153_p;
  wire ffc_153_n;
  wire ffc_154_p;
  wire ffc_154_n;
  wire ffc_155_p;
  wire ffc_155_n;
  wire ffc_156_p;
  wire ffc_156_n;
  wire ffc_157_p;
  wire ffc_157_n;
  wire ffc_158_p;
  wire ffc_158_n;
  wire ffc_159_p;
  wire ffc_159_n;
  wire ffc_160_p;
  wire ffc_160_n;
  wire ffc_161_p;
  wire ffc_161_n;
  wire ffc_162_p;
  wire ffc_162_n;
  wire ffc_163_p;
  wire ffc_163_n;
  wire ffc_164_p;
  wire ffc_164_n;
  wire ffc_165_p;
  wire ffc_165_n;
  wire ffc_166_p;
  wire ffc_166_n;
  wire ffc_167_p;
  wire ffc_167_n;
  wire ffc_168_p;
  wire ffc_168_n;
  wire ffc_169_p;
  wire ffc_169_n;
  wire ffc_170_p;
  wire ffc_170_n;
  wire ffc_171_p;
  wire ffc_171_n;
  wire ffc_172_p;
  wire ffc_172_n;
  wire ffc_173_p;
  wire ffc_173_n;
  wire ffc_174_p;
  wire ffc_174_n;
  wire ffc_175_p;
  wire ffc_175_n;
  wire ffc_176_p;
  wire ffc_176_n;
  wire ffc_177_p;
  wire ffc_177_n;
  wire ffc_178_p;
  wire ffc_178_n;
  wire ffc_179_p;
  wire ffc_179_n;
  wire ffc_180_p;
  wire ffc_180_n;
  wire ffc_181_p;
  wire ffc_181_n;
  wire ffc_182_p;
  wire ffc_182_n;
  wire ffc_183_p;
  wire ffc_183_n;
  wire ffc_184_p;
  wire ffc_184_n;
  wire ffc_185_p;
  wire ffc_185_n;
  wire ffc_186_p;
  wire ffc_186_n;
  wire ffc_187_p;
  wire ffc_187_n;
  wire ffc_188_p;
  wire ffc_188_n;
  wire ffc_189_p;
  wire ffc_189_n;
  wire ffc_190_p;
  wire ffc_190_n;
  wire ffc_191_p;
  wire ffc_191_n;
  wire ffc_192_p;
  wire ffc_192_n;
  wire ffc_193_p;
  wire ffc_193_n;
  wire ffc_194_p;
  wire ffc_194_n;
  wire ffc_195_p;
  wire ffc_195_n;
  wire ffc_196_p;
  wire ffc_196_n;
  wire ffc_197_p;
  wire ffc_197_n;
  wire ffc_198_p;
  wire ffc_198_n;
  wire ffc_199_p;
  wire ffc_199_n;
  wire ffc_200_p;
  wire ffc_200_n;
  wire ffc_201_p;
  wire ffc_201_n;
  wire ffc_202_p;
  wire ffc_202_n;
  wire ffc_203_p;
  wire ffc_203_n;
  wire ffc_204_p;
  wire ffc_204_n;
  wire ffc_205_p;
  wire ffc_205_n;
  wire ffc_206_p;
  wire ffc_206_n;
  wire ffc_207_p;
  wire ffc_207_n;
  wire ffc_208_p;
  wire ffc_208_n;
  wire ffc_209_p;
  wire ffc_209_n;
  wire ffc_210_p;
  wire ffc_210_n;
  wire ffc_211_p;
  wire ffc_211_n;
  wire ffc_212_p;
  wire ffc_212_n;
  wire ffc_213_p;
  wire ffc_213_n;
  wire ffc_214_p;
  wire ffc_214_n;
  wire ffc_215_p;
  wire ffc_215_n;
  wire ffc_216_p;
  wire ffc_216_n;
  wire ffc_217_p;
  wire ffc_217_n;
  wire ffc_218_p;
  wire ffc_218_n;
  wire ffc_219_p;
  wire ffc_219_n;
  wire ffc_220_p;
  wire ffc_220_n;
  wire ffc_221_p;
  wire ffc_221_n;
  wire ffc_222_p;
  wire ffc_222_n;
  wire ffc_223_p;
  wire ffc_223_n;
  wire ffc_224_p;
  wire ffc_224_n;
  wire ffc_225_p;
  wire ffc_225_n;
  wire ffc_226_p;
  wire ffc_226_n;
  wire ffc_227_p;
  wire ffc_227_n;
  wire ffc_228_p;
  wire ffc_228_n;
  wire ffc_229_p;
  wire ffc_229_n;
  wire ffc_230_p;
  wire ffc_230_n;
  wire ffc_231_p;
  wire ffc_231_n;
  wire ffc_232_p;
  wire ffc_232_n;
  wire ffc_233_p;
  wire ffc_233_n;
  wire ffc_234_p;
  wire ffc_234_n;
  wire ffc_235_p;
  wire ffc_235_n;
  wire ffc_236_p;
  wire ffc_236_n;
  wire ffc_237_p;
  wire ffc_237_n;
  wire ffc_238_p;
  wire ffc_238_n;
  wire ffc_239_p;
  wire ffc_239_n;
  wire ffc_240_p;
  wire ffc_240_n;
  wire ffc_241_p;
  wire ffc_241_n;
  wire ffc_242_p;
  wire ffc_242_n;
  wire ffc_243_p;
  wire ffc_243_n;
  wire ffc_244_p;
  wire ffc_244_n;
  wire ffc_245_p;
  wire ffc_245_n;
  wire ffc_246_p;
  wire ffc_246_n;
  wire ffc_247_p;
  wire ffc_247_n;
  wire ffc_248_p;
  wire ffc_248_n;
  wire ffc_249_p;
  wire ffc_249_n;
  wire ffc_250_p;
  wire ffc_250_n;
  wire ffc_251_p;
  wire ffc_251_n;
  wire ffc_252_p;
  wire ffc_252_n;
  wire ffc_253_p;
  wire ffc_253_n;
  wire ffc_254_p;
  wire ffc_254_n;
  wire ffc_255_p;
  wire ffc_255_n;
  wire ffc_256_p;
  wire ffc_256_n;
  wire ffc_257_p;
  wire ffc_257_n;
  wire ffc_258_p;
  wire ffc_258_n;
  wire ffc_259_p;
  wire ffc_259_n;
  wire ffc_260_p;
  wire ffc_260_n;
  wire ffc_261_p;
  wire ffc_261_n;
  wire ffc_262_p;
  wire ffc_262_n;
  wire ffc_263_p;
  wire ffc_263_n;
  wire ffc_264_p;
  wire ffc_264_n;
  wire ffc_265_p;
  wire ffc_265_n;
  wire ffc_266_p;
  wire ffc_266_n;
  wire ffc_267_p;
  wire ffc_267_n;
  wire ffc_268_p;
  wire ffc_268_n;
  wire ffc_269_p;
  wire ffc_269_n;
  wire ffc_270_p;
  wire ffc_270_n;
  wire ffc_271_p;
  wire ffc_271_n;
  wire ffc_272_p;
  wire ffc_272_n;
  wire ffc_273_p;
  wire ffc_273_n;
  wire ffc_274_p;
  wire ffc_274_n;
  wire ffc_275_p;
  wire ffc_275_n;
  wire ffc_276_p;
  wire ffc_276_n;
  wire ffc_277_p;
  wire ffc_277_n;
  wire ffc_278_p;
  wire ffc_278_n;
  wire ffc_279_p;
  wire ffc_279_n;
  wire ffc_280_p;
  wire ffc_280_n;
  wire ffc_281_p;
  wire ffc_281_n;
  wire ffc_282_p;
  wire ffc_282_n;
  wire ffc_283_p;
  wire ffc_283_n;
  wire ffc_284_p;
  wire ffc_284_n;
  wire ffc_285_p;
  wire ffc_285_n;
  wire ffc_286_p;
  wire ffc_286_n;
  wire ffc_287_p;
  wire ffc_287_n;
  wire ffc_288_p;
  wire ffc_288_n;
  wire ffc_289_p;
  wire ffc_289_n;
  wire ffc_290_p;
  wire ffc_290_n;
  wire ffc_291_p;
  wire ffc_291_n;
  wire ffc_292_p;
  wire ffc_292_n;
  wire ffc_293_p;
  wire ffc_293_n;
  wire ffc_294_p;
  wire ffc_294_n;
  wire ffc_295_p;
  wire ffc_295_n;
  wire ffc_296_p;
  wire ffc_296_n;
  wire ffc_297_p;
  wire ffc_297_n;
  wire ffc_298_p;
  wire ffc_298_n;
  wire ffc_299_p;
  wire ffc_299_n;
  wire ffc_300_p;
  wire ffc_300_n;
  wire ffc_301_p;
  wire ffc_301_n;
  wire ffc_302_p;
  wire ffc_302_n;
  wire ffc_303_p;
  wire ffc_303_n;
  wire ffc_304_p;
  wire ffc_304_n;
  wire ffc_305_p;
  wire ffc_305_n;
  wire ffc_306_p;
  wire ffc_306_n;
  wire ffc_307_p;
  wire ffc_307_n;
  wire ffc_308_p;
  wire ffc_308_n;
  wire ffc_309_p;
  wire ffc_309_n;
  wire ffc_310_p;
  wire ffc_310_n;
  wire ffc_311_p;
  wire ffc_311_n;
  wire ffc_312_p;
  wire ffc_312_n;
  wire ffc_313_p;
  wire ffc_313_n;
  wire ffc_314_p;
  wire ffc_314_n;
  wire ffc_315_p;
  wire ffc_315_n;
  wire ffc_316_p;
  wire ffc_316_n;
  wire ffc_317_p;
  wire ffc_317_n;
  wire ffc_318_p;
  wire ffc_318_n;
  wire ffc_319_p;
  wire ffc_319_n;
  wire ffc_320_p;
  wire ffc_320_n;
  wire ffc_321_p;
  wire ffc_321_n;
  wire ffc_322_p;
  wire ffc_322_n;
  wire ffc_323_p;
  wire ffc_323_n;
  wire ffc_324_p;
  wire ffc_324_n;
  wire ffc_325_p;
  wire ffc_325_n;
  wire ffc_326_p;
  wire ffc_326_n;
  wire ffc_327_p;
  wire ffc_327_n;
  wire ffc_328_p;
  wire ffc_328_n;
  wire ffc_329_p;
  wire ffc_329_n;
  wire ffc_330_p;
  wire ffc_330_n;
  wire ffc_331_p;
  wire ffc_331_n;
  wire ffc_332_p;
  wire ffc_332_n;
  wire ffc_333_p;
  wire ffc_333_n;
  wire ffc_334_p;
  wire ffc_334_n;
  wire ffc_335_p;
  wire ffc_335_n;
  wire ffc_336_p;
  wire ffc_336_n;
  wire ffc_337_p;
  wire ffc_337_n;
  wire ffc_338_p;
  wire ffc_338_n;
  wire ffc_339_p;
  wire ffc_339_n;
  wire ffc_340_p;
  wire ffc_340_n;
  wire ffc_341_p;
  wire ffc_341_n;
  wire ffc_342_p;
  wire ffc_342_n;
  wire ffc_343_p;
  wire ffc_343_n;
  wire ffc_344_p;
  wire ffc_344_n;
  wire ffc_345_p;
  wire ffc_345_n;
  wire ffc_346_p;
  wire ffc_346_n;
  wire ffc_347_p;
  wire ffc_347_n;
  wire ffc_348_p;
  wire ffc_348_n;
  wire ffc_349_p;
  wire ffc_349_n;
  wire ffc_350_p;
  wire ffc_350_n;
  wire ffc_351_p;
  wire ffc_351_n;
  wire ffc_352_p;
  wire ffc_352_n;
  wire ffc_353_p;
  wire ffc_353_n;
  wire ffc_354_p;
  wire ffc_354_n;
  wire ffc_355_p;
  wire ffc_355_n;
  wire ffc_356_p;
  wire ffc_356_n;
  wire ffc_357_p;
  wire ffc_357_n;
  wire ffc_358_p;
  wire ffc_358_n;
  wire ffc_359_p;
  wire ffc_359_n;
  wire ffc_360_p;
  wire ffc_360_n;
  wire ffc_361_p;
  wire ffc_361_n;
  wire ffc_362_p;
  wire ffc_362_n;
  wire ffc_363_p;
  wire ffc_363_n;
  wire ffc_364_p;
  wire ffc_364_n;
  wire ffc_365_p;
  wire ffc_365_n;
  wire ffc_366_p;
  wire ffc_366_n;
  wire ffc_367_p;
  wire ffc_367_n;
  wire ffc_368_p;
  wire ffc_368_n;
  wire ffc_369_p;
  wire ffc_369_n;
  wire ffc_370_p;
  wire ffc_370_n;
  wire ffc_371_p;
  wire ffc_371_n;
  wire ffc_372_p;
  wire ffc_372_n;
  wire ffc_373_p;
  wire ffc_373_n;
  wire ffc_374_p;
  wire ffc_374_n;
  wire ffc_375_p;
  wire ffc_375_n;
  wire ffc_376_p;
  wire ffc_376_n;
  wire ffc_377_p;
  wire ffc_377_n;
  wire ffc_378_p;
  wire ffc_378_n;
  wire ffc_379_p;
  wire ffc_379_n;
  wire ffc_380_p;
  wire ffc_380_n;
  wire ffc_381_p;
  wire ffc_381_n;
  wire ffc_382_p;
  wire ffc_382_n;
  wire ffc_383_p;
  wire ffc_383_n;
  wire ffc_384_p;
  wire ffc_384_n;
  wire ffc_385_p;
  wire ffc_385_n;
  wire ffc_386_p;
  wire ffc_386_n;
  wire ffc_387_p;
  wire ffc_387_n;
  wire ffc_388_p;
  wire ffc_388_n;
  wire ffc_389_p;
  wire ffc_389_n;
  wire ffc_390_p;
  wire ffc_390_n;
  wire ffc_391_p;
  wire ffc_391_n;
  wire ffc_392_p;
  wire ffc_392_n;
  wire ffc_393_p;
  wire ffc_393_n;
  wire ffc_394_p;
  wire ffc_394_n;
  wire ffc_395_p;
  wire ffc_395_n;
  wire ffc_396_p;
  wire ffc_396_n;
  wire ffc_397_p;
  wire ffc_397_n;
  wire ffc_398_p;
  wire ffc_398_n;
  wire ffc_399_p;
  wire ffc_399_n;
  wire ffc_400_p;
  wire ffc_400_n;
  wire ffc_401_p;
  wire ffc_401_n;
  wire ffc_402_p;
  wire ffc_402_n;
  wire ffc_403_p;
  wire ffc_403_n;
  wire ffc_404_p;
  wire ffc_404_n;
  wire ffc_405_p;
  wire ffc_405_n;
  wire ffc_406_p;
  wire ffc_406_n;
  wire ffc_407_p;
  wire ffc_407_n;
  wire ffc_408_p;
  wire ffc_408_n;
  wire ffc_409_p;
  wire ffc_409_n;
  wire ffc_410_p;
  wire ffc_410_n;
  wire ffc_411_p;
  wire ffc_411_n;
  wire ffc_412_p;
  wire ffc_412_n;
  wire ffc_413_p;
  wire ffc_413_n;
  wire ffc_414_p;
  wire ffc_414_n;
  wire ffc_415_p;
  wire ffc_415_n;
  wire ffc_416_p;
  wire ffc_416_n;
  wire ffc_417_p;
  wire ffc_417_n;
  wire ffc_418_p;
  wire ffc_418_n;
  wire ffc_419_p;
  wire ffc_419_n;
  wire ffc_420_p;
  wire ffc_420_n;
  wire ffc_421_p;
  wire ffc_421_n;
  wire ffc_422_p;
  wire ffc_422_n;
  wire ffc_423_p;
  wire ffc_423_n;
  wire ffc_424_p;
  wire ffc_424_n;
  wire ffc_425_p;
  wire ffc_425_n;
  wire ffc_426_p;
  wire ffc_426_n;
  wire ffc_427_p;
  wire ffc_427_n;
  wire ffc_428_p;
  wire ffc_428_n;
  wire ffc_429_p;
  wire ffc_429_n;
  wire ffc_430_p;
  wire ffc_430_n;
  wire ffc_431_p;
  wire ffc_431_n;
  wire ffc_432_p;
  wire ffc_432_n;
  wire ffc_433_p;
  wire ffc_433_n;
  wire ffc_434_p;
  wire ffc_434_n;
  wire ffc_435_p;
  wire ffc_435_n;
  wire ffc_436_p;
  wire ffc_436_n;
  wire ffc_437_p;
  wire ffc_437_n;
  wire ffc_438_p;
  wire ffc_438_n;
  wire ffc_439_p;
  wire ffc_439_n;
  wire ffc_440_p;
  wire ffc_440_n;
  wire ffc_441_p;
  wire ffc_441_n;
  wire ffc_442_p;
  wire ffc_442_n;
  wire ffc_443_p;
  wire ffc_443_n;
  wire ffc_444_p;
  wire ffc_444_n;
  wire ffc_445_p;
  wire ffc_445_n;
  wire ffc_446_p;
  wire ffc_446_n;
  wire ffc_447_p;
  wire ffc_447_n;
  wire ffc_448_p;
  wire ffc_448_n;
  wire ffc_449_p;
  wire ffc_449_n;
  wire ffc_450_p;
  wire ffc_450_n;
  wire ffc_451_p;
  wire ffc_451_n;
  wire ffc_452_p;
  wire ffc_452_n;
  wire ffc_453_p;
  wire ffc_453_n;
  wire ffc_454_p;
  wire ffc_454_n;
  wire ffc_455_p;
  wire ffc_455_n;
  wire ffc_456_p;
  wire ffc_456_n;
  wire ffc_457_p;
  wire ffc_457_n;
  wire ffc_458_p;
  wire ffc_458_n;
  wire ffc_459_p;
  wire ffc_459_n;
  wire ffc_460_p;
  wire ffc_460_n;
  wire ffc_461_p;
  wire ffc_461_n;
  wire ffc_462_p;
  wire ffc_462_n;
  wire ffc_463_p;
  wire ffc_463_n;
  wire ffc_464_p;
  wire ffc_464_n;
  wire ffc_465_p;
  wire ffc_465_n;
  wire ffc_466_p;
  wire ffc_466_n;
  wire ffc_467_p;
  wire ffc_467_n;
  wire ffc_468_p;
  wire ffc_468_n;
  wire ffc_469_p;
  wire ffc_469_n;
  wire ffc_470_p;
  wire ffc_470_n;
  wire ffc_471_p;
  wire ffc_471_n;
  wire ffc_472_p;
  wire ffc_472_n;
  wire ffc_473_p;
  wire ffc_473_n;
  wire ffc_474_p;
  wire ffc_474_n;
  wire ffc_475_p;
  wire ffc_475_n;
  wire ffc_476_p;
  wire ffc_476_n;
  wire ffc_477_p;
  wire ffc_477_n;
  wire ffc_478_p;
  wire ffc_478_n;
  wire ffc_479_p;
  wire ffc_479_n;
  wire ffc_480_p;
  wire ffc_480_n;
  wire ffc_481_p;
  wire ffc_481_n;
  wire ffc_482_p;
  wire ffc_482_n;
  wire ffc_483_p;
  wire ffc_483_n;
  wire ffc_484_p;
  wire ffc_484_n;
  wire ffc_485_p;
  wire ffc_485_n;
  wire ffc_486_p;
  wire ffc_486_n;
  wire ffc_487_p;
  wire ffc_487_n;
  wire ffc_488_p;
  wire ffc_488_n;
  wire ffc_489_p;
  wire ffc_489_n;
  wire ffc_490_p;
  wire ffc_490_n;
  wire ffc_491_p;
  wire ffc_491_n;
  wire ffc_492_p;
  wire ffc_492_n;
  wire ffc_493_p;
  wire ffc_493_n;
  wire ffc_494_p;
  wire ffc_494_n;
  wire ffc_495_p;
  wire ffc_495_n;
  wire ffc_496_p;
  wire ffc_496_n;
  wire ffc_497_p;
  wire ffc_497_n;
  wire ffc_498_p;
  wire ffc_498_n;
  wire ffc_499_p;
  wire ffc_499_n;
  wire ffc_500_p;
  wire ffc_500_n;
  wire ffc_501_p;
  wire ffc_501_n;
  wire ffc_502_p;
  wire ffc_502_n;
  wire ffc_503_p;
  wire ffc_503_n;
  wire ffc_504_p;
  wire ffc_504_n;
  wire ffc_505_p;
  wire ffc_505_n;
  wire ffc_506_p;
  wire ffc_506_n;
  wire ffc_507_p;
  wire ffc_507_n;
  wire ffc_508_p;
  wire ffc_508_n;
  wire ffc_509_p;
  wire ffc_509_n;
  wire ffc_510_p;
  wire ffc_510_n;
  wire ffc_511_p;
  wire ffc_511_n;
  wire ffc_512_p;
  wire ffc_512_n;
  wire ffc_513_p;
  wire ffc_513_n;
  wire ffc_514_p;
  wire ffc_514_n;
  wire ffc_515_p;
  wire ffc_515_n;
  wire ffc_516_p;
  wire ffc_516_n;
  wire ffc_517_p;
  wire ffc_517_n;
  wire ffc_518_p;
  wire ffc_518_n;
  wire ffc_519_p;
  wire ffc_519_n;
  wire ffc_520_p;
  wire ffc_520_n;
  wire ffc_521_p;
  wire ffc_521_n;
  wire ffc_522_p;
  wire ffc_522_n;
  wire ffc_523_p;
  wire ffc_523_n;
  wire ffc_524_p;
  wire ffc_524_n;
  wire ffc_525_p;
  wire ffc_525_n;
  wire ffc_526_p;
  wire ffc_526_n;
  wire ffc_527_p;
  wire ffc_527_n;
  wire ffc_528_p;
  wire ffc_528_n;
  wire ffc_529_p;
  wire ffc_529_n;
  wire ffc_530_p;
  wire ffc_530_n;
  wire ffc_531_p;
  wire ffc_531_n;
  wire ffc_532_p;
  wire ffc_532_n;
  wire ffc_533_p;
  wire ffc_533_n;
  wire ffc_534_p;
  wire ffc_534_n;
  wire ffc_535_p;
  wire ffc_535_n;
  wire ffc_536_p;
  wire ffc_536_n;
  wire ffc_537_p;
  wire ffc_537_n;
  wire ffc_538_p;
  wire ffc_538_n;
  wire ffc_539_p;
  wire ffc_539_n;
  wire ffc_540_p;
  wire ffc_540_n;
  wire ffc_541_p;
  wire ffc_541_n;
  wire ffc_542_p;
  wire ffc_542_n;
  wire ffc_543_p;
  wire ffc_543_n;
  wire ffc_544_p;
  wire ffc_544_n;
  wire ffc_545_p;
  wire ffc_545_n;
  wire ffc_546_p;
  wire ffc_546_n;
  wire ffc_547_p;
  wire ffc_547_n;
  wire ffc_548_p;
  wire ffc_548_n;
  wire ffc_549_p;
  wire ffc_549_n;
  wire ffc_550_p;
  wire ffc_550_n;
  wire ffc_551_p;
  wire ffc_551_n;
  wire ffc_552_p;
  wire ffc_552_n;
  wire ffc_553_p;
  wire ffc_553_n;
  wire ffc_554_p;
  wire ffc_554_n;
  wire ffc_555_p;
  wire ffc_555_n;
  wire ffc_556_p;
  wire ffc_556_n;
  wire ffc_557_p;
  wire ffc_557_n;
  wire ffc_558_p;
  wire ffc_558_n;
  wire ffc_559_p;
  wire ffc_559_n;
  wire ffc_560_p;
  wire ffc_560_n;
  wire ffc_561_p;
  wire ffc_561_n;
  wire ffc_562_p;
  wire ffc_562_n;
  wire ffc_563_p;
  wire ffc_563_n;
  wire ffc_564_p;
  wire ffc_564_n;
  wire ffc_565_p;
  wire ffc_565_n;
  wire ffc_566_p;
  wire ffc_566_n;
  wire ffc_567_p;
  wire ffc_567_n;
  wire ffc_568_p;
  wire ffc_568_n;
  wire ffc_569_p;
  wire ffc_569_n;
  wire ffc_570_p;
  wire ffc_570_n;
  wire ffc_571_p;
  wire ffc_571_n;
  wire ffc_572_p;
  wire ffc_572_n;
  wire ffc_573_p;
  wire ffc_573_n;
  wire ffc_574_p;
  wire ffc_574_n;
  wire ffc_575_p;
  wire ffc_575_n;
  wire ffc_576_p;
  wire ffc_576_n;
  wire ffc_577_p;
  wire ffc_577_n;
  wire ffc_578_p;
  wire ffc_578_n;
  wire ffc_579_p;
  wire ffc_579_n;
  wire ffc_580_p;
  wire ffc_580_n;
  wire ffc_581_p;
  wire ffc_581_n;
  wire ffc_582_p;
  wire ffc_582_n;
  wire ffc_583_p;
  wire ffc_583_n;
  wire ffc_584_p;
  wire ffc_584_n;
  wire ffc_585_p;
  wire ffc_585_n;
  wire ffc_586_p;
  wire ffc_586_n;
  wire ffc_587_p;
  wire ffc_587_n;
  wire ffc_588_p;
  wire ffc_588_n;
  wire ffc_589_p;
  wire ffc_589_n;
  wire ffc_590_p;
  wire ffc_590_n;
  wire ffc_591_p;
  wire ffc_591_n;
  wire ffc_592_p;
  wire ffc_592_n;
  wire ffc_593_p;
  wire ffc_593_n;
  wire ffc_594_p;
  wire ffc_594_n;
  wire ffc_595_p;
  wire ffc_595_n;
  wire ffc_596_p;
  wire ffc_596_n;
  wire ffc_597_p;
  wire ffc_597_n;
  wire ffc_598_p;
  wire ffc_598_n;
  wire ffc_599_p;
  wire ffc_599_n;
  wire ffc_600_p;
  wire ffc_600_n;
  wire ffc_601_p;
  wire ffc_601_n;
  wire ffc_602_p;
  wire ffc_602_n;
  wire ffc_603_p;
  wire ffc_603_n;
  wire ffc_604_p;
  wire ffc_604_n;
  wire ffc_605_p;
  wire ffc_605_n;
  wire ffc_606_p;
  wire ffc_606_n;
  wire ffc_607_p;
  wire ffc_607_n;
  wire ffc_608_p;
  wire ffc_608_n;
  wire ffc_609_p;
  wire ffc_609_n;
  wire ffc_610_p;
  wire ffc_610_n;
  wire ffc_611_p;
  wire ffc_611_n;
  wire ffc_612_p;
  wire ffc_612_n;
  wire ffc_613_p;
  wire ffc_613_n;
  wire ffc_614_p;
  wire ffc_614_n;
  wire ffc_615_p;
  wire ffc_615_n;
  wire ffc_616_p;
  wire ffc_616_n;
  wire ffc_617_p;
  wire ffc_617_n;
  wire ffc_618_p;
  wire ffc_618_n;
  wire ffc_619_p;
  wire ffc_619_n;
  wire ffc_620_p;
  wire ffc_620_n;
  wire ffc_621_p;
  wire ffc_621_n;
  wire ffc_622_p;
  wire ffc_622_n;
  wire ffc_623_p;
  wire ffc_623_n;
  wire ffc_624_p;
  wire ffc_624_n;
  wire ffc_625_p;
  wire ffc_625_n;
  wire ffc_626_p;
  wire ffc_626_n;
  wire ffc_627_p;
  wire ffc_627_n;
  wire ffc_628_p;
  wire ffc_628_n;
  wire ffc_629_p;
  wire ffc_629_n;
  wire ffc_630_p;
  wire ffc_630_n;
  wire ffc_631_p;
  wire ffc_631_n;
  wire ffc_632_p;
  wire ffc_632_n;
  wire ffc_633_p;
  wire ffc_633_n;
  wire ffc_634_p;
  wire ffc_634_n;
  wire ffc_635_p;
  wire ffc_635_n;
  wire ffc_636_p;
  wire ffc_636_n;
  wire ffc_637_p;
  wire ffc_637_n;
  wire ffc_638_p;
  wire ffc_638_n;
  wire ffc_639_p;
  wire ffc_639_n;
  wire ffc_640_p;
  wire ffc_640_n;
  wire ffc_641_p;
  wire ffc_641_n;
  wire ffc_642_p;
  wire ffc_642_n;
  wire ffc_643_p;
  wire ffc_643_n;
  wire ffc_644_p;
  wire ffc_644_n;
  wire ffc_645_p;
  wire ffc_645_n;
  wire ffc_646_p;
  wire ffc_646_n;
  wire ffc_647_p;
  wire ffc_647_n;
  wire ffc_648_p;
  wire ffc_648_n;
  wire ffc_649_p;
  wire ffc_649_n;
  wire ffc_650_p;
  wire ffc_650_n;
  wire ffc_651_p;
  wire ffc_651_n;
  wire ffc_652_p;
  wire ffc_652_n;
  wire ffc_653_p;
  wire ffc_653_n;
  wire ffc_654_p;
  wire ffc_654_n;
  wire ffc_655_p;
  wire ffc_655_n;
  wire ffc_656_p;
  wire ffc_656_n;
  wire ffc_657_p;
  wire ffc_657_n;
  wire ffc_658_p;
  wire ffc_658_n;
  wire ffc_659_p;
  wire ffc_659_n;
  wire ffc_660_p;
  wire ffc_660_n;
  wire ffc_661_p;
  wire ffc_661_n;
  wire ffc_662_p;
  wire ffc_662_n;
  wire ffc_663_p;
  wire ffc_663_n;
  wire ffc_664_p;
  wire ffc_664_n;
  wire ffc_665_p;
  wire ffc_665_n;
  wire ffc_666_p;
  wire ffc_666_n;
  wire ffc_667_p;
  wire ffc_667_n;
  wire ffc_668_p;
  wire ffc_668_n;
  wire ffc_669_p;
  wire ffc_669_n;
  wire ffc_670_p;
  wire ffc_670_n;
  wire ffc_671_p;
  wire ffc_671_n;
  wire ffc_672_p;
  wire ffc_672_n;
  wire ffc_673_p;
  wire ffc_673_n;
  wire ffc_674_p;
  wire ffc_674_n;
  wire ffc_675_p;
  wire ffc_675_n;
  wire ffc_676_p;
  wire ffc_676_n;
  wire ffc_677_p;
  wire ffc_677_n;
  wire ffc_678_p;
  wire ffc_678_n;
  wire ffc_679_p;
  wire ffc_679_n;
  wire ffc_680_p;
  wire ffc_680_n;
  wire ffc_681_p;
  wire ffc_681_n;
  wire ffc_682_p;
  wire ffc_682_n;
  wire ffc_683_p;
  wire ffc_683_n;
  wire ffc_684_p;
  wire ffc_684_n;
  wire ffc_685_p;
  wire ffc_685_n;
  wire ffc_686_p;
  wire ffc_686_n;
  wire ffc_687_p;
  wire ffc_687_n;
  wire ffc_688_p;
  wire ffc_688_n;
  wire ffc_689_p;
  wire ffc_689_n;
  wire ffc_690_p;
  wire ffc_690_n;
  wire ffc_691_p;
  wire ffc_691_n;
  wire ffc_692_p;
  wire ffc_692_n;
  wire ffc_693_p;
  wire ffc_693_n;
  wire ffc_694_p;
  wire ffc_694_n;
  wire ffc_695_p;
  wire ffc_695_n;
  wire ffc_696_p;
  wire ffc_696_n;
  wire ffc_697_p;
  wire ffc_697_n;
  wire ffc_698_p;
  wire ffc_698_n;
  wire ffc_699_p;
  wire ffc_699_n;
  wire ffc_700_p;
  wire ffc_700_n;
  wire ffc_701_p;
  wire ffc_701_n;
  wire ffc_702_p;
  wire ffc_702_n;
  wire ffc_703_p;
  wire ffc_703_n;
  wire ffc_704_p;
  wire ffc_704_n;
  wire ffc_705_p;
  wire ffc_705_n;
  wire ffc_706_p;
  wire ffc_706_n;
  wire ffc_707_p;
  wire ffc_707_n;
  wire ffc_708_p;
  wire ffc_708_n;
  wire ffc_709_p;
  wire ffc_709_n;
  wire ffc_710_p;
  wire ffc_710_n;
  wire ffc_711_p;
  wire ffc_711_n;
  wire ffc_712_p;
  wire ffc_712_n;
  wire ffc_713_p;
  wire ffc_713_n;
  wire ffc_714_p;
  wire ffc_714_n;
  wire ffc_715_p;
  wire ffc_715_n;
  wire ffc_716_p;
  wire ffc_716_n;
  wire ffc_717_p;
  wire ffc_717_n;
  wire ffc_718_p;
  wire ffc_718_n;
  wire ffc_719_p;
  wire ffc_719_n;
  wire ffc_720_p;
  wire ffc_720_n;
  wire ffc_721_p;
  wire ffc_721_n;
  wire ffc_722_p;
  wire ffc_722_n;
  wire ffc_723_p;
  wire ffc_723_n;
  wire ffc_724_p;
  wire ffc_724_n;
  wire ffc_725_p;
  wire ffc_725_n;
  wire ffc_726_p;
  wire ffc_726_n;
  wire ffc_727_p;
  wire ffc_727_n;
  wire ffc_728_p;
  wire ffc_728_n;
  wire ffc_729_p;
  wire ffc_729_n;
  wire ffc_730_p;
  wire ffc_730_n;
  wire ffc_731_p;
  wire ffc_731_n;
  wire ffc_732_p;
  wire ffc_732_n;
  wire ffc_733_p;
  wire ffc_733_n;
  wire ffc_734_p;
  wire ffc_734_n;
  wire ffc_735_p;
  wire ffc_735_n;
  wire ffc_736_p;
  wire ffc_736_n;
  wire ffc_737_p;
  wire ffc_737_n;
  wire ffc_738_p;
  wire ffc_738_n;
  wire ffc_739_p;
  wire ffc_739_n;
  wire ffc_740_p;
  wire ffc_740_n;
  wire ffc_741_p;
  wire ffc_741_n;
  wire ffc_742_p;
  wire ffc_742_n;
  wire ffc_743_p;
  wire ffc_743_n;
  wire ffc_744_p;
  wire ffc_744_n;
  wire ffc_745_p;
  wire ffc_745_n;
  wire ffc_746_p;
  wire ffc_746_n;
  wire ffc_747_p;
  wire ffc_747_n;
  wire ffc_748_p;
  wire ffc_748_n;
  wire ffc_749_p;
  wire ffc_749_n;
  wire ffc_750_p;
  wire ffc_750_n;
  wire ffc_751_p;
  wire ffc_751_n;
  wire ffc_752_p;
  wire ffc_752_n;
  wire ffc_753_p;
  wire ffc_753_n;
  wire ffc_754_p;
  wire ffc_754_n;
  wire ffc_755_p;
  wire ffc_755_n;
  wire ffc_756_p;
  wire ffc_756_n;
  wire ffc_757_p;
  wire ffc_757_n;
  wire ffc_758_p;
  wire ffc_758_n;
  wire ffc_759_p;
  wire ffc_759_n;
  wire ffc_760_p;
  wire ffc_760_n;
  wire ffc_761_p;
  wire ffc_761_n;
  wire ffc_762_p;
  wire ffc_762_n;
  wire ffc_763_p;
  wire ffc_763_n;
  wire ffc_764_p;
  wire ffc_764_n;
  wire ffc_765_p;
  wire ffc_765_n;
  wire ffc_766_p;
  wire ffc_766_n;
  wire ffc_767_p;
  wire ffc_767_n;
  wire ffc_768_p;
  wire ffc_768_n;
  wire ffc_769_p;
  wire ffc_769_n;
  wire ffc_770_p;
  wire ffc_770_n;
  wire ffc_771_p;
  wire ffc_771_n;
  wire ffc_772_p;
  wire ffc_772_n;
  wire ffc_773_p;
  wire ffc_773_n;
  wire ffc_774_p;
  wire ffc_774_n;
  wire ffc_775_p;
  wire ffc_775_n;
  wire ffc_776_p;
  wire ffc_776_n;
  wire ffc_777_p;
  wire ffc_777_n;
  wire ffc_778_p;
  wire ffc_778_n;
  wire ffc_779_p;
  wire ffc_779_n;
  wire ffc_780_p;
  wire ffc_780_n;
  wire ffc_781_p;
  wire ffc_781_n;
  wire ffc_782_p;
  wire ffc_782_n;
  wire ffc_783_p;
  wire ffc_783_n;
  wire ffc_784_p;
  wire ffc_784_n;
  wire ffc_785_p;
  wire ffc_785_n;
  wire ffc_786_p;
  wire ffc_786_n;
  wire ffc_787_p;
  wire ffc_787_n;
  wire ffc_788_p;
  wire ffc_788_n;
  wire ffc_789_p;
  wire ffc_789_n;
  wire ffc_790_p;
  wire ffc_790_n;
  wire ffc_791_p;
  wire ffc_791_n;
  wire ffc_792_p;
  wire ffc_792_n;
  wire ffc_793_p;
  wire ffc_793_n;
  wire ffc_794_p;
  wire ffc_794_n;
  wire ffc_795_p;
  wire ffc_795_n;
  wire ffc_796_p;
  wire ffc_796_n;
  wire ffc_797_p;
  wire ffc_797_n;
  wire ffc_798_p;
  wire ffc_798_n;
  wire ffc_799_p;
  wire ffc_799_n;
  wire ffc_800_p;
  wire ffc_800_n;
  wire ffc_801_p;
  wire ffc_801_n;
  wire ffc_802_p;
  wire ffc_802_n;
  wire ffc_803_p;
  wire ffc_803_n;
  wire ffc_804_p;
  wire ffc_804_n;
  wire ffc_805_p;
  wire ffc_805_n;
  wire ffc_806_p;
  wire ffc_806_n;
  wire ffc_807_p;
  wire ffc_807_n;
  wire ffc_808_p;
  wire ffc_808_n;
  wire ffc_809_p;
  wire ffc_809_n;
  wire ffc_810_p;
  wire ffc_810_n;
  wire ffc_811_p;
  wire ffc_811_n;
  wire ffc_812_p;
  wire ffc_812_n;
  wire ffc_813_p;
  wire ffc_813_n;
  wire ffc_814_p;
  wire ffc_814_n;
  wire ffc_815_p;
  wire ffc_815_n;
  wire ffc_816_p;
  wire ffc_816_n;
  wire ffc_817_p;
  wire ffc_817_n;
  wire ffc_818_p;
  wire ffc_818_n;
  wire ffc_819_p;
  wire ffc_819_n;
  wire ffc_820_p;
  wire ffc_820_n;
  wire ffc_821_p;
  wire ffc_821_n;
  wire ffc_822_p;
  wire ffc_822_n;
  wire ffc_823_p;
  wire ffc_823_n;
  wire ffc_824_p;
  wire ffc_824_n;
  wire ffc_825_p;
  wire ffc_825_n;
  wire ffc_826_p;
  wire ffc_826_n;
  wire ffc_827_p;
  wire ffc_827_n;
  wire ffc_828_p;
  wire ffc_828_n;
  wire ffc_829_p;
  wire ffc_829_n;
  wire ffc_830_p;
  wire ffc_830_n;
  wire ffc_831_p;
  wire ffc_831_n;
  wire ffc_832_p;
  wire ffc_832_n;
  wire ffc_833_p;
  wire ffc_833_n;
  wire ffc_834_p;
  wire ffc_834_n;
  wire ffc_835_p;
  wire ffc_835_n;
  wire ffc_836_p;
  wire ffc_836_n;
  wire ffc_837_p;
  wire ffc_837_n;
  wire ffc_838_p;
  wire ffc_838_n;
  wire ffc_839_p;
  wire ffc_839_n;
  wire ffc_840_p;
  wire ffc_840_n;
  wire ffc_841_p;
  wire ffc_841_n;
  wire ffc_842_p;
  wire ffc_842_n;
  wire ffc_843_p;
  wire ffc_843_n;
  wire ffc_844_p;
  wire ffc_844_n;
  wire ffc_845_p;
  wire ffc_845_n;
  wire ffc_846_p;
  wire ffc_846_n;
  wire ffc_847_p;
  wire ffc_847_n;
  wire ffc_848_p;
  wire ffc_848_n;
  wire ffc_849_p;
  wire ffc_849_n;
  wire ffc_850_p;
  wire ffc_850_n;
  wire ffc_851_p;
  wire ffc_851_n;
  wire ffc_852_p;
  wire ffc_852_n;
  wire ffc_853_p;
  wire ffc_853_n;
  wire ffc_854_p;
  wire ffc_854_n;
  wire ffc_855_p;
  wire ffc_855_n;
  wire ffc_856_p;
  wire ffc_856_n;
  wire ffc_857_p;
  wire ffc_857_n;
  wire ffc_858_p;
  wire ffc_858_n;
  wire ffc_859_p;
  wire ffc_859_n;
  wire ffc_860_p;
  wire ffc_860_n;
  wire ffc_861_p;
  wire ffc_861_n;
  wire ffc_862_p;
  wire ffc_862_n;
  wire ffc_863_p;
  wire ffc_863_n;
  wire ffc_864_p;
  wire ffc_864_n;
  wire ffc_865_p;
  wire ffc_865_n;
  wire ffc_866_p;
  wire ffc_866_n;
  wire ffc_867_p;
  wire ffc_867_n;
  wire ffc_868_p;
  wire ffc_868_n;
  wire ffc_869_p;
  wire ffc_869_n;
  wire g1049_p;
  wire g1049_n;
  wire g1050_p;
  wire g1050_n;
  wire g1051_p;
  wire g1051_n;
  wire g1052_p;
  wire g1052_n;
  wire g1053_p;
  wire g1053_n;
  wire g1054_p;
  wire g1054_n;
  wire g1055_p;
  wire g1055_n;
  wire g1056_p;
  wire g1056_n;
  wire g1057_p;
  wire g1057_n;
  wire g1058_p;
  wire g1058_n;
  wire g1059_p;
  wire g1059_n;
  wire g1060_p;
  wire g1060_n;
  wire g1061_p;
  wire g1061_n;
  wire g1062_p;
  wire g1062_n;
  wire g1063_p;
  wire g1063_n;
  wire g1064_p;
  wire g1064_n;
  wire g1065_p;
  wire g1065_n;
  wire g1066_p;
  wire g1066_n;
  wire g1067_p;
  wire g1067_n;
  wire g1068_p;
  wire g1068_n;
  wire g1069_p;
  wire g1069_n;
  wire g1070_p;
  wire g1070_n;
  wire g1071_p;
  wire g1071_n;
  wire g1072_p;
  wire g1072_n;
  wire g1073_p;
  wire g1073_n;
  wire g1074_p;
  wire g1074_n;
  wire g1075_p;
  wire g1075_n;
  wire g1076_p;
  wire g1076_n;
  wire g1077_p;
  wire g1077_n;
  wire g1078_p;
  wire g1078_n;
  wire g1079_p;
  wire g1079_n;
  wire g1080_p;
  wire g1080_n;
  wire g1081_p;
  wire g1081_n;
  wire g1082_p;
  wire g1082_n;
  wire g1083_p;
  wire g1083_n;
  wire g1084_p;
  wire g1084_n;
  wire g1085_p;
  wire g1085_n;
  wire g1086_p;
  wire g1086_n;
  wire g1087_p;
  wire g1087_n;
  wire g1088_p;
  wire g1088_n;
  wire g1089_p;
  wire g1089_n;
  wire g1090_p;
  wire g1090_n;
  wire g1091_p;
  wire g1091_n;
  wire g1092_p;
  wire g1092_n;
  wire g1093_p;
  wire g1093_n;
  wire g1094_p;
  wire g1094_n;
  wire g1095_p;
  wire g1095_n;
  wire g1096_p;
  wire g1096_n;
  wire g1097_p;
  wire g1097_n;
  wire g1098_p;
  wire g1098_n;
  wire g1099_p;
  wire g1099_n;
  wire g1100_p;
  wire g1100_n;
  wire g1101_p;
  wire g1101_n;
  wire g1102_p;
  wire g1102_n;
  wire g1103_p;
  wire g1103_n;
  wire g1104_p;
  wire g1104_n;
  wire g1105_p;
  wire g1105_n;
  wire g1106_p;
  wire g1106_n;
  wire g1107_p;
  wire g1107_n;
  wire g1108_p;
  wire g1108_n;
  wire g1109_p;
  wire g1109_n;
  wire g1110_p;
  wire g1110_n;
  wire g1111_p;
  wire g1111_n;
  wire g1112_p;
  wire g1112_n;
  wire g1113_p;
  wire g1113_n;
  wire g1114_p;
  wire g1114_n;
  wire g1115_p;
  wire g1115_n;
  wire g1116_p;
  wire g1116_n;
  wire g1117_p;
  wire g1117_n;
  wire g1118_p;
  wire g1118_n;
  wire g1119_p;
  wire g1119_n;
  wire g1120_p;
  wire g1120_n;
  wire g1121_p;
  wire g1121_n;
  wire g1122_p;
  wire g1122_n;
  wire g1123_p;
  wire g1123_n;
  wire g1124_p;
  wire g1124_n;
  wire g1125_p;
  wire g1125_n;
  wire g1126_p;
  wire g1126_n;
  wire g1127_p;
  wire g1127_n;
  wire g1128_p;
  wire g1128_n;
  wire g1129_p;
  wire g1129_n;
  wire g1130_p;
  wire g1130_n;
  wire g1131_p;
  wire g1131_n;
  wire g1132_p;
  wire g1132_n;
  wire g1133_p;
  wire g1133_n;
  wire g1134_p;
  wire g1134_n;
  wire g1135_p;
  wire g1135_n;
  wire g1136_p;
  wire g1136_n;
  wire g1137_p;
  wire g1137_n;
  wire g1138_p;
  wire g1138_n;
  wire g1139_p;
  wire g1139_n;
  wire g1140_p;
  wire g1140_n;
  wire g1141_p;
  wire g1141_n;
  wire g1142_p;
  wire g1142_n;
  wire g1143_p;
  wire g1143_n;
  wire g1144_p;
  wire g1144_n;
  wire g1145_p;
  wire g1145_n;
  wire g1146_p;
  wire g1146_n;
  wire g1147_p;
  wire g1147_n;
  wire g1148_p;
  wire g1148_n;
  wire g1149_p;
  wire g1149_n;
  wire g1150_p;
  wire g1150_n;
  wire g1151_p;
  wire g1151_n;
  wire g1152_p;
  wire g1152_n;
  wire g1153_p;
  wire g1153_n;
  wire g1154_p;
  wire g1154_n;
  wire g1155_p;
  wire g1155_n;
  wire g1156_p;
  wire g1156_n;
  wire g1157_p;
  wire g1157_n;
  wire g1158_p;
  wire g1158_n;
  wire g1159_p;
  wire g1159_n;
  wire g1160_p;
  wire g1160_n;
  wire g1161_p;
  wire g1161_n;
  wire g1162_p;
  wire g1162_n;
  wire g1163_p;
  wire g1163_n;
  wire g1164_p;
  wire g1164_n;
  wire g1165_p;
  wire g1165_n;
  wire g1166_p;
  wire g1166_n;
  wire g1167_p;
  wire g1167_n;
  wire g1168_p;
  wire g1168_n;
  wire g1169_p;
  wire g1169_n;
  wire g1170_p;
  wire g1170_n;
  wire g1171_p;
  wire g1171_n;
  wire g1172_p;
  wire g1172_n;
  wire g1173_p;
  wire g1173_n;
  wire g1174_p;
  wire g1174_n;
  wire g1175_p;
  wire g1175_n;
  wire g1176_p;
  wire g1176_n;
  wire g1177_p;
  wire g1177_n;
  wire g1178_p;
  wire g1178_n;
  wire g1179_p;
  wire g1179_n;
  wire g1180_p;
  wire g1180_n;
  wire g1181_p;
  wire g1181_n;
  wire g1182_p;
  wire g1182_n;
  wire g1183_p;
  wire g1183_n;
  wire g1184_p;
  wire g1184_n;
  wire g1185_p;
  wire g1185_n;
  wire g1186_p;
  wire g1186_n;
  wire g1187_p;
  wire g1187_n;
  wire g1188_p;
  wire g1188_n;
  wire g1189_p;
  wire g1189_n;
  wire g1190_p;
  wire g1190_n;
  wire g1191_p;
  wire g1191_n;
  wire g1192_p;
  wire g1192_n;
  wire g1193_p;
  wire g1193_n;
  wire g1194_p;
  wire g1194_n;
  wire g1195_p;
  wire g1195_n;
  wire g1196_p;
  wire g1196_n;
  wire g1197_p;
  wire g1197_n;
  wire g1198_p;
  wire g1198_n;
  wire g1199_p;
  wire g1199_n;
  wire g1200_p;
  wire g1200_n;
  wire g1201_p;
  wire g1201_n;
  wire g1202_p;
  wire g1202_n;
  wire g1203_p;
  wire g1203_n;
  wire g1204_p;
  wire g1204_n;
  wire g1205_p;
  wire g1205_n;
  wire g1206_p;
  wire g1206_n;
  wire g1207_p;
  wire g1207_n;
  wire g1208_p;
  wire g1208_n;
  wire g1209_p;
  wire g1209_n;
  wire g1210_p;
  wire g1210_n;
  wire g1211_p;
  wire g1211_n;
  wire g1212_p;
  wire g1212_n;
  wire g1213_p;
  wire g1213_n;
  wire g1214_p;
  wire g1214_n;
  wire g1215_p;
  wire g1215_n;
  wire g1216_p;
  wire g1216_n;
  wire g1217_p;
  wire g1217_n;
  wire g1218_p;
  wire g1218_n;
  wire g1219_p;
  wire g1219_n;
  wire g1220_p;
  wire g1220_n;
  wire g1221_p;
  wire g1221_n;
  wire g1222_p;
  wire g1222_n;
  wire g1223_p;
  wire g1223_n;
  wire g1224_p;
  wire g1224_n;
  wire g1225_p;
  wire g1225_n;
  wire g1226_p;
  wire g1226_n;
  wire g1227_p;
  wire g1227_n;
  wire g1228_p;
  wire g1228_n;
  wire g1229_p;
  wire g1229_n;
  wire g1230_p;
  wire g1230_n;
  wire g1231_p;
  wire g1231_n;
  wire g1232_p;
  wire g1232_n;
  wire g1233_p;
  wire g1233_n;
  wire g1234_p;
  wire g1234_n;
  wire g1235_p;
  wire g1235_n;
  wire g1236_p;
  wire g1236_n;
  wire g1237_p;
  wire g1237_n;
  wire g1238_p;
  wire g1238_n;
  wire g1239_p;
  wire g1239_n;
  wire g1240_p;
  wire g1240_n;
  wire g1241_p;
  wire g1241_n;
  wire g1242_p;
  wire g1242_n;
  wire g1243_p;
  wire g1243_n;
  wire g1244_p;
  wire g1244_n;
  wire g1245_p;
  wire g1245_n;
  wire g1246_p;
  wire g1246_n;
  wire g1247_p;
  wire g1247_n;
  wire g1248_p;
  wire g1248_n;
  wire g1249_p;
  wire g1249_n;
  wire g1250_p;
  wire g1250_n;
  wire g1251_p;
  wire g1251_n;
  wire g1252_p;
  wire g1252_n;
  wire g1253_p;
  wire g1253_n;
  wire g1254_p;
  wire g1254_n;
  wire g1255_p;
  wire g1255_n;
  wire g1256_p;
  wire g1256_n;
  wire g1257_p;
  wire g1257_n;
  wire g1258_p;
  wire g1258_n;
  wire g1259_p;
  wire g1259_n;
  wire g1260_p;
  wire g1260_n;
  wire g1261_p;
  wire g1261_n;
  wire g1262_p;
  wire g1262_n;
  wire g1263_p;
  wire g1263_n;
  wire g1264_p;
  wire g1264_n;
  wire g1265_p;
  wire g1265_n;
  wire g1266_p;
  wire g1266_n;
  wire g1267_p;
  wire g1267_n;
  wire g1268_p;
  wire g1268_n;
  wire g1269_p;
  wire g1269_n;
  wire g1270_p;
  wire g1270_n;
  wire g1271_p;
  wire g1271_n;
  wire g1272_p;
  wire g1272_n;
  wire g1273_p;
  wire g1273_n;
  wire g1274_p;
  wire g1274_n;
  wire g1275_p;
  wire g1275_n;
  wire g1276_p;
  wire g1276_n;
  wire g1277_p;
  wire g1277_n;
  wire g1278_p;
  wire g1278_n;
  wire g1279_p;
  wire g1279_n;
  wire g1280_p;
  wire g1280_n;
  wire g1281_p;
  wire g1281_n;
  wire g1282_p;
  wire g1282_n;
  wire g1283_p;
  wire g1283_n;
  wire g1284_p;
  wire g1284_n;
  wire g1285_p;
  wire g1285_n;
  wire g1286_p;
  wire g1286_n;
  wire g1287_p;
  wire g1287_n;
  wire g1288_p;
  wire g1288_n;
  wire g1289_p;
  wire g1289_n;
  wire g1290_p;
  wire g1290_n;
  wire g1291_p;
  wire g1291_n;
  wire g1292_p;
  wire g1292_n;
  wire g1293_p;
  wire g1293_n;
  wire g1294_p;
  wire g1294_n;
  wire g1295_p;
  wire g1295_n;
  wire g1296_p;
  wire g1296_n;
  wire g1297_p;
  wire g1297_n;
  wire g1298_p;
  wire g1298_n;
  wire g1299_p;
  wire g1299_n;
  wire g1300_p;
  wire g1300_n;
  wire g1301_p;
  wire g1301_n;
  wire g1302_p;
  wire g1302_n;
  wire g1303_p;
  wire g1303_n;
  wire g1304_p;
  wire g1304_n;
  wire g1305_p;
  wire g1305_n;
  wire g1306_p;
  wire g1306_n;
  wire g1307_p;
  wire g1307_n;
  wire g1308_p;
  wire g1308_n;
  wire g1309_p;
  wire g1309_n;
  wire g1310_p;
  wire g1310_n;
  wire g1311_p;
  wire g1311_n;
  wire g1312_p;
  wire g1312_n;
  wire g1313_p;
  wire g1313_n;
  wire g1314_p;
  wire g1314_n;
  wire g1315_p;
  wire g1315_n;
  wire g1316_p;
  wire g1316_n;
  wire g1317_p;
  wire g1317_n;
  wire g1318_p;
  wire g1318_n;
  wire g1319_p;
  wire g1319_n;
  wire g1320_p;
  wire g1320_n;
  wire g1321_p;
  wire g1321_n;
  wire g1322_p;
  wire g1322_n;
  wire g1323_p;
  wire g1323_n;
  wire g1324_p;
  wire g1324_n;
  wire g1325_p;
  wire g1325_n;
  wire g1326_p;
  wire g1326_n;
  wire g1327_p;
  wire g1327_n;
  wire g1328_p;
  wire g1328_n;
  wire g1329_p;
  wire g1329_n;
  wire g1330_p;
  wire g1330_n;
  wire g1331_p;
  wire g1331_n;
  wire g1332_p;
  wire g1332_n;
  wire g1333_p;
  wire g1333_n;
  wire g1334_p;
  wire g1334_n;
  wire g1335_p;
  wire g1335_n;
  wire g1336_p;
  wire g1336_n;
  wire g1337_p;
  wire g1337_n;
  wire g1338_p;
  wire g1338_n;
  wire g1339_p;
  wire g1339_n;
  wire g1340_p;
  wire g1340_n;
  wire g1341_p;
  wire g1341_n;
  wire g1342_p;
  wire g1342_n;
  wire g1343_p;
  wire g1343_n;
  wire g1344_p;
  wire g1344_n;
  wire g1345_p;
  wire g1345_n;
  wire g1346_p;
  wire g1346_n;
  wire g1347_p;
  wire g1347_n;
  wire g1348_p;
  wire g1348_n;
  wire g1349_p;
  wire g1349_n;
  wire g1350_p;
  wire g1350_n;
  wire g1351_p;
  wire g1351_n;
  wire g1352_p;
  wire g1352_n;
  wire g1353_p;
  wire g1353_n;
  wire g1354_p;
  wire g1354_n;
  wire g1355_p;
  wire g1355_n;
  wire g1356_p;
  wire g1356_n;
  wire g1357_p;
  wire g1357_n;
  wire g1358_p;
  wire g1358_n;
  wire g1359_p;
  wire g1359_n;
  wire g1360_p;
  wire g1360_n;
  wire g1361_p;
  wire g1361_n;
  wire g1362_p;
  wire g1362_n;
  wire g1363_p;
  wire g1363_n;
  wire g1364_p;
  wire g1364_n;
  wire g1365_p;
  wire g1365_n;
  wire g1366_p;
  wire g1366_n;
  wire g1367_p;
  wire g1367_n;
  wire g1368_p;
  wire g1368_n;
  wire g1369_p;
  wire g1369_n;
  wire g1370_p;
  wire g1370_n;
  wire g1371_p;
  wire g1371_n;
  wire g1372_p;
  wire g1372_n;
  wire g1373_p;
  wire g1373_n;
  wire g1374_p;
  wire g1374_n;
  wire g1375_p;
  wire g1375_n;
  wire g1376_p;
  wire g1376_n;
  wire g1377_p;
  wire g1377_n;
  wire g1378_p;
  wire g1378_n;
  wire g1379_p;
  wire g1379_n;
  wire g1380_p;
  wire g1380_n;
  wire g1381_p;
  wire g1381_n;
  wire g1382_p;
  wire g1382_n;
  wire g1383_p;
  wire g1383_n;
  wire g1384_p;
  wire g1384_n;
  wire g1385_p;
  wire g1385_n;
  wire g1386_p;
  wire g1386_n;
  wire g1387_p;
  wire g1387_n;
  wire g1388_p;
  wire g1388_n;
  wire g1389_p;
  wire g1389_n;
  wire g1390_p;
  wire g1390_n;
  wire g1391_p;
  wire g1391_n;
  wire g1392_p;
  wire g1392_n;
  wire g1393_p;
  wire g1393_n;
  wire g1394_p;
  wire g1394_n;
  wire g1395_p;
  wire g1395_n;
  wire g1396_p;
  wire g1396_n;
  wire g1397_p;
  wire g1397_n;
  wire g1398_p;
  wire g1398_n;
  wire g1399_p;
  wire g1399_n;
  wire g1400_p;
  wire g1400_n;
  wire g1401_p;
  wire g1401_n;
  wire g1402_p;
  wire g1402_n;
  wire g1403_p;
  wire g1403_n;
  wire g1404_p;
  wire g1404_n;
  wire g1405_p;
  wire g1405_n;
  wire g1406_p;
  wire g1406_n;
  wire g1407_p;
  wire g1407_n;
  wire g1408_p;
  wire g1408_n;
  wire g1409_p;
  wire g1409_n;
  wire g1410_p;
  wire g1410_n;
  wire g1411_p;
  wire g1411_n;
  wire g1412_p;
  wire g1412_n;
  wire g1413_p;
  wire g1413_n;
  wire g1414_p;
  wire g1414_n;
  wire g1415_p;
  wire g1415_n;
  wire g1416_p;
  wire g1416_n;
  wire g1417_p;
  wire g1417_n;
  wire g1418_p;
  wire g1418_n;
  wire g1419_p;
  wire g1419_n;
  wire g1420_p;
  wire g1420_n;
  wire g1421_p;
  wire g1421_n;
  wire g1422_p;
  wire g1422_n;
  wire g1423_p;
  wire g1423_n;
  wire g1424_p;
  wire g1424_n;
  wire g1425_p;
  wire g1425_n;
  wire g1426_p;
  wire g1426_n;
  wire g1427_p;
  wire g1427_n;
  wire g1428_p;
  wire g1428_n;
  wire g1429_p;
  wire g1429_n;
  wire g1430_p;
  wire g1430_n;
  wire g1431_p;
  wire g1431_n;
  wire g1432_p;
  wire g1432_n;
  wire g1433_p;
  wire g1433_n;
  wire g1434_p;
  wire g1434_n;
  wire g1435_p;
  wire g1435_n;
  wire g1436_p;
  wire g1436_n;
  wire g1437_p;
  wire g1437_n;
  wire g1438_p;
  wire g1438_n;
  wire g1439_p;
  wire g1439_n;
  wire g1440_p;
  wire g1440_n;
  wire g1441_p;
  wire g1441_n;
  wire g1442_p;
  wire g1442_n;
  wire g1443_p;
  wire g1443_n;
  wire g1444_p;
  wire g1444_n;
  wire g1445_p;
  wire g1445_n;
  wire g1446_p;
  wire g1446_n;
  wire g1447_p;
  wire g1447_n;
  wire g1448_p;
  wire g1448_n;
  wire g1449_p;
  wire g1449_n;
  wire g1450_p;
  wire g1450_n;
  wire g1451_p;
  wire g1451_n;
  wire g1452_p;
  wire g1452_n;
  wire g1453_p;
  wire g1453_n;
  wire g1454_p;
  wire g1454_n;
  wire g1455_p;
  wire g1455_n;
  wire g1456_p;
  wire g1456_n;
  wire g1457_p;
  wire g1457_n;
  wire g1458_p;
  wire g1458_n;
  wire g1459_p;
  wire g1459_n;
  wire g1460_p;
  wire g1460_n;
  wire g1461_p;
  wire g1461_n;
  wire g1462_p;
  wire g1462_n;
  wire g1463_p;
  wire g1463_n;
  wire g1464_p;
  wire g1464_n;
  wire g1465_p;
  wire g1465_n;
  wire g1466_p;
  wire g1466_n;
  wire g1467_p;
  wire g1467_n;
  wire g1468_p;
  wire g1468_n;
  wire g1469_p;
  wire g1469_n;
  wire g1470_p;
  wire g1470_n;
  wire g1471_p;
  wire g1471_n;
  wire g1472_p;
  wire g1472_n;
  wire g1473_p;
  wire g1473_n;
  wire g1474_p;
  wire g1474_n;
  wire g1475_p;
  wire g1475_n;
  wire g1476_p;
  wire g1476_n;
  wire g1477_p;
  wire g1477_n;
  wire g1478_p;
  wire g1478_n;
  wire g1479_p;
  wire g1479_n;
  wire g1480_p;
  wire g1480_n;
  wire g1481_p;
  wire g1481_n;
  wire g1482_p;
  wire g1482_n;
  wire g1483_p;
  wire g1483_n;
  wire g1484_p;
  wire g1484_n;
  wire g1485_p;
  wire g1485_n;
  wire g1486_p;
  wire g1486_n;
  wire g1487_p;
  wire g1487_n;
  wire g1488_p;
  wire g1488_n;
  wire g1489_p;
  wire g1489_n;
  wire g1490_p;
  wire g1490_n;
  wire g1491_p;
  wire g1491_n;
  wire g1492_p;
  wire g1492_n;
  wire g1493_p;
  wire g1493_n;
  wire g1494_p;
  wire g1494_n;
  wire g1495_p;
  wire g1495_n;
  wire g1496_p;
  wire g1496_n;
  wire g1497_p;
  wire g1497_n;
  wire g1498_p;
  wire g1498_n;
  wire g1499_p;
  wire g1499_n;
  wire g1500_p;
  wire g1500_n;
  wire g1501_p;
  wire g1501_n;
  wire g1502_p;
  wire g1502_n;
  wire g1503_p;
  wire g1503_n;
  wire g1504_p;
  wire g1504_n;
  wire g1505_p;
  wire g1505_n;
  wire g1506_p;
  wire g1506_n;
  wire g1507_p;
  wire g1507_n;
  wire g1508_p;
  wire g1508_n;
  wire g1509_p;
  wire g1509_n;
  wire g1510_p;
  wire g1510_n;
  wire g1511_p;
  wire g1511_n;
  wire g1512_p;
  wire g1512_n;
  wire g1513_p;
  wire g1513_n;
  wire g1514_p;
  wire g1514_n;
  wire g1515_p;
  wire g1515_n;
  wire g1516_p;
  wire g1516_n;
  wire g1517_p;
  wire g1517_n;
  wire g1518_p;
  wire g1518_n;
  wire g1519_p;
  wire g1519_n;
  wire g1520_p;
  wire g1520_n;
  wire g1521_p;
  wire g1521_n;
  wire g1522_p;
  wire g1522_n;
  wire g1523_p;
  wire g1523_n;
  wire g1524_p;
  wire g1524_n;
  wire g1525_p;
  wire g1525_n;
  wire g1526_p;
  wire g1526_n;
  wire g1527_p;
  wire g1527_n;
  wire g1528_p;
  wire g1528_n;
  wire g1529_p;
  wire g1529_n;
  wire g1530_p;
  wire g1530_n;
  wire g1531_p;
  wire g1531_n;
  wire g1532_p;
  wire g1532_n;
  wire g1533_p;
  wire g1533_n;
  wire g1534_p;
  wire g1534_n;
  wire g1535_p;
  wire g1535_n;
  wire g1536_p;
  wire g1536_n;
  wire g1537_p;
  wire g1537_n;
  wire g1538_p;
  wire g1538_n;
  wire g1539_p;
  wire g1539_n;
  wire g1540_p;
  wire g1540_n;
  wire g1541_p;
  wire g1541_n;
  wire g1542_p;
  wire g1542_n;
  wire g1543_p;
  wire g1543_n;
  wire g1544_p;
  wire g1544_n;
  wire g1545_p;
  wire g1545_n;
  wire g1546_p;
  wire g1546_n;
  wire g1547_p;
  wire g1547_n;
  wire g1548_p;
  wire g1548_n;
  wire g1549_p;
  wire g1549_n;
  wire g1550_p;
  wire g1550_n;
  wire g1551_p;
  wire g1551_n;
  wire g1552_p;
  wire g1552_n;
  wire g1553_p;
  wire g1553_n;
  wire g1554_p;
  wire g1554_n;
  wire g1555_p;
  wire g1555_n;
  wire g1556_p;
  wire g1556_n;
  wire g1557_p;
  wire g1557_n;
  wire g1558_p;
  wire g1558_n;
  wire g1559_p;
  wire g1559_n;
  wire g1560_p;
  wire g1560_n;
  wire g1561_p;
  wire g1561_n;
  wire g1562_p;
  wire g1562_n;
  wire g1563_p;
  wire g1563_n;
  wire g1564_p;
  wire g1564_n;
  wire g1565_p;
  wire g1565_n;
  wire g1566_p;
  wire g1566_n;
  wire g1567_p;
  wire g1567_n;
  wire g1568_p;
  wire g1568_n;
  wire g1569_p;
  wire g1569_n;
  wire g1570_p;
  wire g1570_n;
  wire g1571_p;
  wire g1571_n;
  wire g1572_p;
  wire g1572_n;
  wire g1573_p;
  wire g1573_n;
  wire g1574_p;
  wire g1574_n;
  wire g1575_p;
  wire g1575_n;
  wire g1576_p;
  wire g1576_n;
  wire g1577_p;
  wire g1577_n;
  wire g1578_p;
  wire g1578_n;
  wire g1579_p;
  wire g1579_n;
  wire g1580_p;
  wire g1580_n;
  wire g1581_p;
  wire g1581_n;
  wire g1582_p;
  wire g1582_n;
  wire g1583_p;
  wire g1583_n;
  wire g1584_p;
  wire g1584_n;
  wire g1585_p;
  wire g1585_n;
  wire g1586_p;
  wire g1586_n;
  wire g1587_p;
  wire g1587_n;
  wire g1588_p;
  wire g1588_n;
  wire g1589_p;
  wire g1589_n;
  wire g1590_p;
  wire g1590_n;
  wire g1591_p;
  wire g1591_n;
  wire g1592_p;
  wire g1592_n;
  wire g1593_p;
  wire g1593_n;
  wire g1594_p;
  wire g1594_n;
  wire g1595_p;
  wire g1595_n;
  wire g1596_p;
  wire g1596_n;
  wire g1597_p;
  wire g1597_n;
  wire g1598_p;
  wire g1598_n;
  wire g1599_p;
  wire g1599_n;
  wire g1600_p;
  wire g1600_n;
  wire g1601_p;
  wire g1601_n;
  wire g1602_p;
  wire g1602_n;
  wire g1603_p;
  wire g1603_n;
  wire g1604_p;
  wire g1604_n;
  wire g1605_p;
  wire g1605_n;
  wire g1606_p;
  wire g1606_n;
  wire g1607_p;
  wire g1607_n;
  wire g1608_p;
  wire g1608_n;
  wire g1609_p;
  wire g1609_n;
  wire g1610_p;
  wire g1610_n;
  wire g1611_p;
  wire g1611_n;
  wire g1612_p;
  wire g1612_n;
  wire g1613_p;
  wire g1613_n;
  wire g1614_p;
  wire g1614_n;
  wire g1615_p;
  wire g1615_n;
  wire g1616_p;
  wire g1616_n;
  wire g1617_p;
  wire g1617_n;
  wire g1618_p;
  wire g1618_n;
  wire g1619_p;
  wire g1619_n;
  wire g1620_p;
  wire g1620_n;
  wire g1621_p;
  wire g1621_n;
  wire g1622_p;
  wire g1622_n;
  wire g1623_p;
  wire g1623_n;
  wire g1624_p;
  wire g1624_n;
  wire g1625_p;
  wire g1625_n;
  wire g1626_p;
  wire g1626_n;
  wire g1627_p;
  wire g1627_n;
  wire g1628_p;
  wire g1628_n;
  wire g1629_p;
  wire g1629_n;
  wire g1630_p;
  wire g1630_n;
  wire g1631_p;
  wire g1631_n;
  wire g1632_p;
  wire g1632_n;
  wire g1633_p;
  wire g1633_n;
  wire g1634_p;
  wire g1634_n;
  wire g1635_p;
  wire g1635_n;
  wire g1636_p;
  wire g1636_n;
  wire g1637_p;
  wire g1637_n;
  wire g1638_p;
  wire g1638_n;
  wire g1639_p;
  wire g1639_n;
  wire g1640_p;
  wire g1640_n;
  wire g1641_p;
  wire g1641_n;
  wire g1642_p;
  wire g1642_n;
  wire g1643_p;
  wire g1643_n;
  wire g1644_p;
  wire g1644_n;
  wire g1645_p;
  wire g1645_n;
  wire g1646_p;
  wire g1646_n;
  wire g1647_p;
  wire g1647_n;
  wire g1648_p;
  wire g1648_n;
  wire g1649_p;
  wire g1649_n;
  wire g1650_p;
  wire g1650_n;
  wire g1651_p;
  wire g1651_n;
  wire g1652_p;
  wire g1652_n;
  wire g1653_p;
  wire g1653_n;
  wire g1654_p;
  wire g1654_n;
  wire g1655_p;
  wire g1655_n;
  wire g1656_p;
  wire g1656_n;
  wire g1657_p;
  wire g1657_n;
  wire g1658_p;
  wire g1658_n;
  wire g1659_p;
  wire g1659_n;
  wire g1660_p;
  wire g1660_n;
  wire g1661_p;
  wire g1661_n;
  wire g1662_p;
  wire g1662_n;
  wire g1663_p;
  wire g1663_n;
  wire g1664_p;
  wire g1664_n;
  wire g1665_p;
  wire g1665_n;
  wire g1666_p;
  wire g1666_n;
  wire g1667_p;
  wire g1667_n;
  wire g1668_p;
  wire g1668_n;
  wire g1669_p;
  wire g1669_n;
  wire g1670_p;
  wire g1670_n;
  wire g1671_p;
  wire g1671_n;
  wire g1672_p;
  wire g1672_n;
  wire g1673_p;
  wire g1673_n;
  wire g1674_p;
  wire g1674_n;
  wire g1675_p;
  wire g1675_n;
  wire g1676_p;
  wire g1676_n;
  wire g1677_p;
  wire g1677_n;
  wire g1678_p;
  wire g1678_n;
  wire g1679_p;
  wire g1679_n;
  wire g1680_p;
  wire g1680_n;
  wire g1681_p;
  wire g1681_n;
  wire g1682_p;
  wire g1682_n;
  wire g1683_p;
  wire g1683_n;
  wire g1684_p;
  wire g1684_n;
  wire g1685_p;
  wire g1685_n;
  wire g1686_p;
  wire g1686_n;
  wire g1687_p;
  wire g1687_n;
  wire g1688_p;
  wire g1688_n;
  wire g1689_p;
  wire g1689_n;
  wire g1690_p;
  wire g1690_n;
  wire g1691_p;
  wire g1691_n;
  wire g1692_p;
  wire g1692_n;
  wire g1693_p;
  wire g1693_n;
  wire g1694_p;
  wire g1694_n;
  wire g1695_p;
  wire g1695_n;
  wire g1696_p;
  wire g1696_n;
  wire g1697_p;
  wire g1697_n;
  wire g1698_p;
  wire g1698_n;
  wire g1699_p;
  wire g1699_n;
  wire g1700_p;
  wire g1700_n;
  wire g1701_p;
  wire g1701_n;
  wire g1702_p;
  wire g1702_n;
  wire g1703_p;
  wire g1703_n;
  wire g1704_p;
  wire g1704_n;
  wire g1705_p;
  wire g1705_n;
  wire g1706_p;
  wire g1706_n;
  wire g1707_p;
  wire g1707_n;
  wire g1708_p;
  wire g1708_n;
  wire g1709_p;
  wire g1709_n;
  wire g1710_p;
  wire g1710_n;
  wire g1711_p;
  wire g1711_n;
  wire g1712_p;
  wire g1712_n;
  wire g1713_p;
  wire g1713_n;
  wire g1714_p;
  wire g1714_n;
  wire g1715_p;
  wire g1715_n;
  wire g1716_p;
  wire g1716_n;
  wire g1717_p;
  wire g1717_n;
  wire g1718_p;
  wire g1718_n;
  wire g1719_p;
  wire g1719_n;
  wire g1720_p;
  wire g1720_n;
  wire g1721_p;
  wire g1721_n;
  wire g1722_p;
  wire g1722_n;
  wire g1723_p;
  wire g1723_n;
  wire g1724_p;
  wire g1724_n;
  wire g1725_p;
  wire g1725_n;
  wire g1726_p;
  wire g1726_n;
  wire g1727_p;
  wire g1727_n;
  wire g1728_p;
  wire g1728_n;
  wire g1729_p;
  wire g1729_n;
  wire g1730_p;
  wire g1730_n;
  wire g1731_p;
  wire g1731_n;
  wire g1732_p;
  wire g1732_n;
  wire g1733_p;
  wire g1733_n;
  wire g1734_p;
  wire g1734_n;
  wire g1735_p;
  wire g1735_n;
  wire g1736_p;
  wire g1736_n;
  wire g1737_p;
  wire g1737_n;
  wire g1738_p;
  wire g1738_n;
  wire g1739_p;
  wire g1739_n;
  wire g1740_p;
  wire g1740_n;
  wire g1741_p;
  wire g1741_n;
  wire g1742_p;
  wire g1742_n;
  wire g1743_p;
  wire g1743_n;
  wire g1744_p;
  wire g1744_n;
  wire g1745_p;
  wire g1745_n;
  wire g1746_p;
  wire g1746_n;
  wire g1747_p;
  wire g1747_n;
  wire g1748_p;
  wire g1748_n;
  wire g1749_p;
  wire g1749_n;
  wire g1750_p;
  wire g1750_n;
  wire g1751_p;
  wire g1751_n;
  wire g1752_p;
  wire g1752_n;
  wire g1753_p;
  wire g1753_n;
  wire g1754_p;
  wire g1754_n;
  wire g1755_p;
  wire g1755_n;
  wire g1756_p;
  wire g1756_n;
  wire g1757_p;
  wire g1757_n;
  wire g1758_p;
  wire g1758_n;
  wire g1759_p;
  wire g1759_n;
  wire g1760_p;
  wire g1760_n;
  wire g1761_p;
  wire g1761_n;
  wire g1762_p;
  wire g1762_n;
  wire g1763_p;
  wire g1763_n;
  wire g1764_p;
  wire g1764_n;
  wire g1765_p;
  wire g1765_n;
  wire g1766_p;
  wire g1766_n;
  wire g1767_p;
  wire g1767_n;
  wire g1768_p;
  wire g1768_n;
  wire g1769_p;
  wire g1769_n;
  wire g1770_p;
  wire g1770_n;
  wire g1771_p;
  wire g1771_n;
  wire g1772_p;
  wire g1772_n;
  wire g1773_p;
  wire g1773_n;
  wire g1774_p;
  wire g1774_n;
  wire g1775_p;
  wire g1775_n;
  wire g1776_p;
  wire g1776_n;
  wire g1777_p;
  wire g1777_n;
  wire g1778_p;
  wire g1778_n;
  wire g1779_p;
  wire g1779_n;
  wire g1780_p;
  wire g1780_n;
  wire g1781_p;
  wire g1781_n;
  wire g1782_p;
  wire g1782_n;
  wire g1783_p;
  wire g1783_n;
  wire g1784_p;
  wire g1784_n;
  wire g1785_p;
  wire g1785_n;
  wire g1786_p;
  wire g1786_n;
  wire g1787_p;
  wire g1787_n;
  wire g1788_p;
  wire g1788_n;
  wire g1789_p;
  wire g1789_n;
  wire g1790_p;
  wire g1790_n;
  wire g1791_p;
  wire g1791_n;
  wire g1792_p;
  wire g1792_n;
  wire g1793_p;
  wire g1793_n;
  wire g1794_p;
  wire g1794_n;
  wire g1795_p;
  wire g1795_n;
  wire g1796_p;
  wire g1796_n;
  wire g1797_p;
  wire g1797_n;
  wire g1798_p;
  wire g1798_n;
  wire g1799_p;
  wire g1799_n;
  wire g1800_p;
  wire g1800_n;
  wire g1801_p;
  wire g1801_n;
  wire g1802_p;
  wire g1802_n;
  wire g1803_p;
  wire g1803_n;
  wire g1804_p;
  wire g1804_n;
  wire g1805_p;
  wire g1805_n;
  wire g1806_p;
  wire g1806_n;
  wire g1807_p;
  wire g1807_n;
  wire g1808_p;
  wire g1808_n;
  wire g1809_p;
  wire g1809_n;
  wire g1810_p;
  wire g1810_n;
  wire g1811_p;
  wire g1811_n;
  wire g1812_p;
  wire g1812_n;
  wire g1813_p;
  wire g1813_n;
  wire g1814_p;
  wire g1814_n;
  wire g1815_p;
  wire g1815_n;
  wire g1816_p;
  wire g1816_n;
  wire g1817_p;
  wire g1817_n;
  wire g1818_p;
  wire g1818_n;
  wire g1819_p;
  wire g1819_n;
  wire g1820_p;
  wire g1820_n;
  wire g1821_p;
  wire g1821_n;
  wire g1822_p;
  wire g1822_n;
  wire g1823_p;
  wire g1823_n;
  wire g1824_p;
  wire g1824_n;
  wire g1825_p;
  wire g1825_n;
  wire g1826_p;
  wire g1826_n;
  wire g1827_p;
  wire g1827_n;
  wire g1828_p;
  wire g1828_n;
  wire g1829_p;
  wire g1829_n;
  wire g1830_p;
  wire g1830_n;
  wire g1831_p;
  wire g1831_n;
  wire g1832_p;
  wire g1832_n;
  wire g1833_p;
  wire g1833_n;
  wire g1834_p;
  wire g1834_n;
  wire g1835_p;
  wire g1835_n;
  wire g1836_p;
  wire g1836_n;
  wire g1837_p;
  wire g1837_n;
  wire g1838_p;
  wire g1838_n;
  wire g1839_p;
  wire g1839_n;
  wire g1840_p;
  wire g1840_n;
  wire g1841_p;
  wire g1841_n;
  wire g1842_p;
  wire g1842_n;
  wire g1843_p;
  wire g1843_n;
  wire g1844_p;
  wire g1844_n;
  wire g1845_p;
  wire g1845_n;
  wire g1846_p;
  wire g1846_n;
  wire g1847_p;
  wire g1847_n;
  wire g1848_p;
  wire g1848_n;
  wire g1849_p;
  wire g1849_n;
  wire g1850_p;
  wire g1850_n;
  wire g1851_p;
  wire g1851_n;
  wire g1852_p;
  wire g1852_n;
  wire g1853_p;
  wire g1853_n;
  wire g1854_p;
  wire g1854_n;
  wire g1855_p;
  wire g1855_n;
  wire g1856_p;
  wire g1856_n;
  wire g1857_p;
  wire g1857_n;
  wire g1858_p;
  wire g1858_n;
  wire g1859_p;
  wire g1859_n;
  wire g1860_p;
  wire g1860_n;
  wire g1861_p;
  wire g1861_n;
  wire g1862_p;
  wire g1862_n;
  wire g1863_p;
  wire g1863_n;
  wire g1864_p;
  wire g1864_n;
  wire g1865_p;
  wire g1865_n;
  wire g1866_p;
  wire g1866_n;
  wire g1867_p;
  wire g1867_n;
  wire g1868_p;
  wire g1868_n;
  wire g1869_p;
  wire g1869_n;
  wire g1870_p;
  wire g1870_n;
  wire g1871_p;
  wire g1871_n;
  wire g1872_p;
  wire g1872_n;
  wire g1873_p;
  wire g1873_n;
  wire g1874_p;
  wire g1874_n;
  wire g1875_p;
  wire g1875_n;
  wire g1876_p;
  wire g1876_n;
  wire g1877_p;
  wire g1877_n;
  wire g1878_p;
  wire g1878_n;
  wire g1879_p;
  wire g1879_n;
  wire g1880_p;
  wire g1880_n;
  wire g1881_p;
  wire g1881_n;
  wire g1882_p;
  wire g1882_n;
  wire g1883_p;
  wire g1883_n;
  wire g1884_p;
  wire g1884_n;
  wire g1885_p;
  wire g1885_n;
  wire g1886_p;
  wire g1886_n;
  wire g1887_p;
  wire g1887_n;
  wire g1888_p;
  wire g1888_n;
  wire g1889_p;
  wire g1889_n;
  wire g1890_p;
  wire g1890_n;
  wire g1891_p;
  wire g1891_n;
  wire g1892_p;
  wire g1892_n;
  wire g1893_p;
  wire g1893_n;
  wire g1894_p;
  wire g1894_n;
  wire g1895_p;
  wire g1895_n;
  wire g1896_p;
  wire g1896_n;
  wire g1897_p;
  wire g1897_n;
  wire g1898_p;
  wire g1898_n;
  wire g1899_p;
  wire g1899_n;
  wire g1900_p;
  wire g1900_n;
  wire g1901_p;
  wire g1901_n;
  wire g1902_p;
  wire g1902_n;
  wire g1903_p;
  wire g1903_n;
  wire g1904_p;
  wire g1904_n;
  wire g1905_p;
  wire g1905_n;
  wire g1906_p;
  wire g1906_n;
  wire g1907_p;
  wire g1907_n;
  wire g1908_p;
  wire g1908_n;
  wire g1909_p;
  wire g1909_n;
  wire g1910_p;
  wire g1910_n;
  wire g1911_p;
  wire g1911_n;
  wire g1912_p;
  wire g1912_n;
  wire g1913_p;
  wire g1913_n;
  wire g1914_p;
  wire g1914_n;
  wire g1915_p;
  wire g1915_n;
  wire g1916_p;
  wire g1916_n;
  wire g1917_p;
  wire g1917_n;
  wire g1918_p;
  wire g1918_n;
  wire g1919_p;
  wire g1919_n;
  wire g1920_p;
  wire g1920_n;
  wire g1921_p;
  wire g1921_n;
  wire g1922_p;
  wire g1922_n;
  wire g1923_p;
  wire g1923_n;
  wire g1924_p;
  wire g1924_n;
  wire g1925_p;
  wire g1925_n;
  wire g1926_p;
  wire g1926_n;
  wire g1927_p;
  wire g1927_n;
  wire g1928_p;
  wire g1928_n;
  wire g1929_p;
  wire g1929_n;
  wire g1930_p;
  wire g1930_n;
  wire g1931_p;
  wire g1931_n;
  wire g1932_p;
  wire g1932_n;
  wire g1933_p;
  wire g1933_n;
  wire g1934_p;
  wire g1934_n;
  wire g1935_p;
  wire g1935_n;
  wire g1936_p;
  wire g1936_n;
  wire g1937_p;
  wire g1937_n;
  wire g1938_p;
  wire g1938_n;
  wire g1939_p;
  wire g1939_n;
  wire g1940_p;
  wire g1940_n;
  wire g1941_p;
  wire g1941_n;
  wire g1942_p;
  wire g1942_n;
  wire g1943_p;
  wire g1943_n;
  wire g1944_p;
  wire g1944_n;
  wire g1945_p;
  wire g1945_n;
  wire g1946_p;
  wire g1946_n;
  wire g1947_p;
  wire g1947_n;
  wire g1948_p;
  wire g1948_n;
  wire g1949_p;
  wire g1949_n;
  wire g1950_p;
  wire g1950_n;
  wire g1951_p;
  wire g1951_n;
  wire g1952_p;
  wire g1952_n;
  wire g1953_p;
  wire g1953_n;
  wire g1954_p;
  wire g1954_n;
  wire g1955_p;
  wire g1955_n;
  wire g1956_p;
  wire g1956_n;
  wire g1957_p;
  wire g1957_n;
  wire g1958_p;
  wire g1958_n;
  wire g1959_p;
  wire g1959_n;
  wire g1960_p;
  wire g1960_n;
  wire g1961_p;
  wire g1961_n;
  wire g1962_p;
  wire g1962_n;
  wire g1963_p;
  wire g1963_n;
  wire g1964_p;
  wire g1964_n;
  wire g1965_p;
  wire g1965_n;
  wire g1966_p;
  wire g1966_n;
  wire g1967_p;
  wire g1967_n;
  wire g1968_p;
  wire g1968_n;
  wire g1969_p;
  wire g1969_n;
  wire g1970_p;
  wire g1970_n;
  wire g1971_p;
  wire g1971_n;
  wire g1972_p;
  wire g1972_n;
  wire g1973_p;
  wire g1973_n;
  wire g1974_p;
  wire g1974_n;
  wire g1975_p;
  wire g1975_n;
  wire g1976_p;
  wire g1976_n;
  wire g1977_p;
  wire g1977_n;
  wire g1978_p;
  wire g1978_n;
  wire g1979_p;
  wire g1979_n;
  wire g1980_p;
  wire g1980_n;
  wire g1981_p;
  wire g1981_n;
  wire g1982_p;
  wire g1982_n;
  wire g1983_p;
  wire g1983_n;
  wire g1984_p;
  wire g1984_n;
  wire g1985_p;
  wire g1985_n;
  wire g1986_p;
  wire g1986_n;
  wire g1987_p;
  wire g1987_n;
  wire g1988_p;
  wire g1988_n;
  wire g1989_p;
  wire g1989_n;
  wire g1990_p;
  wire g1990_n;
  wire g1991_p;
  wire g1991_n;
  wire g1992_p;
  wire g1992_n;
  wire g1993_p;
  wire g1993_n;
  wire g1994_p;
  wire g1994_n;
  wire g1995_p;
  wire g1995_n;
  wire g1996_p;
  wire g1996_n;
  wire g1997_p;
  wire g1997_n;
  wire g1998_p;
  wire g1998_n;
  wire g1999_p;
  wire g1999_n;
  wire g2000_p;
  wire g2000_n;
  wire g2001_p;
  wire g2001_n;
  wire g2002_p;
  wire g2002_n;
  wire g2003_p;
  wire g2003_n;
  wire g2004_p;
  wire g2004_n;
  wire g2005_p;
  wire g2005_n;
  wire g2006_p;
  wire g2006_n;
  wire g2007_p;
  wire g2007_n;
  wire g2008_p;
  wire g2008_n;
  wire g2009_p;
  wire g2009_n;
  wire g2010_p;
  wire g2010_n;
  wire g2011_p;
  wire g2011_n;
  wire g2012_p;
  wire g2012_n;
  wire g2013_p;
  wire g2013_n;
  wire g2014_p;
  wire g2014_n;
  wire g2015_p;
  wire g2015_n;
  wire g2016_p;
  wire g2016_n;
  wire g2017_p;
  wire g2017_n;
  wire g2018_p;
  wire g2018_n;
  wire g2019_p;
  wire g2019_n;
  wire g2020_p;
  wire g2020_n;
  wire g2021_p;
  wire g2021_n;
  wire g2022_p;
  wire g2022_n;
  wire g2023_p;
  wire g2023_n;
  wire g2024_p;
  wire g2024_n;
  wire g2025_p;
  wire g2025_n;
  wire g2026_p;
  wire g2026_n;
  wire g2027_p;
  wire g2027_n;
  wire g2028_p;
  wire g2028_n;
  wire g2029_p;
  wire g2029_n;
  wire g2030_p;
  wire g2030_n;
  wire g2031_p;
  wire g2031_n;
  wire g2032_p;
  wire g2032_n;
  wire g2033_p;
  wire g2033_n;
  wire g2034_p;
  wire g2034_n;
  wire g2035_p;
  wire g2035_n;
  wire g2036_p;
  wire g2036_n;
  wire g2037_p;
  wire g2037_n;
  wire g2038_p;
  wire g2038_n;
  wire g2039_p;
  wire g2039_n;
  wire g2040_p;
  wire g2040_n;
  wire g2041_p;
  wire g2041_n;
  wire g2042_p;
  wire g2042_n;
  wire g2043_p;
  wire g2043_n;
  wire g2044_p;
  wire g2044_n;
  wire g2045_p;
  wire g2045_n;
  wire g2046_p;
  wire g2046_n;
  wire g2047_p;
  wire g2047_n;
  wire g2048_p;
  wire g2048_n;
  wire g2049_p;
  wire g2049_n;
  wire g2050_p;
  wire g2050_n;
  wire g2051_p;
  wire g2051_n;
  wire g2052_p;
  wire g2052_n;
  wire g2053_p;
  wire g2053_n;
  wire g2054_p;
  wire g2054_n;
  wire g2055_p;
  wire g2055_n;
  wire g2056_p;
  wire g2056_n;
  wire g2057_p;
  wire g2057_n;
  wire g2058_p;
  wire g2058_n;
  wire g2059_p;
  wire g2059_n;
  wire g2060_p;
  wire g2060_n;
  wire g2061_p;
  wire g2061_n;
  wire g2062_p;
  wire g2062_n;
  wire g2063_p;
  wire g2063_n;
  wire g2064_p;
  wire g2064_n;
  wire g2065_p;
  wire g2065_n;
  wire g2066_p;
  wire g2066_n;
  wire g2067_p;
  wire g2067_n;
  wire g2068_p;
  wire g2068_n;
  wire g2069_p;
  wire g2069_n;
  wire g2070_p;
  wire g2070_n;
  wire g2071_p;
  wire g2071_n;
  wire g2072_p;
  wire g2072_n;
  wire g2073_p;
  wire g2073_n;
  wire g2074_p;
  wire g2074_n;
  wire g2075_p;
  wire g2075_n;
  wire g2076_p;
  wire g2076_n;
  wire g2077_p;
  wire g2077_n;
  wire g2078_p;
  wire g2078_n;
  wire g2079_p;
  wire g2079_n;
  wire g2080_p;
  wire g2080_n;
  wire g2081_p;
  wire g2081_n;
  wire g2082_p;
  wire g2082_n;
  wire g2083_p;
  wire g2083_n;
  wire g2084_p;
  wire g2084_n;
  wire g2085_p;
  wire g2085_n;
  wire g2086_p;
  wire g2086_n;
  wire g2087_p;
  wire g2087_n;
  wire g2088_p;
  wire g2088_n;
  wire g2089_p;
  wire g2089_n;
  wire g2090_p;
  wire g2090_n;
  wire g2091_p;
  wire g2091_n;
  wire g2092_p;
  wire g2092_n;
  wire g2093_p;
  wire g2093_n;
  wire g2094_p;
  wire g2094_n;
  wire g2095_p;
  wire g2095_n;
  wire g2096_p;
  wire g2096_n;
  wire g2097_p;
  wire g2097_n;
  wire g2098_p;
  wire g2098_n;
  wire g2099_p;
  wire g2099_n;
  wire g2100_p;
  wire g2100_n;
  wire g2101_p;
  wire g2101_n;
  wire g2102_p;
  wire g2102_n;
  wire g2103_p;
  wire g2103_n;
  wire g2104_p;
  wire g2104_n;
  wire g2105_p;
  wire g2105_n;
  wire g2106_p;
  wire g2106_n;
  wire g2107_p;
  wire g2107_n;
  wire g2108_p;
  wire g2108_n;
  wire g2109_p;
  wire g2109_n;
  wire g2110_p;
  wire g2110_n;
  wire g2111_p;
  wire g2111_n;
  wire g2112_p;
  wire g2112_n;
  wire g2113_p;
  wire g2113_n;
  wire g2114_p;
  wire g2114_n;
  wire g2115_p;
  wire g2115_n;
  wire g2116_p;
  wire g2116_n;
  wire g2117_p;
  wire g2117_n;
  wire g2118_p;
  wire g2118_n;
  wire g2119_p;
  wire g2119_n;
  wire g2120_p;
  wire g2120_n;
  wire g2121_p;
  wire g2121_n;
  wire g2122_p;
  wire g2122_n;
  wire g2123_p;
  wire g2123_n;
  wire g2124_p;
  wire g2124_n;
  wire g2125_p;
  wire g2125_n;
  wire g2126_p;
  wire g2126_n;
  wire g2127_p;
  wire g2127_n;
  wire g2128_p;
  wire g2128_n;
  wire g2129_p;
  wire g2129_n;
  wire g2130_p;
  wire g2130_n;
  wire g2131_p;
  wire g2131_n;
  wire g2132_p;
  wire g2132_n;
  wire g2133_p;
  wire g2133_n;
  wire g2134_p;
  wire g2134_n;
  wire g2135_p;
  wire g2135_n;
  wire g2136_p;
  wire g2136_n;
  wire g2137_p;
  wire g2137_n;
  wire g2138_p;
  wire g2138_n;
  wire g2139_p;
  wire g2139_n;
  wire g2140_p;
  wire g2140_n;
  wire g2141_p;
  wire g2141_n;
  wire g2142_p;
  wire g2142_n;
  wire g2143_p;
  wire g2143_n;
  wire g2144_p;
  wire g2144_n;
  wire g2145_p;
  wire g2145_n;
  wire g2146_p;
  wire g2146_n;
  wire g2147_p;
  wire g2147_n;
  wire g2148_p;
  wire g2148_n;
  wire g2149_p;
  wire g2149_n;
  wire g2150_p;
  wire g2150_n;
  wire g2151_p;
  wire g2151_n;
  wire g2152_p;
  wire g2152_n;
  wire g2153_p;
  wire g2153_n;
  wire g2154_p;
  wire g2154_n;
  wire g2155_p;
  wire g2155_n;
  wire g2156_p;
  wire g2156_n;
  wire g2157_p;
  wire g2157_n;
  wire g2158_p;
  wire g2158_n;
  wire g2159_p;
  wire g2159_n;
  wire g2160_p;
  wire g2160_n;
  wire g2161_p;
  wire g2161_n;
  wire g2162_p;
  wire g2162_n;
  wire g2163_p;
  wire g2163_n;
  wire g2164_p;
  wire g2164_n;
  wire g2165_p;
  wire g2165_n;
  wire g2166_p;
  wire g2166_n;
  wire g2167_p;
  wire g2167_n;
  wire g2168_p;
  wire g2168_n;
  wire g2169_p;
  wire g2169_n;
  wire g2170_p;
  wire g2170_n;
  wire g2171_p;
  wire g2171_n;
  wire g2172_p;
  wire g2172_n;
  wire g2173_p;
  wire g2173_n;
  wire g2174_p;
  wire g2174_n;
  wire g2175_p;
  wire g2175_n;
  wire g2176_p;
  wire g2176_n;
  wire g2177_p;
  wire g2177_n;
  wire g2178_p;
  wire g2178_n;
  wire g2179_p;
  wire g2179_n;
  wire g2180_p;
  wire g2180_n;
  wire g2181_p;
  wire g2181_n;
  wire g2182_p;
  wire g2182_n;
  wire g2183_p;
  wire g2183_n;
  wire g2184_p;
  wire g2184_n;
  wire g2185_p;
  wire g2185_n;
  wire g2186_p;
  wire g2186_n;
  wire g2187_p;
  wire g2187_n;
  wire g2188_p;
  wire g2188_n;
  wire g2189_p;
  wire g2189_n;
  wire g2190_p;
  wire g2190_n;
  wire g2191_p;
  wire g2191_n;
  wire g2192_p;
  wire g2192_n;
  wire g2193_p;
  wire g2193_n;
  wire g2194_p;
  wire g2194_n;
  wire g2195_p;
  wire g2195_n;
  wire g2196_p;
  wire g2196_n;
  wire g2197_p;
  wire g2197_n;
  wire g2198_p;
  wire g2198_n;
  wire g2199_p;
  wire g2199_n;
  wire g2200_p;
  wire g2200_n;
  wire g2201_p;
  wire g2201_n;
  wire g2202_p;
  wire g2202_n;
  wire g2203_p;
  wire g2203_n;
  wire g2204_p;
  wire g2204_n;
  wire g2205_p;
  wire g2205_n;
  wire g2206_p;
  wire g2206_n;
  wire g2207_p;
  wire g2207_n;
  wire g2208_p;
  wire g2208_n;
  wire g2209_p;
  wire g2209_n;
  wire g2210_p;
  wire g2210_n;
  wire g2211_p;
  wire g2211_n;
  wire g2212_p;
  wire g2212_n;
  wire g2213_p;
  wire g2213_n;
  wire g2214_p;
  wire g2214_n;
  wire g2215_p;
  wire g2215_n;
  wire g2216_p;
  wire g2216_n;
  wire g2217_p;
  wire g2217_n;
  wire g2218_p;
  wire g2218_n;
  wire g2219_p;
  wire g2219_n;
  wire g2220_p;
  wire g2220_n;
  wire g2221_p;
  wire g2221_n;
  wire g2222_p;
  wire g2222_n;
  wire g2223_p;
  wire g2223_n;
  wire g2224_p;
  wire g2224_n;
  wire g2225_p;
  wire g2225_n;
  wire g2226_p;
  wire g2226_n;
  wire g2227_p;
  wire g2227_n;
  wire g2228_p;
  wire g2228_n;
  wire g2229_p;
  wire g2229_n;
  wire g2230_p;
  wire g2230_n;
  wire g2231_p;
  wire g2231_n;
  wire g2232_p;
  wire g2232_n;
  wire g2233_p;
  wire g2233_n;
  wire g2234_p;
  wire g2234_n;
  wire g2235_p;
  wire g2235_n;
  wire g2236_p;
  wire g2236_n;
  wire g2237_p;
  wire g2237_n;
  wire g2238_p;
  wire g2238_n;
  wire g2239_p;
  wire g2239_n;
  wire g2240_p;
  wire g2240_n;
  wire g2241_p;
  wire g2241_n;
  wire g2242_p;
  wire g2242_n;
  wire g2243_p;
  wire g2243_n;
  wire g2244_p;
  wire g2244_n;
  wire g2245_p;
  wire g2245_n;
  wire g2246_p;
  wire g2246_n;
  wire g2247_p;
  wire g2247_n;
  wire g2248_p;
  wire g2248_n;
  wire g2249_p;
  wire g2249_n;
  wire g2250_p;
  wire g2250_n;
  wire g2251_p;
  wire g2251_n;
  wire g2252_p;
  wire g2252_n;
  wire g2253_p;
  wire g2253_n;
  wire g2254_p;
  wire g2254_n;
  wire g2255_p;
  wire g2255_n;
  wire g2256_p;
  wire g2256_n;
  wire g2257_p;
  wire g2257_n;
  wire g2258_p;
  wire g2258_n;
  wire g2259_p;
  wire g2259_n;
  wire g2260_p;
  wire g2260_n;
  wire g2261_p;
  wire g2261_n;
  wire g2262_p;
  wire g2262_n;
  wire g2263_p;
  wire g2263_n;
  wire g2264_p;
  wire g2264_n;
  wire g2265_p;
  wire g2265_n;
  wire g2266_p;
  wire g2266_n;
  wire g2267_p;
  wire g2267_n;
  wire g2268_p;
  wire g2268_n;
  wire g2269_p;
  wire g2269_n;
  wire g2270_p;
  wire g2270_n;
  wire g2271_p;
  wire g2271_n;
  wire g2272_p;
  wire g2272_n;
  wire g2273_p;
  wire g2273_n;
  wire g2274_p;
  wire g2274_n;
  wire g2275_p;
  wire g2275_n;
  wire g2276_p;
  wire g2276_n;
  wire g2277_p;
  wire g2277_n;
  wire g2278_p;
  wire g2278_n;
  wire g2279_p;
  wire g2279_n;
  wire g2280_p;
  wire g2280_n;
  wire g2281_p;
  wire g2281_n;
  wire g2282_p;
  wire g2282_n;
  wire g2283_p;
  wire g2283_n;
  wire g2284_p;
  wire g2284_n;
  wire g2285_p;
  wire g2285_n;
  wire g2286_p;
  wire g2286_n;
  wire g2287_p;
  wire g2287_n;
  wire g2288_p;
  wire g2288_n;
  wire g2289_p;
  wire g2289_n;
  wire g2290_p;
  wire g2290_n;
  wire g2291_p;
  wire g2291_n;
  wire g2292_p;
  wire g2292_n;
  wire g2293_p;
  wire g2293_n;
  wire g2294_p;
  wire g2294_n;
  wire g2295_p;
  wire g2295_n;
  wire g2296_p;
  wire g2296_n;
  wire g2297_p;
  wire g2297_n;
  wire g2298_p;
  wire g2298_n;
  wire g2299_p;
  wire g2299_n;
  wire g2300_p;
  wire g2300_n;
  wire g2301_p;
  wire g2301_n;
  wire g2302_p;
  wire g2302_n;
  wire g2303_p;
  wire g2303_n;
  wire g2304_p;
  wire g2304_n;
  wire g2305_p;
  wire g2305_n;
  wire g2306_p;
  wire g2306_n;
  wire g2307_p;
  wire g2307_n;
  wire g2308_p;
  wire g2308_n;
  wire g2309_p;
  wire g2309_n;
  wire g2310_p;
  wire g2310_n;
  wire g2311_p;
  wire g2311_n;
  wire g2312_p;
  wire g2312_n;
  wire g2313_p;
  wire g2313_n;
  wire g2314_p;
  wire g2314_n;
  wire g2315_p;
  wire g2315_n;
  wire g2316_p;
  wire g2316_n;
  wire g2317_p;
  wire g2317_n;
  wire g2318_p;
  wire g2318_n;
  wire g2319_p;
  wire g2319_n;
  wire g2320_p;
  wire g2320_n;
  wire g2321_p;
  wire g2321_n;
  wire g2322_p;
  wire g2322_n;
  wire g2323_p;
  wire g2323_n;
  wire g2324_p;
  wire g2324_n;
  wire g2325_p;
  wire g2325_n;
  wire g2326_p;
  wire g2326_n;
  wire g2327_p;
  wire g2327_n;
  wire g2328_p;
  wire g2328_n;
  wire g2329_p;
  wire g2329_n;
  wire g2330_p;
  wire g2330_n;
  wire g2331_p;
  wire g2331_n;
  wire g2332_p;
  wire g2332_n;
  wire g2333_p;
  wire g2333_n;
  wire g2334_p;
  wire g2334_n;
  wire g2335_p;
  wire g2335_n;
  wire g2336_p;
  wire g2336_n;
  wire g2337_p;
  wire g2337_n;
  wire g2338_p;
  wire g2338_n;
  wire g2339_p;
  wire g2339_n;
  wire g2340_p;
  wire g2340_n;
  wire g2341_p;
  wire g2341_n;
  wire g2342_p;
  wire g2342_n;
  wire g2343_p;
  wire g2343_n;
  wire g2344_p;
  wire g2344_n;
  wire g2345_p;
  wire g2345_n;
  wire g2346_p;
  wire g2346_n;
  wire g2347_p;
  wire g2347_n;
  wire g2348_p;
  wire g2348_n;
  wire g2349_p;
  wire g2349_n;
  wire g2350_p;
  wire g2350_n;
  wire g2351_p;
  wire g2351_n;
  wire g2352_p;
  wire g2352_n;
  wire g2353_p;
  wire g2353_n;
  wire g2354_p;
  wire g2354_n;
  wire g2355_p;
  wire g2355_n;
  wire g2356_p;
  wire g2356_n;
  wire g2357_p;
  wire g2357_n;
  wire g2358_p;
  wire g2358_n;
  wire g2359_p;
  wire g2359_n;
  wire g2360_p;
  wire g2360_n;
  wire g2361_p;
  wire g2361_n;
  wire g2362_p;
  wire g2362_n;
  wire g2363_p;
  wire g2363_n;
  wire g2364_p;
  wire g2364_n;
  wire g2365_p;
  wire g2365_n;
  wire g2366_p;
  wire g2366_n;
  wire g2367_p;
  wire g2367_n;
  wire g2368_p;
  wire g2368_n;
  wire g2369_p;
  wire g2369_n;
  wire g2370_p;
  wire g2370_n;
  wire g2371_p;
  wire g2371_n;
  wire g2372_p;
  wire g2372_n;
  wire g2373_p;
  wire g2373_n;
  wire g2374_p;
  wire g2374_n;
  wire g2375_p;
  wire g2375_n;
  wire g2376_p;
  wire g2376_n;
  wire g2377_p;
  wire g2377_n;
  wire g2378_p;
  wire g2378_n;
  wire g2379_p;
  wire g2379_n;
  wire g2380_p;
  wire g2380_n;
  wire g2381_p;
  wire g2381_n;
  wire g2382_p;
  wire g2382_n;
  wire g2383_p;
  wire g2383_n;
  wire g2384_p;
  wire g2384_n;
  wire g2385_p;
  wire g2385_n;
  wire g2386_p;
  wire g2386_n;
  wire g2387_p;
  wire g2387_n;
  wire g2388_p;
  wire g2388_n;
  wire g2389_p;
  wire g2389_n;
  wire g2390_p;
  wire g2390_n;
  wire g2391_p;
  wire g2391_n;
  wire g2392_p;
  wire g2392_n;
  wire g2393_p;
  wire g2393_n;
  wire g2394_p;
  wire g2394_n;
  wire ffc_409_n_spl_;
  wire ffc_421_n_spl_;
  wire ffc_249_p_spl_;
  wire ffc_249_p_spl_0;
  wire ffc_249_p_spl_00;
  wire ffc_249_p_spl_01;
  wire ffc_249_p_spl_1;
  wire ffc_3_p_spl_;
  wire ffc_454_n_spl_;
  wire ffc_42_n_spl_;
  wire g1055_n_spl_;
  wire g1055_n_spl_0;
  wire g1055_n_spl_00;
  wire g1055_n_spl_000;
  wire g1055_n_spl_01;
  wire g1055_n_spl_1;
  wire g1055_n_spl_10;
  wire g1055_n_spl_11;
  wire ffc_446_n_spl_;
  wire ffc_446_n_spl_0;
  wire ffc_446_n_spl_00;
  wire ffc_446_n_spl_01;
  wire ffc_446_n_spl_1;
  wire ffc_446_p_spl_;
  wire ffc_446_p_spl_0;
  wire ffc_446_p_spl_00;
  wire ffc_446_p_spl_01;
  wire ffc_446_p_spl_1;
  wire ffc_737_p_spl_;
  wire g1094_n_spl_;
  wire ffc_519_n_spl_;
  wire g1101_n_spl_;
  wire ffc_728_p_spl_;
  wire ffc_729_p_spl_;
  wire ffc_728_n_spl_;
  wire ffc_729_n_spl_;
  wire ffc_730_n_spl_;
  wire ffc_753_n_spl_;
  wire ffc_730_p_spl_;
  wire ffc_753_p_spl_;
  wire ffc_532_p_spl_;
  wire ffc_532_p_spl_0;
  wire ffc_697_p_spl_;
  wire ffc_697_p_spl_0;
  wire ffc_697_p_spl_00;
  wire ffc_697_p_spl_000;
  wire ffc_697_p_spl_001;
  wire ffc_697_p_spl_01;
  wire ffc_697_p_spl_010;
  wire ffc_697_p_spl_011;
  wire ffc_697_p_spl_1;
  wire ffc_697_p_spl_10;
  wire ffc_697_p_spl_100;
  wire ffc_697_p_spl_101;
  wire ffc_697_p_spl_11;
  wire ffc_697_p_spl_110;
  wire ffc_697_p_spl_111;
  wire ffc_498_n_spl_;
  wire ffc_498_n_spl_0;
  wire ffc_498_n_spl_00;
  wire ffc_498_n_spl_000;
  wire ffc_498_n_spl_01;
  wire ffc_498_n_spl_1;
  wire ffc_498_n_spl_10;
  wire ffc_498_n_spl_11;
  wire ffc_494_p_spl_;
  wire ffc_494_p_spl_0;
  wire ffc_494_p_spl_00;
  wire ffc_494_p_spl_000;
  wire ffc_494_p_spl_001;
  wire ffc_494_p_spl_01;
  wire ffc_494_p_spl_010;
  wire ffc_494_p_spl_011;
  wire ffc_494_p_spl_1;
  wire ffc_494_p_spl_10;
  wire ffc_494_p_spl_100;
  wire ffc_494_p_spl_101;
  wire ffc_494_p_spl_11;
  wire ffc_494_p_spl_110;
  wire ffc_697_n_spl_;
  wire ffc_498_p_spl_;
  wire ffc_498_p_spl_0;
  wire ffc_498_p_spl_00;
  wire ffc_498_p_spl_000;
  wire ffc_498_p_spl_01;
  wire ffc_498_p_spl_1;
  wire ffc_498_p_spl_10;
  wire ffc_498_p_spl_11;
  wire ffc_494_n_spl_;
  wire ffc_494_n_spl_0;
  wire ffc_494_n_spl_1;
  wire ffc_723_p_spl_;
  wire ffc_482_n_spl_;
  wire ffc_482_n_spl_0;
  wire ffc_482_n_spl_00;
  wire ffc_482_n_spl_000;
  wire ffc_482_n_spl_0000;
  wire ffc_482_n_spl_0001;
  wire ffc_482_n_spl_001;
  wire ffc_482_n_spl_0010;
  wire ffc_482_n_spl_0011;
  wire ffc_482_n_spl_01;
  wire ffc_482_n_spl_010;
  wire ffc_482_n_spl_011;
  wire ffc_482_n_spl_1;
  wire ffc_482_n_spl_10;
  wire ffc_482_n_spl_100;
  wire ffc_482_n_spl_101;
  wire ffc_482_n_spl_11;
  wire ffc_482_n_spl_110;
  wire ffc_482_n_spl_111;
  wire g1132_n_spl_;
  wire g1132_n_spl_0;
  wire g1132_n_spl_00;
  wire g1132_n_spl_1;
  wire ffc_482_p_spl_;
  wire ffc_482_p_spl_0;
  wire ffc_482_p_spl_00;
  wire ffc_482_p_spl_000;
  wire ffc_482_p_spl_0000;
  wire ffc_482_p_spl_0001;
  wire ffc_482_p_spl_001;
  wire ffc_482_p_spl_0010;
  wire ffc_482_p_spl_0011;
  wire ffc_482_p_spl_01;
  wire ffc_482_p_spl_010;
  wire ffc_482_p_spl_011;
  wire ffc_482_p_spl_1;
  wire ffc_482_p_spl_10;
  wire ffc_482_p_spl_100;
  wire ffc_482_p_spl_101;
  wire ffc_482_p_spl_11;
  wire ffc_482_p_spl_110;
  wire ffc_482_p_spl_111;
  wire g1142_n_spl_;
  wire g1142_n_spl_0;
  wire g1142_n_spl_00;
  wire g1142_n_spl_1;
  wire ffc_478_p_spl_;
  wire ffc_478_p_spl_0;
  wire ffc_478_p_spl_00;
  wire ffc_478_p_spl_000;
  wire ffc_478_p_spl_001;
  wire ffc_478_p_spl_01;
  wire ffc_478_p_spl_1;
  wire ffc_478_p_spl_10;
  wire ffc_478_p_spl_11;
  wire ffc_10_p_spl_;
  wire ffc_84_p_spl_;
  wire ffc_478_n_spl_;
  wire ffc_478_n_spl_0;
  wire ffc_478_n_spl_00;
  wire ffc_478_n_spl_000;
  wire ffc_478_n_spl_001;
  wire ffc_478_n_spl_01;
  wire ffc_478_n_spl_1;
  wire ffc_478_n_spl_10;
  wire ffc_478_n_spl_11;
  wire ffc_523_n_spl_;
  wire ffc_744_n_spl_;
  wire g1159_n_spl_;
  wire ffc_486_n_spl_;
  wire ffc_486_n_spl_0;
  wire ffc_486_n_spl_00;
  wire ffc_486_n_spl_000;
  wire ffc_486_n_spl_0000;
  wire ffc_486_n_spl_0001;
  wire ffc_486_n_spl_001;
  wire ffc_486_n_spl_0010;
  wire ffc_486_n_spl_0011;
  wire ffc_486_n_spl_01;
  wire ffc_486_n_spl_010;
  wire ffc_486_n_spl_011;
  wire ffc_486_n_spl_1;
  wire ffc_486_n_spl_10;
  wire ffc_486_n_spl_100;
  wire ffc_486_n_spl_101;
  wire ffc_486_n_spl_11;
  wire ffc_486_n_spl_110;
  wire ffc_486_n_spl_111;
  wire ffc_486_p_spl_;
  wire ffc_486_p_spl_0;
  wire ffc_486_p_spl_00;
  wire ffc_486_p_spl_000;
  wire ffc_486_p_spl_0000;
  wire ffc_486_p_spl_0001;
  wire ffc_486_p_spl_001;
  wire ffc_486_p_spl_0010;
  wire ffc_486_p_spl_0011;
  wire ffc_486_p_spl_01;
  wire ffc_486_p_spl_010;
  wire ffc_486_p_spl_011;
  wire ffc_486_p_spl_1;
  wire ffc_486_p_spl_10;
  wire ffc_486_p_spl_100;
  wire ffc_486_p_spl_101;
  wire ffc_486_p_spl_11;
  wire ffc_486_p_spl_110;
  wire ffc_486_p_spl_111;
  wire ffc_490_p_spl_;
  wire ffc_490_p_spl_0;
  wire ffc_490_p_spl_00;
  wire ffc_490_p_spl_000;
  wire ffc_490_p_spl_001;
  wire ffc_490_p_spl_01;
  wire ffc_490_p_spl_1;
  wire ffc_490_p_spl_10;
  wire ffc_490_p_spl_11;
  wire ffc_490_n_spl_;
  wire ffc_490_n_spl_0;
  wire ffc_490_n_spl_00;
  wire ffc_490_n_spl_000;
  wire ffc_490_n_spl_001;
  wire ffc_490_n_spl_01;
  wire ffc_490_n_spl_1;
  wire ffc_490_n_spl_10;
  wire ffc_490_n_spl_11;
  wire g1176_n_spl_;
  wire g1183_n_spl_;
  wire g1188_n_spl_;
  wire ffc_561_n_spl_;
  wire ffc_561_n_spl_0;
  wire ffc_561_n_spl_00;
  wire ffc_561_n_spl_1;
  wire g1201_n_spl_;
  wire ffc_561_p_spl_;
  wire ffc_561_p_spl_0;
  wire ffc_561_p_spl_1;
  wire g1201_p_spl_;
  wire g1205_p_spl_;
  wire g1206_n_spl_;
  wire g1205_n_spl_;
  wire g1206_p_spl_;
  wire ffc_504_n_spl_;
  wire ffc_505_p_spl_;
  wire ffc_504_p_spl_;
  wire ffc_505_n_spl_;
  wire ffc_507_n_spl_;
  wire ffc_511_p_spl_;
  wire ffc_507_p_spl_;
  wire ffc_511_n_spl_;
  wire g1215_n_spl_;
  wire g1218_p_spl_;
  wire g1215_p_spl_;
  wire g1218_n_spl_;
  wire ffc_739_n_spl_;
  wire ffc_742_p_spl_;
  wire ffc_739_p_spl_;
  wire ffc_742_n_spl_;
  wire ffc_503_p_spl_;
  wire ffc_506_n_spl_;
  wire ffc_503_n_spl_;
  wire ffc_506_p_spl_;
  wire g1224_n_spl_;
  wire g1227_p_spl_;
  wire g1224_p_spl_;
  wire g1227_n_spl_;
  wire g1234_n_spl_;
  wire ffc_745_n_spl_;
  wire g1243_p_spl_;
  wire g1246_p_spl_;
  wire ffc_746_p_spl_;
  wire g1250_p_spl_;
  wire g1249_p_spl_;
  wire ffc_428_n_spl_;
  wire ffc_428_n_spl_0;
  wire ffc_428_n_spl_00;
  wire ffc_428_n_spl_000;
  wire ffc_428_n_spl_0000;
  wire ffc_428_n_spl_0001;
  wire ffc_428_n_spl_001;
  wire ffc_428_n_spl_0010;
  wire ffc_428_n_spl_0011;
  wire ffc_428_n_spl_01;
  wire ffc_428_n_spl_010;
  wire ffc_428_n_spl_011;
  wire ffc_428_n_spl_1;
  wire ffc_428_n_spl_10;
  wire ffc_428_n_spl_100;
  wire ffc_428_n_spl_101;
  wire ffc_428_n_spl_11;
  wire ffc_428_n_spl_110;
  wire ffc_428_n_spl_111;
  wire ffc_428_p_spl_;
  wire ffc_428_p_spl_0;
  wire ffc_428_p_spl_00;
  wire ffc_428_p_spl_000;
  wire ffc_428_p_spl_0000;
  wire ffc_428_p_spl_0001;
  wire ffc_428_p_spl_001;
  wire ffc_428_p_spl_0010;
  wire ffc_428_p_spl_0011;
  wire ffc_428_p_spl_01;
  wire ffc_428_p_spl_010;
  wire ffc_428_p_spl_011;
  wire ffc_428_p_spl_1;
  wire ffc_428_p_spl_10;
  wire ffc_428_p_spl_100;
  wire ffc_428_p_spl_101;
  wire ffc_428_p_spl_11;
  wire ffc_428_p_spl_110;
  wire ffc_428_p_spl_111;
  wire ffc_432_n_spl_;
  wire ffc_432_n_spl_0;
  wire ffc_432_n_spl_00;
  wire ffc_432_n_spl_000;
  wire ffc_432_n_spl_001;
  wire ffc_432_n_spl_01;
  wire ffc_432_n_spl_1;
  wire ffc_432_n_spl_10;
  wire ffc_432_n_spl_11;
  wire ffc_309_p_spl_;
  wire ffc_305_p_spl_;
  wire ffc_432_p_spl_;
  wire ffc_432_p_spl_0;
  wire ffc_432_p_spl_00;
  wire ffc_432_p_spl_000;
  wire ffc_432_p_spl_001;
  wire ffc_432_p_spl_01;
  wire ffc_432_p_spl_1;
  wire ffc_432_p_spl_10;
  wire ffc_432_p_spl_11;
  wire ffc_241_p_spl_;
  wire ffc_241_p_spl_0;
  wire ffc_241_p_spl_00;
  wire ffc_241_p_spl_000;
  wire ffc_241_p_spl_0000;
  wire ffc_241_p_spl_001;
  wire ffc_241_p_spl_01;
  wire ffc_241_p_spl_010;
  wire ffc_241_p_spl_011;
  wire ffc_241_p_spl_1;
  wire ffc_241_p_spl_10;
  wire ffc_241_p_spl_100;
  wire ffc_241_p_spl_101;
  wire ffc_241_p_spl_11;
  wire ffc_241_p_spl_110;
  wire ffc_241_p_spl_111;
  wire ffc_436_n_spl_;
  wire ffc_436_n_spl_0;
  wire ffc_436_n_spl_00;
  wire ffc_436_n_spl_000;
  wire ffc_436_n_spl_0000;
  wire ffc_436_n_spl_0001;
  wire ffc_436_n_spl_001;
  wire ffc_436_n_spl_0010;
  wire ffc_436_n_spl_0011;
  wire ffc_436_n_spl_01;
  wire ffc_436_n_spl_010;
  wire ffc_436_n_spl_011;
  wire ffc_436_n_spl_1;
  wire ffc_436_n_spl_10;
  wire ffc_436_n_spl_100;
  wire ffc_436_n_spl_101;
  wire ffc_436_n_spl_11;
  wire ffc_436_n_spl_110;
  wire ffc_436_n_spl_111;
  wire ffc_436_p_spl_;
  wire ffc_436_p_spl_0;
  wire ffc_436_p_spl_00;
  wire ffc_436_p_spl_000;
  wire ffc_436_p_spl_0000;
  wire ffc_436_p_spl_0001;
  wire ffc_436_p_spl_001;
  wire ffc_436_p_spl_0010;
  wire ffc_436_p_spl_0011;
  wire ffc_436_p_spl_01;
  wire ffc_436_p_spl_010;
  wire ffc_436_p_spl_011;
  wire ffc_436_p_spl_1;
  wire ffc_436_p_spl_10;
  wire ffc_436_p_spl_100;
  wire ffc_436_p_spl_101;
  wire ffc_436_p_spl_11;
  wire ffc_436_p_spl_110;
  wire ffc_436_p_spl_111;
  wire ffc_440_n_spl_;
  wire ffc_440_n_spl_0;
  wire ffc_440_n_spl_00;
  wire ffc_440_n_spl_000;
  wire ffc_440_n_spl_001;
  wire ffc_440_n_spl_01;
  wire ffc_440_n_spl_1;
  wire ffc_440_n_spl_10;
  wire ffc_440_n_spl_11;
  wire ffc_440_p_spl_;
  wire ffc_440_p_spl_0;
  wire ffc_440_p_spl_00;
  wire ffc_440_p_spl_000;
  wire ffc_440_p_spl_001;
  wire ffc_440_p_spl_01;
  wire ffc_440_p_spl_1;
  wire ffc_440_p_spl_10;
  wire ffc_440_p_spl_11;
  wire ffc_54_p_spl_;
  wire ffc_62_p_spl_;
  wire g1182_n_spl_;
  wire g1182_n_spl_0;
  wire g1182_n_spl_00;
  wire g1182_n_spl_1;
  wire g1155_n_spl_;
  wire g1155_n_spl_0;
  wire g1155_n_spl_00;
  wire g1155_n_spl_1;
  wire ffc_22_p_spl_;
  wire ffc_104_p_spl_;
  wire g1187_n_spl_;
  wire g1187_n_spl_0;
  wire g1187_n_spl_00;
  wire g1187_n_spl_1;
  wire g1158_n_spl_;
  wire g1158_n_spl_0;
  wire g1158_n_spl_00;
  wire g1158_n_spl_1;
  wire ffc_18_p_spl_;
  wire ffc_100_p_spl_;
  wire g1194_n_spl_;
  wire g1194_n_spl_0;
  wire g1194_n_spl_00;
  wire g1194_n_spl_1;
  wire g1164_n_spl_;
  wire g1164_n_spl_0;
  wire g1164_n_spl_00;
  wire g1164_n_spl_1;
  wire ffc_96_n_spl_;
  wire ffc_92_n_spl_;
  wire g1200_p_spl_;
  wire g1200_p_spl_0;
  wire g1200_p_spl_00;
  wire g1200_p_spl_1;
  wire g1137_p_spl_;
  wire g1137_p_spl_0;
  wire g1137_p_spl_00;
  wire g1137_p_spl_1;
  wire ffc_289_p_spl_;
  wire ffc_329_p_spl_;
  wire ffc_273_n_spl_;
  wire ffc_313_n_spl_;
  wire ffc_241_n_spl_;
  wire ffc_241_n_spl_0;
  wire ffc_241_n_spl_1;
  wire ffc_265_p_spl_;
  wire ffc_269_p_spl_;
  wire ffc_257_p_spl_;
  wire ffc_261_p_spl_;
  wire ffc_474_n_spl_;
  wire ffc_474_p_spl_;
  wire ffc_229_n_spl_;
  wire ffc_229_p_spl_;
  wire ffc_532_n_spl_;
  wire g1437_n_spl_;
  wire ffc_342_n_spl_;
  wire ffc_417_n_spl_;
  wire g1049_n_spl_;
  wire g1054_n_spl_;
  wire g1111_n_spl_;
  wire g1120_n_spl_;
  wire g1212_n_spl_;
  wire g1233_n_spl_;
  wire ffc_160_p_spl_;
  wire ffc_164_p_spl_;
  wire g1470_n_spl_;
  wire g1470_n_spl_0;
  wire g1470_n_spl_00;
  wire g1470_n_spl_1;
  wire g1449_n_spl_;
  wire g1449_n_spl_0;
  wire g1449_n_spl_00;
  wire g1449_n_spl_1;
  wire ffc_70_p_spl_;
  wire ffc_66_p_spl_;
  wire g1476_n_spl_;
  wire g1476_n_spl_0;
  wire g1476_n_spl_00;
  wire g1476_n_spl_1;
  wire g1453_n_spl_;
  wire g1453_n_spl_0;
  wire g1453_n_spl_00;
  wire g1453_n_spl_1;
  wire ffc_156_p_spl_;
  wire ffc_152_p_spl_;
  wire g1482_n_spl_;
  wire g1482_n_spl_0;
  wire g1482_n_spl_00;
  wire g1482_n_spl_1;
  wire g1457_n_spl_;
  wire g1457_n_spl_0;
  wire g1457_n_spl_00;
  wire g1457_n_spl_1;
  wire ffc_58_p_spl_;
  wire ffc_140_p_spl_;
  wire g1486_n_spl_;
  wire g1486_n_spl_0;
  wire g1486_n_spl_00;
  wire g1486_n_spl_1;
  wire g1460_n_spl_;
  wire g1460_n_spl_0;
  wire g1460_n_spl_00;
  wire g1460_n_spl_1;
  wire ffc_293_p_spl_;
  wire ffc_333_p_spl_;
  wire ffc_285_p_spl_;
  wire ffc_325_p_spl_;
  wire ffc_281_p_spl_;
  wire ffc_321_p_spl_;
  wire ffc_277_p_spl_;
  wire ffc_317_p_spl_;
  wire g1640_n_spl_;
  wire g1639_n_spl_;
  wire g1645_n_spl_;
  wire ffc_88_n_spl_;
  wire ffc_14_n_spl_;
  wire g1653_p_spl_;
  wire g1653_p_spl_0;
  wire g1653_p_spl_1;
  wire g1656_p_spl_;
  wire g1656_p_spl_0;
  wire g1656_p_spl_1;
  wire ffc_301_n_spl_;
  wire ffc_297_n_spl_;
  wire ffc_610_n_spl_;
  wire ffc_610_n_spl_0;
  wire ffc_610_n_spl_1;
  wire ffc_783_n_spl_;
  wire ffc_610_p_spl_;
  wire ffc_610_p_spl_0;
  wire ffc_783_p_spl_;
  wire ffc_783_p_spl_0;
  wire g1690_n_spl_;
  wire ffc_578_n_spl_;
  wire ffc_578_n_spl_0;
  wire ffc_578_n_spl_00;
  wire ffc_578_n_spl_1;
  wire ffc_624_n_spl_;
  wire ffc_6_p_spl_;
  wire ffc_6_p_spl_0;
  wire ffc_6_p_spl_1;
  wire ffc_587_p_spl_;
  wire g1695_n_spl_;
  wire ffc_842_n_spl_;
  wire ffc_842_p_spl_;
  wire ffc_842_p_spl_0;
  wire ffc_827_n_spl_;
  wire ffc_827_p_spl_;
  wire ffc_840_p_spl_;
  wire ffc_843_p_spl_;
  wire ffc_843_p_spl_0;
  wire ffc_845_p_spl_;
  wire ffc_843_n_spl_;
  wire ffc_770_p_spl_;
  wire ffc_770_p_spl_0;
  wire g1703_p_spl_;
  wire g1703_p_spl_0;
  wire ffc_770_n_spl_;
  wire g1703_n_spl_;
  wire ffc_466_n_spl_;
  wire ffc_466_n_spl_0;
  wire ffc_466_n_spl_00;
  wire ffc_466_n_spl_000;
  wire ffc_466_n_spl_001;
  wire ffc_466_n_spl_01;
  wire ffc_466_n_spl_010;
  wire ffc_466_n_spl_011;
  wire ffc_466_n_spl_1;
  wire ffc_466_n_spl_10;
  wire ffc_466_n_spl_11;
  wire ffc_457_p_spl_;
  wire ffc_457_p_spl_0;
  wire ffc_457_p_spl_00;
  wire ffc_457_p_spl_000;
  wire ffc_457_p_spl_001;
  wire ffc_457_p_spl_01;
  wire ffc_457_p_spl_010;
  wire ffc_457_p_spl_011;
  wire ffc_457_p_spl_1;
  wire ffc_457_p_spl_10;
  wire ffc_457_p_spl_11;
  wire ffc_623_p_spl_;
  wire ffc_623_p_spl_0;
  wire ffc_829_p_spl_;
  wire ffc_829_p_spl_0;
  wire ffc_829_p_spl_00;
  wire ffc_829_p_spl_01;
  wire ffc_829_p_spl_1;
  wire ffc_623_n_spl_;
  wire ffc_829_n_spl_;
  wire ffc_829_n_spl_0;
  wire ffc_829_n_spl_00;
  wire ffc_829_n_spl_1;
  wire ffc_775_p_spl_;
  wire ffc_683_p_spl_;
  wire g1698_n_spl_;
  wire g1698_n_spl_0;
  wire g1698_n_spl_1;
  wire g1698_p_spl_;
  wire g1698_p_spl_0;
  wire ffc_813_n_spl_;
  wire ffc_813_p_spl_;
  wire ffc_795_p_spl_;
  wire ffc_795_p_spl_0;
  wire ffc_795_p_spl_1;
  wire ffc_815_n_spl_;
  wire ffc_795_n_spl_;
  wire ffc_795_n_spl_0;
  wire ffc_815_p_spl_;
  wire ffc_816_p_spl_;
  wire ffc_816_p_spl_0;
  wire ffc_816_p_spl_00;
  wire ffc_816_p_spl_1;
  wire g1700_n_spl_;
  wire g1700_n_spl_0;
  wire ffc_816_n_spl_;
  wire ffc_816_n_spl_0;
  wire ffc_816_n_spl_1;
  wire g1700_p_spl_;
  wire g1717_n_spl_;
  wire g1717_p_spl_;
  wire g1696_p_spl_;
  wire ffc_603_p_spl_;
  wire g1723_n_spl_;
  wire ffc_769_p_spl_;
  wire ffc_769_p_spl_0;
  wire ffc_769_p_spl_1;
  wire ffc_844_p_spl_;
  wire ffc_844_p_spl_0;
  wire ffc_844_p_spl_1;
  wire ffc_769_n_spl_;
  wire ffc_844_n_spl_;
  wire ffc_596_p_spl_;
  wire ffc_596_p_spl_0;
  wire ffc_556_n_spl_;
  wire ffc_556_n_spl_0;
  wire ffc_556_n_spl_1;
  wire ffc_463_n_spl_;
  wire ffc_463_n_spl_0;
  wire ffc_463_n_spl_00;
  wire ffc_463_n_spl_000;
  wire ffc_463_n_spl_001;
  wire ffc_463_n_spl_01;
  wire ffc_463_n_spl_010;
  wire ffc_463_n_spl_1;
  wire ffc_463_n_spl_10;
  wire ffc_463_n_spl_11;
  wire ffc_556_p_spl_;
  wire ffc_556_p_spl_0;
  wire ffc_556_p_spl_1;
  wire ffc_460_p_spl_;
  wire ffc_460_p_spl_0;
  wire ffc_460_p_spl_00;
  wire ffc_460_p_spl_000;
  wire ffc_460_p_spl_001;
  wire ffc_460_p_spl_01;
  wire ffc_460_p_spl_010;
  wire ffc_460_p_spl_1;
  wire ffc_460_p_spl_10;
  wire ffc_460_p_spl_11;
  wire ffc_527_n_spl_;
  wire ffc_527_n_spl_0;
  wire ffc_527_p_spl_;
  wire ffc_527_p_spl_0;
  wire ffc_590_n_spl_;
  wire ffc_590_n_spl_0;
  wire ffc_590_p_spl_;
  wire ffc_590_p_spl_0;
  wire ffc_390_p_spl_;
  wire ffc_390_p_spl_0;
  wire ffc_390_p_spl_00;
  wire ffc_390_p_spl_1;
  wire g1711_n_spl_;
  wire g1711_n_spl_0;
  wire ffc_390_n_spl_;
  wire ffc_390_n_spl_0;
  wire ffc_390_n_spl_1;
  wire g1711_p_spl_;
  wire g1756_p_spl_;
  wire ffc_839_p_spl_;
  wire ffc_839_p_spl_0;
  wire ffc_839_p_spl_00;
  wire ffc_839_p_spl_000;
  wire ffc_839_p_spl_001;
  wire ffc_839_p_spl_01;
  wire ffc_839_p_spl_1;
  wire ffc_839_p_spl_10;
  wire ffc_839_p_spl_11;
  wire ffc_859_p_spl_;
  wire ffc_839_n_spl_;
  wire ffc_839_n_spl_0;
  wire ffc_839_n_spl_00;
  wire ffc_839_n_spl_000;
  wire ffc_839_n_spl_01;
  wire ffc_839_n_spl_1;
  wire ffc_839_n_spl_10;
  wire ffc_839_n_spl_11;
  wire ffc_857_p_spl_;
  wire ffc_857_p_spl_0;
  wire g1721_n_spl_;
  wire g1721_n_spl_0;
  wire ffc_858_p_spl_;
  wire ffc_858_p_spl_0;
  wire g1720_n_spl_;
  wire g1720_n_spl_0;
  wire ffc_861_p_spl_;
  wire ffc_863_p_spl_;
  wire ffc_863_p_spl_0;
  wire ffc_863_p_spl_00;
  wire ffc_863_p_spl_000;
  wire ffc_863_p_spl_001;
  wire ffc_863_p_spl_01;
  wire ffc_863_p_spl_010;
  wire ffc_863_p_spl_011;
  wire ffc_863_p_spl_1;
  wire ffc_863_p_spl_10;
  wire ffc_863_p_spl_11;
  wire ffc_863_n_spl_;
  wire ffc_863_n_spl_0;
  wire ffc_863_n_spl_00;
  wire ffc_863_n_spl_000;
  wire ffc_863_n_spl_001;
  wire ffc_863_n_spl_01;
  wire ffc_863_n_spl_010;
  wire ffc_863_n_spl_1;
  wire ffc_863_n_spl_10;
  wire ffc_863_n_spl_11;
  wire g1704_p_spl_;
  wire g1719_p_spl_;
  wire g1719_p_spl_0;
  wire g1772_n_spl_;
  wire g1719_n_spl_;
  wire g1772_p_spl_;
  wire g1773_n_spl_;
  wire g1773_p_spl_;
  wire ffc_850_p_spl_;
  wire ffc_852_p_spl_;
  wire g1699_p_spl_;
  wire g1699_p_spl_0;
  wire g1781_p_spl_;
  wire g1699_n_spl_;
  wire g1699_n_spl_0;
  wire g1699_n_spl_1;
  wire g1781_n_spl_;
  wire g1712_p_spl_;
  wire g1712_p_spl_0;
  wire g1785_p_spl_;
  wire ffc_854_p_spl_;
  wire ffc_848_p_spl_;
  wire ffc_848_p_spl_0;
  wire g1761_n_spl_;
  wire g1761_n_spl_0;
  wire ffc_856_p_spl_;
  wire ffc_856_p_spl_0;
  wire g1722_n_spl_;
  wire g1722_n_spl_0;
  wire g1763_n_spl_;
  wire g1763_n_spl_0;
  wire g1763_n_spl_1;
  wire ffc_846_p_spl_;
  wire ffc_847_p_spl_;
  wire ffc_388_p_spl_;
  wire ffc_388_p_spl_0;
  wire g1780_n_spl_;
  wire g1780_n_spl_0;
  wire ffc_392_p_spl_;
  wire ffc_392_p_spl_0;
  wire g1777_n_spl_;
  wire g1777_n_spl_0;
  wire ffc_393_p_spl_;
  wire ffc_393_p_spl_0;
  wire g1790_n_spl_;
  wire g1790_n_spl_0;
  wire ffc_849_p_spl_;
  wire ffc_849_p_spl_0;
  wire g1767_n_spl_;
  wire g1767_n_spl_0;
  wire g1807_n_spl_;
  wire g1797_p_spl_;
  wire g1799_p_spl_;
  wire g1799_p_spl_0;
  wire ffc_497_n_spl_;
  wire ffc_497_n_spl_0;
  wire ffc_497_n_spl_00;
  wire ffc_497_n_spl_000;
  wire ffc_497_n_spl_001;
  wire ffc_497_n_spl_01;
  wire ffc_497_n_spl_010;
  wire ffc_497_n_spl_1;
  wire ffc_497_n_spl_10;
  wire ffc_497_n_spl_11;
  wire ffc_497_p_spl_;
  wire ffc_497_p_spl_0;
  wire ffc_497_p_spl_00;
  wire ffc_497_p_spl_000;
  wire ffc_497_p_spl_001;
  wire ffc_497_p_spl_01;
  wire ffc_497_p_spl_010;
  wire ffc_497_p_spl_011;
  wire ffc_497_p_spl_1;
  wire ffc_497_p_spl_10;
  wire ffc_497_p_spl_100;
  wire ffc_497_p_spl_101;
  wire ffc_497_p_spl_11;
  wire ffc_528_n_spl_;
  wire ffc_528_n_spl_0;
  wire ffc_528_p_spl_;
  wire ffc_528_p_spl_0;
  wire ffc_493_n_spl_;
  wire ffc_493_n_spl_0;
  wire ffc_204_p_spl_;
  wire ffc_493_p_spl_;
  wire ffc_493_p_spl_0;
  wire ffc_604_n_spl_;
  wire ffc_604_p_spl_;
  wire ffc_605_p_spl_;
  wire ffc_605_p_spl_0;
  wire ffc_615_p_spl_;
  wire ffc_791_p_spl_;
  wire ffc_811_p_spl_;
  wire ffc_791_n_spl_;
  wire ffc_811_n_spl_;
  wire g1831_p_spl_;
  wire g1834_n_spl_;
  wire g1831_n_spl_;
  wire g1834_p_spl_;
  wire ffc_578_p_spl_;
  wire g1692_p_spl_;
  wire g1692_p_spl_0;
  wire g1840_n_spl_;
  wire g1692_n_spl_;
  wire g1692_n_spl_0;
  wire g1840_p_spl_;
  wire g1755_n_spl_;
  wire g1737_n_spl_;
  wire g1746_n_spl_;
  wire g1854_p_spl_;
  wire g1855_n_spl_;
  wire g1854_n_spl_;
  wire g1855_p_spl_;
  wire ffc_802_p_spl_;
  wire ffc_800_p_spl_;
  wire g1859_p_spl_;
  wire g1860_p_spl_;
  wire g1859_n_spl_;
  wire g1860_n_spl_;
  wire ffc_772_p_spl_;
  wire ffc_772_p_spl_0;
  wire ffc_772_p_spl_1;
  wire ffc_6_n_spl_;
  wire ffc_772_n_spl_;
  wire ffc_772_n_spl_0;
  wire ffc_771_n_spl_;
  wire ffc_771_n_spl_0;
  wire ffc_771_n_spl_1;
  wire ffc_771_p_spl_;
  wire ffc_771_p_spl_0;
  wire ffc_771_p_spl_00;
  wire ffc_771_p_spl_1;
  wire g1872_n_spl_;
  wire g1872_n_spl_0;
  wire g1872_n_spl_00;
  wire g1872_n_spl_1;
  wire g1872_p_spl_;
  wire g1872_p_spl_0;
  wire g1872_p_spl_00;
  wire g1872_p_spl_1;
  wire ffc_659_p_spl_;
  wire ffc_659_n_spl_;
  wire ffc_659_n_spl_0;
  wire g1877_n_spl_;
  wire g1724_p_spl_;
  wire ffc_375_p_spl_;
  wire ffc_375_p_spl_0;
  wire g1884_n_spl_;
  wire ffc_609_p_spl_;
  wire g1693_n_spl_;
  wire g1891_p_spl_;
  wire g1728_n_spl_;
  wire ffc_592_p_spl_;
  wire g1895_n_spl_;
  wire ffc_364_p_spl_;
  wire ffc_790_n_spl_;
  wire ffc_790_n_spl_0;
  wire g1708_n_spl_;
  wire ffc_539_p_spl_;
  wire ffc_539_p_spl_0;
  wire ffc_539_n_spl_;
  wire ffc_539_n_spl_0;
  wire ffc_526_p_spl_;
  wire ffc_526_p_spl_0;
  wire ffc_526_n_spl_;
  wire ffc_526_n_spl_0;
  wire ffc_540_p_spl_;
  wire ffc_540_p_spl_0;
  wire ffc_540_n_spl_;
  wire ffc_540_n_spl_0;
  wire ffc_536_n_spl_;
  wire ffc_536_n_spl_0;
  wire ffc_536_n_spl_1;
  wire ffc_536_p_spl_;
  wire ffc_536_p_spl_0;
  wire ffc_536_p_spl_1;
  wire ffc_598_n_spl_;
  wire ffc_598_n_spl_0;
  wire ffc_598_n_spl_1;
  wire ffc_598_p_spl_;
  wire ffc_598_p_spl_0;
  wire ffc_598_p_spl_1;
  wire ffc_557_n_spl_;
  wire ffc_557_n_spl_0;
  wire ffc_557_p_spl_;
  wire ffc_557_p_spl_0;
  wire ffc_549_n_spl_;
  wire ffc_549_n_spl_0;
  wire ffc_549_p_spl_;
  wire ffc_549_p_spl_0;
  wire ffc_785_n_spl_;
  wire ffc_786_p_spl_;
  wire ffc_785_p_spl_;
  wire ffc_786_n_spl_;
  wire ffc_789_n_spl_;
  wire ffc_789_p_spl_;
  wire ffc_790_p_spl_;
  wire ffc_790_p_spl_0;
  wire g1982_n_spl_;
  wire g1985_p_spl_;
  wire g1982_p_spl_;
  wire g1985_n_spl_;
  wire ffc_784_n_spl_;
  wire ffc_788_p_spl_;
  wire ffc_784_p_spl_;
  wire ffc_788_n_spl_;
  wire ffc_787_n_spl_;
  wire ffc_810_n_spl_;
  wire ffc_787_p_spl_;
  wire ffc_810_p_spl_;
  wire g1991_p_spl_;
  wire g1994_n_spl_;
  wire g1991_n_spl_;
  wire g1994_p_spl_;
  wire ffc_350_p_spl_;
  wire ffc_350_p_spl_0;
  wire ffc_529_p_spl_;
  wire ffc_350_n_spl_;
  wire ffc_350_n_spl_0;
  wire ffc_529_n_spl_;
  wire ffc_608_p_spl_;
  wire ffc_614_p_spl_;
  wire ffc_640_p_spl_;
  wire g2035_n_spl_;
  wire g2038_p_spl_;
  wire ffc_375_n_spl_;
  wire ffc_571_p_spl_;
  wire ffc_571_n_spl_;
  wire g2046_n_spl_;
  wire g2049_p_spl_;
  wire g2054_n_spl_;
  wire g2057_n_spl_;
  wire g2069_p_spl_;
  wire g2070_n_spl_;
  wire g2069_n_spl_;
  wire g2070_p_spl_;
  wire ffc_424_n_spl_;
  wire ffc_424_n_spl_0;
  wire ffc_424_n_spl_1;
  wire ffc_424_p_spl_;
  wire ffc_424_p_spl_0;
  wire ffc_424_p_spl_1;
  wire g2075_p_spl_;
  wire g2076_p_spl_;
  wire g2075_n_spl_;
  wire g2076_n_spl_;
  wire g2082_n_spl_;
  wire g2082_p_spl_;
  wire g2085_p_spl_;
  wire g2085_n_spl_;
  wire g1793_p_spl_;
  wire g1796_p_spl_;
  wire g1796_p_spl_0;
  wire g1762_p_spl_;
  wire ffc_628_n_spl_;
  wire ffc_832_n_spl_;
  wire ffc_832_n_spl_0;
  wire ffc_832_n_spl_00;
  wire ffc_832_n_spl_000;
  wire ffc_832_n_spl_001;
  wire ffc_832_n_spl_01;
  wire ffc_832_n_spl_010;
  wire ffc_832_n_spl_011;
  wire ffc_832_n_spl_1;
  wire ffc_832_n_spl_10;
  wire ffc_832_n_spl_100;
  wire ffc_832_n_spl_101;
  wire ffc_832_n_spl_11;
  wire ffc_832_n_spl_110;
  wire ffc_832_n_spl_111;
  wire ffc_628_p_spl_;
  wire ffc_628_p_spl_0;
  wire ffc_833_n_spl_;
  wire ffc_833_n_spl_0;
  wire ffc_833_n_spl_00;
  wire ffc_833_n_spl_000;
  wire ffc_833_n_spl_001;
  wire ffc_833_n_spl_01;
  wire ffc_833_n_spl_010;
  wire ffc_833_n_spl_011;
  wire ffc_833_n_spl_1;
  wire ffc_833_n_spl_10;
  wire ffc_833_n_spl_100;
  wire ffc_833_n_spl_101;
  wire ffc_833_n_spl_11;
  wire ffc_833_n_spl_110;
  wire ffc_834_p_spl_;
  wire ffc_834_p_spl_0;
  wire ffc_834_p_spl_00;
  wire ffc_834_p_spl_000;
  wire ffc_834_p_spl_001;
  wire ffc_834_p_spl_01;
  wire ffc_834_p_spl_010;
  wire ffc_834_p_spl_011;
  wire ffc_834_p_spl_1;
  wire ffc_834_p_spl_10;
  wire ffc_834_p_spl_100;
  wire ffc_834_p_spl_101;
  wire ffc_834_p_spl_11;
  wire ffc_831_p_spl_;
  wire ffc_831_p_spl_0;
  wire ffc_831_p_spl_00;
  wire ffc_831_p_spl_000;
  wire ffc_831_p_spl_001;
  wire ffc_831_p_spl_01;
  wire ffc_831_p_spl_010;
  wire ffc_831_p_spl_011;
  wire ffc_831_p_spl_1;
  wire ffc_831_p_spl_10;
  wire ffc_831_p_spl_100;
  wire ffc_831_p_spl_101;
  wire ffc_831_p_spl_11;
  wire ffc_831_p_spl_110;
  wire ffc_633_n_spl_;
  wire ffc_633_p_spl_;
  wire ffc_633_p_spl_0;
  wire ffc_677_p_spl_;
  wire ffc_780_p_spl_;
  wire ffc_355_p_spl_;
  wire ffc_355_p_spl_0;
  wire ffc_346_p_spl_;
  wire ffc_366_p_spl_;
  wire ffc_367_p_spl_;
  wire ffc_826_p_spl_;
  wire ffc_826_p_spl_0;
  wire ffc_826_p_spl_1;
  wire ffc_826_n_spl_;
  wire ffc_826_n_spl_0;
  wire ffc_826_n_spl_1;
  wire ffc_812_p_spl_;
  wire g1758_p_spl_;
  wire g1758_p_spl_0;
  wire g2139_n_spl_;
  wire g2139_n_spl_0;
  wire ffc_825_n_spl_;
  wire ffc_825_n_spl_0;
  wire ffc_825_n_spl_1;
  wire g1725_n_spl_;
  wire g1758_n_spl_;
  wire g1758_n_spl_0;
  wire g1758_n_spl_1;
  wire g2142_n_spl_;
  wire ffc_671_n_spl_;
  wire ffc_671_p_spl_;
  wire ffc_671_p_spl_0;
  wire ffc_756_n_spl_;
  wire ffc_756_n_spl_0;
  wire g2146_p_spl_;
  wire ffc_756_p_spl_;
  wire ffc_756_p_spl_0;
  wire ffc_756_p_spl_1;
  wire g2146_n_spl_;
  wire ffc_672_p_spl_;
  wire ffc_778_p_spl_;
  wire ffc_825_p_spl_;
  wire ffc_825_p_spl_0;
  wire ffc_825_p_spl_1;
  wire g2139_p_spl_;
  wire g2139_p_spl_0;
  wire g2151_n_spl_;
  wire g2151_n_spl_0;
  wire g2151_p_spl_;
  wire g2151_p_spl_0;
  wire g2157_n_spl_;
  wire g1702_n_spl_;
  wire g1702_n_spl_0;
  wire g2161_p_spl_;
  wire g1702_p_spl_;
  wire g2161_n_spl_;
  wire ffc_673_n_spl_;
  wire ffc_673_p_spl_;
  wire ffc_673_p_spl_0;
  wire ffc_673_p_spl_1;
  wire g2164_n_spl_;
  wire g2165_p_spl_;
  wire g1705_p_spl_;
  wire ffc_674_p_spl_;
  wire ffc_674_p_spl_0;
  wire g2169_n_spl_;
  wire ffc_674_n_spl_;
  wire g2169_p_spl_;
  wire g2167_n_spl_;
  wire g2172_n_spl_;
  wire g2172_n_spl_0;
  wire g2096_n_spl_;
  wire g1805_p_spl_;
  wire g1808_p_spl_;
  wire ffc_629_p_spl_;
  wire ffc_358_p_spl_;
  wire ffc_622_n_spl_;
  wire ffc_622_p_spl_;
  wire ffc_622_p_spl_0;
  wire ffc_634_p_spl_;
  wire ffc_621_n_spl_;
  wire ffc_621_p_spl_;
  wire ffc_621_p_spl_0;
  wire ffc_635_p_spl_;
  wire ffc_620_n_spl_;
  wire ffc_620_p_spl_;
  wire ffc_620_p_spl_0;
  wire ffc_636_p_spl_;
  wire ffc_627_n_spl_;
  wire ffc_627_p_spl_;
  wire ffc_627_p_spl_0;
  wire ffc_650_p_spl_;
  wire ffc_632_n_spl_;
  wire ffc_632_p_spl_;
  wire ffc_632_p_spl_0;
  wire ffc_663_p_spl_;
  wire ffc_631_n_spl_;
  wire ffc_631_p_spl_;
  wire ffc_631_p_spl_0;
  wire ffc_664_p_spl_;
  wire ffc_675_n_spl_;
  wire ffc_675_p_spl_;
  wire ffc_675_p_spl_0;
  wire g1714_n_spl_;
  wire g1714_n_spl_0;
  wire g1714_p_spl_;
  wire ffc_755_p_spl_;
  wire g2253_n_spl_;
  wire ffc_755_n_spl_;
  wire g2253_p_spl_;
  wire g2250_p_spl_;
  wire g2259_n_spl_;
  wire ffc_334_p_spl_;
  wire g1768_n_spl_;
  wire g2269_p_spl_;
  wire g2272_p_spl_;
  wire g1764_p_spl_;
  wire g1764_p_spl_0;
  wire g1809_p_spl_;
  wire g2099_p_spl_;
  wire g2099_p_spl_0;
  wire g2275_n_spl_;
  wire g2108_n_spl_;
  wire g2108_n_spl_0;
  wire g2123_n_spl_;
  wire g2123_n_spl_0;
  wire g2117_n_spl_;
  wire g2117_n_spl_0;
  wire g2126_p_spl_;
  wire g2126_p_spl_0;
  wire ffc_764_p_spl_;
  wire ffc_764_p_spl_0;
  wire ffc_764_n_spl_;
  wire ffc_832_p_spl_;
  wire ffc_832_p_spl_0;
  wire ffc_832_p_spl_00;
  wire ffc_832_p_spl_1;
  wire ffc_831_n_spl_;
  wire ffc_831_n_spl_0;
  wire ffc_831_n_spl_00;
  wire ffc_831_n_spl_1;
  wire ffc_781_n_spl_;
  wire ffc_781_n_spl_0;
  wire ffc_781_n_spl_1;
  wire ffc_781_p_spl_;
  wire ffc_781_p_spl_0;
  wire ffc_781_p_spl_00;
  wire ffc_781_p_spl_1;
  wire ffc_833_p_spl_;
  wire ffc_833_p_spl_0;
  wire ffc_833_p_spl_1;
  wire ffc_834_n_spl_;
  wire ffc_834_n_spl_0;
  wire ffc_834_n_spl_1;
  wire g2120_n_spl_;
  wire g2120_n_spl_0;
  wire g2295_n_spl_;
  wire ffc_648_n_spl_;
  wire ffc_648_p_spl_;
  wire ffc_648_p_spl_0;
  wire ffc_679_p_spl_;
  wire ffc_661_p_spl_;
  wire ffc_661_p_spl_0;
  wire ffc_661_n_spl_;
  wire ffc_765_p_spl_;
  wire g2306_n_spl_;
  wire g2315_p_spl_;
  wire ffc_779_p_spl_;
  wire g1774_n_spl_;
  wire g1787_n_spl_;
  wire g1697_n_spl_;
  wire g1697_n_spl_0;
  wire g1701_p_spl_;
  wire g1697_p_spl_;
  wire g1701_n_spl_;
  wire g1701_n_spl_0;
  wire ffc_660_n_spl_;
  wire ffc_660_n_spl_0;
  wire ffc_660_n_spl_1;
  wire ffc_660_p_spl_;
  wire ffc_660_p_spl_0;
  wire ffc_660_p_spl_00;
  wire ffc_660_p_spl_1;
  wire ffc_763_p_spl_;
  wire ffc_763_p_spl_0;
  wire ffc_763_n_spl_;
  wire ffc_442_n_spl_;
  wire ffc_442_p_spl_;
  wire g1716_n_spl_;
  wire g1792_p_spl_;
  wire ffc_396_p_spl_;
  wire g2132_n_spl_;
  wire ffc_397_p_spl_;
  wire g1802_n_spl_;
  wire g2133_n_spl_;
  wire ffc_360_p_spl_;
  wire ffc_362_p_spl_;
  wire g2276_n_spl_;
  wire g2276_n_spl_0;
  wire g2137_p_spl_;
  wire g2137_p_spl_0;
  wire g2137_p_spl_1;
  wire g2160_n_spl_;
  wire g2160_n_spl_0;
  wire g2175_p_spl_;
  wire g2098_n_spl_;
  wire g2135_p_spl_;
  wire g1803_p_spl_;
  wire g1804_p_spl_;
  wire g2177_n_spl_;
  wire ffc_391_p_spl_;
  wire ffc_391_p_spl_0;
  wire g2264_n_spl_;
  wire g2264_n_spl_0;
  wire g2267_p_spl_;
  wire g2365_p_spl_;
  wire ffc_395_p_spl_;
  wire g1898_n_spl_;
  wire g2268_n_spl_;
  wire ffc_387_p_spl_;
  wire g2129_n_spl_;
  wire g2361_n_spl_;
  wire g2362_n_spl_;
  wire g2363_n_spl_;
  wire G92_p_spl_;
  wire G124_p_spl_;
  wire G124_p_spl_0;
  wire G124_p_spl_1;
  wire G124_n_spl_;
  wire G124_n_spl_0;
  wire G94_p_spl_;
  wire G107_p_spl_;
  wire ffc_401_n_spl_;
  wire ffc_401_n_spl_0;
  wire ffc_405_p_spl_;
  wire ffc_3_n_spl_;
  wire ffc_3_n_spl_0;
  wire ffc_3_n_spl_1;
  wire ffc_359_n_spl_;
  wire g1064_n_spl_;
  wire g1102_n_spl_;
  wire g1106_p_spl_;
  wire g1126_p_spl_;
  wire g1127_n_spl_;

  FA
  g_g1049_n
  (
    .dout(g1049_n),
    .din1(ffc_409_n_spl_),
    .din2(ffc_421_n_spl_)
  );


  LA
  g_g1050_p
  (
    .dout(g1050_p),
    .din1(ffc_249_p_spl_00),
    .din2(ffc_253_p)
  );


  LA
  g_g1051_p
  (
    .dout(g1051_p),
    .din1(ffc_3_p_spl_),
    .din2(ffc_382_p)
  );


  LA
  g_g1052_p
  (
    .dout(g1052_p),
    .din1(ffc_237_p),
    .din2(ffc_454_n_spl_)
  );


  FA
  g_g1053_n
  (
    .dout(g1053_n),
    .din1(ffc_42_n_spl_),
    .din2(ffc_450_p)
  );


  FA
  g_g1054_n
  (
    .dout(g1054_n),
    .din1(ffc_386_n),
    .din2(ffc_413_n)
  );


  FA
  g_g1055_n
  (
    .dout(g1055_n),
    .din1(ffc_42_n_spl_),
    .din2(ffc_46_n)
  );


  FA
  g_g1056_n
  (
    .dout(g1056_n),
    .din1(ffc_245_n),
    .din2(g1055_n_spl_000)
  );


  FA
  g_g1057_n
  (
    .dout(g1057_n),
    .din1(ffc_132_n),
    .din2(ffc_446_n_spl_00)
  );


  FA
  g_g1058_n
  (
    .dout(g1058_n),
    .din1(ffc_128_n),
    .din2(ffc_446_p_spl_00)
  );


  LA
  g_g1059_p
  (
    .dout(g1059_p),
    .din1(g1057_n),
    .din2(g1058_n)
  );


  FA
  g_g1060_n
  (
    .dout(g1060_n),
    .din1(g1055_n_spl_000),
    .din2(g1059_p)
  );


  FA
  g_g1061_n
  (
    .dout(g1061_n),
    .din1(ffc_50_n),
    .din2(ffc_446_n_spl_00)
  );


  FA
  g_g1062_n
  (
    .dout(g1062_n),
    .din1(ffc_136_n),
    .din2(ffc_446_p_spl_00)
  );


  LA
  g_g1063_p
  (
    .dout(g1063_p),
    .din1(g1061_n),
    .din2(g1062_n)
  );


  FA
  g_g1064_n
  (
    .dout(g1064_n),
    .din1(g1055_n_spl_00),
    .din2(g1063_p)
  );


  FA
  g_g1065_n
  (
    .dout(g1065_n),
    .din1(ffc_124_n),
    .din2(g1055_n_spl_01)
  );


  LA
  g_g1066_p
  (
    .dout(g1066_p),
    .din1(ffc_34_p),
    .din2(ffc_446_n_spl_01)
  );


  LA
  g_g1067_p
  (
    .dout(g1067_p),
    .din1(ffc_30_p),
    .din2(ffc_446_p_spl_01)
  );


  FA
  g_g1068_n
  (
    .dout(g1068_n),
    .din1(g1055_n_spl_01),
    .din2(g1067_p)
  );


  FA
  g_g1069_n
  (
    .dout(g1069_n),
    .din1(g1066_p),
    .din2(g1068_n)
  );


  LA
  g_g1070_p
  (
    .dout(g1070_p),
    .din1(ffc_249_p_spl_00),
    .din2(g1069_n)
  );


  LA
  g_g1071_p
  (
    .dout(g1071_p),
    .din1(ffc_116_p),
    .din2(ffc_446_n_spl_01)
  );


  LA
  g_g1072_p
  (
    .dout(g1072_p),
    .din1(ffc_38_p),
    .din2(ffc_446_p_spl_01)
  );


  FA
  g_g1073_n
  (
    .dout(g1073_n),
    .din1(g1055_n_spl_10),
    .din2(g1072_p)
  );


  FA
  g_g1074_n
  (
    .dout(g1074_n),
    .din1(g1071_p),
    .din2(g1073_n)
  );


  LA
  g_g1075_p
  (
    .dout(g1075_p),
    .din1(ffc_249_p_spl_01),
    .din2(g1074_n)
  );


  LA
  g_g1076_p
  (
    .dout(g1076_p),
    .din1(ffc_26_p),
    .din2(ffc_446_n_spl_1)
  );


  LA
  g_g1077_p
  (
    .dout(g1077_p),
    .din1(ffc_108_p),
    .din2(ffc_446_p_spl_1)
  );


  FA
  g_g1078_n
  (
    .dout(g1078_n),
    .din1(g1055_n_spl_10),
    .din2(g1077_p)
  );


  FA
  g_g1079_n
  (
    .dout(g1079_n),
    .din1(g1076_p),
    .din2(g1078_n)
  );


  LA
  g_g1080_p
  (
    .dout(g1080_p),
    .din1(ffc_249_p_spl_01),
    .din2(g1079_n)
  );


  LA
  g_g1081_p
  (
    .dout(g1081_p),
    .din1(ffc_112_p),
    .din2(ffc_446_n_spl_1)
  );


  LA
  g_g1082_p
  (
    .dout(g1082_p),
    .din1(ffc_120_p),
    .din2(ffc_446_p_spl_1)
  );


  FA
  g_g1083_n
  (
    .dout(g1083_n),
    .din1(g1055_n_spl_11),
    .din2(g1082_p)
  );


  FA
  g_g1084_n
  (
    .dout(g1084_n),
    .din1(g1081_p),
    .din2(g1083_n)
  );


  LA
  g_g1085_p
  (
    .dout(g1085_p),
    .din1(ffc_249_p_spl_1),
    .din2(g1084_n)
  );


  LA
  g_g1086_p
  (
    .dout(g1086_p),
    .din1(ffc_534_p),
    .din2(ffc_535_p)
  );


  LA
  g_g1087_p
  (
    .dout(g1087_p),
    .din1(ffc_525_n),
    .din2(ffc_618_p)
  );


  LA
  g_g1088_p
  (
    .dout(g1088_p),
    .din1(ffc_736_p),
    .din2(g1087_p)
  );


  LA
  g_g1089_p
  (
    .dout(g1089_p),
    .din1(ffc_646_p),
    .din2(ffc_737_p_spl_)
  );


  LA
  g_g1090_p
  (
    .dout(g1090_p),
    .din1(g1088_p),
    .din2(g1089_p)
  );


  LA
  g_g1091_p
  (
    .dout(g1091_p),
    .din1(g1086_p),
    .din2(g1090_p)
  );


  LA
  g_g1092_p
  (
    .dout(g1092_p),
    .din1(ffc_733_p),
    .din2(ffc_734_p)
  );


  LA
  g_g1093_p
  (
    .dout(g1093_p),
    .din1(ffc_732_p),
    .din2(g1092_p)
  );


  FA
  g_g1094_n
  (
    .dout(g1094_n),
    .din1(ffc_695_p),
    .din2(ffc_696_p)
  );


  LA
  g_g1095_p
  (
    .dout(g1095_p),
    .din1(ffc_731_p),
    .din2(g1094_n_spl_)
  );


  LA
  g_g1096_p
  (
    .dout(g1096_p),
    .din1(ffc_533_p),
    .din2(ffc_644_p)
  );


  LA
  g_g1097_p
  (
    .dout(g1097_p),
    .din1(ffc_645_p),
    .din2(ffc_735_p)
  );


  LA
  g_g1098_p
  (
    .dout(g1098_p),
    .din1(g1096_p),
    .din2(g1097_p)
  );


  LA
  g_g1099_p
  (
    .dout(g1099_p),
    .din1(g1095_p),
    .din2(g1098_p)
  );


  LA
  g_g1100_p
  (
    .dout(g1100_p),
    .din1(g1093_p),
    .din2(g1099_p)
  );


  FA
  g_g1101_n
  (
    .dout(g1101_n),
    .din1(ffc_510_n),
    .din2(ffc_519_n_spl_)
  );


  FA
  g_g1102_n
  (
    .dout(g1102_n),
    .din1(ffc_531_n),
    .din2(g1101_n_spl_)
  );


  LA
  g_g1103_p
  (
    .dout(g1103_p),
    .din1(ffc_521_p),
    .din2(ffc_545_n)
  );


  LA
  g_g1104_p
  (
    .dout(g1104_p),
    .din1(ffc_514_p),
    .din2(g1103_p)
  );


  LA
  g_g1105_p
  (
    .dout(g1105_p),
    .din1(ffc_518_p),
    .din2(ffc_599_p)
  );


  LA
  g_g1106_p
  (
    .dout(g1106_p),
    .din1(g1104_p),
    .din2(g1105_p)
  );


  LA
  g_g1107_p
  (
    .dout(g1107_p),
    .din1(ffc_747_n),
    .din2(ffc_748_n)
  );


  FA
  g_g1107_n
  (
    .dout(g1107_n),
    .din1(ffc_747_p),
    .din2(ffc_748_p)
  );


  LA
  g_g1108_p
  (
    .dout(g1108_p),
    .din1(ffc_749_n),
    .din2(ffc_750_n)
  );


  FA
  g_g1108_n
  (
    .dout(g1108_n),
    .din1(ffc_749_p),
    .din2(ffc_750_p)
  );


  LA
  g_g1109_p
  (
    .dout(g1109_p),
    .din1(g1107_n),
    .din2(g1108_p)
  );


  LA
  g_g1110_p
  (
    .dout(g1110_p),
    .din1(g1107_p),
    .din2(g1108_n)
  );


  FA
  g_g1111_n
  (
    .dout(g1111_n),
    .din1(g1109_p),
    .din2(g1110_p)
  );


  LA
  g_g1112_p
  (
    .dout(g1112_p),
    .din1(ffc_728_p_spl_),
    .din2(ffc_729_p_spl_)
  );


  FA
  g_g1112_n
  (
    .dout(g1112_n),
    .din1(ffc_728_n_spl_),
    .din2(ffc_729_n_spl_)
  );


  LA
  g_g1113_p
  (
    .dout(g1113_p),
    .din1(ffc_728_n_spl_),
    .din2(ffc_729_n_spl_)
  );


  FA
  g_g1113_n
  (
    .dout(g1113_n),
    .din1(ffc_728_p_spl_),
    .din2(ffc_729_p_spl_)
  );


  LA
  g_g1114_p
  (
    .dout(g1114_p),
    .din1(g1112_n),
    .din2(g1113_n)
  );


  FA
  g_g1114_n
  (
    .dout(g1114_n),
    .din1(g1112_p),
    .din2(g1113_p)
  );


  LA
  g_g1115_p
  (
    .dout(g1115_p),
    .din1(ffc_730_n_spl_),
    .din2(ffc_753_n_spl_)
  );


  FA
  g_g1115_n
  (
    .dout(g1115_n),
    .din1(ffc_730_p_spl_),
    .din2(ffc_753_p_spl_)
  );


  LA
  g_g1116_p
  (
    .dout(g1116_p),
    .din1(ffc_730_p_spl_),
    .din2(ffc_753_p_spl_)
  );


  FA
  g_g1116_n
  (
    .dout(g1116_n),
    .din1(ffc_730_n_spl_),
    .din2(ffc_753_n_spl_)
  );


  LA
  g_g1117_p
  (
    .dout(g1117_p),
    .din1(g1115_n),
    .din2(g1116_n)
  );


  FA
  g_g1117_n
  (
    .dout(g1117_n),
    .din1(g1115_p),
    .din2(g1116_p)
  );


  LA
  g_g1118_p
  (
    .dout(g1118_p),
    .din1(g1114_n),
    .din2(g1117_p)
  );


  LA
  g_g1119_p
  (
    .dout(g1119_p),
    .din1(g1114_p),
    .din2(g1117_n)
  );


  FA
  g_g1120_n
  (
    .dout(g1120_n),
    .din1(g1118_p),
    .din2(g1119_p)
  );


  FA
  g_g1121_n
  (
    .dout(g1121_n),
    .din1(ffc_530_n),
    .din2(g1101_n_spl_)
  );


  FA
  g_g1122_n
  (
    .dout(g1122_n),
    .din1(ffc_515_n),
    .din2(ffc_519_n_spl_)
  );


  FA
  g_g1123_n
  (
    .dout(g1123_n),
    .din1(ffc_509_n),
    .din2(ffc_517_n)
  );


  LA
  g_g1124_p
  (
    .dout(g1124_p),
    .din1(ffc_513_n),
    .din2(g1123_n)
  );


  LA
  g_g1125_p
  (
    .dout(g1125_p),
    .din1(g1122_n),
    .din2(g1124_p)
  );


  LA
  g_g1126_p
  (
    .dout(g1126_p),
    .din1(g1121_n),
    .din2(g1125_p)
  );


  FA
  g_g1127_n
  (
    .dout(g1127_n),
    .din1(ffc_516_n),
    .din2(ffc_532_p_spl_0)
  );


  LA
  g_g1128_p
  (
    .dout(g1128_p),
    .din1(ffc_643_n),
    .din2(ffc_697_p_spl_000)
  );


  FA
  g_g1129_n
  (
    .dout(g1129_n),
    .din1(ffc_498_n_spl_000),
    .din2(ffc_525_p)
  );


  LA
  g_g1130_p
  (
    .dout(g1130_p),
    .din1(ffc_494_p_spl_000),
    .din2(ffc_694_p)
  );


  LA
  g_g1131_p
  (
    .dout(g1131_p),
    .din1(g1129_n),
    .din2(g1130_p)
  );


  FA
  g_g1132_n
  (
    .dout(g1132_n),
    .din1(g1128_p),
    .din2(g1131_p)
  );


  FA
  g_g1133_n
  (
    .dout(g1133_n),
    .din1(ffc_520_n),
    .din2(ffc_697_n_spl_)
  );


  LA
  g_g1134_p
  (
    .dout(g1134_p),
    .din1(ffc_498_p_spl_000),
    .din2(ffc_737_p_spl_)
  );


  FA
  g_g1135_n
  (
    .dout(g1135_n),
    .din1(ffc_494_n_spl_0),
    .din2(ffc_693_n)
  );


  FA
  g_g1136_n
  (
    .dout(g1136_n),
    .din1(g1134_p),
    .din2(g1135_n)
  );


  LA
  g_g1137_p
  (
    .dout(g1137_p),
    .din1(g1133_n),
    .din2(g1136_n)
  );


  LA
  g_g1138_p
  (
    .dout(g1138_p),
    .din1(ffc_697_p_spl_000),
    .din2(ffc_723_p_spl_)
  );


  FA
  g_g1139_n
  (
    .dout(g1139_n),
    .din1(ffc_498_n_spl_000),
    .din2(ffc_731_n)
  );


  LA
  g_g1140_p
  (
    .dout(g1140_p),
    .din1(ffc_494_p_spl_000),
    .din2(ffc_689_p)
  );


  LA
  g_g1141_p
  (
    .dout(g1141_p),
    .din1(g1139_n),
    .din2(g1140_p)
  );


  FA
  g_g1142_n
  (
    .dout(g1142_n),
    .din1(g1138_p),
    .din2(g1141_p)
  );


  FA
  g_g1143_n
  (
    .dout(g1143_n),
    .din1(ffc_482_n_spl_0000),
    .din2(g1132_n_spl_00)
  );


  FA
  g_g1144_n
  (
    .dout(g1144_n),
    .din1(ffc_482_p_spl_0000),
    .din2(g1142_n_spl_00)
  );


  LA
  g_g1145_p
  (
    .dout(g1145_p),
    .din1(g1143_n),
    .din2(g1144_n)
  );


  LA
  g_g1146_p
  (
    .dout(g1146_p),
    .din1(ffc_478_p_spl_000),
    .din2(g1145_p)
  );


  FA
  g_g1147_n
  (
    .dout(g1147_n),
    .din1(ffc_10_p_spl_),
    .din2(ffc_482_n_spl_0000)
  );


  FA
  g_g1148_n
  (
    .dout(g1148_n),
    .din1(ffc_84_p_spl_),
    .din2(ffc_482_p_spl_0000)
  );


  LA
  g_g1149_p
  (
    .dout(g1149_p),
    .din1(g1147_n),
    .din2(g1148_n)
  );


  LA
  g_g1150_p
  (
    .dout(g1150_p),
    .din1(ffc_478_n_spl_000),
    .din2(g1149_p)
  );


  FA
  g_g1151_n
  (
    .dout(g1151_n),
    .din1(g1146_p),
    .din2(g1150_p)
  );


  LA
  g_g1152_p
  (
    .dout(g1152_p),
    .din1(ffc_523_n_spl_),
    .din2(ffc_697_p_spl_001)
  );


  FA
  g_g1153_n
  (
    .dout(g1153_n),
    .din1(ffc_686_p),
    .din2(ffc_700_p)
  );


  LA
  g_g1154_p
  (
    .dout(g1154_p),
    .din1(ffc_494_p_spl_001),
    .din2(g1153_n)
  );


  FA
  g_g1155_n
  (
    .dout(g1155_n),
    .din1(g1152_p),
    .din2(g1154_p)
  );


  LA
  g_g1156_p
  (
    .dout(g1156_p),
    .din1(ffc_697_p_spl_001),
    .din2(ffc_744_n_spl_)
  );


  LA
  g_g1157_p
  (
    .dout(g1157_p),
    .din1(ffc_494_p_spl_001),
    .din2(ffc_727_p)
  );


  FA
  g_g1158_n
  (
    .dout(g1158_n),
    .din1(g1156_p),
    .din2(g1157_p)
  );


  FA
  g_g1159_n
  (
    .dout(g1159_n),
    .din1(ffc_718_p),
    .din2(ffc_719_n)
  );


  LA
  g_g1160_p
  (
    .dout(g1160_p),
    .din1(ffc_697_p_spl_010),
    .din2(g1159_n_spl_)
  );


  FA
  g_g1161_n
  (
    .dout(g1161_n),
    .din1(ffc_498_n_spl_00),
    .din2(ffc_736_n)
  );


  LA
  g_g1162_p
  (
    .dout(g1162_p),
    .din1(ffc_494_p_spl_010),
    .din2(ffc_690_p)
  );


  LA
  g_g1163_p
  (
    .dout(g1163_p),
    .din1(g1161_n),
    .din2(g1162_p)
  );


  FA
  g_g1164_n
  (
    .dout(g1164_n),
    .din1(g1160_p),
    .din2(g1163_p)
  );


  FA
  g_g1165_n
  (
    .dout(g1165_n),
    .din1(ffc_486_n_spl_0000),
    .din2(g1132_n_spl_00)
  );


  FA
  g_g1166_n
  (
    .dout(g1166_n),
    .din1(ffc_486_p_spl_0000),
    .din2(g1142_n_spl_00)
  );


  LA
  g_g1167_p
  (
    .dout(g1167_p),
    .din1(g1165_n),
    .din2(g1166_n)
  );


  LA
  g_g1168_p
  (
    .dout(g1168_p),
    .din1(ffc_490_p_spl_000),
    .din2(g1167_p)
  );


  FA
  g_g1169_n
  (
    .dout(g1169_n),
    .din1(ffc_10_p_spl_),
    .din2(ffc_486_n_spl_0000)
  );


  FA
  g_g1170_n
  (
    .dout(g1170_n),
    .din1(ffc_84_p_spl_),
    .din2(ffc_486_p_spl_0000)
  );


  LA
  g_g1171_p
  (
    .dout(g1171_p),
    .din1(g1169_n),
    .din2(g1170_n)
  );


  LA
  g_g1172_p
  (
    .dout(g1172_p),
    .din1(ffc_490_n_spl_000),
    .din2(g1171_p)
  );


  FA
  g_g1173_n
  (
    .dout(g1173_n),
    .din1(g1168_p),
    .din2(g1172_p)
  );


  LA
  g_g1174_p
  (
    .dout(g1174_p),
    .din1(ffc_522_n),
    .din2(ffc_714_n)
  );


  LA
  g_g1175_p
  (
    .dout(g1175_p),
    .din1(ffc_522_p),
    .din2(ffc_714_p)
  );


  FA
  g_g1176_n
  (
    .dout(g1176_n),
    .din1(g1174_p),
    .din2(g1175_p)
  );


  LA
  g_g1177_p
  (
    .dout(g1177_p),
    .din1(ffc_697_p_spl_010),
    .din2(g1176_n_spl_)
  );


  LA
  g_g1178_p
  (
    .dout(g1178_p),
    .din1(ffc_201_p),
    .din2(ffc_498_n_spl_01)
  );


  LA
  g_g1179_p
  (
    .dout(g1179_p),
    .din1(ffc_498_p_spl_000),
    .din2(ffc_733_n)
  );


  FA
  g_g1180_n
  (
    .dout(g1180_n),
    .din1(g1178_p),
    .din2(g1179_p)
  );


  LA
  g_g1181_p
  (
    .dout(g1181_p),
    .din1(ffc_494_p_spl_010),
    .din2(g1180_n)
  );


  FA
  g_g1182_n
  (
    .dout(g1182_n),
    .din1(g1177_p),
    .din2(g1181_p)
  );


  FA
  g_g1183_n
  (
    .dout(g1183_n),
    .din1(ffc_641_p),
    .din2(ffc_717_n)
  );


  LA
  g_g1184_p
  (
    .dout(g1184_p),
    .din1(ffc_697_p_spl_011),
    .din2(g1183_n_spl_)
  );


  FA
  g_g1185_n
  (
    .dout(g1185_n),
    .din1(ffc_692_p),
    .din2(ffc_701_p)
  );


  LA
  g_g1186_p
  (
    .dout(g1186_p),
    .din1(ffc_494_p_spl_011),
    .din2(g1185_n)
  );


  FA
  g_g1187_n
  (
    .dout(g1187_n),
    .din1(g1184_p),
    .din2(g1186_p)
  );


  FA
  g_g1188_n
  (
    .dout(g1188_n),
    .din1(ffc_600_p),
    .din2(ffc_713_n)
  );


  LA
  g_g1189_p
  (
    .dout(g1189_p),
    .din1(ffc_697_p_spl_011),
    .din2(g1188_n_spl_)
  );


  LA
  g_g1190_p
  (
    .dout(g1190_p),
    .din1(ffc_213_p),
    .din2(ffc_498_n_spl_01)
  );


  LA
  g_g1191_p
  (
    .dout(g1191_p),
    .din1(ffc_498_p_spl_00),
    .din2(ffc_732_n)
  );


  FA
  g_g1192_n
  (
    .dout(g1192_n),
    .din1(g1190_p),
    .din2(g1191_p)
  );


  LA
  g_g1193_p
  (
    .dout(g1193_p),
    .din1(ffc_494_p_spl_011),
    .din2(g1192_n)
  );


  FA
  g_g1194_n
  (
    .dout(g1194_n),
    .din1(g1189_p),
    .din2(g1193_p)
  );


  FA
  g_g1195_n
  (
    .dout(g1195_n),
    .din1(ffc_697_n_spl_),
    .din2(ffc_741_p)
  );


  LA
  g_g1196_p
  (
    .dout(g1196_p),
    .din1(ffc_498_p_spl_01),
    .din2(g1094_n_spl_)
  );


  LA
  g_g1197_p
  (
    .dout(g1197_p),
    .din1(ffc_209_n),
    .din2(ffc_498_n_spl_10)
  );


  FA
  g_g1198_n
  (
    .dout(g1198_n),
    .din1(ffc_494_n_spl_0),
    .din2(g1197_p)
  );


  FA
  g_g1199_n
  (
    .dout(g1199_n),
    .din1(g1196_p),
    .din2(g1198_n)
  );


  LA
  g_g1200_p
  (
    .dout(g1200_p),
    .din1(g1195_n),
    .din2(g1199_n)
  );


  LA
  g_g1201_p
  (
    .dout(g1201_p),
    .din1(ffc_707_n),
    .din2(ffc_708_n)
  );


  FA
  g_g1201_n
  (
    .dout(g1201_n),
    .din1(ffc_707_p),
    .din2(ffc_708_p)
  );


  LA
  g_g1202_p
  (
    .dout(g1202_p),
    .din1(ffc_561_n_spl_00),
    .din2(g1201_n_spl_)
  );


  FA
  g_g1202_n
  (
    .dout(g1202_n),
    .din1(ffc_561_p_spl_0),
    .din2(g1201_p_spl_)
  );


  LA
  g_g1203_p
  (
    .dout(g1203_p),
    .din1(ffc_561_p_spl_0),
    .din2(g1201_p_spl_)
  );


  FA
  g_g1203_n
  (
    .dout(g1203_n),
    .din1(ffc_561_n_spl_00),
    .din2(g1201_n_spl_)
  );


  LA
  g_g1204_p
  (
    .dout(g1204_p),
    .din1(g1202_n),
    .din2(g1203_n)
  );


  FA
  g_g1204_n
  (
    .dout(g1204_n),
    .din1(g1202_p),
    .din2(g1203_p)
  );


  LA
  g_g1205_p
  (
    .dout(g1205_p),
    .din1(ffc_715_p),
    .din2(ffc_716_n)
  );


  FA
  g_g1205_n
  (
    .dout(g1205_n),
    .din1(ffc_715_n),
    .din2(ffc_716_p)
  );


  LA
  g_g1206_p
  (
    .dout(g1206_p),
    .din1(ffc_751_p),
    .din2(ffc_752_n)
  );


  FA
  g_g1206_n
  (
    .dout(g1206_n),
    .din1(ffc_751_n),
    .din2(ffc_752_p)
  );


  LA
  g_g1207_p
  (
    .dout(g1207_p),
    .din1(g1205_p_spl_),
    .din2(g1206_n_spl_)
  );


  FA
  g_g1207_n
  (
    .dout(g1207_n),
    .din1(g1205_n_spl_),
    .din2(g1206_p_spl_)
  );


  LA
  g_g1208_p
  (
    .dout(g1208_p),
    .din1(g1205_n_spl_),
    .din2(g1206_p_spl_)
  );


  FA
  g_g1208_n
  (
    .dout(g1208_n),
    .din1(g1205_p_spl_),
    .din2(g1206_n_spl_)
  );


  LA
  g_g1209_p
  (
    .dout(g1209_p),
    .din1(g1207_n),
    .din2(g1208_n)
  );


  FA
  g_g1209_n
  (
    .dout(g1209_n),
    .din1(g1207_p),
    .din2(g1208_p)
  );


  LA
  g_g1210_p
  (
    .dout(g1210_p),
    .din1(g1204_n),
    .din2(g1209_p)
  );


  LA
  g_g1211_p
  (
    .dout(g1211_p),
    .din1(g1204_p),
    .din2(g1209_n)
  );


  FA
  g_g1212_n
  (
    .dout(g1212_n),
    .din1(g1210_p),
    .din2(g1211_p)
  );


  LA
  g_g1213_p
  (
    .dout(g1213_p),
    .din1(ffc_504_n_spl_),
    .din2(ffc_505_p_spl_)
  );


  FA
  g_g1213_n
  (
    .dout(g1213_n),
    .din1(ffc_504_p_spl_),
    .din2(ffc_505_n_spl_)
  );


  LA
  g_g1214_p
  (
    .dout(g1214_p),
    .din1(ffc_504_p_spl_),
    .din2(ffc_505_n_spl_)
  );


  FA
  g_g1214_n
  (
    .dout(g1214_n),
    .din1(ffc_504_n_spl_),
    .din2(ffc_505_p_spl_)
  );


  LA
  g_g1215_p
  (
    .dout(g1215_p),
    .din1(g1213_n),
    .din2(g1214_n)
  );


  FA
  g_g1215_n
  (
    .dout(g1215_n),
    .din1(g1213_p),
    .din2(g1214_p)
  );


  LA
  g_g1216_p
  (
    .dout(g1216_p),
    .din1(ffc_507_n_spl_),
    .din2(ffc_511_p_spl_)
  );


  FA
  g_g1216_n
  (
    .dout(g1216_n),
    .din1(ffc_507_p_spl_),
    .din2(ffc_511_n_spl_)
  );


  LA
  g_g1217_p
  (
    .dout(g1217_p),
    .din1(ffc_507_p_spl_),
    .din2(ffc_511_n_spl_)
  );


  FA
  g_g1217_n
  (
    .dout(g1217_n),
    .din1(ffc_507_n_spl_),
    .din2(ffc_511_p_spl_)
  );


  LA
  g_g1218_p
  (
    .dout(g1218_p),
    .din1(g1216_n),
    .din2(g1217_n)
  );


  FA
  g_g1218_n
  (
    .dout(g1218_n),
    .din1(g1216_p),
    .din2(g1217_p)
  );


  LA
  g_g1219_p
  (
    .dout(g1219_p),
    .din1(g1215_n_spl_),
    .din2(g1218_p_spl_)
  );


  FA
  g_g1219_n
  (
    .dout(g1219_n),
    .din1(g1215_p_spl_),
    .din2(g1218_n_spl_)
  );


  LA
  g_g1220_p
  (
    .dout(g1220_p),
    .din1(g1215_p_spl_),
    .din2(g1218_n_spl_)
  );


  FA
  g_g1220_n
  (
    .dout(g1220_n),
    .din1(g1215_n_spl_),
    .din2(g1218_p_spl_)
  );


  LA
  g_g1221_p
  (
    .dout(g1221_p),
    .din1(g1219_n),
    .din2(g1220_n)
  );


  FA
  g_g1221_n
  (
    .dout(g1221_n),
    .din1(g1219_p),
    .din2(g1220_p)
  );


  LA
  g_g1222_p
  (
    .dout(g1222_p),
    .din1(ffc_739_n_spl_),
    .din2(ffc_742_p_spl_)
  );


  FA
  g_g1222_n
  (
    .dout(g1222_n),
    .din1(ffc_739_p_spl_),
    .din2(ffc_742_n_spl_)
  );


  LA
  g_g1223_p
  (
    .dout(g1223_p),
    .din1(ffc_739_p_spl_),
    .din2(ffc_742_n_spl_)
  );


  FA
  g_g1223_n
  (
    .dout(g1223_n),
    .din1(ffc_739_n_spl_),
    .din2(ffc_742_p_spl_)
  );


  LA
  g_g1224_p
  (
    .dout(g1224_p),
    .din1(g1222_n),
    .din2(g1223_n)
  );


  FA
  g_g1224_n
  (
    .dout(g1224_n),
    .din1(g1222_p),
    .din2(g1223_p)
  );


  LA
  g_g1225_p
  (
    .dout(g1225_p),
    .din1(ffc_503_p_spl_),
    .din2(ffc_506_n_spl_)
  );


  FA
  g_g1225_n
  (
    .dout(g1225_n),
    .din1(ffc_503_n_spl_),
    .din2(ffc_506_p_spl_)
  );


  LA
  g_g1226_p
  (
    .dout(g1226_p),
    .din1(ffc_503_n_spl_),
    .din2(ffc_506_p_spl_)
  );


  FA
  g_g1226_n
  (
    .dout(g1226_n),
    .din1(ffc_503_p_spl_),
    .din2(ffc_506_n_spl_)
  );


  LA
  g_g1227_p
  (
    .dout(g1227_p),
    .din1(g1225_n),
    .din2(g1226_n)
  );


  FA
  g_g1227_n
  (
    .dout(g1227_n),
    .din1(g1225_p),
    .din2(g1226_p)
  );


  LA
  g_g1228_p
  (
    .dout(g1228_p),
    .din1(g1224_n_spl_),
    .din2(g1227_p_spl_)
  );


  FA
  g_g1228_n
  (
    .dout(g1228_n),
    .din1(g1224_p_spl_),
    .din2(g1227_n_spl_)
  );


  LA
  g_g1229_p
  (
    .dout(g1229_p),
    .din1(g1224_p_spl_),
    .din2(g1227_n_spl_)
  );


  FA
  g_g1229_n
  (
    .dout(g1229_n),
    .din1(g1224_n_spl_),
    .din2(g1227_p_spl_)
  );


  LA
  g_g1230_p
  (
    .dout(g1230_p),
    .din1(g1228_n),
    .din2(g1229_n)
  );


  FA
  g_g1230_n
  (
    .dout(g1230_n),
    .din1(g1228_p),
    .din2(g1229_p)
  );


  LA
  g_g1231_p
  (
    .dout(g1231_p),
    .din1(g1221_n),
    .din2(g1230_p)
  );


  LA
  g_g1232_p
  (
    .dout(g1232_p),
    .din1(g1221_p),
    .din2(g1230_n)
  );


  FA
  g_g1233_n
  (
    .dout(g1233_n),
    .din1(g1231_p),
    .din2(g1232_p)
  );


  FA
  g_g1234_n
  (
    .dout(g1234_n),
    .din1(ffc_709_p),
    .din2(ffc_710_p)
  );


  FA
  g_g1235_n
  (
    .dout(g1235_n),
    .din1(ffc_723_p_spl_),
    .din2(ffc_741_n)
  );


  FA
  g_g1236_n
  (
    .dout(g1236_n),
    .din1(g1188_n_spl_),
    .din2(g1235_n)
  );


  FA
  g_g1237_n
  (
    .dout(g1237_n),
    .din1(g1183_n_spl_),
    .din2(g1236_n)
  );


  FA
  g_g1238_n
  (
    .dout(g1238_n),
    .din1(g1176_n_spl_),
    .din2(g1237_n)
  );


  FA
  g_g1239_n
  (
    .dout(g1239_n),
    .din1(g1234_n_spl_),
    .din2(g1238_n)
  );


  FA
  g_g1240_n
  (
    .dout(g1240_n),
    .din1(ffc_745_n_spl_),
    .din2(g1239_n)
  );


  FA
  g_g1241_n
  (
    .dout(g1241_n),
    .din1(ffc_512_n),
    .din2(ffc_743_p)
  );


  FA
  g_g1242_n
  (
    .dout(g1242_n),
    .din1(ffc_512_p),
    .din2(ffc_743_n)
  );


  LA
  g_g1243_p
  (
    .dout(g1243_p),
    .din1(g1241_n),
    .din2(g1242_n)
  );


  FA
  g_g1244_n
  (
    .dout(g1244_n),
    .din1(ffc_508_n),
    .din2(ffc_740_n)
  );


  FA
  g_g1245_n
  (
    .dout(g1245_n),
    .din1(ffc_508_p),
    .din2(ffc_740_p)
  );


  LA
  g_g1246_p
  (
    .dout(g1246_p),
    .din1(g1244_n),
    .din2(g1245_n)
  );


  FA
  g_g1247_n
  (
    .dout(g1247_n),
    .din1(g1243_p_spl_),
    .din2(g1246_p_spl_)
  );


  FA
  g_g1248_n
  (
    .dout(g1248_n),
    .din1(g1240_n),
    .din2(g1247_n)
  );


  LA
  g_g1249_p
  (
    .dout(g1249_p),
    .din1(ffc_720_p),
    .din2(ffc_721_n)
  );


  LA
  g_g1250_p
  (
    .dout(g1250_p),
    .din1(ffc_711_n),
    .din2(ffc_712_p)
  );


  FA
  g_g1251_n
  (
    .dout(g1251_n),
    .din1(ffc_520_p),
    .din2(ffc_722_n)
  );


  FA
  g_g1252_n
  (
    .dout(g1252_n),
    .din1(g1159_n_spl_),
    .din2(g1251_n)
  );


  FA
  g_g1253_n
  (
    .dout(g1253_n),
    .din1(ffc_523_n_spl_),
    .din2(g1252_n)
  );


  FA
  g_g1254_n
  (
    .dout(g1254_n),
    .din1(ffc_744_n_spl_),
    .din2(g1253_n)
  );


  FA
  g_g1255_n
  (
    .dout(g1255_n),
    .din1(ffc_746_p_spl_),
    .din2(g1254_n)
  );


  FA
  g_g1256_n
  (
    .dout(g1256_n),
    .din1(g1250_p_spl_),
    .din2(g1255_n)
  );


  FA
  g_g1257_n
  (
    .dout(g1257_n),
    .din1(g1249_p_spl_),
    .din2(g1256_n)
  );


  LA
  g_g1258_p
  (
    .dout(g1258_p),
    .din1(ffc_428_n_spl_0000),
    .din2(g1142_n_spl_0)
  );


  LA
  g_g1259_p
  (
    .dout(g1259_p),
    .din1(ffc_428_p_spl_0000),
    .din2(g1132_n_spl_0)
  );


  FA
  g_g1260_n
  (
    .dout(g1260_n),
    .din1(ffc_432_n_spl_000),
    .din2(g1259_p)
  );


  FA
  g_g1261_n
  (
    .dout(g1261_n),
    .din1(g1258_p),
    .din2(g1260_n)
  );


  LA
  g_g1262_p
  (
    .dout(g1262_p),
    .din1(ffc_309_p_spl_),
    .din2(ffc_428_n_spl_0000)
  );


  LA
  g_g1263_p
  (
    .dout(g1263_p),
    .din1(ffc_305_p_spl_),
    .din2(ffc_428_p_spl_0000)
  );


  FA
  g_g1264_n
  (
    .dout(g1264_n),
    .din1(ffc_432_p_spl_000),
    .din2(g1263_p)
  );


  FA
  g_g1265_n
  (
    .dout(g1265_n),
    .din1(g1262_p),
    .din2(g1264_n)
  );


  LA
  g_g1266_p
  (
    .dout(g1266_p),
    .din1(ffc_241_p_spl_0000),
    .din2(g1265_n)
  );


  LA
  g_g1267_p
  (
    .dout(g1267_p),
    .din1(g1261_n),
    .din2(g1266_p)
  );


  LA
  g_g1268_p
  (
    .dout(g1268_p),
    .din1(ffc_436_n_spl_0000),
    .din2(g1142_n_spl_1)
  );


  LA
  g_g1269_p
  (
    .dout(g1269_p),
    .din1(ffc_436_p_spl_0000),
    .din2(g1132_n_spl_1)
  );


  FA
  g_g1270_n
  (
    .dout(g1270_n),
    .din1(ffc_440_n_spl_000),
    .din2(g1269_p)
  );


  FA
  g_g1271_n
  (
    .dout(g1271_n),
    .din1(g1268_p),
    .din2(g1270_n)
  );


  LA
  g_g1272_p
  (
    .dout(g1272_p),
    .din1(ffc_309_p_spl_),
    .din2(ffc_436_n_spl_0000)
  );


  LA
  g_g1273_p
  (
    .dout(g1273_p),
    .din1(ffc_305_p_spl_),
    .din2(ffc_436_p_spl_0000)
  );


  FA
  g_g1274_n
  (
    .dout(g1274_n),
    .din1(ffc_440_p_spl_000),
    .din2(g1273_p)
  );


  FA
  g_g1275_n
  (
    .dout(g1275_n),
    .din1(g1272_p),
    .din2(g1274_n)
  );


  LA
  g_g1276_p
  (
    .dout(g1276_p),
    .din1(ffc_241_p_spl_0000),
    .din2(g1275_n)
  );


  LA
  g_g1277_p
  (
    .dout(g1277_p),
    .din1(g1271_n),
    .din2(g1276_p)
  );


  FA
  g_g1278_n
  (
    .dout(g1278_n),
    .din1(ffc_54_p_spl_),
    .din2(ffc_482_p_spl_0001)
  );


  FA
  g_g1279_n
  (
    .dout(g1279_n),
    .din1(ffc_62_p_spl_),
    .din2(ffc_482_n_spl_0001)
  );


  LA
  g_g1280_p
  (
    .dout(g1280_p),
    .din1(g1278_n),
    .din2(g1279_n)
  );


  FA
  g_g1281_n
  (
    .dout(g1281_n),
    .din1(ffc_478_p_spl_000),
    .din2(g1280_p)
  );


  LA
  g_g1282_p
  (
    .dout(g1282_p),
    .din1(ffc_482_n_spl_0001),
    .din2(g1182_n_spl_00)
  );


  LA
  g_g1283_p
  (
    .dout(g1283_p),
    .din1(ffc_482_p_spl_0001),
    .din2(g1155_n_spl_00)
  );


  FA
  g_g1284_n
  (
    .dout(g1284_n),
    .din1(ffc_478_n_spl_000),
    .din2(g1283_p)
  );


  FA
  g_g1285_n
  (
    .dout(g1285_n),
    .din1(g1282_p),
    .din2(g1284_n)
  );


  LA
  g_g1286_p
  (
    .dout(g1286_p),
    .din1(g1281_n),
    .din2(g1285_n)
  );


  FA
  g_g1287_n
  (
    .dout(g1287_n),
    .din1(ffc_22_p_spl_),
    .din2(ffc_482_p_spl_0010)
  );


  FA
  g_g1288_n
  (
    .dout(g1288_n),
    .din1(ffc_104_p_spl_),
    .din2(ffc_482_n_spl_0010)
  );


  LA
  g_g1289_p
  (
    .dout(g1289_p),
    .din1(g1287_n),
    .din2(g1288_n)
  );


  FA
  g_g1290_n
  (
    .dout(g1290_n),
    .din1(ffc_478_p_spl_001),
    .din2(g1289_p)
  );


  LA
  g_g1291_p
  (
    .dout(g1291_p),
    .din1(ffc_482_n_spl_0010),
    .din2(g1187_n_spl_00)
  );


  LA
  g_g1292_p
  (
    .dout(g1292_p),
    .din1(ffc_482_p_spl_0010),
    .din2(g1158_n_spl_00)
  );


  FA
  g_g1293_n
  (
    .dout(g1293_n),
    .din1(ffc_478_n_spl_001),
    .din2(g1292_p)
  );


  FA
  g_g1294_n
  (
    .dout(g1294_n),
    .din1(g1291_p),
    .din2(g1293_n)
  );


  LA
  g_g1295_p
  (
    .dout(g1295_p),
    .din1(g1290_n),
    .din2(g1294_n)
  );


  FA
  g_g1296_n
  (
    .dout(g1296_n),
    .din1(ffc_18_p_spl_),
    .din2(ffc_482_p_spl_0011)
  );


  FA
  g_g1297_n
  (
    .dout(g1297_n),
    .din1(ffc_100_p_spl_),
    .din2(ffc_482_n_spl_0011)
  );


  LA
  g_g1298_p
  (
    .dout(g1298_p),
    .din1(g1296_n),
    .din2(g1297_n)
  );


  FA
  g_g1299_n
  (
    .dout(g1299_n),
    .din1(ffc_478_p_spl_001),
    .din2(g1298_p)
  );


  LA
  g_g1300_p
  (
    .dout(g1300_p),
    .din1(ffc_482_n_spl_0011),
    .din2(g1194_n_spl_00)
  );


  LA
  g_g1301_p
  (
    .dout(g1301_p),
    .din1(ffc_482_p_spl_0011),
    .din2(g1164_n_spl_00)
  );


  FA
  g_g1302_n
  (
    .dout(g1302_n),
    .din1(ffc_478_n_spl_001),
    .din2(g1301_p)
  );


  FA
  g_g1303_n
  (
    .dout(g1303_n),
    .din1(g1300_p),
    .din2(g1302_n)
  );


  LA
  g_g1304_p
  (
    .dout(g1304_p),
    .din1(g1299_n),
    .din2(g1303_n)
  );


  FA
  g_g1305_n
  (
    .dout(g1305_n),
    .din1(ffc_96_n_spl_),
    .din2(ffc_482_p_spl_010)
  );


  FA
  g_g1306_n
  (
    .dout(g1306_n),
    .din1(ffc_92_n_spl_),
    .din2(ffc_482_n_spl_010)
  );


  LA
  g_g1307_p
  (
    .dout(g1307_p),
    .din1(g1305_n),
    .din2(g1306_n)
  );


  FA
  g_g1308_n
  (
    .dout(g1308_n),
    .din1(ffc_478_p_spl_01),
    .din2(g1307_p)
  );


  LA
  g_g1309_p
  (
    .dout(g1309_p),
    .din1(ffc_482_n_spl_010),
    .din2(g1200_p_spl_00)
  );


  LA
  g_g1310_p
  (
    .dout(g1310_p),
    .din1(ffc_482_p_spl_010),
    .din2(g1137_p_spl_00)
  );


  FA
  g_g1311_n
  (
    .dout(g1311_n),
    .din1(ffc_478_n_spl_01),
    .din2(g1310_p)
  );


  FA
  g_g1312_n
  (
    .dout(g1312_n),
    .din1(g1309_p),
    .din2(g1311_n)
  );


  LA
  g_g1313_p
  (
    .dout(g1313_p),
    .din1(g1308_n),
    .din2(g1312_n)
  );


  FA
  g_g1314_n
  (
    .dout(g1314_n),
    .din1(ffc_54_p_spl_),
    .din2(ffc_486_p_spl_0001)
  );


  FA
  g_g1315_n
  (
    .dout(g1315_n),
    .din1(ffc_62_p_spl_),
    .din2(ffc_486_n_spl_0001)
  );


  LA
  g_g1316_p
  (
    .dout(g1316_p),
    .din1(g1314_n),
    .din2(g1315_n)
  );


  FA
  g_g1317_n
  (
    .dout(g1317_n),
    .din1(ffc_490_p_spl_000),
    .din2(g1316_p)
  );


  LA
  g_g1318_p
  (
    .dout(g1318_p),
    .din1(ffc_486_n_spl_0001),
    .din2(g1182_n_spl_00)
  );


  LA
  g_g1319_p
  (
    .dout(g1319_p),
    .din1(ffc_486_p_spl_0001),
    .din2(g1155_n_spl_00)
  );


  FA
  g_g1320_n
  (
    .dout(g1320_n),
    .din1(ffc_490_n_spl_000),
    .din2(g1319_p)
  );


  FA
  g_g1321_n
  (
    .dout(g1321_n),
    .din1(g1318_p),
    .din2(g1320_n)
  );


  LA
  g_g1322_p
  (
    .dout(g1322_p),
    .din1(g1317_n),
    .din2(g1321_n)
  );


  FA
  g_g1323_n
  (
    .dout(g1323_n),
    .din1(ffc_22_p_spl_),
    .din2(ffc_486_p_spl_0010)
  );


  FA
  g_g1324_n
  (
    .dout(g1324_n),
    .din1(ffc_104_p_spl_),
    .din2(ffc_486_n_spl_0010)
  );


  LA
  g_g1325_p
  (
    .dout(g1325_p),
    .din1(g1323_n),
    .din2(g1324_n)
  );


  FA
  g_g1326_n
  (
    .dout(g1326_n),
    .din1(ffc_490_p_spl_001),
    .din2(g1325_p)
  );


  LA
  g_g1327_p
  (
    .dout(g1327_p),
    .din1(ffc_486_n_spl_0010),
    .din2(g1187_n_spl_00)
  );


  LA
  g_g1328_p
  (
    .dout(g1328_p),
    .din1(ffc_486_p_spl_0010),
    .din2(g1158_n_spl_00)
  );


  FA
  g_g1329_n
  (
    .dout(g1329_n),
    .din1(ffc_490_n_spl_001),
    .din2(g1328_p)
  );


  FA
  g_g1330_n
  (
    .dout(g1330_n),
    .din1(g1327_p),
    .din2(g1329_n)
  );


  LA
  g_g1331_p
  (
    .dout(g1331_p),
    .din1(g1326_n),
    .din2(g1330_n)
  );


  FA
  g_g1332_n
  (
    .dout(g1332_n),
    .din1(ffc_18_p_spl_),
    .din2(ffc_486_p_spl_0011)
  );


  FA
  g_g1333_n
  (
    .dout(g1333_n),
    .din1(ffc_100_p_spl_),
    .din2(ffc_486_n_spl_0011)
  );


  LA
  g_g1334_p
  (
    .dout(g1334_p),
    .din1(g1332_n),
    .din2(g1333_n)
  );


  FA
  g_g1335_n
  (
    .dout(g1335_n),
    .din1(ffc_490_p_spl_001),
    .din2(g1334_p)
  );


  LA
  g_g1336_p
  (
    .dout(g1336_p),
    .din1(ffc_486_n_spl_0011),
    .din2(g1194_n_spl_00)
  );


  LA
  g_g1337_p
  (
    .dout(g1337_p),
    .din1(ffc_486_p_spl_0011),
    .din2(g1164_n_spl_00)
  );


  FA
  g_g1338_n
  (
    .dout(g1338_n),
    .din1(ffc_490_n_spl_001),
    .din2(g1337_p)
  );


  FA
  g_g1339_n
  (
    .dout(g1339_n),
    .din1(g1336_p),
    .din2(g1338_n)
  );


  LA
  g_g1340_p
  (
    .dout(g1340_p),
    .din1(g1335_n),
    .din2(g1339_n)
  );


  FA
  g_g1341_n
  (
    .dout(g1341_n),
    .din1(ffc_96_n_spl_),
    .din2(ffc_486_p_spl_010)
  );


  FA
  g_g1342_n
  (
    .dout(g1342_n),
    .din1(ffc_92_n_spl_),
    .din2(ffc_486_n_spl_010)
  );


  LA
  g_g1343_p
  (
    .dout(g1343_p),
    .din1(g1341_n),
    .din2(g1342_n)
  );


  FA
  g_g1344_n
  (
    .dout(g1344_n),
    .din1(ffc_490_p_spl_01),
    .din2(g1343_p)
  );


  LA
  g_g1345_p
  (
    .dout(g1345_p),
    .din1(ffc_486_n_spl_010),
    .din2(g1200_p_spl_00)
  );


  LA
  g_g1346_p
  (
    .dout(g1346_p),
    .din1(ffc_486_p_spl_010),
    .din2(g1137_p_spl_00)
  );


  FA
  g_g1347_n
  (
    .dout(g1347_n),
    .din1(ffc_490_n_spl_01),
    .din2(g1346_p)
  );


  FA
  g_g1348_n
  (
    .dout(g1348_n),
    .din1(g1345_p),
    .din2(g1347_n)
  );


  LA
  g_g1349_p
  (
    .dout(g1349_p),
    .din1(g1344_n),
    .din2(g1348_n)
  );


  LA
  g_g1350_p
  (
    .dout(g1350_p),
    .din1(ffc_428_n_spl_0001),
    .din2(g1182_n_spl_0)
  );


  LA
  g_g1351_p
  (
    .dout(g1351_p),
    .din1(ffc_428_p_spl_0001),
    .din2(g1155_n_spl_0)
  );


  FA
  g_g1352_n
  (
    .dout(g1352_n),
    .din1(ffc_432_n_spl_000),
    .din2(g1351_p)
  );


  FA
  g_g1353_n
  (
    .dout(g1353_n),
    .din1(g1350_p),
    .din2(g1352_n)
  );


  LA
  g_g1354_p
  (
    .dout(g1354_p),
    .din1(ffc_289_p_spl_),
    .din2(ffc_428_n_spl_0001)
  );


  LA
  g_g1355_p
  (
    .dout(g1355_p),
    .din1(ffc_329_p_spl_),
    .din2(ffc_428_p_spl_0001)
  );


  FA
  g_g1356_n
  (
    .dout(g1356_n),
    .din1(ffc_432_p_spl_000),
    .din2(g1355_p)
  );


  FA
  g_g1357_n
  (
    .dout(g1357_n),
    .din1(g1354_p),
    .din2(g1356_n)
  );


  LA
  g_g1358_p
  (
    .dout(g1358_p),
    .din1(ffc_241_p_spl_000),
    .din2(g1357_n)
  );


  LA
  g_g1359_p
  (
    .dout(g1359_p),
    .din1(g1353_n),
    .din2(g1358_p)
  );


  FA
  g_g1360_n
  (
    .dout(g1360_n),
    .din1(ffc_428_p_spl_0010),
    .din2(g1200_p_spl_0)
  );


  FA
  g_g1361_n
  (
    .dout(g1361_n),
    .din1(ffc_428_n_spl_0010),
    .din2(g1137_p_spl_0)
  );


  LA
  g_g1362_p
  (
    .dout(g1362_p),
    .din1(ffc_432_p_spl_001),
    .din2(g1361_n)
  );


  LA
  g_g1363_p
  (
    .dout(g1363_p),
    .din1(g1360_n),
    .din2(g1362_p)
  );


  FA
  g_g1364_n
  (
    .dout(g1364_n),
    .din1(ffc_273_n_spl_),
    .din2(ffc_428_p_spl_0010)
  );


  FA
  g_g1365_n
  (
    .dout(g1365_n),
    .din1(ffc_313_n_spl_),
    .din2(ffc_428_n_spl_0010)
  );


  LA
  g_g1366_p
  (
    .dout(g1366_p),
    .din1(ffc_432_n_spl_001),
    .din2(g1365_n)
  );


  LA
  g_g1367_p
  (
    .dout(g1367_p),
    .din1(g1364_n),
    .din2(g1366_p)
  );


  FA
  g_g1368_n
  (
    .dout(g1368_n),
    .din1(ffc_241_n_spl_0),
    .din2(g1367_p)
  );


  FA
  g_g1369_n
  (
    .dout(g1369_n),
    .din1(g1363_p),
    .din2(g1368_n)
  );


  LA
  g_g1370_p
  (
    .dout(g1370_p),
    .din1(ffc_428_n_spl_0011),
    .din2(g1194_n_spl_0)
  );


  LA
  g_g1371_p
  (
    .dout(g1371_p),
    .din1(ffc_428_p_spl_0011),
    .din2(g1164_n_spl_0)
  );


  FA
  g_g1372_n
  (
    .dout(g1372_n),
    .din1(ffc_432_n_spl_001),
    .din2(g1371_p)
  );


  FA
  g_g1373_n
  (
    .dout(g1373_n),
    .din1(g1370_p),
    .din2(g1372_n)
  );


  LA
  g_g1374_p
  (
    .dout(g1374_p),
    .din1(ffc_265_p_spl_),
    .din2(ffc_428_n_spl_0011)
  );


  LA
  g_g1375_p
  (
    .dout(g1375_p),
    .din1(ffc_269_p_spl_),
    .din2(ffc_428_p_spl_0011)
  );


  FA
  g_g1376_n
  (
    .dout(g1376_n),
    .din1(ffc_432_p_spl_001),
    .din2(g1375_p)
  );


  FA
  g_g1377_n
  (
    .dout(g1377_n),
    .din1(g1374_p),
    .din2(g1376_n)
  );


  LA
  g_g1378_p
  (
    .dout(g1378_p),
    .din1(ffc_241_p_spl_001),
    .din2(g1377_n)
  );


  LA
  g_g1379_p
  (
    .dout(g1379_p),
    .din1(g1373_n),
    .din2(g1378_p)
  );


  LA
  g_g1380_p
  (
    .dout(g1380_p),
    .din1(ffc_428_n_spl_010),
    .din2(g1187_n_spl_0)
  );


  LA
  g_g1381_p
  (
    .dout(g1381_p),
    .din1(ffc_428_p_spl_010),
    .din2(g1158_n_spl_0)
  );


  FA
  g_g1382_n
  (
    .dout(g1382_n),
    .din1(ffc_432_n_spl_01),
    .din2(g1381_p)
  );


  FA
  g_g1383_n
  (
    .dout(g1383_n),
    .din1(g1380_p),
    .din2(g1382_n)
  );


  LA
  g_g1384_p
  (
    .dout(g1384_p),
    .din1(ffc_257_p_spl_),
    .din2(ffc_428_n_spl_010)
  );


  LA
  g_g1385_p
  (
    .dout(g1385_p),
    .din1(ffc_261_p_spl_),
    .din2(ffc_428_p_spl_010)
  );


  FA
  g_g1386_n
  (
    .dout(g1386_n),
    .din1(ffc_432_p_spl_01),
    .din2(g1385_p)
  );


  FA
  g_g1387_n
  (
    .dout(g1387_n),
    .din1(g1384_p),
    .din2(g1386_n)
  );


  LA
  g_g1388_p
  (
    .dout(g1388_p),
    .din1(ffc_241_p_spl_001),
    .din2(g1387_n)
  );


  LA
  g_g1389_p
  (
    .dout(g1389_p),
    .din1(g1383_n),
    .din2(g1388_p)
  );


  LA
  g_g1390_p
  (
    .dout(g1390_p),
    .din1(ffc_436_n_spl_0001),
    .din2(g1182_n_spl_1)
  );


  LA
  g_g1391_p
  (
    .dout(g1391_p),
    .din1(ffc_436_p_spl_0001),
    .din2(g1155_n_spl_1)
  );


  FA
  g_g1392_n
  (
    .dout(g1392_n),
    .din1(ffc_440_n_spl_000),
    .din2(g1391_p)
  );


  FA
  g_g1393_n
  (
    .dout(g1393_n),
    .din1(g1390_p),
    .din2(g1392_n)
  );


  LA
  g_g1394_p
  (
    .dout(g1394_p),
    .din1(ffc_289_p_spl_),
    .din2(ffc_436_n_spl_0001)
  );


  LA
  g_g1395_p
  (
    .dout(g1395_p),
    .din1(ffc_329_p_spl_),
    .din2(ffc_436_p_spl_0001)
  );


  FA
  g_g1396_n
  (
    .dout(g1396_n),
    .din1(ffc_440_p_spl_000),
    .din2(g1395_p)
  );


  FA
  g_g1397_n
  (
    .dout(g1397_n),
    .din1(g1394_p),
    .din2(g1396_n)
  );


  LA
  g_g1398_p
  (
    .dout(g1398_p),
    .din1(ffc_241_p_spl_010),
    .din2(g1397_n)
  );


  LA
  g_g1399_p
  (
    .dout(g1399_p),
    .din1(g1393_n),
    .din2(g1398_p)
  );


  FA
  g_g1400_n
  (
    .dout(g1400_n),
    .din1(ffc_436_p_spl_0010),
    .din2(g1200_p_spl_1)
  );


  FA
  g_g1401_n
  (
    .dout(g1401_n),
    .din1(ffc_436_n_spl_0010),
    .din2(g1137_p_spl_1)
  );


  LA
  g_g1402_p
  (
    .dout(g1402_p),
    .din1(ffc_440_p_spl_001),
    .din2(g1401_n)
  );


  LA
  g_g1403_p
  (
    .dout(g1403_p),
    .din1(g1400_n),
    .din2(g1402_p)
  );


  FA
  g_g1404_n
  (
    .dout(g1404_n),
    .din1(ffc_273_n_spl_),
    .din2(ffc_436_p_spl_0010)
  );


  FA
  g_g1405_n
  (
    .dout(g1405_n),
    .din1(ffc_313_n_spl_),
    .din2(ffc_436_n_spl_0010)
  );


  LA
  g_g1406_p
  (
    .dout(g1406_p),
    .din1(ffc_440_n_spl_001),
    .din2(g1405_n)
  );


  LA
  g_g1407_p
  (
    .dout(g1407_p),
    .din1(g1404_n),
    .din2(g1406_p)
  );


  FA
  g_g1408_n
  (
    .dout(g1408_n),
    .din1(ffc_241_n_spl_0),
    .din2(g1407_p)
  );


  FA
  g_g1409_n
  (
    .dout(g1409_n),
    .din1(g1403_p),
    .din2(g1408_n)
  );


  LA
  g_g1410_p
  (
    .dout(g1410_p),
    .din1(ffc_436_n_spl_0011),
    .din2(g1194_n_spl_1)
  );


  LA
  g_g1411_p
  (
    .dout(g1411_p),
    .din1(ffc_436_p_spl_0011),
    .din2(g1164_n_spl_1)
  );


  FA
  g_g1412_n
  (
    .dout(g1412_n),
    .din1(ffc_440_n_spl_001),
    .din2(g1411_p)
  );


  FA
  g_g1413_n
  (
    .dout(g1413_n),
    .din1(g1410_p),
    .din2(g1412_n)
  );


  LA
  g_g1414_p
  (
    .dout(g1414_p),
    .din1(ffc_265_p_spl_),
    .din2(ffc_436_n_spl_0011)
  );


  LA
  g_g1415_p
  (
    .dout(g1415_p),
    .din1(ffc_269_p_spl_),
    .din2(ffc_436_p_spl_0011)
  );


  FA
  g_g1416_n
  (
    .dout(g1416_n),
    .din1(ffc_440_p_spl_001),
    .din2(g1415_p)
  );


  FA
  g_g1417_n
  (
    .dout(g1417_n),
    .din1(g1414_p),
    .din2(g1416_n)
  );


  LA
  g_g1418_p
  (
    .dout(g1418_p),
    .din1(ffc_241_p_spl_010),
    .din2(g1417_n)
  );


  LA
  g_g1419_p
  (
    .dout(g1419_p),
    .din1(g1413_n),
    .din2(g1418_p)
  );


  LA
  g_g1420_p
  (
    .dout(g1420_p),
    .din1(ffc_257_p_spl_),
    .din2(ffc_436_n_spl_010)
  );


  LA
  g_g1421_p
  (
    .dout(g1421_p),
    .din1(ffc_261_p_spl_),
    .din2(ffc_436_p_spl_010)
  );


  FA
  g_g1422_n
  (
    .dout(g1422_n),
    .din1(g1420_p),
    .din2(g1421_p)
  );


  LA
  g_g1423_p
  (
    .dout(g1423_p),
    .din1(ffc_440_n_spl_01),
    .din2(g1422_n)
  );


  FA
  g_g1424_n
  (
    .dout(g1424_n),
    .din1(ffc_436_p_spl_010),
    .din2(g1187_n_spl_1)
  );


  FA
  g_g1425_n
  (
    .dout(g1425_n),
    .din1(ffc_436_n_spl_010),
    .din2(g1158_n_spl_1)
  );


  LA
  g_g1426_p
  (
    .dout(g1426_p),
    .din1(ffc_440_p_spl_01),
    .din2(g1425_n)
  );


  LA
  g_g1427_p
  (
    .dout(g1427_p),
    .din1(g1424_n),
    .din2(g1426_p)
  );


  FA
  g_g1428_n
  (
    .dout(g1428_n),
    .din1(g1423_p),
    .din2(g1427_p)
  );


  LA
  g_g1429_p
  (
    .dout(g1429_p),
    .din1(ffc_241_p_spl_011),
    .din2(g1428_n)
  );


  FA
  g_g1430_n
  (
    .dout(g1430_n),
    .din1(ffc_233_n),
    .din2(ffc_502_n)
  );


  LA
  g_g1431_p
  (
    .dout(g1431_p),
    .din1(ffc_205_p),
    .din2(ffc_474_n_spl_)
  );


  LA
  g_g1432_p
  (
    .dout(g1432_p),
    .din1(ffc_474_p_spl_),
    .din2(ffc_561_n_spl_0)
  );


  FA
  g_g1433_n
  (
    .dout(g1433_n),
    .din1(g1431_p),
    .din2(g1432_p)
  );


  LA
  g_g1434_p
  (
    .dout(g1434_p),
    .din1(ffc_470_p),
    .din2(g1433_n)
  );


  LA
  g_g1435_p
  (
    .dout(g1435_p),
    .din1(ffc_229_n_spl_),
    .din2(ffc_532_p_spl_0)
  );


  FA
  g_g1435_n
  (
    .dout(g1435_n),
    .din1(ffc_229_p_spl_),
    .din2(ffc_532_n_spl_)
  );


  LA
  g_g1436_p
  (
    .dout(g1436_p),
    .din1(ffc_229_p_spl_),
    .din2(ffc_532_n_spl_)
  );


  FA
  g_g1436_n
  (
    .dout(g1436_n),
    .din1(ffc_229_n_spl_),
    .din2(ffc_532_p_spl_)
  );


  LA
  g_g1437_p
  (
    .dout(g1437_p),
    .din1(g1435_n),
    .din2(g1436_n)
  );


  FA
  g_g1437_n
  (
    .dout(g1437_n),
    .din1(g1435_p),
    .din2(g1436_p)
  );


  LA
  g_g1438_p
  (
    .dout(g1438_p),
    .din1(ffc_474_p_spl_),
    .din2(g1437_n_spl_)
  );


  LA
  g_g1439_p
  (
    .dout(g1439_p),
    .din1(ffc_474_n_spl_),
    .din2(ffc_524_p)
  );


  FA
  g_g1440_n
  (
    .dout(g1440_n),
    .din1(g1438_p),
    .din2(g1439_p)
  );


  LA
  g_g1441_p
  (
    .dout(g1441_p),
    .din1(ffc_470_n),
    .din2(g1440_n)
  );


  FA
  g_g1442_n
  (
    .dout(g1442_n),
    .din1(g1434_p),
    .din2(g1441_p)
  );


  LA
  g_g1443_p
  (
    .dout(g1443_p),
    .din1(g1430_n),
    .din2(g1442_n)
  );


  FA
  g_g1444_n
  (
    .dout(g1444_n),
    .din1(ffc_561_p_spl_1),
    .din2(g1437_p)
  );


  FA
  g_g1445_n
  (
    .dout(g1445_n),
    .din1(ffc_561_n_spl_1),
    .din2(g1437_n_spl_)
  );


  LA
  g_g1446_p
  (
    .dout(g1446_p),
    .din1(g1444_n),
    .din2(g1445_n)
  );


  LA
  g_g1447_p
  (
    .dout(g1447_p),
    .din1(ffc_561_n_spl_1),
    .din2(ffc_697_p_spl_100)
  );


  LA
  g_g1448_p
  (
    .dout(g1448_p),
    .din1(ffc_698_p),
    .din2(ffc_702_n)
  );


  FA
  g_g1449_n
  (
    .dout(g1449_n),
    .din1(g1447_p),
    .din2(g1448_p)
  );


  LA
  g_g1450_p
  (
    .dout(g1450_p),
    .din1(ffc_697_p_spl_100),
    .din2(g1249_p_spl_)
  );


  FA
  g_g1451_n
  (
    .dout(g1451_n),
    .din1(ffc_691_p),
    .din2(ffc_703_p)
  );


  LA
  g_g1452_p
  (
    .dout(g1452_p),
    .din1(ffc_494_p_spl_100),
    .din2(g1451_n)
  );


  FA
  g_g1453_n
  (
    .dout(g1453_n),
    .din1(g1450_p),
    .din2(g1452_p)
  );


  LA
  g_g1454_p
  (
    .dout(g1454_p),
    .din1(ffc_697_p_spl_101),
    .din2(g1250_p_spl_)
  );


  FA
  g_g1455_n
  (
    .dout(g1455_n),
    .din1(ffc_688_p),
    .din2(ffc_704_p)
  );


  LA
  g_g1456_p
  (
    .dout(g1456_p),
    .din1(ffc_494_p_spl_100),
    .din2(g1455_n)
  );


  FA
  g_g1457_n
  (
    .dout(g1457_n),
    .din1(g1454_p),
    .din2(g1456_p)
  );


  LA
  g_g1458_p
  (
    .dout(g1458_p),
    .din1(ffc_697_p_spl_101),
    .din2(ffc_746_p_spl_)
  );


  LA
  g_g1459_p
  (
    .dout(g1459_p),
    .din1(ffc_494_p_spl_101),
    .din2(ffc_725_p)
  );


  FA
  g_g1460_n
  (
    .dout(g1460_n),
    .din1(g1458_p),
    .din2(g1459_p)
  );


  FA
  g_g1461_n
  (
    .dout(g1461_n),
    .din1(ffc_342_n_spl_),
    .din2(ffc_417_n_spl_)
  );


  FA
  g_g1462_n
  (
    .dout(g1462_n),
    .din1(g1049_n_spl_),
    .din2(g1461_n)
  );


  FA
  g_g1463_n
  (
    .dout(g1463_n),
    .din1(g1054_n_spl_),
    .din2(g1462_n)
  );


  FA
  g_g1464_n
  (
    .dout(g1464_n),
    .din1(g1111_n_spl_),
    .din2(g1463_n)
  );


  FA
  g_g1465_n
  (
    .dout(g1465_n),
    .din1(g1120_n_spl_),
    .din2(g1464_n)
  );


  FA
  g_g1466_n
  (
    .dout(g1466_n),
    .din1(g1212_n_spl_),
    .din2(g1465_n)
  );


  FA
  g_g1467_n
  (
    .dout(g1467_n),
    .din1(g1233_n_spl_),
    .din2(g1466_n)
  );


  LA
  g_g1468_p
  (
    .dout(g1468_p),
    .din1(ffc_697_p_spl_110),
    .din2(ffc_745_n_spl_)
  );


  LA
  g_g1469_p
  (
    .dout(g1469_p),
    .din1(ffc_494_p_spl_101),
    .din2(ffc_726_p)
  );


  FA
  g_g1470_n
  (
    .dout(g1470_n),
    .din1(g1468_p),
    .din2(g1469_p)
  );


  LA
  g_g1471_p
  (
    .dout(g1471_p),
    .din1(ffc_697_p_spl_110),
    .din2(g1243_p_spl_)
  );


  LA
  g_g1472_p
  (
    .dout(g1472_p),
    .din1(ffc_174_p),
    .din2(ffc_498_n_spl_10)
  );


  LA
  g_g1473_p
  (
    .dout(g1473_p),
    .din1(ffc_498_p_spl_01),
    .din2(ffc_734_n)
  );


  FA
  g_g1474_n
  (
    .dout(g1474_n),
    .din1(g1472_p),
    .din2(g1473_p)
  );


  LA
  g_g1475_p
  (
    .dout(g1475_p),
    .din1(ffc_494_p_spl_110),
    .din2(g1474_n)
  );


  FA
  g_g1476_n
  (
    .dout(g1476_n),
    .din1(g1471_p),
    .din2(g1475_p)
  );


  LA
  g_g1477_p
  (
    .dout(g1477_p),
    .din1(ffc_697_p_spl_111),
    .din2(g1246_p_spl_)
  );


  LA
  g_g1478_p
  (
    .dout(g1478_p),
    .din1(ffc_77_p),
    .din2(ffc_498_n_spl_11)
  );


  LA
  g_g1479_p
  (
    .dout(g1479_p),
    .din1(ffc_498_p_spl_10),
    .din2(ffc_735_n)
  );


  FA
  g_g1480_n
  (
    .dout(g1480_n),
    .din1(g1478_p),
    .din2(g1479_p)
  );


  LA
  g_g1481_p
  (
    .dout(g1481_p),
    .din1(ffc_494_p_spl_110),
    .din2(g1480_n)
  );


  FA
  g_g1482_n
  (
    .dout(g1482_n),
    .din1(g1477_p),
    .din2(g1481_p)
  );


  LA
  g_g1483_p
  (
    .dout(g1483_p),
    .din1(ffc_697_p_spl_111),
    .din2(g1234_n_spl_)
  );


  FA
  g_g1484_n
  (
    .dout(g1484_n),
    .din1(ffc_687_p),
    .din2(ffc_705_p)
  );


  LA
  g_g1485_p
  (
    .dout(g1485_p),
    .din1(ffc_494_p_spl_11),
    .din2(g1484_n)
  );


  FA
  g_g1486_n
  (
    .dout(g1486_n),
    .din1(g1483_p),
    .din2(g1485_p)
  );


  LA
  g_g1487_p
  (
    .dout(g1487_p),
    .din1(ffc_160_p_spl_),
    .din2(ffc_486_n_spl_011)
  );


  LA
  g_g1488_p
  (
    .dout(g1488_p),
    .din1(ffc_164_p_spl_),
    .din2(ffc_486_p_spl_011)
  );


  FA
  g_g1489_n
  (
    .dout(g1489_n),
    .din1(g1487_p),
    .din2(g1488_p)
  );


  LA
  g_g1490_p
  (
    .dout(g1490_p),
    .din1(ffc_490_n_spl_01),
    .din2(g1489_n)
  );


  LA
  g_g1491_p
  (
    .dout(g1491_p),
    .din1(ffc_486_n_spl_011),
    .din2(g1470_n_spl_00)
  );


  LA
  g_g1492_p
  (
    .dout(g1492_p),
    .din1(ffc_486_p_spl_011),
    .din2(g1449_n_spl_00)
  );


  FA
  g_g1493_n
  (
    .dout(g1493_n),
    .din1(g1491_p),
    .din2(g1492_p)
  );


  LA
  g_g1494_p
  (
    .dout(g1494_p),
    .din1(ffc_490_p_spl_01),
    .din2(g1493_n)
  );


  FA
  g_g1495_n
  (
    .dout(g1495_n),
    .din1(g1490_p),
    .din2(g1494_p)
  );


  LA
  g_g1496_p
  (
    .dout(g1496_p),
    .din1(ffc_482_n_spl_011),
    .din2(g1470_n_spl_00)
  );


  LA
  g_g1497_p
  (
    .dout(g1497_p),
    .din1(ffc_482_p_spl_011),
    .din2(g1449_n_spl_00)
  );


  FA
  g_g1498_n
  (
    .dout(g1498_n),
    .din1(ffc_478_n_spl_01),
    .din2(g1497_p)
  );


  FA
  g_g1499_n
  (
    .dout(g1499_n),
    .din1(g1496_p),
    .din2(g1498_n)
  );


  FA
  g_g1500_n
  (
    .dout(g1500_n),
    .din1(ffc_160_p_spl_),
    .din2(ffc_482_p_spl_011)
  );


  FA
  g_g1501_n
  (
    .dout(g1501_n),
    .din1(ffc_164_p_spl_),
    .din2(ffc_482_n_spl_011)
  );


  LA
  g_g1502_p
  (
    .dout(g1502_p),
    .din1(g1500_n),
    .din2(g1501_n)
  );


  FA
  g_g1503_n
  (
    .dout(g1503_n),
    .din1(ffc_478_p_spl_01),
    .din2(g1502_p)
  );


  LA
  g_g1504_p
  (
    .dout(g1504_p),
    .din1(g1499_n),
    .din2(g1503_n)
  );


  FA
  g_g1505_n
  (
    .dout(g1505_n),
    .din1(ffc_70_p_spl_),
    .din2(ffc_482_p_spl_100)
  );


  FA
  g_g1506_n
  (
    .dout(g1506_n),
    .din1(ffc_66_p_spl_),
    .din2(ffc_482_n_spl_100)
  );


  LA
  g_g1507_p
  (
    .dout(g1507_p),
    .din1(g1505_n),
    .din2(g1506_n)
  );


  FA
  g_g1508_n
  (
    .dout(g1508_n),
    .din1(ffc_478_p_spl_10),
    .din2(g1507_p)
  );


  LA
  g_g1509_p
  (
    .dout(g1509_p),
    .din1(ffc_482_n_spl_100),
    .din2(g1476_n_spl_00)
  );


  LA
  g_g1510_p
  (
    .dout(g1510_p),
    .din1(ffc_482_p_spl_100),
    .din2(g1453_n_spl_00)
  );


  FA
  g_g1511_n
  (
    .dout(g1511_n),
    .din1(ffc_478_n_spl_10),
    .din2(g1510_p)
  );


  FA
  g_g1512_n
  (
    .dout(g1512_n),
    .din1(g1509_p),
    .din2(g1511_n)
  );


  LA
  g_g1513_p
  (
    .dout(g1513_p),
    .din1(g1508_n),
    .din2(g1512_n)
  );


  FA
  g_g1514_n
  (
    .dout(g1514_n),
    .din1(ffc_156_p_spl_),
    .din2(ffc_482_p_spl_101)
  );


  FA
  g_g1515_n
  (
    .dout(g1515_n),
    .din1(ffc_152_p_spl_),
    .din2(ffc_482_n_spl_101)
  );


  LA
  g_g1516_p
  (
    .dout(g1516_p),
    .din1(g1514_n),
    .din2(g1515_n)
  );


  FA
  g_g1517_n
  (
    .dout(g1517_n),
    .din1(ffc_478_p_spl_10),
    .din2(g1516_p)
  );


  LA
  g_g1518_p
  (
    .dout(g1518_p),
    .din1(ffc_482_n_spl_101),
    .din2(g1482_n_spl_00)
  );


  LA
  g_g1519_p
  (
    .dout(g1519_p),
    .din1(ffc_482_p_spl_101),
    .din2(g1457_n_spl_00)
  );


  FA
  g_g1520_n
  (
    .dout(g1520_n),
    .din1(ffc_478_n_spl_10),
    .din2(g1519_p)
  );


  FA
  g_g1521_n
  (
    .dout(g1521_n),
    .din1(g1518_p),
    .din2(g1520_n)
  );


  LA
  g_g1522_p
  (
    .dout(g1522_p),
    .din1(g1517_n),
    .din2(g1521_n)
  );


  FA
  g_g1523_n
  (
    .dout(g1523_n),
    .din1(ffc_58_p_spl_),
    .din2(ffc_482_p_spl_110)
  );


  FA
  g_g1524_n
  (
    .dout(g1524_n),
    .din1(ffc_140_p_spl_),
    .din2(ffc_482_n_spl_110)
  );


  LA
  g_g1525_p
  (
    .dout(g1525_p),
    .din1(g1523_n),
    .din2(g1524_n)
  );


  FA
  g_g1526_n
  (
    .dout(g1526_n),
    .din1(ffc_478_p_spl_11),
    .din2(g1525_p)
  );


  LA
  g_g1527_p
  (
    .dout(g1527_p),
    .din1(ffc_482_n_spl_110),
    .din2(g1486_n_spl_00)
  );


  LA
  g_g1528_p
  (
    .dout(g1528_p),
    .din1(ffc_482_p_spl_110),
    .din2(g1460_n_spl_00)
  );


  FA
  g_g1529_n
  (
    .dout(g1529_n),
    .din1(ffc_478_n_spl_11),
    .din2(g1528_p)
  );


  FA
  g_g1530_n
  (
    .dout(g1530_n),
    .din1(g1527_p),
    .din2(g1529_n)
  );


  LA
  g_g1531_p
  (
    .dout(g1531_p),
    .din1(g1526_n),
    .din2(g1530_n)
  );


  FA
  g_g1532_n
  (
    .dout(g1532_n),
    .din1(ffc_70_p_spl_),
    .din2(ffc_486_p_spl_100)
  );


  FA
  g_g1533_n
  (
    .dout(g1533_n),
    .din1(ffc_66_p_spl_),
    .din2(ffc_486_n_spl_100)
  );


  LA
  g_g1534_p
  (
    .dout(g1534_p),
    .din1(g1532_n),
    .din2(g1533_n)
  );


  FA
  g_g1535_n
  (
    .dout(g1535_n),
    .din1(ffc_490_p_spl_10),
    .din2(g1534_p)
  );


  LA
  g_g1536_p
  (
    .dout(g1536_p),
    .din1(ffc_486_n_spl_100),
    .din2(g1476_n_spl_00)
  );


  LA
  g_g1537_p
  (
    .dout(g1537_p),
    .din1(ffc_486_p_spl_100),
    .din2(g1453_n_spl_00)
  );


  FA
  g_g1538_n
  (
    .dout(g1538_n),
    .din1(ffc_490_n_spl_10),
    .din2(g1537_p)
  );


  FA
  g_g1539_n
  (
    .dout(g1539_n),
    .din1(g1536_p),
    .din2(g1538_n)
  );


  LA
  g_g1540_p
  (
    .dout(g1540_p),
    .din1(g1535_n),
    .din2(g1539_n)
  );


  FA
  g_g1541_n
  (
    .dout(g1541_n),
    .din1(ffc_156_p_spl_),
    .din2(ffc_486_p_spl_101)
  );


  FA
  g_g1542_n
  (
    .dout(g1542_n),
    .din1(ffc_152_p_spl_),
    .din2(ffc_486_n_spl_101)
  );


  LA
  g_g1543_p
  (
    .dout(g1543_p),
    .din1(g1541_n),
    .din2(g1542_n)
  );


  FA
  g_g1544_n
  (
    .dout(g1544_n),
    .din1(ffc_490_p_spl_10),
    .din2(g1543_p)
  );


  LA
  g_g1545_p
  (
    .dout(g1545_p),
    .din1(ffc_486_n_spl_101),
    .din2(g1482_n_spl_00)
  );


  LA
  g_g1546_p
  (
    .dout(g1546_p),
    .din1(ffc_486_p_spl_101),
    .din2(g1457_n_spl_00)
  );


  FA
  g_g1547_n
  (
    .dout(g1547_n),
    .din1(ffc_490_n_spl_10),
    .din2(g1546_p)
  );


  FA
  g_g1548_n
  (
    .dout(g1548_n),
    .din1(g1545_p),
    .din2(g1547_n)
  );


  LA
  g_g1549_p
  (
    .dout(g1549_p),
    .din1(g1544_n),
    .din2(g1548_n)
  );


  FA
  g_g1550_n
  (
    .dout(g1550_n),
    .din1(ffc_58_p_spl_),
    .din2(ffc_486_p_spl_110)
  );


  FA
  g_g1551_n
  (
    .dout(g1551_n),
    .din1(ffc_140_p_spl_),
    .din2(ffc_486_n_spl_110)
  );


  LA
  g_g1552_p
  (
    .dout(g1552_p),
    .din1(g1550_n),
    .din2(g1551_n)
  );


  FA
  g_g1553_n
  (
    .dout(g1553_n),
    .din1(ffc_490_p_spl_11),
    .din2(g1552_p)
  );


  LA
  g_g1554_p
  (
    .dout(g1554_p),
    .din1(ffc_486_n_spl_110),
    .din2(g1486_n_spl_00)
  );


  LA
  g_g1555_p
  (
    .dout(g1555_p),
    .din1(ffc_486_p_spl_110),
    .din2(g1460_n_spl_00)
  );


  FA
  g_g1556_n
  (
    .dout(g1556_n),
    .din1(ffc_490_n_spl_11),
    .din2(g1555_p)
  );


  FA
  g_g1557_n
  (
    .dout(g1557_n),
    .din1(g1554_p),
    .din2(g1556_n)
  );


  LA
  g_g1558_p
  (
    .dout(g1558_p),
    .din1(g1553_n),
    .din2(g1557_n)
  );


  LA
  g_g1559_p
  (
    .dout(g1559_p),
    .din1(ffc_428_n_spl_011),
    .din2(g1486_n_spl_0)
  );


  LA
  g_g1560_p
  (
    .dout(g1560_p),
    .din1(ffc_428_p_spl_011),
    .din2(g1460_n_spl_0)
  );


  FA
  g_g1561_n
  (
    .dout(g1561_n),
    .din1(ffc_432_n_spl_01),
    .din2(g1560_p)
  );


  FA
  g_g1562_n
  (
    .dout(g1562_n),
    .din1(g1559_p),
    .din2(g1561_n)
  );


  LA
  g_g1563_p
  (
    .dout(g1563_p),
    .din1(ffc_293_p_spl_),
    .din2(ffc_428_n_spl_011)
  );


  LA
  g_g1564_p
  (
    .dout(g1564_p),
    .din1(ffc_333_p_spl_),
    .din2(ffc_428_p_spl_011)
  );


  FA
  g_g1565_n
  (
    .dout(g1565_n),
    .din1(ffc_432_p_spl_01),
    .din2(g1564_p)
  );


  FA
  g_g1566_n
  (
    .dout(g1566_n),
    .din1(g1563_p),
    .din2(g1565_n)
  );


  LA
  g_g1567_p
  (
    .dout(g1567_p),
    .din1(ffc_241_p_spl_011),
    .din2(g1566_n)
  );


  LA
  g_g1568_p
  (
    .dout(g1568_p),
    .din1(g1562_n),
    .din2(g1567_p)
  );


  LA
  g_g1569_p
  (
    .dout(g1569_p),
    .din1(ffc_428_n_spl_100),
    .din2(g1482_n_spl_0)
  );


  LA
  g_g1570_p
  (
    .dout(g1570_p),
    .din1(ffc_428_p_spl_100),
    .din2(g1457_n_spl_0)
  );


  FA
  g_g1571_n
  (
    .dout(g1571_n),
    .din1(ffc_432_n_spl_10),
    .din2(g1570_p)
  );


  FA
  g_g1572_n
  (
    .dout(g1572_n),
    .din1(g1569_p),
    .din2(g1571_n)
  );


  LA
  g_g1573_p
  (
    .dout(g1573_p),
    .din1(ffc_285_p_spl_),
    .din2(ffc_428_n_spl_100)
  );


  LA
  g_g1574_p
  (
    .dout(g1574_p),
    .din1(ffc_325_p_spl_),
    .din2(ffc_428_p_spl_100)
  );


  FA
  g_g1575_n
  (
    .dout(g1575_n),
    .din1(ffc_432_p_spl_10),
    .din2(g1574_p)
  );


  FA
  g_g1576_n
  (
    .dout(g1576_n),
    .din1(g1573_p),
    .din2(g1575_n)
  );


  LA
  g_g1577_p
  (
    .dout(g1577_p),
    .din1(ffc_241_p_spl_100),
    .din2(g1576_n)
  );


  LA
  g_g1578_p
  (
    .dout(g1578_p),
    .din1(g1572_n),
    .din2(g1577_p)
  );


  LA
  g_g1579_p
  (
    .dout(g1579_p),
    .din1(ffc_428_n_spl_101),
    .din2(g1476_n_spl_0)
  );


  LA
  g_g1580_p
  (
    .dout(g1580_p),
    .din1(ffc_428_p_spl_101),
    .din2(g1453_n_spl_0)
  );


  FA
  g_g1581_n
  (
    .dout(g1581_n),
    .din1(ffc_432_n_spl_10),
    .din2(g1580_p)
  );


  FA
  g_g1582_n
  (
    .dout(g1582_n),
    .din1(g1579_p),
    .din2(g1581_n)
  );


  LA
  g_g1583_p
  (
    .dout(g1583_p),
    .din1(ffc_281_p_spl_),
    .din2(ffc_428_n_spl_101)
  );


  LA
  g_g1584_p
  (
    .dout(g1584_p),
    .din1(ffc_321_p_spl_),
    .din2(ffc_428_p_spl_101)
  );


  FA
  g_g1585_n
  (
    .dout(g1585_n),
    .din1(ffc_432_p_spl_10),
    .din2(g1584_p)
  );


  FA
  g_g1586_n
  (
    .dout(g1586_n),
    .din1(g1583_p),
    .din2(g1585_n)
  );


  LA
  g_g1587_p
  (
    .dout(g1587_p),
    .din1(ffc_241_p_spl_100),
    .din2(g1586_n)
  );


  LA
  g_g1588_p
  (
    .dout(g1588_p),
    .din1(g1582_n),
    .din2(g1587_p)
  );


  LA
  g_g1589_p
  (
    .dout(g1589_p),
    .din1(ffc_277_p_spl_),
    .din2(ffc_428_n_spl_110)
  );


  LA
  g_g1590_p
  (
    .dout(g1590_p),
    .din1(ffc_317_p_spl_),
    .din2(ffc_428_p_spl_110)
  );


  FA
  g_g1591_n
  (
    .dout(g1591_n),
    .din1(g1589_p),
    .din2(g1590_p)
  );


  LA
  g_g1592_p
  (
    .dout(g1592_p),
    .din1(ffc_432_n_spl_11),
    .din2(g1591_n)
  );


  LA
  g_g1593_p
  (
    .dout(g1593_p),
    .din1(ffc_428_n_spl_110),
    .din2(g1470_n_spl_0)
  );


  LA
  g_g1594_p
  (
    .dout(g1594_p),
    .din1(ffc_428_p_spl_110),
    .din2(g1449_n_spl_0)
  );


  FA
  g_g1595_n
  (
    .dout(g1595_n),
    .din1(g1593_p),
    .din2(g1594_p)
  );


  LA
  g_g1596_p
  (
    .dout(g1596_p),
    .din1(ffc_432_p_spl_11),
    .din2(g1595_n)
  );


  FA
  g_g1597_n
  (
    .dout(g1597_n),
    .din1(g1592_p),
    .din2(g1596_p)
  );


  LA
  g_g1598_p
  (
    .dout(g1598_p),
    .din1(ffc_241_p_spl_101),
    .din2(g1597_n)
  );


  LA
  g_g1599_p
  (
    .dout(g1599_p),
    .din1(ffc_293_p_spl_),
    .din2(ffc_436_n_spl_011)
  );


  LA
  g_g1600_p
  (
    .dout(g1600_p),
    .din1(ffc_333_p_spl_),
    .din2(ffc_436_p_spl_011)
  );


  FA
  g_g1601_n
  (
    .dout(g1601_n),
    .din1(g1599_p),
    .din2(g1600_p)
  );


  LA
  g_g1602_p
  (
    .dout(g1602_p),
    .din1(ffc_440_n_spl_01),
    .din2(g1601_n)
  );


  FA
  g_g1603_n
  (
    .dout(g1603_n),
    .din1(ffc_436_p_spl_011),
    .din2(g1486_n_spl_1)
  );


  FA
  g_g1604_n
  (
    .dout(g1604_n),
    .din1(ffc_436_n_spl_011),
    .din2(g1460_n_spl_1)
  );


  LA
  g_g1605_p
  (
    .dout(g1605_p),
    .din1(ffc_440_p_spl_01),
    .din2(g1604_n)
  );


  LA
  g_g1606_p
  (
    .dout(g1606_p),
    .din1(g1603_n),
    .din2(g1605_p)
  );


  FA
  g_g1607_n
  (
    .dout(g1607_n),
    .din1(g1602_p),
    .din2(g1606_p)
  );


  LA
  g_g1608_p
  (
    .dout(g1608_p),
    .din1(ffc_241_p_spl_101),
    .din2(g1607_n)
  );


  LA
  g_g1609_p
  (
    .dout(g1609_p),
    .din1(ffc_436_n_spl_100),
    .din2(g1482_n_spl_1)
  );


  LA
  g_g1610_p
  (
    .dout(g1610_p),
    .din1(ffc_436_p_spl_100),
    .din2(g1457_n_spl_1)
  );


  FA
  g_g1611_n
  (
    .dout(g1611_n),
    .din1(ffc_440_n_spl_10),
    .din2(g1610_p)
  );


  FA
  g_g1612_n
  (
    .dout(g1612_n),
    .din1(g1609_p),
    .din2(g1611_n)
  );


  LA
  g_g1613_p
  (
    .dout(g1613_p),
    .din1(ffc_285_p_spl_),
    .din2(ffc_436_n_spl_100)
  );


  LA
  g_g1614_p
  (
    .dout(g1614_p),
    .din1(ffc_325_p_spl_),
    .din2(ffc_436_p_spl_100)
  );


  FA
  g_g1615_n
  (
    .dout(g1615_n),
    .din1(ffc_440_p_spl_10),
    .din2(g1614_p)
  );


  FA
  g_g1616_n
  (
    .dout(g1616_n),
    .din1(g1613_p),
    .din2(g1615_n)
  );


  LA
  g_g1617_p
  (
    .dout(g1617_p),
    .din1(ffc_241_p_spl_110),
    .din2(g1616_n)
  );


  LA
  g_g1618_p
  (
    .dout(g1618_p),
    .din1(g1612_n),
    .din2(g1617_p)
  );


  LA
  g_g1619_p
  (
    .dout(g1619_p),
    .din1(ffc_436_n_spl_101),
    .din2(g1476_n_spl_1)
  );


  LA
  g_g1620_p
  (
    .dout(g1620_p),
    .din1(ffc_436_p_spl_101),
    .din2(g1453_n_spl_1)
  );


  FA
  g_g1621_n
  (
    .dout(g1621_n),
    .din1(ffc_440_n_spl_10),
    .din2(g1620_p)
  );


  FA
  g_g1622_n
  (
    .dout(g1622_n),
    .din1(g1619_p),
    .din2(g1621_n)
  );


  LA
  g_g1623_p
  (
    .dout(g1623_p),
    .din1(ffc_281_p_spl_),
    .din2(ffc_436_n_spl_101)
  );


  LA
  g_g1624_p
  (
    .dout(g1624_p),
    .din1(ffc_321_p_spl_),
    .din2(ffc_436_p_spl_101)
  );


  FA
  g_g1625_n
  (
    .dout(g1625_n),
    .din1(ffc_440_p_spl_10),
    .din2(g1624_p)
  );


  FA
  g_g1626_n
  (
    .dout(g1626_n),
    .din1(g1623_p),
    .din2(g1625_n)
  );


  LA
  g_g1627_p
  (
    .dout(g1627_p),
    .din1(ffc_241_p_spl_110),
    .din2(g1626_n)
  );


  LA
  g_g1628_p
  (
    .dout(g1628_p),
    .din1(g1622_n),
    .din2(g1627_p)
  );


  LA
  g_g1629_p
  (
    .dout(g1629_p),
    .din1(ffc_436_n_spl_110),
    .din2(g1470_n_spl_1)
  );


  LA
  g_g1630_p
  (
    .dout(g1630_p),
    .din1(ffc_436_p_spl_110),
    .din2(g1449_n_spl_1)
  );


  FA
  g_g1631_n
  (
    .dout(g1631_n),
    .din1(ffc_440_n_spl_11),
    .din2(g1630_p)
  );


  FA
  g_g1632_n
  (
    .dout(g1632_n),
    .din1(g1629_p),
    .din2(g1631_n)
  );


  LA
  g_g1633_p
  (
    .dout(g1633_p),
    .din1(ffc_277_p_spl_),
    .din2(ffc_436_n_spl_110)
  );


  LA
  g_g1634_p
  (
    .dout(g1634_p),
    .din1(ffc_317_p_spl_),
    .din2(ffc_436_p_spl_110)
  );


  FA
  g_g1635_n
  (
    .dout(g1635_n),
    .din1(ffc_440_p_spl_11),
    .din2(g1634_p)
  );


  FA
  g_g1636_n
  (
    .dout(g1636_n),
    .din1(g1633_p),
    .din2(g1635_n)
  );


  LA
  g_g1637_p
  (
    .dout(g1637_p),
    .din1(ffc_241_p_spl_111),
    .din2(g1636_n)
  );


  LA
  g_g1638_p
  (
    .dout(g1638_p),
    .din1(g1632_n),
    .din2(g1637_p)
  );


  FA
  g_g1639_n
  (
    .dout(g1639_n),
    .din1(ffc_699_p),
    .din2(ffc_706_n)
  );


  FA
  g_g1640_n
  (
    .dout(g1640_n),
    .din1(ffc_494_n_spl_1),
    .din2(ffc_498_p_spl_10)
  );


  FA
  g_g1641_n
  (
    .dout(g1641_n),
    .din1(ffc_194_p),
    .din2(g1640_n_spl_)
  );


  LA
  g_g1642_p
  (
    .dout(g1642_p),
    .din1(g1639_n_spl_),
    .din2(g1641_n)
  );


  LA
  g_g1643_p
  (
    .dout(g1643_p),
    .din1(ffc_494_n_spl_1),
    .din2(ffc_754_n)
  );


  FA
  g_g1644_n
  (
    .dout(g1644_n),
    .din1(ffc_498_n_spl_11),
    .din2(ffc_738_p)
  );


  FA
  g_g1645_n
  (
    .dout(g1645_n),
    .din1(g1643_p),
    .din2(g1644_n)
  );


  FA
  g_g1646_n
  (
    .dout(g1646_n),
    .din1(ffc_187_p),
    .din2(g1640_n_spl_)
  );


  LA
  g_g1647_p
  (
    .dout(g1647_p),
    .din1(g1645_n_spl_),
    .din2(g1646_n)
  );


  LA
  g_g1648_p
  (
    .dout(g1648_p),
    .din1(ffc_88_n_spl_),
    .din2(ffc_482_n_spl_111)
  );


  LA
  g_g1649_p
  (
    .dout(g1649_p),
    .din1(ffc_14_n_spl_),
    .din2(ffc_482_p_spl_111)
  );


  FA
  g_g1650_n
  (
    .dout(g1650_n),
    .din1(g1648_p),
    .din2(g1649_p)
  );


  LA
  g_g1651_p
  (
    .dout(g1651_p),
    .din1(ffc_478_n_spl_11),
    .din2(g1650_n)
  );


  FA
  g_g1652_n
  (
    .dout(g1652_n),
    .din1(ffc_148_n),
    .din2(ffc_498_p_spl_11)
  );


  LA
  g_g1653_p
  (
    .dout(g1653_p),
    .din1(g1645_n_spl_),
    .din2(g1652_n)
  );


  FA
  g_g1654_n
  (
    .dout(g1654_n),
    .din1(ffc_482_p_spl_111),
    .din2(g1653_p_spl_0)
  );


  FA
  g_g1655_n
  (
    .dout(g1655_n),
    .din1(ffc_144_n),
    .din2(ffc_498_p_spl_11)
  );


  LA
  g_g1656_p
  (
    .dout(g1656_p),
    .din1(g1639_n_spl_),
    .din2(g1655_n)
  );


  FA
  g_g1657_n
  (
    .dout(g1657_n),
    .din1(ffc_482_n_spl_111),
    .din2(g1656_p_spl_0)
  );


  LA
  g_g1658_p
  (
    .dout(g1658_p),
    .din1(ffc_478_p_spl_11),
    .din2(g1657_n)
  );


  LA
  g_g1659_p
  (
    .dout(g1659_p),
    .din1(g1654_n),
    .din2(g1658_p)
  );


  FA
  g_g1660_n
  (
    .dout(g1660_n),
    .din1(g1651_p),
    .din2(g1659_p)
  );


  LA
  g_g1661_p
  (
    .dout(g1661_p),
    .din1(ffc_88_n_spl_),
    .din2(ffc_486_n_spl_111)
  );


  LA
  g_g1662_p
  (
    .dout(g1662_p),
    .din1(ffc_14_n_spl_),
    .din2(ffc_486_p_spl_111)
  );


  FA
  g_g1663_n
  (
    .dout(g1663_n),
    .din1(g1661_p),
    .din2(g1662_p)
  );


  LA
  g_g1664_p
  (
    .dout(g1664_p),
    .din1(ffc_490_n_spl_11),
    .din2(g1663_n)
  );


  FA
  g_g1665_n
  (
    .dout(g1665_n),
    .din1(ffc_486_p_spl_111),
    .din2(g1653_p_spl_0)
  );


  FA
  g_g1666_n
  (
    .dout(g1666_n),
    .din1(ffc_486_n_spl_111),
    .din2(g1656_p_spl_0)
  );


  LA
  g_g1667_p
  (
    .dout(g1667_p),
    .din1(ffc_490_p_spl_11),
    .din2(g1666_n)
  );


  LA
  g_g1668_p
  (
    .dout(g1668_p),
    .din1(g1665_n),
    .din2(g1667_p)
  );


  FA
  g_g1669_n
  (
    .dout(g1669_n),
    .din1(g1664_p),
    .din2(g1668_p)
  );


  FA
  g_g1670_n
  (
    .dout(g1670_n),
    .din1(ffc_428_p_spl_111),
    .din2(g1653_p_spl_1)
  );


  FA
  g_g1671_n
  (
    .dout(g1671_n),
    .din1(ffc_428_n_spl_111),
    .din2(g1656_p_spl_1)
  );


  LA
  g_g1672_p
  (
    .dout(g1672_p),
    .din1(ffc_432_p_spl_11),
    .din2(g1671_n)
  );


  LA
  g_g1673_p
  (
    .dout(g1673_p),
    .din1(g1670_n),
    .din2(g1672_p)
  );


  FA
  g_g1674_n
  (
    .dout(g1674_n),
    .din1(ffc_301_n_spl_),
    .din2(ffc_428_p_spl_111)
  );


  FA
  g_g1675_n
  (
    .dout(g1675_n),
    .din1(ffc_297_n_spl_),
    .din2(ffc_428_n_spl_111)
  );


  LA
  g_g1676_p
  (
    .dout(g1676_p),
    .din1(ffc_432_n_spl_11),
    .din2(g1675_n)
  );


  LA
  g_g1677_p
  (
    .dout(g1677_p),
    .din1(g1674_n),
    .din2(g1676_p)
  );


  FA
  g_g1678_n
  (
    .dout(g1678_n),
    .din1(ffc_241_n_spl_1),
    .din2(g1677_p)
  );


  FA
  g_g1679_n
  (
    .dout(g1679_n),
    .din1(g1673_p),
    .din2(g1678_n)
  );


  FA
  g_g1680_n
  (
    .dout(g1680_n),
    .din1(ffc_301_n_spl_),
    .din2(ffc_436_p_spl_111)
  );


  FA
  g_g1681_n
  (
    .dout(g1681_n),
    .din1(ffc_297_n_spl_),
    .din2(ffc_436_n_spl_111)
  );


  LA
  g_g1682_p
  (
    .dout(g1682_p),
    .din1(g1680_n),
    .din2(g1681_n)
  );


  FA
  g_g1683_n
  (
    .dout(g1683_n),
    .din1(ffc_440_p_spl_11),
    .din2(g1682_p)
  );


  LA
  g_g1684_p
  (
    .dout(g1684_p),
    .din1(ffc_436_n_spl_111),
    .din2(g1653_p_spl_1)
  );


  LA
  g_g1685_p
  (
    .dout(g1685_p),
    .din1(ffc_436_p_spl_111),
    .din2(g1656_p_spl_1)
  );


  FA
  g_g1686_n
  (
    .dout(g1686_n),
    .din1(ffc_440_n_spl_11),
    .din2(g1685_p)
  );


  FA
  g_g1687_n
  (
    .dout(g1687_n),
    .din1(g1684_p),
    .din2(g1686_n)
  );


  LA
  g_g1688_p
  (
    .dout(g1688_p),
    .din1(g1683_n),
    .din2(g1687_n)
  );


  FA
  g_g1689_n
  (
    .dout(g1689_n),
    .din1(ffc_241_n_spl_1),
    .din2(g1688_p)
  );


  LA
  g_g1690_p
  (
    .dout(g1690_p),
    .din1(ffc_610_n_spl_0),
    .din2(ffc_783_n_spl_)
  );


  FA
  g_g1690_n
  (
    .dout(g1690_n),
    .din1(ffc_610_p_spl_0),
    .din2(ffc_783_p_spl_0)
  );


  LA
  g_g1691_p
  (
    .dout(g1691_p),
    .din1(ffc_610_p_spl_0),
    .din2(ffc_783_p_spl_0)
  );


  FA
  g_g1691_n
  (
    .dout(g1691_n),
    .din1(ffc_610_n_spl_0),
    .din2(ffc_783_n_spl_)
  );


  LA
  g_g1692_p
  (
    .dout(g1692_p),
    .din1(g1690_n_spl_),
    .din2(g1691_n)
  );


  FA
  g_g1692_n
  (
    .dout(g1692_n),
    .din1(g1690_p),
    .din2(g1691_p)
  );


  FA
  g_g1693_n
  (
    .dout(g1693_n),
    .din1(ffc_578_n_spl_00),
    .din2(ffc_624_n_spl_)
  );


  LA
  g_g1694_p
  (
    .dout(g1694_p),
    .din1(ffc_6_p_spl_0),
    .din2(ffc_601_p)
  );


  FA
  g_g1695_n
  (
    .dout(g1695_n),
    .din1(ffc_584_p),
    .din2(g1694_p)
  );


  LA
  g_g1696_p
  (
    .dout(g1696_p),
    .din1(ffc_587_p_spl_),
    .din2(g1695_n_spl_)
  );


  LA
  g_g1697_p
  (
    .dout(g1697_p),
    .din1(ffc_655_n),
    .din2(ffc_757_n)
  );


  FA
  g_g1697_n
  (
    .dout(g1697_n),
    .din1(ffc_655_p),
    .din2(ffc_757_p)
  );


  LA
  g_g1698_p
  (
    .dout(g1698_p),
    .din1(ffc_768_n),
    .din2(ffc_842_n_spl_)
  );


  FA
  g_g1698_n
  (
    .dout(g1698_n),
    .din1(ffc_768_p),
    .din2(ffc_842_p_spl_0)
  );


  LA
  g_g1699_p
  (
    .dout(g1699_p),
    .din1(ffc_817_n),
    .din2(ffc_818_n)
  );


  FA
  g_g1699_n
  (
    .dout(g1699_n),
    .din1(ffc_817_p),
    .din2(ffc_818_p)
  );


  LA
  g_g1700_p
  (
    .dout(g1700_p),
    .din1(ffc_819_n),
    .din2(ffc_820_n)
  );


  FA
  g_g1700_n
  (
    .dout(g1700_n),
    .din1(ffc_819_p),
    .din2(ffc_820_p)
  );


  LA
  g_g1701_p
  (
    .dout(g1701_p),
    .din1(ffc_823_n),
    .din2(ffc_827_n_spl_)
  );


  FA
  g_g1701_n
  (
    .dout(g1701_n),
    .din1(ffc_823_p),
    .din2(ffc_827_p_spl_)
  );


  LA
  g_g1702_p
  (
    .dout(g1702_p),
    .din1(ffc_827_n_spl_),
    .din2(ffc_828_n)
  );


  FA
  g_g1702_n
  (
    .dout(g1702_n),
    .din1(ffc_827_p_spl_),
    .din2(ffc_828_p)
  );


  LA
  g_g1703_p
  (
    .dout(g1703_p),
    .din1(ffc_840_n),
    .din2(ffc_841_p)
  );


  FA
  g_g1703_n
  (
    .dout(g1703_n),
    .din1(ffc_840_p_spl_),
    .din2(ffc_841_n)
  );


  LA
  g_g1704_p
  (
    .dout(g1704_p),
    .din1(ffc_843_p_spl_0),
    .din2(ffc_845_p_spl_)
  );


  FA
  g_g1704_n
  (
    .dout(g1704_n),
    .din1(ffc_843_n_spl_),
    .din2(ffc_845_n)
  );


  LA
  g_g1705_p
  (
    .dout(g1705_p),
    .din1(ffc_770_p_spl_0),
    .din2(g1703_p_spl_0)
  );


  FA
  g_g1705_n
  (
    .dout(g1705_n),
    .din1(ffc_770_n_spl_),
    .din2(g1703_n_spl_)
  );


  LA
  g_g1706_p
  (
    .dout(g1706_p),
    .din1(ffc_466_n_spl_000),
    .din2(ffc_581_p)
  );


  LA
  g_g1707_p
  (
    .dout(g1707_p),
    .din1(ffc_457_p_spl_000),
    .din2(ffc_581_n)
  );


  FA
  g_g1708_n
  (
    .dout(g1708_n),
    .din1(g1706_p),
    .din2(g1707_p)
  );


  LA
  g_g1709_p
  (
    .dout(g1709_p),
    .din1(ffc_623_p_spl_0),
    .din2(ffc_829_p_spl_00)
  );


  FA
  g_g1709_n
  (
    .dout(g1709_n),
    .din1(ffc_623_n_spl_),
    .din2(ffc_829_n_spl_00)
  );


  LA
  g_g1710_p
  (
    .dout(g1710_p),
    .din1(ffc_623_n_spl_),
    .din2(ffc_830_p)
  );


  FA
  g_g1710_n
  (
    .dout(g1710_n),
    .din1(ffc_623_p_spl_0),
    .din2(ffc_830_n)
  );


  LA
  g_g1711_p
  (
    .dout(g1711_p),
    .din1(g1709_n),
    .din2(g1710_n)
  );


  FA
  g_g1711_n
  (
    .dout(g1711_n),
    .din1(g1709_p),
    .din2(g1710_p)
  );


  LA
  g_g1712_p
  (
    .dout(g1712_p),
    .din1(ffc_683_n),
    .din2(ffc_775_p_spl_)
  );


  FA
  g_g1712_n
  (
    .dout(g1712_n),
    .din1(ffc_683_p_spl_),
    .din2(ffc_775_n)
  );


  LA
  g_g1713_p
  (
    .dout(g1713_p),
    .din1(ffc_814_p),
    .din2(g1698_n_spl_0)
  );


  FA
  g_g1713_n
  (
    .dout(g1713_n),
    .din1(ffc_814_n),
    .din2(g1698_p_spl_0)
  );


  LA
  g_g1714_p
  (
    .dout(g1714_p),
    .din1(ffc_813_n_spl_),
    .din2(g1713_n)
  );


  FA
  g_g1714_n
  (
    .dout(g1714_n),
    .din1(ffc_813_p_spl_),
    .din2(g1713_p)
  );


  LA
  g_g1715_p
  (
    .dout(g1715_p),
    .din1(ffc_795_p_spl_0),
    .din2(ffc_815_n_spl_)
  );


  FA
  g_g1715_n
  (
    .dout(g1715_n),
    .din1(ffc_795_n_spl_0),
    .din2(ffc_815_p_spl_)
  );


  LA
  g_g1716_p
  (
    .dout(g1716_p),
    .din1(ffc_842_n_spl_),
    .din2(g1715_n)
  );


  FA
  g_g1716_n
  (
    .dout(g1716_n),
    .din1(ffc_842_p_spl_0),
    .din2(g1715_p)
  );


  LA
  g_g1717_p
  (
    .dout(g1717_p),
    .din1(ffc_816_p_spl_00),
    .din2(g1700_n_spl_0)
  );


  FA
  g_g1717_n
  (
    .dout(g1717_n),
    .din1(ffc_816_n_spl_0),
    .din2(g1700_p_spl_)
  );


  LA
  g_g1718_p
  (
    .dout(g1718_p),
    .din1(ffc_816_n_spl_0),
    .din2(g1700_p_spl_)
  );


  FA
  g_g1718_n
  (
    .dout(g1718_n),
    .din1(ffc_816_p_spl_00),
    .din2(g1700_n_spl_0)
  );


  LA
  g_g1719_p
  (
    .dout(g1719_p),
    .din1(g1717_n_spl_),
    .din2(g1718_n)
  );


  FA
  g_g1719_n
  (
    .dout(g1719_n),
    .din1(g1717_p_spl_),
    .din2(g1718_p)
  );


  LA
  g_g1720_p
  (
    .dout(g1720_p),
    .din1(ffc_864_n),
    .din2(ffc_865_n)
  );


  FA
  g_g1720_n
  (
    .dout(g1720_n),
    .din1(ffc_864_p),
    .din2(ffc_865_p)
  );


  LA
  g_g1721_p
  (
    .dout(g1721_p),
    .din1(ffc_866_n),
    .din2(ffc_867_n)
  );


  FA
  g_g1721_n
  (
    .dout(g1721_n),
    .din1(ffc_866_p),
    .din2(ffc_867_p)
  );


  LA
  g_g1722_p
  (
    .dout(g1722_p),
    .din1(ffc_868_n),
    .din2(ffc_869_n)
  );


  FA
  g_g1722_n
  (
    .dout(g1722_n),
    .din1(ffc_868_p),
    .din2(ffc_869_p)
  );


  FA
  g_g1723_n
  (
    .dout(g1723_n),
    .din1(ffc_574_p),
    .din2(g1696_p_spl_)
  );


  LA
  g_g1724_p
  (
    .dout(g1724_p),
    .din1(ffc_603_p_spl_),
    .din2(g1723_n_spl_)
  );


  LA
  g_g1725_p
  (
    .dout(g1725_p),
    .din1(ffc_769_p_spl_0),
    .din2(ffc_844_p_spl_0)
  );


  FA
  g_g1725_n
  (
    .dout(g1725_n),
    .din1(ffc_769_n_spl_),
    .din2(ffc_844_n_spl_)
  );


  LA
  g_g1726_p
  (
    .dout(g1726_p),
    .din1(ffc_80_p),
    .din2(ffc_596_p_spl_0)
  );


  LA
  g_g1727_p
  (
    .dout(g1727_p),
    .din1(ffc_80_n),
    .din2(ffc_596_n)
  );


  FA
  g_g1728_n
  (
    .dout(g1728_n),
    .din1(g1726_p),
    .din2(g1727_p)
  );


  LA
  g_g1729_p
  (
    .dout(g1729_p),
    .din1(ffc_466_n_spl_000),
    .din2(ffc_556_n_spl_0)
  );


  LA
  g_g1730_p
  (
    .dout(g1730_p),
    .din1(ffc_463_n_spl_000),
    .din2(ffc_556_p_spl_0)
  );


  FA
  g_g1731_n
  (
    .dout(g1731_n),
    .din1(g1729_p),
    .din2(g1730_p)
  );


  LA
  g_g1732_p
  (
    .dout(g1732_p),
    .din1(ffc_580_p),
    .din2(g1731_n)
  );


  LA
  g_g1733_p
  (
    .dout(g1733_p),
    .din1(ffc_460_p_spl_000),
    .din2(ffc_556_p_spl_0)
  );


  LA
  g_g1734_p
  (
    .dout(g1734_p),
    .din1(ffc_457_p_spl_000),
    .din2(ffc_556_n_spl_0)
  );


  FA
  g_g1735_n
  (
    .dout(g1735_n),
    .din1(g1733_p),
    .din2(g1734_p)
  );


  LA
  g_g1736_p
  (
    .dout(g1736_p),
    .din1(ffc_580_n),
    .din2(g1735_n)
  );


  FA
  g_g1737_n
  (
    .dout(g1737_n),
    .din1(g1732_p),
    .din2(g1736_p)
  );


  LA
  g_g1738_p
  (
    .dout(g1738_p),
    .din1(ffc_466_n_spl_001),
    .din2(ffc_527_n_spl_0)
  );


  LA
  g_g1739_p
  (
    .dout(g1739_p),
    .din1(ffc_463_n_spl_000),
    .din2(ffc_527_p_spl_0)
  );


  FA
  g_g1740_n
  (
    .dout(g1740_n),
    .din1(g1738_p),
    .din2(g1739_p)
  );


  LA
  g_g1741_p
  (
    .dout(g1741_p),
    .din1(ffc_543_p),
    .din2(g1740_n)
  );


  LA
  g_g1742_p
  (
    .dout(g1742_p),
    .din1(ffc_460_p_spl_000),
    .din2(ffc_527_p_spl_0)
  );


  LA
  g_g1743_p
  (
    .dout(g1743_p),
    .din1(ffc_457_p_spl_001),
    .din2(ffc_527_n_spl_0)
  );


  FA
  g_g1744_n
  (
    .dout(g1744_n),
    .din1(g1742_p),
    .din2(g1743_p)
  );


  LA
  g_g1745_p
  (
    .dout(g1745_p),
    .din1(ffc_543_n),
    .din2(g1744_n)
  );


  FA
  g_g1746_n
  (
    .dout(g1746_n),
    .din1(g1741_p),
    .din2(g1745_p)
  );


  LA
  g_g1747_p
  (
    .dout(g1747_p),
    .din1(ffc_466_n_spl_001),
    .din2(ffc_590_n_spl_0)
  );


  LA
  g_g1748_p
  (
    .dout(g1748_p),
    .din1(ffc_463_n_spl_001),
    .din2(ffc_590_p_spl_0)
  );


  FA
  g_g1749_n
  (
    .dout(g1749_n),
    .din1(g1747_p),
    .din2(g1748_p)
  );


  LA
  g_g1750_p
  (
    .dout(g1750_p),
    .din1(ffc_607_p),
    .din2(g1749_n)
  );


  LA
  g_g1751_p
  (
    .dout(g1751_p),
    .din1(ffc_460_p_spl_001),
    .din2(ffc_590_p_spl_0)
  );


  LA
  g_g1752_p
  (
    .dout(g1752_p),
    .din1(ffc_457_p_spl_001),
    .din2(ffc_590_n_spl_0)
  );


  FA
  g_g1753_n
  (
    .dout(g1753_n),
    .din1(g1751_p),
    .din2(g1752_p)
  );


  LA
  g_g1754_p
  (
    .dout(g1754_p),
    .din1(ffc_607_n),
    .din2(g1753_n)
  );


  FA
  g_g1755_n
  (
    .dout(g1755_n),
    .din1(g1750_p),
    .din2(g1754_p)
  );


  LA
  g_g1756_p
  (
    .dout(g1756_p),
    .din1(ffc_390_p_spl_00),
    .din2(g1711_n_spl_0)
  );


  FA
  g_g1756_n
  (
    .dout(g1756_n),
    .din1(ffc_390_n_spl_0),
    .din2(g1711_p_spl_)
  );


  LA
  g_g1757_p
  (
    .dout(g1757_p),
    .din1(ffc_390_n_spl_0),
    .din2(g1711_p_spl_)
  );


  FA
  g_g1757_n
  (
    .dout(g1757_n),
    .din1(ffc_390_p_spl_00),
    .din2(g1711_n_spl_0)
  );


  LA
  g_g1758_p
  (
    .dout(g1758_p),
    .din1(g1756_n),
    .din2(g1757_n)
  );


  FA
  g_g1758_n
  (
    .dout(g1758_n),
    .din1(g1756_p_spl_),
    .din2(g1757_p)
  );


  LA
  g_g1759_p
  (
    .dout(g1759_p),
    .din1(ffc_839_p_spl_000),
    .din2(ffc_859_p_spl_)
  );


  FA
  g_g1759_n
  (
    .dout(g1759_n),
    .din1(ffc_839_n_spl_000),
    .din2(ffc_859_n)
  );


  LA
  g_g1760_p
  (
    .dout(g1760_p),
    .din1(ffc_839_n_spl_000),
    .din2(ffc_860_p)
  );


  FA
  g_g1760_n
  (
    .dout(g1760_n),
    .din1(ffc_839_p_spl_000),
    .din2(ffc_860_n)
  );


  LA
  g_g1761_p
  (
    .dout(g1761_p),
    .din1(g1759_n),
    .din2(g1760_n)
  );


  FA
  g_g1761_n
  (
    .dout(g1761_n),
    .din1(g1759_p),
    .din2(g1760_p)
  );


  LA
  g_g1762_p
  (
    .dout(g1762_p),
    .din1(ffc_857_p_spl_0),
    .din2(g1721_n_spl_0)
  );


  FA
  g_g1762_n
  (
    .dout(g1762_n),
    .din1(ffc_857_n),
    .din2(g1721_p)
  );


  FA
  g_g1763_n
  (
    .dout(g1763_n),
    .din1(ffc_857_p_spl_0),
    .din2(g1721_n_spl_0)
  );


  LA
  g_g1764_p
  (
    .dout(g1764_p),
    .din1(ffc_858_p_spl_0),
    .din2(g1720_n_spl_0)
  );


  FA
  g_g1764_n
  (
    .dout(g1764_n),
    .din1(ffc_858_n),
    .din2(g1720_p)
  );


  LA
  g_g1765_p
  (
    .dout(g1765_p),
    .din1(ffc_861_p_spl_),
    .din2(ffc_863_p_spl_000)
  );


  FA
  g_g1765_n
  (
    .dout(g1765_n),
    .din1(ffc_861_n),
    .din2(ffc_863_n_spl_000)
  );


  LA
  g_g1766_p
  (
    .dout(g1766_p),
    .din1(ffc_862_p),
    .din2(ffc_863_n_spl_000)
  );


  FA
  g_g1766_n
  (
    .dout(g1766_n),
    .din1(ffc_862_n),
    .din2(ffc_863_p_spl_000)
  );


  LA
  g_g1767_p
  (
    .dout(g1767_p),
    .din1(g1765_n),
    .din2(g1766_n)
  );


  FA
  g_g1767_n
  (
    .dout(g1767_n),
    .din1(g1765_p),
    .din2(g1766_p)
  );


  FA
  g_g1768_n
  (
    .dout(g1768_n),
    .din1(ffc_769_p_spl_0),
    .din2(ffc_844_p_spl_0)
  );


  LA
  g_g1769_p
  (
    .dout(g1769_p),
    .din1(g1698_n_spl_0),
    .din2(g1704_p_spl_)
  );


  FA
  g_g1769_n
  (
    .dout(g1769_n),
    .din1(g1698_p_spl_0),
    .din2(g1704_n)
  );


  LA
  g_g1770_p
  (
    .dout(g1770_p),
    .din1(ffc_813_p_spl_),
    .din2(ffc_843_p_spl_0)
  );


  FA
  g_g1770_n
  (
    .dout(g1770_n),
    .din1(ffc_813_n_spl_),
    .din2(ffc_843_n_spl_)
  );


  LA
  g_g1771_p
  (
    .dout(g1771_p),
    .din1(ffc_796_n),
    .din2(g1770_n)
  );


  FA
  g_g1771_n
  (
    .dout(g1771_n),
    .din1(ffc_796_p),
    .din2(g1770_p)
  );


  LA
  g_g1772_p
  (
    .dout(g1772_p),
    .din1(g1769_n),
    .din2(g1771_p)
  );


  FA
  g_g1772_n
  (
    .dout(g1772_n),
    .din1(g1769_p),
    .din2(g1771_n)
  );


  LA
  g_g1773_p
  (
    .dout(g1773_p),
    .din1(g1719_p_spl_0),
    .din2(g1772_n_spl_)
  );


  FA
  g_g1773_n
  (
    .dout(g1773_n),
    .din1(g1719_n_spl_),
    .din2(g1772_p_spl_)
  );


  LA
  g_g1774_p
  (
    .dout(g1774_p),
    .din1(g1717_n_spl_),
    .din2(g1773_n_spl_)
  );


  FA
  g_g1774_n
  (
    .dout(g1774_n),
    .din1(g1717_p_spl_),
    .din2(g1773_p_spl_)
  );


  LA
  g_g1775_p
  (
    .dout(g1775_p),
    .din1(ffc_839_p_spl_001),
    .din2(ffc_850_p_spl_)
  );


  FA
  g_g1775_n
  (
    .dout(g1775_n),
    .din1(ffc_839_n_spl_00),
    .din2(ffc_850_n)
  );


  LA
  g_g1776_p
  (
    .dout(g1776_p),
    .din1(ffc_839_n_spl_01),
    .din2(ffc_851_p)
  );


  FA
  g_g1776_n
  (
    .dout(g1776_n),
    .din1(ffc_839_p_spl_001),
    .din2(ffc_851_n)
  );


  LA
  g_g1777_p
  (
    .dout(g1777_p),
    .din1(g1775_n),
    .din2(g1776_n)
  );


  FA
  g_g1777_n
  (
    .dout(g1777_n),
    .din1(g1775_p),
    .din2(g1776_p)
  );


  LA
  g_g1778_p
  (
    .dout(g1778_p),
    .din1(ffc_839_p_spl_01),
    .din2(ffc_852_p_spl_)
  );


  FA
  g_g1778_n
  (
    .dout(g1778_n),
    .din1(ffc_839_n_spl_01),
    .din2(ffc_852_n)
  );


  LA
  g_g1779_p
  (
    .dout(g1779_p),
    .din1(ffc_839_n_spl_10),
    .din2(ffc_853_p)
  );


  FA
  g_g1779_n
  (
    .dout(g1779_n),
    .din1(ffc_839_p_spl_01),
    .din2(ffc_853_n)
  );


  LA
  g_g1780_p
  (
    .dout(g1780_p),
    .din1(g1778_n),
    .din2(g1779_n)
  );


  FA
  g_g1780_n
  (
    .dout(g1780_n),
    .din1(g1778_p),
    .din2(g1779_p)
  );


  LA
  g_g1781_p
  (
    .dout(g1781_p),
    .din1(ffc_824_n),
    .din2(ffc_835_p)
  );


  FA
  g_g1781_n
  (
    .dout(g1781_n),
    .din1(ffc_824_p),
    .din2(ffc_835_n)
  );


  LA
  g_g1782_p
  (
    .dout(g1782_p),
    .din1(g1699_p_spl_0),
    .din2(g1781_p_spl_)
  );


  FA
  g_g1782_n
  (
    .dout(g1782_n),
    .din1(g1699_n_spl_0),
    .din2(g1781_n_spl_)
  );


  LA
  g_g1783_p
  (
    .dout(g1783_p),
    .din1(g1699_n_spl_0),
    .din2(g1781_n_spl_)
  );


  FA
  g_g1783_n
  (
    .dout(g1783_n),
    .din1(g1699_p_spl_0),
    .din2(g1781_p_spl_)
  );


  LA
  g_g1784_p
  (
    .dout(g1784_p),
    .din1(g1782_n),
    .din2(g1783_n)
  );


  FA
  g_g1784_n
  (
    .dout(g1784_n),
    .din1(g1782_p),
    .din2(g1783_p)
  );


  LA
  g_g1785_p
  (
    .dout(g1785_p),
    .din1(g1712_n),
    .din2(g1784_p)
  );


  LA
  g_g1786_p
  (
    .dout(g1786_p),
    .din1(g1712_p_spl_0),
    .din2(g1784_n)
  );


  FA
  g_g1787_n
  (
    .dout(g1787_n),
    .din1(g1785_p_spl_),
    .din2(g1786_p)
  );


  LA
  g_g1788_p
  (
    .dout(g1788_p),
    .din1(ffc_854_p_spl_),
    .din2(ffc_863_p_spl_001)
  );


  LA
  g_g1789_p
  (
    .dout(g1789_p),
    .din1(ffc_855_p),
    .din2(ffc_863_n_spl_001)
  );


  FA
  g_g1790_n
  (
    .dout(g1790_n),
    .din1(g1788_p),
    .din2(g1789_p)
  );


  LA
  g_g1791_p
  (
    .dout(g1791_p),
    .din1(g1719_n_spl_),
    .din2(g1772_p_spl_)
  );


  FA
  g_g1791_n
  (
    .dout(g1791_n),
    .din1(g1719_p_spl_0),
    .din2(g1772_n_spl_)
  );


  LA
  g_g1792_p
  (
    .dout(g1792_p),
    .din1(g1773_n_spl_),
    .din2(g1791_n)
  );


  FA
  g_g1792_n
  (
    .dout(g1792_n),
    .din1(g1773_p_spl_),
    .din2(g1791_p)
  );


  LA
  g_g1793_p
  (
    .dout(g1793_p),
    .din1(ffc_848_p_spl_0),
    .din2(g1761_n_spl_0)
  );


  FA
  g_g1793_n
  (
    .dout(g1793_n),
    .din1(ffc_848_n),
    .din2(g1761_p)
  );


  LA
  g_g1794_p
  (
    .dout(g1794_p),
    .din1(ffc_856_p_spl_0),
    .din2(g1722_n_spl_0)
  );


  FA
  g_g1794_n
  (
    .dout(g1794_n),
    .din1(ffc_856_n),
    .din2(g1722_p)
  );


  FA
  g_g1795_n
  (
    .dout(g1795_n),
    .din1(ffc_856_p_spl_0),
    .din2(g1722_n_spl_0)
  );


  LA
  g_g1796_p
  (
    .dout(g1796_p),
    .din1(g1794_n),
    .din2(g1795_n)
  );


  LA
  g_g1797_p
  (
    .dout(g1797_p),
    .din1(g1762_n),
    .din2(g1763_n_spl_0)
  );


  FA
  g_g1798_n
  (
    .dout(g1798_n),
    .din1(ffc_858_p_spl_0),
    .din2(g1720_n_spl_0)
  );


  LA
  g_g1799_p
  (
    .dout(g1799_p),
    .din1(g1764_n),
    .din2(g1798_n)
  );


  LA
  g_g1800_p
  (
    .dout(g1800_p),
    .din1(ffc_846_p_spl_),
    .din2(ffc_863_p_spl_001)
  );


  FA
  g_g1800_n
  (
    .dout(g1800_n),
    .din1(ffc_846_n),
    .din2(ffc_863_n_spl_001)
  );


  LA
  g_g1801_p
  (
    .dout(g1801_p),
    .din1(ffc_847_p_spl_),
    .din2(ffc_863_n_spl_010)
  );


  FA
  g_g1801_n
  (
    .dout(g1801_n),
    .din1(ffc_847_n),
    .din2(ffc_863_p_spl_010)
  );


  LA
  g_g1802_p
  (
    .dout(g1802_p),
    .din1(g1800_n),
    .din2(g1801_n)
  );


  FA
  g_g1802_n
  (
    .dout(g1802_n),
    .din1(g1800_p),
    .din2(g1801_p)
  );


  LA
  g_g1803_p
  (
    .dout(g1803_p),
    .din1(ffc_388_p_spl_0),
    .din2(g1780_n_spl_0)
  );


  FA
  g_g1803_n
  (
    .dout(g1803_n),
    .din1(ffc_388_n),
    .din2(g1780_p)
  );


  LA
  g_g1804_p
  (
    .dout(g1804_p),
    .din1(ffc_392_p_spl_0),
    .din2(g1777_n_spl_0)
  );


  FA
  g_g1804_n
  (
    .dout(g1804_n),
    .din1(ffc_392_n),
    .din2(g1777_p)
  );


  LA
  g_g1805_p
  (
    .dout(g1805_p),
    .din1(ffc_393_p_spl_0),
    .din2(g1790_n_spl_0)
  );


  LA
  g_g1806_p
  (
    .dout(g1806_p),
    .din1(ffc_849_p_spl_0),
    .din2(g1767_n_spl_0)
  );


  FA
  g_g1806_n
  (
    .dout(g1806_n),
    .din1(ffc_849_n),
    .din2(g1767_p)
  );


  FA
  g_g1807_n
  (
    .dout(g1807_n),
    .din1(ffc_849_p_spl_0),
    .din2(g1767_n_spl_0)
  );


  LA
  g_g1808_p
  (
    .dout(g1808_p),
    .din1(g1806_n),
    .din2(g1807_n_spl_)
  );


  LA
  g_g1809_p
  (
    .dout(g1809_p),
    .din1(g1797_p_spl_),
    .din2(g1799_p_spl_0)
  );


  LA
  g_g1810_p
  (
    .dout(g1810_p),
    .din1(ffc_73_p),
    .din2(ffc_497_n_spl_000)
  );


  LA
  g_g1811_p
  (
    .dout(g1811_p),
    .din1(ffc_170_p),
    .din2(ffc_497_n_spl_000)
  );


  LA
  g_g1812_p
  (
    .dout(g1812_p),
    .din1(ffc_180_p),
    .din2(ffc_497_n_spl_001)
  );


  FA
  g_g1813_n
  (
    .dout(g1813_n),
    .din1(ffc_183_p),
    .din2(ffc_497_p_spl_000)
  );


  FA
  g_g1814_n
  (
    .dout(g1814_n),
    .din1(ffc_190_p),
    .din2(ffc_497_p_spl_000)
  );


  LA
  g_g1815_p
  (
    .dout(g1815_p),
    .din1(ffc_197_p),
    .din2(ffc_497_n_spl_001)
  );


  LA
  g_g1816_p
  (
    .dout(g1816_p),
    .din1(ffc_216_p),
    .din2(ffc_497_n_spl_010)
  );


  FA
  g_g1817_n
  (
    .dout(g1817_n),
    .din1(ffc_219_p),
    .din2(ffc_497_p_spl_001)
  );


  FA
  g_g1818_n
  (
    .dout(g1818_n),
    .din1(ffc_225_p),
    .din2(ffc_497_p_spl_001)
  );


  LA
  g_g1819_p
  (
    .dout(g1819_p),
    .din1(ffc_466_n_spl_010),
    .din2(ffc_528_n_spl_0)
  );


  LA
  g_g1820_p
  (
    .dout(g1820_p),
    .din1(ffc_463_n_spl_001),
    .din2(ffc_528_p_spl_0)
  );


  FA
  g_g1821_n
  (
    .dout(g1821_n),
    .din1(g1819_p),
    .din2(g1820_p)
  );


  LA
  g_g1822_p
  (
    .dout(g1822_p),
    .din1(ffc_542_p),
    .din2(g1821_n)
  );


  LA
  g_g1823_p
  (
    .dout(g1823_p),
    .din1(ffc_460_p_spl_001),
    .din2(ffc_528_p_spl_0)
  );


  LA
  g_g1824_p
  (
    .dout(g1824_p),
    .din1(ffc_457_p_spl_010),
    .din2(ffc_528_n_spl_0)
  );


  FA
  g_g1825_n
  (
    .dout(g1825_n),
    .din1(g1823_p),
    .din2(g1824_p)
  );


  LA
  g_g1826_p
  (
    .dout(g1826_p),
    .din1(ffc_542_n),
    .din2(g1825_n)
  );


  LA
  g_g1827_p
  (
    .dout(g1827_p),
    .din1(ffc_493_n_spl_0),
    .din2(ffc_497_p_spl_010)
  );


  FA
  g_g1828_n
  (
    .dout(g1828_n),
    .din1(ffc_204_p_spl_),
    .din2(ffc_497_p_spl_010)
  );


  LA
  g_g1829_p
  (
    .dout(g1829_p),
    .din1(ffc_493_p_spl_0),
    .din2(g1828_n)
  );


  LA
  g_g1830_p
  (
    .dout(g1830_p),
    .din1(ffc_604_n_spl_),
    .din2(ffc_605_n)
  );


  FA
  g_g1830_n
  (
    .dout(g1830_n),
    .din1(ffc_604_p_spl_),
    .din2(ffc_605_p_spl_0)
  );


  LA
  g_g1831_p
  (
    .dout(g1831_p),
    .din1(ffc_615_n),
    .din2(g1830_n)
  );


  FA
  g_g1831_n
  (
    .dout(g1831_n),
    .din1(ffc_615_p_spl_),
    .din2(g1830_p)
  );


  LA
  g_g1832_p
  (
    .dout(g1832_p),
    .din1(ffc_791_p_spl_),
    .din2(ffc_811_p_spl_)
  );


  FA
  g_g1832_n
  (
    .dout(g1832_n),
    .din1(ffc_791_n_spl_),
    .din2(ffc_811_n_spl_)
  );


  LA
  g_g1833_p
  (
    .dout(g1833_p),
    .din1(ffc_791_n_spl_),
    .din2(ffc_811_n_spl_)
  );


  FA
  g_g1833_n
  (
    .dout(g1833_n),
    .din1(ffc_791_p_spl_),
    .din2(ffc_811_p_spl_)
  );


  LA
  g_g1834_p
  (
    .dout(g1834_p),
    .din1(g1832_n),
    .din2(g1833_n)
  );


  FA
  g_g1834_n
  (
    .dout(g1834_n),
    .din1(g1832_p),
    .din2(g1833_p)
  );


  LA
  g_g1835_p
  (
    .dout(g1835_p),
    .din1(g1831_p_spl_),
    .din2(g1834_n_spl_)
  );


  FA
  g_g1835_n
  (
    .dout(g1835_n),
    .din1(g1831_n_spl_),
    .din2(g1834_p_spl_)
  );


  LA
  g_g1836_p
  (
    .dout(g1836_p),
    .din1(g1831_n_spl_),
    .din2(g1834_p_spl_)
  );


  FA
  g_g1836_n
  (
    .dout(g1836_n),
    .din1(g1831_p_spl_),
    .din2(g1834_n_spl_)
  );


  LA
  g_g1837_p
  (
    .dout(g1837_p),
    .din1(g1835_n),
    .din2(g1836_n)
  );


  FA
  g_g1837_n
  (
    .dout(g1837_n),
    .din1(g1835_p),
    .din2(g1836_p)
  );


  LA
  g_g1838_p
  (
    .dout(g1838_p),
    .din1(ffc_578_p_spl_),
    .din2(ffc_668_p)
  );


  FA
  g_g1838_n
  (
    .dout(g1838_n),
    .din1(ffc_578_n_spl_00),
    .din2(ffc_668_n)
  );


  LA
  g_g1839_p
  (
    .dout(g1839_p),
    .din1(ffc_578_n_spl_0),
    .din2(ffc_808_n)
  );


  FA
  g_g1839_n
  (
    .dout(g1839_n),
    .din1(ffc_578_p_spl_),
    .din2(ffc_808_p)
  );


  LA
  g_g1840_p
  (
    .dout(g1840_p),
    .din1(g1838_n),
    .din2(g1839_n)
  );


  FA
  g_g1840_n
  (
    .dout(g1840_n),
    .din1(g1838_p),
    .din2(g1839_p)
  );


  LA
  g_g1841_p
  (
    .dout(g1841_p),
    .din1(g1692_p_spl_0),
    .din2(g1840_n_spl_)
  );


  FA
  g_g1841_n
  (
    .dout(g1841_n),
    .din1(g1692_n_spl_0),
    .din2(g1840_p_spl_)
  );


  LA
  g_g1842_p
  (
    .dout(g1842_p),
    .din1(g1692_n_spl_0),
    .din2(g1840_p_spl_)
  );


  FA
  g_g1842_n
  (
    .dout(g1842_n),
    .din1(g1692_p_spl_0),
    .din2(g1840_n_spl_)
  );


  LA
  g_g1843_p
  (
    .dout(g1843_p),
    .din1(g1841_n),
    .din2(g1842_n)
  );


  FA
  g_g1843_n
  (
    .dout(g1843_n),
    .din1(g1841_p),
    .din2(g1842_p)
  );


  LA
  g_g1844_p
  (
    .dout(g1844_p),
    .din1(g1837_n),
    .din2(g1843_p)
  );


  LA
  g_g1845_p
  (
    .dout(g1845_p),
    .din1(g1837_p),
    .din2(g1843_n)
  );


  FA
  g_g1846_n
  (
    .dout(g1846_n),
    .din1(g1844_p),
    .din2(g1845_p)
  );


  LA
  g_g1847_p
  (
    .dout(g1847_p),
    .din1(ffc_493_n_spl_0),
    .din2(g1846_n)
  );


  FA
  g_g1848_n
  (
    .dout(g1848_n),
    .din1(ffc_497_n_spl_010),
    .din2(g1755_n_spl_)
  );


  FA
  g_g1849_n
  (
    .dout(g1849_n),
    .din1(ffc_497_n_spl_01),
    .din2(g1737_n_spl_)
  );


  LA
  g_g1850_p
  (
    .dout(g1850_p),
    .din1(ffc_497_p_spl_011),
    .din2(ffc_762_n)
  );


  LA
  g_g1851_p
  (
    .dout(g1851_p),
    .din1(ffc_497_p_spl_011),
    .din2(ffc_761_p)
  );


  LA
  g_g1852_p
  (
    .dout(g1852_p),
    .din1(ffc_497_p_spl_100),
    .din2(ffc_758_n)
  );


  FA
  g_g1853_n
  (
    .dout(g1853_n),
    .din1(ffc_497_n_spl_10),
    .din2(g1746_n_spl_)
  );


  LA
  g_g1854_p
  (
    .dout(g1854_p),
    .din1(ffc_806_n),
    .din2(ffc_807_n)
  );


  FA
  g_g1854_n
  (
    .dout(g1854_n),
    .din1(ffc_806_p),
    .din2(ffc_807_p)
  );


  LA
  g_g1855_p
  (
    .dout(g1855_p),
    .din1(ffc_804_n),
    .din2(ffc_805_n)
  );


  FA
  g_g1855_n
  (
    .dout(g1855_n),
    .din1(ffc_804_p),
    .din2(ffc_805_p)
  );


  LA
  g_g1856_p
  (
    .dout(g1856_p),
    .din1(g1854_p_spl_),
    .din2(g1855_n_spl_)
  );


  FA
  g_g1856_n
  (
    .dout(g1856_n),
    .din1(g1854_n_spl_),
    .din2(g1855_p_spl_)
  );


  LA
  g_g1857_p
  (
    .dout(g1857_p),
    .din1(g1854_n_spl_),
    .din2(g1855_p_spl_)
  );


  FA
  g_g1857_n
  (
    .dout(g1857_n),
    .din1(g1854_p_spl_),
    .din2(g1855_n_spl_)
  );


  LA
  g_g1858_p
  (
    .dout(g1858_p),
    .din1(g1856_n),
    .din2(g1857_n)
  );


  FA
  g_g1858_n
  (
    .dout(g1858_n),
    .din1(g1856_p),
    .din2(g1857_p)
  );


  LA
  g_g1859_p
  (
    .dout(g1859_p),
    .din1(ffc_802_n),
    .din2(ffc_803_p)
  );


  FA
  g_g1859_n
  (
    .dout(g1859_n),
    .din1(ffc_802_p_spl_),
    .din2(ffc_803_n)
  );


  LA
  g_g1860_p
  (
    .dout(g1860_p),
    .din1(ffc_800_n),
    .din2(ffc_801_n)
  );


  FA
  g_g1860_n
  (
    .dout(g1860_n),
    .din1(ffc_800_p_spl_),
    .din2(ffc_801_p)
  );


  LA
  g_g1861_p
  (
    .dout(g1861_p),
    .din1(g1859_p_spl_),
    .din2(g1860_p_spl_)
  );


  FA
  g_g1861_n
  (
    .dout(g1861_n),
    .din1(g1859_n_spl_),
    .din2(g1860_n_spl_)
  );


  LA
  g_g1862_p
  (
    .dout(g1862_p),
    .din1(g1859_n_spl_),
    .din2(g1860_n_spl_)
  );


  FA
  g_g1862_n
  (
    .dout(g1862_n),
    .din1(g1859_p_spl_),
    .din2(g1860_p_spl_)
  );


  LA
  g_g1863_p
  (
    .dout(g1863_p),
    .din1(g1861_n),
    .din2(g1862_n)
  );


  FA
  g_g1863_n
  (
    .dout(g1863_n),
    .din1(g1861_p),
    .din2(g1862_p)
  );


  LA
  g_g1864_p
  (
    .dout(g1864_p),
    .din1(g1858_p),
    .din2(g1863_p)
  );


  LA
  g_g1865_p
  (
    .dout(g1865_p),
    .din1(g1858_n),
    .din2(g1863_n)
  );


  FA
  g_g1866_n
  (
    .dout(g1866_n),
    .din1(ffc_493_n_spl_),
    .din2(g1865_p)
  );


  FA
  g_g1867_n
  (
    .dout(g1867_n),
    .din1(g1864_p),
    .din2(g1866_n)
  );


  LA
  g_g1868_p
  (
    .dout(g1868_p),
    .din1(ffc_497_p_spl_100),
    .din2(g1867_n)
  );


  LA
  g_g1869_p
  (
    .dout(g1869_p),
    .din1(ffc_555_n),
    .din2(ffc_565_p)
  );


  LA
  g_g1870_p
  (
    .dout(g1870_p),
    .din1(ffc_555_p),
    .din2(ffc_565_n)
  );


  LA
  g_g1871_p
  (
    .dout(g1871_p),
    .din1(ffc_6_p_spl_0),
    .din2(ffc_772_p_spl_0)
  );


  FA
  g_g1871_n
  (
    .dout(g1871_n),
    .din1(ffc_6_n_spl_),
    .din2(ffc_772_n_spl_0)
  );


  LA
  g_g1872_p
  (
    .dout(g1872_p),
    .din1(ffc_771_n_spl_0),
    .din2(g1871_n)
  );


  FA
  g_g1872_n
  (
    .dout(g1872_n),
    .din1(ffc_771_p_spl_00),
    .din2(g1871_p)
  );


  LA
  g_g1873_p
  (
    .dout(g1873_p),
    .din1(ffc_567_n),
    .din2(g1872_n_spl_00)
  );


  LA
  g_g1874_p
  (
    .dout(g1874_p),
    .din1(ffc_567_p),
    .din2(g1872_p_spl_00)
  );


  LA
  g_g1875_p
  (
    .dout(g1875_p),
    .din1(ffc_591_p),
    .din2(ffc_659_p_spl_)
  );


  LA
  g_g1876_p
  (
    .dout(g1876_p),
    .din1(ffc_576_n),
    .din2(ffc_659_n_spl_0)
  );


  FA
  g_g1877_n
  (
    .dout(g1877_n),
    .din1(g1875_p),
    .din2(g1876_p)
  );


  FA
  g_g1878_n
  (
    .dout(g1878_n),
    .din1(ffc_578_n_spl_1),
    .din2(g1877_n_spl_)
  );


  LA
  g_g1879_p
  (
    .dout(g1879_p),
    .din1(ffc_578_n_spl_1),
    .din2(g1877_n_spl_)
  );


  FA
  g_g1880_n
  (
    .dout(g1880_n),
    .din1(ffc_587_p_spl_),
    .din2(g1695_n_spl_)
  );


  FA
  g_g1881_n
  (
    .dout(g1881_n),
    .din1(ffc_594_p),
    .din2(g1724_p_spl_)
  );


  LA
  g_g1882_p
  (
    .dout(g1882_p),
    .din1(ffc_375_p_spl_0),
    .din2(ffc_538_p)
  );


  LA
  g_g1883_p
  (
    .dout(g1883_p),
    .din1(ffc_378_p),
    .din2(ffc_538_n)
  );


  FA
  g_g1884_n
  (
    .dout(g1884_n),
    .din1(g1882_p),
    .din2(g1883_p)
  );


  FA
  g_g1885_n
  (
    .dout(g1885_n),
    .din1(ffc_596_p_spl_0),
    .din2(g1884_n_spl_)
  );


  LA
  g_g1886_p
  (
    .dout(g1886_p),
    .din1(ffc_596_p_spl_),
    .din2(g1884_n_spl_)
  );


  FA
  g_g1887_n
  (
    .dout(g1887_n),
    .din1(ffc_603_p_spl_),
    .din2(g1723_n_spl_)
  );


  LA
  g_g1888_p
  (
    .dout(g1888_p),
    .din1(ffc_605_p_spl_0),
    .din2(ffc_609_p_spl_)
  );


  FA
  g_g1889_n
  (
    .dout(g1889_n),
    .din1(ffc_605_p_spl_),
    .din2(ffc_609_p_spl_)
  );


  FA
  g_g1890_n
  (
    .dout(g1890_n),
    .din1(ffc_659_n_spl_0),
    .din2(g1693_n_spl_)
  );


  LA
  g_g1891_p
  (
    .dout(g1891_p),
    .din1(ffc_593_n),
    .din2(g1890_n)
  );


  LA
  g_g1892_p
  (
    .dout(g1892_p),
    .din1(ffc_610_n_spl_1),
    .din2(g1891_p_spl_)
  );


  FA
  g_g1893_n
  (
    .dout(g1893_n),
    .din1(ffc_610_n_spl_1),
    .din2(g1891_p_spl_)
  );


  FA
  g_g1894_n
  (
    .dout(g1894_n),
    .din1(g1692_n_spl_),
    .din2(g1728_n_spl_)
  );


  LA
  g_g1895_p
  (
    .dout(g1895_p),
    .din1(ffc_6_p_spl_1),
    .din2(ffc_592_p_spl_)
  );


  FA
  g_g1895_n
  (
    .dout(g1895_n),
    .din1(ffc_6_n_spl_),
    .din2(ffc_592_n)
  );


  FA
  g_g1896_n
  (
    .dout(g1896_n),
    .din1(ffc_6_p_spl_1),
    .din2(ffc_592_p_spl_)
  );


  LA
  g_g1897_p
  (
    .dout(g1897_p),
    .din1(g1895_n_spl_),
    .din2(g1896_n)
  );


  LA
  g_g1898_p
  (
    .dout(g1898_p),
    .din1(ffc_364_n),
    .din2(ffc_863_n_spl_010)
  );


  FA
  g_g1898_n
  (
    .dout(g1898_n),
    .din1(ffc_364_p_spl_),
    .din2(ffc_863_p_spl_010)
  );


  LA
  g_g1899_p
  (
    .dout(g1899_p),
    .din1(ffc_167_p),
    .din2(ffc_497_n_spl_10)
  );


  LA
  g_g1900_p
  (
    .dout(g1900_p),
    .din1(ffc_497_p_spl_101),
    .din2(ffc_759_n)
  );


  FA
  g_g1901_n
  (
    .dout(g1901_n),
    .din1(g1899_p),
    .din2(g1900_p)
  );


  LA
  g_g1902_p
  (
    .dout(g1902_p),
    .din1(ffc_177_p),
    .din2(ffc_497_n_spl_11)
  );


  LA
  g_g1903_p
  (
    .dout(g1903_p),
    .din1(ffc_497_p_spl_101),
    .din2(ffc_790_n_spl_0)
  );


  FA
  g_g1904_n
  (
    .dout(g1904_n),
    .din1(g1902_p),
    .din2(g1903_p)
  );


  FA
  g_g1905_n
  (
    .dout(g1905_n),
    .din1(ffc_222_n),
    .din2(ffc_497_p_spl_11)
  );


  FA
  g_g1906_n
  (
    .dout(g1906_n),
    .din1(ffc_497_n_spl_11),
    .din2(g1708_n_spl_)
  );


  LA
  g_g1907_p
  (
    .dout(g1907_p),
    .din1(g1905_n),
    .din2(g1906_n)
  );


  FA
  g_g1908_n
  (
    .dout(g1908_n),
    .din1(ffc_539_p_spl_0),
    .din2(ffc_569_p)
  );


  FA
  g_g1909_n
  (
    .dout(g1909_n),
    .din1(ffc_539_n_spl_0),
    .din2(ffc_569_n)
  );


  LA
  g_g1910_p
  (
    .dout(g1910_p),
    .din1(g1908_n),
    .din2(g1909_n)
  );


  LA
  g_g1911_p
  (
    .dout(g1911_p),
    .din1(ffc_526_p_spl_0),
    .din2(ffc_527_n_spl_)
  );


  LA
  g_g1912_p
  (
    .dout(g1912_p),
    .din1(ffc_526_n_spl_0),
    .din2(ffc_527_p_spl_)
  );


  FA
  g_g1913_n
  (
    .dout(g1913_n),
    .din1(g1911_p),
    .din2(g1912_p)
  );


  LA
  g_g1914_p
  (
    .dout(g1914_p),
    .din1(ffc_528_n_spl_),
    .din2(ffc_540_p_spl_0)
  );


  LA
  g_g1915_p
  (
    .dout(g1915_p),
    .din1(ffc_528_p_spl_),
    .din2(ffc_540_n_spl_0)
  );


  FA
  g_g1916_n
  (
    .dout(g1916_n),
    .din1(g1914_p),
    .din2(g1915_p)
  );


  LA
  g_g1917_p
  (
    .dout(g1917_p),
    .din1(ffc_466_n_spl_010),
    .din2(ffc_536_n_spl_0)
  );


  LA
  g_g1918_p
  (
    .dout(g1918_p),
    .din1(ffc_463_n_spl_010),
    .din2(ffc_536_p_spl_0)
  );


  FA
  g_g1919_n
  (
    .dout(g1919_n),
    .din1(g1917_p),
    .din2(g1918_p)
  );


  LA
  g_g1920_p
  (
    .dout(g1920_p),
    .din1(ffc_551_p),
    .din2(g1919_n)
  );


  LA
  g_g1921_p
  (
    .dout(g1921_p),
    .din1(ffc_460_p_spl_010),
    .din2(ffc_536_p_spl_0)
  );


  LA
  g_g1922_p
  (
    .dout(g1922_p),
    .din1(ffc_457_p_spl_010),
    .din2(ffc_536_n_spl_0)
  );


  FA
  g_g1923_n
  (
    .dout(g1923_n),
    .din1(g1921_p),
    .din2(g1922_p)
  );


  LA
  g_g1924_p
  (
    .dout(g1924_p),
    .din1(ffc_551_n),
    .din2(g1923_n)
  );


  FA
  g_g1925_n
  (
    .dout(g1925_n),
    .din1(g1920_p),
    .din2(g1924_p)
  );


  LA
  g_g1926_p
  (
    .dout(g1926_p),
    .din1(ffc_466_n_spl_011),
    .din2(ffc_540_n_spl_0)
  );


  LA
  g_g1927_p
  (
    .dout(g1927_p),
    .din1(ffc_463_n_spl_010),
    .din2(ffc_540_p_spl_0)
  );


  FA
  g_g1928_n
  (
    .dout(g1928_n),
    .din1(g1926_p),
    .din2(g1927_p)
  );


  LA
  g_g1929_p
  (
    .dout(g1929_p),
    .din1(ffc_559_p),
    .din2(g1928_n)
  );


  LA
  g_g1930_p
  (
    .dout(g1930_p),
    .din1(ffc_460_p_spl_010),
    .din2(ffc_540_p_spl_)
  );


  LA
  g_g1931_p
  (
    .dout(g1931_p),
    .din1(ffc_457_p_spl_011),
    .din2(ffc_540_n_spl_)
  );


  FA
  g_g1932_n
  (
    .dout(g1932_n),
    .din1(g1930_p),
    .din2(g1931_p)
  );


  LA
  g_g1933_p
  (
    .dout(g1933_p),
    .din1(ffc_559_n),
    .din2(g1932_n)
  );


  FA
  g_g1934_n
  (
    .dout(g1934_n),
    .din1(g1929_p),
    .din2(g1933_p)
  );


  LA
  g_g1935_p
  (
    .dout(g1935_p),
    .din1(ffc_466_n_spl_011),
    .din2(ffc_598_n_spl_0)
  );


  LA
  g_g1936_p
  (
    .dout(g1936_p),
    .din1(ffc_463_n_spl_01),
    .din2(ffc_598_p_spl_0)
  );


  FA
  g_g1937_n
  (
    .dout(g1937_n),
    .din1(g1935_p),
    .din2(g1936_p)
  );


  LA
  g_g1938_p
  (
    .dout(g1938_p),
    .din1(ffc_616_p),
    .din2(g1937_n)
  );


  LA
  g_g1939_p
  (
    .dout(g1939_p),
    .din1(ffc_460_p_spl_01),
    .din2(ffc_598_p_spl_0)
  );


  LA
  g_g1940_p
  (
    .dout(g1940_p),
    .din1(ffc_457_p_spl_011),
    .din2(ffc_598_n_spl_0)
  );


  FA
  g_g1941_n
  (
    .dout(g1941_n),
    .din1(g1939_p),
    .din2(g1940_p)
  );


  LA
  g_g1942_p
  (
    .dout(g1942_p),
    .din1(ffc_616_n),
    .din2(g1941_n)
  );


  FA
  g_g1943_n
  (
    .dout(g1943_n),
    .din1(g1938_p),
    .din2(g1942_p)
  );


  LA
  g_g1944_p
  (
    .dout(g1944_p),
    .din1(ffc_466_n_spl_10),
    .din2(ffc_539_n_spl_0)
  );


  LA
  g_g1945_p
  (
    .dout(g1945_p),
    .din1(ffc_463_n_spl_10),
    .din2(ffc_539_p_spl_0)
  );


  FA
  g_g1946_n
  (
    .dout(g1946_n),
    .din1(g1944_p),
    .din2(g1945_p)
  );


  LA
  g_g1947_p
  (
    .dout(g1947_p),
    .din1(ffc_560_p),
    .din2(g1946_n)
  );


  LA
  g_g1948_p
  (
    .dout(g1948_p),
    .din1(ffc_460_p_spl_10),
    .din2(ffc_539_p_spl_)
  );


  LA
  g_g1949_p
  (
    .dout(g1949_p),
    .din1(ffc_457_p_spl_10),
    .din2(ffc_539_n_spl_)
  );


  FA
  g_g1950_n
  (
    .dout(g1950_n),
    .din1(g1948_p),
    .din2(g1949_p)
  );


  LA
  g_g1951_p
  (
    .dout(g1951_p),
    .din1(ffc_560_n),
    .din2(g1950_n)
  );


  FA
  g_g1952_n
  (
    .dout(g1952_n),
    .din1(g1947_p),
    .din2(g1951_p)
  );


  LA
  g_g1953_p
  (
    .dout(g1953_p),
    .din1(ffc_466_n_spl_10),
    .din2(ffc_526_n_spl_0)
  );


  LA
  g_g1954_p
  (
    .dout(g1954_p),
    .din1(ffc_463_n_spl_10),
    .din2(ffc_526_p_spl_0)
  );


  FA
  g_g1955_n
  (
    .dout(g1955_n),
    .din1(g1953_p),
    .din2(g1954_p)
  );


  LA
  g_g1956_p
  (
    .dout(g1956_p),
    .din1(ffc_544_p),
    .din2(g1955_n)
  );


  LA
  g_g1957_p
  (
    .dout(g1957_p),
    .din1(ffc_460_p_spl_10),
    .din2(ffc_526_p_spl_)
  );


  LA
  g_g1958_p
  (
    .dout(g1958_p),
    .din1(ffc_457_p_spl_10),
    .din2(ffc_526_n_spl_)
  );


  FA
  g_g1959_n
  (
    .dout(g1959_n),
    .din1(g1957_p),
    .din2(g1958_p)
  );


  LA
  g_g1960_p
  (
    .dout(g1960_p),
    .din1(ffc_544_n),
    .din2(g1959_n)
  );


  FA
  g_g1961_n
  (
    .dout(g1961_n),
    .din1(g1956_p),
    .din2(g1960_p)
  );


  LA
  g_g1962_p
  (
    .dout(g1962_p),
    .din1(ffc_466_n_spl_11),
    .din2(ffc_557_n_spl_0)
  );


  LA
  g_g1963_p
  (
    .dout(g1963_p),
    .din1(ffc_463_n_spl_11),
    .din2(ffc_557_p_spl_0)
  );


  FA
  g_g1964_n
  (
    .dout(g1964_n),
    .din1(g1962_p),
    .din2(g1963_p)
  );


  LA
  g_g1965_p
  (
    .dout(g1965_p),
    .din1(ffc_582_p),
    .din2(g1964_n)
  );


  LA
  g_g1966_p
  (
    .dout(g1966_p),
    .din1(ffc_460_p_spl_11),
    .din2(ffc_557_p_spl_0)
  );


  LA
  g_g1967_p
  (
    .dout(g1967_p),
    .din1(ffc_457_p_spl_11),
    .din2(ffc_557_n_spl_0)
  );


  FA
  g_g1968_n
  (
    .dout(g1968_n),
    .din1(g1966_p),
    .din2(g1967_p)
  );


  LA
  g_g1969_p
  (
    .dout(g1969_p),
    .din1(ffc_582_n),
    .din2(g1968_n)
  );


  FA
  g_g1970_n
  (
    .dout(g1970_n),
    .din1(g1965_p),
    .din2(g1969_p)
  );


  LA
  g_g1971_p
  (
    .dout(g1971_p),
    .din1(ffc_466_n_spl_11),
    .din2(ffc_549_n_spl_0)
  );


  LA
  g_g1972_p
  (
    .dout(g1972_p),
    .din1(ffc_463_n_spl_11),
    .din2(ffc_549_p_spl_0)
  );


  FA
  g_g1973_n
  (
    .dout(g1973_n),
    .din1(g1971_p),
    .din2(g1972_p)
  );


  LA
  g_g1974_p
  (
    .dout(g1974_p),
    .din1(ffc_573_p),
    .din2(g1973_n)
  );


  LA
  g_g1975_p
  (
    .dout(g1975_p),
    .din1(ffc_460_p_spl_11),
    .din2(ffc_549_p_spl_0)
  );


  LA
  g_g1976_p
  (
    .dout(g1976_p),
    .din1(ffc_457_p_spl_11),
    .din2(ffc_549_n_spl_0)
  );


  FA
  g_g1977_n
  (
    .dout(g1977_n),
    .din1(g1975_p),
    .din2(g1976_p)
  );


  LA
  g_g1978_p
  (
    .dout(g1978_p),
    .din1(ffc_573_n),
    .din2(g1977_n)
  );


  FA
  g_g1979_n
  (
    .dout(g1979_n),
    .din1(g1974_p),
    .din2(g1978_p)
  );


  LA
  g_g1980_p
  (
    .dout(g1980_p),
    .din1(ffc_785_n_spl_),
    .din2(ffc_786_p_spl_)
  );


  FA
  g_g1980_n
  (
    .dout(g1980_n),
    .din1(ffc_785_p_spl_),
    .din2(ffc_786_n_spl_)
  );


  LA
  g_g1981_p
  (
    .dout(g1981_p),
    .din1(ffc_785_p_spl_),
    .din2(ffc_786_n_spl_)
  );


  FA
  g_g1981_n
  (
    .dout(g1981_n),
    .din1(ffc_785_n_spl_),
    .din2(ffc_786_p_spl_)
  );


  LA
  g_g1982_p
  (
    .dout(g1982_p),
    .din1(g1980_n),
    .din2(g1981_n)
  );


  FA
  g_g1982_n
  (
    .dout(g1982_n),
    .din1(g1980_p),
    .din2(g1981_p)
  );


  LA
  g_g1983_p
  (
    .dout(g1983_p),
    .din1(ffc_789_n_spl_),
    .din2(ffc_790_n_spl_0)
  );


  FA
  g_g1983_n
  (
    .dout(g1983_n),
    .din1(ffc_789_p_spl_),
    .din2(ffc_790_p_spl_0)
  );


  LA
  g_g1984_p
  (
    .dout(g1984_p),
    .din1(ffc_789_p_spl_),
    .din2(ffc_790_p_spl_0)
  );


  FA
  g_g1984_n
  (
    .dout(g1984_n),
    .din1(ffc_789_n_spl_),
    .din2(ffc_790_n_spl_)
  );


  LA
  g_g1985_p
  (
    .dout(g1985_p),
    .din1(g1983_n),
    .din2(g1984_n)
  );


  FA
  g_g1985_n
  (
    .dout(g1985_n),
    .din1(g1983_p),
    .din2(g1984_p)
  );


  LA
  g_g1986_p
  (
    .dout(g1986_p),
    .din1(g1982_n_spl_),
    .din2(g1985_p_spl_)
  );


  FA
  g_g1986_n
  (
    .dout(g1986_n),
    .din1(g1982_p_spl_),
    .din2(g1985_n_spl_)
  );


  LA
  g_g1987_p
  (
    .dout(g1987_p),
    .din1(g1982_p_spl_),
    .din2(g1985_n_spl_)
  );


  FA
  g_g1987_n
  (
    .dout(g1987_n),
    .din1(g1982_n_spl_),
    .din2(g1985_p_spl_)
  );


  LA
  g_g1988_p
  (
    .dout(g1988_p),
    .din1(g1986_n),
    .din2(g1987_n)
  );


  FA
  g_g1988_n
  (
    .dout(g1988_n),
    .din1(g1986_p),
    .din2(g1987_p)
  );


  LA
  g_g1989_p
  (
    .dout(g1989_p),
    .din1(ffc_784_n_spl_),
    .din2(ffc_788_p_spl_)
  );


  FA
  g_g1989_n
  (
    .dout(g1989_n),
    .din1(ffc_784_p_spl_),
    .din2(ffc_788_n_spl_)
  );


  LA
  g_g1990_p
  (
    .dout(g1990_p),
    .din1(ffc_784_p_spl_),
    .din2(ffc_788_n_spl_)
  );


  FA
  g_g1990_n
  (
    .dout(g1990_n),
    .din1(ffc_784_n_spl_),
    .din2(ffc_788_p_spl_)
  );


  LA
  g_g1991_p
  (
    .dout(g1991_p),
    .din1(g1989_n),
    .din2(g1990_n)
  );


  FA
  g_g1991_n
  (
    .dout(g1991_n),
    .din1(g1989_p),
    .din2(g1990_p)
  );


  LA
  g_g1992_p
  (
    .dout(g1992_p),
    .din1(ffc_787_n_spl_),
    .din2(ffc_810_n_spl_)
  );


  FA
  g_g1992_n
  (
    .dout(g1992_n),
    .din1(ffc_787_p_spl_),
    .din2(ffc_810_p_spl_)
  );


  LA
  g_g1993_p
  (
    .dout(g1993_p),
    .din1(ffc_787_p_spl_),
    .din2(ffc_810_p_spl_)
  );


  FA
  g_g1993_n
  (
    .dout(g1993_n),
    .din1(ffc_787_n_spl_),
    .din2(ffc_810_n_spl_)
  );


  LA
  g_g1994_p
  (
    .dout(g1994_p),
    .din1(g1992_n),
    .din2(g1993_n)
  );


  FA
  g_g1994_n
  (
    .dout(g1994_n),
    .din1(g1992_p),
    .din2(g1993_p)
  );


  LA
  g_g1995_p
  (
    .dout(g1995_p),
    .din1(g1991_p_spl_),
    .din2(g1994_n_spl_)
  );


  FA
  g_g1995_n
  (
    .dout(g1995_n),
    .din1(g1991_n_spl_),
    .din2(g1994_p_spl_)
  );


  LA
  g_g1996_p
  (
    .dout(g1996_p),
    .din1(g1991_n_spl_),
    .din2(g1994_p_spl_)
  );


  FA
  g_g1996_n
  (
    .dout(g1996_n),
    .din1(g1991_p_spl_),
    .din2(g1994_n_spl_)
  );


  LA
  g_g1997_p
  (
    .dout(g1997_p),
    .din1(g1995_n),
    .din2(g1996_n)
  );


  FA
  g_g1997_n
  (
    .dout(g1997_n),
    .din1(g1995_p),
    .din2(g1996_p)
  );


  FA
  g_g1998_n
  (
    .dout(g1998_n),
    .din1(g1988_p),
    .din2(g1997_n)
  );


  FA
  g_g1999_n
  (
    .dout(g1999_n),
    .din1(g1988_n),
    .din2(g1997_p)
  );


  LA
  g_g2000_p
  (
    .dout(g2000_p),
    .din1(ffc_493_p_spl_0),
    .din2(g1999_n)
  );


  LA
  g_g2001_p
  (
    .dout(g2001_p),
    .din1(g1998_n),
    .din2(g2000_p)
  );


  LA
  g_g2002_p
  (
    .dout(g2002_p),
    .din1(ffc_547_n),
    .din2(ffc_619_p)
  );


  LA
  g_g2003_p
  (
    .dout(g2003_p),
    .din1(ffc_547_p),
    .din2(ffc_619_n)
  );


  FA
  g_g2004_n
  (
    .dout(g2004_n),
    .din1(g2002_p),
    .din2(g2003_p)
  );


  FA
  g_g2005_n
  (
    .dout(g2005_n),
    .din1(ffc_553_n),
    .din2(g1872_p_spl_00)
  );


  FA
  g_g2006_n
  (
    .dout(g2006_n),
    .din1(ffc_552_p),
    .din2(g1872_n_spl_00)
  );


  LA
  g_g2007_p
  (
    .dout(g2007_p),
    .din1(g2005_n),
    .din2(g2006_n)
  );


  LA
  g_g2008_p
  (
    .dout(g2008_p),
    .din1(ffc_562_n),
    .din2(g1895_n_spl_)
  );


  FA
  g_g2008_n
  (
    .dout(g2008_n),
    .din1(ffc_562_p),
    .din2(g1895_p)
  );


  FA
  g_g2009_n
  (
    .dout(g2009_n),
    .din1(ffc_566_p),
    .din2(g2008_n)
  );


  FA
  g_g2010_n
  (
    .dout(g2010_n),
    .din1(ffc_566_n),
    .din2(g2008_p)
  );


  LA
  g_g2011_p
  (
    .dout(g2011_p),
    .din1(g2009_n),
    .din2(g2010_n)
  );


  LA
  g_g2012_p
  (
    .dout(g2012_p),
    .din1(ffc_350_p_spl_0),
    .din2(ffc_529_p_spl_)
  );


  FA
  g_g2012_n
  (
    .dout(g2012_n),
    .din1(ffc_350_n_spl_0),
    .din2(ffc_529_n_spl_)
  );


  LA
  g_g2013_p
  (
    .dout(g2013_p),
    .din1(ffc_353_p),
    .din2(ffc_529_n_spl_)
  );


  FA
  g_g2013_n
  (
    .dout(g2013_n),
    .din1(ffc_353_n),
    .din2(ffc_529_p_spl_)
  );


  LA
  g_g2014_p
  (
    .dout(g2014_p),
    .din1(g2012_n),
    .din2(g2013_n)
  );


  FA
  g_g2014_n
  (
    .dout(g2014_n),
    .din1(g2012_p),
    .din2(g2013_p)
  );


  FA
  g_g2015_n
  (
    .dout(g2015_n),
    .din1(ffc_595_p),
    .din2(g2014_n)
  );


  FA
  g_g2016_n
  (
    .dout(g2016_n),
    .din1(ffc_595_n),
    .din2(g2014_p)
  );


  LA
  g_g2017_p
  (
    .dout(g2017_p),
    .din1(g2015_n),
    .din2(g2016_n)
  );


  LA
  g_g2018_p
  (
    .dout(g2018_p),
    .din1(ffc_597_p),
    .din2(g1872_n_spl_0)
  );


  LA
  g_g2019_p
  (
    .dout(g2019_p),
    .din1(ffc_608_p_spl_),
    .din2(g1872_p_spl_0)
  );


  FA
  g_g2020_n
  (
    .dout(g2020_n),
    .din1(g2018_p),
    .din2(g2019_p)
  );


  FA
  g_g2021_n
  (
    .dout(g2021_n),
    .din1(ffc_604_n_spl_),
    .din2(ffc_625_n)
  );


  FA
  g_g2022_n
  (
    .dout(g2022_n),
    .din1(ffc_604_p_spl_),
    .din2(ffc_625_p)
  );


  LA
  g_g2023_p
  (
    .dout(g2023_p),
    .din1(g2021_n),
    .din2(g2022_n)
  );


  LA
  g_g2024_p
  (
    .dout(g2024_p),
    .din1(ffc_613_p),
    .din2(g1872_n_spl_1)
  );


  FA
  g_g2024_n
  (
    .dout(g2024_n),
    .din1(ffc_613_n),
    .din2(g1872_p_spl_1)
  );


  LA
  g_g2025_p
  (
    .dout(g2025_p),
    .din1(ffc_612_p),
    .din2(g1872_p_spl_1)
  );


  FA
  g_g2025_n
  (
    .dout(g2025_n),
    .din1(ffc_612_n),
    .din2(g1872_n_spl_1)
  );


  LA
  g_g2026_p
  (
    .dout(g2026_p),
    .din1(g2024_n),
    .din2(g2025_n)
  );


  FA
  g_g2026_n
  (
    .dout(g2026_n),
    .din1(g2024_p),
    .din2(g2025_p)
  );


  LA
  g_g2027_p
  (
    .dout(g2027_p),
    .din1(ffc_614_p_spl_),
    .din2(g2026_p)
  );


  LA
  g_g2028_p
  (
    .dout(g2028_p),
    .din1(ffc_614_n),
    .din2(g2026_n)
  );


  FA
  g_g2029_n
  (
    .dout(g2029_n),
    .din1(g2027_p),
    .din2(g2028_p)
  );


  LA
  g_g2030_p
  (
    .dout(g2030_p),
    .din1(ffc_624_n_spl_),
    .din2(ffc_659_p_spl_)
  );


  LA
  g_g2031_p
  (
    .dout(g2031_p),
    .din1(ffc_624_p),
    .din2(ffc_659_n_spl_)
  );


  FA
  g_g2032_n
  (
    .dout(g2032_n),
    .din1(g2030_p),
    .din2(g2031_p)
  );


  LA
  g_g2033_p
  (
    .dout(g2033_p),
    .din1(ffc_537_p),
    .din2(ffc_541_n)
  );


  LA
  g_g2034_p
  (
    .dout(g2034_p),
    .din1(ffc_537_n),
    .din2(ffc_541_p)
  );


  FA
  g_g2035_n
  (
    .dout(g2035_n),
    .din1(g2033_p),
    .din2(g2034_p)
  );


  FA
  g_g2036_n
  (
    .dout(g2036_n),
    .din1(ffc_589_p),
    .din2(ffc_640_n)
  );


  FA
  g_g2037_n
  (
    .dout(g2037_n),
    .din1(ffc_589_n),
    .din2(ffc_640_p_spl_)
  );


  LA
  g_g2038_p
  (
    .dout(g2038_p),
    .din1(g2036_n),
    .din2(g2037_n)
  );


  LA
  g_g2039_p
  (
    .dout(g2039_p),
    .din1(g2035_n_spl_),
    .din2(g2038_p_spl_)
  );


  FA
  g_g2040_n
  (
    .dout(g2040_n),
    .din1(g2035_n_spl_),
    .din2(g2038_p_spl_)
  );


  LA
  g_g2041_p
  (
    .dout(g2041_p),
    .din1(ffc_375_n_spl_),
    .din2(ffc_571_p_spl_)
  );


  FA
  g_g2041_n
  (
    .dout(g2041_n),
    .din1(ffc_375_p_spl_0),
    .din2(ffc_571_n_spl_)
  );


  LA
  g_g2042_p
  (
    .dout(g2042_p),
    .din1(ffc_375_p_spl_),
    .din2(ffc_571_n_spl_)
  );


  FA
  g_g2042_n
  (
    .dout(g2042_n),
    .din1(ffc_375_n_spl_),
    .din2(ffc_571_p_spl_)
  );


  LA
  g_g2043_p
  (
    .dout(g2043_p),
    .din1(g2041_n),
    .din2(g2042_n)
  );


  FA
  g_g2043_n
  (
    .dout(g2043_n),
    .din1(g2041_p),
    .din2(g2042_p)
  );


  LA
  g_g2044_p
  (
    .dout(g2044_p),
    .din1(ffc_590_p_spl_),
    .din2(g2043_p)
  );


  LA
  g_g2045_p
  (
    .dout(g2045_p),
    .din1(ffc_590_n_spl_),
    .din2(g2043_n)
  );


  FA
  g_g2046_n
  (
    .dout(g2046_n),
    .din1(g2044_p),
    .din2(g2045_p)
  );


  FA
  g_g2047_n
  (
    .dout(g2047_n),
    .din1(ffc_549_p_spl_),
    .din2(ffc_557_n_spl_)
  );


  FA
  g_g2048_n
  (
    .dout(g2048_n),
    .din1(ffc_549_n_spl_),
    .din2(ffc_557_p_spl_)
  );


  LA
  g_g2049_p
  (
    .dout(g2049_p),
    .din1(g2047_n),
    .din2(g2048_n)
  );


  LA
  g_g2050_p
  (
    .dout(g2050_p),
    .din1(g2046_n_spl_),
    .din2(g2049_p_spl_)
  );


  FA
  g_g2051_n
  (
    .dout(g2051_n),
    .din1(g2046_n_spl_),
    .din2(g2049_p_spl_)
  );


  LA
  g_g2052_p
  (
    .dout(g2052_p),
    .din1(ffc_583_n),
    .din2(ffc_611_p)
  );


  LA
  g_g2053_p
  (
    .dout(g2053_p),
    .din1(ffc_583_p),
    .din2(ffc_611_n)
  );


  FA
  g_g2054_n
  (
    .dout(g2054_n),
    .din1(g2052_p),
    .din2(g2053_p)
  );


  LA
  g_g2055_p
  (
    .dout(g2055_p),
    .din1(ffc_577_n),
    .din2(ffc_586_p)
  );


  LA
  g_g2056_p
  (
    .dout(g2056_p),
    .din1(ffc_577_p),
    .din2(ffc_586_n)
  );


  FA
  g_g2057_n
  (
    .dout(g2057_n),
    .din1(g2055_p),
    .din2(g2056_p)
  );


  FA
  g_g2058_n
  (
    .dout(g2058_n),
    .din1(g2054_n_spl_),
    .din2(g2057_n_spl_)
  );


  LA
  g_g2059_p
  (
    .dout(g2059_p),
    .din1(g2054_n_spl_),
    .din2(g2057_n_spl_)
  );


  LA
  g_g2060_p
  (
    .dout(g2060_p),
    .din1(ffc_556_n_spl_1),
    .din2(ffc_598_p_spl_1)
  );


  FA
  g_g2060_n
  (
    .dout(g2060_n),
    .din1(ffc_556_p_spl_1),
    .din2(ffc_598_n_spl_1)
  );


  LA
  g_g2061_p
  (
    .dout(g2061_p),
    .din1(ffc_556_p_spl_1),
    .din2(ffc_598_n_spl_1)
  );


  FA
  g_g2061_n
  (
    .dout(g2061_n),
    .din1(ffc_556_n_spl_1),
    .din2(ffc_598_p_spl_1)
  );


  LA
  g_g2062_p
  (
    .dout(g2062_p),
    .din1(g2060_n),
    .din2(g2061_n)
  );


  FA
  g_g2062_n
  (
    .dout(g2062_n),
    .din1(g2060_p),
    .din2(g2061_p)
  );


  LA
  g_g2063_p
  (
    .dout(g2063_p),
    .din1(ffc_350_n_spl_0),
    .din2(ffc_536_p_spl_1)
  );


  FA
  g_g2063_n
  (
    .dout(g2063_n),
    .din1(ffc_350_p_spl_0),
    .din2(ffc_536_n_spl_1)
  );


  LA
  g_g2064_p
  (
    .dout(g2064_p),
    .din1(ffc_350_p_spl_),
    .din2(ffc_536_n_spl_1)
  );


  FA
  g_g2064_n
  (
    .dout(g2064_n),
    .din1(ffc_350_n_spl_),
    .din2(ffc_536_p_spl_1)
  );


  LA
  g_g2065_p
  (
    .dout(g2065_p),
    .din1(g2063_n),
    .din2(g2064_n)
  );


  FA
  g_g2065_n
  (
    .dout(g2065_n),
    .din1(g2063_p),
    .din2(g2064_p)
  );


  FA
  g_g2066_n
  (
    .dout(g2066_n),
    .din1(g2062_n),
    .din2(g2065_n)
  );


  FA
  g_g2067_n
  (
    .dout(g2067_n),
    .din1(g2062_p),
    .din2(g2065_p)
  );


  LA
  g_g2068_p
  (
    .dout(g2068_p),
    .din1(g2066_n),
    .din2(g2067_n)
  );


  LA
  g_g2069_p
  (
    .dout(g2069_p),
    .din1(ffc_773_p),
    .din2(ffc_774_n)
  );


  FA
  g_g2069_n
  (
    .dout(g2069_n),
    .din1(ffc_773_n),
    .din2(ffc_774_p)
  );


  LA
  g_g2070_p
  (
    .dout(g2070_p),
    .din1(ffc_642_n),
    .din2(ffc_658_p)
  );


  FA
  g_g2070_n
  (
    .dout(g2070_n),
    .din1(ffc_642_p),
    .din2(ffc_658_n)
  );


  LA
  g_g2071_p
  (
    .dout(g2071_p),
    .din1(g2069_p_spl_),
    .din2(g2070_n_spl_)
  );


  FA
  g_g2071_n
  (
    .dout(g2071_n),
    .din1(g2069_n_spl_),
    .din2(g2070_p_spl_)
  );


  LA
  g_g2072_p
  (
    .dout(g2072_p),
    .din1(g2069_n_spl_),
    .din2(g2070_p_spl_)
  );


  FA
  g_g2072_n
  (
    .dout(g2072_n),
    .din1(g2069_p_spl_),
    .din2(g2070_n_spl_)
  );


  LA
  g_g2073_p
  (
    .dout(g2073_p),
    .din1(g2071_n),
    .din2(g2072_n)
  );


  FA
  g_g2073_n
  (
    .dout(g2073_n),
    .din1(g2071_p),
    .din2(g2072_p)
  );


  LA
  g_g2074_p
  (
    .dout(g2074_p),
    .din1(ffc_424_n_spl_0),
    .din2(g2073_n)
  );


  FA
  g_g2074_n
  (
    .dout(g2074_n),
    .din1(ffc_424_p_spl_0),
    .din2(g2073_p)
  );


  LA
  g_g2075_p
  (
    .dout(g2075_p),
    .din1(ffc_792_n),
    .din2(ffc_793_p)
  );


  FA
  g_g2075_n
  (
    .dout(g2075_n),
    .din1(ffc_792_p),
    .din2(ffc_793_n)
  );


  LA
  g_g2076_p
  (
    .dout(g2076_p),
    .din1(ffc_797_p),
    .din2(ffc_798_n)
  );


  FA
  g_g2076_n
  (
    .dout(g2076_n),
    .din1(ffc_797_n),
    .din2(ffc_798_p)
  );


  LA
  g_g2077_p
  (
    .dout(g2077_p),
    .din1(g2075_p_spl_),
    .din2(g2076_p_spl_)
  );


  FA
  g_g2077_n
  (
    .dout(g2077_n),
    .din1(g2075_n_spl_),
    .din2(g2076_n_spl_)
  );


  LA
  g_g2078_p
  (
    .dout(g2078_p),
    .din1(g2075_n_spl_),
    .din2(g2076_n_spl_)
  );


  FA
  g_g2078_n
  (
    .dout(g2078_n),
    .din1(g2075_p_spl_),
    .din2(g2076_p_spl_)
  );


  LA
  g_g2079_p
  (
    .dout(g2079_p),
    .din1(g2077_n),
    .din2(g2078_n)
  );


  FA
  g_g2079_n
  (
    .dout(g2079_n),
    .din1(g2077_p),
    .din2(g2078_p)
  );


  LA
  g_g2080_p
  (
    .dout(g2080_p),
    .din1(ffc_424_p_spl_0),
    .din2(g2079_p)
  );


  FA
  g_g2080_n
  (
    .dout(g2080_n),
    .din1(ffc_424_n_spl_0),
    .din2(g2079_n)
  );


  LA
  g_g2081_p
  (
    .dout(g2081_p),
    .din1(g2074_n),
    .din2(g2080_n)
  );


  FA
  g_g2081_n
  (
    .dout(g2081_n),
    .din1(g2074_p),
    .din2(g2080_p)
  );


  LA
  g_g2082_p
  (
    .dout(g2082_p),
    .din1(ffc_776_n),
    .din2(ffc_777_p)
  );


  FA
  g_g2082_n
  (
    .dout(g2082_n),
    .din1(ffc_776_p),
    .din2(ffc_777_n)
  );


  LA
  g_g2083_p
  (
    .dout(g2083_p),
    .din1(ffc_771_n_spl_0),
    .din2(ffc_772_n_spl_0)
  );


  FA
  g_g2083_n
  (
    .dout(g2083_n),
    .din1(ffc_771_p_spl_00),
    .din2(ffc_772_p_spl_0)
  );


  LA
  g_g2084_p
  (
    .dout(g2084_p),
    .din1(g2082_n_spl_),
    .din2(g2083_n)
  );


  FA
  g_g2084_n
  (
    .dout(g2084_n),
    .din1(g2082_p_spl_),
    .din2(g2083_p)
  );


  LA
  g_g2085_p
  (
    .dout(g2085_p),
    .din1(ffc_771_n_spl_1),
    .din2(ffc_809_n)
  );


  FA
  g_g2085_n
  (
    .dout(g2085_n),
    .din1(ffc_771_p_spl_0),
    .din2(ffc_809_p)
  );


  LA
  g_g2086_p
  (
    .dout(g2086_p),
    .din1(ffc_772_n_spl_),
    .din2(g2085_p_spl_)
  );


  FA
  g_g2086_n
  (
    .dout(g2086_n),
    .din1(ffc_772_p_spl_1),
    .din2(g2085_n_spl_)
  );


  LA
  g_g2087_p
  (
    .dout(g2087_p),
    .din1(g2084_n),
    .din2(g2086_n)
  );


  FA
  g_g2087_n
  (
    .dout(g2087_n),
    .din1(g2084_p),
    .din2(g2086_p)
  );


  LA
  g_g2088_p
  (
    .dout(g2088_p),
    .din1(ffc_424_p_spl_1),
    .din2(g2087_n)
  );


  FA
  g_g2088_n
  (
    .dout(g2088_n),
    .din1(ffc_424_n_spl_1),
    .din2(g2087_p)
  );


  LA
  g_g2089_p
  (
    .dout(g2089_p),
    .din1(ffc_771_p_spl_1),
    .din2(g2082_n_spl_)
  );


  FA
  g_g2089_n
  (
    .dout(g2089_n),
    .din1(ffc_771_n_spl_1),
    .din2(g2082_p_spl_)
  );


  LA
  g_g2090_p
  (
    .dout(g2090_p),
    .din1(g2085_n_spl_),
    .din2(g2089_n)
  );


  FA
  g_g2090_n
  (
    .dout(g2090_n),
    .din1(g2085_p_spl_),
    .din2(g2089_p)
  );


  LA
  g_g2091_p
  (
    .dout(g2091_p),
    .din1(ffc_424_n_spl_1),
    .din2(g2090_n)
  );


  FA
  g_g2091_n
  (
    .dout(g2091_n),
    .din1(ffc_424_p_spl_1),
    .din2(g2090_p)
  );


  LA
  g_g2092_p
  (
    .dout(g2092_p),
    .din1(g2088_n),
    .din2(g2091_n)
  );


  FA
  g_g2092_n
  (
    .dout(g2092_n),
    .din1(g2088_p),
    .din2(g2091_p)
  );


  FA
  g_g2093_n
  (
    .dout(g2093_n),
    .din1(g2081_p),
    .din2(g2092_n)
  );


  FA
  g_g2094_n
  (
    .dout(g2094_n),
    .din1(g2081_n),
    .din2(g2092_p)
  );


  LA
  g_g2095_p
  (
    .dout(g2095_p),
    .din1(g2093_n),
    .din2(g2094_n)
  );


  FA
  g_g2096_n
  (
    .dout(g2096_n),
    .din1(ffc_848_p_spl_0),
    .din2(g1761_n_spl_0)
  );


  LA
  g_g2097_p
  (
    .dout(g2097_p),
    .din1(g1793_p_spl_),
    .din2(g1796_p_spl_0)
  );


  FA
  g_g2098_n
  (
    .dout(g2098_n),
    .din1(g1794_p),
    .din2(g2097_p)
  );


  LA
  g_g2099_p
  (
    .dout(g2099_p),
    .din1(g1762_p_spl_),
    .din2(g1799_p_spl_0)
  );


  LA
  g_g2100_p
  (
    .dout(g2100_p),
    .din1(ffc_628_n_spl_),
    .din2(ffc_832_n_spl_000)
  );


  LA
  g_g2101_p
  (
    .dout(g2101_p),
    .din1(ffc_628_p_spl_0),
    .din2(ffc_833_n_spl_000)
  );


  FA
  g_g2102_n
  (
    .dout(g2102_n),
    .din1(g2100_p),
    .din2(g2101_p)
  );


  LA
  g_g2103_p
  (
    .dout(g2103_p),
    .din1(ffc_651_p),
    .din2(g2102_n)
  );


  LA
  g_g2104_p
  (
    .dout(g2104_p),
    .din1(ffc_628_p_spl_0),
    .din2(ffc_834_p_spl_000)
  );


  LA
  g_g2105_p
  (
    .dout(g2105_p),
    .din1(ffc_628_n_spl_),
    .din2(ffc_831_p_spl_000)
  );


  FA
  g_g2106_n
  (
    .dout(g2106_n),
    .din1(g2104_p),
    .din2(g2105_p)
  );


  LA
  g_g2107_p
  (
    .dout(g2107_p),
    .din1(ffc_651_n),
    .din2(g2106_n)
  );


  FA
  g_g2108_n
  (
    .dout(g2108_n),
    .din1(g2103_p),
    .din2(g2107_p)
  );


  LA
  g_g2109_p
  (
    .dout(g2109_p),
    .din1(ffc_633_n_spl_),
    .din2(ffc_832_n_spl_000)
  );


  LA
  g_g2110_p
  (
    .dout(g2110_p),
    .din1(ffc_633_p_spl_0),
    .din2(ffc_833_n_spl_000)
  );


  FA
  g_g2111_n
  (
    .dout(g2111_n),
    .din1(g2109_p),
    .din2(g2110_p)
  );


  LA
  g_g2112_p
  (
    .dout(g2112_p),
    .din1(ffc_665_p),
    .din2(g2111_n)
  );


  LA
  g_g2113_p
  (
    .dout(g2113_p),
    .din1(ffc_633_p_spl_0),
    .din2(ffc_834_p_spl_000)
  );


  LA
  g_g2114_p
  (
    .dout(g2114_p),
    .din1(ffc_633_n_spl_),
    .din2(ffc_831_p_spl_000)
  );


  FA
  g_g2115_n
  (
    .dout(g2115_n),
    .din1(g2113_p),
    .din2(g2114_p)
  );


  LA
  g_g2116_p
  (
    .dout(g2116_p),
    .din1(ffc_665_n),
    .din2(g2115_n)
  );


  FA
  g_g2117_n
  (
    .dout(g2117_n),
    .din1(g2112_p),
    .din2(g2116_p)
  );


  LA
  g_g2118_p
  (
    .dout(g2118_p),
    .din1(ffc_677_n),
    .din2(ffc_832_n_spl_001)
  );


  LA
  g_g2119_p
  (
    .dout(g2119_p),
    .din1(ffc_677_p_spl_),
    .din2(ffc_833_n_spl_001)
  );


  FA
  g_g2120_n
  (
    .dout(g2120_n),
    .din1(g2118_p),
    .din2(g2119_p)
  );


  LA
  g_g2121_p
  (
    .dout(g2121_p),
    .din1(ffc_780_n),
    .din2(ffc_832_n_spl_001)
  );


  LA
  g_g2122_p
  (
    .dout(g2122_p),
    .din1(ffc_780_p_spl_),
    .din2(ffc_833_n_spl_001)
  );


  FA
  g_g2123_n
  (
    .dout(g2123_n),
    .din1(g2121_p),
    .din2(g2122_p)
  );


  FA
  g_g2124_n
  (
    .dout(g2124_n),
    .din1(ffc_355_p_spl_0),
    .din2(ffc_831_p_spl_001)
  );


  FA
  g_g2125_n
  (
    .dout(g2125_n),
    .din1(ffc_355_n),
    .din2(ffc_834_p_spl_001)
  );


  LA
  g_g2126_p
  (
    .dout(g2126_p),
    .din1(g2124_n),
    .din2(g2125_n)
  );


  LA
  g_g2127_p
  (
    .dout(g2127_p),
    .din1(ffc_346_p_spl_),
    .din2(ffc_839_p_spl_10)
  );


  FA
  g_g2127_n
  (
    .dout(g2127_n),
    .din1(ffc_346_n),
    .din2(ffc_839_n_spl_10)
  );


  LA
  g_g2128_p
  (
    .dout(g2128_p),
    .din1(ffc_347_p),
    .din2(ffc_839_n_spl_11)
  );


  FA
  g_g2128_n
  (
    .dout(g2128_n),
    .din1(ffc_347_n),
    .din2(ffc_839_p_spl_10)
  );


  LA
  g_g2129_p
  (
    .dout(g2129_p),
    .din1(g2127_n),
    .din2(g2128_n)
  );


  FA
  g_g2129_n
  (
    .dout(g2129_n),
    .din1(g2127_p),
    .din2(g2128_p)
  );


  LA
  g_g2130_p
  (
    .dout(g2130_p),
    .din1(ffc_366_p_spl_),
    .din2(ffc_863_p_spl_011)
  );


  FA
  g_g2130_n
  (
    .dout(g2130_n),
    .din1(ffc_366_n),
    .din2(ffc_863_n_spl_01)
  );


  LA
  g_g2131_p
  (
    .dout(g2131_p),
    .din1(ffc_367_p_spl_),
    .din2(ffc_863_n_spl_10)
  );


  FA
  g_g2131_n
  (
    .dout(g2131_n),
    .din1(ffc_367_n),
    .din2(ffc_863_p_spl_011)
  );


  LA
  g_g2132_p
  (
    .dout(g2132_p),
    .din1(g2130_n),
    .din2(g2131_n)
  );


  FA
  g_g2132_n
  (
    .dout(g2132_n),
    .din1(g2130_p),
    .din2(g2131_p)
  );


  FA
  g_g2133_n
  (
    .dout(g2133_n),
    .din1(ffc_397_n),
    .din2(g1802_p)
  );


  FA
  g_g2134_n
  (
    .dout(g2134_n),
    .din1(ffc_388_p_spl_0),
    .din2(g1780_n_spl_0)
  );


  LA
  g_g2135_p
  (
    .dout(g2135_p),
    .din1(g1803_n),
    .din2(g2134_n)
  );


  FA
  g_g2136_n
  (
    .dout(g2136_n),
    .din1(ffc_392_p_spl_0),
    .din2(g1777_n_spl_0)
  );


  LA
  g_g2137_p
  (
    .dout(g2137_p),
    .din1(g1804_n),
    .din2(g2136_n)
  );


  LA
  g_g2138_p
  (
    .dout(g2138_p),
    .din1(ffc_826_p_spl_0),
    .din2(ffc_844_p_spl_1)
  );


  FA
  g_g2138_n
  (
    .dout(g2138_n),
    .din1(ffc_826_n_spl_0),
    .din2(ffc_844_n_spl_)
  );


  LA
  g_g2139_p
  (
    .dout(g2139_p),
    .din1(ffc_812_n),
    .din2(g2138_n)
  );


  FA
  g_g2139_n
  (
    .dout(g2139_n),
    .din1(ffc_812_p_spl_),
    .din2(g2138_p)
  );


  LA
  g_g2140_p
  (
    .dout(g2140_p),
    .din1(g1758_p_spl_0),
    .din2(g2139_n_spl_0)
  );


  FA
  g_g2141_n
  (
    .dout(g2141_n),
    .din1(g1756_p_spl_),
    .din2(g2140_p)
  );


  FA
  g_g2142_n
  (
    .dout(g2142_n),
    .din1(ffc_825_n_spl_0),
    .din2(g1725_n_spl_)
  );


  FA
  g_g2143_n
  (
    .dout(g2143_n),
    .din1(g1758_n_spl_0),
    .din2(g2142_n_spl_)
  );


  LA
  g_g2144_p
  (
    .dout(g2144_p),
    .din1(ffc_671_n_spl_),
    .din2(ffc_826_p_spl_0)
  );


  FA
  g_g2144_n
  (
    .dout(g2144_n),
    .din1(ffc_671_p_spl_0),
    .din2(ffc_826_n_spl_0)
  );


  LA
  g_g2145_p
  (
    .dout(g2145_p),
    .din1(ffc_671_p_spl_0),
    .din2(ffc_826_n_spl_1)
  );


  FA
  g_g2145_n
  (
    .dout(g2145_n),
    .din1(ffc_671_n_spl_),
    .din2(ffc_826_p_spl_1)
  );


  LA
  g_g2146_p
  (
    .dout(g2146_p),
    .din1(g2144_n),
    .din2(g2145_n)
  );


  FA
  g_g2146_n
  (
    .dout(g2146_n),
    .din1(g2144_p),
    .din2(g2145_p)
  );


  LA
  g_g2147_p
  (
    .dout(g2147_p),
    .din1(ffc_756_n_spl_0),
    .din2(g2146_p_spl_)
  );


  FA
  g_g2147_n
  (
    .dout(g2147_n),
    .din1(ffc_756_p_spl_0),
    .din2(g2146_n_spl_)
  );


  LA
  g_g2148_p
  (
    .dout(g2148_p),
    .din1(ffc_756_p_spl_0),
    .din2(g2146_n_spl_)
  );


  FA
  g_g2148_n
  (
    .dout(g2148_n),
    .din1(ffc_756_n_spl_0),
    .din2(g2146_p_spl_)
  );


  LA
  g_g2149_p
  (
    .dout(g2149_p),
    .din1(g2147_n),
    .din2(g2148_n)
  );


  FA
  g_g2149_n
  (
    .dout(g2149_n),
    .din1(g2147_p),
    .din2(g2148_p)
  );


  LA
  g_g2150_p
  (
    .dout(g2150_p),
    .din1(ffc_672_n),
    .din2(ffc_778_n)
  );


  FA
  g_g2150_n
  (
    .dout(g2150_n),
    .din1(ffc_672_p_spl_),
    .din2(ffc_778_p_spl_)
  );


  LA
  g_g2151_p
  (
    .dout(g2151_p),
    .din1(ffc_825_n_spl_0),
    .din2(g2150_n)
  );


  FA
  g_g2151_n
  (
    .dout(g2151_n),
    .din1(ffc_825_p_spl_0),
    .din2(g2150_p)
  );


  LA
  g_g2152_p
  (
    .dout(g2152_p),
    .din1(g2139_p_spl_0),
    .din2(g2151_n_spl_0)
  );


  FA
  g_g2152_n
  (
    .dout(g2152_n),
    .din1(g2139_n_spl_0),
    .din2(g2151_p_spl_0)
  );


  LA
  g_g2153_p
  (
    .dout(g2153_p),
    .din1(g2139_n_spl_),
    .din2(g2151_p_spl_0)
  );


  FA
  g_g2153_n
  (
    .dout(g2153_n),
    .din1(g2139_p_spl_0),
    .din2(g2151_n_spl_0)
  );


  LA
  g_g2154_p
  (
    .dout(g2154_p),
    .din1(g2152_n),
    .din2(g2153_n)
  );


  FA
  g_g2154_n
  (
    .dout(g2154_n),
    .din1(g2152_p),
    .din2(g2153_p)
  );


  LA
  g_g2155_p
  (
    .dout(g2155_p),
    .din1(g2149_n),
    .din2(g2154_n)
  );


  LA
  g_g2156_p
  (
    .dout(g2156_p),
    .din1(g2149_p),
    .din2(g2154_p)
  );


  FA
  g_g2157_n
  (
    .dout(g2157_n),
    .din1(g2155_p),
    .din2(g2156_p)
  );


  LA
  g_g2158_p
  (
    .dout(g2158_p),
    .din1(g1758_n_spl_0),
    .din2(g2157_n_spl_)
  );


  FA
  g_g2159_n
  (
    .dout(g2159_n),
    .din1(g1758_n_spl_1),
    .din2(g2157_n_spl_)
  );


  FA
  g_g2160_n
  (
    .dout(g2160_n),
    .din1(ffc_393_p_spl_0),
    .din2(g1790_n_spl_0)
  );


  LA
  g_g2161_p
  (
    .dout(g2161_p),
    .din1(ffc_821_n),
    .din2(ffc_822_p)
  );


  FA
  g_g2161_n
  (
    .dout(g2161_n),
    .din1(ffc_821_p),
    .din2(ffc_822_n)
  );


  LA
  g_g2162_p
  (
    .dout(g2162_p),
    .din1(g1702_n_spl_0),
    .din2(g2161_p_spl_)
  );


  FA
  g_g2162_n
  (
    .dout(g2162_n),
    .din1(g1702_p_spl_),
    .din2(g2161_n_spl_)
  );


  LA
  g_g2163_p
  (
    .dout(g2163_p),
    .din1(g1702_p_spl_),
    .din2(g2161_n_spl_)
  );


  FA
  g_g2163_n
  (
    .dout(g2163_n),
    .din1(g1702_n_spl_0),
    .din2(g2161_p_spl_)
  );


  LA
  g_g2164_p
  (
    .dout(g2164_p),
    .din1(g2162_n),
    .din2(g2163_n)
  );


  FA
  g_g2164_n
  (
    .dout(g2164_n),
    .din1(g2162_p),
    .din2(g2163_p)
  );


  LA
  g_g2165_p
  (
    .dout(g2165_p),
    .din1(ffc_673_n_spl_),
    .din2(g2164_p)
  );


  FA
  g_g2165_n
  (
    .dout(g2165_n),
    .din1(ffc_673_p_spl_0),
    .din2(g2164_n_spl_)
  );


  LA
  g_g2166_p
  (
    .dout(g2166_p),
    .din1(ffc_673_p_spl_0),
    .din2(g2164_n_spl_)
  );


  FA
  g_g2167_n
  (
    .dout(g2167_n),
    .din1(g2165_p_spl_),
    .din2(g2166_p)
  );


  LA
  g_g2168_p
  (
    .dout(g2168_p),
    .din1(ffc_770_n_spl_),
    .din2(g1703_n_spl_)
  );


  FA
  g_g2168_n
  (
    .dout(g2168_n),
    .din1(ffc_770_p_spl_0),
    .din2(g1703_p_spl_0)
  );


  LA
  g_g2169_p
  (
    .dout(g2169_p),
    .din1(g1705_n),
    .din2(g2168_n)
  );


  FA
  g_g2169_n
  (
    .dout(g2169_n),
    .din1(g1705_p_spl_),
    .din2(g2168_p)
  );


  LA
  g_g2170_p
  (
    .dout(g2170_p),
    .din1(ffc_674_p_spl_0),
    .din2(g2169_n_spl_)
  );


  FA
  g_g2170_n
  (
    .dout(g2170_n),
    .din1(ffc_674_n_spl_),
    .din2(g2169_p_spl_)
  );


  LA
  g_g2171_p
  (
    .dout(g2171_p),
    .din1(ffc_674_n_spl_),
    .din2(g2169_p_spl_)
  );


  FA
  g_g2171_n
  (
    .dout(g2171_n),
    .din1(ffc_674_p_spl_0),
    .din2(g2169_n_spl_)
  );


  LA
  g_g2172_p
  (
    .dout(g2172_p),
    .din1(g2170_n),
    .din2(g2171_n)
  );


  FA
  g_g2172_n
  (
    .dout(g2172_n),
    .din1(g2170_p),
    .din2(g2171_p)
  );


  LA
  g_g2173_p
  (
    .dout(g2173_p),
    .din1(g2167_n_spl_),
    .din2(g2172_n_spl_0)
  );


  FA
  g_g2174_n
  (
    .dout(g2174_n),
    .din1(g2167_n_spl_),
    .din2(g2172_n_spl_0)
  );


  LA
  g_g2175_p
  (
    .dout(g2175_p),
    .din1(g1793_n),
    .din2(g2096_n_spl_)
  );


  LA
  g_g2176_p
  (
    .dout(g2176_p),
    .din1(g1805_p_spl_),
    .din2(g1808_p_spl_)
  );


  FA
  g_g2177_n
  (
    .dout(g2177_n),
    .din1(g1806_p),
    .din2(g2176_p)
  );


  LA
  g_g2178_p
  (
    .dout(g2178_p),
    .din1(ffc_355_p_spl_0),
    .din2(ffc_629_p_spl_)
  );


  LA
  g_g2179_p
  (
    .dout(g2179_p),
    .din1(ffc_358_p_spl_),
    .din2(ffc_629_n)
  );


  FA
  g_g2180_n
  (
    .dout(g2180_n),
    .din1(g2178_p),
    .din2(g2179_p)
  );


  LA
  g_g2181_p
  (
    .dout(g2181_p),
    .din1(ffc_622_n_spl_),
    .din2(ffc_832_n_spl_010)
  );


  LA
  g_g2182_p
  (
    .dout(g2182_p),
    .din1(ffc_622_p_spl_0),
    .din2(ffc_833_n_spl_010)
  );


  FA
  g_g2183_n
  (
    .dout(g2183_n),
    .din1(g2181_p),
    .din2(g2182_p)
  );


  LA
  g_g2184_p
  (
    .dout(g2184_p),
    .din1(ffc_634_p_spl_),
    .din2(g2183_n)
  );


  LA
  g_g2185_p
  (
    .dout(g2185_p),
    .din1(ffc_622_p_spl_0),
    .din2(ffc_834_p_spl_001)
  );


  LA
  g_g2186_p
  (
    .dout(g2186_p),
    .din1(ffc_622_n_spl_),
    .din2(ffc_831_p_spl_001)
  );


  FA
  g_g2187_n
  (
    .dout(g2187_n),
    .din1(g2185_p),
    .din2(g2186_p)
  );


  LA
  g_g2188_p
  (
    .dout(g2188_p),
    .din1(ffc_634_n),
    .din2(g2187_n)
  );


  FA
  g_g2189_n
  (
    .dout(g2189_n),
    .din1(g2184_p),
    .din2(g2188_p)
  );


  LA
  g_g2190_p
  (
    .dout(g2190_p),
    .din1(ffc_621_n_spl_),
    .din2(ffc_832_n_spl_010)
  );


  LA
  g_g2191_p
  (
    .dout(g2191_p),
    .din1(ffc_621_p_spl_0),
    .din2(ffc_833_n_spl_010)
  );


  FA
  g_g2192_n
  (
    .dout(g2192_n),
    .din1(g2190_p),
    .din2(g2191_p)
  );


  LA
  g_g2193_p
  (
    .dout(g2193_p),
    .din1(ffc_635_p_spl_),
    .din2(g2192_n)
  );


  LA
  g_g2194_p
  (
    .dout(g2194_p),
    .din1(ffc_621_p_spl_0),
    .din2(ffc_834_p_spl_010)
  );


  LA
  g_g2195_p
  (
    .dout(g2195_p),
    .din1(ffc_621_n_spl_),
    .din2(ffc_831_p_spl_010)
  );


  FA
  g_g2196_n
  (
    .dout(g2196_n),
    .din1(g2194_p),
    .din2(g2195_p)
  );


  LA
  g_g2197_p
  (
    .dout(g2197_p),
    .din1(ffc_635_n),
    .din2(g2196_n)
  );


  FA
  g_g2198_n
  (
    .dout(g2198_n),
    .din1(g2193_p),
    .din2(g2197_p)
  );


  LA
  g_g2199_p
  (
    .dout(g2199_p),
    .din1(ffc_620_n_spl_),
    .din2(ffc_832_n_spl_011)
  );


  LA
  g_g2200_p
  (
    .dout(g2200_p),
    .din1(ffc_620_p_spl_0),
    .din2(ffc_833_n_spl_011)
  );


  FA
  g_g2201_n
  (
    .dout(g2201_n),
    .din1(g2199_p),
    .din2(g2200_p)
  );


  LA
  g_g2202_p
  (
    .dout(g2202_p),
    .din1(ffc_636_p_spl_),
    .din2(g2201_n)
  );


  LA
  g_g2203_p
  (
    .dout(g2203_p),
    .din1(ffc_620_p_spl_0),
    .din2(ffc_834_p_spl_010)
  );


  LA
  g_g2204_p
  (
    .dout(g2204_p),
    .din1(ffc_620_n_spl_),
    .din2(ffc_831_p_spl_010)
  );


  FA
  g_g2205_n
  (
    .dout(g2205_n),
    .din1(g2203_p),
    .din2(g2204_p)
  );


  LA
  g_g2206_p
  (
    .dout(g2206_p),
    .din1(ffc_636_n),
    .din2(g2205_n)
  );


  FA
  g_g2207_n
  (
    .dout(g2207_n),
    .din1(g2202_p),
    .din2(g2206_p)
  );


  LA
  g_g2208_p
  (
    .dout(g2208_p),
    .din1(ffc_627_n_spl_),
    .din2(ffc_832_n_spl_011)
  );


  LA
  g_g2209_p
  (
    .dout(g2209_p),
    .din1(ffc_627_p_spl_0),
    .din2(ffc_833_n_spl_011)
  );


  FA
  g_g2210_n
  (
    .dout(g2210_n),
    .din1(g2208_p),
    .din2(g2209_p)
  );


  LA
  g_g2211_p
  (
    .dout(g2211_p),
    .din1(ffc_650_p_spl_),
    .din2(g2210_n)
  );


  LA
  g_g2212_p
  (
    .dout(g2212_p),
    .din1(ffc_627_p_spl_0),
    .din2(ffc_834_p_spl_011)
  );


  LA
  g_g2213_p
  (
    .dout(g2213_p),
    .din1(ffc_627_n_spl_),
    .din2(ffc_831_p_spl_011)
  );


  FA
  g_g2214_n
  (
    .dout(g2214_n),
    .din1(g2212_p),
    .din2(g2213_p)
  );


  LA
  g_g2215_p
  (
    .dout(g2215_p),
    .din1(ffc_650_n),
    .din2(g2214_n)
  );


  FA
  g_g2216_n
  (
    .dout(g2216_n),
    .din1(g2211_p),
    .din2(g2215_p)
  );


  LA
  g_g2217_p
  (
    .dout(g2217_p),
    .din1(ffc_632_n_spl_),
    .din2(ffc_832_n_spl_100)
  );


  LA
  g_g2218_p
  (
    .dout(g2218_p),
    .din1(ffc_632_p_spl_0),
    .din2(ffc_833_n_spl_100)
  );


  FA
  g_g2219_n
  (
    .dout(g2219_n),
    .din1(g2217_p),
    .din2(g2218_p)
  );


  LA
  g_g2220_p
  (
    .dout(g2220_p),
    .din1(ffc_663_p_spl_),
    .din2(g2219_n)
  );


  LA
  g_g2221_p
  (
    .dout(g2221_p),
    .din1(ffc_632_p_spl_0),
    .din2(ffc_834_p_spl_011)
  );


  LA
  g_g2222_p
  (
    .dout(g2222_p),
    .din1(ffc_632_n_spl_),
    .din2(ffc_831_p_spl_011)
  );


  FA
  g_g2223_n
  (
    .dout(g2223_n),
    .din1(g2221_p),
    .din2(g2222_p)
  );


  LA
  g_g2224_p
  (
    .dout(g2224_p),
    .din1(ffc_663_n),
    .din2(g2223_n)
  );


  FA
  g_g2225_n
  (
    .dout(g2225_n),
    .din1(g2220_p),
    .din2(g2224_p)
  );


  LA
  g_g2226_p
  (
    .dout(g2226_p),
    .din1(ffc_631_n_spl_),
    .din2(ffc_832_n_spl_100)
  );


  LA
  g_g2227_p
  (
    .dout(g2227_p),
    .din1(ffc_631_p_spl_0),
    .din2(ffc_833_n_spl_100)
  );


  FA
  g_g2228_n
  (
    .dout(g2228_n),
    .din1(g2226_p),
    .din2(g2227_p)
  );


  LA
  g_g2229_p
  (
    .dout(g2229_p),
    .din1(ffc_664_p_spl_),
    .din2(g2228_n)
  );


  LA
  g_g2230_p
  (
    .dout(g2230_p),
    .din1(ffc_631_p_spl_0),
    .din2(ffc_834_p_spl_100)
  );


  LA
  g_g2231_p
  (
    .dout(g2231_p),
    .din1(ffc_631_n_spl_),
    .din2(ffc_831_p_spl_100)
  );


  FA
  g_g2232_n
  (
    .dout(g2232_n),
    .din1(g2230_p),
    .din2(g2231_p)
  );


  LA
  g_g2233_p
  (
    .dout(g2233_p),
    .din1(ffc_664_n),
    .din2(g2232_n)
  );


  FA
  g_g2234_n
  (
    .dout(g2234_n),
    .din1(g2229_p),
    .din2(g2233_p)
  );


  LA
  g_g2235_p
  (
    .dout(g2235_p),
    .din1(ffc_675_n_spl_),
    .din2(ffc_833_n_spl_101)
  );


  LA
  g_g2236_p
  (
    .dout(g2236_p),
    .din1(ffc_675_p_spl_0),
    .din2(ffc_832_n_spl_101)
  );


  FA
  g_g2237_n
  (
    .dout(g2237_n),
    .din1(g2235_p),
    .din2(g2236_p)
  );


  LA
  g_g2238_p
  (
    .dout(g2238_p),
    .din1(ffc_782_p),
    .din2(g2237_n)
  );


  LA
  g_g2239_p
  (
    .dout(g2239_p),
    .din1(ffc_675_n_spl_),
    .din2(ffc_834_p_spl_100)
  );


  LA
  g_g2240_p
  (
    .dout(g2240_p),
    .din1(ffc_675_p_spl_0),
    .din2(ffc_831_p_spl_100)
  );


  FA
  g_g2241_n
  (
    .dout(g2241_n),
    .din1(g2239_p),
    .din2(g2240_p)
  );


  LA
  g_g2242_p
  (
    .dout(g2242_p),
    .din1(ffc_782_n),
    .din2(g2241_n)
  );


  FA
  g_g2243_n
  (
    .dout(g2243_n),
    .din1(g2238_p),
    .din2(g2242_p)
  );


  LA
  g_g2244_p
  (
    .dout(g2244_p),
    .din1(ffc_795_n_spl_0),
    .din2(g1714_n_spl_0)
  );


  FA
  g_g2244_n
  (
    .dout(g2244_n),
    .din1(ffc_795_p_spl_0),
    .din2(g1714_p_spl_)
  );


  LA
  g_g2245_p
  (
    .dout(g2245_p),
    .din1(ffc_795_p_spl_1),
    .din2(g1714_p_spl_)
  );


  FA
  g_g2245_n
  (
    .dout(g2245_n),
    .din1(ffc_795_n_spl_),
    .din2(g1714_n_spl_0)
  );


  LA
  g_g2246_p
  (
    .dout(g2246_p),
    .din1(g2244_n),
    .din2(g2245_n)
  );


  FA
  g_g2246_n
  (
    .dout(g2246_n),
    .din1(g2244_p),
    .din2(g2245_p)
  );


  LA
  g_g2247_p
  (
    .dout(g2247_p),
    .din1(g1698_p_spl_),
    .din2(g2246_n)
  );


  LA
  g_g2248_p
  (
    .dout(g2248_p),
    .din1(g1698_n_spl_1),
    .din2(g2246_p)
  );


  FA
  g_g2249_n
  (
    .dout(g2249_n),
    .din1(g2247_p),
    .din2(g2248_p)
  );


  LA
  g_g2250_p
  (
    .dout(g2250_p),
    .din1(g2139_p_spl_),
    .din2(g2142_n_spl_)
  );


  LA
  g_g2251_p
  (
    .dout(g2251_p),
    .din1(ffc_756_n_spl_),
    .din2(ffc_825_n_spl_1)
  );


  FA
  g_g2251_n
  (
    .dout(g2251_n),
    .din1(ffc_756_p_spl_1),
    .din2(ffc_825_p_spl_0)
  );


  LA
  g_g2252_p
  (
    .dout(g2252_p),
    .din1(ffc_769_p_spl_1),
    .din2(ffc_825_p_spl_1)
  );


  FA
  g_g2252_n
  (
    .dout(g2252_n),
    .din1(ffc_769_n_spl_),
    .din2(ffc_825_n_spl_1)
  );


  LA
  g_g2253_p
  (
    .dout(g2253_p),
    .din1(ffc_826_n_spl_1),
    .din2(g2252_n)
  );


  FA
  g_g2253_n
  (
    .dout(g2253_n),
    .din1(ffc_826_p_spl_1),
    .din2(g2252_p)
  );


  LA
  g_g2254_p
  (
    .dout(g2254_p),
    .din1(ffc_755_p_spl_),
    .din2(g2253_n_spl_)
  );


  FA
  g_g2254_n
  (
    .dout(g2254_n),
    .din1(ffc_755_n_spl_),
    .din2(g2253_p_spl_)
  );


  LA
  g_g2255_p
  (
    .dout(g2255_p),
    .din1(ffc_755_n_spl_),
    .din2(g2253_p_spl_)
  );


  FA
  g_g2255_n
  (
    .dout(g2255_n),
    .din1(ffc_755_p_spl_),
    .din2(g2253_n_spl_)
  );


  LA
  g_g2256_p
  (
    .dout(g2256_p),
    .din1(g2254_n),
    .din2(g2255_n)
  );


  FA
  g_g2256_n
  (
    .dout(g2256_n),
    .din1(g2254_p),
    .din2(g2255_p)
  );


  LA
  g_g2257_p
  (
    .dout(g2257_p),
    .din1(g2251_n),
    .din2(g2256_p)
  );


  LA
  g_g2258_p
  (
    .dout(g2258_p),
    .din1(g2251_p),
    .din2(g2256_n)
  );


  FA
  g_g2259_n
  (
    .dout(g2259_n),
    .din1(g2257_p),
    .din2(g2258_p)
  );


  FA
  g_g2260_n
  (
    .dout(g2260_n),
    .din1(g2250_p_spl_),
    .din2(g2259_n_spl_)
  );


  LA
  g_g2261_p
  (
    .dout(g2261_p),
    .din1(g2250_p_spl_),
    .din2(g2259_n_spl_)
  );


  LA
  g_g2262_p
  (
    .dout(g2262_p),
    .din1(ffc_334_p_spl_),
    .din2(ffc_839_p_spl_11)
  );


  LA
  g_g2263_p
  (
    .dout(g2263_p),
    .din1(ffc_335_p),
    .din2(ffc_839_n_spl_11)
  );


  FA
  g_g2264_n
  (
    .dout(g2264_n),
    .din1(g2262_p),
    .din2(g2263_p)
  );


  FA
  g_g2265_n
  (
    .dout(g2265_n),
    .din1(ffc_370_n),
    .din2(ffc_863_n_spl_10)
  );


  FA
  g_g2266_n
  (
    .dout(g2266_n),
    .din1(ffc_371_n),
    .din2(ffc_863_p_spl_10)
  );


  LA
  g_g2267_p
  (
    .dout(g2267_p),
    .din1(g2265_n),
    .din2(g2266_n)
  );


  FA
  g_g2268_n
  (
    .dout(g2268_n),
    .din1(ffc_395_n),
    .din2(g1898_p)
  );


  LA
  g_g2269_p
  (
    .dout(g2269_p),
    .din1(g1725_n_spl_),
    .din2(g1768_n_spl_)
  );


  FA
  g_g2270_n
  (
    .dout(g2270_n),
    .din1(g1758_p_spl_0),
    .din2(g2151_p_spl_)
  );


  FA
  g_g2271_n
  (
    .dout(g2271_n),
    .din1(g1758_n_spl_1),
    .din2(g2151_n_spl_)
  );


  LA
  g_g2272_p
  (
    .dout(g2272_p),
    .din1(g2270_n),
    .din2(g2271_n)
  );


  FA
  g_g2273_n
  (
    .dout(g2273_n),
    .din1(g2269_p_spl_),
    .din2(g2272_p_spl_)
  );


  LA
  g_g2274_p
  (
    .dout(g2274_p),
    .din1(g2269_p_spl_),
    .din2(g2272_p_spl_)
  );


  FA
  g_g2275_n
  (
    .dout(g2275_n),
    .din1(g1764_p_spl_0),
    .din2(g1809_p_spl_)
  );


  FA
  g_g2276_n
  (
    .dout(g2276_n),
    .din1(g2099_p_spl_0),
    .din2(g2275_n_spl_)
  );


  LA
  g_g2277_p
  (
    .dout(g2277_p),
    .din1(g2108_n_spl_0),
    .din2(g2123_n_spl_0)
  );


  FA
  g_g2278_n
  (
    .dout(g2278_n),
    .din1(g2108_n_spl_0),
    .din2(g2123_n_spl_0)
  );


  LA
  g_g2279_p
  (
    .dout(g2279_p),
    .din1(g2117_n_spl_0),
    .din2(g2126_p_spl_0)
  );


  FA
  g_g2280_n
  (
    .dout(g2280_n),
    .din1(g2117_n_spl_0),
    .din2(g2126_p_spl_0)
  );


  LA
  g_g2281_p
  (
    .dout(g2281_p),
    .din1(ffc_764_p_spl_0),
    .din2(ffc_832_n_spl_101)
  );


  FA
  g_g2281_n
  (
    .dout(g2281_n),
    .din1(ffc_764_n_spl_),
    .din2(ffc_832_p_spl_00)
  );


  LA
  g_g2282_p
  (
    .dout(g2282_p),
    .din1(ffc_764_n_spl_),
    .din2(ffc_831_p_spl_101)
  );


  FA
  g_g2282_n
  (
    .dout(g2282_n),
    .din1(ffc_764_p_spl_0),
    .din2(ffc_831_n_spl_00)
  );


  LA
  g_g2283_p
  (
    .dout(g2283_p),
    .din1(g2281_n),
    .din2(g2282_n)
  );


  FA
  g_g2283_n
  (
    .dout(g2283_n),
    .din1(g2281_p),
    .din2(g2282_p)
  );


  LA
  g_g2284_p
  (
    .dout(g2284_p),
    .din1(ffc_781_n_spl_0),
    .din2(ffc_832_n_spl_110)
  );


  FA
  g_g2284_n
  (
    .dout(g2284_n),
    .din1(ffc_781_p_spl_00),
    .din2(ffc_832_p_spl_00)
  );


  LA
  g_g2285_p
  (
    .dout(g2285_p),
    .din1(ffc_781_p_spl_00),
    .din2(ffc_833_n_spl_101)
  );


  FA
  g_g2285_n
  (
    .dout(g2285_n),
    .din1(ffc_781_n_spl_0),
    .din2(ffc_833_p_spl_0)
  );


  LA
  g_g2286_p
  (
    .dout(g2286_p),
    .din1(g2284_n),
    .din2(g2285_n)
  );


  FA
  g_g2286_n
  (
    .dout(g2286_n),
    .din1(g2284_p),
    .din2(g2285_p)
  );


  LA
  g_g2287_p
  (
    .dout(g2287_p),
    .din1(ffc_816_p_spl_0),
    .din2(g2286_n)
  );


  FA
  g_g2287_n
  (
    .dout(g2287_n),
    .din1(ffc_816_n_spl_1),
    .din2(g2286_p)
  );


  LA
  g_g2288_p
  (
    .dout(g2288_p),
    .din1(ffc_781_p_spl_0),
    .din2(ffc_834_p_spl_101)
  );


  FA
  g_g2288_n
  (
    .dout(g2288_n),
    .din1(ffc_781_n_spl_1),
    .din2(ffc_834_n_spl_0)
  );


  LA
  g_g2289_p
  (
    .dout(g2289_p),
    .din1(ffc_781_n_spl_1),
    .din2(ffc_831_p_spl_101)
  );


  FA
  g_g2289_n
  (
    .dout(g2289_n),
    .din1(ffc_781_p_spl_1),
    .din2(ffc_831_n_spl_00)
  );


  LA
  g_g2290_p
  (
    .dout(g2290_p),
    .din1(g2288_n),
    .din2(g2289_n)
  );


  FA
  g_g2290_n
  (
    .dout(g2290_n),
    .din1(g2288_p),
    .din2(g2289_p)
  );


  LA
  g_g2291_p
  (
    .dout(g2291_p),
    .din1(ffc_816_n_spl_1),
    .din2(g2290_n)
  );


  FA
  g_g2291_n
  (
    .dout(g2291_n),
    .din1(ffc_816_p_spl_1),
    .din2(g2290_p)
  );


  LA
  g_g2292_p
  (
    .dout(g2292_p),
    .din1(g2287_n),
    .din2(g2291_n)
  );


  FA
  g_g2292_n
  (
    .dout(g2292_n),
    .din1(g2287_p),
    .din2(g2291_p)
  );


  LA
  g_g2293_p
  (
    .dout(g2293_p),
    .din1(g2283_p),
    .din2(g2292_n)
  );


  LA
  g_g2294_p
  (
    .dout(g2294_p),
    .din1(g2283_n),
    .din2(g2292_p)
  );


  FA
  g_g2295_n
  (
    .dout(g2295_n),
    .din1(g2293_p),
    .din2(g2294_p)
  );


  FA
  g_g2296_n
  (
    .dout(g2296_n),
    .din1(g2120_n_spl_0),
    .din2(g2295_n_spl_)
  );


  LA
  g_g2297_p
  (
    .dout(g2297_p),
    .din1(g2120_n_spl_0),
    .din2(g2295_n_spl_)
  );


  LA
  g_g2298_p
  (
    .dout(g2298_p),
    .din1(ffc_648_n_spl_),
    .din2(ffc_832_n_spl_110)
  );


  LA
  g_g2299_p
  (
    .dout(g2299_p),
    .din1(ffc_648_p_spl_0),
    .din2(ffc_833_n_spl_110)
  );


  FA
  g_g2300_n
  (
    .dout(g2300_n),
    .din1(g2298_p),
    .din2(g2299_p)
  );


  LA
  g_g2301_p
  (
    .dout(g2301_p),
    .din1(ffc_679_p_spl_),
    .din2(g2300_n)
  );


  LA
  g_g2302_p
  (
    .dout(g2302_p),
    .din1(ffc_648_p_spl_0),
    .din2(ffc_834_p_spl_101)
  );


  LA
  g_g2303_p
  (
    .dout(g2303_p),
    .din1(ffc_648_n_spl_),
    .din2(ffc_831_p_spl_110)
  );


  FA
  g_g2304_n
  (
    .dout(g2304_n),
    .din1(g2302_p),
    .din2(g2303_p)
  );


  LA
  g_g2305_p
  (
    .dout(g2305_p),
    .din1(ffc_679_n),
    .din2(g2304_n)
  );


  FA
  g_g2306_n
  (
    .dout(g2306_n),
    .din1(g2301_p),
    .din2(g2305_p)
  );


  FA
  g_g2307_n
  (
    .dout(g2307_n),
    .din1(ffc_661_p_spl_0),
    .din2(ffc_832_p_spl_0)
  );


  FA
  g_g2308_n
  (
    .dout(g2308_n),
    .din1(ffc_661_n_spl_),
    .din2(ffc_833_p_spl_0)
  );


  LA
  g_g2309_p
  (
    .dout(g2309_p),
    .din1(g2307_n),
    .din2(g2308_n)
  );


  FA
  g_g2310_n
  (
    .dout(g2310_n),
    .din1(ffc_765_n),
    .din2(g2309_p)
  );


  FA
  g_g2311_n
  (
    .dout(g2311_n),
    .din1(ffc_661_n_spl_),
    .din2(ffc_834_n_spl_0)
  );


  FA
  g_g2312_n
  (
    .dout(g2312_n),
    .din1(ffc_661_p_spl_0),
    .din2(ffc_831_n_spl_0)
  );


  LA
  g_g2313_p
  (
    .dout(g2313_p),
    .din1(g2311_n),
    .din2(g2312_n)
  );


  FA
  g_g2314_n
  (
    .dout(g2314_n),
    .din1(ffc_765_p_spl_),
    .din2(g2313_p)
  );


  LA
  g_g2315_p
  (
    .dout(g2315_p),
    .din1(g2310_n),
    .din2(g2314_n)
  );


  FA
  g_g2316_n
  (
    .dout(g2316_n),
    .din1(g2306_n_spl_),
    .din2(g2315_p_spl_)
  );


  LA
  g_g2317_p
  (
    .dout(g2317_p),
    .din1(g2306_n_spl_),
    .din2(g2315_p_spl_)
  );


  LA
  g_g2318_p
  (
    .dout(g2318_p),
    .din1(ffc_779_n),
    .din2(g1699_n_spl_1)
  );


  LA
  g_g2319_p
  (
    .dout(g2319_p),
    .din1(ffc_779_p_spl_),
    .din2(g1699_p_spl_)
  );


  FA
  g_g2320_n
  (
    .dout(g2320_n),
    .din1(g2318_p),
    .din2(g2319_p)
  );


  LA
  g_g2321_p
  (
    .dout(g2321_p),
    .din1(g1712_p_spl_0),
    .din2(g2320_n)
  );


  FA
  g_g2322_n
  (
    .dout(g2322_n),
    .din1(g1785_p_spl_),
    .din2(g2321_p)
  );


  LA
  g_g2323_p
  (
    .dout(g2323_p),
    .din1(g1774_p),
    .din2(g2322_n)
  );


  LA
  g_g2324_p
  (
    .dout(g2324_p),
    .din1(g1774_n_spl_),
    .din2(g1787_n_spl_)
  );


  FA
  g_g2325_n
  (
    .dout(g2325_n),
    .din1(g2323_p),
    .din2(g2324_p)
  );


  LA
  g_g2326_p
  (
    .dout(g2326_p),
    .din1(g1697_n_spl_0),
    .din2(g1701_p_spl_)
  );


  FA
  g_g2326_n
  (
    .dout(g2326_n),
    .din1(g1697_p_spl_),
    .din2(g1701_n_spl_0)
  );


  LA
  g_g2327_p
  (
    .dout(g2327_p),
    .din1(g1697_p_spl_),
    .din2(g1701_n_spl_0)
  );


  FA
  g_g2327_n
  (
    .dout(g2327_n),
    .din1(g1697_n_spl_0),
    .din2(g1701_p_spl_)
  );


  LA
  g_g2328_p
  (
    .dout(g2328_p),
    .din1(ffc_673_p_spl_1),
    .din2(g2327_n)
  );


  FA
  g_g2328_n
  (
    .dout(g2328_n),
    .din1(ffc_673_n_spl_),
    .din2(g2327_p)
  );


  LA
  g_g2329_p
  (
    .dout(g2329_p),
    .din1(g2326_n),
    .din2(g2328_p)
  );


  FA
  g_g2329_n
  (
    .dout(g2329_n),
    .din1(g2326_p),
    .din2(g2328_n)
  );


  LA
  g_g2330_p
  (
    .dout(g2330_p),
    .din1(g2165_n),
    .din2(g2329_n)
  );


  FA
  g_g2330_n
  (
    .dout(g2330_n),
    .din1(g2165_p_spl_),
    .din2(g2329_p)
  );


  FA
  g_g2331_n
  (
    .dout(g2331_n),
    .din1(g2172_p),
    .din2(g2330_p)
  );


  FA
  g_g2332_n
  (
    .dout(g2332_n),
    .din1(g2172_n_spl_),
    .din2(g2330_n)
  );


  LA
  g_g2333_p
  (
    .dout(g2333_p),
    .din1(g2331_n),
    .din2(g2332_n)
  );


  LA
  g_g2334_p
  (
    .dout(g2334_p),
    .din1(ffc_660_n_spl_0),
    .din2(ffc_832_n_spl_111)
  );


  FA
  g_g2334_n
  (
    .dout(g2334_n),
    .din1(ffc_660_p_spl_00),
    .din2(ffc_832_p_spl_1)
  );


  LA
  g_g2335_p
  (
    .dout(g2335_p),
    .din1(ffc_660_p_spl_00),
    .din2(ffc_833_n_spl_110)
  );


  FA
  g_g2335_n
  (
    .dout(g2335_n),
    .din1(ffc_660_n_spl_0),
    .din2(ffc_833_p_spl_1)
  );


  LA
  g_g2336_p
  (
    .dout(g2336_p),
    .din1(g2334_n),
    .din2(g2335_n)
  );


  FA
  g_g2336_n
  (
    .dout(g2336_n),
    .din1(g2334_p),
    .din2(g2335_p)
  );


  LA
  g_g2337_p
  (
    .dout(g2337_p),
    .din1(ffc_763_p_spl_0),
    .din2(g2336_n)
  );


  FA
  g_g2337_n
  (
    .dout(g2337_n),
    .din1(ffc_763_n_spl_),
    .din2(g2336_p)
  );


  LA
  g_g2338_p
  (
    .dout(g2338_p),
    .din1(ffc_660_p_spl_0),
    .din2(ffc_834_p_spl_11)
  );


  FA
  g_g2338_n
  (
    .dout(g2338_n),
    .din1(ffc_660_n_spl_1),
    .din2(ffc_834_n_spl_1)
  );


  LA
  g_g2339_p
  (
    .dout(g2339_p),
    .din1(ffc_660_n_spl_1),
    .din2(ffc_831_p_spl_110)
  );


  FA
  g_g2339_n
  (
    .dout(g2339_n),
    .din1(ffc_660_p_spl_1),
    .din2(ffc_831_n_spl_1)
  );


  LA
  g_g2340_p
  (
    .dout(g2340_p),
    .din1(g2338_n),
    .din2(g2339_n)
  );


  FA
  g_g2340_n
  (
    .dout(g2340_n),
    .din1(g2338_p),
    .din2(g2339_p)
  );


  LA
  g_g2341_p
  (
    .dout(g2341_p),
    .din1(ffc_763_n_spl_),
    .din2(g2340_n)
  );


  FA
  g_g2341_n
  (
    .dout(g2341_n),
    .din1(ffc_763_p_spl_0),
    .din2(g2340_p)
  );


  LA
  g_g2342_p
  (
    .dout(g2342_p),
    .din1(g2337_n),
    .din2(g2341_n)
  );


  FA
  g_g2342_n
  (
    .dout(g2342_n),
    .din1(g2337_p),
    .din2(g2341_p)
  );


  LA
  g_g2343_p
  (
    .dout(g2343_p),
    .din1(ffc_829_n_spl_00),
    .din2(ffc_832_n_spl_111)
  );


  FA
  g_g2343_n
  (
    .dout(g2343_n),
    .din1(ffc_829_p_spl_00),
    .din2(ffc_832_p_spl_1)
  );


  LA
  g_g2344_p
  (
    .dout(g2344_p),
    .din1(ffc_829_p_spl_01),
    .din2(ffc_833_n_spl_11)
  );


  FA
  g_g2344_n
  (
    .dout(g2344_n),
    .din1(ffc_829_n_spl_0),
    .din2(ffc_833_p_spl_1)
  );


  LA
  g_g2345_p
  (
    .dout(g2345_p),
    .din1(g2343_n),
    .din2(g2344_n)
  );


  FA
  g_g2345_n
  (
    .dout(g2345_n),
    .din1(g2343_p),
    .din2(g2344_p)
  );


  LA
  g_g2346_p
  (
    .dout(g2346_p),
    .din1(ffc_390_p_spl_0),
    .din2(g2345_n)
  );


  FA
  g_g2346_n
  (
    .dout(g2346_n),
    .din1(ffc_390_n_spl_1),
    .din2(g2345_p)
  );


  LA
  g_g2347_p
  (
    .dout(g2347_p),
    .din1(ffc_829_p_spl_01),
    .din2(ffc_834_p_spl_11)
  );


  FA
  g_g2347_n
  (
    .dout(g2347_n),
    .din1(ffc_829_n_spl_1),
    .din2(ffc_834_n_spl_1)
  );


  LA
  g_g2348_p
  (
    .dout(g2348_p),
    .din1(ffc_829_n_spl_1),
    .din2(ffc_831_p_spl_11)
  );


  FA
  g_g2348_n
  (
    .dout(g2348_n),
    .din1(ffc_829_p_spl_1),
    .din2(ffc_831_n_spl_1)
  );


  LA
  g_g2349_p
  (
    .dout(g2349_p),
    .din1(g2347_n),
    .din2(g2348_n)
  );


  FA
  g_g2349_n
  (
    .dout(g2349_n),
    .din1(g2347_p),
    .din2(g2348_p)
  );


  LA
  g_g2350_p
  (
    .dout(g2350_p),
    .din1(ffc_390_n_spl_1),
    .din2(g2349_n)
  );


  FA
  g_g2350_n
  (
    .dout(g2350_n),
    .din1(ffc_390_p_spl_1),
    .din2(g2349_p)
  );


  LA
  g_g2351_p
  (
    .dout(g2351_p),
    .din1(g2346_n),
    .din2(g2350_n)
  );


  FA
  g_g2351_n
  (
    .dout(g2351_n),
    .din1(g2346_p),
    .din2(g2350_p)
  );


  LA
  g_g2352_p
  (
    .dout(g2352_p),
    .din1(g2342_p),
    .din2(g2351_n)
  );


  LA
  g_g2353_p
  (
    .dout(g2353_p),
    .din1(g2342_n),
    .din2(g2351_p)
  );


  FA
  g_g2354_n
  (
    .dout(g2354_n),
    .din1(g2352_p),
    .din2(g2353_p)
  );


  LA
  g_g2355_p
  (
    .dout(g2355_p),
    .din1(ffc_442_n_spl_),
    .din2(g1716_p)
  );


  FA
  g_g2355_n
  (
    .dout(g2355_n),
    .din1(ffc_442_p_spl_),
    .din2(g1716_n_spl_)
  );


  LA
  g_g2356_p
  (
    .dout(g2356_p),
    .din1(ffc_442_p_spl_),
    .din2(ffc_815_n_spl_)
  );


  FA
  g_g2356_n
  (
    .dout(g2356_n),
    .din1(ffc_442_n_spl_),
    .din2(ffc_815_p_spl_)
  );


  LA
  g_g2357_p
  (
    .dout(g2357_p),
    .din1(g2355_n),
    .din2(g2356_n)
  );


  FA
  g_g2357_n
  (
    .dout(g2357_n),
    .din1(g2355_p),
    .din2(g2356_p)
  );


  LA
  g_g2358_p
  (
    .dout(g2358_p),
    .din1(g1792_p_spl_),
    .din2(g2357_n)
  );


  LA
  g_g2359_p
  (
    .dout(g2359_p),
    .din1(g1792_n),
    .din2(g2357_p)
  );


  FA
  g_g2360_n
  (
    .dout(g2360_n),
    .din1(g2358_p),
    .din2(g2359_p)
  );


  FA
  g_g2361_n
  (
    .dout(g2361_n),
    .din1(ffc_387_n),
    .din2(g2129_p)
  );


  FA
  g_g2362_n
  (
    .dout(g2362_n),
    .din1(ffc_396_n),
    .din2(g2132_p)
  );


  FA
  g_g2363_n
  (
    .dout(g2363_n),
    .din1(ffc_396_p_spl_),
    .din2(g2132_n_spl_)
  );


  FA
  g_g2364_n
  (
    .dout(g2364_n),
    .din1(ffc_397_p_spl_),
    .din2(g1802_n_spl_)
  );


  LA
  g_g2365_p
  (
    .dout(g2365_p),
    .din1(g2133_n_spl_),
    .din2(g2364_n)
  );


  LA
  g_g2366_p
  (
    .dout(g2366_p),
    .din1(ffc_360_p_spl_),
    .din2(ffc_863_p_spl_10)
  );


  LA
  g_g2367_p
  (
    .dout(g2367_p),
    .din1(ffc_361_p),
    .din2(ffc_863_n_spl_11)
  );


  LA
  g_g2368_p
  (
    .dout(g2368_p),
    .din1(ffc_362_p_spl_),
    .din2(ffc_863_p_spl_11)
  );


  LA
  g_g2369_p
  (
    .dout(g2369_p),
    .din1(ffc_363_p),
    .din2(ffc_863_n_spl_11)
  );


  LA
  g_g2370_p
  (
    .dout(g2370_p),
    .din1(g1763_n_spl_0),
    .din2(g2276_n_spl_0)
  );


  FA
  g_g2371_n
  (
    .dout(g2371_n),
    .din1(g1763_n_spl_1),
    .din2(g2276_n_spl_0)
  );


  LA
  g_g2372_p
  (
    .dout(g2372_p),
    .din1(g1764_p_spl_0),
    .din2(g2137_p_spl_0)
  );


  LA
  g_g2373_p
  (
    .dout(g2373_p),
    .din1(g1807_n_spl_),
    .din2(g2160_n_spl_0)
  );


  LA
  g_g2374_p
  (
    .dout(g2374_p),
    .din1(g1796_p_spl_0),
    .din2(g2175_p_spl_)
  );


  LA
  g_g2375_p
  (
    .dout(g2375_p),
    .din1(g2098_n_spl_),
    .din2(g2135_p_spl_)
  );


  FA
  g_g2376_n
  (
    .dout(g2376_n),
    .din1(g1803_p_spl_),
    .din2(g2375_p)
  );


  LA
  g_g2377_p
  (
    .dout(g2377_p),
    .din1(g2099_p_spl_0),
    .din2(g2137_p_spl_0)
  );


  FA
  g_g2378_n
  (
    .dout(g2378_n),
    .din1(g1804_p_spl_),
    .din2(g2377_p)
  );


  LA
  g_g2379_p
  (
    .dout(g2379_p),
    .din1(g2137_p_spl_1),
    .din2(g2275_n_spl_)
  );


  FA
  g_g2380_n
  (
    .dout(g2380_n),
    .din1(g2160_n_spl_0),
    .din2(g2177_n_spl_)
  );


  LA
  g_g2381_p
  (
    .dout(g2381_p),
    .din1(ffc_391_p_spl_0),
    .din2(g2264_n_spl_0)
  );


  FA
  g_g2382_n
  (
    .dout(g2382_n),
    .din1(ffc_391_p_spl_0),
    .din2(g2264_n_spl_0)
  );


  LA
  g_g2383_p
  (
    .dout(g2383_p),
    .din1(g2267_p_spl_),
    .din2(g2365_p_spl_)
  );


  FA
  g_g2384_n
  (
    .dout(g2384_n),
    .din1(ffc_395_p_spl_),
    .din2(g1898_n_spl_)
  );


  LA
  g_g2385_p
  (
    .dout(g2385_p),
    .din1(g2268_n_spl_),
    .din2(g2384_n)
  );


  FA
  g_g2386_n
  (
    .dout(g2386_n),
    .din1(ffc_387_p_spl_),
    .din2(g2129_n_spl_)
  );


  LA
  g_g2387_p
  (
    .dout(g2387_p),
    .din1(g2361_n_spl_),
    .din2(g2386_n)
  );


  LA
  g_g2388_p
  (
    .dout(g2388_p),
    .din1(g2362_n_spl_),
    .din2(g2363_n_spl_)
  );


  LA
  g_g2389_p
  (
    .dout(g2389_p),
    .din1(G92_p_spl_),
    .din2(G124_p_spl_0)
  );


  LA
  g_g2390_p
  (
    .dout(g2390_p),
    .din1(G93_p),
    .din2(G124_n_spl_0)
  );


  LA
  g_g2391_p
  (
    .dout(g2391_p),
    .din1(G94_p_spl_),
    .din2(G124_p_spl_0)
  );


  LA
  g_g2392_p
  (
    .dout(g2392_p),
    .din1(G95_p),
    .din2(G124_n_spl_0)
  );


  LA
  g_g2393_p
  (
    .dout(g2393_p),
    .din1(G107_p_spl_),
    .din2(G124_p_spl_1)
  );


  LA
  g_g2394_p
  (
    .dout(g2394_p),
    .din1(G108_p),
    .din2(G124_n_spl_)
  );


  buf

  (
    G5193_p,
    ffc_249_n
  );


  buf

  (
    G5194_p,
    ffc_356_n
  );


  buf

  (
    G5195_p,
    ffc_454_n_spl_
  );


  buf

  (
    G5196_p,
    ffc_401_n_spl_0
  );


  buf

  (
    G5197_p,
    ffc_368_n
  );


  buf

  (
    G5198_p,
    ffc_372_n
  );


  buf

  (
    G5199_n,
    g1049_n_spl_
  );


  buf

  (
    G5200_p,
    ffc_405_n
  );


  buf

  (
    G5201_p,
    ffc_401_n_spl_0
  );


  buf

  (
    G5202_p,
    ffc_401_n_spl_
  );


  buf

  (
    G5203_p,
    ffc_365_n
  );


  buf

  (
    G5204_p,
    ffc_369_n
  );


  buf

  (
    G5205_p,
    g1050_p
  );


  buf

  (
    G5206_p,
    ffc_342_n_spl_
  );


  buf

  (
    G5207_p,
    ffc_409_n_spl_
  );


  buf

  (
    G5208_p,
    ffc_421_n_spl_
  );


  buf

  (
    G5209_p,
    ffc_417_n_spl_
  );


  buf

  (
    G5210_p,
    g1051_p
  );


  buf

  (
    G5211_p,
    g1052_p
  );


  buf

  (
    G5212_p,
    g1053_n
  );


  buf

  (
    G5213_p,
    g1054_n_spl_
  );


  buf

  (
    G5214_p,
    ffc_241_p_spl_111
  );


  buf

  (
    G5215_p,
    ffc_249_p_spl_1
  );


  buf

  (
    G5216_p,
    ffc_3_p_spl_
  );


  buf

  (
    G5217_p,
    ffc_405_p_spl_
  );


  buf

  (
    G5218_p,
    ffc_359_p
  );


  buf

  (
    G5219_p,
    ffc_405_p_spl_
  );


  buf

  (
    G5220_p,
    g1056_n
  );


  buf

  (
    G5221_p,
    g1055_n_spl_11
  );


  buf

  (
    G5222_p,
    ffc_3_n_spl_0
  );


  buf

  (
    G5223_p,
    ffc_3_n_spl_0
  );


  buf

  (
    G5224_p,
    ffc_3_n_spl_1
  );


  buf

  (
    G5225_p,
    ffc_3_n_spl_1
  );


  buf

  (
    G5226_p,
    ffc_359_n_spl_
  );


  buf

  (
    G5227_p,
    ffc_359_n_spl_
  );


  buf

  (
    G5228_p,
    g1060_n
  );


  buf

  (
    G5229_p,
    g1064_n_spl_
  );


  buf

  (
    G5230_p,
    g1064_n_spl_
  );


  buf

  (
    G5231_p,
    g1065_n
  );


  buf

  (
    G5232_p,
    g1070_p
  );


  buf

  (
    G5233_p,
    g1075_p
  );


  buf

  (
    G5234_p,
    g1080_p
  );


  buf

  (
    G5235_p,
    g1085_p
  );


  buf

  (
    G5236_p,
    g1091_p
  );


  buf

  (
    G5237_p,
    g1100_p
  );


  buf

  (
    G5238_n,
    g1102_n_spl_
  );


  buf

  (
    G5239_p,
    g1106_p_spl_
  );


  buf

  (
    G5240_p,
    g1106_p_spl_
  );


  buf

  (
    G5241_n,
    g1102_n_spl_
  );


  buf

  (
    G5242_n,
    g1111_n_spl_
  );


  buf

  (
    G5243_n,
    g1120_n_spl_
  );


  buf

  (
    G5244_n,
    g1126_p_spl_
  );


  buf

  (
    G5245_p,
    g1127_n_spl_
  );


  buf

  (
    G5246_n,
    g1126_p_spl_
  );


  buf

  (
    G5247_p,
    g1127_n_spl_
  );


  buf

  (
    G5248_n,
    g1132_n_spl_1
  );


  buf

  (
    G5249_p,
    g1137_p_spl_1
  );


  buf

  (
    G5250_n,
    g1142_n_spl_1
  );


  buf

  (
    G5251_p,
    ffc_561_p_spl_1
  );


  buf

  (
    G5252_p,
    g1151_n
  );


  buf

  (
    G5253_n,
    g1155_n_spl_1
  );


  buf

  (
    G5254_n,
    g1158_n_spl_1
  );


  buf

  (
    G5255_n,
    g1164_n_spl_1
  );


  buf

  (
    G5256_p,
    g1173_n
  );


  buf

  (
    G5257_n,
    g1182_n_spl_1
  );


  buf

  (
    G5258_n,
    g1187_n_spl_1
  );


  buf

  (
    G5259_n,
    g1194_n_spl_1
  );


  buf

  (
    G5260_p,
    g1200_p_spl_1
  );


  buf

  (
    G5261_n,
    g1212_n_spl_
  );


  buf

  (
    G5262_n,
    g1233_n_spl_
  );


  buf

  (
    G5263_n,
    g1248_n
  );


  buf

  (
    G5264_n,
    g1257_n
  );


  buf

  (
    G5265_p,
    g1267_p
  );


  buf

  (
    G5266_p,
    g1277_p
  );


  buf

  (
    G5267_p,
    g1286_p
  );


  buf

  (
    G5268_p,
    g1295_p
  );


  buf

  (
    G5269_p,
    g1304_p
  );


  buf

  (
    G5270_n,
    g1313_p
  );


  buf

  (
    G5271_p,
    g1322_p
  );


  buf

  (
    G5272_p,
    g1331_p
  );


  buf

  (
    G5273_p,
    g1340_p
  );


  buf

  (
    G5274_n,
    g1349_p
  );


  buf

  (
    G5275_p,
    g1359_p
  );


  buf

  (
    G5276_n,
    g1369_n
  );


  buf

  (
    G5277_p,
    g1379_p
  );


  buf

  (
    G5278_p,
    g1389_p
  );


  buf

  (
    G5279_p,
    g1399_p
  );


  buf

  (
    G5280_n,
    g1409_n
  );


  buf

  (
    G5281_p,
    g1419_p
  );


  buf

  (
    G5282_p,
    g1429_p
  );


  buf

  (
    G5283_p,
    g1443_p
  );


  buf

  (
    G5284_p,
    g1446_p
  );


  buf

  (
    G5285_n,
    g1449_n_spl_1
  );


  buf

  (
    G5286_n,
    g1453_n_spl_1
  );


  buf

  (
    G5287_n,
    g1457_n_spl_1
  );


  buf

  (
    G5288_n,
    g1460_n_spl_1
  );


  buf

  (
    G5289_n,
    g1467_n
  );


  buf

  (
    G5290_n,
    g1470_n_spl_1
  );


  buf

  (
    G5291_n,
    g1476_n_spl_1
  );


  buf

  (
    G5292_n,
    g1482_n_spl_1
  );


  buf

  (
    G5293_n,
    g1486_n_spl_1
  );


  buf

  (
    G5294_p,
    g1495_n
  );


  buf

  (
    G5295_p,
    g1504_p
  );


  buf

  (
    G5296_p,
    g1513_p
  );


  buf

  (
    G5297_p,
    g1522_p
  );


  buf

  (
    G5298_p,
    g1531_p
  );


  buf

  (
    G5299_p,
    g1540_p
  );


  buf

  (
    G5300_p,
    g1549_p
  );


  buf

  (
    G5301_p,
    g1558_p
  );


  buf

  (
    G5302_p,
    g1568_p
  );


  buf

  (
    G5303_p,
    g1578_p
  );


  buf

  (
    G5304_p,
    g1588_p
  );


  buf

  (
    G5305_p,
    g1598_p
  );


  buf

  (
    G5306_p,
    g1608_p
  );


  buf

  (
    G5307_p,
    g1618_p
  );


  buf

  (
    G5308_p,
    g1628_p
  );


  buf

  (
    G5309_p,
    g1638_p
  );


  buf

  (
    G5310_p,
    g1642_p
  );


  buf

  (
    G5311_p,
    g1647_p
  );


  buf

  (
    G5312_n,
    g1660_n
  );


  buf

  (
    G5313_n,
    g1669_n
  );


  buf

  (
    G5314_p,
    g1679_n
  );


  buf

  (
    G5315_p,
    g1689_n
  );


  DROC
  ffc_0_0
  (
    .doutp(ffc_0_p),
    .doutn(ffc_0_n),
    .din(G1_p)
  );


  DROC
  ffc_1_1
  (
    .doutp(ffc_1_p),
    .doutn(ffc_1_n),
    .din(ffc_0_p)
  );


  DROC
  ffc_2_2
  (
    .doutp(ffc_2_p),
    .doutn(ffc_2_n),
    .din(ffc_1_p)
  );


  DROC
  ffc_3_3
  (
    .doutp(ffc_3_p),
    .doutn(ffc_3_n),
    .din(ffc_2_p)
  );


  DROC
  ffc_4_0
  (
    .doutp(ffc_4_p),
    .doutn(ffc_4_n),
    .din(G2_p)
  );


  DROC
  ffc_5_1
  (
    .doutp(ffc_5_p),
    .doutn(ffc_5_n),
    .din(ffc_4_p)
  );


  DROC
  ffc_6_2
  (
    .doutp(ffc_6_p),
    .doutn(ffc_6_n),
    .din(ffc_5_p)
  );


  DROC
  ffc_7_0
  (
    .doutp(ffc_7_p),
    .doutn(ffc_7_n),
    .din(G3_p)
  );


  DROC
  ffc_8_1
  (
    .doutp(ffc_8_p),
    .doutn(ffc_8_n),
    .din(ffc_7_p)
  );


  DROC
  ffc_9_2
  (
    .doutp(ffc_9_p),
    .doutn(ffc_9_n),
    .din(ffc_8_p)
  );


  DROC
  ffc_10_3
  (
    .doutp(ffc_10_p),
    .doutn(ffc_10_n),
    .din(ffc_9_p)
  );


  DROC
  ffc_11_0
  (
    .doutp(ffc_11_p),
    .doutn(ffc_11_n),
    .din(G4_p)
  );


  DROC
  ffc_12_1
  (
    .doutp(ffc_12_p),
    .doutn(ffc_12_n),
    .din(ffc_11_p)
  );


  DROC
  ffc_13_2
  (
    .doutp(ffc_13_p),
    .doutn(ffc_13_n),
    .din(ffc_12_p)
  );


  DROC
  ffc_14_3
  (
    .doutp(ffc_14_p),
    .doutn(ffc_14_n),
    .din(ffc_13_p)
  );


  DROC
  ffc_15_0
  (
    .doutp(ffc_15_p),
    .doutn(ffc_15_n),
    .din(G5_p)
  );


  DROC
  ffc_16_1
  (
    .doutp(ffc_16_p),
    .doutn(ffc_16_n),
    .din(ffc_15_p)
  );


  DROC
  ffc_17_2
  (
    .doutp(ffc_17_p),
    .doutn(ffc_17_n),
    .din(ffc_16_p)
  );


  DROC
  ffc_18_3
  (
    .doutp(ffc_18_p),
    .doutn(ffc_18_n),
    .din(ffc_17_p)
  );


  DROC
  ffc_19_0
  (
    .doutp(ffc_19_p),
    .doutn(ffc_19_n),
    .din(G6_p)
  );


  DROC
  ffc_20_1
  (
    .doutp(ffc_20_p),
    .doutn(ffc_20_n),
    .din(ffc_19_p)
  );


  DROC
  ffc_21_2
  (
    .doutp(ffc_21_p),
    .doutn(ffc_21_n),
    .din(ffc_20_p)
  );


  DROC
  ffc_22_3
  (
    .doutp(ffc_22_p),
    .doutn(ffc_22_n),
    .din(ffc_21_p)
  );


  DROC
  ffc_23_0
  (
    .doutp(ffc_23_p),
    .doutn(ffc_23_n),
    .din(G7_p)
  );


  DROC
  ffc_24_1
  (
    .doutp(ffc_24_p),
    .doutn(ffc_24_n),
    .din(ffc_23_p)
  );


  DROC
  ffc_25_2
  (
    .doutp(ffc_25_p),
    .doutn(ffc_25_n),
    .din(ffc_24_p)
  );


  DROC
  ffc_26_3
  (
    .doutp(ffc_26_p),
    .doutn(ffc_26_n),
    .din(ffc_25_p)
  );


  DROC
  ffc_27_0
  (
    .doutp(ffc_27_p),
    .doutn(ffc_27_n),
    .din(G8_p)
  );


  DROC
  ffc_28_1
  (
    .doutp(ffc_28_p),
    .doutn(ffc_28_n),
    .din(ffc_27_p)
  );


  DROC
  ffc_29_2
  (
    .doutp(ffc_29_p),
    .doutn(ffc_29_n),
    .din(ffc_28_p)
  );


  DROC
  ffc_30_3
  (
    .doutp(ffc_30_p),
    .doutn(ffc_30_n),
    .din(ffc_29_p)
  );


  DROC
  ffc_31_0
  (
    .doutp(ffc_31_p),
    .doutn(ffc_31_n),
    .din(G9_p)
  );


  DROC
  ffc_32_1
  (
    .doutp(ffc_32_p),
    .doutn(ffc_32_n),
    .din(ffc_31_p)
  );


  DROC
  ffc_33_2
  (
    .doutp(ffc_33_p),
    .doutn(ffc_33_n),
    .din(ffc_32_p)
  );


  DROC
  ffc_34_3
  (
    .doutp(ffc_34_p),
    .doutn(ffc_34_n),
    .din(ffc_33_p)
  );


  DROC
  ffc_35_0
  (
    .doutp(ffc_35_p),
    .doutn(ffc_35_n),
    .din(G10_p)
  );


  DROC
  ffc_36_1
  (
    .doutp(ffc_36_p),
    .doutn(ffc_36_n),
    .din(ffc_35_p)
  );


  DROC
  ffc_37_2
  (
    .doutp(ffc_37_p),
    .doutn(ffc_37_n),
    .din(ffc_36_p)
  );


  DROC
  ffc_38_3
  (
    .doutp(ffc_38_p),
    .doutn(ffc_38_n),
    .din(ffc_37_p)
  );


  DROC
  ffc_39_0
  (
    .doutp(ffc_39_p),
    .doutn(ffc_39_n),
    .din(G11_p)
  );


  DROC
  ffc_40_1
  (
    .doutp(ffc_40_p),
    .doutn(ffc_40_n),
    .din(ffc_39_p)
  );


  DROC
  ffc_41_2
  (
    .doutp(ffc_41_p),
    .doutn(ffc_41_n),
    .din(ffc_40_p)
  );


  DROC
  ffc_42_3
  (
    .doutp(ffc_42_p),
    .doutn(ffc_42_n),
    .din(ffc_41_p)
  );


  DROC
  ffc_43_0
  (
    .doutp(ffc_43_p),
    .doutn(ffc_43_n),
    .din(G12_p)
  );


  DROC
  ffc_44_1
  (
    .doutp(ffc_44_p),
    .doutn(ffc_44_n),
    .din(ffc_43_p)
  );


  DROC
  ffc_45_2
  (
    .doutp(ffc_45_p),
    .doutn(ffc_45_n),
    .din(ffc_44_p)
  );


  DROC
  ffc_46_3
  (
    .doutp(ffc_46_p),
    .doutn(ffc_46_n),
    .din(ffc_45_p)
  );


  DROC
  ffc_47_0
  (
    .doutp(ffc_47_p),
    .doutn(ffc_47_n),
    .din(G13_p)
  );


  DROC
  ffc_48_1
  (
    .doutp(ffc_48_p),
    .doutn(ffc_48_n),
    .din(ffc_47_p)
  );


  DROC
  ffc_49_2
  (
    .doutp(ffc_49_p),
    .doutn(ffc_49_n),
    .din(ffc_48_p)
  );


  DROC
  ffc_50_3
  (
    .doutp(ffc_50_p),
    .doutn(ffc_50_n),
    .din(ffc_49_p)
  );


  DROC
  ffc_51_0
  (
    .doutp(ffc_51_p),
    .doutn(ffc_51_n),
    .din(G14_p)
  );


  DROC
  ffc_52_1
  (
    .doutp(ffc_52_p),
    .doutn(ffc_52_n),
    .din(ffc_51_p)
  );


  DROC
  ffc_53_2
  (
    .doutp(ffc_53_p),
    .doutn(ffc_53_n),
    .din(ffc_52_p)
  );


  DROC
  ffc_54_3
  (
    .doutp(ffc_54_p),
    .doutn(ffc_54_n),
    .din(ffc_53_p)
  );


  DROC
  ffc_55_0
  (
    .doutp(ffc_55_p),
    .doutn(ffc_55_n),
    .din(G15_p)
  );


  DROC
  ffc_56_1
  (
    .doutp(ffc_56_p),
    .doutn(ffc_56_n),
    .din(ffc_55_p)
  );


  DROC
  ffc_57_2
  (
    .doutp(ffc_57_p),
    .doutn(ffc_57_n),
    .din(ffc_56_p)
  );


  DROC
  ffc_58_3
  (
    .doutp(ffc_58_p),
    .doutn(ffc_58_n),
    .din(ffc_57_p)
  );


  DROC
  ffc_59_0
  (
    .doutp(ffc_59_p),
    .doutn(ffc_59_n),
    .din(G16_p)
  );


  DROC
  ffc_60_1
  (
    .doutp(ffc_60_p),
    .doutn(ffc_60_n),
    .din(ffc_59_p)
  );


  DROC
  ffc_61_2
  (
    .doutp(ffc_61_p),
    .doutn(ffc_61_n),
    .din(ffc_60_p)
  );


  DROC
  ffc_62_3
  (
    .doutp(ffc_62_p),
    .doutn(ffc_62_n),
    .din(ffc_61_p)
  );


  DROC
  ffc_63_0
  (
    .doutp(ffc_63_p),
    .doutn(ffc_63_n),
    .din(G17_p)
  );


  DROC
  ffc_64_1
  (
    .doutp(ffc_64_p),
    .doutn(ffc_64_n),
    .din(ffc_63_p)
  );


  DROC
  ffc_65_2
  (
    .doutp(ffc_65_p),
    .doutn(ffc_65_n),
    .din(ffc_64_p)
  );


  DROC
  ffc_66_3
  (
    .doutp(ffc_66_p),
    .doutn(ffc_66_n),
    .din(ffc_65_p)
  );


  DROC
  ffc_67_0
  (
    .doutp(ffc_67_p),
    .doutn(ffc_67_n),
    .din(G18_p)
  );


  DROC
  ffc_68_1
  (
    .doutp(ffc_68_p),
    .doutn(ffc_68_n),
    .din(ffc_67_p)
  );


  DROC
  ffc_69_2
  (
    .doutp(ffc_69_p),
    .doutn(ffc_69_n),
    .din(ffc_68_p)
  );


  DROC
  ffc_70_3
  (
    .doutp(ffc_70_p),
    .doutn(ffc_70_n),
    .din(ffc_69_p)
  );


  DROC
  ffc_71_0
  (
    .doutp(ffc_71_p),
    .doutn(ffc_71_n),
    .din(G19_p)
  );


  DROC
  ffc_72_1
  (
    .doutp(ffc_72_p),
    .doutn(ffc_72_n),
    .din(ffc_71_p)
  );


  DROC
  ffc_73_2
  (
    .doutp(ffc_73_p),
    .doutn(ffc_73_n),
    .din(ffc_72_p)
  );


  DROC
  ffc_74_0
  (
    .doutp(ffc_74_p),
    .doutn(ffc_74_n),
    .din(G20_p)
  );


  DROC
  ffc_75_1
  (
    .doutp(ffc_75_p),
    .doutn(ffc_75_n),
    .din(ffc_74_p)
  );


  DROC
  ffc_76_2
  (
    .doutp(ffc_76_p),
    .doutn(ffc_76_n),
    .din(ffc_75_p)
  );


  DROC
  ffc_77_3
  (
    .doutp(ffc_77_p),
    .doutn(ffc_77_n),
    .din(ffc_76_p)
  );


  DROC
  ffc_78_0
  (
    .doutp(ffc_78_p),
    .doutn(ffc_78_n),
    .din(G21_p)
  );


  DROC
  ffc_79_1
  (
    .doutp(ffc_79_p),
    .doutn(ffc_79_n),
    .din(ffc_78_p)
  );


  DROC
  ffc_80_2
  (
    .doutp(ffc_80_p),
    .doutn(ffc_80_n),
    .din(ffc_79_p)
  );


  DROC
  ffc_81_0
  (
    .doutp(ffc_81_p),
    .doutn(ffc_81_n),
    .din(G22_p)
  );


  DROC
  ffc_82_1
  (
    .doutp(ffc_82_p),
    .doutn(ffc_82_n),
    .din(ffc_81_p)
  );


  DROC
  ffc_83_2
  (
    .doutp(ffc_83_p),
    .doutn(ffc_83_n),
    .din(ffc_82_p)
  );


  DROC
  ffc_84_3
  (
    .doutp(ffc_84_p),
    .doutn(ffc_84_n),
    .din(ffc_83_p)
  );


  DROC
  ffc_85_0
  (
    .doutp(ffc_85_p),
    .doutn(ffc_85_n),
    .din(G23_p)
  );


  DROC
  ffc_86_1
  (
    .doutp(ffc_86_p),
    .doutn(ffc_86_n),
    .din(ffc_85_p)
  );


  DROC
  ffc_87_2
  (
    .doutp(ffc_87_p),
    .doutn(ffc_87_n),
    .din(ffc_86_p)
  );


  DROC
  ffc_88_3
  (
    .doutp(ffc_88_p),
    .doutn(ffc_88_n),
    .din(ffc_87_p)
  );


  DROC
  ffc_89_0
  (
    .doutp(ffc_89_p),
    .doutn(ffc_89_n),
    .din(G24_p)
  );


  DROC
  ffc_90_1
  (
    .doutp(ffc_90_p),
    .doutn(ffc_90_n),
    .din(ffc_89_p)
  );


  DROC
  ffc_91_2
  (
    .doutp(ffc_91_p),
    .doutn(ffc_91_n),
    .din(ffc_90_p)
  );


  DROC
  ffc_92_3
  (
    .doutp(ffc_92_p),
    .doutn(ffc_92_n),
    .din(ffc_91_p)
  );


  DROC
  ffc_93_0
  (
    .doutp(ffc_93_p),
    .doutn(ffc_93_n),
    .din(G25_p)
  );


  DROC
  ffc_94_1
  (
    .doutp(ffc_94_p),
    .doutn(ffc_94_n),
    .din(ffc_93_p)
  );


  DROC
  ffc_95_2
  (
    .doutp(ffc_95_p),
    .doutn(ffc_95_n),
    .din(ffc_94_p)
  );


  DROC
  ffc_96_3
  (
    .doutp(ffc_96_p),
    .doutn(ffc_96_n),
    .din(ffc_95_p)
  );


  DROC
  ffc_97_0
  (
    .doutp(ffc_97_p),
    .doutn(ffc_97_n),
    .din(G26_p)
  );


  DROC
  ffc_98_1
  (
    .doutp(ffc_98_p),
    .doutn(ffc_98_n),
    .din(ffc_97_p)
  );


  DROC
  ffc_99_2
  (
    .doutp(ffc_99_p),
    .doutn(ffc_99_n),
    .din(ffc_98_p)
  );


  DROC
  ffc_100_3
  (
    .doutp(ffc_100_p),
    .doutn(ffc_100_n),
    .din(ffc_99_p)
  );


  DROC
  ffc_101_0
  (
    .doutp(ffc_101_p),
    .doutn(ffc_101_n),
    .din(G27_p)
  );


  DROC
  ffc_102_1
  (
    .doutp(ffc_102_p),
    .doutn(ffc_102_n),
    .din(ffc_101_p)
  );


  DROC
  ffc_103_2
  (
    .doutp(ffc_103_p),
    .doutn(ffc_103_n),
    .din(ffc_102_p)
  );


  DROC
  ffc_104_3
  (
    .doutp(ffc_104_p),
    .doutn(ffc_104_n),
    .din(ffc_103_p)
  );


  DROC
  ffc_105_0
  (
    .doutp(ffc_105_p),
    .doutn(ffc_105_n),
    .din(G28_p)
  );


  DROC
  ffc_106_1
  (
    .doutp(ffc_106_p),
    .doutn(ffc_106_n),
    .din(ffc_105_p)
  );


  DROC
  ffc_107_2
  (
    .doutp(ffc_107_p),
    .doutn(ffc_107_n),
    .din(ffc_106_p)
  );


  DROC
  ffc_108_3
  (
    .doutp(ffc_108_p),
    .doutn(ffc_108_n),
    .din(ffc_107_p)
  );


  DROC
  ffc_109_0
  (
    .doutp(ffc_109_p),
    .doutn(ffc_109_n),
    .din(G29_p)
  );


  DROC
  ffc_110_1
  (
    .doutp(ffc_110_p),
    .doutn(ffc_110_n),
    .din(ffc_109_p)
  );


  DROC
  ffc_111_2
  (
    .doutp(ffc_111_p),
    .doutn(ffc_111_n),
    .din(ffc_110_p)
  );


  DROC
  ffc_112_3
  (
    .doutp(ffc_112_p),
    .doutn(ffc_112_n),
    .din(ffc_111_p)
  );


  DROC
  ffc_113_0
  (
    .doutp(ffc_113_p),
    .doutn(ffc_113_n),
    .din(G30_p)
  );


  DROC
  ffc_114_1
  (
    .doutp(ffc_114_p),
    .doutn(ffc_114_n),
    .din(ffc_113_p)
  );


  DROC
  ffc_115_2
  (
    .doutp(ffc_115_p),
    .doutn(ffc_115_n),
    .din(ffc_114_p)
  );


  DROC
  ffc_116_3
  (
    .doutp(ffc_116_p),
    .doutn(ffc_116_n),
    .din(ffc_115_p)
  );


  DROC
  ffc_117_0
  (
    .doutp(ffc_117_p),
    .doutn(ffc_117_n),
    .din(G31_p)
  );


  DROC
  ffc_118_1
  (
    .doutp(ffc_118_p),
    .doutn(ffc_118_n),
    .din(ffc_117_p)
  );


  DROC
  ffc_119_2
  (
    .doutp(ffc_119_p),
    .doutn(ffc_119_n),
    .din(ffc_118_p)
  );


  DROC
  ffc_120_3
  (
    .doutp(ffc_120_p),
    .doutn(ffc_120_n),
    .din(ffc_119_p)
  );


  DROC
  ffc_121_0
  (
    .doutp(ffc_121_p),
    .doutn(ffc_121_n),
    .din(G32_p)
  );


  DROC
  ffc_122_1
  (
    .doutp(ffc_122_p),
    .doutn(ffc_122_n),
    .din(ffc_121_p)
  );


  DROC
  ffc_123_2
  (
    .doutp(ffc_123_p),
    .doutn(ffc_123_n),
    .din(ffc_122_p)
  );


  DROC
  ffc_124_3
  (
    .doutp(ffc_124_p),
    .doutn(ffc_124_n),
    .din(ffc_123_p)
  );


  DROC
  ffc_125_0
  (
    .doutp(ffc_125_p),
    .doutn(ffc_125_n),
    .din(G33_p)
  );


  DROC
  ffc_126_1
  (
    .doutp(ffc_126_p),
    .doutn(ffc_126_n),
    .din(ffc_125_p)
  );


  DROC
  ffc_127_2
  (
    .doutp(ffc_127_p),
    .doutn(ffc_127_n),
    .din(ffc_126_p)
  );


  DROC
  ffc_128_3
  (
    .doutp(ffc_128_p),
    .doutn(ffc_128_n),
    .din(ffc_127_p)
  );


  DROC
  ffc_129_0
  (
    .doutp(ffc_129_p),
    .doutn(ffc_129_n),
    .din(G34_p)
  );


  DROC
  ffc_130_1
  (
    .doutp(ffc_130_p),
    .doutn(ffc_130_n),
    .din(ffc_129_p)
  );


  DROC
  ffc_131_2
  (
    .doutp(ffc_131_p),
    .doutn(ffc_131_n),
    .din(ffc_130_p)
  );


  DROC
  ffc_132_3
  (
    .doutp(ffc_132_p),
    .doutn(ffc_132_n),
    .din(ffc_131_p)
  );


  DROC
  ffc_133_0
  (
    .doutp(ffc_133_p),
    .doutn(ffc_133_n),
    .din(G35_p)
  );


  DROC
  ffc_134_1
  (
    .doutp(ffc_134_p),
    .doutn(ffc_134_n),
    .din(ffc_133_p)
  );


  DROC
  ffc_135_2
  (
    .doutp(ffc_135_p),
    .doutn(ffc_135_n),
    .din(ffc_134_p)
  );


  DROC
  ffc_136_3
  (
    .doutp(ffc_136_p),
    .doutn(ffc_136_n),
    .din(ffc_135_p)
  );


  DROC
  ffc_137_0
  (
    .doutp(ffc_137_p),
    .doutn(ffc_137_n),
    .din(G36_p)
  );


  DROC
  ffc_138_1
  (
    .doutp(ffc_138_p),
    .doutn(ffc_138_n),
    .din(ffc_137_p)
  );


  DROC
  ffc_139_2
  (
    .doutp(ffc_139_p),
    .doutn(ffc_139_n),
    .din(ffc_138_p)
  );


  DROC
  ffc_140_3
  (
    .doutp(ffc_140_p),
    .doutn(ffc_140_n),
    .din(ffc_139_p)
  );


  DROC
  ffc_141_0
  (
    .doutp(ffc_141_p),
    .doutn(ffc_141_n),
    .din(G37_p)
  );


  DROC
  ffc_142_1
  (
    .doutp(ffc_142_p),
    .doutn(ffc_142_n),
    .din(ffc_141_p)
  );


  DROC
  ffc_143_2
  (
    .doutp(ffc_143_p),
    .doutn(ffc_143_n),
    .din(ffc_142_p)
  );


  DROC
  ffc_144_3
  (
    .doutp(ffc_144_p),
    .doutn(ffc_144_n),
    .din(ffc_143_p)
  );


  DROC
  ffc_145_0
  (
    .doutp(ffc_145_p),
    .doutn(ffc_145_n),
    .din(G38_p)
  );


  DROC
  ffc_146_1
  (
    .doutp(ffc_146_p),
    .doutn(ffc_146_n),
    .din(ffc_145_p)
  );


  DROC
  ffc_147_2
  (
    .doutp(ffc_147_p),
    .doutn(ffc_147_n),
    .din(ffc_146_p)
  );


  DROC
  ffc_148_3
  (
    .doutp(ffc_148_p),
    .doutn(ffc_148_n),
    .din(ffc_147_p)
  );


  DROC
  ffc_149_0
  (
    .doutp(ffc_149_p),
    .doutn(ffc_149_n),
    .din(G39_p)
  );


  DROC
  ffc_150_1
  (
    .doutp(ffc_150_p),
    .doutn(ffc_150_n),
    .din(ffc_149_p)
  );


  DROC
  ffc_151_2
  (
    .doutp(ffc_151_p),
    .doutn(ffc_151_n),
    .din(ffc_150_p)
  );


  DROC
  ffc_152_3
  (
    .doutp(ffc_152_p),
    .doutn(ffc_152_n),
    .din(ffc_151_p)
  );


  DROC
  ffc_153_0
  (
    .doutp(ffc_153_p),
    .doutn(ffc_153_n),
    .din(G40_p)
  );


  DROC
  ffc_154_1
  (
    .doutp(ffc_154_p),
    .doutn(ffc_154_n),
    .din(ffc_153_p)
  );


  DROC
  ffc_155_2
  (
    .doutp(ffc_155_p),
    .doutn(ffc_155_n),
    .din(ffc_154_p)
  );


  DROC
  ffc_156_3
  (
    .doutp(ffc_156_p),
    .doutn(ffc_156_n),
    .din(ffc_155_p)
  );


  DROC
  ffc_157_0
  (
    .doutp(ffc_157_p),
    .doutn(ffc_157_n),
    .din(G41_p)
  );


  DROC
  ffc_158_1
  (
    .doutp(ffc_158_p),
    .doutn(ffc_158_n),
    .din(ffc_157_p)
  );


  DROC
  ffc_159_2
  (
    .doutp(ffc_159_p),
    .doutn(ffc_159_n),
    .din(ffc_158_p)
  );


  DROC
  ffc_160_3
  (
    .doutp(ffc_160_p),
    .doutn(ffc_160_n),
    .din(ffc_159_p)
  );


  DROC
  ffc_161_0
  (
    .doutp(ffc_161_p),
    .doutn(ffc_161_n),
    .din(G42_p)
  );


  DROC
  ffc_162_1
  (
    .doutp(ffc_162_p),
    .doutn(ffc_162_n),
    .din(ffc_161_p)
  );


  DROC
  ffc_163_2
  (
    .doutp(ffc_163_p),
    .doutn(ffc_163_n),
    .din(ffc_162_p)
  );


  DROC
  ffc_164_3
  (
    .doutp(ffc_164_p),
    .doutn(ffc_164_n),
    .din(ffc_163_p)
  );


  DROC
  ffc_165_0
  (
    .doutp(ffc_165_p),
    .doutn(ffc_165_n),
    .din(G43_p)
  );


  DROC
  ffc_166_1
  (
    .doutp(ffc_166_p),
    .doutn(ffc_166_n),
    .din(ffc_165_p)
  );


  DROC
  ffc_167_2
  (
    .doutp(ffc_167_p),
    .doutn(ffc_167_n),
    .din(ffc_166_p)
  );


  DROC
  ffc_168_0
  (
    .doutp(ffc_168_p),
    .doutn(ffc_168_n),
    .din(G44_p)
  );


  DROC
  ffc_169_1
  (
    .doutp(ffc_169_p),
    .doutn(ffc_169_n),
    .din(ffc_168_p)
  );


  DROC
  ffc_170_2
  (
    .doutp(ffc_170_p),
    .doutn(ffc_170_n),
    .din(ffc_169_p)
  );


  DROC
  ffc_171_0
  (
    .doutp(ffc_171_p),
    .doutn(ffc_171_n),
    .din(G45_p)
  );


  DROC
  ffc_172_1
  (
    .doutp(ffc_172_p),
    .doutn(ffc_172_n),
    .din(ffc_171_p)
  );


  DROC
  ffc_173_2
  (
    .doutp(ffc_173_p),
    .doutn(ffc_173_n),
    .din(ffc_172_p)
  );


  DROC
  ffc_174_3
  (
    .doutp(ffc_174_p),
    .doutn(ffc_174_n),
    .din(ffc_173_p)
  );


  DROC
  ffc_175_0
  (
    .doutp(ffc_175_p),
    .doutn(ffc_175_n),
    .din(G46_p)
  );


  DROC
  ffc_176_1
  (
    .doutp(ffc_176_p),
    .doutn(ffc_176_n),
    .din(ffc_175_p)
  );


  DROC
  ffc_177_2
  (
    .doutp(ffc_177_p),
    .doutn(ffc_177_n),
    .din(ffc_176_p)
  );


  DROC
  ffc_178_0
  (
    .doutp(ffc_178_p),
    .doutn(ffc_178_n),
    .din(G47_p)
  );


  DROC
  ffc_179_1
  (
    .doutp(ffc_179_p),
    .doutn(ffc_179_n),
    .din(ffc_178_p)
  );


  DROC
  ffc_180_2
  (
    .doutp(ffc_180_p),
    .doutn(ffc_180_n),
    .din(ffc_179_p)
  );


  DROC
  ffc_181_0
  (
    .doutp(ffc_181_p),
    .doutn(ffc_181_n),
    .din(G48_p)
  );


  DROC
  ffc_182_1
  (
    .doutp(ffc_182_p),
    .doutn(ffc_182_n),
    .din(ffc_181_p)
  );


  DROC
  ffc_183_2
  (
    .doutp(ffc_183_p),
    .doutn(ffc_183_n),
    .din(ffc_182_p)
  );


  DROC
  ffc_184_0
  (
    .doutp(ffc_184_p),
    .doutn(ffc_184_n),
    .din(G49_p)
  );


  DROC
  ffc_185_1
  (
    .doutp(ffc_185_p),
    .doutn(ffc_185_n),
    .din(ffc_184_p)
  );


  DROC
  ffc_186_2
  (
    .doutp(ffc_186_p),
    .doutn(ffc_186_n),
    .din(ffc_185_p)
  );


  DROC
  ffc_187_3
  (
    .doutp(ffc_187_p),
    .doutn(ffc_187_n),
    .din(ffc_186_p)
  );


  DROC
  ffc_188_0
  (
    .doutp(ffc_188_p),
    .doutn(ffc_188_n),
    .din(G50_p)
  );


  DROC
  ffc_189_1
  (
    .doutp(ffc_189_p),
    .doutn(ffc_189_n),
    .din(ffc_188_p)
  );


  DROC
  ffc_190_2
  (
    .doutp(ffc_190_p),
    .doutn(ffc_190_n),
    .din(ffc_189_p)
  );


  DROC
  ffc_191_0
  (
    .doutp(ffc_191_p),
    .doutn(ffc_191_n),
    .din(G51_p)
  );


  DROC
  ffc_192_1
  (
    .doutp(ffc_192_p),
    .doutn(ffc_192_n),
    .din(ffc_191_p)
  );


  DROC
  ffc_193_2
  (
    .doutp(ffc_193_p),
    .doutn(ffc_193_n),
    .din(ffc_192_p)
  );


  DROC
  ffc_194_3
  (
    .doutp(ffc_194_p),
    .doutn(ffc_194_n),
    .din(ffc_193_p)
  );


  DROC
  ffc_195_0
  (
    .doutp(ffc_195_p),
    .doutn(ffc_195_n),
    .din(G52_p)
  );


  DROC
  ffc_196_1
  (
    .doutp(ffc_196_p),
    .doutn(ffc_196_n),
    .din(ffc_195_p)
  );


  DROC
  ffc_197_2
  (
    .doutp(ffc_197_p),
    .doutn(ffc_197_n),
    .din(ffc_196_p)
  );


  DROC
  ffc_198_0
  (
    .doutp(ffc_198_p),
    .doutn(ffc_198_n),
    .din(G53_p)
  );


  DROC
  ffc_199_1
  (
    .doutp(ffc_199_p),
    .doutn(ffc_199_n),
    .din(ffc_198_p)
  );


  DROC
  ffc_200_2
  (
    .doutp(ffc_200_p),
    .doutn(ffc_200_n),
    .din(ffc_199_p)
  );


  DROC
  ffc_201_3
  (
    .doutp(ffc_201_p),
    .doutn(ffc_201_n),
    .din(ffc_200_p)
  );


  DROC
  ffc_202_0
  (
    .doutp(ffc_202_p),
    .doutn(ffc_202_n),
    .din(G54_p)
  );


  DROC
  ffc_203_1
  (
    .doutp(ffc_203_p),
    .doutn(ffc_203_n),
    .din(ffc_202_p)
  );


  DROC
  ffc_204_2
  (
    .doutp(ffc_204_p),
    .doutn(ffc_204_n),
    .din(ffc_203_p)
  );


  DROC
  ffc_205_3
  (
    .doutp(ffc_205_p),
    .doutn(ffc_205_n),
    .din(ffc_204_p_spl_)
  );


  DROC
  ffc_206_0
  (
    .doutp(ffc_206_p),
    .doutn(ffc_206_n),
    .din(G55_p)
  );


  DROC
  ffc_207_1
  (
    .doutp(ffc_207_p),
    .doutn(ffc_207_n),
    .din(ffc_206_p)
  );


  DROC
  ffc_208_2
  (
    .doutp(ffc_208_p),
    .doutn(ffc_208_n),
    .din(ffc_207_p)
  );


  DROC
  ffc_209_3
  (
    .doutp(ffc_209_p),
    .doutn(ffc_209_n),
    .din(ffc_208_p)
  );


  DROC
  ffc_210_0
  (
    .doutp(ffc_210_p),
    .doutn(ffc_210_n),
    .din(G56_p)
  );


  DROC
  ffc_211_1
  (
    .doutp(ffc_211_p),
    .doutn(ffc_211_n),
    .din(ffc_210_p)
  );


  DROC
  ffc_212_2
  (
    .doutp(ffc_212_p),
    .doutn(ffc_212_n),
    .din(ffc_211_p)
  );


  DROC
  ffc_213_3
  (
    .doutp(ffc_213_p),
    .doutn(ffc_213_n),
    .din(ffc_212_p)
  );


  DROC
  ffc_214_0
  (
    .doutp(ffc_214_p),
    .doutn(ffc_214_n),
    .din(G57_p)
  );


  DROC
  ffc_215_1
  (
    .doutp(ffc_215_p),
    .doutn(ffc_215_n),
    .din(ffc_214_p)
  );


  DROC
  ffc_216_2
  (
    .doutp(ffc_216_p),
    .doutn(ffc_216_n),
    .din(ffc_215_p)
  );


  DROC
  ffc_217_0
  (
    .doutp(ffc_217_p),
    .doutn(ffc_217_n),
    .din(G58_p)
  );


  DROC
  ffc_218_1
  (
    .doutp(ffc_218_p),
    .doutn(ffc_218_n),
    .din(ffc_217_p)
  );


  DROC
  ffc_219_2
  (
    .doutp(ffc_219_p),
    .doutn(ffc_219_n),
    .din(ffc_218_p)
  );


  DROC
  ffc_220_0
  (
    .doutp(ffc_220_p),
    .doutn(ffc_220_n),
    .din(G59_p)
  );


  DROC
  ffc_221_1
  (
    .doutp(ffc_221_p),
    .doutn(ffc_221_n),
    .din(ffc_220_p)
  );


  DROC
  ffc_222_2
  (
    .doutp(ffc_222_p),
    .doutn(ffc_222_n),
    .din(ffc_221_p)
  );


  DROC
  ffc_223_0
  (
    .doutp(ffc_223_p),
    .doutn(ffc_223_n),
    .din(G60_p)
  );


  DROC
  ffc_224_1
  (
    .doutp(ffc_224_p),
    .doutn(ffc_224_n),
    .din(ffc_223_p)
  );


  DROC
  ffc_225_2
  (
    .doutp(ffc_225_p),
    .doutn(ffc_225_n),
    .din(ffc_224_p)
  );


  DROC
  ffc_226_0
  (
    .doutp(ffc_226_p),
    .doutn(ffc_226_n),
    .din(G61_p)
  );


  DROC
  ffc_227_1
  (
    .doutp(ffc_227_p),
    .doutn(ffc_227_n),
    .din(ffc_226_p)
  );


  DROC
  ffc_228_2
  (
    .doutp(ffc_228_p),
    .doutn(ffc_228_n),
    .din(ffc_227_p)
  );


  DROC
  ffc_229_3
  (
    .doutp(ffc_229_p),
    .doutn(ffc_229_n),
    .din(ffc_228_p)
  );


  DROC
  ffc_230_0
  (
    .doutp(ffc_230_p),
    .doutn(ffc_230_n),
    .din(G62_p)
  );


  DROC
  ffc_231_1
  (
    .doutp(ffc_231_p),
    .doutn(ffc_231_n),
    .din(ffc_230_p)
  );


  DROC
  ffc_232_2
  (
    .doutp(ffc_232_p),
    .doutn(ffc_232_n),
    .din(ffc_231_p)
  );


  DROC
  ffc_233_3
  (
    .doutp(ffc_233_p),
    .doutn(ffc_233_n),
    .din(ffc_232_p)
  );


  DROC
  ffc_234_0
  (
    .doutp(ffc_234_p),
    .doutn(ffc_234_n),
    .din(G63_p)
  );


  DROC
  ffc_235_1
  (
    .doutp(ffc_235_p),
    .doutn(ffc_235_n),
    .din(ffc_234_p)
  );


  DROC
  ffc_236_2
  (
    .doutp(ffc_236_p),
    .doutn(ffc_236_n),
    .din(ffc_235_p)
  );


  DROC
  ffc_237_3
  (
    .doutp(ffc_237_p),
    .doutn(ffc_237_n),
    .din(ffc_236_p)
  );


  DROC
  ffc_238_0
  (
    .doutp(ffc_238_p),
    .doutn(ffc_238_n),
    .din(G64_p)
  );


  DROC
  ffc_239_1
  (
    .doutp(ffc_239_p),
    .doutn(ffc_239_n),
    .din(ffc_238_p)
  );


  DROC
  ffc_240_2
  (
    .doutp(ffc_240_p),
    .doutn(ffc_240_n),
    .din(ffc_239_p)
  );


  DROC
  ffc_241_3
  (
    .doutp(ffc_241_p),
    .doutn(ffc_241_n),
    .din(ffc_240_p)
  );


  DROC
  ffc_242_0
  (
    .doutp(ffc_242_p),
    .doutn(ffc_242_n),
    .din(G65_p)
  );


  DROC
  ffc_243_1
  (
    .doutp(ffc_243_p),
    .doutn(ffc_243_n),
    .din(ffc_242_p)
  );


  DROC
  ffc_244_2
  (
    .doutp(ffc_244_p),
    .doutn(ffc_244_n),
    .din(ffc_243_p)
  );


  DROC
  ffc_245_3
  (
    .doutp(ffc_245_p),
    .doutn(ffc_245_n),
    .din(ffc_244_p)
  );


  DROC
  ffc_246_0
  (
    .doutp(ffc_246_p),
    .doutn(ffc_246_n),
    .din(G66_p)
  );


  DROC
  ffc_247_1
  (
    .doutp(ffc_247_p),
    .doutn(ffc_247_n),
    .din(ffc_246_p)
  );


  DROC
  ffc_248_2
  (
    .doutp(ffc_248_p),
    .doutn(ffc_248_n),
    .din(ffc_247_p)
  );


  DROC
  ffc_249_3
  (
    .doutp(ffc_249_p),
    .doutn(ffc_249_n),
    .din(ffc_248_p)
  );


  DROC
  ffc_250_0
  (
    .doutp(ffc_250_p),
    .doutn(ffc_250_n),
    .din(G67_p)
  );


  DROC
  ffc_251_1
  (
    .doutp(ffc_251_p),
    .doutn(ffc_251_n),
    .din(ffc_250_p)
  );


  DROC
  ffc_252_2
  (
    .doutp(ffc_252_p),
    .doutn(ffc_252_n),
    .din(ffc_251_p)
  );


  DROC
  ffc_253_3
  (
    .doutp(ffc_253_p),
    .doutn(ffc_253_n),
    .din(ffc_252_p)
  );


  DROC
  ffc_254_0
  (
    .doutp(ffc_254_p),
    .doutn(ffc_254_n),
    .din(G68_p)
  );


  DROC
  ffc_255_1
  (
    .doutp(ffc_255_p),
    .doutn(ffc_255_n),
    .din(ffc_254_p)
  );


  DROC
  ffc_256_2
  (
    .doutp(ffc_256_p),
    .doutn(ffc_256_n),
    .din(ffc_255_p)
  );


  DROC
  ffc_257_3
  (
    .doutp(ffc_257_p),
    .doutn(ffc_257_n),
    .din(ffc_256_p)
  );


  DROC
  ffc_258_0
  (
    .doutp(ffc_258_p),
    .doutn(ffc_258_n),
    .din(G69_p)
  );


  DROC
  ffc_259_1
  (
    .doutp(ffc_259_p),
    .doutn(ffc_259_n),
    .din(ffc_258_p)
  );


  DROC
  ffc_260_2
  (
    .doutp(ffc_260_p),
    .doutn(ffc_260_n),
    .din(ffc_259_p)
  );


  DROC
  ffc_261_3
  (
    .doutp(ffc_261_p),
    .doutn(ffc_261_n),
    .din(ffc_260_p)
  );


  DROC
  ffc_262_0
  (
    .doutp(ffc_262_p),
    .doutn(ffc_262_n),
    .din(G70_p)
  );


  DROC
  ffc_263_1
  (
    .doutp(ffc_263_p),
    .doutn(ffc_263_n),
    .din(ffc_262_p)
  );


  DROC
  ffc_264_2
  (
    .doutp(ffc_264_p),
    .doutn(ffc_264_n),
    .din(ffc_263_p)
  );


  DROC
  ffc_265_3
  (
    .doutp(ffc_265_p),
    .doutn(ffc_265_n),
    .din(ffc_264_p)
  );


  DROC
  ffc_266_0
  (
    .doutp(ffc_266_p),
    .doutn(ffc_266_n),
    .din(G71_p)
  );


  DROC
  ffc_267_1
  (
    .doutp(ffc_267_p),
    .doutn(ffc_267_n),
    .din(ffc_266_p)
  );


  DROC
  ffc_268_2
  (
    .doutp(ffc_268_p),
    .doutn(ffc_268_n),
    .din(ffc_267_p)
  );


  DROC
  ffc_269_3
  (
    .doutp(ffc_269_p),
    .doutn(ffc_269_n),
    .din(ffc_268_p)
  );


  DROC
  ffc_270_0
  (
    .doutp(ffc_270_p),
    .doutn(ffc_270_n),
    .din(G72_p)
  );


  DROC
  ffc_271_1
  (
    .doutp(ffc_271_p),
    .doutn(ffc_271_n),
    .din(ffc_270_p)
  );


  DROC
  ffc_272_2
  (
    .doutp(ffc_272_p),
    .doutn(ffc_272_n),
    .din(ffc_271_p)
  );


  DROC
  ffc_273_3
  (
    .doutp(ffc_273_p),
    .doutn(ffc_273_n),
    .din(ffc_272_p)
  );


  DROC
  ffc_274_0
  (
    .doutp(ffc_274_p),
    .doutn(ffc_274_n),
    .din(G73_p)
  );


  DROC
  ffc_275_1
  (
    .doutp(ffc_275_p),
    .doutn(ffc_275_n),
    .din(ffc_274_p)
  );


  DROC
  ffc_276_2
  (
    .doutp(ffc_276_p),
    .doutn(ffc_276_n),
    .din(ffc_275_p)
  );


  DROC
  ffc_277_3
  (
    .doutp(ffc_277_p),
    .doutn(ffc_277_n),
    .din(ffc_276_p)
  );


  DROC
  ffc_278_0
  (
    .doutp(ffc_278_p),
    .doutn(ffc_278_n),
    .din(G74_p)
  );


  DROC
  ffc_279_1
  (
    .doutp(ffc_279_p),
    .doutn(ffc_279_n),
    .din(ffc_278_p)
  );


  DROC
  ffc_280_2
  (
    .doutp(ffc_280_p),
    .doutn(ffc_280_n),
    .din(ffc_279_p)
  );


  DROC
  ffc_281_3
  (
    .doutp(ffc_281_p),
    .doutn(ffc_281_n),
    .din(ffc_280_p)
  );


  DROC
  ffc_282_0
  (
    .doutp(ffc_282_p),
    .doutn(ffc_282_n),
    .din(G75_p)
  );


  DROC
  ffc_283_1
  (
    .doutp(ffc_283_p),
    .doutn(ffc_283_n),
    .din(ffc_282_p)
  );


  DROC
  ffc_284_2
  (
    .doutp(ffc_284_p),
    .doutn(ffc_284_n),
    .din(ffc_283_p)
  );


  DROC
  ffc_285_3
  (
    .doutp(ffc_285_p),
    .doutn(ffc_285_n),
    .din(ffc_284_p)
  );


  DROC
  ffc_286_0
  (
    .doutp(ffc_286_p),
    .doutn(ffc_286_n),
    .din(G76_p)
  );


  DROC
  ffc_287_1
  (
    .doutp(ffc_287_p),
    .doutn(ffc_287_n),
    .din(ffc_286_p)
  );


  DROC
  ffc_288_2
  (
    .doutp(ffc_288_p),
    .doutn(ffc_288_n),
    .din(ffc_287_p)
  );


  DROC
  ffc_289_3
  (
    .doutp(ffc_289_p),
    .doutn(ffc_289_n),
    .din(ffc_288_p)
  );


  DROC
  ffc_290_0
  (
    .doutp(ffc_290_p),
    .doutn(ffc_290_n),
    .din(G77_p)
  );


  DROC
  ffc_291_1
  (
    .doutp(ffc_291_p),
    .doutn(ffc_291_n),
    .din(ffc_290_p)
  );


  DROC
  ffc_292_2
  (
    .doutp(ffc_292_p),
    .doutn(ffc_292_n),
    .din(ffc_291_p)
  );


  DROC
  ffc_293_3
  (
    .doutp(ffc_293_p),
    .doutn(ffc_293_n),
    .din(ffc_292_p)
  );


  DROC
  ffc_294_0
  (
    .doutp(ffc_294_p),
    .doutn(ffc_294_n),
    .din(G78_p)
  );


  DROC
  ffc_295_1
  (
    .doutp(ffc_295_p),
    .doutn(ffc_295_n),
    .din(ffc_294_p)
  );


  DROC
  ffc_296_2
  (
    .doutp(ffc_296_p),
    .doutn(ffc_296_n),
    .din(ffc_295_p)
  );


  DROC
  ffc_297_3
  (
    .doutp(ffc_297_p),
    .doutn(ffc_297_n),
    .din(ffc_296_p)
  );


  DROC
  ffc_298_0
  (
    .doutp(ffc_298_p),
    .doutn(ffc_298_n),
    .din(G79_p)
  );


  DROC
  ffc_299_1
  (
    .doutp(ffc_299_p),
    .doutn(ffc_299_n),
    .din(ffc_298_p)
  );


  DROC
  ffc_300_2
  (
    .doutp(ffc_300_p),
    .doutn(ffc_300_n),
    .din(ffc_299_p)
  );


  DROC
  ffc_301_3
  (
    .doutp(ffc_301_p),
    .doutn(ffc_301_n),
    .din(ffc_300_p)
  );


  DROC
  ffc_302_0
  (
    .doutp(ffc_302_p),
    .doutn(ffc_302_n),
    .din(G80_p)
  );


  DROC
  ffc_303_1
  (
    .doutp(ffc_303_p),
    .doutn(ffc_303_n),
    .din(ffc_302_p)
  );


  DROC
  ffc_304_2
  (
    .doutp(ffc_304_p),
    .doutn(ffc_304_n),
    .din(ffc_303_p)
  );


  DROC
  ffc_305_3
  (
    .doutp(ffc_305_p),
    .doutn(ffc_305_n),
    .din(ffc_304_p)
  );


  DROC
  ffc_306_0
  (
    .doutp(ffc_306_p),
    .doutn(ffc_306_n),
    .din(G81_p)
  );


  DROC
  ffc_307_1
  (
    .doutp(ffc_307_p),
    .doutn(ffc_307_n),
    .din(ffc_306_p)
  );


  DROC
  ffc_308_2
  (
    .doutp(ffc_308_p),
    .doutn(ffc_308_n),
    .din(ffc_307_p)
  );


  DROC
  ffc_309_3
  (
    .doutp(ffc_309_p),
    .doutn(ffc_309_n),
    .din(ffc_308_p)
  );


  DROC
  ffc_310_0
  (
    .doutp(ffc_310_p),
    .doutn(ffc_310_n),
    .din(G82_p)
  );


  DROC
  ffc_311_1
  (
    .doutp(ffc_311_p),
    .doutn(ffc_311_n),
    .din(ffc_310_p)
  );


  DROC
  ffc_312_2
  (
    .doutp(ffc_312_p),
    .doutn(ffc_312_n),
    .din(ffc_311_p)
  );


  DROC
  ffc_313_3
  (
    .doutp(ffc_313_p),
    .doutn(ffc_313_n),
    .din(ffc_312_p)
  );


  DROC
  ffc_314_0
  (
    .doutp(ffc_314_p),
    .doutn(ffc_314_n),
    .din(G83_p)
  );


  DROC
  ffc_315_1
  (
    .doutp(ffc_315_p),
    .doutn(ffc_315_n),
    .din(ffc_314_p)
  );


  DROC
  ffc_316_2
  (
    .doutp(ffc_316_p),
    .doutn(ffc_316_n),
    .din(ffc_315_p)
  );


  DROC
  ffc_317_3
  (
    .doutp(ffc_317_p),
    .doutn(ffc_317_n),
    .din(ffc_316_p)
  );


  DROC
  ffc_318_0
  (
    .doutp(ffc_318_p),
    .doutn(ffc_318_n),
    .din(G84_p)
  );


  DROC
  ffc_319_1
  (
    .doutp(ffc_319_p),
    .doutn(ffc_319_n),
    .din(ffc_318_p)
  );


  DROC
  ffc_320_2
  (
    .doutp(ffc_320_p),
    .doutn(ffc_320_n),
    .din(ffc_319_p)
  );


  DROC
  ffc_321_3
  (
    .doutp(ffc_321_p),
    .doutn(ffc_321_n),
    .din(ffc_320_p)
  );


  DROC
  ffc_322_0
  (
    .doutp(ffc_322_p),
    .doutn(ffc_322_n),
    .din(G85_p)
  );


  DROC
  ffc_323_1
  (
    .doutp(ffc_323_p),
    .doutn(ffc_323_n),
    .din(ffc_322_p)
  );


  DROC
  ffc_324_2
  (
    .doutp(ffc_324_p),
    .doutn(ffc_324_n),
    .din(ffc_323_p)
  );


  DROC
  ffc_325_3
  (
    .doutp(ffc_325_p),
    .doutn(ffc_325_n),
    .din(ffc_324_p)
  );


  DROC
  ffc_326_0
  (
    .doutp(ffc_326_p),
    .doutn(ffc_326_n),
    .din(G86_p)
  );


  DROC
  ffc_327_1
  (
    .doutp(ffc_327_p),
    .doutn(ffc_327_n),
    .din(ffc_326_p)
  );


  DROC
  ffc_328_2
  (
    .doutp(ffc_328_p),
    .doutn(ffc_328_n),
    .din(ffc_327_p)
  );


  DROC
  ffc_329_3
  (
    .doutp(ffc_329_p),
    .doutn(ffc_329_n),
    .din(ffc_328_p)
  );


  DROC
  ffc_330_0
  (
    .doutp(ffc_330_p),
    .doutn(ffc_330_n),
    .din(G87_p)
  );


  DROC
  ffc_331_1
  (
    .doutp(ffc_331_p),
    .doutn(ffc_331_n),
    .din(ffc_330_p)
  );


  DROC
  ffc_332_2
  (
    .doutp(ffc_332_p),
    .doutn(ffc_332_n),
    .din(ffc_331_p)
  );


  DROC
  ffc_333_3
  (
    .doutp(ffc_333_p),
    .doutn(ffc_333_n),
    .din(ffc_332_p)
  );


  DROC
  ffc_334_0
  (
    .doutp(ffc_334_p),
    .doutn(ffc_334_n),
    .din(G88_p)
  );


  DROC
  ffc_335_0
  (
    .doutp(ffc_335_p),
    .doutn(ffc_335_n),
    .din(G89_p)
  );


  DROC
  ffc_336_0
  (
    .doutp(ffc_336_p),
    .doutn(ffc_336_n),
    .din(G96_p)
  );


  DROC
  ffc_337_0
  (
    .doutp(ffc_337_p),
    .doutn(ffc_337_n),
    .din(G97_p)
  );


  DROC
  ffc_338_0
  (
    .doutp(ffc_338_p),
    .doutn(ffc_338_n),
    .din(G98_p)
  );


  DROC
  ffc_339_0
  (
    .doutp(ffc_339_p),
    .doutn(ffc_339_n),
    .din(G99_p)
  );


  DROC
  ffc_340_1
  (
    .doutp(ffc_340_p),
    .doutn(ffc_340_n),
    .din(ffc_339_p)
  );


  DROC
  ffc_341_2
  (
    .doutp(ffc_341_p),
    .doutn(ffc_341_n),
    .din(ffc_340_p)
  );


  DROC
  ffc_342_3
  (
    .doutp(ffc_342_p),
    .doutn(ffc_342_n),
    .din(ffc_341_p)
  );


  DROC
  ffc_343_0
  (
    .doutp(ffc_343_p),
    .doutn(ffc_343_n),
    .din(G100_p)
  );


  DROC
  ffc_344_0
  (
    .doutp(ffc_344_p),
    .doutn(ffc_344_n),
    .din(G101_p)
  );


  DROC
  ffc_345_0
  (
    .doutp(ffc_345_p),
    .doutn(ffc_345_n),
    .din(G102_p)
  );


  DROC
  ffc_346_0
  (
    .doutp(ffc_346_p),
    .doutn(ffc_346_n),
    .din(G103_p)
  );


  DROC
  ffc_347_0
  (
    .doutp(ffc_347_p),
    .doutn(ffc_347_n),
    .din(G104_p)
  );


  DROC
  ffc_348_0
  (
    .doutp(ffc_348_p),
    .doutn(ffc_348_n),
    .din(G111_p)
  );


  DROC
  ffc_349_1
  (
    .doutp(ffc_349_p),
    .doutn(ffc_349_n),
    .din(ffc_348_p)
  );


  DROC
  ffc_350_2
  (
    .doutp(ffc_350_p),
    .doutn(ffc_350_n),
    .din(ffc_349_p)
  );


  DROC
  ffc_351_0
  (
    .doutp(ffc_351_p),
    .doutn(ffc_351_n),
    .din(G112_p)
  );


  DROC
  ffc_352_1
  (
    .doutp(ffc_352_p),
    .doutn(ffc_352_n),
    .din(ffc_351_p)
  );


  DROC
  ffc_353_2
  (
    .doutp(ffc_353_p),
    .doutn(ffc_353_n),
    .din(ffc_352_p)
  );


  DROC
  ffc_354_0
  (
    .doutp(ffc_354_p),
    .doutn(ffc_354_n),
    .din(G113_p)
  );


  DROC
  ffc_355_1
  (
    .doutp(ffc_355_p),
    .doutn(ffc_355_n),
    .din(ffc_354_p)
  );


  DROC
  ffc_356_3
  (
    .doutp(ffc_356_p),
    .doutn(ffc_356_n),
    .din(ffc_640_p_spl_)
  );


  DROC
  ffc_357_0
  (
    .doutp(ffc_357_p),
    .doutn(ffc_357_n),
    .din(G114_p)
  );


  DROC
  ffc_358_1
  (
    .doutp(ffc_358_p),
    .doutn(ffc_358_n),
    .din(ffc_357_p)
  );


  DROC
  ffc_359_3
  (
    .doutp(ffc_359_p),
    .doutn(ffc_359_n),
    .din(ffc_657_p)
  );


  DROC
  ffc_360_0
  (
    .doutp(ffc_360_p),
    .doutn(ffc_360_n),
    .din(G115_p)
  );


  DROC
  ffc_361_0
  (
    .doutp(ffc_361_p),
    .doutn(ffc_361_n),
    .din(G116_p)
  );


  DROC
  ffc_362_0
  (
    .doutp(ffc_362_p),
    .doutn(ffc_362_n),
    .din(G121_p)
  );


  DROC
  ffc_363_0
  (
    .doutp(ffc_363_p),
    .doutn(ffc_363_n),
    .din(G122_p)
  );


  DROC
  ffc_364_0
  (
    .doutp(ffc_364_p),
    .doutn(ffc_364_n),
    .din(G125_p)
  );


  DROC
  ffc_365_3
  (
    .doutp(ffc_365_p),
    .doutn(ffc_365_n),
    .din(ffc_570_p)
  );


  DROC
  ffc_366_0
  (
    .doutp(ffc_366_p),
    .doutn(ffc_366_n),
    .din(G126_p)
  );


  DROC
  ffc_367_0
  (
    .doutp(ffc_367_p),
    .doutn(ffc_367_n),
    .din(G127_p)
  );


  DROC
  ffc_368_3
  (
    .doutp(ffc_368_p),
    .doutn(ffc_368_n),
    .din(ffc_558_p)
  );


  DROC
  ffc_369_3
  (
    .doutp(ffc_369_p),
    .doutn(ffc_369_n),
    .din(ffc_550_p)
  );


  DROC
  ffc_370_0
  (
    .doutp(ffc_370_p),
    .doutn(ffc_370_n),
    .din(G130_p)
  );


  DROC
  ffc_371_0
  (
    .doutp(ffc_371_p),
    .doutn(ffc_371_n),
    .din(G131_p)
  );


  DROC
  ffc_372_3
  (
    .doutp(ffc_372_p),
    .doutn(ffc_372_n),
    .din(ffc_572_p)
  );


  DROC
  ffc_373_0
  (
    .doutp(ffc_373_p),
    .doutn(ffc_373_n),
    .din(G132_p)
  );


  DROC
  ffc_374_1
  (
    .doutp(ffc_374_p),
    .doutn(ffc_374_n),
    .din(ffc_373_p)
  );


  DROC
  ffc_375_2
  (
    .doutp(ffc_375_p),
    .doutn(ffc_375_n),
    .din(ffc_374_p)
  );


  DROC
  ffc_376_0
  (
    .doutp(ffc_376_p),
    .doutn(ffc_376_n),
    .din(G133_p)
  );


  DROC
  ffc_377_1
  (
    .doutp(ffc_377_p),
    .doutn(ffc_377_n),
    .din(ffc_376_p)
  );


  DROC
  ffc_378_2
  (
    .doutp(ffc_378_p),
    .doutn(ffc_378_n),
    .din(ffc_377_p)
  );


  DROC
  ffc_379_0
  (
    .doutp(ffc_379_p),
    .doutn(ffc_379_n),
    .din(G134_p)
  );


  DROC
  ffc_380_1
  (
    .doutp(ffc_380_p),
    .doutn(ffc_380_n),
    .din(ffc_379_p)
  );


  DROC
  ffc_381_2
  (
    .doutp(ffc_381_p),
    .doutn(ffc_381_n),
    .din(ffc_380_p)
  );


  DROC
  ffc_382_3
  (
    .doutp(ffc_382_p),
    .doutn(ffc_382_n),
    .din(ffc_381_p)
  );


  DROC
  ffc_383_0
  (
    .doutp(ffc_383_p),
    .doutn(ffc_383_n),
    .din(G136_p)
  );


  DROC
  ffc_384_1
  (
    .doutp(ffc_384_p),
    .doutn(ffc_384_n),
    .din(ffc_383_p)
  );


  DROC
  ffc_385_2
  (
    .doutp(ffc_385_p),
    .doutn(ffc_385_n),
    .din(ffc_384_p)
  );


  DROC
  ffc_386_3
  (
    .doutp(ffc_386_p),
    .doutn(ffc_386_n),
    .din(ffc_385_p)
  );


  DROC
  ffc_387_0
  (
    .doutp(ffc_387_p),
    .doutn(ffc_387_n),
    .din(G137_p)
  );


  DROC
  ffc_388_0
  (
    .doutp(ffc_388_p),
    .doutn(ffc_388_n),
    .din(G138_p)
  );


  DROC
  ffc_389_0
  (
    .doutp(ffc_389_p),
    .doutn(ffc_389_n),
    .din(G141_p)
  );


  DROC
  ffc_390_1
  (
    .doutp(ffc_390_p),
    .doutn(ffc_390_n),
    .din(ffc_389_p)
  );


  DROC
  ffc_391_0
  (
    .doutp(ffc_391_p),
    .doutn(ffc_391_n),
    .din(G142_p)
  );


  DROC
  ffc_392_0
  (
    .doutp(ffc_392_p),
    .doutn(ffc_392_n),
    .din(G143_p)
  );


  DROC
  ffc_393_0
  (
    .doutp(ffc_393_p),
    .doutn(ffc_393_n),
    .din(G146_p)
  );


  DROC
  ffc_394_0
  (
    .doutp(ffc_394_p),
    .doutn(ffc_394_n),
    .din(G147_p)
  );


  DROC
  ffc_395_0
  (
    .doutp(ffc_395_p),
    .doutn(ffc_395_n),
    .din(G148_p)
  );


  DROC
  ffc_396_0
  (
    .doutp(ffc_396_p),
    .doutn(ffc_396_n),
    .din(G149_p)
  );


  DROC
  ffc_397_0
  (
    .doutp(ffc_397_p),
    .doutn(ffc_397_n),
    .din(G150_p)
  );


  DROC
  ffc_398_0
  (
    .doutp(ffc_398_p),
    .doutn(ffc_398_n),
    .din(G151_p)
  );


  DROC
  ffc_399_1
  (
    .doutp(ffc_399_p),
    .doutn(ffc_399_n),
    .din(ffc_398_p)
  );


  DROC
  ffc_400_2
  (
    .doutp(ffc_400_p),
    .doutn(ffc_400_n),
    .din(ffc_399_p)
  );


  DROC
  ffc_401_3
  (
    .doutp(ffc_401_p),
    .doutn(ffc_401_n),
    .din(ffc_400_p)
  );


  DROC
  ffc_402_0
  (
    .doutp(ffc_402_p),
    .doutn(ffc_402_n),
    .din(G152_p)
  );


  DROC
  ffc_403_1
  (
    .doutp(ffc_403_p),
    .doutn(ffc_403_n),
    .din(ffc_402_p)
  );


  DROC
  ffc_404_2
  (
    .doutp(ffc_404_p),
    .doutn(ffc_404_n),
    .din(ffc_403_p)
  );


  DROC
  ffc_405_3
  (
    .doutp(ffc_405_p),
    .doutn(ffc_405_n),
    .din(ffc_404_p)
  );


  DROC
  ffc_406_0
  (
    .doutp(ffc_406_p),
    .doutn(ffc_406_n),
    .din(G153_p)
  );


  DROC
  ffc_407_1
  (
    .doutp(ffc_407_p),
    .doutn(ffc_407_n),
    .din(ffc_406_p)
  );


  DROC
  ffc_408_2
  (
    .doutp(ffc_408_p),
    .doutn(ffc_408_n),
    .din(ffc_407_p)
  );


  DROC
  ffc_409_3
  (
    .doutp(ffc_409_p),
    .doutn(ffc_409_n),
    .din(ffc_408_p)
  );


  DROC
  ffc_410_0
  (
    .doutp(ffc_410_p),
    .doutn(ffc_410_n),
    .din(G154_p)
  );


  DROC
  ffc_411_1
  (
    .doutp(ffc_411_p),
    .doutn(ffc_411_n),
    .din(ffc_410_p)
  );


  DROC
  ffc_412_2
  (
    .doutp(ffc_412_p),
    .doutn(ffc_412_n),
    .din(ffc_411_p)
  );


  DROC
  ffc_413_3
  (
    .doutp(ffc_413_p),
    .doutn(ffc_413_n),
    .din(ffc_412_p)
  );


  DROC
  ffc_414_0
  (
    .doutp(ffc_414_p),
    .doutn(ffc_414_n),
    .din(G155_p)
  );


  DROC
  ffc_415_1
  (
    .doutp(ffc_415_p),
    .doutn(ffc_415_n),
    .din(ffc_414_p)
  );


  DROC
  ffc_416_2
  (
    .doutp(ffc_416_p),
    .doutn(ffc_416_n),
    .din(ffc_415_p)
  );


  DROC
  ffc_417_3
  (
    .doutp(ffc_417_p),
    .doutn(ffc_417_n),
    .din(ffc_416_p)
  );


  DROC
  ffc_418_0
  (
    .doutp(ffc_418_p),
    .doutn(ffc_418_n),
    .din(G156_p)
  );


  DROC
  ffc_419_1
  (
    .doutp(ffc_419_p),
    .doutn(ffc_419_n),
    .din(ffc_418_p)
  );


  DROC
  ffc_420_2
  (
    .doutp(ffc_420_p),
    .doutn(ffc_420_n),
    .din(ffc_419_p)
  );


  DROC
  ffc_421_3
  (
    .doutp(ffc_421_p),
    .doutn(ffc_421_n),
    .din(ffc_420_p)
  );


  DROC
  ffc_422_0
  (
    .doutp(ffc_422_p),
    .doutn(ffc_422_n),
    .din(G157_p)
  );


  DROC
  ffc_423_1
  (
    .doutp(ffc_423_p),
    .doutn(ffc_423_n),
    .din(ffc_422_p)
  );


  DROC
  ffc_424_2
  (
    .doutp(ffc_424_p),
    .doutn(ffc_424_n),
    .din(ffc_423_p)
  );


  DROC
  ffc_425_0
  (
    .doutp(ffc_425_p),
    .doutn(ffc_425_n),
    .din(G158_p)
  );


  DROC
  ffc_426_1
  (
    .doutp(ffc_426_p),
    .doutn(ffc_426_n),
    .din(ffc_425_p)
  );


  DROC
  ffc_427_2
  (
    .doutp(ffc_427_p),
    .doutn(ffc_427_n),
    .din(ffc_426_p)
  );


  DROC
  ffc_428_3
  (
    .doutp(ffc_428_p),
    .doutn(ffc_428_n),
    .din(ffc_427_p)
  );


  DROC
  ffc_429_0
  (
    .doutp(ffc_429_p),
    .doutn(ffc_429_n),
    .din(G159_p)
  );


  DROC
  ffc_430_1
  (
    .doutp(ffc_430_p),
    .doutn(ffc_430_n),
    .din(ffc_429_p)
  );


  DROC
  ffc_431_2
  (
    .doutp(ffc_431_p),
    .doutn(ffc_431_n),
    .din(ffc_430_p)
  );


  DROC
  ffc_432_3
  (
    .doutp(ffc_432_p),
    .doutn(ffc_432_n),
    .din(ffc_431_p)
  );


  DROC
  ffc_433_0
  (
    .doutp(ffc_433_p),
    .doutn(ffc_433_n),
    .din(G160_p)
  );


  DROC
  ffc_434_1
  (
    .doutp(ffc_434_p),
    .doutn(ffc_434_n),
    .din(ffc_433_p)
  );


  DROC
  ffc_435_2
  (
    .doutp(ffc_435_p),
    .doutn(ffc_435_n),
    .din(ffc_434_p)
  );


  DROC
  ffc_436_3
  (
    .doutp(ffc_436_p),
    .doutn(ffc_436_n),
    .din(ffc_435_p)
  );


  DROC
  ffc_437_0
  (
    .doutp(ffc_437_p),
    .doutn(ffc_437_n),
    .din(G161_p)
  );


  DROC
  ffc_438_1
  (
    .doutp(ffc_438_p),
    .doutn(ffc_438_n),
    .din(ffc_437_p)
  );


  DROC
  ffc_439_2
  (
    .doutp(ffc_439_p),
    .doutn(ffc_439_n),
    .din(ffc_438_p)
  );


  DROC
  ffc_440_3
  (
    .doutp(ffc_440_p),
    .doutn(ffc_440_n),
    .din(ffc_439_p)
  );


  DROC
  ffc_441_0
  (
    .doutp(ffc_441_p),
    .doutn(ffc_441_n),
    .din(G162_p)
  );


  DROC
  ffc_442_1
  (
    .doutp(ffc_442_p),
    .doutn(ffc_442_n),
    .din(ffc_441_p)
  );


  DROC
  ffc_443_0
  (
    .doutp(ffc_443_p),
    .doutn(ffc_443_n),
    .din(G163_p)
  );


  DROC
  ffc_444_1
  (
    .doutp(ffc_444_p),
    .doutn(ffc_444_n),
    .din(ffc_443_p)
  );


  DROC
  ffc_445_2
  (
    .doutp(ffc_445_p),
    .doutn(ffc_445_n),
    .din(ffc_444_p)
  );


  DROC
  ffc_446_3
  (
    .doutp(ffc_446_p),
    .doutn(ffc_446_n),
    .din(ffc_445_p)
  );


  DROC
  ffc_447_0
  (
    .doutp(ffc_447_p),
    .doutn(ffc_447_n),
    .din(G164_p)
  );


  DROC
  ffc_448_1
  (
    .doutp(ffc_448_p),
    .doutn(ffc_448_n),
    .din(ffc_447_p)
  );


  DROC
  ffc_449_2
  (
    .doutp(ffc_449_p),
    .doutn(ffc_449_n),
    .din(ffc_448_p)
  );


  DROC
  ffc_450_3
  (
    .doutp(ffc_450_p),
    .doutn(ffc_450_n),
    .din(ffc_449_p)
  );


  DROC
  ffc_451_0
  (
    .doutp(ffc_451_p),
    .doutn(ffc_451_n),
    .din(G165_p)
  );


  DROC
  ffc_452_1
  (
    .doutp(ffc_452_p),
    .doutn(ffc_452_n),
    .din(ffc_451_p)
  );


  DROC
  ffc_453_2
  (
    .doutp(ffc_453_p),
    .doutn(ffc_453_n),
    .din(ffc_452_p)
  );


  DROC
  ffc_454_3
  (
    .doutp(ffc_454_p),
    .doutn(ffc_454_n),
    .din(ffc_453_p)
  );


  DROC
  ffc_455_0
  (
    .doutp(ffc_455_p),
    .doutn(ffc_455_n),
    .din(G166_p)
  );


  DROC
  ffc_456_1
  (
    .doutp(ffc_456_p),
    .doutn(ffc_456_n),
    .din(ffc_455_p)
  );


  DROC
  ffc_457_2
  (
    .doutp(ffc_457_p),
    .doutn(ffc_457_n),
    .din(ffc_456_p)
  );


  DROC
  ffc_458_0
  (
    .doutp(ffc_458_p),
    .doutn(ffc_458_n),
    .din(G167_p)
  );


  DROC
  ffc_459_1
  (
    .doutp(ffc_459_p),
    .doutn(ffc_459_n),
    .din(ffc_458_p)
  );


  DROC
  ffc_460_2
  (
    .doutp(ffc_460_p),
    .doutn(ffc_460_n),
    .din(ffc_459_p)
  );


  DROC
  ffc_461_0
  (
    .doutp(ffc_461_p),
    .doutn(ffc_461_n),
    .din(G168_p)
  );


  DROC
  ffc_462_1
  (
    .doutp(ffc_462_p),
    .doutn(ffc_462_n),
    .din(ffc_461_p)
  );


  DROC
  ffc_463_2
  (
    .doutp(ffc_463_p),
    .doutn(ffc_463_n),
    .din(ffc_462_p)
  );


  DROC
  ffc_464_0
  (
    .doutp(ffc_464_p),
    .doutn(ffc_464_n),
    .din(G169_p)
  );


  DROC
  ffc_465_1
  (
    .doutp(ffc_465_p),
    .doutn(ffc_465_n),
    .din(ffc_464_p)
  );


  DROC
  ffc_466_2
  (
    .doutp(ffc_466_p),
    .doutn(ffc_466_n),
    .din(ffc_465_p)
  );


  DROC
  ffc_467_0
  (
    .doutp(ffc_467_p),
    .doutn(ffc_467_n),
    .din(G170_p)
  );


  DROC
  ffc_468_1
  (
    .doutp(ffc_468_p),
    .doutn(ffc_468_n),
    .din(ffc_467_p)
  );


  DROC
  ffc_469_2
  (
    .doutp(ffc_469_p),
    .doutn(ffc_469_n),
    .din(ffc_468_p)
  );


  DROC
  ffc_470_3
  (
    .doutp(ffc_470_p),
    .doutn(ffc_470_n),
    .din(ffc_469_p)
  );


  DROC
  ffc_471_0
  (
    .doutp(ffc_471_p),
    .doutn(ffc_471_n),
    .din(G171_p)
  );


  DROC
  ffc_472_1
  (
    .doutp(ffc_472_p),
    .doutn(ffc_472_n),
    .din(ffc_471_p)
  );


  DROC
  ffc_473_2
  (
    .doutp(ffc_473_p),
    .doutn(ffc_473_n),
    .din(ffc_472_p)
  );


  DROC
  ffc_474_3
  (
    .doutp(ffc_474_p),
    .doutn(ffc_474_n),
    .din(ffc_473_p)
  );


  DROC
  ffc_475_0
  (
    .doutp(ffc_475_p),
    .doutn(ffc_475_n),
    .din(G172_p)
  );


  DROC
  ffc_476_1
  (
    .doutp(ffc_476_p),
    .doutn(ffc_476_n),
    .din(ffc_475_p)
  );


  DROC
  ffc_477_2
  (
    .doutp(ffc_477_p),
    .doutn(ffc_477_n),
    .din(ffc_476_p)
  );


  DROC
  ffc_478_3
  (
    .doutp(ffc_478_p),
    .doutn(ffc_478_n),
    .din(ffc_477_p)
  );


  DROC
  ffc_479_0
  (
    .doutp(ffc_479_p),
    .doutn(ffc_479_n),
    .din(G173_p)
  );


  DROC
  ffc_480_1
  (
    .doutp(ffc_480_p),
    .doutn(ffc_480_n),
    .din(ffc_479_p)
  );


  DROC
  ffc_481_2
  (
    .doutp(ffc_481_p),
    .doutn(ffc_481_n),
    .din(ffc_480_p)
  );


  DROC
  ffc_482_3
  (
    .doutp(ffc_482_p),
    .doutn(ffc_482_n),
    .din(ffc_481_p)
  );


  DROC
  ffc_483_0
  (
    .doutp(ffc_483_p),
    .doutn(ffc_483_n),
    .din(G174_p)
  );


  DROC
  ffc_484_1
  (
    .doutp(ffc_484_p),
    .doutn(ffc_484_n),
    .din(ffc_483_p)
  );


  DROC
  ffc_485_2
  (
    .doutp(ffc_485_p),
    .doutn(ffc_485_n),
    .din(ffc_484_p)
  );


  DROC
  ffc_486_3
  (
    .doutp(ffc_486_p),
    .doutn(ffc_486_n),
    .din(ffc_485_p)
  );


  DROC
  ffc_487_0
  (
    .doutp(ffc_487_p),
    .doutn(ffc_487_n),
    .din(G175_p)
  );


  DROC
  ffc_488_1
  (
    .doutp(ffc_488_p),
    .doutn(ffc_488_n),
    .din(ffc_487_p)
  );


  DROC
  ffc_489_2
  (
    .doutp(ffc_489_p),
    .doutn(ffc_489_n),
    .din(ffc_488_p)
  );


  DROC
  ffc_490_3
  (
    .doutp(ffc_490_p),
    .doutn(ffc_490_n),
    .din(ffc_489_p)
  );


  DROC
  ffc_491_0
  (
    .doutp(ffc_491_p),
    .doutn(ffc_491_n),
    .din(G176_p)
  );


  DROC
  ffc_492_1
  (
    .doutp(ffc_492_p),
    .doutn(ffc_492_n),
    .din(ffc_491_p)
  );


  DROC
  ffc_493_2
  (
    .doutp(ffc_493_p),
    .doutn(ffc_493_n),
    .din(ffc_492_p)
  );


  DROC
  ffc_494_3
  (
    .doutp(ffc_494_p),
    .doutn(ffc_494_n),
    .din(ffc_493_p_spl_)
  );


  DROC
  ffc_495_0
  (
    .doutp(ffc_495_p),
    .doutn(ffc_495_n),
    .din(G177_p)
  );


  DROC
  ffc_496_1
  (
    .doutp(ffc_496_p),
    .doutn(ffc_496_n),
    .din(ffc_495_p)
  );


  DROC
  ffc_497_2
  (
    .doutp(ffc_497_p),
    .doutn(ffc_497_n),
    .din(ffc_496_p)
  );


  DROC
  ffc_498_3
  (
    .doutp(ffc_498_p),
    .doutn(ffc_498_n),
    .din(ffc_497_p_spl_11)
  );


  DROC
  ffc_499_0
  (
    .doutp(ffc_499_p),
    .doutn(ffc_499_n),
    .din(G178_p)
  );


  DROC
  ffc_500_1
  (
    .doutp(ffc_500_p),
    .doutn(ffc_500_n),
    .din(ffc_499_p)
  );


  DROC
  ffc_501_2
  (
    .doutp(ffc_501_p),
    .doutn(ffc_501_n),
    .din(ffc_500_p)
  );


  DROC
  ffc_502_3
  (
    .doutp(ffc_502_p),
    .doutn(ffc_502_n),
    .din(ffc_501_p)
  );


  DROC
  ffc_503_3
  (
    .doutp(ffc_503_p),
    .doutn(ffc_503_n),
    .din(ffc_546_p)
  );


  DROC
  ffc_504_3
  (
    .doutp(ffc_504_p),
    .doutn(ffc_504_n),
    .din(ffc_548_p)
  );


  DROC
  ffc_505_3
  (
    .doutp(ffc_505_p),
    .doutn(ffc_505_n),
    .din(ffc_554_p)
  );


  DROC
  ffc_506_3
  (
    .doutp(ffc_506_p),
    .doutn(ffc_506_n),
    .din(ffc_563_p)
  );


  DROC
  ffc_507_3
  (
    .doutp(ffc_507_p),
    .doutn(ffc_507_n),
    .din(ffc_564_p)
  );


  DROC
  ffc_508_3
  (
    .doutp(ffc_508_p),
    .doutn(ffc_508_n),
    .din(ffc_568_p)
  );


  DROC
  ffc_509_3
  (
    .doutp(ffc_509_p),
    .doutn(ffc_509_n),
    .din(ffc_575_p)
  );


  DROC
  ffc_510_3
  (
    .doutp(ffc_510_p),
    .doutn(ffc_510_n),
    .din(ffc_579_p)
  );


  DROC
  ffc_511_3
  (
    .doutp(ffc_511_p),
    .doutn(ffc_511_n),
    .din(ffc_585_p)
  );


  DROC
  ffc_512_3
  (
    .doutp(ffc_512_p),
    .doutn(ffc_512_n),
    .din(ffc_588_p)
  );


  DROC
  ffc_513_3
  (
    .doutp(ffc_513_p),
    .doutn(ffc_513_n),
    .din(ffc_602_p)
  );


  DROC
  ffc_514_3
  (
    .doutp(ffc_514_p),
    .doutn(ffc_514_n),
    .din(ffc_606_p)
  );


  DROC
  ffc_515_3
  (
    .doutp(ffc_515_p),
    .doutn(ffc_515_n),
    .din(ffc_608_p_spl_)
  );


  DROC
  ffc_516_3
  (
    .doutp(ffc_516_p),
    .doutn(ffc_516_n),
    .din(ffc_610_p_spl_)
  );


  DROC
  ffc_517_3
  (
    .doutp(ffc_517_p),
    .doutn(ffc_517_n),
    .din(ffc_614_p_spl_)
  );


  DROC
  ffc_518_3
  (
    .doutp(ffc_518_p),
    .doutn(ffc_518_n),
    .din(ffc_615_p_spl_)
  );


  DROC
  ffc_519_3
  (
    .doutp(ffc_519_p),
    .doutn(ffc_519_n),
    .din(ffc_617_p)
  );


  DROC
  ffc_520_3
  (
    .doutp(ffc_520_p),
    .doutn(ffc_520_n),
    .din(ffc_626_p)
  );


  DROC
  ffc_521_3
  (
    .doutp(ffc_521_p),
    .doutn(ffc_521_n),
    .din(ffc_630_p)
  );


  DROC
  ffc_522_3
  (
    .doutp(ffc_522_p),
    .doutn(ffc_522_n),
    .din(ffc_647_p)
  );


  DROC
  ffc_523_3
  (
    .doutp(ffc_523_p),
    .doutn(ffc_523_n),
    .din(ffc_670_p)
  );


  DROC
  ffc_524_3
  (
    .doutp(ffc_524_p),
    .doutn(ffc_524_n),
    .din(ffc_762_p)
  );


  DROC
  ffc_525_3
  (
    .doutp(ffc_525_p),
    .doutn(ffc_525_n),
    .din(ffc_760_p)
  );


  DROC
  ffc_526_2
  (
    .doutp(ffc_526_p),
    .doutn(ffc_526_n),
    .din(ffc_620_p_spl_)
  );


  DROC
  ffc_527_2
  (
    .doutp(ffc_527_p),
    .doutn(ffc_527_n),
    .din(ffc_621_p_spl_)
  );


  DROC
  ffc_528_2
  (
    .doutp(ffc_528_p),
    .doutn(ffc_528_n),
    .din(ffc_622_p_spl_)
  );


  DROC
  ffc_529_2
  (
    .doutp(ffc_529_p),
    .doutn(ffc_529_n),
    .din(ffc_623_p_spl_)
  );


  DROC
  ffc_530_3
  (
    .doutp(ffc_530_p),
    .doutn(ffc_530_n),
    .din(ffc_771_p_spl_1)
  );


  DROC
  ffc_531_3
  (
    .doutp(ffc_531_p),
    .doutn(ffc_531_n),
    .din(ffc_772_p_spl_1)
  );


  DROC
  ffc_532_3
  (
    .doutp(ffc_532_p),
    .doutn(ffc_532_n),
    .din(ffc_783_p_spl_)
  );


  DROC
  ffc_533_3
  (
    .doutp(ffc_533_p),
    .doutn(ffc_533_n),
    .din(ffc_790_p_spl_)
  );


  DROC
  ffc_534_3
  (
    .doutp(ffc_534_p),
    .doutn(ffc_534_n),
    .din(ffc_802_p_spl_)
  );


  DROC
  ffc_535_3
  (
    .doutp(ffc_535_p),
    .doutn(ffc_535_n),
    .din(ffc_800_p_spl_)
  );


  DROC
  ffc_536_2
  (
    .doutp(ffc_536_p),
    .doutn(ffc_536_n),
    .din(ffc_627_p_spl_)
  );


  DROC
  ffc_537_2
  (
    .doutp(ffc_537_p),
    .doutn(ffc_537_n),
    .din(ffc_628_p_spl_)
  );


  DROC
  ffc_538_2
  (
    .doutp(ffc_538_p),
    .doutn(ffc_538_n),
    .din(ffc_629_p_spl_)
  );


  DROC
  ffc_539_2
  (
    .doutp(ffc_539_p),
    .doutn(ffc_539_n),
    .din(ffc_631_p_spl_)
  );


  DROC
  ffc_540_2
  (
    .doutp(ffc_540_p),
    .doutn(ffc_540_n),
    .din(ffc_632_p_spl_)
  );


  DROC
  ffc_541_2
  (
    .doutp(ffc_541_p),
    .doutn(ffc_541_n),
    .din(ffc_633_p_spl_)
  );


  DROC
  ffc_542_2
  (
    .doutp(ffc_542_p),
    .doutn(ffc_542_n),
    .din(ffc_634_p_spl_)
  );


  DROC
  ffc_543_2
  (
    .doutp(ffc_543_p),
    .doutn(ffc_543_n),
    .din(ffc_635_p_spl_)
  );


  DROC
  ffc_544_2
  (
    .doutp(ffc_544_p),
    .doutn(ffc_544_n),
    .din(ffc_636_p_spl_)
  );


  DROC
  ffc_545_3
  (
    .doutp(ffc_545_p),
    .doutn(ffc_545_n),
    .din(g1690_n_spl_)
  );


  DROC
  ffc_546_2
  (
    .doutp(ffc_546_p),
    .doutn(ffc_546_n),
    .din(ffc_637_p)
  );


  DROC
  ffc_547_2
  (
    .doutp(ffc_547_p),
    .doutn(ffc_547_n),
    .din(ffc_638_p)
  );


  DROC
  ffc_548_2
  (
    .doutp(ffc_548_p),
    .doutn(ffc_548_n),
    .din(ffc_639_p)
  );


  DROC
  ffc_549_2
  (
    .doutp(ffc_549_p),
    .doutn(ffc_549_n),
    .din(ffc_648_p_spl_)
  );


  DROC
  ffc_550_2
  (
    .doutp(ffc_550_p),
    .doutn(ffc_550_n),
    .din(ffc_649_p)
  );


  DROC
  ffc_551_2
  (
    .doutp(ffc_551_p),
    .doutn(ffc_551_n),
    .din(ffc_650_p_spl_)
  );


  DROC
  ffc_552_2
  (
    .doutp(ffc_552_p),
    .doutn(ffc_552_n),
    .din(ffc_653_p)
  );


  DROC
  ffc_553_2
  (
    .doutp(ffc_553_p),
    .doutn(ffc_553_n),
    .din(ffc_654_p)
  );


  DROC
  ffc_554_2
  (
    .doutp(ffc_554_p),
    .doutn(ffc_554_n),
    .din(ffc_652_p)
  );


  DROC
  ffc_555_2
  (
    .doutp(ffc_555_p),
    .doutn(ffc_555_n),
    .din(ffc_656_p)
  );


  DROC
  ffc_556_2
  (
    .doutp(ffc_556_p),
    .doutn(ffc_556_n),
    .din(ffc_660_p_spl_1)
  );


  DROC
  ffc_557_2
  (
    .doutp(ffc_557_p),
    .doutn(ffc_557_n),
    .din(ffc_661_p_spl_)
  );


  DROC
  ffc_558_2
  (
    .doutp(ffc_558_p),
    .doutn(ffc_558_n),
    .din(ffc_662_p)
  );


  DROC
  ffc_559_2
  (
    .doutp(ffc_559_p),
    .doutn(ffc_559_n),
    .din(ffc_663_p_spl_)
  );


  DROC
  ffc_560_2
  (
    .doutp(ffc_560_p),
    .doutn(ffc_560_n),
    .din(ffc_664_p_spl_)
  );


  DROC
  ffc_561_3
  (
    .doutp(ffc_561_p),
    .doutn(ffc_561_n),
    .din(g1692_p_spl_)
  );


  DROC
  ffc_562_2
  (
    .doutp(ffc_562_p),
    .doutn(ffc_562_n),
    .din(ffc_671_p_spl_)
  );


  DROC
  ffc_563_2
  (
    .doutp(ffc_563_p),
    .doutn(ffc_563_n),
    .din(ffc_666_p)
  );


  DROC
  ffc_564_2
  (
    .doutp(ffc_564_p),
    .doutn(ffc_564_n),
    .din(ffc_667_p)
  );


  DROC
  ffc_565_2
  (
    .doutp(ffc_565_p),
    .doutn(ffc_565_n),
    .din(ffc_669_p)
  );


  DROC
  ffc_566_2
  (
    .doutp(ffc_566_p),
    .doutn(ffc_566_n),
    .din(ffc_672_p_spl_)
  );


  DROC
  ffc_567_2
  (
    .doutp(ffc_567_p),
    .doutn(ffc_567_n),
    .din(ffc_673_p_spl_1)
  );


  DROC
  ffc_568_2
  (
    .doutp(ffc_568_p),
    .doutn(ffc_568_n),
    .din(ffc_674_p_spl_)
  );


  DROC
  ffc_569_2
  (
    .doutp(ffc_569_p),
    .doutn(ffc_569_n),
    .din(ffc_675_p_spl_)
  );


  DROC
  ffc_570_2
  (
    .doutp(ffc_570_p),
    .doutn(ffc_570_n),
    .din(ffc_676_p)
  );


  DROC
  ffc_571_2
  (
    .doutp(ffc_571_p),
    .doutn(ffc_571_n),
    .din(ffc_677_p_spl_)
  );


  DROC
  ffc_572_2
  (
    .doutp(ffc_572_p),
    .doutn(ffc_572_n),
    .din(ffc_678_p)
  );


  DROC
  ffc_573_2
  (
    .doutp(ffc_573_p),
    .doutn(ffc_573_n),
    .din(ffc_679_p_spl_)
  );


  DROC
  ffc_574_2
  (
    .doutp(ffc_574_p),
    .doutn(ffc_574_n),
    .din(ffc_681_p)
  );


  DROC
  ffc_575_2
  (
    .doutp(ffc_575_p),
    .doutn(ffc_575_n),
    .din(ffc_682_p)
  );


  DROC
  ffc_576_2
  (
    .doutp(ffc_576_p),
    .doutn(ffc_576_n),
    .din(ffc_683_p_spl_)
  );


  DROC
  ffc_577_2
  (
    .doutp(ffc_577_p),
    .doutn(ffc_577_n),
    .din(ffc_680_p)
  );


  DROC
  ffc_578_2
  (
    .doutp(ffc_578_p),
    .doutn(ffc_578_n),
    .din(ffc_684_p)
  );


  DROC
  ffc_579_2
  (
    .doutp(ffc_579_p),
    .doutn(ffc_579_n),
    .din(ffc_685_p)
  );


  DROC
  ffc_580_2
  (
    .doutp(ffc_580_p),
    .doutn(ffc_580_n),
    .din(ffc_763_p_spl_)
  );


  DROC
  ffc_581_2
  (
    .doutp(ffc_581_p),
    .doutn(ffc_581_n),
    .din(ffc_764_p_spl_)
  );


  DROC
  ffc_582_2
  (
    .doutp(ffc_582_p),
    .doutn(ffc_582_n),
    .din(ffc_765_p_spl_)
  );


  DROC
  ffc_583_2
  (
    .doutp(ffc_583_p),
    .doutn(ffc_583_n),
    .din(ffc_724_p)
  );


  DROC
  ffc_584_2
  (
    .doutp(ffc_584_p),
    .doutn(ffc_584_n),
    .din(ffc_756_p_spl_1)
  );


  DROC
  ffc_585_2
  (
    .doutp(ffc_585_p),
    .doutn(ffc_585_n),
    .din(ffc_766_p)
  );


  DROC
  ffc_586_2
  (
    .doutp(ffc_586_p),
    .doutn(ffc_586_n),
    .din(ffc_767_p)
  );


  DROC
  ffc_587_2
  (
    .doutp(ffc_587_p),
    .doutn(ffc_587_n),
    .din(ffc_769_p_spl_1)
  );


  DROC
  ffc_588_2
  (
    .doutp(ffc_588_p),
    .doutn(ffc_588_n),
    .din(ffc_770_p_spl_)
  );


  DROC
  ffc_589_2
  (
    .doutp(ffc_589_p),
    .doutn(ffc_589_n),
    .din(ffc_780_p_spl_)
  );


  DROC
  ffc_590_2
  (
    .doutp(ffc_590_p),
    .doutn(ffc_590_n),
    .din(ffc_781_p_spl_1)
  );


  DROC
  ffc_591_2
  (
    .doutp(ffc_591_p),
    .doutn(ffc_591_n),
    .din(ffc_775_p_spl_)
  );


  DROC
  ffc_592_2
  (
    .doutp(ffc_592_p),
    .doutn(ffc_592_n),
    .din(ffc_778_p_spl_)
  );


  DROC
  ffc_593_2
  (
    .doutp(ffc_593_p),
    .doutn(ffc_593_n),
    .din(ffc_779_p_spl_)
  );


  DROC
  ffc_594_2
  (
    .doutp(ffc_594_p),
    .doutn(ffc_594_n),
    .din(ffc_812_p_spl_)
  );


  DROC
  ffc_595_2
  (
    .doutp(ffc_595_p),
    .doutn(ffc_595_n),
    .din(ffc_794_p)
  );


  DROC
  ffc_596_2
  (
    .doutp(ffc_596_p),
    .doutn(ffc_596_n),
    .din(ffc_795_p_spl_1)
  );


  DROC
  ffc_597_2
  (
    .doutp(ffc_597_p),
    .doutn(ffc_597_n),
    .din(ffc_799_p)
  );


  DROC
  ffc_598_2
  (
    .doutp(ffc_598_p),
    .doutn(ffc_598_n),
    .din(ffc_829_p_spl_1)
  );


  DROC
  ffc_599_3
  (
    .doutp(ffc_599_n),
    .doutn(ffc_599_p),
    .din(g1693_n_spl_)
  );


  DROC
  ffc_600_3
  (
    .doutp(ffc_600_p),
    .doutn(ffc_600_n),
    .din(g1696_p_spl_)
  );


  DROC
  ffc_601_2
  (
    .doutp(ffc_601_p),
    .doutn(ffc_601_n),
    .din(ffc_825_p_spl_1)
  );


  DROC
  ffc_602_2
  (
    .doutp(ffc_602_p),
    .doutn(ffc_602_n),
    .din(ffc_840_p_spl_)
  );


  DROC
  ffc_603_2
  (
    .doutp(ffc_603_p),
    .doutn(ffc_603_n),
    .din(ffc_844_p_spl_1)
  );


  DROC
  ffc_604_2
  (
    .doutp(ffc_604_p),
    .doutn(ffc_604_n),
    .din(ffc_843_p_spl_)
  );


  DROC
  ffc_605_2
  (
    .doutp(ffc_605_p),
    .doutn(ffc_605_n),
    .din(ffc_845_p_spl_)
  );


  DROC
  ffc_606_2
  (
    .doutp(ffc_606_p),
    .doutn(ffc_606_n),
    .din(ffc_842_p_spl_)
  );


  DROC
  ffc_607_2
  (
    .doutp(ffc_607_p),
    .doutn(ffc_607_n),
    .din(ffc_816_p_spl_1)
  );


  DROC
  ffc_608_2
  (
    .doutp(ffc_608_p),
    .doutn(ffc_608_n),
    .din(g1697_n_spl_)
  );


  DROC
  ffc_609_2
  (
    .doutp(ffc_609_p),
    .doutn(ffc_609_n),
    .din(g1698_n_spl_1)
  );


  DROC
  ffc_610_2
  (
    .doutp(ffc_610_p),
    .doutn(ffc_610_n),
    .din(g1699_n_spl_1)
  );


  DROC
  ffc_611_2
  (
    .doutp(ffc_611_p),
    .doutn(ffc_611_n),
    .din(g1700_n_spl_)
  );


  DROC
  ffc_612_2
  (
    .doutp(ffc_612_p),
    .doutn(ffc_612_n),
    .din(g1701_n_spl_)
  );


  DROC
  ffc_613_2
  (
    .doutp(ffc_613_p),
    .doutn(ffc_613_n),
    .din(g1702_n_spl_)
  );


  DROC
  ffc_614_2
  (
    .doutp(ffc_614_p),
    .doutn(ffc_614_n),
    .din(g1703_p_spl_)
  );


  DROC
  ffc_615_2
  (
    .doutp(ffc_615_p),
    .doutn(ffc_615_n),
    .din(g1704_p_spl_)
  );


  DROC
  ffc_616_2
  (
    .doutp(ffc_616_p),
    .doutn(ffc_616_n),
    .din(ffc_390_p_spl_1)
  );


  DROC
  ffc_617_2
  (
    .doutp(ffc_617_p),
    .doutn(ffc_617_n),
    .din(g1705_p_spl_)
  );


  DROC
  ffc_618_3
  (
    .doutp(ffc_618_p),
    .doutn(ffc_618_n),
    .din(g1708_n_spl_)
  );


  DROC
  ffc_619_2
  (
    .doutp(ffc_619_p),
    .doutn(ffc_619_n),
    .din(g1711_n_spl_)
  );


  DROC
  ffc_620_1
  (
    .doutp(ffc_620_p),
    .doutn(ffc_620_n),
    .din(ffc_836_p)
  );


  DROC
  ffc_621_1
  (
    .doutp(ffc_621_p),
    .doutn(ffc_621_n),
    .din(ffc_837_p)
  );


  DROC
  ffc_622_1
  (
    .doutp(ffc_622_p),
    .doutn(ffc_622_n),
    .din(ffc_838_p)
  );


  DROC
  ffc_623_1
  (
    .doutp(ffc_623_p),
    .doutn(ffc_623_n),
    .din(ffc_839_p_spl_11)
  );


  DROC
  ffc_624_2
  (
    .doutp(ffc_624_p),
    .doutn(ffc_624_n),
    .din(g1712_p_spl_)
  );


  DROC
  ffc_625_2
  (
    .doutp(ffc_625_p),
    .doutn(ffc_625_n),
    .din(g1714_n_spl_)
  );


  DROC
  ffc_626_2
  (
    .doutp(ffc_626_p),
    .doutn(ffc_626_n),
    .din(g1716_n_spl_)
  );


  DROC
  ffc_627_1
  (
    .doutp(ffc_627_p),
    .doutn(ffc_627_n),
    .din(ffc_859_p_spl_)
  );


  DROC
  ffc_628_1
  (
    .doutp(ffc_628_p),
    .doutn(ffc_628_n),
    .din(ffc_861_p_spl_)
  );


  DROC
  ffc_629_1
  (
    .doutp(ffc_629_p),
    .doutn(ffc_629_n),
    .din(ffc_863_p_spl_11)
  );


  DROC
  ffc_630_2
  (
    .doutp(ffc_630_p),
    .doutn(ffc_630_n),
    .din(g1719_p_spl_)
  );


  DROC
  ffc_631_1
  (
    .doutp(ffc_631_p),
    .doutn(ffc_631_n),
    .din(ffc_850_p_spl_)
  );


  DROC
  ffc_632_1
  (
    .doutp(ffc_632_p),
    .doutn(ffc_632_n),
    .din(ffc_852_p_spl_)
  );


  DROC
  ffc_633_1
  (
    .doutp(ffc_633_p),
    .doutn(ffc_633_n),
    .din(ffc_854_p_spl_)
  );


  DROC
  ffc_634_1
  (
    .doutp(ffc_634_p),
    .doutn(ffc_634_n),
    .din(ffc_856_p_spl_)
  );


  DROC
  ffc_635_1
  (
    .doutp(ffc_635_p),
    .doutn(ffc_635_n),
    .din(ffc_857_p_spl_)
  );


  DROC
  ffc_636_1
  (
    .doutp(ffc_636_p),
    .doutn(ffc_636_n),
    .din(ffc_858_p_spl_)
  );


  DROC
  ffc_637_1
  (
    .doutp(ffc_637_p),
    .doutn(ffc_637_n),
    .din(g1720_n_spl_)
  );


  DROC
  ffc_638_1
  (
    .doutp(ffc_638_p),
    .doutn(ffc_638_n),
    .din(g1721_n_spl_)
  );


  DROC
  ffc_639_1
  (
    .doutp(ffc_639_p),
    .doutn(ffc_639_n),
    .din(g1722_n_spl_)
  );


  DROC
  ffc_640_2
  (
    .doutp(ffc_640_p),
    .doutn(ffc_640_n),
    .din(ffc_355_p_spl_)
  );


  DROC
  ffc_641_3
  (
    .doutp(ffc_641_p),
    .doutn(ffc_641_n),
    .din(g1724_p_spl_)
  );


  DROC
  ffc_642_2
  (
    .doutp(ffc_642_p),
    .doutn(ffc_642_n),
    .din(g1725_p)
  );


  DROC
  ffc_643_3
  (
    .doutp(ffc_643_n),
    .doutn(ffc_643_p),
    .din(g1728_n_spl_)
  );


  DROC
  ffc_644_3
  (
    .doutp(ffc_644_p),
    .doutn(ffc_644_n),
    .din(g1737_n_spl_)
  );


  DROC
  ffc_645_3
  (
    .doutp(ffc_645_p),
    .doutn(ffc_645_n),
    .din(g1746_n_spl_)
  );


  DROC
  ffc_646_3
  (
    .doutp(ffc_646_p),
    .doutn(ffc_646_n),
    .din(g1755_n_spl_)
  );


  DROC
  ffc_647_2
  (
    .doutp(ffc_647_p),
    .doutn(ffc_647_n),
    .din(g1758_p_spl_)
  );


  DROC
  ffc_648_1
  (
    .doutp(ffc_648_p),
    .doutn(ffc_648_n),
    .din(ffc_846_p_spl_)
  );


  DROC
  ffc_649_1
  (
    .doutp(ffc_649_p),
    .doutn(ffc_649_n),
    .din(ffc_847_p_spl_)
  );


  DROC
  ffc_650_1
  (
    .doutp(ffc_650_p),
    .doutn(ffc_650_n),
    .din(ffc_848_p_spl_)
  );


  DROC
  ffc_651_1
  (
    .doutp(ffc_651_p),
    .doutn(ffc_651_n),
    .din(ffc_849_p_spl_)
  );


  DROC
  ffc_652_1
  (
    .doutp(ffc_652_p),
    .doutn(ffc_652_n),
    .din(g1761_n_spl_)
  );


  DROC
  ffc_653_1
  (
    .doutp(ffc_653_p),
    .doutn(ffc_653_n),
    .din(g1762_p_spl_)
  );


  DROC
  ffc_654_1
  (
    .doutp(ffc_654_p),
    .doutn(ffc_654_n),
    .din(g1763_n_spl_1)
  );


  DROC
  ffc_655_1
  (
    .doutp(ffc_655_p),
    .doutn(ffc_655_n),
    .din(g1764_p_spl_)
  );


  DROC
  ffc_656_1
  (
    .doutp(ffc_656_p),
    .doutn(ffc_656_n),
    .din(g1767_n_spl_)
  );


  DROC
  ffc_657_2
  (
    .doutp(ffc_657_p),
    .doutn(ffc_657_n),
    .din(ffc_358_p_spl_)
  );


  DROC
  ffc_658_2
  (
    .doutp(ffc_658_p),
    .doutn(ffc_658_n),
    .din(g1768_n_spl_)
  );


  DROC
  ffc_659_2
  (
    .doutp(ffc_659_p),
    .doutn(ffc_659_n),
    .din(g1774_n_spl_)
  );


  DROC
  ffc_660_1
  (
    .doutp(ffc_660_p),
    .doutn(ffc_660_n),
    .din(ffc_346_p_spl_)
  );


  DROC
  ffc_661_1
  (
    .doutp(ffc_661_p),
    .doutn(ffc_661_n),
    .din(ffc_366_p_spl_)
  );


  DROC
  ffc_662_1
  (
    .doutp(ffc_662_p),
    .doutn(ffc_662_n),
    .din(ffc_367_p_spl_)
  );


  DROC
  ffc_663_1
  (
    .doutp(ffc_663_p),
    .doutn(ffc_663_n),
    .din(ffc_388_p_spl_)
  );


  DROC
  ffc_664_1
  (
    .doutp(ffc_664_p),
    .doutn(ffc_664_n),
    .din(ffc_392_p_spl_)
  );


  DROC
  ffc_665_1
  (
    .doutp(ffc_665_p),
    .doutn(ffc_665_n),
    .din(ffc_393_p_spl_)
  );


  DROC
  ffc_666_1
  (
    .doutp(ffc_666_p),
    .doutn(ffc_666_n),
    .din(g1777_n_spl_)
  );


  DROC
  ffc_667_1
  (
    .doutp(ffc_667_p),
    .doutn(ffc_667_n),
    .din(g1780_n_spl_)
  );


  DROC
  ffc_668_2
  (
    .doutp(ffc_668_n),
    .doutn(ffc_668_p),
    .din(g1787_n_spl_)
  );


  DROC
  ffc_669_1
  (
    .doutp(ffc_669_p),
    .doutn(ffc_669_n),
    .din(g1790_n_spl_)
  );


  DROC
  ffc_670_2
  (
    .doutp(ffc_670_p),
    .doutn(ffc_670_n),
    .din(g1792_p_spl_)
  );


  DROC
  ffc_671_1
  (
    .doutp(ffc_671_p),
    .doutn(ffc_671_n),
    .din(g1793_p_spl_)
  );


  DROC
  ffc_672_1
  (
    .doutp(ffc_672_p),
    .doutn(ffc_672_n),
    .din(g1796_p_spl_)
  );


  DROC
  ffc_673_1
  (
    .doutp(ffc_673_p),
    .doutn(ffc_673_n),
    .din(g1797_p_spl_)
  );


  DROC
  ffc_674_1
  (
    .doutp(ffc_674_p),
    .doutn(ffc_674_n),
    .din(g1799_p_spl_)
  );


  DROC
  ffc_675_1
  (
    .doutp(ffc_675_p),
    .doutn(ffc_675_n),
    .din(ffc_334_p_spl_)
  );


  DROC
  ffc_676_1
  (
    .doutp(ffc_676_p),
    .doutn(ffc_676_n),
    .din(ffc_364_p_spl_)
  );


  DROC
  ffc_677_1
  (
    .doutp(ffc_677_p),
    .doutn(ffc_677_n),
    .din(ffc_370_p)
  );


  DROC
  ffc_678_1
  (
    .doutp(ffc_678_p),
    .doutn(ffc_678_n),
    .din(ffc_371_p)
  );


  DROC
  ffc_679_1
  (
    .doutp(ffc_679_p),
    .doutn(ffc_679_n),
    .din(ffc_397_p_spl_)
  );


  DROC
  ffc_680_1
  (
    .doutp(ffc_680_p),
    .doutn(ffc_680_n),
    .din(g1802_n_spl_)
  );


  DROC
  ffc_681_1
  (
    .doutp(ffc_681_p),
    .doutn(ffc_681_n),
    .din(g1803_p_spl_)
  );


  DROC
  ffc_682_1
  (
    .doutp(ffc_682_p),
    .doutn(ffc_682_n),
    .din(g1804_p_spl_)
  );


  DROC
  ffc_683_1
  (
    .doutp(ffc_683_p),
    .doutn(ffc_683_n),
    .din(g1805_p_spl_)
  );


  DROC
  ffc_684_1
  (
    .doutp(ffc_684_p),
    .doutn(ffc_684_n),
    .din(g1808_p_spl_)
  );


  DROC
  ffc_685_1
  (
    .doutp(ffc_685_p),
    .doutn(ffc_685_n),
    .din(g1809_p_spl_)
  );


  DROC
  ffc_686_3
  (
    .doutp(ffc_686_p),
    .doutn(ffc_686_n),
    .din(g1810_p)
  );


  DROC
  ffc_687_3
  (
    .doutp(ffc_687_p),
    .doutn(ffc_687_n),
    .din(g1811_p)
  );


  DROC
  ffc_688_3
  (
    .doutp(ffc_688_p),
    .doutn(ffc_688_n),
    .din(g1812_p)
  );


  DROC
  ffc_689_3
  (
    .doutp(ffc_689_p),
    .doutn(ffc_689_n),
    .din(g1813_n)
  );


  DROC
  ffc_690_3
  (
    .doutp(ffc_690_p),
    .doutn(ffc_690_n),
    .din(g1814_n)
  );


  DROC
  ffc_691_3
  (
    .doutp(ffc_691_p),
    .doutn(ffc_691_n),
    .din(g1815_p)
  );


  DROC
  ffc_692_3
  (
    .doutp(ffc_692_p),
    .doutn(ffc_692_n),
    .din(g1816_p)
  );


  DROC
  ffc_693_3
  (
    .doutp(ffc_693_p),
    .doutn(ffc_693_n),
    .din(g1817_n)
  );


  DROC
  ffc_694_3
  (
    .doutp(ffc_694_p),
    .doutn(ffc_694_n),
    .din(g1818_n)
  );


  DROC
  ffc_695_3
  (
    .doutp(ffc_695_p),
    .doutn(ffc_695_n),
    .din(g1822_p)
  );


  DROC
  ffc_696_3
  (
    .doutp(ffc_696_p),
    .doutn(ffc_696_n),
    .din(g1826_p)
  );


  DROC
  ffc_697_3
  (
    .doutp(ffc_697_p),
    .doutn(ffc_697_n),
    .din(g1827_p)
  );


  DROC
  ffc_698_3
  (
    .doutp(ffc_698_p),
    .doutn(ffc_698_n),
    .din(g1829_p)
  );


  DROC
  ffc_699_3
  (
    .doutp(ffc_699_p),
    .doutn(ffc_699_n),
    .din(g1847_p)
  );


  DROC
  ffc_700_3
  (
    .doutp(ffc_700_n),
    .doutn(ffc_700_p),
    .din(g1848_n)
  );


  DROC
  ffc_701_3
  (
    .doutp(ffc_701_n),
    .doutn(ffc_701_p),
    .din(g1849_n)
  );


  DROC
  ffc_702_3
  (
    .doutp(ffc_702_p),
    .doutn(ffc_702_n),
    .din(g1850_p)
  );


  DROC
  ffc_703_3
  (
    .doutp(ffc_703_p),
    .doutn(ffc_703_n),
    .din(g1851_p)
  );


  DROC
  ffc_704_3
  (
    .doutp(ffc_704_p),
    .doutn(ffc_704_n),
    .din(g1852_p)
  );


  DROC
  ffc_705_3
  (
    .doutp(ffc_705_n),
    .doutn(ffc_705_p),
    .din(g1853_n)
  );


  DROC
  ffc_706_3
  (
    .doutp(ffc_706_p),
    .doutn(ffc_706_n),
    .din(g1868_p)
  );


  DROC
  ffc_707_3
  (
    .doutp(ffc_707_p),
    .doutn(ffc_707_n),
    .din(g1869_p)
  );


  DROC
  ffc_708_3
  (
    .doutp(ffc_708_p),
    .doutn(ffc_708_n),
    .din(g1870_p)
  );


  DROC
  ffc_709_3
  (
    .doutp(ffc_709_p),
    .doutn(ffc_709_n),
    .din(g1873_p)
  );


  DROC
  ffc_710_3
  (
    .doutp(ffc_710_p),
    .doutn(ffc_710_n),
    .din(g1874_p)
  );


  DROC
  ffc_711_3
  (
    .doutp(ffc_711_n),
    .doutn(ffc_711_p),
    .din(g1878_n)
  );


  DROC
  ffc_712_3
  (
    .doutp(ffc_712_n),
    .doutn(ffc_712_p),
    .din(g1879_p)
  );


  DROC
  ffc_713_3
  (
    .doutp(ffc_713_p),
    .doutn(ffc_713_n),
    .din(g1880_n)
  );


  DROC
  ffc_714_3
  (
    .doutp(ffc_714_p),
    .doutn(ffc_714_n),
    .din(g1881_n)
  );


  DROC
  ffc_715_3
  (
    .doutp(ffc_715_p),
    .doutn(ffc_715_n),
    .din(g1885_n)
  );


  DROC
  ffc_716_3
  (
    .doutp(ffc_716_p),
    .doutn(ffc_716_n),
    .din(g1886_p)
  );


  DROC
  ffc_717_3
  (
    .doutp(ffc_717_p),
    .doutn(ffc_717_n),
    .din(g1887_n)
  );


  DROC
  ffc_718_3
  (
    .doutp(ffc_718_p),
    .doutn(ffc_718_n),
    .din(g1888_p)
  );


  DROC
  ffc_719_3
  (
    .doutp(ffc_719_p),
    .doutn(ffc_719_n),
    .din(g1889_n)
  );


  DROC
  ffc_720_3
  (
    .doutp(ffc_720_n),
    .doutn(ffc_720_p),
    .din(g1892_p)
  );


  DROC
  ffc_721_3
  (
    .doutp(ffc_721_n),
    .doutn(ffc_721_p),
    .din(g1893_n)
  );


  DROC
  ffc_722_3
  (
    .doutp(ffc_722_n),
    .doutn(ffc_722_p),
    .din(g1894_n)
  );


  DROC
  ffc_723_3
  (
    .doutp(ffc_723_p),
    .doutn(ffc_723_n),
    .din(g1897_p)
  );


  DROC
  ffc_724_1
  (
    .doutp(ffc_724_p),
    .doutn(ffc_724_n),
    .din(g1898_n_spl_)
  );


  DROC
  ffc_725_3
  (
    .doutp(ffc_725_p),
    .doutn(ffc_725_n),
    .din(g1901_n)
  );


  DROC
  ffc_726_3
  (
    .doutp(ffc_726_p),
    .doutn(ffc_726_n),
    .din(g1904_n)
  );


  DROC
  ffc_727_3
  (
    .doutp(ffc_727_n),
    .doutn(ffc_727_p),
    .din(g1907_p)
  );


  DROC
  ffc_728_3
  (
    .doutp(ffc_728_p),
    .doutn(ffc_728_n),
    .din(g1910_p)
  );


  DROC
  ffc_729_3
  (
    .doutp(ffc_729_p),
    .doutn(ffc_729_n),
    .din(g1913_n)
  );


  DROC
  ffc_730_3
  (
    .doutp(ffc_730_p),
    .doutn(ffc_730_n),
    .din(g1916_n)
  );


  DROC
  ffc_731_3
  (
    .doutp(ffc_731_p),
    .doutn(ffc_731_n),
    .din(g1925_n)
  );


  DROC
  ffc_732_3
  (
    .doutp(ffc_732_p),
    .doutn(ffc_732_n),
    .din(g1934_n)
  );


  DROC
  ffc_733_3
  (
    .doutp(ffc_733_p),
    .doutn(ffc_733_n),
    .din(g1943_n)
  );


  DROC
  ffc_734_3
  (
    .doutp(ffc_734_p),
    .doutn(ffc_734_n),
    .din(g1952_n)
  );


  DROC
  ffc_735_3
  (
    .doutp(ffc_735_p),
    .doutn(ffc_735_n),
    .din(g1961_n)
  );


  DROC
  ffc_736_3
  (
    .doutp(ffc_736_p),
    .doutn(ffc_736_n),
    .din(g1970_n)
  );


  DROC
  ffc_737_3
  (
    .doutp(ffc_737_p),
    .doutn(ffc_737_n),
    .din(g1979_n)
  );


  DROC
  ffc_738_3
  (
    .doutp(ffc_738_p),
    .doutn(ffc_738_n),
    .din(g2001_p)
  );


  DROC
  ffc_739_3
  (
    .doutp(ffc_739_p),
    .doutn(ffc_739_n),
    .din(g2004_n)
  );


  DROC
  ffc_740_3
  (
    .doutp(ffc_740_p),
    .doutn(ffc_740_n),
    .din(g2007_p)
  );


  DROC
  ffc_741_3
  (
    .doutp(ffc_741_p),
    .doutn(ffc_741_n),
    .din(g2011_p)
  );


  DROC
  ffc_742_3
  (
    .doutp(ffc_742_p),
    .doutn(ffc_742_n),
    .din(g2017_p)
  );


  DROC
  ffc_743_3
  (
    .doutp(ffc_743_p),
    .doutn(ffc_743_n),
    .din(g2020_n)
  );


  DROC
  ffc_744_3
  (
    .doutp(ffc_744_p),
    .doutn(ffc_744_n),
    .din(g2023_p)
  );


  DROC
  ffc_745_3
  (
    .doutp(ffc_745_p),
    .doutn(ffc_745_n),
    .din(g2029_n)
  );


  DROC
  ffc_746_3
  (
    .doutp(ffc_746_p),
    .doutn(ffc_746_n),
    .din(g2032_n)
  );


  DROC
  ffc_747_3
  (
    .doutp(ffc_747_p),
    .doutn(ffc_747_n),
    .din(g2039_p)
  );


  DROC
  ffc_748_3
  (
    .doutp(ffc_748_n),
    .doutn(ffc_748_p),
    .din(g2040_n)
  );


  DROC
  ffc_749_3
  (
    .doutp(ffc_749_p),
    .doutn(ffc_749_n),
    .din(g2050_p)
  );


  DROC
  ffc_750_3
  (
    .doutp(ffc_750_n),
    .doutn(ffc_750_p),
    .din(g2051_n)
  );


  DROC
  ffc_751_3
  (
    .doutp(ffc_751_p),
    .doutn(ffc_751_n),
    .din(g2058_n)
  );


  DROC
  ffc_752_3
  (
    .doutp(ffc_752_p),
    .doutn(ffc_752_n),
    .din(g2059_p)
  );


  DROC
  ffc_753_3
  (
    .doutp(ffc_753_p),
    .doutn(ffc_753_n),
    .din(g2068_p)
  );


  DROC
  ffc_754_3
  (
    .doutp(ffc_754_p),
    .doutn(ffc_754_n),
    .din(g2095_p)
  );


  DROC
  ffc_755_1
  (
    .doutp(ffc_755_p),
    .doutn(ffc_755_n),
    .din(g2096_n_spl_)
  );


  DROC
  ffc_756_1
  (
    .doutp(ffc_756_p),
    .doutn(ffc_756_n),
    .din(g2098_n_spl_)
  );


  DROC
  ffc_757_1
  (
    .doutp(ffc_757_p),
    .doutn(ffc_757_n),
    .din(g2099_p_spl_)
  );


  DROC
  ffc_758_2
  (
    .doutp(ffc_758_p),
    .doutn(ffc_758_n),
    .din(g2108_n_spl_)
  );


  DROC
  ffc_759_2
  (
    .doutp(ffc_759_p),
    .doutn(ffc_759_n),
    .din(g2117_n_spl_)
  );


  DROC
  ffc_760_2
  (
    .doutp(ffc_760_n),
    .doutn(ffc_760_p),
    .din(g2120_n_spl_)
  );


  DROC
  ffc_761_2
  (
    .doutp(ffc_761_n),
    .doutn(ffc_761_p),
    .din(g2123_n_spl_)
  );


  DROC
  ffc_762_2
  (
    .doutp(ffc_762_p),
    .doutn(ffc_762_n),
    .din(g2126_p_spl_)
  );


  DROC
  ffc_763_1
  (
    .doutp(ffc_763_p),
    .doutn(ffc_763_n),
    .din(ffc_387_p_spl_)
  );


  DROC
  ffc_764_1
  (
    .doutp(ffc_764_p),
    .doutn(ffc_764_n),
    .din(ffc_395_p_spl_)
  );


  DROC
  ffc_765_1
  (
    .doutp(ffc_765_p),
    .doutn(ffc_765_n),
    .din(ffc_396_p_spl_)
  );


  DROC
  ffc_766_1
  (
    .doutp(ffc_766_p),
    .doutn(ffc_766_n),
    .din(g2129_n_spl_)
  );


  DROC
  ffc_767_1
  (
    .doutp(ffc_767_p),
    .doutn(ffc_767_n),
    .din(g2132_n_spl_)
  );


  DROC
  ffc_768_1
  (
    .doutp(ffc_768_n),
    .doutn(ffc_768_p),
    .din(g2133_n_spl_)
  );


  DROC
  ffc_769_1
  (
    .doutp(ffc_769_p),
    .doutn(ffc_769_n),
    .din(g2135_p_spl_)
  );


  DROC
  ffc_770_1
  (
    .doutp(ffc_770_p),
    .doutn(ffc_770_n),
    .din(g2137_p_spl_1)
  );


  DROC
  ffc_771_2
  (
    .doutp(ffc_771_p),
    .doutn(ffc_771_n),
    .din(g2141_n)
  );


  DROC
  ffc_772_2
  (
    .doutp(ffc_772_n),
    .doutn(ffc_772_p),
    .din(g2143_n)
  );


  DROC
  ffc_773_2
  (
    .doutp(ffc_773_n),
    .doutn(ffc_773_p),
    .din(g2158_p)
  );


  DROC
  ffc_774_2
  (
    .doutp(ffc_774_n),
    .doutn(ffc_774_p),
    .din(g2159_n)
  );


  DROC
  ffc_775_1
  (
    .doutp(ffc_775_p),
    .doutn(ffc_775_n),
    .din(g2160_n_spl_)
  );


  DROC
  ffc_776_2
  (
    .doutp(ffc_776_p),
    .doutn(ffc_776_n),
    .din(g2173_p)
  );


  DROC
  ffc_777_2
  (
    .doutp(ffc_777_p),
    .doutn(ffc_777_n),
    .din(g2174_n)
  );


  DROC
  ffc_778_1
  (
    .doutp(ffc_778_p),
    .doutn(ffc_778_n),
    .din(g2175_p_spl_)
  );


  DROC
  ffc_779_1
  (
    .doutp(ffc_779_p),
    .doutn(ffc_779_n),
    .din(g2177_n_spl_)
  );


  DROC
  ffc_780_1
  (
    .doutp(ffc_780_p),
    .doutn(ffc_780_n),
    .din(ffc_360_p_spl_)
  );


  DROC
  ffc_781_1
  (
    .doutp(ffc_781_p),
    .doutn(ffc_781_n),
    .din(ffc_362_p_spl_)
  );


  DROC
  ffc_782_1
  (
    .doutp(ffc_782_p),
    .doutn(ffc_782_n),
    .din(ffc_391_p_spl_)
  );


  DROC
  ffc_783_2
  (
    .doutp(ffc_783_p),
    .doutn(ffc_783_n),
    .din(g2180_n)
  );


  DROC
  ffc_784_2
  (
    .doutp(ffc_784_p),
    .doutn(ffc_784_n),
    .din(g2189_n)
  );


  DROC
  ffc_785_2
  (
    .doutp(ffc_785_p),
    .doutn(ffc_785_n),
    .din(g2198_n)
  );


  DROC
  ffc_786_2
  (
    .doutp(ffc_786_p),
    .doutn(ffc_786_n),
    .din(g2207_n)
  );


  DROC
  ffc_787_2
  (
    .doutp(ffc_787_p),
    .doutn(ffc_787_n),
    .din(g2216_n)
  );


  DROC
  ffc_788_2
  (
    .doutp(ffc_788_p),
    .doutn(ffc_788_n),
    .din(g2225_n)
  );


  DROC
  ffc_789_2
  (
    .doutp(ffc_789_p),
    .doutn(ffc_789_n),
    .din(g2234_n)
  );


  DROC
  ffc_790_2
  (
    .doutp(ffc_790_p),
    .doutn(ffc_790_n),
    .din(g2243_n)
  );


  DROC
  ffc_791_2
  (
    .doutp(ffc_791_p),
    .doutn(ffc_791_n),
    .din(g2249_n)
  );


  DROC
  ffc_792_2
  (
    .doutp(ffc_792_n),
    .doutn(ffc_792_p),
    .din(g2260_n)
  );


  DROC
  ffc_793_2
  (
    .doutp(ffc_793_n),
    .doutn(ffc_793_p),
    .din(g2261_p)
  );


  DROC
  ffc_794_1
  (
    .doutp(ffc_794_p),
    .doutn(ffc_794_n),
    .din(g2264_n_spl_)
  );


  DROC
  ffc_795_1
  (
    .doutp(ffc_795_n),
    .doutn(ffc_795_p),
    .din(g2267_p_spl_)
  );


  DROC
  ffc_796_1
  (
    .doutp(ffc_796_n),
    .doutn(ffc_796_p),
    .din(g2268_n_spl_)
  );


  DROC
  ffc_797_2
  (
    .doutp(ffc_797_p),
    .doutn(ffc_797_n),
    .din(g2273_n)
  );


  DROC
  ffc_798_2
  (
    .doutp(ffc_798_p),
    .doutn(ffc_798_n),
    .din(g2274_p)
  );


  DROC
  ffc_799_1
  (
    .doutp(ffc_799_p),
    .doutn(ffc_799_n),
    .din(g2276_n_spl_)
  );


  DROC
  ffc_800_2
  (
    .doutp(ffc_800_p),
    .doutn(ffc_800_n),
    .din(g2277_p)
  );


  DROC
  ffc_801_2
  (
    .doutp(ffc_801_n),
    .doutn(ffc_801_p),
    .din(g2278_n)
  );


  DROC
  ffc_802_2
  (
    .doutp(ffc_802_p),
    .doutn(ffc_802_n),
    .din(g2279_p)
  );


  DROC
  ffc_803_2
  (
    .doutp(ffc_803_p),
    .doutn(ffc_803_n),
    .din(g2280_n)
  );


  DROC
  ffc_804_2
  (
    .doutp(ffc_804_n),
    .doutn(ffc_804_p),
    .din(g2296_n)
  );


  DROC
  ffc_805_2
  (
    .doutp(ffc_805_p),
    .doutn(ffc_805_n),
    .din(g2297_p)
  );


  DROC
  ffc_806_2
  (
    .doutp(ffc_806_n),
    .doutn(ffc_806_p),
    .din(g2316_n)
  );


  DROC
  ffc_807_2
  (
    .doutp(ffc_807_p),
    .doutn(ffc_807_n),
    .din(g2317_p)
  );


  DROC
  ffc_808_2
  (
    .doutp(ffc_808_n),
    .doutn(ffc_808_p),
    .din(g2325_n)
  );


  DROC
  ffc_809_2
  (
    .doutp(ffc_809_p),
    .doutn(ffc_809_n),
    .din(g2333_p)
  );


  DROC
  ffc_810_2
  (
    .doutp(ffc_810_p),
    .doutn(ffc_810_n),
    .din(g2354_n)
  );


  DROC
  ffc_811_2
  (
    .doutp(ffc_811_p),
    .doutn(ffc_811_n),
    .din(g2360_n)
  );


  DROC
  ffc_812_1
  (
    .doutp(ffc_812_n),
    .doutn(ffc_812_p),
    .din(g2361_n_spl_)
  );


  DROC
  ffc_813_1
  (
    .doutp(ffc_813_n),
    .doutn(ffc_813_p),
    .din(g2362_n_spl_)
  );


  DROC
  ffc_814_1
  (
    .doutp(ffc_814_p),
    .doutn(ffc_814_n),
    .din(g2363_n_spl_)
  );


  DROC
  ffc_815_1
  (
    .doutp(ffc_815_p),
    .doutn(ffc_815_n),
    .din(g2365_p_spl_)
  );


  DROC
  ffc_816_1
  (
    .doutp(ffc_816_p),
    .doutn(ffc_816_n),
    .din(ffc_394_p)
  );


  DROC
  ffc_817_1
  (
    .doutp(ffc_817_p),
    .doutn(ffc_817_n),
    .din(g2366_p)
  );


  DROC
  ffc_818_1
  (
    .doutp(ffc_818_p),
    .doutn(ffc_818_n),
    .din(g2367_p)
  );


  DROC
  ffc_819_1
  (
    .doutp(ffc_819_p),
    .doutn(ffc_819_n),
    .din(g2368_p)
  );


  DROC
  ffc_820_1
  (
    .doutp(ffc_820_p),
    .doutn(ffc_820_n),
    .din(g2369_p)
  );


  DROC
  ffc_821_1
  (
    .doutp(ffc_821_p),
    .doutn(ffc_821_n),
    .din(g2370_p)
  );


  DROC
  ffc_822_1
  (
    .doutp(ffc_822_p),
    .doutn(ffc_822_n),
    .din(g2371_n)
  );


  DROC
  ffc_823_1
  (
    .doutp(ffc_823_p),
    .doutn(ffc_823_n),
    .din(g2372_p)
  );


  DROC
  ffc_824_1
  (
    .doutp(ffc_824_p),
    .doutn(ffc_824_n),
    .din(g2373_p)
  );


  DROC
  ffc_825_1
  (
    .doutp(ffc_825_p),
    .doutn(ffc_825_n),
    .din(g2374_p)
  );


  DROC
  ffc_826_1
  (
    .doutp(ffc_826_p),
    .doutn(ffc_826_n),
    .din(g2376_n)
  );


  DROC
  ffc_827_1
  (
    .doutp(ffc_827_p),
    .doutn(ffc_827_n),
    .din(g2378_n)
  );


  DROC
  ffc_828_1
  (
    .doutp(ffc_828_p),
    .doutn(ffc_828_n),
    .din(g2379_p)
  );


  DROC
  ffc_829_1
  (
    .doutp(ffc_829_p),
    .doutn(ffc_829_n),
    .din(ffc_336_p)
  );


  DROC
  ffc_830_1
  (
    .doutp(ffc_830_p),
    .doutn(ffc_830_n),
    .din(ffc_337_p)
  );


  DROC
  ffc_831_1
  (
    .doutp(ffc_831_p),
    .doutn(ffc_831_n),
    .din(ffc_338_p)
  );


  DROC
  ffc_832_1
  (
    .doutp(ffc_832_p),
    .doutn(ffc_832_n),
    .din(ffc_343_p)
  );


  DROC
  ffc_833_1
  (
    .doutp(ffc_833_p),
    .doutn(ffc_833_n),
    .din(ffc_344_p)
  );


  DROC
  ffc_834_1
  (
    .doutp(ffc_834_p),
    .doutn(ffc_834_n),
    .din(ffc_345_p)
  );


  DROC
  ffc_835_1
  (
    .doutp(ffc_835_p),
    .doutn(ffc_835_n),
    .din(g2380_n)
  );


  DROC
  ffc_836_0
  (
    .doutp(ffc_836_p),
    .doutn(ffc_836_n),
    .din(G92_p_spl_)
  );


  DROC
  ffc_837_0
  (
    .doutp(ffc_837_p),
    .doutn(ffc_837_n),
    .din(G94_p_spl_)
  );


  DROC
  ffc_838_0
  (
    .doutp(ffc_838_p),
    .doutn(ffc_838_n),
    .din(G107_p_spl_)
  );


  DROC
  ffc_839_0
  (
    .doutp(ffc_839_p),
    .doutn(ffc_839_n),
    .din(G124_p_spl_1)
  );


  DROC
  ffc_840_1
  (
    .doutp(ffc_840_p),
    .doutn(ffc_840_n),
    .din(g2381_p)
  );


  DROC
  ffc_841_1
  (
    .doutp(ffc_841_p),
    .doutn(ffc_841_n),
    .din(g2382_n)
  );


  DROC
  ffc_842_1
  (
    .doutp(ffc_842_p),
    .doutn(ffc_842_n),
    .din(g2383_p)
  );


  DROC
  ffc_843_1
  (
    .doutp(ffc_843_p),
    .doutn(ffc_843_n),
    .din(g2385_p)
  );


  DROC
  ffc_844_1
  (
    .doutp(ffc_844_p),
    .doutn(ffc_844_n),
    .din(g2387_p)
  );


  DROC
  ffc_845_1
  (
    .doutp(ffc_845_p),
    .doutn(ffc_845_n),
    .din(g2388_p)
  );


  DROC
  ffc_846_0
  (
    .doutp(ffc_846_p),
    .doutn(ffc_846_n),
    .din(G128_p)
  );


  DROC
  ffc_847_0
  (
    .doutp(ffc_847_p),
    .doutn(ffc_847_n),
    .din(G129_p)
  );


  DROC
  ffc_848_0
  (
    .doutp(ffc_848_p),
    .doutn(ffc_848_n),
    .din(G135_p)
  );


  DROC
  ffc_849_0
  (
    .doutp(ffc_849_p),
    .doutn(ffc_849_n),
    .din(G145_p)
  );


  DROC
  ffc_850_0
  (
    .doutp(ffc_850_p),
    .doutn(ffc_850_n),
    .din(G90_p)
  );


  DROC
  ffc_851_0
  (
    .doutp(ffc_851_p),
    .doutn(ffc_851_n),
    .din(G91_p)
  );


  DROC
  ffc_852_0
  (
    .doutp(ffc_852_p),
    .doutn(ffc_852_n),
    .din(G105_p)
  );


  DROC
  ffc_853_0
  (
    .doutp(ffc_853_p),
    .doutn(ffc_853_n),
    .din(G106_p)
  );


  DROC
  ffc_854_0
  (
    .doutp(ffc_854_p),
    .doutn(ffc_854_n),
    .din(G119_p)
  );


  DROC
  ffc_855_0
  (
    .doutp(ffc_855_p),
    .doutn(ffc_855_n),
    .din(G120_p)
  );


  DROC
  ffc_856_0
  (
    .doutp(ffc_856_p),
    .doutn(ffc_856_n),
    .din(G139_p)
  );


  DROC
  ffc_857_0
  (
    .doutp(ffc_857_p),
    .doutn(ffc_857_n),
    .din(G140_p)
  );


  DROC
  ffc_858_0
  (
    .doutp(ffc_858_p),
    .doutn(ffc_858_n),
    .din(G144_p)
  );


  DROC
  ffc_859_0
  (
    .doutp(ffc_859_p),
    .doutn(ffc_859_n),
    .din(G109_p)
  );


  DROC
  ffc_860_0
  (
    .doutp(ffc_860_p),
    .doutn(ffc_860_n),
    .din(G110_p)
  );


  DROC
  ffc_861_0
  (
    .doutp(ffc_861_p),
    .doutn(ffc_861_n),
    .din(G117_p)
  );


  DROC
  ffc_862_0
  (
    .doutp(ffc_862_p),
    .doutn(ffc_862_n),
    .din(G118_p)
  );


  DROC
  ffc_863_0
  (
    .doutp(ffc_863_p),
    .doutn(ffc_863_n),
    .din(G123_p)
  );


  DROC
  ffc_864_0
  (
    .doutp(ffc_864_p),
    .doutn(ffc_864_n),
    .din(g2389_p)
  );


  DROC
  ffc_865_0
  (
    .doutp(ffc_865_p),
    .doutn(ffc_865_n),
    .din(g2390_p)
  );


  DROC
  ffc_866_0
  (
    .doutp(ffc_866_p),
    .doutn(ffc_866_n),
    .din(g2391_p)
  );


  DROC
  ffc_867_0
  (
    .doutp(ffc_867_p),
    .doutn(ffc_867_n),
    .din(g2392_p)
  );


  DROC
  ffc_868_0
  (
    .doutp(ffc_868_p),
    .doutn(ffc_868_n),
    .din(g2393_p)
  );


  DROC
  ffc_869_0
  (
    .doutp(ffc_869_p),
    .doutn(ffc_869_n),
    .din(g2394_p)
  );


  buf

  (
    ffc_409_n_spl_,
    ffc_409_n
  );


  buf

  (
    ffc_421_n_spl_,
    ffc_421_n
  );


  buf

  (
    ffc_249_p_spl_,
    ffc_249_p
  );


  buf

  (
    ffc_249_p_spl_0,
    ffc_249_p_spl_
  );


  buf

  (
    ffc_249_p_spl_00,
    ffc_249_p_spl_0
  );


  buf

  (
    ffc_249_p_spl_01,
    ffc_249_p_spl_0
  );


  buf

  (
    ffc_249_p_spl_1,
    ffc_249_p_spl_
  );


  buf

  (
    ffc_3_p_spl_,
    ffc_3_p
  );


  buf

  (
    ffc_454_n_spl_,
    ffc_454_n
  );


  buf

  (
    ffc_42_n_spl_,
    ffc_42_n
  );


  buf

  (
    g1055_n_spl_,
    g1055_n
  );


  buf

  (
    g1055_n_spl_0,
    g1055_n_spl_
  );


  buf

  (
    g1055_n_spl_00,
    g1055_n_spl_0
  );


  buf

  (
    g1055_n_spl_000,
    g1055_n_spl_00
  );


  buf

  (
    g1055_n_spl_01,
    g1055_n_spl_0
  );


  buf

  (
    g1055_n_spl_1,
    g1055_n_spl_
  );


  buf

  (
    g1055_n_spl_10,
    g1055_n_spl_1
  );


  buf

  (
    g1055_n_spl_11,
    g1055_n_spl_1
  );


  buf

  (
    ffc_446_n_spl_,
    ffc_446_n
  );


  buf

  (
    ffc_446_n_spl_0,
    ffc_446_n_spl_
  );


  buf

  (
    ffc_446_n_spl_00,
    ffc_446_n_spl_0
  );


  buf

  (
    ffc_446_n_spl_01,
    ffc_446_n_spl_0
  );


  buf

  (
    ffc_446_n_spl_1,
    ffc_446_n_spl_
  );


  buf

  (
    ffc_446_p_spl_,
    ffc_446_p
  );


  buf

  (
    ffc_446_p_spl_0,
    ffc_446_p_spl_
  );


  buf

  (
    ffc_446_p_spl_00,
    ffc_446_p_spl_0
  );


  buf

  (
    ffc_446_p_spl_01,
    ffc_446_p_spl_0
  );


  buf

  (
    ffc_446_p_spl_1,
    ffc_446_p_spl_
  );


  buf

  (
    ffc_737_p_spl_,
    ffc_737_p
  );


  buf

  (
    g1094_n_spl_,
    g1094_n
  );


  buf

  (
    ffc_519_n_spl_,
    ffc_519_n
  );


  buf

  (
    g1101_n_spl_,
    g1101_n
  );


  buf

  (
    ffc_728_p_spl_,
    ffc_728_p
  );


  buf

  (
    ffc_729_p_spl_,
    ffc_729_p
  );


  buf

  (
    ffc_728_n_spl_,
    ffc_728_n
  );


  buf

  (
    ffc_729_n_spl_,
    ffc_729_n
  );


  buf

  (
    ffc_730_n_spl_,
    ffc_730_n
  );


  buf

  (
    ffc_753_n_spl_,
    ffc_753_n
  );


  buf

  (
    ffc_730_p_spl_,
    ffc_730_p
  );


  buf

  (
    ffc_753_p_spl_,
    ffc_753_p
  );


  buf

  (
    ffc_532_p_spl_,
    ffc_532_p
  );


  buf

  (
    ffc_532_p_spl_0,
    ffc_532_p_spl_
  );


  buf

  (
    ffc_697_p_spl_,
    ffc_697_p
  );


  buf

  (
    ffc_697_p_spl_0,
    ffc_697_p_spl_
  );


  buf

  (
    ffc_697_p_spl_00,
    ffc_697_p_spl_0
  );


  buf

  (
    ffc_697_p_spl_000,
    ffc_697_p_spl_00
  );


  buf

  (
    ffc_697_p_spl_001,
    ffc_697_p_spl_00
  );


  buf

  (
    ffc_697_p_spl_01,
    ffc_697_p_spl_0
  );


  buf

  (
    ffc_697_p_spl_010,
    ffc_697_p_spl_01
  );


  buf

  (
    ffc_697_p_spl_011,
    ffc_697_p_spl_01
  );


  buf

  (
    ffc_697_p_spl_1,
    ffc_697_p_spl_
  );


  buf

  (
    ffc_697_p_spl_10,
    ffc_697_p_spl_1
  );


  buf

  (
    ffc_697_p_spl_100,
    ffc_697_p_spl_10
  );


  buf

  (
    ffc_697_p_spl_101,
    ffc_697_p_spl_10
  );


  buf

  (
    ffc_697_p_spl_11,
    ffc_697_p_spl_1
  );


  buf

  (
    ffc_697_p_spl_110,
    ffc_697_p_spl_11
  );


  buf

  (
    ffc_697_p_spl_111,
    ffc_697_p_spl_11
  );


  buf

  (
    ffc_498_n_spl_,
    ffc_498_n
  );


  buf

  (
    ffc_498_n_spl_0,
    ffc_498_n_spl_
  );


  buf

  (
    ffc_498_n_spl_00,
    ffc_498_n_spl_0
  );


  buf

  (
    ffc_498_n_spl_000,
    ffc_498_n_spl_00
  );


  buf

  (
    ffc_498_n_spl_01,
    ffc_498_n_spl_0
  );


  buf

  (
    ffc_498_n_spl_1,
    ffc_498_n_spl_
  );


  buf

  (
    ffc_498_n_spl_10,
    ffc_498_n_spl_1
  );


  buf

  (
    ffc_498_n_spl_11,
    ffc_498_n_spl_1
  );


  buf

  (
    ffc_494_p_spl_,
    ffc_494_p
  );


  buf

  (
    ffc_494_p_spl_0,
    ffc_494_p_spl_
  );


  buf

  (
    ffc_494_p_spl_00,
    ffc_494_p_spl_0
  );


  buf

  (
    ffc_494_p_spl_000,
    ffc_494_p_spl_00
  );


  buf

  (
    ffc_494_p_spl_001,
    ffc_494_p_spl_00
  );


  buf

  (
    ffc_494_p_spl_01,
    ffc_494_p_spl_0
  );


  buf

  (
    ffc_494_p_spl_010,
    ffc_494_p_spl_01
  );


  buf

  (
    ffc_494_p_spl_011,
    ffc_494_p_spl_01
  );


  buf

  (
    ffc_494_p_spl_1,
    ffc_494_p_spl_
  );


  buf

  (
    ffc_494_p_spl_10,
    ffc_494_p_spl_1
  );


  buf

  (
    ffc_494_p_spl_100,
    ffc_494_p_spl_10
  );


  buf

  (
    ffc_494_p_spl_101,
    ffc_494_p_spl_10
  );


  buf

  (
    ffc_494_p_spl_11,
    ffc_494_p_spl_1
  );


  buf

  (
    ffc_494_p_spl_110,
    ffc_494_p_spl_11
  );


  buf

  (
    ffc_697_n_spl_,
    ffc_697_n
  );


  buf

  (
    ffc_498_p_spl_,
    ffc_498_p
  );


  buf

  (
    ffc_498_p_spl_0,
    ffc_498_p_spl_
  );


  buf

  (
    ffc_498_p_spl_00,
    ffc_498_p_spl_0
  );


  buf

  (
    ffc_498_p_spl_000,
    ffc_498_p_spl_00
  );


  buf

  (
    ffc_498_p_spl_01,
    ffc_498_p_spl_0
  );


  buf

  (
    ffc_498_p_spl_1,
    ffc_498_p_spl_
  );


  buf

  (
    ffc_498_p_spl_10,
    ffc_498_p_spl_1
  );


  buf

  (
    ffc_498_p_spl_11,
    ffc_498_p_spl_1
  );


  buf

  (
    ffc_494_n_spl_,
    ffc_494_n
  );


  buf

  (
    ffc_494_n_spl_0,
    ffc_494_n_spl_
  );


  buf

  (
    ffc_494_n_spl_1,
    ffc_494_n_spl_
  );


  buf

  (
    ffc_723_p_spl_,
    ffc_723_p
  );


  buf

  (
    ffc_482_n_spl_,
    ffc_482_n
  );


  buf

  (
    ffc_482_n_spl_0,
    ffc_482_n_spl_
  );


  buf

  (
    ffc_482_n_spl_00,
    ffc_482_n_spl_0
  );


  buf

  (
    ffc_482_n_spl_000,
    ffc_482_n_spl_00
  );


  buf

  (
    ffc_482_n_spl_0000,
    ffc_482_n_spl_000
  );


  buf

  (
    ffc_482_n_spl_0001,
    ffc_482_n_spl_000
  );


  buf

  (
    ffc_482_n_spl_001,
    ffc_482_n_spl_00
  );


  buf

  (
    ffc_482_n_spl_0010,
    ffc_482_n_spl_001
  );


  buf

  (
    ffc_482_n_spl_0011,
    ffc_482_n_spl_001
  );


  buf

  (
    ffc_482_n_spl_01,
    ffc_482_n_spl_0
  );


  buf

  (
    ffc_482_n_spl_010,
    ffc_482_n_spl_01
  );


  buf

  (
    ffc_482_n_spl_011,
    ffc_482_n_spl_01
  );


  buf

  (
    ffc_482_n_spl_1,
    ffc_482_n_spl_
  );


  buf

  (
    ffc_482_n_spl_10,
    ffc_482_n_spl_1
  );


  buf

  (
    ffc_482_n_spl_100,
    ffc_482_n_spl_10
  );


  buf

  (
    ffc_482_n_spl_101,
    ffc_482_n_spl_10
  );


  buf

  (
    ffc_482_n_spl_11,
    ffc_482_n_spl_1
  );


  buf

  (
    ffc_482_n_spl_110,
    ffc_482_n_spl_11
  );


  buf

  (
    ffc_482_n_spl_111,
    ffc_482_n_spl_11
  );


  buf

  (
    g1132_n_spl_,
    g1132_n
  );


  buf

  (
    g1132_n_spl_0,
    g1132_n_spl_
  );


  buf

  (
    g1132_n_spl_00,
    g1132_n_spl_0
  );


  buf

  (
    g1132_n_spl_1,
    g1132_n_spl_
  );


  buf

  (
    ffc_482_p_spl_,
    ffc_482_p
  );


  buf

  (
    ffc_482_p_spl_0,
    ffc_482_p_spl_
  );


  buf

  (
    ffc_482_p_spl_00,
    ffc_482_p_spl_0
  );


  buf

  (
    ffc_482_p_spl_000,
    ffc_482_p_spl_00
  );


  buf

  (
    ffc_482_p_spl_0000,
    ffc_482_p_spl_000
  );


  buf

  (
    ffc_482_p_spl_0001,
    ffc_482_p_spl_000
  );


  buf

  (
    ffc_482_p_spl_001,
    ffc_482_p_spl_00
  );


  buf

  (
    ffc_482_p_spl_0010,
    ffc_482_p_spl_001
  );


  buf

  (
    ffc_482_p_spl_0011,
    ffc_482_p_spl_001
  );


  buf

  (
    ffc_482_p_spl_01,
    ffc_482_p_spl_0
  );


  buf

  (
    ffc_482_p_spl_010,
    ffc_482_p_spl_01
  );


  buf

  (
    ffc_482_p_spl_011,
    ffc_482_p_spl_01
  );


  buf

  (
    ffc_482_p_spl_1,
    ffc_482_p_spl_
  );


  buf

  (
    ffc_482_p_spl_10,
    ffc_482_p_spl_1
  );


  buf

  (
    ffc_482_p_spl_100,
    ffc_482_p_spl_10
  );


  buf

  (
    ffc_482_p_spl_101,
    ffc_482_p_spl_10
  );


  buf

  (
    ffc_482_p_spl_11,
    ffc_482_p_spl_1
  );


  buf

  (
    ffc_482_p_spl_110,
    ffc_482_p_spl_11
  );


  buf

  (
    ffc_482_p_spl_111,
    ffc_482_p_spl_11
  );


  buf

  (
    g1142_n_spl_,
    g1142_n
  );


  buf

  (
    g1142_n_spl_0,
    g1142_n_spl_
  );


  buf

  (
    g1142_n_spl_00,
    g1142_n_spl_0
  );


  buf

  (
    g1142_n_spl_1,
    g1142_n_spl_
  );


  buf

  (
    ffc_478_p_spl_,
    ffc_478_p
  );


  buf

  (
    ffc_478_p_spl_0,
    ffc_478_p_spl_
  );


  buf

  (
    ffc_478_p_spl_00,
    ffc_478_p_spl_0
  );


  buf

  (
    ffc_478_p_spl_000,
    ffc_478_p_spl_00
  );


  buf

  (
    ffc_478_p_spl_001,
    ffc_478_p_spl_00
  );


  buf

  (
    ffc_478_p_spl_01,
    ffc_478_p_spl_0
  );


  buf

  (
    ffc_478_p_spl_1,
    ffc_478_p_spl_
  );


  buf

  (
    ffc_478_p_spl_10,
    ffc_478_p_spl_1
  );


  buf

  (
    ffc_478_p_spl_11,
    ffc_478_p_spl_1
  );


  buf

  (
    ffc_10_p_spl_,
    ffc_10_p
  );


  buf

  (
    ffc_84_p_spl_,
    ffc_84_p
  );


  buf

  (
    ffc_478_n_spl_,
    ffc_478_n
  );


  buf

  (
    ffc_478_n_spl_0,
    ffc_478_n_spl_
  );


  buf

  (
    ffc_478_n_spl_00,
    ffc_478_n_spl_0
  );


  buf

  (
    ffc_478_n_spl_000,
    ffc_478_n_spl_00
  );


  buf

  (
    ffc_478_n_spl_001,
    ffc_478_n_spl_00
  );


  buf

  (
    ffc_478_n_spl_01,
    ffc_478_n_spl_0
  );


  buf

  (
    ffc_478_n_spl_1,
    ffc_478_n_spl_
  );


  buf

  (
    ffc_478_n_spl_10,
    ffc_478_n_spl_1
  );


  buf

  (
    ffc_478_n_spl_11,
    ffc_478_n_spl_1
  );


  buf

  (
    ffc_523_n_spl_,
    ffc_523_n
  );


  buf

  (
    ffc_744_n_spl_,
    ffc_744_n
  );


  buf

  (
    g1159_n_spl_,
    g1159_n
  );


  buf

  (
    ffc_486_n_spl_,
    ffc_486_n
  );


  buf

  (
    ffc_486_n_spl_0,
    ffc_486_n_spl_
  );


  buf

  (
    ffc_486_n_spl_00,
    ffc_486_n_spl_0
  );


  buf

  (
    ffc_486_n_spl_000,
    ffc_486_n_spl_00
  );


  buf

  (
    ffc_486_n_spl_0000,
    ffc_486_n_spl_000
  );


  buf

  (
    ffc_486_n_spl_0001,
    ffc_486_n_spl_000
  );


  buf

  (
    ffc_486_n_spl_001,
    ffc_486_n_spl_00
  );


  buf

  (
    ffc_486_n_spl_0010,
    ffc_486_n_spl_001
  );


  buf

  (
    ffc_486_n_spl_0011,
    ffc_486_n_spl_001
  );


  buf

  (
    ffc_486_n_spl_01,
    ffc_486_n_spl_0
  );


  buf

  (
    ffc_486_n_spl_010,
    ffc_486_n_spl_01
  );


  buf

  (
    ffc_486_n_spl_011,
    ffc_486_n_spl_01
  );


  buf

  (
    ffc_486_n_spl_1,
    ffc_486_n_spl_
  );


  buf

  (
    ffc_486_n_spl_10,
    ffc_486_n_spl_1
  );


  buf

  (
    ffc_486_n_spl_100,
    ffc_486_n_spl_10
  );


  buf

  (
    ffc_486_n_spl_101,
    ffc_486_n_spl_10
  );


  buf

  (
    ffc_486_n_spl_11,
    ffc_486_n_spl_1
  );


  buf

  (
    ffc_486_n_spl_110,
    ffc_486_n_spl_11
  );


  buf

  (
    ffc_486_n_spl_111,
    ffc_486_n_spl_11
  );


  buf

  (
    ffc_486_p_spl_,
    ffc_486_p
  );


  buf

  (
    ffc_486_p_spl_0,
    ffc_486_p_spl_
  );


  buf

  (
    ffc_486_p_spl_00,
    ffc_486_p_spl_0
  );


  buf

  (
    ffc_486_p_spl_000,
    ffc_486_p_spl_00
  );


  buf

  (
    ffc_486_p_spl_0000,
    ffc_486_p_spl_000
  );


  buf

  (
    ffc_486_p_spl_0001,
    ffc_486_p_spl_000
  );


  buf

  (
    ffc_486_p_spl_001,
    ffc_486_p_spl_00
  );


  buf

  (
    ffc_486_p_spl_0010,
    ffc_486_p_spl_001
  );


  buf

  (
    ffc_486_p_spl_0011,
    ffc_486_p_spl_001
  );


  buf

  (
    ffc_486_p_spl_01,
    ffc_486_p_spl_0
  );


  buf

  (
    ffc_486_p_spl_010,
    ffc_486_p_spl_01
  );


  buf

  (
    ffc_486_p_spl_011,
    ffc_486_p_spl_01
  );


  buf

  (
    ffc_486_p_spl_1,
    ffc_486_p_spl_
  );


  buf

  (
    ffc_486_p_spl_10,
    ffc_486_p_spl_1
  );


  buf

  (
    ffc_486_p_spl_100,
    ffc_486_p_spl_10
  );


  buf

  (
    ffc_486_p_spl_101,
    ffc_486_p_spl_10
  );


  buf

  (
    ffc_486_p_spl_11,
    ffc_486_p_spl_1
  );


  buf

  (
    ffc_486_p_spl_110,
    ffc_486_p_spl_11
  );


  buf

  (
    ffc_486_p_spl_111,
    ffc_486_p_spl_11
  );


  buf

  (
    ffc_490_p_spl_,
    ffc_490_p
  );


  buf

  (
    ffc_490_p_spl_0,
    ffc_490_p_spl_
  );


  buf

  (
    ffc_490_p_spl_00,
    ffc_490_p_spl_0
  );


  buf

  (
    ffc_490_p_spl_000,
    ffc_490_p_spl_00
  );


  buf

  (
    ffc_490_p_spl_001,
    ffc_490_p_spl_00
  );


  buf

  (
    ffc_490_p_spl_01,
    ffc_490_p_spl_0
  );


  buf

  (
    ffc_490_p_spl_1,
    ffc_490_p_spl_
  );


  buf

  (
    ffc_490_p_spl_10,
    ffc_490_p_spl_1
  );


  buf

  (
    ffc_490_p_spl_11,
    ffc_490_p_spl_1
  );


  buf

  (
    ffc_490_n_spl_,
    ffc_490_n
  );


  buf

  (
    ffc_490_n_spl_0,
    ffc_490_n_spl_
  );


  buf

  (
    ffc_490_n_spl_00,
    ffc_490_n_spl_0
  );


  buf

  (
    ffc_490_n_spl_000,
    ffc_490_n_spl_00
  );


  buf

  (
    ffc_490_n_spl_001,
    ffc_490_n_spl_00
  );


  buf

  (
    ffc_490_n_spl_01,
    ffc_490_n_spl_0
  );


  buf

  (
    ffc_490_n_spl_1,
    ffc_490_n_spl_
  );


  buf

  (
    ffc_490_n_spl_10,
    ffc_490_n_spl_1
  );


  buf

  (
    ffc_490_n_spl_11,
    ffc_490_n_spl_1
  );


  buf

  (
    g1176_n_spl_,
    g1176_n
  );


  buf

  (
    g1183_n_spl_,
    g1183_n
  );


  buf

  (
    g1188_n_spl_,
    g1188_n
  );


  buf

  (
    ffc_561_n_spl_,
    ffc_561_n
  );


  buf

  (
    ffc_561_n_spl_0,
    ffc_561_n_spl_
  );


  buf

  (
    ffc_561_n_spl_00,
    ffc_561_n_spl_0
  );


  buf

  (
    ffc_561_n_spl_1,
    ffc_561_n_spl_
  );


  buf

  (
    g1201_n_spl_,
    g1201_n
  );


  buf

  (
    ffc_561_p_spl_,
    ffc_561_p
  );


  buf

  (
    ffc_561_p_spl_0,
    ffc_561_p_spl_
  );


  buf

  (
    ffc_561_p_spl_1,
    ffc_561_p_spl_
  );


  buf

  (
    g1201_p_spl_,
    g1201_p
  );


  buf

  (
    g1205_p_spl_,
    g1205_p
  );


  buf

  (
    g1206_n_spl_,
    g1206_n
  );


  buf

  (
    g1205_n_spl_,
    g1205_n
  );


  buf

  (
    g1206_p_spl_,
    g1206_p
  );


  buf

  (
    ffc_504_n_spl_,
    ffc_504_n
  );


  buf

  (
    ffc_505_p_spl_,
    ffc_505_p
  );


  buf

  (
    ffc_504_p_spl_,
    ffc_504_p
  );


  buf

  (
    ffc_505_n_spl_,
    ffc_505_n
  );


  buf

  (
    ffc_507_n_spl_,
    ffc_507_n
  );


  buf

  (
    ffc_511_p_spl_,
    ffc_511_p
  );


  buf

  (
    ffc_507_p_spl_,
    ffc_507_p
  );


  buf

  (
    ffc_511_n_spl_,
    ffc_511_n
  );


  buf

  (
    g1215_n_spl_,
    g1215_n
  );


  buf

  (
    g1218_p_spl_,
    g1218_p
  );


  buf

  (
    g1215_p_spl_,
    g1215_p
  );


  buf

  (
    g1218_n_spl_,
    g1218_n
  );


  buf

  (
    ffc_739_n_spl_,
    ffc_739_n
  );


  buf

  (
    ffc_742_p_spl_,
    ffc_742_p
  );


  buf

  (
    ffc_739_p_spl_,
    ffc_739_p
  );


  buf

  (
    ffc_742_n_spl_,
    ffc_742_n
  );


  buf

  (
    ffc_503_p_spl_,
    ffc_503_p
  );


  buf

  (
    ffc_506_n_spl_,
    ffc_506_n
  );


  buf

  (
    ffc_503_n_spl_,
    ffc_503_n
  );


  buf

  (
    ffc_506_p_spl_,
    ffc_506_p
  );


  buf

  (
    g1224_n_spl_,
    g1224_n
  );


  buf

  (
    g1227_p_spl_,
    g1227_p
  );


  buf

  (
    g1224_p_spl_,
    g1224_p
  );


  buf

  (
    g1227_n_spl_,
    g1227_n
  );


  buf

  (
    g1234_n_spl_,
    g1234_n
  );


  buf

  (
    ffc_745_n_spl_,
    ffc_745_n
  );


  buf

  (
    g1243_p_spl_,
    g1243_p
  );


  buf

  (
    g1246_p_spl_,
    g1246_p
  );


  buf

  (
    ffc_746_p_spl_,
    ffc_746_p
  );


  buf

  (
    g1250_p_spl_,
    g1250_p
  );


  buf

  (
    g1249_p_spl_,
    g1249_p
  );


  buf

  (
    ffc_428_n_spl_,
    ffc_428_n
  );


  buf

  (
    ffc_428_n_spl_0,
    ffc_428_n_spl_
  );


  buf

  (
    ffc_428_n_spl_00,
    ffc_428_n_spl_0
  );


  buf

  (
    ffc_428_n_spl_000,
    ffc_428_n_spl_00
  );


  buf

  (
    ffc_428_n_spl_0000,
    ffc_428_n_spl_000
  );


  buf

  (
    ffc_428_n_spl_0001,
    ffc_428_n_spl_000
  );


  buf

  (
    ffc_428_n_spl_001,
    ffc_428_n_spl_00
  );


  buf

  (
    ffc_428_n_spl_0010,
    ffc_428_n_spl_001
  );


  buf

  (
    ffc_428_n_spl_0011,
    ffc_428_n_spl_001
  );


  buf

  (
    ffc_428_n_spl_01,
    ffc_428_n_spl_0
  );


  buf

  (
    ffc_428_n_spl_010,
    ffc_428_n_spl_01
  );


  buf

  (
    ffc_428_n_spl_011,
    ffc_428_n_spl_01
  );


  buf

  (
    ffc_428_n_spl_1,
    ffc_428_n_spl_
  );


  buf

  (
    ffc_428_n_spl_10,
    ffc_428_n_spl_1
  );


  buf

  (
    ffc_428_n_spl_100,
    ffc_428_n_spl_10
  );


  buf

  (
    ffc_428_n_spl_101,
    ffc_428_n_spl_10
  );


  buf

  (
    ffc_428_n_spl_11,
    ffc_428_n_spl_1
  );


  buf

  (
    ffc_428_n_spl_110,
    ffc_428_n_spl_11
  );


  buf

  (
    ffc_428_n_spl_111,
    ffc_428_n_spl_11
  );


  buf

  (
    ffc_428_p_spl_,
    ffc_428_p
  );


  buf

  (
    ffc_428_p_spl_0,
    ffc_428_p_spl_
  );


  buf

  (
    ffc_428_p_spl_00,
    ffc_428_p_spl_0
  );


  buf

  (
    ffc_428_p_spl_000,
    ffc_428_p_spl_00
  );


  buf

  (
    ffc_428_p_spl_0000,
    ffc_428_p_spl_000
  );


  buf

  (
    ffc_428_p_spl_0001,
    ffc_428_p_spl_000
  );


  buf

  (
    ffc_428_p_spl_001,
    ffc_428_p_spl_00
  );


  buf

  (
    ffc_428_p_spl_0010,
    ffc_428_p_spl_001
  );


  buf

  (
    ffc_428_p_spl_0011,
    ffc_428_p_spl_001
  );


  buf

  (
    ffc_428_p_spl_01,
    ffc_428_p_spl_0
  );


  buf

  (
    ffc_428_p_spl_010,
    ffc_428_p_spl_01
  );


  buf

  (
    ffc_428_p_spl_011,
    ffc_428_p_spl_01
  );


  buf

  (
    ffc_428_p_spl_1,
    ffc_428_p_spl_
  );


  buf

  (
    ffc_428_p_spl_10,
    ffc_428_p_spl_1
  );


  buf

  (
    ffc_428_p_spl_100,
    ffc_428_p_spl_10
  );


  buf

  (
    ffc_428_p_spl_101,
    ffc_428_p_spl_10
  );


  buf

  (
    ffc_428_p_spl_11,
    ffc_428_p_spl_1
  );


  buf

  (
    ffc_428_p_spl_110,
    ffc_428_p_spl_11
  );


  buf

  (
    ffc_428_p_spl_111,
    ffc_428_p_spl_11
  );


  buf

  (
    ffc_432_n_spl_,
    ffc_432_n
  );


  buf

  (
    ffc_432_n_spl_0,
    ffc_432_n_spl_
  );


  buf

  (
    ffc_432_n_spl_00,
    ffc_432_n_spl_0
  );


  buf

  (
    ffc_432_n_spl_000,
    ffc_432_n_spl_00
  );


  buf

  (
    ffc_432_n_spl_001,
    ffc_432_n_spl_00
  );


  buf

  (
    ffc_432_n_spl_01,
    ffc_432_n_spl_0
  );


  buf

  (
    ffc_432_n_spl_1,
    ffc_432_n_spl_
  );


  buf

  (
    ffc_432_n_spl_10,
    ffc_432_n_spl_1
  );


  buf

  (
    ffc_432_n_spl_11,
    ffc_432_n_spl_1
  );


  buf

  (
    ffc_309_p_spl_,
    ffc_309_p
  );


  buf

  (
    ffc_305_p_spl_,
    ffc_305_p
  );


  buf

  (
    ffc_432_p_spl_,
    ffc_432_p
  );


  buf

  (
    ffc_432_p_spl_0,
    ffc_432_p_spl_
  );


  buf

  (
    ffc_432_p_spl_00,
    ffc_432_p_spl_0
  );


  buf

  (
    ffc_432_p_spl_000,
    ffc_432_p_spl_00
  );


  buf

  (
    ffc_432_p_spl_001,
    ffc_432_p_spl_00
  );


  buf

  (
    ffc_432_p_spl_01,
    ffc_432_p_spl_0
  );


  buf

  (
    ffc_432_p_spl_1,
    ffc_432_p_spl_
  );


  buf

  (
    ffc_432_p_spl_10,
    ffc_432_p_spl_1
  );


  buf

  (
    ffc_432_p_spl_11,
    ffc_432_p_spl_1
  );


  buf

  (
    ffc_241_p_spl_,
    ffc_241_p
  );


  buf

  (
    ffc_241_p_spl_0,
    ffc_241_p_spl_
  );


  buf

  (
    ffc_241_p_spl_00,
    ffc_241_p_spl_0
  );


  buf

  (
    ffc_241_p_spl_000,
    ffc_241_p_spl_00
  );


  buf

  (
    ffc_241_p_spl_0000,
    ffc_241_p_spl_000
  );


  buf

  (
    ffc_241_p_spl_001,
    ffc_241_p_spl_00
  );


  buf

  (
    ffc_241_p_spl_01,
    ffc_241_p_spl_0
  );


  buf

  (
    ffc_241_p_spl_010,
    ffc_241_p_spl_01
  );


  buf

  (
    ffc_241_p_spl_011,
    ffc_241_p_spl_01
  );


  buf

  (
    ffc_241_p_spl_1,
    ffc_241_p_spl_
  );


  buf

  (
    ffc_241_p_spl_10,
    ffc_241_p_spl_1
  );


  buf

  (
    ffc_241_p_spl_100,
    ffc_241_p_spl_10
  );


  buf

  (
    ffc_241_p_spl_101,
    ffc_241_p_spl_10
  );


  buf

  (
    ffc_241_p_spl_11,
    ffc_241_p_spl_1
  );


  buf

  (
    ffc_241_p_spl_110,
    ffc_241_p_spl_11
  );


  buf

  (
    ffc_241_p_spl_111,
    ffc_241_p_spl_11
  );


  buf

  (
    ffc_436_n_spl_,
    ffc_436_n
  );


  buf

  (
    ffc_436_n_spl_0,
    ffc_436_n_spl_
  );


  buf

  (
    ffc_436_n_spl_00,
    ffc_436_n_spl_0
  );


  buf

  (
    ffc_436_n_spl_000,
    ffc_436_n_spl_00
  );


  buf

  (
    ffc_436_n_spl_0000,
    ffc_436_n_spl_000
  );


  buf

  (
    ffc_436_n_spl_0001,
    ffc_436_n_spl_000
  );


  buf

  (
    ffc_436_n_spl_001,
    ffc_436_n_spl_00
  );


  buf

  (
    ffc_436_n_spl_0010,
    ffc_436_n_spl_001
  );


  buf

  (
    ffc_436_n_spl_0011,
    ffc_436_n_spl_001
  );


  buf

  (
    ffc_436_n_spl_01,
    ffc_436_n_spl_0
  );


  buf

  (
    ffc_436_n_spl_010,
    ffc_436_n_spl_01
  );


  buf

  (
    ffc_436_n_spl_011,
    ffc_436_n_spl_01
  );


  buf

  (
    ffc_436_n_spl_1,
    ffc_436_n_spl_
  );


  buf

  (
    ffc_436_n_spl_10,
    ffc_436_n_spl_1
  );


  buf

  (
    ffc_436_n_spl_100,
    ffc_436_n_spl_10
  );


  buf

  (
    ffc_436_n_spl_101,
    ffc_436_n_spl_10
  );


  buf

  (
    ffc_436_n_spl_11,
    ffc_436_n_spl_1
  );


  buf

  (
    ffc_436_n_spl_110,
    ffc_436_n_spl_11
  );


  buf

  (
    ffc_436_n_spl_111,
    ffc_436_n_spl_11
  );


  buf

  (
    ffc_436_p_spl_,
    ffc_436_p
  );


  buf

  (
    ffc_436_p_spl_0,
    ffc_436_p_spl_
  );


  buf

  (
    ffc_436_p_spl_00,
    ffc_436_p_spl_0
  );


  buf

  (
    ffc_436_p_spl_000,
    ffc_436_p_spl_00
  );


  buf

  (
    ffc_436_p_spl_0000,
    ffc_436_p_spl_000
  );


  buf

  (
    ffc_436_p_spl_0001,
    ffc_436_p_spl_000
  );


  buf

  (
    ffc_436_p_spl_001,
    ffc_436_p_spl_00
  );


  buf

  (
    ffc_436_p_spl_0010,
    ffc_436_p_spl_001
  );


  buf

  (
    ffc_436_p_spl_0011,
    ffc_436_p_spl_001
  );


  buf

  (
    ffc_436_p_spl_01,
    ffc_436_p_spl_0
  );


  buf

  (
    ffc_436_p_spl_010,
    ffc_436_p_spl_01
  );


  buf

  (
    ffc_436_p_spl_011,
    ffc_436_p_spl_01
  );


  buf

  (
    ffc_436_p_spl_1,
    ffc_436_p_spl_
  );


  buf

  (
    ffc_436_p_spl_10,
    ffc_436_p_spl_1
  );


  buf

  (
    ffc_436_p_spl_100,
    ffc_436_p_spl_10
  );


  buf

  (
    ffc_436_p_spl_101,
    ffc_436_p_spl_10
  );


  buf

  (
    ffc_436_p_spl_11,
    ffc_436_p_spl_1
  );


  buf

  (
    ffc_436_p_spl_110,
    ffc_436_p_spl_11
  );


  buf

  (
    ffc_436_p_spl_111,
    ffc_436_p_spl_11
  );


  buf

  (
    ffc_440_n_spl_,
    ffc_440_n
  );


  buf

  (
    ffc_440_n_spl_0,
    ffc_440_n_spl_
  );


  buf

  (
    ffc_440_n_spl_00,
    ffc_440_n_spl_0
  );


  buf

  (
    ffc_440_n_spl_000,
    ffc_440_n_spl_00
  );


  buf

  (
    ffc_440_n_spl_001,
    ffc_440_n_spl_00
  );


  buf

  (
    ffc_440_n_spl_01,
    ffc_440_n_spl_0
  );


  buf

  (
    ffc_440_n_spl_1,
    ffc_440_n_spl_
  );


  buf

  (
    ffc_440_n_spl_10,
    ffc_440_n_spl_1
  );


  buf

  (
    ffc_440_n_spl_11,
    ffc_440_n_spl_1
  );


  buf

  (
    ffc_440_p_spl_,
    ffc_440_p
  );


  buf

  (
    ffc_440_p_spl_0,
    ffc_440_p_spl_
  );


  buf

  (
    ffc_440_p_spl_00,
    ffc_440_p_spl_0
  );


  buf

  (
    ffc_440_p_spl_000,
    ffc_440_p_spl_00
  );


  buf

  (
    ffc_440_p_spl_001,
    ffc_440_p_spl_00
  );


  buf

  (
    ffc_440_p_spl_01,
    ffc_440_p_spl_0
  );


  buf

  (
    ffc_440_p_spl_1,
    ffc_440_p_spl_
  );


  buf

  (
    ffc_440_p_spl_10,
    ffc_440_p_spl_1
  );


  buf

  (
    ffc_440_p_spl_11,
    ffc_440_p_spl_1
  );


  buf

  (
    ffc_54_p_spl_,
    ffc_54_p
  );


  buf

  (
    ffc_62_p_spl_,
    ffc_62_p
  );


  buf

  (
    g1182_n_spl_,
    g1182_n
  );


  buf

  (
    g1182_n_spl_0,
    g1182_n_spl_
  );


  buf

  (
    g1182_n_spl_00,
    g1182_n_spl_0
  );


  buf

  (
    g1182_n_spl_1,
    g1182_n_spl_
  );


  buf

  (
    g1155_n_spl_,
    g1155_n
  );


  buf

  (
    g1155_n_spl_0,
    g1155_n_spl_
  );


  buf

  (
    g1155_n_spl_00,
    g1155_n_spl_0
  );


  buf

  (
    g1155_n_spl_1,
    g1155_n_spl_
  );


  buf

  (
    ffc_22_p_spl_,
    ffc_22_p
  );


  buf

  (
    ffc_104_p_spl_,
    ffc_104_p
  );


  buf

  (
    g1187_n_spl_,
    g1187_n
  );


  buf

  (
    g1187_n_spl_0,
    g1187_n_spl_
  );


  buf

  (
    g1187_n_spl_00,
    g1187_n_spl_0
  );


  buf

  (
    g1187_n_spl_1,
    g1187_n_spl_
  );


  buf

  (
    g1158_n_spl_,
    g1158_n
  );


  buf

  (
    g1158_n_spl_0,
    g1158_n_spl_
  );


  buf

  (
    g1158_n_spl_00,
    g1158_n_spl_0
  );


  buf

  (
    g1158_n_spl_1,
    g1158_n_spl_
  );


  buf

  (
    ffc_18_p_spl_,
    ffc_18_p
  );


  buf

  (
    ffc_100_p_spl_,
    ffc_100_p
  );


  buf

  (
    g1194_n_spl_,
    g1194_n
  );


  buf

  (
    g1194_n_spl_0,
    g1194_n_spl_
  );


  buf

  (
    g1194_n_spl_00,
    g1194_n_spl_0
  );


  buf

  (
    g1194_n_spl_1,
    g1194_n_spl_
  );


  buf

  (
    g1164_n_spl_,
    g1164_n
  );


  buf

  (
    g1164_n_spl_0,
    g1164_n_spl_
  );


  buf

  (
    g1164_n_spl_00,
    g1164_n_spl_0
  );


  buf

  (
    g1164_n_spl_1,
    g1164_n_spl_
  );


  buf

  (
    ffc_96_n_spl_,
    ffc_96_n
  );


  buf

  (
    ffc_92_n_spl_,
    ffc_92_n
  );


  buf

  (
    g1200_p_spl_,
    g1200_p
  );


  buf

  (
    g1200_p_spl_0,
    g1200_p_spl_
  );


  buf

  (
    g1200_p_spl_00,
    g1200_p_spl_0
  );


  buf

  (
    g1200_p_spl_1,
    g1200_p_spl_
  );


  buf

  (
    g1137_p_spl_,
    g1137_p
  );


  buf

  (
    g1137_p_spl_0,
    g1137_p_spl_
  );


  buf

  (
    g1137_p_spl_00,
    g1137_p_spl_0
  );


  buf

  (
    g1137_p_spl_1,
    g1137_p_spl_
  );


  buf

  (
    ffc_289_p_spl_,
    ffc_289_p
  );


  buf

  (
    ffc_329_p_spl_,
    ffc_329_p
  );


  buf

  (
    ffc_273_n_spl_,
    ffc_273_n
  );


  buf

  (
    ffc_313_n_spl_,
    ffc_313_n
  );


  buf

  (
    ffc_241_n_spl_,
    ffc_241_n
  );


  buf

  (
    ffc_241_n_spl_0,
    ffc_241_n_spl_
  );


  buf

  (
    ffc_241_n_spl_1,
    ffc_241_n_spl_
  );


  buf

  (
    ffc_265_p_spl_,
    ffc_265_p
  );


  buf

  (
    ffc_269_p_spl_,
    ffc_269_p
  );


  buf

  (
    ffc_257_p_spl_,
    ffc_257_p
  );


  buf

  (
    ffc_261_p_spl_,
    ffc_261_p
  );


  buf

  (
    ffc_474_n_spl_,
    ffc_474_n
  );


  buf

  (
    ffc_474_p_spl_,
    ffc_474_p
  );


  buf

  (
    ffc_229_n_spl_,
    ffc_229_n
  );


  buf

  (
    ffc_229_p_spl_,
    ffc_229_p
  );


  buf

  (
    ffc_532_n_spl_,
    ffc_532_n
  );


  buf

  (
    g1437_n_spl_,
    g1437_n
  );


  buf

  (
    ffc_342_n_spl_,
    ffc_342_n
  );


  buf

  (
    ffc_417_n_spl_,
    ffc_417_n
  );


  buf

  (
    g1049_n_spl_,
    g1049_n
  );


  buf

  (
    g1054_n_spl_,
    g1054_n
  );


  buf

  (
    g1111_n_spl_,
    g1111_n
  );


  buf

  (
    g1120_n_spl_,
    g1120_n
  );


  buf

  (
    g1212_n_spl_,
    g1212_n
  );


  buf

  (
    g1233_n_spl_,
    g1233_n
  );


  buf

  (
    ffc_160_p_spl_,
    ffc_160_p
  );


  buf

  (
    ffc_164_p_spl_,
    ffc_164_p
  );


  buf

  (
    g1470_n_spl_,
    g1470_n
  );


  buf

  (
    g1470_n_spl_0,
    g1470_n_spl_
  );


  buf

  (
    g1470_n_spl_00,
    g1470_n_spl_0
  );


  buf

  (
    g1470_n_spl_1,
    g1470_n_spl_
  );


  buf

  (
    g1449_n_spl_,
    g1449_n
  );


  buf

  (
    g1449_n_spl_0,
    g1449_n_spl_
  );


  buf

  (
    g1449_n_spl_00,
    g1449_n_spl_0
  );


  buf

  (
    g1449_n_spl_1,
    g1449_n_spl_
  );


  buf

  (
    ffc_70_p_spl_,
    ffc_70_p
  );


  buf

  (
    ffc_66_p_spl_,
    ffc_66_p
  );


  buf

  (
    g1476_n_spl_,
    g1476_n
  );


  buf

  (
    g1476_n_spl_0,
    g1476_n_spl_
  );


  buf

  (
    g1476_n_spl_00,
    g1476_n_spl_0
  );


  buf

  (
    g1476_n_spl_1,
    g1476_n_spl_
  );


  buf

  (
    g1453_n_spl_,
    g1453_n
  );


  buf

  (
    g1453_n_spl_0,
    g1453_n_spl_
  );


  buf

  (
    g1453_n_spl_00,
    g1453_n_spl_0
  );


  buf

  (
    g1453_n_spl_1,
    g1453_n_spl_
  );


  buf

  (
    ffc_156_p_spl_,
    ffc_156_p
  );


  buf

  (
    ffc_152_p_spl_,
    ffc_152_p
  );


  buf

  (
    g1482_n_spl_,
    g1482_n
  );


  buf

  (
    g1482_n_spl_0,
    g1482_n_spl_
  );


  buf

  (
    g1482_n_spl_00,
    g1482_n_spl_0
  );


  buf

  (
    g1482_n_spl_1,
    g1482_n_spl_
  );


  buf

  (
    g1457_n_spl_,
    g1457_n
  );


  buf

  (
    g1457_n_spl_0,
    g1457_n_spl_
  );


  buf

  (
    g1457_n_spl_00,
    g1457_n_spl_0
  );


  buf

  (
    g1457_n_spl_1,
    g1457_n_spl_
  );


  buf

  (
    ffc_58_p_spl_,
    ffc_58_p
  );


  buf

  (
    ffc_140_p_spl_,
    ffc_140_p
  );


  buf

  (
    g1486_n_spl_,
    g1486_n
  );


  buf

  (
    g1486_n_spl_0,
    g1486_n_spl_
  );


  buf

  (
    g1486_n_spl_00,
    g1486_n_spl_0
  );


  buf

  (
    g1486_n_spl_1,
    g1486_n_spl_
  );


  buf

  (
    g1460_n_spl_,
    g1460_n
  );


  buf

  (
    g1460_n_spl_0,
    g1460_n_spl_
  );


  buf

  (
    g1460_n_spl_00,
    g1460_n_spl_0
  );


  buf

  (
    g1460_n_spl_1,
    g1460_n_spl_
  );


  buf

  (
    ffc_293_p_spl_,
    ffc_293_p
  );


  buf

  (
    ffc_333_p_spl_,
    ffc_333_p
  );


  buf

  (
    ffc_285_p_spl_,
    ffc_285_p
  );


  buf

  (
    ffc_325_p_spl_,
    ffc_325_p
  );


  buf

  (
    ffc_281_p_spl_,
    ffc_281_p
  );


  buf

  (
    ffc_321_p_spl_,
    ffc_321_p
  );


  buf

  (
    ffc_277_p_spl_,
    ffc_277_p
  );


  buf

  (
    ffc_317_p_spl_,
    ffc_317_p
  );


  buf

  (
    g1640_n_spl_,
    g1640_n
  );


  buf

  (
    g1639_n_spl_,
    g1639_n
  );


  buf

  (
    g1645_n_spl_,
    g1645_n
  );


  buf

  (
    ffc_88_n_spl_,
    ffc_88_n
  );


  buf

  (
    ffc_14_n_spl_,
    ffc_14_n
  );


  buf

  (
    g1653_p_spl_,
    g1653_p
  );


  buf

  (
    g1653_p_spl_0,
    g1653_p_spl_
  );


  buf

  (
    g1653_p_spl_1,
    g1653_p_spl_
  );


  buf

  (
    g1656_p_spl_,
    g1656_p
  );


  buf

  (
    g1656_p_spl_0,
    g1656_p_spl_
  );


  buf

  (
    g1656_p_spl_1,
    g1656_p_spl_
  );


  buf

  (
    ffc_301_n_spl_,
    ffc_301_n
  );


  buf

  (
    ffc_297_n_spl_,
    ffc_297_n
  );


  buf

  (
    ffc_610_n_spl_,
    ffc_610_n
  );


  buf

  (
    ffc_610_n_spl_0,
    ffc_610_n_spl_
  );


  buf

  (
    ffc_610_n_spl_1,
    ffc_610_n_spl_
  );


  buf

  (
    ffc_783_n_spl_,
    ffc_783_n
  );


  buf

  (
    ffc_610_p_spl_,
    ffc_610_p
  );


  buf

  (
    ffc_610_p_spl_0,
    ffc_610_p_spl_
  );


  buf

  (
    ffc_783_p_spl_,
    ffc_783_p
  );


  buf

  (
    ffc_783_p_spl_0,
    ffc_783_p_spl_
  );


  buf

  (
    g1690_n_spl_,
    g1690_n
  );


  buf

  (
    ffc_578_n_spl_,
    ffc_578_n
  );


  buf

  (
    ffc_578_n_spl_0,
    ffc_578_n_spl_
  );


  buf

  (
    ffc_578_n_spl_00,
    ffc_578_n_spl_0
  );


  buf

  (
    ffc_578_n_spl_1,
    ffc_578_n_spl_
  );


  buf

  (
    ffc_624_n_spl_,
    ffc_624_n
  );


  buf

  (
    ffc_6_p_spl_,
    ffc_6_p
  );


  buf

  (
    ffc_6_p_spl_0,
    ffc_6_p_spl_
  );


  buf

  (
    ffc_6_p_spl_1,
    ffc_6_p_spl_
  );


  buf

  (
    ffc_587_p_spl_,
    ffc_587_p
  );


  buf

  (
    g1695_n_spl_,
    g1695_n
  );


  buf

  (
    ffc_842_n_spl_,
    ffc_842_n
  );


  buf

  (
    ffc_842_p_spl_,
    ffc_842_p
  );


  buf

  (
    ffc_842_p_spl_0,
    ffc_842_p_spl_
  );


  buf

  (
    ffc_827_n_spl_,
    ffc_827_n
  );


  buf

  (
    ffc_827_p_spl_,
    ffc_827_p
  );


  buf

  (
    ffc_840_p_spl_,
    ffc_840_p
  );


  buf

  (
    ffc_843_p_spl_,
    ffc_843_p
  );


  buf

  (
    ffc_843_p_spl_0,
    ffc_843_p_spl_
  );


  buf

  (
    ffc_845_p_spl_,
    ffc_845_p
  );


  buf

  (
    ffc_843_n_spl_,
    ffc_843_n
  );


  buf

  (
    ffc_770_p_spl_,
    ffc_770_p
  );


  buf

  (
    ffc_770_p_spl_0,
    ffc_770_p_spl_
  );


  buf

  (
    g1703_p_spl_,
    g1703_p
  );


  buf

  (
    g1703_p_spl_0,
    g1703_p_spl_
  );


  buf

  (
    ffc_770_n_spl_,
    ffc_770_n
  );


  buf

  (
    g1703_n_spl_,
    g1703_n
  );


  buf

  (
    ffc_466_n_spl_,
    ffc_466_n
  );


  buf

  (
    ffc_466_n_spl_0,
    ffc_466_n_spl_
  );


  buf

  (
    ffc_466_n_spl_00,
    ffc_466_n_spl_0
  );


  buf

  (
    ffc_466_n_spl_000,
    ffc_466_n_spl_00
  );


  buf

  (
    ffc_466_n_spl_001,
    ffc_466_n_spl_00
  );


  buf

  (
    ffc_466_n_spl_01,
    ffc_466_n_spl_0
  );


  buf

  (
    ffc_466_n_spl_010,
    ffc_466_n_spl_01
  );


  buf

  (
    ffc_466_n_spl_011,
    ffc_466_n_spl_01
  );


  buf

  (
    ffc_466_n_spl_1,
    ffc_466_n_spl_
  );


  buf

  (
    ffc_466_n_spl_10,
    ffc_466_n_spl_1
  );


  buf

  (
    ffc_466_n_spl_11,
    ffc_466_n_spl_1
  );


  buf

  (
    ffc_457_p_spl_,
    ffc_457_p
  );


  buf

  (
    ffc_457_p_spl_0,
    ffc_457_p_spl_
  );


  buf

  (
    ffc_457_p_spl_00,
    ffc_457_p_spl_0
  );


  buf

  (
    ffc_457_p_spl_000,
    ffc_457_p_spl_00
  );


  buf

  (
    ffc_457_p_spl_001,
    ffc_457_p_spl_00
  );


  buf

  (
    ffc_457_p_spl_01,
    ffc_457_p_spl_0
  );


  buf

  (
    ffc_457_p_spl_010,
    ffc_457_p_spl_01
  );


  buf

  (
    ffc_457_p_spl_011,
    ffc_457_p_spl_01
  );


  buf

  (
    ffc_457_p_spl_1,
    ffc_457_p_spl_
  );


  buf

  (
    ffc_457_p_spl_10,
    ffc_457_p_spl_1
  );


  buf

  (
    ffc_457_p_spl_11,
    ffc_457_p_spl_1
  );


  buf

  (
    ffc_623_p_spl_,
    ffc_623_p
  );


  buf

  (
    ffc_623_p_spl_0,
    ffc_623_p_spl_
  );


  buf

  (
    ffc_829_p_spl_,
    ffc_829_p
  );


  buf

  (
    ffc_829_p_spl_0,
    ffc_829_p_spl_
  );


  buf

  (
    ffc_829_p_spl_00,
    ffc_829_p_spl_0
  );


  buf

  (
    ffc_829_p_spl_01,
    ffc_829_p_spl_0
  );


  buf

  (
    ffc_829_p_spl_1,
    ffc_829_p_spl_
  );


  buf

  (
    ffc_623_n_spl_,
    ffc_623_n
  );


  buf

  (
    ffc_829_n_spl_,
    ffc_829_n
  );


  buf

  (
    ffc_829_n_spl_0,
    ffc_829_n_spl_
  );


  buf

  (
    ffc_829_n_spl_00,
    ffc_829_n_spl_0
  );


  buf

  (
    ffc_829_n_spl_1,
    ffc_829_n_spl_
  );


  buf

  (
    ffc_775_p_spl_,
    ffc_775_p
  );


  buf

  (
    ffc_683_p_spl_,
    ffc_683_p
  );


  buf

  (
    g1698_n_spl_,
    g1698_n
  );


  buf

  (
    g1698_n_spl_0,
    g1698_n_spl_
  );


  buf

  (
    g1698_n_spl_1,
    g1698_n_spl_
  );


  buf

  (
    g1698_p_spl_,
    g1698_p
  );


  buf

  (
    g1698_p_spl_0,
    g1698_p_spl_
  );


  buf

  (
    ffc_813_n_spl_,
    ffc_813_n
  );


  buf

  (
    ffc_813_p_spl_,
    ffc_813_p
  );


  buf

  (
    ffc_795_p_spl_,
    ffc_795_p
  );


  buf

  (
    ffc_795_p_spl_0,
    ffc_795_p_spl_
  );


  buf

  (
    ffc_795_p_spl_1,
    ffc_795_p_spl_
  );


  buf

  (
    ffc_815_n_spl_,
    ffc_815_n
  );


  buf

  (
    ffc_795_n_spl_,
    ffc_795_n
  );


  buf

  (
    ffc_795_n_spl_0,
    ffc_795_n_spl_
  );


  buf

  (
    ffc_815_p_spl_,
    ffc_815_p
  );


  buf

  (
    ffc_816_p_spl_,
    ffc_816_p
  );


  buf

  (
    ffc_816_p_spl_0,
    ffc_816_p_spl_
  );


  buf

  (
    ffc_816_p_spl_00,
    ffc_816_p_spl_0
  );


  buf

  (
    ffc_816_p_spl_1,
    ffc_816_p_spl_
  );


  buf

  (
    g1700_n_spl_,
    g1700_n
  );


  buf

  (
    g1700_n_spl_0,
    g1700_n_spl_
  );


  buf

  (
    ffc_816_n_spl_,
    ffc_816_n
  );


  buf

  (
    ffc_816_n_spl_0,
    ffc_816_n_spl_
  );


  buf

  (
    ffc_816_n_spl_1,
    ffc_816_n_spl_
  );


  buf

  (
    g1700_p_spl_,
    g1700_p
  );


  buf

  (
    g1717_n_spl_,
    g1717_n
  );


  buf

  (
    g1717_p_spl_,
    g1717_p
  );


  buf

  (
    g1696_p_spl_,
    g1696_p
  );


  buf

  (
    ffc_603_p_spl_,
    ffc_603_p
  );


  buf

  (
    g1723_n_spl_,
    g1723_n
  );


  buf

  (
    ffc_769_p_spl_,
    ffc_769_p
  );


  buf

  (
    ffc_769_p_spl_0,
    ffc_769_p_spl_
  );


  buf

  (
    ffc_769_p_spl_1,
    ffc_769_p_spl_
  );


  buf

  (
    ffc_844_p_spl_,
    ffc_844_p
  );


  buf

  (
    ffc_844_p_spl_0,
    ffc_844_p_spl_
  );


  buf

  (
    ffc_844_p_spl_1,
    ffc_844_p_spl_
  );


  buf

  (
    ffc_769_n_spl_,
    ffc_769_n
  );


  buf

  (
    ffc_844_n_spl_,
    ffc_844_n
  );


  buf

  (
    ffc_596_p_spl_,
    ffc_596_p
  );


  buf

  (
    ffc_596_p_spl_0,
    ffc_596_p_spl_
  );


  buf

  (
    ffc_556_n_spl_,
    ffc_556_n
  );


  buf

  (
    ffc_556_n_spl_0,
    ffc_556_n_spl_
  );


  buf

  (
    ffc_556_n_spl_1,
    ffc_556_n_spl_
  );


  buf

  (
    ffc_463_n_spl_,
    ffc_463_n
  );


  buf

  (
    ffc_463_n_spl_0,
    ffc_463_n_spl_
  );


  buf

  (
    ffc_463_n_spl_00,
    ffc_463_n_spl_0
  );


  buf

  (
    ffc_463_n_spl_000,
    ffc_463_n_spl_00
  );


  buf

  (
    ffc_463_n_spl_001,
    ffc_463_n_spl_00
  );


  buf

  (
    ffc_463_n_spl_01,
    ffc_463_n_spl_0
  );


  buf

  (
    ffc_463_n_spl_010,
    ffc_463_n_spl_01
  );


  buf

  (
    ffc_463_n_spl_1,
    ffc_463_n_spl_
  );


  buf

  (
    ffc_463_n_spl_10,
    ffc_463_n_spl_1
  );


  buf

  (
    ffc_463_n_spl_11,
    ffc_463_n_spl_1
  );


  buf

  (
    ffc_556_p_spl_,
    ffc_556_p
  );


  buf

  (
    ffc_556_p_spl_0,
    ffc_556_p_spl_
  );


  buf

  (
    ffc_556_p_spl_1,
    ffc_556_p_spl_
  );


  buf

  (
    ffc_460_p_spl_,
    ffc_460_p
  );


  buf

  (
    ffc_460_p_spl_0,
    ffc_460_p_spl_
  );


  buf

  (
    ffc_460_p_spl_00,
    ffc_460_p_spl_0
  );


  buf

  (
    ffc_460_p_spl_000,
    ffc_460_p_spl_00
  );


  buf

  (
    ffc_460_p_spl_001,
    ffc_460_p_spl_00
  );


  buf

  (
    ffc_460_p_spl_01,
    ffc_460_p_spl_0
  );


  buf

  (
    ffc_460_p_spl_010,
    ffc_460_p_spl_01
  );


  buf

  (
    ffc_460_p_spl_1,
    ffc_460_p_spl_
  );


  buf

  (
    ffc_460_p_spl_10,
    ffc_460_p_spl_1
  );


  buf

  (
    ffc_460_p_spl_11,
    ffc_460_p_spl_1
  );


  buf

  (
    ffc_527_n_spl_,
    ffc_527_n
  );


  buf

  (
    ffc_527_n_spl_0,
    ffc_527_n_spl_
  );


  buf

  (
    ffc_527_p_spl_,
    ffc_527_p
  );


  buf

  (
    ffc_527_p_spl_0,
    ffc_527_p_spl_
  );


  buf

  (
    ffc_590_n_spl_,
    ffc_590_n
  );


  buf

  (
    ffc_590_n_spl_0,
    ffc_590_n_spl_
  );


  buf

  (
    ffc_590_p_spl_,
    ffc_590_p
  );


  buf

  (
    ffc_590_p_spl_0,
    ffc_590_p_spl_
  );


  buf

  (
    ffc_390_p_spl_,
    ffc_390_p
  );


  buf

  (
    ffc_390_p_spl_0,
    ffc_390_p_spl_
  );


  buf

  (
    ffc_390_p_spl_00,
    ffc_390_p_spl_0
  );


  buf

  (
    ffc_390_p_spl_1,
    ffc_390_p_spl_
  );


  buf

  (
    g1711_n_spl_,
    g1711_n
  );


  buf

  (
    g1711_n_spl_0,
    g1711_n_spl_
  );


  buf

  (
    ffc_390_n_spl_,
    ffc_390_n
  );


  buf

  (
    ffc_390_n_spl_0,
    ffc_390_n_spl_
  );


  buf

  (
    ffc_390_n_spl_1,
    ffc_390_n_spl_
  );


  buf

  (
    g1711_p_spl_,
    g1711_p
  );


  buf

  (
    g1756_p_spl_,
    g1756_p
  );


  buf

  (
    ffc_839_p_spl_,
    ffc_839_p
  );


  buf

  (
    ffc_839_p_spl_0,
    ffc_839_p_spl_
  );


  buf

  (
    ffc_839_p_spl_00,
    ffc_839_p_spl_0
  );


  buf

  (
    ffc_839_p_spl_000,
    ffc_839_p_spl_00
  );


  buf

  (
    ffc_839_p_spl_001,
    ffc_839_p_spl_00
  );


  buf

  (
    ffc_839_p_spl_01,
    ffc_839_p_spl_0
  );


  buf

  (
    ffc_839_p_spl_1,
    ffc_839_p_spl_
  );


  buf

  (
    ffc_839_p_spl_10,
    ffc_839_p_spl_1
  );


  buf

  (
    ffc_839_p_spl_11,
    ffc_839_p_spl_1
  );


  buf

  (
    ffc_859_p_spl_,
    ffc_859_p
  );


  buf

  (
    ffc_839_n_spl_,
    ffc_839_n
  );


  buf

  (
    ffc_839_n_spl_0,
    ffc_839_n_spl_
  );


  buf

  (
    ffc_839_n_spl_00,
    ffc_839_n_spl_0
  );


  buf

  (
    ffc_839_n_spl_000,
    ffc_839_n_spl_00
  );


  buf

  (
    ffc_839_n_spl_01,
    ffc_839_n_spl_0
  );


  buf

  (
    ffc_839_n_spl_1,
    ffc_839_n_spl_
  );


  buf

  (
    ffc_839_n_spl_10,
    ffc_839_n_spl_1
  );


  buf

  (
    ffc_839_n_spl_11,
    ffc_839_n_spl_1
  );


  buf

  (
    ffc_857_p_spl_,
    ffc_857_p
  );


  buf

  (
    ffc_857_p_spl_0,
    ffc_857_p_spl_
  );


  buf

  (
    g1721_n_spl_,
    g1721_n
  );


  buf

  (
    g1721_n_spl_0,
    g1721_n_spl_
  );


  buf

  (
    ffc_858_p_spl_,
    ffc_858_p
  );


  buf

  (
    ffc_858_p_spl_0,
    ffc_858_p_spl_
  );


  buf

  (
    g1720_n_spl_,
    g1720_n
  );


  buf

  (
    g1720_n_spl_0,
    g1720_n_spl_
  );


  buf

  (
    ffc_861_p_spl_,
    ffc_861_p
  );


  buf

  (
    ffc_863_p_spl_,
    ffc_863_p
  );


  buf

  (
    ffc_863_p_spl_0,
    ffc_863_p_spl_
  );


  buf

  (
    ffc_863_p_spl_00,
    ffc_863_p_spl_0
  );


  buf

  (
    ffc_863_p_spl_000,
    ffc_863_p_spl_00
  );


  buf

  (
    ffc_863_p_spl_001,
    ffc_863_p_spl_00
  );


  buf

  (
    ffc_863_p_spl_01,
    ffc_863_p_spl_0
  );


  buf

  (
    ffc_863_p_spl_010,
    ffc_863_p_spl_01
  );


  buf

  (
    ffc_863_p_spl_011,
    ffc_863_p_spl_01
  );


  buf

  (
    ffc_863_p_spl_1,
    ffc_863_p_spl_
  );


  buf

  (
    ffc_863_p_spl_10,
    ffc_863_p_spl_1
  );


  buf

  (
    ffc_863_p_spl_11,
    ffc_863_p_spl_1
  );


  buf

  (
    ffc_863_n_spl_,
    ffc_863_n
  );


  buf

  (
    ffc_863_n_spl_0,
    ffc_863_n_spl_
  );


  buf

  (
    ffc_863_n_spl_00,
    ffc_863_n_spl_0
  );


  buf

  (
    ffc_863_n_spl_000,
    ffc_863_n_spl_00
  );


  buf

  (
    ffc_863_n_spl_001,
    ffc_863_n_spl_00
  );


  buf

  (
    ffc_863_n_spl_01,
    ffc_863_n_spl_0
  );


  buf

  (
    ffc_863_n_spl_010,
    ffc_863_n_spl_01
  );


  buf

  (
    ffc_863_n_spl_1,
    ffc_863_n_spl_
  );


  buf

  (
    ffc_863_n_spl_10,
    ffc_863_n_spl_1
  );


  buf

  (
    ffc_863_n_spl_11,
    ffc_863_n_spl_1
  );


  buf

  (
    g1704_p_spl_,
    g1704_p
  );


  buf

  (
    g1719_p_spl_,
    g1719_p
  );


  buf

  (
    g1719_p_spl_0,
    g1719_p_spl_
  );


  buf

  (
    g1772_n_spl_,
    g1772_n
  );


  buf

  (
    g1719_n_spl_,
    g1719_n
  );


  buf

  (
    g1772_p_spl_,
    g1772_p
  );


  buf

  (
    g1773_n_spl_,
    g1773_n
  );


  buf

  (
    g1773_p_spl_,
    g1773_p
  );


  buf

  (
    ffc_850_p_spl_,
    ffc_850_p
  );


  buf

  (
    ffc_852_p_spl_,
    ffc_852_p
  );


  buf

  (
    g1699_p_spl_,
    g1699_p
  );


  buf

  (
    g1699_p_spl_0,
    g1699_p_spl_
  );


  buf

  (
    g1781_p_spl_,
    g1781_p
  );


  buf

  (
    g1699_n_spl_,
    g1699_n
  );


  buf

  (
    g1699_n_spl_0,
    g1699_n_spl_
  );


  buf

  (
    g1699_n_spl_1,
    g1699_n_spl_
  );


  buf

  (
    g1781_n_spl_,
    g1781_n
  );


  buf

  (
    g1712_p_spl_,
    g1712_p
  );


  buf

  (
    g1712_p_spl_0,
    g1712_p_spl_
  );


  buf

  (
    g1785_p_spl_,
    g1785_p
  );


  buf

  (
    ffc_854_p_spl_,
    ffc_854_p
  );


  buf

  (
    ffc_848_p_spl_,
    ffc_848_p
  );


  buf

  (
    ffc_848_p_spl_0,
    ffc_848_p_spl_
  );


  buf

  (
    g1761_n_spl_,
    g1761_n
  );


  buf

  (
    g1761_n_spl_0,
    g1761_n_spl_
  );


  buf

  (
    ffc_856_p_spl_,
    ffc_856_p
  );


  buf

  (
    ffc_856_p_spl_0,
    ffc_856_p_spl_
  );


  buf

  (
    g1722_n_spl_,
    g1722_n
  );


  buf

  (
    g1722_n_spl_0,
    g1722_n_spl_
  );


  buf

  (
    g1763_n_spl_,
    g1763_n
  );


  buf

  (
    g1763_n_spl_0,
    g1763_n_spl_
  );


  buf

  (
    g1763_n_spl_1,
    g1763_n_spl_
  );


  buf

  (
    ffc_846_p_spl_,
    ffc_846_p
  );


  buf

  (
    ffc_847_p_spl_,
    ffc_847_p
  );


  buf

  (
    ffc_388_p_spl_,
    ffc_388_p
  );


  buf

  (
    ffc_388_p_spl_0,
    ffc_388_p_spl_
  );


  buf

  (
    g1780_n_spl_,
    g1780_n
  );


  buf

  (
    g1780_n_spl_0,
    g1780_n_spl_
  );


  buf

  (
    ffc_392_p_spl_,
    ffc_392_p
  );


  buf

  (
    ffc_392_p_spl_0,
    ffc_392_p_spl_
  );


  buf

  (
    g1777_n_spl_,
    g1777_n
  );


  buf

  (
    g1777_n_spl_0,
    g1777_n_spl_
  );


  buf

  (
    ffc_393_p_spl_,
    ffc_393_p
  );


  buf

  (
    ffc_393_p_spl_0,
    ffc_393_p_spl_
  );


  buf

  (
    g1790_n_spl_,
    g1790_n
  );


  buf

  (
    g1790_n_spl_0,
    g1790_n_spl_
  );


  buf

  (
    ffc_849_p_spl_,
    ffc_849_p
  );


  buf

  (
    ffc_849_p_spl_0,
    ffc_849_p_spl_
  );


  buf

  (
    g1767_n_spl_,
    g1767_n
  );


  buf

  (
    g1767_n_spl_0,
    g1767_n_spl_
  );


  buf

  (
    g1807_n_spl_,
    g1807_n
  );


  buf

  (
    g1797_p_spl_,
    g1797_p
  );


  buf

  (
    g1799_p_spl_,
    g1799_p
  );


  buf

  (
    g1799_p_spl_0,
    g1799_p_spl_
  );


  buf

  (
    ffc_497_n_spl_,
    ffc_497_n
  );


  buf

  (
    ffc_497_n_spl_0,
    ffc_497_n_spl_
  );


  buf

  (
    ffc_497_n_spl_00,
    ffc_497_n_spl_0
  );


  buf

  (
    ffc_497_n_spl_000,
    ffc_497_n_spl_00
  );


  buf

  (
    ffc_497_n_spl_001,
    ffc_497_n_spl_00
  );


  buf

  (
    ffc_497_n_spl_01,
    ffc_497_n_spl_0
  );


  buf

  (
    ffc_497_n_spl_010,
    ffc_497_n_spl_01
  );


  buf

  (
    ffc_497_n_spl_1,
    ffc_497_n_spl_
  );


  buf

  (
    ffc_497_n_spl_10,
    ffc_497_n_spl_1
  );


  buf

  (
    ffc_497_n_spl_11,
    ffc_497_n_spl_1
  );


  buf

  (
    ffc_497_p_spl_,
    ffc_497_p
  );


  buf

  (
    ffc_497_p_spl_0,
    ffc_497_p_spl_
  );


  buf

  (
    ffc_497_p_spl_00,
    ffc_497_p_spl_0
  );


  buf

  (
    ffc_497_p_spl_000,
    ffc_497_p_spl_00
  );


  buf

  (
    ffc_497_p_spl_001,
    ffc_497_p_spl_00
  );


  buf

  (
    ffc_497_p_spl_01,
    ffc_497_p_spl_0
  );


  buf

  (
    ffc_497_p_spl_010,
    ffc_497_p_spl_01
  );


  buf

  (
    ffc_497_p_spl_011,
    ffc_497_p_spl_01
  );


  buf

  (
    ffc_497_p_spl_1,
    ffc_497_p_spl_
  );


  buf

  (
    ffc_497_p_spl_10,
    ffc_497_p_spl_1
  );


  buf

  (
    ffc_497_p_spl_100,
    ffc_497_p_spl_10
  );


  buf

  (
    ffc_497_p_spl_101,
    ffc_497_p_spl_10
  );


  buf

  (
    ffc_497_p_spl_11,
    ffc_497_p_spl_1
  );


  buf

  (
    ffc_528_n_spl_,
    ffc_528_n
  );


  buf

  (
    ffc_528_n_spl_0,
    ffc_528_n_spl_
  );


  buf

  (
    ffc_528_p_spl_,
    ffc_528_p
  );


  buf

  (
    ffc_528_p_spl_0,
    ffc_528_p_spl_
  );


  buf

  (
    ffc_493_n_spl_,
    ffc_493_n
  );


  buf

  (
    ffc_493_n_spl_0,
    ffc_493_n_spl_
  );


  buf

  (
    ffc_204_p_spl_,
    ffc_204_p
  );


  buf

  (
    ffc_493_p_spl_,
    ffc_493_p
  );


  buf

  (
    ffc_493_p_spl_0,
    ffc_493_p_spl_
  );


  buf

  (
    ffc_604_n_spl_,
    ffc_604_n
  );


  buf

  (
    ffc_604_p_spl_,
    ffc_604_p
  );


  buf

  (
    ffc_605_p_spl_,
    ffc_605_p
  );


  buf

  (
    ffc_605_p_spl_0,
    ffc_605_p_spl_
  );


  buf

  (
    ffc_615_p_spl_,
    ffc_615_p
  );


  buf

  (
    ffc_791_p_spl_,
    ffc_791_p
  );


  buf

  (
    ffc_811_p_spl_,
    ffc_811_p
  );


  buf

  (
    ffc_791_n_spl_,
    ffc_791_n
  );


  buf

  (
    ffc_811_n_spl_,
    ffc_811_n
  );


  buf

  (
    g1831_p_spl_,
    g1831_p
  );


  buf

  (
    g1834_n_spl_,
    g1834_n
  );


  buf

  (
    g1831_n_spl_,
    g1831_n
  );


  buf

  (
    g1834_p_spl_,
    g1834_p
  );


  buf

  (
    ffc_578_p_spl_,
    ffc_578_p
  );


  buf

  (
    g1692_p_spl_,
    g1692_p
  );


  buf

  (
    g1692_p_spl_0,
    g1692_p_spl_
  );


  buf

  (
    g1840_n_spl_,
    g1840_n
  );


  buf

  (
    g1692_n_spl_,
    g1692_n
  );


  buf

  (
    g1692_n_spl_0,
    g1692_n_spl_
  );


  buf

  (
    g1840_p_spl_,
    g1840_p
  );


  buf

  (
    g1755_n_spl_,
    g1755_n
  );


  buf

  (
    g1737_n_spl_,
    g1737_n
  );


  buf

  (
    g1746_n_spl_,
    g1746_n
  );


  buf

  (
    g1854_p_spl_,
    g1854_p
  );


  buf

  (
    g1855_n_spl_,
    g1855_n
  );


  buf

  (
    g1854_n_spl_,
    g1854_n
  );


  buf

  (
    g1855_p_spl_,
    g1855_p
  );


  buf

  (
    ffc_802_p_spl_,
    ffc_802_p
  );


  buf

  (
    ffc_800_p_spl_,
    ffc_800_p
  );


  buf

  (
    g1859_p_spl_,
    g1859_p
  );


  buf

  (
    g1860_p_spl_,
    g1860_p
  );


  buf

  (
    g1859_n_spl_,
    g1859_n
  );


  buf

  (
    g1860_n_spl_,
    g1860_n
  );


  buf

  (
    ffc_772_p_spl_,
    ffc_772_p
  );


  buf

  (
    ffc_772_p_spl_0,
    ffc_772_p_spl_
  );


  buf

  (
    ffc_772_p_spl_1,
    ffc_772_p_spl_
  );


  buf

  (
    ffc_6_n_spl_,
    ffc_6_n
  );


  buf

  (
    ffc_772_n_spl_,
    ffc_772_n
  );


  buf

  (
    ffc_772_n_spl_0,
    ffc_772_n_spl_
  );


  buf

  (
    ffc_771_n_spl_,
    ffc_771_n
  );


  buf

  (
    ffc_771_n_spl_0,
    ffc_771_n_spl_
  );


  buf

  (
    ffc_771_n_spl_1,
    ffc_771_n_spl_
  );


  buf

  (
    ffc_771_p_spl_,
    ffc_771_p
  );


  buf

  (
    ffc_771_p_spl_0,
    ffc_771_p_spl_
  );


  buf

  (
    ffc_771_p_spl_00,
    ffc_771_p_spl_0
  );


  buf

  (
    ffc_771_p_spl_1,
    ffc_771_p_spl_
  );


  buf

  (
    g1872_n_spl_,
    g1872_n
  );


  buf

  (
    g1872_n_spl_0,
    g1872_n_spl_
  );


  buf

  (
    g1872_n_spl_00,
    g1872_n_spl_0
  );


  buf

  (
    g1872_n_spl_1,
    g1872_n_spl_
  );


  buf

  (
    g1872_p_spl_,
    g1872_p
  );


  buf

  (
    g1872_p_spl_0,
    g1872_p_spl_
  );


  buf

  (
    g1872_p_spl_00,
    g1872_p_spl_0
  );


  buf

  (
    g1872_p_spl_1,
    g1872_p_spl_
  );


  buf

  (
    ffc_659_p_spl_,
    ffc_659_p
  );


  buf

  (
    ffc_659_n_spl_,
    ffc_659_n
  );


  buf

  (
    ffc_659_n_spl_0,
    ffc_659_n_spl_
  );


  buf

  (
    g1877_n_spl_,
    g1877_n
  );


  buf

  (
    g1724_p_spl_,
    g1724_p
  );


  buf

  (
    ffc_375_p_spl_,
    ffc_375_p
  );


  buf

  (
    ffc_375_p_spl_0,
    ffc_375_p_spl_
  );


  buf

  (
    g1884_n_spl_,
    g1884_n
  );


  buf

  (
    ffc_609_p_spl_,
    ffc_609_p
  );


  buf

  (
    g1693_n_spl_,
    g1693_n
  );


  buf

  (
    g1891_p_spl_,
    g1891_p
  );


  buf

  (
    g1728_n_spl_,
    g1728_n
  );


  buf

  (
    ffc_592_p_spl_,
    ffc_592_p
  );


  buf

  (
    g1895_n_spl_,
    g1895_n
  );


  buf

  (
    ffc_364_p_spl_,
    ffc_364_p
  );


  buf

  (
    ffc_790_n_spl_,
    ffc_790_n
  );


  buf

  (
    ffc_790_n_spl_0,
    ffc_790_n_spl_
  );


  buf

  (
    g1708_n_spl_,
    g1708_n
  );


  buf

  (
    ffc_539_p_spl_,
    ffc_539_p
  );


  buf

  (
    ffc_539_p_spl_0,
    ffc_539_p_spl_
  );


  buf

  (
    ffc_539_n_spl_,
    ffc_539_n
  );


  buf

  (
    ffc_539_n_spl_0,
    ffc_539_n_spl_
  );


  buf

  (
    ffc_526_p_spl_,
    ffc_526_p
  );


  buf

  (
    ffc_526_p_spl_0,
    ffc_526_p_spl_
  );


  buf

  (
    ffc_526_n_spl_,
    ffc_526_n
  );


  buf

  (
    ffc_526_n_spl_0,
    ffc_526_n_spl_
  );


  buf

  (
    ffc_540_p_spl_,
    ffc_540_p
  );


  buf

  (
    ffc_540_p_spl_0,
    ffc_540_p_spl_
  );


  buf

  (
    ffc_540_n_spl_,
    ffc_540_n
  );


  buf

  (
    ffc_540_n_spl_0,
    ffc_540_n_spl_
  );


  buf

  (
    ffc_536_n_spl_,
    ffc_536_n
  );


  buf

  (
    ffc_536_n_spl_0,
    ffc_536_n_spl_
  );


  buf

  (
    ffc_536_n_spl_1,
    ffc_536_n_spl_
  );


  buf

  (
    ffc_536_p_spl_,
    ffc_536_p
  );


  buf

  (
    ffc_536_p_spl_0,
    ffc_536_p_spl_
  );


  buf

  (
    ffc_536_p_spl_1,
    ffc_536_p_spl_
  );


  buf

  (
    ffc_598_n_spl_,
    ffc_598_n
  );


  buf

  (
    ffc_598_n_spl_0,
    ffc_598_n_spl_
  );


  buf

  (
    ffc_598_n_spl_1,
    ffc_598_n_spl_
  );


  buf

  (
    ffc_598_p_spl_,
    ffc_598_p
  );


  buf

  (
    ffc_598_p_spl_0,
    ffc_598_p_spl_
  );


  buf

  (
    ffc_598_p_spl_1,
    ffc_598_p_spl_
  );


  buf

  (
    ffc_557_n_spl_,
    ffc_557_n
  );


  buf

  (
    ffc_557_n_spl_0,
    ffc_557_n_spl_
  );


  buf

  (
    ffc_557_p_spl_,
    ffc_557_p
  );


  buf

  (
    ffc_557_p_spl_0,
    ffc_557_p_spl_
  );


  buf

  (
    ffc_549_n_spl_,
    ffc_549_n
  );


  buf

  (
    ffc_549_n_spl_0,
    ffc_549_n_spl_
  );


  buf

  (
    ffc_549_p_spl_,
    ffc_549_p
  );


  buf

  (
    ffc_549_p_spl_0,
    ffc_549_p_spl_
  );


  buf

  (
    ffc_785_n_spl_,
    ffc_785_n
  );


  buf

  (
    ffc_786_p_spl_,
    ffc_786_p
  );


  buf

  (
    ffc_785_p_spl_,
    ffc_785_p
  );


  buf

  (
    ffc_786_n_spl_,
    ffc_786_n
  );


  buf

  (
    ffc_789_n_spl_,
    ffc_789_n
  );


  buf

  (
    ffc_789_p_spl_,
    ffc_789_p
  );


  buf

  (
    ffc_790_p_spl_,
    ffc_790_p
  );


  buf

  (
    ffc_790_p_spl_0,
    ffc_790_p_spl_
  );


  buf

  (
    g1982_n_spl_,
    g1982_n
  );


  buf

  (
    g1985_p_spl_,
    g1985_p
  );


  buf

  (
    g1982_p_spl_,
    g1982_p
  );


  buf

  (
    g1985_n_spl_,
    g1985_n
  );


  buf

  (
    ffc_784_n_spl_,
    ffc_784_n
  );


  buf

  (
    ffc_788_p_spl_,
    ffc_788_p
  );


  buf

  (
    ffc_784_p_spl_,
    ffc_784_p
  );


  buf

  (
    ffc_788_n_spl_,
    ffc_788_n
  );


  buf

  (
    ffc_787_n_spl_,
    ffc_787_n
  );


  buf

  (
    ffc_810_n_spl_,
    ffc_810_n
  );


  buf

  (
    ffc_787_p_spl_,
    ffc_787_p
  );


  buf

  (
    ffc_810_p_spl_,
    ffc_810_p
  );


  buf

  (
    g1991_p_spl_,
    g1991_p
  );


  buf

  (
    g1994_n_spl_,
    g1994_n
  );


  buf

  (
    g1991_n_spl_,
    g1991_n
  );


  buf

  (
    g1994_p_spl_,
    g1994_p
  );


  buf

  (
    ffc_350_p_spl_,
    ffc_350_p
  );


  buf

  (
    ffc_350_p_spl_0,
    ffc_350_p_spl_
  );


  buf

  (
    ffc_529_p_spl_,
    ffc_529_p
  );


  buf

  (
    ffc_350_n_spl_,
    ffc_350_n
  );


  buf

  (
    ffc_350_n_spl_0,
    ffc_350_n_spl_
  );


  buf

  (
    ffc_529_n_spl_,
    ffc_529_n
  );


  buf

  (
    ffc_608_p_spl_,
    ffc_608_p
  );


  buf

  (
    ffc_614_p_spl_,
    ffc_614_p
  );


  buf

  (
    ffc_640_p_spl_,
    ffc_640_p
  );


  buf

  (
    g2035_n_spl_,
    g2035_n
  );


  buf

  (
    g2038_p_spl_,
    g2038_p
  );


  buf

  (
    ffc_375_n_spl_,
    ffc_375_n
  );


  buf

  (
    ffc_571_p_spl_,
    ffc_571_p
  );


  buf

  (
    ffc_571_n_spl_,
    ffc_571_n
  );


  buf

  (
    g2046_n_spl_,
    g2046_n
  );


  buf

  (
    g2049_p_spl_,
    g2049_p
  );


  buf

  (
    g2054_n_spl_,
    g2054_n
  );


  buf

  (
    g2057_n_spl_,
    g2057_n
  );


  buf

  (
    g2069_p_spl_,
    g2069_p
  );


  buf

  (
    g2070_n_spl_,
    g2070_n
  );


  buf

  (
    g2069_n_spl_,
    g2069_n
  );


  buf

  (
    g2070_p_spl_,
    g2070_p
  );


  buf

  (
    ffc_424_n_spl_,
    ffc_424_n
  );


  buf

  (
    ffc_424_n_spl_0,
    ffc_424_n_spl_
  );


  buf

  (
    ffc_424_n_spl_1,
    ffc_424_n_spl_
  );


  buf

  (
    ffc_424_p_spl_,
    ffc_424_p
  );


  buf

  (
    ffc_424_p_spl_0,
    ffc_424_p_spl_
  );


  buf

  (
    ffc_424_p_spl_1,
    ffc_424_p_spl_
  );


  buf

  (
    g2075_p_spl_,
    g2075_p
  );


  buf

  (
    g2076_p_spl_,
    g2076_p
  );


  buf

  (
    g2075_n_spl_,
    g2075_n
  );


  buf

  (
    g2076_n_spl_,
    g2076_n
  );


  buf

  (
    g2082_n_spl_,
    g2082_n
  );


  buf

  (
    g2082_p_spl_,
    g2082_p
  );


  buf

  (
    g2085_p_spl_,
    g2085_p
  );


  buf

  (
    g2085_n_spl_,
    g2085_n
  );


  buf

  (
    g1793_p_spl_,
    g1793_p
  );


  buf

  (
    g1796_p_spl_,
    g1796_p
  );


  buf

  (
    g1796_p_spl_0,
    g1796_p_spl_
  );


  buf

  (
    g1762_p_spl_,
    g1762_p
  );


  buf

  (
    ffc_628_n_spl_,
    ffc_628_n
  );


  buf

  (
    ffc_832_n_spl_,
    ffc_832_n
  );


  buf

  (
    ffc_832_n_spl_0,
    ffc_832_n_spl_
  );


  buf

  (
    ffc_832_n_spl_00,
    ffc_832_n_spl_0
  );


  buf

  (
    ffc_832_n_spl_000,
    ffc_832_n_spl_00
  );


  buf

  (
    ffc_832_n_spl_001,
    ffc_832_n_spl_00
  );


  buf

  (
    ffc_832_n_spl_01,
    ffc_832_n_spl_0
  );


  buf

  (
    ffc_832_n_spl_010,
    ffc_832_n_spl_01
  );


  buf

  (
    ffc_832_n_spl_011,
    ffc_832_n_spl_01
  );


  buf

  (
    ffc_832_n_spl_1,
    ffc_832_n_spl_
  );


  buf

  (
    ffc_832_n_spl_10,
    ffc_832_n_spl_1
  );


  buf

  (
    ffc_832_n_spl_100,
    ffc_832_n_spl_10
  );


  buf

  (
    ffc_832_n_spl_101,
    ffc_832_n_spl_10
  );


  buf

  (
    ffc_832_n_spl_11,
    ffc_832_n_spl_1
  );


  buf

  (
    ffc_832_n_spl_110,
    ffc_832_n_spl_11
  );


  buf

  (
    ffc_832_n_spl_111,
    ffc_832_n_spl_11
  );


  buf

  (
    ffc_628_p_spl_,
    ffc_628_p
  );


  buf

  (
    ffc_628_p_spl_0,
    ffc_628_p_spl_
  );


  buf

  (
    ffc_833_n_spl_,
    ffc_833_n
  );


  buf

  (
    ffc_833_n_spl_0,
    ffc_833_n_spl_
  );


  buf

  (
    ffc_833_n_spl_00,
    ffc_833_n_spl_0
  );


  buf

  (
    ffc_833_n_spl_000,
    ffc_833_n_spl_00
  );


  buf

  (
    ffc_833_n_spl_001,
    ffc_833_n_spl_00
  );


  buf

  (
    ffc_833_n_spl_01,
    ffc_833_n_spl_0
  );


  buf

  (
    ffc_833_n_spl_010,
    ffc_833_n_spl_01
  );


  buf

  (
    ffc_833_n_spl_011,
    ffc_833_n_spl_01
  );


  buf

  (
    ffc_833_n_spl_1,
    ffc_833_n_spl_
  );


  buf

  (
    ffc_833_n_spl_10,
    ffc_833_n_spl_1
  );


  buf

  (
    ffc_833_n_spl_100,
    ffc_833_n_spl_10
  );


  buf

  (
    ffc_833_n_spl_101,
    ffc_833_n_spl_10
  );


  buf

  (
    ffc_833_n_spl_11,
    ffc_833_n_spl_1
  );


  buf

  (
    ffc_833_n_spl_110,
    ffc_833_n_spl_11
  );


  buf

  (
    ffc_834_p_spl_,
    ffc_834_p
  );


  buf

  (
    ffc_834_p_spl_0,
    ffc_834_p_spl_
  );


  buf

  (
    ffc_834_p_spl_00,
    ffc_834_p_spl_0
  );


  buf

  (
    ffc_834_p_spl_000,
    ffc_834_p_spl_00
  );


  buf

  (
    ffc_834_p_spl_001,
    ffc_834_p_spl_00
  );


  buf

  (
    ffc_834_p_spl_01,
    ffc_834_p_spl_0
  );


  buf

  (
    ffc_834_p_spl_010,
    ffc_834_p_spl_01
  );


  buf

  (
    ffc_834_p_spl_011,
    ffc_834_p_spl_01
  );


  buf

  (
    ffc_834_p_spl_1,
    ffc_834_p_spl_
  );


  buf

  (
    ffc_834_p_spl_10,
    ffc_834_p_spl_1
  );


  buf

  (
    ffc_834_p_spl_100,
    ffc_834_p_spl_10
  );


  buf

  (
    ffc_834_p_spl_101,
    ffc_834_p_spl_10
  );


  buf

  (
    ffc_834_p_spl_11,
    ffc_834_p_spl_1
  );


  buf

  (
    ffc_831_p_spl_,
    ffc_831_p
  );


  buf

  (
    ffc_831_p_spl_0,
    ffc_831_p_spl_
  );


  buf

  (
    ffc_831_p_spl_00,
    ffc_831_p_spl_0
  );


  buf

  (
    ffc_831_p_spl_000,
    ffc_831_p_spl_00
  );


  buf

  (
    ffc_831_p_spl_001,
    ffc_831_p_spl_00
  );


  buf

  (
    ffc_831_p_spl_01,
    ffc_831_p_spl_0
  );


  buf

  (
    ffc_831_p_spl_010,
    ffc_831_p_spl_01
  );


  buf

  (
    ffc_831_p_spl_011,
    ffc_831_p_spl_01
  );


  buf

  (
    ffc_831_p_spl_1,
    ffc_831_p_spl_
  );


  buf

  (
    ffc_831_p_spl_10,
    ffc_831_p_spl_1
  );


  buf

  (
    ffc_831_p_spl_100,
    ffc_831_p_spl_10
  );


  buf

  (
    ffc_831_p_spl_101,
    ffc_831_p_spl_10
  );


  buf

  (
    ffc_831_p_spl_11,
    ffc_831_p_spl_1
  );


  buf

  (
    ffc_831_p_spl_110,
    ffc_831_p_spl_11
  );


  buf

  (
    ffc_633_n_spl_,
    ffc_633_n
  );


  buf

  (
    ffc_633_p_spl_,
    ffc_633_p
  );


  buf

  (
    ffc_633_p_spl_0,
    ffc_633_p_spl_
  );


  buf

  (
    ffc_677_p_spl_,
    ffc_677_p
  );


  buf

  (
    ffc_780_p_spl_,
    ffc_780_p
  );


  buf

  (
    ffc_355_p_spl_,
    ffc_355_p
  );


  buf

  (
    ffc_355_p_spl_0,
    ffc_355_p_spl_
  );


  buf

  (
    ffc_346_p_spl_,
    ffc_346_p
  );


  buf

  (
    ffc_366_p_spl_,
    ffc_366_p
  );


  buf

  (
    ffc_367_p_spl_,
    ffc_367_p
  );


  buf

  (
    ffc_826_p_spl_,
    ffc_826_p
  );


  buf

  (
    ffc_826_p_spl_0,
    ffc_826_p_spl_
  );


  buf

  (
    ffc_826_p_spl_1,
    ffc_826_p_spl_
  );


  buf

  (
    ffc_826_n_spl_,
    ffc_826_n
  );


  buf

  (
    ffc_826_n_spl_0,
    ffc_826_n_spl_
  );


  buf

  (
    ffc_826_n_spl_1,
    ffc_826_n_spl_
  );


  buf

  (
    ffc_812_p_spl_,
    ffc_812_p
  );


  buf

  (
    g1758_p_spl_,
    g1758_p
  );


  buf

  (
    g1758_p_spl_0,
    g1758_p_spl_
  );


  buf

  (
    g2139_n_spl_,
    g2139_n
  );


  buf

  (
    g2139_n_spl_0,
    g2139_n_spl_
  );


  buf

  (
    ffc_825_n_spl_,
    ffc_825_n
  );


  buf

  (
    ffc_825_n_spl_0,
    ffc_825_n_spl_
  );


  buf

  (
    ffc_825_n_spl_1,
    ffc_825_n_spl_
  );


  buf

  (
    g1725_n_spl_,
    g1725_n
  );


  buf

  (
    g1758_n_spl_,
    g1758_n
  );


  buf

  (
    g1758_n_spl_0,
    g1758_n_spl_
  );


  buf

  (
    g1758_n_spl_1,
    g1758_n_spl_
  );


  buf

  (
    g2142_n_spl_,
    g2142_n
  );


  buf

  (
    ffc_671_n_spl_,
    ffc_671_n
  );


  buf

  (
    ffc_671_p_spl_,
    ffc_671_p
  );


  buf

  (
    ffc_671_p_spl_0,
    ffc_671_p_spl_
  );


  buf

  (
    ffc_756_n_spl_,
    ffc_756_n
  );


  buf

  (
    ffc_756_n_spl_0,
    ffc_756_n_spl_
  );


  buf

  (
    g2146_p_spl_,
    g2146_p
  );


  buf

  (
    ffc_756_p_spl_,
    ffc_756_p
  );


  buf

  (
    ffc_756_p_spl_0,
    ffc_756_p_spl_
  );


  buf

  (
    ffc_756_p_spl_1,
    ffc_756_p_spl_
  );


  buf

  (
    g2146_n_spl_,
    g2146_n
  );


  buf

  (
    ffc_672_p_spl_,
    ffc_672_p
  );


  buf

  (
    ffc_778_p_spl_,
    ffc_778_p
  );


  buf

  (
    ffc_825_p_spl_,
    ffc_825_p
  );


  buf

  (
    ffc_825_p_spl_0,
    ffc_825_p_spl_
  );


  buf

  (
    ffc_825_p_spl_1,
    ffc_825_p_spl_
  );


  buf

  (
    g2139_p_spl_,
    g2139_p
  );


  buf

  (
    g2139_p_spl_0,
    g2139_p_spl_
  );


  buf

  (
    g2151_n_spl_,
    g2151_n
  );


  buf

  (
    g2151_n_spl_0,
    g2151_n_spl_
  );


  buf

  (
    g2151_p_spl_,
    g2151_p
  );


  buf

  (
    g2151_p_spl_0,
    g2151_p_spl_
  );


  buf

  (
    g2157_n_spl_,
    g2157_n
  );


  buf

  (
    g1702_n_spl_,
    g1702_n
  );


  buf

  (
    g1702_n_spl_0,
    g1702_n_spl_
  );


  buf

  (
    g2161_p_spl_,
    g2161_p
  );


  buf

  (
    g1702_p_spl_,
    g1702_p
  );


  buf

  (
    g2161_n_spl_,
    g2161_n
  );


  buf

  (
    ffc_673_n_spl_,
    ffc_673_n
  );


  buf

  (
    ffc_673_p_spl_,
    ffc_673_p
  );


  buf

  (
    ffc_673_p_spl_0,
    ffc_673_p_spl_
  );


  buf

  (
    ffc_673_p_spl_1,
    ffc_673_p_spl_
  );


  buf

  (
    g2164_n_spl_,
    g2164_n
  );


  buf

  (
    g2165_p_spl_,
    g2165_p
  );


  buf

  (
    g1705_p_spl_,
    g1705_p
  );


  buf

  (
    ffc_674_p_spl_,
    ffc_674_p
  );


  buf

  (
    ffc_674_p_spl_0,
    ffc_674_p_spl_
  );


  buf

  (
    g2169_n_spl_,
    g2169_n
  );


  buf

  (
    ffc_674_n_spl_,
    ffc_674_n
  );


  buf

  (
    g2169_p_spl_,
    g2169_p
  );


  buf

  (
    g2167_n_spl_,
    g2167_n
  );


  buf

  (
    g2172_n_spl_,
    g2172_n
  );


  buf

  (
    g2172_n_spl_0,
    g2172_n_spl_
  );


  buf

  (
    g2096_n_spl_,
    g2096_n
  );


  buf

  (
    g1805_p_spl_,
    g1805_p
  );


  buf

  (
    g1808_p_spl_,
    g1808_p
  );


  buf

  (
    ffc_629_p_spl_,
    ffc_629_p
  );


  buf

  (
    ffc_358_p_spl_,
    ffc_358_p
  );


  buf

  (
    ffc_622_n_spl_,
    ffc_622_n
  );


  buf

  (
    ffc_622_p_spl_,
    ffc_622_p
  );


  buf

  (
    ffc_622_p_spl_0,
    ffc_622_p_spl_
  );


  buf

  (
    ffc_634_p_spl_,
    ffc_634_p
  );


  buf

  (
    ffc_621_n_spl_,
    ffc_621_n
  );


  buf

  (
    ffc_621_p_spl_,
    ffc_621_p
  );


  buf

  (
    ffc_621_p_spl_0,
    ffc_621_p_spl_
  );


  buf

  (
    ffc_635_p_spl_,
    ffc_635_p
  );


  buf

  (
    ffc_620_n_spl_,
    ffc_620_n
  );


  buf

  (
    ffc_620_p_spl_,
    ffc_620_p
  );


  buf

  (
    ffc_620_p_spl_0,
    ffc_620_p_spl_
  );


  buf

  (
    ffc_636_p_spl_,
    ffc_636_p
  );


  buf

  (
    ffc_627_n_spl_,
    ffc_627_n
  );


  buf

  (
    ffc_627_p_spl_,
    ffc_627_p
  );


  buf

  (
    ffc_627_p_spl_0,
    ffc_627_p_spl_
  );


  buf

  (
    ffc_650_p_spl_,
    ffc_650_p
  );


  buf

  (
    ffc_632_n_spl_,
    ffc_632_n
  );


  buf

  (
    ffc_632_p_spl_,
    ffc_632_p
  );


  buf

  (
    ffc_632_p_spl_0,
    ffc_632_p_spl_
  );


  buf

  (
    ffc_663_p_spl_,
    ffc_663_p
  );


  buf

  (
    ffc_631_n_spl_,
    ffc_631_n
  );


  buf

  (
    ffc_631_p_spl_,
    ffc_631_p
  );


  buf

  (
    ffc_631_p_spl_0,
    ffc_631_p_spl_
  );


  buf

  (
    ffc_664_p_spl_,
    ffc_664_p
  );


  buf

  (
    ffc_675_n_spl_,
    ffc_675_n
  );


  buf

  (
    ffc_675_p_spl_,
    ffc_675_p
  );


  buf

  (
    ffc_675_p_spl_0,
    ffc_675_p_spl_
  );


  buf

  (
    g1714_n_spl_,
    g1714_n
  );


  buf

  (
    g1714_n_spl_0,
    g1714_n_spl_
  );


  buf

  (
    g1714_p_spl_,
    g1714_p
  );


  buf

  (
    ffc_755_p_spl_,
    ffc_755_p
  );


  buf

  (
    g2253_n_spl_,
    g2253_n
  );


  buf

  (
    ffc_755_n_spl_,
    ffc_755_n
  );


  buf

  (
    g2253_p_spl_,
    g2253_p
  );


  buf

  (
    g2250_p_spl_,
    g2250_p
  );


  buf

  (
    g2259_n_spl_,
    g2259_n
  );


  buf

  (
    ffc_334_p_spl_,
    ffc_334_p
  );


  buf

  (
    g1768_n_spl_,
    g1768_n
  );


  buf

  (
    g2269_p_spl_,
    g2269_p
  );


  buf

  (
    g2272_p_spl_,
    g2272_p
  );


  buf

  (
    g1764_p_spl_,
    g1764_p
  );


  buf

  (
    g1764_p_spl_0,
    g1764_p_spl_
  );


  buf

  (
    g1809_p_spl_,
    g1809_p
  );


  buf

  (
    g2099_p_spl_,
    g2099_p
  );


  buf

  (
    g2099_p_spl_0,
    g2099_p_spl_
  );


  buf

  (
    g2275_n_spl_,
    g2275_n
  );


  buf

  (
    g2108_n_spl_,
    g2108_n
  );


  buf

  (
    g2108_n_spl_0,
    g2108_n_spl_
  );


  buf

  (
    g2123_n_spl_,
    g2123_n
  );


  buf

  (
    g2123_n_spl_0,
    g2123_n_spl_
  );


  buf

  (
    g2117_n_spl_,
    g2117_n
  );


  buf

  (
    g2117_n_spl_0,
    g2117_n_spl_
  );


  buf

  (
    g2126_p_spl_,
    g2126_p
  );


  buf

  (
    g2126_p_spl_0,
    g2126_p_spl_
  );


  buf

  (
    ffc_764_p_spl_,
    ffc_764_p
  );


  buf

  (
    ffc_764_p_spl_0,
    ffc_764_p_spl_
  );


  buf

  (
    ffc_764_n_spl_,
    ffc_764_n
  );


  buf

  (
    ffc_832_p_spl_,
    ffc_832_p
  );


  buf

  (
    ffc_832_p_spl_0,
    ffc_832_p_spl_
  );


  buf

  (
    ffc_832_p_spl_00,
    ffc_832_p_spl_0
  );


  buf

  (
    ffc_832_p_spl_1,
    ffc_832_p_spl_
  );


  buf

  (
    ffc_831_n_spl_,
    ffc_831_n
  );


  buf

  (
    ffc_831_n_spl_0,
    ffc_831_n_spl_
  );


  buf

  (
    ffc_831_n_spl_00,
    ffc_831_n_spl_0
  );


  buf

  (
    ffc_831_n_spl_1,
    ffc_831_n_spl_
  );


  buf

  (
    ffc_781_n_spl_,
    ffc_781_n
  );


  buf

  (
    ffc_781_n_spl_0,
    ffc_781_n_spl_
  );


  buf

  (
    ffc_781_n_spl_1,
    ffc_781_n_spl_
  );


  buf

  (
    ffc_781_p_spl_,
    ffc_781_p
  );


  buf

  (
    ffc_781_p_spl_0,
    ffc_781_p_spl_
  );


  buf

  (
    ffc_781_p_spl_00,
    ffc_781_p_spl_0
  );


  buf

  (
    ffc_781_p_spl_1,
    ffc_781_p_spl_
  );


  buf

  (
    ffc_833_p_spl_,
    ffc_833_p
  );


  buf

  (
    ffc_833_p_spl_0,
    ffc_833_p_spl_
  );


  buf

  (
    ffc_833_p_spl_1,
    ffc_833_p_spl_
  );


  buf

  (
    ffc_834_n_spl_,
    ffc_834_n
  );


  buf

  (
    ffc_834_n_spl_0,
    ffc_834_n_spl_
  );


  buf

  (
    ffc_834_n_spl_1,
    ffc_834_n_spl_
  );


  buf

  (
    g2120_n_spl_,
    g2120_n
  );


  buf

  (
    g2120_n_spl_0,
    g2120_n_spl_
  );


  buf

  (
    g2295_n_spl_,
    g2295_n
  );


  buf

  (
    ffc_648_n_spl_,
    ffc_648_n
  );


  buf

  (
    ffc_648_p_spl_,
    ffc_648_p
  );


  buf

  (
    ffc_648_p_spl_0,
    ffc_648_p_spl_
  );


  buf

  (
    ffc_679_p_spl_,
    ffc_679_p
  );


  buf

  (
    ffc_661_p_spl_,
    ffc_661_p
  );


  buf

  (
    ffc_661_p_spl_0,
    ffc_661_p_spl_
  );


  buf

  (
    ffc_661_n_spl_,
    ffc_661_n
  );


  buf

  (
    ffc_765_p_spl_,
    ffc_765_p
  );


  buf

  (
    g2306_n_spl_,
    g2306_n
  );


  buf

  (
    g2315_p_spl_,
    g2315_p
  );


  buf

  (
    ffc_779_p_spl_,
    ffc_779_p
  );


  buf

  (
    g1774_n_spl_,
    g1774_n
  );


  buf

  (
    g1787_n_spl_,
    g1787_n
  );


  buf

  (
    g1697_n_spl_,
    g1697_n
  );


  buf

  (
    g1697_n_spl_0,
    g1697_n_spl_
  );


  buf

  (
    g1701_p_spl_,
    g1701_p
  );


  buf

  (
    g1697_p_spl_,
    g1697_p
  );


  buf

  (
    g1701_n_spl_,
    g1701_n
  );


  buf

  (
    g1701_n_spl_0,
    g1701_n_spl_
  );


  buf

  (
    ffc_660_n_spl_,
    ffc_660_n
  );


  buf

  (
    ffc_660_n_spl_0,
    ffc_660_n_spl_
  );


  buf

  (
    ffc_660_n_spl_1,
    ffc_660_n_spl_
  );


  buf

  (
    ffc_660_p_spl_,
    ffc_660_p
  );


  buf

  (
    ffc_660_p_spl_0,
    ffc_660_p_spl_
  );


  buf

  (
    ffc_660_p_spl_00,
    ffc_660_p_spl_0
  );


  buf

  (
    ffc_660_p_spl_1,
    ffc_660_p_spl_
  );


  buf

  (
    ffc_763_p_spl_,
    ffc_763_p
  );


  buf

  (
    ffc_763_p_spl_0,
    ffc_763_p_spl_
  );


  buf

  (
    ffc_763_n_spl_,
    ffc_763_n
  );


  buf

  (
    ffc_442_n_spl_,
    ffc_442_n
  );


  buf

  (
    ffc_442_p_spl_,
    ffc_442_p
  );


  buf

  (
    g1716_n_spl_,
    g1716_n
  );


  buf

  (
    g1792_p_spl_,
    g1792_p
  );


  buf

  (
    ffc_396_p_spl_,
    ffc_396_p
  );


  buf

  (
    g2132_n_spl_,
    g2132_n
  );


  buf

  (
    ffc_397_p_spl_,
    ffc_397_p
  );


  buf

  (
    g1802_n_spl_,
    g1802_n
  );


  buf

  (
    g2133_n_spl_,
    g2133_n
  );


  buf

  (
    ffc_360_p_spl_,
    ffc_360_p
  );


  buf

  (
    ffc_362_p_spl_,
    ffc_362_p
  );


  buf

  (
    g2276_n_spl_,
    g2276_n
  );


  buf

  (
    g2276_n_spl_0,
    g2276_n_spl_
  );


  buf

  (
    g2137_p_spl_,
    g2137_p
  );


  buf

  (
    g2137_p_spl_0,
    g2137_p_spl_
  );


  buf

  (
    g2137_p_spl_1,
    g2137_p_spl_
  );


  buf

  (
    g2160_n_spl_,
    g2160_n
  );


  buf

  (
    g2160_n_spl_0,
    g2160_n_spl_
  );


  buf

  (
    g2175_p_spl_,
    g2175_p
  );


  buf

  (
    g2098_n_spl_,
    g2098_n
  );


  buf

  (
    g2135_p_spl_,
    g2135_p
  );


  buf

  (
    g1803_p_spl_,
    g1803_p
  );


  buf

  (
    g1804_p_spl_,
    g1804_p
  );


  buf

  (
    g2177_n_spl_,
    g2177_n
  );


  buf

  (
    ffc_391_p_spl_,
    ffc_391_p
  );


  buf

  (
    ffc_391_p_spl_0,
    ffc_391_p_spl_
  );


  buf

  (
    g2264_n_spl_,
    g2264_n
  );


  buf

  (
    g2264_n_spl_0,
    g2264_n_spl_
  );


  buf

  (
    g2267_p_spl_,
    g2267_p
  );


  buf

  (
    g2365_p_spl_,
    g2365_p
  );


  buf

  (
    ffc_395_p_spl_,
    ffc_395_p
  );


  buf

  (
    g1898_n_spl_,
    g1898_n
  );


  buf

  (
    g2268_n_spl_,
    g2268_n
  );


  buf

  (
    ffc_387_p_spl_,
    ffc_387_p
  );


  buf

  (
    g2129_n_spl_,
    g2129_n
  );


  buf

  (
    g2361_n_spl_,
    g2361_n
  );


  buf

  (
    g2362_n_spl_,
    g2362_n
  );


  buf

  (
    g2363_n_spl_,
    g2363_n
  );


  buf

  (
    G92_p_spl_,
    G92_p
  );


  buf

  (
    G124_p_spl_,
    G124_p
  );


  buf

  (
    G124_p_spl_0,
    G124_p_spl_
  );


  buf

  (
    G124_p_spl_1,
    G124_p_spl_
  );


  buf

  (
    G124_n_spl_,
    G124_n
  );


  buf

  (
    G124_n_spl_0,
    G124_n_spl_
  );


  buf

  (
    G94_p_spl_,
    G94_p
  );


  buf

  (
    G107_p_spl_,
    G107_p
  );


  buf

  (
    ffc_401_n_spl_,
    ffc_401_n
  );


  buf

  (
    ffc_401_n_spl_0,
    ffc_401_n_spl_
  );


  buf

  (
    ffc_405_p_spl_,
    ffc_405_p
  );


  buf

  (
    ffc_3_n_spl_,
    ffc_3_n
  );


  buf

  (
    ffc_3_n_spl_0,
    ffc_3_n_spl_
  );


  buf

  (
    ffc_3_n_spl_1,
    ffc_3_n_spl_
  );


  buf

  (
    ffc_359_n_spl_,
    ffc_359_n
  );


  buf

  (
    g1064_n_spl_,
    g1064_n
  );


  buf

  (
    g1102_n_spl_,
    g1102_n
  );


  buf

  (
    g1106_p_spl_,
    g1106_p
  );


  buf

  (
    g1126_p_spl_,
    g1126_p
  );


  buf

  (
    g1127_n_spl_,
    g1127_n
  );


endmodule
