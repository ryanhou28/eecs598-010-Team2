// Benchmark "c3540" written by ABC on Sun Oct 29 19:31:55 2023

module c3540 (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50,
    G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528,
    G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538,
    G3539, G3540  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50;
  output G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528,
    G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538,
    G3539, G3540;
  reg n1743_lo, n1746_lo, n1749_lo, n1752_lo, n1755_lo, n1758_lo, n1761_lo,
    n1764_lo, n1767_lo, n1770_lo, n1773_lo, n1776_lo, n1779_lo, n1782_lo,
    n1785_lo, n1788_lo, n1791_lo, n1794_lo, n1797_lo, n1800_lo, n1803_lo,
    n1806_lo, n1809_lo, n1812_lo, n1815_lo, n1818_lo, n1821_lo, n1824_lo,
    n1827_lo, n1830_lo, n1833_lo, n1836_lo, n1839_lo, n1842_lo, n1845_lo,
    n1848_lo, n1851_lo, n1854_lo, n1857_lo, n1860_lo, n1863_lo, n1866_lo,
    n1869_lo, n1872_lo, n1875_lo, n1878_lo, n1881_lo, n1884_lo, n1887_lo,
    n1890_lo, n1893_lo, n1896_lo, n1899_lo, n1902_lo, n1905_lo, n1908_lo,
    n1911_lo, n1914_lo, n1917_lo, n1920_lo, n1923_lo, n1926_lo, n1929_lo,
    n1932_lo, n1935_lo, n1938_lo, n1941_lo, n1944_lo, n1947_lo, n1950_lo,
    n1953_lo, n1956_lo, n1959_lo, n1962_lo, n1965_lo, n1968_lo, n1971_lo,
    n1974_lo, n1977_lo, n1980_lo, n1983_lo, n1986_lo, n1989_lo, n1992_lo,
    n1995_lo, n1998_lo, n2001_lo, n2004_lo, n2007_lo, n2010_lo, n2013_lo,
    n2016_lo, n2019_lo, n2022_lo, n2025_lo, n2028_lo, n2031_lo, n2034_lo,
    n2037_lo, n2040_lo, n2043_lo, n2046_lo, n2049_lo, n2052_lo, n2055_lo,
    n2058_lo, n2061_lo, n2064_lo, n2067_lo, n2070_lo, n2073_lo, n2076_lo,
    n2079_lo, n2082_lo, n2085_lo, n2088_lo, n2091_lo, n2094_lo, n2097_lo,
    n2100_lo, n2103_lo, n2106_lo, n2109_lo, n2112_lo, n2115_lo, n2118_lo,
    n2121_lo, n2124_lo, n2127_lo, n2130_lo, n2133_lo, n2136_lo, n2139_lo,
    n2142_lo, n2145_lo, n2148_lo, n2151_lo, n2154_lo, n2157_lo, n2160_lo,
    n2163_lo, n2166_lo, n2169_lo, n2172_lo, n2175_lo, n2178_lo, n2181_lo,
    n2184_lo, n2187_lo, n2190_lo, n2193_lo, n2196_lo, n2199_lo, n2202_lo,
    n2205_lo, n2208_lo, n2211_lo, n2214_lo, n2217_lo, n2220_lo, n2223_lo,
    n2226_lo, n2229_lo, n2232_lo, n2235_lo, n2238_lo, n2241_lo, n2244_lo,
    n2247_lo, n2250_lo, n2253_lo, n2256_lo, n2259_lo, n2262_lo, n2265_lo,
    n2268_lo, n2271_lo, n2274_lo, n2277_lo, n2280_lo, n2283_lo, n2286_lo,
    n2289_lo, n2292_lo, n2295_lo, n2298_lo, n2301_lo, n2304_lo, n2307_lo,
    n2310_lo, n2313_lo, n2316_lo, n2319_lo, n2322_lo, n2325_lo, n2328_lo,
    n2331_lo, n2334_lo, n2337_lo, n2340_lo;
  wire new_G353_, new_G363_, new_G368_, new_G377_, new_G381_, new_G384_,
    new_G388_, new_G397_, new_G400_, new_G404_, new_G413_, new_G422_,
    new_G425_, new_G434_, new_G438_, new_G447_, new_G451_, new_G461_,
    new_G466_, new_G467_, new_G470_, new_G477_, new_G480_, new_G484_,
    new_G491_, new_G492_, new_G496_, new_G501_, new_G518_, new_G519_,
    new_G523_, new_G527_, new_G530_, new_G533_, new_G534_, new_G537_,
    new_G540_, new_G543_, new_G546_, new_G549_, new_G552_, new_G556_,
    new_G559_, new_G562_, new_G565_, new_G568_, new_G572_, new_G575_,
    new_G578_, new_G581_, new_G584_, new_G587_, new_G588_, new_G589_,
    new_G590_, new_G593_, new_G594_, new_G611_, new_G612_, new_G613_,
    new_G614_, new_G615_, new_G618_, new_G621_, new_G624_, new_G627_,
    new_G630_, new_G633_, new_G636_, new_G639_, new_G642_, new_G645_,
    new_G648_, new_G651_, new_G654_, new_G657_, new_G660_, new_G663_,
    new_G666_, new_G667_, new_G684_, new_G685_, new_G686_, new_G691_,
    new_G708_, new_G713_, new_G714_, new_G715_, new_G716_, new_G717_,
    new_G718_, new_G719_, new_G720_, new_G721_, new_G722_, new_G723_,
    new_G724_, new_G725_, new_G726_, new_G727_, new_G730_, new_G731_,
    new_G734_, new_G735_, new_G736_, new_G739_, new_G742_, new_G745_,
    new_G749_, new_G753_, new_G762_, new_G769_, new_G772_, new_G775_,
    new_G778_, new_G781_, new_G784_, new_G785_, new_G786_, new_G787_,
    new_G790_, new_G791_, new_G792_, new_G793_, new_G794_, new_G795_,
    new_G796_, new_G797_, new_G798_, new_G799_, new_G800_, new_G805_,
    new_G810_, new_G813_, new_G816_, new_G831_, new_G848_, new_G849_,
    new_G850_, new_G851_, new_G852_, new_G853_, new_G854_, new_G855_,
    new_G856_, new_G873_, new_G874_, new_G875_, new_G882_, new_G883_,
    new_G884_, new_G887_, new_G890_, new_G891_, new_G892_, new_G893_,
    new_G894_, new_G897_, new_G898_, new_G901_, new_G904_, new_G907_,
    new_G910_, new_G913_, new_G916_, new_G919_, new_G922_, new_G925_,
    new_G928_, new_G929_, new_G930_, new_G931_, new_G932_, new_G933_,
    new_G934_, new_G935_, new_G939_, new_G956_, new_G957_, new_G958_,
    new_G959_, new_G960_, new_G961_, new_G962_, new_G963_, new_G964_,
    new_G965_, new_G966_, new_G967_, new_G968_, new_G969_, new_G970_,
    new_G971_, new_G972_, new_G973_, new_G974_, new_G975_, new_G976_,
    new_G977_, new_G978_, new_G979_, new_G980_, new_G981_, new_G982_,
    new_G983_, new_G984_, new_G985_, new_G986_, new_G989_, new_G992_,
    new_G993_, new_G994_, new_G995_, new_G996_, new_G997_, new_G998_,
    new_G999_, new_G1000_, new_G1001_, new_G1002_, new_G1003_, new_G1004_,
    new_G1005_, new_G1008_, new_G1011_, new_G1012_, new_G1015_, new_G1016_,
    new_G1017_, new_G1018_, new_G1019_, new_G1020_, new_G1021_, new_G1022_,
    new_G1023_, new_G1024_, new_G1025_, new_G1034_, new_G1043_, new_G1048_,
    new_G1051_, new_G1052_, new_G1053_, new_G1054_, new_G1055_, new_G1056_,
    new_G1057_, new_G1058_, new_G1059_, new_G1060_, new_G1061_, new_G1062_,
    new_G1063_, new_G1064_, new_G1065_, new_G1066_, new_G1067_, new_G1068_,
    new_G1069_, new_G1070_, new_G1071_, new_G1072_, new_G1073_, new_G1074_,
    new_G1077_, new_G1080_, new_G1083_, new_G1086_, new_G1089_, new_G1092_,
    new_G1095_, new_G1104_, new_G1113_, new_G1114_, new_G1115_, new_G1116_,
    new_G1117_, new_G1118_, new_G1119_, new_G1120_, new_G1121_, new_G1122_,
    new_G1123_, new_G1124_, new_G1125_, new_G1126_, new_G1127_, new_G1128_,
    new_G1129_, new_G1130_, new_G1131_, new_G1132_, new_G1133_, new_G1134_,
    new_G1135_, new_G1136_, new_G1137_, new_G1140_, new_G1141_, new_G1142_,
    new_G1145_, new_G1146_, new_G1147_, new_G1150_, new_G1151_, new_G1152_,
    new_G1155_, new_G1156_, new_G1157_, new_G1160_, new_G1161_, new_G1162_,
    new_G1165_, new_G1166_, new_G1167_, new_G1170_, new_G1171_, new_G1172_,
    new_G1175_, new_G1176_, new_G1179_, new_G1180_, new_G1184_, new_G1189_,
    new_G1193_, new_G1197_, new_G1200_, new_G1203_, new_G1206_, new_G1207_,
    new_G1208_, new_G1209_, new_G1210_, new_G1211_, new_G1212_, new_G1213_,
    new_G1214_, new_G1215_, new_G1216_, new_G1217_, new_G1218_, new_G1219_,
    new_G1222_, new_G1223_, new_G1224_, new_G1225_, new_G1226_, new_G1227_,
    new_G1228_, new_G1229_, new_G1230_, new_G1231_, new_G1232_, new_G1233_,
    new_G1234_, new_G1235_, new_G1236_, new_G1237_, new_G1238_, new_G1239_,
    new_G1240_, new_G1241_, new_G1242_, new_G1243_, new_G1244_, new_G1249_,
    new_G1258_, new_G1263_, new_G1272_, new_G1275_, new_G1278_, new_G1281_,
    new_G1284_, new_G1287_, new_G1290_, new_G1293_, new_G1296_, new_G1297_,
    new_G1298_, new_G1299_, new_G1300_, new_G1301_, new_G1302_, new_G1303_,
    new_G1304_, new_G1305_, new_G1306_, new_G1307_, new_G1308_, new_G1309_,
    new_G1310_, new_G1311_, new_G1312_, new_G1313_, new_G1314_, new_G1315_,
    new_G1316_, new_G1317_, new_G1318_, new_G1319_, new_G1320_, new_G1321_,
    new_G1322_, new_G1323_, new_G1324_, new_G1325_, new_G1326_, new_G1327_,
    new_G1328_, new_G1345_, new_G1348_, new_G1349_, new_G1350_, new_G1351_,
    new_G1352_, new_G1353_, new_G1354_, new_G1357_, new_G1360_, new_G1363_,
    new_G1366_, new_G1369_, new_G1372_, new_G1375_, new_G1378_, new_G1379_,
    new_G1380_, new_G1381_, new_G1390_, new_G1399_, new_G1400_, new_G1401_,
    new_G1402_, new_G1403_, new_G1404_, new_G1405_, new_G1406_, new_G1407_,
    new_G1408_, new_G1409_, new_G1410_, new_G1411_, new_G1412_, new_G1413_,
    new_G1414_, new_G1415_, new_G1418_, new_G1421_, new_G1424_, new_G1427_,
    new_G1430_, new_G1433_, new_G1436_, new_G1439_, new_G1442_, new_G1445_,
    new_G1448_, new_G1451_, new_G1454_, new_G1457_, new_G1460_, new_G1463_,
    new_G1466_, new_G1467_, new_G1468_, new_G1469_, new_G1470_, new_G1471_,
    new_G1472_, new_G1473_, new_G1474_, new_G1475_, new_G1476_, new_G1477_,
    new_G1478_, new_G1479_, new_G1482_, new_G1485_, new_G1486_, new_G1487_,
    new_G1488_, new_G1489_, new_G1490_, new_G1491_, new_G1492_, new_G1493_,
    new_G1494_, new_G1495_, new_G1496_, new_G1497_, new_G1498_, new_G1499_,
    new_G1500_, new_G1501_, new_G1502_, new_G1503_, new_G1504_, new_G1505_,
    new_G1506_, new_G1507_, new_G1508_, new_G1509_, new_G1510_, new_G1511_,
    new_G1512_, new_G1513_, new_G1514_, new_G1517_, new_G1518_, new_G1519_,
    new_G1520_, new_G1521_, new_G1522_, new_G1523_, new_G1524_, new_G1527_,
    new_G1528_, new_G1529_, new_G1538_, new_G1547_, new_G1556_, new_G1565_,
    new_G1574_, new_G1583_, new_G1592_, new_G1601_, new_G1610_, new_G1619_,
    new_G1628_, new_G1637_, new_G1646_, new_G1655_, new_G1664_, new_G1673_,
    new_G1674_, new_G1675_, new_G1676_, new_G1677_, new_G1678_, new_G1679_,
    new_G1680_, new_G1681_, new_G1682_, new_G1683_, new_G1684_, new_G1685_,
    new_G1686_, new_G1687_, new_G1688_, new_G1689_, new_G1693_, new_G1697_,
    new_G1700_, new_G1703_, new_G1707_, new_G1711_, new_G1714_, new_G1718_,
    new_G1722_, new_G1725_, new_G1729_, new_G1733_, new_G1738_, new_G1743_,
    new_G1747_, new_G1751_, new_G1756_, new_G1760_, new_G1764_, new_G1769_,
    new_G1770_, new_G1771_, new_G1772_, new_G1773_, new_G1774_, new_G1775_,
    new_G1776_, new_G1777_, new_G1778_, new_G1779_, new_G1780_, new_G1781_,
    new_G1782_, new_G1783_, new_G1784_, new_G1785_, new_G1786_, new_G1787_,
    new_G1788_, new_G1789_, new_G1790_, new_G1791_, new_G1792_, new_G1793_,
    new_G1794_, new_G1795_, new_G1796_, new_G1799_, new_G1802_, new_G1805_,
    new_G1806_, new_G1807_, new_G1808_, new_G1809_, new_G1810_, new_G1811_,
    new_G1812_, new_G1813_, new_G1816_, new_G1819_, new_G1823_, new_G1826_,
    new_G1827_, new_G1828_, new_G1829_, new_G1830_, new_G1831_, new_G1832_,
    new_G1833_, new_G1834_, new_G1835_, new_G1836_, new_G1837_, new_G1838_,
    new_G1839_, new_G1840_, new_G1841_, new_G1842_, new_G1843_, new_G1844_,
    new_G1845_, new_G1846_, new_G1847_, new_G1848_, new_G1849_, new_G1850_,
    new_G1851_, new_G1852_, new_G1853_, new_G1854_, new_G1855_, new_G1856_,
    new_G1857_, new_G1858_, new_G1859_, new_G1860_, new_G1861_, new_G1862_,
    new_G1863_, new_G1864_, new_G1865_, new_G1866_, new_G1867_, new_G1868_,
    new_G1869_, new_G1870_, new_G1871_, new_G1872_, new_G1873_, new_G1874_,
    new_G1875_, new_G1876_, new_G1877_, new_G1878_, new_G1879_, new_G1880_,
    new_G1881_, new_G1882_, new_G1883_, new_G1884_, new_G1885_, new_G1886_,
    new_G1887_, new_G1888_, new_G1889_, new_G1890_, new_G1891_, new_G1892_,
    new_G1893_, new_G1894_, new_G1895_, new_G1896_, new_G1897_, new_G1898_,
    new_G1899_, new_G1900_, new_G1901_, new_G1902_, new_G1903_, new_G1904_,
    new_G1905_, new_G1906_, new_G1907_, new_G1908_, new_G1909_, new_G1910_,
    new_G1911_, new_G1912_, new_G1913_, new_G1914_, new_G1915_, new_G1916_,
    new_G1917_, new_G1918_, new_G1919_, new_G1920_, new_G1921_, new_G1922_,
    new_G1923_, new_G1924_, new_G1925_, new_G1926_, new_G1927_, new_G1928_,
    new_G1929_, new_G1930_, new_G1931_, new_G1932_, new_G1933_, new_G1934_,
    new_G1935_, new_G1936_, new_G1937_, new_G1938_, new_G1939_, new_G1940_,
    new_G1941_, new_G1942_, new_G1943_, new_G1944_, new_G1945_, new_G1946_,
    new_G1947_, new_G1948_, new_G1949_, new_G1950_, new_G1951_, new_G1952_,
    new_G1953_, new_G1954_, new_G1955_, new_G1958_, new_G1961_, new_G1962_,
    new_G1965_, new_G1968_, new_G1971_, new_G1974_, new_G1977_, new_G1978_,
    new_G1981_, new_G1984_, new_G1985_, new_G1988_, new_G1991_, new_G1992_,
    new_G1995_, new_G1998_, new_G2001_, new_G2004_, new_G2007_, new_G2008_,
    new_G2011_, new_G2014_, new_G2015_, new_G2018_, new_G2021_, new_G2024_,
    new_G2027_, new_G2030_, new_G2033_, new_G2034_, new_G2035_, new_G2036_,
    new_G2037_, new_G2038_, new_G2039_, new_G2040_, new_G2041_, new_G2042_,
    new_G2043_, new_G2044_, new_G2045_, new_G2046_, new_G2047_, new_G2048_,
    new_G2049_, new_G2050_, new_G2051_, new_G2052_, new_G2053_, new_G2054_,
    new_G2055_, new_G2056_, new_G2057_, new_G2058_, new_G2059_, new_G2060_,
    new_G2061_, new_G2062_, new_G2063_, new_G2064_, new_G2065_, new_G2066_,
    new_G2067_, new_G2068_, new_G2069_, new_G2070_, new_G2071_, new_G2072_,
    new_G2073_, new_G2074_, new_G2075_, new_G2076_, new_G2077_, new_G2078_,
    new_G2079_, new_G2080_, new_G2081_, new_G2082_, new_G2083_, new_G2084_,
    new_G2085_, new_G2086_, new_G2087_, new_G2088_, new_G2089_, new_G2090_,
    new_G2091_, new_G2092_, new_G2093_, new_G2094_, new_G2095_, new_G2096_,
    new_G2097_, new_G2098_, new_G2099_, new_G2100_, new_G2101_, new_G2102_,
    new_G2103_, new_G2104_, new_G2105_, new_G2106_, new_G2107_, new_G2108_,
    new_G2109_, new_G2110_, new_G2111_, new_G2112_, new_G2113_, new_G2114_,
    new_G2115_, new_G2116_, new_G2117_, new_G2118_, new_G2119_, new_G2120_,
    new_G2121_, new_G2122_, new_G2123_, new_G2124_, new_G2125_, new_G2126_,
    new_G2127_, new_G2128_, new_G2129_, new_G2130_, new_G2131_, new_G2132_,
    new_G2133_, new_G2134_, new_G2135_, new_G2136_, new_G2137_, new_G2138_,
    new_G2139_, new_G2140_, new_G2141_, new_G2142_, new_G2143_, new_G2144_,
    new_G2145_, new_G2146_, new_G2147_, new_G2148_, new_G2149_, new_G2150_,
    new_G2151_, new_G2152_, new_G2153_, new_G2154_, new_G2155_, new_G2156_,
    new_G2157_, new_G2158_, new_G2159_, new_G2160_, new_G2161_, new_G2162_,
    new_G2163_, new_G2164_, new_G2165_, new_G2166_, new_G2167_, new_G2168_,
    new_G2169_, new_G2172_, new_G2173_, new_G2174_, new_G2175_, new_G2176_,
    new_G2177_, new_G2178_, new_G2179_, new_G2180_, new_G2181_, new_G2182_,
    new_G2183_, new_G2184_, new_G2185_, new_G2186_, new_G2187_, new_G2188_,
    new_G2189_, new_G2190_, new_G2191_, new_G2192_, new_G2195_, new_G2198_,
    new_G2199_, new_G2200_, new_G2204_, new_G2208_, new_G2211_, new_G2214_,
    new_G2215_, new_G2216_, new_G2219_, new_G2222_, new_G2223_, new_G2224_,
    new_G2227_, new_G2230_, new_G2231_, new_G2232_, new_G2236_, new_G2240_,
    new_G2243_, new_G2246_, new_G2247_, new_G2248_, new_G2251_, new_G2254_,
    new_G2255_, new_G2256_, new_G2257_, new_G2260_, new_G2263_, new_G2266_,
    new_G2269_, new_G2272_, new_G2275_, new_G2278_, new_G2281_, new_G2284_,
    new_G2287_, new_G2290_, new_G2293_, new_G2296_, new_G2299_, new_G2302_,
    new_G2305_, new_G2308_, new_G2311_, new_G2312_, new_G2313_, new_G2314_,
    new_G2315_, new_G2316_, new_G2317_, new_G2318_, new_G2319_, new_G2320_,
    new_G2321_, new_G2322_, new_G2323_, new_G2324_, new_G2325_, new_G2326_,
    new_G2327_, new_G2328_, new_G2329_, new_G2330_, new_G2331_, new_G2332_,
    new_G2333_, new_G2334_, new_G2335_, new_G2336_, new_G2337_, new_G2338_,
    new_G2339_, new_G2340_, new_G2341_, new_G2342_, new_G2343_, new_G2344_,
    new_G2345_, new_G2346_, new_G2347_, new_G2348_, new_G2349_, new_G2350_,
    new_G2351_, new_G2352_, new_G2353_, new_G2354_, new_G2355_, new_G2356_,
    new_G2359_, new_G2362_, new_G2363_, new_G2364_, new_G2365_, new_G2368_,
    new_G2369_, new_G2372_, new_G2373_, new_G2374_, new_G2375_, new_G2378_,
    new_G2381_, new_G2382_, new_G2383_, new_G2384_, new_G2387_, new_G2388_,
    new_G2391_, new_G2392_, new_G2393_, new_G2396_, new_G2397_, new_G2398_,
    new_G2399_, new_G2400_, new_G2401_, new_G2404_, new_G2405_, new_G2406_,
    new_G2407_, new_G2408_, new_G2411_, new_G2414_, new_G2415_, new_G2416_,
    new_G2417_, new_G2418_, new_G2419_, new_G2420_, new_G2421_, new_G2422_,
    new_G2423_, new_G2424_, new_G2425_, new_G2426_, new_G2427_, new_G2428_,
    new_G2429_, new_G2430_, new_G2436_, new_G2437_, new_G2441_, new_G2444_,
    new_G2450_, new_G2451_, new_G2455_, new_G2458_, new_G2459_, new_G2460_,
    new_G2461_, new_G2462_, new_G2463_, new_G2464_, new_G2465_, new_G2466_,
    new_G2467_, new_G2468_, new_G2471_, new_G2472_, new_G2475_, new_G2476_,
    new_G2479_, new_G2482_, new_G2485_, new_G2488_, new_G2491_, new_G2494_,
    new_G2497_, new_G2500_, new_G2501_, new_G2502_, new_G2507_, new_G2512_,
    new_G2515_, new_G2518_, new_G2521_, new_G2524_, new_G2527_, new_G2530_,
    new_G2531_, new_G2532_, new_G2533_, new_G2534_, new_G2535_, new_G2536_,
    new_G2537_, new_G2538_, new_G2539_, new_G2542_, new_G2543_, new_G2546_,
    new_G2547_, new_G2550_, new_G2551_, new_G2552_, new_G2556_, new_G2557_,
    new_G2558_, new_G2561_, new_G2562_, new_G2563_, new_G2566_, new_G2569_,
    new_G2570_, new_G2571_, new_G2574_, new_G2577_, new_G2580_, new_G2583_,
    new_G2586_, new_G2589_, new_G2592_, new_G2595_, new_G2598_, new_G2601_,
    new_G2604_, new_G2607_, new_G2610_, new_G2613_, new_G2614_, new_G2615_,
    new_G2616_, new_G2617_, new_G2618_, new_G2619_, new_G2620_, new_G2623_,
    new_G2624_, new_G2625_, new_G2626_, new_G2627_, new_G2628_, new_G2629_,
    new_G2630_, new_G2631_, new_G2632_, new_G2633_, new_G2634_, new_G2635_,
    new_G2636_, new_G2637_, new_G2638_, new_G2639_, new_G2640_, new_G2643_,
    new_G2646_, new_G2647_, new_G2648_, new_G2651_, new_G2654_, new_G2655_,
    new_G2656_, new_G2657_, new_G2658_, new_G2659_, new_G2660_, new_G2661_,
    new_G2662_, new_G2663_, new_G2664_, new_G2665_, new_G2666_, new_G2669_,
    new_G2673_, new_G2674_, new_G2675_, new_G2676_, new_G2677_, new_G2678_,
    new_G2679_, new_G2680_, new_G2681_, new_G2682_, new_G2683_, new_G2684_,
    new_G2685_, new_G2686_, new_G2687_, new_G2690_, new_G2693_, new_G2694_,
    new_G2697_, new_G2698_, new_G2699_, new_G2705_, new_G2708_, new_G2711_,
    new_G2712_, new_G2713_, new_G2714_, new_G2715_, new_G2716_, new_G2717_,
    new_G2718_, new_G2719_, new_G2720_, new_G2721_, new_G2728_, new_G2733_,
    new_G2736_, new_G2739_, new_G2740_, new_G2741_, new_G2742_, new_G2743_,
    new_G2744_, new_G2745_, new_G2746_, new_G2747_, new_G2750_, new_G2753_,
    new_G2759_, new_G2763_, new_G2768_, new_G2773_, new_G2778_, new_G2779_,
    new_G2780_, new_G2781_, new_G2784_, new_G2787_, new_G2788_, new_G2789_,
    new_G2790_, new_G2791_, new_G2792_, new_G2793_, new_G2794_, new_G2795_,
    new_G2796_, new_G2799_, new_G2803_, new_G2804_, new_G2805_, new_G2808_,
    new_G2809_, new_G2810_, new_G2811_, new_G2816_, new_G2820_, new_G2821_,
    new_G2822_, new_G2823_, new_G2826_, new_G2827_, new_G2828_, new_G2829_,
    new_G2830_, new_G2831_, new_G2832_, new_G2833_, new_G2836_, new_G2839_,
    new_G2842_, new_G2845_, new_G2848_, new_G2851_, new_G2854_, new_G2857_,
    new_G2860_, new_G2863_, new_G2866_, new_G2869_, new_G2872_, new_G2875_,
    new_G2876_, new_G2877_, new_G2880_, new_G2883_, new_G2884_, new_G2887_,
    new_G2890_, new_G2893_, new_G2896_, new_G2899_, new_G2902_, new_G2905_,
    new_G2906_, new_G2909_, new_G2910_, new_G2911_, new_G2912_, new_G2913_,
    new_G2916_, new_G2917_, new_G2918_, new_G2919_, new_G2920_, new_G2923_,
    new_G2926_, new_G2929_, new_G2932_, new_G2935_, new_G2936_, new_G2937_,
    new_G2938_, new_G2939_, new_G2942_, new_G2943_, new_G2944_, new_G2947_,
    new_G2950_, new_G2951_, new_G2952_, new_G2953_, new_G2954_, new_G2955_,
    new_G2956_, new_G2957_, new_G2958_, new_G2959_, new_G2960_, new_G2961_,
    new_G2962_, new_G2965_, new_G2968_, new_G2971_, new_G2974_, new_G2975_,
    new_G2978_, new_G2979_, new_G2980_, new_G2981_, new_G2984_, new_G2985_,
    new_G2986_, new_G2990_, new_G2991_, new_G2994_, new_G2995_, new_G2996_,
    new_G2999_, new_G3002_, new_G3005_, new_G3006_, new_G3007_, new_G3010_,
    new_G3011_, new_G3012_, new_G3015_, new_G3016_, new_G3017_, new_G3018_,
    new_G3021_, new_G3024_, new_G3027_, new_G3030_, new_G3031_, new_G3032_,
    new_G3033_, new_G3034_, new_G3035_, new_G3036_, new_G3037_, new_G3038_,
    new_G3039_, new_G3042_, new_G3045_, new_G3048_, new_G3051_, new_G3054_,
    new_G3057_, new_G3058_, new_G3059_, new_G3060_, new_G3061_, new_G3062_,
    new_G3063_, new_G3064_, new_G3065_, new_G3066_, new_G3067_, new_G3068_,
    new_G3069_, new_G3072_, new_G3075_, new_G3078_, new_G3081_, new_G3082_,
    new_G3083_, new_G3084_, new_G3085_, new_G3086_, new_G3089_, new_G3090_,
    new_G3094_, new_G3095_, new_G3099_, new_G3100_, new_G3103_, new_G3106_,
    new_G3107_, new_G3110_, new_G3114_, new_G3115_, new_G3116_, new_G3117_,
    new_G3118_, new_G3119_, new_G3120_, new_G3121_, new_G3122_, new_G3126_,
    new_G3129_, new_G3132_, new_G3135_, new_G3136_, new_G3137_, new_G3138_,
    new_G3139_, new_G3140_, new_G3143_, new_G3146_, new_G3149_, new_G3152_,
    new_G3155_, new_G3158_, new_G3159_, new_G3160_, new_G3164_, new_G3165_,
    new_G3168_, new_G3169_, new_G3170_, new_G3171_, new_G3174_, new_G3177_,
    new_G3180_, new_G3183_, new_G3186_, new_G3189_, new_G3190_, new_G3191_,
    new_G3192_, new_G3193_, new_G3194_, new_G3195_, new_G3199_, new_G3202_,
    new_G3203_, new_G3206_, new_G3207_, new_G3208_, new_G3209_, new_G3210_,
    new_G3211_, new_G3212_, new_G3213_, new_G3214_, new_G3215_, new_G3216_,
    new_G3217_, new_G3220_, new_G3223_, new_G3226_, new_G3227_, new_G3230_,
    new_G3231_, new_G3232_, new_G3233_, new_G3234_, new_G3235_, new_G3236_,
    new_G3237_, new_G3240_, new_G3243_, new_G3246_, new_G3247_, new_G3248_,
    new_G3249_, new_G3250_, new_G3251_, new_G3254_, new_G3257_, new_G3258_,
    new_G3259_, new_G3260_, new_G3261_, new_G3262_, new_G3265_, new_G3266_,
    new_G3267_, new_G3268_, new_G3269_, new_G3270_, new_G3271_, new_G3272_,
    new_G3275_, new_G3278_, new_G3281_, new_G3284_, new_G3287_, new_G3288_,
    new_G3291_, new_G3294_, new_G3297_, new_G3300_, new_G3301_, new_G3302_,
    new_G3305_, new_G3308_, new_G3311_, new_G3312_, new_G3317_, new_G3320_,
    new_G3323_, new_G3326_, new_G3329_, new_G3332_, new_G3337_, new_G3340_,
    new_G3341_, new_G3342_, new_G3343_, new_G3344_, new_G3345_, new_G3346_,
    new_G3347_, new_G3350_, new_G3353_, new_G3356_, new_G3359_, new_G3360_,
    new_G3363_, new_G3366_, new_G3367_, new_G3370_, new_G3373_, new_G3376_,
    new_G3379_, new_G3380_, new_G3383_, new_G3386_, new_G3387_, new_G3388_,
    new_G3391_, new_G3394_, new_G3395_, new_G3396_, new_G3399_, new_G3402_,
    new_G3403_, new_G3404_, new_G3405_, new_G3406_, new_G3407_, new_G3408_,
    new_G3409_, new_G3412_, new_G3415_, new_G3416_, new_G3417_, new_G3418_,
    new_G3419_, new_G3420_, new_G3421_, new_G3422_, new_G3423_, new_G3424_,
    new_G3425_, new_G3428_, new_G3429_, new_G3430_, new_G3431_, new_G3432_,
    new_G3436_, new_G3437_, new_G3438_, new_G3439_, new_G3440_, new_G3441_,
    new_G3444_, new_G3445_, new_G3448_, new_G3449_, new_G3452_, new_G3453_,
    new_G3456_, new_G3459_, new_G3460_, new_G3461_, new_G3464_, new_G3465_,
    new_G3466_, new_G3467_, new_G3468_, new_G3471_, new_G3474_, new_G3475_,
    new_G3478_, new_G3481_, new_G3484_, new_G3487_, new_G3488_, new_G3489_,
    new_G3490_, new_G3491_, new_G3494_, new_G3497_, new_G3500_, new_G3503_,
    new_G3504_, new_G3505_, new_G3506_, new_G3507_, new_G3508_, new_G3509_,
    new_G3510_, new_G3511_, new_G3512_, new_G3513_, new_G3514_, new_G3515_,
    new_G3516_, new_G3517_, new_G3518_, n1743_li, n1746_li, n1749_li,
    n1752_li, n1755_li, n1758_li, n1761_li, n1764_li, n1767_li, n1770_li,
    n1773_li, n1776_li, n1779_li, n1782_li, n1785_li, n1788_li, n1791_li,
    n1794_li, n1797_li, n1800_li, n1803_li, n1806_li, n1809_li, n1812_li,
    n1815_li, n1818_li, n1821_li, n1824_li, n1827_li, n1830_li, n1833_li,
    n1836_li, n1839_li, n1842_li, n1845_li, n1848_li, n1851_li, n1854_li,
    n1857_li, n1860_li, n1863_li, n1866_li, n1869_li, n1872_li, n1875_li,
    n1878_li, n1881_li, n1884_li, n1887_li, n1890_li, n1893_li, n1896_li,
    n1899_li, n1902_li, n1905_li, n1908_li, n1911_li, n1914_li, n1917_li,
    n1920_li, n1923_li, n1926_li, n1929_li, n1932_li, n1935_li, n1938_li,
    n1941_li, n1944_li, n1947_li, n1950_li, n1953_li, n1956_li, n1959_li,
    n1962_li, n1965_li, n1968_li, n1971_li, n1974_li, n1977_li, n1980_li,
    n1983_li, n1986_li, n1989_li, n1992_li, n1995_li, n1998_li, n2001_li,
    n2004_li, n2007_li, n2010_li, n2013_li, n2016_li, n2019_li, n2022_li,
    n2025_li, n2028_li, n2031_li, n2034_li, n2037_li, n2040_li, n2043_li,
    n2046_li, n2049_li, n2052_li, n2055_li, n2058_li, n2061_li, n2064_li,
    n2067_li, n2070_li, n2073_li, n2076_li, n2079_li, n2082_li, n2085_li,
    n2088_li, n2091_li, n2094_li, n2097_li, n2100_li, n2103_li, n2106_li,
    n2109_li, n2112_li, n2115_li, n2118_li, n2121_li, n2124_li, n2127_li,
    n2130_li, n2133_li, n2136_li, n2139_li, n2142_li, n2145_li, n2148_li,
    n2151_li, n2154_li, n2157_li, n2160_li, n2163_li, n2166_li, n2169_li,
    n2172_li, n2175_li, n2178_li, n2181_li, n2184_li, n2187_li, n2190_li,
    n2193_li, n2196_li, n2199_li, n2202_li, n2205_li, n2208_li, n2211_li,
    n2214_li, n2217_li, n2220_li, n2223_li, n2226_li, n2229_li, n2232_li,
    n2235_li, n2238_li, n2241_li, n2244_li, n2247_li, n2250_li, n2253_li,
    n2256_li, n2259_li, n2262_li, n2265_li, n2268_li, n2271_li, n2274_li,
    n2277_li, n2280_li, n2283_li, n2286_li, n2289_li, n2292_li, n2295_li,
    n2298_li, n2301_li, n2304_li, n2307_li, n2310_li, n2313_li, n2316_li,
    n2319_li, n2322_li, n2325_li, n2328_li, n2331_li, n2334_li, n2337_li,
    n2340_li;
  assign new_G353_ = ~n1824_lo;
  assign new_G363_ = ~n1824_lo;
  assign new_G368_ = ~n1836_lo;
  assign new_G377_ = ~n1836_lo;
  assign new_G381_ = ~n1848_lo;
  assign new_G384_ = ~n1848_lo;
  assign new_G388_ = ~n1848_lo;
  assign new_G397_ = ~n1860_lo;
  assign new_G400_ = ~n1860_lo;
  assign new_G404_ = ~n1860_lo;
  assign new_G413_ = ~n1872_lo;
  assign new_G422_ = ~n1872_lo;
  assign new_G425_ = ~n1884_lo;
  assign new_G434_ = ~n1884_lo;
  assign new_G438_ = ~n1896_lo;
  assign new_G447_ = ~n1896_lo;
  assign new_G451_ = ~n1908_lo;
  assign new_G461_ = ~n1908_lo;
  assign new_G466_ = n2160_lo | n2172_lo;
  assign new_G467_ = ~n1752_lo;
  assign new_G470_ = ~n1752_lo;
  assign new_G477_ = ~n1752_lo;
  assign new_G480_ = ~n1764_lo;
  assign new_G484_ = ~n1764_lo;
  assign new_G491_ = n1764_lo & n1776_lo;
  assign new_G492_ = ~n1776_lo;
  assign new_G496_ = ~n1776_lo;
  assign new_G501_ = ~n1776_lo;
  assign new_G518_ = ~n1788_lo;
  assign new_G519_ = ~n1788_lo;
  assign new_G523_ = ~n1788_lo;
  assign new_G527_ = n1788_lo & n1800_lo;
  assign new_G530_ = ~n1800_lo;
  assign new_G533_ = n1800_lo | n1812_lo;
  assign new_G534_ = ~n1812_lo;
  assign new_G537_ = ~n1812_lo;
  assign new_G540_ = ~n1824_lo;
  assign new_G543_ = ~n1836_lo;
  assign new_G546_ = ~n1836_lo;
  assign new_G549_ = ~n1848_lo;
  assign new_G552_ = ~n1848_lo;
  assign new_G556_ = ~n1872_lo;
  assign new_G559_ = ~n1872_lo;
  assign new_G562_ = ~n1884_lo;
  assign new_G565_ = ~n1884_lo;
  assign new_G568_ = ~n1896_lo;
  assign new_G572_ = ~n1752_lo;
  assign new_G575_ = ~n1848_lo;
  assign new_G578_ = ~n1896_lo;
  assign new_G581_ = ~n1776_lo;
  assign new_G584_ = ~n2040_lo;
  assign new_G587_ = ~n2052_lo;
  assign new_G588_ = n1776_lo & n2052_lo;
  assign new_G589_ = ~n1776_lo | ~n2052_lo;
  assign new_G590_ = n1776_lo & n2028_lo;
  assign new_G593_ = ~n1776_lo;
  assign new_G594_ = n2328_lo | n1788_lo;
  assign new_G611_ = ~n1752_lo | ~n1764_lo;
  assign new_G612_ = ~n1752_lo | ~n1776_lo | ~n1788_lo;
  assign new_G613_ = ~n1776_lo;
  assign new_G614_ = ~n1788_lo;
  assign new_G615_ = ~n2028_lo;
  assign new_G618_ = ~n2064_lo;
  assign new_G621_ = ~n2316_lo;
  assign new_G624_ = ~n2100_lo;
  assign new_G627_ = ~n2112_lo;
  assign new_G630_ = ~n2124_lo;
  assign new_G633_ = ~n2136_lo;
  assign new_G636_ = ~n2148_lo;
  assign new_G639_ = ~n2160_lo;
  assign new_G642_ = ~n2172_lo;
  assign new_G645_ = ~n2184_lo;
  assign new_G648_ = ~n1824_lo;
  assign new_G651_ = ~n1836_lo;
  assign new_G654_ = ~n1836_lo;
  assign new_G657_ = ~n1884_lo;
  assign new_G660_ = ~n1884_lo;
  assign new_G663_ = ~n2304_lo;
  assign new_G666_ = n2148_lo & new_G466_;
  assign new_G667_ = new_G518_ | n1776_lo;
  assign new_G684_ = new_G593_ | n2016_lo;
  assign new_G685_ = ~new_G491_;
  assign new_G686_ = new_G613_ | n1752_lo;
  assign new_G691_ = new_G611_ & new_G612_;
  assign new_G708_ = new_G614_ | n1752_lo;
  assign new_G713_ = new_G540_ & new_G546_ & new_G552_;
  assign new_G714_ = ~n2100_lo | ~new_G353_;
  assign new_G715_ = ~n2112_lo | ~new_G368_;
  assign new_G716_ = ~n2124_lo | ~new_G388_;
  assign new_G717_ = ~n2136_lo | ~new_G404_;
  assign new_G718_ = ~n2148_lo | ~new_G413_;
  assign new_G719_ = ~n2160_lo | ~new_G425_;
  assign new_G720_ = ~n2172_lo | ~new_G438_;
  assign new_G721_ = ~n2184_lo | ~new_G451_;
  assign new_G722_ = ~new_G624_;
  assign new_G723_ = ~new_G627_;
  assign new_G724_ = ~new_G630_;
  assign new_G725_ = ~new_G633_;
  assign new_G726_ = ~new_G377_ | ~new_G384_;
  assign new_G727_ = ~new_G434_ | ~new_G447_;
  assign new_G730_ = ~new_G381_ | ~new_G397_;
  assign new_G731_ = ~new_G363_;
  assign new_G734_ = ~new_G651_;
  assign new_G735_ = ~new_G657_;
  assign new_G736_ = ~new_G537_;
  assign new_G739_ = ~new_G537_;
  assign new_G742_ = ~new_G480_;
  assign new_G745_ = ~new_G523_;
  assign new_G749_ = ~new_G530_;
  assign new_G753_ = new_G477_ & new_G533_;
  assign new_G762_ = new_G477_ & new_G534_ & new_G530_;
  assign new_G769_ = new_G467_ & new_G534_;
  assign new_G772_ = new_G470_ & new_G484_ & new_G496_;
  assign new_G775_ = ~new_G470_ | ~new_G484_ | ~new_G496_;
  assign new_G778_ = ~new_G470_ | ~new_G484_;
  assign new_G781_ = ~new_G572_;
  assign new_G784_ = ~new_G480_ | ~new_G492_ | ~n1812_lo;
  assign new_G785_ = ~new_G540_ | ~new_G546_ | ~new_G552_;
  assign new_G786_ = ~new_G654_;
  assign new_G787_ = new_G559_ & new_G565_ & new_G568_;
  assign new_G790_ = ~new_G559_ | ~new_G565_ | ~new_G568_;
  assign new_G791_ = ~new_G660_;
  assign new_G792_ = ~new_G501_;
  assign new_G793_ = ~new_G501_;
  assign new_G794_ = ~new_G501_;
  assign new_G795_ = ~new_G501_;
  assign new_G796_ = ~new_G501_;
  assign new_G797_ = ~new_G501_;
  assign new_G798_ = ~new_G501_;
  assign new_G799_ = ~new_G501_;
  assign new_G800_ = new_G581_ | new_G584_;
  assign new_G805_ = ~new_G581_ & ~new_G584_;
  assign new_G810_ = ~new_G590_;
  assign new_G813_ = ~new_G590_;
  assign new_G816_ = ~new_G519_;
  assign new_G831_ = ~new_G523_;
  assign new_G848_ = ~new_G594_;
  assign new_G849_ = ~new_G594_;
  assign new_G850_ = ~new_G594_;
  assign new_G851_ = ~new_G594_;
  assign new_G852_ = ~new_G594_;
  assign new_G853_ = ~new_G594_;
  assign new_G854_ = ~new_G594_;
  assign new_G855_ = ~new_G594_;
  assign new_G856_ = n1752_lo | new_G685_;
  assign new_G873_ = ~new_G527_;
  assign new_G874_ = ~new_G527_;
  assign new_G875_ = new_G467_ & new_G480_ & new_G492_;
  assign new_G882_ = ~new_G615_;
  assign new_G883_ = ~new_G663_;
  assign new_G884_ = new_G618_ | new_G621_;
  assign new_G887_ = ~new_G618_ & ~new_G621_;
  assign new_G890_ = ~new_G636_;
  assign new_G891_ = ~new_G639_;
  assign new_G892_ = ~new_G642_;
  assign new_G893_ = ~new_G645_;
  assign new_G894_ = ~new_G377_;
  assign new_G897_ = ~new_G648_;
  assign new_G898_ = ~new_G384_;
  assign new_G901_ = ~new_G400_;
  assign new_G904_ = ~new_G422_;
  assign new_G907_ = ~new_G434_;
  assign new_G910_ = ~new_G447_;
  assign new_G913_ = ~new_G461_;
  assign new_G916_ = ~new_G575_;
  assign new_G919_ = ~new_G575_;
  assign new_G922_ = ~new_G578_;
  assign new_G925_ = ~new_G578_;
  assign new_G928_ = ~new_G400_ | ~new_G713_;
  assign new_G929_ = new_G714_ & new_G715_ & new_G716_ & new_G717_;
  assign new_G930_ = new_G718_ & new_G719_ & new_G720_ & new_G721_;
  assign new_G931_ = ~new_G627_ | ~new_G722_;
  assign new_G932_ = ~new_G624_ | ~new_G723_;
  assign new_G933_ = ~new_G633_ | ~new_G724_;
  assign new_G934_ = ~new_G630_ | ~new_G725_;
  assign new_G935_ = new_G353_ & new_G726_;
  assign new_G939_ = new_G572_ & new_G784_;
  assign new_G956_ = ~new_G667_;
  assign new_G957_ = new_G501_ & new_G667_;
  assign new_G958_ = new_G785_ & new_G792_;
  assign new_G959_ = ~new_G667_;
  assign new_G960_ = new_G501_ & new_G667_;
  assign new_G961_ = ~new_G667_;
  assign new_G962_ = new_G501_ & new_G667_;
  assign new_G963_ = new_G552_ & new_G794_;
  assign new_G964_ = ~new_G667_;
  assign new_G965_ = new_G501_ & new_G667_;
  assign new_G966_ = n1860_lo & new_G795_;
  assign new_G967_ = ~new_G667_;
  assign new_G968_ = new_G501_ & new_G667_;
  assign new_G969_ = new_G790_ & new_G796_;
  assign new_G970_ = ~new_G667_;
  assign new_G971_ = new_G501_ & new_G667_;
  assign new_G972_ = ~new_G667_;
  assign new_G973_ = new_G501_ & new_G667_;
  assign new_G974_ = new_G568_ & new_G798_;
  assign new_G975_ = ~new_G667_;
  assign new_G976_ = new_G501_ & new_G667_;
  assign new_G977_ = n1908_lo & new_G799_;
  assign new_G978_ = n2076_lo & new_G848_;
  assign new_G979_ = n2088_lo & new_G849_;
  assign new_G980_ = n2100_lo & new_G850_;
  assign new_G981_ = n2112_lo & new_G851_;
  assign new_G982_ = n2124_lo & new_G852_;
  assign new_G983_ = n2136_lo & new_G853_;
  assign new_G984_ = n2148_lo & new_G854_;
  assign new_G985_ = n2160_lo & new_G855_;
  assign new_G986_ = n1752_lo & n1764_lo & new_G873_;
  assign new_G989_ = n1752_lo & n1764_lo & new_G874_;
  assign new_G992_ = ~new_G691_;
  assign new_G993_ = ~new_G691_;
  assign new_G994_ = ~new_G691_;
  assign new_G995_ = ~new_G691_;
  assign new_G996_ = ~new_G691_;
  assign new_G997_ = ~new_G691_;
  assign new_G998_ = ~new_G691_;
  assign new_G999_ = ~new_G691_;
  assign new_G1000_ = ~new_G639_ | ~new_G890_;
  assign new_G1001_ = ~new_G636_ | ~new_G891_;
  assign new_G1002_ = ~new_G645_ | ~new_G892_;
  assign new_G1003_ = ~new_G642_ | ~new_G893_;
  assign new_G1004_ = n1872_lo & new_G727_;
  assign new_G1005_ = ~new_G931_ | ~new_G932_;
  assign new_G1008_ = ~new_G933_ | ~new_G934_;
  assign new_G1011_ = ~new_G929_ | ~new_G930_;
  assign new_G1012_ = new_G461_ & new_G787_;
  assign new_G1015_ = ~new_G461_ | ~new_G787_;
  assign new_G1016_ = ~new_G731_;
  assign new_G1017_ = ~new_G916_ | ~new_G734_;
  assign new_G1018_ = ~new_G916_;
  assign new_G1019_ = new_G381_ & new_G731_;
  assign new_G1020_ = ~new_G922_ | ~new_G735_;
  assign new_G1021_ = ~new_G922_;
  assign new_G1022_ = ~n1872_lo | ~new_G727_;
  assign new_G1023_ = ~new_G736_;
  assign new_G1024_ = ~new_G739_;
  assign new_G1025_ = ~new_G772_ | ~new_G519_;
  assign new_G1034_ = ~new_G772_ | ~new_G523_;
  assign new_G1043_ = ~new_G470_ | ~new_G742_ | ~new_G496_;
  assign new_G1048_ = ~new_G470_ | ~new_G484_ | ~new_G496_ | ~new_G749_;
  assign new_G1051_ = ~new_G919_ | ~new_G786_;
  assign new_G1052_ = ~new_G919_;
  assign new_G1053_ = ~new_G925_ | ~new_G791_;
  assign new_G1054_ = ~new_G925_;
  assign new_G1055_ = ~new_G775_;
  assign new_G1056_ = ~new_G781_;
  assign new_G1057_ = ~new_G778_;
  assign new_G1058_ = new_G543_ & new_G956_;
  assign new_G1059_ = n1992_lo & new_G957_;
  assign new_G1060_ = new_G549_ & new_G959_;
  assign new_G1061_ = n2004_lo & new_G960_;
  assign new_G1062_ = n1860_lo & new_G961_;
  assign new_G1063_ = n1824_lo & new_G962_;
  assign new_G1064_ = new_G556_ & new_G964_;
  assign new_G1065_ = new_G543_ & new_G965_;
  assign new_G1066_ = new_G562_ & new_G967_;
  assign new_G1067_ = new_G549_ & new_G968_;
  assign new_G1068_ = n1896_lo & new_G970_;
  assign new_G1069_ = n1860_lo & new_G971_;
  assign new_G1070_ = n1908_lo & new_G972_;
  assign new_G1071_ = new_G556_ & new_G973_;
  assign new_G1072_ = n2208_lo & new_G975_;
  assign new_G1073_ = new_G562_ & new_G976_;
  assign new_G1074_ = n2052_lo & new_G810_;
  assign new_G1077_ = new_G587_ & new_G810_;
  assign new_G1080_ = new_G588_ & new_G813_;
  assign new_G1083_ = new_G589_ & new_G813_;
  assign new_G1086_ = ~new_G745_ | ~new_G749_;
  assign new_G1089_ = ~new_G519_ | ~new_G749_;
  assign new_G1092_ = ~new_G470_ | ~new_G742_ | ~new_G684_;
  assign new_G1095_ = ~new_G484_ | ~new_G492_ | ~new_G745_;
  assign new_G1104_ = ~new_G484_ | ~new_G745_;
  assign new_G1113_ = ~new_G816_;
  assign new_G1114_ = ~new_G816_;
  assign new_G1115_ = ~new_G816_;
  assign new_G1116_ = ~new_G816_;
  assign new_G1117_ = ~new_G816_;
  assign new_G1118_ = ~new_G816_;
  assign new_G1119_ = ~new_G816_;
  assign new_G1120_ = ~new_G831_;
  assign new_G1121_ = new_G831_ & new_G594_;
  assign new_G1122_ = ~new_G831_;
  assign new_G1123_ = new_G831_ & new_G594_;
  assign new_G1124_ = ~new_G831_;
  assign new_G1125_ = new_G831_ & new_G594_;
  assign new_G1126_ = ~new_G831_;
  assign new_G1127_ = new_G831_ & new_G594_;
  assign new_G1128_ = ~new_G831_;
  assign new_G1129_ = new_G831_ & new_G594_;
  assign new_G1130_ = ~new_G831_;
  assign new_G1131_ = new_G831_ & new_G594_;
  assign new_G1132_ = ~new_G831_;
  assign new_G1133_ = new_G831_ & new_G594_;
  assign new_G1134_ = ~new_G831_;
  assign new_G1135_ = new_G831_ & new_G594_;
  assign new_G1136_ = new_G691_ & new_G856_;
  assign new_G1137_ = ~n1824_lo & ~new_G856_;
  assign new_G1140_ = ~new_G753_;
  assign new_G1141_ = new_G691_ & new_G856_;
  assign new_G1142_ = ~n1836_lo & ~new_G856_;
  assign new_G1145_ = ~new_G753_;
  assign new_G1146_ = new_G691_ & new_G856_;
  assign new_G1147_ = ~n1848_lo & ~new_G856_;
  assign new_G1150_ = ~new_G753_;
  assign new_G1151_ = new_G691_ & new_G856_;
  assign new_G1152_ = ~n1860_lo & ~new_G856_;
  assign new_G1155_ = ~new_G753_;
  assign new_G1156_ = new_G691_ & new_G856_;
  assign new_G1157_ = ~n1872_lo & ~new_G856_;
  assign new_G1160_ = ~new_G769_;
  assign new_G1161_ = new_G691_ & new_G856_;
  assign new_G1162_ = ~n1884_lo & ~new_G856_;
  assign new_G1165_ = ~new_G762_;
  assign new_G1166_ = new_G691_ & new_G856_;
  assign new_G1167_ = ~n1896_lo & ~new_G856_;
  assign new_G1170_ = ~new_G762_;
  assign new_G1171_ = new_G691_ & new_G856_;
  assign new_G1172_ = ~n1908_lo & ~new_G856_;
  assign new_G1175_ = ~new_G762_;
  assign new_G1176_ = new_G875_ & n2064_lo;
  assign new_G1179_ = ~new_G875_ | ~n2064_lo;
  assign new_G1180_ = new_G875_ & n2064_lo & n2316_lo;
  assign new_G1184_ = ~new_G875_ | ~n2064_lo | ~n2316_lo;
  assign new_G1189_ = new_G875_ & n2064_lo & n2316_lo;
  assign new_G1193_ = ~new_G875_ | ~n2064_lo | ~n2316_lo;
  assign new_G1197_ = ~new_G887_;
  assign new_G1200_ = ~new_G1000_ | ~new_G1001_;
  assign new_G1203_ = ~new_G1002_ | ~new_G1003_;
  assign new_G1206_ = ~new_G894_;
  assign new_G1207_ = ~new_G894_ | ~new_G897_;
  assign new_G1208_ = ~new_G898_;
  assign new_G1209_ = ~new_G901_;
  assign new_G1210_ = ~new_G904_;
  assign new_G1211_ = ~new_G907_;
  assign new_G1212_ = ~new_G910_;
  assign new_G1213_ = ~new_G913_;
  assign new_G1214_ = ~new_G651_ | ~new_G1018_;
  assign new_G1215_ = ~new_G657_ | ~new_G1021_;
  assign new_G1216_ = new_G935_ & new_G739_;
  assign new_G1217_ = ~new_G654_ | ~new_G1052_;
  assign new_G1218_ = ~new_G660_ | ~new_G1054_;
  assign new_G1219_ = new_G666_ & new_G1055_;
  assign new_G1222_ = new_G958_ | new_G1058_ | new_G1059_;
  assign new_G1223_ = new_G963_ | new_G1062_ | new_G1063_;
  assign new_G1224_ = new_G966_ | new_G1064_ | new_G1065_;
  assign new_G1225_ = new_G969_ | new_G1066_ | new_G1067_;
  assign new_G1226_ = new_G974_ | new_G1070_ | new_G1071_;
  assign new_G1227_ = new_G977_ | new_G1072_ | new_G1073_;
  assign new_G1228_ = n1860_lo & new_G1120_;
  assign new_G1229_ = n2088_lo & new_G1121_;
  assign new_G1230_ = n1872_lo & new_G1122_;
  assign new_G1231_ = n2100_lo & new_G1123_;
  assign new_G1232_ = n1884_lo & new_G1124_;
  assign new_G1233_ = n2112_lo & new_G1125_;
  assign new_G1234_ = n1896_lo & new_G1126_;
  assign new_G1235_ = n2124_lo & new_G1127_;
  assign new_G1236_ = n1908_lo & new_G1128_;
  assign new_G1237_ = n2136_lo & new_G1129_;
  assign new_G1238_ = n2208_lo & new_G1130_;
  assign new_G1239_ = n2148_lo & new_G1131_;
  assign new_G1240_ = n2220_lo & new_G1132_;
  assign new_G1241_ = n2160_lo & new_G1133_;
  assign new_G1242_ = n2232_lo & new_G1134_;
  assign new_G1243_ = n2172_lo & new_G1135_;
  assign new_G1244_ = ~new_G986_;
  assign new_G1249_ = ~new_G986_;
  assign new_G1258_ = ~new_G989_;
  assign new_G1263_ = ~new_G989_;
  assign new_G1272_ = n1824_lo & new_G686_ & new_G1136_;
  assign new_G1275_ = n1836_lo & new_G686_ & new_G1141_;
  assign new_G1278_ = n1848_lo & new_G686_ & new_G1146_;
  assign new_G1281_ = n1860_lo & new_G686_ & new_G1151_;
  assign new_G1284_ = n1872_lo & new_G708_ & new_G1156_;
  assign new_G1287_ = n1884_lo & new_G708_ & new_G1161_;
  assign new_G1290_ = n1896_lo & new_G708_ & new_G1166_;
  assign new_G1293_ = n1908_lo & new_G708_ & new_G1171_;
  assign new_G1296_ = ~new_G939_;
  assign new_G1297_ = ~new_G939_;
  assign new_G1298_ = ~new_G939_;
  assign new_G1299_ = ~new_G939_;
  assign new_G1300_ = ~new_G939_;
  assign new_G1301_ = ~new_G939_;
  assign new_G1302_ = ~new_G939_;
  assign new_G1303_ = ~new_G939_;
  assign new_G1304_ = ~new_G648_ | ~new_G1206_;
  assign new_G1305_ = ~new_G901_ | ~new_G1208_;
  assign new_G1306_ = ~new_G898_ | ~new_G1209_;
  assign new_G1307_ = ~new_G907_ | ~new_G1210_;
  assign new_G1308_ = ~new_G904_ | ~new_G1211_;
  assign new_G1309_ = ~new_G913_ | ~new_G1212_;
  assign new_G1310_ = ~new_G910_ | ~new_G1213_;
  assign new_G1311_ = ~new_G1200_;
  assign new_G1312_ = ~new_G1203_;
  assign new_G1313_ = ~new_G1025_;
  assign new_G1314_ = new_G1025_ & new_G1034_;
  assign new_G1315_ = ~new_G1034_;
  assign new_G1316_ = ~new_G1017_ | ~new_G1214_;
  assign new_G1317_ = ~new_G1020_ | ~new_G1215_;
  assign new_G1318_ = new_G1012_ & new_G730_ & new_G363_ & n1836_lo;
  assign new_G1319_ = ~new_G1025_;
  assign new_G1320_ = new_G1025_ & new_G1034_;
  assign new_G1321_ = ~new_G1034_;
  assign new_G1322_ = ~new_G1025_;
  assign new_G1323_ = ~new_G1034_;
  assign new_G1324_ = new_G1025_ & new_G1034_;
  assign new_G1325_ = ~new_G1025_;
  assign new_G1326_ = ~new_G1034_;
  assign new_G1327_ = new_G1025_ & new_G1034_;
  assign new_G1328_ = ~new_G1048_;
  assign new_G1345_ = ~new_G1048_;
  assign new_G1348_ = ~new_G1051_ | ~new_G1217_;
  assign new_G1349_ = ~new_G1053_ | ~new_G1218_;
  assign new_G1350_ = ~new_G1043_;
  assign new_G1351_ = new_G1043_ & new_G775_;
  assign new_G1352_ = ~new_G1043_;
  assign new_G1353_ = new_G778_ & new_G1043_;
  assign new_G1354_ = ~new_G805_ | ~new_G1083_;
  assign new_G1357_ = ~new_G805_ | ~new_G1080_;
  assign new_G1360_ = ~new_G800_ | ~new_G1083_;
  assign new_G1363_ = ~new_G800_ | ~new_G1080_;
  assign new_G1366_ = ~new_G805_ | ~new_G1077_;
  assign new_G1369_ = ~new_G805_ | ~new_G1074_;
  assign new_G1372_ = ~new_G800_ | ~new_G1077_;
  assign new_G1375_ = ~new_G800_ | ~new_G1074_;
  assign new_G1378_ = ~new_G1086_;
  assign new_G1379_ = ~new_G1089_;
  assign new_G1380_ = new_G1086_ & new_G1089_;
  assign new_G1381_ = ~new_G1092_;
  assign new_G1390_ = ~new_G1092_;
  assign new_G1399_ = ~new_G1104_;
  assign new_G1400_ = ~new_G1104_;
  assign new_G1401_ = ~new_G1104_;
  assign new_G1402_ = ~new_G1104_;
  assign new_G1403_ = ~new_G1095_;
  assign new_G1404_ = ~new_G1095_;
  assign new_G1405_ = ~new_G1095_;
  assign new_G1406_ = ~new_G1095_;
  assign new_G1407_ = new_G1228_ | new_G978_ | new_G1229_;
  assign new_G1408_ = new_G1230_ | new_G979_ | new_G1231_;
  assign new_G1409_ = new_G1232_ | new_G980_ | new_G1233_;
  assign new_G1410_ = new_G1234_ | new_G981_ | new_G1235_;
  assign new_G1411_ = new_G1236_ | new_G982_ | new_G1237_;
  assign new_G1412_ = new_G1238_ | new_G983_ | new_G1239_;
  assign new_G1413_ = new_G1240_ | new_G984_ | new_G1241_;
  assign new_G1414_ = new_G1242_ | new_G985_ | new_G1243_;
  assign new_G1415_ = new_G1222_ & new_G992_;
  assign new_G1418_ = new_G1223_ & new_G994_;
  assign new_G1421_ = new_G1224_ & new_G995_;
  assign new_G1424_ = new_G1225_ & new_G996_;
  assign new_G1427_ = new_G1226_ & new_G998_;
  assign new_G1430_ = new_G1227_ & new_G999_;
  assign new_G1433_ = ~new_G1184_;
  assign new_G1436_ = new_G1197_ & n2340_lo;
  assign new_G1439_ = ~new_G1197_ | ~n2340_lo;
  assign new_G1442_ = ~new_G1005_;
  assign new_G1445_ = ~new_G1008_;
  assign new_G1448_ = ~new_G1005_;
  assign new_G1451_ = ~new_G1008_;
  assign new_G1454_ = ~new_G1207_ | ~new_G1304_;
  assign new_G1457_ = ~new_G1305_ | ~new_G1306_;
  assign new_G1460_ = ~new_G1307_ | ~new_G1308_;
  assign new_G1463_ = ~new_G1309_ | ~new_G1310_;
  assign new_G1466_ = ~new_G1203_ | ~new_G1311_;
  assign new_G1467_ = ~new_G1200_ | ~new_G1312_;
  assign new_G1468_ = new_G422_ & new_G1314_;
  assign new_G1469_ = new_G1316_ & new_G397_ & new_G1016_;
  assign new_G1470_ = new_G451_ & new_G1317_;
  assign new_G1471_ = new_G1318_ & new_G736_;
  assign new_G1472_ = new_G434_ & new_G1320_;
  assign new_G1473_ = new_G1022_ & new_G1323_;
  assign new_G1474_ = new_G461_ & new_G1324_;
  assign new_G1475_ = new_G1015_ & new_G1326_;
  assign new_G1476_ = new_G447_ & new_G1327_;
  assign new_G1477_ = ~new_G1348_;
  assign new_G1478_ = ~new_G1349_;
  assign new_G1479_ = new_G935_ & new_G1350_;
  assign new_G1482_ = new_G1011_ & new_G1351_;
  assign new_G1485_ = new_G363_ & new_G1380_;
  assign new_G1486_ = new_G1263_ & n2100_lo & new_G1140_;
  assign new_G1487_ = new_G1263_ & n2196_lo & new_G753_;
  assign new_G1488_ = new_G1258_ & new_G1407_;
  assign new_G1489_ = new_G1263_ & n2112_lo & new_G1145_;
  assign new_G1490_ = new_G1263_ & n2196_lo & new_G753_;
  assign new_G1491_ = new_G1258_ & new_G1408_;
  assign new_G1492_ = new_G1263_ & n2124_lo & new_G1150_;
  assign new_G1493_ = new_G1263_ & n2196_lo & new_G753_;
  assign new_G1494_ = new_G1258_ & new_G1409_;
  assign new_G1495_ = new_G1263_ & n2136_lo & new_G1155_;
  assign new_G1496_ = new_G1263_ & n2196_lo & new_G753_;
  assign new_G1497_ = new_G1258_ & new_G1410_;
  assign new_G1498_ = new_G1249_ & n2148_lo & new_G1160_;
  assign new_G1499_ = new_G1249_ & n2196_lo & new_G769_;
  assign new_G1500_ = new_G1244_ & new_G1411_;
  assign new_G1501_ = new_G1249_ & n2160_lo & new_G1165_;
  assign new_G1502_ = new_G1249_ & n2196_lo & new_G762_;
  assign new_G1503_ = new_G1244_ & new_G1412_;
  assign new_G1504_ = new_G1249_ & n2172_lo & new_G1170_;
  assign new_G1505_ = new_G1249_ & n2196_lo & new_G762_;
  assign new_G1506_ = new_G1244_ & new_G1413_;
  assign new_G1507_ = new_G1249_ & n2184_lo & new_G1175_;
  assign new_G1508_ = new_G1249_ & n2196_lo & new_G762_;
  assign new_G1509_ = new_G1244_ & new_G1414_;
  assign new_G1510_ = ~new_G1442_;
  assign new_G1511_ = ~new_G1445_;
  assign new_G1512_ = ~new_G1448_;
  assign new_G1513_ = ~new_G1451_;
  assign new_G1514_ = ~new_G1466_ | ~new_G1467_;
  assign new_G1517_ = ~new_G1454_;
  assign new_G1518_ = ~new_G1457_;
  assign new_G1519_ = ~new_G1460_;
  assign new_G1520_ = ~new_G1463_;
  assign new_G1521_ = new_G1469_ | new_G1019_;
  assign new_G1522_ = ~new_G1345_;
  assign new_G1523_ = new_G1345_ & new_G781_;
  assign new_G1524_ = new_G1470_ & new_G1352_;
  assign new_G1527_ = new_G1477_ & new_G793_;
  assign new_G1528_ = new_G1478_ & new_G797_;
  assign new_G1529_ = ~new_G1354_;
  assign new_G1538_ = ~new_G1357_;
  assign new_G1547_ = ~new_G1360_;
  assign new_G1556_ = ~new_G1363_;
  assign new_G1565_ = ~new_G1366_;
  assign new_G1574_ = ~new_G1369_;
  assign new_G1583_ = ~new_G1372_;
  assign new_G1592_ = ~new_G1375_;
  assign new_G1601_ = ~new_G1354_;
  assign new_G1610_ = ~new_G1357_;
  assign new_G1619_ = ~new_G1360_;
  assign new_G1628_ = ~new_G1363_;
  assign new_G1637_ = ~new_G1366_;
  assign new_G1646_ = ~new_G1369_;
  assign new_G1655_ = ~new_G1372_;
  assign new_G1664_ = ~new_G1375_;
  assign new_G1673_ = ~new_G1381_;
  assign new_G1674_ = new_G1381_ & new_G1104_;
  assign new_G1675_ = ~new_G1381_;
  assign new_G1676_ = new_G1381_ & new_G1104_;
  assign new_G1677_ = ~new_G1381_;
  assign new_G1678_ = new_G1381_ & new_G1104_;
  assign new_G1679_ = ~new_G1381_;
  assign new_G1680_ = new_G1381_ & new_G1104_;
  assign new_G1681_ = ~new_G1390_;
  assign new_G1682_ = new_G1390_ & new_G1095_;
  assign new_G1683_ = ~new_G1390_;
  assign new_G1684_ = new_G1390_ & new_G1095_;
  assign new_G1685_ = ~new_G1390_;
  assign new_G1686_ = new_G1390_ & new_G1095_;
  assign new_G1687_ = ~new_G1390_;
  assign new_G1688_ = new_G1390_ & new_G1095_;
  assign new_G1689_ = new_G1415_ | new_G1137_ | new_G1272_;
  assign new_G1693_ = ~new_G1415_ & ~new_G1137_ & ~new_G1272_;
  assign new_G1697_ = new_G1486_ | new_G1487_ | new_G1488_;
  assign new_G1700_ = new_G1489_ | new_G1490_ | new_G1491_;
  assign new_G1703_ = new_G1418_ | new_G1147_ | new_G1278_;
  assign new_G1707_ = ~new_G1418_ & ~new_G1147_ & ~new_G1278_;
  assign new_G1711_ = new_G1492_ | new_G1493_ | new_G1494_;
  assign new_G1714_ = new_G1421_ | new_G1152_ | new_G1281_;
  assign new_G1718_ = ~new_G1421_ & ~new_G1152_ & ~new_G1281_;
  assign new_G1722_ = new_G1495_ | new_G1496_ | new_G1497_;
  assign new_G1725_ = new_G1424_ | new_G1157_ | new_G1284_;
  assign new_G1729_ = ~new_G1424_ & ~new_G1157_ & ~new_G1284_;
  assign new_G1733_ = new_G1498_ | new_G1499_ | new_G1500_;
  assign new_G1738_ = new_G1501_ | new_G1502_ | new_G1503_;
  assign new_G1743_ = new_G1427_ | new_G1167_ | new_G1290_;
  assign new_G1747_ = ~new_G1427_ & ~new_G1167_ & ~new_G1290_;
  assign new_G1751_ = new_G1504_ | new_G1505_ | new_G1506_;
  assign new_G1756_ = new_G1430_ | new_G1172_ | new_G1293_;
  assign new_G1760_ = ~new_G1430_ & ~new_G1172_ & ~new_G1293_;
  assign new_G1764_ = new_G1507_ | new_G1508_ | new_G1509_;
  assign new_G1769_ = ~new_G1433_;
  assign new_G1770_ = ~new_G1328_;
  assign new_G1771_ = new_G939_ & new_G1328_;
  assign new_G1772_ = ~new_G1328_;
  assign new_G1773_ = new_G939_ & new_G1328_;
  assign new_G1774_ = ~new_G1328_;
  assign new_G1775_ = new_G939_ & new_G1328_;
  assign new_G1776_ = ~new_G1328_;
  assign new_G1777_ = new_G939_ & new_G1328_;
  assign new_G1778_ = ~new_G1328_;
  assign new_G1779_ = new_G939_ & new_G1328_;
  assign new_G1780_ = ~new_G1328_;
  assign new_G1781_ = new_G939_ & new_G1328_;
  assign new_G1782_ = ~new_G1328_;
  assign new_G1783_ = new_G939_ & new_G1328_;
  assign new_G1784_ = ~new_G1328_;
  assign new_G1785_ = new_G939_ & new_G1328_;
  assign new_G1786_ = new_G1479_ | new_G1219_ | new_G1482_;
  assign new_G1787_ = ~new_G1479_ & ~new_G1219_ & ~new_G1482_;
  assign new_G1788_ = ~new_G1445_ | ~new_G1510_;
  assign new_G1789_ = ~new_G1442_ | ~new_G1511_;
  assign new_G1790_ = ~new_G1451_ | ~new_G1512_;
  assign new_G1791_ = ~new_G1448_ | ~new_G1513_;
  assign new_G1792_ = ~new_G1457_ | ~new_G1517_;
  assign new_G1793_ = ~new_G1454_ | ~new_G1518_;
  assign new_G1794_ = ~new_G1463_ | ~new_G1519_;
  assign new_G1795_ = ~new_G1460_ | ~new_G1520_;
  assign new_G1796_ = new_G935_ & new_G1522_;
  assign new_G1799_ = new_G1012_ & new_G1523_;
  assign new_G1802_ = new_G1521_ & new_G1057_;
  assign new_G1805_ = new_G1527_ | new_G1060_ | new_G1061_;
  assign new_G1806_ = new_G1528_ | new_G1068_ | new_G1069_;
  assign new_G1807_ = new_G363_ & new_G1674_;
  assign new_G1808_ = new_G377_ & new_G1676_;
  assign new_G1809_ = new_G384_ & new_G1678_;
  assign new_G1810_ = new_G400_ & new_G1680_;
  assign new_G1811_ = ~new_G1787_;
  assign new_G1812_ = ~new_G1788_ | ~new_G1789_;
  assign new_G1813_ = ~new_G1790_ | ~new_G1791_;
  assign new_G1816_ = ~new_G1514_;
  assign new_G1819_ = ~new_G1792_ | ~new_G1793_;
  assign new_G1823_ = ~new_G1794_ | ~new_G1795_;
  assign new_G1826_ = new_G1514_ & new_G1313_;
  assign new_G1827_ = ~new_G1529_;
  assign new_G1828_ = ~new_G1538_;
  assign new_G1829_ = ~new_G1547_;
  assign new_G1830_ = ~new_G1556_;
  assign new_G1831_ = ~new_G1565_;
  assign new_G1832_ = ~new_G1574_;
  assign new_G1833_ = ~new_G1583_;
  assign new_G1834_ = ~new_G1592_;
  assign new_G1835_ = ~new_G1529_;
  assign new_G1836_ = ~new_G1538_;
  assign new_G1837_ = ~new_G1547_;
  assign new_G1838_ = ~new_G1556_;
  assign new_G1839_ = ~new_G1565_;
  assign new_G1840_ = ~new_G1574_;
  assign new_G1841_ = ~new_G1583_;
  assign new_G1842_ = ~new_G1592_;
  assign new_G1843_ = ~new_G1529_;
  assign new_G1844_ = ~new_G1538_;
  assign new_G1845_ = ~new_G1547_;
  assign new_G1846_ = ~new_G1556_;
  assign new_G1847_ = ~new_G1565_;
  assign new_G1848_ = ~new_G1574_;
  assign new_G1849_ = ~new_G1583_;
  assign new_G1850_ = ~new_G1592_;
  assign new_G1851_ = ~new_G1529_;
  assign new_G1852_ = ~new_G1538_;
  assign new_G1853_ = ~new_G1547_;
  assign new_G1854_ = ~new_G1556_;
  assign new_G1855_ = ~new_G1565_;
  assign new_G1856_ = ~new_G1574_;
  assign new_G1857_ = ~new_G1583_;
  assign new_G1858_ = ~new_G1592_;
  assign new_G1859_ = ~new_G1529_;
  assign new_G1860_ = ~new_G1538_;
  assign new_G1861_ = ~new_G1547_;
  assign new_G1862_ = ~new_G1556_;
  assign new_G1863_ = ~new_G1565_;
  assign new_G1864_ = ~new_G1574_;
  assign new_G1865_ = ~new_G1583_;
  assign new_G1866_ = ~new_G1592_;
  assign new_G1867_ = ~new_G1529_;
  assign new_G1868_ = ~new_G1538_;
  assign new_G1869_ = ~new_G1547_;
  assign new_G1870_ = ~new_G1556_;
  assign new_G1871_ = ~new_G1565_;
  assign new_G1872_ = ~new_G1574_;
  assign new_G1873_ = ~new_G1583_;
  assign new_G1874_ = ~new_G1592_;
  assign new_G1875_ = ~new_G1529_;
  assign new_G1876_ = ~new_G1538_;
  assign new_G1877_ = ~new_G1547_;
  assign new_G1878_ = ~new_G1556_;
  assign new_G1879_ = ~new_G1565_;
  assign new_G1880_ = ~new_G1574_;
  assign new_G1881_ = ~new_G1583_;
  assign new_G1882_ = ~new_G1592_;
  assign new_G1883_ = ~new_G1529_;
  assign new_G1884_ = ~new_G1538_;
  assign new_G1885_ = ~new_G1547_;
  assign new_G1886_ = ~new_G1556_;
  assign new_G1887_ = ~new_G1565_;
  assign new_G1888_ = ~new_G1574_;
  assign new_G1889_ = ~new_G1583_;
  assign new_G1890_ = ~new_G1592_;
  assign new_G1891_ = ~new_G1601_;
  assign new_G1892_ = ~new_G1610_;
  assign new_G1893_ = ~new_G1619_;
  assign new_G1894_ = ~new_G1628_;
  assign new_G1895_ = ~new_G1637_;
  assign new_G1896_ = ~new_G1646_;
  assign new_G1897_ = ~new_G1655_;
  assign new_G1898_ = ~new_G1664_;
  assign new_G1899_ = ~new_G1601_;
  assign new_G1900_ = ~new_G1610_;
  assign new_G1901_ = ~new_G1619_;
  assign new_G1902_ = ~new_G1628_;
  assign new_G1903_ = ~new_G1637_;
  assign new_G1904_ = ~new_G1646_;
  assign new_G1905_ = ~new_G1655_;
  assign new_G1906_ = ~new_G1664_;
  assign new_G1907_ = ~new_G1601_;
  assign new_G1908_ = ~new_G1610_;
  assign new_G1909_ = ~new_G1619_;
  assign new_G1910_ = ~new_G1628_;
  assign new_G1911_ = ~new_G1637_;
  assign new_G1912_ = ~new_G1646_;
  assign new_G1913_ = ~new_G1655_;
  assign new_G1914_ = ~new_G1664_;
  assign new_G1915_ = ~new_G1601_;
  assign new_G1916_ = ~new_G1610_;
  assign new_G1917_ = ~new_G1619_;
  assign new_G1918_ = ~new_G1628_;
  assign new_G1919_ = ~new_G1637_;
  assign new_G1920_ = ~new_G1646_;
  assign new_G1921_ = ~new_G1655_;
  assign new_G1922_ = ~new_G1664_;
  assign new_G1923_ = ~new_G1601_;
  assign new_G1924_ = ~new_G1610_;
  assign new_G1925_ = ~new_G1619_;
  assign new_G1926_ = ~new_G1628_;
  assign new_G1927_ = ~new_G1637_;
  assign new_G1928_ = ~new_G1646_;
  assign new_G1929_ = ~new_G1655_;
  assign new_G1930_ = ~new_G1664_;
  assign new_G1931_ = ~new_G1601_;
  assign new_G1932_ = ~new_G1610_;
  assign new_G1933_ = ~new_G1619_;
  assign new_G1934_ = ~new_G1628_;
  assign new_G1935_ = ~new_G1637_;
  assign new_G1936_ = ~new_G1646_;
  assign new_G1937_ = ~new_G1655_;
  assign new_G1938_ = ~new_G1664_;
  assign new_G1939_ = ~new_G1601_;
  assign new_G1940_ = ~new_G1610_;
  assign new_G1941_ = ~new_G1619_;
  assign new_G1942_ = ~new_G1628_;
  assign new_G1943_ = ~new_G1637_;
  assign new_G1944_ = ~new_G1646_;
  assign new_G1945_ = ~new_G1655_;
  assign new_G1946_ = ~new_G1664_;
  assign new_G1947_ = ~new_G1601_;
  assign new_G1948_ = ~new_G1610_;
  assign new_G1949_ = ~new_G1619_;
  assign new_G1950_ = ~new_G1628_;
  assign new_G1951_ = ~new_G1637_;
  assign new_G1952_ = ~new_G1646_;
  assign new_G1953_ = ~new_G1655_;
  assign new_G1954_ = ~new_G1664_;
  assign new_G1955_ = ~new_G1697_;
  assign new_G1958_ = ~new_G1697_;
  assign new_G1961_ = ~new_G1693_;
  assign new_G1962_ = new_G1805_ & new_G993_;
  assign new_G1965_ = ~new_G1700_;
  assign new_G1968_ = ~new_G1700_;
  assign new_G1971_ = ~new_G1711_;
  assign new_G1974_ = ~new_G1711_;
  assign new_G1977_ = ~new_G1707_;
  assign new_G1978_ = ~new_G1722_;
  assign new_G1981_ = ~new_G1722_;
  assign new_G1984_ = ~new_G1718_;
  assign new_G1985_ = ~new_G1733_;
  assign new_G1988_ = ~new_G1733_;
  assign new_G1991_ = ~new_G1729_;
  assign new_G1992_ = new_G1806_ & new_G997_;
  assign new_G1995_ = ~new_G1738_;
  assign new_G1998_ = ~new_G1738_;
  assign new_G2001_ = ~new_G1751_;
  assign new_G2004_ = ~new_G1751_;
  assign new_G2007_ = ~new_G1747_;
  assign new_G2008_ = ~new_G1764_;
  assign new_G2011_ = ~new_G1764_;
  assign new_G2014_ = ~new_G1760_;
  assign new_G2015_ = new_G1176_ & new_G1689_;
  assign new_G2018_ = new_G1180_ & new_G1703_;
  assign new_G2021_ = new_G1180_ & new_G1714_;
  assign new_G2024_ = new_G1180_ & new_G1725_;
  assign new_G2027_ = new_G1189_ & new_G1743_;
  assign new_G2030_ = new_G1189_ & new_G1756_;
  assign new_G2033_ = ~new_G1733_;
  assign new_G2034_ = ~new_G1738_;
  assign new_G2035_ = ~new_G1751_;
  assign new_G2036_ = ~new_G1764_;
  assign new_G2037_ = new_G1733_ & new_G1738_ & new_G1751_ & new_G1764_ & new_G882_;
  assign new_G2038_ = ~new_G1812_;
  assign new_G2039_ = new_G1826_ | new_G1315_ | new_G1468_;
  assign new_G2040_ = n1920_lo & new_G1827_;
  assign new_G2041_ = n2004_lo & new_G1828_;
  assign new_G2042_ = n1992_lo & new_G1829_;
  assign new_G2043_ = n1980_lo & new_G1830_;
  assign new_G2044_ = n1968_lo & new_G1831_;
  assign new_G2045_ = n1956_lo & new_G1832_;
  assign new_G2046_ = n1944_lo & new_G1833_;
  assign new_G2047_ = n1932_lo & new_G1834_;
  assign new_G2048_ = n1932_lo & new_G1835_;
  assign new_G2049_ = new_G353_ & new_G1836_;
  assign new_G2050_ = n2004_lo & new_G1837_;
  assign new_G2051_ = n1992_lo & new_G1838_;
  assign new_G2052_ = n1980_lo & new_G1839_;
  assign new_G2053_ = n1968_lo & new_G1840_;
  assign new_G2054_ = n1956_lo & new_G1841_;
  assign new_G2055_ = n1944_lo & new_G1842_;
  assign new_G2056_ = n1944_lo & new_G1843_;
  assign new_G2057_ = new_G368_ & new_G1844_;
  assign new_G2058_ = new_G353_ & new_G1845_;
  assign new_G2059_ = n2004_lo & new_G1846_;
  assign new_G2060_ = n1992_lo & new_G1847_;
  assign new_G2061_ = n1980_lo & new_G1848_;
  assign new_G2062_ = n1968_lo & new_G1849_;
  assign new_G2063_ = n1956_lo & new_G1850_;
  assign new_G2064_ = n1956_lo & new_G1851_;
  assign new_G2065_ = new_G388_ & new_G1852_;
  assign new_G2066_ = new_G368_ & new_G1853_;
  assign new_G2067_ = new_G353_ & new_G1854_;
  assign new_G2068_ = n2004_lo & new_G1855_;
  assign new_G2069_ = n1992_lo & new_G1856_;
  assign new_G2070_ = n1980_lo & new_G1857_;
  assign new_G2071_ = n1968_lo & new_G1858_;
  assign new_G2072_ = n1968_lo & new_G1859_;
  assign new_G2073_ = new_G404_ & new_G1860_;
  assign new_G2074_ = new_G388_ & new_G1861_;
  assign new_G2075_ = new_G368_ & new_G1862_;
  assign new_G2076_ = new_G353_ & new_G1863_;
  assign new_G2077_ = n2004_lo & new_G1864_;
  assign new_G2078_ = n1992_lo & new_G1865_;
  assign new_G2079_ = n1980_lo & new_G1866_;
  assign new_G2080_ = n1980_lo & new_G1867_;
  assign new_G2081_ = new_G413_ & new_G1868_;
  assign new_G2082_ = new_G404_ & new_G1869_;
  assign new_G2083_ = new_G388_ & new_G1870_;
  assign new_G2084_ = new_G368_ & new_G1871_;
  assign new_G2085_ = new_G353_ & new_G1872_;
  assign new_G2086_ = n2004_lo & new_G1873_;
  assign new_G2087_ = n1992_lo & new_G1874_;
  assign new_G2088_ = n1992_lo & new_G1875_;
  assign new_G2089_ = new_G425_ & new_G1876_;
  assign new_G2090_ = new_G413_ & new_G1877_;
  assign new_G2091_ = new_G404_ & new_G1878_;
  assign new_G2092_ = new_G388_ & new_G1879_;
  assign new_G2093_ = new_G368_ & new_G1880_;
  assign new_G2094_ = new_G353_ & new_G1881_;
  assign new_G2095_ = n2004_lo & new_G1882_;
  assign new_G2096_ = n2004_lo & new_G1883_;
  assign new_G2097_ = new_G438_ & new_G1884_;
  assign new_G2098_ = new_G425_ & new_G1885_;
  assign new_G2099_ = new_G413_ & new_G1886_;
  assign new_G2100_ = new_G404_ & new_G1887_;
  assign new_G2101_ = new_G388_ & new_G1888_;
  assign new_G2102_ = new_G368_ & new_G1889_;
  assign new_G2103_ = new_G353_ & new_G1890_;
  assign new_G2104_ = n2208_lo & new_G1891_;
  assign new_G2105_ = new_G368_ & new_G1892_;
  assign new_G2106_ = new_G388_ & new_G1893_;
  assign new_G2107_ = new_G404_ & new_G1894_;
  assign new_G2108_ = new_G413_ & new_G1895_;
  assign new_G2109_ = new_G425_ & new_G1896_;
  assign new_G2110_ = new_G438_ & new_G1897_;
  assign new_G2111_ = new_G451_ & new_G1898_;
  assign new_G2112_ = n2220_lo & new_G1899_;
  assign new_G2113_ = new_G388_ & new_G1900_;
  assign new_G2114_ = new_G404_ & new_G1901_;
  assign new_G2115_ = new_G413_ & new_G1902_;
  assign new_G2116_ = new_G425_ & new_G1903_;
  assign new_G2117_ = new_G438_ & new_G1904_;
  assign new_G2118_ = new_G451_ & new_G1905_;
  assign new_G2119_ = n2208_lo & new_G1906_;
  assign new_G2120_ = n2232_lo & new_G1907_;
  assign new_G2121_ = new_G404_ & new_G1908_;
  assign new_G2122_ = new_G413_ & new_G1909_;
  assign new_G2123_ = new_G425_ & new_G1910_;
  assign new_G2124_ = new_G438_ & new_G1911_;
  assign new_G2125_ = new_G451_ & new_G1912_;
  assign new_G2126_ = n2208_lo & new_G1913_;
  assign new_G2127_ = n2220_lo & new_G1914_;
  assign new_G2128_ = n2244_lo & new_G1915_;
  assign new_G2129_ = new_G413_ & new_G1916_;
  assign new_G2130_ = new_G425_ & new_G1917_;
  assign new_G2131_ = new_G438_ & new_G1918_;
  assign new_G2132_ = new_G451_ & new_G1919_;
  assign new_G2133_ = n2208_lo & new_G1920_;
  assign new_G2134_ = n2220_lo & new_G1921_;
  assign new_G2135_ = n2232_lo & new_G1922_;
  assign new_G2136_ = n2256_lo & new_G1923_;
  assign new_G2137_ = new_G425_ & new_G1924_;
  assign new_G2138_ = new_G438_ & new_G1925_;
  assign new_G2139_ = new_G451_ & new_G1926_;
  assign new_G2140_ = n2208_lo & new_G1927_;
  assign new_G2141_ = n2220_lo & new_G1928_;
  assign new_G2142_ = n2232_lo & new_G1929_;
  assign new_G2143_ = n2244_lo & new_G1930_;
  assign new_G2144_ = n2268_lo & new_G1931_;
  assign new_G2145_ = new_G438_ & new_G1932_;
  assign new_G2146_ = new_G451_ & new_G1933_;
  assign new_G2147_ = n2208_lo & new_G1934_;
  assign new_G2148_ = n2220_lo & new_G1935_;
  assign new_G2149_ = n2232_lo & new_G1936_;
  assign new_G2150_ = n2244_lo & new_G1937_;
  assign new_G2151_ = n2256_lo & new_G1938_;
  assign new_G2152_ = n2280_lo & new_G1939_;
  assign new_G2153_ = new_G451_ & new_G1940_;
  assign new_G2154_ = n2208_lo & new_G1941_;
  assign new_G2155_ = n2220_lo & new_G1942_;
  assign new_G2156_ = n2232_lo & new_G1943_;
  assign new_G2157_ = n2244_lo & new_G1944_;
  assign new_G2158_ = n2256_lo & new_G1945_;
  assign new_G2159_ = n2268_lo & new_G1946_;
  assign new_G2160_ = n2292_lo & new_G1947_;
  assign new_G2161_ = n2208_lo & new_G1948_;
  assign new_G2162_ = n2220_lo & new_G1949_;
  assign new_G2163_ = n2232_lo & new_G1950_;
  assign new_G2164_ = n2244_lo & new_G1951_;
  assign new_G2165_ = n2256_lo & new_G1952_;
  assign new_G2166_ = n2268_lo & new_G1953_;
  assign new_G2167_ = n2280_lo & new_G1954_;
  assign new_G2168_ = new_G2033_ & new_G2034_ & new_G2035_ & new_G2036_ & new_G615_;
  assign new_G2169_ = ~new_G1823_;
  assign new_G2172_ = new_G2038_ & new_G1023_;
  assign new_G2173_ = new_G1823_ & new_G1319_;
  assign new_G2174_ = new_G1819_ & new_G1024_;
  assign new_G2175_ = ~new_G2047_ & ~new_G2046_ & ~new_G2045_ & ~new_G2044_ & ~new_G2043_ & ~new_G2040_ & ~new_G2041_ & ~new_G2042_;
  assign new_G2176_ = ~new_G2055_ & ~new_G2054_ & ~new_G2053_ & ~new_G2052_ & ~new_G2051_ & ~new_G2048_ & ~new_G2049_ & ~new_G2050_;
  assign new_G2177_ = ~new_G2063_ & ~new_G2062_ & ~new_G2061_ & ~new_G2060_ & ~new_G2059_ & ~new_G2056_ & ~new_G2057_ & ~new_G2058_;
  assign new_G2178_ = ~new_G2071_ & ~new_G2070_ & ~new_G2069_ & ~new_G2068_ & ~new_G2067_ & ~new_G2064_ & ~new_G2065_ & ~new_G2066_;
  assign new_G2179_ = ~new_G2079_ & ~new_G2078_ & ~new_G2077_ & ~new_G2076_ & ~new_G2075_ & ~new_G2072_ & ~new_G2073_ & ~new_G2074_;
  assign new_G2180_ = ~new_G2087_ & ~new_G2086_ & ~new_G2085_ & ~new_G2084_ & ~new_G2083_ & ~new_G2080_ & ~new_G2081_ & ~new_G2082_;
  assign new_G2181_ = ~new_G2095_ & ~new_G2094_ & ~new_G2093_ & ~new_G2092_ & ~new_G2091_ & ~new_G2088_ & ~new_G2089_ & ~new_G2090_;
  assign new_G2182_ = ~new_G2103_ & ~new_G2102_ & ~new_G2101_ & ~new_G2100_ & ~new_G2099_ & ~new_G2096_ & ~new_G2097_ & ~new_G2098_;
  assign new_G2183_ = ~new_G2111_ & ~new_G2110_ & ~new_G2109_ & ~new_G2108_ & ~new_G2107_ & ~new_G2104_ & ~new_G2105_ & ~new_G2106_;
  assign new_G2184_ = ~new_G2119_ & ~new_G2118_ & ~new_G2117_ & ~new_G2116_ & ~new_G2115_ & ~new_G2112_ & ~new_G2113_ & ~new_G2114_;
  assign new_G2185_ = ~new_G2127_ & ~new_G2126_ & ~new_G2125_ & ~new_G2124_ & ~new_G2123_ & ~new_G2120_ & ~new_G2121_ & ~new_G2122_;
  assign new_G2186_ = ~new_G2135_ & ~new_G2134_ & ~new_G2133_ & ~new_G2132_ & ~new_G2131_ & ~new_G2128_ & ~new_G2129_ & ~new_G2130_;
  assign new_G2187_ = ~new_G2143_ & ~new_G2142_ & ~new_G2141_ & ~new_G2140_ & ~new_G2139_ & ~new_G2136_ & ~new_G2137_ & ~new_G2138_;
  assign new_G2188_ = ~new_G2151_ & ~new_G2150_ & ~new_G2149_ & ~new_G2148_ & ~new_G2147_ & ~new_G2144_ & ~new_G2145_ & ~new_G2146_;
  assign new_G2189_ = ~new_G2159_ & ~new_G2158_ & ~new_G2157_ & ~new_G2156_ & ~new_G2155_ & ~new_G2152_ & ~new_G2153_ & ~new_G2154_;
  assign new_G2190_ = ~new_G2167_ & ~new_G2166_ & ~new_G2165_ & ~new_G2164_ & ~new_G2163_ & ~new_G2160_ & ~new_G2161_ & ~new_G2162_;
  assign new_G2191_ = new_G2039_ & new_G1682_;
  assign new_G2192_ = n2016_lo & new_G1689_ & new_G1955_;
  assign new_G2195_ = n2028_lo & new_G1689_ & new_G1958_;
  assign new_G2198_ = n2040_lo & new_G1693_ & new_G1958_;
  assign new_G2199_ = n2052_lo & new_G1693_ & new_G1955_;
  assign new_G2200_ = new_G1962_ | new_G1142_ | new_G1275_;
  assign new_G2204_ = ~new_G1962_ & ~new_G1142_ & ~new_G1275_;
  assign new_G2208_ = n2016_lo & new_G1703_ & new_G1971_;
  assign new_G2211_ = n2028_lo & new_G1703_ & new_G1974_;
  assign new_G2214_ = n2040_lo & new_G1707_ & new_G1974_;
  assign new_G2215_ = n2052_lo & new_G1707_ & new_G1971_;
  assign new_G2216_ = n2016_lo & new_G1714_ & new_G1978_;
  assign new_G2219_ = n2028_lo & new_G1714_ & new_G1981_;
  assign new_G2222_ = n2040_lo & new_G1718_ & new_G1981_;
  assign new_G2223_ = n2052_lo & new_G1718_ & new_G1978_;
  assign new_G2224_ = n2016_lo & new_G1725_ & new_G1985_;
  assign new_G2227_ = n2028_lo & new_G1725_ & new_G1988_;
  assign new_G2230_ = n2040_lo & new_G1729_ & new_G1988_;
  assign new_G2231_ = n2052_lo & new_G1729_ & new_G1985_;
  assign new_G2232_ = new_G1992_ | new_G1162_ | new_G1287_;
  assign new_G2236_ = ~new_G1992_ & ~new_G1162_ & ~new_G1287_;
  assign new_G2240_ = n2016_lo & new_G1743_ & new_G2001_;
  assign new_G2243_ = n2028_lo & new_G1743_ & new_G2004_;
  assign new_G2246_ = n2040_lo & new_G1747_ & new_G2004_;
  assign new_G2247_ = n2052_lo & new_G1747_ & new_G2001_;
  assign new_G2248_ = n2016_lo & new_G1756_ & new_G2008_;
  assign new_G2251_ = n2028_lo & new_G1756_ & new_G2011_;
  assign new_G2254_ = n2040_lo & new_G1760_ & new_G2011_;
  assign new_G2255_ = n2052_lo & new_G1760_ & new_G2008_;
  assign new_G2256_ = new_G2037_ | new_G2168_;
  assign new_G2257_ = ~new_G1813_;
  assign new_G2260_ = ~new_G1816_;
  assign new_G2263_ = ~new_G1813_;
  assign new_G2266_ = ~new_G1816_;
  assign new_G2269_ = ~new_G1819_;
  assign new_G2272_ = ~new_G1819_;
  assign new_G2275_ = ~new_G2015_;
  assign new_G2278_ = ~new_G2015_;
  assign new_G2281_ = ~new_G2018_;
  assign new_G2284_ = ~new_G2018_;
  assign new_G2287_ = ~new_G2021_;
  assign new_G2290_ = ~new_G2021_;
  assign new_G2293_ = ~new_G2024_;
  assign new_G2296_ = ~new_G2024_;
  assign new_G2299_ = ~new_G2027_;
  assign new_G2302_ = ~new_G2027_;
  assign new_G2305_ = ~new_G2030_;
  assign new_G2308_ = ~new_G2030_;
  assign new_G2311_ = ~new_G2172_ & ~new_G1471_;
  assign new_G2312_ = new_G2173_ | new_G1321_ | new_G1472_;
  assign new_G2313_ = ~new_G2174_ & ~new_G1216_;
  assign new_G2314_ = new_G2175_ & new_G1378_;
  assign new_G2315_ = new_G2183_ & new_G1379_;
  assign new_G2316_ = new_G2176_ & new_G1113_;
  assign new_G2317_ = new_G2184_ & new_G816_;
  assign new_G2318_ = new_G2177_ & new_G1114_;
  assign new_G2319_ = new_G2185_ & new_G816_;
  assign new_G2320_ = new_G2178_ & new_G1115_;
  assign new_G2321_ = new_G2186_ & new_G816_;
  assign new_G2322_ = new_G2179_ & new_G1116_;
  assign new_G2323_ = new_G2187_ & new_G816_;
  assign new_G2324_ = new_G2180_ & new_G1117_;
  assign new_G2325_ = new_G2188_ & new_G816_;
  assign new_G2326_ = new_G2181_ & new_G1118_;
  assign new_G2327_ = new_G2189_ & new_G816_;
  assign new_G2328_ = new_G2182_ & new_G1119_;
  assign new_G2329_ = new_G2190_ & new_G816_;
  assign new_G2330_ = new_G2198_ | new_G2199_ | new_G1961_;
  assign new_G2331_ = new_G2214_ | new_G2215_ | new_G1977_;
  assign new_G2332_ = new_G2222_ | new_G2223_ | new_G1984_;
  assign new_G2333_ = new_G2230_ | new_G2231_ | new_G1991_;
  assign new_G2334_ = new_G2246_ | new_G2247_ | new_G2007_;
  assign new_G2335_ = new_G2254_ | new_G2255_ | new_G2014_;
  assign new_G2336_ = new_G2256_ & new_G1769_;
  assign new_G2337_ = ~new_G2263_;
  assign new_G2338_ = ~new_G2266_;
  assign new_G2339_ = ~new_G2272_;
  assign new_G2340_ = ~new_G2269_;
  assign new_G2341_ = ~new_G2257_;
  assign new_G2342_ = ~new_G2260_;
  assign new_G2343_ = new_G2313_ & new_G1322_;
  assign new_G2344_ = new_G2311_ & new_G1325_;
  assign new_G2345_ = new_G2314_ | new_G2315_ | new_G1485_;
  assign new_G2346_ = new_G2316_ | new_G2317_;
  assign new_G2347_ = new_G2318_ | new_G2319_;
  assign new_G2348_ = new_G2320_ | new_G2321_;
  assign new_G2349_ = new_G2322_ | new_G2323_;
  assign new_G2350_ = new_G2324_ | new_G2325_;
  assign new_G2351_ = new_G2326_ | new_G2327_;
  assign new_G2352_ = new_G2328_ | new_G2329_;
  assign new_G2353_ = new_G2312_ & new_G1684_;
  assign new_G2354_ = new_G2192_ | new_G2195_;
  assign new_G2355_ = ~new_G2192_ & ~new_G2195_;
  assign new_G2356_ = n2016_lo & new_G2200_ & new_G1965_;
  assign new_G2359_ = n2028_lo & new_G2200_ & new_G1968_;
  assign new_G2362_ = n2040_lo & new_G2204_ & new_G1968_;
  assign new_G2363_ = n2052_lo & new_G2204_ & new_G1965_;
  assign new_G2364_ = ~new_G2204_;
  assign new_G2365_ = new_G2208_ | new_G2211_;
  assign new_G2368_ = ~new_G2208_ & ~new_G2211_;
  assign new_G2369_ = new_G2216_ | new_G2219_;
  assign new_G2372_ = ~new_G2216_ & ~new_G2219_;
  assign new_G2373_ = new_G2224_ | new_G2227_;
  assign new_G2374_ = ~new_G2224_ & ~new_G2227_;
  assign new_G2375_ = n2016_lo & new_G2232_ & new_G1995_;
  assign new_G2378_ = n2028_lo & new_G2232_ & new_G1998_;
  assign new_G2381_ = n2040_lo & new_G2236_ & new_G1998_;
  assign new_G2382_ = n2052_lo & new_G2236_ & new_G1995_;
  assign new_G2383_ = ~new_G2236_;
  assign new_G2384_ = new_G2240_ | new_G2243_;
  assign new_G2387_ = ~new_G2240_ & ~new_G2243_;
  assign new_G2388_ = new_G2248_ | new_G2251_;
  assign new_G2391_ = ~new_G2248_ & ~new_G2251_;
  assign new_G2392_ = ~new_G2278_;
  assign new_G2393_ = new_G1176_ & new_G2200_;
  assign new_G2396_ = ~new_G2281_;
  assign new_G2397_ = ~new_G2284_;
  assign new_G2398_ = ~new_G2287_;
  assign new_G2399_ = ~new_G2290_;
  assign new_G2400_ = ~new_G2296_;
  assign new_G2401_ = new_G1189_ & new_G2232_;
  assign new_G2404_ = ~new_G2302_;
  assign new_G2405_ = ~new_G2305_;
  assign new_G2406_ = ~new_G2308_;
  assign new_G2407_ = ~new_G2299_;
  assign new_G2408_ = ~new_G2169_;
  assign new_G2411_ = ~new_G2169_;
  assign new_G2414_ = ~new_G2275_;
  assign new_G2415_ = ~new_G2293_;
  assign new_G2416_ = ~new_G2260_ | ~new_G2341_;
  assign new_G2417_ = ~new_G2257_ | ~new_G2342_;
  assign new_G2418_ = ~new_G2266_ | ~new_G2337_;
  assign new_G2419_ = ~new_G2263_ | ~new_G2338_;
  assign new_G2420_ = new_G2343_ | new_G1473_ | new_G1474_;
  assign new_G2421_ = new_G2344_ | new_G1475_ | new_G1476_;
  assign new_G2422_ = new_G2345_ & new_G1673_;
  assign new_G2423_ = new_G2346_ & new_G1675_;
  assign new_G2424_ = new_G2347_ & new_G1677_;
  assign new_G2425_ = new_G2348_ & new_G1679_;
  assign new_G2426_ = new_G2349_ & new_G1681_;
  assign new_G2427_ = new_G2350_ & new_G1683_;
  assign new_G2428_ = new_G2351_ & new_G1685_;
  assign new_G2429_ = new_G2352_ & new_G1687_;
  assign new_G2430_ = new_G2355_ & new_G2330_;
  assign new_G2436_ = new_G2362_ | new_G2363_ | new_G2364_;
  assign new_G2437_ = new_G2368_ & new_G2331_;
  assign new_G2441_ = new_G2372_ & new_G2332_;
  assign new_G2444_ = new_G2374_ & new_G2333_;
  assign new_G2450_ = new_G2381_ | new_G2382_ | new_G2383_;
  assign new_G2451_ = new_G2387_ & new_G2334_;
  assign new_G2455_ = new_G2391_ & new_G2335_;
  assign new_G2458_ = ~new_G2354_;
  assign new_G2459_ = ~new_G2373_;
  assign new_G2460_ = ~new_G2416_ | ~new_G2417_;
  assign new_G2461_ = ~new_G2418_ | ~new_G2419_;
  assign new_G2462_ = ~new_G2411_ | ~new_G2339_;
  assign new_G2463_ = ~new_G2411_;
  assign new_G2464_ = ~new_G2408_ | ~new_G2340_;
  assign new_G2465_ = ~new_G2408_;
  assign new_G2466_ = new_G2421_ & new_G1686_;
  assign new_G2467_ = new_G2420_ & new_G1688_;
  assign new_G2468_ = new_G2356_ | new_G2359_;
  assign new_G2471_ = ~new_G2356_ & ~new_G2359_;
  assign new_G2472_ = new_G2375_ | new_G2378_;
  assign new_G2475_ = ~new_G2375_ & ~new_G2378_;
  assign new_G2476_ = new_G2365_ & new_G1184_;
  assign new_G2479_ = new_G2369_ & new_G1184_;
  assign new_G2482_ = new_G2384_ & new_G1193_;
  assign new_G2485_ = new_G2388_ & new_G1193_;
  assign new_G2488_ = ~new_G2393_;
  assign new_G2491_ = ~new_G2393_;
  assign new_G2494_ = ~new_G2401_;
  assign new_G2497_ = ~new_G2401_;
  assign new_G2500_ = ~new_G2272_ | ~new_G2463_;
  assign new_G2501_ = ~new_G2269_ | ~new_G2465_;
  assign new_G2502_ = new_G2471_ & new_G2436_;
  assign new_G2507_ = new_G2475_ & new_G2450_;
  assign new_G2512_ = ~new_G2430_;
  assign new_G2515_ = ~new_G2437_;
  assign new_G2518_ = ~new_G2441_;
  assign new_G2521_ = ~new_G2444_;
  assign new_G2524_ = ~new_G2451_;
  assign new_G2527_ = ~new_G2455_;
  assign new_G2530_ = ~new_G2462_ | ~new_G2500_;
  assign new_G2531_ = ~new_G2464_ | ~new_G2501_;
  assign new_G2532_ = ~new_G2430_ | ~new_G2468_;
  assign new_G2533_ = ~new_G2444_ | ~new_G2472_;
  assign new_G2534_ = ~new_G2488_;
  assign new_G2535_ = ~new_G2491_;
  assign new_G2536_ = ~new_G2497_;
  assign new_G2537_ = ~new_G2494_;
  assign new_G2538_ = new_G2468_ & new_G1179_;
  assign new_G2539_ = ~new_G2479_;
  assign new_G2542_ = new_G2472_ & new_G1184_;
  assign new_G2543_ = ~new_G2485_;
  assign new_G2546_ = ~new_G2476_;
  assign new_G2547_ = ~new_G2485_;
  assign new_G2550_ = ~new_G2530_;
  assign new_G2551_ = ~new_G2531_;
  assign new_G2552_ = new_G2430_ & new_G2502_ & new_G2437_ & new_G2441_;
  assign new_G2556_ = ~new_G2430_ | ~new_G2502_ | ~new_G2365_;
  assign new_G2557_ = ~new_G2369_ | ~new_G2502_ | ~new_G2437_ | ~new_G2430_;
  assign new_G2558_ = new_G2444_ & new_G2507_ & new_G2451_ & new_G2455_;
  assign new_G2561_ = ~new_G2444_ | ~new_G2507_ | ~new_G2384_;
  assign new_G2562_ = ~new_G2388_ | ~new_G2507_ | ~new_G2451_ | ~new_G2444_;
  assign new_G2563_ = ~new_G2502_;
  assign new_G2566_ = ~new_G2507_;
  assign new_G2569_ = ~new_G2538_;
  assign new_G2570_ = ~new_G2542_;
  assign new_G2571_ = ~new_G2512_;
  assign new_G2574_ = ~new_G2512_;
  assign new_G2577_ = ~new_G2515_;
  assign new_G2580_ = ~new_G2515_;
  assign new_G2583_ = ~new_G2518_;
  assign new_G2586_ = ~new_G2518_;
  assign new_G2589_ = ~new_G2521_;
  assign new_G2592_ = ~new_G2521_;
  assign new_G2595_ = ~new_G2524_;
  assign new_G2598_ = ~new_G2524_;
  assign new_G2601_ = ~new_G2527_;
  assign new_G2604_ = ~new_G2527_;
  assign new_G2607_ = ~new_G2458_ | ~new_G2532_ | ~new_G2556_ | ~new_G2557_;
  assign new_G2610_ = ~new_G2459_ | ~new_G2533_ | ~new_G2561_ | ~new_G2562_;
  assign new_G2613_ = ~new_G2547_;
  assign new_G2614_ = ~new_G2574_ | ~new_G2392_;
  assign new_G2615_ = ~new_G2580_ | ~new_G2397_;
  assign new_G2616_ = ~new_G2586_ | ~new_G2399_;
  assign new_G2617_ = ~new_G2592_ | ~new_G2400_;
  assign new_G2618_ = ~new_G2598_ | ~new_G2404_;
  assign new_G2619_ = ~new_G2604_ | ~new_G2406_;
  assign new_G2620_ = ~new_G2552_;
  assign new_G2623_ = ~new_G2574_;
  assign new_G2624_ = ~new_G2577_;
  assign new_G2625_ = ~new_G2577_ | ~new_G2396_;
  assign new_G2626_ = ~new_G2580_;
  assign new_G2627_ = ~new_G2583_;
  assign new_G2628_ = ~new_G2583_ | ~new_G2398_;
  assign new_G2629_ = ~new_G2586_;
  assign new_G2630_ = ~new_G2592_;
  assign new_G2631_ = ~new_G2598_;
  assign new_G2632_ = ~new_G2601_;
  assign new_G2633_ = ~new_G2601_ | ~new_G2405_;
  assign new_G2634_ = ~new_G2604_;
  assign new_G2635_ = ~new_G2595_;
  assign new_G2636_ = ~new_G2595_ | ~new_G2407_;
  assign new_G2637_ = new_G2558_ & new_G1433_;
  assign new_G2638_ = ~new_G2571_;
  assign new_G2639_ = ~new_G2571_ | ~new_G2414_;
  assign new_G2640_ = ~new_G2563_;
  assign new_G2643_ = ~new_G2563_;
  assign new_G2646_ = ~new_G2589_;
  assign new_G2647_ = ~new_G2589_ | ~new_G2415_;
  assign new_G2648_ = ~new_G2566_;
  assign new_G2651_ = ~new_G2566_;
  assign new_G2654_ = ~new_G2552_ | ~new_G2610_;
  assign new_G2655_ = ~new_G2607_;
  assign new_G2656_ = ~new_G2278_ | ~new_G2623_;
  assign new_G2657_ = ~new_G2284_ | ~new_G2626_;
  assign new_G2658_ = ~new_G2290_ | ~new_G2629_;
  assign new_G2659_ = ~new_G2296_ | ~new_G2630_;
  assign new_G2660_ = ~new_G2302_ | ~new_G2631_;
  assign new_G2661_ = ~new_G2308_ | ~new_G2634_;
  assign new_G2662_ = ~new_G2281_ | ~new_G2624_;
  assign new_G2663_ = ~new_G2287_ | ~new_G2627_;
  assign new_G2664_ = ~new_G2305_ | ~new_G2632_;
  assign new_G2665_ = ~new_G2299_ | ~new_G2635_;
  assign new_G2666_ = new_G2610_ & new_G1193_;
  assign new_G2669_ = new_G2336_ | new_G2637_;
  assign new_G2673_ = ~new_G2275_ | ~new_G2638_;
  assign new_G2674_ = ~new_G2293_ | ~new_G2646_;
  assign new_G2675_ = new_G2654_ & new_G2655_;
  assign new_G2676_ = ~new_G2656_ | ~new_G2614_;
  assign new_G2677_ = ~new_G2643_ | ~new_G2535_;
  assign new_G2678_ = ~new_G2657_ | ~new_G2615_;
  assign new_G2679_ = ~new_G2658_ | ~new_G2616_;
  assign new_G2680_ = ~new_G2659_ | ~new_G2617_;
  assign new_G2681_ = ~new_G2651_ | ~new_G2536_;
  assign new_G2682_ = ~new_G2660_ | ~new_G2618_;
  assign new_G2683_ = ~new_G2661_ | ~new_G2619_;
  assign new_G2684_ = ~new_G2640_;
  assign new_G2685_ = ~new_G2640_ | ~new_G2534_;
  assign new_G2686_ = ~new_G2643_;
  assign new_G2687_ = ~new_G2662_ | ~new_G2625_;
  assign new_G2690_ = ~new_G2663_ | ~new_G2628_;
  assign new_G2693_ = ~new_G2651_;
  assign new_G2694_ = ~new_G2664_ | ~new_G2633_;
  assign new_G2697_ = ~new_G2648_;
  assign new_G2698_ = ~new_G2648_ | ~new_G2537_;
  assign new_G2699_ = ~new_G2665_ | ~new_G2636_;
  assign new_G2705_ = ~new_G2673_ | ~new_G2639_;
  assign new_G2708_ = ~new_G2674_ | ~new_G2647_;
  assign new_G2711_ = ~new_G2676_;
  assign new_G2712_ = ~new_G2491_ | ~new_G2686_;
  assign new_G2713_ = ~new_G2678_;
  assign new_G2714_ = ~new_G2679_;
  assign new_G2715_ = ~new_G2680_;
  assign new_G2716_ = ~new_G2497_ | ~new_G2693_;
  assign new_G2717_ = ~new_G2682_;
  assign new_G2718_ = ~new_G2683_;
  assign new_G2719_ = ~new_G2488_ | ~new_G2684_;
  assign new_G2720_ = ~new_G2494_ | ~new_G2697_;
  assign new_G2721_ = ~new_G2666_;
  assign new_G2728_ = ~new_G2669_;
  assign new_G2733_ = ~new_G2666_;
  assign new_G2736_ = n2304_lo & new_G2669_;
  assign new_G2739_ = new_G2711_ & new_G1399_;
  assign new_G2740_ = ~new_G2712_ | ~new_G2677_;
  assign new_G2741_ = new_G2713_ & new_G1401_;
  assign new_G2742_ = new_G2714_ & new_G1402_;
  assign new_G2743_ = new_G2715_ & new_G1403_;
  assign new_G2744_ = ~new_G2716_ | ~new_G2681_;
  assign new_G2745_ = new_G2717_ & new_G1405_;
  assign new_G2746_ = new_G2718_ & new_G1406_;
  assign new_G2747_ = ~new_G2719_ | ~new_G2685_;
  assign new_G2750_ = ~new_G2687_;
  assign new_G2753_ = ~new_G2687_;
  assign new_G2759_ = ~new_G2690_;
  assign new_G2763_ = ~new_G2690_;
  assign new_G2768_ = ~new_G2720_ | ~new_G2698_;
  assign new_G2773_ = ~new_G2694_;
  assign new_G2778_ = new_G2699_ & new_G2543_;
  assign new_G2779_ = ~new_G2705_;
  assign new_G2780_ = ~new_G2708_;
  assign new_G2781_ = n2304_lo & new_G2694_;
  assign new_G2784_ = ~new_G2699_;
  assign new_G2787_ = ~new_G2422_ & ~new_G2739_ & ~new_G1807_;
  assign new_G2788_ = ~new_G2740_;
  assign new_G2789_ = ~new_G2424_ & ~new_G2741_ & ~new_G1809_;
  assign new_G2790_ = ~new_G2425_ & ~new_G2742_ & ~new_G1810_;
  assign new_G2791_ = ~new_G2426_ & ~new_G2743_ & ~new_G2191_;
  assign new_G2792_ = ~new_G2744_;
  assign new_G2793_ = ~new_G2428_ & ~new_G2745_ & ~new_G2466_;
  assign new_G2794_ = ~new_G2429_ & ~new_G2746_ & ~new_G2467_;
  assign new_G2795_ = new_G2721_ & new_G2620_;
  assign new_G2796_ = new_G2728_ & new_G2620_;
  assign new_G2799_ = new_G2482_ | new_G2778_;
  assign new_G2803_ = ~new_G2736_;
  assign new_G2804_ = ~new_G2721_;
  assign new_G2805_ = ~new_G2721_;
  assign new_G2808_ = ~new_G2733_;
  assign new_G2809_ = new_G2788_ & new_G1400_;
  assign new_G2810_ = new_G2792_ & new_G1404_;
  assign new_G2811_ = ~new_G2747_;
  assign new_G2816_ = new_G2607_ | new_G2795_;
  assign new_G2820_ = new_G2728_ & new_G2763_ & new_G2753_;
  assign new_G2821_ = new_G2728_ & new_G2759_;
  assign new_G2822_ = new_G2773_ & new_G2699_ & new_G2768_;
  assign new_G2823_ = new_G2773_ & new_G2699_;
  assign new_G2826_ = new_G2721_ & new_G2759_;
  assign new_G2827_ = ~new_G2753_ | ~new_G2539_;
  assign new_G2828_ = ~new_G2753_ | ~new_G2763_ | ~new_G2721_;
  assign new_G2829_ = ~new_G2768_ | ~new_G2482_;
  assign new_G2830_ = ~new_G2768_ | ~new_G2699_ | ~new_G2543_;
  assign new_G2831_ = ~new_G2784_ | ~new_G2613_;
  assign new_G2832_ = ~new_G2784_;
  assign new_G2833_ = n2304_lo & new_G2669_ & new_G2804_;
  assign new_G2836_ = new_G2787_ & new_G1771_;
  assign new_G2839_ = new_G2789_ & new_G1775_;
  assign new_G2842_ = new_G2790_ & new_G1777_;
  assign new_G2845_ = new_G2791_ & new_G1779_;
  assign new_G2848_ = new_G2793_ & new_G1783_;
  assign new_G2851_ = new_G2794_ & new_G1785_;
  assign new_G2854_ = ~new_G2747_;
  assign new_G2857_ = ~new_G2753_;
  assign new_G2860_ = ~new_G2759_;
  assign new_G2863_ = ~new_G2768_;
  assign new_G2866_ = ~new_G2781_;
  assign new_G2869_ = ~new_G2781_;
  assign new_G2872_ = new_G2773_ & new_G2773_;
  assign new_G2875_ = ~new_G2423_ & ~new_G2809_ & ~new_G1808_;
  assign new_G2876_ = ~new_G2427_ & ~new_G2810_ & ~new_G2353_;
  assign new_G2877_ = n2304_lo & new_G2821_;
  assign new_G2880_ = n2304_lo & new_G2822_;
  assign new_G2883_ = ~new_G2547_ | ~new_G2832_;
  assign new_G2884_ = ~new_G2799_;
  assign new_G2887_ = ~new_G2796_;
  assign new_G2890_ = ~new_G2546_ | ~new_G2827_ | ~new_G2828_;
  assign new_G2893_ = new_G2479_ | new_G2826_;
  assign new_G2896_ = ~new_G2570_ | ~new_G2829_ | ~new_G2830_;
  assign new_G2899_ = ~new_G2799_;
  assign new_G2902_ = n2304_lo & new_G2820_;
  assign new_G2905_ = new_G2833_ | new_G2805_;
  assign new_G2906_ = new_G2728_ & new_G2811_ & new_G2753_ & new_G2763_;
  assign new_G2909_ = ~new_G2811_ | ~new_G2476_;
  assign new_G2910_ = ~new_G2811_ | ~new_G2750_ | ~new_G2539_;
  assign new_G2911_ = ~new_G2811_ | ~new_G2750_ | ~new_G2763_ | ~new_G2721_;
  assign new_G2912_ = ~new_G2857_;
  assign new_G2913_ = ~new_G2831_ | ~new_G2883_;
  assign new_G2916_ = ~new_G2866_;
  assign new_G2917_ = ~new_G2869_;
  assign new_G2918_ = ~new_G2872_ | ~new_G883_;
  assign new_G2919_ = ~new_G2872_;
  assign new_G2920_ = ~new_G2816_;
  assign new_G2923_ = ~new_G2833_ & ~new_G2805_;
  assign new_G2926_ = new_G2875_ & new_G1773_;
  assign new_G2929_ = new_G2876_ & new_G1781_;
  assign new_G2932_ = ~new_G2816_;
  assign new_G2935_ = ~new_G2854_;
  assign new_G2936_ = ~new_G2860_;
  assign new_G2937_ = ~new_G2860_ | ~new_G2808_;
  assign new_G2938_ = ~new_G2863_;
  assign new_G2939_ = n2304_lo & new_G2823_;
  assign new_G2942_ = ~new_G2884_;
  assign new_G2943_ = new_G2799_ & new_G2884_;
  assign new_G2944_ = new_G2905_ & new_G1056_;
  assign new_G2947_ = ~new_G2569_ | ~new_G2909_ | ~new_G2910_ | ~new_G2911_;
  assign new_G2950_ = ~new_G2887_;
  assign new_G2951_ = ~new_G2902_;
  assign new_G2952_ = ~new_G2893_;
  assign new_G2953_ = ~new_G2893_ | ~new_G2912_;
  assign new_G2954_ = ~new_G2896_;
  assign new_G2955_ = ~new_G2896_ | ~new_G2780_;
  assign new_G2956_ = ~new_G663_ | ~new_G2919_;
  assign new_G2957_ = ~new_G2890_;
  assign new_G2958_ = ~new_G2890_ | ~new_G2935_;
  assign new_G2959_ = ~new_G2733_ | ~new_G2936_;
  assign new_G2960_ = ~new_G2899_;
  assign new_G2961_ = ~new_G2899_ | ~new_G2938_;
  assign new_G2962_ = ~new_G2877_;
  assign new_G2965_ = ~new_G2877_;
  assign new_G2968_ = ~new_G2880_;
  assign new_G2971_ = ~new_G2880_;
  assign new_G2974_ = n2304_lo & new_G2823_ & new_G2942_;
  assign new_G2975_ = n2304_lo & new_G2906_;
  assign new_G2978_ = ~new_G2857_ | ~new_G2952_;
  assign new_G2979_ = ~new_G2708_ | ~new_G2954_;
  assign new_G2980_ = ~new_G2939_;
  assign new_G2981_ = ~new_G2918_ | ~new_G2956_;
  assign new_G2984_ = ~new_G2920_;
  assign new_G2985_ = new_G2816_ & new_G2920_;
  assign new_G2986_ = ~new_G2923_;
  assign new_G2990_ = ~new_G2932_;
  assign new_G2991_ = ~new_G2906_;
  assign new_G2994_ = ~new_G2854_ | ~new_G2957_;
  assign new_G2995_ = ~new_G2863_ | ~new_G2960_;
  assign new_G2996_ = ~new_G2937_ | ~new_G2959_;
  assign new_G2999_ = ~new_G2913_;
  assign new_G3002_ = ~new_G2913_;
  assign new_G3005_ = new_G1796_ | new_G2944_ | new_G1799_;
  assign new_G3006_ = ~new_G1796_ & ~new_G2944_ & ~new_G1799_;
  assign new_G3007_ = ~new_G2978_ | ~new_G2953_;
  assign new_G3010_ = ~new_G2962_;
  assign new_G3011_ = ~new_G2965_;
  assign new_G3012_ = ~new_G2979_ | ~new_G2955_;
  assign new_G3015_ = ~new_G2968_;
  assign new_G3016_ = ~new_G2971_;
  assign new_G3017_ = n2304_lo & new_G2796_ & new_G2984_;
  assign new_G3018_ = ~new_G2947_;
  assign new_G3021_ = ~new_G2947_;
  assign new_G3024_ = ~new_G2994_ | ~new_G2958_;
  assign new_G3027_ = ~new_G2995_ | ~new_G2961_;
  assign new_G3030_ = ~new_G3006_;
  assign new_G3031_ = ~new_G2991_ | ~new_G2950_;
  assign new_G3032_ = ~new_G2991_;
  assign new_G3033_ = ~new_G2996_;
  assign new_G3034_ = ~new_G2996_ | ~new_G2803_;
  assign new_G3035_ = ~new_G2999_;
  assign new_G3036_ = ~new_G2999_ | ~new_G2916_;
  assign new_G3037_ = ~new_G3002_;
  assign new_G3038_ = ~new_G3002_ | ~new_G2917_;
  assign new_G3039_ = ~new_G3017_ & ~new_G2985_;
  assign new_G3042_ = new_G2981_ & new_G1303_;
  assign new_G3045_ = new_G2981_ & new_G1784_;
  assign new_G3048_ = ~new_G2975_;
  assign new_G3051_ = ~new_G2975_;
  assign new_G3054_ = ~new_G2986_;
  assign new_G3057_ = ~new_G2887_ | ~new_G3032_;
  assign new_G3058_ = ~new_G3021_;
  assign new_G3059_ = ~new_G3021_ | ~new_G2779_;
  assign new_G3060_ = ~new_G3024_;
  assign new_G3061_ = ~new_G3024_ | ~new_G2951_;
  assign new_G3062_ = ~new_G2736_ | ~new_G3033_;
  assign new_G3063_ = ~new_G3027_;
  assign new_G3064_ = ~new_G3027_ | ~new_G2980_;
  assign new_G3065_ = ~new_G2866_ | ~new_G3035_;
  assign new_G3066_ = ~new_G2869_ | ~new_G3037_;
  assign new_G3067_ = ~new_G3018_;
  assign new_G3068_ = ~new_G3018_ | ~new_G2990_;
  assign new_G3069_ = ~new_G3007_;
  assign new_G3072_ = ~new_G3007_;
  assign new_G3075_ = ~new_G3012_;
  assign new_G3078_ = ~new_G3012_;
  assign new_G3081_ = ~new_G3031_ | ~new_G3057_;
  assign new_G3082_ = ~new_G2705_ | ~new_G3058_;
  assign new_G3083_ = ~new_G3048_;
  assign new_G3084_ = ~new_G3051_;
  assign new_G3085_ = ~new_G2902_ | ~new_G3060_;
  assign new_G3086_ = ~new_G3062_ | ~new_G3034_;
  assign new_G3089_ = ~new_G2939_ | ~new_G3063_;
  assign new_G3090_ = ~new_G3065_ | ~new_G3036_;
  assign new_G3094_ = ~new_G3066_ | ~new_G3038_;
  assign new_G3095_ = ~new_G3039_;
  assign new_G3099_ = ~new_G3054_;
  assign new_G3100_ = new_G3042_ | new_G3045_ | new_G2851_;
  assign new_G3103_ = ~new_G3042_ & ~new_G3045_ & ~new_G2851_;
  assign new_G3106_ = ~new_G2932_ | ~new_G3067_;
  assign new_G3107_ = ~new_G3082_ | ~new_G3059_;
  assign new_G3110_ = ~new_G3085_ | ~new_G3061_;
  assign new_G3114_ = ~new_G3069_;
  assign new_G3115_ = ~new_G3069_ | ~new_G3010_;
  assign new_G3116_ = ~new_G3072_;
  assign new_G3117_ = ~new_G3072_ | ~new_G3011_;
  assign new_G3118_ = ~new_G3075_;
  assign new_G3119_ = ~new_G3075_ | ~new_G3015_;
  assign new_G3120_ = ~new_G3078_;
  assign new_G3121_ = ~new_G3078_ | ~new_G3016_;
  assign new_G3122_ = ~new_G3089_ | ~new_G3064_;
  assign new_G3126_ = ~new_G3106_ | ~new_G3068_;
  assign new_G3129_ = n2304_lo & new_G3081_;
  assign new_G3132_ = ~new_G3094_;
  assign new_G3135_ = ~new_G3103_;
  assign new_G3136_ = ~new_G2962_ | ~new_G3114_;
  assign new_G3137_ = ~new_G2965_ | ~new_G3116_;
  assign new_G3138_ = ~new_G2968_ | ~new_G3118_;
  assign new_G3139_ = ~new_G2971_ | ~new_G3120_;
  assign new_G3140_ = new_G3086_ & new_G1299_;
  assign new_G3143_ = new_G3086_ & new_G1776_;
  assign new_G3146_ = new_G3090_ & new_G1302_;
  assign new_G3149_ = ~new_G3095_;
  assign new_G3152_ = new_G3090_ & new_G2923_;
  assign new_G3155_ = ~new_G3100_;
  assign new_G3158_ = ~new_G3126_;
  assign new_G3159_ = ~new_G3129_;
  assign new_G3160_ = ~new_G3136_ | ~new_G3115_;
  assign new_G3164_ = ~new_G3137_ | ~new_G3117_;
  assign new_G3165_ = ~new_G3138_ | ~new_G3119_;
  assign new_G3168_ = ~new_G3139_ | ~new_G3121_;
  assign new_G3169_ = ~new_G3132_ | ~new_G3099_;
  assign new_G3170_ = ~new_G3132_;
  assign new_G3171_ = new_G3110_ & new_G1297_;
  assign new_G3174_ = new_G3122_ & new_G1301_;
  assign new_G3177_ = ~new_G3107_;
  assign new_G3180_ = ~new_G3107_;
  assign new_G3183_ = ~new_G3110_;
  assign new_G3186_ = ~new_G3122_;
  assign new_G3189_ = ~new_G3129_ | ~new_G3158_;
  assign new_G3190_ = ~new_G3126_ | ~new_G3159_;
  assign new_G3191_ = ~new_G3168_;
  assign new_G3192_ = ~new_G3149_;
  assign new_G3193_ = ~new_G3152_;
  assign new_G3194_ = ~new_G3054_ | ~new_G3170_;
  assign new_G3195_ = new_G3140_ | new_G3143_ | new_G2842_;
  assign new_G3199_ = ~new_G3140_ & ~new_G3143_ & ~new_G2842_;
  assign new_G3202_ = ~new_G3155_;
  assign new_G3203_ = ~new_G3164_;
  assign new_G3206_ = ~new_G3189_ | ~new_G3190_;
  assign new_G3207_ = ~new_G3177_;
  assign new_G3208_ = ~new_G3177_ | ~new_G3083_;
  assign new_G3209_ = ~new_G3180_;
  assign new_G3210_ = ~new_G3180_ | ~new_G3084_;
  assign new_G3211_ = ~new_G3191_ & ~new_G2986_;
  assign new_G3212_ = new_G3090_ & new_G3122_ & new_G3165_ & new_G2986_;
  assign new_G3213_ = ~new_G3183_;
  assign new_G3214_ = ~new_G3186_;
  assign new_G3215_ = ~new_G3186_ | ~new_G3193_;
  assign new_G3216_ = ~new_G3194_ | ~new_G3169_;
  assign new_G3217_ = new_G3160_ & new_G1298_;
  assign new_G3220_ = new_G3165_ & new_G1300_;
  assign new_G3223_ = new_G3160_ & new_G3039_;
  assign new_G3226_ = ~new_G3199_;
  assign new_G3227_ = new_G3206_ & new_G1353_;
  assign new_G3230_ = ~new_G3048_ | ~new_G3207_;
  assign new_G3231_ = ~new_G3051_ | ~new_G3209_;
  assign new_G3232_ = new_G3211_ | new_G3212_;
  assign new_G3233_ = ~new_G3203_ | ~new_G3192_;
  assign new_G3234_ = ~new_G3203_;
  assign new_G3235_ = ~new_G3152_ | ~new_G3214_;
  assign new_G3236_ = ~new_G3216_;
  assign new_G3237_ = ~new_G3195_;
  assign new_G3240_ = ~new_G3195_;
  assign new_G3243_ = ~new_G3230_ | ~new_G3208_;
  assign new_G3246_ = ~new_G3231_ | ~new_G3210_;
  assign new_G3247_ = ~new_G3223_ | ~new_G3213_;
  assign new_G3248_ = ~new_G3223_;
  assign new_G3249_ = ~new_G3149_ | ~new_G3234_;
  assign new_G3250_ = ~new_G3235_ | ~new_G3215_;
  assign new_G3251_ = new_G3232_ & new_G1778_;
  assign new_G3254_ = new_G3236_ & new_G1782_;
  assign new_G3257_ = new_G1802_ | new_G1524_ | new_G3227_;
  assign new_G3258_ = ~new_G1802_ & ~new_G1524_ & ~new_G3227_;
  assign new_G3259_ = ~new_G3246_;
  assign new_G3260_ = ~new_G3183_ | ~new_G3248_;
  assign new_G3261_ = ~new_G3249_ | ~new_G3233_;
  assign new_G3262_ = new_G3250_ & new_G1780_;
  assign new_G3265_ = ~new_G3237_;
  assign new_G3266_ = ~new_G3240_;
  assign new_G3267_ = ~new_G3258_;
  assign new_G3268_ = ~new_G3259_ & ~new_G3095_;
  assign new_G3269_ = new_G3160_ & new_G3110_ & new_G3243_ & new_G3095_;
  assign new_G3270_ = ~new_G3247_ | ~new_G3260_;
  assign new_G3271_ = ~new_G3261_;
  assign new_G3272_ = new_G3243_ & new_G1296_;
  assign new_G3275_ = new_G3220_ | new_G3251_ | new_G2845_;
  assign new_G3278_ = ~new_G3220_ & ~new_G3251_ & ~new_G2845_;
  assign new_G3281_ = new_G3146_ | new_G3254_ | new_G2848_;
  assign new_G3284_ = ~new_G3146_ & ~new_G3254_ & ~new_G2848_;
  assign new_G3287_ = new_G3268_ | new_G3269_;
  assign new_G3288_ = new_G3270_ & new_G1772_;
  assign new_G3291_ = new_G3271_ & new_G1774_;
  assign new_G3294_ = new_G3174_ | new_G3262_ | new_G2929_;
  assign new_G3297_ = ~new_G3174_ & ~new_G3262_ & ~new_G2929_;
  assign new_G3300_ = ~new_G3278_;
  assign new_G3301_ = ~new_G3284_;
  assign new_G3302_ = new_G3287_ & new_G1770_;
  assign new_G3305_ = ~new_G3281_;
  assign new_G3308_ = ~new_G3275_;
  assign new_G3311_ = ~new_G3297_;
  assign new_G3312_ = new_G3171_ | new_G3288_ | new_G2926_;
  assign new_G3317_ = ~new_G3171_ & ~new_G3288_ & ~new_G2926_;
  assign new_G3320_ = new_G3217_ | new_G3291_ | new_G2839_;
  assign new_G3323_ = ~new_G3217_ & ~new_G3291_ & ~new_G2839_;
  assign new_G3326_ = new_G3103_ & new_G3284_ & new_G3297_ & new_G3278_;
  assign new_G3329_ = ~new_G3294_;
  assign new_G3332_ = new_G3272_ | new_G3302_ | new_G2836_;
  assign new_G3337_ = ~new_G3272_ & ~new_G3302_ & ~new_G2836_;
  assign new_G3340_ = ~new_G3305_ | ~new_G3202_;
  assign new_G3341_ = ~new_G3305_;
  assign new_G3342_ = ~new_G3308_;
  assign new_G3343_ = ~new_G3323_;
  assign new_G3344_ = ~new_G3155_ | ~new_G3341_;
  assign new_G3345_ = ~new_G3329_;
  assign new_G3346_ = ~new_G3329_ | ~new_G3342_;
  assign new_G3347_ = ~new_G3320_;
  assign new_G3350_ = new_G3312_ & new_G884_;
  assign new_G3353_ = ~new_G3312_;
  assign new_G3356_ = ~new_G3340_ | ~new_G3344_;
  assign new_G3359_ = ~new_G3308_ | ~new_G3345_;
  assign new_G3360_ = new_G884_ & new_G3332_;
  assign new_G3363_ = new_G3199_ & new_G3323_ & new_G3317_ & new_G3337_;
  assign new_G3366_ = new_G3317_ & new_G3337_ & new_G887_;
  assign new_G3367_ = ~new_G3332_;
  assign new_G3370_ = ~new_G3359_ | ~new_G3346_;
  assign new_G3373_ = ~new_G3347_;
  assign new_G3376_ = ~new_G3347_;
  assign new_G3379_ = ~new_G3353_;
  assign new_G3380_ = ~new_G3350_;
  assign new_G3383_ = ~new_G3350_;
  assign new_G3386_ = new_G3326_ & new_G3363_;
  assign new_G3387_ = new_G3326_ & new_G3363_;
  assign new_G3388_ = ~new_G3356_;
  assign new_G3391_ = ~new_G3356_;
  assign new_G3394_ = ~new_G3367_;
  assign new_G3395_ = ~new_G3367_ | ~new_G3379_;
  assign new_G3396_ = ~new_G3360_;
  assign new_G3399_ = ~new_G3360_;
  assign new_G3402_ = ~new_G3366_ & ~new_G3387_;
  assign new_G3403_ = ~new_G3373_ | ~new_G3265_;
  assign new_G3404_ = ~new_G3373_;
  assign new_G3405_ = ~new_G3376_ | ~new_G3266_;
  assign new_G3406_ = ~new_G3376_;
  assign new_G3407_ = ~new_G3380_;
  assign new_G3408_ = ~new_G3383_;
  assign new_G3409_ = ~new_G3370_;
  assign new_G3412_ = ~new_G3370_;
  assign new_G3415_ = ~new_G3353_ | ~new_G3394_;
  assign new_G3416_ = n2064_lo & new_G3402_;
  assign new_G3417_ = ~new_G3388_;
  assign new_G3418_ = ~new_G3391_;
  assign new_G3419_ = ~new_G3237_ | ~new_G3404_;
  assign new_G3420_ = ~new_G3240_ | ~new_G3406_;
  assign new_G3421_ = ~new_G3396_;
  assign new_G3422_ = ~new_G3396_ | ~new_G3407_;
  assign new_G3423_ = ~new_G3399_ | ~new_G3408_;
  assign new_G3424_ = ~new_G3399_;
  assign new_G3425_ = ~new_G3395_ | ~new_G3415_;
  assign new_G3428_ = ~new_G3409_ | ~new_G3417_;
  assign new_G3429_ = ~new_G3409_;
  assign new_G3430_ = ~new_G3412_ | ~new_G3418_;
  assign new_G3431_ = ~new_G3412_;
  assign new_G3432_ = ~new_G3403_ | ~new_G3419_;
  assign new_G3436_ = ~new_G3405_ | ~new_G3420_;
  assign new_G3437_ = ~new_G3380_ | ~new_G3421_;
  assign new_G3438_ = ~new_G3383_ | ~new_G3424_;
  assign new_G3439_ = ~new_G3388_ | ~new_G3429_;
  assign new_G3440_ = ~new_G3391_ | ~new_G3431_;
  assign new_G3441_ = ~new_G3436_;
  assign new_G3444_ = ~new_G3425_;
  assign new_G3445_ = ~new_G3437_ | ~new_G3422_;
  assign new_G3448_ = ~new_G3438_ | ~new_G3423_;
  assign new_G3449_ = ~new_G3428_ | ~new_G3439_;
  assign new_G3452_ = ~new_G3430_ | ~new_G3440_;
  assign new_G3453_ = ~new_G3448_;
  assign new_G3456_ = ~new_G3432_;
  assign new_G3459_ = new_G3432_ & new_G3445_ & new_G1436_;
  assign new_G3460_ = new_G3441_ & new_G3445_ & new_G1439_;
  assign new_G3461_ = ~new_G3452_;
  assign new_G3464_ = ~new_G3456_;
  assign new_G3465_ = ~new_G3456_ | ~new_G3444_;
  assign new_G3466_ = new_G3432_ & new_G3453_ & new_G1439_;
  assign new_G3467_ = new_G3441_ & new_G3453_ & new_G1436_;
  assign new_G3468_ = ~new_G3449_;
  assign new_G3471_ = ~new_G3449_;
  assign new_G3474_ = ~new_G3425_ | ~new_G3464_;
  assign new_G3475_ = new_G3467_ | new_G3459_ | new_G3466_ | new_G3460_;
  assign new_G3478_ = ~new_G3461_;
  assign new_G3481_ = ~new_G3461_;
  assign new_G3484_ = ~new_G3474_ | ~new_G3465_;
  assign new_G3487_ = ~new_G3471_;
  assign new_G3488_ = ~new_G3468_;
  assign new_G3489_ = ~new_G3481_;
  assign new_G3490_ = ~new_G3478_;
  assign new_G3491_ = ~new_G3475_;
  assign new_G3494_ = ~new_G3475_;
  assign new_G3497_ = ~new_G3484_;
  assign new_G3500_ = ~new_G3484_;
  assign new_G3503_ = ~new_G3491_ | ~new_G3490_;
  assign new_G3504_ = ~new_G3494_ | ~new_G3489_;
  assign new_G3505_ = ~new_G3494_;
  assign new_G3506_ = ~new_G3491_;
  assign new_G3507_ = ~new_G3497_ | ~new_G3488_;
  assign new_G3508_ = ~new_G3500_ | ~new_G3487_;
  assign new_G3509_ = ~new_G3478_ | ~new_G3506_;
  assign new_G3510_ = ~new_G3481_ | ~new_G3505_;
  assign new_G3511_ = ~new_G3500_;
  assign new_G3512_ = ~new_G3497_;
  assign new_G3513_ = ~new_G3468_ | ~new_G3512_;
  assign new_G3514_ = ~new_G3471_ | ~new_G3511_;
  assign new_G3515_ = ~new_G3509_ | ~new_G3503_;
  assign new_G3516_ = ~new_G3510_ | ~new_G3504_;
  assign new_G3517_ = ~new_G3507_ | ~new_G3513_;
  assign new_G3518_ = ~new_G3508_ | ~new_G3514_;
  assign G3519 = ~new_G928_;
  assign G3520 = ~new_G1004_;
  assign G3521 = ~new_G1786_ | ~new_G1811_;
  assign G3522 = ~new_G2460_ | ~new_G2461_;
  assign G3523 = ~new_G2550_ | ~new_G2551_;
  assign G3524 = new_G2558_ & new_G2552_;
  assign G3525 = ~new_G2675_;
  assign G3526 = new_G2974_ | new_G2943_;
  assign G3527 = new_G3005_ & new_G3030_;
  assign G3528 = new_G3100_ & new_G3135_;
  assign G3529 = new_G3195_ & new_G3226_;
  assign G3530 = new_G3257_ & new_G3267_;
  assign G3531 = new_G3275_ & new_G3300_;
  assign G3532 = new_G3281_ & new_G3301_;
  assign G3533 = new_G3294_ & new_G3311_;
  assign G3534 = new_G3312_ & new_G3312_;
  assign G3535 = new_G3332_ & new_G3332_;
  assign G3536 = new_G3320_ & new_G3343_;
  assign G3537 = ~new_G3386_;
  assign G3538 = ~new_G3416_;
  assign G3539 = new_G3515_ & new_G3516_;
  assign G3540 = ~new_G3517_ | ~new_G3518_;
  assign n1743_li = G1;
  assign n1746_li = n1743_lo;
  assign n1749_li = n1746_lo;
  assign n1752_li = n1749_lo;
  assign n1755_li = G2;
  assign n1758_li = n1755_lo;
  assign n1761_li = n1758_lo;
  assign n1764_li = n1761_lo;
  assign n1767_li = G3;
  assign n1770_li = n1767_lo;
  assign n1773_li = n1770_lo;
  assign n1776_li = n1773_lo;
  assign n1779_li = G4;
  assign n1782_li = n1779_lo;
  assign n1785_li = n1782_lo;
  assign n1788_li = n1785_lo;
  assign n1791_li = G5;
  assign n1794_li = n1791_lo;
  assign n1797_li = n1794_lo;
  assign n1800_li = n1797_lo;
  assign n1803_li = G6;
  assign n1806_li = n1803_lo;
  assign n1809_li = n1806_lo;
  assign n1812_li = n1809_lo;
  assign n1815_li = G7;
  assign n1818_li = n1815_lo;
  assign n1821_li = n1818_lo;
  assign n1824_li = n1821_lo;
  assign n1827_li = G8;
  assign n1830_li = n1827_lo;
  assign n1833_li = n1830_lo;
  assign n1836_li = n1833_lo;
  assign n1839_li = G9;
  assign n1842_li = n1839_lo;
  assign n1845_li = n1842_lo;
  assign n1848_li = n1845_lo;
  assign n1851_li = G10;
  assign n1854_li = n1851_lo;
  assign n1857_li = n1854_lo;
  assign n1860_li = n1857_lo;
  assign n1863_li = G11;
  assign n1866_li = n1863_lo;
  assign n1869_li = n1866_lo;
  assign n1872_li = n1869_lo;
  assign n1875_li = G12;
  assign n1878_li = n1875_lo;
  assign n1881_li = n1878_lo;
  assign n1884_li = n1881_lo;
  assign n1887_li = G13;
  assign n1890_li = n1887_lo;
  assign n1893_li = n1890_lo;
  assign n1896_li = n1893_lo;
  assign n1899_li = G14;
  assign n1902_li = n1899_lo;
  assign n1905_li = n1902_lo;
  assign n1908_li = n1905_lo;
  assign n1911_li = G15;
  assign n1914_li = n1911_lo;
  assign n1917_li = n1914_lo;
  assign n1920_li = n1917_lo;
  assign n1923_li = G16;
  assign n1926_li = n1923_lo;
  assign n1929_li = n1926_lo;
  assign n1932_li = n1929_lo;
  assign n1935_li = G17;
  assign n1938_li = n1935_lo;
  assign n1941_li = n1938_lo;
  assign n1944_li = n1941_lo;
  assign n1947_li = G18;
  assign n1950_li = n1947_lo;
  assign n1953_li = n1950_lo;
  assign n1956_li = n1953_lo;
  assign n1959_li = G19;
  assign n1962_li = n1959_lo;
  assign n1965_li = n1962_lo;
  assign n1968_li = n1965_lo;
  assign n1971_li = G20;
  assign n1974_li = n1971_lo;
  assign n1977_li = n1974_lo;
  assign n1980_li = n1977_lo;
  assign n1983_li = G21;
  assign n1986_li = n1983_lo;
  assign n1989_li = n1986_lo;
  assign n1992_li = n1989_lo;
  assign n1995_li = G22;
  assign n1998_li = n1995_lo;
  assign n2001_li = n1998_lo;
  assign n2004_li = n2001_lo;
  assign n2007_li = G23;
  assign n2010_li = n2007_lo;
  assign n2013_li = n2010_lo;
  assign n2016_li = n2013_lo;
  assign n2019_li = G24;
  assign n2022_li = n2019_lo;
  assign n2025_li = n2022_lo;
  assign n2028_li = n2025_lo;
  assign n2031_li = G25;
  assign n2034_li = n2031_lo;
  assign n2037_li = n2034_lo;
  assign n2040_li = n2037_lo;
  assign n2043_li = G26;
  assign n2046_li = n2043_lo;
  assign n2049_li = n2046_lo;
  assign n2052_li = n2049_lo;
  assign n2055_li = G27;
  assign n2058_li = n2055_lo;
  assign n2061_li = n2058_lo;
  assign n2064_li = n2061_lo;
  assign n2067_li = G28;
  assign n2070_li = n2067_lo;
  assign n2073_li = n2070_lo;
  assign n2076_li = n2073_lo;
  assign n2079_li = G29;
  assign n2082_li = n2079_lo;
  assign n2085_li = n2082_lo;
  assign n2088_li = n2085_lo;
  assign n2091_li = G30;
  assign n2094_li = n2091_lo;
  assign n2097_li = n2094_lo;
  assign n2100_li = n2097_lo;
  assign n2103_li = G31;
  assign n2106_li = n2103_lo;
  assign n2109_li = n2106_lo;
  assign n2112_li = n2109_lo;
  assign n2115_li = G32;
  assign n2118_li = n2115_lo;
  assign n2121_li = n2118_lo;
  assign n2124_li = n2121_lo;
  assign n2127_li = G33;
  assign n2130_li = n2127_lo;
  assign n2133_li = n2130_lo;
  assign n2136_li = n2133_lo;
  assign n2139_li = G34;
  assign n2142_li = n2139_lo;
  assign n2145_li = n2142_lo;
  assign n2148_li = n2145_lo;
  assign n2151_li = G35;
  assign n2154_li = n2151_lo;
  assign n2157_li = n2154_lo;
  assign n2160_li = n2157_lo;
  assign n2163_li = G36;
  assign n2166_li = n2163_lo;
  assign n2169_li = n2166_lo;
  assign n2172_li = n2169_lo;
  assign n2175_li = G37;
  assign n2178_li = n2175_lo;
  assign n2181_li = n2178_lo;
  assign n2184_li = n2181_lo;
  assign n2187_li = G38;
  assign n2190_li = n2187_lo;
  assign n2193_li = n2190_lo;
  assign n2196_li = n2193_lo;
  assign n2199_li = G39;
  assign n2202_li = n2199_lo;
  assign n2205_li = n2202_lo;
  assign n2208_li = n2205_lo;
  assign n2211_li = G40;
  assign n2214_li = n2211_lo;
  assign n2217_li = n2214_lo;
  assign n2220_li = n2217_lo;
  assign n2223_li = G41;
  assign n2226_li = n2223_lo;
  assign n2229_li = n2226_lo;
  assign n2232_li = n2229_lo;
  assign n2235_li = G42;
  assign n2238_li = n2235_lo;
  assign n2241_li = n2238_lo;
  assign n2244_li = n2241_lo;
  assign n2247_li = G43;
  assign n2250_li = n2247_lo;
  assign n2253_li = n2250_lo;
  assign n2256_li = n2253_lo;
  assign n2259_li = G44;
  assign n2262_li = n2259_lo;
  assign n2265_li = n2262_lo;
  assign n2268_li = n2265_lo;
  assign n2271_li = G45;
  assign n2274_li = n2271_lo;
  assign n2277_li = n2274_lo;
  assign n2280_li = n2277_lo;
  assign n2283_li = G46;
  assign n2286_li = n2283_lo;
  assign n2289_li = n2286_lo;
  assign n2292_li = n2289_lo;
  assign n2295_li = G47;
  assign n2298_li = n2295_lo;
  assign n2301_li = n2298_lo;
  assign n2304_li = n2301_lo;
  assign n2307_li = G48;
  assign n2310_li = n2307_lo;
  assign n2313_li = n2310_lo;
  assign n2316_li = n2313_lo;
  assign n2319_li = G49;
  assign n2322_li = n2319_lo;
  assign n2325_li = n2322_lo;
  assign n2328_li = n2325_lo;
  assign n2331_li = G50;
  assign n2334_li = n2331_lo;
  assign n2337_li = n2334_lo;
  assign n2340_li = n2337_lo;
  always @ (posedge clock) begin
    n1743_lo <= n1743_li;
    n1746_lo <= n1746_li;
    n1749_lo <= n1749_li;
    n1752_lo <= n1752_li;
    n1755_lo <= n1755_li;
    n1758_lo <= n1758_li;
    n1761_lo <= n1761_li;
    n1764_lo <= n1764_li;
    n1767_lo <= n1767_li;
    n1770_lo <= n1770_li;
    n1773_lo <= n1773_li;
    n1776_lo <= n1776_li;
    n1779_lo <= n1779_li;
    n1782_lo <= n1782_li;
    n1785_lo <= n1785_li;
    n1788_lo <= n1788_li;
    n1791_lo <= n1791_li;
    n1794_lo <= n1794_li;
    n1797_lo <= n1797_li;
    n1800_lo <= n1800_li;
    n1803_lo <= n1803_li;
    n1806_lo <= n1806_li;
    n1809_lo <= n1809_li;
    n1812_lo <= n1812_li;
    n1815_lo <= n1815_li;
    n1818_lo <= n1818_li;
    n1821_lo <= n1821_li;
    n1824_lo <= n1824_li;
    n1827_lo <= n1827_li;
    n1830_lo <= n1830_li;
    n1833_lo <= n1833_li;
    n1836_lo <= n1836_li;
    n1839_lo <= n1839_li;
    n1842_lo <= n1842_li;
    n1845_lo <= n1845_li;
    n1848_lo <= n1848_li;
    n1851_lo <= n1851_li;
    n1854_lo <= n1854_li;
    n1857_lo <= n1857_li;
    n1860_lo <= n1860_li;
    n1863_lo <= n1863_li;
    n1866_lo <= n1866_li;
    n1869_lo <= n1869_li;
    n1872_lo <= n1872_li;
    n1875_lo <= n1875_li;
    n1878_lo <= n1878_li;
    n1881_lo <= n1881_li;
    n1884_lo <= n1884_li;
    n1887_lo <= n1887_li;
    n1890_lo <= n1890_li;
    n1893_lo <= n1893_li;
    n1896_lo <= n1896_li;
    n1899_lo <= n1899_li;
    n1902_lo <= n1902_li;
    n1905_lo <= n1905_li;
    n1908_lo <= n1908_li;
    n1911_lo <= n1911_li;
    n1914_lo <= n1914_li;
    n1917_lo <= n1917_li;
    n1920_lo <= n1920_li;
    n1923_lo <= n1923_li;
    n1926_lo <= n1926_li;
    n1929_lo <= n1929_li;
    n1932_lo <= n1932_li;
    n1935_lo <= n1935_li;
    n1938_lo <= n1938_li;
    n1941_lo <= n1941_li;
    n1944_lo <= n1944_li;
    n1947_lo <= n1947_li;
    n1950_lo <= n1950_li;
    n1953_lo <= n1953_li;
    n1956_lo <= n1956_li;
    n1959_lo <= n1959_li;
    n1962_lo <= n1962_li;
    n1965_lo <= n1965_li;
    n1968_lo <= n1968_li;
    n1971_lo <= n1971_li;
    n1974_lo <= n1974_li;
    n1977_lo <= n1977_li;
    n1980_lo <= n1980_li;
    n1983_lo <= n1983_li;
    n1986_lo <= n1986_li;
    n1989_lo <= n1989_li;
    n1992_lo <= n1992_li;
    n1995_lo <= n1995_li;
    n1998_lo <= n1998_li;
    n2001_lo <= n2001_li;
    n2004_lo <= n2004_li;
    n2007_lo <= n2007_li;
    n2010_lo <= n2010_li;
    n2013_lo <= n2013_li;
    n2016_lo <= n2016_li;
    n2019_lo <= n2019_li;
    n2022_lo <= n2022_li;
    n2025_lo <= n2025_li;
    n2028_lo <= n2028_li;
    n2031_lo <= n2031_li;
    n2034_lo <= n2034_li;
    n2037_lo <= n2037_li;
    n2040_lo <= n2040_li;
    n2043_lo <= n2043_li;
    n2046_lo <= n2046_li;
    n2049_lo <= n2049_li;
    n2052_lo <= n2052_li;
    n2055_lo <= n2055_li;
    n2058_lo <= n2058_li;
    n2061_lo <= n2061_li;
    n2064_lo <= n2064_li;
    n2067_lo <= n2067_li;
    n2070_lo <= n2070_li;
    n2073_lo <= n2073_li;
    n2076_lo <= n2076_li;
    n2079_lo <= n2079_li;
    n2082_lo <= n2082_li;
    n2085_lo <= n2085_li;
    n2088_lo <= n2088_li;
    n2091_lo <= n2091_li;
    n2094_lo <= n2094_li;
    n2097_lo <= n2097_li;
    n2100_lo <= n2100_li;
    n2103_lo <= n2103_li;
    n2106_lo <= n2106_li;
    n2109_lo <= n2109_li;
    n2112_lo <= n2112_li;
    n2115_lo <= n2115_li;
    n2118_lo <= n2118_li;
    n2121_lo <= n2121_li;
    n2124_lo <= n2124_li;
    n2127_lo <= n2127_li;
    n2130_lo <= n2130_li;
    n2133_lo <= n2133_li;
    n2136_lo <= n2136_li;
    n2139_lo <= n2139_li;
    n2142_lo <= n2142_li;
    n2145_lo <= n2145_li;
    n2148_lo <= n2148_li;
    n2151_lo <= n2151_li;
    n2154_lo <= n2154_li;
    n2157_lo <= n2157_li;
    n2160_lo <= n2160_li;
    n2163_lo <= n2163_li;
    n2166_lo <= n2166_li;
    n2169_lo <= n2169_li;
    n2172_lo <= n2172_li;
    n2175_lo <= n2175_li;
    n2178_lo <= n2178_li;
    n2181_lo <= n2181_li;
    n2184_lo <= n2184_li;
    n2187_lo <= n2187_li;
    n2190_lo <= n2190_li;
    n2193_lo <= n2193_li;
    n2196_lo <= n2196_li;
    n2199_lo <= n2199_li;
    n2202_lo <= n2202_li;
    n2205_lo <= n2205_li;
    n2208_lo <= n2208_li;
    n2211_lo <= n2211_li;
    n2214_lo <= n2214_li;
    n2217_lo <= n2217_li;
    n2220_lo <= n2220_li;
    n2223_lo <= n2223_li;
    n2226_lo <= n2226_li;
    n2229_lo <= n2229_li;
    n2232_lo <= n2232_li;
    n2235_lo <= n2235_li;
    n2238_lo <= n2238_li;
    n2241_lo <= n2241_li;
    n2244_lo <= n2244_li;
    n2247_lo <= n2247_li;
    n2250_lo <= n2250_li;
    n2253_lo <= n2253_li;
    n2256_lo <= n2256_li;
    n2259_lo <= n2259_li;
    n2262_lo <= n2262_li;
    n2265_lo <= n2265_li;
    n2268_lo <= n2268_li;
    n2271_lo <= n2271_li;
    n2274_lo <= n2274_li;
    n2277_lo <= n2277_li;
    n2280_lo <= n2280_li;
    n2283_lo <= n2283_li;
    n2286_lo <= n2286_li;
    n2289_lo <= n2289_li;
    n2292_lo <= n2292_li;
    n2295_lo <= n2295_li;
    n2298_lo <= n2298_li;
    n2301_lo <= n2301_li;
    n2304_lo <= n2304_li;
    n2307_lo <= n2307_li;
    n2310_lo <= n2310_li;
    n2313_lo <= n2313_li;
    n2316_lo <= n2316_li;
    n2319_lo <= n2319_li;
    n2322_lo <= n2322_li;
    n2325_lo <= n2325_li;
    n2328_lo <= n2328_li;
    n2331_lo <= n2331_li;
    n2334_lo <= n2334_li;
    n2337_lo <= n2337_li;
    n2340_lo <= n2340_li;
  end
  initial begin
    n1743_lo <= 1'b0;
    n1746_lo <= 1'b0;
    n1749_lo <= 1'b0;
    n1752_lo <= 1'b0;
    n1755_lo <= 1'b0;
    n1758_lo <= 1'b0;
    n1761_lo <= 1'b0;
    n1764_lo <= 1'b0;
    n1767_lo <= 1'b0;
    n1770_lo <= 1'b0;
    n1773_lo <= 1'b0;
    n1776_lo <= 1'b0;
    n1779_lo <= 1'b0;
    n1782_lo <= 1'b0;
    n1785_lo <= 1'b0;
    n1788_lo <= 1'b0;
    n1791_lo <= 1'b0;
    n1794_lo <= 1'b0;
    n1797_lo <= 1'b0;
    n1800_lo <= 1'b0;
    n1803_lo <= 1'b0;
    n1806_lo <= 1'b0;
    n1809_lo <= 1'b0;
    n1812_lo <= 1'b0;
    n1815_lo <= 1'b0;
    n1818_lo <= 1'b0;
    n1821_lo <= 1'b0;
    n1824_lo <= 1'b0;
    n1827_lo <= 1'b0;
    n1830_lo <= 1'b0;
    n1833_lo <= 1'b0;
    n1836_lo <= 1'b0;
    n1839_lo <= 1'b0;
    n1842_lo <= 1'b0;
    n1845_lo <= 1'b0;
    n1848_lo <= 1'b0;
    n1851_lo <= 1'b0;
    n1854_lo <= 1'b0;
    n1857_lo <= 1'b0;
    n1860_lo <= 1'b0;
    n1863_lo <= 1'b0;
    n1866_lo <= 1'b0;
    n1869_lo <= 1'b0;
    n1872_lo <= 1'b0;
    n1875_lo <= 1'b0;
    n1878_lo <= 1'b0;
    n1881_lo <= 1'b0;
    n1884_lo <= 1'b0;
    n1887_lo <= 1'b0;
    n1890_lo <= 1'b0;
    n1893_lo <= 1'b0;
    n1896_lo <= 1'b0;
    n1899_lo <= 1'b0;
    n1902_lo <= 1'b0;
    n1905_lo <= 1'b0;
    n1908_lo <= 1'b0;
    n1911_lo <= 1'b0;
    n1914_lo <= 1'b0;
    n1917_lo <= 1'b0;
    n1920_lo <= 1'b0;
    n1923_lo <= 1'b0;
    n1926_lo <= 1'b0;
    n1929_lo <= 1'b0;
    n1932_lo <= 1'b0;
    n1935_lo <= 1'b0;
    n1938_lo <= 1'b0;
    n1941_lo <= 1'b0;
    n1944_lo <= 1'b0;
    n1947_lo <= 1'b0;
    n1950_lo <= 1'b0;
    n1953_lo <= 1'b0;
    n1956_lo <= 1'b0;
    n1959_lo <= 1'b0;
    n1962_lo <= 1'b0;
    n1965_lo <= 1'b0;
    n1968_lo <= 1'b0;
    n1971_lo <= 1'b0;
    n1974_lo <= 1'b0;
    n1977_lo <= 1'b0;
    n1980_lo <= 1'b0;
    n1983_lo <= 1'b0;
    n1986_lo <= 1'b0;
    n1989_lo <= 1'b0;
    n1992_lo <= 1'b0;
    n1995_lo <= 1'b0;
    n1998_lo <= 1'b0;
    n2001_lo <= 1'b0;
    n2004_lo <= 1'b0;
    n2007_lo <= 1'b0;
    n2010_lo <= 1'b0;
    n2013_lo <= 1'b0;
    n2016_lo <= 1'b0;
    n2019_lo <= 1'b0;
    n2022_lo <= 1'b0;
    n2025_lo <= 1'b0;
    n2028_lo <= 1'b0;
    n2031_lo <= 1'b0;
    n2034_lo <= 1'b0;
    n2037_lo <= 1'b0;
    n2040_lo <= 1'b0;
    n2043_lo <= 1'b0;
    n2046_lo <= 1'b0;
    n2049_lo <= 1'b0;
    n2052_lo <= 1'b0;
    n2055_lo <= 1'b0;
    n2058_lo <= 1'b0;
    n2061_lo <= 1'b0;
    n2064_lo <= 1'b0;
    n2067_lo <= 1'b0;
    n2070_lo <= 1'b0;
    n2073_lo <= 1'b0;
    n2076_lo <= 1'b0;
    n2079_lo <= 1'b0;
    n2082_lo <= 1'b0;
    n2085_lo <= 1'b0;
    n2088_lo <= 1'b0;
    n2091_lo <= 1'b0;
    n2094_lo <= 1'b0;
    n2097_lo <= 1'b0;
    n2100_lo <= 1'b0;
    n2103_lo <= 1'b0;
    n2106_lo <= 1'b0;
    n2109_lo <= 1'b0;
    n2112_lo <= 1'b0;
    n2115_lo <= 1'b0;
    n2118_lo <= 1'b0;
    n2121_lo <= 1'b0;
    n2124_lo <= 1'b0;
    n2127_lo <= 1'b0;
    n2130_lo <= 1'b0;
    n2133_lo <= 1'b0;
    n2136_lo <= 1'b0;
    n2139_lo <= 1'b0;
    n2142_lo <= 1'b0;
    n2145_lo <= 1'b0;
    n2148_lo <= 1'b0;
    n2151_lo <= 1'b0;
    n2154_lo <= 1'b0;
    n2157_lo <= 1'b0;
    n2160_lo <= 1'b0;
    n2163_lo <= 1'b0;
    n2166_lo <= 1'b0;
    n2169_lo <= 1'b0;
    n2172_lo <= 1'b0;
    n2175_lo <= 1'b0;
    n2178_lo <= 1'b0;
    n2181_lo <= 1'b0;
    n2184_lo <= 1'b0;
    n2187_lo <= 1'b0;
    n2190_lo <= 1'b0;
    n2193_lo <= 1'b0;
    n2196_lo <= 1'b0;
    n2199_lo <= 1'b0;
    n2202_lo <= 1'b0;
    n2205_lo <= 1'b0;
    n2208_lo <= 1'b0;
    n2211_lo <= 1'b0;
    n2214_lo <= 1'b0;
    n2217_lo <= 1'b0;
    n2220_lo <= 1'b0;
    n2223_lo <= 1'b0;
    n2226_lo <= 1'b0;
    n2229_lo <= 1'b0;
    n2232_lo <= 1'b0;
    n2235_lo <= 1'b0;
    n2238_lo <= 1'b0;
    n2241_lo <= 1'b0;
    n2244_lo <= 1'b0;
    n2247_lo <= 1'b0;
    n2250_lo <= 1'b0;
    n2253_lo <= 1'b0;
    n2256_lo <= 1'b0;
    n2259_lo <= 1'b0;
    n2262_lo <= 1'b0;
    n2265_lo <= 1'b0;
    n2268_lo <= 1'b0;
    n2271_lo <= 1'b0;
    n2274_lo <= 1'b0;
    n2277_lo <= 1'b0;
    n2280_lo <= 1'b0;
    n2283_lo <= 1'b0;
    n2286_lo <= 1'b0;
    n2289_lo <= 1'b0;
    n2292_lo <= 1'b0;
    n2295_lo <= 1'b0;
    n2298_lo <= 1'b0;
    n2301_lo <= 1'b0;
    n2304_lo <= 1'b0;
    n2307_lo <= 1'b0;
    n2310_lo <= 1'b0;
    n2313_lo <= 1'b0;
    n2316_lo <= 1'b0;
    n2319_lo <= 1'b0;
    n2322_lo <= 1'b0;
    n2325_lo <= 1'b0;
    n2328_lo <= 1'b0;
    n2331_lo <= 1'b0;
    n2334_lo <= 1'b0;
    n2337_lo <= 1'b0;
    n2340_lo <= 1'b0;
  end
endmodule


