// Benchmark "mymod" written by ABC on Sun Oct 29 19:31:56 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50,
    G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528,
    G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538,
    G3539, G3540  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50;
  output G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528,
    G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538,
    G3539, G3540;
  reg n1836_lo, n1872_lo, n1884_lo, n1911_lo, n1914_lo, n1917_lo, n1923_lo,
    n1926_lo, n1929_lo, n1935_lo, n1938_lo, n1947_lo, n1950_lo, n1959_lo,
    n1962_lo, n1971_lo, n1974_lo, n1983_lo, n1995_lo, n2007_lo, n2019_lo,
    n2031_lo, n2043_lo, n2055_lo, n2064_lo, n2067_lo, n2100_lo, n2112_lo,
    n2124_lo, n2136_lo, n2148_lo, n2160_lo, n2163_lo, n2172_lo, n2175_lo,
    n2184_lo, n2223_lo, n2235_lo, n2238_lo, n2247_lo, n2250_lo, n2259_lo,
    n2262_lo, n2271_lo, n2274_lo, n2283_lo, n2286_lo, n2295_lo, n2298_lo,
    n2304_lo, n2307_lo, n2331_lo, n2334_lo, n2337_lo, n2340_lo, n3241_o2,
    n3242_o2, n3610_o2, n3980_o2, n3968_o2, n4298_o2, n4371_o2, n4413_o2,
    n4418_o2, n4628_o2, n4629_o2, n4633_o2, n4634_o2, n4732_o2, n4733_o2,
    n4884_o2, n4886_o2, n4890_o2, n5011_o2, n5012_o2, n5013_o2, n5014_o2,
    n5015_o2, n5021_o2, n5016_o2, n5026_o2, n4377_o2, n4378_o2, n4389_o2,
    n327_inv, n330_inv, n4398_o2, n4401_o2, n5117_o2, n5115_o2, n5122_o2,
    n5121_o2, n5119_o2, n5116_o2, n5123_o2, n5156_o2, n5167_o2, n4454_o2,
    n4455_o2, n4456_o2, n4505_o2, G742_o2, G727_o2, n4567_o2, n4568_o2,
    n4569_o2, n4571_o2, n4572_o2, n399_inv, n4539_o2, n4651_o2, n4652_o2,
    n4653_o2, G1514_o2, G1823_o2, n4783_o2, n4787_o2, n426_inv, n429_inv,
    n4816_o2, n435_inv, G572_o2, n4919_o2, n4920_o2, n4921_o2, G1048_o2,
    n5041_o2, n5094_o2, n5278_o2, n5301_o2, G2610_o2, G3174_o2, G3146_o2,
    G3217_o2, G3220_o2, G2839_o2, G3251_o2, G3042_o2, G3045_o2, G3262_o2,
    G2845_o2, G2929_o2, G2848_o2, G2851_o2, G3291_o2, G3254_o2, G2666_o2,
    n5099_o2, n5100_o2, n5101_o2, G2558_o2, n5266_o2, n5267_o2, G2759_o2,
    n537_inv, n540_inv, n543_inv, n5292_o2, n5293_o2, n5294_o2, n5295_o2,
    G618_o2, G621_o2, G384_o2, G377_o2, n570_inv, G3171_o2, G2552_o2,
    G3272_o2, G2015_o2, G3294_o2, G3281_o2, G3320_o2, G3275_o2, G3140_o2,
    G2836_o2, G2926_o2, G2842_o2, G3302_o2, G3288_o2, G3143_o2, G3100_o2,
    G2512_o2, n5325_o2, n5326_o2, n5327_o2, n1857_lo_buf_o2,
    n2097_lo_buf_o2, G2669_o2, n642_inv, G568_o2, n648_inv, G565_o2,
    G559_o2, n1821_lo_buf_o2, n1905_lo_buf_o2, n2133_lo_buf_o2,
    n2145_lo_buf_o2, n2157_lo_buf_o2, n2205_lo_buf_o2, n2217_lo_buf_o2,
    G447_o2, G434_o2, G422_o2, G461_o2, G3312_o2, G3332_o2, G3195_o2,
    G2607_o2, n702_inv, G1005_o2, G1008_o2, n2001_lo_buf_o2,
    n2169_lo_buf_o2, n2229_lo_buf_o2, n2301_lo_buf_o2, n723_inv, G2947_o2,
    n2013_lo_buf_o2, n2025_lo_buf_o2, n2037_lo_buf_o2, n2049_lo_buf_o2,
    n2181_lo_buf_o2, n744_inv, n747_inv, n750_inv, n753_inv, G3350_o2,
    G3360_o2, G3373_o2, G3237_o2, G2773_o2, G1733_o2, G1738_o2, G1751_o2,
    G2216_o2, G2219_o2, n786_inv, n789_inv, G787_o2, G2823_o2, G2796_o2,
    G875_o2, G2208_o2, G2211_o2, n1989_lo_buf_o2, n2061_lo_buf_o2,
    n2313_lo_buf_o2, G2232_o2, G1725_o2, G1764_o2, G2356_o2, G2359_o2,
    G1180_o2, G1756_o2, G2441_o2, G2887_o2, G2991_o2, n849_inv, n852_inv,
    n855_inv, n858_inv, n861_inv, G2805_o2, G2906_o2, G2833_o2, n873_inv,
    G3353_o2, G3367_o2, G3346_o2, G3340_o2, G3376_o2, G3359_o2, G3240_o2,
    G3344_o2, G2880_o2, G2939_o2, G2248_o2, G2251_o2, G2021_o2, G3383_o2,
    G3399_o2, G3404_o2, G3265_o2, G2866_o2, G2999_o2, G736_o2, G739_o2,
    G1200_o2, G1203_o2, G3027_o2, G1463_o2, G1460_o2, G3012_o2, G1574_o2,
    G1646_o2, G1592_o2, G1664_o2, G1547_o2, G1619_o2, G1556_o2, G1628_o2,
    G1583_o2, G1655_o2, G1529_o2, G1601_o2, G1538_o2, G1610_o2, G1565_o2,
    G1637_o2, G2437_o2, n1008_inv, n1785_lo_buf_o2, n1845_lo_buf_o2,
    n1893_lo_buf_o2, n1941_lo_buf_o2, n1953_lo_buf_o2, n1965_lo_buf_o2,
    n1977_lo_buf_o2, n2241_lo_buf_o2, n2253_lo_buf_o2, n2265_lo_buf_o2,
    n2277_lo_buf_o2, n2289_lo_buf_o2, G519_o2, n1050_inv, n1053_inv,
    n1056_inv, G1318_o2, n1062_inv, G593_o2, n1068_inv, n1071_inv,
    n1074_inv, G2284_o2, G2580_o2, G2302_o2, G2598_o2, G2497_o2, G2651_o2,
    G2296_o2, G2308_o2, G2592_o2, G2604_o2, G2902_o2, G2975_o2, G2962_o2,
    G3069_o2, G2018_o2, G1176_o2, G1189_o2, G3066_o2, G3137_o2, G3038_o2,
    G3117_o2, G2384_o2, G2472_o2, G772_o2, G935_o2, G2923_o2, G2971_o2,
    G2980_o2, G3039_o2, G2388_o2, G2287_o2, G3024_o2, G2916_o2, n1176_inv,
    G3035_o2, G3107_o2, G1023_o2, G1024_o2, G1311_o2, G1312_o2, G3063_o2,
    G1520_o2, G1519_o2, G3078_o2, G2038_o2, G1848_o2, G1864_o2, G1872_o2,
    G1880_o2, G1888_o2, G1912_o2, G1928_o2, G1936_o2, G1944_o2, G1952_o2,
    G1850_o2, G1866_o2, G1874_o2, G1882_o2, G1890_o2, G1914_o2, G1930_o2,
    G1938_o2, G1946_o2, G1954_o2, G1845_o2, G1861_o2, G1869_o2, G1877_o2,
    G1885_o2, G1909_o2, G1925_o2, G1933_o2, G1941_o2, G1949_o2, G1846_o2,
    G1862_o2, G1870_o2, G1878_o2, G1886_o2, G1910_o2, G1926_o2, G1934_o2,
    G1942_o2, G1950_o2, G1849_o2, G1865_o2, G1873_o2, G1881_o2, G1889_o2,
    G1913_o2, G1929_o2, G1937_o2, G1945_o2, G1953_o2, G1843_o2, G1859_o2,
    G1867_o2, G1875_o2, G1883_o2, G1907_o2, G1923_o2, G1931_o2, G1939_o2,
    G1947_o2, G1844_o2, G1860_o2, G1868_o2, G1876_o2, G1884_o2, G1908_o2,
    G1924_o2, G1932_o2, G1940_o2, G1948_o2, G1847_o2, G1863_o2, G1871_o2,
    G1879_o2, G1887_o2, G1911_o2, G1927_o2, G1935_o2, G1943_o2, G1951_o2,
    G2444_o2, G2451_o2, G2502_o2, G2507_o2, n1464_inv, G2583_o2,
    n1797_lo_buf_o2, n1833_lo_buf_o2, n1881_lo_buf_o2, n1479_inv,
    n1482_inv, n1485_inv, G615_o2, G2254_o2, G2255_o2, G2027_o2, G2393_o2,
    G527_o2, G594_o2, G1689_o2, G1693_o2, G2281_o2, G2014_o2, G2459_o2,
    G2561_o2, G2533_o2, n1749_lo_buf_o2, n1761_lo_buf_o2, n1773_lo_buf_o2,
    n1809_lo_buf_o2, G1955_o2, G1958_o2, G2562_o2, G2398_o2, n1554_inv,
    n1557_inv, G2577_o2, G2627_o2, G654_o2, G660_o2, G831_o2, G919_o2,
    G925_o2, n1815_lo_buf_o2, n1899_lo_buf_o2, n2079_lo_buf_o2,
    n2127_lo_buf_o2, n2139_lo_buf_o2, n2151_lo_buf_o2, n2187_lo_buf_o2,
    n2199_lo_buf_o2, n2211_lo_buf_o2, G533_o2, n1854_lo_buf_o2,
    n2094_lo_buf_o2, G667_o2, G874_o2, G851_o2, G1127_o2, n1869_lo_buf_o2,
    n2109_lo_buf_o2, n2121_lo_buf_o2, G477_o2, G491_o2, G501_o2, G786_o2,
    G791_o2, G1126_o2, G1052_o2, G1054_o2;
  wire new_n1131_, new_n1133_, new_n1135_, new_n1136_, new_n1137_,
    new_n1139_, new_n1141_, new_n1143_, new_n1145_, new_n1147_, new_n1149_,
    new_n1151_, new_n1153_, new_n1155_, new_n1157_, new_n1159_, new_n1161_,
    new_n1163_, new_n1165_, new_n1167_, new_n1169_, new_n1171_, new_n1173_,
    new_n1175_, new_n1177_, new_n1179_, new_n1181_, new_n1183_, new_n1185_,
    new_n1187_, new_n1189_, new_n1191_, new_n1193_, new_n1195_, new_n1197_,
    new_n1199_, new_n1201_, new_n1203_, new_n1205_, new_n1207_, new_n1209_,
    new_n1211_, new_n1213_, new_n1215_, new_n1217_, new_n1219_, new_n1221_,
    new_n1223_, new_n1225_, new_n1227_, new_n1229_, new_n1231_, new_n1232_,
    new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1239_, new_n1242_,
    new_n1243_, new_n1245_, new_n1248_, new_n1249_, new_n1251_, new_n1253_,
    new_n1255_, new_n1257_, new_n1259_, new_n1261_, new_n1263_, new_n1265_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1281_, new_n1284_, new_n1286_, new_n1288_, new_n1290_,
    new_n1292_, new_n1294_, new_n1295_, new_n1296_, new_n1298_, new_n1299_,
    new_n1302_, new_n1303_, new_n1305_, new_n1307_, new_n1309_, new_n1311_,
    new_n1313_, new_n1315_, new_n1317_, new_n1319_, new_n1321_, new_n1323_,
    new_n1325_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1335_, new_n1337_, new_n1339_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1346_, new_n1348_,
    new_n1350_, new_n1351_, new_n1353_, new_n1356_, new_n1357_, new_n1359_,
    new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_,
    new_n1368_, new_n1369_, new_n1370_, new_n1372_, new_n1374_, new_n1375_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1385_, new_n1386_, new_n1387_, new_n1389_, new_n1392_,
    new_n1393_, new_n1395_, new_n1397_, new_n1398_, new_n1399_, new_n1401_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1409_,
    new_n1411_, new_n1413_, new_n1415_, new_n1417_, new_n1419_, new_n1420_,
    new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1427_,
    new_n1429_, new_n1431_, new_n1433_, new_n1434_, new_n1436_, new_n1437_,
    new_n1439_, new_n1441_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1465_, new_n1467_, new_n1468_,
    new_n1469_, new_n1470_, new_n1471_, new_n1473_, new_n1474_, new_n1475_,
    new_n1476_, new_n1477_, new_n1479_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1493_, new_n1495_, new_n1497_, new_n1499_,
    new_n1501_, new_n1503_, new_n1505_, new_n1508_, new_n1509_, new_n1511_,
    new_n1513_, new_n1515_, new_n1517_, new_n1519_, new_n1521_, new_n1523_,
    new_n1524_, new_n1525_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_,
    new_n1538_, new_n1539_, new_n1541_, new_n1543_, new_n1545_, new_n1547_,
    new_n1549_, new_n1550_, new_n1551_, new_n1553_, new_n1554_, new_n1555_,
    new_n1556_, new_n1558_, new_n1560_, new_n1561_, new_n1562_, new_n1563_,
    new_n1565_, new_n1567_, new_n1569_, new_n1570_, new_n1571_, new_n1573_,
    new_n1575_, new_n1577_, new_n1579_, new_n1581_, new_n1583_, new_n1585_,
    new_n1587_, new_n1589_, new_n1591_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1611_, new_n1613_, new_n1615_, new_n1617_, new_n1619_,
    new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_,
    new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1631_, new_n1633_,
    new_n1634_, new_n1635_, new_n1638_, new_n1639_, new_n1641_, new_n1643_,
    new_n1645_, new_n1647_, new_n1649_, new_n1651_, new_n1653_, new_n1655_,
    new_n1657_, new_n1658_, new_n1659_, new_n1661_, new_n1662_, new_n1663_,
    new_n1665_, new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_,
    new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_,
    new_n1679_, new_n1681_, new_n1683_, new_n1685_, new_n1686_, new_n1687_,
    new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_,
    new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_,
    new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_,
    new_n1707_, new_n1709_, new_n1711_, new_n1713_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1723_,
    new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_,
    new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_,
    new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_,
    new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_,
    new_n1755_, new_n1756_, new_n1757_, new_n1759_, new_n1761_, new_n1763_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_,
    new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_,
    new_n1802_, new_n1804_, new_n1805_, new_n1807_, new_n1809_, new_n1811_,
    new_n1812_, new_n1814_, new_n1816_, new_n1817_, new_n1818_, new_n1819_,
    new_n1821_, new_n1823_, new_n1825_, new_n1828_, new_n1830_, new_n1831_,
    new_n1833_, new_n1836_, new_n1838_, new_n1839_, new_n1841_, new_n1843_,
    new_n1845_, new_n1847_, new_n1849_, new_n1851_, new_n1852_, new_n1853_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1862_, new_n1864_, new_n1866_, new_n1867_, new_n1868_, new_n1869_,
    new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_,
    new_n1876_, new_n1877_, new_n1879_, new_n1880_, new_n1881_, new_n1882_,
    new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1888_, new_n1889_,
    new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_,
    new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_,
    new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_,
    new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_,
    new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_,
    new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_,
    new_n1926_, new_n1927_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1949_, new_n1950_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1974_, new_n1976_, new_n1978_, new_n1979_,
    new_n1980_, new_n1981_, new_n1983_, new_n1985_, new_n1986_, new_n1987_,
    new_n1989_, new_n1991_, new_n1994_, new_n1995_, new_n1998_, new_n1999_,
    new_n2001_, new_n2004_, new_n2005_, new_n2008_, new_n2009_, new_n2011_,
    new_n2014_, new_n2015_, new_n2018_, new_n2019_, new_n2021_, new_n2024_,
    new_n2025_, new_n2028_, new_n2030_, new_n2032_, new_n2033_, new_n2036_,
    new_n2037_, new_n2040_, new_n2042_, new_n2043_, new_n2046_, new_n2047_,
    new_n2049_, new_n2051_, new_n2054_, new_n2055_, new_n2058_, new_n2059_,
    new_n2061_, new_n2064_, new_n2065_, new_n2068_, new_n2070_, new_n2072_,
    new_n2073_, new_n2076_, new_n2077_, new_n2080_, new_n2082_, new_n2083_,
    new_n2086_, new_n2087_, new_n2089_, new_n2091_, new_n2094_, new_n2095_,
    new_n2098_, new_n2099_, new_n2101_, new_n2104_, new_n2105_, new_n2108_,
    new_n2109_, new_n2111_, new_n2114_, new_n2115_, new_n2118_, new_n2119_,
    new_n2121_, new_n2124_, new_n2125_, new_n2128_, new_n2129_, new_n2131_,
    new_n2134_, new_n2135_, new_n2138_, new_n2139_, new_n2141_, new_n2144_,
    new_n2145_, new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_,
    new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2159_,
    new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_,
    new_n2166_, new_n2167_, new_n2169_, new_n2171_, new_n2173_, new_n2174_,
    new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_,
    new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_,
    new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_,
    new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_,
    new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_,
    new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_,
    new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_,
    new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_,
    new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_,
    new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_,
    new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_,
    new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_, new_n2246_,
    new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_,
    new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_,
    new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_,
    new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_,
    new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_,
    new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_,
    new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_,
    new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_,
    new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_,
    new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_,
    new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_,
    new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_,
    new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_,
    new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_,
    new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_,
    new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_,
    new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_,
    new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_, new_n2360_,
    new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_,
    new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_,
    new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_,
    new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_,
    new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_,
    new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_,
    new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_,
    new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_,
    new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_,
    new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_,
    new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_,
    new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_,
    new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_,
    new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_,
    new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_,
    new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_,
    new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_,
    new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_,
    new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_,
    new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_,
    new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_,
    new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_,
    new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_,
    new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_, new_n2504_,
    new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_, new_n2510_,
    new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_, new_n2516_,
    new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_, new_n2522_,
    new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_, new_n2528_,
    new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_, new_n2534_,
    new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_, new_n2540_,
    new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_, new_n2546_,
    new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_, new_n2552_,
    new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_, new_n2558_,
    new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_, new_n2564_,
    new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_,
    new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_,
    new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_,
    new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_,
    new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_,
    new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_, new_n2600_,
    new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_, new_n2606_,
    new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_, new_n2612_,
    new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_,
    new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2623_, new_n2624_,
    new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_, new_n2630_,
    new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_, new_n2636_,
    new_n2637_, new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_,
    new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_,
    new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2654_,
    new_n2655_, new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_,
    new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_,
    new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_,
    new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_,
    new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_,
    new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_,
    new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_,
    new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_,
    new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_,
    new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_,
    new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_,
    new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_,
    new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_,
    new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_,
    new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_,
    new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_,
    new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_,
    new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_,
    new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_,
    new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_,
    new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_,
    new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_,
    new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_,
    new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_,
    new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_,
    new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_,
    new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_,
    new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_,
    new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_,
    new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_,
    new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_,
    new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_,
    new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_,
    new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_,
    new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_,
    new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_,
    new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_,
    new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_,
    new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_,
    new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_,
    new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_,
    new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_,
    new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_,
    new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_,
    new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_,
    new_n2925_, new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_,
    new_n2931_, new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_,
    new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_,
    new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_,
    new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_,
    new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_,
    new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_,
    new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_,
    new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_,
    new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_,
    new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_,
    new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_,
    new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_,
    new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_,
    new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_,
    new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3019_, new_n3020_,
    new_n3021_, new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_,
    new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_,
    new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_,
    new_n3039_, new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_,
    new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_,
    new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_,
    new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_,
    new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_,
    new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_,
    new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_,
    new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_,
    new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_,
    new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_,
    new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_,
    new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_,
    new_n3111_, new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_,
    new_n3117_, new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_,
    new_n3123_, new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_,
    new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_,
    new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_,
    new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_,
    new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_,
    new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_,
    new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_,
    new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_,
    new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_,
    new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_,
    new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_,
    new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_,
    new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_,
    new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_,
    new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_,
    new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_,
    new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_,
    new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_,
    new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_,
    new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_,
    new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_,
    new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_,
    new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_,
    new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_,
    new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_,
    new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_,
    new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_,
    new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_,
    new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_,
    new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_,
    new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_,
    new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_,
    new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_,
    new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_,
    new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_,
    new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_,
    new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_,
    new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_,
    new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_,
    new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_,
    new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_,
    new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_,
    new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_,
    new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_,
    new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_,
    new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_,
    new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_,
    new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_,
    new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_,
    new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_,
    new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_,
    new_n3429_, new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_,
    new_n3435_, new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_,
    new_n3441_, new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_,
    new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_,
    new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_,
    new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_,
    new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_,
    new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_,
    new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_,
    new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_,
    new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_,
    new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_,
    new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_,
    new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_,
    new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_,
    new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_,
    new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_,
    new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_,
    new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_,
    new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_, new_n3548_,
    new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_,
    new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_,
    new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_,
    new_n3567_, new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_,
    new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_,
    new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_,
    new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_,
    new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_,
    new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_,
    new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_,
    new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_,
    new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_,
    new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_,
    new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_,
    new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_,
    new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_,
    new_n3645_, new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_,
    new_n3651_, new_n3652_, new_n3653_, new_n3654_, new_n3655_, new_n3656_,
    new_n3657_, new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_,
    new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_,
    new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_,
    new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_,
    new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_,
    new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_,
    new_n3693_, new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_,
    new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_,
    new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_, new_n3710_,
    new_n3711_, new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_,
    new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_,
    new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_,
    new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_,
    new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3739_, new_n3740_,
    new_n3741_, new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_,
    new_n3747_, new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_,
    new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_,
    new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_,
    new_n3765_, new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_,
    new_n3771_, new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_,
    new_n3777_, new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_,
    new_n3783_, new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_,
    new_n3789_, new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_,
    new_n3795_, new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_,
    new_n3801_, new_n3802_, new_n3803_, new_n3804_, new_n3805_, new_n3806_,
    new_n3807_, new_n3808_, new_n3809_, new_n3810_, new_n3811_, new_n4363_,
    new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_,
    new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_, new_n4375_,
    new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_, new_n4381_,
    new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_,
    new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_, new_n4393_,
    new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_, new_n4399_,
    new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_, new_n4405_,
    new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_,
    new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_,
    new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_,
    new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_,
    new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_,
    new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_,
    new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_,
    new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_,
    new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_,
    new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_,
    new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_,
    new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_,
    new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_,
    new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_,
    new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_,
    new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_,
    new_n4502_, new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_,
    new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_,
    new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_,
    new_n4520_, new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_,
    new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_,
    new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_,
    new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_,
    new_n4544_, new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_,
    new_n4550_, new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_,
    new_n4556_, new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_,
    new_n4562_, new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_,
    new_n4568_, new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_,
    new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_,
    new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_,
    new_n4586_, new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_,
    new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_,
    new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4603_,
    new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4609_,
    new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_,
    new_n4616_, new_n4617_, new_n4618_, new_n4619_, new_n4620_, new_n4621_,
    new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_, new_n4627_,
    new_n4628_, new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_,
    new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_,
    new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_,
    new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_,
    new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_,
    new_n4658_, new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_,
    new_n4664_, new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_,
    new_n4670_, new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_,
    new_n4676_, new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_,
    new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_, new_n4687_,
    new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_, new_n4693_,
    new_n4694_, new_n4695_, new_n4696_, new_n4697_, new_n4698_, new_n4699_,
    new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_, new_n4705_,
    new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_,
    new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_,
    new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4722_, new_n4723_,
    new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_,
    new_n4730_, new_n4731_, new_n4732_, new_n4733_, new_n4734_, new_n4735_,
    new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_,
    new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_,
    new_n4748_, new_n4749_, new_n4750_, new_n4751_, new_n4752_, new_n4753_,
    new_n4754_, new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_,
    new_n4760_, new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_,
    new_n4766_, new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_,
    new_n4772_, new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_,
    new_n4778_, new_n4779_, new_n4780_, new_n4781_, new_n4782_, new_n4783_,
    new_n4784_, new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_,
    new_n4790_, new_n4791_, new_n4792_, new_n4793_, new_n4794_, new_n4795_,
    new_n4796_, new_n4797_, new_n4798_, new_n4799_, new_n4800_, new_n4801_,
    new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_,
    new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_, new_n4813_,
    new_n4814_, new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_,
    new_n4820_, new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_,
    new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_,
    new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_,
    new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_, new_n4843_,
    new_n4844_, new_n4845_, new_n4846_, new_n4847_, new_n4848_, new_n4849_,
    new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_, new_n4855_,
    new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_,
    new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_,
    new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_,
    new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4879_,
    new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_,
    new_n4886_, new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_,
    new_n4892_, new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_,
    new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_,
    new_n4904_, new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_,
    new_n4910_, new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_,
    new_n4916_, new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_,
    new_n4922_, new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_,
    new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_,
    new_n4934_, new_n4935_, new_n4936_, new_n4937_, new_n4938_, new_n4939_,
    new_n4940_, new_n4941_, new_n4942_, new_n4943_, new_n4944_, new_n4945_,
    new_n4946_, new_n4947_, new_n4948_, new_n4949_, new_n4950_, new_n4951_,
    new_n4952_, new_n4953_, new_n4954_, new_n4955_, new_n4956_, new_n4957_,
    new_n4958_, new_n4959_, new_n4960_, new_n4961_, new_n4962_, new_n4963_,
    new_n4964_, new_n4965_, new_n4966_, new_n4967_, new_n4968_, new_n4969_,
    new_n4970_, new_n4971_, new_n4972_, new_n4973_, new_n4974_, new_n4975_,
    new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_, new_n4981_,
    new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_, new_n4987_,
    new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_, new_n4993_,
    new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_, new_n4999_,
    new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_, new_n5005_,
    new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_, new_n5011_,
    new_n5012_, new_n5013_, new_n5014_, new_n5015_, new_n5016_, new_n5017_,
    new_n5018_, new_n5019_, new_n5020_, new_n5021_, new_n5022_, new_n5023_,
    new_n5024_, new_n5025_, new_n5026_, new_n5027_, new_n5028_, new_n5029_,
    new_n5030_, new_n5031_, new_n5032_, new_n5033_, new_n5034_, new_n5035_,
    new_n5036_, new_n5037_, new_n5038_, new_n5039_, new_n5040_, new_n5041_,
    new_n5042_, new_n5043_, new_n5044_, new_n5045_, new_n5046_, new_n5047_,
    new_n5048_, new_n5049_, new_n5050_, new_n5051_, new_n5052_, new_n5053_,
    new_n5054_, new_n5055_, new_n5056_, new_n5057_, new_n5058_, new_n5059_,
    new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_, new_n5065_,
    new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5070_, new_n5071_,
    new_n5072_, new_n5073_, new_n5074_, new_n5075_, new_n5076_, new_n5077_,
    new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_, new_n5083_,
    new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_, new_n5089_,
    new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_, new_n5095_,
    new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_, new_n5101_,
    new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_,
    new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_, new_n5113_,
    new_n5114_, new_n5115_, new_n5116_, new_n5117_, new_n5118_, new_n5119_,
    new_n5120_, new_n5121_, new_n5122_, new_n5123_, new_n5124_, new_n5125_,
    new_n5126_, new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_,
    new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_, new_n5137_,
    new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_, new_n5143_,
    new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_, new_n5149_,
    new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_, new_n5155_,
    new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_, new_n5161_,
    new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_, new_n5167_,
    new_n5168_, new_n5169_, new_n5170_, new_n5171_, new_n5172_, new_n5173_,
    new_n5174_, new_n5175_, new_n5176_, new_n5177_, new_n5178_, new_n5179_,
    new_n5180_, new_n5181_, new_n5182_, new_n5183_, new_n5184_, new_n5185_,
    new_n5186_, new_n5187_, new_n5188_, new_n5189_, new_n5190_, new_n5191_,
    new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_, new_n5197_,
    new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_, new_n5203_,
    new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_, new_n5209_,
    new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_, new_n5215_,
    new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_, new_n5221_,
    new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_, new_n5227_,
    new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_, new_n5233_,
    new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_, new_n5239_,
    new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_, new_n5245_,
    new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_, new_n5251_,
    new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_, new_n5257_,
    new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_, new_n5263_,
    new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_, new_n5269_,
    new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_, new_n5275_,
    new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_, new_n5281_,
    new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_, new_n5287_,
    new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_, new_n5293_,
    new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_, new_n5299_,
    new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_, new_n5305_,
    new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_, new_n5311_,
    new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_, new_n5317_,
    new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_, new_n5323_,
    new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_, new_n5329_,
    new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_, new_n5335_,
    new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_, new_n5341_,
    new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_, new_n5347_,
    new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_, new_n5353_,
    new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_,
    new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_,
    new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_, new_n5371_,
    new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_,
    new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_,
    new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_,
    new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_,
    new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_,
    new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_,
    new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_,
    new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_, new_n5419_,
    new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_,
    new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_,
    new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_, new_n5437_,
    new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_,
    new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_,
    new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_, new_n5455_,
    new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_,
    new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_,
    new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_,
    new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_, new_n5479_,
    new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_,
    new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_,
    new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_, new_n5497_,
    new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_,
    new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_,
    new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_, new_n5515_,
    new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_, new_n5521_,
    new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_, new_n5527_,
    new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_, new_n5533_,
    new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_,
    new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_, new_n5545_,
    new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_,
    new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_,
    new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_,
    new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_,
    new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_,
    new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_,
    new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_,
    new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_,
    new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_,
    new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_,
    new_n5606_, new_n5607_, new_n5608_, new_n5609_, n1836_li, n1872_li,
    n1884_li, n1911_li, n1914_li, n1917_li, n1923_li, n1926_li, n1929_li,
    n1935_li, n1938_li, n1947_li, n1950_li, n1959_li, n1962_li, n1971_li,
    n1974_li, n1983_li, n1995_li, n2007_li, n2019_li, n2031_li, n2043_li,
    n2055_li, n2064_li, n2067_li, n2100_li, n2112_li, n2124_li, n2136_li,
    n2148_li, n2160_li, n2163_li, n2172_li, n2175_li, n2184_li, n2223_li,
    n2235_li, n2238_li, n2247_li, n2250_li, n2259_li, n2262_li, n2271_li,
    n2274_li, n2283_li, n2286_li, n2295_li, n2298_li, n2304_li, n2307_li,
    n2331_li, n2334_li, n2337_li, n2340_li, n3241_i2, n3242_i2, n3610_i2,
    n3980_i2, n3968_i2, n4298_i2, n4371_i2, n4413_i2, n4418_i2, n4628_i2,
    n4629_i2, n4633_i2, n4634_i2, n4732_i2, n4733_i2, n4884_i2, n4886_i2,
    n4890_i2, n5011_i2, n5012_i2, n5013_i2, n5014_i2, n5015_i2, n5021_i2,
    n5016_i2, n5026_i2, n4377_i2, n4378_i2, n4389_i2, n4390_i2, n4391_i2,
    n4398_i2, n4401_i2, n5117_i2, n5115_i2, n5122_i2, n5121_i2, n5119_i2,
    n5116_i2, n5123_i2, n5156_i2, n5167_i2, n4454_i2, n4455_i2, n4456_i2,
    n4505_i2, G742_i2, G727_i2, n4567_i2, n4568_i2, n4569_i2, n4571_i2,
    n4572_i2, n4537_i2, n4539_i2, n4651_i2, n4652_i2, n4653_i2, G1514_i2,
    G1823_i2, n4783_i2, n4787_i2, n4808_i2, n4815_i2, n4816_i2, n4822_i2,
    G572_i2, n4919_i2, n4920_i2, n4921_i2, G1048_i2, n5041_i2, n5094_i2,
    n5278_i2, n5301_i2, G2610_i2, G3174_i2, G3146_i2, G3217_i2, G3220_i2,
    G2839_i2, G3251_i2, G3042_i2, G3045_i2, G3262_i2, G2845_i2, G2929_i2,
    G2848_i2, G2851_i2, G3291_i2, G3254_i2, G2666_i2, n5099_i2, n5100_i2,
    n5101_i2, G2558_i2, n5266_i2, n5267_i2, G2759_i2, n5269_i2, n5270_i2,
    n5271_i2, n5292_i2, n5293_i2, n5294_i2, n5295_i2, G618_i2, G621_i2,
    G384_i2, G377_i2, G400_i2, G3171_i2, G2552_i2, G3272_i2, G2015_i2,
    G3294_i2, G3281_i2, G3320_i2, G3275_i2, G3140_i2, G2836_i2, G2926_i2,
    G2842_i2, G3302_i2, G3288_i2, G3143_i2, G3100_i2, G2512_i2, n5325_i2,
    n5326_i2, n5327_i2, n1857_lo_buf_i2, n2097_lo_buf_i2, G2669_i2,
    G552_i2, G568_i2, G530_i2, G565_i2, G559_i2, n1821_lo_buf_i2,
    n1905_lo_buf_i2, n2133_lo_buf_i2, n2145_lo_buf_i2, n2157_lo_buf_i2,
    n2205_lo_buf_i2, n2217_lo_buf_i2, G447_i2, G434_i2, G422_i2, G461_i2,
    G3312_i2, G3332_i2, G3195_i2, G2607_i2, G2799_i2, G1005_i2, G1008_i2,
    n2001_lo_buf_i2, n2169_lo_buf_i2, n2229_lo_buf_i2, n2301_lo_buf_i2,
    G2816_i2, G2947_i2, n2013_lo_buf_i2, n2025_lo_buf_i2, n2037_lo_buf_i2,
    n2049_lo_buf_i2, n2181_lo_buf_i2, G546_i2, G480_i2, G492_i2, G540_i2,
    G3350_i2, G3360_i2, G3373_i2, G3237_i2, G2773_i2, G1733_i2, G1738_i2,
    G1751_i2, G2216_i2, G2219_i2, G381_i2, G397_i2, G787_i2, G2823_i2,
    G2796_i2, G875_i2, G2208_i2, G2211_i2, n1989_lo_buf_i2,
    n2061_lo_buf_i2, n2313_lo_buf_i2, G2232_i2, G1725_i2, G1764_i2,
    G2356_i2, G2359_i2, G1180_i2, G1756_i2, G2441_i2, G2887_i2, G2991_i2,
    G470_i2, G484_i2, G496_i2, G353_i2, G363_i2, G2805_i2, G2906_i2,
    G2833_i2, G1012_i2, G3353_i2, G3367_i2, G3346_i2, G3340_i2, G3376_i2,
    G3359_i2, G3240_i2, G3344_i2, G2880_i2, G2939_i2, G2248_i2, G2251_i2,
    G2021_i2, G3383_i2, G3399_i2, G3404_i2, G3265_i2, G2866_i2, G2999_i2,
    G736_i2, G739_i2, G1200_i2, G1203_i2, G3027_i2, G1463_i2, G1460_i2,
    G3012_i2, G1574_i2, G1646_i2, G1592_i2, G1664_i2, G1547_i2, G1619_i2,
    G1556_i2, G1628_i2, G1583_i2, G1655_i2, G1529_i2, G1601_i2, G1538_i2,
    G1610_i2, G1565_i2, G1637_i2, G2437_i2, G2518_i2, n1785_lo_buf_i2,
    n1845_lo_buf_i2, n1893_lo_buf_i2, n1941_lo_buf_i2, n1953_lo_buf_i2,
    n1965_lo_buf_i2, n1977_lo_buf_i2, n2241_lo_buf_i2, n2253_lo_buf_i2,
    n2265_lo_buf_i2, n2277_lo_buf_i2, n2289_lo_buf_i2, G519_i2, G388_i2,
    G438_i2, G368_i2, G1318_i2, G425_i2, G593_i2, G413_i2, G404_i2,
    G451_i2, G2284_i2, G2580_i2, G2302_i2, G2598_i2, G2497_i2, G2651_i2,
    G2296_i2, G2308_i2, G2592_i2, G2604_i2, G2902_i2, G2975_i2, G2962_i2,
    G3069_i2, G2018_i2, G1176_i2, G1189_i2, G3066_i2, G3137_i2, G3038_i2,
    G3117_i2, G2384_i2, G2472_i2, G772_i2, G935_i2, G2923_i2, G2971_i2,
    G2980_i2, G3039_i2, G2388_i2, G2287_i2, G3024_i2, G2916_i2, G1819_i2,
    G3035_i2, G3107_i2, G1023_i2, G1024_i2, G1311_i2, G1312_i2, G3063_i2,
    G1520_i2, G1519_i2, G3078_i2, G2038_i2, G1848_i2, G1864_i2, G1872_i2,
    G1880_i2, G1888_i2, G1912_i2, G1928_i2, G1936_i2, G1944_i2, G1952_i2,
    G1850_i2, G1866_i2, G1874_i2, G1882_i2, G1890_i2, G1914_i2, G1930_i2,
    G1938_i2, G1946_i2, G1954_i2, G1845_i2, G1861_i2, G1869_i2, G1877_i2,
    G1885_i2, G1909_i2, G1925_i2, G1933_i2, G1941_i2, G1949_i2, G1846_i2,
    G1862_i2, G1870_i2, G1878_i2, G1886_i2, G1910_i2, G1926_i2, G1934_i2,
    G1942_i2, G1950_i2, G1849_i2, G1865_i2, G1873_i2, G1881_i2, G1889_i2,
    G1913_i2, G1929_i2, G1937_i2, G1945_i2, G1953_i2, G1843_i2, G1859_i2,
    G1867_i2, G1875_i2, G1883_i2, G1907_i2, G1923_i2, G1931_i2, G1939_i2,
    G1947_i2, G1844_i2, G1860_i2, G1868_i2, G1876_i2, G1884_i2, G1908_i2,
    G1924_i2, G1932_i2, G1940_i2, G1948_i2, G1847_i2, G1863_i2, G1871_i2,
    G1879_i2, G1887_i2, G1911_i2, G1927_i2, G1935_i2, G1943_i2, G1951_i2,
    G2444_i2, G2451_i2, G2502_i2, G2507_i2, G2515_i2, G2583_i2,
    n1797_lo_buf_i2, n1833_lo_buf_i2, n1881_lo_buf_i2, G523_i2, G575_i2,
    G578_i2, G615_i2, G2254_i2, G2255_i2, G2027_i2, G2393_i2, G527_i2,
    G594_i2, G1689_i2, G1693_i2, G2281_i2, G2014_i2, G2459_i2, G2561_i2,
    G2533_i2, n1749_lo_buf_i2, n1761_lo_buf_i2, n1773_lo_buf_i2,
    n1809_lo_buf_i2, G1955_i2, G1958_i2, G2562_i2, G2398_i2, G2524_i2,
    G2563_i2, G2577_i2, G2627_i2, G654_i2, G660_i2, G831_i2, G919_i2,
    G925_i2, n1815_lo_buf_i2, n1899_lo_buf_i2, n2079_lo_buf_i2,
    n2127_lo_buf_i2, n2139_lo_buf_i2, n2151_lo_buf_i2, n2187_lo_buf_i2,
    n2199_lo_buf_i2, n2211_lo_buf_i2, G533_i2, n1854_lo_buf_i2,
    n2094_lo_buf_i2, G667_i2, G874_i2, G851_i2, G1127_i2, n1869_lo_buf_i2,
    n2109_lo_buf_i2, n2121_lo_buf_i2, G477_i2, G491_i2, G501_i2, G786_i2,
    G791_i2, G1126_i2, G1052_i2, G1054_i2;
  assign new_n1131_ = G1;
  assign new_n1133_ = G2;
  assign new_n1135_ = G3;
  assign new_n1136_ = ~G3;
  assign new_n1137_ = G4;
  assign new_n1139_ = G5;
  assign new_n1141_ = G6;
  assign new_n1143_ = G7;
  assign new_n1145_ = G8;
  assign new_n1147_ = G9;
  assign new_n1149_ = G10;
  assign new_n1151_ = G11;
  assign new_n1153_ = G12;
  assign new_n1155_ = G13;
  assign new_n1157_ = G14;
  assign new_n1159_ = G15;
  assign new_n1161_ = G16;
  assign new_n1163_ = G17;
  assign new_n1165_ = G18;
  assign new_n1167_ = G19;
  assign new_n1169_ = G20;
  assign new_n1171_ = G21;
  assign new_n1173_ = G22;
  assign new_n1175_ = G23;
  assign new_n1177_ = G24;
  assign new_n1179_ = G25;
  assign new_n1181_ = G26;
  assign new_n1183_ = G27;
  assign new_n1185_ = G28;
  assign new_n1187_ = G29;
  assign new_n1189_ = G30;
  assign new_n1191_ = G31;
  assign new_n1193_ = G32;
  assign new_n1195_ = G33;
  assign new_n1197_ = G34;
  assign new_n1199_ = G35;
  assign new_n1201_ = G36;
  assign new_n1203_ = G37;
  assign new_n1205_ = G38;
  assign new_n1207_ = G39;
  assign new_n1209_ = G40;
  assign new_n1211_ = G41;
  assign new_n1213_ = G42;
  assign new_n1215_ = G43;
  assign new_n1217_ = G44;
  assign new_n1219_ = G45;
  assign new_n1221_ = G46;
  assign new_n1223_ = G47;
  assign new_n1225_ = G48;
  assign new_n1227_ = G49;
  assign new_n1229_ = G50;
  assign new_n1231_ = n1836_lo;
  assign new_n1232_ = ~n1836_lo;
  assign new_n1234_ = ~n1872_lo;
  assign new_n1235_ = n1884_lo;
  assign new_n1236_ = ~n1884_lo;
  assign new_n1237_ = n1911_lo;
  assign new_n1239_ = n1914_lo;
  assign new_n1242_ = ~n1917_lo;
  assign new_n1243_ = n1923_lo;
  assign new_n1245_ = n1926_lo;
  assign new_n1248_ = ~n1929_lo;
  assign new_n1249_ = n1935_lo;
  assign new_n1251_ = n1938_lo;
  assign new_n1253_ = n1947_lo;
  assign new_n1255_ = n1950_lo;
  assign new_n1257_ = n1959_lo;
  assign new_n1259_ = n1962_lo;
  assign new_n1261_ = n1971_lo;
  assign new_n1263_ = n1974_lo;
  assign new_n1265_ = n1983_lo;
  assign new_n1267_ = n1995_lo;
  assign new_n1268_ = ~n1995_lo;
  assign new_n1269_ = n2007_lo;
  assign new_n1270_ = ~n2007_lo;
  assign new_n1271_ = n2019_lo;
  assign new_n1272_ = ~n2019_lo;
  assign new_n1273_ = n2031_lo;
  assign new_n1274_ = ~n2031_lo;
  assign new_n1275_ = n2043_lo;
  assign new_n1276_ = ~n2043_lo;
  assign new_n1277_ = n2055_lo;
  assign new_n1278_ = ~n2055_lo;
  assign new_n1279_ = n2064_lo;
  assign new_n1281_ = n2067_lo;
  assign new_n1284_ = ~n2100_lo;
  assign new_n1286_ = ~n2112_lo;
  assign new_n1288_ = ~n2124_lo;
  assign new_n1290_ = ~n2136_lo;
  assign new_n1292_ = ~n2148_lo;
  assign new_n1294_ = ~n2160_lo;
  assign new_n1295_ = n2163_lo;
  assign new_n1296_ = ~n2163_lo;
  assign new_n1298_ = ~n2172_lo;
  assign new_n1299_ = n2175_lo;
  assign new_n1302_ = ~n2184_lo;
  assign new_n1303_ = n2223_lo;
  assign new_n1305_ = n2235_lo;
  assign new_n1307_ = n2238_lo;
  assign new_n1309_ = n2247_lo;
  assign new_n1311_ = n2250_lo;
  assign new_n1313_ = n2259_lo;
  assign new_n1315_ = n2262_lo;
  assign new_n1317_ = n2271_lo;
  assign new_n1319_ = n2274_lo;
  assign new_n1321_ = n2283_lo;
  assign new_n1323_ = n2286_lo;
  assign new_n1325_ = n2295_lo;
  assign new_n1327_ = n2298_lo;
  assign new_n1328_ = ~n2298_lo;
  assign new_n1329_ = n2304_lo;
  assign new_n1330_ = ~n2304_lo;
  assign new_n1331_ = n2307_lo;
  assign new_n1332_ = ~n2307_lo;
  assign new_n1333_ = n2331_lo;
  assign new_n1335_ = n2334_lo;
  assign new_n1337_ = n2337_lo;
  assign new_n1339_ = n2340_lo;
  assign new_n1340_ = ~n2340_lo;
  assign new_n1341_ = n3241_o2;
  assign new_n1342_ = ~n3241_o2;
  assign new_n1343_ = n3242_o2;
  assign new_n1344_ = ~n3242_o2;
  assign new_n1346_ = ~n3610_o2;
  assign new_n1348_ = ~n3980_o2;
  assign new_n1350_ = ~n3968_o2;
  assign new_n1351_ = n4298_o2;
  assign new_n1353_ = n4371_o2;
  assign new_n1356_ = ~n4413_o2;
  assign new_n1357_ = n4418_o2;
  assign new_n1359_ = n4628_o2;
  assign new_n1362_ = ~n4629_o2;
  assign new_n1363_ = n4633_o2;
  assign new_n1364_ = ~n4633_o2;
  assign new_n1365_ = n4634_o2;
  assign new_n1366_ = ~n4634_o2;
  assign new_n1367_ = n4732_o2;
  assign new_n1368_ = ~n4732_o2;
  assign new_n1369_ = n4733_o2;
  assign new_n1370_ = ~n4733_o2;
  assign new_n1372_ = ~n4884_o2;
  assign new_n1374_ = ~n4886_o2;
  assign new_n1375_ = n4890_o2;
  assign new_n1377_ = n5011_o2;
  assign new_n1378_ = ~n5011_o2;
  assign new_n1379_ = n5012_o2;
  assign new_n1380_ = ~n5012_o2;
  assign new_n1381_ = n5013_o2;
  assign new_n1382_ = ~n5013_o2;
  assign new_n1383_ = n5014_o2;
  assign new_n1385_ = n5015_o2;
  assign new_n1386_ = ~n5015_o2;
  assign new_n1387_ = n5021_o2;
  assign new_n1389_ = n5016_o2;
  assign new_n1392_ = ~n5026_o2;
  assign new_n1393_ = n4377_o2;
  assign new_n1395_ = n4378_o2;
  assign new_n1397_ = n4389_o2;
  assign new_n1398_ = ~n4389_o2;
  assign new_n1399_ = n327_inv;
  assign new_n1401_ = n330_inv;
  assign new_n1403_ = n4398_o2;
  assign new_n1404_ = ~n4398_o2;
  assign new_n1405_ = n4401_o2;
  assign new_n1406_ = ~n4401_o2;
  assign new_n1407_ = n5117_o2;
  assign new_n1409_ = n5115_o2;
  assign new_n1411_ = n5122_o2;
  assign new_n1413_ = n5121_o2;
  assign new_n1415_ = n5119_o2;
  assign new_n1417_ = n5116_o2;
  assign new_n1419_ = n5123_o2;
  assign new_n1420_ = ~n5123_o2;
  assign new_n1421_ = n5156_o2;
  assign new_n1422_ = ~n5156_o2;
  assign new_n1423_ = n5167_o2;
  assign new_n1424_ = ~n5167_o2;
  assign new_n1425_ = n4454_o2;
  assign new_n1427_ = n4455_o2;
  assign new_n1429_ = n4456_o2;
  assign new_n1431_ = n4505_o2;
  assign new_n1433_ = G742_o2;
  assign new_n1434_ = ~G742_o2;
  assign new_n1436_ = ~G727_o2;
  assign new_n1437_ = n4567_o2;
  assign new_n1439_ = n4568_o2;
  assign new_n1441_ = n4569_o2;
  assign new_n1443_ = n4571_o2;
  assign new_n1444_ = ~n4571_o2;
  assign new_n1445_ = n4572_o2;
  assign new_n1446_ = ~n4572_o2;
  assign new_n1447_ = n399_inv;
  assign new_n1449_ = n4539_o2;
  assign new_n1450_ = ~n4539_o2;
  assign new_n1451_ = n4651_o2;
  assign new_n1452_ = ~n4651_o2;
  assign new_n1453_ = n4652_o2;
  assign new_n1455_ = n4653_o2;
  assign new_n1456_ = ~n4653_o2;
  assign new_n1457_ = G1514_o2;
  assign new_n1458_ = ~G1514_o2;
  assign new_n1459_ = G1823_o2;
  assign new_n1460_ = ~G1823_o2;
  assign new_n1461_ = n4783_o2;
  assign new_n1462_ = ~n4783_o2;
  assign new_n1463_ = n4787_o2;
  assign new_n1465_ = n426_inv;
  assign new_n1467_ = n429_inv;
  assign new_n1468_ = ~n429_inv;
  assign new_n1469_ = n4816_o2;
  assign new_n1470_ = ~n4816_o2;
  assign new_n1471_ = n435_inv;
  assign new_n1473_ = G572_o2;
  assign new_n1474_ = ~G572_o2;
  assign new_n1475_ = n4919_o2;
  assign new_n1476_ = ~n4919_o2;
  assign new_n1477_ = n4920_o2;
  assign new_n1479_ = n4921_o2;
  assign new_n1481_ = G1048_o2;
  assign new_n1482_ = ~G1048_o2;
  assign new_n1483_ = n5041_o2;
  assign new_n1484_ = ~n5041_o2;
  assign new_n1485_ = n5094_o2;
  assign new_n1486_ = ~n5094_o2;
  assign new_n1487_ = n5278_o2;
  assign new_n1488_ = ~n5278_o2;
  assign new_n1489_ = n5301_o2;
  assign new_n1490_ = ~n5301_o2;
  assign new_n1491_ = G2610_o2;
  assign new_n1493_ = G3174_o2;
  assign new_n1495_ = G3146_o2;
  assign new_n1497_ = G3217_o2;
  assign new_n1499_ = G3220_o2;
  assign new_n1501_ = G2839_o2;
  assign new_n1503_ = G3251_o2;
  assign new_n1505_ = G3042_o2;
  assign new_n1508_ = ~G3045_o2;
  assign new_n1509_ = G3262_o2;
  assign new_n1511_ = G2845_o2;
  assign new_n1513_ = G2929_o2;
  assign new_n1515_ = G2848_o2;
  assign new_n1517_ = G2851_o2;
  assign new_n1519_ = G3291_o2;
  assign new_n1521_ = G3254_o2;
  assign new_n1523_ = G2666_o2;
  assign new_n1524_ = ~G2666_o2;
  assign new_n1525_ = n5099_o2;
  assign new_n1527_ = n5100_o2;
  assign new_n1528_ = ~n5100_o2;
  assign new_n1529_ = n5101_o2;
  assign new_n1530_ = ~n5101_o2;
  assign new_n1531_ = G2558_o2;
  assign new_n1533_ = n5266_o2;
  assign new_n1534_ = ~n5266_o2;
  assign new_n1535_ = n5267_o2;
  assign new_n1536_ = ~n5267_o2;
  assign new_n1537_ = G2759_o2;
  assign new_n1538_ = ~G2759_o2;
  assign new_n1539_ = n537_inv;
  assign new_n1541_ = n540_inv;
  assign new_n1543_ = n543_inv;
  assign new_n1545_ = n5292_o2;
  assign new_n1547_ = n5293_o2;
  assign new_n1549_ = n5294_o2;
  assign new_n1550_ = ~n5294_o2;
  assign new_n1551_ = n5295_o2;
  assign new_n1553_ = G618_o2;
  assign new_n1554_ = ~G618_o2;
  assign new_n1555_ = G621_o2;
  assign new_n1556_ = ~G621_o2;
  assign new_n1558_ = ~G384_o2;
  assign new_n1560_ = ~G377_o2;
  assign new_n1561_ = n570_inv;
  assign new_n1562_ = ~n570_inv;
  assign new_n1563_ = G3171_o2;
  assign new_n1565_ = G2552_o2;
  assign new_n1567_ = G3272_o2;
  assign new_n1569_ = G2015_o2;
  assign new_n1570_ = ~G2015_o2;
  assign new_n1571_ = G3294_o2;
  assign new_n1573_ = G3281_o2;
  assign new_n1575_ = G3320_o2;
  assign new_n1577_ = G3275_o2;
  assign new_n1579_ = G3140_o2;
  assign new_n1581_ = G2836_o2;
  assign new_n1583_ = G2926_o2;
  assign new_n1585_ = G2842_o2;
  assign new_n1587_ = G3302_o2;
  assign new_n1589_ = G3288_o2;
  assign new_n1591_ = G3143_o2;
  assign new_n1594_ = ~G3100_o2;
  assign new_n1595_ = G2512_o2;
  assign new_n1596_ = ~G2512_o2;
  assign new_n1597_ = n5325_o2;
  assign new_n1598_ = ~n5325_o2;
  assign new_n1599_ = n5326_o2;
  assign new_n1600_ = ~n5326_o2;
  assign new_n1601_ = n5327_o2;
  assign new_n1602_ = ~n5327_o2;
  assign new_n1603_ = n1857_lo_buf_o2;
  assign new_n1604_ = ~n1857_lo_buf_o2;
  assign new_n1605_ = n2097_lo_buf_o2;
  assign new_n1606_ = ~n2097_lo_buf_o2;
  assign new_n1607_ = G2669_o2;
  assign new_n1608_ = ~G2669_o2;
  assign new_n1609_ = n642_inv;
  assign new_n1611_ = G568_o2;
  assign new_n1613_ = n648_inv;
  assign new_n1615_ = G565_o2;
  assign new_n1617_ = G559_o2;
  assign new_n1619_ = n1821_lo_buf_o2;
  assign new_n1620_ = ~n1821_lo_buf_o2;
  assign new_n1621_ = n1905_lo_buf_o2;
  assign new_n1622_ = ~n1905_lo_buf_o2;
  assign new_n1623_ = n2133_lo_buf_o2;
  assign new_n1624_ = ~n2133_lo_buf_o2;
  assign new_n1625_ = n2145_lo_buf_o2;
  assign new_n1626_ = ~n2145_lo_buf_o2;
  assign new_n1627_ = n2157_lo_buf_o2;
  assign new_n1628_ = ~n2157_lo_buf_o2;
  assign new_n1629_ = n2205_lo_buf_o2;
  assign new_n1631_ = n2217_lo_buf_o2;
  assign new_n1633_ = G447_o2;
  assign new_n1634_ = ~G447_o2;
  assign new_n1635_ = G434_o2;
  assign new_n1638_ = ~G422_o2;
  assign new_n1639_ = G461_o2;
  assign new_n1641_ = G3312_o2;
  assign new_n1643_ = G3332_o2;
  assign new_n1645_ = G3195_o2;
  assign new_n1647_ = G2607_o2;
  assign new_n1649_ = n702_inv;
  assign new_n1651_ = G1005_o2;
  assign new_n1653_ = G1008_o2;
  assign new_n1655_ = n2001_lo_buf_o2;
  assign new_n1657_ = n2169_lo_buf_o2;
  assign new_n1658_ = ~n2169_lo_buf_o2;
  assign new_n1659_ = n2229_lo_buf_o2;
  assign new_n1661_ = n2301_lo_buf_o2;
  assign new_n1662_ = ~n2301_lo_buf_o2;
  assign new_n1663_ = n723_inv;
  assign new_n1665_ = G2947_o2;
  assign new_n1667_ = n2013_lo_buf_o2;
  assign new_n1668_ = ~n2013_lo_buf_o2;
  assign new_n1669_ = n2025_lo_buf_o2;
  assign new_n1670_ = ~n2025_lo_buf_o2;
  assign new_n1671_ = n2037_lo_buf_o2;
  assign new_n1672_ = ~n2037_lo_buf_o2;
  assign new_n1673_ = n2049_lo_buf_o2;
  assign new_n1674_ = ~n2049_lo_buf_o2;
  assign new_n1675_ = n2181_lo_buf_o2;
  assign new_n1676_ = ~n2181_lo_buf_o2;
  assign new_n1677_ = n744_inv;
  assign new_n1679_ = n747_inv;
  assign new_n1681_ = n750_inv;
  assign new_n1683_ = n753_inv;
  assign new_n1685_ = G3350_o2;
  assign new_n1686_ = ~G3350_o2;
  assign new_n1687_ = G3360_o2;
  assign new_n1688_ = ~G3360_o2;
  assign new_n1689_ = G3373_o2;
  assign new_n1690_ = ~G3373_o2;
  assign new_n1691_ = G3237_o2;
  assign new_n1692_ = ~G3237_o2;
  assign new_n1693_ = G2773_o2;
  assign new_n1694_ = ~G2773_o2;
  assign new_n1695_ = G1733_o2;
  assign new_n1696_ = ~G1733_o2;
  assign new_n1697_ = G1738_o2;
  assign new_n1698_ = ~G1738_o2;
  assign new_n1699_ = G1751_o2;
  assign new_n1700_ = ~G1751_o2;
  assign new_n1701_ = G2216_o2;
  assign new_n1702_ = ~G2216_o2;
  assign new_n1703_ = G2219_o2;
  assign new_n1704_ = ~G2219_o2;
  assign new_n1705_ = n786_inv;
  assign new_n1707_ = n789_inv;
  assign new_n1709_ = G787_o2;
  assign new_n1711_ = G2823_o2;
  assign new_n1713_ = G2796_o2;
  assign new_n1715_ = G875_o2;
  assign new_n1716_ = ~G875_o2;
  assign new_n1717_ = G2208_o2;
  assign new_n1718_ = ~G2208_o2;
  assign new_n1719_ = G2211_o2;
  assign new_n1720_ = ~G2211_o2;
  assign new_n1721_ = n1989_lo_buf_o2;
  assign new_n1723_ = n2061_lo_buf_o2;
  assign new_n1724_ = ~n2061_lo_buf_o2;
  assign new_n1725_ = n2313_lo_buf_o2;
  assign new_n1726_ = ~n2313_lo_buf_o2;
  assign new_n1727_ = G2232_o2;
  assign new_n1728_ = ~G2232_o2;
  assign new_n1729_ = G1725_o2;
  assign new_n1730_ = ~G1725_o2;
  assign new_n1731_ = G1764_o2;
  assign new_n1732_ = ~G1764_o2;
  assign new_n1733_ = G2356_o2;
  assign new_n1734_ = ~G2356_o2;
  assign new_n1735_ = G2359_o2;
  assign new_n1736_ = ~G2359_o2;
  assign new_n1737_ = G1180_o2;
  assign new_n1738_ = ~G1180_o2;
  assign new_n1739_ = G1756_o2;
  assign new_n1740_ = ~G1756_o2;
  assign new_n1742_ = ~G2441_o2;
  assign new_n1743_ = G2887_o2;
  assign new_n1744_ = ~G2887_o2;
  assign new_n1745_ = G2991_o2;
  assign new_n1746_ = ~G2991_o2;
  assign new_n1747_ = n849_inv;
  assign new_n1748_ = ~n849_inv;
  assign new_n1749_ = n852_inv;
  assign new_n1750_ = ~n852_inv;
  assign new_n1751_ = n855_inv;
  assign new_n1752_ = ~n855_inv;
  assign new_n1753_ = n858_inv;
  assign new_n1754_ = ~n858_inv;
  assign new_n1755_ = n861_inv;
  assign new_n1756_ = ~n861_inv;
  assign new_n1757_ = G2805_o2;
  assign new_n1759_ = G2906_o2;
  assign new_n1761_ = G2833_o2;
  assign new_n1763_ = n873_inv;
  assign new_n1765_ = G3353_o2;
  assign new_n1766_ = ~G3353_o2;
  assign new_n1767_ = G3367_o2;
  assign new_n1768_ = ~G3367_o2;
  assign new_n1769_ = G3346_o2;
  assign new_n1770_ = ~G3346_o2;
  assign new_n1771_ = G3340_o2;
  assign new_n1772_ = ~G3340_o2;
  assign new_n1773_ = G3376_o2;
  assign new_n1774_ = ~G3376_o2;
  assign new_n1775_ = G3359_o2;
  assign new_n1776_ = ~G3359_o2;
  assign new_n1777_ = G3240_o2;
  assign new_n1778_ = ~G3240_o2;
  assign new_n1779_ = G3344_o2;
  assign new_n1780_ = ~G3344_o2;
  assign new_n1781_ = G2880_o2;
  assign new_n1782_ = ~G2880_o2;
  assign new_n1783_ = G2939_o2;
  assign new_n1784_ = ~G2939_o2;
  assign new_n1785_ = G2248_o2;
  assign new_n1786_ = ~G2248_o2;
  assign new_n1787_ = G2251_o2;
  assign new_n1788_ = ~G2251_o2;
  assign new_n1789_ = G2021_o2;
  assign new_n1791_ = G3383_o2;
  assign new_n1792_ = ~G3383_o2;
  assign new_n1793_ = G3399_o2;
  assign new_n1794_ = ~G3399_o2;
  assign new_n1795_ = G3404_o2;
  assign new_n1796_ = ~G3404_o2;
  assign new_n1797_ = G3265_o2;
  assign new_n1798_ = ~G3265_o2;
  assign new_n1799_ = G2866_o2;
  assign new_n1800_ = ~G2866_o2;
  assign new_n1801_ = G2999_o2;
  assign new_n1802_ = ~G2999_o2;
  assign new_n1804_ = ~G736_o2;
  assign new_n1805_ = G739_o2;
  assign new_n1807_ = G1200_o2;
  assign new_n1809_ = G1203_o2;
  assign new_n1811_ = G3027_o2;
  assign new_n1812_ = ~G3027_o2;
  assign new_n1814_ = ~G1463_o2;
  assign new_n1816_ = ~G1460_o2;
  assign new_n1817_ = G3012_o2;
  assign new_n1818_ = ~G3012_o2;
  assign new_n1819_ = G1574_o2;
  assign new_n1821_ = G1646_o2;
  assign new_n1823_ = G1592_o2;
  assign new_n1825_ = G1664_o2;
  assign new_n1828_ = ~G1547_o2;
  assign new_n1830_ = ~G1619_o2;
  assign new_n1831_ = G1556_o2;
  assign new_n1833_ = G1628_o2;
  assign new_n1836_ = ~G1583_o2;
  assign new_n1838_ = ~G1655_o2;
  assign new_n1839_ = G1529_o2;
  assign new_n1841_ = G1601_o2;
  assign new_n1843_ = G1538_o2;
  assign new_n1845_ = G1610_o2;
  assign new_n1847_ = G1565_o2;
  assign new_n1849_ = G1637_o2;
  assign new_n1851_ = G2437_o2;
  assign new_n1852_ = ~G2437_o2;
  assign new_n1853_ = n1008_inv;
  assign new_n1855_ = n1785_lo_buf_o2;
  assign new_n1856_ = ~n1785_lo_buf_o2;
  assign new_n1857_ = n1845_lo_buf_o2;
  assign new_n1858_ = ~n1845_lo_buf_o2;
  assign new_n1859_ = n1893_lo_buf_o2;
  assign new_n1860_ = ~n1893_lo_buf_o2;
  assign new_n1862_ = ~n1941_lo_buf_o2;
  assign new_n1864_ = ~n1953_lo_buf_o2;
  assign new_n1866_ = ~n1965_lo_buf_o2;
  assign new_n1867_ = n1977_lo_buf_o2;
  assign new_n1868_ = ~n1977_lo_buf_o2;
  assign new_n1869_ = n2241_lo_buf_o2;
  assign new_n1870_ = ~n2241_lo_buf_o2;
  assign new_n1871_ = n2253_lo_buf_o2;
  assign new_n1872_ = ~n2253_lo_buf_o2;
  assign new_n1873_ = n2265_lo_buf_o2;
  assign new_n1874_ = ~n2265_lo_buf_o2;
  assign new_n1875_ = n2277_lo_buf_o2;
  assign new_n1876_ = ~n2277_lo_buf_o2;
  assign new_n1877_ = n2289_lo_buf_o2;
  assign new_n1879_ = G519_o2;
  assign new_n1880_ = ~G519_o2;
  assign new_n1881_ = n1050_inv;
  assign new_n1882_ = ~n1050_inv;
  assign new_n1883_ = n1053_inv;
  assign new_n1884_ = ~n1053_inv;
  assign new_n1885_ = n1056_inv;
  assign new_n1886_ = ~n1056_inv;
  assign new_n1888_ = ~G1318_o2;
  assign new_n1889_ = n1062_inv;
  assign new_n1890_ = ~n1062_inv;
  assign new_n1891_ = G593_o2;
  assign new_n1892_ = ~G593_o2;
  assign new_n1893_ = n1068_inv;
  assign new_n1894_ = ~n1068_inv;
  assign new_n1895_ = n1071_inv;
  assign new_n1896_ = ~n1071_inv;
  assign new_n1897_ = n1074_inv;
  assign new_n1898_ = ~n1074_inv;
  assign new_n1899_ = G2284_o2;
  assign new_n1900_ = ~G2284_o2;
  assign new_n1901_ = G2580_o2;
  assign new_n1902_ = ~G2580_o2;
  assign new_n1903_ = G2302_o2;
  assign new_n1904_ = ~G2302_o2;
  assign new_n1905_ = G2598_o2;
  assign new_n1906_ = ~G2598_o2;
  assign new_n1907_ = G2497_o2;
  assign new_n1908_ = ~G2497_o2;
  assign new_n1909_ = G2651_o2;
  assign new_n1910_ = ~G2651_o2;
  assign new_n1911_ = G2296_o2;
  assign new_n1912_ = ~G2296_o2;
  assign new_n1913_ = G2308_o2;
  assign new_n1914_ = ~G2308_o2;
  assign new_n1915_ = G2592_o2;
  assign new_n1916_ = ~G2592_o2;
  assign new_n1917_ = G2604_o2;
  assign new_n1918_ = ~G2604_o2;
  assign new_n1919_ = G2902_o2;
  assign new_n1920_ = ~G2902_o2;
  assign new_n1921_ = G2975_o2;
  assign new_n1922_ = ~G2975_o2;
  assign new_n1923_ = G2962_o2;
  assign new_n1924_ = ~G2962_o2;
  assign new_n1925_ = G3069_o2;
  assign new_n1926_ = ~G3069_o2;
  assign new_n1927_ = G2018_o2;
  assign new_n1929_ = G1176_o2;
  assign new_n1930_ = ~G1176_o2;
  assign new_n1931_ = G1189_o2;
  assign new_n1932_ = ~G1189_o2;
  assign new_n1933_ = G3066_o2;
  assign new_n1934_ = ~G3066_o2;
  assign new_n1935_ = G3137_o2;
  assign new_n1936_ = ~G3137_o2;
  assign new_n1937_ = G3038_o2;
  assign new_n1938_ = ~G3038_o2;
  assign new_n1939_ = G3117_o2;
  assign new_n1940_ = ~G3117_o2;
  assign new_n1941_ = G2384_o2;
  assign new_n1942_ = ~G2384_o2;
  assign new_n1943_ = G2472_o2;
  assign new_n1944_ = ~G2472_o2;
  assign new_n1945_ = G772_o2;
  assign new_n1946_ = ~G772_o2;
  assign new_n1947_ = G935_o2;
  assign new_n1949_ = G2923_o2;
  assign new_n1950_ = ~G2923_o2;
  assign new_n1951_ = G2971_o2;
  assign new_n1952_ = ~G2971_o2;
  assign new_n1953_ = G2980_o2;
  assign new_n1954_ = ~G2980_o2;
  assign new_n1955_ = G3039_o2;
  assign new_n1956_ = ~G3039_o2;
  assign new_n1957_ = G2388_o2;
  assign new_n1958_ = ~G2388_o2;
  assign new_n1959_ = G2287_o2;
  assign new_n1960_ = ~G2287_o2;
  assign new_n1961_ = G3024_o2;
  assign new_n1962_ = ~G3024_o2;
  assign new_n1963_ = G2916_o2;
  assign new_n1964_ = ~G2916_o2;
  assign new_n1965_ = n1176_inv;
  assign new_n1966_ = ~n1176_inv;
  assign new_n1967_ = G3035_o2;
  assign new_n1968_ = ~G3035_o2;
  assign new_n1969_ = G3107_o2;
  assign new_n1970_ = ~G3107_o2;
  assign new_n1971_ = G1023_o2;
  assign new_n1974_ = ~G1024_o2;
  assign new_n1976_ = ~G1311_o2;
  assign new_n1978_ = ~G1312_o2;
  assign new_n1979_ = G3063_o2;
  assign new_n1980_ = ~G3063_o2;
  assign new_n1981_ = G1520_o2;
  assign new_n1983_ = G1519_o2;
  assign new_n1985_ = G3078_o2;
  assign new_n1986_ = ~G3078_o2;
  assign new_n1987_ = G2038_o2;
  assign new_n1989_ = G1848_o2;
  assign new_n1991_ = G1864_o2;
  assign new_n1994_ = ~G1872_o2;
  assign new_n1995_ = G1880_o2;
  assign new_n1998_ = ~G1888_o2;
  assign new_n1999_ = G1912_o2;
  assign new_n2001_ = G1928_o2;
  assign new_n2004_ = ~G1936_o2;
  assign new_n2005_ = G1944_o2;
  assign new_n2008_ = ~G1952_o2;
  assign new_n2009_ = G1850_o2;
  assign new_n2011_ = G1866_o2;
  assign new_n2014_ = ~G1874_o2;
  assign new_n2015_ = G1882_o2;
  assign new_n2018_ = ~G1890_o2;
  assign new_n2019_ = G1914_o2;
  assign new_n2021_ = G1930_o2;
  assign new_n2024_ = ~G1938_o2;
  assign new_n2025_ = G1946_o2;
  assign new_n2028_ = ~G1954_o2;
  assign new_n2030_ = ~G1845_o2;
  assign new_n2032_ = ~G1861_o2;
  assign new_n2033_ = G1869_o2;
  assign new_n2036_ = ~G1877_o2;
  assign new_n2037_ = G1885_o2;
  assign new_n2040_ = ~G1909_o2;
  assign new_n2042_ = ~G1925_o2;
  assign new_n2043_ = G1933_o2;
  assign new_n2046_ = ~G1941_o2;
  assign new_n2047_ = G1949_o2;
  assign new_n2049_ = G1846_o2;
  assign new_n2051_ = G1862_o2;
  assign new_n2054_ = ~G1870_o2;
  assign new_n2055_ = G1878_o2;
  assign new_n2058_ = ~G1886_o2;
  assign new_n2059_ = G1910_o2;
  assign new_n2061_ = G1926_o2;
  assign new_n2064_ = ~G1934_o2;
  assign new_n2065_ = G1942_o2;
  assign new_n2068_ = ~G1950_o2;
  assign new_n2070_ = ~G1849_o2;
  assign new_n2072_ = ~G1865_o2;
  assign new_n2073_ = G1873_o2;
  assign new_n2076_ = ~G1881_o2;
  assign new_n2077_ = G1889_o2;
  assign new_n2080_ = ~G1913_o2;
  assign new_n2082_ = ~G1929_o2;
  assign new_n2083_ = G1937_o2;
  assign new_n2086_ = ~G1945_o2;
  assign new_n2087_ = G1953_o2;
  assign new_n2089_ = G1843_o2;
  assign new_n2091_ = G1859_o2;
  assign new_n2094_ = ~G1867_o2;
  assign new_n2095_ = G1875_o2;
  assign new_n2098_ = ~G1883_o2;
  assign new_n2099_ = G1907_o2;
  assign new_n2101_ = G1923_o2;
  assign new_n2104_ = ~G1931_o2;
  assign new_n2105_ = G1939_o2;
  assign new_n2108_ = ~G1947_o2;
  assign new_n2109_ = G1844_o2;
  assign new_n2111_ = G1860_o2;
  assign new_n2114_ = ~G1868_o2;
  assign new_n2115_ = G1876_o2;
  assign new_n2118_ = ~G1884_o2;
  assign new_n2119_ = G1908_o2;
  assign new_n2121_ = G1924_o2;
  assign new_n2124_ = ~G1932_o2;
  assign new_n2125_ = G1940_o2;
  assign new_n2128_ = ~G1948_o2;
  assign new_n2129_ = G1847_o2;
  assign new_n2131_ = G1863_o2;
  assign new_n2134_ = ~G1871_o2;
  assign new_n2135_ = G1879_o2;
  assign new_n2138_ = ~G1887_o2;
  assign new_n2139_ = G1911_o2;
  assign new_n2141_ = G1927_o2;
  assign new_n2144_ = ~G1935_o2;
  assign new_n2145_ = G1943_o2;
  assign new_n2148_ = ~G1951_o2;
  assign new_n2149_ = G2444_o2;
  assign new_n2150_ = ~G2444_o2;
  assign new_n2151_ = G2451_o2;
  assign new_n2152_ = ~G2451_o2;
  assign new_n2153_ = G2502_o2;
  assign new_n2154_ = ~G2502_o2;
  assign new_n2155_ = G2507_o2;
  assign new_n2156_ = ~G2507_o2;
  assign new_n2157_ = n1464_inv;
  assign new_n2159_ = G2583_o2;
  assign new_n2160_ = ~G2583_o2;
  assign new_n2161_ = n1797_lo_buf_o2;
  assign new_n2162_ = ~n1797_lo_buf_o2;
  assign new_n2163_ = n1833_lo_buf_o2;
  assign new_n2164_ = ~n1833_lo_buf_o2;
  assign new_n2165_ = n1881_lo_buf_o2;
  assign new_n2166_ = ~n1881_lo_buf_o2;
  assign new_n2167_ = n1479_inv;
  assign new_n2169_ = n1482_inv;
  assign new_n2171_ = n1485_inv;
  assign new_n2173_ = G615_o2;
  assign new_n2174_ = ~G615_o2;
  assign new_n2175_ = G2254_o2;
  assign new_n2176_ = ~G2254_o2;
  assign new_n2177_ = G2255_o2;
  assign new_n2178_ = ~G2255_o2;
  assign new_n2179_ = G2027_o2;
  assign new_n2180_ = ~G2027_o2;
  assign new_n2181_ = G2393_o2;
  assign new_n2182_ = ~G2393_o2;
  assign new_n2183_ = G527_o2;
  assign new_n2184_ = ~G527_o2;
  assign new_n2185_ = G594_o2;
  assign new_n2186_ = ~G594_o2;
  assign new_n2187_ = G1689_o2;
  assign new_n2188_ = ~G1689_o2;
  assign new_n2189_ = G1693_o2;
  assign new_n2190_ = ~G1693_o2;
  assign new_n2191_ = G2281_o2;
  assign new_n2192_ = ~G2281_o2;
  assign new_n2193_ = G2014_o2;
  assign new_n2194_ = ~G2014_o2;
  assign new_n2195_ = G2459_o2;
  assign new_n2196_ = ~G2459_o2;
  assign new_n2197_ = G2561_o2;
  assign new_n2198_ = ~G2561_o2;
  assign new_n2199_ = G2533_o2;
  assign new_n2200_ = ~G2533_o2;
  assign new_n2201_ = n1749_lo_buf_o2;
  assign new_n2202_ = ~n1749_lo_buf_o2;
  assign new_n2203_ = n1761_lo_buf_o2;
  assign new_n2204_ = ~n1761_lo_buf_o2;
  assign new_n2205_ = n1773_lo_buf_o2;
  assign new_n2206_ = ~n1773_lo_buf_o2;
  assign new_n2207_ = n1809_lo_buf_o2;
  assign new_n2208_ = ~n1809_lo_buf_o2;
  assign new_n2209_ = G1955_o2;
  assign new_n2210_ = ~G1955_o2;
  assign new_n2211_ = G1958_o2;
  assign new_n2212_ = ~G1958_o2;
  assign new_n2213_ = G2562_o2;
  assign new_n2214_ = ~G2562_o2;
  assign new_n2215_ = G2398_o2;
  assign new_n2216_ = ~G2398_o2;
  assign new_n2217_ = n1554_inv;
  assign new_n2218_ = ~n1554_inv;
  assign new_n2219_ = n1557_inv;
  assign new_n2220_ = ~n1557_inv;
  assign new_n2221_ = G2577_o2;
  assign new_n2222_ = ~G2577_o2;
  assign new_n2223_ = G2627_o2;
  assign new_n2224_ = ~G2627_o2;
  assign new_n2225_ = G654_o2;
  assign new_n2226_ = ~G654_o2;
  assign new_n2227_ = G660_o2;
  assign new_n2228_ = ~G660_o2;
  assign new_n2229_ = G831_o2;
  assign new_n2230_ = ~G831_o2;
  assign new_n2231_ = G919_o2;
  assign new_n2232_ = ~G919_o2;
  assign new_n2233_ = G925_o2;
  assign new_n2234_ = ~G925_o2;
  assign new_n2235_ = n1815_lo_buf_o2;
  assign new_n2236_ = ~n1815_lo_buf_o2;
  assign new_n2237_ = n1899_lo_buf_o2;
  assign new_n2238_ = ~n1899_lo_buf_o2;
  assign new_n2239_ = n2079_lo_buf_o2;
  assign new_n2240_ = ~n2079_lo_buf_o2;
  assign new_n2241_ = n2127_lo_buf_o2;
  assign new_n2242_ = ~n2127_lo_buf_o2;
  assign new_n2243_ = n2139_lo_buf_o2;
  assign new_n2244_ = ~n2139_lo_buf_o2;
  assign new_n2245_ = n2151_lo_buf_o2;
  assign new_n2246_ = ~n2151_lo_buf_o2;
  assign new_n2247_ = n2187_lo_buf_o2;
  assign new_n2248_ = ~n2187_lo_buf_o2;
  assign new_n2249_ = n2199_lo_buf_o2;
  assign new_n2250_ = ~n2199_lo_buf_o2;
  assign new_n2251_ = n2211_lo_buf_o2;
  assign new_n2252_ = ~n2211_lo_buf_o2;
  assign new_n2253_ = G533_o2;
  assign new_n2254_ = ~G533_o2;
  assign new_n2255_ = n1854_lo_buf_o2;
  assign new_n2256_ = ~n1854_lo_buf_o2;
  assign new_n2257_ = n2094_lo_buf_o2;
  assign new_n2258_ = ~n2094_lo_buf_o2;
  assign new_n2259_ = G667_o2;
  assign new_n2260_ = ~G667_o2;
  assign new_n2261_ = G874_o2;
  assign new_n2262_ = ~G874_o2;
  assign new_n2263_ = G851_o2;
  assign new_n2264_ = ~G851_o2;
  assign new_n2265_ = G1127_o2;
  assign new_n2266_ = ~G1127_o2;
  assign new_n2267_ = n1869_lo_buf_o2;
  assign new_n2268_ = ~n1869_lo_buf_o2;
  assign new_n2269_ = n2109_lo_buf_o2;
  assign new_n2270_ = ~n2109_lo_buf_o2;
  assign new_n2271_ = n2121_lo_buf_o2;
  assign new_n2272_ = ~n2121_lo_buf_o2;
  assign new_n2273_ = G477_o2;
  assign new_n2274_ = ~G477_o2;
  assign new_n2275_ = G491_o2;
  assign new_n2276_ = ~G491_o2;
  assign new_n2277_ = G501_o2;
  assign new_n2278_ = ~G501_o2;
  assign new_n2279_ = G786_o2;
  assign new_n2280_ = ~G786_o2;
  assign new_n2281_ = G791_o2;
  assign new_n2282_ = ~G791_o2;
  assign new_n2283_ = G1126_o2;
  assign new_n2284_ = ~G1126_o2;
  assign new_n2285_ = G1052_o2;
  assign new_n2286_ = ~G1052_o2;
  assign new_n2287_ = G1054_o2;
  assign new_n2288_ = ~G1054_o2;
  assign new_n2289_ = new_n1350_ & new_n1348_;
  assign new_n2290_ = new_n2289_ & new_n1346_;
  assign new_n2291_ = new_n2290_ & new_n1356_;
  assign new_n2292_ = new_n1436_ | new_n1234_;
  assign new_n2293_ = new_n1433_ & new_n4363_;
  assign new_n2294_ = new_n1434_ | new_n4364_;
  assign new_n2295_ = new_n2293_ & new_n4365_;
  assign new_n2296_ = new_n2294_ | new_n4366_;
  assign new_n2297_ = new_n4367_ | new_n1422_;
  assign new_n2298_ = new_n4368_ & new_n4369_;
  assign new_n2299_ = new_n2298_ | new_n4370_;
  assign new_n2300_ = new_n1380_ & new_n4363_;
  assign new_n2301_ = new_n1379_ | new_n4364_;
  assign new_n2302_ = new_n4371_ & new_n4365_;
  assign new_n2303_ = new_n4372_ | new_n4366_;
  assign new_n2304_ = new_n2303_ | new_n2299_;
  assign new_n2305_ = new_n1383_ | new_n1284_;
  assign new_n2306_ = new_n1407_ | new_n1286_;
  assign new_n2307_ = new_n1409_ | new_n1288_;
  assign new_n2308_ = new_n1411_ | new_n1290_;
  assign new_n2309_ = new_n2306_ & new_n2305_;
  assign new_n2310_ = new_n2309_ & new_n2307_;
  assign new_n2311_ = new_n2310_ & new_n2308_;
  assign new_n2312_ = new_n1413_ | new_n4370_;
  assign new_n2313_ = new_n1415_ | new_n4369_;
  assign new_n2314_ = new_n1417_ | new_n4368_;
  assign new_n2315_ = new_n1419_ | new_n1302_;
  assign new_n2316_ = new_n2313_ & new_n2312_;
  assign new_n2317_ = new_n2316_ & new_n2314_;
  assign new_n2318_ = new_n2317_ & new_n2315_;
  assign new_n2319_ = new_n2318_ & new_n2311_;
  assign new_n2320_ = new_n2302_ | new_n4373_;
  assign new_n2321_ = new_n2320_ | new_n2319_;
  assign new_n2322_ = new_n2304_ & new_n2297_;
  assign new_n2323_ = new_n2322_ & new_n2321_;
  assign new_n2324_ = new_n4374_ & new_n4375_;
  assign new_n2325_ = new_n4376_ | new_n4377_;
  assign new_n2326_ = new_n4376_ & new_n4377_;
  assign new_n2327_ = new_n4374_ | new_n4375_;
  assign new_n2328_ = new_n2327_ & new_n2325_;
  assign new_n2329_ = new_n2326_ | new_n2324_;
  assign new_n2330_ = new_n2328_ | new_n1458_;
  assign new_n2331_ = new_n2329_ | new_n1457_;
  assign new_n2332_ = new_n2331_ & new_n2330_;
  assign new_n2333_ = new_n1459_ & new_n1424_;
  assign new_n2334_ = new_n1460_ & new_n1423_;
  assign new_n2335_ = new_n2334_ | new_n2333_;
  assign new_n2336_ = new_n4378_ & new_n1353_;
  assign new_n2337_ = new_n4378_ & new_n1351_;
  assign new_n2338_ = new_n2337_ | new_n1359_;
  assign new_n2339_ = new_n1375_ & new_n4379_;
  assign new_n2340_ = new_n2339_ & new_n1362_;
  assign new_n2341_ = new_n1482_ & new_n1421_;
  assign new_n2342_ = new_n1389_ | new_n1387_;
  assign new_n2343_ = new_n2342_ & new_n1474_;
  assign new_n2344_ = new_n1481_ & new_n1473_;
  assign new_n2345_ = new_n2344_ & new_n1392_;
  assign new_n2346_ = new_n2343_ | new_n2341_;
  assign new_n2347_ = new_n2346_ | new_n2345_;
  assign new_n2348_ = new_n1508_ | new_n1505_;
  assign new_n2349_ = new_n2348_ | new_n1517_;
  assign new_n2350_ = new_n4380_ & new_n1594_;
  assign new_n2351_ = new_n1591_ | new_n1579_;
  assign new_n2352_ = new_n2351_ | new_n1585_;
  assign new_n2353_ = new_n4381_ & new_n1645_;
  assign new_n2354_ = new_n1341_ & new_n1231_;
  assign new_n2355_ = new_n1342_ & new_n1232_;
  assign new_n2356_ = new_n2355_ | new_n2354_;
  assign new_n2357_ = new_n2356_ & new_n1374_;
  assign new_n2358_ = new_n2357_ & new_n1386_;
  assign new_n2359_ = new_n1385_ & new_n1372_;
  assign new_n2360_ = new_n2359_ | new_n2358_;
  assign new_n2361_ = new_n2360_ & new_n4371_;
  assign new_n2362_ = new_n1343_ & new_n1235_;
  assign new_n2363_ = new_n1344_ & new_n1236_;
  assign new_n2364_ = new_n2363_ | new_n2362_;
  assign new_n2365_ = new_n2364_ & new_n1420_;
  assign new_n2366_ = new_n2365_ & new_n4373_;
  assign new_n2367_ = new_n4382_ & new_n4383_;
  assign new_n2368_ = new_n4384_ | new_n4385_;
  assign new_n2369_ = new_n4384_ & new_n4385_;
  assign new_n2370_ = new_n4382_ | new_n4383_;
  assign new_n2371_ = new_n2370_ & new_n2368_;
  assign new_n2372_ = new_n2369_ | new_n2367_;
  assign new_n2373_ = new_n2372_ & new_n4379_;
  assign new_n2374_ = new_n2371_ | new_n1330_;
  assign new_n2375_ = new_n4386_ & new_n4387_;
  assign new_n2376_ = new_n4388_ | new_n4389_;
  assign new_n2377_ = new_n4388_ & new_n4389_;
  assign new_n2378_ = new_n4386_ | new_n4387_;
  assign new_n2379_ = new_n2378_ & new_n2376_;
  assign new_n2380_ = new_n2377_ | new_n2375_;
  assign new_n2381_ = new_n2379_ & new_n2373_;
  assign new_n2382_ = new_n2380_ & new_n2374_;
  assign new_n2383_ = new_n2382_ | new_n2381_;
  assign new_n2384_ = new_n4372_ & new_n4367_;
  assign new_n2385_ = new_n2384_ & new_n2383_;
  assign new_n2386_ = new_n2366_ | new_n2361_;
  assign new_n2387_ = new_n2386_ | new_n2385_;
  assign new_n2388_ = new_n1503_ | new_n1499_;
  assign new_n2389_ = new_n2388_ | new_n1511_;
  assign new_n2390_ = new_n4390_ & new_n1577_;
  assign new_n2391_ = new_n1521_ | new_n1495_;
  assign new_n2392_ = new_n2391_ | new_n1515_;
  assign new_n2393_ = new_n4391_ & new_n1573_;
  assign new_n2394_ = new_n1509_ | new_n1493_;
  assign new_n2395_ = new_n2394_ | new_n1513_;
  assign new_n2396_ = new_n4392_ & new_n1571_;
  assign new_n2397_ = new_n1519_ | new_n1497_;
  assign new_n2398_ = new_n2397_ | new_n1501_;
  assign new_n2399_ = new_n4393_ & new_n1575_;
  assign new_n2400_ = new_n4391_ | new_n4380_;
  assign new_n2401_ = new_n2400_ | new_n4392_;
  assign new_n2402_ = new_n2401_ | new_n4390_;
  assign new_n2403_ = new_n1589_ | new_n1563_;
  assign new_n2404_ = new_n2403_ | new_n1583_;
  assign new_n2405_ = new_n1587_ | new_n1567_;
  assign new_n2406_ = new_n2405_ | new_n1581_;
  assign new_n2407_ = new_n4393_ | new_n4381_;
  assign new_n2408_ = new_n2407_ | new_n4394_;
  assign new_n2409_ = new_n2408_ | new_n4395_;
  assign new_n2410_ = new_n2409_ | new_n2402_;
  assign new_n2411_ = new_n1555_ & new_n1553_;
  assign new_n2412_ = new_n1556_ | new_n1554_;
  assign new_n2413_ = new_n4395_ | new_n4394_;
  assign new_n2414_ = new_n2413_ | new_n4396_;
  assign new_n2415_ = new_n2414_ & new_n4397_;
  assign new_n2416_ = new_n2415_ & new_n1279_;
  assign new_n2417_ = new_n1776_ & new_n1770_;
  assign new_n2418_ = new_n1775_ | new_n1769_;
  assign new_n2419_ = new_n1780_ & new_n1771_;
  assign new_n2420_ = new_n1779_ | new_n1772_;
  assign new_n2421_ = new_n4398_ & new_n4399_;
  assign new_n2422_ = new_n4400_ | new_n4401_;
  assign new_n2423_ = new_n4400_ & new_n4401_;
  assign new_n2424_ = new_n4398_ | new_n4399_;
  assign new_n2425_ = new_n2424_ & new_n2422_;
  assign new_n2426_ = new_n2423_ | new_n2421_;
  assign new_n2427_ = new_n1797_ & new_n1689_;
  assign new_n2428_ = new_n1798_ | new_n1690_;
  assign new_n2429_ = new_n1796_ & new_n1692_;
  assign new_n2430_ = new_n1795_ | new_n1691_;
  assign new_n2431_ = new_n2430_ & new_n2428_;
  assign new_n2432_ = new_n2429_ | new_n2427_;
  assign new_n2433_ = new_n4402_ & new_n4403_;
  assign new_n2434_ = new_n4404_ | new_n4405_;
  assign new_n2435_ = new_n4404_ & new_n4405_;
  assign new_n2436_ = new_n4402_ | new_n4403_;
  assign new_n2437_ = new_n2436_ & new_n2434_;
  assign new_n2438_ = new_n2435_ | new_n2433_;
  assign new_n2439_ = new_n4396_ & new_n1339_;
  assign new_n2440_ = new_n2411_ | new_n1340_;
  assign new_n2441_ = new_n4406_ & new_n4408_;
  assign new_n2442_ = new_n4410_ | new_n4412_;
  assign new_n2443_ = new_n2441_ & new_n4415_;
  assign new_n2444_ = new_n2442_ | new_n4418_;
  assign new_n2445_ = new_n4420_ & new_n4421_;
  assign new_n2446_ = new_n4422_ | new_n4423_;
  assign new_n2447_ = new_n4422_ & new_n4423_;
  assign new_n2448_ = new_n4420_ | new_n4421_;
  assign new_n2449_ = new_n2448_ & new_n2446_;
  assign new_n2450_ = new_n2447_ | new_n2445_;
  assign new_n2451_ = new_n4424_ & new_n4408_;
  assign new_n2452_ = new_n4425_ | new_n4412_;
  assign new_n2453_ = new_n2451_ & new_n4418_;
  assign new_n2454_ = new_n2452_ | new_n4415_;
  assign new_n2455_ = new_n4426_ & new_n4427_;
  assign new_n2456_ = new_n4428_ | new_n4429_;
  assign new_n2457_ = new_n4428_ & new_n4429_;
  assign new_n2458_ = new_n4426_ | new_n4427_;
  assign new_n2459_ = new_n2458_ & new_n2456_;
  assign new_n2460_ = new_n2457_ | new_n2455_;
  assign new_n2461_ = new_n4430_ & new_n4406_;
  assign new_n2462_ = new_n4431_ | new_n4410_;
  assign new_n2463_ = new_n2461_ & new_n4419_;
  assign new_n2464_ = new_n2462_ | new_n4416_;
  assign new_n2465_ = new_n4430_ & new_n4424_;
  assign new_n2466_ = new_n4431_ | new_n4425_;
  assign new_n2467_ = new_n2465_ & new_n4416_;
  assign new_n2468_ = new_n2466_ | new_n4419_;
  assign new_n2469_ = new_n2454_ & new_n2444_;
  assign new_n2470_ = new_n2453_ | new_n2443_;
  assign new_n2471_ = new_n2469_ & new_n2464_;
  assign new_n2472_ = new_n2470_ | new_n2463_;
  assign new_n2473_ = new_n2471_ & new_n2468_;
  assign new_n2474_ = new_n2472_ | new_n2467_;
  assign new_n2475_ = new_n2474_ & new_n4432_;
  assign new_n2476_ = new_n2473_ & new_n4433_;
  assign new_n2477_ = new_n2476_ | new_n2475_;
  assign new_n2478_ = new_n4434_ & new_n4435_;
  assign new_n2479_ = new_n4436_ | new_n4437_;
  assign new_n2480_ = new_n4436_ & new_n4437_;
  assign new_n2481_ = new_n4434_ | new_n4435_;
  assign new_n2482_ = new_n2481_ & new_n2479_;
  assign new_n2483_ = new_n2480_ | new_n2478_;
  assign new_n2484_ = new_n4438_ & new_n4409_;
  assign new_n2485_ = new_n4439_ | new_n4413_;
  assign new_n2486_ = new_n4439_ & new_n4413_;
  assign new_n2487_ = new_n4438_ | new_n4409_;
  assign new_n2488_ = new_n2487_ & new_n2485_;
  assign new_n2489_ = new_n2486_ | new_n2484_;
  assign new_n2490_ = new_n2489_ | new_n4433_;
  assign new_n2491_ = new_n2488_ | new_n4432_;
  assign new_n2492_ = new_n2491_ & new_n2490_;
  assign new_n2493_ = new_n4440_ | new_n1633_;
  assign new_n2494_ = new_n1976_ & new_n1809_;
  assign new_n2495_ = new_n1978_ & new_n1807_;
  assign new_n2496_ = new_n2495_ | new_n2494_;
  assign new_n2497_ = new_n1983_ | new_n1814_;
  assign new_n2498_ = new_n1981_ | new_n1816_;
  assign new_n2499_ = new_n2498_ & new_n2497_;
  assign new_n2500_ = new_n4442_ & new_n4443_;
  assign new_n2501_ = new_n4445_ | new_n4448_;
  assign new_n2502_ = new_n2500_ & new_n1752_;
  assign new_n2503_ = new_n2501_ | new_n4449_;
  assign new_n2504_ = new_n2502_ & new_n4451_;
  assign new_n2505_ = new_n2503_ | new_n4453_;
  assign new_n2506_ = new_n2200_ & new_n2196_;
  assign new_n2507_ = new_n2199_ | new_n2195_;
  assign new_n2508_ = new_n2506_ & new_n2198_;
  assign new_n2509_ = new_n2507_ | new_n2197_;
  assign new_n2510_ = new_n2508_ & new_n2214_;
  assign new_n2511_ = new_n2509_ | new_n2213_;
  assign new_n2512_ = new_n1980_ & new_n1783_;
  assign new_n2513_ = new_n1979_ | new_n1784_;
  assign new_n2514_ = new_n1954_ & new_n1811_;
  assign new_n2515_ = new_n1953_ | new_n1812_;
  assign new_n2516_ = new_n2515_ & new_n2513_;
  assign new_n2517_ = new_n2514_ | new_n2512_;
  assign new_n2518_ = new_n4454_ & new_n4455_;
  assign new_n2519_ = new_n4456_ | new_n4458_;
  assign new_n2520_ = new_n2518_ & new_n1405_;
  assign new_n2521_ = new_n2519_ | new_n1406_;
  assign new_n2522_ = new_n2521_ & new_n1404_;
  assign new_n2523_ = new_n2520_ | new_n4459_;
  assign new_n2524_ = new_n4461_ & new_n4462_;
  assign new_n2525_ = new_n1968_ & new_n1800_;
  assign new_n2526_ = new_n1967_ | new_n1799_;
  assign new_n2527_ = new_n1963_ & new_n1801_;
  assign new_n2528_ = new_n1964_ | new_n1802_;
  assign new_n2529_ = new_n2528_ & new_n2526_;
  assign new_n2530_ = new_n2527_ | new_n2525_;
  assign new_n2531_ = new_n4464_ | new_n4467_;
  assign new_n2532_ = new_n4471_ & new_n4472_;
  assign new_n2533_ = new_n4473_ | new_n4474_;
  assign new_n2534_ = new_n4473_ & new_n4474_;
  assign new_n2535_ = new_n4471_ | new_n4472_;
  assign new_n2536_ = new_n2535_ & new_n2533_;
  assign new_n2537_ = new_n2534_ | new_n2532_;
  assign new_n2538_ = new_n4476_ | new_n4467_;
  assign new_n2539_ = new_n1818_ | new_n1781_;
  assign new_n2540_ = new_n1817_ | new_n1782_;
  assign new_n2541_ = new_n2540_ & new_n2539_;
  assign new_n2542_ = new_n4477_ | new_n4468_;
  assign new_n2543_ = new_n2089_ | new_n4479_;
  assign new_n2544_ = new_n2109_ | new_n4482_;
  assign new_n2545_ = new_n2030_ | new_n4487_;
  assign new_n2546_ = new_n2049_ | new_n4492_;
  assign new_n2547_ = new_n2129_ | new_n4497_;
  assign new_n2548_ = new_n1989_ | new_n4502_;
  assign new_n2549_ = new_n2070_ | new_n4506_;
  assign new_n2550_ = new_n2009_ | new_n4509_;
  assign new_n2551_ = new_n2544_ & new_n2543_;
  assign new_n2552_ = new_n2551_ & new_n2545_;
  assign new_n2553_ = new_n2552_ & new_n2546_;
  assign new_n2554_ = new_n2553_ & new_n2547_;
  assign new_n2555_ = new_n2554_ & new_n2548_;
  assign new_n2556_ = new_n2555_ & new_n2549_;
  assign new_n2557_ = new_n2556_ & new_n2550_;
  assign new_n2558_ = new_n2557_ & new_n4514_;
  assign new_n2559_ = new_n2099_ | new_n4520_;
  assign new_n2560_ = new_n2119_ | new_n4524_;
  assign new_n2561_ = new_n2040_ | new_n4529_;
  assign new_n2562_ = new_n2059_ | new_n4534_;
  assign new_n2563_ = new_n2139_ | new_n4540_;
  assign new_n2564_ = new_n1999_ | new_n4545_;
  assign new_n2565_ = new_n2080_ | new_n4551_;
  assign new_n2566_ = new_n2019_ | new_n4556_;
  assign new_n2567_ = new_n2560_ & new_n2559_;
  assign new_n2568_ = new_n2567_ & new_n2561_;
  assign new_n2569_ = new_n2568_ & new_n2562_;
  assign new_n2570_ = new_n2569_ & new_n2563_;
  assign new_n2571_ = new_n2570_ & new_n2564_;
  assign new_n2572_ = new_n2571_ & new_n2565_;
  assign new_n2573_ = new_n2572_ & new_n2566_;
  assign new_n2574_ = new_n2573_ & new_n4561_;
  assign new_n2575_ = new_n2574_ | new_n2558_;
  assign new_n2576_ = new_n1891_ & new_n1462_;
  assign new_n2577_ = new_n1892_ | new_n1461_;
  assign new_n2578_ = new_n4443_ & new_n4458_;
  assign new_n2579_ = new_n4448_ | new_n4455_;
  assign new_n2580_ = new_n2578_ & new_n2577_;
  assign new_n2581_ = new_n2579_ | new_n2576_;
  assign new_n2582_ = new_n4568_ & new_n2575_;
  assign new_n2583_ = new_n1901_ | new_n1899_;
  assign new_n2584_ = new_n1902_ | new_n1900_;
  assign new_n2585_ = new_n2584_ & new_n2583_;
  assign new_n2586_ = new_n4442_ & new_n4573_;
  assign new_n2587_ = new_n4445_ | new_n4576_;
  assign new_n2588_ = new_n4579_ & new_n2585_;
  assign new_n2589_ = new_n2587_ & new_n4582_;
  assign new_n2590_ = new_n4585_ & new_n1558_;
  assign new_n2591_ = new_n2588_ | new_n2582_;
  assign new_n2592_ = new_n2591_ | new_n2590_;
  assign new_n2593_ = new_n4468_ & new_n4589_;
  assign new_n2594_ = new_n4461_ | new_n4595_;
  assign new_n2595_ = new_n4598_ | new_n2592_;
  assign new_n2596_ = new_n1986_ | new_n1951_;
  assign new_n2597_ = new_n1985_ | new_n1952_;
  assign new_n2598_ = new_n2597_ & new_n2596_;
  assign new_n2599_ = new_n2598_ | new_n4602_;
  assign new_n2600_ = new_n4464_ | new_n4603_;
  assign new_n2601_ = new_n2600_ | new_n4477_;
  assign new_n2602_ = new_n2601_ | new_n4605_;
  assign new_n2603_ = new_n2602_ & new_n2599_;
  assign new_n2604_ = new_n2603_ | new_n4589_;
  assign new_n2605_ = new_n1693_ & new_n4607_;
  assign new_n2606_ = new_n1694_ & new_n4608_;
  assign new_n2607_ = new_n2606_ | new_n2605_;
  assign new_n2608_ = new_n4609_ & new_n4460_;
  assign new_n2609_ = new_n4609_ & new_n4595_;
  assign new_n2610_ = new_n2530_ & new_n4605_;
  assign new_n2611_ = new_n4463_ | new_n4602_;
  assign new_n2612_ = new_n2610_ & new_n4462_;
  assign new_n2613_ = new_n2611_ & new_n4603_;
  assign new_n2614_ = new_n2613_ | new_n2612_;
  assign new_n2615_ = new_n2614_ & new_n4594_;
  assign new_n2616_ = new_n2091_ | new_n4506_;
  assign new_n2617_ = new_n2111_ | new_n4524_;
  assign new_n2618_ = new_n2032_ | new_n4612_;
  assign new_n2619_ = new_n2051_ | new_n4482_;
  assign new_n2620_ = new_n2131_ | new_n4487_;
  assign new_n2621_ = new_n1991_ | new_n4492_;
  assign new_n2622_ = new_n2072_ | new_n4497_;
  assign new_n2623_ = new_n2011_ | new_n4502_;
  assign new_n2624_ = new_n2617_ & new_n2616_;
  assign new_n2625_ = new_n2624_ & new_n2618_;
  assign new_n2626_ = new_n2625_ & new_n2619_;
  assign new_n2627_ = new_n2626_ & new_n2620_;
  assign new_n2628_ = new_n2627_ & new_n2621_;
  assign new_n2629_ = new_n2628_ & new_n2622_;
  assign new_n2630_ = new_n2629_ & new_n2623_;
  assign new_n2631_ = new_n2630_ & new_n4514_;
  assign new_n2632_ = new_n2101_ | new_n4615_;
  assign new_n2633_ = new_n2121_ | new_n4534_;
  assign new_n2634_ = new_n2042_ | new_n4540_;
  assign new_n2635_ = new_n2061_ | new_n4545_;
  assign new_n2636_ = new_n2141_ | new_n4551_;
  assign new_n2637_ = new_n2001_ | new_n4556_;
  assign new_n2638_ = new_n2082_ | new_n4520_;
  assign new_n2639_ = new_n2021_ | new_n4617_;
  assign new_n2640_ = new_n2633_ & new_n2632_;
  assign new_n2641_ = new_n2640_ & new_n2634_;
  assign new_n2642_ = new_n2641_ & new_n2635_;
  assign new_n2643_ = new_n2642_ & new_n2636_;
  assign new_n2644_ = new_n2643_ & new_n2637_;
  assign new_n2645_ = new_n2644_ & new_n2638_;
  assign new_n2646_ = new_n2645_ & new_n2639_;
  assign new_n2647_ = new_n2646_ & new_n4561_;
  assign new_n2648_ = new_n2647_ | new_n2631_;
  assign new_n2649_ = new_n2648_ & new_n4568_;
  assign new_n2650_ = new_n1915_ | new_n1911_;
  assign new_n2651_ = new_n1916_ | new_n1912_;
  assign new_n2652_ = new_n2651_ & new_n2650_;
  assign new_n2653_ = new_n4441_ & new_n4454_;
  assign new_n2654_ = new_n4446_ | new_n4456_;
  assign new_n2655_ = new_n2653_ & new_n4573_;
  assign new_n2656_ = new_n2654_ | new_n4576_;
  assign new_n2657_ = new_n4619_ & new_n2652_;
  assign new_n2658_ = new_n4620_ & new_n4513_;
  assign new_n2659_ = new_n4621_ | new_n4560_;
  assign new_n2660_ = new_n4623_ & new_n4624_;
  assign new_n2661_ = new_n4620_ & new_n4577_;
  assign new_n2662_ = new_n4621_ | new_n4574_;
  assign new_n2663_ = new_n4626_ & new_n4628_;
  assign new_n2664_ = new_n4630_ | new_n4623_;
  assign new_n2665_ = new_n4631_ & new_n1638_;
  assign new_n2666_ = new_n4630_ | new_n2660_;
  assign new_n2667_ = new_n2666_ | new_n2665_;
  assign new_n2668_ = new_n4633_ & new_n4582_;
  assign new_n2669_ = new_n4619_ | new_n4569_;
  assign new_n2670_ = new_n4634_ & new_n2667_;
  assign new_n2671_ = new_n2657_ | new_n2649_;
  assign new_n2672_ = new_n2671_ | new_n2670_;
  assign new_n2673_ = new_n2672_ | new_n4598_;
  assign new_n2674_ = new_n2094_ & new_n1867_;
  assign new_n2675_ = new_n2114_ & new_n4635_;
  assign new_n2676_ = new_n2033_ & new_n4636_;
  assign new_n2677_ = new_n2054_ & new_n4637_;
  assign new_n2678_ = new_n2134_ & new_n4638_;
  assign new_n2679_ = new_n1994_ & new_n4639_;
  assign new_n2680_ = new_n2073_ & new_n4640_;
  assign new_n2681_ = new_n2014_ & new_n1475_;
  assign new_n2682_ = new_n2675_ | new_n2674_;
  assign new_n2683_ = new_n2682_ | new_n2676_;
  assign new_n2684_ = new_n2683_ | new_n2677_;
  assign new_n2685_ = new_n2684_ | new_n2678_;
  assign new_n2686_ = new_n2685_ | new_n2679_;
  assign new_n2687_ = new_n2686_ | new_n2680_;
  assign new_n2688_ = new_n2687_ | new_n2681_;
  assign new_n2689_ = new_n2688_ | new_n4562_;
  assign new_n2690_ = new_n2104_ & new_n4641_;
  assign new_n2691_ = new_n2124_ & new_n4642_;
  assign new_n2692_ = new_n2043_ & new_n1898_;
  assign new_n2693_ = new_n2064_ & new_n4643_;
  assign new_n2694_ = new_n2144_ & new_n4644_;
  assign new_n2695_ = new_n2004_ & new_n4645_;
  assign new_n2696_ = new_n2083_ & new_n4646_;
  assign new_n2697_ = new_n2024_ & new_n4647_;
  assign new_n2698_ = new_n2691_ | new_n2690_;
  assign new_n2699_ = new_n2698_ | new_n2692_;
  assign new_n2700_ = new_n2699_ | new_n2693_;
  assign new_n2701_ = new_n2700_ | new_n2694_;
  assign new_n2702_ = new_n2701_ | new_n2695_;
  assign new_n2703_ = new_n2702_ | new_n2696_;
  assign new_n2704_ = new_n2703_ | new_n2697_;
  assign new_n2705_ = new_n2704_ | new_n4515_;
  assign new_n2706_ = new_n2705_ & new_n2689_;
  assign new_n2707_ = new_n2706_ | new_n4583_;
  assign new_n2708_ = new_n1910_ & new_n1908_;
  assign new_n2709_ = new_n1909_ & new_n1907_;
  assign new_n2710_ = new_n2709_ | new_n2708_;
  assign new_n2711_ = new_n2710_ | new_n4633_;
  assign new_n2712_ = new_n4628_ | new_n4648_;
  assign new_n2713_ = new_n4649_ | new_n4440_;
  assign new_n2714_ = new_n2712_ & new_n4626_;
  assign new_n2715_ = new_n2714_ & new_n2713_;
  assign new_n2716_ = new_n2715_ | new_n4650_;
  assign new_n2717_ = new_n2711_ & new_n2707_;
  assign new_n2718_ = new_n2717_ & new_n2716_;
  assign new_n2719_ = new_n2718_ & new_n4651_;
  assign new_n2720_ = new_n2095_ | new_n4498_;
  assign new_n2721_ = new_n2115_ | new_n4535_;
  assign new_n2722_ = new_n2036_ | new_n4529_;
  assign new_n2723_ = new_n2055_ | new_n4525_;
  assign new_n2724_ = new_n2135_ | new_n4612_;
  assign new_n2725_ = new_n1995_ | new_n4483_;
  assign new_n2726_ = new_n2076_ | new_n4488_;
  assign new_n2727_ = new_n2015_ | new_n4493_;
  assign new_n2728_ = new_n2721_ & new_n2720_;
  assign new_n2729_ = new_n2728_ & new_n2722_;
  assign new_n2730_ = new_n2729_ & new_n2723_;
  assign new_n2731_ = new_n2730_ & new_n2724_;
  assign new_n2732_ = new_n2731_ & new_n2725_;
  assign new_n2733_ = new_n2732_ & new_n2726_;
  assign new_n2734_ = new_n2733_ & new_n2727_;
  assign new_n2735_ = new_n2734_ & new_n4515_;
  assign new_n2736_ = new_n2105_ | new_n1876_;
  assign new_n2737_ = new_n2125_ | new_n4546_;
  assign new_n2738_ = new_n2046_ | new_n4552_;
  assign new_n2739_ = new_n2065_ | new_n4555_;
  assign new_n2740_ = new_n2145_ | new_n4521_;
  assign new_n2741_ = new_n2005_ | new_n4617_;
  assign new_n2742_ = new_n2086_ | new_n4615_;
  assign new_n2743_ = new_n2025_ | new_n1874_;
  assign new_n2744_ = new_n2737_ & new_n2736_;
  assign new_n2745_ = new_n2744_ & new_n2738_;
  assign new_n2746_ = new_n2745_ & new_n2739_;
  assign new_n2747_ = new_n2746_ & new_n2740_;
  assign new_n2748_ = new_n2747_ & new_n2741_;
  assign new_n2749_ = new_n2748_ & new_n2742_;
  assign new_n2750_ = new_n2749_ & new_n2743_;
  assign new_n2751_ = new_n2750_ & new_n4562_;
  assign new_n2752_ = new_n2751_ | new_n2735_;
  assign new_n2753_ = new_n2752_ & new_n4569_;
  assign new_n2754_ = new_n1905_ | new_n1903_;
  assign new_n2755_ = new_n1906_ | new_n1904_;
  assign new_n2756_ = new_n2755_ & new_n2754_;
  assign new_n2757_ = new_n2756_ & new_n4618_;
  assign new_n2758_ = new_n1987_ | new_n1971_;
  assign new_n2759_ = new_n1888_ | new_n1804_;
  assign new_n2760_ = new_n2759_ & new_n2758_;
  assign new_n2761_ = new_n2760_ & new_n4622_;
  assign new_n2762_ = new_n1709_ | new_n4652_;
  assign new_n2763_ = new_n2762_ & new_n4629_;
  assign new_n2764_ = new_n4631_ & new_n1634_;
  assign new_n2765_ = new_n2763_ | new_n2761_;
  assign new_n2766_ = new_n2765_ | new_n2764_;
  assign new_n2767_ = new_n2766_ & new_n4634_;
  assign new_n2768_ = new_n2757_ | new_n2753_;
  assign new_n2769_ = new_n2768_ | new_n2767_;
  assign new_n2770_ = new_n2769_ | new_n4599_;
  assign new_n2771_ = new_n2098_ & new_n4640_;
  assign new_n2772_ = new_n2118_ & new_n4642_;
  assign new_n2773_ = new_n2037_ & new_n1890_;
  assign new_n2774_ = new_n2058_ & new_n4635_;
  assign new_n2775_ = new_n2138_ & new_n4636_;
  assign new_n2776_ = new_n1998_ & new_n4637_;
  assign new_n2777_ = new_n2077_ & new_n4638_;
  assign new_n2778_ = new_n2018_ & new_n4639_;
  assign new_n2779_ = new_n2772_ | new_n2771_;
  assign new_n2780_ = new_n2779_ | new_n2773_;
  assign new_n2781_ = new_n2780_ | new_n2774_;
  assign new_n2782_ = new_n2781_ | new_n2775_;
  assign new_n2783_ = new_n2782_ | new_n2776_;
  assign new_n2784_ = new_n2783_ | new_n2777_;
  assign new_n2785_ = new_n2784_ | new_n2778_;
  assign new_n2786_ = new_n2785_ | new_n4564_;
  assign new_n2787_ = new_n2108_ & new_n1877_;
  assign new_n2788_ = new_n2128_ & new_n4643_;
  assign new_n2789_ = new_n2047_ & new_n4644_;
  assign new_n2790_ = new_n2068_ & new_n4645_;
  assign new_n2791_ = new_n2148_ & new_n4646_;
  assign new_n2792_ = new_n2008_ & new_n4647_;
  assign new_n2793_ = new_n2087_ & new_n4641_;
  assign new_n2794_ = new_n2028_ & new_n1875_;
  assign new_n2795_ = new_n2788_ | new_n2787_;
  assign new_n2796_ = new_n2795_ | new_n2789_;
  assign new_n2797_ = new_n2796_ | new_n2790_;
  assign new_n2798_ = new_n2797_ | new_n2791_;
  assign new_n2799_ = new_n2798_ | new_n2792_;
  assign new_n2800_ = new_n2799_ | new_n2793_;
  assign new_n2801_ = new_n2800_ | new_n2794_;
  assign new_n2802_ = new_n2801_ | new_n4517_;
  assign new_n2803_ = new_n2802_ & new_n2786_;
  assign new_n2804_ = new_n2803_ | new_n4583_;
  assign new_n2805_ = new_n1918_ & new_n1914_;
  assign new_n2806_ = new_n1917_ & new_n1913_;
  assign new_n2807_ = new_n2806_ | new_n2805_;
  assign new_n2808_ = new_n2807_ | new_n4632_;
  assign new_n2809_ = new_n1974_ & new_n1966_;
  assign new_n2810_ = new_n4653_ & new_n1805_;
  assign new_n2811_ = new_n2810_ | new_n2809_;
  assign new_n2812_ = new_n2811_ | new_n4627_;
  assign new_n2813_ = new_n4654_ & new_n4655_;
  assign new_n2814_ = new_n2813_ | new_n4625_;
  assign new_n2815_ = new_n4649_ | new_n4652_;
  assign new_n2816_ = new_n2814_ & new_n2812_;
  assign new_n2817_ = new_n2816_ & new_n2815_;
  assign new_n2818_ = new_n2817_ | new_n4650_;
  assign new_n2819_ = new_n2808_ & new_n2804_;
  assign new_n2820_ = new_n2819_ & new_n2818_;
  assign new_n2821_ = new_n2820_ & new_n4651_;
  assign new_n2822_ = new_n1940_ & new_n1935_;
  assign new_n2823_ = new_n1939_ | new_n1936_;
  assign new_n2824_ = new_n2823_ & new_n4657_;
  assign new_n2825_ = new_n2822_ & new_n4659_;
  assign new_n2826_ = new_n2825_ | new_n2824_;
  assign new_n2827_ = new_n2826_ | new_n4590_;
  assign new_n2828_ = new_n1938_ & new_n1933_;
  assign new_n2829_ = new_n1937_ | new_n1934_;
  assign new_n2830_ = new_n2829_ & new_n4604_;
  assign new_n2831_ = new_n2828_ & new_n4601_;
  assign new_n2832_ = new_n2831_ | new_n2830_;
  assign new_n2833_ = new_n2832_ | new_n4590_;
  assign new_n2834_ = new_n4660_ & new_n1716_;
  assign new_n2835_ = new_n1724_ | new_n1715_;
  assign new_n2836_ = new_n4661_ & new_n4662_;
  assign new_n2837_ = new_n4663_ | new_n1726_;
  assign new_n2838_ = new_n4666_ & new_n4671_;
  assign new_n2839_ = new_n4674_ | new_n2510_;
  assign new_n2840_ = new_n1788_ & new_n1786_;
  assign new_n2841_ = new_n1787_ | new_n1785_;
  assign new_n2842_ = new_n2178_ & new_n2176_;
  assign new_n2843_ = new_n2177_ | new_n2175_;
  assign new_n2844_ = new_n2842_ & new_n2194_;
  assign new_n2845_ = new_n2843_ | new_n2193_;
  assign new_n2846_ = new_n2845_ & new_n2840_;
  assign new_n2847_ = new_n2844_ | new_n2841_;
  assign new_n2848_ = new_n4680_ & new_n4683_;
  assign new_n2849_ = new_n4686_ | new_n4688_;
  assign new_n2850_ = new_n2848_ & new_n2151_;
  assign new_n2851_ = new_n2849_ | new_n2152_;
  assign new_n2852_ = new_n2850_ & new_n4690_;
  assign new_n2853_ = new_n2851_ | new_n4693_;
  assign new_n2854_ = new_n2224_ & new_n1960_;
  assign new_n2855_ = new_n2223_ | new_n1959_;
  assign new_n2856_ = new_n2215_ & new_n2159_;
  assign new_n2857_ = new_n2216_ | new_n2160_;
  assign new_n2858_ = new_n2857_ & new_n2855_;
  assign new_n2859_ = new_n2856_ | new_n2854_;
  assign new_n2860_ = new_n4694_ & new_n4695_;
  assign new_n2861_ = new_n4696_ | new_n4697_;
  assign new_n2862_ = new_n4696_ & new_n4697_;
  assign new_n2863_ = new_n4694_ | new_n4695_;
  assign new_n2864_ = new_n2863_ & new_n2861_;
  assign new_n2865_ = new_n2862_ | new_n2860_;
  assign new_n2866_ = new_n4699_ | new_n4470_;
  assign new_n2867_ = new_n4701_ & new_n4702_;
  assign new_n2868_ = new_n4704_ | new_n1668_;
  assign new_n2869_ = new_n2867_ & new_n4705_;
  assign new_n2870_ = new_n2868_ | new_n4706_;
  assign new_n2871_ = new_n4701_ & new_n4707_;
  assign new_n2872_ = new_n4704_ | new_n4708_;
  assign new_n2873_ = new_n2871_ & new_n4709_;
  assign new_n2874_ = new_n2872_ | new_n4710_;
  assign new_n2875_ = new_n2874_ & new_n2870_;
  assign new_n2876_ = new_n2873_ | new_n2869_;
  assign new_n2877_ = new_n4712_ & new_n4713_;
  assign new_n2878_ = new_n4715_ | new_n4716_;
  assign new_n2879_ = new_n2877_ & new_n4709_;
  assign new_n2880_ = new_n2878_ | new_n4710_;
  assign new_n2881_ = new_n4712_ & new_n4717_;
  assign new_n2882_ = new_n4715_ | new_n4719_;
  assign new_n2883_ = new_n2881_ & new_n4705_;
  assign new_n2884_ = new_n2882_ | new_n4706_;
  assign new_n2885_ = new_n2884_ & new_n2880_;
  assign new_n2886_ = new_n2883_ | new_n2879_;
  assign new_n2887_ = new_n2885_ & new_n4711_;
  assign new_n2888_ = new_n2886_ | new_n4714_;
  assign new_n2889_ = new_n2888_ & new_n2875_;
  assign new_n2890_ = new_n2887_ | new_n4720_;
  assign new_n2891_ = new_n4723_ & new_n4726_;
  assign new_n2892_ = new_n4728_ | new_n2154_;
  assign new_n2893_ = new_n2892_ | new_n1852_;
  assign new_n2894_ = new_n2893_ | new_n1742_;
  assign new_n2895_ = new_n1970_ | new_n1921_;
  assign new_n2896_ = new_n1969_ | new_n1922_;
  assign new_n2897_ = new_n2896_ & new_n2895_;
  assign new_n2898_ = new_n4730_ | new_n4470_;
  assign new_n2899_ = new_n4700_ & new_n1929_;
  assign new_n2900_ = new_n4703_ | new_n1930_;
  assign new_n2901_ = new_n4731_ | new_n4732_;
  assign new_n2902_ = new_n2901_ | new_n4733_;
  assign new_n2903_ = new_n4734_ & new_n4735_;
  assign new_n2904_ = new_n2903_ & new_n4736_;
  assign new_n2905_ = new_n4737_ & new_n4738_;
  assign new_n2906_ = new_n2905_ & new_n4739_;
  assign new_n2907_ = new_n4740_ & new_n4741_;
  assign new_n2908_ = new_n2907_ & new_n4742_;
  assign new_n2909_ = new_n4607_ & new_n1608_;
  assign new_n2910_ = new_n4608_ | new_n1607_;
  assign new_n2911_ = new_n4743_ & new_n4744_;
  assign new_n2912_ = new_n4745_ | new_n4746_;
  assign new_n2913_ = new_n4745_ & new_n4746_;
  assign new_n2914_ = new_n4743_ | new_n4744_;
  assign new_n2915_ = new_n2914_ & new_n2912_;
  assign new_n2916_ = new_n2913_ | new_n2911_;
  assign new_n2917_ = new_n2916_ | new_n2910_;
  assign new_n2918_ = new_n2915_ | new_n2909_;
  assign new_n2919_ = new_n2918_ & new_n2917_;
  assign new_n2920_ = new_n4747_ | new_n4469_;
  assign new_n2921_ = new_n4749_ | new_n1242_;
  assign new_n2922_ = new_n4751_ | new_n4493_;
  assign new_n2923_ = new_n4753_ | new_n4498_;
  assign new_n2924_ = new_n4501_ | new_n4755_;
  assign new_n2925_ = new_n4505_ | new_n4757_;
  assign new_n2926_ = new_n4509_ | new_n4759_;
  assign new_n2927_ = new_n4479_ | new_n4761_;
  assign new_n2928_ = new_n4763_ | new_n4764_;
  assign new_n2929_ = new_n2922_ & new_n2921_;
  assign new_n2930_ = new_n2929_ & new_n2923_;
  assign new_n2931_ = new_n2930_ & new_n2924_;
  assign new_n2932_ = new_n2931_ & new_n2925_;
  assign new_n2933_ = new_n2932_ & new_n2926_;
  assign new_n2934_ = new_n2933_ & new_n2927_;
  assign new_n2935_ = new_n2934_ & new_n2928_;
  assign new_n2936_ = new_n4451_ & new_n4574_;
  assign new_n2937_ = new_n4453_ | new_n4577_;
  assign new_n2938_ = new_n2936_ & new_n2935_;
  assign new_n2939_ = new_n4766_ | new_n4552_;
  assign new_n2940_ = new_n4483_ | new_n4768_;
  assign new_n2941_ = new_n4613_ | new_n4770_;
  assign new_n2942_ = new_n4525_ | new_n4772_;
  assign new_n2943_ = new_n4530_ | new_n4774_;
  assign new_n2944_ = new_n4535_ | new_n4776_;
  assign new_n2945_ = new_n4541_ | new_n4778_;
  assign new_n2946_ = new_n4546_ | new_n4780_;
  assign new_n2947_ = new_n2940_ & new_n2939_;
  assign new_n2948_ = new_n2947_ & new_n2941_;
  assign new_n2949_ = new_n2948_ & new_n2942_;
  assign new_n2950_ = new_n2949_ & new_n2943_;
  assign new_n2951_ = new_n2950_ & new_n2944_;
  assign new_n2952_ = new_n2951_ & new_n2945_;
  assign new_n2953_ = new_n2952_ & new_n2946_;
  assign new_n2954_ = new_n4517_ & new_n4450_;
  assign new_n2955_ = new_n4564_ | new_n4452_;
  assign new_n2956_ = new_n2954_ & new_n2953_;
  assign new_n2957_ = new_n2955_ & new_n2937_;
  assign new_n2958_ = new_n2957_ & new_n4781_;
  assign new_n2959_ = new_n2956_ | new_n2938_;
  assign new_n2960_ = new_n2959_ | new_n2958_;
  assign new_n2961_ = new_n2960_ & new_n4571_;
  assign new_n2962_ = new_n1595_ | new_n1569_;
  assign new_n2963_ = new_n1596_ | new_n1570_;
  assign new_n2964_ = new_n2963_ & new_n2962_;
  assign new_n2965_ = new_n2964_ & new_n4579_;
  assign new_n2966_ = new_n4585_ & new_n4781_;
  assign new_n2967_ = new_n2965_ | new_n2961_;
  assign new_n2968_ = new_n2967_ | new_n2966_;
  assign new_n2969_ = new_n2968_ | new_n4599_;
  assign new_n2970_ = new_n4749_ | new_n4764_;
  assign new_n2971_ = new_n4751_ | new_n4488_;
  assign new_n2972_ = new_n4753_ | new_n4494_;
  assign new_n2973_ = new_n4755_ | new_n4499_;
  assign new_n2974_ = new_n4503_ | new_n4757_;
  assign new_n2975_ = new_n4507_ | new_n4759_;
  assign new_n2976_ = new_n4510_ | new_n4761_;
  assign new_n2977_ = new_n4478_ | new_n4763_;
  assign new_n2978_ = new_n2971_ & new_n2970_;
  assign new_n2979_ = new_n2978_ & new_n2972_;
  assign new_n2980_ = new_n2979_ & new_n2973_;
  assign new_n2981_ = new_n2980_ & new_n2974_;
  assign new_n2982_ = new_n2981_ & new_n2975_;
  assign new_n2983_ = new_n2982_ & new_n2976_;
  assign new_n2984_ = new_n2983_ & new_n2977_;
  assign new_n2985_ = new_n2984_ & new_n4518_;
  assign new_n2986_ = new_n4766_ | new_n4557_;
  assign new_n2987_ = new_n4613_ | new_n4768_;
  assign new_n2988_ = new_n4526_ | new_n4770_;
  assign new_n2989_ = new_n4530_ | new_n4772_;
  assign new_n2990_ = new_n4537_ | new_n4774_;
  assign new_n2991_ = new_n4541_ | new_n4776_;
  assign new_n2992_ = new_n4548_ | new_n4778_;
  assign new_n2993_ = new_n4780_ | new_n4553_;
  assign new_n2994_ = new_n2987_ & new_n2986_;
  assign new_n2995_ = new_n2994_ & new_n2988_;
  assign new_n2996_ = new_n2995_ & new_n2989_;
  assign new_n2997_ = new_n2996_ & new_n2990_;
  assign new_n2998_ = new_n2997_ & new_n2991_;
  assign new_n2999_ = new_n2998_ & new_n2992_;
  assign new_n3000_ = new_n2999_ & new_n2993_;
  assign new_n3001_ = new_n3000_ & new_n4565_;
  assign new_n3002_ = new_n3001_ | new_n2985_;
  assign new_n3003_ = new_n3002_ & new_n4571_;
  assign new_n3004_ = new_n1489_ | new_n1487_;
  assign new_n3005_ = new_n1490_ | new_n1488_;
  assign new_n3006_ = new_n3005_ & new_n3004_;
  assign new_n3007_ = new_n3006_ & new_n4580_;
  assign new_n3008_ = new_n4586_ & new_n1560_;
  assign new_n3009_ = new_n3007_ | new_n3003_;
  assign new_n3010_ = new_n3009_ | new_n3008_;
  assign new_n3011_ = new_n3010_ | new_n4600_;
  assign new_n3012_ = new_n4510_ | new_n4748_;
  assign new_n3013_ = new_n4614_ | new_n4750_;
  assign new_n3014_ = new_n4484_ | new_n4752_;
  assign new_n3015_ = new_n4754_ | new_n4489_;
  assign new_n3016_ = new_n4756_ | new_n4494_;
  assign new_n3017_ = new_n4758_ | new_n4499_;
  assign new_n3018_ = new_n4503_ | new_n4760_;
  assign new_n3019_ = new_n4507_ | new_n4762_;
  assign new_n3020_ = new_n3013_ & new_n3012_;
  assign new_n3021_ = new_n3020_ & new_n3014_;
  assign new_n3022_ = new_n3021_ & new_n3015_;
  assign new_n3023_ = new_n3022_ & new_n3016_;
  assign new_n3024_ = new_n3023_ & new_n3017_;
  assign new_n3025_ = new_n3024_ & new_n3018_;
  assign new_n3026_ = new_n3025_ & new_n3019_;
  assign new_n3027_ = new_n3026_ & new_n4518_;
  assign new_n3028_ = new_n4616_ | new_n4765_;
  assign new_n3029_ = new_n4531_ | new_n4767_;
  assign new_n3030_ = new_n4537_ | new_n4769_;
  assign new_n3031_ = new_n4542_ | new_n4771_;
  assign new_n3032_ = new_n4548_ | new_n4773_;
  assign new_n3033_ = new_n4775_ | new_n4553_;
  assign new_n3034_ = new_n4777_ | new_n4557_;
  assign new_n3035_ = new_n4779_ | new_n4521_;
  assign new_n3036_ = new_n3029_ & new_n3028_;
  assign new_n3037_ = new_n3036_ & new_n3030_;
  assign new_n3038_ = new_n3037_ & new_n3031_;
  assign new_n3039_ = new_n3038_ & new_n3032_;
  assign new_n3040_ = new_n3039_ & new_n3033_;
  assign new_n3041_ = new_n3040_ & new_n3034_;
  assign new_n3042_ = new_n3041_ & new_n3035_;
  assign new_n3043_ = new_n3042_ & new_n4565_;
  assign new_n3044_ = new_n3043_ | new_n3027_;
  assign new_n3045_ = new_n3044_ & new_n4570_;
  assign new_n3046_ = new_n1485_ | new_n1483_;
  assign new_n3047_ = new_n1486_ | new_n1484_;
  assign new_n3048_ = new_n3047_ & new_n3046_;
  assign new_n3049_ = new_n3048_ & new_n4580_;
  assign new_n3050_ = new_n4586_ & new_n1562_;
  assign new_n3051_ = new_n3049_ | new_n3045_;
  assign new_n3052_ = new_n3051_ | new_n3050_;
  assign new_n3053_ = new_n3052_ | new_n4600_;
  assign new_n3054_ = new_n4730_ | new_n4659_;
  assign new_n3055_ = new_n4699_ | new_n4476_;
  assign new_n3056_ = new_n3055_ | new_n4729_;
  assign new_n3057_ = new_n3056_ | new_n4657_;
  assign new_n3058_ = new_n3057_ & new_n3054_;
  assign new_n3059_ = new_n3058_ | new_n4592_;
  assign new_n3060_ = new_n2537_ & new_n4656_;
  assign new_n3061_ = new_n4475_ | new_n4658_;
  assign new_n3062_ = new_n3061_ | new_n4698_;
  assign new_n3063_ = new_n3060_ | new_n2865_;
  assign new_n3064_ = new_n3063_ & new_n3062_;
  assign new_n3065_ = new_n3064_ | new_n4592_;
  assign new_n3066_ = new_n4747_ | new_n4593_;
  assign new_n3067_ = new_n4782_ | new_n4783_;
  assign new_n3068_ = new_n3067_ | new_n4784_;
  assign new_n3069_ = new_n4785_ & new_n4786_;
  assign new_n3070_ = new_n4787_ | new_n4788_;
  assign new_n3071_ = new_n3069_ & new_n4789_;
  assign new_n3072_ = new_n3070_ | new_n4790_;
  assign new_n3073_ = new_n3071_ & new_n4791_;
  assign new_n3074_ = new_n3072_ | new_n4792_;
  assign new_n3075_ = new_n3073_ & new_n4793_;
  assign new_n3076_ = new_n3074_ | new_n4794_;
  assign new_n3077_ = new_n4787_ & new_n4788_;
  assign new_n3078_ = new_n4785_ | new_n4786_;
  assign new_n3079_ = new_n3077_ & new_n4790_;
  assign new_n3080_ = new_n3078_ | new_n4789_;
  assign new_n3081_ = new_n3079_ & new_n4792_;
  assign new_n3082_ = new_n3080_ | new_n4791_;
  assign new_n3083_ = new_n3081_ & new_n4794_;
  assign new_n3084_ = new_n3082_ | new_n4793_;
  assign new_n3085_ = new_n3084_ & new_n3076_;
  assign new_n3086_ = new_n3083_ | new_n3075_;
  assign new_n3087_ = new_n3086_ & new_n4666_;
  assign new_n3088_ = new_n3085_ | new_n4674_;
  assign new_n3089_ = new_n4795_ & new_n4675_;
  assign new_n3090_ = new_n2853_ | new_n4667_;
  assign new_n3091_ = new_n3090_ & new_n3088_;
  assign new_n3092_ = new_n3089_ | new_n3087_;
  assign new_n3093_ = new_n4796_ & new_n4797_;
  assign new_n3094_ = new_n3093_ & new_n4798_;
  assign new_n3095_ = new_n4799_ & new_n4800_;
  assign new_n3096_ = new_n3095_ & new_n4801_;
  assign new_n3097_ = new_n4802_ & new_n4803_;
  assign new_n3098_ = new_n3097_ & new_n4804_;
  assign new_n3099_ = new_n1736_ & new_n1734_;
  assign new_n3100_ = new_n1735_ | new_n1733_;
  assign new_n3101_ = new_n4805_ & new_n4723_;
  assign new_n3102_ = new_n1720_ & new_n1718_;
  assign new_n3103_ = new_n1719_ | new_n1717_;
  assign new_n3104_ = new_n4806_ & new_n2891_;
  assign new_n3105_ = new_n1704_ & new_n1702_;
  assign new_n3106_ = new_n1703_ | new_n1701_;
  assign new_n3107_ = new_n4807_ & new_n4726_;
  assign new_n3108_ = new_n3107_ & new_n1851_;
  assign new_n3109_ = new_n3108_ & new_n4724_;
  assign new_n3110_ = new_n3101_ | new_n4720_;
  assign new_n3111_ = new_n3110_ | new_n3104_;
  assign new_n3112_ = new_n3111_ | new_n3109_;
  assign new_n3113_ = new_n4667_ & new_n1941_;
  assign new_n3114_ = new_n4675_ | new_n1942_;
  assign new_n3115_ = new_n4808_ & new_n4809_;
  assign new_n3116_ = new_n4811_ | new_n4813_;
  assign new_n3117_ = new_n4811_ & new_n4813_;
  assign new_n3118_ = new_n4808_ | new_n4809_;
  assign new_n3119_ = new_n3118_ & new_n3116_;
  assign new_n3120_ = new_n3117_ | new_n3115_;
  assign new_n3121_ = new_n4669_ & new_n1957_;
  assign new_n3122_ = new_n4677_ | new_n1958_;
  assign new_n3123_ = new_n4814_ & new_n4815_;
  assign new_n3124_ = new_n4817_ | new_n4819_;
  assign new_n3125_ = new_n3124_ & new_n4821_;
  assign new_n3126_ = new_n4822_ | new_n4823_;
  assign new_n3127_ = new_n4825_ & new_n4826_;
  assign new_n3128_ = new_n4827_ | new_n4829_;
  assign new_n3129_ = new_n4827_ & new_n4829_;
  assign new_n3130_ = new_n4825_ | new_n4826_;
  assign new_n3131_ = new_n3130_ & new_n3128_;
  assign new_n3132_ = new_n3129_ | new_n3127_;
  assign new_n3133_ = new_n4830_ & new_n4832_;
  assign new_n3134_ = new_n4834_ | new_n4835_;
  assign new_n3135_ = new_n4834_ & new_n4835_;
  assign new_n3136_ = new_n4830_ | new_n4832_;
  assign new_n3137_ = new_n3136_ & new_n3134_;
  assign new_n3138_ = new_n3135_ | new_n3133_;
  assign new_n3139_ = new_n4837_ & new_n4840_;
  assign new_n3140_ = new_n3139_ | new_n4843_;
  assign new_n3141_ = new_n4805_ & new_n4663_;
  assign new_n3142_ = new_n3099_ | new_n4661_;
  assign new_n3143_ = new_n4844_ & new_n4845_;
  assign new_n3144_ = new_n4847_ | new_n4849_;
  assign new_n3145_ = new_n4847_ & new_n4849_;
  assign new_n3146_ = new_n4844_ | new_n4845_;
  assign new_n3147_ = new_n3146_ & new_n3144_;
  assign new_n3148_ = new_n3145_ | new_n3143_;
  assign new_n3149_ = new_n4806_ & new_n4669_;
  assign new_n3150_ = new_n3102_ | new_n4677_;
  assign new_n3151_ = new_n4850_ & new_n4852_;
  assign new_n3152_ = new_n4853_ | new_n4855_;
  assign new_n3153_ = new_n4857_ & new_n4858_;
  assign new_n3154_ = new_n4859_ | new_n4860_;
  assign new_n3155_ = new_n4859_ & new_n4860_;
  assign new_n3156_ = new_n4857_ | new_n4858_;
  assign new_n3157_ = new_n3156_ & new_n3154_;
  assign new_n3158_ = new_n3155_ | new_n3153_;
  assign new_n3159_ = new_n4807_ & new_n4670_;
  assign new_n3160_ = new_n3105_ | new_n4678_;
  assign new_n3161_ = new_n4862_ & new_n4852_;
  assign new_n3162_ = new_n4866_ | new_n4855_;
  assign new_n3163_ = new_n4869_ & new_n4871_;
  assign new_n3164_ = new_n4872_ | new_n4874_;
  assign new_n3165_ = new_n4869_ & new_n4876_;
  assign new_n3166_ = new_n4872_ | new_n4880_;
  assign new_n3167_ = new_n3165_ & new_n4840_;
  assign new_n3168_ = new_n3166_ | new_n4884_;
  assign new_n3169_ = new_n3152_ & new_n3142_;
  assign new_n3170_ = new_n3151_ | new_n3141_;
  assign new_n3171_ = new_n3169_ & new_n3164_;
  assign new_n3172_ = new_n3170_ | new_n3163_;
  assign new_n3173_ = new_n3171_ & new_n3168_;
  assign new_n3174_ = new_n3172_ | new_n3167_;
  assign new_n3175_ = new_n4886_ & new_n4888_;
  assign new_n3176_ = new_n4889_ | new_n4891_;
  assign new_n3177_ = new_n4889_ | new_n4893_;
  assign new_n3178_ = new_n4894_ & new_n1739_;
  assign new_n3179_ = new_n4895_ | new_n1740_;
  assign new_n3180_ = new_n4896_ & new_n4693_;
  assign new_n3181_ = new_n4898_ | new_n4690_;
  assign new_n3182_ = new_n4898_ & new_n4691_;
  assign new_n3183_ = new_n4896_ | new_n4692_;
  assign new_n3184_ = new_n3183_ & new_n3181_;
  assign new_n3185_ = new_n3182_ | new_n3180_;
  assign new_n3186_ = new_n4900_ & new_n4904_;
  assign new_n3187_ = new_n2204_ | new_n4911_;
  assign new_n3188_ = new_n4915_ & new_n2184_;
  assign new_n3189_ = new_n4917_ | new_n2183_;
  assign new_n3190_ = new_n4918_ & new_n4911_;
  assign new_n3191_ = new_n4920_ | new_n4904_;
  assign new_n3192_ = new_n4924_ & new_n4930_;
  assign new_n3193_ = new_n4934_ | new_n4939_;
  assign new_n3194_ = new_n3192_ & new_n4940_;
  assign new_n3195_ = new_n3193_ | new_n4941_;
  assign new_n3196_ = new_n4924_ & new_n4942_;
  assign new_n3197_ = new_n4934_ | new_n4943_;
  assign new_n3198_ = new_n4944_ & new_n4941_;
  assign new_n3199_ = new_n4945_ | new_n4940_;
  assign new_n3200_ = new_n4948_ & new_n4953_;
  assign new_n3201_ = new_n4960_ | new_n4964_;
  assign new_n3202_ = new_n4968_ & new_n4972_;
  assign new_n3203_ = new_n4978_ | new_n4981_;
  assign new_n3204_ = new_n4964_ & new_n4981_;
  assign new_n3205_ = new_n4953_ | new_n4972_;
  assign new_n3206_ = new_n4986_ & new_n4991_;
  assign new_n3207_ = new_n4995_ | new_n4998_;
  assign new_n3208_ = new_n3203_ & new_n3201_;
  assign new_n3209_ = new_n3202_ | new_n3200_;
  assign new_n3210_ = new_n3208_ & new_n3207_;
  assign new_n3211_ = new_n3209_ | new_n3206_;
  assign new_n3212_ = new_n3211_ & new_n4923_;
  assign new_n3213_ = new_n3210_ | new_n4935_;
  assign new_n3214_ = new_n3199_ & new_n3195_;
  assign new_n3215_ = new_n3198_ | new_n3194_;
  assign new_n3216_ = new_n3214_ & new_n3213_;
  assign new_n3217_ = new_n3215_ | new_n3212_;
  assign new_n3218_ = new_n4999_ & new_n4918_;
  assign new_n3219_ = new_n5000_ | new_n4920_;
  assign new_n3220_ = new_n3218_ & new_n2162_;
  assign new_n3221_ = new_n3219_ | new_n5001_;
  assign new_n3222_ = new_n4925_ & new_n5003_;
  assign new_n3223_ = new_n4935_ | new_n5005_;
  assign new_n3224_ = new_n3222_ & new_n5007_;
  assign new_n3225_ = new_n3223_ | new_n5010_;
  assign new_n3226_ = new_n5010_ & new_n4944_;
  assign new_n3227_ = new_n5007_ | new_n4945_;
  assign new_n3228_ = new_n5012_ & new_n4954_;
  assign new_n3229_ = new_n5013_ | new_n4965_;
  assign new_n3230_ = new_n4991_ & new_n4973_;
  assign new_n3231_ = new_n4998_ | new_n4982_;
  assign new_n3232_ = new_n4986_ & new_n4930_;
  assign new_n3233_ = new_n4995_ | new_n4939_;
  assign new_n3234_ = new_n3231_ & new_n3229_;
  assign new_n3235_ = new_n3230_ | new_n3228_;
  assign new_n3236_ = new_n3234_ & new_n3233_;
  assign new_n3237_ = new_n3235_ | new_n3232_;
  assign new_n3238_ = new_n3237_ & new_n4925_;
  assign new_n3239_ = new_n3236_ | new_n4937_;
  assign new_n3240_ = new_n5014_ & new_n3225_;
  assign new_n3241_ = new_n5016_ | new_n3224_;
  assign new_n3242_ = new_n3240_ & new_n3239_;
  assign new_n3243_ = new_n3241_ | new_n3238_;
  assign new_n3244_ = new_n4927_ & new_n5018_;
  assign new_n3245_ = new_n4937_ | new_n1296_;
  assign new_n3246_ = new_n3244_ & new_n5008_;
  assign new_n3247_ = new_n3245_ | new_n5009_;
  assign new_n3248_ = new_n5019_ & new_n4954_;
  assign new_n3249_ = new_n2252_ | new_n4965_;
  assign new_n3250_ = new_n4931_ & new_n4973_;
  assign new_n3251_ = new_n4938_ | new_n4982_;
  assign new_n3252_ = new_n4987_ & new_n5003_;
  assign new_n3253_ = new_n4994_ | new_n5005_;
  assign new_n3254_ = new_n3251_ & new_n3249_;
  assign new_n3255_ = new_n3250_ | new_n3248_;
  assign new_n3256_ = new_n3254_ & new_n3253_;
  assign new_n3257_ = new_n3255_ | new_n3252_;
  assign new_n3258_ = new_n3257_ & new_n4927_;
  assign new_n3259_ = new_n3256_ | new_n4936_;
  assign new_n3260_ = new_n3247_ & new_n5014_;
  assign new_n3261_ = new_n3246_ | new_n5016_;
  assign new_n3262_ = new_n3260_ & new_n3259_;
  assign new_n3263_ = new_n3261_ | new_n3258_;
  assign new_n3264_ = new_n5023_ & new_n5030_;
  assign new_n3265_ = new_n5036_ | new_n5043_;
  assign new_n3266_ = new_n5047_ & new_n5053_;
  assign new_n3267_ = new_n5060_ | new_n5067_;
  assign new_n3268_ = new_n5036_ & new_n5067_;
  assign new_n3269_ = new_n5023_ | new_n5053_;
  assign new_n3270_ = new_n5074_ & new_n5080_;
  assign new_n3271_ = new_n5084_ | new_n5090_;
  assign new_n3272_ = new_n3267_ & new_n3265_;
  assign new_n3273_ = new_n3266_ | new_n3264_;
  assign new_n3274_ = new_n3272_ & new_n3271_;
  assign new_n3275_ = new_n3273_ | new_n3270_;
  assign new_n3276_ = new_n5095_ & new_n4905_;
  assign new_n3277_ = new_n5097_ | new_n4912_;
  assign new_n3278_ = new_n3276_ & new_n5099_;
  assign new_n3279_ = new_n3277_ | new_n5100_;
  assign new_n3280_ = new_n3279_ & new_n4917_;
  assign new_n3281_ = new_n3278_ | new_n4915_;
  assign new_n3282_ = new_n5104_ & new_n3275_;
  assign new_n3283_ = new_n5111_ | new_n3274_;
  assign new_n3284_ = new_n2275_ & new_n4912_;
  assign new_n3285_ = new_n2276_ | new_n4905_;
  assign new_n3286_ = new_n5119_ & new_n5043_;
  assign new_n3287_ = new_n5126_ | new_n5030_;
  assign new_n3288_ = new_n5095_ & new_n4913_;
  assign new_n3289_ = new_n5097_ | new_n4907_;
  assign new_n3290_ = new_n5126_ & new_n5111_;
  assign new_n3291_ = new_n5119_ | new_n5104_;
  assign new_n3292_ = new_n5132_ & new_n5031_;
  assign new_n3293_ = new_n5135_ | new_n5042_;
  assign new_n3294_ = new_n3292_ & new_n5138_;
  assign new_n3295_ = new_n3293_ | new_n5145_;
  assign new_n3296_ = new_n3287_ & new_n3283_;
  assign new_n3297_ = new_n3286_ | new_n3282_;
  assign new_n3298_ = new_n3296_ & new_n3295_;
  assign new_n3299_ = new_n3297_ | new_n3294_;
  assign new_n3300_ = new_n4914_ & new_n2262_;
  assign new_n3301_ = new_n4916_ | new_n2261_;
  assign new_n3302_ = new_n4999_ & new_n2253_;
  assign new_n3303_ = new_n5000_ | new_n2254_;
  assign new_n3304_ = new_n5152_ & new_n4992_;
  assign new_n3305_ = new_n5159_ | new_n4997_;
  assign new_n3306_ = new_n3304_ & new_n5165_;
  assign new_n3307_ = new_n3305_ | new_n5168_;
  assign new_n3308_ = new_n5152_ & new_n4942_;
  assign new_n3309_ = new_n5159_ | new_n4943_;
  assign new_n3310_ = new_n3308_ & new_n5168_;
  assign new_n3311_ = new_n3309_ | new_n5165_;
  assign new_n3312_ = new_n2284_ & new_n5172_;
  assign new_n3313_ = new_n2283_ | new_n5179_;
  assign new_n3314_ = new_n5183_ & new_n2264_;
  assign new_n3315_ = new_n5186_ | new_n2263_;
  assign new_n3316_ = new_n4968_ & new_n2265_;
  assign new_n3317_ = new_n4978_ | new_n2266_;
  assign new_n3318_ = new_n3315_ & new_n3313_;
  assign new_n3319_ = new_n3314_ | new_n3312_;
  assign new_n3320_ = new_n3318_ & new_n3317_;
  assign new_n3321_ = new_n3319_ | new_n3316_;
  assign new_n3322_ = new_n3321_ & new_n5151_;
  assign new_n3323_ = new_n3320_ | new_n5160_;
  assign new_n3324_ = new_n5188_ & new_n3307_;
  assign new_n3325_ = new_n5190_ | new_n3306_;
  assign new_n3326_ = new_n3324_ & new_n3323_;
  assign new_n3327_ = new_n3325_ | new_n3322_;
  assign new_n3328_ = new_n5194_ | new_n5198_;
  assign new_n3329_ = new_n3328_ | new_n5201_;
  assign new_n3330_ = new_n5194_ | new_n5204_;
  assign new_n3331_ = new_n3330_ | new_n5201_;
  assign new_n3332_ = new_n1617_ | new_n1615_;
  assign new_n3333_ = new_n3332_ | new_n1611_;
  assign new_n3334_ = new_n3185_ | new_n4819_;
  assign new_n3335_ = new_n5208_ & new_n4837_;
  assign new_n3336_ = new_n4900_ | new_n4907_;
  assign new_n3337_ = new_n3336_ | new_n5094_;
  assign new_n3338_ = new_n5022_ & new_n5211_;
  assign new_n3339_ = new_n5037_ | new_n5215_;
  assign new_n3340_ = new_n5052_ & new_n5031_;
  assign new_n3341_ = new_n5068_ | new_n5044_;
  assign new_n3342_ = new_n5074_ & new_n5222_;
  assign new_n3343_ = new_n5084_ | new_n5224_;
  assign new_n3344_ = new_n3341_ & new_n3339_;
  assign new_n3345_ = new_n3340_ | new_n3338_;
  assign new_n3346_ = new_n3344_ & new_n3343_;
  assign new_n3347_ = new_n3345_ | new_n3342_;
  assign new_n3348_ = new_n3347_ & new_n5103_;
  assign new_n3349_ = new_n3346_ | new_n5112_;
  assign new_n3350_ = new_n5118_ & new_n5211_;
  assign new_n3351_ = new_n5127_ | new_n5215_;
  assign new_n3352_ = new_n5132_ & new_n5216_;
  assign new_n3353_ = new_n5135_ | new_n5210_;
  assign new_n3354_ = new_n3352_ & new_n5138_;
  assign new_n3355_ = new_n3353_ | new_n5145_;
  assign new_n3356_ = new_n3351_ & new_n3349_;
  assign new_n3357_ = new_n3350_ | new_n3348_;
  assign new_n3358_ = new_n3356_ & new_n3355_;
  assign new_n3359_ = new_n3357_ | new_n3354_;
  assign new_n3360_ = new_n5153_ & new_n4969_;
  assign new_n3361_ = new_n5160_ | new_n4977_;
  assign new_n3362_ = new_n3360_ & new_n5164_;
  assign new_n3363_ = new_n3361_ | new_n5169_;
  assign new_n3364_ = new_n4956_ & new_n5227_;
  assign new_n3365_ = new_n4966_ | new_n5234_;
  assign new_n3366_ = new_n5238_ & new_n4975_;
  assign new_n3367_ = new_n5240_ | new_n4983_;
  assign new_n3368_ = new_n4987_ & new_n5183_;
  assign new_n3369_ = new_n4996_ | new_n5186_;
  assign new_n3370_ = new_n3367_ & new_n3365_;
  assign new_n3371_ = new_n3366_ | new_n3364_;
  assign new_n3372_ = new_n3370_ & new_n3369_;
  assign new_n3373_ = new_n3371_ | new_n3368_;
  assign new_n3374_ = new_n3373_ & new_n5153_;
  assign new_n3375_ = new_n3372_ | new_n5162_;
  assign new_n3376_ = new_n3363_ & new_n5188_;
  assign new_n3377_ = new_n3362_ | new_n5190_;
  assign new_n3378_ = new_n3376_ & new_n3375_;
  assign new_n3379_ = new_n3377_ | new_n3374_;
  assign new_n3380_ = new_n5243_ | new_n5198_;
  assign new_n3381_ = new_n3380_ | new_n5245_;
  assign new_n3382_ = new_n5243_ | new_n5204_;
  assign new_n3383_ = new_n3382_ | new_n5245_;
  assign new_n3384_ = new_n2281_ & new_n2233_;
  assign new_n3385_ = new_n2282_ | new_n2234_;
  assign new_n3386_ = new_n2288_ & new_n2228_;
  assign new_n3387_ = new_n2287_ | new_n2227_;
  assign new_n3388_ = new_n3387_ & new_n3385_;
  assign new_n3389_ = new_n3386_ | new_n3384_;
  assign new_n3390_ = new_n3388_ & new_n5024_;
  assign new_n3391_ = new_n3389_ | new_n5037_;
  assign new_n3392_ = new_n5054_ & new_n5172_;
  assign new_n3393_ = new_n5068_ | new_n5179_;
  assign new_n3394_ = new_n5075_ & new_n5033_;
  assign new_n3395_ = new_n5085_ | new_n5044_;
  assign new_n3396_ = new_n3393_ & new_n3391_;
  assign new_n3397_ = new_n3392_ | new_n3390_;
  assign new_n3398_ = new_n3396_ & new_n3395_;
  assign new_n3399_ = new_n3397_ | new_n3394_;
  assign new_n3400_ = new_n3399_ & new_n5105_;
  assign new_n3401_ = new_n3398_ | new_n5112_;
  assign new_n3402_ = new_n5120_ & new_n5234_;
  assign new_n3403_ = new_n5127_ | new_n5227_;
  assign new_n3404_ = new_n4913_ & new_n5099_;
  assign new_n3405_ = new_n4908_ | new_n5100_;
  assign new_n3406_ = new_n5247_ & new_n5228_;
  assign new_n3407_ = new_n5250_ | new_n5235_;
  assign new_n3408_ = new_n3406_ & new_n5139_;
  assign new_n3409_ = new_n3407_ | new_n5146_;
  assign new_n3410_ = new_n3403_ & new_n3401_;
  assign new_n3411_ = new_n3402_ | new_n3400_;
  assign new_n3412_ = new_n3410_ & new_n3409_;
  assign new_n3413_ = new_n3411_ | new_n3408_;
  assign new_n3414_ = new_n5047_ & new_n5235_;
  assign new_n3415_ = new_n5060_ | new_n5228_;
  assign new_n3416_ = new_n3414_ & new_n5180_;
  assign new_n3417_ = new_n3415_ | new_n5173_;
  assign new_n3418_ = new_n3417_ & new_n5024_;
  assign new_n3419_ = new_n3416_ | new_n5039_;
  assign new_n3420_ = new_n5054_ & new_n5236_;
  assign new_n3421_ = new_n5070_ | new_n5230_;
  assign new_n3422_ = new_n5075_ & new_n5212_;
  assign new_n3423_ = new_n5085_ | new_n5216_;
  assign new_n3424_ = new_n3421_ & new_n3419_;
  assign new_n3425_ = new_n3420_ | new_n3418_;
  assign new_n3426_ = new_n3424_ & new_n3423_;
  assign new_n3427_ = new_n3425_ | new_n3422_;
  assign new_n3428_ = new_n3427_ & new_n5105_;
  assign new_n3429_ = new_n3426_ | new_n5114_;
  assign new_n3430_ = new_n5120_ & new_n5048_;
  assign new_n3431_ = new_n5129_ | new_n5061_;
  assign new_n3432_ = new_n5247_ & new_n5061_;
  assign new_n3433_ = new_n5250_ | new_n5048_;
  assign new_n3434_ = new_n3432_ & new_n5139_;
  assign new_n3435_ = new_n3433_ | new_n5146_;
  assign new_n3436_ = new_n3431_ & new_n3429_;
  assign new_n3437_ = new_n3430_ | new_n3428_;
  assign new_n3438_ = new_n3436_ & new_n3435_;
  assign new_n3439_ = new_n3437_ | new_n3434_;
  assign new_n3440_ = new_n4928_ & new_n5252_;
  assign new_n3441_ = new_n3440_ & new_n5008_;
  assign new_n3442_ = new_n4956_ & new_n5253_;
  assign new_n3443_ = new_n5004_ & new_n4975_;
  assign new_n3444_ = new_n4989_ & new_n5018_;
  assign new_n3445_ = new_n3443_ | new_n3442_;
  assign new_n3446_ = new_n3445_ | new_n3444_;
  assign new_n3447_ = new_n3446_ & new_n4928_;
  assign new_n3448_ = new_n3441_ | new_n5015_;
  assign new_n3449_ = new_n3448_ | new_n3447_;
  assign new_n3450_ = new_n2279_ & new_n2231_;
  assign new_n3451_ = new_n2280_ | new_n2232_;
  assign new_n3452_ = new_n2286_ & new_n2226_;
  assign new_n3453_ = new_n2285_ | new_n2225_;
  assign new_n3454_ = new_n3453_ & new_n3451_;
  assign new_n3455_ = new_n3452_ | new_n3450_;
  assign new_n3456_ = new_n3454_ & new_n5026_;
  assign new_n3457_ = new_n3455_ | new_n5039_;
  assign new_n3458_ = new_n5056_ & new_n5212_;
  assign new_n3459_ = new_n5070_ | new_n5218_;
  assign new_n3460_ = new_n5077_ & new_n5254_;
  assign new_n3461_ = new_n5087_ | new_n1268_;
  assign new_n3462_ = new_n3459_ & new_n3457_;
  assign new_n3463_ = new_n3458_ | new_n3456_;
  assign new_n3464_ = new_n3462_ & new_n3461_;
  assign new_n3465_ = new_n3463_ | new_n3460_;
  assign new_n3466_ = new_n3465_ & new_n5107_;
  assign new_n3467_ = new_n3464_ | new_n5114_;
  assign new_n3468_ = new_n5122_ & new_n5080_;
  assign new_n3469_ = new_n5129_ | new_n5090_;
  assign new_n3470_ = new_n5133_ & new_n5091_;
  assign new_n3471_ = new_n5134_ | new_n5081_;
  assign new_n3472_ = new_n3470_ & new_n5141_;
  assign new_n3473_ = new_n3471_ | new_n5148_;
  assign new_n3474_ = new_n3469_ & new_n3467_;
  assign new_n3475_ = new_n3468_ | new_n3466_;
  assign new_n3476_ = new_n3474_ & new_n3473_;
  assign new_n3477_ = new_n3475_ | new_n3472_;
  assign new_n3478_ = new_n5155_ & new_n5184_;
  assign new_n3479_ = new_n5162_ | new_n5185_;
  assign new_n3480_ = new_n3478_ & new_n5166_;
  assign new_n3481_ = new_n3479_ | new_n5169_;
  assign new_n3482_ = new_n5063_ & new_n4957_;
  assign new_n3483_ = new_n5049_ | new_n4966_;
  assign new_n3484_ = new_n5255_ & new_n4976_;
  assign new_n3485_ = new_n2240_ | new_n4983_;
  assign new_n3486_ = new_n4989_ & new_n5238_;
  assign new_n3487_ = new_n4996_ | new_n5240_;
  assign new_n3488_ = new_n3485_ & new_n3483_;
  assign new_n3489_ = new_n3484_ | new_n3482_;
  assign new_n3490_ = new_n3488_ & new_n3487_;
  assign new_n3491_ = new_n3489_ | new_n3486_;
  assign new_n3492_ = new_n3491_ & new_n5155_;
  assign new_n3493_ = new_n3490_ | new_n5161_;
  assign new_n3494_ = new_n3481_ & new_n5187_;
  assign new_n3495_ = new_n3480_ | new_n5191_;
  assign new_n3496_ = new_n3494_ & new_n3493_;
  assign new_n3497_ = new_n3495_ | new_n3492_;
  assign new_n3498_ = new_n5258_ | new_n5199_;
  assign new_n3499_ = new_n3498_ | new_n5260_;
  assign new_n3500_ = new_n5258_ | new_n5205_;
  assign new_n3501_ = new_n3500_ | new_n5260_;
  assign new_n3502_ = new_n5261_ | new_n1278_;
  assign new_n3503_ = new_n5263_ | new_n1332_;
  assign new_n3504_ = new_n5026_ & new_n4948_;
  assign new_n3505_ = new_n5040_ | new_n4960_;
  assign new_n3506_ = new_n5056_ & new_n5012_;
  assign new_n3507_ = new_n5071_ | new_n5013_;
  assign new_n3508_ = new_n5077_ & new_n5236_;
  assign new_n3509_ = new_n5087_ | new_n5230_;
  assign new_n3510_ = new_n3507_ & new_n3505_;
  assign new_n3511_ = new_n3506_ | new_n3504_;
  assign new_n3512_ = new_n3510_ & new_n3509_;
  assign new_n3513_ = new_n3511_ | new_n3508_;
  assign new_n3514_ = new_n3513_ & new_n5107_;
  assign new_n3515_ = new_n3512_ | new_n5115_;
  assign new_n3516_ = new_n5122_ & new_n4959_;
  assign new_n3517_ = new_n5130_ | new_n4949_;
  assign new_n3518_ = new_n5248_ & new_n4949_;
  assign new_n3519_ = new_n5251_ | new_n4961_;
  assign new_n3520_ = new_n3518_ & new_n5141_;
  assign new_n3521_ = new_n3519_ | new_n5148_;
  assign new_n3522_ = new_n3517_ & new_n3515_;
  assign new_n3523_ = new_n3516_ | new_n3514_;
  assign new_n3524_ = new_n3522_ & new_n3521_;
  assign new_n3525_ = new_n3523_ | new_n3520_;
  assign new_n3526_ = new_n5264_ & new_n5265_;
  assign new_n3527_ = new_n5193_ & new_n5267_;
  assign new_n3528_ = new_n3527_ & new_n5269_;
  assign new_n3529_ = new_n5195_ & new_n5271_;
  assign new_n3530_ = new_n3529_ & new_n5269_;
  assign new_n3531_ = new_n3530_ | new_n3528_;
  assign new_n3532_ = new_n3531_ | new_n3299_;
  assign new_n3533_ = new_n3532_ & new_n3526_;
  assign new_n3534_ = new_n4856_ | new_n5273_;
  assign new_n3535_ = new_n3534_ | new_n4866_;
  assign new_n3536_ = new_n3535_ | new_n4880_;
  assign new_n3537_ = new_n5208_ | new_n5276_;
  assign new_n3538_ = new_n3537_ | new_n4841_;
  assign new_n3539_ = new_n5280_ | new_n5282_;
  assign new_n3540_ = new_n5285_ | new_n5287_;
  assign new_n3541_ = new_n5289_ & new_n5291_;
  assign new_n3542_ = new_n5285_ & new_n5287_;
  assign new_n3543_ = new_n5289_ | new_n5291_;
  assign new_n3544_ = new_n4894_ & new_n1727_;
  assign new_n3545_ = new_n4895_ | new_n1728_;
  assign new_n3546_ = new_n5292_ & new_n4686_;
  assign new_n3547_ = new_n5294_ | new_n4680_;
  assign new_n3548_ = new_n5294_ & new_n4681_;
  assign new_n3549_ = new_n5292_ | new_n4685_;
  assign new_n3550_ = new_n3549_ & new_n3547_;
  assign new_n3551_ = new_n3548_ | new_n3546_;
  assign new_n3552_ = new_n5296_ | new_n5299_;
  assign new_n3553_ = new_n3552_ | new_n5276_;
  assign new_n3554_ = new_n5299_ | new_n5277_;
  assign new_n3555_ = new_n5300_ | new_n5199_;
  assign new_n3556_ = new_n3555_ | new_n5303_;
  assign new_n3557_ = new_n5300_ | new_n5205_;
  assign new_n3558_ = new_n3557_ | new_n5303_;
  assign new_n3559_ = new_n5307_ | new_n5195_;
  assign new_n3560_ = new_n5309_ | new_n5277_;
  assign new_n3561_ = new_n4817_ & new_n4820_;
  assign new_n3562_ = new_n3561_ | new_n4822_;
  assign new_n3563_ = new_n1628_ & new_n5310_;
  assign new_n3564_ = new_n5311_ & new_n1626_;
  assign new_n3565_ = new_n3564_ | new_n3563_;
  assign new_n3566_ = new_n1676_ & new_n5312_;
  assign new_n3567_ = new_n5313_ & new_n1658_;
  assign new_n3568_ = new_n3567_ | new_n3566_;
  assign new_n3569_ = new_n5296_ & new_n3126_;
  assign new_n3570_ = new_n5315_ & new_n5316_;
  assign new_n3571_ = new_n3570_ | new_n3569_;
  assign new_n3572_ = new_n5282_ & new_n1530_;
  assign new_n3573_ = new_n1622_ & new_n5318_;
  assign new_n3574_ = new_n3573_ | new_n3572_;
  assign new_n3575_ = new_n1598_ & new_n5320_;
  assign new_n3576_ = new_n5323_ & new_n1536_;
  assign new_n3577_ = new_n3576_ | new_n3575_;
  assign new_n3578_ = new_n1737_ & new_n1729_;
  assign new_n3579_ = new_n1738_ | new_n1730_;
  assign new_n3580_ = new_n5325_ & new_n4688_;
  assign new_n3581_ = new_n5327_ | new_n4683_;
  assign new_n3582_ = new_n5327_ & new_n4684_;
  assign new_n3583_ = new_n5325_ | new_n4687_;
  assign new_n3584_ = new_n3583_ & new_n3581_;
  assign new_n3585_ = new_n3582_ | new_n3580_;
  assign new_n3586_ = new_n4670_ & new_n1943_;
  assign new_n3587_ = new_n4678_ | new_n1944_;
  assign new_n3588_ = new_n5315_ & new_n4823_;
  assign new_n3589_ = new_n5297_ | new_n4821_;
  assign new_n3590_ = new_n5314_ & new_n4815_;
  assign new_n3591_ = new_n5297_ | new_n4820_;
  assign new_n3592_ = new_n3590_ & new_n4814_;
  assign new_n3593_ = new_n3591_ | new_n4816_;
  assign new_n3594_ = new_n3589_ & new_n3587_;
  assign new_n3595_ = new_n3588_ | new_n3586_;
  assign new_n3596_ = new_n3594_ & new_n3593_;
  assign new_n3597_ = new_n3595_ | new_n3592_;
  assign new_n3598_ = new_n3596_ & new_n3585_;
  assign new_n3599_ = new_n3597_ & new_n3584_;
  assign new_n3600_ = new_n3599_ | new_n3598_;
  assign new_n3601_ = new_n4713_ & new_n5330_;
  assign new_n3602_ = new_n4716_ | new_n5333_;
  assign new_n3603_ = new_n4707_ & new_n5330_;
  assign new_n3604_ = new_n4708_ | new_n5333_;
  assign new_n3605_ = new_n5335_ | new_n4719_;
  assign new_n3606_ = new_n5336_ | new_n5338_;
  assign new_n3607_ = new_n5336_ | new_n5341_;
  assign new_n3608_ = new_n4718_ | new_n5332_;
  assign new_n3609_ = new_n5343_ & new_n3604_;
  assign new_n3610_ = new_n5344_ & new_n5338_;
  assign new_n3611_ = new_n5343_ | new_n5335_;
  assign new_n3612_ = new_n5345_ | new_n5341_;
  assign new_n3613_ = new_n5334_ | new_n4717_;
  assign new_n3614_ = new_n5346_ | new_n5342_;
  assign new_n3615_ = new_n5344_ & new_n5342_;
  assign new_n3616_ = new_n5345_ | new_n5339_;
  assign new_n3617_ = new_n5346_ | new_n5339_;
  assign new_n3618_ = new_n5347_ & new_n5348_;
  assign new_n3619_ = new_n5242_ & new_n5267_;
  assign new_n3620_ = new_n3619_ & new_n5349_;
  assign new_n3621_ = new_n5244_ & new_n5271_;
  assign new_n3622_ = new_n3621_ & new_n5349_;
  assign new_n3623_ = new_n3622_ | new_n3620_;
  assign new_n3624_ = new_n3623_ | new_n3359_;
  assign new_n3625_ = new_n3624_ & new_n3618_;
  assign new_n3626_ = new_n5351_ & new_n5353_;
  assign new_n3627_ = new_n3626_ | new_n5354_;
  assign new_n3628_ = new_n3627_ | new_n5357_;
  assign new_n3629_ = new_n3628_ | new_n5360_;
  assign new_n3630_ = new_n5273_ | new_n4879_;
  assign new_n3631_ = new_n5361_ | new_n4867_;
  assign new_n3632_ = new_n3631_ | new_n5279_;
  assign new_n3633_ = new_n5362_ | new_n5279_;
  assign new_n3634_ = new_n5361_ | new_n5278_;
  assign new_n3635_ = new_n4876_ & new_n4841_;
  assign new_n3636_ = new_n4881_ | new_n4884_;
  assign new_n3637_ = new_n3636_ & new_n4871_;
  assign new_n3638_ = new_n3635_ | new_n4874_;
  assign new_n3639_ = new_n3637_ & new_n4867_;
  assign new_n3640_ = new_n3638_ & new_n4862_;
  assign new_n3641_ = new_n3640_ | new_n3639_;
  assign new_n3642_ = new_n5307_ | new_n5244_;
  assign new_n3643_ = new_n5364_ & new_n5367_;
  assign new_n3644_ = new_n5370_ & new_n5372_;
  assign new_n3645_ = new_n5364_ | new_n5367_;
  assign new_n3646_ = new_n5370_ | new_n5372_;
  assign new_n3647_ = new_n5027_ & new_n5180_;
  assign new_n3648_ = new_n5040_ | new_n5173_;
  assign new_n3649_ = new_n5057_ & new_n4950_;
  assign new_n3650_ = new_n5071_ | new_n4961_;
  assign new_n3651_ = new_n5078_ & new_n5049_;
  assign new_n3652_ = new_n5086_ | new_n5063_;
  assign new_n3653_ = new_n3650_ & new_n3648_;
  assign new_n3654_ = new_n3649_ | new_n3647_;
  assign new_n3655_ = new_n3653_ & new_n3652_;
  assign new_n3656_ = new_n3654_ | new_n3651_;
  assign new_n3657_ = new_n3656_ & new_n5108_;
  assign new_n3658_ = new_n3655_ | new_n5115_;
  assign new_n3659_ = new_n5123_ & new_n5181_;
  assign new_n3660_ = new_n5130_ | new_n5175_;
  assign new_n3661_ = new_n5248_ & new_n5175_;
  assign new_n3662_ = new_n5251_ | new_n5181_;
  assign new_n3663_ = new_n3661_ & new_n5142_;
  assign new_n3664_ = new_n3662_ | new_n5147_;
  assign new_n3665_ = new_n3660_ & new_n3658_;
  assign new_n3666_ = new_n3659_ | new_n3657_;
  assign new_n3667_ = new_n3665_ & new_n3664_;
  assign new_n3668_ = new_n3666_ | new_n3663_;
  assign new_n3669_ = new_n5374_ & new_n5377_;
  assign new_n3670_ = new_n5380_ | new_n5200_;
  assign new_n3671_ = new_n3669_ & new_n5382_;
  assign new_n3672_ = new_n3670_ | new_n5385_;
  assign new_n3673_ = new_n5374_ & new_n5389_;
  assign new_n3674_ = new_n5380_ | new_n5206_;
  assign new_n3675_ = new_n3673_ & new_n5382_;
  assign new_n3676_ = new_n3674_ | new_n5385_;
  assign new_n3677_ = new_n3676_ & new_n3672_;
  assign new_n3678_ = new_n3675_ | new_n3671_;
  assign new_n3679_ = new_n5393_ & new_n5377_;
  assign new_n3680_ = new_n5396_ | new_n5200_;
  assign new_n3681_ = new_n3679_ & new_n5397_;
  assign new_n3682_ = new_n3680_ | new_n5400_;
  assign new_n3683_ = new_n5393_ & new_n5389_;
  assign new_n3684_ = new_n5396_ | new_n5206_;
  assign new_n3685_ = new_n3683_ & new_n5397_;
  assign new_n3686_ = new_n3684_ | new_n5400_;
  assign new_n3687_ = new_n3686_ & new_n3682_;
  assign new_n3688_ = new_n3685_ | new_n3681_;
  assign new_n3689_ = new_n5402_ | new_n5404_;
  assign new_n3690_ = new_n3689_ | new_n5329_;
  assign new_n3691_ = new_n5407_ | new_n5412_;
  assign new_n3692_ = new_n3691_ & new_n5416_;
  assign new_n3693_ = new_n5417_ & new_n4842_;
  assign new_n3694_ = new_n5418_ & new_n5419_;
  assign new_n3695_ = new_n3694_ & new_n5420_;
  assign new_n3696_ = new_n5421_ & new_n5422_;
  assign new_n3697_ = new_n4870_ & new_n4863_;
  assign new_n3698_ = new_n4873_ | new_n4868_;
  assign new_n3699_ = new_n4863_ & new_n4877_;
  assign new_n3700_ = new_n4868_ | new_n4881_;
  assign new_n3701_ = new_n3699_ & new_n4842_;
  assign new_n3702_ = new_n3700_ | new_n4883_;
  assign new_n3703_ = new_n3698_ & new_n4853_;
  assign new_n3704_ = new_n3697_ | new_n4850_;
  assign new_n3705_ = new_n3703_ & new_n3702_;
  assign new_n3706_ = new_n3704_ | new_n3701_;
  assign new_n3707_ = new_n3705_ & new_n4851_;
  assign new_n3708_ = new_n3706_ & new_n4856_;
  assign new_n3709_ = new_n3708_ | new_n3707_;
  assign new_n3710_ = new_n5425_ & new_n5353_;
  assign new_n3711_ = new_n5351_ | new_n5412_;
  assign new_n3712_ = new_n5350_ & new_n5413_;
  assign new_n3713_ = new_n5425_ | new_n5352_;
  assign new_n3714_ = new_n3713_ & new_n3711_;
  assign new_n3715_ = new_n3712_ | new_n3710_;
  assign new_n3716_ = new_n5357_ & new_n5407_;
  assign new_n3717_ = new_n5416_ | new_n5360_;
  assign new_n3718_ = new_n5415_ & new_n5359_;
  assign new_n3719_ = new_n5356_ | new_n5408_;
  assign new_n3720_ = new_n3719_ & new_n3717_;
  assign new_n3721_ = new_n3718_ | new_n3716_;
  assign new_n3722_ = new_n3721_ | new_n3714_;
  assign new_n3723_ = new_n3720_ | new_n3715_;
  assign new_n3724_ = new_n3723_ & new_n3722_;
  assign new_n3725_ = new_n5427_ & new_n4728_;
  assign new_n3726_ = new_n5429_ | new_n4724_;
  assign new_n3727_ = new_n5429_ & new_n4725_;
  assign new_n3728_ = new_n5427_ | new_n4727_;
  assign new_n3729_ = new_n3728_ & new_n3726_;
  assign new_n3730_ = new_n3727_ | new_n3725_;
  assign new_n3731_ = new_n3730_ & new_n5430_;
  assign new_n3732_ = new_n3729_ & new_n3173_;
  assign new_n3733_ = new_n3732_ | new_n3731_;
  assign new_n3734_ = new_n3137_ & new_n5431_;
  assign new_n3735_ = new_n5432_ & new_n3131_;
  assign new_n3736_ = new_n3735_ | new_n3734_;
  assign new_n3737_ = new_n5435_ & new_n5378_;
  assign new_n3738_ = new_n3737_ & new_n5437_;
  assign new_n3739_ = new_n5435_ & new_n5388_;
  assign new_n3740_ = new_n3739_ & new_n5437_;
  assign new_n3741_ = new_n3740_ | new_n3738_;
  assign new_n3742_ = new_n5434_ | new_n5439_;
  assign new_n3743_ = new_n3742_ | new_n5442_;
  assign new_n3744_ = new_n5436_ | new_n5444_;
  assign new_n3745_ = new_n3744_ | new_n5442_;
  assign new_n3746_ = new_n3745_ & new_n3743_;
  assign new_n3747_ = new_n3746_ & new_n3438_;
  assign new_n3748_ = new_n3747_ | new_n5446_;
  assign new_n3749_ = new_n5375_ | new_n5439_;
  assign new_n3750_ = new_n3749_ | new_n5384_;
  assign new_n3751_ = new_n5375_ | new_n5444_;
  assign new_n3752_ = new_n3751_ | new_n5386_;
  assign new_n3753_ = new_n3752_ & new_n3750_;
  assign new_n3754_ = new_n3753_ & new_n5381_;
  assign new_n3755_ = new_n3754_ | new_n5447_;
  assign new_n3756_ = new_n5448_ & new_n5449_;
  assign new_n3757_ = new_n5257_ & new_n5268_;
  assign new_n3758_ = new_n3757_ & new_n5450_;
  assign new_n3759_ = new_n5259_ & new_n5272_;
  assign new_n3760_ = new_n3759_ & new_n5450_;
  assign new_n3761_ = new_n3760_ | new_n3758_;
  assign new_n3762_ = new_n3761_ | new_n3477_;
  assign new_n3763_ = new_n3762_ & new_n3756_;
  assign new_n3764_ = new_n5392_ | new_n5440_;
  assign new_n3765_ = new_n3764_ | new_n5399_;
  assign new_n3766_ = new_n5394_ | new_n5445_;
  assign new_n3767_ = new_n3766_ | new_n5401_;
  assign new_n3768_ = new_n3767_ & new_n3765_;
  assign new_n3769_ = new_n3768_ & new_n5395_;
  assign new_n3770_ = new_n3769_ | new_n5451_;
  assign new_n3771_ = new_n5453_ | new_n5440_;
  assign new_n3772_ = new_n3771_ | new_n5302_;
  assign new_n3773_ = new_n5453_ | new_n5445_;
  assign new_n3774_ = new_n3773_ | new_n5304_;
  assign new_n3775_ = new_n5381_ | new_n5306_;
  assign new_n3776_ = new_n5263_ | new_n5259_;
  assign new_n3777_ = new_n5456_ & new_n5459_;
  assign new_n3778_ = new_n1227_ | new_n5459_;
  assign new_n3779_ = new_n5222_ | new_n5091_;
  assign new_n3780_ = new_n3779_ | new_n5218_;
  assign new_n3781_ = new_n3780_ & new_n5027_;
  assign new_n3782_ = new_n5057_ & new_n5081_;
  assign new_n3783_ = new_n5078_ & new_n5464_;
  assign new_n3784_ = new_n3782_ | new_n3781_;
  assign new_n3785_ = new_n3784_ | new_n3783_;
  assign new_n3786_ = new_n3785_ & new_n5108_;
  assign new_n3787_ = new_n5123_ & new_n5224_;
  assign new_n3788_ = new_n5133_ & new_n5221_;
  assign new_n3789_ = new_n3788_ & new_n5142_;
  assign new_n3790_ = new_n3787_ | new_n3786_;
  assign new_n3791_ = new_n3790_ | new_n3789_;
  assign new_n3792_ = new_n5466_ | new_n5468_;
  assign new_n3793_ = new_n3792_ | new_n3677_;
  assign new_n3794_ = new_n5468_ | new_n3687_;
  assign new_n3795_ = new_n5156_ & new_n5239_;
  assign new_n3796_ = new_n3795_ & new_n5166_;
  assign new_n3797_ = new_n5033_ & new_n4957_;
  assign new_n3798_ = new_n4976_ & new_n1281_;
  assign new_n3799_ = new_n4988_ & new_n5255_;
  assign new_n3800_ = new_n3798_ | new_n3797_;
  assign new_n3801_ = new_n3800_ | new_n3799_;
  assign new_n3802_ = new_n3801_ & new_n5156_;
  assign new_n3803_ = new_n3796_ | new_n5191_;
  assign new_n3804_ = new_n3803_ | new_n3802_;
  assign new_n3805_ = new_n5466_ | new_n5470_;
  assign new_n3806_ = new_n3805_ | new_n5472_;
  assign new_n3807_ = new_n3806_ | new_n5469_;
  assign new_n3808_ = new_n5473_ | new_n5456_;
  assign new_n3809_ = new_n5460_ & new_n1136_;
  assign new_n3810_ = new_n5475_ & new_n5460_;
  assign new_n3811_ = new_n5477_ & new_n5478_;
  assign G3519 = new_n2291_;
  assign G3520 = new_n2292_;
  assign G3521 = new_n2323_;
  assign G3522 = new_n2332_;
  assign G3523 = new_n2335_;
  assign G3524 = new_n2336_;
  assign G3525 = new_n2338_;
  assign G3526 = new_n2340_;
  assign G3527 = new_n2347_;
  assign G3528 = new_n2350_;
  assign G3529 = new_n2353_;
  assign G3530 = new_n2387_;
  assign G3531 = new_n2390_;
  assign G3532 = new_n2393_;
  assign G3533 = new_n2396_;
  assign G3534 = new_n1641_;
  assign G3535 = new_n1643_;
  assign G3536 = new_n2399_;
  assign G3537 = new_n4397_;
  assign G3538 = ~new_n2416_;
  assign G3539 = new_n2477_;
  assign G3540 = new_n2492_;
  assign n1836_li = new_n1393_;
  assign n1872_li = new_n4655_;
  assign n1884_li = new_n1395_;
  assign n1911_li = new_n1159_;
  assign n1914_li = new_n1237_;
  assign n1917_li = new_n1239_;
  assign n1923_li = new_n1161_;
  assign n1926_li = new_n1243_;
  assign n1929_li = new_n1245_;
  assign n1935_li = new_n1163_;
  assign n1938_li = new_n1249_;
  assign n1947_li = new_n1165_;
  assign n1950_li = new_n1253_;
  assign n1959_li = new_n1167_;
  assign n1962_li = new_n1257_;
  assign n1971_li = new_n1169_;
  assign n1974_li = new_n1261_;
  assign n1983_li = new_n1171_;
  assign n1995_li = new_n1173_;
  assign n2007_li = new_n1175_;
  assign n2019_li = new_n1177_;
  assign n2031_li = new_n1179_;
  assign n2043_li = new_n1181_;
  assign n2055_li = new_n1183_;
  assign n2064_li = new_n4888_;
  assign n2067_li = new_n1185_;
  assign n2100_li = new_n1431_;
  assign n2112_li = new_n1427_;
  assign n2124_li = new_n1429_;
  assign n2136_li = new_n1437_;
  assign n2148_li = new_n1439_;
  assign n2160_li = new_n1441_;
  assign n2163_li = new_n1201_;
  assign n2172_li = new_n1453_;
  assign n2175_li = new_n1203_;
  assign n2184_li = new_n1463_;
  assign n2223_li = new_n1211_;
  assign n2235_li = new_n1213_;
  assign n2238_li = new_n1305_;
  assign n2247_li = new_n1215_;
  assign n2250_li = new_n1309_;
  assign n2259_li = new_n1217_;
  assign n2262_li = new_n1313_;
  assign n2271_li = new_n1219_;
  assign n2274_li = new_n1317_;
  assign n2283_li = new_n1221_;
  assign n2286_li = new_n1321_;
  assign n2295_li = new_n1223_;
  assign n2298_li = new_n1325_;
  assign n2304_li = new_n4606_;
  assign n2307_li = new_n1225_;
  assign n2331_li = new_n1229_;
  assign n2334_li = new_n1333_;
  assign n2337_li = new_n1335_;
  assign n2340_li = new_n1337_;
  assign n3241_i2 = new_n1399_;
  assign n3242_i2 = new_n1401_;
  assign n3610_i2 = new_n1447_;
  assign n3980_i2 = new_n1471_;
  assign n3968_i2 = new_n1465_;
  assign n4298_i2 = new_n1491_;
  assign n4371_i2 = new_n1531_;
  assign n4413_i2 = new_n1561_;
  assign n4418_i2 = new_n1565_;
  assign n4628_i2 = new_n1647_;
  assign n4629_i2 = new_n1649_;
  assign n4633_i2 = new_n1651_;
  assign n4634_i2 = new_n1653_;
  assign n4732_i2 = new_n1663_;
  assign n4733_i2 = new_n1665_;
  assign n4884_i2 = new_n1705_;
  assign n4886_i2 = new_n1707_;
  assign n4890_i2 = new_n1711_;
  assign n5011_i2 = new_n4447_;
  assign n5012_i2 = new_n4446_;
  assign n5013_i2 = new_n4449_;
  assign n5014_i2 = new_n4489_;
  assign n5015_i2 = new_n1755_;
  assign n5021_i2 = new_n1761_;
  assign n5016_i2 = new_n1757_;
  assign n5026_i2 = new_n1763_;
  assign n4377_i2 = new_n5408_;
  assign n4378_i2 = new_n5320_;
  assign n4389_i2 = new_n1539_;
  assign n4390_i2 = new_n1541_;
  assign n4391_i2 = new_n1543_;
  assign n4398_i2 = new_n5404_;
  assign n4401_i2 = new_n5481_;
  assign n5117_i2 = new_n4484_;
  assign n5115_i2 = new_n4614_;
  assign n5122_i2 = new_n4526_;
  assign n5121_i2 = new_n4531_;
  assign n5119_i2 = new_n4536_;
  assign n5116_i2 = new_n4542_;
  assign n5123_i2 = new_n4547_;
  assign n5156_i2 = new_n4653_;
  assign n5167_i2 = new_n1965_;
  assign n4454_i2 = new_n5323_;
  assign n4455_i2 = new_n4828_;
  assign n4456_i2 = new_n4831_;
  assign n4505_i2 = new_n4824_;
  assign G742_i2 = new_n4457_;
  assign G727_i2 = new_n4654_;
  assign n4567_i2 = new_n4833_;
  assign n4568_i2 = new_n5310_;
  assign n4569_i2 = new_n5311_;
  assign n4571_i2 = new_n1629_;
  assign n4572_i2 = new_n1631_;
  assign n4537_i2 = new_n1609_;
  assign n4539_i2 = new_n1613_;
  assign n4651_i2 = new_n1655_;
  assign n4652_i2 = new_n5312_;
  assign n4653_i2 = new_n1659_;
  assign G1514_i2 = new_n4624_;
  assign G1823_i2 = ~new_n4648_;
  assign n4783_i2 = new_n4702_;
  assign n4787_i2 = new_n5313_;
  assign n4808_i2 = new_n1677_;
  assign n4815_i2 = new_n1679_;
  assign n4816_i2 = new_n1681_;
  assign n4822_i2 = new_n1683_;
  assign G572_i2 = new_n4459_;
  assign n4919_i2 = new_n1721_;
  assign n4920_i2 = new_n4660_;
  assign n4921_i2 = new_n4662_;
  assign G1048_i2 = new_n4593_;
  assign n5041_i2 = new_n1789_;
  assign n5094_i2 = new_n1853_;
  assign n5278_i2 = new_n4848_;
  assign n5301_i2 = new_n4846_;
  assign G2610_i2 = new_n4671_;
  assign G3174_i2 = new_n4732_;
  assign G3146_i2 = ~new_n4735_;
  assign G3217_i2 = ~new_n4738_;
  assign G3220_i2 = ~new_n4741_;
  assign G2839_i2 = ~new_n4739_;
  assign G3251_i2 = ~new_n4740_;
  assign G3042_i2 = new_n4783_;
  assign G3045_i2 = ~new_n4782_;
  assign G3262_i2 = new_n4731_;
  assign G2845_i2 = ~new_n4742_;
  assign G2929_i2 = new_n4733_;
  assign G2848_i2 = ~new_n4736_;
  assign G2851_i2 = new_n4784_;
  assign G3291_i2 = ~new_n4737_;
  assign G3254_i2 = ~new_n4734_;
  assign G2666_i2 = new_n4885_;
  assign n5099_i2 = new_n5098_;
  assign n5100_i2 = new_n5219_;
  assign n5101_i2 = new_n5176_;
  assign G2558_i2 = new_n4795_;
  assign n5266_i2 = new_n5092_;
  assign n5267_i2 = new_n5231_;
  assign G2759_i2 = new_n4877_;
  assign n5269_i2 = new_n2167_;
  assign n5270_i2 = new_n2169_;
  assign n5271_i2 = new_n2171_;
  assign n5292_i2 = new_n4908_;
  assign n5293_i2 = new_n4901_;
  assign n5294_i2 = new_n5096_;
  assign n5295_i2 = new_n4919_;
  assign G618_i2 = new_n4887_;
  assign G621_i2 = new_n4886_;
  assign G384_i2 = new_n5413_;
  assign G377_i2 = new_n5409_;
  assign G400_i2 = new_n5424_;
  assign G3171_i2 = ~new_n4797_;
  assign G2552_i2 = ~new_n4836_;
  assign G3272_i2 = ~new_n4800_;
  assign G2015_i2 = new_n5428_;
  assign G3294_i2 = new_n5286_;
  assign G3281_i2 = ~new_n5290_;
  assign G3320_i2 = ~new_n5484_;
  assign G3275_i2 = ~new_n5284_;
  assign G3140_i2 = ~new_n4803_;
  assign G2836_i2 = ~new_n4801_;
  assign G2926_i2 = ~new_n4798_;
  assign G2842_i2 = ~new_n4804_;
  assign G3302_i2 = ~new_n4799_;
  assign G3288_i2 = ~new_n4796_;
  assign G3143_i2 = ~new_n4802_;
  assign G3100_i2 = ~new_n5288_;
  assign G2512_i2 = new_n4725_;
  assign n5325_i2 = new_n5064_;
  assign n5326_i2 = new_n5184_;
  assign n5327_i2 = new_n4969_;
  assign n1857_lo_buf_i2 = new_n5032_;
  assign n2097_lo_buf_i2 = new_n5239_;
  assign G2669_i2 = new_n5207_;
  assign G552_i2 = n5100_i2;
  assign G568_i2 = n5101_i2;
  assign G530_i2 = new_n5001_;
  assign G565_i2 = n5267_i2;
  assign G559_i2 = n5325_i2;
  assign n1821_lo_buf_i2 = new_n5223_;
  assign n1905_lo_buf_i2 = new_n4950_;
  assign n2133_lo_buf_i2 = new_n4992_;
  assign n2145_lo_buf_i2 = new_n4931_;
  assign n2157_lo_buf_i2 = new_n5004_;
  assign n2205_lo_buf_i2 = new_n5011_;
  assign n2217_lo_buf_i2 = new_n5019_;
  assign G447_i2 = new_n5318_;
  assign G434_i2 = new_n5321_;
  assign G422_i2 = new_n5324_;
  assign G461_i2 = new_n5283_;
  assign G3312_i2 = ~new_n4891_;
  assign G3332_i2 = ~new_n4893_;
  assign G3195_i2 = ~new_n5487_;
  assign G2607_i2 = new_n4843_;
  assign G2799_i2 = new_n5316_;
  assign G1005_i2 = new_n5431_;
  assign G1008_i2 = new_n5432_;
  assign n2001_lo_buf_i2 = new_n5254_;
  assign n2169_lo_buf_i2 = new_n5017_;
  assign n2229_lo_buf_i2 = new_n5253_;
  assign n2301_lo_buf_i2 = new_n5419_;
  assign G2816_i2 = ~new_n5420_;
  assign G2947_i2 = new_n5430_;
  assign n2013_lo_buf_i2 = new_n5378_;
  assign n2025_lo_buf_i2 = new_n5390_;
  assign n2037_lo_buf_i2 = new_n5268_;
  assign n2049_lo_buf_i2 = new_n5272_;
  assign n2181_lo_buf_i2 = new_n5252_;
  assign G546_i2 = n5266_i2;
  assign G480_i2 = n5293_i2;
  assign G492_i2 = n5294_i2;
  assign G540_i2 = n1821_lo_buf_i2;
  assign G3350_i2 = ~new_n5489_;
  assign G3360_i2 = ~new_n5490_;
  assign G3373_i2 = G3320_i2;
  assign G3237_i2 = G3195_i2;
  assign G2773_i2 = new_n5309_;
  assign G1733_i2 = new_n5441_;
  assign G1738_i2 = new_n5401_;
  assign G1751_i2 = new_n5386_;
  assign G2216_i2 = ~new_n5265_;
  assign G2219_i2 = ~new_n5264_;
  assign G381_i2 = new_n5414_;
  assign G397_i2 = new_n5426_;
  assign G787_i2 = new_n5280_;
  assign G2823_i2 = ~new_n5298_;
  assign G2796_i2 = new_n5418_;
  assign G875_i2 = new_n5261_;
  assign G2208_i2 = ~new_n5348_;
  assign G2211_i2 = ~new_n5347_;
  assign n1989_lo_buf_i2 = new_n5464_;
  assign n2061_lo_buf_i2 = new_n1277_;
  assign n2313_lo_buf_i2 = new_n1331_;
  assign G2232_i2 = new_n5394_;
  assign G1725_i2 = new_n5436_;
  assign G1764_i2 = new_n5304_;
  assign G2356_i2 = ~new_n5449_;
  assign G2359_i2 = ~new_n5448_;
  assign G1180_i2 = ~new_n5308_;
  assign G1756_i2 = new_n5454_;
  assign G2441_i2 = new_n5492_;
  assign G2887_i2 = new_n1713_;
  assign G2991_i2 = new_n1759_;
  assign G470_i2 = new_n5403_;
  assign G484_i2 = new_n5402_;
  assign G496_i2 = new_n5331_;
  assign G353_i2 = new_n5358_;
  assign G363_i2 = G353_i2;
  assign G2805_i2 = G2666_i2;
  assign G2906_i2 = ~new_n5362_;
  assign G2833_i2 = ~new_n5417_;
  assign G1012_i2 = new_n5354_;
  assign G3353_i2 = ~new_n4890_;
  assign G3367_i2 = ~new_n4892_;
  assign G3346_i2 = ~new_n3540_;
  assign G3340_i2 = ~new_n3541_;
  assign G3376_i2 = ~new_n5485_;
  assign G3359_i2 = new_n3542_;
  assign G3240_i2 = ~new_n5488_;
  assign G3344_i2 = ~new_n3543_;
  assign G2880_i2 = ~new_n5494_;
  assign G2939_i2 = ~new_n5495_;
  assign G2248_i2 = ~new_n5422_;
  assign G2251_i2 = ~new_n5421_;
  assign G2021_i2 = ~new_n5497_;
  assign G3383_i2 = G3350_i2;
  assign G3399_i2 = G3360_i2;
  assign G3404_i2 = G3376_i2;
  assign G3265_i2 = G3240_i2;
  assign G2866_i2 = ~new_n5368_;
  assign G2999_i2 = ~new_n5365_;
  assign G736_i2 = n4401_i2;
  assign G739_i2 = new_n5480_;
  assign G1200_i2 = new_n5498_;
  assign G1203_i2 = new_n5499_;
  assign G3027_i2 = new_n5500_;
  assign G1463_i2 = new_n5501_;
  assign G1460_i2 = new_n5502_;
  assign G3012_i2 = new_n5503_;
  assign G1574_i2 = ~new_n5507_;
  assign G1646_i2 = G1574_i2;
  assign G1592_i2 = ~new_n5518_;
  assign G1664_i2 = G1592_i2;
  assign G1547_i2 = ~new_n5529_;
  assign G1619_i2 = G1547_i2;
  assign G1556_i2 = ~new_n5540_;
  assign G1628_i2 = G1556_i2;
  assign G1583_i2 = new_n5551_;
  assign G1655_i2 = G1583_i2;
  assign G1529_i2 = new_n5562_;
  assign G1601_i2 = G1529_i2;
  assign G1538_i2 = ~new_n5573_;
  assign G1610_i2 = G1538_i2;
  assign G1565_i2 = ~new_n5584_;
  assign G1637_i2 = G1565_i2;
  assign G2437_i2 = new_n5593_;
  assign G2518_i2 = G2441_i2;
  assign n1785_lo_buf_i2 = new_n5462_;
  assign n1845_lo_buf_i2 = new_n5595_;
  assign n1893_lo_buf_i2 = new_n5598_;
  assign n1941_lo_buf_i2 = new_n1251_;
  assign n1953_lo_buf_i2 = new_n1255_;
  assign n1965_lo_buf_i2 = new_n1259_;
  assign n1977_lo_buf_i2 = new_n1263_;
  assign n2241_lo_buf_i2 = new_n1307_;
  assign n2253_lo_buf_i2 = new_n1311_;
  assign n2265_lo_buf_i2 = new_n1315_;
  assign n2277_lo_buf_i2 = new_n1319_;
  assign n2289_lo_buf_i2 = new_n1323_;
  assign G519_i2 = new_n1525_;
  assign G388_i2 = G381_i2;
  assign G438_i2 = new_n5317_;
  assign G368_i2 = G377_i2;
  assign G1318_i2 = ~new_n3629_;
  assign G425_i2 = G434_i2;
  assign G593_i2 = G496_i2;
  assign G413_i2 = G422_i2;
  assign G404_i2 = G397_i2;
  assign G451_i2 = G461_i2;
  assign G2284_i2 = new_n1927_;
  assign G2580_i2 = new_n2157_;
  assign G2302_i2 = new_n4812_;
  assign G2598_i2 = new_n4810_;
  assign G2497_i2 = new_n5293_;
  assign G2651_i2 = new_n4681_;
  assign G2296_i2 = new_n5326_;
  assign G2308_i2 = new_n4897_;
  assign G2592_i2 = new_n4684_;
  assign G2604_i2 = new_n4691_;
  assign G2902_i2 = ~new_n3632_;
  assign G2975_i2 = ~new_n3633_;
  assign G2962_i2 = ~new_n5371_;
  assign G3069_i2 = ~new_n5369_;
  assign G2018_i2 = ~new_n5600_;
  assign G1176_i2 = ~new_n5262_;
  assign G1189_i2 = G1180_i2;
  assign G3066_i2 = ~new_n3643_;
  assign G3137_i2 = ~new_n3644_;
  assign G3038_i2 = ~new_n3645_;
  assign G3117_i2 = ~new_n3646_;
  assign G2384_i2 = new_n5447_;
  assign G2472_i2 = new_n5451_;
  assign G772_i2 = new_n3690_;
  assign G935_i2 = new_n3692_;
  assign G2923_i2 = ~new_n3693_;
  assign G2971_i2 = G2880_i2;
  assign G2980_i2 = G2939_i2;
  assign G3039_i2 = new_n3695_;
  assign G2388_i2 = ~new_n5470_;
  assign G2287_i2 = G2021_i2;
  assign G3024_i2 = new_n3709_;
  assign G2916_i2 = G2866_i2;
  assign G1819_i2 = new_n3724_;
  assign G3035_i2 = G2999_i2;
  assign G3107_i2 = new_n3733_;
  assign G1023_i2 = new_n5482_;
  assign G1024_i2 = G1023_i2;
  assign G1311_i2 = G1200_i2;
  assign G1312_i2 = G1203_i2;
  assign G3063_i2 = G3027_i2;
  assign G1520_i2 = G1463_i2;
  assign G1519_i2 = G1460_i2;
  assign G3078_i2 = G3012_i2;
  assign G2038_i2 = new_n3736_;
  assign G1848_i2 = ~new_n5508_;
  assign G1864_i2 = G1848_i2;
  assign G1872_i2 = ~new_n5510_;
  assign G1880_i2 = G1872_i2;
  assign G1888_i2 = ~new_n5511_;
  assign G1912_i2 = G1888_i2;
  assign G1928_i2 = ~new_n5513_;
  assign G1936_i2 = G1928_i2;
  assign G1944_i2 = ~new_n5514_;
  assign G1952_i2 = G1944_i2;
  assign G1850_i2 = ~new_n5519_;
  assign G1866_i2 = G1850_i2;
  assign G1874_i2 = ~new_n5521_;
  assign G1882_i2 = G1874_i2;
  assign G1890_i2 = ~new_n5522_;
  assign G1914_i2 = G1890_i2;
  assign G1930_i2 = ~new_n5524_;
  assign G1938_i2 = G1930_i2;
  assign G1946_i2 = ~new_n5525_;
  assign G1954_i2 = G1946_i2;
  assign G1845_i2 = ~new_n5530_;
  assign G1861_i2 = G1845_i2;
  assign G1869_i2 = ~new_n5532_;
  assign G1877_i2 = G1869_i2;
  assign G1885_i2 = ~new_n5533_;
  assign G1909_i2 = G1885_i2;
  assign G1925_i2 = ~new_n5535_;
  assign G1933_i2 = G1925_i2;
  assign G1941_i2 = ~new_n5536_;
  assign G1949_i2 = G1941_i2;
  assign G1846_i2 = ~new_n5541_;
  assign G1862_i2 = G1846_i2;
  assign G1870_i2 = ~new_n5543_;
  assign G1878_i2 = G1870_i2;
  assign G1886_i2 = ~new_n5544_;
  assign G1910_i2 = G1886_i2;
  assign G1926_i2 = ~new_n5546_;
  assign G1934_i2 = G1926_i2;
  assign G1942_i2 = ~new_n5547_;
  assign G1950_i2 = G1942_i2;
  assign G1849_i2 = new_n5552_;
  assign G1865_i2 = G1849_i2;
  assign G1873_i2 = new_n5554_;
  assign G1881_i2 = G1873_i2;
  assign G1889_i2 = new_n5555_;
  assign G1913_i2 = G1889_i2;
  assign G1929_i2 = new_n5557_;
  assign G1937_i2 = G1929_i2;
  assign G1945_i2 = new_n5558_;
  assign G1953_i2 = G1945_i2;
  assign G1843_i2 = new_n5563_;
  assign G1859_i2 = G1843_i2;
  assign G1867_i2 = new_n5565_;
  assign G1875_i2 = G1867_i2;
  assign G1883_i2 = new_n5566_;
  assign G1907_i2 = G1883_i2;
  assign G1923_i2 = new_n5568_;
  assign G1931_i2 = G1923_i2;
  assign G1939_i2 = new_n5569_;
  assign G1947_i2 = G1939_i2;
  assign G1844_i2 = ~new_n5574_;
  assign G1860_i2 = G1844_i2;
  assign G1868_i2 = ~new_n5576_;
  assign G1876_i2 = G1868_i2;
  assign G1884_i2 = ~new_n5577_;
  assign G1908_i2 = G1884_i2;
  assign G1924_i2 = ~new_n5579_;
  assign G1932_i2 = G1924_i2;
  assign G1940_i2 = ~new_n5580_;
  assign G1948_i2 = G1940_i2;
  assign G1847_i2 = ~new_n5585_;
  assign G1863_i2 = G1847_i2;
  assign G1871_i2 = ~new_n5587_;
  assign G1879_i2 = G1871_i2;
  assign G1887_i2 = ~new_n5588_;
  assign G1911_i2 = G1887_i2;
  assign G1927_i2 = ~new_n5590_;
  assign G1935_i2 = G1927_i2;
  assign G1943_i2 = ~new_n5591_;
  assign G1951_i2 = G1943_i2;
  assign G2444_i2 = ~new_n5469_;
  assign G2451_i2 = ~new_n5472_;
  assign G2502_i2 = new_n5601_;
  assign G2507_i2 = ~new_n5465_;
  assign G2515_i2 = G2437_i2;
  assign G2583_i2 = new_n5493_;
  assign n1797_lo_buf_i2 = new_n5455_;
  assign n1833_lo_buf_i2 = new_n5603_;
  assign n1881_lo_buf_i2 = new_n5605_;
  assign G523_i2 = n1785_lo_buf_i2;
  assign G575_i2 = n1845_lo_buf_i2;
  assign G578_i2 = n1893_lo_buf_i2;
  assign G615_i2 = n2025_lo_buf_i2;
  assign G2254_i2 = ~new_n3772_;
  assign G2255_i2 = ~new_n3774_;
  assign G2027_i2 = ~new_n3775_;
  assign G2393_i2 = ~new_n3776_;
  assign G527_i2 = new_n5606_;
  assign G594_i2 = new_n5475_;
  assign G1689_i2 = new_n5607_;
  assign G1693_i2 = G1689_i2;
  assign G2281_i2 = G2018_i2;
  assign G2014_i2 = G1756_i2;
  assign G2459_i2 = new_n5446_;
  assign G2561_i2 = ~new_n3793_;
  assign G2533_i2 = ~new_n3794_;
  assign n1749_lo_buf_i2 = new_n5608_;
  assign n1761_lo_buf_i2 = new_n5478_;
  assign n1773_lo_buf_i2 = new_n5477_;
  assign n1809_lo_buf_i2 = new_n5473_;
  assign G1955_i2 = new_n5609_;
  assign G1958_i2 = G1955_i2;
  assign G2562_i2 = ~new_n3807_;
  assign G2398_i2 = ~new_n5496_;
  assign G2524_i2 = ~new_n5471_;
  assign G2563_i2 = G2502_i2;
  assign G2577_i2 = new_n5592_;
  assign G2627_i2 = G2583_i2;
  assign G654_i2 = n1833_lo_buf_i2;
  assign G660_i2 = n1881_lo_buf_i2;
  assign G831_i2 = new_n5463_;
  assign G919_i2 = new_n5596_;
  assign G925_i2 = new_n5599_;
  assign n1815_lo_buf_i2 = new_n1143_;
  assign n1899_lo_buf_i2 = new_n1157_;
  assign n2079_lo_buf_i2 = new_n1187_;
  assign n2127_lo_buf_i2 = new_n1195_;
  assign n2139_lo_buf_i2 = new_n1197_;
  assign n2151_lo_buf_i2 = new_n1199_;
  assign n2187_lo_buf_i2 = new_n1205_;
  assign n2199_lo_buf_i2 = new_n1207_;
  assign n2211_lo_buf_i2 = new_n1209_;
  assign G533_i2 = new_n3808_;
  assign n1854_lo_buf_i2 = new_n1149_;
  assign n2094_lo_buf_i2 = new_n1189_;
  assign G667_i2 = new_n3809_;
  assign G874_i2 = G527_i2;
  assign G851_i2 = new_n5474_;
  assign G1127_i2 = new_n3810_;
  assign n1869_lo_buf_i2 = new_n1151_;
  assign n2109_lo_buf_i2 = new_n1191_;
  assign n2121_lo_buf_i2 = new_n1193_;
  assign G477_i2 = n1749_lo_buf_i2;
  assign G491_i2 = new_n3811_;
  assign G501_i2 = new_n5476_;
  assign G786_i2 = new_n5602_;
  assign G791_i2 = new_n5604_;
  assign G1126_i2 = G831_i2;
  assign G1052_i2 = G919_i2;
  assign G1054_i2 = G925_i2;
  assign new_n4363_ = new_n1378_;
  assign new_n4364_ = new_n1377_;
  assign new_n4365_ = new_n1382_;
  assign new_n4366_ = new_n1381_;
  assign new_n4367_ = new_n2296_;
  assign new_n4368_ = new_n1298_;
  assign new_n4369_ = new_n1294_;
  assign new_n4370_ = new_n1292_;
  assign new_n4371_ = new_n2300_;
  assign new_n4372_ = new_n2301_;
  assign new_n4373_ = new_n2295_;
  assign new_n4374_ = new_n1366_;
  assign new_n4375_ = new_n1363_;
  assign new_n4376_ = new_n1365_;
  assign new_n4377_ = new_n1364_;
  assign new_n4378_ = new_n1357_;
  assign new_n4379_ = new_n1329_;
  assign new_n4380_ = new_n2349_;
  assign new_n4381_ = new_n2352_;
  assign new_n4382_ = new_n1746_;
  assign new_n4383_ = new_n1743_;
  assign new_n4384_ = new_n1745_;
  assign new_n4385_ = new_n1744_;
  assign new_n4386_ = new_n1369_;
  assign new_n4387_ = new_n1367_;
  assign new_n4388_ = new_n1370_;
  assign new_n4389_ = new_n1368_;
  assign new_n4390_ = new_n2389_;
  assign new_n4391_ = new_n2392_;
  assign new_n4392_ = new_n2395_;
  assign new_n4393_ = new_n2398_;
  assign new_n4394_ = new_n2404_;
  assign new_n4395_ = new_n2406_;
  assign new_n4396_ = new_n2412_;
  assign new_n4397_ = new_n2410_;
  assign new_n4398_ = new_n2420_;
  assign new_n4399_ = new_n2417_;
  assign new_n4400_ = new_n2419_;
  assign new_n4401_ = new_n2418_;
  assign new_n4402_ = new_n1687_;
  assign new_n4403_ = new_n1686_;
  assign new_n4404_ = new_n1688_;
  assign new_n4405_ = new_n1685_;
  assign new_n4406_ = new_n2438_;
  assign new_n4407_ = new_n2432_;
  assign new_n4408_ = new_n4407_;
  assign new_n4409_ = new_n4407_;
  assign new_n4410_ = new_n2437_;
  assign new_n4411_ = new_n2431_;
  assign new_n4412_ = new_n4411_;
  assign new_n4413_ = new_n4411_;
  assign new_n4414_ = new_n2439_;
  assign new_n4415_ = new_n4414_;
  assign new_n4416_ = new_n4414_;
  assign new_n4417_ = new_n2440_;
  assign new_n4418_ = new_n4417_;
  assign new_n4419_ = new_n4417_;
  assign new_n4420_ = new_n1793_;
  assign new_n4421_ = new_n1792_;
  assign new_n4422_ = new_n1794_;
  assign new_n4423_ = new_n1791_;
  assign new_n4424_ = new_n2449_;
  assign new_n4425_ = new_n2450_;
  assign new_n4426_ = new_n1777_;
  assign new_n4427_ = new_n1773_;
  assign new_n4428_ = new_n1778_;
  assign new_n4429_ = new_n1774_;
  assign new_n4430_ = new_n2459_;
  assign new_n4431_ = new_n2460_;
  assign new_n4432_ = new_n2426_;
  assign new_n4433_ = new_n2425_;
  assign new_n4434_ = new_n1768_;
  assign new_n4435_ = new_n1765_;
  assign new_n4436_ = new_n1767_;
  assign new_n4437_ = new_n1766_;
  assign new_n4438_ = new_n2483_;
  assign new_n4439_ = new_n2482_;
  assign new_n4440_ = new_n1635_;
  assign new_n4441_ = new_n1750_;
  assign new_n4442_ = new_n4441_;
  assign new_n4443_ = new_n1748_;
  assign new_n4444_ = new_n1749_;
  assign new_n4445_ = new_n4444_;
  assign new_n4446_ = new_n4444_;
  assign new_n4447_ = new_n1747_;
  assign new_n4448_ = new_n4447_;
  assign new_n4449_ = new_n1751_;
  assign new_n4450_ = new_n1449_;
  assign new_n4451_ = new_n4450_;
  assign new_n4452_ = new_n1450_;
  assign new_n4453_ = new_n4452_;
  assign new_n4454_ = new_n1470_;
  assign new_n4455_ = new_n1468_;
  assign new_n4456_ = new_n1469_;
  assign new_n4457_ = new_n1467_;
  assign new_n4458_ = new_n4457_;
  assign new_n4459_ = new_n1403_;
  assign new_n4460_ = new_n2523_;
  assign new_n4461_ = new_n4460_;
  assign new_n4462_ = new_n2517_;
  assign new_n4463_ = new_n2529_;
  assign new_n4464_ = new_n4463_;
  assign new_n4465_ = new_n2522_;
  assign new_n4466_ = new_n4465_;
  assign new_n4467_ = new_n4466_;
  assign new_n4468_ = new_n4466_;
  assign new_n4469_ = new_n4465_;
  assign new_n4470_ = new_n4469_;
  assign new_n4471_ = new_n1926_;
  assign new_n4472_ = new_n1924_;
  assign new_n4473_ = new_n1925_;
  assign new_n4474_ = new_n1923_;
  assign new_n4475_ = new_n2536_;
  assign new_n4476_ = new_n4475_;
  assign new_n4477_ = new_n2541_;
  assign new_n4478_ = new_n1862_;
  assign new_n4479_ = new_n4478_;
  assign new_n4480_ = new_n1885_;
  assign new_n4481_ = new_n4480_;
  assign new_n4482_ = new_n4481_;
  assign new_n4483_ = new_n4481_;
  assign new_n4484_ = new_n4480_;
  assign new_n4485_ = new_n1753_;
  assign new_n4486_ = new_n4485_;
  assign new_n4487_ = new_n4486_;
  assign new_n4488_ = new_n4486_;
  assign new_n4489_ = new_n4485_;
  assign new_n4490_ = new_n1452_;
  assign new_n4491_ = new_n4490_;
  assign new_n4492_ = new_n4491_;
  assign new_n4493_ = new_n4491_;
  assign new_n4494_ = new_n4490_;
  assign new_n4495_ = new_n1476_;
  assign new_n4496_ = new_n4495_;
  assign new_n4497_ = new_n4496_;
  assign new_n4498_ = new_n4496_;
  assign new_n4499_ = new_n4495_;
  assign new_n4500_ = new_n1868_;
  assign new_n4501_ = new_n4500_;
  assign new_n4502_ = new_n4501_;
  assign new_n4503_ = new_n4500_;
  assign new_n4504_ = new_n1866_;
  assign new_n4505_ = new_n4504_;
  assign new_n4506_ = new_n4505_;
  assign new_n4507_ = new_n4504_;
  assign new_n4508_ = new_n1864_;
  assign new_n4509_ = new_n4508_;
  assign new_n4510_ = new_n4508_;
  assign new_n4511_ = new_n1880_;
  assign new_n4512_ = new_n4511_;
  assign new_n4513_ = new_n4512_;
  assign new_n4514_ = new_n4513_;
  assign new_n4515_ = new_n4512_;
  assign new_n4516_ = new_n4511_;
  assign new_n4517_ = new_n4516_;
  assign new_n4518_ = new_n4516_;
  assign new_n4519_ = new_n1456_;
  assign new_n4520_ = new_n4519_;
  assign new_n4521_ = new_n4519_;
  assign new_n4522_ = new_n1895_;
  assign new_n4523_ = new_n4522_;
  assign new_n4524_ = new_n4523_;
  assign new_n4525_ = new_n4523_;
  assign new_n4526_ = new_n4522_;
  assign new_n4527_ = new_n1893_;
  assign new_n4528_ = new_n4527_;
  assign new_n4529_ = new_n4528_;
  assign new_n4530_ = new_n4528_;
  assign new_n4531_ = new_n4527_;
  assign new_n4532_ = new_n1889_;
  assign new_n4533_ = new_n4532_;
  assign new_n4534_ = new_n4533_;
  assign new_n4535_ = new_n4533_;
  assign new_n4536_ = new_n4532_;
  assign new_n4537_ = new_n4536_;
  assign new_n4538_ = new_n1883_;
  assign new_n4539_ = new_n4538_;
  assign new_n4540_ = new_n4539_;
  assign new_n4541_ = new_n4539_;
  assign new_n4542_ = new_n4538_;
  assign new_n4543_ = new_n1897_;
  assign new_n4544_ = new_n4543_;
  assign new_n4545_ = new_n4544_;
  assign new_n4546_ = new_n4544_;
  assign new_n4547_ = new_n4543_;
  assign new_n4548_ = new_n4547_;
  assign new_n4549_ = new_n1444_;
  assign new_n4550_ = new_n4549_;
  assign new_n4551_ = new_n4550_;
  assign new_n4552_ = new_n4550_;
  assign new_n4553_ = new_n4549_;
  assign new_n4554_ = new_n1446_;
  assign new_n4555_ = new_n4554_;
  assign new_n4556_ = new_n4555_;
  assign new_n4557_ = new_n4554_;
  assign new_n4558_ = new_n1879_;
  assign new_n4559_ = new_n4558_;
  assign new_n4560_ = new_n4559_;
  assign new_n4561_ = new_n4560_;
  assign new_n4562_ = new_n4559_;
  assign new_n4563_ = new_n4558_;
  assign new_n4564_ = new_n4563_;
  assign new_n4565_ = new_n4563_;
  assign new_n4566_ = new_n2581_;
  assign new_n4567_ = new_n4566_;
  assign new_n4568_ = new_n4567_;
  assign new_n4569_ = new_n4567_;
  assign new_n4570_ = new_n4566_;
  assign new_n4571_ = new_n4570_;
  assign new_n4572_ = new_n1397_;
  assign new_n4573_ = new_n4572_;
  assign new_n4574_ = new_n4572_;
  assign new_n4575_ = new_n1398_;
  assign new_n4576_ = new_n4575_;
  assign new_n4577_ = new_n4575_;
  assign new_n4578_ = new_n2586_;
  assign new_n4579_ = new_n4578_;
  assign new_n4580_ = new_n4578_;
  assign new_n4581_ = new_n2580_;
  assign new_n4582_ = new_n4581_;
  assign new_n4583_ = new_n4581_;
  assign new_n4584_ = new_n2589_;
  assign new_n4585_ = new_n4584_;
  assign new_n4586_ = new_n4584_;
  assign new_n4587_ = new_n2504_;
  assign new_n4588_ = new_n4587_;
  assign new_n4589_ = new_n4588_;
  assign new_n4590_ = new_n4588_;
  assign new_n4591_ = new_n4587_;
  assign new_n4592_ = new_n4591_;
  assign new_n4593_ = new_n4591_;
  assign new_n4594_ = new_n2505_;
  assign new_n4595_ = new_n4594_;
  assign new_n4596_ = new_n2594_;
  assign new_n4597_ = new_n4596_;
  assign new_n4598_ = new_n4597_;
  assign new_n4599_ = new_n4597_;
  assign new_n4600_ = new_n4596_;
  assign new_n4601_ = new_n1949_;
  assign new_n4602_ = new_n4601_;
  assign new_n4603_ = new_n2516_;
  assign new_n4604_ = new_n1950_;
  assign new_n4605_ = new_n4604_;
  assign new_n4606_ = new_n1661_;
  assign new_n4607_ = new_n4606_;
  assign new_n4608_ = new_n1662_;
  assign new_n4609_ = new_n2607_;
  assign new_n4610_ = new_n1881_;
  assign new_n4611_ = new_n4610_;
  assign new_n4612_ = new_n4611_;
  assign new_n4613_ = new_n4611_;
  assign new_n4614_ = new_n4610_;
  assign new_n4615_ = new_n1872_;
  assign new_n4616_ = new_n1870_;
  assign new_n4617_ = new_n4616_;
  assign new_n4618_ = new_n2655_;
  assign new_n4619_ = new_n4618_;
  assign new_n4620_ = new_n1946_;
  assign new_n4621_ = new_n1945_;
  assign new_n4622_ = new_n2658_;
  assign new_n4623_ = new_n4622_;
  assign new_n4624_ = new_n2496_;
  assign new_n4625_ = new_n2662_;
  assign new_n4626_ = new_n4625_;
  assign new_n4627_ = new_n2659_;
  assign new_n4628_ = new_n4627_;
  assign new_n4629_ = new_n2661_;
  assign new_n4630_ = new_n4629_;
  assign new_n4631_ = new_n2663_;
  assign new_n4632_ = new_n2656_;
  assign new_n4633_ = new_n4632_;
  assign new_n4634_ = new_n2668_;
  assign new_n4635_ = new_n1894_;
  assign new_n4636_ = new_n1896_;
  assign new_n4637_ = new_n1882_;
  assign new_n4638_ = new_n1886_;
  assign new_n4639_ = new_n1754_;
  assign new_n4640_ = new_n1451_;
  assign new_n4641_ = new_n1873_;
  assign new_n4642_ = new_n1884_;
  assign new_n4643_ = new_n1443_;
  assign new_n4644_ = new_n1445_;
  assign new_n4645_ = new_n1455_;
  assign new_n4646_ = new_n1869_;
  assign new_n4647_ = new_n1871_;
  assign new_n4648_ = new_n2499_;
  assign new_n4649_ = new_n2664_;
  assign new_n4650_ = new_n2669_;
  assign new_n4651_ = new_n2593_;
  assign new_n4652_ = new_n1639_;
  assign new_n4653_ = new_n1947_;
  assign new_n4654_ = new_n2493_;
  assign new_n4655_ = new_n1425_;
  assign new_n4656_ = new_n1956_;
  assign new_n4657_ = new_n4656_;
  assign new_n4658_ = new_n1955_;
  assign new_n4659_ = new_n4658_;
  assign new_n4660_ = new_n1723_;
  assign new_n4661_ = new_n2834_;
  assign new_n4662_ = new_n1725_;
  assign new_n4663_ = new_n2835_;
  assign new_n4664_ = new_n2837_;
  assign new_n4665_ = new_n4664_;
  assign new_n4666_ = new_n4665_;
  assign new_n4667_ = new_n4665_;
  assign new_n4668_ = new_n4664_;
  assign new_n4669_ = new_n4668_;
  assign new_n4670_ = new_n4668_;
  assign new_n4671_ = new_n2511_;
  assign new_n4672_ = new_n2836_;
  assign new_n4673_ = new_n4672_;
  assign new_n4674_ = new_n4673_;
  assign new_n4675_ = new_n4673_;
  assign new_n4676_ = new_n4672_;
  assign new_n4677_ = new_n4676_;
  assign new_n4678_ = new_n4676_;
  assign new_n4679_ = new_n2155_;
  assign new_n4680_ = new_n4679_;
  assign new_n4681_ = new_n4679_;
  assign new_n4682_ = new_n2149_;
  assign new_n4683_ = new_n4682_;
  assign new_n4684_ = new_n4682_;
  assign new_n4685_ = new_n2156_;
  assign new_n4686_ = new_n4685_;
  assign new_n4687_ = new_n2150_;
  assign new_n4688_ = new_n4687_;
  assign new_n4689_ = new_n2846_;
  assign new_n4690_ = new_n4689_;
  assign new_n4691_ = new_n4689_;
  assign new_n4692_ = new_n2847_;
  assign new_n4693_ = new_n4692_;
  assign new_n4694_ = new_n1962_;
  assign new_n4695_ = new_n1919_;
  assign new_n4696_ = new_n1961_;
  assign new_n4697_ = new_n1920_;
  assign new_n4698_ = new_n2864_;
  assign new_n4699_ = new_n4698_;
  assign new_n4700_ = new_n2187_;
  assign new_n4701_ = new_n4700_;
  assign new_n4702_ = new_n1667_;
  assign new_n4703_ = new_n2188_;
  assign new_n4704_ = new_n4703_;
  assign new_n4705_ = new_n2210_;
  assign new_n4706_ = new_n2209_;
  assign new_n4707_ = new_n1669_;
  assign new_n4708_ = new_n1670_;
  assign new_n4709_ = new_n2212_;
  assign new_n4710_ = new_n2211_;
  assign new_n4711_ = new_n2190_;
  assign new_n4712_ = new_n4711_;
  assign new_n4713_ = new_n1671_;
  assign new_n4714_ = new_n2189_;
  assign new_n4715_ = new_n4714_;
  assign new_n4716_ = new_n1672_;
  assign new_n4717_ = new_n1673_;
  assign new_n4718_ = new_n1674_;
  assign new_n4719_ = new_n4718_;
  assign new_n4720_ = new_n2876_;
  assign new_n4721_ = new_n2889_;
  assign new_n4722_ = new_n4721_;
  assign new_n4723_ = new_n4722_;
  assign new_n4724_ = new_n4722_;
  assign new_n4725_ = new_n4721_;
  assign new_n4726_ = new_n2153_;
  assign new_n4727_ = new_n2890_;
  assign new_n4728_ = new_n4727_;
  assign new_n4729_ = new_n2897_;
  assign new_n4730_ = new_n4729_;
  assign new_n4731_ = new_n2615_;
  assign new_n4732_ = new_n2524_;
  assign new_n4733_ = new_n2719_;
  assign new_n4734_ = new_n2833_;
  assign new_n4735_ = new_n2531_;
  assign new_n4736_ = new_n2770_;
  assign new_n4737_ = new_n2827_;
  assign new_n4738_ = new_n2538_;
  assign new_n4739_ = new_n2595_;
  assign new_n4740_ = new_n2604_;
  assign new_n4741_ = new_n2542_;
  assign new_n4742_ = new_n2673_;
  assign new_n4743_ = new_n1538_;
  assign new_n4744_ = new_n1523_;
  assign new_n4745_ = new_n1537_;
  assign new_n4746_ = new_n1524_;
  assign new_n4747_ = new_n2919_;
  assign new_n4748_ = new_n1839_;
  assign new_n4749_ = new_n4748_;
  assign new_n4750_ = new_n1843_;
  assign new_n4751_ = new_n4750_;
  assign new_n4752_ = new_n1828_;
  assign new_n4753_ = new_n4752_;
  assign new_n4754_ = new_n1831_;
  assign new_n4755_ = new_n4754_;
  assign new_n4756_ = new_n1847_;
  assign new_n4757_ = new_n4756_;
  assign new_n4758_ = new_n1819_;
  assign new_n4759_ = new_n4758_;
  assign new_n4760_ = new_n1836_;
  assign new_n4761_ = new_n4760_;
  assign new_n4762_ = new_n1823_;
  assign new_n4763_ = new_n4762_;
  assign new_n4764_ = new_n1248_;
  assign new_n4765_ = new_n1841_;
  assign new_n4766_ = new_n4765_;
  assign new_n4767_ = new_n1845_;
  assign new_n4768_ = new_n4767_;
  assign new_n4769_ = new_n1830_;
  assign new_n4770_ = new_n4769_;
  assign new_n4771_ = new_n1833_;
  assign new_n4772_ = new_n4771_;
  assign new_n4773_ = new_n1849_;
  assign new_n4774_ = new_n4773_;
  assign new_n4775_ = new_n1821_;
  assign new_n4776_ = new_n4775_;
  assign new_n4777_ = new_n1838_;
  assign new_n4778_ = new_n4777_;
  assign new_n4779_ = new_n1825_;
  assign new_n4780_ = new_n4779_;
  assign new_n4781_ = new_n1756_;
  assign new_n4782_ = new_n2609_;
  assign new_n4783_ = new_n2608_;
  assign new_n4784_ = new_n2821_;
  assign new_n4785_ = new_n1697_;
  assign new_n4786_ = new_n1695_;
  assign new_n4787_ = new_n1698_;
  assign new_n4788_ = new_n1696_;
  assign new_n4789_ = new_n1699_;
  assign new_n4790_ = new_n1700_;
  assign new_n4791_ = new_n1731_;
  assign new_n4792_ = new_n1732_;
  assign new_n4793_ = new_n2173_;
  assign new_n4794_ = new_n2174_;
  assign new_n4795_ = new_n2852_;
  assign new_n4796_ = new_n3065_;
  assign new_n4797_ = new_n2866_;
  assign new_n4798_ = new_n3011_;
  assign new_n4799_ = new_n3059_;
  assign new_n4800_ = new_n2898_;
  assign new_n4801_ = new_n2969_;
  assign new_n4802_ = new_n3066_;
  assign new_n4803_ = new_n2920_;
  assign new_n4804_ = new_n3053_;
  assign new_n4805_ = new_n3100_;
  assign new_n4806_ = new_n3103_;
  assign new_n4807_ = new_n3106_;
  assign new_n4808_ = new_n2218_;
  assign new_n4809_ = new_n2180_;
  assign new_n4810_ = new_n2217_;
  assign new_n4811_ = new_n4810_;
  assign new_n4812_ = new_n2179_;
  assign new_n4813_ = new_n4812_;
  assign new_n4814_ = new_n3122_;
  assign new_n4815_ = new_n3120_;
  assign new_n4816_ = new_n3121_;
  assign new_n4817_ = new_n4816_;
  assign new_n4818_ = new_n3119_;
  assign new_n4819_ = new_n4818_;
  assign new_n4820_ = new_n4818_;
  assign new_n4821_ = new_n3114_;
  assign new_n4822_ = new_n3123_;
  assign new_n4823_ = new_n3113_;
  assign new_n4824_ = new_n1605_;
  assign new_n4825_ = new_n4824_;
  assign new_n4826_ = new_n1600_;
  assign new_n4827_ = new_n1606_;
  assign new_n4828_ = new_n1599_;
  assign new_n4829_ = new_n4828_;
  assign new_n4830_ = new_n1624_;
  assign new_n4831_ = new_n1601_;
  assign new_n4832_ = new_n4831_;
  assign new_n4833_ = new_n1623_;
  assign new_n4834_ = new_n4833_;
  assign new_n4835_ = new_n1602_;
  assign new_n4836_ = new_n2894_;
  assign new_n4837_ = new_n4836_;
  assign new_n4838_ = new_n2839_;
  assign new_n4839_ = new_n4838_;
  assign new_n4840_ = new_n4839_;
  assign new_n4841_ = new_n4839_;
  assign new_n4842_ = new_n4838_;
  assign new_n4843_ = new_n3112_;
  assign new_n4844_ = new_n2220_;
  assign new_n4845_ = new_n2182_;
  assign new_n4846_ = new_n2219_;
  assign new_n4847_ = new_n4846_;
  assign new_n4848_ = new_n2181_;
  assign new_n4849_ = new_n4848_;
  assign new_n4850_ = new_n3149_;
  assign new_n4851_ = new_n3147_;
  assign new_n4852_ = new_n4851_;
  assign new_n4853_ = new_n3150_;
  assign new_n4854_ = new_n3148_;
  assign new_n4855_ = new_n4854_;
  assign new_n4856_ = new_n4854_;
  assign new_n4857_ = new_n2222_;
  assign new_n4858_ = new_n2192_;
  assign new_n4859_ = new_n2221_;
  assign new_n4860_ = new_n2191_;
  assign new_n4861_ = new_n3157_;
  assign new_n4862_ = new_n4861_;
  assign new_n4863_ = new_n4861_;
  assign new_n4864_ = new_n3158_;
  assign new_n4865_ = new_n4864_;
  assign new_n4866_ = new_n4865_;
  assign new_n4867_ = new_n4865_;
  assign new_n4868_ = new_n4864_;
  assign new_n4869_ = new_n3161_;
  assign new_n4870_ = new_n3160_;
  assign new_n4871_ = new_n4870_;
  assign new_n4872_ = new_n3162_;
  assign new_n4873_ = new_n3159_;
  assign new_n4874_ = new_n4873_;
  assign new_n4875_ = new_n2858_;
  assign new_n4876_ = new_n4875_;
  assign new_n4877_ = new_n4875_;
  assign new_n4878_ = new_n2859_;
  assign new_n4879_ = new_n4878_;
  assign new_n4880_ = new_n4879_;
  assign new_n4881_ = new_n4878_;
  assign new_n4882_ = new_n2838_;
  assign new_n4883_ = new_n4882_;
  assign new_n4884_ = new_n4883_;
  assign new_n4885_ = new_n4882_;
  assign new_n4886_ = new_n1479_;
  assign new_n4887_ = new_n1477_;
  assign new_n4888_ = new_n4887_;
  assign new_n4889_ = new_n3175_;
  assign new_n4890_ = new_n3094_;
  assign new_n4891_ = new_n4890_;
  assign new_n4892_ = new_n3096_;
  assign new_n4893_ = new_n4892_;
  assign new_n4894_ = new_n1931_;
  assign new_n4895_ = new_n1932_;
  assign new_n4896_ = new_n3179_;
  assign new_n4897_ = new_n3178_;
  assign new_n4898_ = new_n4897_;
  assign new_n4899_ = new_n2203_;
  assign new_n4900_ = new_n4899_;
  assign new_n4901_ = new_n4899_;
  assign new_n4902_ = new_n2201_;
  assign new_n4903_ = new_n4902_;
  assign new_n4904_ = new_n4903_;
  assign new_n4905_ = new_n4903_;
  assign new_n4906_ = new_n4902_;
  assign new_n4907_ = new_n4906_;
  assign new_n4908_ = new_n4906_;
  assign new_n4909_ = new_n2202_;
  assign new_n4910_ = new_n4909_;
  assign new_n4911_ = new_n4910_;
  assign new_n4912_ = new_n4910_;
  assign new_n4913_ = new_n4909_;
  assign new_n4914_ = new_n3186_;
  assign new_n4915_ = new_n4914_;
  assign new_n4916_ = new_n3187_;
  assign new_n4917_ = new_n4916_;
  assign new_n4918_ = new_n2208_;
  assign new_n4919_ = new_n2207_;
  assign new_n4920_ = new_n4919_;
  assign new_n4921_ = new_n3189_;
  assign new_n4922_ = new_n4921_;
  assign new_n4923_ = new_n4922_;
  assign new_n4924_ = new_n4923_;
  assign new_n4925_ = new_n4922_;
  assign new_n4926_ = new_n4921_;
  assign new_n4927_ = new_n4926_;
  assign new_n4928_ = new_n4926_;
  assign new_n4929_ = new_n2243_;
  assign new_n4930_ = new_n4929_;
  assign new_n4931_ = new_n4929_;
  assign new_n4932_ = new_n3188_;
  assign new_n4933_ = new_n4932_;
  assign new_n4934_ = new_n4933_;
  assign new_n4935_ = new_n4933_;
  assign new_n4936_ = new_n4932_;
  assign new_n4937_ = new_n4936_;
  assign new_n4938_ = new_n2244_;
  assign new_n4939_ = new_n4938_;
  assign new_n4940_ = new_n3191_;
  assign new_n4941_ = new_n3190_;
  assign new_n4942_ = new_n2247_;
  assign new_n4943_ = new_n2248_;
  assign new_n4944_ = new_n3196_;
  assign new_n4945_ = new_n3197_;
  assign new_n4946_ = new_n2237_;
  assign new_n4947_ = new_n4946_;
  assign new_n4948_ = new_n4947_;
  assign new_n4949_ = new_n4947_;
  assign new_n4950_ = new_n4946_;
  assign new_n4951_ = new_n2230_;
  assign new_n4952_ = new_n4951_;
  assign new_n4953_ = new_n4952_;
  assign new_n4954_ = new_n4952_;
  assign new_n4955_ = new_n4951_;
  assign new_n4956_ = new_n4955_;
  assign new_n4957_ = new_n4955_;
  assign new_n4958_ = new_n2238_;
  assign new_n4959_ = new_n4958_;
  assign new_n4960_ = new_n4959_;
  assign new_n4961_ = new_n4958_;
  assign new_n4962_ = new_n2229_;
  assign new_n4963_ = new_n4962_;
  assign new_n4964_ = new_n4963_;
  assign new_n4965_ = new_n4963_;
  assign new_n4966_ = new_n4962_;
  assign new_n4967_ = new_n2271_;
  assign new_n4968_ = new_n4967_;
  assign new_n4969_ = new_n4967_;
  assign new_n4970_ = new_n2186_;
  assign new_n4971_ = new_n4970_;
  assign new_n4972_ = new_n4971_;
  assign new_n4973_ = new_n4971_;
  assign new_n4974_ = new_n4970_;
  assign new_n4975_ = new_n4974_;
  assign new_n4976_ = new_n4974_;
  assign new_n4977_ = new_n2272_;
  assign new_n4978_ = new_n4977_;
  assign new_n4979_ = new_n2185_;
  assign new_n4980_ = new_n4979_;
  assign new_n4981_ = new_n4980_;
  assign new_n4982_ = new_n4980_;
  assign new_n4983_ = new_n4979_;
  assign new_n4984_ = new_n3204_;
  assign new_n4985_ = new_n4984_;
  assign new_n4986_ = new_n4985_;
  assign new_n4987_ = new_n4985_;
  assign new_n4988_ = new_n4984_;
  assign new_n4989_ = new_n4988_;
  assign new_n4990_ = new_n2241_;
  assign new_n4991_ = new_n4990_;
  assign new_n4992_ = new_n4990_;
  assign new_n4993_ = new_n3205_;
  assign new_n4994_ = new_n4993_;
  assign new_n4995_ = new_n4994_;
  assign new_n4996_ = new_n4993_;
  assign new_n4997_ = new_n2242_;
  assign new_n4998_ = new_n4997_;
  assign new_n4999_ = new_n2274_;
  assign new_n5000_ = new_n2273_;
  assign new_n5001_ = new_n2161_;
  assign new_n5002_ = new_n2245_;
  assign new_n5003_ = new_n5002_;
  assign new_n5004_ = new_n5002_;
  assign new_n5005_ = new_n2246_;
  assign new_n5006_ = new_n3221_;
  assign new_n5007_ = new_n5006_;
  assign new_n5008_ = new_n5006_;
  assign new_n5009_ = new_n3220_;
  assign new_n5010_ = new_n5009_;
  assign new_n5011_ = new_n2249_;
  assign new_n5012_ = new_n5011_;
  assign new_n5013_ = new_n2250_;
  assign new_n5014_ = new_n3227_;
  assign new_n5015_ = new_n3226_;
  assign new_n5016_ = new_n5015_;
  assign new_n5017_ = new_n1295_;
  assign new_n5018_ = new_n5017_;
  assign new_n5019_ = new_n2251_;
  assign new_n5020_ = new_n2277_;
  assign new_n5021_ = new_n5020_;
  assign new_n5022_ = new_n5021_;
  assign new_n5023_ = new_n5022_;
  assign new_n5024_ = new_n5021_;
  assign new_n5025_ = new_n5020_;
  assign new_n5026_ = new_n5025_;
  assign new_n5027_ = new_n5025_;
  assign new_n5028_ = new_n2255_;
  assign new_n5029_ = new_n5028_;
  assign new_n5030_ = new_n5029_;
  assign new_n5031_ = new_n5029_;
  assign new_n5032_ = new_n5028_;
  assign new_n5033_ = new_n5032_;
  assign new_n5034_ = new_n2278_;
  assign new_n5035_ = new_n5034_;
  assign new_n5036_ = new_n5035_;
  assign new_n5037_ = new_n5035_;
  assign new_n5038_ = new_n5034_;
  assign new_n5039_ = new_n5038_;
  assign new_n5040_ = new_n5038_;
  assign new_n5041_ = new_n2256_;
  assign new_n5042_ = new_n5041_;
  assign new_n5043_ = new_n5042_;
  assign new_n5044_ = new_n5041_;
  assign new_n5045_ = new_n2268_;
  assign new_n5046_ = new_n5045_;
  assign new_n5047_ = new_n5046_;
  assign new_n5048_ = new_n5046_;
  assign new_n5049_ = new_n5045_;
  assign new_n5050_ = new_n2259_;
  assign new_n5051_ = new_n5050_;
  assign new_n5052_ = new_n5051_;
  assign new_n5053_ = new_n5052_;
  assign new_n5054_ = new_n5051_;
  assign new_n5055_ = new_n5050_;
  assign new_n5056_ = new_n5055_;
  assign new_n5057_ = new_n5055_;
  assign new_n5058_ = new_n2267_;
  assign new_n5059_ = new_n5058_;
  assign new_n5060_ = new_n5059_;
  assign new_n5061_ = new_n5059_;
  assign new_n5062_ = new_n5058_;
  assign new_n5063_ = new_n5062_;
  assign new_n5064_ = new_n5062_;
  assign new_n5065_ = new_n2260_;
  assign new_n5066_ = new_n5065_;
  assign new_n5067_ = new_n5066_;
  assign new_n5068_ = new_n5066_;
  assign new_n5069_ = new_n5065_;
  assign new_n5070_ = new_n5069_;
  assign new_n5071_ = new_n5069_;
  assign new_n5072_ = new_n3268_;
  assign new_n5073_ = new_n5072_;
  assign new_n5074_ = new_n5073_;
  assign new_n5075_ = new_n5073_;
  assign new_n5076_ = new_n5072_;
  assign new_n5077_ = new_n5076_;
  assign new_n5078_ = new_n5076_;
  assign new_n5079_ = new_n2164_;
  assign new_n5080_ = new_n5079_;
  assign new_n5081_ = new_n5079_;
  assign new_n5082_ = new_n3269_;
  assign new_n5083_ = new_n5082_;
  assign new_n5084_ = new_n5083_;
  assign new_n5085_ = new_n5083_;
  assign new_n5086_ = new_n5082_;
  assign new_n5087_ = new_n5086_;
  assign new_n5088_ = new_n2163_;
  assign new_n5089_ = new_n5088_;
  assign new_n5090_ = new_n5089_;
  assign new_n5091_ = new_n5089_;
  assign new_n5092_ = new_n5088_;
  assign new_n5093_ = new_n2205_;
  assign new_n5094_ = new_n5093_;
  assign new_n5095_ = new_n5094_;
  assign new_n5096_ = new_n5093_;
  assign new_n5097_ = new_n2206_;
  assign new_n5098_ = new_n1855_;
  assign new_n5099_ = new_n5098_;
  assign new_n5100_ = new_n1856_;
  assign new_n5101_ = new_n3281_;
  assign new_n5102_ = new_n5101_;
  assign new_n5103_ = new_n5102_;
  assign new_n5104_ = new_n5103_;
  assign new_n5105_ = new_n5102_;
  assign new_n5106_ = new_n5101_;
  assign new_n5107_ = new_n5106_;
  assign new_n5108_ = new_n5106_;
  assign new_n5109_ = new_n3280_;
  assign new_n5110_ = new_n5109_;
  assign new_n5111_ = new_n5110_;
  assign new_n5112_ = new_n5110_;
  assign new_n5113_ = new_n5109_;
  assign new_n5114_ = new_n5113_;
  assign new_n5115_ = new_n5113_;
  assign new_n5116_ = new_n3284_;
  assign new_n5117_ = new_n5116_;
  assign new_n5118_ = new_n5117_;
  assign new_n5119_ = new_n5118_;
  assign new_n5120_ = new_n5117_;
  assign new_n5121_ = new_n5116_;
  assign new_n5122_ = new_n5121_;
  assign new_n5123_ = new_n5121_;
  assign new_n5124_ = new_n3285_;
  assign new_n5125_ = new_n5124_;
  assign new_n5126_ = new_n5125_;
  assign new_n5127_ = new_n5125_;
  assign new_n5128_ = new_n5124_;
  assign new_n5129_ = new_n5128_;
  assign new_n5130_ = new_n5128_;
  assign new_n5131_ = new_n3289_;
  assign new_n5132_ = new_n5131_;
  assign new_n5133_ = new_n5131_;
  assign new_n5134_ = new_n3288_;
  assign new_n5135_ = new_n5134_;
  assign new_n5136_ = new_n3290_;
  assign new_n5137_ = new_n5136_;
  assign new_n5138_ = new_n5137_;
  assign new_n5139_ = new_n5137_;
  assign new_n5140_ = new_n5136_;
  assign new_n5141_ = new_n5140_;
  assign new_n5142_ = new_n5140_;
  assign new_n5143_ = new_n3291_;
  assign new_n5144_ = new_n5143_;
  assign new_n5145_ = new_n5144_;
  assign new_n5146_ = new_n5144_;
  assign new_n5147_ = new_n5143_;
  assign new_n5148_ = new_n5147_;
  assign new_n5149_ = new_n3301_;
  assign new_n5150_ = new_n5149_;
  assign new_n5151_ = new_n5150_;
  assign new_n5152_ = new_n5151_;
  assign new_n5153_ = new_n5150_;
  assign new_n5154_ = new_n5149_;
  assign new_n5155_ = new_n5154_;
  assign new_n5156_ = new_n5154_;
  assign new_n5157_ = new_n3300_;
  assign new_n5158_ = new_n5157_;
  assign new_n5159_ = new_n5158_;
  assign new_n5160_ = new_n5158_;
  assign new_n5161_ = new_n5157_;
  assign new_n5162_ = new_n5161_;
  assign new_n5163_ = new_n3303_;
  assign new_n5164_ = new_n5163_;
  assign new_n5165_ = new_n5164_;
  assign new_n5166_ = new_n5163_;
  assign new_n5167_ = new_n3302_;
  assign new_n5168_ = new_n5167_;
  assign new_n5169_ = new_n5167_;
  assign new_n5170_ = new_n1859_;
  assign new_n5171_ = new_n5170_;
  assign new_n5172_ = new_n5171_;
  assign new_n5173_ = new_n5171_;
  assign new_n5174_ = new_n5170_;
  assign new_n5175_ = new_n5174_;
  assign new_n5176_ = new_n5174_;
  assign new_n5177_ = new_n1860_;
  assign new_n5178_ = new_n5177_;
  assign new_n5179_ = new_n5178_;
  assign new_n5180_ = new_n5178_;
  assign new_n5181_ = new_n5177_;
  assign new_n5182_ = new_n2269_;
  assign new_n5183_ = new_n5182_;
  assign new_n5184_ = new_n5182_;
  assign new_n5185_ = new_n2270_;
  assign new_n5186_ = new_n5185_;
  assign new_n5187_ = new_n3311_;
  assign new_n5188_ = new_n5187_;
  assign new_n5189_ = new_n3310_;
  assign new_n5190_ = new_n5189_;
  assign new_n5191_ = new_n5189_;
  assign new_n5192_ = new_n3298_;
  assign new_n5193_ = new_n5192_;
  assign new_n5194_ = new_n5193_;
  assign new_n5195_ = new_n5192_;
  assign new_n5196_ = new_n1270_;
  assign new_n5197_ = new_n5196_;
  assign new_n5198_ = new_n5197_;
  assign new_n5199_ = new_n5197_;
  assign new_n5200_ = new_n5196_;
  assign new_n5201_ = new_n3327_;
  assign new_n5202_ = new_n1272_;
  assign new_n5203_ = new_n5202_;
  assign new_n5204_ = new_n5203_;
  assign new_n5205_ = new_n5203_;
  assign new_n5206_ = new_n5202_;
  assign new_n5207_ = new_n3091_;
  assign new_n5208_ = new_n5207_;
  assign new_n5209_ = new_n1858_;
  assign new_n5210_ = new_n5209_;
  assign new_n5211_ = new_n5210_;
  assign new_n5212_ = new_n5209_;
  assign new_n5213_ = new_n1857_;
  assign new_n5214_ = new_n5213_;
  assign new_n5215_ = new_n5214_;
  assign new_n5216_ = new_n5214_;
  assign new_n5217_ = new_n5213_;
  assign new_n5218_ = new_n5217_;
  assign new_n5219_ = new_n5217_;
  assign new_n5220_ = new_n2235_;
  assign new_n5221_ = new_n5220_;
  assign new_n5222_ = new_n5221_;
  assign new_n5223_ = new_n5220_;
  assign new_n5224_ = new_n2236_;
  assign new_n5225_ = new_n2165_;
  assign new_n5226_ = new_n5225_;
  assign new_n5227_ = new_n5226_;
  assign new_n5228_ = new_n5226_;
  assign new_n5229_ = new_n5225_;
  assign new_n5230_ = new_n5229_;
  assign new_n5231_ = new_n5229_;
  assign new_n5232_ = new_n2166_;
  assign new_n5233_ = new_n5232_;
  assign new_n5234_ = new_n5233_;
  assign new_n5235_ = new_n5233_;
  assign new_n5236_ = new_n5232_;
  assign new_n5237_ = new_n2257_;
  assign new_n5238_ = new_n5237_;
  assign new_n5239_ = new_n5237_;
  assign new_n5240_ = new_n2258_;
  assign new_n5241_ = new_n3358_;
  assign new_n5242_ = new_n5241_;
  assign new_n5243_ = new_n5242_;
  assign new_n5244_ = new_n5241_;
  assign new_n5245_ = new_n3379_;
  assign new_n5246_ = new_n3405_;
  assign new_n5247_ = new_n5246_;
  assign new_n5248_ = new_n5246_;
  assign new_n5249_ = new_n3404_;
  assign new_n5250_ = new_n5249_;
  assign new_n5251_ = new_n5249_;
  assign new_n5252_ = new_n1299_;
  assign new_n5253_ = new_n1303_;
  assign new_n5254_ = new_n1267_;
  assign new_n5255_ = new_n2239_;
  assign new_n5256_ = new_n3476_;
  assign new_n5257_ = new_n5256_;
  assign new_n5258_ = new_n5257_;
  assign new_n5259_ = new_n5256_;
  assign new_n5260_ = new_n3497_;
  assign new_n5261_ = new_n3337_;
  assign new_n5262_ = new_n3502_;
  assign new_n5263_ = new_n5262_;
  assign new_n5264_ = new_n3331_;
  assign new_n5265_ = new_n3329_;
  assign new_n5266_ = new_n1273_;
  assign new_n5267_ = new_n5266_;
  assign new_n5268_ = new_n5266_;
  assign new_n5269_ = new_n3326_;
  assign new_n5270_ = new_n1275_;
  assign new_n5271_ = new_n5270_;
  assign new_n5272_ = new_n5270_;
  assign new_n5273_ = new_n3092_;
  assign new_n5274_ = new_n1328_;
  assign new_n5275_ = new_n5274_;
  assign new_n5276_ = new_n5275_;
  assign new_n5277_ = new_n5275_;
  assign new_n5278_ = new_n5274_;
  assign new_n5279_ = new_n5278_;
  assign new_n5280_ = new_n3333_;
  assign new_n5281_ = new_n1621_;
  assign new_n5282_ = new_n5281_;
  assign new_n5283_ = new_n5281_;
  assign new_n5284_ = new_n2908_;
  assign new_n5285_ = new_n5284_;
  assign new_n5286_ = new_n2902_;
  assign new_n5287_ = new_n5286_;
  assign new_n5288_ = new_n3068_;
  assign new_n5289_ = new_n5288_;
  assign new_n5290_ = new_n2904_;
  assign new_n5291_ = new_n5290_;
  assign new_n5292_ = new_n3545_;
  assign new_n5293_ = new_n3544_;
  assign new_n5294_ = new_n5293_;
  assign new_n5295_ = new_n3550_;
  assign new_n5296_ = new_n5295_;
  assign new_n5297_ = new_n5295_;
  assign new_n5298_ = new_n3334_;
  assign new_n5299_ = new_n5298_;
  assign new_n5300_ = new_n3524_;
  assign new_n5301_ = new_n3449_;
  assign new_n5302_ = new_n5301_;
  assign new_n5303_ = new_n5302_;
  assign new_n5304_ = new_n5301_;
  assign new_n5305_ = new_n3503_;
  assign new_n5306_ = new_n5305_;
  assign new_n5307_ = new_n5306_;
  assign new_n5308_ = new_n5305_;
  assign new_n5309_ = new_n3184_;
  assign new_n5310_ = new_n1625_;
  assign new_n5311_ = new_n1627_;
  assign new_n5312_ = new_n1657_;
  assign new_n5313_ = new_n1675_;
  assign new_n5314_ = new_n3551_;
  assign new_n5315_ = new_n5314_;
  assign new_n5316_ = new_n3125_;
  assign new_n5317_ = new_n1529_;
  assign new_n5318_ = new_n5317_;
  assign new_n5319_ = new_n1535_;
  assign new_n5320_ = new_n5319_;
  assign new_n5321_ = new_n5319_;
  assign new_n5322_ = new_n1597_;
  assign new_n5323_ = new_n5322_;
  assign new_n5324_ = new_n5322_;
  assign new_n5325_ = new_n3579_;
  assign new_n5326_ = new_n3578_;
  assign new_n5327_ = new_n5326_;
  assign new_n5328_ = new_n1549_;
  assign new_n5329_ = new_n5328_;
  assign new_n5330_ = new_n5329_;
  assign new_n5331_ = new_n5328_;
  assign new_n5332_ = new_n1550_;
  assign new_n5333_ = new_n5332_;
  assign new_n5334_ = new_n3603_;
  assign new_n5335_ = new_n5334_;
  assign new_n5336_ = new_n3605_;
  assign new_n5337_ = new_n3602_;
  assign new_n5338_ = new_n5337_;
  assign new_n5339_ = new_n5337_;
  assign new_n5340_ = new_n3601_;
  assign new_n5341_ = new_n5340_;
  assign new_n5342_ = new_n5340_;
  assign new_n5343_ = new_n3608_;
  assign new_n5344_ = new_n3609_;
  assign new_n5345_ = new_n3611_;
  assign new_n5346_ = new_n3613_;
  assign new_n5347_ = new_n3383_;
  assign new_n5348_ = new_n3381_;
  assign new_n5349_ = new_n3378_;
  assign new_n5350_ = new_n1604_;
  assign new_n5351_ = new_n5350_;
  assign new_n5352_ = new_n1528_;
  assign new_n5353_ = new_n5352_;
  assign new_n5354_ = new_n3539_;
  assign new_n5355_ = new_n1619_;
  assign new_n5356_ = new_n5355_;
  assign new_n5357_ = new_n5356_;
  assign new_n5358_ = new_n5355_;
  assign new_n5359_ = new_n1534_;
  assign new_n5360_ = new_n5359_;
  assign new_n5361_ = new_n3630_;
  assign new_n5362_ = new_n3536_;
  assign new_n5363_ = new_n3562_;
  assign new_n5364_ = new_n5363_;
  assign new_n5365_ = new_n5363_;
  assign new_n5366_ = new_n3560_;
  assign new_n5367_ = new_n5366_;
  assign new_n5368_ = new_n5366_;
  assign new_n5369_ = new_n3641_;
  assign new_n5370_ = new_n5369_;
  assign new_n5371_ = new_n3634_;
  assign new_n5372_ = new_n5371_;
  assign new_n5373_ = new_n3668_;
  assign new_n5374_ = new_n5373_;
  assign new_n5375_ = new_n5373_;
  assign new_n5376_ = new_n1269_;
  assign new_n5377_ = new_n5376_;
  assign new_n5378_ = new_n5376_;
  assign new_n5379_ = new_n3667_;
  assign new_n5380_ = new_n5379_;
  assign new_n5381_ = new_n5379_;
  assign new_n5382_ = new_n3262_;
  assign new_n5383_ = new_n3263_;
  assign new_n5384_ = new_n5383_;
  assign new_n5385_ = new_n5384_;
  assign new_n5386_ = new_n5383_;
  assign new_n5387_ = new_n1271_;
  assign new_n5388_ = new_n5387_;
  assign new_n5389_ = new_n5388_;
  assign new_n5390_ = new_n5387_;
  assign new_n5391_ = new_n3413_;
  assign new_n5392_ = new_n5391_;
  assign new_n5393_ = new_n5392_;
  assign new_n5394_ = new_n5391_;
  assign new_n5395_ = new_n3412_;
  assign new_n5396_ = new_n5395_;
  assign new_n5397_ = new_n3242_;
  assign new_n5398_ = new_n3243_;
  assign new_n5399_ = new_n5398_;
  assign new_n5400_ = new_n5399_;
  assign new_n5401_ = new_n5398_;
  assign new_n5402_ = new_n1547_;
  assign new_n5403_ = new_n1545_;
  assign new_n5404_ = new_n5403_;
  assign new_n5405_ = new_n1533_;
  assign new_n5406_ = new_n5405_;
  assign new_n5407_ = new_n5406_;
  assign new_n5408_ = new_n5406_;
  assign new_n5409_ = new_n5405_;
  assign new_n5410_ = new_n1527_;
  assign new_n5411_ = new_n5410_;
  assign new_n5412_ = new_n5411_;
  assign new_n5413_ = new_n5411_;
  assign new_n5414_ = new_n5410_;
  assign new_n5415_ = new_n1620_;
  assign new_n5416_ = new_n5415_;
  assign new_n5417_ = new_n3538_;
  assign new_n5418_ = new_n3335_;
  assign new_n5419_ = new_n1327_;
  assign new_n5420_ = new_n3140_;
  assign new_n5421_ = new_n3558_;
  assign new_n5422_ = new_n3556_;
  assign new_n5423_ = new_n1603_;
  assign new_n5424_ = new_n5423_;
  assign new_n5425_ = new_n5424_;
  assign new_n5426_ = new_n5423_;
  assign new_n5427_ = new_n2900_;
  assign new_n5428_ = new_n2899_;
  assign new_n5429_ = new_n5428_;
  assign new_n5430_ = new_n3174_;
  assign new_n5431_ = new_n3132_;
  assign new_n5432_ = new_n3138_;
  assign new_n5433_ = new_n3439_;
  assign new_n5434_ = new_n5433_;
  assign new_n5435_ = new_n5434_;
  assign new_n5436_ = new_n5433_;
  assign new_n5437_ = new_n3216_;
  assign new_n5438_ = new_n1274_;
  assign new_n5439_ = new_n5438_;
  assign new_n5440_ = new_n5438_;
  assign new_n5441_ = new_n3217_;
  assign new_n5442_ = new_n5441_;
  assign new_n5443_ = new_n1276_;
  assign new_n5444_ = new_n5443_;
  assign new_n5445_ = new_n5443_;
  assign new_n5446_ = new_n3741_;
  assign new_n5447_ = new_n3678_;
  assign new_n5448_ = new_n3501_;
  assign new_n5449_ = new_n3499_;
  assign new_n5450_ = new_n3496_;
  assign new_n5451_ = new_n3688_;
  assign new_n5452_ = new_n3525_;
  assign new_n5453_ = new_n5452_;
  assign new_n5454_ = new_n5452_;
  assign new_n5455_ = new_n1139_;
  assign new_n5456_ = new_n5455_;
  assign new_n5457_ = new_n1137_;
  assign new_n5458_ = new_n5457_;
  assign new_n5459_ = new_n5458_;
  assign new_n5460_ = new_n5458_;
  assign new_n5461_ = new_n5457_;
  assign new_n5462_ = new_n5461_;
  assign new_n5463_ = new_n5461_;
  assign new_n5464_ = new_n1265_;
  assign new_n5465_ = new_n3770_;
  assign new_n5466_ = new_n5465_;
  assign new_n5467_ = new_n3748_;
  assign new_n5468_ = new_n5467_;
  assign new_n5469_ = new_n5467_;
  assign new_n5470_ = new_n3696_;
  assign new_n5471_ = new_n3755_;
  assign new_n5472_ = new_n5471_;
  assign new_n5473_ = new_n1141_;
  assign new_n5474_ = new_n3778_;
  assign new_n5475_ = new_n5474_;
  assign new_n5476_ = new_n1135_;
  assign new_n5477_ = new_n5476_;
  assign new_n5478_ = new_n1133_;
  assign new_n5479_ = new_n1551_;
  assign new_n5480_ = new_n5479_;
  assign new_n5481_ = new_n5480_;
  assign new_n5482_ = new_n5479_;
  assign new_n5483_ = new_n2906_;
  assign new_n5484_ = new_n5483_;
  assign new_n5485_ = new_n5483_;
  assign new_n5486_ = new_n3098_;
  assign new_n5487_ = new_n5486_;
  assign new_n5488_ = new_n5486_;
  assign new_n5489_ = new_n3176_;
  assign new_n5490_ = new_n3177_;
  assign new_n5491_ = new_n3533_;
  assign new_n5492_ = new_n5491_;
  assign new_n5493_ = new_n5491_;
  assign new_n5494_ = new_n3553_;
  assign new_n5495_ = new_n3554_;
  assign new_n5496_ = new_n3559_;
  assign new_n5497_ = new_n5496_;
  assign new_n5498_ = new_n3565_;
  assign new_n5499_ = new_n3568_;
  assign new_n5500_ = new_n3571_;
  assign new_n5501_ = new_n3574_;
  assign new_n5502_ = new_n3577_;
  assign new_n5503_ = new_n3600_;
  assign new_n5504_ = new_n3606_;
  assign new_n5505_ = new_n5504_;
  assign new_n5506_ = new_n5505_;
  assign new_n5507_ = new_n5506_;
  assign new_n5508_ = new_n5506_;
  assign new_n5509_ = new_n5505_;
  assign new_n5510_ = new_n5509_;
  assign new_n5511_ = new_n5509_;
  assign new_n5512_ = new_n5504_;
  assign new_n5513_ = new_n5512_;
  assign new_n5514_ = new_n5512_;
  assign new_n5515_ = new_n3607_;
  assign new_n5516_ = new_n5515_;
  assign new_n5517_ = new_n5516_;
  assign new_n5518_ = new_n5517_;
  assign new_n5519_ = new_n5517_;
  assign new_n5520_ = new_n5516_;
  assign new_n5521_ = new_n5520_;
  assign new_n5522_ = new_n5520_;
  assign new_n5523_ = new_n5515_;
  assign new_n5524_ = new_n5523_;
  assign new_n5525_ = new_n5523_;
  assign new_n5526_ = new_n3610_;
  assign new_n5527_ = new_n5526_;
  assign new_n5528_ = new_n5527_;
  assign new_n5529_ = new_n5528_;
  assign new_n5530_ = new_n5528_;
  assign new_n5531_ = new_n5527_;
  assign new_n5532_ = new_n5531_;
  assign new_n5533_ = new_n5531_;
  assign new_n5534_ = new_n5526_;
  assign new_n5535_ = new_n5534_;
  assign new_n5536_ = new_n5534_;
  assign new_n5537_ = new_n3612_;
  assign new_n5538_ = new_n5537_;
  assign new_n5539_ = new_n5538_;
  assign new_n5540_ = new_n5539_;
  assign new_n5541_ = new_n5539_;
  assign new_n5542_ = new_n5538_;
  assign new_n5543_ = new_n5542_;
  assign new_n5544_ = new_n5542_;
  assign new_n5545_ = new_n5537_;
  assign new_n5546_ = new_n5545_;
  assign new_n5547_ = new_n5545_;
  assign new_n5548_ = new_n3614_;
  assign new_n5549_ = new_n5548_;
  assign new_n5550_ = new_n5549_;
  assign new_n5551_ = new_n5550_;
  assign new_n5552_ = new_n5550_;
  assign new_n5553_ = new_n5549_;
  assign new_n5554_ = new_n5553_;
  assign new_n5555_ = new_n5553_;
  assign new_n5556_ = new_n5548_;
  assign new_n5557_ = new_n5556_;
  assign new_n5558_ = new_n5556_;
  assign new_n5559_ = new_n3615_;
  assign new_n5560_ = new_n5559_;
  assign new_n5561_ = new_n5560_;
  assign new_n5562_ = new_n5561_;
  assign new_n5563_ = new_n5561_;
  assign new_n5564_ = new_n5560_;
  assign new_n5565_ = new_n5564_;
  assign new_n5566_ = new_n5564_;
  assign new_n5567_ = new_n5559_;
  assign new_n5568_ = new_n5567_;
  assign new_n5569_ = new_n5567_;
  assign new_n5570_ = new_n3616_;
  assign new_n5571_ = new_n5570_;
  assign new_n5572_ = new_n5571_;
  assign new_n5573_ = new_n5572_;
  assign new_n5574_ = new_n5572_;
  assign new_n5575_ = new_n5571_;
  assign new_n5576_ = new_n5575_;
  assign new_n5577_ = new_n5575_;
  assign new_n5578_ = new_n5570_;
  assign new_n5579_ = new_n5578_;
  assign new_n5580_ = new_n5578_;
  assign new_n5581_ = new_n3617_;
  assign new_n5582_ = new_n5581_;
  assign new_n5583_ = new_n5582_;
  assign new_n5584_ = new_n5583_;
  assign new_n5585_ = new_n5583_;
  assign new_n5586_ = new_n5582_;
  assign new_n5587_ = new_n5586_;
  assign new_n5588_ = new_n5586_;
  assign new_n5589_ = new_n5581_;
  assign new_n5590_ = new_n5589_;
  assign new_n5591_ = new_n5589_;
  assign new_n5592_ = new_n3625_;
  assign new_n5593_ = new_n5592_;
  assign new_n5594_ = new_n1147_;
  assign new_n5595_ = new_n5594_;
  assign new_n5596_ = new_n5594_;
  assign new_n5597_ = new_n1155_;
  assign new_n5598_ = new_n5597_;
  assign new_n5599_ = new_n5597_;
  assign new_n5600_ = new_n3642_;
  assign new_n5601_ = new_n3763_;
  assign new_n5602_ = new_n1145_;
  assign new_n5603_ = new_n5602_;
  assign new_n5604_ = new_n1153_;
  assign new_n5605_ = new_n5604_;
  assign new_n5606_ = new_n3777_;
  assign new_n5607_ = new_n3791_;
  assign new_n5608_ = new_n1131_;
  assign new_n5609_ = new_n3804_;
  always @ (posedge clock) begin
    n1836_lo <= n1836_li;
    n1872_lo <= n1872_li;
    n1884_lo <= n1884_li;
    n1911_lo <= n1911_li;
    n1914_lo <= n1914_li;
    n1917_lo <= n1917_li;
    n1923_lo <= n1923_li;
    n1926_lo <= n1926_li;
    n1929_lo <= n1929_li;
    n1935_lo <= n1935_li;
    n1938_lo <= n1938_li;
    n1947_lo <= n1947_li;
    n1950_lo <= n1950_li;
    n1959_lo <= n1959_li;
    n1962_lo <= n1962_li;
    n1971_lo <= n1971_li;
    n1974_lo <= n1974_li;
    n1983_lo <= n1983_li;
    n1995_lo <= n1995_li;
    n2007_lo <= n2007_li;
    n2019_lo <= n2019_li;
    n2031_lo <= n2031_li;
    n2043_lo <= n2043_li;
    n2055_lo <= n2055_li;
    n2064_lo <= n2064_li;
    n2067_lo <= n2067_li;
    n2100_lo <= n2100_li;
    n2112_lo <= n2112_li;
    n2124_lo <= n2124_li;
    n2136_lo <= n2136_li;
    n2148_lo <= n2148_li;
    n2160_lo <= n2160_li;
    n2163_lo <= n2163_li;
    n2172_lo <= n2172_li;
    n2175_lo <= n2175_li;
    n2184_lo <= n2184_li;
    n2223_lo <= n2223_li;
    n2235_lo <= n2235_li;
    n2238_lo <= n2238_li;
    n2247_lo <= n2247_li;
    n2250_lo <= n2250_li;
    n2259_lo <= n2259_li;
    n2262_lo <= n2262_li;
    n2271_lo <= n2271_li;
    n2274_lo <= n2274_li;
    n2283_lo <= n2283_li;
    n2286_lo <= n2286_li;
    n2295_lo <= n2295_li;
    n2298_lo <= n2298_li;
    n2304_lo <= n2304_li;
    n2307_lo <= n2307_li;
    n2331_lo <= n2331_li;
    n2334_lo <= n2334_li;
    n2337_lo <= n2337_li;
    n2340_lo <= n2340_li;
    n3241_o2 <= n3241_i2;
    n3242_o2 <= n3242_i2;
    n3610_o2 <= n3610_i2;
    n3980_o2 <= n3980_i2;
    n3968_o2 <= n3968_i2;
    n4298_o2 <= n4298_i2;
    n4371_o2 <= n4371_i2;
    n4413_o2 <= n4413_i2;
    n4418_o2 <= n4418_i2;
    n4628_o2 <= n4628_i2;
    n4629_o2 <= n4629_i2;
    n4633_o2 <= n4633_i2;
    n4634_o2 <= n4634_i2;
    n4732_o2 <= n4732_i2;
    n4733_o2 <= n4733_i2;
    n4884_o2 <= n4884_i2;
    n4886_o2 <= n4886_i2;
    n4890_o2 <= n4890_i2;
    n5011_o2 <= n5011_i2;
    n5012_o2 <= n5012_i2;
    n5013_o2 <= n5013_i2;
    n5014_o2 <= n5014_i2;
    n5015_o2 <= n5015_i2;
    n5021_o2 <= n5021_i2;
    n5016_o2 <= n5016_i2;
    n5026_o2 <= n5026_i2;
    n4377_o2 <= n4377_i2;
    n4378_o2 <= n4378_i2;
    n4389_o2 <= n4389_i2;
    n327_inv <= n4390_i2;
    n330_inv <= n4391_i2;
    n4398_o2 <= n4398_i2;
    n4401_o2 <= n4401_i2;
    n5117_o2 <= n5117_i2;
    n5115_o2 <= n5115_i2;
    n5122_o2 <= n5122_i2;
    n5121_o2 <= n5121_i2;
    n5119_o2 <= n5119_i2;
    n5116_o2 <= n5116_i2;
    n5123_o2 <= n5123_i2;
    n5156_o2 <= n5156_i2;
    n5167_o2 <= n5167_i2;
    n4454_o2 <= n4454_i2;
    n4455_o2 <= n4455_i2;
    n4456_o2 <= n4456_i2;
    n4505_o2 <= n4505_i2;
    G742_o2 <= G742_i2;
    G727_o2 <= G727_i2;
    n4567_o2 <= n4567_i2;
    n4568_o2 <= n4568_i2;
    n4569_o2 <= n4569_i2;
    n4571_o2 <= n4571_i2;
    n4572_o2 <= n4572_i2;
    n399_inv <= n4537_i2;
    n4539_o2 <= n4539_i2;
    n4651_o2 <= n4651_i2;
    n4652_o2 <= n4652_i2;
    n4653_o2 <= n4653_i2;
    G1514_o2 <= G1514_i2;
    G1823_o2 <= G1823_i2;
    n4783_o2 <= n4783_i2;
    n4787_o2 <= n4787_i2;
    n426_inv <= n4808_i2;
    n429_inv <= n4815_i2;
    n4816_o2 <= n4816_i2;
    n435_inv <= n4822_i2;
    G572_o2 <= G572_i2;
    n4919_o2 <= n4919_i2;
    n4920_o2 <= n4920_i2;
    n4921_o2 <= n4921_i2;
    G1048_o2 <= G1048_i2;
    n5041_o2 <= n5041_i2;
    n5094_o2 <= n5094_i2;
    n5278_o2 <= n5278_i2;
    n5301_o2 <= n5301_i2;
    G2610_o2 <= G2610_i2;
    G3174_o2 <= G3174_i2;
    G3146_o2 <= G3146_i2;
    G3217_o2 <= G3217_i2;
    G3220_o2 <= G3220_i2;
    G2839_o2 <= G2839_i2;
    G3251_o2 <= G3251_i2;
    G3042_o2 <= G3042_i2;
    G3045_o2 <= G3045_i2;
    G3262_o2 <= G3262_i2;
    G2845_o2 <= G2845_i2;
    G2929_o2 <= G2929_i2;
    G2848_o2 <= G2848_i2;
    G2851_o2 <= G2851_i2;
    G3291_o2 <= G3291_i2;
    G3254_o2 <= G3254_i2;
    G2666_o2 <= G2666_i2;
    n5099_o2 <= n5099_i2;
    n5100_o2 <= n5100_i2;
    n5101_o2 <= n5101_i2;
    G2558_o2 <= G2558_i2;
    n5266_o2 <= n5266_i2;
    n5267_o2 <= n5267_i2;
    G2759_o2 <= G2759_i2;
    n537_inv <= n5269_i2;
    n540_inv <= n5270_i2;
    n543_inv <= n5271_i2;
    n5292_o2 <= n5292_i2;
    n5293_o2 <= n5293_i2;
    n5294_o2 <= n5294_i2;
    n5295_o2 <= n5295_i2;
    G618_o2 <= G618_i2;
    G621_o2 <= G621_i2;
    G384_o2 <= G384_i2;
    G377_o2 <= G377_i2;
    n570_inv <= G400_i2;
    G3171_o2 <= G3171_i2;
    G2552_o2 <= G2552_i2;
    G3272_o2 <= G3272_i2;
    G2015_o2 <= G2015_i2;
    G3294_o2 <= G3294_i2;
    G3281_o2 <= G3281_i2;
    G3320_o2 <= G3320_i2;
    G3275_o2 <= G3275_i2;
    G3140_o2 <= G3140_i2;
    G2836_o2 <= G2836_i2;
    G2926_o2 <= G2926_i2;
    G2842_o2 <= G2842_i2;
    G3302_o2 <= G3302_i2;
    G3288_o2 <= G3288_i2;
    G3143_o2 <= G3143_i2;
    G3100_o2 <= G3100_i2;
    G2512_o2 <= G2512_i2;
    n5325_o2 <= n5325_i2;
    n5326_o2 <= n5326_i2;
    n5327_o2 <= n5327_i2;
    n1857_lo_buf_o2 <= n1857_lo_buf_i2;
    n2097_lo_buf_o2 <= n2097_lo_buf_i2;
    G2669_o2 <= G2669_i2;
    n642_inv <= G552_i2;
    G568_o2 <= G568_i2;
    n648_inv <= G530_i2;
    G565_o2 <= G565_i2;
    G559_o2 <= G559_i2;
    n1821_lo_buf_o2 <= n1821_lo_buf_i2;
    n1905_lo_buf_o2 <= n1905_lo_buf_i2;
    n2133_lo_buf_o2 <= n2133_lo_buf_i2;
    n2145_lo_buf_o2 <= n2145_lo_buf_i2;
    n2157_lo_buf_o2 <= n2157_lo_buf_i2;
    n2205_lo_buf_o2 <= n2205_lo_buf_i2;
    n2217_lo_buf_o2 <= n2217_lo_buf_i2;
    G447_o2 <= G447_i2;
    G434_o2 <= G434_i2;
    G422_o2 <= G422_i2;
    G461_o2 <= G461_i2;
    G3312_o2 <= G3312_i2;
    G3332_o2 <= G3332_i2;
    G3195_o2 <= G3195_i2;
    G2607_o2 <= G2607_i2;
    n702_inv <= G2799_i2;
    G1005_o2 <= G1005_i2;
    G1008_o2 <= G1008_i2;
    n2001_lo_buf_o2 <= n2001_lo_buf_i2;
    n2169_lo_buf_o2 <= n2169_lo_buf_i2;
    n2229_lo_buf_o2 <= n2229_lo_buf_i2;
    n2301_lo_buf_o2 <= n2301_lo_buf_i2;
    n723_inv <= G2816_i2;
    G2947_o2 <= G2947_i2;
    n2013_lo_buf_o2 <= n2013_lo_buf_i2;
    n2025_lo_buf_o2 <= n2025_lo_buf_i2;
    n2037_lo_buf_o2 <= n2037_lo_buf_i2;
    n2049_lo_buf_o2 <= n2049_lo_buf_i2;
    n2181_lo_buf_o2 <= n2181_lo_buf_i2;
    n744_inv <= G546_i2;
    n747_inv <= G480_i2;
    n750_inv <= G492_i2;
    n753_inv <= G540_i2;
    G3350_o2 <= G3350_i2;
    G3360_o2 <= G3360_i2;
    G3373_o2 <= G3373_i2;
    G3237_o2 <= G3237_i2;
    G2773_o2 <= G2773_i2;
    G1733_o2 <= G1733_i2;
    G1738_o2 <= G1738_i2;
    G1751_o2 <= G1751_i2;
    G2216_o2 <= G2216_i2;
    G2219_o2 <= G2219_i2;
    n786_inv <= G381_i2;
    n789_inv <= G397_i2;
    G787_o2 <= G787_i2;
    G2823_o2 <= G2823_i2;
    G2796_o2 <= G2796_i2;
    G875_o2 <= G875_i2;
    G2208_o2 <= G2208_i2;
    G2211_o2 <= G2211_i2;
    n1989_lo_buf_o2 <= n1989_lo_buf_i2;
    n2061_lo_buf_o2 <= n2061_lo_buf_i2;
    n2313_lo_buf_o2 <= n2313_lo_buf_i2;
    G2232_o2 <= G2232_i2;
    G1725_o2 <= G1725_i2;
    G1764_o2 <= G1764_i2;
    G2356_o2 <= G2356_i2;
    G2359_o2 <= G2359_i2;
    G1180_o2 <= G1180_i2;
    G1756_o2 <= G1756_i2;
    G2441_o2 <= G2441_i2;
    G2887_o2 <= G2887_i2;
    G2991_o2 <= G2991_i2;
    n849_inv <= G470_i2;
    n852_inv <= G484_i2;
    n855_inv <= G496_i2;
    n858_inv <= G353_i2;
    n861_inv <= G363_i2;
    G2805_o2 <= G2805_i2;
    G2906_o2 <= G2906_i2;
    G2833_o2 <= G2833_i2;
    n873_inv <= G1012_i2;
    G3353_o2 <= G3353_i2;
    G3367_o2 <= G3367_i2;
    G3346_o2 <= G3346_i2;
    G3340_o2 <= G3340_i2;
    G3376_o2 <= G3376_i2;
    G3359_o2 <= G3359_i2;
    G3240_o2 <= G3240_i2;
    G3344_o2 <= G3344_i2;
    G2880_o2 <= G2880_i2;
    G2939_o2 <= G2939_i2;
    G2248_o2 <= G2248_i2;
    G2251_o2 <= G2251_i2;
    G2021_o2 <= G2021_i2;
    G3383_o2 <= G3383_i2;
    G3399_o2 <= G3399_i2;
    G3404_o2 <= G3404_i2;
    G3265_o2 <= G3265_i2;
    G2866_o2 <= G2866_i2;
    G2999_o2 <= G2999_i2;
    G736_o2 <= G736_i2;
    G739_o2 <= G739_i2;
    G1200_o2 <= G1200_i2;
    G1203_o2 <= G1203_i2;
    G3027_o2 <= G3027_i2;
    G1463_o2 <= G1463_i2;
    G1460_o2 <= G1460_i2;
    G3012_o2 <= G3012_i2;
    G1574_o2 <= G1574_i2;
    G1646_o2 <= G1646_i2;
    G1592_o2 <= G1592_i2;
    G1664_o2 <= G1664_i2;
    G1547_o2 <= G1547_i2;
    G1619_o2 <= G1619_i2;
    G1556_o2 <= G1556_i2;
    G1628_o2 <= G1628_i2;
    G1583_o2 <= G1583_i2;
    G1655_o2 <= G1655_i2;
    G1529_o2 <= G1529_i2;
    G1601_o2 <= G1601_i2;
    G1538_o2 <= G1538_i2;
    G1610_o2 <= G1610_i2;
    G1565_o2 <= G1565_i2;
    G1637_o2 <= G1637_i2;
    G2437_o2 <= G2437_i2;
    n1008_inv <= G2518_i2;
    n1785_lo_buf_o2 <= n1785_lo_buf_i2;
    n1845_lo_buf_o2 <= n1845_lo_buf_i2;
    n1893_lo_buf_o2 <= n1893_lo_buf_i2;
    n1941_lo_buf_o2 <= n1941_lo_buf_i2;
    n1953_lo_buf_o2 <= n1953_lo_buf_i2;
    n1965_lo_buf_o2 <= n1965_lo_buf_i2;
    n1977_lo_buf_o2 <= n1977_lo_buf_i2;
    n2241_lo_buf_o2 <= n2241_lo_buf_i2;
    n2253_lo_buf_o2 <= n2253_lo_buf_i2;
    n2265_lo_buf_o2 <= n2265_lo_buf_i2;
    n2277_lo_buf_o2 <= n2277_lo_buf_i2;
    n2289_lo_buf_o2 <= n2289_lo_buf_i2;
    G519_o2 <= G519_i2;
    n1050_inv <= G388_i2;
    n1053_inv <= G438_i2;
    n1056_inv <= G368_i2;
    G1318_o2 <= G1318_i2;
    n1062_inv <= G425_i2;
    G593_o2 <= G593_i2;
    n1068_inv <= G413_i2;
    n1071_inv <= G404_i2;
    n1074_inv <= G451_i2;
    G2284_o2 <= G2284_i2;
    G2580_o2 <= G2580_i2;
    G2302_o2 <= G2302_i2;
    G2598_o2 <= G2598_i2;
    G2497_o2 <= G2497_i2;
    G2651_o2 <= G2651_i2;
    G2296_o2 <= G2296_i2;
    G2308_o2 <= G2308_i2;
    G2592_o2 <= G2592_i2;
    G2604_o2 <= G2604_i2;
    G2902_o2 <= G2902_i2;
    G2975_o2 <= G2975_i2;
    G2962_o2 <= G2962_i2;
    G3069_o2 <= G3069_i2;
    G2018_o2 <= G2018_i2;
    G1176_o2 <= G1176_i2;
    G1189_o2 <= G1189_i2;
    G3066_o2 <= G3066_i2;
    G3137_o2 <= G3137_i2;
    G3038_o2 <= G3038_i2;
    G3117_o2 <= G3117_i2;
    G2384_o2 <= G2384_i2;
    G2472_o2 <= G2472_i2;
    G772_o2 <= G772_i2;
    G935_o2 <= G935_i2;
    G2923_o2 <= G2923_i2;
    G2971_o2 <= G2971_i2;
    G2980_o2 <= G2980_i2;
    G3039_o2 <= G3039_i2;
    G2388_o2 <= G2388_i2;
    G2287_o2 <= G2287_i2;
    G3024_o2 <= G3024_i2;
    G2916_o2 <= G2916_i2;
    n1176_inv <= G1819_i2;
    G3035_o2 <= G3035_i2;
    G3107_o2 <= G3107_i2;
    G1023_o2 <= G1023_i2;
    G1024_o2 <= G1024_i2;
    G1311_o2 <= G1311_i2;
    G1312_o2 <= G1312_i2;
    G3063_o2 <= G3063_i2;
    G1520_o2 <= G1520_i2;
    G1519_o2 <= G1519_i2;
    G3078_o2 <= G3078_i2;
    G2038_o2 <= G2038_i2;
    G1848_o2 <= G1848_i2;
    G1864_o2 <= G1864_i2;
    G1872_o2 <= G1872_i2;
    G1880_o2 <= G1880_i2;
    G1888_o2 <= G1888_i2;
    G1912_o2 <= G1912_i2;
    G1928_o2 <= G1928_i2;
    G1936_o2 <= G1936_i2;
    G1944_o2 <= G1944_i2;
    G1952_o2 <= G1952_i2;
    G1850_o2 <= G1850_i2;
    G1866_o2 <= G1866_i2;
    G1874_o2 <= G1874_i2;
    G1882_o2 <= G1882_i2;
    G1890_o2 <= G1890_i2;
    G1914_o2 <= G1914_i2;
    G1930_o2 <= G1930_i2;
    G1938_o2 <= G1938_i2;
    G1946_o2 <= G1946_i2;
    G1954_o2 <= G1954_i2;
    G1845_o2 <= G1845_i2;
    G1861_o2 <= G1861_i2;
    G1869_o2 <= G1869_i2;
    G1877_o2 <= G1877_i2;
    G1885_o2 <= G1885_i2;
    G1909_o2 <= G1909_i2;
    G1925_o2 <= G1925_i2;
    G1933_o2 <= G1933_i2;
    G1941_o2 <= G1941_i2;
    G1949_o2 <= G1949_i2;
    G1846_o2 <= G1846_i2;
    G1862_o2 <= G1862_i2;
    G1870_o2 <= G1870_i2;
    G1878_o2 <= G1878_i2;
    G1886_o2 <= G1886_i2;
    G1910_o2 <= G1910_i2;
    G1926_o2 <= G1926_i2;
    G1934_o2 <= G1934_i2;
    G1942_o2 <= G1942_i2;
    G1950_o2 <= G1950_i2;
    G1849_o2 <= G1849_i2;
    G1865_o2 <= G1865_i2;
    G1873_o2 <= G1873_i2;
    G1881_o2 <= G1881_i2;
    G1889_o2 <= G1889_i2;
    G1913_o2 <= G1913_i2;
    G1929_o2 <= G1929_i2;
    G1937_o2 <= G1937_i2;
    G1945_o2 <= G1945_i2;
    G1953_o2 <= G1953_i2;
    G1843_o2 <= G1843_i2;
    G1859_o2 <= G1859_i2;
    G1867_o2 <= G1867_i2;
    G1875_o2 <= G1875_i2;
    G1883_o2 <= G1883_i2;
    G1907_o2 <= G1907_i2;
    G1923_o2 <= G1923_i2;
    G1931_o2 <= G1931_i2;
    G1939_o2 <= G1939_i2;
    G1947_o2 <= G1947_i2;
    G1844_o2 <= G1844_i2;
    G1860_o2 <= G1860_i2;
    G1868_o2 <= G1868_i2;
    G1876_o2 <= G1876_i2;
    G1884_o2 <= G1884_i2;
    G1908_o2 <= G1908_i2;
    G1924_o2 <= G1924_i2;
    G1932_o2 <= G1932_i2;
    G1940_o2 <= G1940_i2;
    G1948_o2 <= G1948_i2;
    G1847_o2 <= G1847_i2;
    G1863_o2 <= G1863_i2;
    G1871_o2 <= G1871_i2;
    G1879_o2 <= G1879_i2;
    G1887_o2 <= G1887_i2;
    G1911_o2 <= G1911_i2;
    G1927_o2 <= G1927_i2;
    G1935_o2 <= G1935_i2;
    G1943_o2 <= G1943_i2;
    G1951_o2 <= G1951_i2;
    G2444_o2 <= G2444_i2;
    G2451_o2 <= G2451_i2;
    G2502_o2 <= G2502_i2;
    G2507_o2 <= G2507_i2;
    n1464_inv <= G2515_i2;
    G2583_o2 <= G2583_i2;
    n1797_lo_buf_o2 <= n1797_lo_buf_i2;
    n1833_lo_buf_o2 <= n1833_lo_buf_i2;
    n1881_lo_buf_o2 <= n1881_lo_buf_i2;
    n1479_inv <= G523_i2;
    n1482_inv <= G575_i2;
    n1485_inv <= G578_i2;
    G615_o2 <= G615_i2;
    G2254_o2 <= G2254_i2;
    G2255_o2 <= G2255_i2;
    G2027_o2 <= G2027_i2;
    G2393_o2 <= G2393_i2;
    G527_o2 <= G527_i2;
    G594_o2 <= G594_i2;
    G1689_o2 <= G1689_i2;
    G1693_o2 <= G1693_i2;
    G2281_o2 <= G2281_i2;
    G2014_o2 <= G2014_i2;
    G2459_o2 <= G2459_i2;
    G2561_o2 <= G2561_i2;
    G2533_o2 <= G2533_i2;
    n1749_lo_buf_o2 <= n1749_lo_buf_i2;
    n1761_lo_buf_o2 <= n1761_lo_buf_i2;
    n1773_lo_buf_o2 <= n1773_lo_buf_i2;
    n1809_lo_buf_o2 <= n1809_lo_buf_i2;
    G1955_o2 <= G1955_i2;
    G1958_o2 <= G1958_i2;
    G2562_o2 <= G2562_i2;
    G2398_o2 <= G2398_i2;
    n1554_inv <= G2524_i2;
    n1557_inv <= G2563_i2;
    G2577_o2 <= G2577_i2;
    G2627_o2 <= G2627_i2;
    G654_o2 <= G654_i2;
    G660_o2 <= G660_i2;
    G831_o2 <= G831_i2;
    G919_o2 <= G919_i2;
    G925_o2 <= G925_i2;
    n1815_lo_buf_o2 <= n1815_lo_buf_i2;
    n1899_lo_buf_o2 <= n1899_lo_buf_i2;
    n2079_lo_buf_o2 <= n2079_lo_buf_i2;
    n2127_lo_buf_o2 <= n2127_lo_buf_i2;
    n2139_lo_buf_o2 <= n2139_lo_buf_i2;
    n2151_lo_buf_o2 <= n2151_lo_buf_i2;
    n2187_lo_buf_o2 <= n2187_lo_buf_i2;
    n2199_lo_buf_o2 <= n2199_lo_buf_i2;
    n2211_lo_buf_o2 <= n2211_lo_buf_i2;
    G533_o2 <= G533_i2;
    n1854_lo_buf_o2 <= n1854_lo_buf_i2;
    n2094_lo_buf_o2 <= n2094_lo_buf_i2;
    G667_o2 <= G667_i2;
    G874_o2 <= G874_i2;
    G851_o2 <= G851_i2;
    G1127_o2 <= G1127_i2;
    n1869_lo_buf_o2 <= n1869_lo_buf_i2;
    n2109_lo_buf_o2 <= n2109_lo_buf_i2;
    n2121_lo_buf_o2 <= n2121_lo_buf_i2;
    G477_o2 <= G477_i2;
    G491_o2 <= G491_i2;
    G501_o2 <= G501_i2;
    G786_o2 <= G786_i2;
    G791_o2 <= G791_i2;
    G1126_o2 <= G1126_i2;
    G1052_o2 <= G1052_i2;
    G1054_o2 <= G1054_i2;
  end
  initial begin
    n1836_lo <= 1'b0;
    n1872_lo <= 1'b0;
    n1884_lo <= 1'b0;
    n1911_lo <= 1'b0;
    n1914_lo <= 1'b0;
    n1917_lo <= 1'b0;
    n1923_lo <= 1'b0;
    n1926_lo <= 1'b0;
    n1929_lo <= 1'b0;
    n1935_lo <= 1'b0;
    n1938_lo <= 1'b0;
    n1947_lo <= 1'b0;
    n1950_lo <= 1'b0;
    n1959_lo <= 1'b0;
    n1962_lo <= 1'b0;
    n1971_lo <= 1'b0;
    n1974_lo <= 1'b0;
    n1983_lo <= 1'b0;
    n1995_lo <= 1'b0;
    n2007_lo <= 1'b0;
    n2019_lo <= 1'b0;
    n2031_lo <= 1'b0;
    n2043_lo <= 1'b0;
    n2055_lo <= 1'b0;
    n2064_lo <= 1'b0;
    n2067_lo <= 1'b0;
    n2100_lo <= 1'b0;
    n2112_lo <= 1'b0;
    n2124_lo <= 1'b0;
    n2136_lo <= 1'b0;
    n2148_lo <= 1'b0;
    n2160_lo <= 1'b0;
    n2163_lo <= 1'b0;
    n2172_lo <= 1'b0;
    n2175_lo <= 1'b0;
    n2184_lo <= 1'b0;
    n2223_lo <= 1'b0;
    n2235_lo <= 1'b0;
    n2238_lo <= 1'b0;
    n2247_lo <= 1'b0;
    n2250_lo <= 1'b0;
    n2259_lo <= 1'b0;
    n2262_lo <= 1'b0;
    n2271_lo <= 1'b0;
    n2274_lo <= 1'b0;
    n2283_lo <= 1'b0;
    n2286_lo <= 1'b0;
    n2295_lo <= 1'b0;
    n2298_lo <= 1'b0;
    n2304_lo <= 1'b0;
    n2307_lo <= 1'b0;
    n2331_lo <= 1'b0;
    n2334_lo <= 1'b0;
    n2337_lo <= 1'b0;
    n2340_lo <= 1'b0;
    n3241_o2 <= 1'b0;
    n3242_o2 <= 1'b0;
    n3610_o2 <= 1'b0;
    n3980_o2 <= 1'b0;
    n3968_o2 <= 1'b0;
    n4298_o2 <= 1'b0;
    n4371_o2 <= 1'b0;
    n4413_o2 <= 1'b0;
    n4418_o2 <= 1'b0;
    n4628_o2 <= 1'b0;
    n4629_o2 <= 1'b0;
    n4633_o2 <= 1'b0;
    n4634_o2 <= 1'b0;
    n4732_o2 <= 1'b0;
    n4733_o2 <= 1'b0;
    n4884_o2 <= 1'b0;
    n4886_o2 <= 1'b0;
    n4890_o2 <= 1'b0;
    n5011_o2 <= 1'b0;
    n5012_o2 <= 1'b0;
    n5013_o2 <= 1'b0;
    n5014_o2 <= 1'b0;
    n5015_o2 <= 1'b0;
    n5021_o2 <= 1'b0;
    n5016_o2 <= 1'b0;
    n5026_o2 <= 1'b0;
    n4377_o2 <= 1'b0;
    n4378_o2 <= 1'b0;
    n4389_o2 <= 1'b0;
    n327_inv <= 1'b0;
    n330_inv <= 1'b0;
    n4398_o2 <= 1'b0;
    n4401_o2 <= 1'b0;
    n5117_o2 <= 1'b0;
    n5115_o2 <= 1'b0;
    n5122_o2 <= 1'b0;
    n5121_o2 <= 1'b0;
    n5119_o2 <= 1'b0;
    n5116_o2 <= 1'b0;
    n5123_o2 <= 1'b0;
    n5156_o2 <= 1'b0;
    n5167_o2 <= 1'b0;
    n4454_o2 <= 1'b0;
    n4455_o2 <= 1'b0;
    n4456_o2 <= 1'b0;
    n4505_o2 <= 1'b0;
    G742_o2 <= 1'b0;
    G727_o2 <= 1'b0;
    n4567_o2 <= 1'b0;
    n4568_o2 <= 1'b0;
    n4569_o2 <= 1'b0;
    n4571_o2 <= 1'b0;
    n4572_o2 <= 1'b0;
    n399_inv <= 1'b0;
    n4539_o2 <= 1'b0;
    n4651_o2 <= 1'b0;
    n4652_o2 <= 1'b0;
    n4653_o2 <= 1'b0;
    G1514_o2 <= 1'b0;
    G1823_o2 <= 1'b0;
    n4783_o2 <= 1'b0;
    n4787_o2 <= 1'b0;
    n426_inv <= 1'b0;
    n429_inv <= 1'b0;
    n4816_o2 <= 1'b0;
    n435_inv <= 1'b0;
    G572_o2 <= 1'b0;
    n4919_o2 <= 1'b0;
    n4920_o2 <= 1'b0;
    n4921_o2 <= 1'b0;
    G1048_o2 <= 1'b0;
    n5041_o2 <= 1'b0;
    n5094_o2 <= 1'b0;
    n5278_o2 <= 1'b0;
    n5301_o2 <= 1'b0;
    G2610_o2 <= 1'b0;
    G3174_o2 <= 1'b0;
    G3146_o2 <= 1'b0;
    G3217_o2 <= 1'b0;
    G3220_o2 <= 1'b0;
    G2839_o2 <= 1'b0;
    G3251_o2 <= 1'b0;
    G3042_o2 <= 1'b0;
    G3045_o2 <= 1'b0;
    G3262_o2 <= 1'b0;
    G2845_o2 <= 1'b0;
    G2929_o2 <= 1'b0;
    G2848_o2 <= 1'b0;
    G2851_o2 <= 1'b0;
    G3291_o2 <= 1'b0;
    G3254_o2 <= 1'b0;
    G2666_o2 <= 1'b0;
    n5099_o2 <= 1'b0;
    n5100_o2 <= 1'b0;
    n5101_o2 <= 1'b0;
    G2558_o2 <= 1'b0;
    n5266_o2 <= 1'b0;
    n5267_o2 <= 1'b0;
    G2759_o2 <= 1'b0;
    n537_inv <= 1'b0;
    n540_inv <= 1'b0;
    n543_inv <= 1'b0;
    n5292_o2 <= 1'b0;
    n5293_o2 <= 1'b0;
    n5294_o2 <= 1'b0;
    n5295_o2 <= 1'b0;
    G618_o2 <= 1'b0;
    G621_o2 <= 1'b0;
    G384_o2 <= 1'b0;
    G377_o2 <= 1'b0;
    n570_inv <= 1'b0;
    G3171_o2 <= 1'b0;
    G2552_o2 <= 1'b0;
    G3272_o2 <= 1'b0;
    G2015_o2 <= 1'b0;
    G3294_o2 <= 1'b0;
    G3281_o2 <= 1'b0;
    G3320_o2 <= 1'b0;
    G3275_o2 <= 1'b0;
    G3140_o2 <= 1'b0;
    G2836_o2 <= 1'b0;
    G2926_o2 <= 1'b0;
    G2842_o2 <= 1'b0;
    G3302_o2 <= 1'b0;
    G3288_o2 <= 1'b0;
    G3143_o2 <= 1'b0;
    G3100_o2 <= 1'b0;
    G2512_o2 <= 1'b0;
    n5325_o2 <= 1'b0;
    n5326_o2 <= 1'b0;
    n5327_o2 <= 1'b0;
    n1857_lo_buf_o2 <= 1'b0;
    n2097_lo_buf_o2 <= 1'b0;
    G2669_o2 <= 1'b0;
    n642_inv <= 1'b0;
    G568_o2 <= 1'b0;
    n648_inv <= 1'b0;
    G565_o2 <= 1'b0;
    G559_o2 <= 1'b0;
    n1821_lo_buf_o2 <= 1'b0;
    n1905_lo_buf_o2 <= 1'b0;
    n2133_lo_buf_o2 <= 1'b0;
    n2145_lo_buf_o2 <= 1'b0;
    n2157_lo_buf_o2 <= 1'b0;
    n2205_lo_buf_o2 <= 1'b0;
    n2217_lo_buf_o2 <= 1'b0;
    G447_o2 <= 1'b0;
    G434_o2 <= 1'b0;
    G422_o2 <= 1'b0;
    G461_o2 <= 1'b0;
    G3312_o2 <= 1'b0;
    G3332_o2 <= 1'b0;
    G3195_o2 <= 1'b0;
    G2607_o2 <= 1'b0;
    n702_inv <= 1'b0;
    G1005_o2 <= 1'b0;
    G1008_o2 <= 1'b0;
    n2001_lo_buf_o2 <= 1'b0;
    n2169_lo_buf_o2 <= 1'b0;
    n2229_lo_buf_o2 <= 1'b0;
    n2301_lo_buf_o2 <= 1'b0;
    n723_inv <= 1'b0;
    G2947_o2 <= 1'b0;
    n2013_lo_buf_o2 <= 1'b0;
    n2025_lo_buf_o2 <= 1'b0;
    n2037_lo_buf_o2 <= 1'b0;
    n2049_lo_buf_o2 <= 1'b0;
    n2181_lo_buf_o2 <= 1'b0;
    n744_inv <= 1'b0;
    n747_inv <= 1'b0;
    n750_inv <= 1'b0;
    n753_inv <= 1'b0;
    G3350_o2 <= 1'b0;
    G3360_o2 <= 1'b0;
    G3373_o2 <= 1'b0;
    G3237_o2 <= 1'b0;
    G2773_o2 <= 1'b0;
    G1733_o2 <= 1'b0;
    G1738_o2 <= 1'b0;
    G1751_o2 <= 1'b0;
    G2216_o2 <= 1'b0;
    G2219_o2 <= 1'b0;
    n786_inv <= 1'b0;
    n789_inv <= 1'b0;
    G787_o2 <= 1'b0;
    G2823_o2 <= 1'b0;
    G2796_o2 <= 1'b0;
    G875_o2 <= 1'b0;
    G2208_o2 <= 1'b0;
    G2211_o2 <= 1'b0;
    n1989_lo_buf_o2 <= 1'b0;
    n2061_lo_buf_o2 <= 1'b0;
    n2313_lo_buf_o2 <= 1'b0;
    G2232_o2 <= 1'b0;
    G1725_o2 <= 1'b0;
    G1764_o2 <= 1'b0;
    G2356_o2 <= 1'b0;
    G2359_o2 <= 1'b0;
    G1180_o2 <= 1'b0;
    G1756_o2 <= 1'b0;
    G2441_o2 <= 1'b0;
    G2887_o2 <= 1'b0;
    G2991_o2 <= 1'b0;
    n849_inv <= 1'b0;
    n852_inv <= 1'b0;
    n855_inv <= 1'b0;
    n858_inv <= 1'b0;
    n861_inv <= 1'b0;
    G2805_o2 <= 1'b0;
    G2906_o2 <= 1'b0;
    G2833_o2 <= 1'b0;
    n873_inv <= 1'b0;
    G3353_o2 <= 1'b0;
    G3367_o2 <= 1'b0;
    G3346_o2 <= 1'b0;
    G3340_o2 <= 1'b0;
    G3376_o2 <= 1'b0;
    G3359_o2 <= 1'b0;
    G3240_o2 <= 1'b0;
    G3344_o2 <= 1'b0;
    G2880_o2 <= 1'b0;
    G2939_o2 <= 1'b0;
    G2248_o2 <= 1'b0;
    G2251_o2 <= 1'b0;
    G2021_o2 <= 1'b0;
    G3383_o2 <= 1'b0;
    G3399_o2 <= 1'b0;
    G3404_o2 <= 1'b0;
    G3265_o2 <= 1'b0;
    G2866_o2 <= 1'b0;
    G2999_o2 <= 1'b0;
    G736_o2 <= 1'b0;
    G739_o2 <= 1'b0;
    G1200_o2 <= 1'b0;
    G1203_o2 <= 1'b0;
    G3027_o2 <= 1'b0;
    G1463_o2 <= 1'b0;
    G1460_o2 <= 1'b0;
    G3012_o2 <= 1'b0;
    G1574_o2 <= 1'b0;
    G1646_o2 <= 1'b0;
    G1592_o2 <= 1'b0;
    G1664_o2 <= 1'b0;
    G1547_o2 <= 1'b0;
    G1619_o2 <= 1'b0;
    G1556_o2 <= 1'b0;
    G1628_o2 <= 1'b0;
    G1583_o2 <= 1'b0;
    G1655_o2 <= 1'b0;
    G1529_o2 <= 1'b0;
    G1601_o2 <= 1'b0;
    G1538_o2 <= 1'b0;
    G1610_o2 <= 1'b0;
    G1565_o2 <= 1'b0;
    G1637_o2 <= 1'b0;
    G2437_o2 <= 1'b0;
    n1008_inv <= 1'b0;
    n1785_lo_buf_o2 <= 1'b0;
    n1845_lo_buf_o2 <= 1'b0;
    n1893_lo_buf_o2 <= 1'b0;
    n1941_lo_buf_o2 <= 1'b0;
    n1953_lo_buf_o2 <= 1'b0;
    n1965_lo_buf_o2 <= 1'b0;
    n1977_lo_buf_o2 <= 1'b0;
    n2241_lo_buf_o2 <= 1'b0;
    n2253_lo_buf_o2 <= 1'b0;
    n2265_lo_buf_o2 <= 1'b0;
    n2277_lo_buf_o2 <= 1'b0;
    n2289_lo_buf_o2 <= 1'b0;
    G519_o2 <= 1'b0;
    n1050_inv <= 1'b0;
    n1053_inv <= 1'b0;
    n1056_inv <= 1'b0;
    G1318_o2 <= 1'b0;
    n1062_inv <= 1'b0;
    G593_o2 <= 1'b0;
    n1068_inv <= 1'b0;
    n1071_inv <= 1'b0;
    n1074_inv <= 1'b0;
    G2284_o2 <= 1'b0;
    G2580_o2 <= 1'b0;
    G2302_o2 <= 1'b0;
    G2598_o2 <= 1'b0;
    G2497_o2 <= 1'b0;
    G2651_o2 <= 1'b0;
    G2296_o2 <= 1'b0;
    G2308_o2 <= 1'b0;
    G2592_o2 <= 1'b0;
    G2604_o2 <= 1'b0;
    G2902_o2 <= 1'b0;
    G2975_o2 <= 1'b0;
    G2962_o2 <= 1'b0;
    G3069_o2 <= 1'b0;
    G2018_o2 <= 1'b0;
    G1176_o2 <= 1'b0;
    G1189_o2 <= 1'b0;
    G3066_o2 <= 1'b0;
    G3137_o2 <= 1'b0;
    G3038_o2 <= 1'b0;
    G3117_o2 <= 1'b0;
    G2384_o2 <= 1'b0;
    G2472_o2 <= 1'b0;
    G772_o2 <= 1'b0;
    G935_o2 <= 1'b0;
    G2923_o2 <= 1'b0;
    G2971_o2 <= 1'b0;
    G2980_o2 <= 1'b0;
    G3039_o2 <= 1'b0;
    G2388_o2 <= 1'b0;
    G2287_o2 <= 1'b0;
    G3024_o2 <= 1'b0;
    G2916_o2 <= 1'b0;
    n1176_inv <= 1'b0;
    G3035_o2 <= 1'b0;
    G3107_o2 <= 1'b0;
    G1023_o2 <= 1'b0;
    G1024_o2 <= 1'b0;
    G1311_o2 <= 1'b0;
    G1312_o2 <= 1'b0;
    G3063_o2 <= 1'b0;
    G1520_o2 <= 1'b0;
    G1519_o2 <= 1'b0;
    G3078_o2 <= 1'b0;
    G2038_o2 <= 1'b0;
    G1848_o2 <= 1'b0;
    G1864_o2 <= 1'b0;
    G1872_o2 <= 1'b0;
    G1880_o2 <= 1'b0;
    G1888_o2 <= 1'b0;
    G1912_o2 <= 1'b0;
    G1928_o2 <= 1'b0;
    G1936_o2 <= 1'b0;
    G1944_o2 <= 1'b0;
    G1952_o2 <= 1'b0;
    G1850_o2 <= 1'b0;
    G1866_o2 <= 1'b0;
    G1874_o2 <= 1'b0;
    G1882_o2 <= 1'b0;
    G1890_o2 <= 1'b0;
    G1914_o2 <= 1'b0;
    G1930_o2 <= 1'b0;
    G1938_o2 <= 1'b0;
    G1946_o2 <= 1'b0;
    G1954_o2 <= 1'b0;
    G1845_o2 <= 1'b0;
    G1861_o2 <= 1'b0;
    G1869_o2 <= 1'b0;
    G1877_o2 <= 1'b0;
    G1885_o2 <= 1'b0;
    G1909_o2 <= 1'b0;
    G1925_o2 <= 1'b0;
    G1933_o2 <= 1'b0;
    G1941_o2 <= 1'b0;
    G1949_o2 <= 1'b0;
    G1846_o2 <= 1'b0;
    G1862_o2 <= 1'b0;
    G1870_o2 <= 1'b0;
    G1878_o2 <= 1'b0;
    G1886_o2 <= 1'b0;
    G1910_o2 <= 1'b0;
    G1926_o2 <= 1'b0;
    G1934_o2 <= 1'b0;
    G1942_o2 <= 1'b0;
    G1950_o2 <= 1'b0;
    G1849_o2 <= 1'b0;
    G1865_o2 <= 1'b0;
    G1873_o2 <= 1'b0;
    G1881_o2 <= 1'b0;
    G1889_o2 <= 1'b0;
    G1913_o2 <= 1'b0;
    G1929_o2 <= 1'b0;
    G1937_o2 <= 1'b0;
    G1945_o2 <= 1'b0;
    G1953_o2 <= 1'b0;
    G1843_o2 <= 1'b0;
    G1859_o2 <= 1'b0;
    G1867_o2 <= 1'b0;
    G1875_o2 <= 1'b0;
    G1883_o2 <= 1'b0;
    G1907_o2 <= 1'b0;
    G1923_o2 <= 1'b0;
    G1931_o2 <= 1'b0;
    G1939_o2 <= 1'b0;
    G1947_o2 <= 1'b0;
    G1844_o2 <= 1'b0;
    G1860_o2 <= 1'b0;
    G1868_o2 <= 1'b0;
    G1876_o2 <= 1'b0;
    G1884_o2 <= 1'b0;
    G1908_o2 <= 1'b0;
    G1924_o2 <= 1'b0;
    G1932_o2 <= 1'b0;
    G1940_o2 <= 1'b0;
    G1948_o2 <= 1'b0;
    G1847_o2 <= 1'b0;
    G1863_o2 <= 1'b0;
    G1871_o2 <= 1'b0;
    G1879_o2 <= 1'b0;
    G1887_o2 <= 1'b0;
    G1911_o2 <= 1'b0;
    G1927_o2 <= 1'b0;
    G1935_o2 <= 1'b0;
    G1943_o2 <= 1'b0;
    G1951_o2 <= 1'b0;
    G2444_o2 <= 1'b0;
    G2451_o2 <= 1'b0;
    G2502_o2 <= 1'b0;
    G2507_o2 <= 1'b0;
    n1464_inv <= 1'b0;
    G2583_o2 <= 1'b0;
    n1797_lo_buf_o2 <= 1'b0;
    n1833_lo_buf_o2 <= 1'b0;
    n1881_lo_buf_o2 <= 1'b0;
    n1479_inv <= 1'b0;
    n1482_inv <= 1'b0;
    n1485_inv <= 1'b0;
    G615_o2 <= 1'b0;
    G2254_o2 <= 1'b0;
    G2255_o2 <= 1'b0;
    G2027_o2 <= 1'b0;
    G2393_o2 <= 1'b0;
    G527_o2 <= 1'b0;
    G594_o2 <= 1'b0;
    G1689_o2 <= 1'b0;
    G1693_o2 <= 1'b0;
    G2281_o2 <= 1'b0;
    G2014_o2 <= 1'b0;
    G2459_o2 <= 1'b0;
    G2561_o2 <= 1'b0;
    G2533_o2 <= 1'b0;
    n1749_lo_buf_o2 <= 1'b0;
    n1761_lo_buf_o2 <= 1'b0;
    n1773_lo_buf_o2 <= 1'b0;
    n1809_lo_buf_o2 <= 1'b0;
    G1955_o2 <= 1'b0;
    G1958_o2 <= 1'b0;
    G2562_o2 <= 1'b0;
    G2398_o2 <= 1'b0;
    n1554_inv <= 1'b0;
    n1557_inv <= 1'b0;
    G2577_o2 <= 1'b0;
    G2627_o2 <= 1'b0;
    G654_o2 <= 1'b0;
    G660_o2 <= 1'b0;
    G831_o2 <= 1'b0;
    G919_o2 <= 1'b0;
    G925_o2 <= 1'b0;
    n1815_lo_buf_o2 <= 1'b0;
    n1899_lo_buf_o2 <= 1'b0;
    n2079_lo_buf_o2 <= 1'b0;
    n2127_lo_buf_o2 <= 1'b0;
    n2139_lo_buf_o2 <= 1'b0;
    n2151_lo_buf_o2 <= 1'b0;
    n2187_lo_buf_o2 <= 1'b0;
    n2199_lo_buf_o2 <= 1'b0;
    n2211_lo_buf_o2 <= 1'b0;
    G533_o2 <= 1'b0;
    n1854_lo_buf_o2 <= 1'b0;
    n2094_lo_buf_o2 <= 1'b0;
    G667_o2 <= 1'b0;
    G874_o2 <= 1'b0;
    G851_o2 <= 1'b0;
    G1127_o2 <= 1'b0;
    n1869_lo_buf_o2 <= 1'b0;
    n2109_lo_buf_o2 <= 1'b0;
    n2121_lo_buf_o2 <= 1'b0;
    G477_o2 <= 1'b0;
    G491_o2 <= 1'b0;
    G501_o2 <= 1'b0;
    G786_o2 <= 1'b0;
    G791_o2 <= 1'b0;
    G1126_o2 <= 1'b0;
    G1052_o2 <= 1'b0;
    G1054_o2 <= 1'b0;
  end
endmodule


