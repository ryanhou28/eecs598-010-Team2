
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  G42,
  G43,
  G44,
  G45,
  G46,
  G47,
  G48,
  G49,
  G50,
  n1752_lo,
  n1776_lo,
  n1824_lo,
  n1836_lo,
  n1848_lo,
  n1860_lo,
  n1872_lo,
  n1884_lo,
  n1896_lo,
  n1908_lo,
  n1911_lo,
  n1914_lo,
  n1923_lo,
  n1926_lo,
  n1935_lo,
  n1938_lo,
  n1947_lo,
  n1950_lo,
  n1959_lo,
  n1962_lo,
  n1971_lo,
  n1974_lo,
  n1983_lo,
  n1995_lo,
  n2055_lo,
  n2064_lo,
  n2067_lo,
  n2079_lo,
  n2100_lo,
  n2112_lo,
  n2124_lo,
  n2136_lo,
  n2148_lo,
  n2160_lo,
  n2172_lo,
  n2184_lo,
  n2235_lo,
  n2238_lo,
  n2247_lo,
  n2250_lo,
  n2259_lo,
  n2262_lo,
  n2271_lo,
  n2274_lo,
  n2283_lo,
  n2286_lo,
  n2289_lo,
  n2295_lo,
  n2298_lo,
  n2304_lo,
  n2307_lo,
  n2316_lo,
  n2331_lo,
  n2334_lo,
  n2337_lo,
  n2340_lo,
  n2071_o2,
  n2080_o2,
  n2137_o2,
  n2368_o2,
  n2383_o2,
  n2405_o2,
  n2471_o2,
  n2617_o2,
  n2765_o2,
  n2775_o2,
  n2829_o2,
  n2579_o2,
  n2580_o2,
  n2618_o2,
  n2619_o2,
  n2620_o2,
  n2621_o2,
  n2622_o2,
  n2623_o2,
  n2624_o2,
  n2625_o2,
  n2626_o2,
  n2627_o2,
  n3029_o2,
  n3035_o2,
  n2643_o2,
  n2644_o2,
  n2645_o2,
  n327_inv,
  n2658_o2,
  n2659_o2,
  n2674_o2,
  n2675_o2,
  n2676_o2,
  n3119_o2,
  n3153_o2,
  n351_inv,
  n2729_o2,
  n2730_o2,
  n2731_o2,
  n698_o2,
  n366_inv,
  n2757_o2,
  n2758_o2,
  n1000_o2,
  n1160_o2,
  n1153_o2,
  n2793_o2,
  n2794_o2,
  n2795_o2,
  n1001_o2,
  n2859_o2,
  n744_o2,
  n402_inv,
  n2926_o2,
  n408_inv,
  n2966_o2,
  n2967_o2,
  n2947_o2,
  n1010_o2,
  n2976_o2,
  n3069_o2,
  n3028_o2,
  n3081_o2,
  n3082_o2,
  n3142_o2,
  n3214_o2,
  n2992_o2,
  n2993_o2,
  n870_o2,
  n3086_o2,
  n3087_o2,
  n3088_o2,
  n3089_o2,
  n3090_o2,
  n3091_o2,
  n3092_o2,
  n3093_o2,
  n3094_o2,
  n3095_o2,
  n483_inv,
  n3170_o2,
  n3171_o2,
  n3172_o2,
  n3179_o2,
  n498_inv,
  n3193_o2,
  n3211_o2,
  n3212_o2,
  n3213_o2,
  n513_inv,
  n1125_o2,
  n1081_o2,
  n1139_o2,
  n3245_o2,
  n3246_o2,
  n3247_o2,
  lo074_buf_o2,
  lo078_buf_o2,
  lo186_buf_o2,
  lo118_buf_o2,
  lo146_buf_o2,
  n1038_o2,
  n1044_o2,
  n555_inv,
  n558_inv,
  lo026_buf_o2,
  lo030_buf_o2,
  lo090_buf_o2,
  lo094_buf_o2,
  lo098_buf_o2,
  lo102_buf_o2,
  lo066_buf_o2,
  lo070_buf_o2,
  n1202_o2,
  n1003_o2,
  n1031_o2,
  n1034_o2,
  n1040_o2,
  n1046_o2,
  n1380_o2,
  n1425_o2,
  n697_o2,
  n1143_o2,
  n673_o2,
  n789_o2,
  n786_o2,
  n1047_o2,
  n1036_o2,
  n1307_o2,
  n1035_o2,
  n1297_o2,
  n1099_o2,
  n1128_o2,
  n645_inv,
  n826_o2,
  n853_o2,
  n654_inv,
  n700_o2,
  n884_o2,
  lo082_buf_o2,
  lo086_buf_o2,
  n801_o2,
  n840_o2,
  n675_inv,
  lo002_buf_o2,
  lo010_buf_o2,
  lo166_buf_o2,
  lo170_buf_o2,
  n1426_o2,
  n1082_o2,
  n1310_o2,
  n1015_o2,
  n1206_o2,
  n1262_o2,
  n1456_o2,
  n1244_o2,
  n1280_o2,
  n1290_o2,
  n1012_o2,
  n1074_o2,
  n1112_o2,
  n1212_o2,
  n1454_o2,
  n1182_o2,
  n1220_o2,
  n701_o2,
  n744_inv,
  n1282_o2,
  n1144_o2,
  n1278_o2,
  n1459_o2,
  n1324_o2,
  n1288_o2,
  n1271_o2,
  n1132_o2,
  n1231_o2,
  n1462_o2,
  n1482_o2,
  n994_o2,
  n998_o2,
  lo106_buf_o2,
  n769_o2,
  n814_o2,
  n841_o2,
  n867_o2,
  lo006_buf_o2,
  lo014_buf_o2,
  lo022_buf_o2,
  lo042_buf_o2,
  lo046_buf_o2,
  lo050_buf_o2,
  lo054_buf_o2,
  lo130_buf_o2,
  lo134_buf_o2,
  lo154_buf_o2,
  lo174_buf_o2,
  lo178_buf_o2,
  n1007_o2,
  n1294_o2,
  n1084_o2,
  n1399_o2,
  n1311_o2,
  n1392_o2,
  n1102_o2,
  n1041_o2,
  n1298_o2,
  n738_o2,
  n1214_o2,
  n1222_o2,
  n1155_o2,
  n1147_o2,
  n1393_o2,
  n999_o2,
  n1306_o2,
  n1312_o2,
  n1382_o2,
  n1383_o2,
  n1152_o2,
  n1334_o2,
  n1335_o2,
  n906_inv,
  n773_o2,
  lo190_buf_o2,
  n1368_o2,
  n1362_o2,
  n1406_o2,
  n1403_o2,
  n741_o2,
  n1407_o2,
  n1395_o2,
  n1359_o2,
  n1159_o2,
  n1221_o2,
  n945_inv,
  n989_o2,
  n881_o2,
  n1340_o2,
  n1341_o2,
  n906_o2,
  n1388_o2,
  n791_o2,
  n1372_o2,
  n815_o2,
  n868_o2,
  lo018_buf_o2,
  lo138_buf_o2,
  lo158_buf_o2,
  n780_o2,
  n728_o2,
  n993_inv,
  n929_o2,
  n955_o2,
  n938_o2,
  n1117_o2,
  n1121_o2,
  n965_o2,
  n752_o2,
  n753_o2,
  n760_o2,
  n770_o2,
  n923_o2,
  n947_o2,
  n897_o2,
  n919_o2,
  n895_o2,
  n917_o2,
  n751_o2,
  n774_o2,
  lo126_buf_o2,
  lo142_buf_o2,
  lo162_buf_o2,
  n1059_inv,
  n792_o2,
  n869_o2,
  n1068_inv,
  lo024_buf_o2,
  lo028_buf_o2,
  lo088_buf_o2,
  lo092_buf_o2,
  lo096_buf_o2,
  lo100_buf_o2,
  n763_o2,
  n754_o2,
  n755_o2,
  n822_o2,
  n849_o2,
  n777_o2,
  n778_o2,
  n820_o2,
  n846_o2,
  n806_o2,
  n771_o2,
  n854_o2,
  n828_o2,
  lo117_buf_o2,
  lo145_buf_o2,
  n762_o2,
  n805_o2,
  n859_o2,
  n833_o2,
  lo034_buf_o2,
  lo038_buf_o2,
  lo122_buf_o2,
  lo150_buf_o2,
  G3519,
  G3520,
  G3521,
  G3522,
  G3523,
  G3524,
  G3525,
  G3526,
  G3527,
  G3528,
  G3529,
  G3530,
  G3531,
  G3532,
  G3533,
  G3534,
  G3535,
  G3536,
  G3537,
  G3538,
  G3539,
  G3540,
  n4070_li003_li003,
  n4094_li011_li011,
  n4142_li027_li027,
  n4154_li031_li031,
  n4166_li035_li035,
  n4178_li039_li039,
  n4190_li043_li043,
  n4202_li047_li047,
  n4214_li051_li051,
  n4226_li055_li055,
  n4229_li056_li056,
  n4232_li057_li057,
  n4241_li060_li060,
  n4244_li061_li061,
  n4253_li064_li064,
  n4256_li065_li065,
  n4265_li068_li068,
  n4268_li069_li069,
  n4277_li072_li072,
  n4280_li073_li073,
  n4289_li076_li076,
  n4292_li077_li077,
  n4301_li080_li080,
  n4313_li084_li084,
  n4373_li104_li104,
  n4382_li107_li107,
  n4385_li108_li108,
  n4397_li112_li112,
  n4418_li119_li119,
  n4430_li123_li123,
  n4442_li127_li127,
  n4454_li131_li131,
  n4466_li135_li135,
  n4478_li139_li139,
  n4490_li143_li143,
  n4502_li147_li147,
  n4553_li164_li164,
  n4556_li165_li165,
  n4565_li168_li168,
  n4568_li169_li169,
  n4577_li172_li172,
  n4580_li173_li173,
  n4589_li176_li176,
  n4592_li177_li177,
  n4601_li180_li180,
  n4604_li181_li181,
  n4607_li182_li182,
  n4613_li184_li184,
  n4616_li185_li185,
  n4622_li187_li187,
  n4625_li188_li188,
  n4634_li191_li191,
  n4649_li196_li196,
  n4652_li197_li197,
  n4655_li198_li198,
  n4658_li199_li199,
  n2071_i2,
  n2080_i2,
  n2137_i2,
  n2368_i2,
  n2383_i2,
  n2405_i2,
  n2471_i2,
  n2617_i2,
  n2765_i2,
  n2775_i2,
  n2829_i2,
  n2579_i2,
  n2580_i2,
  n2618_i2,
  n2619_i2,
  n2620_i2,
  n2621_i2,
  n2622_i2,
  n2623_i2,
  n2624_i2,
  n2625_i2,
  n2626_i2,
  n2627_i2,
  n3029_i2,
  n3035_i2,
  n2643_i2,
  n2644_i2,
  n2645_i2,
  n2640_i2,
  n2658_i2,
  n2659_i2,
  n2674_i2,
  n2675_i2,
  n2676_i2,
  n3119_i2,
  n3153_i2,
  n2681_i2,
  n2729_i2,
  n2730_i2,
  n2731_i2,
  n698_i2,
  n677_i2,
  n2757_i2,
  n2758_i2,
  n1000_i2,
  n1160_i2,
  n1153_i2,
  n2793_i2,
  n2794_i2,
  n2795_i2,
  n1001_i2,
  n2859_i2,
  n744_i2,
  n2908_i2,
  n2926_i2,
  n2928_i2,
  n2966_i2,
  n2967_i2,
  n2947_i2,
  n1010_i2,
  n2976_i2,
  n3069_i2,
  n3028_i2,
  n3081_i2,
  n3082_i2,
  n3142_i2,
  n3214_i2,
  n2992_i2,
  n2993_i2,
  n870_i2,
  n3086_i2,
  n3087_i2,
  n3088_i2,
  n3089_i2,
  n3090_i2,
  n3091_i2,
  n3092_i2,
  n3093_i2,
  n3094_i2,
  n3095_i2,
  n3136_i2,
  n3170_i2,
  n3171_i2,
  n3172_i2,
  n3179_i2,
  n3180_i2,
  n3193_i2,
  n3211_i2,
  n3212_i2,
  n3213_i2,
  n3219_i2,
  n1125_i2,
  n1081_i2,
  n1139_i2,
  n3245_i2,
  n3246_i2,
  n3247_i2,
  lo074_buf_i2,
  lo078_buf_i2,
  lo186_buf_i2,
  lo118_buf_i2,
  lo146_buf_i2,
  n1038_i2,
  n1044_i2,
  n980_i2,
  n1145_i2,
  lo026_buf_i2,
  lo030_buf_i2,
  lo090_buf_i2,
  lo094_buf_i2,
  lo098_buf_i2,
  lo102_buf_i2,
  lo066_buf_i2,
  lo070_buf_i2,
  n1202_i2,
  n1003_i2,
  n1031_i2,
  n1034_i2,
  n1040_i2,
  n1046_i2,
  n1380_i2,
  n1425_i2,
  n697_i2,
  n1143_i2,
  n673_i2,
  n789_i2,
  n786_i2,
  n1047_i2,
  n1036_i2,
  n1307_i2,
  n1035_i2,
  n1297_i2,
  n1099_i2,
  n1128_i2,
  n674_i2,
  n826_i2,
  n853_i2,
  n951_i2,
  n700_i2,
  n884_i2,
  lo082_buf_i2,
  lo086_buf_i2,
  n801_i2,
  n840_i2,
  n866_i2,
  lo002_buf_i2,
  lo010_buf_i2,
  lo166_buf_i2,
  lo170_buf_i2,
  n1426_i2,
  n1082_i2,
  n1310_i2,
  n1015_i2,
  n1206_i2,
  n1262_i2,
  n1456_i2,
  n1244_i2,
  n1280_i2,
  n1290_i2,
  n1012_i2,
  n1074_i2,
  n1112_i2,
  n1212_i2,
  n1454_i2,
  n1182_i2,
  n1220_i2,
  n701_i2,
  n973_i2,
  n1282_i2,
  n1144_i2,
  n1278_i2,
  n1459_i2,
  n1324_i2,
  n1288_i2,
  n1271_i2,
  n1132_i2,
  n1231_i2,
  n1462_i2,
  n1482_i2,
  n994_i2,
  n998_i2,
  lo106_buf_i2,
  n769_i2,
  n814_i2,
  n841_i2,
  n867_i2,
  lo006_buf_i2,
  lo014_buf_i2,
  lo022_buf_i2,
  lo042_buf_i2,
  lo046_buf_i2,
  lo050_buf_i2,
  lo054_buf_i2,
  lo130_buf_i2,
  lo134_buf_i2,
  lo154_buf_i2,
  lo174_buf_i2,
  lo178_buf_i2,
  n1007_i2,
  n1294_i2,
  n1084_i2,
  n1399_i2,
  n1311_i2,
  n1392_i2,
  n1102_i2,
  n1041_i2,
  n1298_i2,
  n738_i2,
  n1214_i2,
  n1222_i2,
  n1155_i2,
  n1147_i2,
  n1393_i2,
  n999_i2,
  n1306_i2,
  n1312_i2,
  n1382_i2,
  n1383_i2,
  n1152_i2,
  n1334_i2,
  n1335_i2,
  n695_i2,
  n773_i2,
  lo190_buf_i2,
  n1368_i2,
  n1362_i2,
  n1406_i2,
  n1403_i2,
  n741_i2,
  n1407_i2,
  n1395_i2,
  n1359_i2,
  n1159_i2,
  n1221_i2,
  n987_i2,
  n989_i2,
  n881_i2,
  n1340_i2,
  n1341_i2,
  n906_i2,
  n1388_i2,
  n791_i2,
  n1372_i2,
  n815_i2,
  n868_i2,
  lo018_buf_i2,
  lo138_buf_i2,
  lo158_buf_i2,
  n780_i2,
  n728_i2,
  n676_i2,
  n929_i2,
  n955_i2,
  n938_i2,
  n1117_i2,
  n1121_i2,
  n965_i2,
  n752_i2,
  n753_i2,
  n760_i2,
  n770_i2,
  n923_i2,
  n947_i2,
  n897_i2,
  n919_i2,
  n895_i2,
  n917_i2,
  n751_i2,
  n774_i2,
  lo126_buf_i2,
  lo142_buf_i2,
  lo162_buf_i2,
  n990_i2,
  n792_i2,
  n869_i2,
  n848_i2,
  lo024_buf_i2,
  lo028_buf_i2,
  lo088_buf_i2,
  lo092_buf_i2,
  lo096_buf_i2,
  lo100_buf_i2,
  n763_i2,
  n754_i2,
  n755_i2,
  n822_i2,
  n849_i2,
  n777_i2,
  n778_i2,
  n820_i2,
  n846_i2,
  n806_i2,
  n771_i2,
  n854_i2,
  n828_i2,
  lo117_buf_i2,
  lo145_buf_i2,
  n762_i2,
  n805_i2,
  n859_i2,
  n833_i2,
  lo034_buf_i2,
  lo038_buf_i2,
  lo122_buf_i2,
  lo150_buf_i2
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input G42;input G43;input G44;input G45;input G46;input G47;input G48;input G49;input G50;input n1752_lo;input n1776_lo;input n1824_lo;input n1836_lo;input n1848_lo;input n1860_lo;input n1872_lo;input n1884_lo;input n1896_lo;input n1908_lo;input n1911_lo;input n1914_lo;input n1923_lo;input n1926_lo;input n1935_lo;input n1938_lo;input n1947_lo;input n1950_lo;input n1959_lo;input n1962_lo;input n1971_lo;input n1974_lo;input n1983_lo;input n1995_lo;input n2055_lo;input n2064_lo;input n2067_lo;input n2079_lo;input n2100_lo;input n2112_lo;input n2124_lo;input n2136_lo;input n2148_lo;input n2160_lo;input n2172_lo;input n2184_lo;input n2235_lo;input n2238_lo;input n2247_lo;input n2250_lo;input n2259_lo;input n2262_lo;input n2271_lo;input n2274_lo;input n2283_lo;input n2286_lo;input n2289_lo;input n2295_lo;input n2298_lo;input n2304_lo;input n2307_lo;input n2316_lo;input n2331_lo;input n2334_lo;input n2337_lo;input n2340_lo;input n2071_o2;input n2080_o2;input n2137_o2;input n2368_o2;input n2383_o2;input n2405_o2;input n2471_o2;input n2617_o2;input n2765_o2;input n2775_o2;input n2829_o2;input n2579_o2;input n2580_o2;input n2618_o2;input n2619_o2;input n2620_o2;input n2621_o2;input n2622_o2;input n2623_o2;input n2624_o2;input n2625_o2;input n2626_o2;input n2627_o2;input n3029_o2;input n3035_o2;input n2643_o2;input n2644_o2;input n2645_o2;input n327_inv;input n2658_o2;input n2659_o2;input n2674_o2;input n2675_o2;input n2676_o2;input n3119_o2;input n3153_o2;input n351_inv;input n2729_o2;input n2730_o2;input n2731_o2;input n698_o2;input n366_inv;input n2757_o2;input n2758_o2;input n1000_o2;input n1160_o2;input n1153_o2;input n2793_o2;input n2794_o2;input n2795_o2;input n1001_o2;input n2859_o2;input n744_o2;input n402_inv;input n2926_o2;input n408_inv;input n2966_o2;input n2967_o2;input n2947_o2;input n1010_o2;input n2976_o2;input n3069_o2;input n3028_o2;input n3081_o2;input n3082_o2;input n3142_o2;input n3214_o2;input n2992_o2;input n2993_o2;input n870_o2;input n3086_o2;input n3087_o2;input n3088_o2;input n3089_o2;input n3090_o2;input n3091_o2;input n3092_o2;input n3093_o2;input n3094_o2;input n3095_o2;input n483_inv;input n3170_o2;input n3171_o2;input n3172_o2;input n3179_o2;input n498_inv;input n3193_o2;input n3211_o2;input n3212_o2;input n3213_o2;input n513_inv;input n1125_o2;input n1081_o2;input n1139_o2;input n3245_o2;input n3246_o2;input n3247_o2;input lo074_buf_o2;input lo078_buf_o2;input lo186_buf_o2;input lo118_buf_o2;input lo146_buf_o2;input n1038_o2;input n1044_o2;input n555_inv;input n558_inv;input lo026_buf_o2;input lo030_buf_o2;input lo090_buf_o2;input lo094_buf_o2;input lo098_buf_o2;input lo102_buf_o2;input lo066_buf_o2;input lo070_buf_o2;input n1202_o2;input n1003_o2;input n1031_o2;input n1034_o2;input n1040_o2;input n1046_o2;input n1380_o2;input n1425_o2;input n697_o2;input n1143_o2;input n673_o2;input n789_o2;input n786_o2;input n1047_o2;input n1036_o2;input n1307_o2;input n1035_o2;input n1297_o2;input n1099_o2;input n1128_o2;input n645_inv;input n826_o2;input n853_o2;input n654_inv;input n700_o2;input n884_o2;input lo082_buf_o2;input lo086_buf_o2;input n801_o2;input n840_o2;input n675_inv;input lo002_buf_o2;input lo010_buf_o2;input lo166_buf_o2;input lo170_buf_o2;input n1426_o2;input n1082_o2;input n1310_o2;input n1015_o2;input n1206_o2;input n1262_o2;input n1456_o2;input n1244_o2;input n1280_o2;input n1290_o2;input n1012_o2;input n1074_o2;input n1112_o2;input n1212_o2;input n1454_o2;input n1182_o2;input n1220_o2;input n701_o2;input n744_inv;input n1282_o2;input n1144_o2;input n1278_o2;input n1459_o2;input n1324_o2;input n1288_o2;input n1271_o2;input n1132_o2;input n1231_o2;input n1462_o2;input n1482_o2;input n994_o2;input n998_o2;input lo106_buf_o2;input n769_o2;input n814_o2;input n841_o2;input n867_o2;input lo006_buf_o2;input lo014_buf_o2;input lo022_buf_o2;input lo042_buf_o2;input lo046_buf_o2;input lo050_buf_o2;input lo054_buf_o2;input lo130_buf_o2;input lo134_buf_o2;input lo154_buf_o2;input lo174_buf_o2;input lo178_buf_o2;input n1007_o2;input n1294_o2;input n1084_o2;input n1399_o2;input n1311_o2;input n1392_o2;input n1102_o2;input n1041_o2;input n1298_o2;input n738_o2;input n1214_o2;input n1222_o2;input n1155_o2;input n1147_o2;input n1393_o2;input n999_o2;input n1306_o2;input n1312_o2;input n1382_o2;input n1383_o2;input n1152_o2;input n1334_o2;input n1335_o2;input n906_inv;input n773_o2;input lo190_buf_o2;input n1368_o2;input n1362_o2;input n1406_o2;input n1403_o2;input n741_o2;input n1407_o2;input n1395_o2;input n1359_o2;input n1159_o2;input n1221_o2;input n945_inv;input n989_o2;input n881_o2;input n1340_o2;input n1341_o2;input n906_o2;input n1388_o2;input n791_o2;input n1372_o2;input n815_o2;input n868_o2;input lo018_buf_o2;input lo138_buf_o2;input lo158_buf_o2;input n780_o2;input n728_o2;input n993_inv;input n929_o2;input n955_o2;input n938_o2;input n1117_o2;input n1121_o2;input n965_o2;input n752_o2;input n753_o2;input n760_o2;input n770_o2;input n923_o2;input n947_o2;input n897_o2;input n919_o2;input n895_o2;input n917_o2;input n751_o2;input n774_o2;input lo126_buf_o2;input lo142_buf_o2;input lo162_buf_o2;input n1059_inv;input n792_o2;input n869_o2;input n1068_inv;input lo024_buf_o2;input lo028_buf_o2;input lo088_buf_o2;input lo092_buf_o2;input lo096_buf_o2;input lo100_buf_o2;input n763_o2;input n754_o2;input n755_o2;input n822_o2;input n849_o2;input n777_o2;input n778_o2;input n820_o2;input n846_o2;input n806_o2;input n771_o2;input n854_o2;input n828_o2;input lo117_buf_o2;input lo145_buf_o2;input n762_o2;input n805_o2;input n859_o2;input n833_o2;input lo034_buf_o2;input lo038_buf_o2;input lo122_buf_o2;input lo150_buf_o2;
  output G3519;output G3520;output G3521;output G3522;output G3523;output G3524;output G3525;output G3526;output G3527;output G3528;output G3529;output G3530;output G3531;output G3532;output G3533;output G3534;output G3535;output G3536;output G3537;output G3538;output G3539;output G3540;output n4070_li003_li003;output n4094_li011_li011;output n4142_li027_li027;output n4154_li031_li031;output n4166_li035_li035;output n4178_li039_li039;output n4190_li043_li043;output n4202_li047_li047;output n4214_li051_li051;output n4226_li055_li055;output n4229_li056_li056;output n4232_li057_li057;output n4241_li060_li060;output n4244_li061_li061;output n4253_li064_li064;output n4256_li065_li065;output n4265_li068_li068;output n4268_li069_li069;output n4277_li072_li072;output n4280_li073_li073;output n4289_li076_li076;output n4292_li077_li077;output n4301_li080_li080;output n4313_li084_li084;output n4373_li104_li104;output n4382_li107_li107;output n4385_li108_li108;output n4397_li112_li112;output n4418_li119_li119;output n4430_li123_li123;output n4442_li127_li127;output n4454_li131_li131;output n4466_li135_li135;output n4478_li139_li139;output n4490_li143_li143;output n4502_li147_li147;output n4553_li164_li164;output n4556_li165_li165;output n4565_li168_li168;output n4568_li169_li169;output n4577_li172_li172;output n4580_li173_li173;output n4589_li176_li176;output n4592_li177_li177;output n4601_li180_li180;output n4604_li181_li181;output n4607_li182_li182;output n4613_li184_li184;output n4616_li185_li185;output n4622_li187_li187;output n4625_li188_li188;output n4634_li191_li191;output n4649_li196_li196;output n4652_li197_li197;output n4655_li198_li198;output n4658_li199_li199;output n2071_i2;output n2080_i2;output n2137_i2;output n2368_i2;output n2383_i2;output n2405_i2;output n2471_i2;output n2617_i2;output n2765_i2;output n2775_i2;output n2829_i2;output n2579_i2;output n2580_i2;output n2618_i2;output n2619_i2;output n2620_i2;output n2621_i2;output n2622_i2;output n2623_i2;output n2624_i2;output n2625_i2;output n2626_i2;output n2627_i2;output n3029_i2;output n3035_i2;output n2643_i2;output n2644_i2;output n2645_i2;output n2640_i2;output n2658_i2;output n2659_i2;output n2674_i2;output n2675_i2;output n2676_i2;output n3119_i2;output n3153_i2;output n2681_i2;output n2729_i2;output n2730_i2;output n2731_i2;output n698_i2;output n677_i2;output n2757_i2;output n2758_i2;output n1000_i2;output n1160_i2;output n1153_i2;output n2793_i2;output n2794_i2;output n2795_i2;output n1001_i2;output n2859_i2;output n744_i2;output n2908_i2;output n2926_i2;output n2928_i2;output n2966_i2;output n2967_i2;output n2947_i2;output n1010_i2;output n2976_i2;output n3069_i2;output n3028_i2;output n3081_i2;output n3082_i2;output n3142_i2;output n3214_i2;output n2992_i2;output n2993_i2;output n870_i2;output n3086_i2;output n3087_i2;output n3088_i2;output n3089_i2;output n3090_i2;output n3091_i2;output n3092_i2;output n3093_i2;output n3094_i2;output n3095_i2;output n3136_i2;output n3170_i2;output n3171_i2;output n3172_i2;output n3179_i2;output n3180_i2;output n3193_i2;output n3211_i2;output n3212_i2;output n3213_i2;output n3219_i2;output n1125_i2;output n1081_i2;output n1139_i2;output n3245_i2;output n3246_i2;output n3247_i2;output lo074_buf_i2;output lo078_buf_i2;output lo186_buf_i2;output lo118_buf_i2;output lo146_buf_i2;output n1038_i2;output n1044_i2;output n980_i2;output n1145_i2;output lo026_buf_i2;output lo030_buf_i2;output lo090_buf_i2;output lo094_buf_i2;output lo098_buf_i2;output lo102_buf_i2;output lo066_buf_i2;output lo070_buf_i2;output n1202_i2;output n1003_i2;output n1031_i2;output n1034_i2;output n1040_i2;output n1046_i2;output n1380_i2;output n1425_i2;output n697_i2;output n1143_i2;output n673_i2;output n789_i2;output n786_i2;output n1047_i2;output n1036_i2;output n1307_i2;output n1035_i2;output n1297_i2;output n1099_i2;output n1128_i2;output n674_i2;output n826_i2;output n853_i2;output n951_i2;output n700_i2;output n884_i2;output lo082_buf_i2;output lo086_buf_i2;output n801_i2;output n840_i2;output n866_i2;output lo002_buf_i2;output lo010_buf_i2;output lo166_buf_i2;output lo170_buf_i2;output n1426_i2;output n1082_i2;output n1310_i2;output n1015_i2;output n1206_i2;output n1262_i2;output n1456_i2;output n1244_i2;output n1280_i2;output n1290_i2;output n1012_i2;output n1074_i2;output n1112_i2;output n1212_i2;output n1454_i2;output n1182_i2;output n1220_i2;output n701_i2;output n973_i2;output n1282_i2;output n1144_i2;output n1278_i2;output n1459_i2;output n1324_i2;output n1288_i2;output n1271_i2;output n1132_i2;output n1231_i2;output n1462_i2;output n1482_i2;output n994_i2;output n998_i2;output lo106_buf_i2;output n769_i2;output n814_i2;output n841_i2;output n867_i2;output lo006_buf_i2;output lo014_buf_i2;output lo022_buf_i2;output lo042_buf_i2;output lo046_buf_i2;output lo050_buf_i2;output lo054_buf_i2;output lo130_buf_i2;output lo134_buf_i2;output lo154_buf_i2;output lo174_buf_i2;output lo178_buf_i2;output n1007_i2;output n1294_i2;output n1084_i2;output n1399_i2;output n1311_i2;output n1392_i2;output n1102_i2;output n1041_i2;output n1298_i2;output n738_i2;output n1214_i2;output n1222_i2;output n1155_i2;output n1147_i2;output n1393_i2;output n999_i2;output n1306_i2;output n1312_i2;output n1382_i2;output n1383_i2;output n1152_i2;output n1334_i2;output n1335_i2;output n695_i2;output n773_i2;output lo190_buf_i2;output n1368_i2;output n1362_i2;output n1406_i2;output n1403_i2;output n741_i2;output n1407_i2;output n1395_i2;output n1359_i2;output n1159_i2;output n1221_i2;output n987_i2;output n989_i2;output n881_i2;output n1340_i2;output n1341_i2;output n906_i2;output n1388_i2;output n791_i2;output n1372_i2;output n815_i2;output n868_i2;output lo018_buf_i2;output lo138_buf_i2;output lo158_buf_i2;output n780_i2;output n728_i2;output n676_i2;output n929_i2;output n955_i2;output n938_i2;output n1117_i2;output n1121_i2;output n965_i2;output n752_i2;output n753_i2;output n760_i2;output n770_i2;output n923_i2;output n947_i2;output n897_i2;output n919_i2;output n895_i2;output n917_i2;output n751_i2;output n774_i2;output lo126_buf_i2;output lo142_buf_i2;output lo162_buf_i2;output n990_i2;output n792_i2;output n869_i2;output n848_i2;output lo024_buf_i2;output lo028_buf_i2;output lo088_buf_i2;output lo092_buf_i2;output lo096_buf_i2;output lo100_buf_i2;output n763_i2;output n754_i2;output n755_i2;output n822_i2;output n849_i2;output n777_i2;output n778_i2;output n820_i2;output n846_i2;output n806_i2;output n771_i2;output n854_i2;output n828_i2;output lo117_buf_i2;output lo145_buf_i2;output n762_i2;output n805_i2;output n859_i2;output n833_i2;output lo034_buf_i2;output lo038_buf_i2;output lo122_buf_i2;output lo150_buf_i2;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire n1752_lo_p;
  wire n1752_lo_n;
  wire n1776_lo_p;
  wire n1776_lo_n;
  wire n1824_lo_p;
  wire n1824_lo_n;
  wire n1836_lo_p;
  wire n1836_lo_n;
  wire n1848_lo_p;
  wire n1848_lo_n;
  wire n1860_lo_p;
  wire n1860_lo_n;
  wire n1872_lo_p;
  wire n1872_lo_n;
  wire n1884_lo_p;
  wire n1884_lo_n;
  wire n1896_lo_p;
  wire n1896_lo_n;
  wire n1908_lo_p;
  wire n1908_lo_n;
  wire n1911_lo_p;
  wire n1911_lo_n;
  wire n1914_lo_p;
  wire n1914_lo_n;
  wire n1923_lo_p;
  wire n1923_lo_n;
  wire n1926_lo_p;
  wire n1926_lo_n;
  wire n1935_lo_p;
  wire n1935_lo_n;
  wire n1938_lo_p;
  wire n1938_lo_n;
  wire n1947_lo_p;
  wire n1947_lo_n;
  wire n1950_lo_p;
  wire n1950_lo_n;
  wire n1959_lo_p;
  wire n1959_lo_n;
  wire n1962_lo_p;
  wire n1962_lo_n;
  wire n1971_lo_p;
  wire n1971_lo_n;
  wire n1974_lo_p;
  wire n1974_lo_n;
  wire n1983_lo_p;
  wire n1983_lo_n;
  wire n1995_lo_p;
  wire n1995_lo_n;
  wire n2055_lo_p;
  wire n2055_lo_n;
  wire n2064_lo_p;
  wire n2064_lo_n;
  wire n2067_lo_p;
  wire n2067_lo_n;
  wire n2079_lo_p;
  wire n2079_lo_n;
  wire n2100_lo_p;
  wire n2100_lo_n;
  wire n2112_lo_p;
  wire n2112_lo_n;
  wire n2124_lo_p;
  wire n2124_lo_n;
  wire n2136_lo_p;
  wire n2136_lo_n;
  wire n2148_lo_p;
  wire n2148_lo_n;
  wire n2160_lo_p;
  wire n2160_lo_n;
  wire n2172_lo_p;
  wire n2172_lo_n;
  wire n2184_lo_p;
  wire n2184_lo_n;
  wire n2235_lo_p;
  wire n2235_lo_n;
  wire n2238_lo_p;
  wire n2238_lo_n;
  wire n2247_lo_p;
  wire n2247_lo_n;
  wire n2250_lo_p;
  wire n2250_lo_n;
  wire n2259_lo_p;
  wire n2259_lo_n;
  wire n2262_lo_p;
  wire n2262_lo_n;
  wire n2271_lo_p;
  wire n2271_lo_n;
  wire n2274_lo_p;
  wire n2274_lo_n;
  wire n2283_lo_p;
  wire n2283_lo_n;
  wire n2286_lo_p;
  wire n2286_lo_n;
  wire n2289_lo_p;
  wire n2289_lo_n;
  wire n2295_lo_p;
  wire n2295_lo_n;
  wire n2298_lo_p;
  wire n2298_lo_n;
  wire n2304_lo_p;
  wire n2304_lo_n;
  wire n2307_lo_p;
  wire n2307_lo_n;
  wire n2316_lo_p;
  wire n2316_lo_n;
  wire n2331_lo_p;
  wire n2331_lo_n;
  wire n2334_lo_p;
  wire n2334_lo_n;
  wire n2337_lo_p;
  wire n2337_lo_n;
  wire n2340_lo_p;
  wire n2340_lo_n;
  wire n2071_o2_p;
  wire n2071_o2_n;
  wire n2080_o2_p;
  wire n2080_o2_n;
  wire n2137_o2_p;
  wire n2137_o2_n;
  wire n2368_o2_p;
  wire n2368_o2_n;
  wire n2383_o2_p;
  wire n2383_o2_n;
  wire n2405_o2_p;
  wire n2405_o2_n;
  wire n2471_o2_p;
  wire n2471_o2_n;
  wire n2617_o2_p;
  wire n2617_o2_n;
  wire n2765_o2_p;
  wire n2765_o2_n;
  wire n2775_o2_p;
  wire n2775_o2_n;
  wire n2829_o2_p;
  wire n2829_o2_n;
  wire n2579_o2_p;
  wire n2579_o2_n;
  wire n2580_o2_p;
  wire n2580_o2_n;
  wire n2618_o2_p;
  wire n2618_o2_n;
  wire n2619_o2_p;
  wire n2619_o2_n;
  wire n2620_o2_p;
  wire n2620_o2_n;
  wire n2621_o2_p;
  wire n2621_o2_n;
  wire n2622_o2_p;
  wire n2622_o2_n;
  wire n2623_o2_p;
  wire n2623_o2_n;
  wire n2624_o2_p;
  wire n2624_o2_n;
  wire n2625_o2_p;
  wire n2625_o2_n;
  wire n2626_o2_p;
  wire n2626_o2_n;
  wire n2627_o2_p;
  wire n2627_o2_n;
  wire n3029_o2_p;
  wire n3029_o2_n;
  wire n3035_o2_p;
  wire n3035_o2_n;
  wire n2643_o2_p;
  wire n2643_o2_n;
  wire n2644_o2_p;
  wire n2644_o2_n;
  wire n2645_o2_p;
  wire n2645_o2_n;
  wire n327_inv_p;
  wire n327_inv_n;
  wire n2658_o2_p;
  wire n2658_o2_n;
  wire n2659_o2_p;
  wire n2659_o2_n;
  wire n2674_o2_p;
  wire n2674_o2_n;
  wire n2675_o2_p;
  wire n2675_o2_n;
  wire n2676_o2_p;
  wire n2676_o2_n;
  wire n3119_o2_p;
  wire n3119_o2_n;
  wire n3153_o2_p;
  wire n3153_o2_n;
  wire n351_inv_p;
  wire n351_inv_n;
  wire n2729_o2_p;
  wire n2729_o2_n;
  wire n2730_o2_p;
  wire n2730_o2_n;
  wire n2731_o2_p;
  wire n2731_o2_n;
  wire n698_o2_p;
  wire n698_o2_n;
  wire n366_inv_p;
  wire n366_inv_n;
  wire n2757_o2_p;
  wire n2757_o2_n;
  wire n2758_o2_p;
  wire n2758_o2_n;
  wire n1000_o2_p;
  wire n1000_o2_n;
  wire n1160_o2_p;
  wire n1160_o2_n;
  wire n1153_o2_p;
  wire n1153_o2_n;
  wire n2793_o2_p;
  wire n2793_o2_n;
  wire n2794_o2_p;
  wire n2794_o2_n;
  wire n2795_o2_p;
  wire n2795_o2_n;
  wire n1001_o2_p;
  wire n1001_o2_n;
  wire n2859_o2_p;
  wire n2859_o2_n;
  wire n744_o2_p;
  wire n744_o2_n;
  wire n402_inv_p;
  wire n402_inv_n;
  wire n2926_o2_p;
  wire n2926_o2_n;
  wire n408_inv_p;
  wire n408_inv_n;
  wire n2966_o2_p;
  wire n2966_o2_n;
  wire n2967_o2_p;
  wire n2967_o2_n;
  wire n2947_o2_p;
  wire n2947_o2_n;
  wire n1010_o2_p;
  wire n1010_o2_n;
  wire n2976_o2_p;
  wire n2976_o2_n;
  wire n3069_o2_p;
  wire n3069_o2_n;
  wire n3028_o2_p;
  wire n3028_o2_n;
  wire n3081_o2_p;
  wire n3081_o2_n;
  wire n3082_o2_p;
  wire n3082_o2_n;
  wire n3142_o2_p;
  wire n3142_o2_n;
  wire n3214_o2_p;
  wire n3214_o2_n;
  wire n2992_o2_p;
  wire n2992_o2_n;
  wire n2993_o2_p;
  wire n2993_o2_n;
  wire n870_o2_p;
  wire n870_o2_n;
  wire n3086_o2_p;
  wire n3086_o2_n;
  wire n3087_o2_p;
  wire n3087_o2_n;
  wire n3088_o2_p;
  wire n3088_o2_n;
  wire n3089_o2_p;
  wire n3089_o2_n;
  wire n3090_o2_p;
  wire n3090_o2_n;
  wire n3091_o2_p;
  wire n3091_o2_n;
  wire n3092_o2_p;
  wire n3092_o2_n;
  wire n3093_o2_p;
  wire n3093_o2_n;
  wire n3094_o2_p;
  wire n3094_o2_n;
  wire n3095_o2_p;
  wire n3095_o2_n;
  wire n483_inv_p;
  wire n483_inv_n;
  wire n3170_o2_p;
  wire n3170_o2_n;
  wire n3171_o2_p;
  wire n3171_o2_n;
  wire n3172_o2_p;
  wire n3172_o2_n;
  wire n3179_o2_p;
  wire n3179_o2_n;
  wire n498_inv_p;
  wire n498_inv_n;
  wire n3193_o2_p;
  wire n3193_o2_n;
  wire n3211_o2_p;
  wire n3211_o2_n;
  wire n3212_o2_p;
  wire n3212_o2_n;
  wire n3213_o2_p;
  wire n3213_o2_n;
  wire n513_inv_p;
  wire n513_inv_n;
  wire n1125_o2_p;
  wire n1125_o2_n;
  wire n1081_o2_p;
  wire n1081_o2_n;
  wire n1139_o2_p;
  wire n1139_o2_n;
  wire n3245_o2_p;
  wire n3245_o2_n;
  wire n3246_o2_p;
  wire n3246_o2_n;
  wire n3247_o2_p;
  wire n3247_o2_n;
  wire lo074_buf_o2_p;
  wire lo074_buf_o2_n;
  wire lo078_buf_o2_p;
  wire lo078_buf_o2_n;
  wire lo186_buf_o2_p;
  wire lo186_buf_o2_n;
  wire lo118_buf_o2_p;
  wire lo118_buf_o2_n;
  wire lo146_buf_o2_p;
  wire lo146_buf_o2_n;
  wire n1038_o2_p;
  wire n1038_o2_n;
  wire n1044_o2_p;
  wire n1044_o2_n;
  wire n555_inv_p;
  wire n555_inv_n;
  wire n558_inv_p;
  wire n558_inv_n;
  wire lo026_buf_o2_p;
  wire lo026_buf_o2_n;
  wire lo030_buf_o2_p;
  wire lo030_buf_o2_n;
  wire lo090_buf_o2_p;
  wire lo090_buf_o2_n;
  wire lo094_buf_o2_p;
  wire lo094_buf_o2_n;
  wire lo098_buf_o2_p;
  wire lo098_buf_o2_n;
  wire lo102_buf_o2_p;
  wire lo102_buf_o2_n;
  wire lo066_buf_o2_p;
  wire lo066_buf_o2_n;
  wire lo070_buf_o2_p;
  wire lo070_buf_o2_n;
  wire n1202_o2_p;
  wire n1202_o2_n;
  wire n1003_o2_p;
  wire n1003_o2_n;
  wire n1031_o2_p;
  wire n1031_o2_n;
  wire n1034_o2_p;
  wire n1034_o2_n;
  wire n1040_o2_p;
  wire n1040_o2_n;
  wire n1046_o2_p;
  wire n1046_o2_n;
  wire n1380_o2_p;
  wire n1380_o2_n;
  wire n1425_o2_p;
  wire n1425_o2_n;
  wire n697_o2_p;
  wire n697_o2_n;
  wire n1143_o2_p;
  wire n1143_o2_n;
  wire n673_o2_p;
  wire n673_o2_n;
  wire n789_o2_p;
  wire n789_o2_n;
  wire n786_o2_p;
  wire n786_o2_n;
  wire n1047_o2_p;
  wire n1047_o2_n;
  wire n1036_o2_p;
  wire n1036_o2_n;
  wire n1307_o2_p;
  wire n1307_o2_n;
  wire n1035_o2_p;
  wire n1035_o2_n;
  wire n1297_o2_p;
  wire n1297_o2_n;
  wire n1099_o2_p;
  wire n1099_o2_n;
  wire n1128_o2_p;
  wire n1128_o2_n;
  wire n645_inv_p;
  wire n645_inv_n;
  wire n826_o2_p;
  wire n826_o2_n;
  wire n853_o2_p;
  wire n853_o2_n;
  wire n654_inv_p;
  wire n654_inv_n;
  wire n700_o2_p;
  wire n700_o2_n;
  wire n884_o2_p;
  wire n884_o2_n;
  wire lo082_buf_o2_p;
  wire lo082_buf_o2_n;
  wire lo086_buf_o2_p;
  wire lo086_buf_o2_n;
  wire n801_o2_p;
  wire n801_o2_n;
  wire n840_o2_p;
  wire n840_o2_n;
  wire n675_inv_p;
  wire n675_inv_n;
  wire lo002_buf_o2_p;
  wire lo002_buf_o2_n;
  wire lo010_buf_o2_p;
  wire lo010_buf_o2_n;
  wire lo166_buf_o2_p;
  wire lo166_buf_o2_n;
  wire lo170_buf_o2_p;
  wire lo170_buf_o2_n;
  wire n1426_o2_p;
  wire n1426_o2_n;
  wire n1082_o2_p;
  wire n1082_o2_n;
  wire n1310_o2_p;
  wire n1310_o2_n;
  wire n1015_o2_p;
  wire n1015_o2_n;
  wire n1206_o2_p;
  wire n1206_o2_n;
  wire n1262_o2_p;
  wire n1262_o2_n;
  wire n1456_o2_p;
  wire n1456_o2_n;
  wire n1244_o2_p;
  wire n1244_o2_n;
  wire n1280_o2_p;
  wire n1280_o2_n;
  wire n1290_o2_p;
  wire n1290_o2_n;
  wire n1012_o2_p;
  wire n1012_o2_n;
  wire n1074_o2_p;
  wire n1074_o2_n;
  wire n1112_o2_p;
  wire n1112_o2_n;
  wire n1212_o2_p;
  wire n1212_o2_n;
  wire n1454_o2_p;
  wire n1454_o2_n;
  wire n1182_o2_p;
  wire n1182_o2_n;
  wire n1220_o2_p;
  wire n1220_o2_n;
  wire n701_o2_p;
  wire n701_o2_n;
  wire n744_inv_p;
  wire n744_inv_n;
  wire n1282_o2_p;
  wire n1282_o2_n;
  wire n1144_o2_p;
  wire n1144_o2_n;
  wire n1278_o2_p;
  wire n1278_o2_n;
  wire n1459_o2_p;
  wire n1459_o2_n;
  wire n1324_o2_p;
  wire n1324_o2_n;
  wire n1288_o2_p;
  wire n1288_o2_n;
  wire n1271_o2_p;
  wire n1271_o2_n;
  wire n1132_o2_p;
  wire n1132_o2_n;
  wire n1231_o2_p;
  wire n1231_o2_n;
  wire n1462_o2_p;
  wire n1462_o2_n;
  wire n1482_o2_p;
  wire n1482_o2_n;
  wire n994_o2_p;
  wire n994_o2_n;
  wire n998_o2_p;
  wire n998_o2_n;
  wire lo106_buf_o2_p;
  wire lo106_buf_o2_n;
  wire n769_o2_p;
  wire n769_o2_n;
  wire n814_o2_p;
  wire n814_o2_n;
  wire n841_o2_p;
  wire n841_o2_n;
  wire n867_o2_p;
  wire n867_o2_n;
  wire lo006_buf_o2_p;
  wire lo006_buf_o2_n;
  wire lo014_buf_o2_p;
  wire lo014_buf_o2_n;
  wire lo022_buf_o2_p;
  wire lo022_buf_o2_n;
  wire lo042_buf_o2_p;
  wire lo042_buf_o2_n;
  wire lo046_buf_o2_p;
  wire lo046_buf_o2_n;
  wire lo050_buf_o2_p;
  wire lo050_buf_o2_n;
  wire lo054_buf_o2_p;
  wire lo054_buf_o2_n;
  wire lo130_buf_o2_p;
  wire lo130_buf_o2_n;
  wire lo134_buf_o2_p;
  wire lo134_buf_o2_n;
  wire lo154_buf_o2_p;
  wire lo154_buf_o2_n;
  wire lo174_buf_o2_p;
  wire lo174_buf_o2_n;
  wire lo178_buf_o2_p;
  wire lo178_buf_o2_n;
  wire n1007_o2_p;
  wire n1007_o2_n;
  wire n1294_o2_p;
  wire n1294_o2_n;
  wire n1084_o2_p;
  wire n1084_o2_n;
  wire n1399_o2_p;
  wire n1399_o2_n;
  wire n1311_o2_p;
  wire n1311_o2_n;
  wire n1392_o2_p;
  wire n1392_o2_n;
  wire n1102_o2_p;
  wire n1102_o2_n;
  wire n1041_o2_p;
  wire n1041_o2_n;
  wire n1298_o2_p;
  wire n1298_o2_n;
  wire n738_o2_p;
  wire n738_o2_n;
  wire n1214_o2_p;
  wire n1214_o2_n;
  wire n1222_o2_p;
  wire n1222_o2_n;
  wire n1155_o2_p;
  wire n1155_o2_n;
  wire n1147_o2_p;
  wire n1147_o2_n;
  wire n1393_o2_p;
  wire n1393_o2_n;
  wire n999_o2_p;
  wire n999_o2_n;
  wire n1306_o2_p;
  wire n1306_o2_n;
  wire n1312_o2_p;
  wire n1312_o2_n;
  wire n1382_o2_p;
  wire n1382_o2_n;
  wire n1383_o2_p;
  wire n1383_o2_n;
  wire n1152_o2_p;
  wire n1152_o2_n;
  wire n1334_o2_p;
  wire n1334_o2_n;
  wire n1335_o2_p;
  wire n1335_o2_n;
  wire n906_inv_p;
  wire n906_inv_n;
  wire n773_o2_p;
  wire n773_o2_n;
  wire lo190_buf_o2_p;
  wire lo190_buf_o2_n;
  wire n1368_o2_p;
  wire n1368_o2_n;
  wire n1362_o2_p;
  wire n1362_o2_n;
  wire n1406_o2_p;
  wire n1406_o2_n;
  wire n1403_o2_p;
  wire n1403_o2_n;
  wire n741_o2_p;
  wire n741_o2_n;
  wire n1407_o2_p;
  wire n1407_o2_n;
  wire n1395_o2_p;
  wire n1395_o2_n;
  wire n1359_o2_p;
  wire n1359_o2_n;
  wire n1159_o2_p;
  wire n1159_o2_n;
  wire n1221_o2_p;
  wire n1221_o2_n;
  wire n945_inv_p;
  wire n945_inv_n;
  wire n989_o2_p;
  wire n989_o2_n;
  wire n881_o2_p;
  wire n881_o2_n;
  wire n1340_o2_p;
  wire n1340_o2_n;
  wire n1341_o2_p;
  wire n1341_o2_n;
  wire n906_o2_p;
  wire n906_o2_n;
  wire n1388_o2_p;
  wire n1388_o2_n;
  wire n791_o2_p;
  wire n791_o2_n;
  wire n1372_o2_p;
  wire n1372_o2_n;
  wire n815_o2_p;
  wire n815_o2_n;
  wire n868_o2_p;
  wire n868_o2_n;
  wire lo018_buf_o2_p;
  wire lo018_buf_o2_n;
  wire lo138_buf_o2_p;
  wire lo138_buf_o2_n;
  wire lo158_buf_o2_p;
  wire lo158_buf_o2_n;
  wire n780_o2_p;
  wire n780_o2_n;
  wire n728_o2_p;
  wire n728_o2_n;
  wire n993_inv_p;
  wire n993_inv_n;
  wire n929_o2_p;
  wire n929_o2_n;
  wire n955_o2_p;
  wire n955_o2_n;
  wire n938_o2_p;
  wire n938_o2_n;
  wire n1117_o2_p;
  wire n1117_o2_n;
  wire n1121_o2_p;
  wire n1121_o2_n;
  wire n965_o2_p;
  wire n965_o2_n;
  wire n752_o2_p;
  wire n752_o2_n;
  wire n753_o2_p;
  wire n753_o2_n;
  wire n760_o2_p;
  wire n760_o2_n;
  wire n770_o2_p;
  wire n770_o2_n;
  wire n923_o2_p;
  wire n923_o2_n;
  wire n947_o2_p;
  wire n947_o2_n;
  wire n897_o2_p;
  wire n897_o2_n;
  wire n919_o2_p;
  wire n919_o2_n;
  wire n895_o2_p;
  wire n895_o2_n;
  wire n917_o2_p;
  wire n917_o2_n;
  wire n751_o2_p;
  wire n751_o2_n;
  wire n774_o2_p;
  wire n774_o2_n;
  wire lo126_buf_o2_p;
  wire lo126_buf_o2_n;
  wire lo142_buf_o2_p;
  wire lo142_buf_o2_n;
  wire lo162_buf_o2_p;
  wire lo162_buf_o2_n;
  wire n1059_inv_p;
  wire n1059_inv_n;
  wire n792_o2_p;
  wire n792_o2_n;
  wire n869_o2_p;
  wire n869_o2_n;
  wire n1068_inv_p;
  wire n1068_inv_n;
  wire lo024_buf_o2_p;
  wire lo024_buf_o2_n;
  wire lo028_buf_o2_p;
  wire lo028_buf_o2_n;
  wire lo088_buf_o2_p;
  wire lo088_buf_o2_n;
  wire lo092_buf_o2_p;
  wire lo092_buf_o2_n;
  wire lo096_buf_o2_p;
  wire lo096_buf_o2_n;
  wire lo100_buf_o2_p;
  wire lo100_buf_o2_n;
  wire n763_o2_p;
  wire n763_o2_n;
  wire n754_o2_p;
  wire n754_o2_n;
  wire n755_o2_p;
  wire n755_o2_n;
  wire n822_o2_p;
  wire n822_o2_n;
  wire n849_o2_p;
  wire n849_o2_n;
  wire n777_o2_p;
  wire n777_o2_n;
  wire n778_o2_p;
  wire n778_o2_n;
  wire n820_o2_p;
  wire n820_o2_n;
  wire n846_o2_p;
  wire n846_o2_n;
  wire n806_o2_p;
  wire n806_o2_n;
  wire n771_o2_p;
  wire n771_o2_n;
  wire n854_o2_p;
  wire n854_o2_n;
  wire n828_o2_p;
  wire n828_o2_n;
  wire lo117_buf_o2_p;
  wire lo117_buf_o2_n;
  wire lo145_buf_o2_p;
  wire lo145_buf_o2_n;
  wire n762_o2_p;
  wire n762_o2_n;
  wire n805_o2_p;
  wire n805_o2_n;
  wire n859_o2_p;
  wire n859_o2_n;
  wire n833_o2_p;
  wire n833_o2_n;
  wire lo034_buf_o2_p;
  wire lo034_buf_o2_n;
  wire lo038_buf_o2_p;
  wire lo038_buf_o2_n;
  wire lo122_buf_o2_p;
  wire lo122_buf_o2_n;
  wire lo150_buf_o2_p;
  wire lo150_buf_o2_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire g686_p;
  wire g686_n;
  wire g687_p;
  wire g687_n;
  wire g688_p;
  wire g688_n;
  wire g689_p;
  wire g689_n;
  wire g690_p;
  wire g690_n;
  wire g691_p;
  wire g691_n;
  wire g692_p;
  wire g692_n;
  wire g693_p;
  wire g693_n;
  wire g694_p;
  wire g694_n;
  wire g695_p;
  wire g695_n;
  wire g696_p;
  wire g696_n;
  wire g697_p;
  wire g697_n;
  wire g698_p;
  wire g698_n;
  wire g699_p;
  wire g699_n;
  wire g700_p;
  wire g700_n;
  wire g701_p;
  wire g701_n;
  wire g702_p;
  wire g702_n;
  wire g703_p;
  wire g703_n;
  wire g704_p;
  wire g704_n;
  wire g705_p;
  wire g705_n;
  wire g706_p;
  wire g706_n;
  wire g707_p;
  wire g707_n;
  wire g708_p;
  wire g708_n;
  wire g709_p;
  wire g709_n;
  wire g710_p;
  wire g710_n;
  wire g711_p;
  wire g711_n;
  wire g712_p;
  wire g712_n;
  wire g713_p;
  wire g713_n;
  wire g714_p;
  wire g714_n;
  wire g715_p;
  wire g715_n;
  wire g716_p;
  wire g716_n;
  wire g717_p;
  wire g717_n;
  wire g718_p;
  wire g718_n;
  wire g719_p;
  wire g719_n;
  wire g720_p;
  wire g720_n;
  wire g721_p;
  wire g721_n;
  wire g722_p;
  wire g722_n;
  wire g723_p;
  wire g723_n;
  wire g724_p;
  wire g724_n;
  wire g725_p;
  wire g725_n;
  wire g726_p;
  wire g726_n;
  wire g727_p;
  wire g727_n;
  wire g728_p;
  wire g728_n;
  wire g729_p;
  wire g729_n;
  wire g730_p;
  wire g730_n;
  wire g731_p;
  wire g731_n;
  wire g732_p;
  wire g732_n;
  wire g733_p;
  wire g733_n;
  wire g734_p;
  wire g734_n;
  wire g735_p;
  wire g735_n;
  wire g736_p;
  wire g736_n;
  wire g737_p;
  wire g737_n;
  wire g738_p;
  wire g738_n;
  wire g739_p;
  wire g739_n;
  wire g740_p;
  wire g740_n;
  wire g741_p;
  wire g741_n;
  wire g742_p;
  wire g742_n;
  wire g743_p;
  wire g743_n;
  wire g744_p;
  wire g744_n;
  wire g745_p;
  wire g745_n;
  wire g746_p;
  wire g746_n;
  wire g747_p;
  wire g747_n;
  wire g748_p;
  wire g748_n;
  wire g749_p;
  wire g749_n;
  wire g750_p;
  wire g750_n;
  wire g751_p;
  wire g751_n;
  wire g752_p;
  wire g752_n;
  wire g753_p;
  wire g753_n;
  wire g754_p;
  wire g754_n;
  wire g755_p;
  wire g755_n;
  wire g756_p;
  wire g756_n;
  wire g757_p;
  wire g757_n;
  wire g758_p;
  wire g758_n;
  wire g759_p;
  wire g759_n;
  wire g760_p;
  wire g760_n;
  wire g761_p;
  wire g761_n;
  wire g762_p;
  wire g762_n;
  wire g763_p;
  wire g763_n;
  wire g764_p;
  wire g764_n;
  wire g765_p;
  wire g765_n;
  wire g766_p;
  wire g766_n;
  wire g767_p;
  wire g767_n;
  wire g768_p;
  wire g768_n;
  wire g769_p;
  wire g769_n;
  wire g770_p;
  wire g770_n;
  wire g771_p;
  wire g771_n;
  wire g772_p;
  wire g772_n;
  wire g773_p;
  wire g773_n;
  wire g774_p;
  wire g774_n;
  wire g775_p;
  wire g775_n;
  wire g776_p;
  wire g776_n;
  wire g777_p;
  wire g777_n;
  wire g778_p;
  wire g778_n;
  wire g779_p;
  wire g779_n;
  wire g780_p;
  wire g780_n;
  wire g781_p;
  wire g781_n;
  wire g782_p;
  wire g782_n;
  wire g783_p;
  wire g783_n;
  wire g784_p;
  wire g784_n;
  wire g785_p;
  wire g785_n;
  wire g786_p;
  wire g786_n;
  wire g787_p;
  wire g787_n;
  wire g788_p;
  wire g788_n;
  wire g789_p;
  wire g789_n;
  wire g790_p;
  wire g790_n;
  wire g791_p;
  wire g791_n;
  wire g792_p;
  wire g792_n;
  wire g793_p;
  wire g793_n;
  wire g794_p;
  wire g794_n;
  wire g795_p;
  wire g795_n;
  wire g796_p;
  wire g796_n;
  wire g797_p;
  wire g797_n;
  wire g798_p;
  wire g798_n;
  wire g799_p;
  wire g799_n;
  wire g800_p;
  wire g800_n;
  wire g801_p;
  wire g801_n;
  wire g802_p;
  wire g802_n;
  wire g803_p;
  wire g803_n;
  wire g804_p;
  wire g804_n;
  wire g805_p;
  wire g805_n;
  wire g806_p;
  wire g806_n;
  wire g807_p;
  wire g807_n;
  wire g808_p;
  wire g808_n;
  wire g809_p;
  wire g809_n;
  wire g810_p;
  wire g810_n;
  wire g811_p;
  wire g811_n;
  wire g812_p;
  wire g812_n;
  wire g813_p;
  wire g813_n;
  wire g814_p;
  wire g814_n;
  wire g815_p;
  wire g815_n;
  wire g816_p;
  wire g816_n;
  wire g817_p;
  wire g817_n;
  wire g818_p;
  wire g818_n;
  wire g819_p;
  wire g819_n;
  wire g820_p;
  wire g820_n;
  wire g821_p;
  wire g821_n;
  wire g822_p;
  wire g822_n;
  wire g823_p;
  wire g823_n;
  wire g824_p;
  wire g824_n;
  wire g825_p;
  wire g825_n;
  wire g826_p;
  wire g826_n;
  wire g827_p;
  wire g827_n;
  wire g828_p;
  wire g828_n;
  wire g829_p;
  wire g829_n;
  wire g830_p;
  wire g830_n;
  wire g831_p;
  wire g831_n;
  wire g832_p;
  wire g832_n;
  wire g833_p;
  wire g833_n;
  wire g834_p;
  wire g834_n;
  wire g835_p;
  wire g835_n;
  wire g836_p;
  wire g836_n;
  wire g837_p;
  wire g837_n;
  wire g838_p;
  wire g838_n;
  wire g839_p;
  wire g839_n;
  wire g840_p;
  wire g840_n;
  wire g841_p;
  wire g841_n;
  wire g842_p;
  wire g842_n;
  wire g843_p;
  wire g843_n;
  wire g844_p;
  wire g844_n;
  wire g845_p;
  wire g845_n;
  wire g846_p;
  wire g846_n;
  wire g847_p;
  wire g847_n;
  wire g848_p;
  wire g848_n;
  wire g849_p;
  wire g849_n;
  wire g850_p;
  wire g850_n;
  wire g851_p;
  wire g851_n;
  wire g852_p;
  wire g852_n;
  wire g853_p;
  wire g853_n;
  wire g854_p;
  wire g854_n;
  wire g855_p;
  wire g855_n;
  wire g856_p;
  wire g856_n;
  wire g857_p;
  wire g857_n;
  wire g858_p;
  wire g858_n;
  wire g859_p;
  wire g859_n;
  wire g860_p;
  wire g860_n;
  wire g861_p;
  wire g861_n;
  wire g862_p;
  wire g862_n;
  wire g863_p;
  wire g863_n;
  wire g864_p;
  wire g864_n;
  wire g865_p;
  wire g865_n;
  wire g866_p;
  wire g866_n;
  wire g867_p;
  wire g867_n;
  wire g868_p;
  wire g868_n;
  wire g869_p;
  wire g869_n;
  wire g870_p;
  wire g870_n;
  wire g871_p;
  wire g871_n;
  wire g872_p;
  wire g872_n;
  wire g873_p;
  wire g873_n;
  wire g874_p;
  wire g874_n;
  wire g875_p;
  wire g875_n;
  wire g876_p;
  wire g876_n;
  wire g877_p;
  wire g877_n;
  wire g878_p;
  wire g878_n;
  wire g879_p;
  wire g879_n;
  wire g880_p;
  wire g880_n;
  wire g881_p;
  wire g881_n;
  wire g882_p;
  wire g882_n;
  wire g883_p;
  wire g883_n;
  wire g884_p;
  wire g884_n;
  wire g885_p;
  wire g885_n;
  wire g886_p;
  wire g886_n;
  wire g887_p;
  wire g887_n;
  wire g888_p;
  wire g888_n;
  wire g889_p;
  wire g889_n;
  wire g890_p;
  wire g890_n;
  wire g891_p;
  wire g891_n;
  wire g892_p;
  wire g892_n;
  wire g893_p;
  wire g893_n;
  wire g894_p;
  wire g894_n;
  wire g895_p;
  wire g895_n;
  wire g896_p;
  wire g896_n;
  wire g897_p;
  wire g897_n;
  wire g898_p;
  wire g898_n;
  wire g899_p;
  wire g899_n;
  wire g900_p;
  wire g900_n;
  wire g901_p;
  wire g901_n;
  wire g902_p;
  wire g902_n;
  wire g903_p;
  wire g903_n;
  wire g904_p;
  wire g904_n;
  wire g905_p;
  wire g905_n;
  wire g906_p;
  wire g906_n;
  wire g907_p;
  wire g907_n;
  wire g908_p;
  wire g908_n;
  wire g909_p;
  wire g909_n;
  wire g910_p;
  wire g910_n;
  wire g911_p;
  wire g911_n;
  wire g912_p;
  wire g912_n;
  wire g913_p;
  wire g913_n;
  wire g914_p;
  wire g914_n;
  wire g915_p;
  wire g915_n;
  wire g916_p;
  wire g916_n;
  wire g917_p;
  wire g917_n;
  wire g918_p;
  wire g918_n;
  wire g919_p;
  wire g919_n;
  wire g920_p;
  wire g920_n;
  wire g921_p;
  wire g921_n;
  wire g922_p;
  wire g922_n;
  wire g923_p;
  wire g923_n;
  wire g924_p;
  wire g924_n;
  wire g925_p;
  wire g925_n;
  wire g926_p;
  wire g926_n;
  wire g927_p;
  wire g927_n;
  wire g928_p;
  wire g928_n;
  wire g929_p;
  wire g929_n;
  wire g930_p;
  wire g930_n;
  wire g931_p;
  wire g931_n;
  wire g932_p;
  wire g932_n;
  wire g933_p;
  wire g933_n;
  wire g934_p;
  wire g934_n;
  wire g935_p;
  wire g935_n;
  wire g936_p;
  wire g936_n;
  wire g937_p;
  wire g937_n;
  wire g938_p;
  wire g938_n;
  wire g939_p;
  wire g939_n;
  wire g940_p;
  wire g940_n;
  wire g941_p;
  wire g941_n;
  wire g942_p;
  wire g942_n;
  wire g943_p;
  wire g943_n;
  wire g944_p;
  wire g944_n;
  wire g945_p;
  wire g945_n;
  wire g946_p;
  wire g946_n;
  wire g947_p;
  wire g947_n;
  wire g948_p;
  wire g948_n;
  wire g949_p;
  wire g949_n;
  wire g950_p;
  wire g950_n;
  wire g951_p;
  wire g951_n;
  wire g952_p;
  wire g952_n;
  wire g953_p;
  wire g953_n;
  wire g954_p;
  wire g954_n;
  wire g955_p;
  wire g955_n;
  wire g956_p;
  wire g956_n;
  wire g957_p;
  wire g957_n;
  wire g958_p;
  wire g958_n;
  wire g959_p;
  wire g959_n;
  wire g960_p;
  wire g960_n;
  wire g961_p;
  wire g961_n;
  wire g962_p;
  wire g962_n;
  wire g963_p;
  wire g963_n;
  wire g964_p;
  wire g964_n;
  wire g965_p;
  wire g965_n;
  wire g966_p;
  wire g966_n;
  wire g967_p;
  wire g967_n;
  wire g968_p;
  wire g968_n;
  wire g969_p;
  wire g969_n;
  wire g970_p;
  wire g970_n;
  wire g971_p;
  wire g971_n;
  wire g972_p;
  wire g972_n;
  wire g973_p;
  wire g973_n;
  wire g974_p;
  wire g974_n;
  wire g975_p;
  wire g975_n;
  wire g976_p;
  wire g976_n;
  wire g977_p;
  wire g977_n;
  wire g978_p;
  wire g978_n;
  wire g979_p;
  wire g979_n;
  wire g980_p;
  wire g980_n;
  wire g981_p;
  wire g981_n;
  wire g982_p;
  wire g982_n;
  wire g983_p;
  wire g983_n;
  wire g984_p;
  wire g984_n;
  wire g985_p;
  wire g985_n;
  wire g986_p;
  wire g986_n;
  wire g987_p;
  wire g987_n;
  wire g988_p;
  wire g988_n;
  wire g989_p;
  wire g989_n;
  wire g990_p;
  wire g990_n;
  wire g991_p;
  wire g991_n;
  wire g992_p;
  wire g992_n;
  wire g993_p;
  wire g993_n;
  wire g994_p;
  wire g994_n;
  wire g995_p;
  wire g995_n;
  wire g996_p;
  wire g996_n;
  wire g997_p;
  wire g997_n;
  wire g998_p;
  wire g998_n;
  wire g999_p;
  wire g999_n;
  wire g1000_p;
  wire g1000_n;
  wire g1001_p;
  wire g1001_n;
  wire g1002_p;
  wire g1002_n;
  wire g1003_p;
  wire g1003_n;
  wire g1004_p;
  wire g1004_n;
  wire g1005_p;
  wire g1005_n;
  wire g1006_p;
  wire g1006_n;
  wire g1007_p;
  wire g1007_n;
  wire g1008_p;
  wire g1008_n;
  wire g1009_p;
  wire g1009_n;
  wire g1010_p;
  wire g1010_n;
  wire g1011_p;
  wire g1011_n;
  wire g1012_p;
  wire g1012_n;
  wire g1013_p;
  wire g1013_n;
  wire g1014_p;
  wire g1014_n;
  wire g1015_p;
  wire g1015_n;
  wire g1016_p;
  wire g1016_n;
  wire g1017_p;
  wire g1017_n;
  wire g1018_p;
  wire g1018_n;
  wire g1019_p;
  wire g1019_n;
  wire g1020_p;
  wire g1020_n;
  wire g1021_p;
  wire g1021_n;
  wire g1022_p;
  wire g1022_n;
  wire g1023_p;
  wire g1023_n;
  wire g1024_p;
  wire g1024_n;
  wire g1025_p;
  wire g1025_n;
  wire g1026_p;
  wire g1026_n;
  wire g1027_p;
  wire g1027_n;
  wire g1028_p;
  wire g1028_n;
  wire g1029_p;
  wire g1029_n;
  wire g1030_p;
  wire g1030_n;
  wire g1031_p;
  wire g1031_n;
  wire g1032_p;
  wire g1032_n;
  wire g1033_p;
  wire g1033_n;
  wire g1034_p;
  wire g1034_n;
  wire g1035_p;
  wire g1035_n;
  wire g1036_p;
  wire g1036_n;
  wire g1037_p;
  wire g1037_n;
  wire g1038_p;
  wire g1038_n;
  wire g1039_p;
  wire g1039_n;
  wire g1040_p;
  wire g1040_n;
  wire g1041_p;
  wire g1041_n;
  wire g1042_p;
  wire g1042_n;
  wire g1043_p;
  wire g1043_n;
  wire g1044_p;
  wire g1044_n;
  wire g1045_p;
  wire g1045_n;
  wire g1046_p;
  wire g1046_n;
  wire g1047_p;
  wire g1047_n;
  wire g1048_p;
  wire g1048_n;
  wire g1049_p;
  wire g1049_n;
  wire g1050_p;
  wire g1050_n;
  wire g1051_p;
  wire g1051_n;
  wire g1052_p;
  wire g1052_n;
  wire g1053_p;
  wire g1053_n;
  wire g1054_p;
  wire g1054_n;
  wire g1055_p;
  wire g1055_n;
  wire g1056_p;
  wire g1056_n;
  wire g1057_p;
  wire g1057_n;
  wire g1058_p;
  wire g1058_n;
  wire g1059_p;
  wire g1059_n;
  wire g1060_p;
  wire g1060_n;
  wire g1061_p;
  wire g1061_n;
  wire g1062_p;
  wire g1062_n;
  wire g1063_p;
  wire g1063_n;
  wire g1064_p;
  wire g1064_n;
  wire g1065_p;
  wire g1065_n;
  wire g1066_p;
  wire g1066_n;
  wire g1067_p;
  wire g1067_n;
  wire g1068_p;
  wire g1068_n;
  wire g1069_p;
  wire g1069_n;
  wire g1070_p;
  wire g1070_n;
  wire g1071_p;
  wire g1071_n;
  wire g1072_p;
  wire g1072_n;
  wire g1073_p;
  wire g1073_n;
  wire g1074_p;
  wire g1074_n;
  wire g1075_p;
  wire g1075_n;
  wire g1076_p;
  wire g1076_n;
  wire g1077_p;
  wire g1077_n;
  wire g1078_p;
  wire g1078_n;
  wire g1079_p;
  wire g1079_n;
  wire g1080_p;
  wire g1080_n;
  wire g1081_p;
  wire g1081_n;
  wire g1082_p;
  wire g1082_n;
  wire g1083_p;
  wire g1083_n;
  wire g1084_p;
  wire g1084_n;
  wire g1085_p;
  wire g1085_n;
  wire g1086_p;
  wire g1086_n;
  wire g1087_p;
  wire g1087_n;
  wire g1088_p;
  wire g1088_n;
  wire g1089_p;
  wire g1089_n;
  wire g1090_p;
  wire g1090_n;
  wire g1091_p;
  wire g1091_n;
  wire g1092_p;
  wire g1092_n;
  wire g1093_p;
  wire g1093_n;
  wire g1094_p;
  wire g1094_n;
  wire g1095_p;
  wire g1095_n;
  wire g1096_p;
  wire g1096_n;
  wire g1097_p;
  wire g1097_n;
  wire g1098_p;
  wire g1098_n;
  wire g1099_p;
  wire g1099_n;
  wire g1100_p;
  wire g1100_n;
  wire g1101_p;
  wire g1101_n;
  wire g1102_p;
  wire g1102_n;
  wire g1103_p;
  wire g1103_n;
  wire g1104_p;
  wire g1104_n;
  wire g1105_p;
  wire g1105_n;
  wire g1106_p;
  wire g1106_n;
  wire g1107_p;
  wire g1107_n;
  wire g1108_p;
  wire g1108_n;
  wire g1109_p;
  wire g1109_n;
  wire g1110_p;
  wire g1110_n;
  wire g1111_p;
  wire g1111_n;
  wire g1112_p;
  wire g1112_n;
  wire g1113_p;
  wire g1113_n;
  wire g1114_p;
  wire g1114_n;
  wire g1115_p;
  wire g1115_n;
  wire g1116_p;
  wire g1116_n;
  wire g1117_p;
  wire g1117_n;
  wire g1118_p;
  wire g1118_n;
  wire g1119_p;
  wire g1119_n;
  wire g1120_p;
  wire g1120_n;
  wire g1121_p;
  wire g1121_n;
  wire g1122_p;
  wire g1122_n;
  wire g1123_p;
  wire g1123_n;
  wire g1124_p;
  wire g1124_n;
  wire g1125_p;
  wire g1125_n;
  wire g1126_p;
  wire g1126_n;
  wire g1127_p;
  wire g1127_n;
  wire g1128_p;
  wire g1128_n;
  wire g1129_p;
  wire g1129_n;
  wire g1130_p;
  wire g1130_n;
  wire g1131_p;
  wire g1131_n;
  wire g1132_p;
  wire g1132_n;
  wire g1133_p;
  wire g1133_n;
  wire g1134_p;
  wire g1134_n;
  wire g1135_p;
  wire g1135_n;
  wire g1136_p;
  wire g1136_n;
  wire g1137_p;
  wire g1137_n;
  wire g1138_p;
  wire g1138_n;
  wire g1139_p;
  wire g1139_n;
  wire g1140_p;
  wire g1140_n;
  wire g1141_p;
  wire g1141_n;
  wire g1142_p;
  wire g1142_n;
  wire g1143_p;
  wire g1143_n;
  wire g1144_p;
  wire g1144_n;
  wire g1145_p;
  wire g1145_n;
  wire g1146_p;
  wire g1146_n;
  wire g1147_p;
  wire g1147_n;
  wire g1148_p;
  wire g1148_n;
  wire g1149_p;
  wire g1149_n;
  wire g1150_p;
  wire g1150_n;
  wire g1151_p;
  wire g1151_n;
  wire g1152_p;
  wire g1152_n;
  wire g1153_p;
  wire g1153_n;
  wire g1154_p;
  wire g1154_n;
  wire g1155_p;
  wire g1155_n;
  wire g1156_p;
  wire g1156_n;
  wire g1157_p;
  wire g1157_n;
  wire g1158_p;
  wire g1158_n;
  wire g1159_p;
  wire g1159_n;
  wire g1160_p;
  wire g1160_n;
  wire g1161_p;
  wire g1161_n;
  wire g1162_p;
  wire g1162_n;
  wire g1163_p;
  wire g1163_n;
  wire g1164_p;
  wire g1164_n;
  wire g1165_p;
  wire g1165_n;
  wire g1166_p;
  wire g1166_n;
  wire g1167_p;
  wire g1167_n;
  wire g1168_p;
  wire g1168_n;
  wire g1169_p;
  wire g1169_n;
  wire g1170_p;
  wire g1170_n;
  wire g1171_p;
  wire g1171_n;
  wire g1172_p;
  wire g1172_n;
  wire g1173_p;
  wire g1173_n;
  wire g1174_p;
  wire g1174_n;
  wire g1175_p;
  wire g1175_n;
  wire g1176_p;
  wire g1176_n;
  wire g1177_p;
  wire g1177_n;
  wire g1178_p;
  wire g1178_n;
  wire g1179_p;
  wire g1179_n;
  wire g1180_p;
  wire g1180_n;
  wire g1181_p;
  wire g1181_n;
  wire g1182_p;
  wire g1182_n;
  wire g1183_p;
  wire g1183_n;
  wire g1184_p;
  wire g1184_n;
  wire g1185_p;
  wire g1185_n;
  wire g1186_p;
  wire g1186_n;
  wire g1187_p;
  wire g1187_n;
  wire g1188_p;
  wire g1188_n;
  wire g1189_p;
  wire g1189_n;
  wire g1190_p;
  wire g1190_n;
  wire g1191_p;
  wire g1191_n;
  wire g1192_p;
  wire g1192_n;
  wire g1193_p;
  wire g1193_n;
  wire g1194_p;
  wire g1194_n;
  wire g1195_p;
  wire g1195_n;
  wire g1196_p;
  wire g1196_n;
  wire g1197_p;
  wire g1197_n;
  wire g1198_p;
  wire g1198_n;
  wire g1199_p;
  wire g1199_n;
  wire g1200_p;
  wire g1200_n;
  wire g1201_p;
  wire g1201_n;
  wire g1202_p;
  wire g1202_n;
  wire g1203_p;
  wire g1203_n;
  wire g1204_p;
  wire g1204_n;
  wire g1205_p;
  wire g1205_n;
  wire g1206_p;
  wire g1206_n;
  wire g1207_p;
  wire g1207_n;
  wire g1208_p;
  wire g1208_n;
  wire g1209_p;
  wire g1209_n;
  wire g1210_p;
  wire g1210_n;
  wire g1211_p;
  wire g1211_n;
  wire g1212_p;
  wire g1212_n;
  wire g1213_p;
  wire g1213_n;
  wire g1214_p;
  wire g1214_n;
  wire g1215_p;
  wire g1215_n;
  wire g1216_p;
  wire g1216_n;
  wire g1217_p;
  wire g1217_n;
  wire g1218_p;
  wire g1218_n;
  wire g1219_p;
  wire g1219_n;
  wire g1220_p;
  wire g1220_n;
  wire g1221_p;
  wire g1221_n;
  wire g1222_p;
  wire g1222_n;
  wire g1223_p;
  wire g1223_n;
  wire g1224_p;
  wire g1224_n;
  wire g1225_p;
  wire g1225_n;
  wire g1226_p;
  wire g1226_n;
  wire g1227_p;
  wire g1227_n;
  wire g1228_p;
  wire g1228_n;
  wire g1229_p;
  wire g1229_n;
  wire g1230_p;
  wire g1230_n;
  wire g1231_p;
  wire g1231_n;
  wire g1232_p;
  wire g1232_n;
  wire g1233_p;
  wire g1233_n;
  wire g1234_p;
  wire g1234_n;
  wire g1235_p;
  wire g1235_n;
  wire n1860_lo_n_spl_;
  wire n1776_lo_n_spl_;
  wire n1752_lo_n_spl_;
  wire n2148_lo_n_spl_;
  wire n2148_lo_n_spl_0;
  wire n2148_lo_n_spl_1;
  wire n1872_lo_p_spl_;
  wire n2124_lo_n_spl_;
  wire n2124_lo_n_spl_0;
  wire n2100_lo_n_spl_;
  wire n2100_lo_n_spl_0;
  wire n1824_lo_p_spl_;
  wire n2136_lo_n_spl_;
  wire n2136_lo_n_spl_0;
  wire n2184_lo_n_spl_;
  wire n2184_lo_n_spl_0;
  wire n1908_lo_p_spl_;
  wire n1908_lo_p_spl_0;
  wire n2112_lo_n_spl_;
  wire n2112_lo_n_spl_0;
  wire n2160_lo_n_spl_;
  wire n2160_lo_n_spl_0;
  wire n2160_lo_n_spl_1;
  wire n1884_lo_p_spl_;
  wire n2172_lo_n_spl_;
  wire n2172_lo_n_spl_0;
  wire n2172_lo_n_spl_1;
  wire n1896_lo_p_spl_;
  wire n1896_lo_p_spl_0;
  wire g430_n_spl_;
  wire n2172_lo_p_spl_;
  wire n2184_lo_p_spl_;
  wire n2148_lo_p_spl_;
  wire n2160_lo_p_spl_;
  wire g442_p_spl_;
  wire g439_n_spl_;
  wire g442_n_spl_;
  wire g439_p_spl_;
  wire n2124_lo_p_spl_;
  wire n2136_lo_p_spl_;
  wire n2100_lo_p_spl_;
  wire n2112_lo_p_spl_;
  wire g451_n_spl_;
  wire g448_p_spl_;
  wire g451_p_spl_;
  wire g448_n_spl_;
  wire n1908_lo_n_spl_;
  wire n1908_lo_n_spl_0;
  wire n1896_lo_n_spl_;
  wire g462_p_spl_;
  wire g459_p_spl_;
  wire g462_n_spl_;
  wire g459_n_spl_;
  wire n3029_o2_p_spl_;
  wire n1001_o2_n_spl_;
  wire n1001_o2_n_spl_0;
  wire n1010_o2_n_spl_;
  wire n1010_o2_p_spl_;
  wire g481_n_spl_;
  wire n3119_o2_p_spl_;
  wire g481_p_spl_;
  wire n3119_o2_n_spl_;
  wire n1153_o2_p_spl_;
  wire n1160_o2_p_spl_;
  wire n1153_o2_n_spl_;
  wire n1160_o2_n_spl_;
  wire n1001_o2_p_spl_;
  wire g514_p_spl_;
  wire g480_p_spl_;
  wire g514_n_spl_;
  wire g514_n_spl_0;
  wire g480_n_spl_;
  wire g480_n_spl_0;
  wire g511_p_spl_;
  wire g505_p_spl_;
  wire g511_n_spl_;
  wire g511_n_spl_0;
  wire g505_n_spl_;
  wire g505_n_spl_0;
  wire g508_p_spl_;
  wire g477_p_spl_;
  wire g508_n_spl_;
  wire g508_n_spl_0;
  wire g477_n_spl_;
  wire g477_n_spl_0;
  wire g517_n_spl_;
  wire g516_n_spl_;
  wire g515_n_spl_;
  wire n1462_o2_p_spl_;
  wire n1462_o2_p_spl_0;
  wire n2064_lo_p_spl_;
  wire g521_n_spl_;
  wire g520_n_spl_;
  wire g528_n_spl_;
  wire g526_p_spl_;
  wire g528_p_spl_;
  wire g526_n_spl_;
  wire g534_n_spl_;
  wire g534_n_spl_0;
  wire g534_n_spl_1;
  wire n2340_lo_p_spl_;
  wire g534_p_spl_;
  wire g534_p_spl_0;
  wire g534_p_spl_1;
  wire n2340_lo_n_spl_;
  wire g538_p_spl_;
  wire g533_p_spl_;
  wire g533_p_spl_0;
  wire g533_p_spl_1;
  wire g538_n_spl_;
  wire g533_n_spl_;
  wire g533_n_spl_0;
  wire g533_n_spl_1;
  wire g531_n_spl_;
  wire g531_p_spl_;
  wire n2793_o2_p_spl_;
  wire n2793_o2_p_spl_0;
  wire n2793_o2_p_spl_1;
  wire n2621_o2_n_spl_;
  wire n994_o2_n_spl_;
  wire n994_o2_n_spl_0;
  wire n994_o2_p_spl_;
  wire n945_inv_p_spl_;
  wire n3028_o2_n_spl_;
  wire n3028_o2_p_spl_;
  wire n3028_o2_p_spl_0;
  wire n2620_o2_p_spl_;
  wire n1007_o2_p_spl_;
  wire n2620_o2_n_spl_;
  wire n2579_o2_p_spl_;
  wire g561_p_spl_;
  wire g556_p_spl_;
  wire g556_p_spl_0;
  wire g561_n_spl_;
  wire g561_n_spl_0;
  wire g561_n_spl_00;
  wire g561_n_spl_01;
  wire g561_n_spl_1;
  wire g556_n_spl_;
  wire g556_n_spl_0;
  wire g556_n_spl_1;
  wire n869_o2_p_spl_;
  wire n792_o2_p_spl_;
  wire n869_o2_n_spl_;
  wire n792_o2_n_spl_;
  wire n1059_inv_n_spl_;
  wire n1059_inv_n_spl_0;
  wire n1059_inv_n_spl_00;
  wire n1059_inv_n_spl_000;
  wire n1059_inv_n_spl_001;
  wire n1059_inv_n_spl_01;
  wire n1059_inv_n_spl_1;
  wire n1059_inv_n_spl_10;
  wire n1059_inv_n_spl_11;
  wire n1059_inv_p_spl_;
  wire n1059_inv_p_spl_0;
  wire n1059_inv_p_spl_00;
  wire n1059_inv_p_spl_000;
  wire n1059_inv_p_spl_001;
  wire n1059_inv_p_spl_01;
  wire n1059_inv_p_spl_010;
  wire n1059_inv_p_spl_011;
  wire n1059_inv_p_spl_1;
  wire n1059_inv_p_spl_10;
  wire n1059_inv_p_spl_11;
  wire g563_p_spl_;
  wire n897_o2_n_spl_;
  wire n897_o2_n_spl_0;
  wire n897_o2_p_spl_;
  wire g569_n_spl_;
  wire g568_n_spl_;
  wire g568_n_spl_0;
  wire g569_p_spl_;
  wire g568_p_spl_;
  wire n919_o2_n_spl_;
  wire n919_o2_n_spl_0;
  wire n919_o2_p_spl_;
  wire g574_n_spl_;
  wire g573_n_spl_;
  wire g573_n_spl_0;
  wire g574_p_spl_;
  wire g573_p_spl_;
  wire n2993_o2_p_spl_;
  wire n2993_o2_p_spl_0;
  wire n2993_o2_p_spl_00;
  wire n2993_o2_p_spl_1;
  wire n2993_o2_n_spl_;
  wire n2993_o2_n_spl_0;
  wire g579_p_spl_;
  wire g579_p_spl_0;
  wire g579_p_spl_00;
  wire g579_p_spl_01;
  wire g579_p_spl_1;
  wire lo102_buf_o2_n_spl_;
  wire g578_p_spl_;
  wire g578_p_spl_0;
  wire g578_p_spl_1;
  wire lo102_buf_o2_p_spl_;
  wire n791_o2_n_spl_;
  wire n814_o2_p_spl_;
  wire n841_o2_p_spl_;
  wire n675_inv_p_spl_;
  wire g572_p_spl_;
  wire g572_p_spl_0;
  wire g567_p_spl_;
  wire g567_p_spl_0;
  wire lo026_buf_o2_n_spl_;
  wire n1962_lo_p_spl_;
  wire n1962_lo_p_spl_0;
  wire g589_n_spl_;
  wire g593_n_spl_;
  wire g578_n_spl_;
  wire g593_p_spl_;
  wire g594_p_spl_;
  wire g579_n_spl_;
  wire g579_n_spl_0;
  wire g579_n_spl_1;
  wire g594_n_spl_;
  wire g596_p_spl_;
  wire g596_n_spl_;
  wire n1334_o2_n_spl_;
  wire n1334_o2_p_spl_;
  wire n1147_o2_p_spl_;
  wire lo186_buf_o2_p_spl_;
  wire lo186_buf_o2_p_spl_0;
  wire lo186_buf_o2_p_spl_1;
  wire lo186_buf_o2_n_spl_;
  wire lo186_buf_o2_n_spl_0;
  wire lo186_buf_o2_n_spl_1;
  wire g555_p_spl_;
  wire g603_n_spl_;
  wire g601_n_spl_;
  wire g601_n_spl_0;
  wire g603_p_spl_;
  wire g601_p_spl_;
  wire g604_n_spl_;
  wire g600_n_spl_;
  wire g600_n_spl_0;
  wire n2619_o2_n_spl_;
  wire n2619_o2_n_spl_0;
  wire n2619_o2_n_spl_00;
  wire n2619_o2_n_spl_01;
  wire n2619_o2_n_spl_1;
  wire n2619_o2_n_spl_10;
  wire g609_n_spl_;
  wire g609_n_spl_0;
  wire g609_n_spl_1;
  wire n2580_o2_p_spl_;
  wire n327_inv_p_spl_;
  wire g612_p_spl_;
  wire g612_p_spl_0;
  wire g612_p_spl_00;
  wire g612_p_spl_01;
  wire g612_p_spl_1;
  wire g612_p_spl_10;
  wire g562_p_spl_;
  wire g562_p_spl_0;
  wire g562_p_spl_00;
  wire g562_p_spl_01;
  wire g562_p_spl_1;
  wire g562_p_spl_10;
  wire g622_n_spl_;
  wire g622_n_spl_0;
  wire g554_n_spl_;
  wire g554_n_spl_0;
  wire g622_p_spl_;
  wire g554_p_spl_;
  wire lo034_buf_o2_p_spl_;
  wire lo034_buf_o2_p_spl_0;
  wire lo034_buf_o2_p_spl_00;
  wire lo034_buf_o2_p_spl_1;
  wire lo028_buf_o2_p_spl_;
  wire lo028_buf_o2_p_spl_0;
  wire lo028_buf_o2_p_spl_1;
  wire n965_o2_n_spl_;
  wire n965_o2_p_spl_;
  wire n786_o2_n_spl_;
  wire g648_p_spl_;
  wire g648_p_spl_0;
  wire g648_n_spl_;
  wire g648_n_spl_0;
  wire n789_o2_p_spl_;
  wire n789_o2_n_spl_;
  wire g651_n_spl_;
  wire g651_p_spl_;
  wire n989_o2_n_spl_;
  wire n989_o2_n_spl_0;
  wire g653_n_spl_;
  wire g652_n_spl_;
  wire g652_n_spl_0;
  wire g653_p_spl_;
  wire g652_p_spl_;
  wire lo024_buf_o2_p_spl_;
  wire lo024_buf_o2_p_spl_0;
  wire lo024_buf_o2_p_spl_1;
  wire lo092_buf_o2_n_spl_;
  wire lo092_buf_o2_p_spl_;
  wire lo092_buf_o2_p_spl_0;
  wire lo088_buf_o2_p_spl_;
  wire lo100_buf_o2_p_spl_;
  wire lo096_buf_o2_p_spl_;
  wire g599_n_spl_;
  wire g599_n_spl_0;
  wire n3089_o2_n_spl_;
  wire g597_p_spl_;
  wire g597_p_spl_0;
  wire n3091_o2_p_spl_;
  wire g598_p_spl_;
  wire g597_n_spl_;
  wire g597_n_spl_0;
  wire g597_n_spl_1;
  wire n3245_o2_n_spl_;
  wire g595_p_spl_;
  wire n3246_o2_p_spl_;
  wire n3246_o2_p_spl_0;
  wire n3246_o2_p_spl_00;
  wire n3246_o2_p_spl_1;
  wire lo086_buf_o2_p_spl_;
  wire lo086_buf_o2_p_spl_0;
  wire n1950_lo_p_spl_;
  wire n1950_lo_p_spl_0;
  wire g592_n_spl_;
  wire g657_n_spl_;
  wire n762_o2_n_spl_;
  wire g668_n_spl_;
  wire g668_n_spl_0;
  wire g668_n_spl_1;
  wire lo042_buf_o2_p_spl_;
  wire lo042_buf_o2_p_spl_0;
  wire lo042_buf_o2_p_spl_00;
  wire lo042_buf_o2_p_spl_1;
  wire g668_p_spl_;
  wire g668_p_spl_0;
  wire g668_p_spl_1;
  wire lo042_buf_o2_n_spl_;
  wire lo042_buf_o2_n_spl_0;
  wire lo042_buf_o2_n_spl_1;
  wire n760_o2_n_spl_;
  wire n760_o2_n_spl_0;
  wire n760_o2_n_spl_1;
  wire n760_o2_p_spl_;
  wire n760_o2_p_spl_0;
  wire n760_o2_p_spl_00;
  wire n760_o2_p_spl_01;
  wire n760_o2_p_spl_1;
  wire n760_o2_p_spl_10;
  wire lo034_buf_o2_n_spl_;
  wire lo034_buf_o2_n_spl_0;
  wire lo034_buf_o2_n_spl_1;
  wire n754_o2_n_spl_;
  wire n754_o2_n_spl_0;
  wire n754_o2_n_spl_1;
  wire n754_o2_p_spl_;
  wire n754_o2_p_spl_0;
  wire n751_o2_p_spl_;
  wire n751_o2_p_spl_0;
  wire n751_o2_p_spl_00;
  wire n751_o2_p_spl_000;
  wire n751_o2_p_spl_01;
  wire n751_o2_p_spl_1;
  wire n751_o2_p_spl_10;
  wire n751_o2_p_spl_11;
  wire n751_o2_n_spl_;
  wire n751_o2_n_spl_0;
  wire n751_o2_n_spl_00;
  wire n751_o2_n_spl_1;
  wire lo046_buf_o2_p_spl_;
  wire lo046_buf_o2_p_spl_0;
  wire lo046_buf_o2_p_spl_1;
  wire lo046_buf_o2_n_spl_;
  wire lo046_buf_o2_n_spl_0;
  wire lo046_buf_o2_n_spl_1;
  wire lo038_buf_o2_p_spl_;
  wire lo038_buf_o2_p_spl_0;
  wire lo038_buf_o2_p_spl_00;
  wire lo038_buf_o2_p_spl_1;
  wire n755_o2_n_spl_;
  wire n755_o2_n_spl_0;
  wire n755_o2_n_spl_1;
  wire lo038_buf_o2_n_spl_;
  wire lo028_buf_o2_n_spl_;
  wire lo028_buf_o2_n_spl_0;
  wire lo028_buf_o2_n_spl_1;
  wire g646_n_spl_;
  wire lo006_buf_o2_p_spl_;
  wire lo002_buf_o2_p_spl_;
  wire lo002_buf_o2_p_spl_0;
  wire lo002_buf_o2_p_spl_1;
  wire n771_o2_n_spl_;
  wire n771_o2_n_spl_0;
  wire n771_o2_n_spl_00;
  wire n771_o2_n_spl_01;
  wire n771_o2_n_spl_1;
  wire n771_o2_n_spl_10;
  wire n771_o2_p_spl_;
  wire n771_o2_p_spl_0;
  wire n771_o2_p_spl_00;
  wire n771_o2_p_spl_01;
  wire n771_o2_p_spl_1;
  wire n771_o2_p_spl_10;
  wire lo018_buf_o2_p_spl_;
  wire lo022_buf_o2_p_spl_;
  wire g690_p_spl_;
  wire g690_p_spl_0;
  wire g688_p_spl_;
  wire g688_p_spl_0;
  wire g690_n_spl_;
  wire g690_n_spl_0;
  wire g688_n_spl_;
  wire g688_n_spl_0;
  wire lo010_buf_o2_p_spl_;
  wire lo010_buf_o2_p_spl_0;
  wire lo010_buf_o2_p_spl_00;
  wire lo010_buf_o2_p_spl_1;
  wire lo010_buf_o2_n_spl_;
  wire g692_n_spl_;
  wire g692_p_spl_;
  wire g692_p_spl_0;
  wire g693_n_spl_;
  wire lo050_buf_o2_n_spl_;
  wire lo050_buf_o2_n_spl_0;
  wire lo050_buf_o2_p_spl_;
  wire lo050_buf_o2_p_spl_0;
  wire n753_o2_p_spl_;
  wire n753_o2_p_spl_0;
  wire lo054_buf_o2_p_spl_;
  wire lo054_buf_o2_p_spl_0;
  wire lo054_buf_o2_p_spl_1;
  wire n753_o2_n_spl_;
  wire lo054_buf_o2_n_spl_;
  wire lo054_buf_o2_n_spl_0;
  wire g705_n_spl_;
  wire g658_p_spl_;
  wire g658_p_spl_0;
  wire g658_p_spl_1;
  wire n774_o2_n_spl_;
  wire n774_o2_n_spl_0;
  wire n774_o2_p_spl_;
  wire n774_o2_p_spl_0;
  wire g708_n_spl_;
  wire g708_n_spl_0;
  wire g708_p_spl_;
  wire g708_p_spl_0;
  wire g711_n_spl_;
  wire n1081_o2_n_spl_;
  wire g661_n_spl_;
  wire n3087_o2_p_spl_;
  wire n3087_o2_p_spl_0;
  wire g717_n_spl_;
  wire g717_n_spl_0;
  wire g717_n_spl_1;
  wire n998_o2_n_spl_;
  wire n3245_o2_p_spl_;
  wire n3245_o2_p_spl_0;
  wire n3245_o2_p_spl_1;
  wire g599_p_spl_;
  wire n998_o2_p_spl_;
  wire n1221_o2_p_spl_;
  wire n1221_o2_n_spl_;
  wire g724_n_spl_;
  wire g722_n_spl_;
  wire g724_p_spl_;
  wire g722_p_spl_;
  wire g722_p_spl_0;
  wire n1214_o2_n_spl_;
  wire n3082_o2_n_spl_;
  wire n1214_o2_p_spl_;
  wire n3082_o2_p_spl_;
  wire g731_n_spl_;
  wire g553_n_spl_;
  wire g731_p_spl_;
  wire g553_p_spl_;
  wire g553_p_spl_0;
  wire g732_p_spl_;
  wire g730_p_spl_;
  wire g730_p_spl_0;
  wire g730_p_spl_1;
  wire g732_n_spl_;
  wire g730_n_spl_;
  wire g730_n_spl_0;
  wire g730_n_spl_00;
  wire g730_n_spl_1;
  wire g735_p_spl_;
  wire g727_p_spl_;
  wire n1003_o2_p_spl_;
  wire n1003_o2_p_spl_0;
  wire n1003_o2_p_spl_1;
  wire g727_n_spl_;
  wire g727_n_spl_0;
  wire g735_n_spl_;
  wire n2619_o2_p_spl_;
  wire n2619_o2_p_spl_0;
  wire n2619_o2_p_spl_00;
  wire n2619_o2_p_spl_01;
  wire n2619_o2_p_spl_1;
  wire n2619_o2_p_spl_10;
  wire n2624_o2_n_spl_;
  wire n2624_o2_n_spl_0;
  wire n2624_o2_n_spl_1;
  wire g559_n_spl_;
  wire g551_n_spl_;
  wire g552_n_spl_;
  wire g612_n_spl_;
  wire n1040_o2_p_spl_;
  wire n1040_o2_p_spl_0;
  wire n1040_o2_p_spl_00;
  wire n1040_o2_p_spl_1;
  wire n1044_o2_n_spl_;
  wire n1044_o2_n_spl_0;
  wire n1044_o2_n_spl_1;
  wire n1034_o2_p_spl_;
  wire n1034_o2_p_spl_0;
  wire n1034_o2_p_spl_1;
  wire n1046_o2_p_spl_;
  wire n1046_o2_p_spl_0;
  wire n2676_o2_n_spl_;
  wire n1038_o2_p_spl_;
  wire n1038_o2_p_spl_0;
  wire n1038_o2_p_spl_1;
  wire n1031_o2_n_spl_;
  wire n1031_o2_n_spl_0;
  wire n2645_o2_n_spl_;
  wire g760_p_spl_;
  wire n2794_o2_p_spl_;
  wire n2794_o2_p_spl_0;
  wire n2622_o2_p_spl_;
  wire g771_n_spl_;
  wire g562_n_spl_;
  wire n2624_o2_p_spl_;
  wire n2621_o2_p_spl_;
  wire n2623_o2_p_spl_;
  wire n1031_o2_p_spl_;
  wire n1031_o2_p_spl_0;
  wire n1031_o2_p_spl_00;
  wire n1031_o2_p_spl_1;
  wire n2623_o2_n_spl_;
  wire n1038_o2_n_spl_;
  wire n1038_o2_n_spl_0;
  wire n1038_o2_n_spl_00;
  wire n1038_o2_n_spl_01;
  wire n1038_o2_n_spl_1;
  wire n1038_o2_n_spl_10;
  wire lo170_buf_o2_p_spl_;
  wire n2627_o2_p_spl_;
  wire n2627_o2_p_spl_0;
  wire n2627_o2_p_spl_1;
  wire n1040_o2_n_spl_;
  wire n1040_o2_n_spl_0;
  wire n1040_o2_n_spl_00;
  wire n1040_o2_n_spl_000;
  wire n1040_o2_n_spl_01;
  wire n1040_o2_n_spl_1;
  wire n1040_o2_n_spl_10;
  wire n1040_o2_n_spl_11;
  wire n2645_o2_p_spl_;
  wire n2645_o2_p_spl_0;
  wire n2622_o2_n_spl_;
  wire n1034_o2_n_spl_;
  wire n1034_o2_n_spl_0;
  wire n1034_o2_n_spl_00;
  wire n1034_o2_n_spl_01;
  wire n1034_o2_n_spl_1;
  wire n1046_o2_n_spl_;
  wire n1046_o2_n_spl_0;
  wire n1046_o2_n_spl_00;
  wire n1046_o2_n_spl_01;
  wire n1046_o2_n_spl_1;
  wire n1046_o2_n_spl_10;
  wire n1044_o2_p_spl_;
  wire n1044_o2_p_spl_0;
  wire n1044_o2_p_spl_00;
  wire n1044_o2_p_spl_01;
  wire n1044_o2_p_spl_1;
  wire n1044_o2_p_spl_10;
  wire n2676_o2_p_spl_;
  wire n2966_o2_p_spl_;
  wire n2966_o2_p_spl_0;
  wire g849_p_spl_;
  wire g848_n_spl_;
  wire n2967_o2_p_spl_;
  wire n2967_o2_p_spl_0;
  wire n1298_o2_n_spl_;
  wire n2793_o2_n_spl_;
  wire n3214_o2_p_spl_;
  wire n3214_o2_n_spl_;
  wire g870_n_spl_;
  wire n3081_o2_n_spl_;
  wire g870_p_spl_;
  wire n3081_o2_p_spl_;
  wire g873_n_spl_;
  wire g873_n_spl_0;
  wire g687_n_spl_;
  wire g878_n_spl_;
  wire g877_p_spl_;
  wire g877_p_spl_0;
  wire g883_n_spl_;
  wire g883_n_spl_0;
  wire g883_n_spl_1;
  wire g884_n_spl_;
  wire g885_n_spl_;
  wire n1003_o2_n_spl_;
  wire n1003_o2_n_spl_0;
  wire g888_n_spl_;
  wire g656_n_spl_;
  wire g577_n_spl_;
  wire g577_n_spl_0;
  wire lo174_buf_o2_p_spl_;
  wire lo030_buf_o2_p_spl_;
  wire lo030_buf_o2_p_spl_0;
  wire n3090_o2_p_spl_;
  wire g960_p_spl_;
  wire g960_n_spl_;
  wire g873_p_spl_;
  wire g645_n_spl_;
  wire g645_n_spl_0;
  wire g621_n_spl_;
  wire g621_n_spl_0;
  wire lo154_buf_o2_p_spl_;
  wire lo142_buf_o2_p_spl_;
  wire g990_n_spl_;
  wire g705_p_spl_;
  wire g659_n_spl_;
  wire g659_n_spl_0;
  wire g659_n_spl_00;
  wire g659_n_spl_01;
  wire g659_n_spl_1;
  wire g659_n_spl_10;
  wire g676_n_spl_;
  wire g707_n_spl_;
  wire g711_p_spl_;
  wire g684_n_spl_;
  wire g713_n_spl_;
  wire n3086_o2_p_spl_;
  wire lo026_buf_o2_p_spl_;
  wire n3089_o2_p_spl_;
  wire n3092_o2_p_spl_;
  wire g581_n_spl_;
  wire g581_n_spl_0;
  wire g581_n_spl_00;
  wire g581_n_spl_01;
  wire g581_n_spl_1;
  wire n3092_o2_n_spl_;
  wire n3213_o2_p_spl_;
  wire g583_n_spl_;
  wire g583_n_spl_0;
  wire g583_n_spl_00;
  wire g583_n_spl_01;
  wire g583_n_spl_1;
  wire n1938_lo_p_spl_;
  wire n1938_lo_p_spl_0;
  wire g1013_p_spl_;
  wire g1013_p_spl_0;
  wire g890_n_spl_;
  wire g886_n_spl_;
  wire g886_n_spl_0;
  wire n1926_lo_p_spl_;
  wire g976_n_spl_;
  wire n2298_lo_n_spl_;
  wire n2250_lo_p_spl_;
  wire n2238_lo_p_spl_;
  wire g1020_n_spl_;
  wire g590_p_spl_;
  wire n2298_lo_p_spl_;
  wire g577_p_spl_;
  wire g577_p_spl_0;
  wire g1026_p_spl_;
  wire g656_p_spl_;
  wire g656_p_spl_0;
  wire g1031_n_spl_;
  wire g1025_n_spl_;
  wire g1025_n_spl_0;
  wire G2_n_spl_;
  wire G1_p_spl_;
  wire G1_p_spl_0;
  wire G6_p_spl_;
  wire g664_n_spl_;
  wire g662_n_spl_;
  wire g716_p_spl_;
  wire lo082_buf_o2_p_spl_;
  wire lo082_buf_o2_p_spl_0;
  wire g591_n_spl_;
  wire n1974_lo_p_spl_;
  wire n1974_lo_p_spl_0;
  wire g598_n_spl_;
  wire g598_n_spl_0;
  wire g598_n_spl_1;
  wire n3170_o2_p_spl_;
  wire g719_n_spl_;
  wire n3095_o2_p_spl_;
  wire n3095_o2_p_spl_0;
  wire g950_n_spl_;
  wire g720_n_spl_;
  wire g595_n_spl_;
  wire g595_n_spl_0;
  wire g972_n_spl_;
  wire g875_n_spl_;
  wire g876_n_spl_;
  wire n752_o2_p_spl_;
  wire n752_o2_p_spl_0;
  wire g1082_p_spl_;
  wire g1082_p_spl_0;
  wire g1082_p_spl_1;
  wire g666_p_spl_;
  wire g1088_p_spl_;
  wire g1086_n_spl_;
  wire g665_n_spl_;
  wire lo145_buf_o2_p_spl_;
  wire n780_o2_n_spl_;
  wire n780_o2_n_spl_0;
  wire lo138_buf_o2_p_spl_;
  wire n780_o2_p_spl_;
  wire n780_o2_p_spl_0;
  wire g1108_n_spl_;
  wire g663_p_spl_;
  wire g660_p_spl_;
  wire g990_p_spl_;
  wire g701_n_spl_;
  wire g992_n_spl_;
  wire g998_p_spl_;
  wire g995_p_spl_;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_00;
  wire G4_p_spl_000;
  wire G4_p_spl_001;
  wire G4_p_spl_01;
  wire G4_p_spl_1;
  wire G4_p_spl_10;
  wire G4_p_spl_11;
  wire G12_p_spl_;
  wire G12_p_spl_0;
  wire G12_p_spl_1;
  wire G11_p_spl_;
  wire G13_p_spl_;
  wire G13_p_spl_0;
  wire n1983_lo_p_spl_;
  wire g667_n_spl_;
  wire n1995_lo_p_spl_;
  wire g686_p_spl_;
  wire lo117_buf_o2_p_spl_;
  wire lo117_buf_o2_p_spl_0;
  wire lo014_buf_o2_p_spl_;
  wire lo014_buf_o2_p_spl_0;
  wire lo014_buf_o2_p_spl_00;
  wire lo014_buf_o2_p_spl_1;
  wire lo014_buf_o2_n_spl_;
  wire lo014_buf_o2_n_spl_0;
  wire lo014_buf_o2_n_spl_1;
  wire n2079_lo_p_spl_;
  wire g1108_p_spl_;
  wire lo122_buf_o2_p_spl_;
  wire g691_p_spl_;
  wire G4_n_spl_;
  wire G4_n_spl_0;
  wire G4_n_spl_00;
  wire G4_n_spl_1;
  wire G3_p_spl_;
  wire G3_p_spl_0;
  wire G3_p_spl_00;
  wire G3_p_spl_1;
  wire g1034_n_spl_;
  wire G3_n_spl_;
  wire G5_p_spl_;
  wire G5_p_spl_0;
  wire lo126_buf_o2_n_spl_;
  wire lo122_buf_o2_n_spl_;
  wire g691_n_spl_;
  wire g1179_p_spl_;
  wire g658_n_spl_;
  wire g658_n_spl_0;
  wire g1085_n_spl_;
  wire g1085_n_spl_0;
  wire g1190_p_spl_;
  wire g1098_n_spl_;
  wire g1098_n_spl_0;
  wire G1_n_spl_;
  wire G1_n_spl_0;
  wire g1197_n_spl_;
  wire g1035_n_spl_;
  wire g1035_n_spl_0;
  wire g1074_n_spl_;
  wire g985_n_spl_;
  wire g1110_n_spl_;
  wire g1121_p_spl_;
  wire g1120_p_spl_;
  wire G13_n_spl_;
  wire g1124_n_spl_;
  wire g1123_n_spl_;
  wire g1208_p_spl_;
  wire G41_p_spl_;
  wire g1162_n_spl_;
  wire g1162_n_spl_0;
  wire g1162_n_spl_1;
  wire g1122_n_spl_;
  wire g1122_n_spl_0;
  wire g1122_n_spl_1;
  wire G34_n_spl_;
  wire g1164_p_spl_;
  wire g1201_n_spl_;
  wire G35_p_spl_;
  wire G35_p_spl_0;
  wire g1200_p_spl_;
  wire g1163_n_spl_;
  wire G40_p_spl_;
  wire G33_p_spl_;
  wire G14_p_spl_;
  wire G34_p_spl_;
  wire g1210_n_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    G37_p,
    G37
  );


  not

  (
    G37_n,
    G37
  );


  buf

  (
    G38_p,
    G38
  );


  not

  (
    G38_n,
    G38
  );


  buf

  (
    G39_p,
    G39
  );


  not

  (
    G39_n,
    G39
  );


  buf

  (
    G40_p,
    G40
  );


  not

  (
    G40_n,
    G40
  );


  buf

  (
    G41_p,
    G41
  );


  not

  (
    G41_n,
    G41
  );


  buf

  (
    G42_p,
    G42
  );


  not

  (
    G42_n,
    G42
  );


  buf

  (
    G43_p,
    G43
  );


  not

  (
    G43_n,
    G43
  );


  buf

  (
    G44_p,
    G44
  );


  not

  (
    G44_n,
    G44
  );


  buf

  (
    G45_p,
    G45
  );


  not

  (
    G45_n,
    G45
  );


  buf

  (
    G46_p,
    G46
  );


  not

  (
    G46_n,
    G46
  );


  buf

  (
    G47_p,
    G47
  );


  not

  (
    G47_n,
    G47
  );


  buf

  (
    G48_p,
    G48
  );


  not

  (
    G48_n,
    G48
  );


  buf

  (
    G49_p,
    G49
  );


  not

  (
    G49_n,
    G49
  );


  buf

  (
    G50_p,
    G50
  );


  not

  (
    G50_n,
    G50
  );


  buf

  (
    n1752_lo_p,
    n1752_lo
  );


  not

  (
    n1752_lo_n,
    n1752_lo
  );


  buf

  (
    n1776_lo_p,
    n1776_lo
  );


  not

  (
    n1776_lo_n,
    n1776_lo
  );


  buf

  (
    n1824_lo_p,
    n1824_lo
  );


  not

  (
    n1824_lo_n,
    n1824_lo
  );


  buf

  (
    n1836_lo_p,
    n1836_lo
  );


  not

  (
    n1836_lo_n,
    n1836_lo
  );


  buf

  (
    n1848_lo_p,
    n1848_lo
  );


  not

  (
    n1848_lo_n,
    n1848_lo
  );


  buf

  (
    n1860_lo_p,
    n1860_lo
  );


  not

  (
    n1860_lo_n,
    n1860_lo
  );


  buf

  (
    n1872_lo_p,
    n1872_lo
  );


  not

  (
    n1872_lo_n,
    n1872_lo
  );


  buf

  (
    n1884_lo_p,
    n1884_lo
  );


  not

  (
    n1884_lo_n,
    n1884_lo
  );


  buf

  (
    n1896_lo_p,
    n1896_lo
  );


  not

  (
    n1896_lo_n,
    n1896_lo
  );


  buf

  (
    n1908_lo_p,
    n1908_lo
  );


  not

  (
    n1908_lo_n,
    n1908_lo
  );


  buf

  (
    n1911_lo_p,
    n1911_lo
  );


  not

  (
    n1911_lo_n,
    n1911_lo
  );


  buf

  (
    n1914_lo_p,
    n1914_lo
  );


  not

  (
    n1914_lo_n,
    n1914_lo
  );


  buf

  (
    n1923_lo_p,
    n1923_lo
  );


  not

  (
    n1923_lo_n,
    n1923_lo
  );


  buf

  (
    n1926_lo_p,
    n1926_lo
  );


  not

  (
    n1926_lo_n,
    n1926_lo
  );


  buf

  (
    n1935_lo_p,
    n1935_lo
  );


  not

  (
    n1935_lo_n,
    n1935_lo
  );


  buf

  (
    n1938_lo_p,
    n1938_lo
  );


  not

  (
    n1938_lo_n,
    n1938_lo
  );


  buf

  (
    n1947_lo_p,
    n1947_lo
  );


  not

  (
    n1947_lo_n,
    n1947_lo
  );


  buf

  (
    n1950_lo_p,
    n1950_lo
  );


  not

  (
    n1950_lo_n,
    n1950_lo
  );


  buf

  (
    n1959_lo_p,
    n1959_lo
  );


  not

  (
    n1959_lo_n,
    n1959_lo
  );


  buf

  (
    n1962_lo_p,
    n1962_lo
  );


  not

  (
    n1962_lo_n,
    n1962_lo
  );


  buf

  (
    n1971_lo_p,
    n1971_lo
  );


  not

  (
    n1971_lo_n,
    n1971_lo
  );


  buf

  (
    n1974_lo_p,
    n1974_lo
  );


  not

  (
    n1974_lo_n,
    n1974_lo
  );


  buf

  (
    n1983_lo_p,
    n1983_lo
  );


  not

  (
    n1983_lo_n,
    n1983_lo
  );


  buf

  (
    n1995_lo_p,
    n1995_lo
  );


  not

  (
    n1995_lo_n,
    n1995_lo
  );


  buf

  (
    n2055_lo_p,
    n2055_lo
  );


  not

  (
    n2055_lo_n,
    n2055_lo
  );


  buf

  (
    n2064_lo_p,
    n2064_lo
  );


  not

  (
    n2064_lo_n,
    n2064_lo
  );


  buf

  (
    n2067_lo_p,
    n2067_lo
  );


  not

  (
    n2067_lo_n,
    n2067_lo
  );


  buf

  (
    n2079_lo_p,
    n2079_lo
  );


  not

  (
    n2079_lo_n,
    n2079_lo
  );


  buf

  (
    n2100_lo_p,
    n2100_lo
  );


  not

  (
    n2100_lo_n,
    n2100_lo
  );


  buf

  (
    n2112_lo_p,
    n2112_lo
  );


  not

  (
    n2112_lo_n,
    n2112_lo
  );


  buf

  (
    n2124_lo_p,
    n2124_lo
  );


  not

  (
    n2124_lo_n,
    n2124_lo
  );


  buf

  (
    n2136_lo_p,
    n2136_lo
  );


  not

  (
    n2136_lo_n,
    n2136_lo
  );


  buf

  (
    n2148_lo_p,
    n2148_lo
  );


  not

  (
    n2148_lo_n,
    n2148_lo
  );


  buf

  (
    n2160_lo_p,
    n2160_lo
  );


  not

  (
    n2160_lo_n,
    n2160_lo
  );


  buf

  (
    n2172_lo_p,
    n2172_lo
  );


  not

  (
    n2172_lo_n,
    n2172_lo
  );


  buf

  (
    n2184_lo_p,
    n2184_lo
  );


  not

  (
    n2184_lo_n,
    n2184_lo
  );


  buf

  (
    n2235_lo_p,
    n2235_lo
  );


  not

  (
    n2235_lo_n,
    n2235_lo
  );


  buf

  (
    n2238_lo_p,
    n2238_lo
  );


  not

  (
    n2238_lo_n,
    n2238_lo
  );


  buf

  (
    n2247_lo_p,
    n2247_lo
  );


  not

  (
    n2247_lo_n,
    n2247_lo
  );


  buf

  (
    n2250_lo_p,
    n2250_lo
  );


  not

  (
    n2250_lo_n,
    n2250_lo
  );


  buf

  (
    n2259_lo_p,
    n2259_lo
  );


  not

  (
    n2259_lo_n,
    n2259_lo
  );


  buf

  (
    n2262_lo_p,
    n2262_lo
  );


  not

  (
    n2262_lo_n,
    n2262_lo
  );


  buf

  (
    n2271_lo_p,
    n2271_lo
  );


  not

  (
    n2271_lo_n,
    n2271_lo
  );


  buf

  (
    n2274_lo_p,
    n2274_lo
  );


  not

  (
    n2274_lo_n,
    n2274_lo
  );


  buf

  (
    n2283_lo_p,
    n2283_lo
  );


  not

  (
    n2283_lo_n,
    n2283_lo
  );


  buf

  (
    n2286_lo_p,
    n2286_lo
  );


  not

  (
    n2286_lo_n,
    n2286_lo
  );


  buf

  (
    n2289_lo_p,
    n2289_lo
  );


  not

  (
    n2289_lo_n,
    n2289_lo
  );


  buf

  (
    n2295_lo_p,
    n2295_lo
  );


  not

  (
    n2295_lo_n,
    n2295_lo
  );


  buf

  (
    n2298_lo_p,
    n2298_lo
  );


  not

  (
    n2298_lo_n,
    n2298_lo
  );


  buf

  (
    n2304_lo_p,
    n2304_lo
  );


  not

  (
    n2304_lo_n,
    n2304_lo
  );


  buf

  (
    n2307_lo_p,
    n2307_lo
  );


  not

  (
    n2307_lo_n,
    n2307_lo
  );


  buf

  (
    n2316_lo_p,
    n2316_lo
  );


  not

  (
    n2316_lo_n,
    n2316_lo
  );


  buf

  (
    n2331_lo_p,
    n2331_lo
  );


  not

  (
    n2331_lo_n,
    n2331_lo
  );


  buf

  (
    n2334_lo_p,
    n2334_lo
  );


  not

  (
    n2334_lo_n,
    n2334_lo
  );


  buf

  (
    n2337_lo_p,
    n2337_lo
  );


  not

  (
    n2337_lo_n,
    n2337_lo
  );


  buf

  (
    n2340_lo_p,
    n2340_lo
  );


  not

  (
    n2340_lo_n,
    n2340_lo
  );


  buf

  (
    n2071_o2_p,
    n2071_o2
  );


  not

  (
    n2071_o2_n,
    n2071_o2
  );


  buf

  (
    n2080_o2_p,
    n2080_o2
  );


  not

  (
    n2080_o2_n,
    n2080_o2
  );


  buf

  (
    n2137_o2_p,
    n2137_o2
  );


  not

  (
    n2137_o2_n,
    n2137_o2
  );


  buf

  (
    n2368_o2_p,
    n2368_o2
  );


  not

  (
    n2368_o2_n,
    n2368_o2
  );


  buf

  (
    n2383_o2_p,
    n2383_o2
  );


  not

  (
    n2383_o2_n,
    n2383_o2
  );


  buf

  (
    n2405_o2_p,
    n2405_o2
  );


  not

  (
    n2405_o2_n,
    n2405_o2
  );


  buf

  (
    n2471_o2_p,
    n2471_o2
  );


  not

  (
    n2471_o2_n,
    n2471_o2
  );


  buf

  (
    n2617_o2_p,
    n2617_o2
  );


  not

  (
    n2617_o2_n,
    n2617_o2
  );


  buf

  (
    n2765_o2_p,
    n2765_o2
  );


  not

  (
    n2765_o2_n,
    n2765_o2
  );


  buf

  (
    n2775_o2_p,
    n2775_o2
  );


  not

  (
    n2775_o2_n,
    n2775_o2
  );


  buf

  (
    n2829_o2_p,
    n2829_o2
  );


  not

  (
    n2829_o2_n,
    n2829_o2
  );


  buf

  (
    n2579_o2_p,
    n2579_o2
  );


  not

  (
    n2579_o2_n,
    n2579_o2
  );


  buf

  (
    n2580_o2_p,
    n2580_o2
  );


  not

  (
    n2580_o2_n,
    n2580_o2
  );


  buf

  (
    n2618_o2_p,
    n2618_o2
  );


  not

  (
    n2618_o2_n,
    n2618_o2
  );


  buf

  (
    n2619_o2_p,
    n2619_o2
  );


  not

  (
    n2619_o2_n,
    n2619_o2
  );


  buf

  (
    n2620_o2_p,
    n2620_o2
  );


  not

  (
    n2620_o2_n,
    n2620_o2
  );


  buf

  (
    n2621_o2_p,
    n2621_o2
  );


  not

  (
    n2621_o2_n,
    n2621_o2
  );


  buf

  (
    n2622_o2_p,
    n2622_o2
  );


  not

  (
    n2622_o2_n,
    n2622_o2
  );


  buf

  (
    n2623_o2_p,
    n2623_o2
  );


  not

  (
    n2623_o2_n,
    n2623_o2
  );


  buf

  (
    n2624_o2_p,
    n2624_o2
  );


  not

  (
    n2624_o2_n,
    n2624_o2
  );


  buf

  (
    n2625_o2_p,
    n2625_o2
  );


  not

  (
    n2625_o2_n,
    n2625_o2
  );


  buf

  (
    n2626_o2_p,
    n2626_o2
  );


  not

  (
    n2626_o2_n,
    n2626_o2
  );


  buf

  (
    n2627_o2_p,
    n2627_o2
  );


  not

  (
    n2627_o2_n,
    n2627_o2
  );


  buf

  (
    n3029_o2_p,
    n3029_o2
  );


  not

  (
    n3029_o2_n,
    n3029_o2
  );


  buf

  (
    n3035_o2_p,
    n3035_o2
  );


  not

  (
    n3035_o2_n,
    n3035_o2
  );


  buf

  (
    n2643_o2_p,
    n2643_o2
  );


  not

  (
    n2643_o2_n,
    n2643_o2
  );


  buf

  (
    n2644_o2_p,
    n2644_o2
  );


  not

  (
    n2644_o2_n,
    n2644_o2
  );


  buf

  (
    n2645_o2_p,
    n2645_o2
  );


  not

  (
    n2645_o2_n,
    n2645_o2
  );


  buf

  (
    n327_inv_p,
    n327_inv
  );


  not

  (
    n327_inv_n,
    n327_inv
  );


  buf

  (
    n2658_o2_p,
    n2658_o2
  );


  not

  (
    n2658_o2_n,
    n2658_o2
  );


  buf

  (
    n2659_o2_p,
    n2659_o2
  );


  not

  (
    n2659_o2_n,
    n2659_o2
  );


  buf

  (
    n2674_o2_p,
    n2674_o2
  );


  not

  (
    n2674_o2_n,
    n2674_o2
  );


  buf

  (
    n2675_o2_p,
    n2675_o2
  );


  not

  (
    n2675_o2_n,
    n2675_o2
  );


  buf

  (
    n2676_o2_p,
    n2676_o2
  );


  not

  (
    n2676_o2_n,
    n2676_o2
  );


  buf

  (
    n3119_o2_p,
    n3119_o2
  );


  not

  (
    n3119_o2_n,
    n3119_o2
  );


  buf

  (
    n3153_o2_p,
    n3153_o2
  );


  not

  (
    n3153_o2_n,
    n3153_o2
  );


  buf

  (
    n351_inv_p,
    n351_inv
  );


  not

  (
    n351_inv_n,
    n351_inv
  );


  buf

  (
    n2729_o2_p,
    n2729_o2
  );


  not

  (
    n2729_o2_n,
    n2729_o2
  );


  buf

  (
    n2730_o2_p,
    n2730_o2
  );


  not

  (
    n2730_o2_n,
    n2730_o2
  );


  buf

  (
    n2731_o2_p,
    n2731_o2
  );


  not

  (
    n2731_o2_n,
    n2731_o2
  );


  buf

  (
    n698_o2_p,
    n698_o2
  );


  not

  (
    n698_o2_n,
    n698_o2
  );


  buf

  (
    n366_inv_p,
    n366_inv
  );


  not

  (
    n366_inv_n,
    n366_inv
  );


  buf

  (
    n2757_o2_p,
    n2757_o2
  );


  not

  (
    n2757_o2_n,
    n2757_o2
  );


  buf

  (
    n2758_o2_p,
    n2758_o2
  );


  not

  (
    n2758_o2_n,
    n2758_o2
  );


  buf

  (
    n1000_o2_p,
    n1000_o2
  );


  not

  (
    n1000_o2_n,
    n1000_o2
  );


  buf

  (
    n1160_o2_p,
    n1160_o2
  );


  not

  (
    n1160_o2_n,
    n1160_o2
  );


  buf

  (
    n1153_o2_p,
    n1153_o2
  );


  not

  (
    n1153_o2_n,
    n1153_o2
  );


  buf

  (
    n2793_o2_p,
    n2793_o2
  );


  not

  (
    n2793_o2_n,
    n2793_o2
  );


  buf

  (
    n2794_o2_p,
    n2794_o2
  );


  not

  (
    n2794_o2_n,
    n2794_o2
  );


  buf

  (
    n2795_o2_p,
    n2795_o2
  );


  not

  (
    n2795_o2_n,
    n2795_o2
  );


  buf

  (
    n1001_o2_p,
    n1001_o2
  );


  not

  (
    n1001_o2_n,
    n1001_o2
  );


  buf

  (
    n2859_o2_p,
    n2859_o2
  );


  not

  (
    n2859_o2_n,
    n2859_o2
  );


  buf

  (
    n744_o2_p,
    n744_o2
  );


  not

  (
    n744_o2_n,
    n744_o2
  );


  buf

  (
    n402_inv_p,
    n402_inv
  );


  not

  (
    n402_inv_n,
    n402_inv
  );


  buf

  (
    n2926_o2_p,
    n2926_o2
  );


  not

  (
    n2926_o2_n,
    n2926_o2
  );


  buf

  (
    n408_inv_p,
    n408_inv
  );


  not

  (
    n408_inv_n,
    n408_inv
  );


  buf

  (
    n2966_o2_p,
    n2966_o2
  );


  not

  (
    n2966_o2_n,
    n2966_o2
  );


  buf

  (
    n2967_o2_p,
    n2967_o2
  );


  not

  (
    n2967_o2_n,
    n2967_o2
  );


  buf

  (
    n2947_o2_p,
    n2947_o2
  );


  not

  (
    n2947_o2_n,
    n2947_o2
  );


  buf

  (
    n1010_o2_p,
    n1010_o2
  );


  not

  (
    n1010_o2_n,
    n1010_o2
  );


  buf

  (
    n2976_o2_p,
    n2976_o2
  );


  not

  (
    n2976_o2_n,
    n2976_o2
  );


  buf

  (
    n3069_o2_p,
    n3069_o2
  );


  not

  (
    n3069_o2_n,
    n3069_o2
  );


  buf

  (
    n3028_o2_p,
    n3028_o2
  );


  not

  (
    n3028_o2_n,
    n3028_o2
  );


  buf

  (
    n3081_o2_p,
    n3081_o2
  );


  not

  (
    n3081_o2_n,
    n3081_o2
  );


  buf

  (
    n3082_o2_p,
    n3082_o2
  );


  not

  (
    n3082_o2_n,
    n3082_o2
  );


  buf

  (
    n3142_o2_p,
    n3142_o2
  );


  not

  (
    n3142_o2_n,
    n3142_o2
  );


  buf

  (
    n3214_o2_p,
    n3214_o2
  );


  not

  (
    n3214_o2_n,
    n3214_o2
  );


  buf

  (
    n2992_o2_p,
    n2992_o2
  );


  not

  (
    n2992_o2_n,
    n2992_o2
  );


  buf

  (
    n2993_o2_p,
    n2993_o2
  );


  not

  (
    n2993_o2_n,
    n2993_o2
  );


  buf

  (
    n870_o2_p,
    n870_o2
  );


  not

  (
    n870_o2_n,
    n870_o2
  );


  buf

  (
    n3086_o2_p,
    n3086_o2
  );


  not

  (
    n3086_o2_n,
    n3086_o2
  );


  buf

  (
    n3087_o2_p,
    n3087_o2
  );


  not

  (
    n3087_o2_n,
    n3087_o2
  );


  buf

  (
    n3088_o2_p,
    n3088_o2
  );


  not

  (
    n3088_o2_n,
    n3088_o2
  );


  buf

  (
    n3089_o2_p,
    n3089_o2
  );


  not

  (
    n3089_o2_n,
    n3089_o2
  );


  buf

  (
    n3090_o2_p,
    n3090_o2
  );


  not

  (
    n3090_o2_n,
    n3090_o2
  );


  buf

  (
    n3091_o2_p,
    n3091_o2
  );


  not

  (
    n3091_o2_n,
    n3091_o2
  );


  buf

  (
    n3092_o2_p,
    n3092_o2
  );


  not

  (
    n3092_o2_n,
    n3092_o2
  );


  buf

  (
    n3093_o2_p,
    n3093_o2
  );


  not

  (
    n3093_o2_n,
    n3093_o2
  );


  buf

  (
    n3094_o2_p,
    n3094_o2
  );


  not

  (
    n3094_o2_n,
    n3094_o2
  );


  buf

  (
    n3095_o2_p,
    n3095_o2
  );


  not

  (
    n3095_o2_n,
    n3095_o2
  );


  buf

  (
    n483_inv_p,
    n483_inv
  );


  not

  (
    n483_inv_n,
    n483_inv
  );


  buf

  (
    n3170_o2_p,
    n3170_o2
  );


  not

  (
    n3170_o2_n,
    n3170_o2
  );


  buf

  (
    n3171_o2_p,
    n3171_o2
  );


  not

  (
    n3171_o2_n,
    n3171_o2
  );


  buf

  (
    n3172_o2_p,
    n3172_o2
  );


  not

  (
    n3172_o2_n,
    n3172_o2
  );


  buf

  (
    n3179_o2_p,
    n3179_o2
  );


  not

  (
    n3179_o2_n,
    n3179_o2
  );


  buf

  (
    n498_inv_p,
    n498_inv
  );


  not

  (
    n498_inv_n,
    n498_inv
  );


  buf

  (
    n3193_o2_p,
    n3193_o2
  );


  not

  (
    n3193_o2_n,
    n3193_o2
  );


  buf

  (
    n3211_o2_p,
    n3211_o2
  );


  not

  (
    n3211_o2_n,
    n3211_o2
  );


  buf

  (
    n3212_o2_p,
    n3212_o2
  );


  not

  (
    n3212_o2_n,
    n3212_o2
  );


  buf

  (
    n3213_o2_p,
    n3213_o2
  );


  not

  (
    n3213_o2_n,
    n3213_o2
  );


  buf

  (
    n513_inv_p,
    n513_inv
  );


  not

  (
    n513_inv_n,
    n513_inv
  );


  buf

  (
    n1125_o2_p,
    n1125_o2
  );


  not

  (
    n1125_o2_n,
    n1125_o2
  );


  buf

  (
    n1081_o2_p,
    n1081_o2
  );


  not

  (
    n1081_o2_n,
    n1081_o2
  );


  buf

  (
    n1139_o2_p,
    n1139_o2
  );


  not

  (
    n1139_o2_n,
    n1139_o2
  );


  buf

  (
    n3245_o2_p,
    n3245_o2
  );


  not

  (
    n3245_o2_n,
    n3245_o2
  );


  buf

  (
    n3246_o2_p,
    n3246_o2
  );


  not

  (
    n3246_o2_n,
    n3246_o2
  );


  buf

  (
    n3247_o2_p,
    n3247_o2
  );


  not

  (
    n3247_o2_n,
    n3247_o2
  );


  buf

  (
    lo074_buf_o2_p,
    lo074_buf_o2
  );


  not

  (
    lo074_buf_o2_n,
    lo074_buf_o2
  );


  buf

  (
    lo078_buf_o2_p,
    lo078_buf_o2
  );


  not

  (
    lo078_buf_o2_n,
    lo078_buf_o2
  );


  buf

  (
    lo186_buf_o2_p,
    lo186_buf_o2
  );


  not

  (
    lo186_buf_o2_n,
    lo186_buf_o2
  );


  buf

  (
    lo118_buf_o2_p,
    lo118_buf_o2
  );


  not

  (
    lo118_buf_o2_n,
    lo118_buf_o2
  );


  buf

  (
    lo146_buf_o2_p,
    lo146_buf_o2
  );


  not

  (
    lo146_buf_o2_n,
    lo146_buf_o2
  );


  buf

  (
    n1038_o2_p,
    n1038_o2
  );


  not

  (
    n1038_o2_n,
    n1038_o2
  );


  buf

  (
    n1044_o2_p,
    n1044_o2
  );


  not

  (
    n1044_o2_n,
    n1044_o2
  );


  buf

  (
    n555_inv_p,
    n555_inv
  );


  not

  (
    n555_inv_n,
    n555_inv
  );


  buf

  (
    n558_inv_p,
    n558_inv
  );


  not

  (
    n558_inv_n,
    n558_inv
  );


  buf

  (
    lo026_buf_o2_p,
    lo026_buf_o2
  );


  not

  (
    lo026_buf_o2_n,
    lo026_buf_o2
  );


  buf

  (
    lo030_buf_o2_p,
    lo030_buf_o2
  );


  not

  (
    lo030_buf_o2_n,
    lo030_buf_o2
  );


  buf

  (
    lo090_buf_o2_p,
    lo090_buf_o2
  );


  not

  (
    lo090_buf_o2_n,
    lo090_buf_o2
  );


  buf

  (
    lo094_buf_o2_p,
    lo094_buf_o2
  );


  not

  (
    lo094_buf_o2_n,
    lo094_buf_o2
  );


  buf

  (
    lo098_buf_o2_p,
    lo098_buf_o2
  );


  not

  (
    lo098_buf_o2_n,
    lo098_buf_o2
  );


  buf

  (
    lo102_buf_o2_p,
    lo102_buf_o2
  );


  not

  (
    lo102_buf_o2_n,
    lo102_buf_o2
  );


  buf

  (
    lo066_buf_o2_p,
    lo066_buf_o2
  );


  not

  (
    lo066_buf_o2_n,
    lo066_buf_o2
  );


  buf

  (
    lo070_buf_o2_p,
    lo070_buf_o2
  );


  not

  (
    lo070_buf_o2_n,
    lo070_buf_o2
  );


  buf

  (
    n1202_o2_p,
    n1202_o2
  );


  not

  (
    n1202_o2_n,
    n1202_o2
  );


  buf

  (
    n1003_o2_p,
    n1003_o2
  );


  not

  (
    n1003_o2_n,
    n1003_o2
  );


  buf

  (
    n1031_o2_p,
    n1031_o2
  );


  not

  (
    n1031_o2_n,
    n1031_o2
  );


  buf

  (
    n1034_o2_p,
    n1034_o2
  );


  not

  (
    n1034_o2_n,
    n1034_o2
  );


  buf

  (
    n1040_o2_p,
    n1040_o2
  );


  not

  (
    n1040_o2_n,
    n1040_o2
  );


  buf

  (
    n1046_o2_p,
    n1046_o2
  );


  not

  (
    n1046_o2_n,
    n1046_o2
  );


  buf

  (
    n1380_o2_p,
    n1380_o2
  );


  not

  (
    n1380_o2_n,
    n1380_o2
  );


  buf

  (
    n1425_o2_p,
    n1425_o2
  );


  not

  (
    n1425_o2_n,
    n1425_o2
  );


  buf

  (
    n697_o2_p,
    n697_o2
  );


  not

  (
    n697_o2_n,
    n697_o2
  );


  buf

  (
    n1143_o2_p,
    n1143_o2
  );


  not

  (
    n1143_o2_n,
    n1143_o2
  );


  buf

  (
    n673_o2_p,
    n673_o2
  );


  not

  (
    n673_o2_n,
    n673_o2
  );


  buf

  (
    n789_o2_p,
    n789_o2
  );


  not

  (
    n789_o2_n,
    n789_o2
  );


  buf

  (
    n786_o2_p,
    n786_o2
  );


  not

  (
    n786_o2_n,
    n786_o2
  );


  buf

  (
    n1047_o2_p,
    n1047_o2
  );


  not

  (
    n1047_o2_n,
    n1047_o2
  );


  buf

  (
    n1036_o2_p,
    n1036_o2
  );


  not

  (
    n1036_o2_n,
    n1036_o2
  );


  buf

  (
    n1307_o2_p,
    n1307_o2
  );


  not

  (
    n1307_o2_n,
    n1307_o2
  );


  buf

  (
    n1035_o2_p,
    n1035_o2
  );


  not

  (
    n1035_o2_n,
    n1035_o2
  );


  buf

  (
    n1297_o2_p,
    n1297_o2
  );


  not

  (
    n1297_o2_n,
    n1297_o2
  );


  buf

  (
    n1099_o2_p,
    n1099_o2
  );


  not

  (
    n1099_o2_n,
    n1099_o2
  );


  buf

  (
    n1128_o2_p,
    n1128_o2
  );


  not

  (
    n1128_o2_n,
    n1128_o2
  );


  buf

  (
    n645_inv_p,
    n645_inv
  );


  not

  (
    n645_inv_n,
    n645_inv
  );


  buf

  (
    n826_o2_p,
    n826_o2
  );


  not

  (
    n826_o2_n,
    n826_o2
  );


  buf

  (
    n853_o2_p,
    n853_o2
  );


  not

  (
    n853_o2_n,
    n853_o2
  );


  buf

  (
    n654_inv_p,
    n654_inv
  );


  not

  (
    n654_inv_n,
    n654_inv
  );


  buf

  (
    n700_o2_p,
    n700_o2
  );


  not

  (
    n700_o2_n,
    n700_o2
  );


  buf

  (
    n884_o2_p,
    n884_o2
  );


  not

  (
    n884_o2_n,
    n884_o2
  );


  buf

  (
    lo082_buf_o2_p,
    lo082_buf_o2
  );


  not

  (
    lo082_buf_o2_n,
    lo082_buf_o2
  );


  buf

  (
    lo086_buf_o2_p,
    lo086_buf_o2
  );


  not

  (
    lo086_buf_o2_n,
    lo086_buf_o2
  );


  buf

  (
    n801_o2_p,
    n801_o2
  );


  not

  (
    n801_o2_n,
    n801_o2
  );


  buf

  (
    n840_o2_p,
    n840_o2
  );


  not

  (
    n840_o2_n,
    n840_o2
  );


  buf

  (
    n675_inv_p,
    n675_inv
  );


  not

  (
    n675_inv_n,
    n675_inv
  );


  buf

  (
    lo002_buf_o2_p,
    lo002_buf_o2
  );


  not

  (
    lo002_buf_o2_n,
    lo002_buf_o2
  );


  buf

  (
    lo010_buf_o2_p,
    lo010_buf_o2
  );


  not

  (
    lo010_buf_o2_n,
    lo010_buf_o2
  );


  buf

  (
    lo166_buf_o2_p,
    lo166_buf_o2
  );


  not

  (
    lo166_buf_o2_n,
    lo166_buf_o2
  );


  buf

  (
    lo170_buf_o2_p,
    lo170_buf_o2
  );


  not

  (
    lo170_buf_o2_n,
    lo170_buf_o2
  );


  buf

  (
    n1426_o2_p,
    n1426_o2
  );


  not

  (
    n1426_o2_n,
    n1426_o2
  );


  buf

  (
    n1082_o2_p,
    n1082_o2
  );


  not

  (
    n1082_o2_n,
    n1082_o2
  );


  buf

  (
    n1310_o2_p,
    n1310_o2
  );


  not

  (
    n1310_o2_n,
    n1310_o2
  );


  buf

  (
    n1015_o2_p,
    n1015_o2
  );


  not

  (
    n1015_o2_n,
    n1015_o2
  );


  buf

  (
    n1206_o2_p,
    n1206_o2
  );


  not

  (
    n1206_o2_n,
    n1206_o2
  );


  buf

  (
    n1262_o2_p,
    n1262_o2
  );


  not

  (
    n1262_o2_n,
    n1262_o2
  );


  buf

  (
    n1456_o2_p,
    n1456_o2
  );


  not

  (
    n1456_o2_n,
    n1456_o2
  );


  buf

  (
    n1244_o2_p,
    n1244_o2
  );


  not

  (
    n1244_o2_n,
    n1244_o2
  );


  buf

  (
    n1280_o2_p,
    n1280_o2
  );


  not

  (
    n1280_o2_n,
    n1280_o2
  );


  buf

  (
    n1290_o2_p,
    n1290_o2
  );


  not

  (
    n1290_o2_n,
    n1290_o2
  );


  buf

  (
    n1012_o2_p,
    n1012_o2
  );


  not

  (
    n1012_o2_n,
    n1012_o2
  );


  buf

  (
    n1074_o2_p,
    n1074_o2
  );


  not

  (
    n1074_o2_n,
    n1074_o2
  );


  buf

  (
    n1112_o2_p,
    n1112_o2
  );


  not

  (
    n1112_o2_n,
    n1112_o2
  );


  buf

  (
    n1212_o2_p,
    n1212_o2
  );


  not

  (
    n1212_o2_n,
    n1212_o2
  );


  buf

  (
    n1454_o2_p,
    n1454_o2
  );


  not

  (
    n1454_o2_n,
    n1454_o2
  );


  buf

  (
    n1182_o2_p,
    n1182_o2
  );


  not

  (
    n1182_o2_n,
    n1182_o2
  );


  buf

  (
    n1220_o2_p,
    n1220_o2
  );


  not

  (
    n1220_o2_n,
    n1220_o2
  );


  buf

  (
    n701_o2_p,
    n701_o2
  );


  not

  (
    n701_o2_n,
    n701_o2
  );


  buf

  (
    n744_inv_p,
    n744_inv
  );


  not

  (
    n744_inv_n,
    n744_inv
  );


  buf

  (
    n1282_o2_p,
    n1282_o2
  );


  not

  (
    n1282_o2_n,
    n1282_o2
  );


  buf

  (
    n1144_o2_p,
    n1144_o2
  );


  not

  (
    n1144_o2_n,
    n1144_o2
  );


  buf

  (
    n1278_o2_p,
    n1278_o2
  );


  not

  (
    n1278_o2_n,
    n1278_o2
  );


  buf

  (
    n1459_o2_p,
    n1459_o2
  );


  not

  (
    n1459_o2_n,
    n1459_o2
  );


  buf

  (
    n1324_o2_p,
    n1324_o2
  );


  not

  (
    n1324_o2_n,
    n1324_o2
  );


  buf

  (
    n1288_o2_p,
    n1288_o2
  );


  not

  (
    n1288_o2_n,
    n1288_o2
  );


  buf

  (
    n1271_o2_p,
    n1271_o2
  );


  not

  (
    n1271_o2_n,
    n1271_o2
  );


  buf

  (
    n1132_o2_p,
    n1132_o2
  );


  not

  (
    n1132_o2_n,
    n1132_o2
  );


  buf

  (
    n1231_o2_p,
    n1231_o2
  );


  not

  (
    n1231_o2_n,
    n1231_o2
  );


  buf

  (
    n1462_o2_p,
    n1462_o2
  );


  not

  (
    n1462_o2_n,
    n1462_o2
  );


  buf

  (
    n1482_o2_p,
    n1482_o2
  );


  not

  (
    n1482_o2_n,
    n1482_o2
  );


  buf

  (
    n994_o2_p,
    n994_o2
  );


  not

  (
    n994_o2_n,
    n994_o2
  );


  buf

  (
    n998_o2_p,
    n998_o2
  );


  not

  (
    n998_o2_n,
    n998_o2
  );


  buf

  (
    lo106_buf_o2_p,
    lo106_buf_o2
  );


  not

  (
    lo106_buf_o2_n,
    lo106_buf_o2
  );


  buf

  (
    n769_o2_p,
    n769_o2
  );


  not

  (
    n769_o2_n,
    n769_o2
  );


  buf

  (
    n814_o2_p,
    n814_o2
  );


  not

  (
    n814_o2_n,
    n814_o2
  );


  buf

  (
    n841_o2_p,
    n841_o2
  );


  not

  (
    n841_o2_n,
    n841_o2
  );


  buf

  (
    n867_o2_p,
    n867_o2
  );


  not

  (
    n867_o2_n,
    n867_o2
  );


  buf

  (
    lo006_buf_o2_p,
    lo006_buf_o2
  );


  not

  (
    lo006_buf_o2_n,
    lo006_buf_o2
  );


  buf

  (
    lo014_buf_o2_p,
    lo014_buf_o2
  );


  not

  (
    lo014_buf_o2_n,
    lo014_buf_o2
  );


  buf

  (
    lo022_buf_o2_p,
    lo022_buf_o2
  );


  not

  (
    lo022_buf_o2_n,
    lo022_buf_o2
  );


  buf

  (
    lo042_buf_o2_p,
    lo042_buf_o2
  );


  not

  (
    lo042_buf_o2_n,
    lo042_buf_o2
  );


  buf

  (
    lo046_buf_o2_p,
    lo046_buf_o2
  );


  not

  (
    lo046_buf_o2_n,
    lo046_buf_o2
  );


  buf

  (
    lo050_buf_o2_p,
    lo050_buf_o2
  );


  not

  (
    lo050_buf_o2_n,
    lo050_buf_o2
  );


  buf

  (
    lo054_buf_o2_p,
    lo054_buf_o2
  );


  not

  (
    lo054_buf_o2_n,
    lo054_buf_o2
  );


  buf

  (
    lo130_buf_o2_p,
    lo130_buf_o2
  );


  not

  (
    lo130_buf_o2_n,
    lo130_buf_o2
  );


  buf

  (
    lo134_buf_o2_p,
    lo134_buf_o2
  );


  not

  (
    lo134_buf_o2_n,
    lo134_buf_o2
  );


  buf

  (
    lo154_buf_o2_p,
    lo154_buf_o2
  );


  not

  (
    lo154_buf_o2_n,
    lo154_buf_o2
  );


  buf

  (
    lo174_buf_o2_p,
    lo174_buf_o2
  );


  not

  (
    lo174_buf_o2_n,
    lo174_buf_o2
  );


  buf

  (
    lo178_buf_o2_p,
    lo178_buf_o2
  );


  not

  (
    lo178_buf_o2_n,
    lo178_buf_o2
  );


  buf

  (
    n1007_o2_p,
    n1007_o2
  );


  not

  (
    n1007_o2_n,
    n1007_o2
  );


  buf

  (
    n1294_o2_p,
    n1294_o2
  );


  not

  (
    n1294_o2_n,
    n1294_o2
  );


  buf

  (
    n1084_o2_p,
    n1084_o2
  );


  not

  (
    n1084_o2_n,
    n1084_o2
  );


  buf

  (
    n1399_o2_p,
    n1399_o2
  );


  not

  (
    n1399_o2_n,
    n1399_o2
  );


  buf

  (
    n1311_o2_p,
    n1311_o2
  );


  not

  (
    n1311_o2_n,
    n1311_o2
  );


  buf

  (
    n1392_o2_p,
    n1392_o2
  );


  not

  (
    n1392_o2_n,
    n1392_o2
  );


  buf

  (
    n1102_o2_p,
    n1102_o2
  );


  not

  (
    n1102_o2_n,
    n1102_o2
  );


  buf

  (
    n1041_o2_p,
    n1041_o2
  );


  not

  (
    n1041_o2_n,
    n1041_o2
  );


  buf

  (
    n1298_o2_p,
    n1298_o2
  );


  not

  (
    n1298_o2_n,
    n1298_o2
  );


  buf

  (
    n738_o2_p,
    n738_o2
  );


  not

  (
    n738_o2_n,
    n738_o2
  );


  buf

  (
    n1214_o2_p,
    n1214_o2
  );


  not

  (
    n1214_o2_n,
    n1214_o2
  );


  buf

  (
    n1222_o2_p,
    n1222_o2
  );


  not

  (
    n1222_o2_n,
    n1222_o2
  );


  buf

  (
    n1155_o2_p,
    n1155_o2
  );


  not

  (
    n1155_o2_n,
    n1155_o2
  );


  buf

  (
    n1147_o2_p,
    n1147_o2
  );


  not

  (
    n1147_o2_n,
    n1147_o2
  );


  buf

  (
    n1393_o2_p,
    n1393_o2
  );


  not

  (
    n1393_o2_n,
    n1393_o2
  );


  buf

  (
    n999_o2_p,
    n999_o2
  );


  not

  (
    n999_o2_n,
    n999_o2
  );


  buf

  (
    n1306_o2_p,
    n1306_o2
  );


  not

  (
    n1306_o2_n,
    n1306_o2
  );


  buf

  (
    n1312_o2_p,
    n1312_o2
  );


  not

  (
    n1312_o2_n,
    n1312_o2
  );


  buf

  (
    n1382_o2_p,
    n1382_o2
  );


  not

  (
    n1382_o2_n,
    n1382_o2
  );


  buf

  (
    n1383_o2_p,
    n1383_o2
  );


  not

  (
    n1383_o2_n,
    n1383_o2
  );


  buf

  (
    n1152_o2_p,
    n1152_o2
  );


  not

  (
    n1152_o2_n,
    n1152_o2
  );


  buf

  (
    n1334_o2_p,
    n1334_o2
  );


  not

  (
    n1334_o2_n,
    n1334_o2
  );


  buf

  (
    n1335_o2_p,
    n1335_o2
  );


  not

  (
    n1335_o2_n,
    n1335_o2
  );


  buf

  (
    n906_inv_p,
    n906_inv
  );


  not

  (
    n906_inv_n,
    n906_inv
  );


  buf

  (
    n773_o2_p,
    n773_o2
  );


  not

  (
    n773_o2_n,
    n773_o2
  );


  buf

  (
    lo190_buf_o2_p,
    lo190_buf_o2
  );


  not

  (
    lo190_buf_o2_n,
    lo190_buf_o2
  );


  buf

  (
    n1368_o2_p,
    n1368_o2
  );


  not

  (
    n1368_o2_n,
    n1368_o2
  );


  buf

  (
    n1362_o2_p,
    n1362_o2
  );


  not

  (
    n1362_o2_n,
    n1362_o2
  );


  buf

  (
    n1406_o2_p,
    n1406_o2
  );


  not

  (
    n1406_o2_n,
    n1406_o2
  );


  buf

  (
    n1403_o2_p,
    n1403_o2
  );


  not

  (
    n1403_o2_n,
    n1403_o2
  );


  buf

  (
    n741_o2_p,
    n741_o2
  );


  not

  (
    n741_o2_n,
    n741_o2
  );


  buf

  (
    n1407_o2_p,
    n1407_o2
  );


  not

  (
    n1407_o2_n,
    n1407_o2
  );


  buf

  (
    n1395_o2_p,
    n1395_o2
  );


  not

  (
    n1395_o2_n,
    n1395_o2
  );


  buf

  (
    n1359_o2_p,
    n1359_o2
  );


  not

  (
    n1359_o2_n,
    n1359_o2
  );


  buf

  (
    n1159_o2_p,
    n1159_o2
  );


  not

  (
    n1159_o2_n,
    n1159_o2
  );


  buf

  (
    n1221_o2_p,
    n1221_o2
  );


  not

  (
    n1221_o2_n,
    n1221_o2
  );


  buf

  (
    n945_inv_p,
    n945_inv
  );


  not

  (
    n945_inv_n,
    n945_inv
  );


  buf

  (
    n989_o2_p,
    n989_o2
  );


  not

  (
    n989_o2_n,
    n989_o2
  );


  buf

  (
    n881_o2_p,
    n881_o2
  );


  not

  (
    n881_o2_n,
    n881_o2
  );


  buf

  (
    n1340_o2_p,
    n1340_o2
  );


  not

  (
    n1340_o2_n,
    n1340_o2
  );


  buf

  (
    n1341_o2_p,
    n1341_o2
  );


  not

  (
    n1341_o2_n,
    n1341_o2
  );


  buf

  (
    n906_o2_p,
    n906_o2
  );


  not

  (
    n906_o2_n,
    n906_o2
  );


  buf

  (
    n1388_o2_p,
    n1388_o2
  );


  not

  (
    n1388_o2_n,
    n1388_o2
  );


  buf

  (
    n791_o2_p,
    n791_o2
  );


  not

  (
    n791_o2_n,
    n791_o2
  );


  buf

  (
    n1372_o2_p,
    n1372_o2
  );


  not

  (
    n1372_o2_n,
    n1372_o2
  );


  buf

  (
    n815_o2_p,
    n815_o2
  );


  not

  (
    n815_o2_n,
    n815_o2
  );


  buf

  (
    n868_o2_p,
    n868_o2
  );


  not

  (
    n868_o2_n,
    n868_o2
  );


  buf

  (
    lo018_buf_o2_p,
    lo018_buf_o2
  );


  not

  (
    lo018_buf_o2_n,
    lo018_buf_o2
  );


  buf

  (
    lo138_buf_o2_p,
    lo138_buf_o2
  );


  not

  (
    lo138_buf_o2_n,
    lo138_buf_o2
  );


  buf

  (
    lo158_buf_o2_p,
    lo158_buf_o2
  );


  not

  (
    lo158_buf_o2_n,
    lo158_buf_o2
  );


  buf

  (
    n780_o2_p,
    n780_o2
  );


  not

  (
    n780_o2_n,
    n780_o2
  );


  buf

  (
    n728_o2_p,
    n728_o2
  );


  not

  (
    n728_o2_n,
    n728_o2
  );


  buf

  (
    n993_inv_p,
    n993_inv
  );


  not

  (
    n993_inv_n,
    n993_inv
  );


  buf

  (
    n929_o2_p,
    n929_o2
  );


  not

  (
    n929_o2_n,
    n929_o2
  );


  buf

  (
    n955_o2_p,
    n955_o2
  );


  not

  (
    n955_o2_n,
    n955_o2
  );


  buf

  (
    n938_o2_p,
    n938_o2
  );


  not

  (
    n938_o2_n,
    n938_o2
  );


  buf

  (
    n1117_o2_p,
    n1117_o2
  );


  not

  (
    n1117_o2_n,
    n1117_o2
  );


  buf

  (
    n1121_o2_p,
    n1121_o2
  );


  not

  (
    n1121_o2_n,
    n1121_o2
  );


  buf

  (
    n965_o2_p,
    n965_o2
  );


  not

  (
    n965_o2_n,
    n965_o2
  );


  buf

  (
    n752_o2_p,
    n752_o2
  );


  not

  (
    n752_o2_n,
    n752_o2
  );


  buf

  (
    n753_o2_p,
    n753_o2
  );


  not

  (
    n753_o2_n,
    n753_o2
  );


  buf

  (
    n760_o2_p,
    n760_o2
  );


  not

  (
    n760_o2_n,
    n760_o2
  );


  buf

  (
    n770_o2_p,
    n770_o2
  );


  not

  (
    n770_o2_n,
    n770_o2
  );


  buf

  (
    n923_o2_p,
    n923_o2
  );


  not

  (
    n923_o2_n,
    n923_o2
  );


  buf

  (
    n947_o2_p,
    n947_o2
  );


  not

  (
    n947_o2_n,
    n947_o2
  );


  buf

  (
    n897_o2_p,
    n897_o2
  );


  not

  (
    n897_o2_n,
    n897_o2
  );


  buf

  (
    n919_o2_p,
    n919_o2
  );


  not

  (
    n919_o2_n,
    n919_o2
  );


  buf

  (
    n895_o2_p,
    n895_o2
  );


  not

  (
    n895_o2_n,
    n895_o2
  );


  buf

  (
    n917_o2_p,
    n917_o2
  );


  not

  (
    n917_o2_n,
    n917_o2
  );


  buf

  (
    n751_o2_p,
    n751_o2
  );


  not

  (
    n751_o2_n,
    n751_o2
  );


  buf

  (
    n774_o2_p,
    n774_o2
  );


  not

  (
    n774_o2_n,
    n774_o2
  );


  buf

  (
    lo126_buf_o2_p,
    lo126_buf_o2
  );


  not

  (
    lo126_buf_o2_n,
    lo126_buf_o2
  );


  buf

  (
    lo142_buf_o2_p,
    lo142_buf_o2
  );


  not

  (
    lo142_buf_o2_n,
    lo142_buf_o2
  );


  buf

  (
    lo162_buf_o2_p,
    lo162_buf_o2
  );


  not

  (
    lo162_buf_o2_n,
    lo162_buf_o2
  );


  buf

  (
    n1059_inv_p,
    n1059_inv
  );


  not

  (
    n1059_inv_n,
    n1059_inv
  );


  buf

  (
    n792_o2_p,
    n792_o2
  );


  not

  (
    n792_o2_n,
    n792_o2
  );


  buf

  (
    n869_o2_p,
    n869_o2
  );


  not

  (
    n869_o2_n,
    n869_o2
  );


  buf

  (
    n1068_inv_p,
    n1068_inv
  );


  not

  (
    n1068_inv_n,
    n1068_inv
  );


  buf

  (
    lo024_buf_o2_p,
    lo024_buf_o2
  );


  not

  (
    lo024_buf_o2_n,
    lo024_buf_o2
  );


  buf

  (
    lo028_buf_o2_p,
    lo028_buf_o2
  );


  not

  (
    lo028_buf_o2_n,
    lo028_buf_o2
  );


  buf

  (
    lo088_buf_o2_p,
    lo088_buf_o2
  );


  not

  (
    lo088_buf_o2_n,
    lo088_buf_o2
  );


  buf

  (
    lo092_buf_o2_p,
    lo092_buf_o2
  );


  not

  (
    lo092_buf_o2_n,
    lo092_buf_o2
  );


  buf

  (
    lo096_buf_o2_p,
    lo096_buf_o2
  );


  not

  (
    lo096_buf_o2_n,
    lo096_buf_o2
  );


  buf

  (
    lo100_buf_o2_p,
    lo100_buf_o2
  );


  not

  (
    lo100_buf_o2_n,
    lo100_buf_o2
  );


  buf

  (
    n763_o2_p,
    n763_o2
  );


  not

  (
    n763_o2_n,
    n763_o2
  );


  buf

  (
    n754_o2_p,
    n754_o2
  );


  not

  (
    n754_o2_n,
    n754_o2
  );


  buf

  (
    n755_o2_p,
    n755_o2
  );


  not

  (
    n755_o2_n,
    n755_o2
  );


  buf

  (
    n822_o2_p,
    n822_o2
  );


  not

  (
    n822_o2_n,
    n822_o2
  );


  buf

  (
    n849_o2_p,
    n849_o2
  );


  not

  (
    n849_o2_n,
    n849_o2
  );


  buf

  (
    n777_o2_p,
    n777_o2
  );


  not

  (
    n777_o2_n,
    n777_o2
  );


  buf

  (
    n778_o2_p,
    n778_o2
  );


  not

  (
    n778_o2_n,
    n778_o2
  );


  buf

  (
    n820_o2_p,
    n820_o2
  );


  not

  (
    n820_o2_n,
    n820_o2
  );


  buf

  (
    n846_o2_p,
    n846_o2
  );


  not

  (
    n846_o2_n,
    n846_o2
  );


  buf

  (
    n806_o2_p,
    n806_o2
  );


  not

  (
    n806_o2_n,
    n806_o2
  );


  buf

  (
    n771_o2_p,
    n771_o2
  );


  not

  (
    n771_o2_n,
    n771_o2
  );


  buf

  (
    n854_o2_p,
    n854_o2
  );


  not

  (
    n854_o2_n,
    n854_o2
  );


  buf

  (
    n828_o2_p,
    n828_o2
  );


  not

  (
    n828_o2_n,
    n828_o2
  );


  buf

  (
    lo117_buf_o2_p,
    lo117_buf_o2
  );


  not

  (
    lo117_buf_o2_n,
    lo117_buf_o2
  );


  buf

  (
    lo145_buf_o2_p,
    lo145_buf_o2
  );


  not

  (
    lo145_buf_o2_n,
    lo145_buf_o2
  );


  buf

  (
    n762_o2_p,
    n762_o2
  );


  not

  (
    n762_o2_n,
    n762_o2
  );


  buf

  (
    n805_o2_p,
    n805_o2
  );


  not

  (
    n805_o2_n,
    n805_o2
  );


  buf

  (
    n859_o2_p,
    n859_o2
  );


  not

  (
    n859_o2_n,
    n859_o2
  );


  buf

  (
    n833_o2_p,
    n833_o2
  );


  not

  (
    n833_o2_n,
    n833_o2
  );


  buf

  (
    lo034_buf_o2_p,
    lo034_buf_o2
  );


  not

  (
    lo034_buf_o2_n,
    lo034_buf_o2
  );


  buf

  (
    lo038_buf_o2_p,
    lo038_buf_o2
  );


  not

  (
    lo038_buf_o2_n,
    lo038_buf_o2
  );


  buf

  (
    lo122_buf_o2_p,
    lo122_buf_o2
  );


  not

  (
    lo122_buf_o2_n,
    lo122_buf_o2
  );


  buf

  (
    lo150_buf_o2_p,
    lo150_buf_o2
  );


  not

  (
    lo150_buf_o2_n,
    lo150_buf_o2
  );


  and

  (
    g412_p,
    n2368_o2_n,
    n1860_lo_n_spl_
  );


  and

  (
    g413_p,
    n1776_lo_n_spl_,
    n1752_lo_n_spl_
  );


  or

  (
    g414_n,
    n2148_lo_n_spl_0,
    n1872_lo_p_spl_
  );


  or

  (
    g415_n,
    n2124_lo_n_spl_0,
    n1848_lo_p
  );


  and

  (
    g416_p,
    g415_n,
    g414_n
  );


  or

  (
    g417_n,
    n2100_lo_n_spl_0,
    n1824_lo_p_spl_
  );


  or

  (
    g418_n,
    n2136_lo_n_spl_0,
    n1860_lo_p
  );


  and

  (
    g419_p,
    g418_n,
    g417_n
  );


  and

  (
    g420_p,
    g419_p,
    g416_p
  );


  or

  (
    g421_n,
    n2184_lo_n_spl_0,
    n1908_lo_p_spl_0
  );


  or

  (
    g422_n,
    n2112_lo_n_spl_0,
    n1836_lo_p
  );


  and

  (
    g423_p,
    g422_n,
    g421_n
  );


  or

  (
    g424_n,
    n2160_lo_n_spl_0,
    n1884_lo_p_spl_
  );


  or

  (
    g425_n,
    n2172_lo_n_spl_0,
    n1896_lo_p_spl_0
  );


  and

  (
    g426_p,
    g425_n,
    g424_n
  );


  and

  (
    g427_p,
    g426_p,
    g423_p
  );


  and

  (
    g428_p,
    g427_p,
    g420_p
  );


  or

  (
    g429_n,
    g428_p,
    g413_p
  );


  and

  (
    g430_p,
    n2071_o2_p,
    n1776_lo_n_spl_
  );


  or

  (
    g430_n,
    n2071_o2_n,
    n1776_lo_p
  );


  or

  (
    g431_n,
    g430_n_spl_,
    n698_o2_n
  );


  and

  (
    g432_p,
    n2172_lo_n_spl_0,
    n2160_lo_n_spl_0
  );


  or

  (
    g433_n,
    g432_p,
    n2148_lo_n_spl_0
  );


  or

  (
    g434_n,
    g433_n,
    n2471_o2_p
  );


  and

  (
    g435_p,
    g434_n,
    g431_n
  );


  and

  (
    g436_p,
    g435_p,
    g429_n
  );


  and

  (
    g437_p,
    n2184_lo_n_spl_0,
    n2172_lo_p_spl_
  );


  or

  (
    g437_n,
    n2184_lo_p_spl_,
    n2172_lo_n_spl_1
  );


  and

  (
    g438_p,
    n2184_lo_p_spl_,
    n2172_lo_n_spl_1
  );


  or

  (
    g438_n,
    n2184_lo_n_spl_,
    n2172_lo_p_spl_
  );


  and

  (
    g439_p,
    g438_n,
    g437_n
  );


  or

  (
    g439_n,
    g438_p,
    g437_p
  );


  and

  (
    g440_p,
    n2160_lo_n_spl_1,
    n2148_lo_p_spl_
  );


  or

  (
    g440_n,
    n2160_lo_p_spl_,
    n2148_lo_n_spl_1
  );


  and

  (
    g441_p,
    n2160_lo_p_spl_,
    n2148_lo_n_spl_1
  );


  or

  (
    g441_n,
    n2160_lo_n_spl_1,
    n2148_lo_p_spl_
  );


  and

  (
    g442_p,
    g441_n,
    g440_n
  );


  or

  (
    g442_n,
    g441_p,
    g440_p
  );


  and

  (
    g443_p,
    g442_p_spl_,
    g439_n_spl_
  );


  or

  (
    g443_n,
    g442_n_spl_,
    g439_p_spl_
  );


  and

  (
    g444_p,
    g442_n_spl_,
    g439_p_spl_
  );


  or

  (
    g444_n,
    g442_p_spl_,
    g439_n_spl_
  );


  and

  (
    g445_p,
    g444_n,
    g443_n
  );


  or

  (
    g445_n,
    g444_p,
    g443_p
  );


  and

  (
    g446_p,
    n2136_lo_n_spl_0,
    n2124_lo_p_spl_
  );


  or

  (
    g446_n,
    n2136_lo_p_spl_,
    n2124_lo_n_spl_0
  );


  and

  (
    g447_p,
    n2136_lo_p_spl_,
    n2124_lo_n_spl_
  );


  or

  (
    g447_n,
    n2136_lo_n_spl_,
    n2124_lo_p_spl_
  );


  and

  (
    g448_p,
    g447_n,
    g446_n
  );


  or

  (
    g448_n,
    g447_p,
    g446_p
  );


  and

  (
    g449_p,
    n2112_lo_n_spl_0,
    n2100_lo_p_spl_
  );


  or

  (
    g449_n,
    n2112_lo_p_spl_,
    n2100_lo_n_spl_0
  );


  and

  (
    g450_p,
    n2112_lo_p_spl_,
    n2100_lo_n_spl_
  );


  or

  (
    g450_n,
    n2112_lo_n_spl_,
    n2100_lo_p_spl_
  );


  and

  (
    g451_p,
    g450_n,
    g449_n
  );


  or

  (
    g451_n,
    g450_p,
    g449_p
  );


  and

  (
    g452_p,
    g451_n_spl_,
    g448_p_spl_
  );


  or

  (
    g452_n,
    g451_p_spl_,
    g448_n_spl_
  );


  and

  (
    g453_p,
    g451_p_spl_,
    g448_n_spl_
  );


  or

  (
    g453_n,
    g451_n_spl_,
    g448_p_spl_
  );


  and

  (
    g454_p,
    g453_n,
    g452_n
  );


  or

  (
    g454_n,
    g453_p,
    g452_p
  );


  or

  (
    g455_n,
    g454_p,
    g445_p
  );


  or

  (
    g456_n,
    g454_n,
    g445_n
  );


  and

  (
    g457_p,
    g456_n,
    g455_n
  );


  and

  (
    g458_p,
    n1884_lo_p_spl_,
    n1872_lo_p_spl_
  );


  or

  (
    g458_n,
    n1884_lo_n,
    n1872_lo_n
  );


  and

  (
    g459_p,
    g458_n,
    n2080_o2_p
  );


  or

  (
    g459_n,
    g458_p,
    n2080_o2_n
  );


  and

  (
    g460_p,
    n1908_lo_n_spl_0,
    n1896_lo_p_spl_0
  );


  or

  (
    g460_n,
    n1908_lo_p_spl_0,
    n1896_lo_n_spl_
  );


  and

  (
    g461_p,
    n1908_lo_p_spl_,
    n1896_lo_n_spl_
  );


  or

  (
    g461_n,
    n1908_lo_n_spl_0,
    n1896_lo_p_spl_
  );


  and

  (
    g462_p,
    g461_n,
    g460_n
  );


  or

  (
    g462_n,
    g461_p,
    g460_p
  );


  and

  (
    g463_p,
    g462_p_spl_,
    g459_p_spl_
  );


  or

  (
    g463_n,
    g462_n_spl_,
    g459_n_spl_
  );


  and

  (
    g464_p,
    g462_n_spl_,
    g459_n_spl_
  );


  or

  (
    g464_n,
    g462_p_spl_,
    g459_p_spl_
  );


  and

  (
    g465_p,
    g464_n,
    g463_n
  );


  or

  (
    g465_n,
    g464_p,
    g463_p
  );


  and

  (
    g466_p,
    g465_n,
    n744_o2_n
  );


  and

  (
    g467_p,
    g465_p,
    n744_o2_p
  );


  or

  (
    g468_n,
    g467_p,
    g466_p
  );


  and

  (
    g469_p,
    n3029_o2_p_spl_,
    n2617_o2_p
  );


  and

  (
    g470_p,
    n3029_o2_p_spl_,
    n2765_o2_p
  );


  or

  (
    g471_n,
    g470_p,
    n3153_o2_p
  );


  and

  (
    g472_p,
    n1001_o2_n_spl_0,
    n698_o2_p
  );


  and

  (
    g473_p,
    n2829_o2_p,
    n1752_lo_n_spl_
  );


  or

  (
    g474_n,
    g473_p,
    g472_p
  );


  and

  (
    g475_p,
    n1012_o2_n,
    n1010_o2_n_spl_
  );


  or

  (
    g475_n,
    n1012_o2_p,
    n1010_o2_p_spl_
  );


  and

  (
    g476_p,
    n1074_o2_p,
    n1015_o2_n
  );


  or

  (
    g476_n,
    n1074_o2_n,
    n1015_o2_p
  );


  and

  (
    g477_p,
    g476_n,
    g475_n
  );


  or

  (
    g477_n,
    g476_p,
    g475_p
  );


  and

  (
    g478_p,
    n1112_o2_p,
    n1082_o2_n
  );


  or

  (
    g478_n,
    n1112_o2_n,
    n1082_o2_p
  );


  and

  (
    g479_p,
    n1132_o2_p,
    n1010_o2_n_spl_
  );


  or

  (
    g479_n,
    n1132_o2_n,
    n1010_o2_p_spl_
  );


  and

  (
    g480_p,
    g479_n,
    g478_n
  );


  or

  (
    g480_n,
    g479_p,
    g478_p
  );


  and

  (
    g481_p,
    n3035_o2_p,
    n2775_o2_p
  );


  or

  (
    g481_n,
    n3035_o2_n,
    n2775_o2_n
  );


  and

  (
    g482_p,
    g481_n_spl_,
    n3119_o2_p_spl_
  );


  or

  (
    g482_n,
    g481_p_spl_,
    n3119_o2_n_spl_
  );


  and

  (
    g483_p,
    g481_p_spl_,
    n3119_o2_n_spl_
  );


  or

  (
    g483_n,
    g481_n_spl_,
    n3119_o2_p_spl_
  );


  and

  (
    g484_p,
    g483_n,
    g482_n
  );


  or

  (
    g484_n,
    g483_p,
    g482_p
  );


  and

  (
    g485_p,
    g484_n,
    n2304_lo_p
  );


  or

  (
    g485_n,
    g484_p,
    n2304_lo_n
  );


  and

  (
    g486_p,
    n1153_o2_p_spl_,
    n1160_o2_p_spl_
  );


  or

  (
    g486_n,
    n1153_o2_n_spl_,
    n1160_o2_n_spl_
  );


  and

  (
    g487_p,
    n1153_o2_n_spl_,
    n1160_o2_n_spl_
  );


  or

  (
    g487_n,
    n1153_o2_p_spl_,
    n1160_o2_p_spl_
  );


  and

  (
    g488_p,
    g487_n,
    g486_n
  );


  or

  (
    g488_n,
    g487_p,
    g486_p
  );


  and

  (
    g489_p,
    g488_p,
    g485_p
  );


  and

  (
    g490_p,
    g488_n,
    g485_n
  );


  or

  (
    g491_n,
    g490_p,
    g489_p
  );


  and

  (
    g492_p,
    g430_n_spl_,
    n2405_o2_p
  );


  and

  (
    g493_p,
    g492_p,
    g491_n
  );


  and

  (
    g494_p,
    g430_p,
    n1908_lo_n_spl_
  );


  and

  (
    g495_p,
    g494_p,
    n2137_o2_n
  );


  and

  (
    g496_p,
    n2383_o2_n,
    n1860_lo_n_spl_
  );


  or

  (
    g497_n,
    g496_p,
    n1824_lo_p_spl_
  );


  or

  (
    g498_n,
    n1848_lo_n,
    n1824_lo_n
  );


  and

  (
    g499_p,
    g498_n,
    n2405_o2_n
  );


  and

  (
    g500_p,
    g499_p,
    g497_n
  );


  or

  (
    g501_n,
    g500_p,
    g495_p
  );


  or

  (
    g502_n,
    g501_n,
    g493_p
  );


  and

  (
    g503_p,
    n1182_o2_n,
    n1212_o2_p
  );


  or

  (
    g503_n,
    n1182_o2_p,
    n1212_o2_n
  );


  and

  (
    g504_p,
    n1231_o2_p,
    n1244_o2_n
  );


  or

  (
    g504_n,
    n1231_o2_n,
    n1244_o2_p
  );


  and

  (
    g505_p,
    g504_n,
    g503_n
  );


  or

  (
    g505_n,
    g504_p,
    g503_p
  );


  and

  (
    g506_p,
    n1282_o2_p,
    n1001_o2_n_spl_0
  );


  or

  (
    g506_n,
    n1282_o2_n,
    n1001_o2_p_spl_
  );


  and

  (
    g507_p,
    n1278_o2_n,
    n1280_o2_n
  );


  or

  (
    g507_n,
    n1278_o2_p,
    n1280_o2_p
  );


  and

  (
    g508_p,
    g507_p,
    g506_n
  );


  or

  (
    g508_n,
    g507_n,
    g506_p
  );


  and

  (
    g509_p,
    n1288_o2_p,
    n1001_o2_n_spl_
  );


  or

  (
    g509_n,
    n1288_o2_n,
    n1001_o2_p_spl_
  );


  and

  (
    g510_p,
    n1324_o2_n,
    n1290_o2_n
  );


  or

  (
    g510_n,
    n1324_o2_p,
    n1290_o2_p
  );


  and

  (
    g511_p,
    g510_p,
    g509_n
  );


  or

  (
    g511_n,
    g510_n,
    g509_p
  );


  and

  (
    g512_p,
    n1454_o2_p,
    n1426_o2_n
  );


  or

  (
    g512_n,
    n1454_o2_n,
    n1426_o2_p
  );


  and

  (
    g513_p,
    n1459_o2_p,
    n1456_o2_n
  );


  or

  (
    g513_n,
    n1459_o2_n,
    n1456_o2_p
  );


  and

  (
    g514_p,
    g513_n,
    g512_n
  );


  or

  (
    g514_n,
    g513_p,
    g512_p
  );


  and

  (
    g515_p,
    g514_p_spl_,
    g480_p_spl_
  );


  or

  (
    g515_n,
    g514_n_spl_0,
    g480_n_spl_0
  );


  and

  (
    g516_p,
    g511_p_spl_,
    g505_p_spl_
  );


  or

  (
    g516_n,
    g511_n_spl_0,
    g505_n_spl_0
  );


  and

  (
    g517_p,
    g508_p_spl_,
    g477_p_spl_
  );


  or

  (
    g517_n,
    g508_n_spl_0,
    g477_n_spl_0
  );


  or

  (
    g518_n,
    g517_n_spl_,
    g516_n_spl_
  );


  or

  (
    g519_n,
    g518_n,
    g515_n_spl_
  );


  or

  (
    g520_n,
    g519_n,
    n1462_o2_p_spl_0
  );


  and

  (
    g521_p,
    n2316_lo_p,
    n2064_lo_p_spl_
  );


  or

  (
    g521_n,
    n2316_lo_n,
    n2064_lo_n
  );


  or

  (
    g522_n,
    g521_n_spl_,
    n1462_o2_p_spl_0
  );


  and

  (
    g523_p,
    g522_n,
    n2064_lo_p_spl_
  );


  and

  (
    g524_p,
    g523_p,
    g520_n_spl_
  );


  and

  (
    g525_p,
    g508_n_spl_0,
    g477_n_spl_0
  );


  or

  (
    g525_n,
    g508_p_spl_,
    g477_p_spl_
  );


  and

  (
    g526_p,
    g525_n,
    g517_n_spl_
  );


  or

  (
    g526_n,
    g525_p,
    g517_p
  );


  and

  (
    g527_p,
    g511_n_spl_0,
    g505_n_spl_0
  );


  or

  (
    g527_n,
    g511_p_spl_,
    g505_p_spl_
  );


  and

  (
    g528_p,
    g527_n,
    g516_n_spl_
  );


  or

  (
    g528_n,
    g527_p,
    g516_p
  );


  and

  (
    g529_p,
    g528_n_spl_,
    g526_p_spl_
  );


  or

  (
    g529_n,
    g528_p_spl_,
    g526_n_spl_
  );


  and

  (
    g530_p,
    g528_p_spl_,
    g526_n_spl_
  );


  or

  (
    g530_n,
    g528_n_spl_,
    g526_p_spl_
  );


  and

  (
    g531_p,
    g530_n,
    g529_n
  );


  or

  (
    g531_n,
    g530_p,
    g529_p
  );


  and

  (
    g532_p,
    g514_n_spl_0,
    g480_n_spl_0
  );


  or

  (
    g532_n,
    g514_p_spl_,
    g480_p_spl_
  );


  and

  (
    g533_p,
    g532_n,
    g515_n_spl_
  );


  or

  (
    g533_n,
    g532_p,
    g515_p
  );


  and

  (
    g534_p,
    n1482_o2_n,
    n1462_o2_p_spl_
  );


  or

  (
    g534_n,
    n1482_o2_p,
    n1462_o2_n
  );


  and

  (
    g535_p,
    g534_n_spl_0,
    n2340_lo_p_spl_
  );


  or

  (
    g535_n,
    g534_p_spl_0,
    n2340_lo_n_spl_
  );


  and

  (
    g536_p,
    g534_p_spl_0,
    n2340_lo_n_spl_
  );


  or

  (
    g536_n,
    g534_n_spl_0,
    n2340_lo_p_spl_
  );


  and

  (
    g537_p,
    g536_n,
    g535_n
  );


  or

  (
    g537_n,
    g536_p,
    g535_p
  );


  and

  (
    g538_p,
    g537_n,
    g521_n_spl_
  );


  or

  (
    g538_n,
    g537_p,
    g521_p
  );


  and

  (
    g539_p,
    g538_p_spl_,
    g533_p_spl_0
  );


  or

  (
    g539_n,
    g538_n_spl_,
    g533_n_spl_0
  );


  and

  (
    g540_p,
    g538_n_spl_,
    g533_n_spl_0
  );


  or

  (
    g540_n,
    g538_p_spl_,
    g533_p_spl_0
  );


  and

  (
    g541_p,
    g540_n,
    g539_n
  );


  or

  (
    g541_n,
    g540_p,
    g539_p
  );


  and

  (
    g542_p,
    g541_n,
    g531_n_spl_
  );


  and

  (
    g543_p,
    g541_p,
    g531_p_spl_
  );


  or

  (
    g544_n,
    g543_p,
    g542_p
  );


  and

  (
    g545_p,
    g534_n_spl_1,
    g533_n_spl_1
  );


  or

  (
    g545_n,
    g534_p_spl_1,
    g533_p_spl_1
  );


  and

  (
    g546_p,
    g534_p_spl_1,
    g533_p_spl_1
  );


  or

  (
    g546_n,
    g534_n_spl_1,
    g533_n_spl_1
  );


  and

  (
    g547_p,
    g546_n,
    g545_n
  );


  or

  (
    g547_n,
    g546_p,
    g545_p
  );


  or

  (
    g548_n,
    g547_p,
    g531_p_spl_
  );


  or

  (
    g549_n,
    g547_n,
    g531_n_spl_
  );


  and

  (
    g550_p,
    g549_n,
    g548_n
  );


  or

  (
    g551_n,
    n2859_o2_n,
    n2793_o2_p_spl_0
  );


  or

  (
    g552_n,
    n2659_o2_n,
    n2621_o2_n_spl_
  );


  and

  (
    g553_p,
    n999_o2_p,
    n994_o2_n_spl_0
  );


  or

  (
    g553_n,
    n999_o2_n,
    n994_o2_p_spl_
  );


  and

  (
    g554_p,
    n1159_o2_n,
    n1155_o2_n
  );


  or

  (
    g554_n,
    n1159_o2_p,
    n1155_o2_p
  );


  and

  (
    g555_p,
    n945_inv_n,
    n1152_o2_p
  );


  or

  (
    g555_n,
    n945_inv_p_spl_,
    n1152_o2_n
  );


  and

  (
    g556_p,
    n3028_o2_n_spl_,
    n2643_o2_p
  );


  or

  (
    g556_n,
    n3028_o2_p_spl_0,
    n2643_o2_n
  );


  and

  (
    g557_p,
    n741_o2_n,
    n738_o2_p
  );


  and

  (
    g558_p,
    n741_o2_p,
    n738_o2_n
  );


  or

  (
    g559_n,
    g558_p,
    g557_p
  );


  and

  (
    g560_p,
    n1007_o2_n,
    n2620_o2_p_spl_
  );


  or

  (
    g560_n,
    n1007_o2_p_spl_,
    n2620_o2_n_spl_
  );


  and

  (
    g561_p,
    g560_n,
    n2579_o2_n
  );


  or

  (
    g561_n,
    g560_p,
    n2579_o2_p_spl_
  );


  and

  (
    g562_p,
    g561_p_spl_,
    g556_p_spl_0
  );


  or

  (
    g562_n,
    g561_n_spl_00,
    g556_n_spl_0
  );


  and

  (
    g563_p,
    n869_o2_p_spl_,
    n792_o2_p_spl_
  );


  or

  (
    g563_n,
    n869_o2_n_spl_,
    n792_o2_n_spl_
  );


  and

  (
    g564_p,
    n1121_o2_n,
    n1117_o2_n
  );


  or

  (
    g564_n,
    n1121_o2_p,
    n1117_o2_p
  );


  and

  (
    g565_p,
    g564_p,
    n1059_inv_n_spl_000
  );


  or

  (
    g565_n,
    g564_n,
    n1059_inv_p_spl_000
  );


  and

  (
    g566_p,
    g563_p_spl_,
    n1059_inv_p_spl_000
  );


  or

  (
    g566_n,
    g563_n,
    n1059_inv_n_spl_000
  );


  and

  (
    g567_p,
    g566_n,
    g565_n
  );


  or

  (
    g567_n,
    g566_p,
    g565_p
  );


  and

  (
    g568_p,
    n895_o2_p,
    n897_o2_n_spl_0
  );


  or

  (
    g568_n,
    n895_o2_n,
    n897_o2_p_spl_
  );


  and

  (
    g569_p,
    n1059_inv_p_spl_001,
    n881_o2_p
  );


  or

  (
    g569_n,
    n1059_inv_n_spl_001,
    n881_o2_n
  );


  and

  (
    g570_p,
    g569_n_spl_,
    g568_n_spl_0
  );


  or

  (
    g570_n,
    g569_p_spl_,
    g568_p_spl_
  );


  and

  (
    g571_p,
    g569_p_spl_,
    g568_p_spl_
  );


  or

  (
    g571_n,
    g569_n_spl_,
    g568_n_spl_0
  );


  and

  (
    g572_p,
    g571_n,
    g570_n
  );


  or

  (
    g572_n,
    g571_p,
    g570_p
  );


  and

  (
    g573_p,
    n917_o2_p,
    n919_o2_n_spl_0
  );


  or

  (
    g573_n,
    n917_o2_n,
    n919_o2_p_spl_
  );


  and

  (
    g574_p,
    n1059_inv_p_spl_001,
    n906_o2_p
  );


  or

  (
    g574_n,
    n1059_inv_n_spl_001,
    n906_o2_n
  );


  and

  (
    g575_p,
    g574_n_spl_,
    g573_n_spl_0
  );


  or

  (
    g575_n,
    g574_p_spl_,
    g573_p_spl_
  );


  and

  (
    g576_p,
    g574_p_spl_,
    g573_p_spl_
  );


  or

  (
    g576_n,
    g574_n_spl_,
    g573_n_spl_0
  );


  and

  (
    g577_p,
    g576_n,
    g575_n
  );


  or

  (
    g577_n,
    g576_p,
    g575_p
  );


  and

  (
    g578_p,
    lo094_buf_o2_p,
    n2993_o2_p_spl_00
  );


  or

  (
    g578_n,
    lo094_buf_o2_n,
    n2993_o2_n_spl_0
  );


  and

  (
    g579_p,
    lo098_buf_o2_p,
    n2993_o2_p_spl_00
  );


  or

  (
    g579_n,
    lo098_buf_o2_n,
    n2993_o2_n_spl_0
  );


  or

  (
    g580_n,
    g579_p_spl_00,
    lo102_buf_o2_n_spl_
  );


  or

  (
    g581_n,
    g580_n,
    g578_p_spl_0
  );


  or

  (
    g582_n,
    g579_p_spl_00,
    lo102_buf_o2_p_spl_
  );


  or

  (
    g583_n,
    g582_n,
    g578_p_spl_0
  );


  and

  (
    g584_p,
    n869_o2_p_spl_,
    n791_o2_p
  );


  or

  (
    g584_n,
    n869_o2_n_spl_,
    n791_o2_n_spl_
  );


  and

  (
    g585_p,
    n868_o2_p,
    n814_o2_p_spl_
  );


  or

  (
    g585_n,
    n868_o2_n,
    n814_o2_n
  );


  and

  (
    g586_p,
    n841_o2_p_spl_,
    n675_inv_p_spl_
  );


  or

  (
    g586_n,
    n841_o2_n,
    n675_inv_n
  );


  and

  (
    g587_p,
    g586_n,
    n840_o2_n
  );


  or

  (
    g587_n,
    g586_p,
    n840_o2_p
  );


  and

  (
    g588_p,
    g587_p,
    g585_n
  );


  or

  (
    g588_n,
    g587_n,
    g585_p
  );


  and

  (
    g589_p,
    g588_p,
    g584_n
  );


  or

  (
    g589_n,
    g588_n,
    g584_p
  );


  and

  (
    g590_p,
    g572_p_spl_0,
    g567_p_spl_0
  );


  or

  (
    g590_n,
    g572_n,
    g567_n
  );


  or

  (
    g591_n,
    lo026_buf_o2_n_spl_,
    n1962_lo_p_spl_0
  );


  and

  (
    g592_p,
    g589_n_spl_,
    n1059_inv_n_spl_01
  );


  or

  (
    g592_n,
    g589_p,
    n1059_inv_p_spl_010
  );


  and

  (
    g593_p,
    lo102_buf_o2_p_spl_,
    n2993_o2_p_spl_0
  );


  or

  (
    g593_n,
    lo102_buf_o2_n_spl_,
    n2993_o2_n_spl_
  );


  and

  (
    g594_p,
    g593_n_spl_,
    g578_n_spl_
  );


  or

  (
    g594_n,
    g593_p_spl_,
    g578_p_spl_1
  );


  and

  (
    g595_p,
    g594_p_spl_,
    g579_n_spl_0
  );


  or

  (
    g595_n,
    g594_n_spl_,
    g579_p_spl_01
  );


  and

  (
    g596_p,
    g593_p_spl_,
    g578_n_spl_
  );


  or

  (
    g596_n,
    g593_n_spl_,
    g578_p_spl_1
  );


  and

  (
    g597_p,
    g596_p_spl_,
    g579_p_spl_01
  );


  or

  (
    g597_n,
    g596_n_spl_,
    g579_n_spl_0
  );


  and

  (
    g598_p,
    g594_p_spl_,
    g579_p_spl_1
  );


  or

  (
    g598_n,
    g594_n_spl_,
    g579_n_spl_1
  );


  and

  (
    g599_p,
    g596_p_spl_,
    g579_n_spl_1
  );


  or

  (
    g599_n,
    g596_n_spl_,
    g579_p_spl_1
  );


  and

  (
    g600_p,
    n1335_o2_n,
    n1334_o2_n_spl_
  );


  or

  (
    g600_n,
    n1335_o2_p,
    n1334_o2_p_spl_
  );


  and

  (
    g601_p,
    n1341_o2_n,
    n1340_o2_p
  );


  or

  (
    g601_n,
    n1341_o2_p,
    n1340_o2_n
  );


  and

  (
    g602_p,
    n1147_o2_p_spl_,
    lo186_buf_o2_p_spl_0
  );


  or

  (
    g602_n,
    n1147_o2_n,
    lo186_buf_o2_n_spl_0
  );


  and

  (
    g603_p,
    g602_p,
    g555_n
  );


  or

  (
    g603_n,
    g602_n,
    g555_p_spl_
  );


  and

  (
    g604_p,
    g603_n_spl_,
    g601_n_spl_0
  );


  or

  (
    g604_n,
    g603_p_spl_,
    g601_p_spl_
  );


  and

  (
    g605_p,
    g604_n_spl_,
    g600_p
  );


  and

  (
    g606_p,
    g604_p,
    g600_n_spl_0
  );


  or

  (
    g607_n,
    g606_p,
    g605_p
  );


  and

  (
    g608_p,
    g607_n,
    g556_n_spl_0
  );


  or

  (
    g609_n,
    n2619_o2_n_spl_00,
    n2618_o2_p
  );


  or

  (
    g610_n,
    g609_n_spl_0,
    n1143_o2_n
  );


  and

  (
    g611_p,
    n2795_o2_n,
    n2580_o2_p_spl_
  );


  or

  (
    g611_n,
    n2795_o2_p,
    n2580_o2_n
  );


  and

  (
    g612_p,
    g611_n,
    n327_inv_p_spl_
  );


  or

  (
    g612_n,
    g611_p,
    n327_inv_n
  );


  or

  (
    g613_n,
    n1359_o2_p,
    n1362_o2_n
  );


  or

  (
    g614_n,
    n1372_o2_n,
    n1368_o2_n
  );


  and

  (
    g615_p,
    g614_n,
    g613_n
  );


  or

  (
    g616_n,
    g615_p,
    g612_p_spl_00
  );


  and

  (
    g617_p,
    g616_n,
    g562_p_spl_00
  );


  and

  (
    g618_p,
    g617_p,
    g610_n
  );


  and

  (
    g619_p,
    g600_n_spl_0,
    g561_n_spl_00
  );


  or

  (
    g620_n,
    g619_p,
    g618_p
  );


  or

  (
    g621_n,
    g620_n,
    g608_p
  );


  and

  (
    g622_p,
    n1383_o2_n,
    n1382_o2_p
  );


  or

  (
    g622_n,
    n1383_o2_p,
    n1382_o2_n
  );


  or

  (
    g623_n,
    g622_n_spl_0,
    g609_n_spl_0
  );


  or

  (
    g624_n,
    n1388_o2_p,
    n1393_o2_p
  );


  or

  (
    g625_n,
    n1395_o2_p,
    n1392_o2_n
  );


  or

  (
    g626_n,
    g625_n,
    g624_n
  );


  or

  (
    g627_n,
    n1403_o2_n,
    n1399_o2_n
  );


  or

  (
    g628_n,
    n1407_o2_n,
    n1406_o2_n
  );


  or

  (
    g629_n,
    g628_n,
    g627_n
  );


  and

  (
    g630_p,
    g629_n,
    g626_n
  );


  or

  (
    g631_n,
    g630_p,
    g612_p_spl_00
  );


  and

  (
    g632_p,
    g631_n,
    g562_p_spl_00
  );


  and

  (
    g633_p,
    g632_p,
    g623_n
  );


  and

  (
    g634_p,
    g622_n_spl_0,
    g554_n_spl_0
  );


  or

  (
    g634_n,
    g622_p_spl_,
    g554_p_spl_
  );


  and

  (
    g635_p,
    g622_p_spl_,
    g554_p_spl_
  );


  or

  (
    g635_n,
    g622_n_spl_,
    g554_n_spl_0
  );


  and

  (
    g636_p,
    g635_n,
    g634_n
  );


  or

  (
    g636_n,
    g635_p,
    g634_p
  );


  and

  (
    g637_p,
    g636_n,
    n1334_o2_n_spl_
  );


  and

  (
    g638_p,
    g636_p,
    n1334_o2_p_spl_
  );


  or

  (
    g639_n,
    g638_p,
    g637_p
  );


  and

  (
    g640_p,
    g601_n_spl_0,
    g600_n_spl_
  );


  or

  (
    g641_n,
    g640_p,
    g603_n_spl_
  );


  and

  (
    g642_p,
    g641_n,
    g556_n_spl_1
  );


  or

  (
    g643_n,
    g642_p,
    g561_n_spl_01
  );


  and

  (
    g644_p,
    g643_n,
    g639_n
  );


  or

  (
    g645_n,
    g644_p,
    g633_p
  );


  or

  (
    g646_n,
    lo034_buf_o2_p_spl_00,
    lo028_buf_o2_p_spl_0
  );


  and

  (
    g647_p,
    n965_o2_n_spl_,
    n786_o2_p
  );


  or

  (
    g647_n,
    n965_o2_p_spl_,
    n786_o2_n_spl_
  );


  and

  (
    g648_p,
    n947_o2_n,
    n955_o2_n
  );


  or

  (
    g648_n,
    n947_o2_p,
    n955_o2_p
  );


  and

  (
    g649_p,
    g648_p_spl_0,
    g647_n
  );


  or

  (
    g649_n,
    g648_n_spl_0,
    g647_p
  );


  and

  (
    g650_p,
    n965_o2_n_spl_,
    n789_o2_p_spl_
  );


  or

  (
    g650_n,
    n965_o2_p_spl_,
    n789_o2_n_spl_
  );


  and

  (
    g651_p,
    g650_p,
    g648_n_spl_0
  );


  or

  (
    g651_n,
    g650_n,
    g648_p_spl_0
  );


  and

  (
    g652_p,
    g651_n_spl_,
    g649_n
  );


  or

  (
    g652_n,
    g651_p_spl_,
    g649_p
  );


  and

  (
    g653_p,
    g648_n_spl_,
    n989_o2_p
  );


  or

  (
    g653_n,
    g648_p_spl_,
    n989_o2_n_spl_0
  );


  and

  (
    g654_p,
    g653_n_spl_,
    g652_n_spl_0
  );


  or

  (
    g654_n,
    g653_p_spl_,
    g652_p_spl_
  );


  and

  (
    g655_p,
    g653_p_spl_,
    g652_p_spl_
  );


  or

  (
    g655_n,
    g653_n_spl_,
    g652_n_spl_0
  );


  and

  (
    g656_p,
    g655_n,
    g654_n
  );


  or

  (
    g656_n,
    g655_p,
    g654_p
  );


  or

  (
    g657_n,
    lo028_buf_o2_p_spl_0,
    lo024_buf_o2_p_spl_0
  );


  and

  (
    g658_p,
    lo092_buf_o2_n_spl_,
    lo088_buf_o2_n
  );


  or

  (
    g658_n,
    lo092_buf_o2_p_spl_0,
    lo088_buf_o2_p_spl_
  );


  or

  (
    g659_n,
    lo100_buf_o2_p_spl_,
    lo096_buf_o2_p_spl_
  );


  and

  (
    g660_p,
    g599_n_spl_0,
    n3089_o2_n_spl_
  );


  or

  (
    g661_n,
    g597_p_spl_0,
    n3091_o2_p_spl_
  );


  or

  (
    g662_n,
    g598_p_spl_,
    n3172_o2_n
  );


  and

  (
    g663_p,
    g597_n_spl_0,
    n3245_o2_n_spl_
  );


  or

  (
    g664_n,
    g595_p_spl_,
    n3246_o2_p_spl_00
  );


  or

  (
    g665_n,
    lo086_buf_o2_p_spl_0,
    n1950_lo_p_spl_0
  );


  and

  (
    g666_p,
    g592_n_spl_,
    g572_p_spl_0
  );


  or

  (
    g667_n,
    g657_n_spl_,
    lo034_buf_o2_p_spl_00
  );


  and

  (
    g668_p,
    n762_o2_n_spl_,
    n763_o2_n
  );


  or

  (
    g668_n,
    n762_o2_p,
    n763_o2_p
  );


  and

  (
    g669_p,
    g668_n_spl_0,
    lo042_buf_o2_p_spl_00
  );


  or

  (
    g669_n,
    g668_p_spl_0,
    lo042_buf_o2_n_spl_0
  );


  and

  (
    g670_p,
    n760_o2_n_spl_0,
    lo042_buf_o2_n_spl_0
  );


  or

  (
    g670_n,
    n760_o2_p_spl_00,
    lo042_buf_o2_p_spl_00
  );


  and

  (
    g671_p,
    g670_n,
    g669_n
  );


  or

  (
    g671_n,
    g670_p,
    g669_p
  );


  and

  (
    g672_p,
    lo034_buf_o2_n_spl_0,
    n754_o2_n_spl_0
  );


  or

  (
    g672_n,
    lo034_buf_o2_p_spl_0,
    n754_o2_p_spl_0
  );


  and

  (
    g673_p,
    n820_o2_n,
    n822_o2_n
  );


  or

  (
    g673_n,
    n820_o2_p,
    n822_o2_p
  );


  and

  (
    g674_p,
    g673_p,
    g672_n
  );


  or

  (
    g674_n,
    g673_n,
    g672_p
  );


  and

  (
    g675_p,
    g674_n,
    n751_o2_p_spl_000
  );


  or

  (
    g675_n,
    g674_p,
    n751_o2_n_spl_00
  );


  and

  (
    g676_p,
    g675_n,
    g671_n
  );


  or

  (
    g676_n,
    g675_p,
    g671_p
  );


  and

  (
    g677_p,
    g668_n_spl_0,
    lo046_buf_o2_p_spl_0
  );


  or

  (
    g677_n,
    g668_p_spl_0,
    lo046_buf_o2_n_spl_0
  );


  and

  (
    g678_p,
    n760_o2_n_spl_0,
    lo046_buf_o2_n_spl_0
  );


  or

  (
    g678_n,
    n760_o2_p_spl_00,
    lo046_buf_o2_p_spl_0
  );


  and

  (
    g679_p,
    g678_n,
    g677_n
  );


  or

  (
    g679_n,
    g678_p,
    g677_p
  );


  and

  (
    g680_p,
    lo038_buf_o2_p_spl_00,
    n755_o2_n_spl_0
  );


  or

  (
    g680_n,
    lo038_buf_o2_n_spl_,
    n755_o2_p
  );


  and

  (
    g681_p,
    n846_o2_n,
    n849_o2_n
  );


  or

  (
    g681_n,
    n846_o2_p,
    n849_o2_p
  );


  and

  (
    g682_p,
    g681_p,
    g680_n
  );


  or

  (
    g682_n,
    g681_n,
    g680_p
  );


  and

  (
    g683_p,
    g682_n,
    n751_o2_p_spl_000
  );


  or

  (
    g683_n,
    g682_p,
    n751_o2_n_spl_00
  );


  and

  (
    g684_p,
    g683_n,
    g679_n
  );


  or

  (
    g684_n,
    g683_p,
    g679_p
  );


  or

  (
    g685_n,
    lo034_buf_o2_n_spl_0,
    lo028_buf_o2_n_spl_0
  );


  and

  (
    g686_p,
    g685_n,
    g646_n_spl_
  );


  or

  (
    g687_n,
    lo006_buf_o2_p_spl_,
    lo002_buf_o2_p_spl_0
  );


  and

  (
    g688_p,
    lo150_buf_o2_p,
    n771_o2_n_spl_00
  );


  or

  (
    g688_n,
    lo150_buf_o2_n,
    n771_o2_p_spl_00
  );


  and

  (
    g689_p,
    lo018_buf_o2_n,
    lo022_buf_o2_n
  );


  or

  (
    g689_n,
    lo018_buf_o2_p_spl_,
    lo022_buf_o2_p_spl_
  );


  and

  (
    g690_p,
    g689_n,
    lo002_buf_o2_n
  );


  or

  (
    g690_n,
    g689_p,
    lo002_buf_o2_p_spl_0
  );


  and

  (
    g691_p,
    g690_p_spl_0,
    g688_p_spl_0
  );


  or

  (
    g691_n,
    g690_n_spl_0,
    g688_n_spl_0
  );


  and

  (
    g692_p,
    n751_o2_p_spl_00,
    lo010_buf_o2_p_spl_00
  );


  or

  (
    g692_n,
    n751_o2_n_spl_0,
    lo010_buf_o2_n_spl_
  );


  and

  (
    g693_p,
    g692_n_spl_,
    n760_o2_n_spl_1
  );


  or

  (
    g693_n,
    g692_p_spl_0,
    n760_o2_p_spl_01
  );


  and

  (
    g694_p,
    g693_n_spl_,
    lo050_buf_o2_n_spl_0
  );


  or

  (
    g694_n,
    g693_p,
    lo050_buf_o2_p_spl_0
  );


  and

  (
    g695_p,
    n754_o2_n_spl_0,
    lo042_buf_o2_n_spl_1
  );


  or

  (
    g695_n,
    n754_o2_p_spl_0,
    lo042_buf_o2_p_spl_0
  );


  and

  (
    g696_p,
    n753_o2_p_spl_0,
    lo054_buf_o2_p_spl_0
  );


  or

  (
    g696_n,
    n753_o2_n_spl_,
    lo054_buf_o2_n_spl_0
  );


  and

  (
    g697_p,
    g696_n,
    g695_n
  );


  or

  (
    g697_n,
    g696_p,
    g695_p
  );


  and

  (
    g698_p,
    g697_n,
    n751_o2_p_spl_01
  );


  or

  (
    g698_n,
    g697_p,
    n751_o2_n_spl_1
  );


  and

  (
    g699_p,
    g668_p_spl_1,
    lo050_buf_o2_p_spl_0
  );


  or

  (
    g699_n,
    g668_n_spl_1,
    lo050_buf_o2_n_spl_0
  );


  and

  (
    g700_p,
    g699_n,
    g698_n
  );


  or

  (
    g700_n,
    g699_p,
    g698_p
  );


  and

  (
    g701_p,
    g700_p,
    g694_n
  );


  or

  (
    g701_n,
    g700_n,
    g694_p
  );


  and

  (
    g702_p,
    g688_p_spl_0,
    n773_o2_n
  );


  or

  (
    g702_n,
    g688_n_spl_0,
    n773_o2_p
  );


  and

  (
    g703_p,
    n833_o2_n,
    n828_o2_n
  );


  or

  (
    g703_n,
    n833_o2_p,
    n828_o2_p
  );


  and

  (
    g704_p,
    g703_n,
    n771_o2_n_spl_00
  );


  or

  (
    g704_n,
    g703_p,
    n771_o2_p_spl_00
  );


  and

  (
    g705_p,
    g704_n,
    g702_n
  );


  or

  (
    g705_n,
    g704_p,
    g702_p
  );


  or

  (
    g706_n,
    g705_n_spl_,
    g658_p_spl_0
  );


  or

  (
    g707_n,
    g706_n,
    g676_p
  );


  and

  (
    g708_p,
    g688_p_spl_,
    n774_o2_n_spl_0
  );


  or

  (
    g708_n,
    g688_n_spl_,
    n774_o2_p_spl_0
  );


  and

  (
    g709_p,
    n859_o2_n,
    n854_o2_n
  );


  or

  (
    g709_n,
    n859_o2_p,
    n854_o2_p
  );


  and

  (
    g710_p,
    g709_n,
    n771_o2_n_spl_01
  );


  or

  (
    g710_n,
    g709_p,
    n771_o2_p_spl_01
  );


  and

  (
    g711_p,
    g710_n,
    g708_n_spl_0
  );


  or

  (
    g711_n,
    g710_p,
    g708_p_spl_0
  );


  or

  (
    g712_n,
    g711_n_spl_,
    g658_p_spl_0
  );


  or

  (
    g713_n,
    g712_n,
    g684_p
  );


  or

  (
    g714_n,
    g609_n_spl_1,
    n1139_o2_n
  );


  or

  (
    g715_n,
    g609_n_spl_1,
    n1081_o2_n_spl_
  );


  and

  (
    g716_p,
    g661_n_spl_,
    n3087_o2_p_spl_0
  );


  or

  (
    g717_n,
    n1007_o2_p_spl_,
    n2619_o2_n_spl_00
  );


  or

  (
    g718_n,
    g717_n_spl_0,
    n998_o2_n_spl_
  );


  or

  (
    g719_n,
    g595_p_spl_,
    n3245_o2_p_spl_0
  );


  or

  (
    g720_n,
    g599_p_spl_,
    n3246_o2_p_spl_00
  );


  and

  (
    g721_p,
    g603_p_spl_,
    g601_p_spl_
  );


  and

  (
    g722_p,
    n998_o2_n_spl_,
    lo186_buf_o2_p_spl_0
  );


  or

  (
    g722_n,
    n998_o2_p_spl_,
    lo186_buf_o2_n_spl_0
  );


  and

  (
    g723_p,
    n994_o2_p_spl_,
    n1220_o2_p
  );


  or

  (
    g723_n,
    n994_o2_n_spl_0,
    n1220_o2_n
  );


  and

  (
    g724_p,
    g723_n,
    n1221_o2_p_spl_
  );


  or

  (
    g724_n,
    g723_p,
    n1221_o2_n_spl_
  );


  and

  (
    g725_p,
    g724_n_spl_,
    g722_n_spl_
  );


  or

  (
    g725_n,
    g724_p_spl_,
    g722_p_spl_0
  );


  and

  (
    g726_p,
    g724_p_spl_,
    g722_p_spl_0
  );


  or

  (
    g726_n,
    g724_n_spl_,
    g722_n_spl_
  );


  and

  (
    g727_p,
    g726_n,
    g725_n
  );


  or

  (
    g727_n,
    g726_p,
    g725_p
  );


  and

  (
    g728_p,
    n1214_o2_n_spl_,
    n3082_o2_n_spl_
  );


  or

  (
    g728_n,
    n1214_o2_p_spl_,
    n3082_o2_p_spl_
  );


  and

  (
    g729_p,
    n1214_o2_p_spl_,
    n3082_o2_p_spl_
  );


  or

  (
    g729_n,
    n1214_o2_n_spl_,
    n3082_o2_n_spl_
  );


  and

  (
    g730_p,
    g729_n,
    g728_n
  );


  or

  (
    g730_n,
    g729_p,
    g728_p
  );


  and

  (
    g731_p,
    n1221_o2_p_spl_,
    n1222_o2_n
  );


  or

  (
    g731_n,
    n1221_o2_n_spl_,
    n1222_o2_p
  );


  and

  (
    g732_p,
    g731_n_spl_,
    g553_n_spl_
  );


  or

  (
    g732_n,
    g731_p_spl_,
    g553_p_spl_0
  );


  and

  (
    g733_p,
    g732_p_spl_,
    g730_p_spl_0
  );


  or

  (
    g733_n,
    g732_n_spl_,
    g730_n_spl_00
  );


  and

  (
    g734_p,
    g732_n_spl_,
    g730_n_spl_00
  );


  or

  (
    g734_n,
    g732_p_spl_,
    g730_p_spl_0
  );


  and

  (
    g735_p,
    g734_n,
    g733_n
  );


  or

  (
    g735_n,
    g734_p,
    g733_p
  );


  or

  (
    g736_n,
    g735_p_spl_,
    g727_p_spl_
  );


  and

  (
    g737_p,
    g736_n,
    n1003_o2_p_spl_0
  );


  or

  (
    g738_n,
    g737_p,
    g556_p_spl_0
  );


  and

  (
    g739_p,
    g738_n,
    g561_p_spl_
  );


  and

  (
    g740_p,
    g727_n_spl_0,
    g561_n_spl_01
  );


  and

  (
    g741_p,
    g735_n_spl_,
    g561_n_spl_1
  );


  and

  (
    g742_p,
    n998_o2_p_spl_,
    lo186_buf_o2_n_spl_1
  );


  or

  (
    g743_n,
    g742_p,
    g722_p_spl_
  );


  and

  (
    g744_p,
    n3028_o2_n_spl_,
    n2619_o2_n_spl_01
  );


  or

  (
    g744_n,
    n3028_o2_p_spl_0,
    n2619_o2_p_spl_00
  );


  or

  (
    g745_n,
    g744_p,
    n2624_o2_n_spl_0
  );


  and

  (
    g746_p,
    g559_n_spl_,
    n2620_o2_n_spl_
  );


  and

  (
    g747_p,
    g551_n_spl_,
    n2620_o2_p_spl_
  );


  or

  (
    g748_n,
    g744_n,
    g552_n_spl_
  );


  or

  (
    g749_n,
    g748_n,
    g747_p
  );


  or

  (
    g750_n,
    g749_n,
    g746_p
  );


  and

  (
    g751_p,
    g750_n,
    g745_n
  );


  or

  (
    g752_n,
    g751_p,
    g612_n_spl_
  );


  or

  (
    g753_n,
    n1040_o2_p_spl_00,
    n2289_lo_n
  );


  or

  (
    g754_n,
    lo174_buf_o2_n,
    n1044_o2_n_spl_0
  );


  or

  (
    g755_n,
    lo170_buf_o2_n,
    n1034_o2_p_spl_0
  );


  and

  (
    g756_p,
    g755_n,
    g754_n
  );


  and

  (
    g757_p,
    g756_p,
    g753_n
  );


  or

  (
    g758_n,
    n1034_o2_p_spl_0,
    n2627_o2_n
  );


  or

  (
    g759_n,
    lo166_buf_o2_n,
    n1040_o2_p_spl_00
  );


  and

  (
    g760_p,
    g759_n,
    g758_n
  );


  or

  (
    g761_n,
    n1046_o2_p_spl_0,
    n2676_o2_n_spl_
  );


  and

  (
    g762_p,
    g761_n,
    n2619_o2_p_spl_00
  );


  or

  (
    g763_n,
    lo178_buf_o2_n,
    n1038_o2_p_spl_0
  );


  or

  (
    g764_n,
    n1031_o2_n_spl_0,
    n2645_o2_n_spl_
  );


  and

  (
    g765_p,
    g764_n,
    g763_n
  );


  and

  (
    g766_p,
    g765_p,
    g762_p
  );


  and

  (
    g767_p,
    g766_p,
    g760_p_spl_
  );


  and

  (
    g768_p,
    g767_p,
    g757_p
  );


  or

  (
    g769_n,
    n1044_o2_n_spl_0,
    n2794_o2_p_spl_0
  );


  and

  (
    g770_p,
    g769_n,
    n1035_o2_p
  );


  or

  (
    g771_n,
    n1031_o2_n_spl_0,
    n2622_o2_p_spl_
  );


  and

  (
    g772_p,
    g771_n_spl_,
    n1036_o2_p
  );


  and

  (
    g773_p,
    g772_p,
    g770_p
  );


  or

  (
    g774_n,
    n1041_o2_p,
    n1040_o2_p_spl_0
  );


  and

  (
    g775_p,
    g774_n,
    n2619_o2_n_spl_01
  );


  or

  (
    g776_n,
    n1038_o2_p_spl_0,
    n2793_o2_p_spl_0
  );


  and

  (
    g777_p,
    g776_n,
    n1047_o2_p
  );


  and

  (
    g778_p,
    g777_p,
    g775_p
  );


  and

  (
    g779_p,
    g778_p,
    g773_p
  );


  or

  (
    g780_n,
    g779_p,
    g612_p_spl_01
  );


  or

  (
    g781_n,
    g780_n,
    g768_p
  );


  and

  (
    g782_p,
    g781_n,
    g752_n
  );


  or

  (
    g783_n,
    g782_p,
    g562_n_spl_
  );


  or

  (
    g784_n,
    n1040_o2_p_spl_1,
    n2624_o2_p_spl_
  );


  or

  (
    g785_n,
    n1034_o2_p_spl_1,
    n2621_o2_p_spl_
  );


  or

  (
    g786_n,
    n1038_o2_p_spl_1,
    n2676_o2_n_spl_
  );


  and

  (
    g787_p,
    g786_n,
    g785_n
  );


  and

  (
    g788_p,
    g787_p,
    g784_n
  );


  and

  (
    g789_p,
    g771_n_spl_,
    n2619_o2_p_spl_01
  );


  or

  (
    g790_n,
    n1046_o2_p_spl_0,
    n2623_o2_p_spl_
  );


  or

  (
    g791_n,
    n1044_o2_n_spl_1,
    n2645_o2_n_spl_
  );


  and

  (
    g792_p,
    g791_n,
    g790_n
  );


  and

  (
    g793_p,
    g792_p,
    g789_p
  );


  and

  (
    g794_p,
    g793_p,
    g760_p_spl_
  );


  and

  (
    g795_p,
    g794_p,
    g788_p
  );


  or

  (
    g796_n,
    n1031_o2_n_spl_,
    n2794_o2_p_spl_0
  );


  or

  (
    g797_n,
    n1038_o2_p_spl_1,
    lo074_buf_o2_n
  );


  or

  (
    g798_n,
    n1044_o2_n_spl_1,
    lo078_buf_o2_n
  );


  and

  (
    g799_p,
    g798_n,
    g797_n
  );


  and

  (
    g800_p,
    g799_p,
    g796_n
  );


  or

  (
    g801_n,
    n1099_o2_n,
    n1040_o2_p_spl_1
  );


  and

  (
    g802_p,
    g801_n,
    n2619_o2_n_spl_10
  );


  or

  (
    g803_n,
    n1046_o2_p_spl_,
    n2793_o2_p_spl_1
  );


  or

  (
    g804_n,
    n1102_o2_p,
    n1034_o2_p_spl_1
  );


  and

  (
    g805_p,
    g804_n,
    g803_n
  );


  and

  (
    g806_p,
    g805_p,
    g802_p
  );


  and

  (
    g807_p,
    g806_p,
    g800_p
  );


  or

  (
    g808_n,
    g807_p,
    g795_p
  );


  and

  (
    g809_p,
    g808_n,
    g612_n_spl_
  );


  or

  (
    g810_n,
    g809_p,
    g562_n_spl_
  );


  and

  (
    g811_p,
    n1031_o2_p_spl_00,
    n2623_o2_n_spl_
  );


  and

  (
    g812_p,
    lo166_buf_o2_p,
    n1038_o2_n_spl_00
  );


  or

  (
    g813_n,
    lo170_buf_o2_p_spl_,
    n2627_o2_p_spl_0
  );


  and

  (
    g814_p,
    g813_n,
    n1040_o2_n_spl_000
  );


  or

  (
    g815_n,
    g814_p,
    g812_p
  );


  or

  (
    g816_n,
    g815_n,
    g811_p
  );


  or

  (
    g817_n,
    n2645_o2_p_spl_0,
    n2622_o2_n_spl_
  );


  and

  (
    g818_p,
    g817_n,
    n1034_o2_n_spl_00
  );


  or

  (
    g819_n,
    g818_p,
    n2619_o2_n_spl_10
  );


  and

  (
    g820_p,
    n1046_o2_n_spl_00,
    n2624_o2_n_spl_0
  );


  and

  (
    g821_p,
    n1044_o2_p_spl_00,
    n2676_o2_p_spl_
  );


  or

  (
    g822_n,
    g821_p,
    g820_p
  );


  or

  (
    g823_n,
    g822_n,
    g819_n
  );


  or

  (
    g824_n,
    g823_n,
    g816_n
  );


  and

  (
    g825_p,
    n1044_o2_p_spl_00,
    n2966_o2_p_spl_0
  );


  and

  (
    g826_p,
    n1038_o2_n_spl_00,
    lo078_buf_o2_p
  );


  and

  (
    g827_p,
    n1041_o2_n,
    n1034_o2_n_spl_00
  );


  or

  (
    g828_n,
    g827_p,
    g826_p
  );


  or

  (
    g829_n,
    g828_n,
    g825_p
  );


  and

  (
    g830_p,
    n1040_o2_n_spl_000,
    n1202_o2_n
  );


  or

  (
    g831_n,
    g830_p,
    n2619_o2_p_spl_01
  );


  and

  (
    g832_p,
    n1046_o2_n_spl_00,
    n2794_o2_n
  );


  or

  (
    g833_n,
    g832_p,
    n1206_o2_p
  );


  or

  (
    g834_n,
    g833_n,
    g831_n
  );


  or

  (
    g835_n,
    g834_n,
    g829_n
  );


  and

  (
    g836_p,
    g835_n,
    g824_n
  );


  or

  (
    g837_n,
    g836_p,
    g612_p_spl_01
  );


  and

  (
    g838_p,
    g837_n,
    g562_p_spl_01
  );


  and

  (
    g839_p,
    n1040_o2_n_spl_00,
    n2623_o2_n_spl_
  );


  and

  (
    g840_p,
    n1044_o2_p_spl_01,
    n2627_o2_p_spl_0
  );


  or

  (
    g841_n,
    g840_p,
    g839_p
  );


  and

  (
    g842_p,
    n1038_o2_n_spl_01,
    n2645_o2_p_spl_0
  );


  or

  (
    g843_n,
    n2730_o2_n,
    n2624_o2_n_spl_1
  );


  and

  (
    g844_p,
    g843_n,
    n1034_o2_n_spl_01
  );


  or

  (
    g845_n,
    g844_p,
    g842_p
  );


  or

  (
    g846_n,
    g845_n,
    g841_n
  );


  and

  (
    g847_p,
    n1040_o2_n_spl_01,
    n2676_o2_p_spl_
  );


  or

  (
    g848_n,
    g847_p,
    n2619_o2_n_spl_1
  );


  and

  (
    g849_p,
    n1031_o2_p_spl_00,
    n2621_o2_n_spl_
  );


  and

  (
    g850_p,
    n1046_o2_n_spl_01,
    n2622_o2_n_spl_
  );


  or

  (
    g851_n,
    g850_p,
    g849_p_spl_
  );


  or

  (
    g852_n,
    g851_n,
    g848_n_spl_
  );


  or

  (
    g853_n,
    g852_n,
    g846_n
  );


  or

  (
    g854_n,
    lo066_buf_o2_p,
    n2966_o2_p_spl_0
  );


  and

  (
    g855_p,
    g854_n,
    n1040_o2_n_spl_01
  );


  and

  (
    g856_p,
    n1046_o2_n_spl_01,
    n2967_o2_p_spl_0
  );


  and

  (
    g857_p,
    n1298_o2_n_spl_,
    n1034_o2_n_spl_01
  );


  or

  (
    g858_n,
    g857_p,
    g856_p
  );


  or

  (
    g859_n,
    g858_n,
    g855_p
  );


  and

  (
    g860_p,
    n1031_o2_p_spl_0,
    n2793_o2_n_spl_
  );


  and

  (
    g861_p,
    n1044_o2_p_spl_01,
    lo074_buf_o2_p
  );


  or

  (
    g862_n,
    g861_p,
    g860_p
  );


  and

  (
    g863_p,
    lo070_buf_o2_p,
    n1038_o2_n_spl_01
  );


  or

  (
    g864_n,
    g863_p,
    n2619_o2_p_spl_10
  );


  or

  (
    g865_n,
    g864_n,
    g862_n
  );


  or

  (
    g866_n,
    g865_n,
    g859_n
  );


  and

  (
    g867_p,
    g866_n,
    g853_n
  );


  or

  (
    g868_n,
    g867_p,
    g612_p_spl_10
  );


  and

  (
    g869_p,
    g868_n,
    g562_p_spl_01
  );


  and

  (
    g870_p,
    n3214_o2_p_spl_,
    n2926_o2_p
  );


  or

  (
    g870_n,
    n3214_o2_n_spl_,
    n2926_o2_n
  );


  and

  (
    g871_p,
    g870_n_spl_,
    n3081_o2_n_spl_
  );


  or

  (
    g871_n,
    g870_p_spl_,
    n3081_o2_p_spl_
  );


  and

  (
    g872_p,
    g870_p_spl_,
    n3081_o2_p_spl_
  );


  or

  (
    g872_n,
    g870_n_spl_,
    n3081_o2_n_spl_
  );


  and

  (
    g873_p,
    g872_n,
    g871_n
  );


  or

  (
    g873_n,
    g872_p,
    g871_p
  );


  or

  (
    g874_n,
    g873_n_spl_0,
    g717_n_spl_0
  );


  or

  (
    g875_n,
    n1059_inv_p_spl_010,
    n791_o2_n_spl_
  );


  or

  (
    g876_n,
    g687_n_spl_,
    lo010_buf_o2_p_spl_00
  );


  and

  (
    g877_p,
    n923_o2_n,
    n929_o2_n
  );


  or

  (
    g877_n,
    n923_o2_p,
    n929_o2_p
  );


  and

  (
    g878_p,
    n938_o2_n,
    n884_o2_n
  );


  or

  (
    g878_n,
    n938_o2_p,
    n884_o2_p
  );


  or

  (
    g879_n,
    g878_n_spl_,
    n786_o2_n_spl_
  );


  and

  (
    g880_p,
    g879_n,
    g877_p_spl_0
  );


  and

  (
    g881_p,
    g877_n,
    n789_o2_p_spl_
  );


  or

  (
    g881_n,
    g877_p_spl_0,
    n789_o2_n_spl_
  );


  and

  (
    g882_p,
    g881_p,
    g878_p
  );


  or

  (
    g882_n,
    g881_n,
    g878_n_spl_
  );


  or

  (
    g883_n,
    g882_p,
    g880_p
  );


  or

  (
    g884_n,
    g883_n_spl_0,
    g652_n_spl_
  );


  or

  (
    g885_n,
    g884_n_spl_,
    g573_n_spl_
  );


  or

  (
    g886_n,
    g885_n_spl_,
    g568_n_spl_
  );


  or

  (
    g887_n,
    g727_n_spl_0,
    n1003_o2_n_spl_0
  );


  and

  (
    g888_p,
    g727_n_spl_,
    n1003_o2_n_spl_0
  );


  or

  (
    g888_n,
    g727_p_spl_,
    n1003_o2_p_spl_0
  );


  and

  (
    g889_p,
    g888_n_spl_,
    g887_n
  );


  or

  (
    g890_n,
    g656_n_spl_,
    g577_n_spl_0
  );


  or

  (
    g891_n,
    g717_n_spl_1,
    n994_o2_n_spl_
  );


  and

  (
    g892_p,
    lo174_buf_o2_p_spl_,
    n1038_o2_n_spl_10
  );


  and

  (
    g893_p,
    n1031_o2_p_spl_1,
    n2627_o2_p_spl_1
  );


  or

  (
    g894_n,
    g893_p,
    g892_p
  );


  and

  (
    g895_p,
    n1084_o2_n,
    n1034_o2_n_spl_1
  );


  and

  (
    g896_p,
    lo170_buf_o2_p_spl_,
    n1044_o2_p_spl_10
  );


  or

  (
    g897_n,
    g896_p,
    g895_p
  );


  or

  (
    g898_n,
    g897_n,
    g894_n
  );


  and

  (
    g899_p,
    n1046_o2_n_spl_10,
    n2645_o2_p_spl_
  );


  and

  (
    g900_p,
    lo178_buf_o2_p,
    n1040_o2_n_spl_10
  );


  or

  (
    g901_n,
    g900_p,
    g899_p
  );


  or

  (
    g902_n,
    g901_n,
    g848_n_spl_
  );


  or

  (
    g903_n,
    g902_n,
    g898_n
  );


  and

  (
    g904_p,
    n1038_o2_n_spl_10,
    n2967_o2_p_spl_0
  );


  and

  (
    g905_p,
    n1102_o2_n,
    n1040_o2_n_spl_10
  );


  or

  (
    g906_n,
    g905_p,
    g904_p
  );


  or

  (
    g907_n,
    g906_n,
    n1262_o2_n
  );


  and

  (
    g908_p,
    n1044_o2_p_spl_10,
    n2793_o2_n_spl_
  );


  or

  (
    g909_n,
    g908_p,
    g849_p_spl_
  );


  or

  (
    g910_n,
    n1271_o2_n,
    n2619_o2_p_spl_10
  );


  or

  (
    g911_n,
    g910_n,
    g909_n
  );


  or

  (
    g912_n,
    g911_n,
    g907_n
  );


  and

  (
    g913_p,
    g912_n,
    g903_n
  );


  or

  (
    g914_n,
    g913_p,
    g612_p_spl_10
  );


  and

  (
    g915_p,
    g914_n,
    g562_p_spl_10
  );


  and

  (
    g916_p,
    g915_p,
    g891_n
  );


  and

  (
    g917_p,
    g601_n_spl_,
    g561_n_spl_1
  );


  and

  (
    g918_p,
    g604_n_spl_,
    g556_n_spl_1
  );


  or

  (
    g919_n,
    g918_p,
    g917_p
  );


  or

  (
    g920_n,
    g730_n_spl_0,
    g717_n_spl_1
  );


  and

  (
    g921_p,
    n1046_o2_n_spl_10,
    n2729_o2_n
  );


  and

  (
    g922_p,
    n1038_o2_n_spl_1,
    n2966_o2_p_spl_
  );


  and

  (
    g923_p,
    n1044_o2_p_spl_1,
    n2967_o2_p_spl_
  );


  or

  (
    g924_n,
    g923_p,
    g922_p
  );


  or

  (
    g925_n,
    g924_n,
    g921_p
  );


  and

  (
    g926_p,
    n1298_o2_n_spl_,
    n1040_o2_n_spl_11
  );


  or

  (
    g927_n,
    g926_p,
    n2619_o2_p_spl_1
  );


  and

  (
    g928_p,
    n1294_o2_n,
    n1034_o2_n_spl_1
  );


  or

  (
    g929_n,
    g928_p,
    n1297_o2_p
  );


  or

  (
    g930_n,
    g929_n,
    g927_n
  );


  or

  (
    g931_n,
    g930_n,
    g925_n
  );


  and

  (
    g932_p,
    n1046_o2_n_spl_1,
    n2627_o2_p_spl_1
  );


  and

  (
    g933_p,
    lo174_buf_o2_p_spl_,
    n1040_o2_n_spl_11
  );


  and

  (
    g934_p,
    n1031_o2_p_spl_1,
    n2624_o2_n_spl_1
  );


  or

  (
    g935_n,
    g934_p,
    g933_p
  );


  or

  (
    g936_n,
    g935_n,
    g932_p
  );


  or

  (
    g937_n,
    n1306_o2_p,
    n1307_o2_p
  );


  or

  (
    g938_n,
    n1312_o2_p,
    n1311_o2_p
  );


  or

  (
    g939_n,
    g938_n,
    g937_n
  );


  or

  (
    g940_n,
    g939_n,
    n1310_o2_n
  );


  or

  (
    g941_n,
    g940_n,
    g936_n
  );


  and

  (
    g942_p,
    g941_n,
    g931_n
  );


  or

  (
    g943_n,
    g942_p,
    g612_p_spl_1
  );


  and

  (
    g944_p,
    g943_n,
    g562_p_spl_10
  );


  and

  (
    g945_p,
    g944_p,
    g920_n
  );


  and

  (
    g946_p,
    g888_n_spl_,
    g735_p_spl_
  );


  and

  (
    g947_p,
    g888_p,
    g735_n_spl_
  );


  or

  (
    g948_n,
    g947_p,
    g946_p
  );


  and

  (
    g949_p,
    lo030_buf_o2_p_spl_0,
    n3090_o2_p_spl_
  );


  or

  (
    g950_n,
    g949_p,
    g597_p_spl_0
  );


  and

  (
    g951_p,
    lo186_buf_o2_p_spl_1,
    n1125_o2_n
  );


  or

  (
    g951_n,
    lo186_buf_o2_n_spl_1,
    n1125_o2_p
  );


  and

  (
    g952_p,
    n1003_o2_p_spl_1,
    n1081_o2_n_spl_
  );


  or

  (
    g952_n,
    n1003_o2_n_spl_,
    n1081_o2_p
  );


  and

  (
    g953_p,
    g952_n,
    n1128_o2_n
  );


  or

  (
    g953_n,
    g952_p,
    n1128_o2_p
  );


  and

  (
    g954_p,
    g953_p,
    g951_p
  );


  and

  (
    g955_p,
    g953_n,
    g951_n
  );


  or

  (
    g956_n,
    g955_p,
    g954_p
  );


  and

  (
    g957_p,
    g730_n_spl_1,
    g553_p_spl_0
  );


  or

  (
    g957_n,
    g730_p_spl_1,
    g553_n_spl_
  );


  and

  (
    g958_p,
    n3214_o2_n_spl_,
    n2976_o2_p
  );


  or

  (
    g958_n,
    n3214_o2_p_spl_,
    n2976_o2_n
  );


  and

  (
    g959_p,
    g731_n_spl_,
    g730_n_spl_1
  );


  or

  (
    g959_n,
    g731_p_spl_,
    g730_p_spl_1
  );


  and

  (
    g960_p,
    g959_n,
    g958_n
  );


  or

  (
    g960_n,
    g959_p,
    g958_p
  );


  and

  (
    g961_p,
    g960_p_spl_,
    g873_n_spl_0
  );


  or

  (
    g961_n,
    g960_n_spl_,
    g873_p_spl_
  );


  and

  (
    g962_p,
    g960_n_spl_,
    g873_p_spl_
  );


  or

  (
    g962_n,
    g960_p_spl_,
    g873_n_spl_
  );


  and

  (
    g963_p,
    g962_n,
    g961_n
  );


  or

  (
    g963_n,
    g962_p,
    g961_p
  );


  and

  (
    g964_p,
    g963_n,
    g957_n
  );


  and

  (
    g965_p,
    g963_p,
    g957_p
  );


  or

  (
    g966_n,
    g965_p,
    g964_p
  );


  or

  (
    g967_n,
    g645_n_spl_0,
    g621_n_spl_0
  );


  and

  (
    g968_p,
    g645_n_spl_0,
    g621_n_spl_0
  );


  and

  (
    g969_p,
    n1059_inv_p_spl_011,
    n801_o2_p
  );


  or

  (
    g969_n,
    n1059_inv_n_spl_01,
    n801_o2_n
  );


  and

  (
    g970_p,
    g969_n,
    n815_o2_n
  );


  and

  (
    g971_p,
    g969_p,
    n815_o2_p
  );


  or

  (
    g972_n,
    g971_p,
    g970_p
  );


  and

  (
    g973_p,
    n1059_inv_p_spl_011,
    n769_o2_p
  );


  or

  (
    g973_n,
    n1059_inv_n_spl_10,
    n769_o2_n
  );


  and

  (
    g974_p,
    g973_n,
    n792_o2_n_spl_
  );


  and

  (
    g975_p,
    g973_p,
    n792_o2_p_spl_
  );


  or

  (
    g976_n,
    g975_p,
    g974_p
  );


  and

  (
    g977_p,
    n754_o2_n_spl_1,
    lo046_buf_o2_n_spl_1
  );


  or

  (
    g977_n,
    n754_o2_p_spl_,
    lo046_buf_o2_p_spl_1
  );


  and

  (
    g978_p,
    n753_o2_p_spl_0,
    lo154_buf_o2_p_spl_
  );


  or

  (
    g978_n,
    n753_o2_n_spl_,
    lo154_buf_o2_n
  );


  and

  (
    g979_p,
    g978_n,
    g977_n
  );


  or

  (
    g979_n,
    g978_p,
    g977_p
  );


  and

  (
    g980_p,
    g979_n,
    n751_o2_p_spl_01
  );


  or

  (
    g980_n,
    g979_p,
    n751_o2_n_spl_1
  );


  and

  (
    g981_p,
    n760_o2_n_spl_1,
    lo054_buf_o2_n_spl_0
  );


  or

  (
    g981_n,
    n760_o2_p_spl_01,
    lo054_buf_o2_p_spl_0
  );


  and

  (
    g982_p,
    g692_n_spl_,
    lo054_buf_o2_p_spl_1
  );


  or

  (
    g982_n,
    g692_p_spl_0,
    lo054_buf_o2_n_spl_
  );


  and

  (
    g983_p,
    g982_p,
    g668_n_spl_1
  );


  or

  (
    g983_n,
    g982_n,
    g668_p_spl_1
  );


  and

  (
    g984_p,
    g983_n,
    g981_n
  );


  or

  (
    g984_n,
    g983_p,
    g981_p
  );


  and

  (
    g985_p,
    g984_n,
    g980_n
  );


  or

  (
    g985_n,
    g984_p,
    g980_p
  );


  and

  (
    g986_p,
    lo142_buf_o2_p_spl_,
    n774_o2_p_spl_0
  );


  or

  (
    g986_n,
    lo142_buf_o2_n,
    n774_o2_n_spl_0
  );


  and

  (
    g987_p,
    n805_o2_n,
    n806_o2_n
  );


  or

  (
    g987_n,
    n805_o2_p,
    n806_o2_p
  );


  and

  (
    g988_p,
    g987_p,
    g986_n
  );


  or

  (
    g988_n,
    g987_n,
    g986_p
  );


  and

  (
    g989_p,
    g988_n,
    n771_o2_n_spl_01
  );


  or

  (
    g989_n,
    g988_p,
    n771_o2_p_spl_01
  );


  and

  (
    g990_p,
    g989_n,
    g708_n_spl_0
  );


  or

  (
    g990_n,
    g989_p,
    g708_p_spl_0
  );


  or

  (
    g991_n,
    g990_n_spl_,
    g658_p_spl_1
  );


  or

  (
    g992_n,
    g991_n,
    g701_p
  );


  and

  (
    g993_p,
    g705_p_spl_,
    g659_n_spl_00
  );


  or

  (
    g994_n,
    g993_p,
    g676_n_spl_
  );


  and

  (
    g995_p,
    g994_n,
    g707_n_spl_
  );


  and

  (
    g996_p,
    g711_p_spl_,
    g659_n_spl_00
  );


  or

  (
    g997_n,
    g996_p,
    g684_n_spl_
  );


  and

  (
    g998_p,
    g997_n,
    g713_n_spl_
  );


  or

  (
    g999_n,
    n3086_o2_p_spl_,
    n2993_o2_p_spl_1
  );


  and

  (
    g1000_p,
    lo026_buf_o2_p_spl_,
    n3089_o2_p_spl_
  );


  and

  (
    g1001_p,
    n3092_o2_p_spl_,
    n2238_lo_n
  );


  and

  (
    g1002_p,
    g581_n_spl_00,
    n3092_o2_n_spl_
  );


  and

  (
    g1003_p,
    g597_n_spl_0,
    n3213_o2_p_spl_
  );


  and

  (
    g1004_p,
    g583_n_spl_00,
    n1938_lo_p_spl_0
  );


  or

  (
    g1005_n,
    g1004_p,
    n3193_o2_n
  );


  and

  (
    g1006_p,
    lo082_buf_o2_n,
    n3245_o2_p_spl_0
  );


  and

  (
    g1007_p,
    lo086_buf_o2_n,
    n3246_o2_p_spl_0
  );


  and

  (
    g1008_p,
    lo030_buf_o2_p_spl_0,
    n1974_lo_n
  );


  or

  (
    g1009_n,
    lo030_buf_o2_n,
    lo026_buf_o2_n_spl_
  );


  and

  (
    g1010_p,
    g1009_n,
    n673_o2_p
  );


  and

  (
    g1011_p,
    n1059_inv_p_spl_10,
    n853_o2_p
  );


  and

  (
    g1012_p,
    n1059_inv_n_spl_10,
    n814_o2_p_spl_
  );


  and

  (
    g1013_p,
    n1059_inv_n_spl_11,
    n897_o2_p_spl_
  );


  or

  (
    g1013_n,
    n1059_inv_p_spl_10,
    n897_o2_n_spl_0
  );


  or

  (
    g1014_n,
    g1013_p_spl_0,
    g890_n_spl_
  );


  and

  (
    g1015_p,
    g886_n_spl_0,
    g567_p_spl_0
  );


  and

  (
    g1016_p,
    g581_n_spl_00,
    n1926_lo_p_spl_
  );


  or

  (
    g1017_n,
    g976_n_spl_,
    n2298_lo_n_spl_
  );


  and

  (
    g1018_p,
    g581_n_spl_01,
    n2250_lo_p_spl_
  );


  and

  (
    g1019_p,
    g583_n_spl_00,
    n2238_lo_p_spl_
  );


  or

  (
    g1020_n,
    g877_p_spl_,
    n989_o2_n_spl_0
  );


  and

  (
    g1021_p,
    g1020_n_spl_,
    g883_n_spl_0
  );


  or

  (
    g1022_n,
    g1020_n_spl_,
    g883_n_spl_1
  );


  and

  (
    g1023_p,
    g886_n_spl_0,
    g592_n_spl_
  );


  and

  (
    g1024_p,
    g590_p_spl_,
    n2298_lo_p_spl_
  );


  or

  (
    g1024_n,
    g590_n,
    n2298_lo_n_spl_
  );


  or

  (
    g1025_n,
    g1024_n,
    g577_n_spl_0
  );


  and

  (
    g1026_p,
    n1059_inv_n_spl_11,
    n919_o2_p_spl_
  );


  or

  (
    g1026_n,
    n1059_inv_p_spl_11,
    n919_o2_n_spl_0
  );


  and

  (
    g1027_p,
    g1013_n,
    g577_p_spl_0
  );


  or

  (
    g1027_n,
    g1013_p_spl_0,
    g577_n_spl_
  );


  and

  (
    g1028_p,
    g1027_n,
    g1026_n
  );


  or

  (
    g1028_n,
    g1027_p,
    g1026_p_spl_
  );


  and

  (
    g1029_p,
    g1028_p,
    g656_p_spl_0
  );


  and

  (
    g1030_p,
    g1028_n,
    g656_n_spl_
  );


  or

  (
    g1031_n,
    g1030_p,
    g1029_p
  );


  or

  (
    g1032_n,
    g1031_n_spl_,
    g1025_n_spl_0
  );


  and

  (
    g1033_p,
    g1031_n_spl_,
    g1025_n_spl_0
  );


  or

  (
    g1034_n,
    G2_n_spl_,
    G1_p_spl_0
  );


  or

  (
    g1035_n,
    G6_p_spl_,
    G1_p_spl_0
  );


  and

  (
    g1036_p,
    g664_n_spl_,
    g662_n_spl_
  );


  and

  (
    g1037_p,
    g1036_p,
    g716_p_spl_
  );


  and

  (
    g1038_p,
    g599_n_spl_0,
    lo082_buf_o2_p_spl_0
  );


  and

  (
    g1039_p,
    g597_n_spl_1,
    g591_n_spl_
  );


  or

  (
    g1040_n,
    g1039_p,
    g1038_p
  );


  or

  (
    g1041_n,
    n1974_lo_p_spl_0,
    n1926_lo_p_spl_
  );


  and

  (
    g1042_p,
    g1041_n,
    g598_n_spl_0
  );


  or

  (
    g1043_n,
    g1042_p,
    n3087_o2_p_spl_0
  );


  or

  (
    g1044_n,
    g1043_n,
    g1040_n
  );


  and

  (
    g1045_p,
    n3170_o2_p_spl_,
    n3087_o2_n
  );


  and

  (
    g1046_p,
    g1045_p,
    g719_n_spl_
  );


  and

  (
    g1047_p,
    g583_n_spl_01,
    n3091_o2_n
  );


  or

  (
    g1048_n,
    n3095_o2_p_spl_0,
    n3089_o2_n_spl_
  );


  and

  (
    g1049_p,
    g1048_n,
    g598_n_spl_0
  );


  or

  (
    g1050_n,
    g1049_p,
    g1047_p
  );


  or

  (
    g1051_n,
    n3246_o2_p_spl_1,
    n3245_o2_p_spl_1
  );


  or

  (
    g1052_n,
    n3246_o2_n,
    n3245_o2_n_spl_
  );


  and

  (
    g1053_p,
    g1052_n,
    g1051_n
  );


  and

  (
    g1054_p,
    g950_n_spl_,
    g720_n_spl_
  );


  or

  (
    g1055_n,
    n1962_lo_p_spl_0,
    n1914_lo_p
  );


  and

  (
    g1056_p,
    g1055_n,
    g598_n_spl_1
  );


  and

  (
    g1057_p,
    g595_n_spl_0,
    lo082_buf_o2_p_spl_0
  );


  or

  (
    g1058_n,
    g1057_p,
    g1056_p
  );


  and

  (
    g1059_p,
    g595_n_spl_0,
    lo086_buf_o2_p_spl_0
  );


  and

  (
    g1060_p,
    g581_n_spl_01,
    n1938_lo_p_spl_0
  );


  and

  (
    g1061_p,
    g583_n_spl_01,
    n1950_lo_p_spl_0
  );


  or

  (
    g1062_n,
    g1061_p,
    g1060_p
  );


  or

  (
    g1063_n,
    g1062_n,
    g1059_p
  );


  and

  (
    g1064_p,
    g1026_p_spl_,
    g656_p_spl_0
  );


  and

  (
    g1065_p,
    g651_p_spl_,
    n989_o2_n_spl_
  );


  or

  (
    g1066_n,
    g1065_p,
    g1064_p
  );


  and

  (
    g1067_p,
    g972_n_spl_,
    g875_n_spl_
  );


  or

  (
    g1068_n,
    g885_n_spl_,
    n897_o2_n_spl_
  );


  or

  (
    g1069_n,
    g884_n_spl_,
    n919_o2_n_spl_
  );


  or

  (
    g1070_n,
    g883_n_spl_1,
    g651_n_spl_
  );


  and

  (
    g1071_p,
    g1070_n,
    g882_n
  );


  and

  (
    g1072_p,
    g1071_p,
    g1069_n
  );


  and

  (
    g1073_p,
    g1072_p,
    g1068_n
  );


  or

  (
    g1074_n,
    g876_n_spl_,
    n2055_lo_n
  );


  and

  (
    g1075_p,
    n754_o2_n_spl_1,
    lo028_buf_o2_n_spl_0
  );


  and

  (
    g1076_p,
    n752_o2_p_spl_0,
    lo042_buf_o2_n_spl_1
  );


  or

  (
    g1077_n,
    g1076_p,
    g1075_p
  );


  and

  (
    g1078_p,
    g1077_n,
    n751_o2_p_spl_10
  );


  or

  (
    g1079_n,
    lo038_buf_o2_p_spl_00,
    n760_o2_p_spl_10
  );


  or

  (
    g1080_n,
    g692_p_spl_,
    lo038_buf_o2_n_spl_
  );


  or

  (
    g1081_n,
    lo010_buf_o2_n_spl_,
    lo002_buf_o2_p_spl_1
  );


  and

  (
    g1082_p,
    g1081_n,
    n762_o2_n_spl_
  );


  or

  (
    g1083_n,
    g1082_p_spl_0,
    g1080_n
  );


  and

  (
    g1084_p,
    g1083_n,
    g1079_n
  );


  or

  (
    g1085_n,
    g1084_p,
    g1078_p
  );


  or

  (
    g1086_n,
    g1013_p_spl_,
    g666_p_spl_
  );


  or

  (
    g1087_n,
    g1024_p,
    g577_p_spl_0
  );


  and

  (
    g1088_p,
    g1087_n,
    g1025_n_spl_
  );


  or

  (
    g1089_n,
    g1088_p_spl_,
    g1086_n_spl_
  );


  and

  (
    g1090_p,
    g1088_p_spl_,
    g1086_n_spl_
  );


  and

  (
    g1091_p,
    g693_n_spl_,
    lo034_buf_o2_n_spl_1
  );


  and

  (
    g1092_p,
    n755_o2_n_spl_0,
    lo024_buf_o2_p_spl_0
  );


  and

  (
    g1093_p,
    lo038_buf_o2_p_spl_0,
    n753_o2_p_spl_
  );


  or

  (
    g1094_n,
    g1093_p,
    g1092_p
  );


  and

  (
    g1095_p,
    g1094_n,
    n751_o2_p_spl_10
  );


  and

  (
    g1096_p,
    g1082_p_spl_0,
    lo034_buf_o2_p_spl_1
  );


  or

  (
    g1097_n,
    g1096_p,
    g1095_p
  );


  or

  (
    g1098_n,
    g1097_n,
    g1091_p
  );


  and

  (
    g1099_p,
    g599_n_spl_,
    n1974_lo_p_spl_0
  );


  and

  (
    g1100_p,
    g665_n_spl_,
    g597_n_spl_1
  );


  or

  (
    g1101_n,
    g1100_p,
    g1099_p
  );


  and

  (
    g1102_p,
    lo145_buf_o2_p_spl_,
    n774_o2_p_spl_
  );


  or

  (
    g1102_n,
    lo145_buf_o2_n,
    n774_o2_n_spl_
  );


  and

  (
    g1103_p,
    n778_o2_n,
    n777_o2_p
  );


  or

  (
    g1103_n,
    n778_o2_p,
    n777_o2_n
  );


  and

  (
    g1104_p,
    n780_o2_n_spl_0,
    lo138_buf_o2_p_spl_
  );


  or

  (
    g1104_n,
    n780_o2_p_spl_0,
    lo138_buf_o2_n
  );


  and

  (
    g1105_p,
    g1104_n,
    g1103_n
  );


  or

  (
    g1105_n,
    g1104_p,
    g1103_p
  );


  and

  (
    g1106_p,
    g1105_p,
    g1102_n
  );


  or

  (
    g1106_n,
    g1105_n,
    g1102_p
  );


  and

  (
    g1107_p,
    g1106_n,
    n771_o2_n_spl_10
  );


  or

  (
    g1107_n,
    g1106_p,
    n771_o2_p_spl_10
  );


  and

  (
    g1108_p,
    g1107_n,
    g708_n_spl_
  );


  or

  (
    g1108_n,
    g1107_p,
    g708_p_spl_
  );


  or

  (
    g1109_n,
    g1108_n_spl_,
    g658_p_spl_1
  );


  or

  (
    g1110_n,
    g1109_n,
    g985_p
  );


  and

  (
    g1111_p,
    g598_n_spl_1,
    n3090_o2_n
  );


  or

  (
    g1112_n,
    g1111_p,
    g663_p_spl_
  );


  and

  (
    g1113_p,
    g581_n_spl_1,
    n3095_o2_p_spl_0
  );


  and

  (
    g1114_p,
    g583_n_spl_1,
    n3092_o2_n_spl_
  );


  or

  (
    g1115_n,
    g1114_p,
    g1113_p
  );


  or

  (
    g1116_n,
    g1115_n,
    g660_p_spl_
  );


  or

  (
    g1117_n,
    g1116_n,
    g1112_n
  );


  and

  (
    g1118_p,
    g990_p_spl_,
    g659_n_spl_01
  );


  or

  (
    g1119_n,
    g1118_p,
    g701_n_spl_
  );


  and

  (
    g1120_p,
    g1119_n,
    g992_n_spl_
  );


  and

  (
    g1121_p,
    g998_p_spl_,
    g995_p_spl_
  );


  or

  (
    g1122_n,
    G49_p,
    G4_p_spl_000
  );


  or

  (
    g1123_n,
    G12_p_spl_0,
    G11_p_spl_
  );


  or

  (
    g1124_n,
    G13_p_spl_0,
    G12_p_spl_0
  );


  and

  (
    g1125_p,
    n755_o2_n_spl_1,
    n1983_lo_p_spl_
  );


  and

  (
    g1126_p,
    lo028_buf_o2_n_spl_1,
    n752_o2_p_spl_0
  );


  and

  (
    g1127_p,
    g667_n_spl_,
    lo010_buf_o2_p_spl_0
  );


  or

  (
    g1128_n,
    g1127_p,
    g1126_p
  );


  or

  (
    g1129_n,
    g1128_n,
    g1125_p
  );


  and

  (
    g1130_p,
    g1129_n,
    n751_o2_p_spl_11
  );


  and

  (
    g1131_p,
    n755_o2_n_spl_1,
    n1995_lo_p_spl_
  );


  and

  (
    g1132_p,
    lo034_buf_o2_n_spl_1,
    n752_o2_p_spl_
  );


  and

  (
    g1133_p,
    g686_p_spl_,
    lo010_buf_o2_p_spl_1
  );


  or

  (
    g1134_n,
    g1133_p,
    g1132_p
  );


  or

  (
    g1135_n,
    g1134_n,
    g1131_p
  );


  and

  (
    g1136_p,
    g1135_n,
    n751_o2_p_spl_11
  );


  and

  (
    g1137_p,
    g690_n_spl_0,
    lo117_buf_o2_p_spl_0
  );


  or

  (
    g1138_n,
    lo038_buf_o2_p_spl_1,
    lo014_buf_o2_p_spl_00
  );


  or

  (
    g1139_n,
    lo014_buf_o2_n_spl_0,
    n2079_lo_p_spl_
  );


  and

  (
    g1140_p,
    g1139_n,
    g1138_n
  );


  and

  (
    g1141_p,
    n780_o2_n_spl_0,
    n2067_lo_p
  );


  or

  (
    g1142_n,
    g1141_p,
    g1140_p
  );


  or

  (
    g1143_n,
    g1142_n,
    g1137_p
  );


  and

  (
    g1144_p,
    g1143_n,
    n771_o2_n_spl_10
  );


  or

  (
    g1145_n,
    g1108_p_spl_,
    g990_p_spl_
  );


  or

  (
    g1146_n,
    g711_p_spl_,
    g705_p_spl_
  );


  or

  (
    g1147_n,
    g1146_n,
    g1145_n
  );


  and

  (
    g1148_p,
    g1147_n,
    lo092_buf_o2_p_spl_0
  );


  or

  (
    g1149_n,
    g1108_n_spl_,
    g990_n_spl_
  );


  or

  (
    g1150_n,
    g711_n_spl_,
    g705_n_spl_
  );


  or

  (
    g1151_n,
    g1150_n,
    g1149_n
  );


  and

  (
    g1152_p,
    g1151_n,
    lo092_buf_o2_n_spl_
  );


  and

  (
    g1153_p,
    g690_n_spl_,
    lo122_buf_o2_p_spl_
  );


  or

  (
    g1154_n,
    lo042_buf_o2_p_spl_1,
    lo014_buf_o2_p_spl_00
  );


  or

  (
    g1155_n,
    lo117_buf_o2_p_spl_0,
    lo014_buf_o2_n_spl_0
  );


  and

  (
    g1156_p,
    g1155_n,
    g1154_n
  );


  and

  (
    g1157_p,
    n780_o2_n_spl_,
    n2079_lo_p_spl_
  );


  or

  (
    g1158_n,
    g1157_p,
    g1156_p
  );


  or

  (
    g1159_n,
    g1158_n,
    g1153_p
  );


  and

  (
    g1160_p,
    g1159_n,
    n771_o2_n_spl_1
  );


  or

  (
    g1161_n,
    g1160_p,
    g691_p_spl_
  );


  or

  (
    g1162_n,
    G4_n_spl_00,
    G3_p_spl_00
  );


  or

  (
    g1163_n,
    g1034_n_spl_,
    G3_n_spl_
  );


  and

  (
    g1164_p,
    G5_p_spl_0,
    G4_p_spl_000
  );


  or

  (
    g1165_n,
    g1082_p_spl_1,
    lo024_buf_o2_n
  );


  or

  (
    g1166_n,
    lo024_buf_o2_p_spl_1,
    n760_o2_p_spl_10
  );


  and

  (
    g1167_p,
    g1166_n,
    g1165_n
  );


  or

  (
    g1168_n,
    g1082_p_spl_1,
    lo028_buf_o2_n_spl_1
  );


  or

  (
    g1169_n,
    lo028_buf_o2_p_spl_1,
    n760_o2_p_spl_1
  );


  and

  (
    g1170_p,
    g1169_n,
    g1168_n
  );


  or

  (
    g1171_n,
    g690_p_spl_0,
    lo130_buf_o2_n
  );


  and

  (
    g1172_p,
    lo050_buf_o2_n_spl_,
    lo014_buf_o2_n_spl_1
  );


  and

  (
    g1173_p,
    lo126_buf_o2_n_spl_,
    lo014_buf_o2_p_spl_0
  );


  or

  (
    g1174_n,
    g1173_p,
    g1172_p
  );


  or

  (
    g1175_n,
    lo122_buf_o2_n_spl_,
    n780_o2_p_spl_0
  );


  and

  (
    g1176_p,
    g1175_n,
    g1174_n
  );


  and

  (
    g1177_p,
    g1176_p,
    g1171_n
  );


  or

  (
    g1178_n,
    g1177_p,
    n771_o2_p_spl_10
  );


  and

  (
    g1179_p,
    g1178_n,
    g691_n_spl_
  );


  and

  (
    g1180_p,
    g1179_p_spl_,
    g658_n_spl_0
  );


  and

  (
    g1181_p,
    g1180_p,
    g1085_n_spl_0
  );


  or

  (
    g1182_n,
    g690_p_spl_,
    lo126_buf_o2_n_spl_
  );


  and

  (
    g1183_p,
    lo046_buf_o2_n_spl_1,
    lo014_buf_o2_n_spl_1
  );


  and

  (
    g1184_p,
    lo122_buf_o2_n_spl_,
    lo014_buf_o2_p_spl_1
  );


  or

  (
    g1185_n,
    g1184_p,
    g1183_p
  );


  or

  (
    g1186_n,
    lo117_buf_o2_n,
    n780_o2_p_spl_
  );


  and

  (
    g1187_p,
    g1186_n,
    g1185_n
  );


  and

  (
    g1188_p,
    g1187_p,
    g1182_n
  );


  or

  (
    g1189_n,
    g1188_p,
    n771_o2_p_spl_1
  );


  and

  (
    g1190_p,
    g1189_n,
    g691_n_spl_
  );


  and

  (
    g1191_p,
    g1190_p_spl_,
    g658_n_spl_0
  );


  and

  (
    g1192_p,
    g1191_p,
    g1098_n_spl_0
  );


  and

  (
    g1193_p,
    g1179_p_spl_,
    g659_n_spl_01
  );


  or

  (
    g1194_n,
    g1193_p,
    g1085_n_spl_0
  );


  and

  (
    g1195_p,
    g1190_p_spl_,
    g659_n_spl_10
  );


  or

  (
    g1196_n,
    g1195_p,
    g1098_n_spl_0
  );


  or

  (
    g1197_n,
    G2_n_spl_,
    G1_n_spl_0
  );


  or

  (
    g1198_n,
    G3_n_spl_,
    G1_n_spl_0
  );


  or

  (
    g1199_n,
    g1198_n,
    G4_n_spl_00
  );


  and

  (
    g1200_p,
    g1199_n,
    g1197_n_spl_
  );


  or

  (
    g1201_n,
    g1035_n_spl_0,
    G5_p_spl_0
  );


  or

  (
    g1202_n,
    g1074_n_spl_,
    n2307_lo_n
  );


  and

  (
    g1203_p,
    g1108_p_spl_,
    g659_n_spl_10
  );


  or

  (
    g1204_n,
    g1203_p,
    g985_n_spl_
  );


  and

  (
    g1205_p,
    g1204_n,
    g1110_n_spl_
  );


  and

  (
    g1206_p,
    g1121_p_spl_,
    g1120_p_spl_
  );


  or

  (
    g1207_n,
    G13_n_spl_,
    G12_n
  );


  and

  (
    g1208_p,
    g1207_n,
    g1124_n_spl_
  );


  and

  (
    g1209_p,
    G4_p_spl_001,
    G1_n_spl_
  );


  or

  (
    g1210_n,
    G4_p_spl_001,
    G3_p_spl_00
  );


  or

  (
    g1211_n,
    g1123_n_spl_,
    G13_p_spl_0
  );


  and

  (
    g1212_p,
    g1211_n,
    G3_p_spl_0
  );


  and

  (
    g1213_p,
    g1208_p_spl_,
    G3_p_spl_1
  );


  or

  (
    g1214_n,
    G41_p_spl_,
    G4_p_spl_01
  );


  and

  (
    g1215_p,
    G36_n,
    G4_p_spl_01
  );


  or

  (
    g1216_n,
    g1162_n_spl_0,
    G12_p_spl_1
  );


  or

  (
    g1217_n,
    g1162_n_spl_0,
    G13_n_spl_
  );


  or

  (
    g1218_n,
    g1122_n_spl_0,
    G34_n_spl_
  );


  or

  (
    g1219_n,
    g1197_n_spl_,
    g1164_p_spl_
  );


  and

  (
    g1220_p,
    g1201_n_spl_,
    G35_p_spl_0
  );


  or

  (
    g1221_n,
    g1122_n_spl_0,
    G32_n
  );


  and

  (
    g1222_p,
    g1200_p_spl_,
    g1163_n_spl_
  );


  or

  (
    g1223_n,
    G40_p_spl_,
    G4_p_spl_10
  );


  or

  (
    g1224_n,
    G35_p_spl_0,
    G4_n_spl_0
  );


  and

  (
    g1225_p,
    g1224_n,
    g1223_n
  );


  and

  (
    g1226_p,
    G39_n,
    G4_n_spl_1
  );


  and

  (
    g1227_p,
    G34_n_spl_,
    G4_p_spl_10
  );


  or

  (
    g1228_n,
    g1227_p,
    g1226_p
  );


  or

  (
    g1229_n,
    g1122_n_spl_1,
    G33_n
  );


  and

  (
    g1230_p,
    g1229_n,
    g1228_n
  );


  and

  (
    g1231_p,
    G33_p_spl_,
    G4_p_spl_11
  );


  and

  (
    g1232_p,
    G14_p_spl_,
    G4_n_spl_1
  );


  or

  (
    g1233_n,
    g1232_p,
    g1231_p
  );


  and

  (
    g1234_p,
    g1035_n_spl_0,
    G34_p_spl_
  );


  or

  (
    g1235_n,
    g1234_p,
    g1233_n
  );


  buf

  (
    G3519,
    g412_p
  );


  buf

  (
    G3520,
    n366_inv_n
  );


  buf

  (
    G3521,
    g436_p
  );


  buf

  (
    G3522,
    g457_p
  );


  buf

  (
    G3523,
    g468_n
  );


  buf

  (
    G3524,
    g469_p
  );


  buf

  (
    G3525,
    g471_n
  );


  buf

  (
    G3526,
    n1000_o2_p
  );


  buf

  (
    G3527,
    g474_n
  );


  buf

  (
    G3528,
    g477_n_spl_
  );


  buf

  (
    G3529,
    g480_n_spl_
  );


  buf

  (
    G3530,
    g502_n
  );


  buf

  (
    G3531,
    g505_n_spl_
  );


  buf

  (
    G3532,
    g508_n_spl_
  );


  buf

  (
    G3533,
    g511_n_spl_
  );


  buf

  (
    G3534,
    n1380_o2_p
  );


  buf

  (
    G3535,
    n1425_o2_p
  );


  buf

  (
    G3536,
    g514_n_spl_
  );


  buf

  (
    G3537,
    g520_n_spl_
  );


  not

  (
    G3538,
    g524_p
  );


  buf

  (
    G3539,
    g544_n
  );


  buf

  (
    G3540,
    g550_p
  );


  buf

  (
    n4070_li003_li003,
    n2579_o2_p_spl_
  );


  buf

  (
    n4094_li011_li011,
    n2580_o2_p_spl_
  );


  buf

  (
    n4142_li027_li027,
    n2793_o2_p_spl_1
  );


  buf

  (
    n4154_li031_li031,
    n2794_o2_p_spl_
  );


  buf

  (
    n4166_li035_li035,
    n2729_o2_p
  );


  buf

  (
    n4178_li039_li039,
    n2730_o2_p
  );


  buf

  (
    n4190_li043_li043,
    n2621_o2_p_spl_
  );


  buf

  (
    n4202_li047_li047,
    n2622_o2_p_spl_
  );


  buf

  (
    n4214_li051_li051,
    n2623_o2_p_spl_
  );


  buf

  (
    n4226_li055_li055,
    n2624_o2_p_spl_
  );


  buf

  (
    n4229_li056_li056,
    G15_p
  );


  buf

  (
    n4232_li057_li057,
    n1911_lo_p
  );


  buf

  (
    n4241_li060_li060,
    G16_p
  );


  buf

  (
    n4244_li061_li061,
    n1923_lo_p
  );


  buf

  (
    n4253_li064_li064,
    G17_p
  );


  buf

  (
    n4256_li065_li065,
    n1935_lo_p
  );


  buf

  (
    n4265_li068_li068,
    G18_p
  );


  buf

  (
    n4268_li069_li069,
    n1947_lo_p
  );


  buf

  (
    n4277_li072_li072,
    G19_p
  );


  buf

  (
    n4280_li073_li073,
    n1959_lo_p
  );


  buf

  (
    n4289_li076_li076,
    G20_p
  );


  buf

  (
    n4292_li077_li077,
    n1971_lo_p
  );


  buf

  (
    n4301_li080_li080,
    G21_p
  );


  buf

  (
    n4313_li084_li084,
    G22_p
  );


  buf

  (
    n4373_li104_li104,
    G27_p
  );


  buf

  (
    n4382_li107_li107,
    n3069_o2_p
  );


  buf

  (
    n4385_li108_li108,
    G28_p
  );


  buf

  (
    n4397_li112_li112,
    G29_p
  );


  buf

  (
    n4418_li119_li119,
    n2757_o2_p
  );


  buf

  (
    n4430_li123_li123,
    n2731_o2_p
  );


  buf

  (
    n4442_li127_li127,
    n2674_o2_p
  );


  buf

  (
    n4454_li131_li131,
    n2625_o2_p
  );


  buf

  (
    n4466_li135_li135,
    n2626_o2_p
  );


  buf

  (
    n4478_li139_li139,
    n2644_o2_p
  );


  buf

  (
    n4490_li143_li143,
    n2675_o2_p
  );


  buf

  (
    n4502_li147_li147,
    n2758_o2_p
  );


  buf

  (
    n4553_li164_li164,
    G42_p
  );


  buf

  (
    n4556_li165_li165,
    n2235_lo_p
  );


  buf

  (
    n4565_li168_li168,
    G43_p
  );


  buf

  (
    n4568_li169_li169,
    n2247_lo_p
  );


  buf

  (
    n4577_li172_li172,
    G44_p
  );


  buf

  (
    n4580_li173_li173,
    n2259_lo_p
  );


  buf

  (
    n4589_li176_li176,
    G45_p
  );


  buf

  (
    n4592_li177_li177,
    n2271_lo_p
  );


  buf

  (
    n4601_li180_li180,
    G46_p
  );


  buf

  (
    n4604_li181_li181,
    n2283_lo_p
  );


  buf

  (
    n4607_li182_li182,
    n2286_lo_p
  );


  buf

  (
    n4613_li184_li184,
    G47_p
  );


  buf

  (
    n4616_li185_li185,
    n2295_lo_p
  );


  buf

  (
    n4622_li187_li187,
    lo186_buf_o2_p_spl_1
  );


  buf

  (
    n4625_li188_li188,
    G48_p
  );


  buf

  (
    n4634_li191_li191,
    n3142_o2_p
  );


  buf

  (
    n4649_li196_li196,
    G50_p
  );


  buf

  (
    n4652_li197_li197,
    n2331_lo_p
  );


  buf

  (
    n4655_li198_li198,
    n2334_lo_p
  );


  buf

  (
    n4658_li199_li199,
    n2337_lo_p
  );


  buf

  (
    n2071_i2,
    n327_inv_p_spl_
  );


  buf

  (
    n2080_i2,
    n2658_o2_p
  );


  buf

  (
    n2137_i2,
    n351_inv_p
  );


  buf

  (
    n2368_i2,
    n402_inv_p
  );


  buf

  (
    n2383_i2,
    n408_inv_p
  );


  buf

  (
    n2405_i2,
    n2947_o2_p
  );


  buf

  (
    n2471_i2,
    n3028_o2_p_spl_
  );


  buf

  (
    n2617_i2,
    n870_o2_p
  );


  buf

  (
    n2765_i2,
    n555_inv_p
  );


  buf

  (
    n2775_i2,
    n558_inv_p
  );


  buf

  (
    n2829_i2,
    n1003_o2_p_spl_1
  );


  buf

  (
    n2579_i2,
    n2992_o2_p
  );


  buf

  (
    n2580_i2,
    n2993_o2_p_spl_1
  );


  buf

  (
    n2618_i2,
    n3086_o2_p_spl_
  );


  buf

  (
    n2619_i2,
    n3087_o2_p_spl_
  );


  buf

  (
    n2620_i2,
    n3088_o2_p
  );


  buf

  (
    n2621_i2,
    n3089_o2_p_spl_
  );


  buf

  (
    n2622_i2,
    n3090_o2_p_spl_
  );


  buf

  (
    n2623_i2,
    n3091_o2_p_spl_
  );


  buf

  (
    n2624_i2,
    n3092_o2_p_spl_
  );


  buf

  (
    n2625_i2,
    n3093_o2_p
  );


  buf

  (
    n2626_i2,
    n3094_o2_p
  );


  buf

  (
    n2627_i2,
    n3095_o2_p_spl_
  );


  buf

  (
    n3029_i2,
    n744_inv_p
  );


  buf

  (
    n3035_i2,
    n1144_o2_p
  );


  buf

  (
    n2643_i2,
    n3170_o2_p_spl_
  );


  buf

  (
    n2644_i2,
    n3171_o2_p
  );


  buf

  (
    n2645_i2,
    n3172_o2_p
  );


  buf

  (
    n2640_i2,
    n483_inv_p
  );


  buf

  (
    n2658_i2,
    n3179_o2_p
  );


  buf

  (
    n2659_i2,
    n498_inv_p
  );


  buf

  (
    n2674_i2,
    n3211_o2_p
  );


  buf

  (
    n2675_i2,
    n3212_o2_p
  );


  buf

  (
    n2676_i2,
    n3213_o2_p_spl_
  );


  buf

  (
    n3119_i2,
    n1147_o2_p_spl_
  );


  buf

  (
    n3153_i2,
    n945_inv_p_spl_
  );


  buf

  (
    n2681_i2,
    n513_inv_p
  );


  buf

  (
    n2729_i2,
    n3245_o2_p_spl_1
  );


  buf

  (
    n2730_i2,
    n3246_o2_p_spl_1
  );


  buf

  (
    n2731_i2,
    n3247_o2_p
  );


  not

  (
    n698_i2,
    g551_n_spl_
  );


  not

  (
    n677_i2,
    g552_n_spl_
  );


  buf

  (
    n2757_i2,
    lo118_buf_o2_p
  );


  buf

  (
    n2758_i2,
    lo146_buf_o2_p
  );


  buf

  (
    n1000_i2,
    g553_p_spl_
  );


  buf

  (
    n1160_i2,
    g554_n_spl_
  );


  buf

  (
    n1153_i2,
    g555_p_spl_
  );


  buf

  (
    n2793_i2,
    lo026_buf_o2_p_spl_
  );


  buf

  (
    n2794_i2,
    lo030_buf_o2_p_spl_
  );


  buf

  (
    n2795_i2,
    lo090_buf_o2_p
  );


  buf

  (
    n1001_i2,
    g556_p_spl_
  );


  buf

  (
    n2859_i2,
    n697_o2_p
  );


  buf

  (
    n744_i2,
    g559_n_spl_
  );


  buf

  (
    n2908_i2,
    n645_inv_p
  );


  buf

  (
    n2926_i2,
    n826_o2_p
  );


  buf

  (
    n2928_i2,
    n654_inv_p
  );


  buf

  (
    n2966_i2,
    lo082_buf_o2_p_spl_
  );


  buf

  (
    n2967_i2,
    lo086_buf_o2_p_spl_
  );


  buf

  (
    n2947_i2,
    n700_o2_p
  );


  buf

  (
    n1010_i2,
    g562_p_spl_1
  );


  buf

  (
    n2976_i2,
    n675_inv_p_spl_
  );


  buf

  (
    n3069_i2,
    lo106_buf_o2_p
  );


  buf

  (
    n3028_i2,
    n701_o2_p
  );


  buf

  (
    n3081_i2,
    n841_o2_p_spl_
  );


  buf

  (
    n3082_i2,
    n867_o2_p
  );


  buf

  (
    n3142_i2,
    lo190_buf_o2_p
  );


  buf

  (
    n3214_i2,
    n1059_inv_p_spl_11
  );


  buf

  (
    n2992_i2,
    lo002_buf_o2_p_spl_1
  );


  buf

  (
    n2993_i2,
    lo010_buf_o2_p_spl_1
  );


  buf

  (
    n870_i2,
    g563_p_spl_
  );


  buf

  (
    n3086_i2,
    lo006_buf_o2_p_spl_
  );


  buf

  (
    n3087_i2,
    lo014_buf_o2_p_spl_1
  );


  buf

  (
    n3088_i2,
    lo022_buf_o2_p_spl_
  );


  buf

  (
    n3089_i2,
    lo042_buf_o2_p_spl_1
  );


  buf

  (
    n3090_i2,
    lo046_buf_o2_p_spl_1
  );


  buf

  (
    n3091_i2,
    lo050_buf_o2_p_spl_
  );


  buf

  (
    n3092_i2,
    lo054_buf_o2_p_spl_1
  );


  buf

  (
    n3093_i2,
    lo130_buf_o2_p
  );


  buf

  (
    n3094_i2,
    lo134_buf_o2_p
  );


  buf

  (
    n3095_i2,
    lo154_buf_o2_p_spl_
  );


  buf

  (
    n3136_i2,
    n906_inv_p
  );


  buf

  (
    n3170_i2,
    lo018_buf_o2_p_spl_
  );


  buf

  (
    n3171_i2,
    lo138_buf_o2_p_spl_
  );


  buf

  (
    n3172_i2,
    lo158_buf_o2_p
  );


  buf

  (
    n3179_i2,
    n728_o2_p
  );


  buf

  (
    n3180_i2,
    n993_inv_p
  );


  buf

  (
    n3193_i2,
    n770_o2_p
  );


  buf

  (
    n3211_i2,
    lo126_buf_o2_p
  );


  buf

  (
    n3212_i2,
    lo142_buf_o2_p_spl_
  );


  buf

  (
    n3213_i2,
    lo162_buf_o2_p
  );


  buf

  (
    n3219_i2,
    n1068_inv_p
  );


  buf

  (
    n1125_i2,
    g567_p_spl_
  );


  buf

  (
    n1081_i2,
    g572_p_spl_
  );


  buf

  (
    n1139_i2,
    g577_p_spl_
  );


  buf

  (
    n3245_i2,
    lo034_buf_o2_p_spl_1
  );


  buf

  (
    n3246_i2,
    lo038_buf_o2_p_spl_1
  );


  buf

  (
    n3247_i2,
    lo122_buf_o2_p_spl_
  );


  buf

  (
    lo074_buf_i2,
    n1962_lo_p_spl_
  );


  buf

  (
    lo078_buf_i2,
    n1974_lo_p_spl_
  );


  buf

  (
    lo186_buf_i2,
    n2298_lo_p_spl_
  );


  buf

  (
    lo118_buf_i2,
    lo117_buf_o2_p_spl_
  );


  buf

  (
    lo146_buf_i2,
    lo145_buf_o2_p_spl_
  );


  not

  (
    n1038_i2,
    g581_n_spl_1
  );


  buf

  (
    n1044_i2,
    g583_n_spl_1
  );


  buf

  (
    n980_i2,
    g589_n_spl_
  );


  buf

  (
    n1145_i2,
    g590_p_spl_
  );


  buf

  (
    lo026_buf_i2,
    lo024_buf_o2_p_spl_1
  );


  buf

  (
    lo030_buf_i2,
    lo028_buf_o2_p_spl_1
  );


  buf

  (
    lo090_buf_i2,
    lo088_buf_o2_p_spl_
  );


  buf

  (
    lo094_buf_i2,
    lo092_buf_o2_p_spl_
  );


  buf

  (
    lo098_buf_i2,
    lo096_buf_o2_p_spl_
  );


  buf

  (
    lo102_buf_i2,
    lo100_buf_o2_p_spl_
  );


  buf

  (
    lo066_buf_i2,
    n1938_lo_p_spl_
  );


  buf

  (
    lo070_buf_i2,
    n1950_lo_p_spl_
  );


  not

  (
    n1202_i2,
    g591_n_spl_
  );


  buf

  (
    n1003_i2,
    g592_p
  );


  buf

  (
    n1031_i2,
    g595_n_spl_
  );


  buf

  (
    n1034_i2,
    g597_p_spl_
  );


  buf

  (
    n1040_i2,
    g598_p_spl_
  );


  buf

  (
    n1046_i2,
    g599_p_spl_
  );


  buf

  (
    n1380_i2,
    g621_n_spl_
  );


  buf

  (
    n1425_i2,
    g645_n_spl_
  );


  buf

  (
    n697_i2,
    g646_n_spl_
  );


  buf

  (
    n1143_i2,
    g656_p_spl_
  );


  buf

  (
    n673_i2,
    g657_n_spl_
  );


  buf

  (
    n789_i2,
    g658_n_spl_
  );


  buf

  (
    n786_i2,
    g659_n_spl_1
  );


  not

  (
    n1047_i2,
    g660_p_spl_
  );


  buf

  (
    n1036_i2,
    g661_n_spl_
  );


  not

  (
    n1307_i2,
    g662_n_spl_
  );


  not

  (
    n1035_i2,
    g663_p_spl_
  );


  not

  (
    n1297_i2,
    g664_n_spl_
  );


  buf

  (
    n1099_i2,
    g665_n_spl_
  );


  buf

  (
    n1128_i2,
    g666_p_spl_
  );


  buf

  (
    n674_i2,
    g667_n_spl_
  );


  buf

  (
    n826_i2,
    g676_n_spl_
  );


  buf

  (
    n853_i2,
    g684_n_spl_
  );


  buf

  (
    n951_i2,
    g686_p_spl_
  );


  buf

  (
    n700_i2,
    g687_n_spl_
  );


  buf

  (
    n884_i2,
    g691_p_spl_
  );


  buf

  (
    lo082_buf_i2,
    n1983_lo_p_spl_
  );


  buf

  (
    lo086_buf_i2,
    n1995_lo_p_spl_
  );


  buf

  (
    n801_i2,
    g701_n_spl_
  );


  not

  (
    n840_i2,
    g707_n_spl_
  );


  not

  (
    n866_i2,
    g713_n_spl_
  );


  buf

  (
    lo002_buf_i2,
    G1_p_spl_
  );


  buf

  (
    lo010_buf_i2,
    G3_p_spl_1
  );


  buf

  (
    lo166_buf_i2,
    n2238_lo_p_spl_
  );


  buf

  (
    lo170_buf_i2,
    n2250_lo_p_spl_
  );


  not

  (
    n1426_i2,
    g714_n
  );


  not

  (
    n1082_i2,
    g715_n
  );


  buf

  (
    n1310_i2,
    g716_p_spl_
  );


  not

  (
    n1015_i2,
    g718_n
  );


  not

  (
    n1206_i2,
    g719_n_spl_
  );


  buf

  (
    n1262_i2,
    g720_n_spl_
  );


  buf

  (
    n1456_i2,
    g721_p
  );


  buf

  (
    n1244_i2,
    g739_p
  );


  buf

  (
    n1280_i2,
    g740_p
  );


  buf

  (
    n1290_i2,
    g741_p
  );


  buf

  (
    n1012_i2,
    g743_n
  );


  not

  (
    n1074_i2,
    g783_n
  );


  not

  (
    n1112_i2,
    g810_n
  );


  buf

  (
    n1212_i2,
    g838_p
  );


  buf

  (
    n1454_i2,
    g869_p
  );


  not

  (
    n1182_i2,
    g874_n
  );


  not

  (
    n1220_i2,
    g875_n_spl_
  );


  buf

  (
    n701_i2,
    g876_n_spl_
  );


  not

  (
    n973_i2,
    g886_n_spl_
  );


  buf

  (
    n1282_i2,
    g889_p
  );


  not

  (
    n1144_i2,
    g890_n_spl_
  );


  buf

  (
    n1278_i2,
    g916_p
  );


  buf

  (
    n1459_i2,
    g919_n
  );


  buf

  (
    n1324_i2,
    g945_p
  );


  buf

  (
    n1288_i2,
    g948_n
  );


  buf

  (
    n1271_i2,
    g950_n_spl_
  );


  buf

  (
    n1132_i2,
    g956_n
  );


  buf

  (
    n1231_i2,
    g966_n
  );


  buf

  (
    n1462_i2,
    g967_n
  );


  buf

  (
    n1482_i2,
    g968_p
  );


  not

  (
    n994_i2,
    g972_n_spl_
  );


  not

  (
    n998_i2,
    g976_n_spl_
  );


  buf

  (
    lo106_buf_i2,
    n2055_lo_p
  );


  buf

  (
    n769_i2,
    g985_n_spl_
  );


  not

  (
    n814_i2,
    g992_n_spl_
  );


  buf

  (
    n841_i2,
    g995_p_spl_
  );


  buf

  (
    n867_i2,
    g998_p_spl_
  );


  buf

  (
    lo006_buf_i2,
    G2_p
  );


  buf

  (
    lo014_buf_i2,
    G4_p_spl_11
  );


  buf

  (
    lo022_buf_i2,
    G6_p_spl_
  );


  buf

  (
    lo042_buf_i2,
    G11_p_spl_
  );


  buf

  (
    lo046_buf_i2,
    G12_p_spl_1
  );


  buf

  (
    lo050_buf_i2,
    G13_p_spl_
  );


  buf

  (
    lo054_buf_i2,
    G14_p_spl_
  );


  buf

  (
    lo130_buf_i2,
    G33_p_spl_
  );


  buf

  (
    lo134_buf_i2,
    G34_p_spl_
  );


  buf

  (
    lo154_buf_i2,
    G39_p
  );


  buf

  (
    lo174_buf_i2,
    n2262_lo_p
  );


  buf

  (
    lo178_buf_i2,
    n2274_lo_p
  );


  buf

  (
    n1007_i2,
    g999_n
  );


  buf

  (
    n1294_i2,
    g1000_p
  );


  buf

  (
    n1084_i2,
    g1001_p
  );


  not

  (
    n1399_i2,
    g1002_p
  );


  buf

  (
    n1311_i2,
    g1003_p
  );


  not

  (
    n1392_i2,
    g1005_n
  );


  buf

  (
    n1102_i2,
    g1006_p
  );


  buf

  (
    n1041_i2,
    g1007_p
  );


  buf

  (
    n1298_i2,
    g1008_p
  );


  buf

  (
    n738_i2,
    g1010_p
  );


  buf

  (
    n1214_i2,
    g1011_p
  );


  buf

  (
    n1222_i2,
    g1012_p
  );


  not

  (
    n1155_i2,
    g1014_n
  );


  buf

  (
    n1147_i2,
    g1015_p
  );


  buf

  (
    n1393_i2,
    g1016_p
  );


  not

  (
    n999_i2,
    g1017_n
  );


  buf

  (
    n1306_i2,
    g1018_p
  );


  buf

  (
    n1312_i2,
    g1019_p
  );


  not

  (
    n1382_i2,
    g1021_p
  );


  not

  (
    n1383_i2,
    g1022_n
  );


  not

  (
    n1152_i2,
    g1023_p
  );


  not

  (
    n1334_i2,
    g1032_n
  );


  buf

  (
    n1335_i2,
    g1033_p
  );


  not

  (
    n695_i2,
    g1034_n_spl_
  );


  buf

  (
    n773_i2,
    g1035_n_spl_
  );


  buf

  (
    lo190_buf_i2,
    n2307_lo_p
  );


  buf

  (
    n1368_i2,
    g1037_p
  );


  not

  (
    n1362_i2,
    g1044_n
  );


  buf

  (
    n1406_i2,
    g1046_p
  );


  not

  (
    n1403_i2,
    g1050_n
  );


  buf

  (
    n741_i2,
    g1053_p
  );


  buf

  (
    n1407_i2,
    g1054_p
  );


  buf

  (
    n1395_i2,
    g1058_n
  );


  buf

  (
    n1359_i2,
    g1063_n
  );


  buf

  (
    n1159_i2,
    g1066_n
  );


  not

  (
    n1221_i2,
    g1067_p
  );


  not

  (
    n987_i2,
    g1073_p
  );


  not

  (
    n989_i2,
    g1074_n_spl_
  );


  buf

  (
    n881_i2,
    g1085_n_spl_
  );


  buf

  (
    n1340_i2,
    g1089_n
  );


  buf

  (
    n1341_i2,
    g1090_p
  );


  buf

  (
    n906_i2,
    g1098_n_spl_
  );


  buf

  (
    n1388_i2,
    g1101_n
  );


  not

  (
    n791_i2,
    g1110_n_spl_
  );


  not

  (
    n1372_i2,
    g1117_n
  );


  buf

  (
    n815_i2,
    g1120_p_spl_
  );


  buf

  (
    n868_i2,
    g1121_p_spl_
  );


  buf

  (
    lo018_buf_i2,
    G5_p_spl_
  );


  buf

  (
    lo138_buf_i2,
    G35_p_spl_
  );


  buf

  (
    lo158_buf_i2,
    G40_p_spl_
  );


  buf

  (
    n780_i2,
    g1122_n_spl_1
  );


  buf

  (
    n728_i2,
    g1123_n_spl_
  );


  buf

  (
    n676_i2,
    g1124_n_spl_
  );


  buf

  (
    n929_i2,
    g1130_p
  );


  buf

  (
    n955_i2,
    g1136_p
  );


  buf

  (
    n938_i2,
    g1144_p
  );


  buf

  (
    n1117_i2,
    g1148_p
  );


  buf

  (
    n1121_i2,
    g1152_p
  );


  buf

  (
    n965_i2,
    g1161_n
  );


  not

  (
    n752_i2,
    g1162_n_spl_1
  );


  not

  (
    n753_i2,
    g1162_n_spl_1
  );


  not

  (
    n760_i2,
    g1163_n_spl_
  );


  buf

  (
    n770_i2,
    g1164_p_spl_
  );


  buf

  (
    n923_i2,
    g1167_p
  );


  buf

  (
    n947_i2,
    g1170_p
  );


  buf

  (
    n897_i2,
    g1181_p
  );


  buf

  (
    n919_i2,
    g1192_p
  );


  buf

  (
    n895_i2,
    g1194_n
  );


  buf

  (
    n917_i2,
    g1196_n
  );


  not

  (
    n751_i2,
    g1200_p_spl_
  );


  buf

  (
    n774_i2,
    g1201_n_spl_
  );


  buf

  (
    lo126_buf_i2,
    G32_p
  );


  buf

  (
    lo142_buf_i2,
    G36_p
  );


  buf

  (
    lo162_buf_i2,
    G41_p_spl_
  );


  not

  (
    n990_i2,
    g1202_n
  );


  buf

  (
    n792_i2,
    g1205_p
  );


  buf

  (
    n869_i2,
    g1206_p
  );


  buf

  (
    n848_i2,
    g1208_p_spl_
  );


  buf

  (
    lo024_buf_i2,
    G7_p
  );


  buf

  (
    lo028_buf_i2,
    G8_p
  );


  buf

  (
    lo088_buf_i2,
    G23_p
  );


  buf

  (
    lo092_buf_i2,
    G24_p
  );


  buf

  (
    lo096_buf_i2,
    G25_p
  );


  buf

  (
    lo100_buf_i2,
    G26_p
  );


  buf

  (
    n763_i2,
    g1209_p
  );


  buf

  (
    n754_i2,
    g1210_n_spl_
  );


  buf

  (
    n755_i2,
    g1210_n_spl_
  );


  buf

  (
    n822_i2,
    g1212_p
  );


  buf

  (
    n849_i2,
    g1213_p
  );


  buf

  (
    n777_i2,
    g1214_n
  );


  buf

  (
    n778_i2,
    g1215_p
  );


  not

  (
    n820_i2,
    g1216_n
  );


  not

  (
    n846_i2,
    g1217_n
  );


  not

  (
    n806_i2,
    g1218_n
  );


  not

  (
    n771_i2,
    g1219_n
  );


  buf

  (
    n854_i2,
    g1220_p
  );


  not

  (
    n828_i2,
    g1221_n
  );


  buf

  (
    lo117_buf_i2,
    G30_p
  );


  buf

  (
    lo145_buf_i2,
    G37_p
  );


  not

  (
    n762_i2,
    g1222_p
  );


  buf

  (
    n805_i2,
    g1225_p
  );


  not

  (
    n859_i2,
    g1230_p
  );


  buf

  (
    n833_i2,
    g1235_n
  );


  buf

  (
    lo034_buf_i2,
    G9_p
  );


  buf

  (
    lo038_buf_i2,
    G10_p
  );


  buf

  (
    lo122_buf_i2,
    G31_p
  );


  buf

  (
    lo150_buf_i2,
    G38_p
  );


  buf

  (
    n1860_lo_n_spl_,
    n1860_lo_n
  );


  buf

  (
    n1776_lo_n_spl_,
    n1776_lo_n
  );


  buf

  (
    n1752_lo_n_spl_,
    n1752_lo_n
  );


  buf

  (
    n2148_lo_n_spl_,
    n2148_lo_n
  );


  buf

  (
    n2148_lo_n_spl_0,
    n2148_lo_n_spl_
  );


  buf

  (
    n2148_lo_n_spl_1,
    n2148_lo_n_spl_
  );


  buf

  (
    n1872_lo_p_spl_,
    n1872_lo_p
  );


  buf

  (
    n2124_lo_n_spl_,
    n2124_lo_n
  );


  buf

  (
    n2124_lo_n_spl_0,
    n2124_lo_n_spl_
  );


  buf

  (
    n2100_lo_n_spl_,
    n2100_lo_n
  );


  buf

  (
    n2100_lo_n_spl_0,
    n2100_lo_n_spl_
  );


  buf

  (
    n1824_lo_p_spl_,
    n1824_lo_p
  );


  buf

  (
    n2136_lo_n_spl_,
    n2136_lo_n
  );


  buf

  (
    n2136_lo_n_spl_0,
    n2136_lo_n_spl_
  );


  buf

  (
    n2184_lo_n_spl_,
    n2184_lo_n
  );


  buf

  (
    n2184_lo_n_spl_0,
    n2184_lo_n_spl_
  );


  buf

  (
    n1908_lo_p_spl_,
    n1908_lo_p
  );


  buf

  (
    n1908_lo_p_spl_0,
    n1908_lo_p_spl_
  );


  buf

  (
    n2112_lo_n_spl_,
    n2112_lo_n
  );


  buf

  (
    n2112_lo_n_spl_0,
    n2112_lo_n_spl_
  );


  buf

  (
    n2160_lo_n_spl_,
    n2160_lo_n
  );


  buf

  (
    n2160_lo_n_spl_0,
    n2160_lo_n_spl_
  );


  buf

  (
    n2160_lo_n_spl_1,
    n2160_lo_n_spl_
  );


  buf

  (
    n1884_lo_p_spl_,
    n1884_lo_p
  );


  buf

  (
    n2172_lo_n_spl_,
    n2172_lo_n
  );


  buf

  (
    n2172_lo_n_spl_0,
    n2172_lo_n_spl_
  );


  buf

  (
    n2172_lo_n_spl_1,
    n2172_lo_n_spl_
  );


  buf

  (
    n1896_lo_p_spl_,
    n1896_lo_p
  );


  buf

  (
    n1896_lo_p_spl_0,
    n1896_lo_p_spl_
  );


  buf

  (
    g430_n_spl_,
    g430_n
  );


  buf

  (
    n2172_lo_p_spl_,
    n2172_lo_p
  );


  buf

  (
    n2184_lo_p_spl_,
    n2184_lo_p
  );


  buf

  (
    n2148_lo_p_spl_,
    n2148_lo_p
  );


  buf

  (
    n2160_lo_p_spl_,
    n2160_lo_p
  );


  buf

  (
    g442_p_spl_,
    g442_p
  );


  buf

  (
    g439_n_spl_,
    g439_n
  );


  buf

  (
    g442_n_spl_,
    g442_n
  );


  buf

  (
    g439_p_spl_,
    g439_p
  );


  buf

  (
    n2124_lo_p_spl_,
    n2124_lo_p
  );


  buf

  (
    n2136_lo_p_spl_,
    n2136_lo_p
  );


  buf

  (
    n2100_lo_p_spl_,
    n2100_lo_p
  );


  buf

  (
    n2112_lo_p_spl_,
    n2112_lo_p
  );


  buf

  (
    g451_n_spl_,
    g451_n
  );


  buf

  (
    g448_p_spl_,
    g448_p
  );


  buf

  (
    g451_p_spl_,
    g451_p
  );


  buf

  (
    g448_n_spl_,
    g448_n
  );


  buf

  (
    n1908_lo_n_spl_,
    n1908_lo_n
  );


  buf

  (
    n1908_lo_n_spl_0,
    n1908_lo_n_spl_
  );


  buf

  (
    n1896_lo_n_spl_,
    n1896_lo_n
  );


  buf

  (
    g462_p_spl_,
    g462_p
  );


  buf

  (
    g459_p_spl_,
    g459_p
  );


  buf

  (
    g462_n_spl_,
    g462_n
  );


  buf

  (
    g459_n_spl_,
    g459_n
  );


  buf

  (
    n3029_o2_p_spl_,
    n3029_o2_p
  );


  buf

  (
    n1001_o2_n_spl_,
    n1001_o2_n
  );


  buf

  (
    n1001_o2_n_spl_0,
    n1001_o2_n_spl_
  );


  buf

  (
    n1010_o2_n_spl_,
    n1010_o2_n
  );


  buf

  (
    n1010_o2_p_spl_,
    n1010_o2_p
  );


  buf

  (
    g481_n_spl_,
    g481_n
  );


  buf

  (
    n3119_o2_p_spl_,
    n3119_o2_p
  );


  buf

  (
    g481_p_spl_,
    g481_p
  );


  buf

  (
    n3119_o2_n_spl_,
    n3119_o2_n
  );


  buf

  (
    n1153_o2_p_spl_,
    n1153_o2_p
  );


  buf

  (
    n1160_o2_p_spl_,
    n1160_o2_p
  );


  buf

  (
    n1153_o2_n_spl_,
    n1153_o2_n
  );


  buf

  (
    n1160_o2_n_spl_,
    n1160_o2_n
  );


  buf

  (
    n1001_o2_p_spl_,
    n1001_o2_p
  );


  buf

  (
    g514_p_spl_,
    g514_p
  );


  buf

  (
    g480_p_spl_,
    g480_p
  );


  buf

  (
    g514_n_spl_,
    g514_n
  );


  buf

  (
    g514_n_spl_0,
    g514_n_spl_
  );


  buf

  (
    g480_n_spl_,
    g480_n
  );


  buf

  (
    g480_n_spl_0,
    g480_n_spl_
  );


  buf

  (
    g511_p_spl_,
    g511_p
  );


  buf

  (
    g505_p_spl_,
    g505_p
  );


  buf

  (
    g511_n_spl_,
    g511_n
  );


  buf

  (
    g511_n_spl_0,
    g511_n_spl_
  );


  buf

  (
    g505_n_spl_,
    g505_n
  );


  buf

  (
    g505_n_spl_0,
    g505_n_spl_
  );


  buf

  (
    g508_p_spl_,
    g508_p
  );


  buf

  (
    g477_p_spl_,
    g477_p
  );


  buf

  (
    g508_n_spl_,
    g508_n
  );


  buf

  (
    g508_n_spl_0,
    g508_n_spl_
  );


  buf

  (
    g477_n_spl_,
    g477_n
  );


  buf

  (
    g477_n_spl_0,
    g477_n_spl_
  );


  buf

  (
    g517_n_spl_,
    g517_n
  );


  buf

  (
    g516_n_spl_,
    g516_n
  );


  buf

  (
    g515_n_spl_,
    g515_n
  );


  buf

  (
    n1462_o2_p_spl_,
    n1462_o2_p
  );


  buf

  (
    n1462_o2_p_spl_0,
    n1462_o2_p_spl_
  );


  buf

  (
    n2064_lo_p_spl_,
    n2064_lo_p
  );


  buf

  (
    g521_n_spl_,
    g521_n
  );


  buf

  (
    g520_n_spl_,
    g520_n
  );


  buf

  (
    g528_n_spl_,
    g528_n
  );


  buf

  (
    g526_p_spl_,
    g526_p
  );


  buf

  (
    g528_p_spl_,
    g528_p
  );


  buf

  (
    g526_n_spl_,
    g526_n
  );


  buf

  (
    g534_n_spl_,
    g534_n
  );


  buf

  (
    g534_n_spl_0,
    g534_n_spl_
  );


  buf

  (
    g534_n_spl_1,
    g534_n_spl_
  );


  buf

  (
    n2340_lo_p_spl_,
    n2340_lo_p
  );


  buf

  (
    g534_p_spl_,
    g534_p
  );


  buf

  (
    g534_p_spl_0,
    g534_p_spl_
  );


  buf

  (
    g534_p_spl_1,
    g534_p_spl_
  );


  buf

  (
    n2340_lo_n_spl_,
    n2340_lo_n
  );


  buf

  (
    g538_p_spl_,
    g538_p
  );


  buf

  (
    g533_p_spl_,
    g533_p
  );


  buf

  (
    g533_p_spl_0,
    g533_p_spl_
  );


  buf

  (
    g533_p_spl_1,
    g533_p_spl_
  );


  buf

  (
    g538_n_spl_,
    g538_n
  );


  buf

  (
    g533_n_spl_,
    g533_n
  );


  buf

  (
    g533_n_spl_0,
    g533_n_spl_
  );


  buf

  (
    g533_n_spl_1,
    g533_n_spl_
  );


  buf

  (
    g531_n_spl_,
    g531_n
  );


  buf

  (
    g531_p_spl_,
    g531_p
  );


  buf

  (
    n2793_o2_p_spl_,
    n2793_o2_p
  );


  buf

  (
    n2793_o2_p_spl_0,
    n2793_o2_p_spl_
  );


  buf

  (
    n2793_o2_p_spl_1,
    n2793_o2_p_spl_
  );


  buf

  (
    n2621_o2_n_spl_,
    n2621_o2_n
  );


  buf

  (
    n994_o2_n_spl_,
    n994_o2_n
  );


  buf

  (
    n994_o2_n_spl_0,
    n994_o2_n_spl_
  );


  buf

  (
    n994_o2_p_spl_,
    n994_o2_p
  );


  buf

  (
    n945_inv_p_spl_,
    n945_inv_p
  );


  buf

  (
    n3028_o2_n_spl_,
    n3028_o2_n
  );


  buf

  (
    n3028_o2_p_spl_,
    n3028_o2_p
  );


  buf

  (
    n3028_o2_p_spl_0,
    n3028_o2_p_spl_
  );


  buf

  (
    n2620_o2_p_spl_,
    n2620_o2_p
  );


  buf

  (
    n1007_o2_p_spl_,
    n1007_o2_p
  );


  buf

  (
    n2620_o2_n_spl_,
    n2620_o2_n
  );


  buf

  (
    n2579_o2_p_spl_,
    n2579_o2_p
  );


  buf

  (
    g561_p_spl_,
    g561_p
  );


  buf

  (
    g556_p_spl_,
    g556_p
  );


  buf

  (
    g556_p_spl_0,
    g556_p_spl_
  );


  buf

  (
    g561_n_spl_,
    g561_n
  );


  buf

  (
    g561_n_spl_0,
    g561_n_spl_
  );


  buf

  (
    g561_n_spl_00,
    g561_n_spl_0
  );


  buf

  (
    g561_n_spl_01,
    g561_n_spl_0
  );


  buf

  (
    g561_n_spl_1,
    g561_n_spl_
  );


  buf

  (
    g556_n_spl_,
    g556_n
  );


  buf

  (
    g556_n_spl_0,
    g556_n_spl_
  );


  buf

  (
    g556_n_spl_1,
    g556_n_spl_
  );


  buf

  (
    n869_o2_p_spl_,
    n869_o2_p
  );


  buf

  (
    n792_o2_p_spl_,
    n792_o2_p
  );


  buf

  (
    n869_o2_n_spl_,
    n869_o2_n
  );


  buf

  (
    n792_o2_n_spl_,
    n792_o2_n
  );


  buf

  (
    n1059_inv_n_spl_,
    n1059_inv_n
  );


  buf

  (
    n1059_inv_n_spl_0,
    n1059_inv_n_spl_
  );


  buf

  (
    n1059_inv_n_spl_00,
    n1059_inv_n_spl_0
  );


  buf

  (
    n1059_inv_n_spl_000,
    n1059_inv_n_spl_00
  );


  buf

  (
    n1059_inv_n_spl_001,
    n1059_inv_n_spl_00
  );


  buf

  (
    n1059_inv_n_spl_01,
    n1059_inv_n_spl_0
  );


  buf

  (
    n1059_inv_n_spl_1,
    n1059_inv_n_spl_
  );


  buf

  (
    n1059_inv_n_spl_10,
    n1059_inv_n_spl_1
  );


  buf

  (
    n1059_inv_n_spl_11,
    n1059_inv_n_spl_1
  );


  buf

  (
    n1059_inv_p_spl_,
    n1059_inv_p
  );


  buf

  (
    n1059_inv_p_spl_0,
    n1059_inv_p_spl_
  );


  buf

  (
    n1059_inv_p_spl_00,
    n1059_inv_p_spl_0
  );


  buf

  (
    n1059_inv_p_spl_000,
    n1059_inv_p_spl_00
  );


  buf

  (
    n1059_inv_p_spl_001,
    n1059_inv_p_spl_00
  );


  buf

  (
    n1059_inv_p_spl_01,
    n1059_inv_p_spl_0
  );


  buf

  (
    n1059_inv_p_spl_010,
    n1059_inv_p_spl_01
  );


  buf

  (
    n1059_inv_p_spl_011,
    n1059_inv_p_spl_01
  );


  buf

  (
    n1059_inv_p_spl_1,
    n1059_inv_p_spl_
  );


  buf

  (
    n1059_inv_p_spl_10,
    n1059_inv_p_spl_1
  );


  buf

  (
    n1059_inv_p_spl_11,
    n1059_inv_p_spl_1
  );


  buf

  (
    g563_p_spl_,
    g563_p
  );


  buf

  (
    n897_o2_n_spl_,
    n897_o2_n
  );


  buf

  (
    n897_o2_n_spl_0,
    n897_o2_n_spl_
  );


  buf

  (
    n897_o2_p_spl_,
    n897_o2_p
  );


  buf

  (
    g569_n_spl_,
    g569_n
  );


  buf

  (
    g568_n_spl_,
    g568_n
  );


  buf

  (
    g568_n_spl_0,
    g568_n_spl_
  );


  buf

  (
    g569_p_spl_,
    g569_p
  );


  buf

  (
    g568_p_spl_,
    g568_p
  );


  buf

  (
    n919_o2_n_spl_,
    n919_o2_n
  );


  buf

  (
    n919_o2_n_spl_0,
    n919_o2_n_spl_
  );


  buf

  (
    n919_o2_p_spl_,
    n919_o2_p
  );


  buf

  (
    g574_n_spl_,
    g574_n
  );


  buf

  (
    g573_n_spl_,
    g573_n
  );


  buf

  (
    g573_n_spl_0,
    g573_n_spl_
  );


  buf

  (
    g574_p_spl_,
    g574_p
  );


  buf

  (
    g573_p_spl_,
    g573_p
  );


  buf

  (
    n2993_o2_p_spl_,
    n2993_o2_p
  );


  buf

  (
    n2993_o2_p_spl_0,
    n2993_o2_p_spl_
  );


  buf

  (
    n2993_o2_p_spl_00,
    n2993_o2_p_spl_0
  );


  buf

  (
    n2993_o2_p_spl_1,
    n2993_o2_p_spl_
  );


  buf

  (
    n2993_o2_n_spl_,
    n2993_o2_n
  );


  buf

  (
    n2993_o2_n_spl_0,
    n2993_o2_n_spl_
  );


  buf

  (
    g579_p_spl_,
    g579_p
  );


  buf

  (
    g579_p_spl_0,
    g579_p_spl_
  );


  buf

  (
    g579_p_spl_00,
    g579_p_spl_0
  );


  buf

  (
    g579_p_spl_01,
    g579_p_spl_0
  );


  buf

  (
    g579_p_spl_1,
    g579_p_spl_
  );


  buf

  (
    lo102_buf_o2_n_spl_,
    lo102_buf_o2_n
  );


  buf

  (
    g578_p_spl_,
    g578_p
  );


  buf

  (
    g578_p_spl_0,
    g578_p_spl_
  );


  buf

  (
    g578_p_spl_1,
    g578_p_spl_
  );


  buf

  (
    lo102_buf_o2_p_spl_,
    lo102_buf_o2_p
  );


  buf

  (
    n791_o2_n_spl_,
    n791_o2_n
  );


  buf

  (
    n814_o2_p_spl_,
    n814_o2_p
  );


  buf

  (
    n841_o2_p_spl_,
    n841_o2_p
  );


  buf

  (
    n675_inv_p_spl_,
    n675_inv_p
  );


  buf

  (
    g572_p_spl_,
    g572_p
  );


  buf

  (
    g572_p_spl_0,
    g572_p_spl_
  );


  buf

  (
    g567_p_spl_,
    g567_p
  );


  buf

  (
    g567_p_spl_0,
    g567_p_spl_
  );


  buf

  (
    lo026_buf_o2_n_spl_,
    lo026_buf_o2_n
  );


  buf

  (
    n1962_lo_p_spl_,
    n1962_lo_p
  );


  buf

  (
    n1962_lo_p_spl_0,
    n1962_lo_p_spl_
  );


  buf

  (
    g589_n_spl_,
    g589_n
  );


  buf

  (
    g593_n_spl_,
    g593_n
  );


  buf

  (
    g578_n_spl_,
    g578_n
  );


  buf

  (
    g593_p_spl_,
    g593_p
  );


  buf

  (
    g594_p_spl_,
    g594_p
  );


  buf

  (
    g579_n_spl_,
    g579_n
  );


  buf

  (
    g579_n_spl_0,
    g579_n_spl_
  );


  buf

  (
    g579_n_spl_1,
    g579_n_spl_
  );


  buf

  (
    g594_n_spl_,
    g594_n
  );


  buf

  (
    g596_p_spl_,
    g596_p
  );


  buf

  (
    g596_n_spl_,
    g596_n
  );


  buf

  (
    n1334_o2_n_spl_,
    n1334_o2_n
  );


  buf

  (
    n1334_o2_p_spl_,
    n1334_o2_p
  );


  buf

  (
    n1147_o2_p_spl_,
    n1147_o2_p
  );


  buf

  (
    lo186_buf_o2_p_spl_,
    lo186_buf_o2_p
  );


  buf

  (
    lo186_buf_o2_p_spl_0,
    lo186_buf_o2_p_spl_
  );


  buf

  (
    lo186_buf_o2_p_spl_1,
    lo186_buf_o2_p_spl_
  );


  buf

  (
    lo186_buf_o2_n_spl_,
    lo186_buf_o2_n
  );


  buf

  (
    lo186_buf_o2_n_spl_0,
    lo186_buf_o2_n_spl_
  );


  buf

  (
    lo186_buf_o2_n_spl_1,
    lo186_buf_o2_n_spl_
  );


  buf

  (
    g555_p_spl_,
    g555_p
  );


  buf

  (
    g603_n_spl_,
    g603_n
  );


  buf

  (
    g601_n_spl_,
    g601_n
  );


  buf

  (
    g601_n_spl_0,
    g601_n_spl_
  );


  buf

  (
    g603_p_spl_,
    g603_p
  );


  buf

  (
    g601_p_spl_,
    g601_p
  );


  buf

  (
    g604_n_spl_,
    g604_n
  );


  buf

  (
    g600_n_spl_,
    g600_n
  );


  buf

  (
    g600_n_spl_0,
    g600_n_spl_
  );


  buf

  (
    n2619_o2_n_spl_,
    n2619_o2_n
  );


  buf

  (
    n2619_o2_n_spl_0,
    n2619_o2_n_spl_
  );


  buf

  (
    n2619_o2_n_spl_00,
    n2619_o2_n_spl_0
  );


  buf

  (
    n2619_o2_n_spl_01,
    n2619_o2_n_spl_0
  );


  buf

  (
    n2619_o2_n_spl_1,
    n2619_o2_n_spl_
  );


  buf

  (
    n2619_o2_n_spl_10,
    n2619_o2_n_spl_1
  );


  buf

  (
    g609_n_spl_,
    g609_n
  );


  buf

  (
    g609_n_spl_0,
    g609_n_spl_
  );


  buf

  (
    g609_n_spl_1,
    g609_n_spl_
  );


  buf

  (
    n2580_o2_p_spl_,
    n2580_o2_p
  );


  buf

  (
    n327_inv_p_spl_,
    n327_inv_p
  );


  buf

  (
    g612_p_spl_,
    g612_p
  );


  buf

  (
    g612_p_spl_0,
    g612_p_spl_
  );


  buf

  (
    g612_p_spl_00,
    g612_p_spl_0
  );


  buf

  (
    g612_p_spl_01,
    g612_p_spl_0
  );


  buf

  (
    g612_p_spl_1,
    g612_p_spl_
  );


  buf

  (
    g612_p_spl_10,
    g612_p_spl_1
  );


  buf

  (
    g562_p_spl_,
    g562_p
  );


  buf

  (
    g562_p_spl_0,
    g562_p_spl_
  );


  buf

  (
    g562_p_spl_00,
    g562_p_spl_0
  );


  buf

  (
    g562_p_spl_01,
    g562_p_spl_0
  );


  buf

  (
    g562_p_spl_1,
    g562_p_spl_
  );


  buf

  (
    g562_p_spl_10,
    g562_p_spl_1
  );


  buf

  (
    g622_n_spl_,
    g622_n
  );


  buf

  (
    g622_n_spl_0,
    g622_n_spl_
  );


  buf

  (
    g554_n_spl_,
    g554_n
  );


  buf

  (
    g554_n_spl_0,
    g554_n_spl_
  );


  buf

  (
    g622_p_spl_,
    g622_p
  );


  buf

  (
    g554_p_spl_,
    g554_p
  );


  buf

  (
    lo034_buf_o2_p_spl_,
    lo034_buf_o2_p
  );


  buf

  (
    lo034_buf_o2_p_spl_0,
    lo034_buf_o2_p_spl_
  );


  buf

  (
    lo034_buf_o2_p_spl_00,
    lo034_buf_o2_p_spl_0
  );


  buf

  (
    lo034_buf_o2_p_spl_1,
    lo034_buf_o2_p_spl_
  );


  buf

  (
    lo028_buf_o2_p_spl_,
    lo028_buf_o2_p
  );


  buf

  (
    lo028_buf_o2_p_spl_0,
    lo028_buf_o2_p_spl_
  );


  buf

  (
    lo028_buf_o2_p_spl_1,
    lo028_buf_o2_p_spl_
  );


  buf

  (
    n965_o2_n_spl_,
    n965_o2_n
  );


  buf

  (
    n965_o2_p_spl_,
    n965_o2_p
  );


  buf

  (
    n786_o2_n_spl_,
    n786_o2_n
  );


  buf

  (
    g648_p_spl_,
    g648_p
  );


  buf

  (
    g648_p_spl_0,
    g648_p_spl_
  );


  buf

  (
    g648_n_spl_,
    g648_n
  );


  buf

  (
    g648_n_spl_0,
    g648_n_spl_
  );


  buf

  (
    n789_o2_p_spl_,
    n789_o2_p
  );


  buf

  (
    n789_o2_n_spl_,
    n789_o2_n
  );


  buf

  (
    g651_n_spl_,
    g651_n
  );


  buf

  (
    g651_p_spl_,
    g651_p
  );


  buf

  (
    n989_o2_n_spl_,
    n989_o2_n
  );


  buf

  (
    n989_o2_n_spl_0,
    n989_o2_n_spl_
  );


  buf

  (
    g653_n_spl_,
    g653_n
  );


  buf

  (
    g652_n_spl_,
    g652_n
  );


  buf

  (
    g652_n_spl_0,
    g652_n_spl_
  );


  buf

  (
    g653_p_spl_,
    g653_p
  );


  buf

  (
    g652_p_spl_,
    g652_p
  );


  buf

  (
    lo024_buf_o2_p_spl_,
    lo024_buf_o2_p
  );


  buf

  (
    lo024_buf_o2_p_spl_0,
    lo024_buf_o2_p_spl_
  );


  buf

  (
    lo024_buf_o2_p_spl_1,
    lo024_buf_o2_p_spl_
  );


  buf

  (
    lo092_buf_o2_n_spl_,
    lo092_buf_o2_n
  );


  buf

  (
    lo092_buf_o2_p_spl_,
    lo092_buf_o2_p
  );


  buf

  (
    lo092_buf_o2_p_spl_0,
    lo092_buf_o2_p_spl_
  );


  buf

  (
    lo088_buf_o2_p_spl_,
    lo088_buf_o2_p
  );


  buf

  (
    lo100_buf_o2_p_spl_,
    lo100_buf_o2_p
  );


  buf

  (
    lo096_buf_o2_p_spl_,
    lo096_buf_o2_p
  );


  buf

  (
    g599_n_spl_,
    g599_n
  );


  buf

  (
    g599_n_spl_0,
    g599_n_spl_
  );


  buf

  (
    n3089_o2_n_spl_,
    n3089_o2_n
  );


  buf

  (
    g597_p_spl_,
    g597_p
  );


  buf

  (
    g597_p_spl_0,
    g597_p_spl_
  );


  buf

  (
    n3091_o2_p_spl_,
    n3091_o2_p
  );


  buf

  (
    g598_p_spl_,
    g598_p
  );


  buf

  (
    g597_n_spl_,
    g597_n
  );


  buf

  (
    g597_n_spl_0,
    g597_n_spl_
  );


  buf

  (
    g597_n_spl_1,
    g597_n_spl_
  );


  buf

  (
    n3245_o2_n_spl_,
    n3245_o2_n
  );


  buf

  (
    g595_p_spl_,
    g595_p
  );


  buf

  (
    n3246_o2_p_spl_,
    n3246_o2_p
  );


  buf

  (
    n3246_o2_p_spl_0,
    n3246_o2_p_spl_
  );


  buf

  (
    n3246_o2_p_spl_00,
    n3246_o2_p_spl_0
  );


  buf

  (
    n3246_o2_p_spl_1,
    n3246_o2_p_spl_
  );


  buf

  (
    lo086_buf_o2_p_spl_,
    lo086_buf_o2_p
  );


  buf

  (
    lo086_buf_o2_p_spl_0,
    lo086_buf_o2_p_spl_
  );


  buf

  (
    n1950_lo_p_spl_,
    n1950_lo_p
  );


  buf

  (
    n1950_lo_p_spl_0,
    n1950_lo_p_spl_
  );


  buf

  (
    g592_n_spl_,
    g592_n
  );


  buf

  (
    g657_n_spl_,
    g657_n
  );


  buf

  (
    n762_o2_n_spl_,
    n762_o2_n
  );


  buf

  (
    g668_n_spl_,
    g668_n
  );


  buf

  (
    g668_n_spl_0,
    g668_n_spl_
  );


  buf

  (
    g668_n_spl_1,
    g668_n_spl_
  );


  buf

  (
    lo042_buf_o2_p_spl_,
    lo042_buf_o2_p
  );


  buf

  (
    lo042_buf_o2_p_spl_0,
    lo042_buf_o2_p_spl_
  );


  buf

  (
    lo042_buf_o2_p_spl_00,
    lo042_buf_o2_p_spl_0
  );


  buf

  (
    lo042_buf_o2_p_spl_1,
    lo042_buf_o2_p_spl_
  );


  buf

  (
    g668_p_spl_,
    g668_p
  );


  buf

  (
    g668_p_spl_0,
    g668_p_spl_
  );


  buf

  (
    g668_p_spl_1,
    g668_p_spl_
  );


  buf

  (
    lo042_buf_o2_n_spl_,
    lo042_buf_o2_n
  );


  buf

  (
    lo042_buf_o2_n_spl_0,
    lo042_buf_o2_n_spl_
  );


  buf

  (
    lo042_buf_o2_n_spl_1,
    lo042_buf_o2_n_spl_
  );


  buf

  (
    n760_o2_n_spl_,
    n760_o2_n
  );


  buf

  (
    n760_o2_n_spl_0,
    n760_o2_n_spl_
  );


  buf

  (
    n760_o2_n_spl_1,
    n760_o2_n_spl_
  );


  buf

  (
    n760_o2_p_spl_,
    n760_o2_p
  );


  buf

  (
    n760_o2_p_spl_0,
    n760_o2_p_spl_
  );


  buf

  (
    n760_o2_p_spl_00,
    n760_o2_p_spl_0
  );


  buf

  (
    n760_o2_p_spl_01,
    n760_o2_p_spl_0
  );


  buf

  (
    n760_o2_p_spl_1,
    n760_o2_p_spl_
  );


  buf

  (
    n760_o2_p_spl_10,
    n760_o2_p_spl_1
  );


  buf

  (
    lo034_buf_o2_n_spl_,
    lo034_buf_o2_n
  );


  buf

  (
    lo034_buf_o2_n_spl_0,
    lo034_buf_o2_n_spl_
  );


  buf

  (
    lo034_buf_o2_n_spl_1,
    lo034_buf_o2_n_spl_
  );


  buf

  (
    n754_o2_n_spl_,
    n754_o2_n
  );


  buf

  (
    n754_o2_n_spl_0,
    n754_o2_n_spl_
  );


  buf

  (
    n754_o2_n_spl_1,
    n754_o2_n_spl_
  );


  buf

  (
    n754_o2_p_spl_,
    n754_o2_p
  );


  buf

  (
    n754_o2_p_spl_0,
    n754_o2_p_spl_
  );


  buf

  (
    n751_o2_p_spl_,
    n751_o2_p
  );


  buf

  (
    n751_o2_p_spl_0,
    n751_o2_p_spl_
  );


  buf

  (
    n751_o2_p_spl_00,
    n751_o2_p_spl_0
  );


  buf

  (
    n751_o2_p_spl_000,
    n751_o2_p_spl_00
  );


  buf

  (
    n751_o2_p_spl_01,
    n751_o2_p_spl_0
  );


  buf

  (
    n751_o2_p_spl_1,
    n751_o2_p_spl_
  );


  buf

  (
    n751_o2_p_spl_10,
    n751_o2_p_spl_1
  );


  buf

  (
    n751_o2_p_spl_11,
    n751_o2_p_spl_1
  );


  buf

  (
    n751_o2_n_spl_,
    n751_o2_n
  );


  buf

  (
    n751_o2_n_spl_0,
    n751_o2_n_spl_
  );


  buf

  (
    n751_o2_n_spl_00,
    n751_o2_n_spl_0
  );


  buf

  (
    n751_o2_n_spl_1,
    n751_o2_n_spl_
  );


  buf

  (
    lo046_buf_o2_p_spl_,
    lo046_buf_o2_p
  );


  buf

  (
    lo046_buf_o2_p_spl_0,
    lo046_buf_o2_p_spl_
  );


  buf

  (
    lo046_buf_o2_p_spl_1,
    lo046_buf_o2_p_spl_
  );


  buf

  (
    lo046_buf_o2_n_spl_,
    lo046_buf_o2_n
  );


  buf

  (
    lo046_buf_o2_n_spl_0,
    lo046_buf_o2_n_spl_
  );


  buf

  (
    lo046_buf_o2_n_spl_1,
    lo046_buf_o2_n_spl_
  );


  buf

  (
    lo038_buf_o2_p_spl_,
    lo038_buf_o2_p
  );


  buf

  (
    lo038_buf_o2_p_spl_0,
    lo038_buf_o2_p_spl_
  );


  buf

  (
    lo038_buf_o2_p_spl_00,
    lo038_buf_o2_p_spl_0
  );


  buf

  (
    lo038_buf_o2_p_spl_1,
    lo038_buf_o2_p_spl_
  );


  buf

  (
    n755_o2_n_spl_,
    n755_o2_n
  );


  buf

  (
    n755_o2_n_spl_0,
    n755_o2_n_spl_
  );


  buf

  (
    n755_o2_n_spl_1,
    n755_o2_n_spl_
  );


  buf

  (
    lo038_buf_o2_n_spl_,
    lo038_buf_o2_n
  );


  buf

  (
    lo028_buf_o2_n_spl_,
    lo028_buf_o2_n
  );


  buf

  (
    lo028_buf_o2_n_spl_0,
    lo028_buf_o2_n_spl_
  );


  buf

  (
    lo028_buf_o2_n_spl_1,
    lo028_buf_o2_n_spl_
  );


  buf

  (
    g646_n_spl_,
    g646_n
  );


  buf

  (
    lo006_buf_o2_p_spl_,
    lo006_buf_o2_p
  );


  buf

  (
    lo002_buf_o2_p_spl_,
    lo002_buf_o2_p
  );


  buf

  (
    lo002_buf_o2_p_spl_0,
    lo002_buf_o2_p_spl_
  );


  buf

  (
    lo002_buf_o2_p_spl_1,
    lo002_buf_o2_p_spl_
  );


  buf

  (
    n771_o2_n_spl_,
    n771_o2_n
  );


  buf

  (
    n771_o2_n_spl_0,
    n771_o2_n_spl_
  );


  buf

  (
    n771_o2_n_spl_00,
    n771_o2_n_spl_0
  );


  buf

  (
    n771_o2_n_spl_01,
    n771_o2_n_spl_0
  );


  buf

  (
    n771_o2_n_spl_1,
    n771_o2_n_spl_
  );


  buf

  (
    n771_o2_n_spl_10,
    n771_o2_n_spl_1
  );


  buf

  (
    n771_o2_p_spl_,
    n771_o2_p
  );


  buf

  (
    n771_o2_p_spl_0,
    n771_o2_p_spl_
  );


  buf

  (
    n771_o2_p_spl_00,
    n771_o2_p_spl_0
  );


  buf

  (
    n771_o2_p_spl_01,
    n771_o2_p_spl_0
  );


  buf

  (
    n771_o2_p_spl_1,
    n771_o2_p_spl_
  );


  buf

  (
    n771_o2_p_spl_10,
    n771_o2_p_spl_1
  );


  buf

  (
    lo018_buf_o2_p_spl_,
    lo018_buf_o2_p
  );


  buf

  (
    lo022_buf_o2_p_spl_,
    lo022_buf_o2_p
  );


  buf

  (
    g690_p_spl_,
    g690_p
  );


  buf

  (
    g690_p_spl_0,
    g690_p_spl_
  );


  buf

  (
    g688_p_spl_,
    g688_p
  );


  buf

  (
    g688_p_spl_0,
    g688_p_spl_
  );


  buf

  (
    g690_n_spl_,
    g690_n
  );


  buf

  (
    g690_n_spl_0,
    g690_n_spl_
  );


  buf

  (
    g688_n_spl_,
    g688_n
  );


  buf

  (
    g688_n_spl_0,
    g688_n_spl_
  );


  buf

  (
    lo010_buf_o2_p_spl_,
    lo010_buf_o2_p
  );


  buf

  (
    lo010_buf_o2_p_spl_0,
    lo010_buf_o2_p_spl_
  );


  buf

  (
    lo010_buf_o2_p_spl_00,
    lo010_buf_o2_p_spl_0
  );


  buf

  (
    lo010_buf_o2_p_spl_1,
    lo010_buf_o2_p_spl_
  );


  buf

  (
    lo010_buf_o2_n_spl_,
    lo010_buf_o2_n
  );


  buf

  (
    g692_n_spl_,
    g692_n
  );


  buf

  (
    g692_p_spl_,
    g692_p
  );


  buf

  (
    g692_p_spl_0,
    g692_p_spl_
  );


  buf

  (
    g693_n_spl_,
    g693_n
  );


  buf

  (
    lo050_buf_o2_n_spl_,
    lo050_buf_o2_n
  );


  buf

  (
    lo050_buf_o2_n_spl_0,
    lo050_buf_o2_n_spl_
  );


  buf

  (
    lo050_buf_o2_p_spl_,
    lo050_buf_o2_p
  );


  buf

  (
    lo050_buf_o2_p_spl_0,
    lo050_buf_o2_p_spl_
  );


  buf

  (
    n753_o2_p_spl_,
    n753_o2_p
  );


  buf

  (
    n753_o2_p_spl_0,
    n753_o2_p_spl_
  );


  buf

  (
    lo054_buf_o2_p_spl_,
    lo054_buf_o2_p
  );


  buf

  (
    lo054_buf_o2_p_spl_0,
    lo054_buf_o2_p_spl_
  );


  buf

  (
    lo054_buf_o2_p_spl_1,
    lo054_buf_o2_p_spl_
  );


  buf

  (
    n753_o2_n_spl_,
    n753_o2_n
  );


  buf

  (
    lo054_buf_o2_n_spl_,
    lo054_buf_o2_n
  );


  buf

  (
    lo054_buf_o2_n_spl_0,
    lo054_buf_o2_n_spl_
  );


  buf

  (
    g705_n_spl_,
    g705_n
  );


  buf

  (
    g658_p_spl_,
    g658_p
  );


  buf

  (
    g658_p_spl_0,
    g658_p_spl_
  );


  buf

  (
    g658_p_spl_1,
    g658_p_spl_
  );


  buf

  (
    n774_o2_n_spl_,
    n774_o2_n
  );


  buf

  (
    n774_o2_n_spl_0,
    n774_o2_n_spl_
  );


  buf

  (
    n774_o2_p_spl_,
    n774_o2_p
  );


  buf

  (
    n774_o2_p_spl_0,
    n774_o2_p_spl_
  );


  buf

  (
    g708_n_spl_,
    g708_n
  );


  buf

  (
    g708_n_spl_0,
    g708_n_spl_
  );


  buf

  (
    g708_p_spl_,
    g708_p
  );


  buf

  (
    g708_p_spl_0,
    g708_p_spl_
  );


  buf

  (
    g711_n_spl_,
    g711_n
  );


  buf

  (
    n1081_o2_n_spl_,
    n1081_o2_n
  );


  buf

  (
    g661_n_spl_,
    g661_n
  );


  buf

  (
    n3087_o2_p_spl_,
    n3087_o2_p
  );


  buf

  (
    n3087_o2_p_spl_0,
    n3087_o2_p_spl_
  );


  buf

  (
    g717_n_spl_,
    g717_n
  );


  buf

  (
    g717_n_spl_0,
    g717_n_spl_
  );


  buf

  (
    g717_n_spl_1,
    g717_n_spl_
  );


  buf

  (
    n998_o2_n_spl_,
    n998_o2_n
  );


  buf

  (
    n3245_o2_p_spl_,
    n3245_o2_p
  );


  buf

  (
    n3245_o2_p_spl_0,
    n3245_o2_p_spl_
  );


  buf

  (
    n3245_o2_p_spl_1,
    n3245_o2_p_spl_
  );


  buf

  (
    g599_p_spl_,
    g599_p
  );


  buf

  (
    n998_o2_p_spl_,
    n998_o2_p
  );


  buf

  (
    n1221_o2_p_spl_,
    n1221_o2_p
  );


  buf

  (
    n1221_o2_n_spl_,
    n1221_o2_n
  );


  buf

  (
    g724_n_spl_,
    g724_n
  );


  buf

  (
    g722_n_spl_,
    g722_n
  );


  buf

  (
    g724_p_spl_,
    g724_p
  );


  buf

  (
    g722_p_spl_,
    g722_p
  );


  buf

  (
    g722_p_spl_0,
    g722_p_spl_
  );


  buf

  (
    n1214_o2_n_spl_,
    n1214_o2_n
  );


  buf

  (
    n3082_o2_n_spl_,
    n3082_o2_n
  );


  buf

  (
    n1214_o2_p_spl_,
    n1214_o2_p
  );


  buf

  (
    n3082_o2_p_spl_,
    n3082_o2_p
  );


  buf

  (
    g731_n_spl_,
    g731_n
  );


  buf

  (
    g553_n_spl_,
    g553_n
  );


  buf

  (
    g731_p_spl_,
    g731_p
  );


  buf

  (
    g553_p_spl_,
    g553_p
  );


  buf

  (
    g553_p_spl_0,
    g553_p_spl_
  );


  buf

  (
    g732_p_spl_,
    g732_p
  );


  buf

  (
    g730_p_spl_,
    g730_p
  );


  buf

  (
    g730_p_spl_0,
    g730_p_spl_
  );


  buf

  (
    g730_p_spl_1,
    g730_p_spl_
  );


  buf

  (
    g732_n_spl_,
    g732_n
  );


  buf

  (
    g730_n_spl_,
    g730_n
  );


  buf

  (
    g730_n_spl_0,
    g730_n_spl_
  );


  buf

  (
    g730_n_spl_00,
    g730_n_spl_0
  );


  buf

  (
    g730_n_spl_1,
    g730_n_spl_
  );


  buf

  (
    g735_p_spl_,
    g735_p
  );


  buf

  (
    g727_p_spl_,
    g727_p
  );


  buf

  (
    n1003_o2_p_spl_,
    n1003_o2_p
  );


  buf

  (
    n1003_o2_p_spl_0,
    n1003_o2_p_spl_
  );


  buf

  (
    n1003_o2_p_spl_1,
    n1003_o2_p_spl_
  );


  buf

  (
    g727_n_spl_,
    g727_n
  );


  buf

  (
    g727_n_spl_0,
    g727_n_spl_
  );


  buf

  (
    g735_n_spl_,
    g735_n
  );


  buf

  (
    n2619_o2_p_spl_,
    n2619_o2_p
  );


  buf

  (
    n2619_o2_p_spl_0,
    n2619_o2_p_spl_
  );


  buf

  (
    n2619_o2_p_spl_00,
    n2619_o2_p_spl_0
  );


  buf

  (
    n2619_o2_p_spl_01,
    n2619_o2_p_spl_0
  );


  buf

  (
    n2619_o2_p_spl_1,
    n2619_o2_p_spl_
  );


  buf

  (
    n2619_o2_p_spl_10,
    n2619_o2_p_spl_1
  );


  buf

  (
    n2624_o2_n_spl_,
    n2624_o2_n
  );


  buf

  (
    n2624_o2_n_spl_0,
    n2624_o2_n_spl_
  );


  buf

  (
    n2624_o2_n_spl_1,
    n2624_o2_n_spl_
  );


  buf

  (
    g559_n_spl_,
    g559_n
  );


  buf

  (
    g551_n_spl_,
    g551_n
  );


  buf

  (
    g552_n_spl_,
    g552_n
  );


  buf

  (
    g612_n_spl_,
    g612_n
  );


  buf

  (
    n1040_o2_p_spl_,
    n1040_o2_p
  );


  buf

  (
    n1040_o2_p_spl_0,
    n1040_o2_p_spl_
  );


  buf

  (
    n1040_o2_p_spl_00,
    n1040_o2_p_spl_0
  );


  buf

  (
    n1040_o2_p_spl_1,
    n1040_o2_p_spl_
  );


  buf

  (
    n1044_o2_n_spl_,
    n1044_o2_n
  );


  buf

  (
    n1044_o2_n_spl_0,
    n1044_o2_n_spl_
  );


  buf

  (
    n1044_o2_n_spl_1,
    n1044_o2_n_spl_
  );


  buf

  (
    n1034_o2_p_spl_,
    n1034_o2_p
  );


  buf

  (
    n1034_o2_p_spl_0,
    n1034_o2_p_spl_
  );


  buf

  (
    n1034_o2_p_spl_1,
    n1034_o2_p_spl_
  );


  buf

  (
    n1046_o2_p_spl_,
    n1046_o2_p
  );


  buf

  (
    n1046_o2_p_spl_0,
    n1046_o2_p_spl_
  );


  buf

  (
    n2676_o2_n_spl_,
    n2676_o2_n
  );


  buf

  (
    n1038_o2_p_spl_,
    n1038_o2_p
  );


  buf

  (
    n1038_o2_p_spl_0,
    n1038_o2_p_spl_
  );


  buf

  (
    n1038_o2_p_spl_1,
    n1038_o2_p_spl_
  );


  buf

  (
    n1031_o2_n_spl_,
    n1031_o2_n
  );


  buf

  (
    n1031_o2_n_spl_0,
    n1031_o2_n_spl_
  );


  buf

  (
    n2645_o2_n_spl_,
    n2645_o2_n
  );


  buf

  (
    g760_p_spl_,
    g760_p
  );


  buf

  (
    n2794_o2_p_spl_,
    n2794_o2_p
  );


  buf

  (
    n2794_o2_p_spl_0,
    n2794_o2_p_spl_
  );


  buf

  (
    n2622_o2_p_spl_,
    n2622_o2_p
  );


  buf

  (
    g771_n_spl_,
    g771_n
  );


  buf

  (
    g562_n_spl_,
    g562_n
  );


  buf

  (
    n2624_o2_p_spl_,
    n2624_o2_p
  );


  buf

  (
    n2621_o2_p_spl_,
    n2621_o2_p
  );


  buf

  (
    n2623_o2_p_spl_,
    n2623_o2_p
  );


  buf

  (
    n1031_o2_p_spl_,
    n1031_o2_p
  );


  buf

  (
    n1031_o2_p_spl_0,
    n1031_o2_p_spl_
  );


  buf

  (
    n1031_o2_p_spl_00,
    n1031_o2_p_spl_0
  );


  buf

  (
    n1031_o2_p_spl_1,
    n1031_o2_p_spl_
  );


  buf

  (
    n2623_o2_n_spl_,
    n2623_o2_n
  );


  buf

  (
    n1038_o2_n_spl_,
    n1038_o2_n
  );


  buf

  (
    n1038_o2_n_spl_0,
    n1038_o2_n_spl_
  );


  buf

  (
    n1038_o2_n_spl_00,
    n1038_o2_n_spl_0
  );


  buf

  (
    n1038_o2_n_spl_01,
    n1038_o2_n_spl_0
  );


  buf

  (
    n1038_o2_n_spl_1,
    n1038_o2_n_spl_
  );


  buf

  (
    n1038_o2_n_spl_10,
    n1038_o2_n_spl_1
  );


  buf

  (
    lo170_buf_o2_p_spl_,
    lo170_buf_o2_p
  );


  buf

  (
    n2627_o2_p_spl_,
    n2627_o2_p
  );


  buf

  (
    n2627_o2_p_spl_0,
    n2627_o2_p_spl_
  );


  buf

  (
    n2627_o2_p_spl_1,
    n2627_o2_p_spl_
  );


  buf

  (
    n1040_o2_n_spl_,
    n1040_o2_n
  );


  buf

  (
    n1040_o2_n_spl_0,
    n1040_o2_n_spl_
  );


  buf

  (
    n1040_o2_n_spl_00,
    n1040_o2_n_spl_0
  );


  buf

  (
    n1040_o2_n_spl_000,
    n1040_o2_n_spl_00
  );


  buf

  (
    n1040_o2_n_spl_01,
    n1040_o2_n_spl_0
  );


  buf

  (
    n1040_o2_n_spl_1,
    n1040_o2_n_spl_
  );


  buf

  (
    n1040_o2_n_spl_10,
    n1040_o2_n_spl_1
  );


  buf

  (
    n1040_o2_n_spl_11,
    n1040_o2_n_spl_1
  );


  buf

  (
    n2645_o2_p_spl_,
    n2645_o2_p
  );


  buf

  (
    n2645_o2_p_spl_0,
    n2645_o2_p_spl_
  );


  buf

  (
    n2622_o2_n_spl_,
    n2622_o2_n
  );


  buf

  (
    n1034_o2_n_spl_,
    n1034_o2_n
  );


  buf

  (
    n1034_o2_n_spl_0,
    n1034_o2_n_spl_
  );


  buf

  (
    n1034_o2_n_spl_00,
    n1034_o2_n_spl_0
  );


  buf

  (
    n1034_o2_n_spl_01,
    n1034_o2_n_spl_0
  );


  buf

  (
    n1034_o2_n_spl_1,
    n1034_o2_n_spl_
  );


  buf

  (
    n1046_o2_n_spl_,
    n1046_o2_n
  );


  buf

  (
    n1046_o2_n_spl_0,
    n1046_o2_n_spl_
  );


  buf

  (
    n1046_o2_n_spl_00,
    n1046_o2_n_spl_0
  );


  buf

  (
    n1046_o2_n_spl_01,
    n1046_o2_n_spl_0
  );


  buf

  (
    n1046_o2_n_spl_1,
    n1046_o2_n_spl_
  );


  buf

  (
    n1046_o2_n_spl_10,
    n1046_o2_n_spl_1
  );


  buf

  (
    n1044_o2_p_spl_,
    n1044_o2_p
  );


  buf

  (
    n1044_o2_p_spl_0,
    n1044_o2_p_spl_
  );


  buf

  (
    n1044_o2_p_spl_00,
    n1044_o2_p_spl_0
  );


  buf

  (
    n1044_o2_p_spl_01,
    n1044_o2_p_spl_0
  );


  buf

  (
    n1044_o2_p_spl_1,
    n1044_o2_p_spl_
  );


  buf

  (
    n1044_o2_p_spl_10,
    n1044_o2_p_spl_1
  );


  buf

  (
    n2676_o2_p_spl_,
    n2676_o2_p
  );


  buf

  (
    n2966_o2_p_spl_,
    n2966_o2_p
  );


  buf

  (
    n2966_o2_p_spl_0,
    n2966_o2_p_spl_
  );


  buf

  (
    g849_p_spl_,
    g849_p
  );


  buf

  (
    g848_n_spl_,
    g848_n
  );


  buf

  (
    n2967_o2_p_spl_,
    n2967_o2_p
  );


  buf

  (
    n2967_o2_p_spl_0,
    n2967_o2_p_spl_
  );


  buf

  (
    n1298_o2_n_spl_,
    n1298_o2_n
  );


  buf

  (
    n2793_o2_n_spl_,
    n2793_o2_n
  );


  buf

  (
    n3214_o2_p_spl_,
    n3214_o2_p
  );


  buf

  (
    n3214_o2_n_spl_,
    n3214_o2_n
  );


  buf

  (
    g870_n_spl_,
    g870_n
  );


  buf

  (
    n3081_o2_n_spl_,
    n3081_o2_n
  );


  buf

  (
    g870_p_spl_,
    g870_p
  );


  buf

  (
    n3081_o2_p_spl_,
    n3081_o2_p
  );


  buf

  (
    g873_n_spl_,
    g873_n
  );


  buf

  (
    g873_n_spl_0,
    g873_n_spl_
  );


  buf

  (
    g687_n_spl_,
    g687_n
  );


  buf

  (
    g878_n_spl_,
    g878_n
  );


  buf

  (
    g877_p_spl_,
    g877_p
  );


  buf

  (
    g877_p_spl_0,
    g877_p_spl_
  );


  buf

  (
    g883_n_spl_,
    g883_n
  );


  buf

  (
    g883_n_spl_0,
    g883_n_spl_
  );


  buf

  (
    g883_n_spl_1,
    g883_n_spl_
  );


  buf

  (
    g884_n_spl_,
    g884_n
  );


  buf

  (
    g885_n_spl_,
    g885_n
  );


  buf

  (
    n1003_o2_n_spl_,
    n1003_o2_n
  );


  buf

  (
    n1003_o2_n_spl_0,
    n1003_o2_n_spl_
  );


  buf

  (
    g888_n_spl_,
    g888_n
  );


  buf

  (
    g656_n_spl_,
    g656_n
  );


  buf

  (
    g577_n_spl_,
    g577_n
  );


  buf

  (
    g577_n_spl_0,
    g577_n_spl_
  );


  buf

  (
    lo174_buf_o2_p_spl_,
    lo174_buf_o2_p
  );


  buf

  (
    lo030_buf_o2_p_spl_,
    lo030_buf_o2_p
  );


  buf

  (
    lo030_buf_o2_p_spl_0,
    lo030_buf_o2_p_spl_
  );


  buf

  (
    n3090_o2_p_spl_,
    n3090_o2_p
  );


  buf

  (
    g960_p_spl_,
    g960_p
  );


  buf

  (
    g960_n_spl_,
    g960_n
  );


  buf

  (
    g873_p_spl_,
    g873_p
  );


  buf

  (
    g645_n_spl_,
    g645_n
  );


  buf

  (
    g645_n_spl_0,
    g645_n_spl_
  );


  buf

  (
    g621_n_spl_,
    g621_n
  );


  buf

  (
    g621_n_spl_0,
    g621_n_spl_
  );


  buf

  (
    lo154_buf_o2_p_spl_,
    lo154_buf_o2_p
  );


  buf

  (
    lo142_buf_o2_p_spl_,
    lo142_buf_o2_p
  );


  buf

  (
    g990_n_spl_,
    g990_n
  );


  buf

  (
    g705_p_spl_,
    g705_p
  );


  buf

  (
    g659_n_spl_,
    g659_n
  );


  buf

  (
    g659_n_spl_0,
    g659_n_spl_
  );


  buf

  (
    g659_n_spl_00,
    g659_n_spl_0
  );


  buf

  (
    g659_n_spl_01,
    g659_n_spl_0
  );


  buf

  (
    g659_n_spl_1,
    g659_n_spl_
  );


  buf

  (
    g659_n_spl_10,
    g659_n_spl_1
  );


  buf

  (
    g676_n_spl_,
    g676_n
  );


  buf

  (
    g707_n_spl_,
    g707_n
  );


  buf

  (
    g711_p_spl_,
    g711_p
  );


  buf

  (
    g684_n_spl_,
    g684_n
  );


  buf

  (
    g713_n_spl_,
    g713_n
  );


  buf

  (
    n3086_o2_p_spl_,
    n3086_o2_p
  );


  buf

  (
    lo026_buf_o2_p_spl_,
    lo026_buf_o2_p
  );


  buf

  (
    n3089_o2_p_spl_,
    n3089_o2_p
  );


  buf

  (
    n3092_o2_p_spl_,
    n3092_o2_p
  );


  buf

  (
    g581_n_spl_,
    g581_n
  );


  buf

  (
    g581_n_spl_0,
    g581_n_spl_
  );


  buf

  (
    g581_n_spl_00,
    g581_n_spl_0
  );


  buf

  (
    g581_n_spl_01,
    g581_n_spl_0
  );


  buf

  (
    g581_n_spl_1,
    g581_n_spl_
  );


  buf

  (
    n3092_o2_n_spl_,
    n3092_o2_n
  );


  buf

  (
    n3213_o2_p_spl_,
    n3213_o2_p
  );


  buf

  (
    g583_n_spl_,
    g583_n
  );


  buf

  (
    g583_n_spl_0,
    g583_n_spl_
  );


  buf

  (
    g583_n_spl_00,
    g583_n_spl_0
  );


  buf

  (
    g583_n_spl_01,
    g583_n_spl_0
  );


  buf

  (
    g583_n_spl_1,
    g583_n_spl_
  );


  buf

  (
    n1938_lo_p_spl_,
    n1938_lo_p
  );


  buf

  (
    n1938_lo_p_spl_0,
    n1938_lo_p_spl_
  );


  buf

  (
    g1013_p_spl_,
    g1013_p
  );


  buf

  (
    g1013_p_spl_0,
    g1013_p_spl_
  );


  buf

  (
    g890_n_spl_,
    g890_n
  );


  buf

  (
    g886_n_spl_,
    g886_n
  );


  buf

  (
    g886_n_spl_0,
    g886_n_spl_
  );


  buf

  (
    n1926_lo_p_spl_,
    n1926_lo_p
  );


  buf

  (
    g976_n_spl_,
    g976_n
  );


  buf

  (
    n2298_lo_n_spl_,
    n2298_lo_n
  );


  buf

  (
    n2250_lo_p_spl_,
    n2250_lo_p
  );


  buf

  (
    n2238_lo_p_spl_,
    n2238_lo_p
  );


  buf

  (
    g1020_n_spl_,
    g1020_n
  );


  buf

  (
    g590_p_spl_,
    g590_p
  );


  buf

  (
    n2298_lo_p_spl_,
    n2298_lo_p
  );


  buf

  (
    g577_p_spl_,
    g577_p
  );


  buf

  (
    g577_p_spl_0,
    g577_p_spl_
  );


  buf

  (
    g1026_p_spl_,
    g1026_p
  );


  buf

  (
    g656_p_spl_,
    g656_p
  );


  buf

  (
    g656_p_spl_0,
    g656_p_spl_
  );


  buf

  (
    g1031_n_spl_,
    g1031_n
  );


  buf

  (
    g1025_n_spl_,
    g1025_n
  );


  buf

  (
    g1025_n_spl_0,
    g1025_n_spl_
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G1_p_spl_0,
    G1_p_spl_
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    g664_n_spl_,
    g664_n
  );


  buf

  (
    g662_n_spl_,
    g662_n
  );


  buf

  (
    g716_p_spl_,
    g716_p
  );


  buf

  (
    lo082_buf_o2_p_spl_,
    lo082_buf_o2_p
  );


  buf

  (
    lo082_buf_o2_p_spl_0,
    lo082_buf_o2_p_spl_
  );


  buf

  (
    g591_n_spl_,
    g591_n
  );


  buf

  (
    n1974_lo_p_spl_,
    n1974_lo_p
  );


  buf

  (
    n1974_lo_p_spl_0,
    n1974_lo_p_spl_
  );


  buf

  (
    g598_n_spl_,
    g598_n
  );


  buf

  (
    g598_n_spl_0,
    g598_n_spl_
  );


  buf

  (
    g598_n_spl_1,
    g598_n_spl_
  );


  buf

  (
    n3170_o2_p_spl_,
    n3170_o2_p
  );


  buf

  (
    g719_n_spl_,
    g719_n
  );


  buf

  (
    n3095_o2_p_spl_,
    n3095_o2_p
  );


  buf

  (
    n3095_o2_p_spl_0,
    n3095_o2_p_spl_
  );


  buf

  (
    g950_n_spl_,
    g950_n
  );


  buf

  (
    g720_n_spl_,
    g720_n
  );


  buf

  (
    g595_n_spl_,
    g595_n
  );


  buf

  (
    g595_n_spl_0,
    g595_n_spl_
  );


  buf

  (
    g972_n_spl_,
    g972_n
  );


  buf

  (
    g875_n_spl_,
    g875_n
  );


  buf

  (
    g876_n_spl_,
    g876_n
  );


  buf

  (
    n752_o2_p_spl_,
    n752_o2_p
  );


  buf

  (
    n752_o2_p_spl_0,
    n752_o2_p_spl_
  );


  buf

  (
    g1082_p_spl_,
    g1082_p
  );


  buf

  (
    g1082_p_spl_0,
    g1082_p_spl_
  );


  buf

  (
    g1082_p_spl_1,
    g1082_p_spl_
  );


  buf

  (
    g666_p_spl_,
    g666_p
  );


  buf

  (
    g1088_p_spl_,
    g1088_p
  );


  buf

  (
    g1086_n_spl_,
    g1086_n
  );


  buf

  (
    g665_n_spl_,
    g665_n
  );


  buf

  (
    lo145_buf_o2_p_spl_,
    lo145_buf_o2_p
  );


  buf

  (
    n780_o2_n_spl_,
    n780_o2_n
  );


  buf

  (
    n780_o2_n_spl_0,
    n780_o2_n_spl_
  );


  buf

  (
    lo138_buf_o2_p_spl_,
    lo138_buf_o2_p
  );


  buf

  (
    n780_o2_p_spl_,
    n780_o2_p
  );


  buf

  (
    n780_o2_p_spl_0,
    n780_o2_p_spl_
  );


  buf

  (
    g1108_n_spl_,
    g1108_n
  );


  buf

  (
    g663_p_spl_,
    g663_p
  );


  buf

  (
    g660_p_spl_,
    g660_p
  );


  buf

  (
    g990_p_spl_,
    g990_p
  );


  buf

  (
    g701_n_spl_,
    g701_n
  );


  buf

  (
    g992_n_spl_,
    g992_n
  );


  buf

  (
    g998_p_spl_,
    g998_p
  );


  buf

  (
    g995_p_spl_,
    g995_p
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_00,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_000,
    G4_p_spl_00
  );


  buf

  (
    G4_p_spl_001,
    G4_p_spl_00
  );


  buf

  (
    G4_p_spl_01,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_10,
    G4_p_spl_1
  );


  buf

  (
    G4_p_spl_11,
    G4_p_spl_1
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G12_p_spl_0,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_1,
    G12_p_spl_
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    G13_p_spl_,
    G13_p
  );


  buf

  (
    G13_p_spl_0,
    G13_p_spl_
  );


  buf

  (
    n1983_lo_p_spl_,
    n1983_lo_p
  );


  buf

  (
    g667_n_spl_,
    g667_n
  );


  buf

  (
    n1995_lo_p_spl_,
    n1995_lo_p
  );


  buf

  (
    g686_p_spl_,
    g686_p
  );


  buf

  (
    lo117_buf_o2_p_spl_,
    lo117_buf_o2_p
  );


  buf

  (
    lo117_buf_o2_p_spl_0,
    lo117_buf_o2_p_spl_
  );


  buf

  (
    lo014_buf_o2_p_spl_,
    lo014_buf_o2_p
  );


  buf

  (
    lo014_buf_o2_p_spl_0,
    lo014_buf_o2_p_spl_
  );


  buf

  (
    lo014_buf_o2_p_spl_00,
    lo014_buf_o2_p_spl_0
  );


  buf

  (
    lo014_buf_o2_p_spl_1,
    lo014_buf_o2_p_spl_
  );


  buf

  (
    lo014_buf_o2_n_spl_,
    lo014_buf_o2_n
  );


  buf

  (
    lo014_buf_o2_n_spl_0,
    lo014_buf_o2_n_spl_
  );


  buf

  (
    lo014_buf_o2_n_spl_1,
    lo014_buf_o2_n_spl_
  );


  buf

  (
    n2079_lo_p_spl_,
    n2079_lo_p
  );


  buf

  (
    g1108_p_spl_,
    g1108_p
  );


  buf

  (
    lo122_buf_o2_p_spl_,
    lo122_buf_o2_p
  );


  buf

  (
    g691_p_spl_,
    g691_p
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    G4_n_spl_0,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_00,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_1,
    G4_n_spl_
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G3_p_spl_0,
    G3_p_spl_
  );


  buf

  (
    G3_p_spl_00,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_1,
    G3_p_spl_
  );


  buf

  (
    g1034_n_spl_,
    g1034_n
  );


  buf

  (
    G3_n_spl_,
    G3_n
  );


  buf

  (
    G5_p_spl_,
    G5_p
  );


  buf

  (
    G5_p_spl_0,
    G5_p_spl_
  );


  buf

  (
    lo126_buf_o2_n_spl_,
    lo126_buf_o2_n
  );


  buf

  (
    lo122_buf_o2_n_spl_,
    lo122_buf_o2_n
  );


  buf

  (
    g691_n_spl_,
    g691_n
  );


  buf

  (
    g1179_p_spl_,
    g1179_p
  );


  buf

  (
    g658_n_spl_,
    g658_n
  );


  buf

  (
    g658_n_spl_0,
    g658_n_spl_
  );


  buf

  (
    g1085_n_spl_,
    g1085_n
  );


  buf

  (
    g1085_n_spl_0,
    g1085_n_spl_
  );


  buf

  (
    g1190_p_spl_,
    g1190_p
  );


  buf

  (
    g1098_n_spl_,
    g1098_n
  );


  buf

  (
    g1098_n_spl_0,
    g1098_n_spl_
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G1_n_spl_0,
    G1_n_spl_
  );


  buf

  (
    g1197_n_spl_,
    g1197_n
  );


  buf

  (
    g1035_n_spl_,
    g1035_n
  );


  buf

  (
    g1035_n_spl_0,
    g1035_n_spl_
  );


  buf

  (
    g1074_n_spl_,
    g1074_n
  );


  buf

  (
    g985_n_spl_,
    g985_n
  );


  buf

  (
    g1110_n_spl_,
    g1110_n
  );


  buf

  (
    g1121_p_spl_,
    g1121_p
  );


  buf

  (
    g1120_p_spl_,
    g1120_p
  );


  buf

  (
    G13_n_spl_,
    G13_n
  );


  buf

  (
    g1124_n_spl_,
    g1124_n
  );


  buf

  (
    g1123_n_spl_,
    g1123_n
  );


  buf

  (
    g1208_p_spl_,
    g1208_p
  );


  buf

  (
    G41_p_spl_,
    G41_p
  );


  buf

  (
    g1162_n_spl_,
    g1162_n
  );


  buf

  (
    g1162_n_spl_0,
    g1162_n_spl_
  );


  buf

  (
    g1162_n_spl_1,
    g1162_n_spl_
  );


  buf

  (
    g1122_n_spl_,
    g1122_n
  );


  buf

  (
    g1122_n_spl_0,
    g1122_n_spl_
  );


  buf

  (
    g1122_n_spl_1,
    g1122_n_spl_
  );


  buf

  (
    G34_n_spl_,
    G34_n
  );


  buf

  (
    g1164_p_spl_,
    g1164_p
  );


  buf

  (
    g1201_n_spl_,
    g1201_n
  );


  buf

  (
    G35_p_spl_,
    G35_p
  );


  buf

  (
    G35_p_spl_0,
    G35_p_spl_
  );


  buf

  (
    g1200_p_spl_,
    g1200_p
  );


  buf

  (
    g1163_n_spl_,
    g1163_n
  );


  buf

  (
    G40_p_spl_,
    G40_p
  );


  buf

  (
    G33_p_spl_,
    G33_p
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G34_p_spl_,
    G34_p
  );


  buf

  (
    g1210_n_spl_,
    g1210_n
  );


endmodule
