// Benchmark "mymod" written by ABC on Sun Oct 29 19:31:51 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41,
    G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
    G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
    G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
    G1354, G1355  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
    G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
    G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
    G1354, G1355;
  reg n630_lo, n642_lo, n654_lo, n666_lo, n678_lo, n690_lo, n702_lo,
    n714_lo, n726_lo, n738_lo, n750_lo, n762_lo, n774_lo, n786_lo, n798_lo,
    n810_lo, n822_lo, n834_lo, n846_lo, n858_lo, n870_lo, n882_lo, n894_lo,
    n906_lo, n918_lo, n930_lo, n942_lo, n954_lo, n966_lo, n978_lo, n990_lo,
    n1002_lo, n1005_lo, n1008_lo, n1017_lo, n1020_lo, n1029_lo, n1032_lo,
    n1041_lo, n1044_lo, n1053_lo, n1056_lo, n1065_lo, n1068_lo, n1077_lo,
    n1080_lo, n1089_lo, n1092_lo, n1101_lo, n1104_lo, n1837_o2, n1838_o2,
    n1839_o2, n1840_o2, n1841_o2, n1842_o2, n1843_o2, n1844_o2, n1845_o2,
    n1846_o2, n1847_o2, n1848_o2, n1849_o2, n1850_o2, n1851_o2, n1852_o2,
    n1853_o2, n1854_o2, n1855_o2, n1856_o2, n1857_o2, n1858_o2, n1859_o2,
    n1860_o2, n1861_o2, n1862_o2, n1863_o2, n1864_o2, n1865_o2, n1866_o2,
    n1867_o2, n1868_o2, G834_o2, G847_o2, G860_o2, G873_o2, G925_o2,
    G886_o2, G912_o2, G899_o2, n2151_o2, n2152_o2, n2153_o2, n2154_o2,
    n2155_o2, n2156_o2, n2157_o2, n2158_o2, n2159_o2, n2160_o2, n2161_o2,
    n2162_o2, n2163_o2, n2164_o2, n2165_o2, n2166_o2, n2167_o2, n2168_o2,
    n2169_o2, n2170_o2, n2171_o2, n2172_o2, n2173_o2, n2174_o2, n2175_o2,
    n2176_o2, n2177_o2, n2178_o2, n2179_o2, n2180_o2, n2181_o2, n2182_o2,
    G974_o2, G976_o2, G970_o2, G972_o2, G973_o2, G977_o2, G971_o2, G975_o2,
    G954_o2, G956_o2, G950_o2, G952_o2, G953_o2, G957_o2, G951_o2, G955_o2,
    G986_o2, G991_o2, G770_o2, G773_o2, G776_o2, G779_o2, G782_o2, G785_o2,
    G788_o2, G791_o2, G642_o2, G645_o2, G648_o2, G651_o2, G654_o2, G657_o2,
    G660_o2, G663_o2, G602_o2, G607_o2, G612_o2, G617_o2, G622_o2, G627_o2,
    G632_o2, G637_o2, n627_lo_buf_o2, n639_lo_buf_o2, n651_lo_buf_o2,
    n663_lo_buf_o2, n675_lo_buf_o2, n687_lo_buf_o2, n699_lo_buf_o2,
    n711_lo_buf_o2, n723_lo_buf_o2, n735_lo_buf_o2, n747_lo_buf_o2,
    n759_lo_buf_o2, n771_lo_buf_o2, n783_lo_buf_o2, n795_lo_buf_o2,
    n807_lo_buf_o2, n819_lo_buf_o2, n831_lo_buf_o2, n843_lo_buf_o2,
    n855_lo_buf_o2, n867_lo_buf_o2, n879_lo_buf_o2, n891_lo_buf_o2,
    n903_lo_buf_o2, n915_lo_buf_o2, n927_lo_buf_o2, n939_lo_buf_o2,
    n951_lo_buf_o2, n963_lo_buf_o2, n975_lo_buf_o2, n987_lo_buf_o2,
    n999_lo_buf_o2;
  wire new_new_n467__, new_new_n469__, new_new_n471__, new_new_n473__,
    new_new_n475__, new_new_n477__, new_new_n479__, new_new_n481__,
    new_new_n483__, new_new_n485__, new_new_n487__, new_new_n489__,
    new_new_n491__, new_new_n493__, new_new_n495__, new_new_n497__,
    new_new_n499__, new_new_n501__, new_new_n503__, new_new_n505__,
    new_new_n507__, new_new_n509__, new_new_n511__, new_new_n513__,
    new_new_n515__, new_new_n517__, new_new_n519__, new_new_n521__,
    new_new_n523__, new_new_n525__, new_new_n527__, new_new_n529__,
    new_new_n531__, new_new_n533__, new_new_n535__, new_new_n537__,
    new_new_n539__, new_new_n541__, new_new_n543__, new_new_n545__,
    new_new_n547__, new_new_n548__, new_new_n549__, new_new_n550__,
    new_new_n551__, new_new_n552__, new_new_n553__, new_new_n554__,
    new_new_n555__, new_new_n556__, new_new_n557__, new_new_n558__,
    new_new_n559__, new_new_n560__, new_new_n561__, new_new_n562__,
    new_new_n563__, new_new_n564__, new_new_n565__, new_new_n566__,
    new_new_n567__, new_new_n568__, new_new_n569__, new_new_n570__,
    new_new_n571__, new_new_n572__, new_new_n573__, new_new_n574__,
    new_new_n575__, new_new_n576__, new_new_n577__, new_new_n578__,
    new_new_n579__, new_new_n580__, new_new_n581__, new_new_n582__,
    new_new_n583__, new_new_n584__, new_new_n585__, new_new_n586__,
    new_new_n587__, new_new_n588__, new_new_n589__, new_new_n590__,
    new_new_n591__, new_new_n592__, new_new_n593__, new_new_n594__,
    new_new_n595__, new_new_n596__, new_new_n597__, new_new_n598__,
    new_new_n599__, new_new_n600__, new_new_n601__, new_new_n602__,
    new_new_n603__, new_new_n604__, new_new_n605__, new_new_n606__,
    new_new_n607__, new_new_n608__, new_new_n609__, new_new_n610__,
    new_new_n611__, new_new_n613__, new_new_n614__, new_new_n615__,
    new_new_n617__, new_new_n618__, new_new_n619__, new_new_n621__,
    new_new_n622__, new_new_n623__, new_new_n625__, new_new_n626__,
    new_new_n627__, new_new_n629__, new_new_n630__, new_new_n631__,
    new_new_n633__, new_new_n634__, new_new_n635__, new_new_n637__,
    new_new_n638__, new_new_n639__, new_new_n641__, new_new_n642__,
    new_new_n643__, new_new_n645__, new_new_n646__, new_new_n647__,
    new_new_n649__, new_new_n651__, new_new_n653__, new_new_n655__,
    new_new_n657__, new_new_n659__, new_new_n661__, new_new_n663__,
    new_new_n665__, new_new_n667__, new_new_n669__, new_new_n671__,
    new_new_n673__, new_new_n675__, new_new_n677__, new_new_n679__,
    new_new_n681__, new_new_n683__, new_new_n685__, new_new_n687__,
    new_new_n689__, new_new_n691__, new_new_n693__, new_new_n695__,
    new_new_n697__, new_new_n699__, new_new_n701__, new_new_n703__,
    new_new_n705__, new_new_n707__, new_new_n709__, new_new_n711__,
    new_new_n712__, new_new_n713__, new_new_n714__, new_new_n715__,
    new_new_n716__, new_new_n717__, new_new_n718__, new_new_n719__,
    new_new_n720__, new_new_n721__, new_new_n722__, new_new_n723__,
    new_new_n724__, new_new_n725__, new_new_n726__, new_new_n727__,
    new_new_n728__, new_new_n729__, new_new_n730__, new_new_n731__,
    new_new_n732__, new_new_n733__, new_new_n734__, new_new_n735__,
    new_new_n736__, new_new_n737__, new_new_n738__, new_new_n739__,
    new_new_n740__, new_new_n741__, new_new_n742__, new_new_n743__,
    new_new_n744__, new_new_n745__, new_new_n746__, new_new_n747__,
    new_new_n748__, new_new_n749__, new_new_n750__, new_new_n751__,
    new_new_n752__, new_new_n753__, new_new_n754__, new_new_n755__,
    new_new_n756__, new_new_n757__, new_new_n758__, new_new_n759__,
    new_new_n760__, new_new_n761__, new_new_n762__, new_new_n763__,
    new_new_n764__, new_new_n765__, new_new_n766__, new_new_n767__,
    new_new_n768__, new_new_n769__, new_new_n770__, new_new_n771__,
    new_new_n772__, new_new_n773__, new_new_n774__, new_new_n775__,
    new_new_n776__, new_new_n777__, new_new_n778__, new_new_n779__,
    new_new_n780__, new_new_n781__, new_new_n782__, new_new_n783__,
    new_new_n784__, new_new_n785__, new_new_n786__, new_new_n787__,
    new_new_n788__, new_new_n789__, new_new_n790__, new_new_n791__,
    new_new_n792__, new_new_n793__, new_new_n794__, new_new_n795__,
    new_new_n796__, new_new_n797__, new_new_n798__, new_new_n799__,
    new_new_n800__, new_new_n801__, new_new_n802__, new_new_n803__,
    new_new_n804__, new_new_n805__, new_new_n806__, new_new_n807__,
    new_new_n808__, new_new_n809__, new_new_n810__, new_new_n811__,
    new_new_n812__, new_new_n813__, new_new_n814__, new_new_n815__,
    new_new_n816__, new_new_n817__, new_new_n818__, new_new_n819__,
    new_new_n820__, new_new_n821__, new_new_n822__, new_new_n823__,
    new_new_n824__, new_new_n825__, new_new_n826__, new_new_n827__,
    new_new_n828__, new_new_n829__, new_new_n830__, new_new_n831__,
    new_new_n832__, new_new_n833__, new_new_n834__, new_new_n835__,
    new_new_n836__, new_new_n837__, new_new_n838__, new_new_n839__,
    new_new_n840__, new_new_n841__, new_new_n842__, new_new_n843__,
    new_new_n844__, new_new_n845__, new_new_n846__, new_new_n847__,
    new_new_n848__, new_new_n849__, new_new_n850__, new_new_n851__,
    new_new_n852__, new_new_n853__, new_new_n854__, new_new_n855__,
    new_new_n856__, new_new_n857__, new_new_n858__, new_new_n859__,
    new_new_n860__, new_new_n861__, new_new_n862__, new_new_n863__,
    new_new_n864__, new_new_n865__, new_new_n866__, new_new_n867__,
    new_new_n868__, new_new_n869__, new_new_n870__, new_new_n871__,
    new_new_n872__, new_new_n873__, new_new_n874__, new_new_n875__,
    new_new_n876__, new_new_n877__, new_new_n878__, new_new_n879__,
    new_new_n880__, new_new_n881__, new_new_n882__, new_new_n883__,
    new_new_n884__, new_new_n885__, new_new_n886__, new_new_n887__,
    new_new_n888__, new_new_n889__, new_new_n890__, new_new_n891__,
    new_new_n892__, new_new_n893__, new_new_n894__, new_new_n895__,
    new_new_n896__, new_new_n897__, new_new_n898__, new_new_n899__,
    new_new_n900__, new_new_n901__, new_new_n902__, new_new_n903__,
    new_new_n904__, new_new_n905__, new_new_n906__, new_new_n907__,
    new_new_n908__, new_new_n909__, new_new_n910__, new_new_n911__,
    new_new_n912__, new_new_n913__, new_new_n914__, new_new_n915__,
    new_new_n916__, new_new_n917__, new_new_n918__, new_new_n919__,
    new_new_n920__, new_new_n921__, new_new_n922__, new_new_n923__,
    new_new_n924__, new_new_n925__, new_new_n926__, new_new_n927__,
    new_new_n928__, new_new_n929__, new_new_n930__, new_new_n931__,
    new_new_n932__, new_new_n933__, new_new_n934__, new_new_n935__,
    new_new_n936__, new_new_n937__, new_new_n938__, new_new_n939__,
    new_new_n940__, new_new_n941__, new_new_n942__, new_new_n943__,
    new_new_n944__, new_new_n945__, new_new_n946__, new_new_n947__,
    new_new_n948__, new_new_n949__, new_new_n950__, new_new_n951__,
    new_new_n952__, new_new_n953__, new_new_n954__, new_new_n955__,
    new_new_n956__, new_new_n957__, new_new_n958__, new_new_n959__,
    new_new_n960__, new_new_n961__, new_new_n962__, new_new_n963__,
    new_new_n964__, new_new_n965__, new_new_n966__, new_new_n967__,
    new_new_n968__, new_new_n969__, new_new_n970__, new_new_n971__,
    new_new_n972__, new_new_n973__, new_new_n974__, new_new_n975__,
    new_new_n976__, new_new_n977__, new_new_n978__, new_new_n979__,
    new_new_n980__, new_new_n981__, new_new_n982__, new_new_n983__,
    new_new_n984__, new_new_n985__, new_new_n986__, new_new_n987__,
    new_new_n988__, new_new_n989__, new_new_n990__, new_new_n991__,
    new_new_n992__, new_new_n993__, new_new_n994__, new_new_n995__,
    new_new_n996__, new_new_n997__, new_new_n998__, new_new_n999__,
    new_new_n1000__, new_new_n1001__, new_new_n1002__, new_new_n1003__,
    new_new_n1004__, new_new_n1005__, new_new_n1006__, new_new_n1007__,
    new_new_n1008__, new_new_n1009__, new_new_n1010__, new_new_n1011__,
    new_new_n1012__, new_new_n1013__, new_new_n1014__, new_new_n1015__,
    new_new_n1016__, new_new_n1017__, new_new_n1018__, new_new_n1019__,
    new_new_n1020__, new_new_n1021__, new_new_n1022__, new_new_n1023__,
    new_new_n1024__, new_new_n1025__, new_new_n1026__, new_new_n1027__,
    new_new_n1028__, new_new_n1029__, new_new_n1030__, new_new_n1031__,
    new_new_n1032__, new_new_n1033__, new_new_n1034__, new_new_n1035__,
    new_new_n1036__, new_new_n1037__, new_new_n1038__, new_new_n1039__,
    new_new_n1040__, new_new_n1041__, new_new_n1042__, new_new_n1043__,
    new_new_n1044__, new_new_n1045__, new_new_n1046__, new_new_n1047__,
    new_new_n1048__, new_new_n1049__, new_new_n1050__, new_new_n1051__,
    new_new_n1052__, new_new_n1053__, new_new_n1054__, new_new_n1055__,
    new_new_n1056__, new_new_n1057__, new_new_n1058__, new_new_n1059__,
    new_new_n1060__, new_new_n1061__, new_new_n1062__, new_new_n1063__,
    new_new_n1064__, new_new_n1065__, new_new_n1066__, new_new_n1067__,
    new_new_n1068__, new_new_n1069__, new_new_n1070__, new_new_n1071__,
    new_new_n1072__, new_new_n1073__, new_new_n1074__, new_new_n1075__,
    new_new_n1076__, new_new_n1077__, new_new_n1078__, new_new_n1079__,
    new_new_n1080__, new_new_n1081__, new_new_n1082__, new_new_n1083__,
    new_new_n1084__, new_new_n1085__, new_new_n1086__, new_new_n1087__,
    new_new_n1088__, new_new_n1089__, new_new_n1090__, new_new_n1091__,
    new_new_n1092__, new_new_n1093__, new_new_n1094__, new_new_n1095__,
    new_new_n1096__, new_new_n1097__, new_new_n1098__, new_new_n1099__,
    new_new_n1100__, new_new_n1101__, new_new_n1102__, new_new_n1103__,
    new_new_n1104__, new_new_n1105__, new_new_n1106__, new_new_n1107__,
    new_new_n1108__, new_new_n1109__, new_new_n1110__, new_new_n1111__,
    new_new_n1112__, new_new_n1113__, new_new_n1114__, new_new_n1115__,
    new_new_n1116__, new_new_n1117__, new_new_n1118__, new_new_n1119__,
    new_new_n1120__, new_new_n1121__, new_new_n1122__, new_new_n1123__,
    new_new_n1124__, new_new_n1125__, new_new_n1126__, new_new_n1127__,
    new_new_n1128__, new_new_n1129__, new_new_n1130__, new_new_n1131__,
    new_new_n1132__, new_new_n1133__, new_new_n1134__, new_new_n1135__,
    new_new_n1136__, new_new_n1137__, new_new_n1138__, new_new_n1139__,
    new_new_n1140__, new_new_n1141__, new_new_n1142__, new_new_n1143__,
    new_new_n1144__, new_new_n1145__, new_new_n1146__, new_new_n1147__,
    new_new_n1148__, new_new_n1149__, new_new_n1150__, new_new_n1151__,
    new_new_n1152__, new_new_n1153__, new_new_n1154__, new_new_n1155__,
    new_new_n1156__, new_new_n1157__, new_new_n1158__, new_new_n1159__,
    new_new_n1160__, new_new_n1161__, new_new_n1162__, new_new_n1163__,
    new_new_n1164__, new_new_n1165__, new_new_n1166__, new_new_n1167__,
    new_new_n1168__, new_new_n1169__, new_new_n1170__, new_new_n1171__,
    new_new_n1172__, new_new_n1173__, new_new_n1174__, new_new_n1175__,
    new_new_n1176__, new_new_n1177__, new_new_n1178__, new_new_n1179__,
    new_new_n1180__, new_new_n1181__, new_new_n1182__, new_new_n1183__,
    new_new_n1184__, new_new_n1185__, new_new_n1186__, new_new_n1187__,
    new_new_n1188__, new_new_n1189__, new_new_n1190__, new_new_n1191__,
    new_new_n1192__, new_new_n1193__, new_new_n1194__, new_new_n1195__,
    new_new_n1196__, new_new_n1197__, new_new_n1198__, new_new_n1199__,
    new_new_n1200__, new_new_n1201__, new_new_n1202__, new_new_n1203__,
    new_new_n1204__, new_new_n1205__, new_new_n1206__, new_new_n1207__,
    new_new_n1208__, new_new_n1209__, new_new_n1210__, new_new_n1211__,
    new_new_n1212__, new_new_n1213__, new_new_n1214__, new_new_n1215__,
    new_new_n1216__, new_new_n1217__, new_new_n1218__, new_new_n1219__,
    new_new_n1220__, new_new_n1221__, new_new_n1222__, new_new_n1223__,
    new_new_n1224__, new_new_n1225__, new_new_n1226__, new_new_n1227__,
    new_new_n1228__, new_new_n1229__, new_new_n1230__, new_new_n1231__,
    new_new_n1232__, new_new_n1233__, new_new_n1234__, new_new_n1235__,
    new_new_n1236__, new_new_n1237__, new_new_n1238__, new_new_n1239__,
    new_new_n1240__, new_new_n1241__, new_new_n1242__, new_new_n1243__,
    new_new_n1244__, new_new_n1245__, new_new_n1246__, new_new_n1247__,
    new_new_n1248__, new_new_n1249__, new_new_n1250__, new_new_n1251__,
    new_new_n1252__, new_new_n1253__, new_new_n1254__, new_new_n1255__,
    new_new_n1256__, new_new_n1257__, new_new_n1258__, new_new_n1259__,
    new_new_n1260__, new_new_n1261__, new_new_n1262__, new_new_n1263__,
    new_new_n1264__, new_new_n1265__, new_new_n1266__, new_new_n1267__,
    new_new_n1268__, new_new_n1269__, new_new_n1270__, new_new_n1271__,
    new_new_n1272__, new_new_n1273__, new_new_n1274__, new_new_n1275__,
    new_new_n1276__, new_new_n1277__, new_new_n1278__, new_new_n1279__,
    new_new_n1280__, new_new_n1281__, new_new_n1282__, new_new_n1283__,
    new_new_n1284__, new_new_n1285__, new_new_n1286__, new_new_n1287__,
    new_new_n1288__, new_new_n1289__, new_new_n1290__, new_new_n1291__,
    new_new_n1292__, new_new_n1293__, new_new_n1294__, new_new_n1295__,
    new_new_n1296__, new_new_n1297__, new_new_n1298__, new_new_n1299__,
    new_new_n1300__, new_new_n1301__, new_new_n1302__, new_new_n1303__,
    new_new_n1304__, new_new_n1305__, new_new_n1306__, new_new_n1307__,
    new_new_n1308__, new_new_n1309__, new_new_n1310__, new_new_n1311__,
    new_new_n1312__, new_new_n1313__, new_new_n1314__, new_new_n1315__,
    new_new_n1316__, new_new_n1317__, new_new_n1318__, new_new_n1319__,
    new_new_n1320__, new_new_n1321__, new_new_n1322__, new_new_n1323__,
    new_new_n1324__, new_new_n1325__, new_new_n1326__, new_new_n1327__,
    new_new_n1328__, new_new_n1329__, new_new_n1330__, new_new_n1331__,
    new_new_n1332__, new_new_n1333__, new_new_n1334__, new_new_n1335__,
    new_new_n1336__, new_new_n1337__, new_new_n1338__, new_new_n1339__,
    new_new_n1340__, new_new_n1341__, new_new_n1342__, new_new_n1343__,
    new_new_n1344__, new_new_n1345__, new_new_n1346__, new_new_n1347__,
    new_new_n1348__, new_new_n1349__, new_new_n1350__, new_new_n1351__,
    new_new_n1352__, new_new_n1353__, new_new_n1354__, new_new_n1355__,
    new_new_n1356__, new_new_n1357__, new_new_n1358__, new_new_n1359__,
    new_new_n1360__, new_new_n1361__, new_new_n1362__, new_new_n1363__,
    new_new_n1364__, new_new_n1365__, new_new_n1366__, new_new_n1367__,
    new_new_n1368__, new_new_n1369__, new_new_n1370__, new_new_n1371__,
    new_new_n1372__, new_new_n1373__, new_new_n1374__, new_new_n1375__,
    new_new_n1376__, new_new_n1377__, new_new_n1378__, new_new_n1379__,
    new_new_n1380__, new_new_n1381__, new_new_n1382__, new_new_n1383__,
    new_new_n1384__, new_new_n1385__, new_new_n1386__, new_new_n1387__,
    new_new_n1388__, new_new_n1389__, new_new_n1390__, new_new_n1391__,
    new_new_n1392__, new_new_n1393__, new_new_n1394__, new_new_n1395__,
    new_new_n1396__, new_new_n1397__, new_new_n1398__, new_new_n1399__,
    new_new_n1400__, new_new_n1401__, new_new_n1402__, new_new_n1403__,
    new_new_n1404__, new_new_n1405__, new_new_n1406__, new_new_n1407__,
    new_new_n1408__, new_new_n1409__, new_new_n1410__, new_new_n1411__,
    new_new_n1412__, new_new_n1413__, new_new_n1414__, new_new_n1415__,
    new_new_n1416__, new_new_n1417__, new_new_n1418__, new_new_n1419__,
    new_new_n1420__, new_new_n1421__, new_new_n1422__, new_new_n1423__,
    new_new_n1424__, new_new_n1425__, new_new_n1426__, new_new_n1427__,
    new_new_n1428__, new_new_n1429__, new_new_n1430__, new_new_n1431__,
    new_new_n1432__, new_new_n1433__, new_new_n1434__, new_new_n1435__,
    new_new_n1436__, new_new_n1437__, new_new_n1438__, new_new_n1439__,
    new_new_n1440__, new_new_n1441__, new_new_n1442__, new_new_n1443__,
    new_new_n1444__, new_new_n1445__, new_new_n1446__, new_new_n1447__,
    new_new_n1448__, new_new_n1449__, new_new_n1450__, new_new_n1451__,
    new_new_n1452__, new_new_n1453__, new_new_n1454__, new_new_n1455__,
    new_new_n1456__, new_new_n1457__, new_new_n1458__, new_new_n1459__,
    new_new_n1460__, new_new_n1461__, new_new_n1462__, new_new_n1463__,
    new_new_n1464__, new_new_n1465__, new_new_n1466__, new_new_n1467__,
    new_new_n1468__, new_new_n1469__, new_new_n1470__, new_new_n1471__,
    new_new_n1472__, new_new_n1473__, new_new_n1474__, new_new_n1475__,
    new_new_n1476__, new_new_n1477__, new_new_n1478__, new_new_n1479__,
    new_new_n1480__, new_new_n1481__, new_new_n1482__, new_new_n1483__,
    new_new_n1484__, new_new_n1485__, new_new_n1486__, new_new_n1487__,
    new_new_n1488__, new_new_n1489__, new_new_n1490__, new_new_n1491__,
    new_new_n1492__, new_new_n1493__, new_new_n1494__, new_new_n1495__,
    new_new_n1496__, new_new_n1497__, new_new_n1498__, new_new_n1499__,
    new_new_n1500__, new_new_n1501__, new_new_n1502__, new_new_n1503__,
    new_new_n1504__, new_new_n1505__, new_new_n1506__, new_new_n1507__,
    new_new_n1508__, new_new_n1509__, new_new_n1510__, new_new_n1511__,
    new_new_n1512__, new_new_n1513__, new_new_n1514__, new_new_n1515__,
    new_new_n1516__, new_new_n1517__, new_new_n1518__, new_new_n1519__,
    new_new_n1520__, new_new_n1521__, new_new_n1522__, new_new_n1523__,
    new_new_n1524__, new_new_n1525__, new_new_n1526__, new_new_n1527__,
    new_new_n1528__, new_new_n1529__, new_new_n1530__, new_new_n1531__,
    new_new_n1532__, new_new_n1533__, new_new_n1534__, new_new_n1535__,
    new_new_n1536__, new_new_n1537__, new_new_n1538__, new_new_n1539__,
    new_new_n1540__, new_new_n1541__, new_new_n1542__, new_new_n1543__,
    new_new_n1544__, new_new_n1545__, new_new_n1546__, new_new_n1547__,
    new_new_n1548__, new_new_n1549__, new_new_n1550__, new_new_n1551__,
    new_new_n1552__, new_new_n1553__, new_new_n1554__, new_new_n1555__,
    new_new_n1556__, new_new_n1557__, new_new_n1558__, new_new_n1559__,
    new_new_n1560__, new_new_n1561__, new_new_n1562__, new_new_n1563__,
    new_new_n1564__, new_new_n1565__, new_new_n1566__, new_new_n1567__,
    new_new_n1568__, new_new_n1569__, new_new_n1570__, new_new_n1571__,
    new_new_n1572__, new_new_n1573__, new_new_n1574__, new_new_n1575__,
    new_new_n1576__, new_new_n1577__, new_new_n1578__, new_new_n1579__,
    new_new_n1580__, new_new_n1581__, new_new_n1582__, new_new_n1583__,
    new_new_n1584__, new_new_n1585__, new_new_n1586__, new_new_n1587__,
    new_new_n1588__, new_new_n1589__, new_new_n1590__, new_new_n1591__,
    new_new_n1592__, new_new_n1593__, new_new_n1594__, new_new_n1595__,
    new_new_n1596__, new_new_n1597__, new_new_n1598__, new_new_n1599__,
    new_new_n1600__, new_new_n1601__, new_new_n1602__, new_new_n1603__,
    new_new_n1604__, new_new_n1605__, new_new_n1606__, new_new_n1607__,
    new_new_n1608__, new_new_n1609__, new_new_n1610__, new_new_n1611__,
    new_new_n1612__, new_new_n1613__, new_new_n1614__, new_new_n1615__,
    new_new_n1616__, new_new_n1617__, new_new_n1618__, new_new_n1619__,
    new_new_n1620__, new_new_n1621__, new_new_n1622__, new_new_n1623__,
    new_new_n1624__, new_new_n1625__, new_new_n1626__, new_new_n1627__,
    new_new_n1628__, new_new_n1629__, new_new_n1630__, new_new_n1631__,
    new_new_n1632__, new_new_n1633__, new_new_n1634__, new_new_n1635__,
    new_new_n1636__, new_new_n1637__, new_new_n1638__, new_new_n1639__,
    new_new_n1640__, new_new_n1641__, new_new_n1642__, new_new_n1643__,
    new_new_n1644__, new_new_n1645__, new_new_n1646__, new_new_n1647__,
    new_new_n1648__, new_new_n1649__, new_new_n1650__, new_new_n1651__,
    new_new_n1652__, new_new_n1653__, new_new_n1654__, new_new_n1655__,
    new_new_n1656__, new_new_n1657__, new_new_n1658__, new_new_n1659__,
    new_new_n1660__, new_new_n1661__, new_new_n1662__, new_new_n1663__,
    new_new_n1664__, new_new_n1665__, new_new_n1666__, new_new_n1667__,
    new_new_n1668__, new_new_n1669__, new_new_n1670__, new_new_n1671__,
    new_new_n1672__, new_new_n1673__, new_new_n1674__, new_new_n1675__,
    new_new_n1676__, new_new_n1677__, new_new_n1678__, new_new_n1679__,
    new_new_n1680__, new_new_n1681__, new_new_n1682__, new_new_n1683__,
    new_new_n1684__, new_new_n1685__, new_new_n1686__, new_new_n1687__,
    new_new_n1688__, new_new_n1689__, new_new_n1690__, new_new_n1691__,
    new_new_n1692__, new_new_n1693__, new_new_n1694__, new_new_n1695__,
    new_new_n1696__, new_new_n1697__, new_new_n1698__, new_new_n1699__,
    new_new_n1700__, new_new_n1701__, new_new_n1702__, new_new_n1703__,
    new_new_n1704__, new_new_n1705__, new_new_n1706__, new_new_n1707__,
    new_new_n1708__, new_new_n1709__, new_new_n1710__, new_new_n1711__,
    new_new_n1712__, new_new_n1713__, new_new_n1714__, new_new_n1715__,
    new_new_n1716__, new_new_n1717__, new_new_n1718__, new_new_n1719__,
    new_new_n1948__, new_new_n1949__, new_new_n1950__, new_new_n1951__,
    new_new_n1952__, new_new_n1953__, new_new_n1954__, new_new_n1955__,
    new_new_n1956__, new_new_n1957__, new_new_n1958__, new_new_n1959__,
    new_new_n1960__, new_new_n1961__, new_new_n1962__, new_new_n1963__,
    new_new_n1964__, new_new_n1965__, new_new_n1966__, new_new_n1967__,
    new_new_n1968__, new_new_n1969__, new_new_n1970__, new_new_n1971__,
    new_new_n1972__, new_new_n1973__, new_new_n1974__, new_new_n1975__,
    new_new_n1976__, new_new_n1977__, new_new_n1978__, new_new_n1979__,
    new_new_n1980__, new_new_n1981__, new_new_n1982__, new_new_n1983__,
    new_new_n1984__, new_new_n1985__, new_new_n1986__, new_new_n1987__,
    new_new_n1988__, new_new_n1989__, new_new_n1990__, new_new_n1991__,
    new_new_n1992__, new_new_n1993__, new_new_n1994__, new_new_n1995__,
    new_new_n1996__, new_new_n1997__, new_new_n1998__, new_new_n1999__,
    new_new_n2000__, new_new_n2001__, new_new_n2002__, new_new_n2003__,
    new_new_n2004__, new_new_n2005__, new_new_n2006__, new_new_n2007__,
    new_new_n2008__, new_new_n2009__, new_new_n2010__, new_new_n2011__,
    new_new_n2012__, new_new_n2013__, new_new_n2014__, new_new_n2015__,
    new_new_n2016__, new_new_n2017__, new_new_n2018__, new_new_n2019__,
    new_new_n2020__, new_new_n2021__, new_new_n2022__, new_new_n2023__,
    new_new_n2024__, new_new_n2025__, new_new_n2026__, new_new_n2027__,
    new_new_n2028__, new_new_n2029__, new_new_n2030__, new_new_n2031__,
    new_new_n2032__, new_new_n2033__, new_new_n2034__, new_new_n2035__,
    new_new_n2036__, new_new_n2037__, new_new_n2038__, new_new_n2039__,
    new_new_n2040__, new_new_n2041__, new_new_n2042__, new_new_n2043__,
    new_new_n2044__, new_new_n2045__, new_new_n2046__, new_new_n2047__,
    new_new_n2048__, new_new_n2049__, new_new_n2050__, new_new_n2051__,
    new_new_n2052__, new_new_n2053__, new_new_n2054__, new_new_n2055__,
    new_new_n2056__, new_new_n2057__, new_new_n2058__, new_new_n2059__,
    new_new_n2060__, new_new_n2061__, new_new_n2062__, new_new_n2063__,
    new_new_n2064__, new_new_n2065__, new_new_n2066__, new_new_n2067__,
    new_new_n2068__, new_new_n2069__, new_new_n2070__, new_new_n2071__,
    new_new_n2072__, new_new_n2073__, new_new_n2074__, new_new_n2075__,
    new_new_n2076__, new_new_n2077__, new_new_n2078__, new_new_n2079__,
    new_new_n2080__, new_new_n2081__, new_new_n2082__, new_new_n2083__,
    new_new_n2084__, new_new_n2085__, new_new_n2086__, new_new_n2087__,
    new_new_n2088__, new_new_n2089__, new_new_n2090__, new_new_n2091__,
    new_new_n2092__, new_new_n2093__, new_new_n2094__, new_new_n2095__,
    new_new_n2096__, new_new_n2097__, new_new_n2098__, new_new_n2099__,
    new_new_n2100__, new_new_n2101__, new_new_n2102__, new_new_n2103__,
    new_new_n2104__, new_new_n2105__, new_new_n2106__, new_new_n2107__,
    new_new_n2108__, new_new_n2109__, new_new_n2110__, new_new_n2111__,
    new_new_n2112__, new_new_n2113__, new_new_n2114__, new_new_n2115__,
    new_new_n2116__, new_new_n2117__, new_new_n2118__, new_new_n2119__,
    new_new_n2120__, new_new_n2121__, new_new_n2122__, new_new_n2123__,
    new_new_n2124__, new_new_n2125__, new_new_n2126__, new_new_n2127__,
    new_new_n2128__, new_new_n2129__, new_new_n2130__, new_new_n2131__,
    new_new_n2132__, new_new_n2133__, new_new_n2134__, new_new_n2135__,
    new_new_n2136__, new_new_n2137__, new_new_n2138__, new_new_n2139__,
    new_new_n2140__, new_new_n2141__, new_new_n2142__, new_new_n2143__,
    new_new_n2144__, new_new_n2145__, new_new_n2146__, new_new_n2147__,
    new_new_n2148__, new_new_n2149__, new_new_n2150__, new_new_n2151__,
    new_new_n2152__, new_new_n2153__, new_new_n2154__, new_new_n2155__,
    new_new_n2156__, new_new_n2157__, new_new_n2158__, new_new_n2159__,
    new_new_n2160__, new_new_n2161__, new_new_n2162__, new_new_n2163__,
    new_new_n2164__, new_new_n2165__, new_new_n2166__, new_new_n2167__,
    new_new_n2168__, new_new_n2169__, new_new_n2170__, new_new_n2171__,
    new_new_n2172__, new_new_n2173__, new_new_n2174__, new_new_n2175__,
    new_new_n2176__, new_new_n2177__, new_new_n2178__, new_new_n2179__,
    new_new_n2180__, new_new_n2181__, new_new_n2182__, new_new_n2183__,
    new_new_n2184__, new_new_n2185__, new_new_n2186__, new_new_n2187__,
    new_new_n2188__, new_new_n2189__, new_new_n2190__, new_new_n2191__,
    new_new_n2192__, new_new_n2193__, new_new_n2194__, new_new_n2195__,
    new_new_n2196__, new_new_n2197__, new_new_n2198__, new_new_n2199__,
    new_new_n2200__, new_new_n2201__, new_new_n2202__, new_new_n2203__,
    new_new_n2204__, new_new_n2205__, new_new_n2206__, new_new_n2207__,
    new_new_n2208__, new_new_n2209__, new_new_n2210__, new_new_n2211__,
    new_new_n2212__, new_new_n2213__, new_new_n2214__, new_new_n2215__,
    new_new_n2216__, new_new_n2217__, new_new_n2218__, new_new_n2219__,
    new_new_n2220__, new_new_n2221__, new_new_n2222__, new_new_n2223__,
    new_new_n2224__, new_new_n2225__, new_new_n2226__, new_new_n2227__,
    new_new_n2228__, new_new_n2229__, new_new_n2230__, new_new_n2231__,
    new_new_n2232__, new_new_n2233__, new_new_n2234__, new_new_n2235__,
    new_new_n2236__, new_new_n2237__, new_new_n2238__, new_new_n2239__,
    new_new_n2240__, new_new_n2241__, new_new_n2242__, new_new_n2243__,
    new_new_n2244__, new_new_n2245__, new_new_n2246__, new_new_n2247__,
    new_new_n2248__, new_new_n2249__, new_new_n2250__, new_new_n2251__,
    new_new_n2252__, new_new_n2253__, new_new_n2254__, new_new_n2255__,
    new_new_n2256__, new_new_n2257__, new_new_n2258__, new_new_n2259__,
    new_new_n2260__, new_new_n2261__, new_new_n2262__, new_new_n2263__,
    new_new_n2264__, new_new_n2265__, new_new_n2266__, new_new_n2267__,
    new_new_n2268__, new_new_n2269__, new_new_n2270__, new_new_n2271__,
    new_new_n2272__, new_new_n2273__, new_new_n2274__, new_new_n2275__,
    new_new_n2276__, new_new_n2277__, new_new_n2278__, new_new_n2279__,
    new_new_n2280__, new_new_n2281__, new_new_n2282__, new_new_n2283__,
    new_new_n2284__, new_new_n2285__, new_new_n2286__, new_new_n2287__,
    new_new_n2288__, new_new_n2289__, new_new_n2290__, new_new_n2291__,
    new_new_n2292__, new_new_n2293__, new_new_n2294__, new_new_n2295__,
    new_new_n2296__, new_new_n2297__, new_new_n2298__, new_new_n2299__,
    new_new_n2300__, new_new_n2301__, new_new_n2302__, new_new_n2303__,
    new_new_n2304__, new_new_n2305__, new_new_n2306__, new_new_n2307__,
    new_new_n2308__, new_new_n2309__, new_new_n2310__, new_new_n2311__,
    new_new_n2312__, new_new_n2313__, new_new_n2314__, new_new_n2315__,
    new_new_n2316__, new_new_n2317__, new_new_n2318__, new_new_n2319__,
    new_new_n2320__, new_new_n2321__, new_new_n2322__, new_new_n2323__,
    new_new_n2324__, new_new_n2325__, new_new_n2326__, new_new_n2327__,
    new_new_n2328__, new_new_n2329__, new_new_n2330__, new_new_n2331__,
    new_new_n2332__, new_new_n2333__, new_new_n2334__, new_new_n2335__,
    new_new_n2336__, new_new_n2337__, new_new_n2338__, new_new_n2339__,
    new_new_n2340__, new_new_n2341__, new_new_n2342__, new_new_n2343__,
    new_new_n2344__, new_new_n2345__, new_new_n2346__, new_new_n2347__,
    new_new_n2348__, new_new_n2349__, new_new_n2350__, new_new_n2351__,
    new_new_n2352__, new_new_n2353__, new_new_n2354__, new_new_n2355__,
    new_new_n2356__, new_new_n2357__, new_new_n2358__, new_new_n2359__,
    new_new_n2360__, new_new_n2361__, new_new_n2362__, new_new_n2363__,
    new_new_n2364__, new_new_n2365__, new_new_n2366__, new_new_n2367__,
    new_new_n2368__, new_new_n2369__, new_new_n2370__, new_new_n2371__,
    new_new_n2372__, new_new_n2373__, new_new_n2374__, new_new_n2375__,
    new_new_n2376__, new_new_n2377__, new_new_n2378__, new_new_n2379__,
    new_new_n2380__, new_new_n2381__, new_new_n2382__, new_new_n2383__,
    new_new_n2384__, new_new_n2385__, new_new_n2386__, new_new_n2387__,
    new_new_n2388__, new_new_n2389__, new_new_n2390__, new_new_n2391__,
    new_new_n2392__, new_new_n2393__, new_new_n2394__, new_new_n2395__,
    new_new_n2396__, new_new_n2397__, new_new_n2398__, new_new_n2399__,
    new_new_n2400__, new_new_n2401__, new_new_n2402__, new_new_n2403__,
    new_new_n2404__, new_new_n2405__, new_new_n2406__, new_new_n2407__,
    new_new_n2408__, new_new_n2409__, new_new_n2410__, new_new_n2411__,
    new_new_n2412__, new_new_n2413__, new_new_n2414__, new_new_n2415__,
    new_new_n2416__, new_new_n2417__, new_new_n2418__, new_new_n2419__,
    new_new_n2420__, new_new_n2421__, new_new_n2422__, new_new_n2423__,
    new_new_n2424__, new_new_n2425__, new_new_n2426__, new_new_n2427__,
    new_new_n2428__, new_new_n2429__, new_new_n2430__, new_new_n2431__,
    new_new_n2432__, new_new_n2433__, new_new_n2434__, new_new_n2435__,
    new_new_n2436__, new_new_n2437__, new_new_n2438__, new_new_n2439__,
    new_new_n2440__, new_new_n2441__, new_new_n2442__, new_new_n2443__,
    new_new_n2444__, new_new_n2445__, new_new_n2446__, new_new_n2447__,
    new_new_n2448__, new_new_n2449__, new_new_n2450__, new_new_n2451__,
    new_new_n2452__, new_new_n2453__, new_new_n2454__, new_new_n2455__,
    new_new_n2456__, new_new_n2457__, new_new_n2458__, new_new_n2459__,
    new_new_n2460__, new_new_n2461__, new_new_n2462__, new_new_n2463__,
    new_new_n2464__, new_new_n2465__, new_new_n2466__, new_new_n2467__,
    new_new_n2468__, new_new_n2469__, new_new_n2470__, new_new_n2471__,
    new_new_n2472__, new_new_n2473__, new_new_n2474__, new_new_n2475__,
    new_new_n2476__, new_new_n2477__, new_new_n2478__, new_new_n2479__,
    new_new_n2480__, new_new_n2481__, new_new_n2482__, new_new_n2483__,
    new_new_n2484__, new_new_n2485__, new_new_n2486__, new_new_n2487__,
    new_new_n2488__, new_new_n2489__, new_new_n2490__, new_new_n2491__,
    new_new_n2492__, new_new_n2493__, new_new_n2494__, new_new_n2495__,
    new_new_n2496__, new_new_n2497__, new_new_n2498__, new_new_n2499__,
    new_new_n2500__, new_new_n2501__, new_new_n2502__, new_new_n2503__,
    new_new_n2504__, new_new_n2505__, new_new_n2506__, new_new_n2507__,
    new_new_n2508__, new_new_n2509__, new_new_n2510__, new_new_n2511__,
    new_new_n2512__, new_new_n2513__, new_new_n2514__, new_new_n2515__,
    new_new_n2516__, new_new_n2517__, new_new_n2518__, new_new_n2519__,
    new_new_n2520__, new_new_n2521__, new_new_n2522__, new_new_n2523__,
    new_new_n2524__, new_new_n2525__, new_new_n2526__, new_new_n2527__,
    new_new_n2528__, new_new_n2529__, new_new_n2530__, new_new_n2531__,
    new_new_n2532__, new_new_n2533__, new_new_n2534__, new_new_n2535__,
    new_new_n2536__, new_new_n2537__, new_new_n2538__, new_new_n2539__,
    new_new_n2540__, new_new_n2541__, new_new_n2542__, new_new_n2543__,
    new_new_n2544__, new_new_n2545__, new_new_n2546__, new_new_n2547__,
    new_new_n2548__, new_new_n2549__, new_new_n2550__, new_new_n2551__,
    new_new_n2552__, new_new_n2553__, new_new_n2554__, new_new_n2555__,
    new_new_n2556__, new_new_n2557__, new_new_n2558__, new_new_n2559__,
    new_new_n2560__, new_new_n2561__, new_new_n2562__, new_new_n2563__,
    n4343, n4346, n4349, n4352, n4355, n4358, n4361, n4364, n4367, n4370,
    n4373, n4376, n4379, n4382, n4385, n4388, n4391, n4394, n4397, n4400,
    n4403, n4406, n4409, n4412, n4415, n4418, n4421, n4424, n4427, n4430,
    n4433, n4436, n4439, n4442, n4445, n4448, n4451, n4454, n4457, n4460,
    n4463, n4466, n4469, n4472, n4475, n4478, n4481, n4484, n4487, n4490,
    n4493, n4496, n4499, n4502, n4505, n4508, n4511, n4514, n4517, n4520,
    n4523, n4526, n4529, n4532, n4535, n4538, n4541, n4544, n4547, n4550,
    n4553, n4556, n4559, n4562, n4565, n4568, n4571, n4574, n4577, n4580,
    n4583, n4586, n4589, n4592, n4595, n4598, n4601, n4604, n4607, n4610,
    n4613, n4616, n4619, n4622, n4625, n4628, n4631, n4634, n4637, n4640,
    n4643, n4646, n4649, n4652, n4655, n4658, n4661, n4664, n4667, n4670,
    n4673, n4676, n4679, n4682, n4685, n4688, n4691, n4694, n4697, n4700,
    n4703, n4706, n4709, n4712, n4715, n4718, n4721, n4724, n4727, n4730,
    n4733, n4736, n4739, n4742, n4745, n4748, n4751, n4754, n4757, n4760,
    n4763, n4766, n4769, n4772, n4775, n4778, n4781, n4784, n4787, n4790,
    n4793, n4796, n4799, n4802, n4805, n4808, n4811, n4814, n4817, n4820,
    n4823, n4826, n4829, n4832, n4835, n4838, n4841, n4844, n4847, n4850,
    n4853, n4856, n4859, n4862, n4865, n4868, n4871, n4874, n4877, n4880,
    n4883, n4886, n4889, n4892, n4895, n4898, n4901, n4904, n4907, n4910,
    n4913, n4916, n4919, n4922, n4925, n4928;
  not1  g0000(.din(G1), .dout(new_new_n467__));
  not1  g0001(.din(G2), .dout(new_new_n469__));
  not1  g0002(.din(G3), .dout(new_new_n471__));
  not1  g0003(.din(G4), .dout(new_new_n473__));
  not1  g0004(.din(G5), .dout(new_new_n475__));
  not1  g0005(.din(G6), .dout(new_new_n477__));
  not1  g0006(.din(G7), .dout(new_new_n479__));
  not1  g0007(.din(G8), .dout(new_new_n481__));
  not1  g0008(.din(G9), .dout(new_new_n483__));
  not1  g0009(.din(G10), .dout(new_new_n485__));
  not1  g0010(.din(G11), .dout(new_new_n487__));
  not1  g0011(.din(G12), .dout(new_new_n489__));
  not1  g0012(.din(G13), .dout(new_new_n491__));
  not1  g0013(.din(G14), .dout(new_new_n493__));
  not1  g0014(.din(G15), .dout(new_new_n495__));
  not1  g0015(.din(G16), .dout(new_new_n497__));
  not1  g0016(.din(G17), .dout(new_new_n499__));
  not1  g0017(.din(G18), .dout(new_new_n501__));
  not1  g0018(.din(G19), .dout(new_new_n503__));
  not1  g0019(.din(G20), .dout(new_new_n505__));
  not1  g0020(.din(G21), .dout(new_new_n507__));
  not1  g0021(.din(G22), .dout(new_new_n509__));
  not1  g0022(.din(G23), .dout(new_new_n511__));
  not1  g0023(.din(G24), .dout(new_new_n513__));
  not1  g0024(.din(G25), .dout(new_new_n515__));
  not1  g0025(.din(G26), .dout(new_new_n517__));
  not1  g0026(.din(G27), .dout(new_new_n519__));
  not1  g0027(.din(G28), .dout(new_new_n521__));
  not1  g0028(.din(G29), .dout(new_new_n523__));
  not1  g0029(.din(G30), .dout(new_new_n525__));
  not1  g0030(.din(G31), .dout(new_new_n527__));
  not1  g0031(.din(G32), .dout(new_new_n529__));
  not1  g0032(.din(G33), .dout(new_new_n531__));
  not1  g0033(.din(G34), .dout(new_new_n533__));
  not1  g0034(.din(G35), .dout(new_new_n535__));
  not1  g0035(.din(G36), .dout(new_new_n537__));
  not1  g0036(.din(G37), .dout(new_new_n539__));
  not1  g0037(.din(G38), .dout(new_new_n541__));
  not1  g0038(.din(G39), .dout(new_new_n543__));
  not1  g0039(.din(G40), .dout(new_new_n545__));
  not1  g0040(.din(G41), .dout(new_new_n547__));
  buf1  g0041(.din(n630_lo), .dout(new_new_n548__));
  not1  g0042(.din(n630_lo), .dout(new_new_n549__));
  buf1  g0043(.din(n642_lo), .dout(new_new_n550__));
  not1  g0044(.din(n642_lo), .dout(new_new_n551__));
  buf1  g0045(.din(n654_lo), .dout(new_new_n552__));
  not1  g0046(.din(n654_lo), .dout(new_new_n553__));
  buf1  g0047(.din(n666_lo), .dout(new_new_n554__));
  not1  g0048(.din(n666_lo), .dout(new_new_n555__));
  buf1  g0049(.din(n678_lo), .dout(new_new_n556__));
  not1  g0050(.din(n678_lo), .dout(new_new_n557__));
  buf1  g0051(.din(n690_lo), .dout(new_new_n558__));
  not1  g0052(.din(n690_lo), .dout(new_new_n559__));
  buf1  g0053(.din(n702_lo), .dout(new_new_n560__));
  not1  g0054(.din(n702_lo), .dout(new_new_n561__));
  buf1  g0055(.din(n714_lo), .dout(new_new_n562__));
  not1  g0056(.din(n714_lo), .dout(new_new_n563__));
  buf1  g0057(.din(n726_lo), .dout(new_new_n564__));
  not1  g0058(.din(n726_lo), .dout(new_new_n565__));
  buf1  g0059(.din(n738_lo), .dout(new_new_n566__));
  not1  g0060(.din(n738_lo), .dout(new_new_n567__));
  buf1  g0061(.din(n750_lo), .dout(new_new_n568__));
  not1  g0062(.din(n750_lo), .dout(new_new_n569__));
  buf1  g0063(.din(n762_lo), .dout(new_new_n570__));
  not1  g0064(.din(n762_lo), .dout(new_new_n571__));
  buf1  g0065(.din(n774_lo), .dout(new_new_n572__));
  not1  g0066(.din(n774_lo), .dout(new_new_n573__));
  buf1  g0067(.din(n786_lo), .dout(new_new_n574__));
  not1  g0068(.din(n786_lo), .dout(new_new_n575__));
  buf1  g0069(.din(n798_lo), .dout(new_new_n576__));
  not1  g0070(.din(n798_lo), .dout(new_new_n577__));
  buf1  g0071(.din(n810_lo), .dout(new_new_n578__));
  not1  g0072(.din(n810_lo), .dout(new_new_n579__));
  buf1  g0073(.din(n822_lo), .dout(new_new_n580__));
  not1  g0074(.din(n822_lo), .dout(new_new_n581__));
  buf1  g0075(.din(n834_lo), .dout(new_new_n582__));
  not1  g0076(.din(n834_lo), .dout(new_new_n583__));
  buf1  g0077(.din(n846_lo), .dout(new_new_n584__));
  not1  g0078(.din(n846_lo), .dout(new_new_n585__));
  buf1  g0079(.din(n858_lo), .dout(new_new_n586__));
  not1  g0080(.din(n858_lo), .dout(new_new_n587__));
  buf1  g0081(.din(n870_lo), .dout(new_new_n588__));
  not1  g0082(.din(n870_lo), .dout(new_new_n589__));
  buf1  g0083(.din(n882_lo), .dout(new_new_n590__));
  not1  g0084(.din(n882_lo), .dout(new_new_n591__));
  buf1  g0085(.din(n894_lo), .dout(new_new_n592__));
  not1  g0086(.din(n894_lo), .dout(new_new_n593__));
  buf1  g0087(.din(n906_lo), .dout(new_new_n594__));
  not1  g0088(.din(n906_lo), .dout(new_new_n595__));
  buf1  g0089(.din(n918_lo), .dout(new_new_n596__));
  not1  g0090(.din(n918_lo), .dout(new_new_n597__));
  buf1  g0091(.din(n930_lo), .dout(new_new_n598__));
  not1  g0092(.din(n930_lo), .dout(new_new_n599__));
  buf1  g0093(.din(n942_lo), .dout(new_new_n600__));
  not1  g0094(.din(n942_lo), .dout(new_new_n601__));
  buf1  g0095(.din(n954_lo), .dout(new_new_n602__));
  not1  g0096(.din(n954_lo), .dout(new_new_n603__));
  buf1  g0097(.din(n966_lo), .dout(new_new_n604__));
  not1  g0098(.din(n966_lo), .dout(new_new_n605__));
  buf1  g0099(.din(n978_lo), .dout(new_new_n606__));
  not1  g0100(.din(n978_lo), .dout(new_new_n607__));
  buf1  g0101(.din(n990_lo), .dout(new_new_n608__));
  not1  g0102(.din(n990_lo), .dout(new_new_n609__));
  buf1  g0103(.din(n1002_lo), .dout(new_new_n610__));
  not1  g0104(.din(n1002_lo), .dout(new_new_n611__));
  not1  g0105(.din(n1005_lo), .dout(new_new_n613__));
  buf1  g0106(.din(n1008_lo), .dout(new_new_n614__));
  not1  g0107(.din(n1008_lo), .dout(new_new_n615__));
  not1  g0108(.din(n1017_lo), .dout(new_new_n617__));
  buf1  g0109(.din(n1020_lo), .dout(new_new_n618__));
  not1  g0110(.din(n1020_lo), .dout(new_new_n619__));
  not1  g0111(.din(n1029_lo), .dout(new_new_n621__));
  buf1  g0112(.din(n1032_lo), .dout(new_new_n622__));
  not1  g0113(.din(n1032_lo), .dout(new_new_n623__));
  not1  g0114(.din(n1041_lo), .dout(new_new_n625__));
  buf1  g0115(.din(n1044_lo), .dout(new_new_n626__));
  not1  g0116(.din(n1044_lo), .dout(new_new_n627__));
  not1  g0117(.din(n1053_lo), .dout(new_new_n629__));
  buf1  g0118(.din(n1056_lo), .dout(new_new_n630__));
  not1  g0119(.din(n1056_lo), .dout(new_new_n631__));
  not1  g0120(.din(n1065_lo), .dout(new_new_n633__));
  buf1  g0121(.din(n1068_lo), .dout(new_new_n634__));
  not1  g0122(.din(n1068_lo), .dout(new_new_n635__));
  not1  g0123(.din(n1077_lo), .dout(new_new_n637__));
  buf1  g0124(.din(n1080_lo), .dout(new_new_n638__));
  not1  g0125(.din(n1080_lo), .dout(new_new_n639__));
  not1  g0126(.din(n1089_lo), .dout(new_new_n641__));
  buf1  g0127(.din(n1092_lo), .dout(new_new_n642__));
  not1  g0128(.din(n1092_lo), .dout(new_new_n643__));
  not1  g0129(.din(n1101_lo), .dout(new_new_n645__));
  buf1  g0130(.din(n1104_lo), .dout(new_new_n646__));
  not1  g0131(.din(n1104_lo), .dout(new_new_n647__));
  not1  g0132(.din(n1837_o2), .dout(new_new_n649__));
  not1  g0133(.din(n1838_o2), .dout(new_new_n651__));
  not1  g0134(.din(n1839_o2), .dout(new_new_n653__));
  not1  g0135(.din(n1840_o2), .dout(new_new_n655__));
  not1  g0136(.din(n1841_o2), .dout(new_new_n657__));
  not1  g0137(.din(n1842_o2), .dout(new_new_n659__));
  not1  g0138(.din(n1843_o2), .dout(new_new_n661__));
  not1  g0139(.din(n1844_o2), .dout(new_new_n663__));
  not1  g0140(.din(n1845_o2), .dout(new_new_n665__));
  not1  g0141(.din(n1846_o2), .dout(new_new_n667__));
  not1  g0142(.din(n1847_o2), .dout(new_new_n669__));
  not1  g0143(.din(n1848_o2), .dout(new_new_n671__));
  not1  g0144(.din(n1849_o2), .dout(new_new_n673__));
  not1  g0145(.din(n1850_o2), .dout(new_new_n675__));
  not1  g0146(.din(n1851_o2), .dout(new_new_n677__));
  not1  g0147(.din(n1852_o2), .dout(new_new_n679__));
  not1  g0148(.din(n1853_o2), .dout(new_new_n681__));
  not1  g0149(.din(n1854_o2), .dout(new_new_n683__));
  not1  g0150(.din(n1855_o2), .dout(new_new_n685__));
  not1  g0151(.din(n1856_o2), .dout(new_new_n687__));
  not1  g0152(.din(n1857_o2), .dout(new_new_n689__));
  not1  g0153(.din(n1858_o2), .dout(new_new_n691__));
  not1  g0154(.din(n1859_o2), .dout(new_new_n693__));
  not1  g0155(.din(n1860_o2), .dout(new_new_n695__));
  not1  g0156(.din(n1861_o2), .dout(new_new_n697__));
  not1  g0157(.din(n1862_o2), .dout(new_new_n699__));
  not1  g0158(.din(n1863_o2), .dout(new_new_n701__));
  not1  g0159(.din(n1864_o2), .dout(new_new_n703__));
  not1  g0160(.din(n1865_o2), .dout(new_new_n705__));
  not1  g0161(.din(n1866_o2), .dout(new_new_n707__));
  not1  g0162(.din(n1867_o2), .dout(new_new_n709__));
  not1  g0163(.din(n1868_o2), .dout(new_new_n711__));
  buf1  g0164(.din(G834_o2), .dout(new_new_n712__));
  not1  g0165(.din(G834_o2), .dout(new_new_n713__));
  buf1  g0166(.din(G847_o2), .dout(new_new_n714__));
  not1  g0167(.din(G847_o2), .dout(new_new_n715__));
  buf1  g0168(.din(G860_o2), .dout(new_new_n716__));
  not1  g0169(.din(G860_o2), .dout(new_new_n717__));
  buf1  g0170(.din(G873_o2), .dout(new_new_n718__));
  not1  g0171(.din(G873_o2), .dout(new_new_n719__));
  buf1  g0172(.din(G925_o2), .dout(new_new_n720__));
  not1  g0173(.din(G925_o2), .dout(new_new_n721__));
  buf1  g0174(.din(G886_o2), .dout(new_new_n722__));
  not1  g0175(.din(G886_o2), .dout(new_new_n723__));
  buf1  g0176(.din(G912_o2), .dout(new_new_n724__));
  not1  g0177(.din(G912_o2), .dout(new_new_n725__));
  buf1  g0178(.din(G899_o2), .dout(new_new_n726__));
  not1  g0179(.din(G899_o2), .dout(new_new_n727__));
  buf1  g0180(.din(n2151_o2), .dout(new_new_n728__));
  not1  g0181(.din(n2151_o2), .dout(new_new_n729__));
  buf1  g0182(.din(n2152_o2), .dout(new_new_n730__));
  not1  g0183(.din(n2152_o2), .dout(new_new_n731__));
  buf1  g0184(.din(n2153_o2), .dout(new_new_n732__));
  not1  g0185(.din(n2153_o2), .dout(new_new_n733__));
  buf1  g0186(.din(n2154_o2), .dout(new_new_n734__));
  not1  g0187(.din(n2154_o2), .dout(new_new_n735__));
  buf1  g0188(.din(n2155_o2), .dout(new_new_n736__));
  not1  g0189(.din(n2155_o2), .dout(new_new_n737__));
  buf1  g0190(.din(n2156_o2), .dout(new_new_n738__));
  not1  g0191(.din(n2156_o2), .dout(new_new_n739__));
  buf1  g0192(.din(n2157_o2), .dout(new_new_n740__));
  not1  g0193(.din(n2157_o2), .dout(new_new_n741__));
  buf1  g0194(.din(n2158_o2), .dout(new_new_n742__));
  not1  g0195(.din(n2158_o2), .dout(new_new_n743__));
  buf1  g0196(.din(n2159_o2), .dout(new_new_n744__));
  not1  g0197(.din(n2159_o2), .dout(new_new_n745__));
  buf1  g0198(.din(n2160_o2), .dout(new_new_n746__));
  not1  g0199(.din(n2160_o2), .dout(new_new_n747__));
  buf1  g0200(.din(n2161_o2), .dout(new_new_n748__));
  not1  g0201(.din(n2161_o2), .dout(new_new_n749__));
  buf1  g0202(.din(n2162_o2), .dout(new_new_n750__));
  not1  g0203(.din(n2162_o2), .dout(new_new_n751__));
  buf1  g0204(.din(n2163_o2), .dout(new_new_n752__));
  not1  g0205(.din(n2163_o2), .dout(new_new_n753__));
  buf1  g0206(.din(n2164_o2), .dout(new_new_n754__));
  not1  g0207(.din(n2164_o2), .dout(new_new_n755__));
  buf1  g0208(.din(n2165_o2), .dout(new_new_n756__));
  not1  g0209(.din(n2165_o2), .dout(new_new_n757__));
  buf1  g0210(.din(n2166_o2), .dout(new_new_n758__));
  not1  g0211(.din(n2166_o2), .dout(new_new_n759__));
  buf1  g0212(.din(n2167_o2), .dout(new_new_n760__));
  not1  g0213(.din(n2167_o2), .dout(new_new_n761__));
  buf1  g0214(.din(n2168_o2), .dout(new_new_n762__));
  not1  g0215(.din(n2168_o2), .dout(new_new_n763__));
  buf1  g0216(.din(n2169_o2), .dout(new_new_n764__));
  not1  g0217(.din(n2169_o2), .dout(new_new_n765__));
  buf1  g0218(.din(n2170_o2), .dout(new_new_n766__));
  not1  g0219(.din(n2170_o2), .dout(new_new_n767__));
  buf1  g0220(.din(n2171_o2), .dout(new_new_n768__));
  not1  g0221(.din(n2171_o2), .dout(new_new_n769__));
  buf1  g0222(.din(n2172_o2), .dout(new_new_n770__));
  not1  g0223(.din(n2172_o2), .dout(new_new_n771__));
  buf1  g0224(.din(n2173_o2), .dout(new_new_n772__));
  not1  g0225(.din(n2173_o2), .dout(new_new_n773__));
  buf1  g0226(.din(n2174_o2), .dout(new_new_n774__));
  not1  g0227(.din(n2174_o2), .dout(new_new_n775__));
  buf1  g0228(.din(n2175_o2), .dout(new_new_n776__));
  not1  g0229(.din(n2175_o2), .dout(new_new_n777__));
  buf1  g0230(.din(n2176_o2), .dout(new_new_n778__));
  not1  g0231(.din(n2176_o2), .dout(new_new_n779__));
  buf1  g0232(.din(n2177_o2), .dout(new_new_n780__));
  not1  g0233(.din(n2177_o2), .dout(new_new_n781__));
  buf1  g0234(.din(n2178_o2), .dout(new_new_n782__));
  not1  g0235(.din(n2178_o2), .dout(new_new_n783__));
  buf1  g0236(.din(n2179_o2), .dout(new_new_n784__));
  not1  g0237(.din(n2179_o2), .dout(new_new_n785__));
  buf1  g0238(.din(n2180_o2), .dout(new_new_n786__));
  not1  g0239(.din(n2180_o2), .dout(new_new_n787__));
  buf1  g0240(.din(n2181_o2), .dout(new_new_n788__));
  not1  g0241(.din(n2181_o2), .dout(new_new_n789__));
  buf1  g0242(.din(n2182_o2), .dout(new_new_n790__));
  not1  g0243(.din(n2182_o2), .dout(new_new_n791__));
  buf1  g0244(.din(G974_o2), .dout(new_new_n792__));
  not1  g0245(.din(G974_o2), .dout(new_new_n793__));
  buf1  g0246(.din(G976_o2), .dout(new_new_n794__));
  not1  g0247(.din(G976_o2), .dout(new_new_n795__));
  buf1  g0248(.din(G970_o2), .dout(new_new_n796__));
  not1  g0249(.din(G970_o2), .dout(new_new_n797__));
  buf1  g0250(.din(G972_o2), .dout(new_new_n798__));
  not1  g0251(.din(G972_o2), .dout(new_new_n799__));
  buf1  g0252(.din(G973_o2), .dout(new_new_n800__));
  not1  g0253(.din(G973_o2), .dout(new_new_n801__));
  buf1  g0254(.din(G977_o2), .dout(new_new_n802__));
  not1  g0255(.din(G977_o2), .dout(new_new_n803__));
  buf1  g0256(.din(G971_o2), .dout(new_new_n804__));
  not1  g0257(.din(G971_o2), .dout(new_new_n805__));
  buf1  g0258(.din(G975_o2), .dout(new_new_n806__));
  not1  g0259(.din(G975_o2), .dout(new_new_n807__));
  buf1  g0260(.din(G954_o2), .dout(new_new_n808__));
  not1  g0261(.din(G954_o2), .dout(new_new_n809__));
  buf1  g0262(.din(G956_o2), .dout(new_new_n810__));
  not1  g0263(.din(G956_o2), .dout(new_new_n811__));
  buf1  g0264(.din(G950_o2), .dout(new_new_n812__));
  not1  g0265(.din(G950_o2), .dout(new_new_n813__));
  buf1  g0266(.din(G952_o2), .dout(new_new_n814__));
  not1  g0267(.din(G952_o2), .dout(new_new_n815__));
  buf1  g0268(.din(G953_o2), .dout(new_new_n816__));
  not1  g0269(.din(G953_o2), .dout(new_new_n817__));
  buf1  g0270(.din(G957_o2), .dout(new_new_n818__));
  not1  g0271(.din(G957_o2), .dout(new_new_n819__));
  buf1  g0272(.din(G951_o2), .dout(new_new_n820__));
  not1  g0273(.din(G951_o2), .dout(new_new_n821__));
  buf1  g0274(.din(G955_o2), .dout(new_new_n822__));
  not1  g0275(.din(G955_o2), .dout(new_new_n823__));
  buf1  g0276(.din(G986_o2), .dout(new_new_n824__));
  not1  g0277(.din(G986_o2), .dout(new_new_n825__));
  buf1  g0278(.din(G991_o2), .dout(new_new_n826__));
  not1  g0279(.din(G991_o2), .dout(new_new_n827__));
  buf1  g0280(.din(G770_o2), .dout(new_new_n828__));
  not1  g0281(.din(G770_o2), .dout(new_new_n829__));
  buf1  g0282(.din(G773_o2), .dout(new_new_n830__));
  not1  g0283(.din(G773_o2), .dout(new_new_n831__));
  buf1  g0284(.din(G776_o2), .dout(new_new_n832__));
  not1  g0285(.din(G776_o2), .dout(new_new_n833__));
  buf1  g0286(.din(G779_o2), .dout(new_new_n834__));
  not1  g0287(.din(G779_o2), .dout(new_new_n835__));
  buf1  g0288(.din(G782_o2), .dout(new_new_n836__));
  not1  g0289(.din(G782_o2), .dout(new_new_n837__));
  buf1  g0290(.din(G785_o2), .dout(new_new_n838__));
  not1  g0291(.din(G785_o2), .dout(new_new_n839__));
  buf1  g0292(.din(G788_o2), .dout(new_new_n840__));
  not1  g0293(.din(G788_o2), .dout(new_new_n841__));
  buf1  g0294(.din(G791_o2), .dout(new_new_n842__));
  not1  g0295(.din(G791_o2), .dout(new_new_n843__));
  buf1  g0296(.din(G642_o2), .dout(new_new_n844__));
  not1  g0297(.din(G642_o2), .dout(new_new_n845__));
  buf1  g0298(.din(G645_o2), .dout(new_new_n846__));
  not1  g0299(.din(G645_o2), .dout(new_new_n847__));
  buf1  g0300(.din(G648_o2), .dout(new_new_n848__));
  not1  g0301(.din(G648_o2), .dout(new_new_n849__));
  buf1  g0302(.din(G651_o2), .dout(new_new_n850__));
  not1  g0303(.din(G651_o2), .dout(new_new_n851__));
  buf1  g0304(.din(G654_o2), .dout(new_new_n852__));
  not1  g0305(.din(G654_o2), .dout(new_new_n853__));
  buf1  g0306(.din(G657_o2), .dout(new_new_n854__));
  not1  g0307(.din(G657_o2), .dout(new_new_n855__));
  buf1  g0308(.din(G660_o2), .dout(new_new_n856__));
  not1  g0309(.din(G660_o2), .dout(new_new_n857__));
  buf1  g0310(.din(G663_o2), .dout(new_new_n858__));
  not1  g0311(.din(G663_o2), .dout(new_new_n859__));
  buf1  g0312(.din(G602_o2), .dout(new_new_n860__));
  not1  g0313(.din(G602_o2), .dout(new_new_n861__));
  buf1  g0314(.din(G607_o2), .dout(new_new_n862__));
  not1  g0315(.din(G607_o2), .dout(new_new_n863__));
  buf1  g0316(.din(G612_o2), .dout(new_new_n864__));
  not1  g0317(.din(G612_o2), .dout(new_new_n865__));
  buf1  g0318(.din(G617_o2), .dout(new_new_n866__));
  not1  g0319(.din(G617_o2), .dout(new_new_n867__));
  buf1  g0320(.din(G622_o2), .dout(new_new_n868__));
  not1  g0321(.din(G622_o2), .dout(new_new_n869__));
  buf1  g0322(.din(G627_o2), .dout(new_new_n870__));
  not1  g0323(.din(G627_o2), .dout(new_new_n871__));
  buf1  g0324(.din(G632_o2), .dout(new_new_n872__));
  not1  g0325(.din(G632_o2), .dout(new_new_n873__));
  buf1  g0326(.din(G637_o2), .dout(new_new_n874__));
  not1  g0327(.din(G637_o2), .dout(new_new_n875__));
  buf1  g0328(.din(n627_lo_buf_o2), .dout(new_new_n876__));
  not1  g0329(.din(n627_lo_buf_o2), .dout(new_new_n877__));
  buf1  g0330(.din(n639_lo_buf_o2), .dout(new_new_n878__));
  not1  g0331(.din(n639_lo_buf_o2), .dout(new_new_n879__));
  buf1  g0332(.din(n651_lo_buf_o2), .dout(new_new_n880__));
  not1  g0333(.din(n651_lo_buf_o2), .dout(new_new_n881__));
  buf1  g0334(.din(n663_lo_buf_o2), .dout(new_new_n882__));
  not1  g0335(.din(n663_lo_buf_o2), .dout(new_new_n883__));
  buf1  g0336(.din(n675_lo_buf_o2), .dout(new_new_n884__));
  not1  g0337(.din(n675_lo_buf_o2), .dout(new_new_n885__));
  buf1  g0338(.din(n687_lo_buf_o2), .dout(new_new_n886__));
  not1  g0339(.din(n687_lo_buf_o2), .dout(new_new_n887__));
  buf1  g0340(.din(n699_lo_buf_o2), .dout(new_new_n888__));
  not1  g0341(.din(n699_lo_buf_o2), .dout(new_new_n889__));
  buf1  g0342(.din(n711_lo_buf_o2), .dout(new_new_n890__));
  not1  g0343(.din(n711_lo_buf_o2), .dout(new_new_n891__));
  buf1  g0344(.din(n723_lo_buf_o2), .dout(new_new_n892__));
  not1  g0345(.din(n723_lo_buf_o2), .dout(new_new_n893__));
  buf1  g0346(.din(n735_lo_buf_o2), .dout(new_new_n894__));
  not1  g0347(.din(n735_lo_buf_o2), .dout(new_new_n895__));
  buf1  g0348(.din(n747_lo_buf_o2), .dout(new_new_n896__));
  not1  g0349(.din(n747_lo_buf_o2), .dout(new_new_n897__));
  buf1  g0350(.din(n759_lo_buf_o2), .dout(new_new_n898__));
  not1  g0351(.din(n759_lo_buf_o2), .dout(new_new_n899__));
  buf1  g0352(.din(n771_lo_buf_o2), .dout(new_new_n900__));
  not1  g0353(.din(n771_lo_buf_o2), .dout(new_new_n901__));
  buf1  g0354(.din(n783_lo_buf_o2), .dout(new_new_n902__));
  not1  g0355(.din(n783_lo_buf_o2), .dout(new_new_n903__));
  buf1  g0356(.din(n795_lo_buf_o2), .dout(new_new_n904__));
  not1  g0357(.din(n795_lo_buf_o2), .dout(new_new_n905__));
  buf1  g0358(.din(n807_lo_buf_o2), .dout(new_new_n906__));
  not1  g0359(.din(n807_lo_buf_o2), .dout(new_new_n907__));
  buf1  g0360(.din(n819_lo_buf_o2), .dout(new_new_n908__));
  not1  g0361(.din(n819_lo_buf_o2), .dout(new_new_n909__));
  buf1  g0362(.din(n831_lo_buf_o2), .dout(new_new_n910__));
  not1  g0363(.din(n831_lo_buf_o2), .dout(new_new_n911__));
  buf1  g0364(.din(n843_lo_buf_o2), .dout(new_new_n912__));
  not1  g0365(.din(n843_lo_buf_o2), .dout(new_new_n913__));
  buf1  g0366(.din(n855_lo_buf_o2), .dout(new_new_n914__));
  not1  g0367(.din(n855_lo_buf_o2), .dout(new_new_n915__));
  buf1  g0368(.din(n867_lo_buf_o2), .dout(new_new_n916__));
  not1  g0369(.din(n867_lo_buf_o2), .dout(new_new_n917__));
  buf1  g0370(.din(n879_lo_buf_o2), .dout(new_new_n918__));
  not1  g0371(.din(n879_lo_buf_o2), .dout(new_new_n919__));
  buf1  g0372(.din(n891_lo_buf_o2), .dout(new_new_n920__));
  not1  g0373(.din(n891_lo_buf_o2), .dout(new_new_n921__));
  buf1  g0374(.din(n903_lo_buf_o2), .dout(new_new_n922__));
  not1  g0375(.din(n903_lo_buf_o2), .dout(new_new_n923__));
  buf1  g0376(.din(n915_lo_buf_o2), .dout(new_new_n924__));
  not1  g0377(.din(n915_lo_buf_o2), .dout(new_new_n925__));
  buf1  g0378(.din(n927_lo_buf_o2), .dout(new_new_n926__));
  not1  g0379(.din(n927_lo_buf_o2), .dout(new_new_n927__));
  buf1  g0380(.din(n939_lo_buf_o2), .dout(new_new_n928__));
  not1  g0381(.din(n939_lo_buf_o2), .dout(new_new_n929__));
  buf1  g0382(.din(n951_lo_buf_o2), .dout(new_new_n930__));
  not1  g0383(.din(n951_lo_buf_o2), .dout(new_new_n931__));
  buf1  g0384(.din(n963_lo_buf_o2), .dout(new_new_n932__));
  not1  g0385(.din(n963_lo_buf_o2), .dout(new_new_n933__));
  buf1  g0386(.din(n975_lo_buf_o2), .dout(new_new_n934__));
  not1  g0387(.din(n975_lo_buf_o2), .dout(new_new_n935__));
  buf1  g0388(.din(n987_lo_buf_o2), .dout(new_new_n936__));
  not1  g0389(.din(n987_lo_buf_o2), .dout(new_new_n937__));
  buf1  g0390(.din(n999_lo_buf_o2), .dout(new_new_n938__));
  not1  g0391(.din(n999_lo_buf_o2), .dout(new_new_n939__));
  and1  g0392(.dina(new_new_n813__), .dinb(new_new_n1950__), .dout(new_new_n940__));
  or1   g0393(.dina(new_new_n812__), .dinb(new_new_n1955__), .dout(new_new_n941__));
  and1  g0394(.dina(new_new_n940__), .dinb(new_new_n1960__), .dout(new_new_n942__));
  or1   g0395(.dina(new_new_n941__), .dinb(new_new_n1965__), .dout(new_new_n943__));
  and1  g0396(.dina(new_new_n942__), .dinb(new_new_n821__), .dout(new_new_n944__));
  or1   g0397(.dina(new_new_n943__), .dinb(new_new_n820__), .dout(new_new_n945__));
  and1  g0398(.dina(new_new_n944__), .dinb(new_new_n1969__), .dout(new_new_n946__));
  or1   g0399(.dina(new_new_n945__), .dinb(new_new_n1972__), .dout(new_new_n947__));
  and1  g0400(.dina(new_new_n1975__), .dinb(new_new_n1979__), .dout(new_new_n948__));
  or1   g0401(.dina(new_new_n1983__), .dinb(new_new_n1987__), .dout(new_new_n949__));
  or1   g0402(.dina(new_new_n949__), .dinb(new_new_n549__), .dout(new_new_n950__));
  and1  g0403(.dina(new_new_n1990__), .dinb(new_new_n548__), .dout(new_new_n951__));
  and1  g0404(.dina(new_new_n1990__), .dinb(new_new_n948__), .dout(new_new_n952__));
  or1   g0405(.dina(new_new_n952__), .dinb(new_new_n951__), .dout(new_new_n953__));
  and1  g0406(.dina(new_new_n1975__), .dinb(new_new_n1993__), .dout(new_new_n954__));
  or1   g0407(.dina(new_new_n1983__), .dinb(new_new_n1998__), .dout(new_new_n955__));
  or1   g0408(.dina(new_new_n955__), .dinb(new_new_n551__), .dout(new_new_n956__));
  and1  g0409(.dina(new_new_n2001__), .dinb(new_new_n550__), .dout(new_new_n957__));
  and1  g0410(.dina(new_new_n2001__), .dinb(new_new_n954__), .dout(new_new_n958__));
  or1   g0411(.dina(new_new_n958__), .dinb(new_new_n957__), .dout(new_new_n959__));
  and1  g0412(.dina(new_new_n1976__), .dinb(new_new_n2004__), .dout(new_new_n960__));
  or1   g0413(.dina(new_new_n1984__), .dinb(new_new_n2009__), .dout(new_new_n961__));
  or1   g0414(.dina(new_new_n961__), .dinb(new_new_n553__), .dout(new_new_n962__));
  and1  g0415(.dina(new_new_n2012__), .dinb(new_new_n552__), .dout(new_new_n963__));
  and1  g0416(.dina(new_new_n2012__), .dinb(new_new_n960__), .dout(new_new_n964__));
  or1   g0417(.dina(new_new_n964__), .dinb(new_new_n963__), .dout(new_new_n965__));
  and1  g0418(.dina(new_new_n1976__), .dinb(new_new_n2015__), .dout(new_new_n966__));
  or1   g0419(.dina(new_new_n1984__), .dinb(new_new_n2020__), .dout(new_new_n967__));
  or1   g0420(.dina(new_new_n967__), .dinb(new_new_n555__), .dout(new_new_n968__));
  and1  g0421(.dina(new_new_n2023__), .dinb(new_new_n554__), .dout(new_new_n969__));
  and1  g0422(.dina(new_new_n2023__), .dinb(new_new_n966__), .dout(new_new_n970__));
  or1   g0423(.dina(new_new_n970__), .dinb(new_new_n969__), .dout(new_new_n971__));
  and1  g0424(.dina(new_new_n815__), .dinb(new_new_n1950__), .dout(new_new_n972__));
  or1   g0425(.dina(new_new_n814__), .dinb(new_new_n1955__), .dout(new_new_n973__));
  and1  g0426(.dina(new_new_n972__), .dinb(new_new_n817__), .dout(new_new_n974__));
  or1   g0427(.dina(new_new_n973__), .dinb(new_new_n816__), .dout(new_new_n975__));
  and1  g0428(.dina(new_new_n974__), .dinb(new_new_n2026__), .dout(new_new_n976__));
  or1   g0429(.dina(new_new_n975__), .dinb(new_new_n2031__), .dout(new_new_n977__));
  and1  g0430(.dina(new_new_n976__), .dinb(new_new_n1969__), .dout(new_new_n978__));
  or1   g0431(.dina(new_new_n977__), .dinb(new_new_n1972__), .dout(new_new_n979__));
  and1  g0432(.dina(new_new_n2035__), .dinb(new_new_n1979__), .dout(new_new_n980__));
  or1   g0433(.dina(new_new_n2038__), .dinb(new_new_n1987__), .dout(new_new_n981__));
  or1   g0434(.dina(new_new_n981__), .dinb(new_new_n557__), .dout(new_new_n982__));
  and1  g0435(.dina(new_new_n2040__), .dinb(new_new_n556__), .dout(new_new_n983__));
  and1  g0436(.dina(new_new_n2040__), .dinb(new_new_n980__), .dout(new_new_n984__));
  or1   g0437(.dina(new_new_n984__), .dinb(new_new_n983__), .dout(new_new_n985__));
  and1  g0438(.dina(new_new_n2035__), .dinb(new_new_n1993__), .dout(new_new_n986__));
  or1   g0439(.dina(new_new_n2038__), .dinb(new_new_n1998__), .dout(new_new_n987__));
  or1   g0440(.dina(new_new_n987__), .dinb(new_new_n559__), .dout(new_new_n988__));
  and1  g0441(.dina(new_new_n2041__), .dinb(new_new_n558__), .dout(new_new_n989__));
  and1  g0442(.dina(new_new_n2041__), .dinb(new_new_n986__), .dout(new_new_n990__));
  or1   g0443(.dina(new_new_n990__), .dinb(new_new_n989__), .dout(new_new_n991__));
  and1  g0444(.dina(new_new_n2036__), .dinb(new_new_n2004__), .dout(new_new_n992__));
  or1   g0445(.dina(new_new_n2039__), .dinb(new_new_n2009__), .dout(new_new_n993__));
  or1   g0446(.dina(new_new_n993__), .dinb(new_new_n561__), .dout(new_new_n994__));
  and1  g0447(.dina(new_new_n2042__), .dinb(new_new_n560__), .dout(new_new_n995__));
  and1  g0448(.dina(new_new_n2042__), .dinb(new_new_n992__), .dout(new_new_n996__));
  or1   g0449(.dina(new_new_n996__), .dinb(new_new_n995__), .dout(new_new_n997__));
  and1  g0450(.dina(new_new_n2036__), .dinb(new_new_n2015__), .dout(new_new_n998__));
  or1   g0451(.dina(new_new_n2039__), .dinb(new_new_n2020__), .dout(new_new_n999__));
  or1   g0452(.dina(new_new_n999__), .dinb(new_new_n563__), .dout(new_new_n1000__));
  and1  g0453(.dina(new_new_n2043__), .dinb(new_new_n562__), .dout(new_new_n1001__));
  and1  g0454(.dina(new_new_n2043__), .dinb(new_new_n998__), .dout(new_new_n1002__));
  or1   g0455(.dina(new_new_n1002__), .dinb(new_new_n1001__), .dout(new_new_n1003__));
  and1  g0456(.dina(new_new_n809__), .dinb(new_new_n2046__), .dout(new_new_n1004__));
  or1   g0457(.dina(new_new_n808__), .dinb(new_new_n2051__), .dout(new_new_n1005__));
  and1  g0458(.dina(new_new_n1004__), .dinb(new_new_n1960__), .dout(new_new_n1006__));
  or1   g0459(.dina(new_new_n1005__), .dinb(new_new_n1965__), .dout(new_new_n1007__));
  and1  g0460(.dina(new_new_n1006__), .dinb(new_new_n823__), .dout(new_new_n1008__));
  or1   g0461(.dina(new_new_n1007__), .dinb(new_new_n822__), .dout(new_new_n1009__));
  and1  g0462(.dina(new_new_n1008__), .dinb(new_new_n1970__), .dout(new_new_n1010__));
  or1   g0463(.dina(new_new_n1009__), .dinb(new_new_n1973__), .dout(new_new_n1011__));
  and1  g0464(.dina(new_new_n2055__), .dinb(new_new_n1980__), .dout(new_new_n1012__));
  or1   g0465(.dina(new_new_n2058__), .dinb(new_new_n1988__), .dout(new_new_n1013__));
  or1   g0466(.dina(new_new_n1013__), .dinb(new_new_n565__), .dout(new_new_n1014__));
  and1  g0467(.dina(new_new_n2060__), .dinb(new_new_n564__), .dout(new_new_n1015__));
  and1  g0468(.dina(new_new_n2060__), .dinb(new_new_n1012__), .dout(new_new_n1016__));
  or1   g0469(.dina(new_new_n1016__), .dinb(new_new_n1015__), .dout(new_new_n1017__));
  and1  g0470(.dina(new_new_n2055__), .dinb(new_new_n1994__), .dout(new_new_n1018__));
  or1   g0471(.dina(new_new_n2058__), .dinb(new_new_n1999__), .dout(new_new_n1019__));
  or1   g0472(.dina(new_new_n1019__), .dinb(new_new_n567__), .dout(new_new_n1020__));
  and1  g0473(.dina(new_new_n2061__), .dinb(new_new_n566__), .dout(new_new_n1021__));
  and1  g0474(.dina(new_new_n2061__), .dinb(new_new_n1018__), .dout(new_new_n1022__));
  or1   g0475(.dina(new_new_n1022__), .dinb(new_new_n1021__), .dout(new_new_n1023__));
  and1  g0476(.dina(new_new_n2056__), .dinb(new_new_n2005__), .dout(new_new_n1024__));
  or1   g0477(.dina(new_new_n2059__), .dinb(new_new_n2010__), .dout(new_new_n1025__));
  or1   g0478(.dina(new_new_n1025__), .dinb(new_new_n569__), .dout(new_new_n1026__));
  and1  g0479(.dina(new_new_n2062__), .dinb(new_new_n568__), .dout(new_new_n1027__));
  and1  g0480(.dina(new_new_n2062__), .dinb(new_new_n1024__), .dout(new_new_n1028__));
  or1   g0481(.dina(new_new_n1028__), .dinb(new_new_n1027__), .dout(new_new_n1029__));
  and1  g0482(.dina(new_new_n2056__), .dinb(new_new_n2016__), .dout(new_new_n1030__));
  or1   g0483(.dina(new_new_n2059__), .dinb(new_new_n2021__), .dout(new_new_n1031__));
  or1   g0484(.dina(new_new_n1031__), .dinb(new_new_n571__), .dout(new_new_n1032__));
  and1  g0485(.dina(new_new_n2063__), .dinb(new_new_n570__), .dout(new_new_n1033__));
  and1  g0486(.dina(new_new_n2063__), .dinb(new_new_n1030__), .dout(new_new_n1034__));
  or1   g0487(.dina(new_new_n1034__), .dinb(new_new_n1033__), .dout(new_new_n1035__));
  and1  g0488(.dina(new_new_n811__), .dinb(new_new_n2046__), .dout(new_new_n1036__));
  or1   g0489(.dina(new_new_n810__), .dinb(new_new_n2051__), .dout(new_new_n1037__));
  and1  g0490(.dina(new_new_n1036__), .dinb(new_new_n819__), .dout(new_new_n1038__));
  or1   g0491(.dina(new_new_n1037__), .dinb(new_new_n818__), .dout(new_new_n1039__));
  and1  g0492(.dina(new_new_n1038__), .dinb(new_new_n2026__), .dout(new_new_n1040__));
  or1   g0493(.dina(new_new_n1039__), .dinb(new_new_n2031__), .dout(new_new_n1041__));
  and1  g0494(.dina(new_new_n1040__), .dinb(new_new_n1970__), .dout(new_new_n1042__));
  or1   g0495(.dina(new_new_n1041__), .dinb(new_new_n1973__), .dout(new_new_n1043__));
  and1  g0496(.dina(new_new_n2065__), .dinb(new_new_n1980__), .dout(new_new_n1044__));
  or1   g0497(.dina(new_new_n2068__), .dinb(new_new_n1988__), .dout(new_new_n1045__));
  or1   g0498(.dina(new_new_n1045__), .dinb(new_new_n573__), .dout(new_new_n1046__));
  and1  g0499(.dina(new_new_n2070__), .dinb(new_new_n572__), .dout(new_new_n1047__));
  and1  g0500(.dina(new_new_n2070__), .dinb(new_new_n1044__), .dout(new_new_n1048__));
  or1   g0501(.dina(new_new_n1048__), .dinb(new_new_n1047__), .dout(new_new_n1049__));
  and1  g0502(.dina(new_new_n2065__), .dinb(new_new_n1994__), .dout(new_new_n1050__));
  or1   g0503(.dina(new_new_n2068__), .dinb(new_new_n1999__), .dout(new_new_n1051__));
  or1   g0504(.dina(new_new_n1051__), .dinb(new_new_n575__), .dout(new_new_n1052__));
  and1  g0505(.dina(new_new_n2071__), .dinb(new_new_n574__), .dout(new_new_n1053__));
  and1  g0506(.dina(new_new_n2071__), .dinb(new_new_n1050__), .dout(new_new_n1054__));
  or1   g0507(.dina(new_new_n1054__), .dinb(new_new_n1053__), .dout(new_new_n1055__));
  and1  g0508(.dina(new_new_n2066__), .dinb(new_new_n2005__), .dout(new_new_n1056__));
  or1   g0509(.dina(new_new_n2069__), .dinb(new_new_n2010__), .dout(new_new_n1057__));
  or1   g0510(.dina(new_new_n1057__), .dinb(new_new_n577__), .dout(new_new_n1058__));
  and1  g0511(.dina(new_new_n2072__), .dinb(new_new_n576__), .dout(new_new_n1059__));
  and1  g0512(.dina(new_new_n2072__), .dinb(new_new_n1056__), .dout(new_new_n1060__));
  or1   g0513(.dina(new_new_n1060__), .dinb(new_new_n1059__), .dout(new_new_n1061__));
  and1  g0514(.dina(new_new_n2066__), .dinb(new_new_n2016__), .dout(new_new_n1062__));
  or1   g0515(.dina(new_new_n2069__), .dinb(new_new_n2021__), .dout(new_new_n1063__));
  or1   g0516(.dina(new_new_n1063__), .dinb(new_new_n579__), .dout(new_new_n1064__));
  and1  g0517(.dina(new_new_n2073__), .dinb(new_new_n578__), .dout(new_new_n1065__));
  and1  g0518(.dina(new_new_n2073__), .dinb(new_new_n1062__), .dout(new_new_n1066__));
  or1   g0519(.dina(new_new_n1066__), .dinb(new_new_n1065__), .dout(new_new_n1067__));
  and1  g0520(.dina(new_new_n797__), .dinb(new_new_n1981__), .dout(new_new_n1068__));
  or1   g0521(.dina(new_new_n796__), .dinb(new_new_n1989__), .dout(new_new_n1069__));
  and1  g0522(.dina(new_new_n1068__), .dinb(new_new_n2006__), .dout(new_new_n1070__));
  or1   g0523(.dina(new_new_n1069__), .dinb(new_new_n2011__), .dout(new_new_n1071__));
  and1  g0524(.dina(new_new_n1070__), .dinb(new_new_n805__), .dout(new_new_n1072__));
  or1   g0525(.dina(new_new_n1071__), .dinb(new_new_n804__), .dout(new_new_n1073__));
  and1  g0526(.dina(new_new_n1072__), .dinb(new_new_n2075__), .dout(new_new_n1074__));
  or1   g0527(.dina(new_new_n1073__), .dinb(new_new_n2078__), .dout(new_new_n1075__));
  and1  g0528(.dina(new_new_n2081__), .dinb(new_new_n1951__), .dout(new_new_n1076__));
  or1   g0529(.dina(new_new_n2084__), .dinb(new_new_n1956__), .dout(new_new_n1077__));
  or1   g0530(.dina(new_new_n1077__), .dinb(new_new_n581__), .dout(new_new_n1078__));
  and1  g0531(.dina(new_new_n2086__), .dinb(new_new_n580__), .dout(new_new_n1079__));
  and1  g0532(.dina(new_new_n2086__), .dinb(new_new_n1076__), .dout(new_new_n1080__));
  or1   g0533(.dina(new_new_n1080__), .dinb(new_new_n1079__), .dout(new_new_n1081__));
  and1  g0534(.dina(new_new_n2081__), .dinb(new_new_n2047__), .dout(new_new_n1082__));
  or1   g0535(.dina(new_new_n2084__), .dinb(new_new_n2052__), .dout(new_new_n1083__));
  or1   g0536(.dina(new_new_n1083__), .dinb(new_new_n583__), .dout(new_new_n1084__));
  and1  g0537(.dina(new_new_n2087__), .dinb(new_new_n582__), .dout(new_new_n1085__));
  and1  g0538(.dina(new_new_n2087__), .dinb(new_new_n1082__), .dout(new_new_n1086__));
  or1   g0539(.dina(new_new_n1086__), .dinb(new_new_n1085__), .dout(new_new_n1087__));
  and1  g0540(.dina(new_new_n2082__), .dinb(new_new_n1961__), .dout(new_new_n1088__));
  or1   g0541(.dina(new_new_n2085__), .dinb(new_new_n1966__), .dout(new_new_n1089__));
  or1   g0542(.dina(new_new_n1089__), .dinb(new_new_n585__), .dout(new_new_n1090__));
  and1  g0543(.dina(new_new_n2088__), .dinb(new_new_n584__), .dout(new_new_n1091__));
  and1  g0544(.dina(new_new_n2088__), .dinb(new_new_n1088__), .dout(new_new_n1092__));
  or1   g0545(.dina(new_new_n1092__), .dinb(new_new_n1091__), .dout(new_new_n1093__));
  and1  g0546(.dina(new_new_n2082__), .dinb(new_new_n2027__), .dout(new_new_n1094__));
  or1   g0547(.dina(new_new_n2085__), .dinb(new_new_n2032__), .dout(new_new_n1095__));
  or1   g0548(.dina(new_new_n1095__), .dinb(new_new_n587__), .dout(new_new_n1096__));
  and1  g0549(.dina(new_new_n2089__), .dinb(new_new_n586__), .dout(new_new_n1097__));
  and1  g0550(.dina(new_new_n2089__), .dinb(new_new_n1094__), .dout(new_new_n1098__));
  or1   g0551(.dina(new_new_n1098__), .dinb(new_new_n1097__), .dout(new_new_n1099__));
  and1  g0552(.dina(new_new_n799__), .dinb(new_new_n1981__), .dout(new_new_n1100__));
  or1   g0553(.dina(new_new_n798__), .dinb(new_new_n1989__), .dout(new_new_n1101__));
  and1  g0554(.dina(new_new_n1100__), .dinb(new_new_n801__), .dout(new_new_n1102__));
  or1   g0555(.dina(new_new_n1101__), .dinb(new_new_n800__), .dout(new_new_n1103__));
  and1  g0556(.dina(new_new_n1102__), .dinb(new_new_n2017__), .dout(new_new_n1104__));
  or1   g0557(.dina(new_new_n1103__), .dinb(new_new_n2022__), .dout(new_new_n1105__));
  and1  g0558(.dina(new_new_n1104__), .dinb(new_new_n2075__), .dout(new_new_n1106__));
  or1   g0559(.dina(new_new_n1105__), .dinb(new_new_n2078__), .dout(new_new_n1107__));
  and1  g0560(.dina(new_new_n2091__), .dinb(new_new_n1951__), .dout(new_new_n1108__));
  or1   g0561(.dina(new_new_n2094__), .dinb(new_new_n1956__), .dout(new_new_n1109__));
  or1   g0562(.dina(new_new_n1109__), .dinb(new_new_n589__), .dout(new_new_n1110__));
  and1  g0563(.dina(new_new_n2096__), .dinb(new_new_n588__), .dout(new_new_n1111__));
  and1  g0564(.dina(new_new_n2096__), .dinb(new_new_n1108__), .dout(new_new_n1112__));
  or1   g0565(.dina(new_new_n1112__), .dinb(new_new_n1111__), .dout(new_new_n1113__));
  and1  g0566(.dina(new_new_n2091__), .dinb(new_new_n2047__), .dout(new_new_n1114__));
  or1   g0567(.dina(new_new_n2094__), .dinb(new_new_n2052__), .dout(new_new_n1115__));
  or1   g0568(.dina(new_new_n1115__), .dinb(new_new_n591__), .dout(new_new_n1116__));
  and1  g0569(.dina(new_new_n2097__), .dinb(new_new_n590__), .dout(new_new_n1117__));
  and1  g0570(.dina(new_new_n2097__), .dinb(new_new_n1114__), .dout(new_new_n1118__));
  or1   g0571(.dina(new_new_n1118__), .dinb(new_new_n1117__), .dout(new_new_n1119__));
  and1  g0572(.dina(new_new_n2092__), .dinb(new_new_n1961__), .dout(new_new_n1120__));
  or1   g0573(.dina(new_new_n2095__), .dinb(new_new_n1966__), .dout(new_new_n1121__));
  or1   g0574(.dina(new_new_n1121__), .dinb(new_new_n593__), .dout(new_new_n1122__));
  and1  g0575(.dina(new_new_n2098__), .dinb(new_new_n592__), .dout(new_new_n1123__));
  and1  g0576(.dina(new_new_n2098__), .dinb(new_new_n1120__), .dout(new_new_n1124__));
  or1   g0577(.dina(new_new_n1124__), .dinb(new_new_n1123__), .dout(new_new_n1125__));
  and1  g0578(.dina(new_new_n2092__), .dinb(new_new_n2027__), .dout(new_new_n1126__));
  or1   g0579(.dina(new_new_n2095__), .dinb(new_new_n2032__), .dout(new_new_n1127__));
  or1   g0580(.dina(new_new_n1127__), .dinb(new_new_n595__), .dout(new_new_n1128__));
  and1  g0581(.dina(new_new_n2099__), .dinb(new_new_n594__), .dout(new_new_n1129__));
  and1  g0582(.dina(new_new_n2099__), .dinb(new_new_n1126__), .dout(new_new_n1130__));
  or1   g0583(.dina(new_new_n1130__), .dinb(new_new_n1129__), .dout(new_new_n1131__));
  and1  g0584(.dina(new_new_n793__), .dinb(new_new_n1995__), .dout(new_new_n1132__));
  or1   g0585(.dina(new_new_n792__), .dinb(new_new_n2000__), .dout(new_new_n1133__));
  and1  g0586(.dina(new_new_n1132__), .dinb(new_new_n2006__), .dout(new_new_n1134__));
  or1   g0587(.dina(new_new_n1133__), .dinb(new_new_n2011__), .dout(new_new_n1135__));
  and1  g0588(.dina(new_new_n1134__), .dinb(new_new_n807__), .dout(new_new_n1136__));
  or1   g0589(.dina(new_new_n1135__), .dinb(new_new_n806__), .dout(new_new_n1137__));
  and1  g0590(.dina(new_new_n1136__), .dinb(new_new_n2076__), .dout(new_new_n1138__));
  or1   g0591(.dina(new_new_n1137__), .dinb(new_new_n2079__), .dout(new_new_n1139__));
  and1  g0592(.dina(new_new_n2101__), .dinb(new_new_n1952__), .dout(new_new_n1140__));
  or1   g0593(.dina(new_new_n2104__), .dinb(new_new_n1957__), .dout(new_new_n1141__));
  or1   g0594(.dina(new_new_n1141__), .dinb(new_new_n597__), .dout(new_new_n1142__));
  and1  g0595(.dina(new_new_n2106__), .dinb(new_new_n596__), .dout(new_new_n1143__));
  and1  g0596(.dina(new_new_n2106__), .dinb(new_new_n1140__), .dout(new_new_n1144__));
  or1   g0597(.dina(new_new_n1144__), .dinb(new_new_n1143__), .dout(new_new_n1145__));
  and1  g0598(.dina(new_new_n2101__), .dinb(new_new_n2048__), .dout(new_new_n1146__));
  or1   g0599(.dina(new_new_n2104__), .dinb(new_new_n2053__), .dout(new_new_n1147__));
  or1   g0600(.dina(new_new_n1147__), .dinb(new_new_n599__), .dout(new_new_n1148__));
  and1  g0601(.dina(new_new_n2107__), .dinb(new_new_n598__), .dout(new_new_n1149__));
  and1  g0602(.dina(new_new_n2107__), .dinb(new_new_n1146__), .dout(new_new_n1150__));
  or1   g0603(.dina(new_new_n1150__), .dinb(new_new_n1149__), .dout(new_new_n1151__));
  and1  g0604(.dina(new_new_n2102__), .dinb(new_new_n1962__), .dout(new_new_n1152__));
  or1   g0605(.dina(new_new_n2105__), .dinb(new_new_n1967__), .dout(new_new_n1153__));
  or1   g0606(.dina(new_new_n1153__), .dinb(new_new_n601__), .dout(new_new_n1154__));
  and1  g0607(.dina(new_new_n2108__), .dinb(new_new_n600__), .dout(new_new_n1155__));
  and1  g0608(.dina(new_new_n2108__), .dinb(new_new_n1152__), .dout(new_new_n1156__));
  or1   g0609(.dina(new_new_n1156__), .dinb(new_new_n1155__), .dout(new_new_n1157__));
  and1  g0610(.dina(new_new_n2102__), .dinb(new_new_n2028__), .dout(new_new_n1158__));
  or1   g0611(.dina(new_new_n2105__), .dinb(new_new_n2033__), .dout(new_new_n1159__));
  or1   g0612(.dina(new_new_n1159__), .dinb(new_new_n603__), .dout(new_new_n1160__));
  and1  g0613(.dina(new_new_n2109__), .dinb(new_new_n602__), .dout(new_new_n1161__));
  and1  g0614(.dina(new_new_n2109__), .dinb(new_new_n1158__), .dout(new_new_n1162__));
  or1   g0615(.dina(new_new_n1162__), .dinb(new_new_n1161__), .dout(new_new_n1163__));
  and1  g0616(.dina(new_new_n795__), .dinb(new_new_n1995__), .dout(new_new_n1164__));
  or1   g0617(.dina(new_new_n794__), .dinb(new_new_n2000__), .dout(new_new_n1165__));
  and1  g0618(.dina(new_new_n1164__), .dinb(new_new_n803__), .dout(new_new_n1166__));
  or1   g0619(.dina(new_new_n1165__), .dinb(new_new_n802__), .dout(new_new_n1167__));
  and1  g0620(.dina(new_new_n1166__), .dinb(new_new_n2017__), .dout(new_new_n1168__));
  or1   g0621(.dina(new_new_n1167__), .dinb(new_new_n2022__), .dout(new_new_n1169__));
  and1  g0622(.dina(new_new_n1168__), .dinb(new_new_n2076__), .dout(new_new_n1170__));
  or1   g0623(.dina(new_new_n1169__), .dinb(new_new_n2079__), .dout(new_new_n1171__));
  and1  g0624(.dina(new_new_n2111__), .dinb(new_new_n1952__), .dout(new_new_n1172__));
  or1   g0625(.dina(new_new_n2114__), .dinb(new_new_n1957__), .dout(new_new_n1173__));
  or1   g0626(.dina(new_new_n1173__), .dinb(new_new_n605__), .dout(new_new_n1174__));
  and1  g0627(.dina(new_new_n2116__), .dinb(new_new_n604__), .dout(new_new_n1175__));
  and1  g0628(.dina(new_new_n2116__), .dinb(new_new_n1172__), .dout(new_new_n1176__));
  or1   g0629(.dina(new_new_n1176__), .dinb(new_new_n1175__), .dout(new_new_n1177__));
  and1  g0630(.dina(new_new_n2111__), .dinb(new_new_n2048__), .dout(new_new_n1178__));
  or1   g0631(.dina(new_new_n2114__), .dinb(new_new_n2053__), .dout(new_new_n1179__));
  or1   g0632(.dina(new_new_n1179__), .dinb(new_new_n607__), .dout(new_new_n1180__));
  and1  g0633(.dina(new_new_n2117__), .dinb(new_new_n606__), .dout(new_new_n1181__));
  and1  g0634(.dina(new_new_n2117__), .dinb(new_new_n1178__), .dout(new_new_n1182__));
  or1   g0635(.dina(new_new_n1182__), .dinb(new_new_n1181__), .dout(new_new_n1183__));
  and1  g0636(.dina(new_new_n2112__), .dinb(new_new_n1962__), .dout(new_new_n1184__));
  or1   g0637(.dina(new_new_n2115__), .dinb(new_new_n1967__), .dout(new_new_n1185__));
  or1   g0638(.dina(new_new_n1185__), .dinb(new_new_n609__), .dout(new_new_n1186__));
  and1  g0639(.dina(new_new_n2118__), .dinb(new_new_n608__), .dout(new_new_n1187__));
  and1  g0640(.dina(new_new_n2118__), .dinb(new_new_n1184__), .dout(new_new_n1188__));
  or1   g0641(.dina(new_new_n1188__), .dinb(new_new_n1187__), .dout(new_new_n1189__));
  and1  g0642(.dina(new_new_n2112__), .dinb(new_new_n2028__), .dout(new_new_n1190__));
  or1   g0643(.dina(new_new_n2115__), .dinb(new_new_n2033__), .dout(new_new_n1191__));
  or1   g0644(.dina(new_new_n1191__), .dinb(new_new_n611__), .dout(new_new_n1192__));
  and1  g0645(.dina(new_new_n2119__), .dinb(new_new_n610__), .dout(new_new_n1193__));
  and1  g0646(.dina(new_new_n2119__), .dinb(new_new_n1190__), .dout(new_new_n1194__));
  or1   g0647(.dina(new_new_n1194__), .dinb(new_new_n1193__), .dout(new_new_n1195__));
  and1  g0648(.dina(new_new_n2120__), .dinb(new_new_n2121__), .dout(new_new_n1196__));
  or1   g0649(.dina(new_new_n2122__), .dinb(new_new_n2123__), .dout(new_new_n1197__));
  and1  g0650(.dina(new_new_n2124__), .dinb(new_new_n2120__), .dout(new_new_n1198__));
  or1   g0651(.dina(new_new_n2125__), .dinb(new_new_n2122__), .dout(new_new_n1199__));
  and1  g0652(.dina(new_new_n2124__), .dinb(new_new_n2121__), .dout(new_new_n1200__));
  or1   g0653(.dina(new_new_n2125__), .dinb(new_new_n2123__), .dout(new_new_n1201__));
  and1  g0654(.dina(new_new_n1201__), .dinb(new_new_n1199__), .dout(new_new_n1202__));
  or1   g0655(.dina(new_new_n1200__), .dinb(new_new_n1198__), .dout(new_new_n1203__));
  and1  g0656(.dina(new_new_n2126__), .dinb(new_new_n2127__), .dout(new_new_n1204__));
  or1   g0657(.dina(new_new_n2128__), .dinb(new_new_n2129__), .dout(new_new_n1205__));
  and1  g0658(.dina(new_new_n2130__), .dinb(new_new_n2126__), .dout(new_new_n1206__));
  or1   g0659(.dina(new_new_n2131__), .dinb(new_new_n2128__), .dout(new_new_n1207__));
  and1  g0660(.dina(new_new_n2130__), .dinb(new_new_n2127__), .dout(new_new_n1208__));
  or1   g0661(.dina(new_new_n2131__), .dinb(new_new_n2129__), .dout(new_new_n1209__));
  and1  g0662(.dina(new_new_n1209__), .dinb(new_new_n1207__), .dout(new_new_n1210__));
  or1   g0663(.dina(new_new_n1208__), .dinb(new_new_n1206__), .dout(new_new_n1211__));
  and1  g0664(.dina(new_new_n2132__), .dinb(new_new_n2133__), .dout(new_new_n1212__));
  or1   g0665(.dina(new_new_n2134__), .dinb(new_new_n2135__), .dout(new_new_n1213__));
  and1  g0666(.dina(new_new_n2136__), .dinb(new_new_n2132__), .dout(new_new_n1214__));
  or1   g0667(.dina(new_new_n2137__), .dinb(new_new_n2134__), .dout(new_new_n1215__));
  and1  g0668(.dina(new_new_n2136__), .dinb(new_new_n2133__), .dout(new_new_n1216__));
  or1   g0669(.dina(new_new_n2137__), .dinb(new_new_n2135__), .dout(new_new_n1217__));
  and1  g0670(.dina(new_new_n1217__), .dinb(new_new_n1215__), .dout(new_new_n1218__));
  or1   g0671(.dina(new_new_n1216__), .dinb(new_new_n1214__), .dout(new_new_n1219__));
  and1  g0672(.dina(new_new_n2138__), .dinb(new_new_n2139__), .dout(new_new_n1220__));
  or1   g0673(.dina(new_new_n2140__), .dinb(new_new_n2141__), .dout(new_new_n1221__));
  and1  g0674(.dina(new_new_n2142__), .dinb(new_new_n2138__), .dout(new_new_n1222__));
  or1   g0675(.dina(new_new_n2143__), .dinb(new_new_n2140__), .dout(new_new_n1223__));
  and1  g0676(.dina(new_new_n2142__), .dinb(new_new_n2139__), .dout(new_new_n1224__));
  or1   g0677(.dina(new_new_n2143__), .dinb(new_new_n2141__), .dout(new_new_n1225__));
  and1  g0678(.dina(new_new_n1225__), .dinb(new_new_n1223__), .dout(new_new_n1226__));
  or1   g0679(.dina(new_new_n1224__), .dinb(new_new_n1222__), .dout(new_new_n1227__));
  and1  g0680(.dina(new_new_n2144__), .dinb(new_new_n2145__), .dout(new_new_n1228__));
  or1   g0681(.dina(new_new_n2146__), .dinb(new_new_n2147__), .dout(new_new_n1229__));
  and1  g0682(.dina(new_new_n2148__), .dinb(new_new_n2144__), .dout(new_new_n1230__));
  or1   g0683(.dina(new_new_n2149__), .dinb(new_new_n2146__), .dout(new_new_n1231__));
  and1  g0684(.dina(new_new_n2148__), .dinb(new_new_n2145__), .dout(new_new_n1232__));
  or1   g0685(.dina(new_new_n2149__), .dinb(new_new_n2147__), .dout(new_new_n1233__));
  and1  g0686(.dina(new_new_n1233__), .dinb(new_new_n1231__), .dout(new_new_n1234__));
  or1   g0687(.dina(new_new_n1232__), .dinb(new_new_n1230__), .dout(new_new_n1235__));
  and1  g0688(.dina(new_new_n2150__), .dinb(new_new_n2151__), .dout(new_new_n1236__));
  or1   g0689(.dina(new_new_n2152__), .dinb(new_new_n2153__), .dout(new_new_n1237__));
  and1  g0690(.dina(new_new_n2154__), .dinb(new_new_n2150__), .dout(new_new_n1238__));
  or1   g0691(.dina(new_new_n2155__), .dinb(new_new_n2152__), .dout(new_new_n1239__));
  and1  g0692(.dina(new_new_n2154__), .dinb(new_new_n2151__), .dout(new_new_n1240__));
  or1   g0693(.dina(new_new_n2155__), .dinb(new_new_n2153__), .dout(new_new_n1241__));
  and1  g0694(.dina(new_new_n1241__), .dinb(new_new_n1239__), .dout(new_new_n1242__));
  or1   g0695(.dina(new_new_n1240__), .dinb(new_new_n1238__), .dout(new_new_n1243__));
  and1  g0696(.dina(new_new_n2156__), .dinb(new_new_n2157__), .dout(new_new_n1244__));
  or1   g0697(.dina(new_new_n2158__), .dinb(new_new_n2159__), .dout(new_new_n1245__));
  and1  g0698(.dina(new_new_n2160__), .dinb(new_new_n2156__), .dout(new_new_n1246__));
  or1   g0699(.dina(new_new_n2161__), .dinb(new_new_n2158__), .dout(new_new_n1247__));
  and1  g0700(.dina(new_new_n2160__), .dinb(new_new_n2157__), .dout(new_new_n1248__));
  or1   g0701(.dina(new_new_n2161__), .dinb(new_new_n2159__), .dout(new_new_n1249__));
  and1  g0702(.dina(new_new_n1249__), .dinb(new_new_n1247__), .dout(new_new_n1250__));
  or1   g0703(.dina(new_new_n1248__), .dinb(new_new_n1246__), .dout(new_new_n1251__));
  and1  g0704(.dina(new_new_n2162__), .dinb(new_new_n2163__), .dout(new_new_n1252__));
  or1   g0705(.dina(new_new_n2164__), .dinb(new_new_n2165__), .dout(new_new_n1253__));
  and1  g0706(.dina(new_new_n2166__), .dinb(new_new_n2162__), .dout(new_new_n1254__));
  or1   g0707(.dina(new_new_n2167__), .dinb(new_new_n2164__), .dout(new_new_n1255__));
  and1  g0708(.dina(new_new_n2166__), .dinb(new_new_n2163__), .dout(new_new_n1256__));
  or1   g0709(.dina(new_new_n2167__), .dinb(new_new_n2165__), .dout(new_new_n1257__));
  and1  g0710(.dina(new_new_n1257__), .dinb(new_new_n1255__), .dout(new_new_n1258__));
  or1   g0711(.dina(new_new_n1256__), .dinb(new_new_n1254__), .dout(new_new_n1259__));
  or1   g0712(.dina(new_new_n2168__), .dinb(new_new_n2169__), .dout(new_new_n1260__));
  or1   g0713(.dina(new_new_n2170__), .dinb(new_new_n2172__), .dout(new_new_n1261__));
  or1   g0714(.dina(new_new_n1261__), .dinb(new_new_n2174__), .dout(new_new_n1262__));
  or1   g0715(.dina(new_new_n2170__), .dinb(new_new_n2177__), .dout(new_new_n1263__));
  or1   g0716(.dina(new_new_n1263__), .dinb(new_new_n2180__), .dout(new_new_n1264__));
  or1   g0717(.dina(new_new_n2182__), .dinb(new_new_n2169__), .dout(new_new_n1265__));
  or1   g0718(.dina(new_new_n1265__), .dinb(new_new_n2172__), .dout(new_new_n1266__));
  or1   g0719(.dina(new_new_n1266__), .dinb(new_new_n2180__), .dout(new_new_n1267__));
  or1   g0720(.dina(new_new_n2168__), .dinb(new_new_n2185__), .dout(new_new_n1268__));
  or1   g0721(.dina(new_new_n1268__), .dinb(new_new_n2171__), .dout(new_new_n1269__));
  or1   g0722(.dina(new_new_n1269__), .dinb(new_new_n2179__), .dout(new_new_n1270__));
  and1  g0723(.dina(new_new_n1264__), .dinb(new_new_n1262__), .dout(new_new_n1271__));
  and1  g0724(.dina(new_new_n1271__), .dinb(new_new_n1267__), .dout(new_new_n1272__));
  and1  g0725(.dina(new_new_n1272__), .dinb(new_new_n1270__), .dout(new_new_n1273__));
  or1   g0726(.dina(new_new_n2187__), .dinb(new_new_n2188__), .dout(new_new_n1274__));
  or1   g0727(.dina(new_new_n2189__), .dinb(new_new_n2191__), .dout(new_new_n1275__));
  or1   g0728(.dina(new_new_n1275__), .dinb(new_new_n2193__), .dout(new_new_n1276__));
  or1   g0729(.dina(new_new_n2189__), .dinb(new_new_n2196__), .dout(new_new_n1277__));
  or1   g0730(.dina(new_new_n1277__), .dinb(new_new_n2199__), .dout(new_new_n1278__));
  or1   g0731(.dina(new_new_n2201__), .dinb(new_new_n2188__), .dout(new_new_n1279__));
  or1   g0732(.dina(new_new_n1279__), .dinb(new_new_n2191__), .dout(new_new_n1280__));
  or1   g0733(.dina(new_new_n1280__), .dinb(new_new_n2199__), .dout(new_new_n1281__));
  or1   g0734(.dina(new_new_n2187__), .dinb(new_new_n2204__), .dout(new_new_n1282__));
  or1   g0735(.dina(new_new_n1282__), .dinb(new_new_n2190__), .dout(new_new_n1283__));
  or1   g0736(.dina(new_new_n1283__), .dinb(new_new_n2198__), .dout(new_new_n1284__));
  and1  g0737(.dina(new_new_n1278__), .dinb(new_new_n1276__), .dout(new_new_n1285__));
  and1  g0738(.dina(new_new_n1285__), .dinb(new_new_n1281__), .dout(new_new_n1286__));
  and1  g0739(.dina(new_new_n1286__), .dinb(new_new_n1284__), .dout(new_new_n1287__));
  and1  g0740(.dina(new_new_n2208__), .dinb(new_new_n614__), .dout(new_new_n1288__));
  or1   g0741(.dina(new_new_n2215__), .dinb(new_new_n615__), .dout(new_new_n1289__));
  and1  g0742(.dina(new_new_n2221__), .dinb(new_new_n2224__), .dout(new_new_n1290__));
  or1   g0743(.dina(new_new_n2227__), .dinb(new_new_n2230__), .dout(new_new_n1291__));
  and1  g0744(.dina(new_new_n2232__), .dinb(new_new_n2224__), .dout(new_new_n1292__));
  or1   g0745(.dina(new_new_n2233__), .dinb(new_new_n2230__), .dout(new_new_n1293__));
  and1  g0746(.dina(new_new_n2232__), .dinb(new_new_n2221__), .dout(new_new_n1294__));
  or1   g0747(.dina(new_new_n2233__), .dinb(new_new_n2227__), .dout(new_new_n1295__));
  and1  g0748(.dina(new_new_n1295__), .dinb(new_new_n1293__), .dout(new_new_n1296__));
  or1   g0749(.dina(new_new_n1294__), .dinb(new_new_n1292__), .dout(new_new_n1297__));
  and1  g0750(.dina(new_new_n1297__), .dinb(new_new_n1288__), .dout(new_new_n1298__));
  or1   g0751(.dina(new_new_n2234__), .dinb(new_new_n1289__), .dout(new_new_n1299__));
  or1   g0752(.dina(new_new_n2234__), .dinb(new_new_n1296__), .dout(new_new_n1300__));
  and1  g0753(.dina(new_new_n1300__), .dinb(new_new_n1299__), .dout(new_new_n1301__));
  and1  g0754(.dina(new_new_n2208__), .dinb(new_new_n618__), .dout(new_new_n1302__));
  or1   g0755(.dina(new_new_n2215__), .dinb(new_new_n619__), .dout(new_new_n1303__));
  and1  g0756(.dina(new_new_n2236__), .dinb(new_new_n2239__), .dout(new_new_n1304__));
  or1   g0757(.dina(new_new_n2242__), .dinb(new_new_n2245__), .dout(new_new_n1305__));
  and1  g0758(.dina(new_new_n2247__), .dinb(new_new_n2239__), .dout(new_new_n1306__));
  or1   g0759(.dina(new_new_n2248__), .dinb(new_new_n2245__), .dout(new_new_n1307__));
  and1  g0760(.dina(new_new_n2247__), .dinb(new_new_n2236__), .dout(new_new_n1308__));
  or1   g0761(.dina(new_new_n2248__), .dinb(new_new_n2242__), .dout(new_new_n1309__));
  and1  g0762(.dina(new_new_n1309__), .dinb(new_new_n1307__), .dout(new_new_n1310__));
  or1   g0763(.dina(new_new_n1308__), .dinb(new_new_n1306__), .dout(new_new_n1311__));
  and1  g0764(.dina(new_new_n1311__), .dinb(new_new_n1302__), .dout(new_new_n1312__));
  or1   g0765(.dina(new_new_n2249__), .dinb(new_new_n1303__), .dout(new_new_n1313__));
  or1   g0766(.dina(new_new_n2249__), .dinb(new_new_n1310__), .dout(new_new_n1314__));
  and1  g0767(.dina(new_new_n1314__), .dinb(new_new_n1313__), .dout(new_new_n1315__));
  and1  g0768(.dina(new_new_n2209__), .dinb(new_new_n622__), .dout(new_new_n1316__));
  or1   g0769(.dina(new_new_n2216__), .dinb(new_new_n623__), .dout(new_new_n1317__));
  and1  g0770(.dina(new_new_n2240__), .dinb(new_new_n2225__), .dout(new_new_n1318__));
  or1   g0771(.dina(new_new_n2246__), .dinb(new_new_n2231__), .dout(new_new_n1319__));
  and1  g0772(.dina(new_new_n2250__), .dinb(new_new_n2225__), .dout(new_new_n1320__));
  or1   g0773(.dina(new_new_n2251__), .dinb(new_new_n2231__), .dout(new_new_n1321__));
  and1  g0774(.dina(new_new_n2250__), .dinb(new_new_n2240__), .dout(new_new_n1322__));
  or1   g0775(.dina(new_new_n2251__), .dinb(new_new_n2246__), .dout(new_new_n1323__));
  and1  g0776(.dina(new_new_n1323__), .dinb(new_new_n1321__), .dout(new_new_n1324__));
  or1   g0777(.dina(new_new_n1322__), .dinb(new_new_n1320__), .dout(new_new_n1325__));
  and1  g0778(.dina(new_new_n1325__), .dinb(new_new_n1316__), .dout(new_new_n1326__));
  or1   g0779(.dina(new_new_n2252__), .dinb(new_new_n1317__), .dout(new_new_n1327__));
  or1   g0780(.dina(new_new_n2252__), .dinb(new_new_n1324__), .dout(new_new_n1328__));
  and1  g0781(.dina(new_new_n1328__), .dinb(new_new_n1327__), .dout(new_new_n1329__));
  and1  g0782(.dina(new_new_n2209__), .dinb(new_new_n626__), .dout(new_new_n1330__));
  or1   g0783(.dina(new_new_n2216__), .dinb(new_new_n627__), .dout(new_new_n1331__));
  and1  g0784(.dina(new_new_n2237__), .dinb(new_new_n2222__), .dout(new_new_n1332__));
  or1   g0785(.dina(new_new_n2243__), .dinb(new_new_n2228__), .dout(new_new_n1333__));
  and1  g0786(.dina(new_new_n2253__), .dinb(new_new_n2222__), .dout(new_new_n1334__));
  or1   g0787(.dina(new_new_n2254__), .dinb(new_new_n2228__), .dout(new_new_n1335__));
  and1  g0788(.dina(new_new_n2253__), .dinb(new_new_n2237__), .dout(new_new_n1336__));
  or1   g0789(.dina(new_new_n2254__), .dinb(new_new_n2243__), .dout(new_new_n1337__));
  and1  g0790(.dina(new_new_n1337__), .dinb(new_new_n1335__), .dout(new_new_n1338__));
  or1   g0791(.dina(new_new_n1336__), .dinb(new_new_n1334__), .dout(new_new_n1339__));
  and1  g0792(.dina(new_new_n1339__), .dinb(new_new_n1330__), .dout(new_new_n1340__));
  or1   g0793(.dina(new_new_n2255__), .dinb(new_new_n1331__), .dout(new_new_n1341__));
  or1   g0794(.dina(new_new_n2255__), .dinb(new_new_n1338__), .dout(new_new_n1342__));
  and1  g0795(.dina(new_new_n1342__), .dinb(new_new_n1341__), .dout(new_new_n1343__));
  and1  g0796(.dina(new_new_n2211__), .dinb(new_new_n630__), .dout(new_new_n1344__));
  or1   g0797(.dina(new_new_n2218__), .dinb(new_new_n631__), .dout(new_new_n1345__));
  and1  g0798(.dina(new_new_n2257__), .dinb(new_new_n2260__), .dout(new_new_n1346__));
  or1   g0799(.dina(new_new_n2263__), .dinb(new_new_n2266__), .dout(new_new_n1347__));
  and1  g0800(.dina(new_new_n2268__), .dinb(new_new_n2260__), .dout(new_new_n1348__));
  or1   g0801(.dina(new_new_n2269__), .dinb(new_new_n2266__), .dout(new_new_n1349__));
  and1  g0802(.dina(new_new_n2268__), .dinb(new_new_n2257__), .dout(new_new_n1350__));
  or1   g0803(.dina(new_new_n2269__), .dinb(new_new_n2263__), .dout(new_new_n1351__));
  and1  g0804(.dina(new_new_n1351__), .dinb(new_new_n1349__), .dout(new_new_n1352__));
  or1   g0805(.dina(new_new_n1350__), .dinb(new_new_n1348__), .dout(new_new_n1353__));
  and1  g0806(.dina(new_new_n1353__), .dinb(new_new_n1344__), .dout(new_new_n1354__));
  or1   g0807(.dina(new_new_n2270__), .dinb(new_new_n1345__), .dout(new_new_n1355__));
  or1   g0808(.dina(new_new_n2270__), .dinb(new_new_n1352__), .dout(new_new_n1356__));
  and1  g0809(.dina(new_new_n1356__), .dinb(new_new_n1355__), .dout(new_new_n1357__));
  and1  g0810(.dina(new_new_n2211__), .dinb(new_new_n634__), .dout(new_new_n1358__));
  or1   g0811(.dina(new_new_n2218__), .dinb(new_new_n635__), .dout(new_new_n1359__));
  and1  g0812(.dina(new_new_n2272__), .dinb(new_new_n2275__), .dout(new_new_n1360__));
  or1   g0813(.dina(new_new_n2278__), .dinb(new_new_n2281__), .dout(new_new_n1361__));
  and1  g0814(.dina(new_new_n2283__), .dinb(new_new_n2275__), .dout(new_new_n1362__));
  or1   g0815(.dina(new_new_n2284__), .dinb(new_new_n2281__), .dout(new_new_n1363__));
  and1  g0816(.dina(new_new_n2283__), .dinb(new_new_n2272__), .dout(new_new_n1364__));
  or1   g0817(.dina(new_new_n2284__), .dinb(new_new_n2278__), .dout(new_new_n1365__));
  and1  g0818(.dina(new_new_n1365__), .dinb(new_new_n1363__), .dout(new_new_n1366__));
  or1   g0819(.dina(new_new_n1364__), .dinb(new_new_n1362__), .dout(new_new_n1367__));
  and1  g0820(.dina(new_new_n1367__), .dinb(new_new_n1358__), .dout(new_new_n1368__));
  or1   g0821(.dina(new_new_n2285__), .dinb(new_new_n1359__), .dout(new_new_n1369__));
  or1   g0822(.dina(new_new_n2285__), .dinb(new_new_n1366__), .dout(new_new_n1370__));
  and1  g0823(.dina(new_new_n1370__), .dinb(new_new_n1369__), .dout(new_new_n1371__));
  and1  g0824(.dina(new_new_n2212__), .dinb(new_new_n638__), .dout(new_new_n1372__));
  or1   g0825(.dina(new_new_n2219__), .dinb(new_new_n639__), .dout(new_new_n1373__));
  and1  g0826(.dina(new_new_n2276__), .dinb(new_new_n2261__), .dout(new_new_n1374__));
  or1   g0827(.dina(new_new_n2282__), .dinb(new_new_n2267__), .dout(new_new_n1375__));
  and1  g0828(.dina(new_new_n2286__), .dinb(new_new_n2261__), .dout(new_new_n1376__));
  or1   g0829(.dina(new_new_n2287__), .dinb(new_new_n2267__), .dout(new_new_n1377__));
  and1  g0830(.dina(new_new_n2286__), .dinb(new_new_n2276__), .dout(new_new_n1378__));
  or1   g0831(.dina(new_new_n2287__), .dinb(new_new_n2282__), .dout(new_new_n1379__));
  and1  g0832(.dina(new_new_n1379__), .dinb(new_new_n1377__), .dout(new_new_n1380__));
  or1   g0833(.dina(new_new_n1378__), .dinb(new_new_n1376__), .dout(new_new_n1381__));
  and1  g0834(.dina(new_new_n1381__), .dinb(new_new_n1372__), .dout(new_new_n1382__));
  or1   g0835(.dina(new_new_n2288__), .dinb(new_new_n1373__), .dout(new_new_n1383__));
  or1   g0836(.dina(new_new_n2288__), .dinb(new_new_n1380__), .dout(new_new_n1384__));
  and1  g0837(.dina(new_new_n1384__), .dinb(new_new_n1383__), .dout(new_new_n1385__));
  and1  g0838(.dina(new_new_n2212__), .dinb(new_new_n642__), .dout(new_new_n1386__));
  or1   g0839(.dina(new_new_n2219__), .dinb(new_new_n643__), .dout(new_new_n1387__));
  and1  g0840(.dina(new_new_n2273__), .dinb(new_new_n2258__), .dout(new_new_n1388__));
  or1   g0841(.dina(new_new_n2279__), .dinb(new_new_n2264__), .dout(new_new_n1389__));
  and1  g0842(.dina(new_new_n2289__), .dinb(new_new_n2258__), .dout(new_new_n1390__));
  or1   g0843(.dina(new_new_n2290__), .dinb(new_new_n2264__), .dout(new_new_n1391__));
  and1  g0844(.dina(new_new_n2289__), .dinb(new_new_n2273__), .dout(new_new_n1392__));
  or1   g0845(.dina(new_new_n2290__), .dinb(new_new_n2279__), .dout(new_new_n1393__));
  and1  g0846(.dina(new_new_n1393__), .dinb(new_new_n1391__), .dout(new_new_n1394__));
  or1   g0847(.dina(new_new_n1392__), .dinb(new_new_n1390__), .dout(new_new_n1395__));
  and1  g0848(.dina(new_new_n1395__), .dinb(new_new_n1386__), .dout(new_new_n1396__));
  or1   g0849(.dina(new_new_n2291__), .dinb(new_new_n1387__), .dout(new_new_n1397__));
  or1   g0850(.dina(new_new_n2291__), .dinb(new_new_n1394__), .dout(new_new_n1398__));
  and1  g0851(.dina(new_new_n1398__), .dinb(new_new_n1397__), .dout(new_new_n1399__));
  and1  g0852(.dina(new_new_n2292__), .dinb(new_new_n2293__), .dout(new_new_n1400__));
  or1   g0853(.dina(new_new_n2295__), .dinb(new_new_n2297__), .dout(new_new_n1401__));
  and1  g0854(.dina(new_new_n2298__), .dinb(new_new_n2293__), .dout(new_new_n1402__));
  or1   g0855(.dina(new_new_n2299__), .dinb(new_new_n2297__), .dout(new_new_n1403__));
  and1  g0856(.dina(new_new_n2298__), .dinb(new_new_n2292__), .dout(new_new_n1404__));
  or1   g0857(.dina(new_new_n2299__), .dinb(new_new_n2295__), .dout(new_new_n1405__));
  and1  g0858(.dina(new_new_n1405__), .dinb(new_new_n1403__), .dout(new_new_n1406__));
  or1   g0859(.dina(new_new_n1404__), .dinb(new_new_n1402__), .dout(new_new_n1407__));
  and1  g0860(.dina(new_new_n2300__), .dinb(new_new_n2301__), .dout(new_new_n1408__));
  or1   g0861(.dina(new_new_n2303__), .dinb(new_new_n2305__), .dout(new_new_n1409__));
  and1  g0862(.dina(new_new_n2306__), .dinb(new_new_n2301__), .dout(new_new_n1410__));
  or1   g0863(.dina(new_new_n2307__), .dinb(new_new_n2305__), .dout(new_new_n1411__));
  and1  g0864(.dina(new_new_n2306__), .dinb(new_new_n2300__), .dout(new_new_n1412__));
  or1   g0865(.dina(new_new_n2307__), .dinb(new_new_n2303__), .dout(new_new_n1413__));
  and1  g0866(.dina(new_new_n1413__), .dinb(new_new_n1411__), .dout(new_new_n1414__));
  or1   g0867(.dina(new_new_n1412__), .dinb(new_new_n1410__), .dout(new_new_n1415__));
  and1  g0868(.dina(new_new_n1415__), .dinb(new_new_n1407__), .dout(new_new_n1416__));
  or1   g0869(.dina(new_new_n2308__), .dinb(new_new_n1406__), .dout(new_new_n1417__));
  or1   g0870(.dina(new_new_n2308__), .dinb(new_new_n1414__), .dout(new_new_n1418__));
  and1  g0871(.dina(new_new_n1418__), .dinb(new_new_n1417__), .dout(new_new_n1419__));
  and1  g0872(.dina(new_new_n2309__), .dinb(new_new_n2310__), .dout(new_new_n1420__));
  or1   g0873(.dina(new_new_n2312__), .dinb(new_new_n2314__), .dout(new_new_n1421__));
  and1  g0874(.dina(new_new_n2315__), .dinb(new_new_n2310__), .dout(new_new_n1422__));
  or1   g0875(.dina(new_new_n2316__), .dinb(new_new_n2314__), .dout(new_new_n1423__));
  and1  g0876(.dina(new_new_n2315__), .dinb(new_new_n2309__), .dout(new_new_n1424__));
  or1   g0877(.dina(new_new_n2316__), .dinb(new_new_n2312__), .dout(new_new_n1425__));
  and1  g0878(.dina(new_new_n1425__), .dinb(new_new_n1423__), .dout(new_new_n1426__));
  or1   g0879(.dina(new_new_n1424__), .dinb(new_new_n1422__), .dout(new_new_n1427__));
  and1  g0880(.dina(new_new_n2317__), .dinb(new_new_n2318__), .dout(new_new_n1428__));
  or1   g0881(.dina(new_new_n2320__), .dinb(new_new_n2322__), .dout(new_new_n1429__));
  and1  g0882(.dina(new_new_n2323__), .dinb(new_new_n2318__), .dout(new_new_n1430__));
  or1   g0883(.dina(new_new_n2324__), .dinb(new_new_n2322__), .dout(new_new_n1431__));
  and1  g0884(.dina(new_new_n2323__), .dinb(new_new_n2317__), .dout(new_new_n1432__));
  or1   g0885(.dina(new_new_n2324__), .dinb(new_new_n2320__), .dout(new_new_n1433__));
  and1  g0886(.dina(new_new_n1433__), .dinb(new_new_n1431__), .dout(new_new_n1434__));
  or1   g0887(.dina(new_new_n1432__), .dinb(new_new_n1430__), .dout(new_new_n1435__));
  and1  g0888(.dina(new_new_n1435__), .dinb(new_new_n1427__), .dout(new_new_n1436__));
  or1   g0889(.dina(new_new_n2325__), .dinb(new_new_n1426__), .dout(new_new_n1437__));
  or1   g0890(.dina(new_new_n2325__), .dinb(new_new_n1434__), .dout(new_new_n1438__));
  and1  g0891(.dina(new_new_n1438__), .dinb(new_new_n1437__), .dout(new_new_n1439__));
  and1  g0892(.dina(new_new_n2326__), .dinb(new_new_n2327__), .dout(new_new_n1440__));
  or1   g0893(.dina(new_new_n2329__), .dinb(new_new_n2331__), .dout(new_new_n1441__));
  and1  g0894(.dina(new_new_n2332__), .dinb(new_new_n2327__), .dout(new_new_n1442__));
  or1   g0895(.dina(new_new_n2333__), .dinb(new_new_n2331__), .dout(new_new_n1443__));
  and1  g0896(.dina(new_new_n2332__), .dinb(new_new_n2326__), .dout(new_new_n1444__));
  or1   g0897(.dina(new_new_n2333__), .dinb(new_new_n2329__), .dout(new_new_n1445__));
  and1  g0898(.dina(new_new_n1445__), .dinb(new_new_n1443__), .dout(new_new_n1446__));
  or1   g0899(.dina(new_new_n1444__), .dinb(new_new_n1442__), .dout(new_new_n1447__));
  and1  g0900(.dina(new_new_n2334__), .dinb(new_new_n2335__), .dout(new_new_n1448__));
  or1   g0901(.dina(new_new_n2337__), .dinb(new_new_n2339__), .dout(new_new_n1449__));
  and1  g0902(.dina(new_new_n2340__), .dinb(new_new_n2335__), .dout(new_new_n1450__));
  or1   g0903(.dina(new_new_n2341__), .dinb(new_new_n2339__), .dout(new_new_n1451__));
  and1  g0904(.dina(new_new_n2340__), .dinb(new_new_n2334__), .dout(new_new_n1452__));
  or1   g0905(.dina(new_new_n2341__), .dinb(new_new_n2337__), .dout(new_new_n1453__));
  and1  g0906(.dina(new_new_n1453__), .dinb(new_new_n1451__), .dout(new_new_n1454__));
  or1   g0907(.dina(new_new_n1452__), .dinb(new_new_n1450__), .dout(new_new_n1455__));
  and1  g0908(.dina(new_new_n1455__), .dinb(new_new_n1447__), .dout(new_new_n1456__));
  or1   g0909(.dina(new_new_n2342__), .dinb(new_new_n1446__), .dout(new_new_n1457__));
  or1   g0910(.dina(new_new_n2342__), .dinb(new_new_n1454__), .dout(new_new_n1458__));
  and1  g0911(.dina(new_new_n1458__), .dinb(new_new_n1457__), .dout(new_new_n1459__));
  and1  g0912(.dina(new_new_n2343__), .dinb(new_new_n2344__), .dout(new_new_n1460__));
  or1   g0913(.dina(new_new_n2346__), .dinb(new_new_n2348__), .dout(new_new_n1461__));
  and1  g0914(.dina(new_new_n2349__), .dinb(new_new_n2344__), .dout(new_new_n1462__));
  or1   g0915(.dina(new_new_n2350__), .dinb(new_new_n2348__), .dout(new_new_n1463__));
  and1  g0916(.dina(new_new_n2349__), .dinb(new_new_n2343__), .dout(new_new_n1464__));
  or1   g0917(.dina(new_new_n2350__), .dinb(new_new_n2346__), .dout(new_new_n1465__));
  and1  g0918(.dina(new_new_n1465__), .dinb(new_new_n1463__), .dout(new_new_n1466__));
  or1   g0919(.dina(new_new_n1464__), .dinb(new_new_n1462__), .dout(new_new_n1467__));
  and1  g0920(.dina(new_new_n2351__), .dinb(new_new_n2352__), .dout(new_new_n1468__));
  or1   g0921(.dina(new_new_n2354__), .dinb(new_new_n2356__), .dout(new_new_n1469__));
  and1  g0922(.dina(new_new_n2357__), .dinb(new_new_n2352__), .dout(new_new_n1470__));
  or1   g0923(.dina(new_new_n2358__), .dinb(new_new_n2356__), .dout(new_new_n1471__));
  and1  g0924(.dina(new_new_n2357__), .dinb(new_new_n2351__), .dout(new_new_n1472__));
  or1   g0925(.dina(new_new_n2358__), .dinb(new_new_n2354__), .dout(new_new_n1473__));
  and1  g0926(.dina(new_new_n1473__), .dinb(new_new_n1471__), .dout(new_new_n1474__));
  or1   g0927(.dina(new_new_n1472__), .dinb(new_new_n1470__), .dout(new_new_n1475__));
  and1  g0928(.dina(new_new_n1475__), .dinb(new_new_n1467__), .dout(new_new_n1476__));
  or1   g0929(.dina(new_new_n2359__), .dinb(new_new_n1466__), .dout(new_new_n1477__));
  or1   g0930(.dina(new_new_n2359__), .dinb(new_new_n1474__), .dout(new_new_n1478__));
  and1  g0931(.dina(new_new_n1478__), .dinb(new_new_n1477__), .dout(new_new_n1479__));
  and1  g0932(.dina(new_new_n2360__), .dinb(new_new_n2361__), .dout(new_new_n1480__));
  or1   g0933(.dina(new_new_n2363__), .dinb(new_new_n2365__), .dout(new_new_n1481__));
  and1  g0934(.dina(new_new_n2366__), .dinb(new_new_n2361__), .dout(new_new_n1482__));
  or1   g0935(.dina(new_new_n2367__), .dinb(new_new_n2365__), .dout(new_new_n1483__));
  and1  g0936(.dina(new_new_n2366__), .dinb(new_new_n2360__), .dout(new_new_n1484__));
  or1   g0937(.dina(new_new_n2367__), .dinb(new_new_n2363__), .dout(new_new_n1485__));
  and1  g0938(.dina(new_new_n1485__), .dinb(new_new_n1483__), .dout(new_new_n1486__));
  or1   g0939(.dina(new_new_n1484__), .dinb(new_new_n1482__), .dout(new_new_n1487__));
  and1  g0940(.dina(new_new_n2368__), .dinb(new_new_n2369__), .dout(new_new_n1488__));
  or1   g0941(.dina(new_new_n2371__), .dinb(new_new_n2373__), .dout(new_new_n1489__));
  and1  g0942(.dina(new_new_n2374__), .dinb(new_new_n2369__), .dout(new_new_n1490__));
  or1   g0943(.dina(new_new_n2375__), .dinb(new_new_n2373__), .dout(new_new_n1491__));
  and1  g0944(.dina(new_new_n2374__), .dinb(new_new_n2368__), .dout(new_new_n1492__));
  or1   g0945(.dina(new_new_n2375__), .dinb(new_new_n2371__), .dout(new_new_n1493__));
  and1  g0946(.dina(new_new_n1493__), .dinb(new_new_n1491__), .dout(new_new_n1494__));
  or1   g0947(.dina(new_new_n1492__), .dinb(new_new_n1490__), .dout(new_new_n1495__));
  and1  g0948(.dina(new_new_n1495__), .dinb(new_new_n1487__), .dout(new_new_n1496__));
  or1   g0949(.dina(new_new_n2376__), .dinb(new_new_n1486__), .dout(new_new_n1497__));
  or1   g0950(.dina(new_new_n2376__), .dinb(new_new_n1494__), .dout(new_new_n1498__));
  and1  g0951(.dina(new_new_n1498__), .dinb(new_new_n1497__), .dout(new_new_n1499__));
  and1  g0952(.dina(new_new_n2377__), .dinb(new_new_n2378__), .dout(new_new_n1500__));
  or1   g0953(.dina(new_new_n2380__), .dinb(new_new_n2382__), .dout(new_new_n1501__));
  and1  g0954(.dina(new_new_n2383__), .dinb(new_new_n2378__), .dout(new_new_n1502__));
  or1   g0955(.dina(new_new_n2384__), .dinb(new_new_n2382__), .dout(new_new_n1503__));
  and1  g0956(.dina(new_new_n2383__), .dinb(new_new_n2377__), .dout(new_new_n1504__));
  or1   g0957(.dina(new_new_n2384__), .dinb(new_new_n2380__), .dout(new_new_n1505__));
  and1  g0958(.dina(new_new_n1505__), .dinb(new_new_n1503__), .dout(new_new_n1506__));
  or1   g0959(.dina(new_new_n1504__), .dinb(new_new_n1502__), .dout(new_new_n1507__));
  and1  g0960(.dina(new_new_n2385__), .dinb(new_new_n2386__), .dout(new_new_n1508__));
  or1   g0961(.dina(new_new_n2388__), .dinb(new_new_n2390__), .dout(new_new_n1509__));
  and1  g0962(.dina(new_new_n2391__), .dinb(new_new_n2386__), .dout(new_new_n1510__));
  or1   g0963(.dina(new_new_n2392__), .dinb(new_new_n2390__), .dout(new_new_n1511__));
  and1  g0964(.dina(new_new_n2391__), .dinb(new_new_n2385__), .dout(new_new_n1512__));
  or1   g0965(.dina(new_new_n2392__), .dinb(new_new_n2388__), .dout(new_new_n1513__));
  and1  g0966(.dina(new_new_n1513__), .dinb(new_new_n1511__), .dout(new_new_n1514__));
  or1   g0967(.dina(new_new_n1512__), .dinb(new_new_n1510__), .dout(new_new_n1515__));
  and1  g0968(.dina(new_new_n1515__), .dinb(new_new_n1507__), .dout(new_new_n1516__));
  or1   g0969(.dina(new_new_n2393__), .dinb(new_new_n1506__), .dout(new_new_n1517__));
  or1   g0970(.dina(new_new_n2393__), .dinb(new_new_n1514__), .dout(new_new_n1518__));
  and1  g0971(.dina(new_new_n1518__), .dinb(new_new_n1517__), .dout(new_new_n1519__));
  and1  g0972(.dina(new_new_n2394__), .dinb(new_new_n2395__), .dout(new_new_n1520__));
  or1   g0973(.dina(new_new_n2397__), .dinb(new_new_n2399__), .dout(new_new_n1521__));
  and1  g0974(.dina(new_new_n2400__), .dinb(new_new_n2395__), .dout(new_new_n1522__));
  or1   g0975(.dina(new_new_n2401__), .dinb(new_new_n2399__), .dout(new_new_n1523__));
  and1  g0976(.dina(new_new_n2400__), .dinb(new_new_n2394__), .dout(new_new_n1524__));
  or1   g0977(.dina(new_new_n2401__), .dinb(new_new_n2397__), .dout(new_new_n1525__));
  and1  g0978(.dina(new_new_n1525__), .dinb(new_new_n1523__), .dout(new_new_n1526__));
  or1   g0979(.dina(new_new_n1524__), .dinb(new_new_n1522__), .dout(new_new_n1527__));
  and1  g0980(.dina(new_new_n2402__), .dinb(new_new_n2403__), .dout(new_new_n1528__));
  or1   g0981(.dina(new_new_n2405__), .dinb(new_new_n2407__), .dout(new_new_n1529__));
  and1  g0982(.dina(new_new_n2408__), .dinb(new_new_n2403__), .dout(new_new_n1530__));
  or1   g0983(.dina(new_new_n2409__), .dinb(new_new_n2407__), .dout(new_new_n1531__));
  and1  g0984(.dina(new_new_n2408__), .dinb(new_new_n2402__), .dout(new_new_n1532__));
  or1   g0985(.dina(new_new_n2409__), .dinb(new_new_n2405__), .dout(new_new_n1533__));
  and1  g0986(.dina(new_new_n1533__), .dinb(new_new_n1531__), .dout(new_new_n1534__));
  or1   g0987(.dina(new_new_n1532__), .dinb(new_new_n1530__), .dout(new_new_n1535__));
  and1  g0988(.dina(new_new_n1535__), .dinb(new_new_n1527__), .dout(new_new_n1536__));
  or1   g0989(.dina(new_new_n2410__), .dinb(new_new_n1526__), .dout(new_new_n1537__));
  or1   g0990(.dina(new_new_n2410__), .dinb(new_new_n1534__), .dout(new_new_n1538__));
  and1  g0991(.dina(new_new_n1538__), .dinb(new_new_n1537__), .dout(new_new_n1539__));
  and1  g0992(.dina(new_new_n2411__), .dinb(new_new_n2412__), .dout(new_new_n1540__));
  or1   g0993(.dina(new_new_n2414__), .dinb(new_new_n2416__), .dout(new_new_n1541__));
  and1  g0994(.dina(new_new_n2417__), .dinb(new_new_n2412__), .dout(new_new_n1542__));
  or1   g0995(.dina(new_new_n2418__), .dinb(new_new_n2416__), .dout(new_new_n1543__));
  and1  g0996(.dina(new_new_n2417__), .dinb(new_new_n2411__), .dout(new_new_n1544__));
  or1   g0997(.dina(new_new_n2418__), .dinb(new_new_n2414__), .dout(new_new_n1545__));
  and1  g0998(.dina(new_new_n1545__), .dinb(new_new_n1543__), .dout(new_new_n1546__));
  or1   g0999(.dina(new_new_n1544__), .dinb(new_new_n1542__), .dout(new_new_n1547__));
  and1  g1000(.dina(new_new_n2419__), .dinb(new_new_n2420__), .dout(new_new_n1548__));
  or1   g1001(.dina(new_new_n2422__), .dinb(new_new_n2424__), .dout(new_new_n1549__));
  and1  g1002(.dina(new_new_n2425__), .dinb(new_new_n2420__), .dout(new_new_n1550__));
  or1   g1003(.dina(new_new_n2426__), .dinb(new_new_n2424__), .dout(new_new_n1551__));
  and1  g1004(.dina(new_new_n2425__), .dinb(new_new_n2419__), .dout(new_new_n1552__));
  or1   g1005(.dina(new_new_n2426__), .dinb(new_new_n2422__), .dout(new_new_n1553__));
  and1  g1006(.dina(new_new_n1553__), .dinb(new_new_n1551__), .dout(new_new_n1554__));
  or1   g1007(.dina(new_new_n1552__), .dinb(new_new_n1550__), .dout(new_new_n1555__));
  and1  g1008(.dina(new_new_n1555__), .dinb(new_new_n1547__), .dout(new_new_n1556__));
  or1   g1009(.dina(new_new_n2427__), .dinb(new_new_n1546__), .dout(new_new_n1557__));
  or1   g1010(.dina(new_new_n2427__), .dinb(new_new_n1554__), .dout(new_new_n1558__));
  and1  g1011(.dina(new_new_n1558__), .dinb(new_new_n1557__), .dout(new_new_n1559__));
  and1  g1012(.dina(new_new_n2428__), .dinb(new_new_n2429__), .dout(new_new_n1560__));
  or1   g1013(.dina(new_new_n2431__), .dinb(new_new_n2433__), .dout(new_new_n1561__));
  and1  g1014(.dina(new_new_n2434__), .dinb(new_new_n2429__), .dout(new_new_n1562__));
  or1   g1015(.dina(new_new_n2435__), .dinb(new_new_n2433__), .dout(new_new_n1563__));
  and1  g1016(.dina(new_new_n2434__), .dinb(new_new_n2428__), .dout(new_new_n1564__));
  or1   g1017(.dina(new_new_n2435__), .dinb(new_new_n2431__), .dout(new_new_n1565__));
  and1  g1018(.dina(new_new_n1565__), .dinb(new_new_n1563__), .dout(new_new_n1566__));
  or1   g1019(.dina(new_new_n1564__), .dinb(new_new_n1562__), .dout(new_new_n1567__));
  and1  g1020(.dina(new_new_n2436__), .dinb(new_new_n2437__), .dout(new_new_n1568__));
  or1   g1021(.dina(new_new_n2439__), .dinb(new_new_n2441__), .dout(new_new_n1569__));
  and1  g1022(.dina(new_new_n2442__), .dinb(new_new_n2437__), .dout(new_new_n1570__));
  or1   g1023(.dina(new_new_n2443__), .dinb(new_new_n2441__), .dout(new_new_n1571__));
  and1  g1024(.dina(new_new_n2442__), .dinb(new_new_n2436__), .dout(new_new_n1572__));
  or1   g1025(.dina(new_new_n2443__), .dinb(new_new_n2439__), .dout(new_new_n1573__));
  and1  g1026(.dina(new_new_n1573__), .dinb(new_new_n1571__), .dout(new_new_n1574__));
  or1   g1027(.dina(new_new_n1572__), .dinb(new_new_n1570__), .dout(new_new_n1575__));
  and1  g1028(.dina(new_new_n1575__), .dinb(new_new_n1567__), .dout(new_new_n1576__));
  or1   g1029(.dina(new_new_n2444__), .dinb(new_new_n1566__), .dout(new_new_n1577__));
  or1   g1030(.dina(new_new_n2444__), .dinb(new_new_n1574__), .dout(new_new_n1578__));
  and1  g1031(.dina(new_new_n1578__), .dinb(new_new_n1577__), .dout(new_new_n1579__));
  and1  g1032(.dina(new_new_n2445__), .dinb(new_new_n2446__), .dout(new_new_n1580__));
  or1   g1033(.dina(new_new_n2448__), .dinb(new_new_n2450__), .dout(new_new_n1581__));
  and1  g1034(.dina(new_new_n2451__), .dinb(new_new_n2446__), .dout(new_new_n1582__));
  or1   g1035(.dina(new_new_n2452__), .dinb(new_new_n2450__), .dout(new_new_n1583__));
  and1  g1036(.dina(new_new_n2451__), .dinb(new_new_n2445__), .dout(new_new_n1584__));
  or1   g1037(.dina(new_new_n2452__), .dinb(new_new_n2448__), .dout(new_new_n1585__));
  and1  g1038(.dina(new_new_n1585__), .dinb(new_new_n1583__), .dout(new_new_n1586__));
  or1   g1039(.dina(new_new_n1584__), .dinb(new_new_n1582__), .dout(new_new_n1587__));
  and1  g1040(.dina(new_new_n2453__), .dinb(new_new_n2454__), .dout(new_new_n1588__));
  or1   g1041(.dina(new_new_n2456__), .dinb(new_new_n2458__), .dout(new_new_n1589__));
  and1  g1042(.dina(new_new_n2459__), .dinb(new_new_n2454__), .dout(new_new_n1590__));
  or1   g1043(.dina(new_new_n2460__), .dinb(new_new_n2458__), .dout(new_new_n1591__));
  and1  g1044(.dina(new_new_n2459__), .dinb(new_new_n2453__), .dout(new_new_n1592__));
  or1   g1045(.dina(new_new_n2460__), .dinb(new_new_n2456__), .dout(new_new_n1593__));
  and1  g1046(.dina(new_new_n1593__), .dinb(new_new_n1591__), .dout(new_new_n1594__));
  or1   g1047(.dina(new_new_n1592__), .dinb(new_new_n1590__), .dout(new_new_n1595__));
  and1  g1048(.dina(new_new_n1595__), .dinb(new_new_n1587__), .dout(new_new_n1596__));
  or1   g1049(.dina(new_new_n2461__), .dinb(new_new_n1586__), .dout(new_new_n1597__));
  or1   g1050(.dina(new_new_n2461__), .dinb(new_new_n1594__), .dout(new_new_n1598__));
  and1  g1051(.dina(new_new_n1598__), .dinb(new_new_n1597__), .dout(new_new_n1599__));
  and1  g1052(.dina(new_new_n2462__), .dinb(new_new_n2463__), .dout(new_new_n1600__));
  or1   g1053(.dina(new_new_n2465__), .dinb(new_new_n2467__), .dout(new_new_n1601__));
  and1  g1054(.dina(new_new_n2468__), .dinb(new_new_n2463__), .dout(new_new_n1602__));
  or1   g1055(.dina(new_new_n2469__), .dinb(new_new_n2467__), .dout(new_new_n1603__));
  and1  g1056(.dina(new_new_n2468__), .dinb(new_new_n2462__), .dout(new_new_n1604__));
  or1   g1057(.dina(new_new_n2469__), .dinb(new_new_n2465__), .dout(new_new_n1605__));
  and1  g1058(.dina(new_new_n1605__), .dinb(new_new_n1603__), .dout(new_new_n1606__));
  or1   g1059(.dina(new_new_n1604__), .dinb(new_new_n1602__), .dout(new_new_n1607__));
  and1  g1060(.dina(new_new_n2470__), .dinb(new_new_n2471__), .dout(new_new_n1608__));
  or1   g1061(.dina(new_new_n2473__), .dinb(new_new_n2475__), .dout(new_new_n1609__));
  and1  g1062(.dina(new_new_n2476__), .dinb(new_new_n2471__), .dout(new_new_n1610__));
  or1   g1063(.dina(new_new_n2477__), .dinb(new_new_n2475__), .dout(new_new_n1611__));
  and1  g1064(.dina(new_new_n2476__), .dinb(new_new_n2470__), .dout(new_new_n1612__));
  or1   g1065(.dina(new_new_n2477__), .dinb(new_new_n2473__), .dout(new_new_n1613__));
  and1  g1066(.dina(new_new_n1613__), .dinb(new_new_n1611__), .dout(new_new_n1614__));
  or1   g1067(.dina(new_new_n1612__), .dinb(new_new_n1610__), .dout(new_new_n1615__));
  and1  g1068(.dina(new_new_n1615__), .dinb(new_new_n1607__), .dout(new_new_n1616__));
  or1   g1069(.dina(new_new_n2478__), .dinb(new_new_n1606__), .dout(new_new_n1617__));
  or1   g1070(.dina(new_new_n2478__), .dinb(new_new_n1614__), .dout(new_new_n1618__));
  and1  g1071(.dina(new_new_n1618__), .dinb(new_new_n1617__), .dout(new_new_n1619__));
  and1  g1072(.dina(new_new_n2479__), .dinb(new_new_n2480__), .dout(new_new_n1620__));
  or1   g1073(.dina(new_new_n2482__), .dinb(new_new_n2484__), .dout(new_new_n1621__));
  and1  g1074(.dina(new_new_n2485__), .dinb(new_new_n2480__), .dout(new_new_n1622__));
  or1   g1075(.dina(new_new_n2486__), .dinb(new_new_n2484__), .dout(new_new_n1623__));
  and1  g1076(.dina(new_new_n2485__), .dinb(new_new_n2479__), .dout(new_new_n1624__));
  or1   g1077(.dina(new_new_n2486__), .dinb(new_new_n2482__), .dout(new_new_n1625__));
  and1  g1078(.dina(new_new_n1625__), .dinb(new_new_n1623__), .dout(new_new_n1626__));
  or1   g1079(.dina(new_new_n1624__), .dinb(new_new_n1622__), .dout(new_new_n1627__));
  and1  g1080(.dina(new_new_n2487__), .dinb(new_new_n2488__), .dout(new_new_n1628__));
  or1   g1081(.dina(new_new_n2490__), .dinb(new_new_n2492__), .dout(new_new_n1629__));
  and1  g1082(.dina(new_new_n2493__), .dinb(new_new_n2488__), .dout(new_new_n1630__));
  or1   g1083(.dina(new_new_n2494__), .dinb(new_new_n2492__), .dout(new_new_n1631__));
  and1  g1084(.dina(new_new_n2493__), .dinb(new_new_n2487__), .dout(new_new_n1632__));
  or1   g1085(.dina(new_new_n2494__), .dinb(new_new_n2490__), .dout(new_new_n1633__));
  and1  g1086(.dina(new_new_n1633__), .dinb(new_new_n1631__), .dout(new_new_n1634__));
  or1   g1087(.dina(new_new_n1632__), .dinb(new_new_n1630__), .dout(new_new_n1635__));
  and1  g1088(.dina(new_new_n1635__), .dinb(new_new_n1627__), .dout(new_new_n1636__));
  or1   g1089(.dina(new_new_n2495__), .dinb(new_new_n1626__), .dout(new_new_n1637__));
  or1   g1090(.dina(new_new_n2495__), .dinb(new_new_n1634__), .dout(new_new_n1638__));
  and1  g1091(.dina(new_new_n1638__), .dinb(new_new_n1637__), .dout(new_new_n1639__));
  and1  g1092(.dina(new_new_n2496__), .dinb(new_new_n2497__), .dout(new_new_n1640__));
  or1   g1093(.dina(new_new_n2499__), .dinb(new_new_n2501__), .dout(new_new_n1641__));
  and1  g1094(.dina(new_new_n2502__), .dinb(new_new_n2497__), .dout(new_new_n1642__));
  or1   g1095(.dina(new_new_n2503__), .dinb(new_new_n2501__), .dout(new_new_n1643__));
  and1  g1096(.dina(new_new_n2502__), .dinb(new_new_n2496__), .dout(new_new_n1644__));
  or1   g1097(.dina(new_new_n2503__), .dinb(new_new_n2499__), .dout(new_new_n1645__));
  and1  g1098(.dina(new_new_n1645__), .dinb(new_new_n1643__), .dout(new_new_n1646__));
  or1   g1099(.dina(new_new_n1644__), .dinb(new_new_n1642__), .dout(new_new_n1647__));
  and1  g1100(.dina(new_new_n2504__), .dinb(new_new_n2505__), .dout(new_new_n1648__));
  or1   g1101(.dina(new_new_n2507__), .dinb(new_new_n2509__), .dout(new_new_n1649__));
  and1  g1102(.dina(new_new_n2510__), .dinb(new_new_n2505__), .dout(new_new_n1650__));
  or1   g1103(.dina(new_new_n2511__), .dinb(new_new_n2509__), .dout(new_new_n1651__));
  and1  g1104(.dina(new_new_n2510__), .dinb(new_new_n2504__), .dout(new_new_n1652__));
  or1   g1105(.dina(new_new_n2511__), .dinb(new_new_n2507__), .dout(new_new_n1653__));
  and1  g1106(.dina(new_new_n1653__), .dinb(new_new_n1651__), .dout(new_new_n1654__));
  or1   g1107(.dina(new_new_n1652__), .dinb(new_new_n1650__), .dout(new_new_n1655__));
  and1  g1108(.dina(new_new_n1655__), .dinb(new_new_n1647__), .dout(new_new_n1656__));
  or1   g1109(.dina(new_new_n2512__), .dinb(new_new_n1646__), .dout(new_new_n1657__));
  or1   g1110(.dina(new_new_n2512__), .dinb(new_new_n1654__), .dout(new_new_n1658__));
  and1  g1111(.dina(new_new_n1658__), .dinb(new_new_n1657__), .dout(new_new_n1659__));
  and1  g1112(.dina(new_new_n2513__), .dinb(new_new_n2514__), .dout(new_new_n1660__));
  or1   g1113(.dina(new_new_n2516__), .dinb(new_new_n2518__), .dout(new_new_n1661__));
  and1  g1114(.dina(new_new_n2519__), .dinb(new_new_n2514__), .dout(new_new_n1662__));
  or1   g1115(.dina(new_new_n2520__), .dinb(new_new_n2518__), .dout(new_new_n1663__));
  and1  g1116(.dina(new_new_n2519__), .dinb(new_new_n2513__), .dout(new_new_n1664__));
  or1   g1117(.dina(new_new_n2520__), .dinb(new_new_n2516__), .dout(new_new_n1665__));
  and1  g1118(.dina(new_new_n1665__), .dinb(new_new_n1663__), .dout(new_new_n1666__));
  or1   g1119(.dina(new_new_n1664__), .dinb(new_new_n1662__), .dout(new_new_n1667__));
  and1  g1120(.dina(new_new_n2521__), .dinb(new_new_n2522__), .dout(new_new_n1668__));
  or1   g1121(.dina(new_new_n2524__), .dinb(new_new_n2526__), .dout(new_new_n1669__));
  and1  g1122(.dina(new_new_n2527__), .dinb(new_new_n2522__), .dout(new_new_n1670__));
  or1   g1123(.dina(new_new_n2528__), .dinb(new_new_n2526__), .dout(new_new_n1671__));
  and1  g1124(.dina(new_new_n2527__), .dinb(new_new_n2521__), .dout(new_new_n1672__));
  or1   g1125(.dina(new_new_n2528__), .dinb(new_new_n2524__), .dout(new_new_n1673__));
  and1  g1126(.dina(new_new_n1673__), .dinb(new_new_n1671__), .dout(new_new_n1674__));
  or1   g1127(.dina(new_new_n1672__), .dinb(new_new_n1670__), .dout(new_new_n1675__));
  and1  g1128(.dina(new_new_n1675__), .dinb(new_new_n1667__), .dout(new_new_n1676__));
  or1   g1129(.dina(new_new_n2529__), .dinb(new_new_n1666__), .dout(new_new_n1677__));
  or1   g1130(.dina(new_new_n2529__), .dinb(new_new_n1674__), .dout(new_new_n1678__));
  and1  g1131(.dina(new_new_n1678__), .dinb(new_new_n1677__), .dout(new_new_n1679__));
  and1  g1132(.dina(new_new_n2530__), .dinb(new_new_n2531__), .dout(new_new_n1680__));
  or1   g1133(.dina(new_new_n2533__), .dinb(new_new_n2535__), .dout(new_new_n1681__));
  and1  g1134(.dina(new_new_n2536__), .dinb(new_new_n2531__), .dout(new_new_n1682__));
  or1   g1135(.dina(new_new_n2537__), .dinb(new_new_n2535__), .dout(new_new_n1683__));
  and1  g1136(.dina(new_new_n2536__), .dinb(new_new_n2530__), .dout(new_new_n1684__));
  or1   g1137(.dina(new_new_n2537__), .dinb(new_new_n2533__), .dout(new_new_n1685__));
  and1  g1138(.dina(new_new_n1685__), .dinb(new_new_n1683__), .dout(new_new_n1686__));
  or1   g1139(.dina(new_new_n1684__), .dinb(new_new_n1682__), .dout(new_new_n1687__));
  and1  g1140(.dina(new_new_n2538__), .dinb(new_new_n2539__), .dout(new_new_n1688__));
  or1   g1141(.dina(new_new_n2541__), .dinb(new_new_n2543__), .dout(new_new_n1689__));
  and1  g1142(.dina(new_new_n2544__), .dinb(new_new_n2539__), .dout(new_new_n1690__));
  or1   g1143(.dina(new_new_n2545__), .dinb(new_new_n2543__), .dout(new_new_n1691__));
  and1  g1144(.dina(new_new_n2544__), .dinb(new_new_n2538__), .dout(new_new_n1692__));
  or1   g1145(.dina(new_new_n2545__), .dinb(new_new_n2541__), .dout(new_new_n1693__));
  and1  g1146(.dina(new_new_n1693__), .dinb(new_new_n1691__), .dout(new_new_n1694__));
  or1   g1147(.dina(new_new_n1692__), .dinb(new_new_n1690__), .dout(new_new_n1695__));
  and1  g1148(.dina(new_new_n1695__), .dinb(new_new_n1687__), .dout(new_new_n1696__));
  or1   g1149(.dina(new_new_n2546__), .dinb(new_new_n1686__), .dout(new_new_n1697__));
  or1   g1150(.dina(new_new_n2546__), .dinb(new_new_n1694__), .dout(new_new_n1698__));
  and1  g1151(.dina(new_new_n1698__), .dinb(new_new_n1697__), .dout(new_new_n1699__));
  and1  g1152(.dina(new_new_n2547__), .dinb(new_new_n2548__), .dout(new_new_n1700__));
  or1   g1153(.dina(new_new_n2550__), .dinb(new_new_n2552__), .dout(new_new_n1701__));
  and1  g1154(.dina(new_new_n2553__), .dinb(new_new_n2548__), .dout(new_new_n1702__));
  or1   g1155(.dina(new_new_n2554__), .dinb(new_new_n2552__), .dout(new_new_n1703__));
  and1  g1156(.dina(new_new_n2553__), .dinb(new_new_n2547__), .dout(new_new_n1704__));
  or1   g1157(.dina(new_new_n2554__), .dinb(new_new_n2550__), .dout(new_new_n1705__));
  and1  g1158(.dina(new_new_n1705__), .dinb(new_new_n1703__), .dout(new_new_n1706__));
  or1   g1159(.dina(new_new_n1704__), .dinb(new_new_n1702__), .dout(new_new_n1707__));
  and1  g1160(.dina(new_new_n2555__), .dinb(new_new_n2556__), .dout(new_new_n1708__));
  or1   g1161(.dina(new_new_n2558__), .dinb(new_new_n2560__), .dout(new_new_n1709__));
  and1  g1162(.dina(new_new_n2561__), .dinb(new_new_n2556__), .dout(new_new_n1710__));
  or1   g1163(.dina(new_new_n2562__), .dinb(new_new_n2560__), .dout(new_new_n1711__));
  and1  g1164(.dina(new_new_n2561__), .dinb(new_new_n2555__), .dout(new_new_n1712__));
  or1   g1165(.dina(new_new_n2562__), .dinb(new_new_n2558__), .dout(new_new_n1713__));
  and1  g1166(.dina(new_new_n1713__), .dinb(new_new_n1711__), .dout(new_new_n1714__));
  or1   g1167(.dina(new_new_n1712__), .dinb(new_new_n1710__), .dout(new_new_n1715__));
  and1  g1168(.dina(new_new_n1715__), .dinb(new_new_n1707__), .dout(new_new_n1716__));
  or1   g1169(.dina(new_new_n2563__), .dinb(new_new_n1706__), .dout(new_new_n1717__));
  or1   g1170(.dina(new_new_n2563__), .dinb(new_new_n1714__), .dout(new_new_n1718__));
  and1  g1171(.dina(new_new_n1718__), .dinb(new_new_n1717__), .dout(new_new_n1719__));
  not1  g1172(.din(new_new_n953__), .dout(G1324));
  not1  g1173(.din(new_new_n959__), .dout(G1325));
  not1  g1174(.din(new_new_n965__), .dout(G1326));
  not1  g1175(.din(new_new_n971__), .dout(G1327));
  not1  g1176(.din(new_new_n985__), .dout(G1328));
  not1  g1177(.din(new_new_n991__), .dout(G1329));
  not1  g1178(.din(new_new_n997__), .dout(G1330));
  not1  g1179(.din(new_new_n1003__), .dout(G1331));
  not1  g1180(.din(new_new_n1017__), .dout(G1332));
  not1  g1181(.din(new_new_n1023__), .dout(G1333));
  not1  g1182(.din(new_new_n1029__), .dout(G1334));
  not1  g1183(.din(new_new_n1035__), .dout(G1335));
  not1  g1184(.din(new_new_n1049__), .dout(G1336));
  not1  g1185(.din(new_new_n1055__), .dout(G1337));
  not1  g1186(.din(new_new_n1061__), .dout(G1338));
  not1  g1187(.din(new_new_n1067__), .dout(G1339));
  not1  g1188(.din(new_new_n1081__), .dout(G1340));
  not1  g1189(.din(new_new_n1087__), .dout(G1341));
  not1  g1190(.din(new_new_n1093__), .dout(G1342));
  not1  g1191(.din(new_new_n1099__), .dout(G1343));
  not1  g1192(.din(new_new_n1113__), .dout(G1344));
  not1  g1193(.din(new_new_n1119__), .dout(G1345));
  not1  g1194(.din(new_new_n1125__), .dout(G1346));
  not1  g1195(.din(new_new_n1131__), .dout(G1347));
  not1  g1196(.din(new_new_n1145__), .dout(G1348));
  not1  g1197(.din(new_new_n1151__), .dout(G1349));
  not1  g1198(.din(new_new_n1157__), .dout(G1350));
  not1  g1199(.din(new_new_n1163__), .dout(G1351));
  not1  g1200(.din(new_new_n1177__), .dout(G1352));
  not1  g1201(.din(new_new_n1183__), .dout(G1353));
  not1  g1202(.din(new_new_n1189__), .dout(G1354));
  not1  g1203(.din(new_new_n1195__), .dout(G1355));
  not1  g1204(.din(new_new_n649__), .dout(n4343));
  not1  g1205(.din(new_new_n651__), .dout(n4346));
  not1  g1206(.din(new_new_n653__), .dout(n4349));
  not1  g1207(.din(new_new_n655__), .dout(n4352));
  not1  g1208(.din(new_new_n657__), .dout(n4355));
  not1  g1209(.din(new_new_n659__), .dout(n4358));
  not1  g1210(.din(new_new_n661__), .dout(n4361));
  not1  g1211(.din(new_new_n663__), .dout(n4364));
  not1  g1212(.din(new_new_n665__), .dout(n4367));
  not1  g1213(.din(new_new_n667__), .dout(n4370));
  not1  g1214(.din(new_new_n669__), .dout(n4373));
  not1  g1215(.din(new_new_n671__), .dout(n4376));
  not1  g1216(.din(new_new_n673__), .dout(n4379));
  not1  g1217(.din(new_new_n675__), .dout(n4382));
  not1  g1218(.din(new_new_n677__), .dout(n4385));
  not1  g1219(.din(new_new_n679__), .dout(n4388));
  not1  g1220(.din(new_new_n681__), .dout(n4391));
  not1  g1221(.din(new_new_n683__), .dout(n4394));
  not1  g1222(.din(new_new_n685__), .dout(n4397));
  not1  g1223(.din(new_new_n687__), .dout(n4400));
  not1  g1224(.din(new_new_n689__), .dout(n4403));
  not1  g1225(.din(new_new_n691__), .dout(n4406));
  not1  g1226(.din(new_new_n693__), .dout(n4409));
  not1  g1227(.din(new_new_n695__), .dout(n4412));
  not1  g1228(.din(new_new_n697__), .dout(n4415));
  not1  g1229(.din(new_new_n699__), .dout(n4418));
  not1  g1230(.din(new_new_n701__), .dout(n4421));
  not1  g1231(.din(new_new_n703__), .dout(n4424));
  not1  g1232(.din(new_new_n705__), .dout(n4427));
  not1  g1233(.din(new_new_n707__), .dout(n4430));
  not1  g1234(.din(new_new_n709__), .dout(n4433));
  not1  g1235(.din(new_new_n711__), .dout(n4436));
  not1  g1236(.din(new_new_n531__), .dout(n4439));
  not1  g1237(.din(new_new_n613__), .dout(n4442));
  not1  g1238(.din(new_new_n533__), .dout(n4445));
  not1  g1239(.din(new_new_n617__), .dout(n4448));
  not1  g1240(.din(new_new_n535__), .dout(n4451));
  not1  g1241(.din(new_new_n621__), .dout(n4454));
  not1  g1242(.din(new_new_n537__), .dout(n4457));
  not1  g1243(.din(new_new_n625__), .dout(n4460));
  not1  g1244(.din(new_new_n539__), .dout(n4463));
  not1  g1245(.din(new_new_n629__), .dout(n4466));
  not1  g1246(.din(new_new_n541__), .dout(n4469));
  not1  g1247(.din(new_new_n633__), .dout(n4472));
  not1  g1248(.din(new_new_n543__), .dout(n4475));
  not1  g1249(.din(new_new_n637__), .dout(n4478));
  not1  g1250(.din(new_new_n545__), .dout(n4481));
  not1  g1251(.din(new_new_n641__), .dout(n4484));
  not1  g1252(.din(new_new_n547__), .dout(n4487));
  not1  g1253(.din(new_new_n645__), .dout(n4490));
  not1  g1254(.din(new_new_n2296__), .dout(n4493));
  not1  g1255(.din(new_new_n2313__), .dout(n4496));
  not1  g1256(.din(new_new_n2330__), .dout(n4499));
  not1  g1257(.din(new_new_n2347__), .dout(n4502));
  not1  g1258(.din(new_new_n2294__), .dout(n4505));
  not1  g1259(.din(new_new_n2311__), .dout(n4508));
  not1  g1260(.din(new_new_n2328__), .dout(n4511));
  not1  g1261(.din(new_new_n2345__), .dout(n4514));
  not1  g1262(.din(new_new_n2304__), .dout(n4517));
  not1  g1263(.din(new_new_n2321__), .dout(n4520));
  not1  g1264(.din(new_new_n2338__), .dout(n4523));
  not1  g1265(.din(new_new_n2355__), .dout(n4526));
  not1  g1266(.din(new_new_n2302__), .dout(n4529));
  not1  g1267(.din(new_new_n2319__), .dout(n4532));
  not1  g1268(.din(new_new_n2336__), .dout(n4535));
  not1  g1269(.din(new_new_n2353__), .dout(n4538));
  not1  g1270(.din(new_new_n2364__), .dout(n4541));
  not1  g1271(.din(new_new_n2381__), .dout(n4544));
  not1  g1272(.din(new_new_n2398__), .dout(n4547));
  not1  g1273(.din(new_new_n2415__), .dout(n4550));
  not1  g1274(.din(new_new_n2362__), .dout(n4553));
  not1  g1275(.din(new_new_n2379__), .dout(n4556));
  not1  g1276(.din(new_new_n2396__), .dout(n4559));
  not1  g1277(.din(new_new_n2413__), .dout(n4562));
  not1  g1278(.din(new_new_n2372__), .dout(n4565));
  not1  g1279(.din(new_new_n2389__), .dout(n4568));
  not1  g1280(.din(new_new_n2406__), .dout(n4571));
  not1  g1281(.din(new_new_n2423__), .dout(n4574));
  not1  g1282(.din(new_new_n2370__), .dout(n4577));
  not1  g1283(.din(new_new_n2387__), .dout(n4580));
  not1  g1284(.din(new_new_n2404__), .dout(n4583));
  not1  g1285(.din(new_new_n2421__), .dout(n4586));
  not1  g1286(.din(new_new_n2185__), .dout(n4589));
  not1  g1287(.din(new_new_n2182__), .dout(n4592));
  not1  g1288(.din(new_new_n2177__), .dout(n4595));
  not1  g1289(.din(new_new_n2174__), .dout(n4598));
  not1  g1290(.din(new_new_n2204__), .dout(n4601));
  not1  g1291(.din(new_new_n2201__), .dout(n4604));
  not1  g1292(.din(new_new_n2196__), .dout(n4607));
  not1  g1293(.din(new_new_n2193__), .dout(n4610));
  not1  g1294(.din(new_new_n2432__), .dout(n4613));
  not1  g1295(.din(new_new_n2430__), .dout(n4616));
  not1  g1296(.din(new_new_n2440__), .dout(n4619));
  not1  g1297(.din(new_new_n2438__), .dout(n4622));
  not1  g1298(.din(new_new_n2449__), .dout(n4625));
  not1  g1299(.din(new_new_n2447__), .dout(n4628));
  not1  g1300(.din(new_new_n2457__), .dout(n4631));
  not1  g1301(.din(new_new_n2455__), .dout(n4634));
  not1  g1302(.din(new_new_n2466__), .dout(n4637));
  not1  g1303(.din(new_new_n2464__), .dout(n4640));
  not1  g1304(.din(new_new_n2474__), .dout(n4643));
  not1  g1305(.din(new_new_n2472__), .dout(n4646));
  not1  g1306(.din(new_new_n2483__), .dout(n4649));
  not1  g1307(.din(new_new_n2481__), .dout(n4652));
  not1  g1308(.din(new_new_n2491__), .dout(n4655));
  not1  g1309(.din(new_new_n2489__), .dout(n4658));
  not1  g1310(.din(new_new_n2500__), .dout(n4661));
  not1  g1311(.din(new_new_n2498__), .dout(n4664));
  not1  g1312(.din(new_new_n2508__), .dout(n4667));
  not1  g1313(.din(new_new_n2506__), .dout(n4670));
  not1  g1314(.din(new_new_n2517__), .dout(n4673));
  not1  g1315(.din(new_new_n2515__), .dout(n4676));
  not1  g1316(.din(new_new_n2525__), .dout(n4679));
  not1  g1317(.din(new_new_n2523__), .dout(n4682));
  not1  g1318(.din(new_new_n2534__), .dout(n4685));
  not1  g1319(.din(new_new_n2532__), .dout(n4688));
  not1  g1320(.din(new_new_n2542__), .dout(n4691));
  not1  g1321(.din(new_new_n2540__), .dout(n4694));
  not1  g1322(.din(new_new_n2551__), .dout(n4697));
  not1  g1323(.din(new_new_n2549__), .dout(n4700));
  not1  g1324(.din(new_new_n2559__), .dout(n4703));
  not1  g1325(.din(new_new_n2557__), .dout(n4706));
  not1  g1326(.din(new_new_n2186__), .dout(n4709));
  buf1  g1327(.din(n4709), .dout(n4712));
  not1  g1328(.din(new_new_n2183__), .dout(n4715));
  buf1  g1329(.din(n4715), .dout(n4718));
  not1  g1330(.din(new_new_n2178__), .dout(n4721));
  buf1  g1331(.din(n4721), .dout(n4724));
  not1  g1332(.din(new_new_n2175__), .dout(n4727));
  buf1  g1333(.din(n4727), .dout(n4730));
  not1  g1334(.din(new_new_n2205__), .dout(n4733));
  buf1  g1335(.din(n4733), .dout(n4736));
  not1  g1336(.din(new_new_n2202__), .dout(n4739));
  buf1  g1337(.din(n4739), .dout(n4742));
  not1  g1338(.din(new_new_n2197__), .dout(n4745));
  buf1  g1339(.din(n4745), .dout(n4748));
  not1  g1340(.din(new_new_n2194__), .dout(n4751));
  buf1  g1341(.din(n4751), .dout(n4754));
  not1  g1342(.din(new_new_n1273__), .dout(n4757));
  not1  g1343(.din(new_new_n1287__), .dout(n4760));
  not1  g1344(.din(new_new_n1301__), .dout(n4763));
  not1  g1345(.din(new_new_n1315__), .dout(n4766));
  not1  g1346(.din(new_new_n1329__), .dout(n4769));
  not1  g1347(.din(new_new_n1343__), .dout(n4772));
  not1  g1348(.din(new_new_n1357__), .dout(n4775));
  not1  g1349(.din(new_new_n1371__), .dout(n4778));
  not1  g1350(.din(new_new_n1385__), .dout(n4781));
  not1  g1351(.din(new_new_n1399__), .dout(n4784));
  not1  g1352(.din(new_new_n1419__), .dout(n4787));
  not1  g1353(.din(new_new_n1439__), .dout(n4790));
  not1  g1354(.din(new_new_n1459__), .dout(n4793));
  not1  g1355(.din(new_new_n1479__), .dout(n4796));
  not1  g1356(.din(new_new_n1499__), .dout(n4799));
  not1  g1357(.din(new_new_n1519__), .dout(n4802));
  not1  g1358(.din(new_new_n1539__), .dout(n4805));
  not1  g1359(.din(new_new_n1559__), .dout(n4808));
  not1  g1360(.din(new_new_n1579__), .dout(n4811));
  not1  g1361(.din(new_new_n1599__), .dout(n4814));
  not1  g1362(.din(new_new_n1619__), .dout(n4817));
  not1  g1363(.din(new_new_n1639__), .dout(n4820));
  not1  g1364(.din(new_new_n1659__), .dout(n4823));
  not1  g1365(.din(new_new_n1679__), .dout(n4826));
  not1  g1366(.din(new_new_n1699__), .dout(n4829));
  not1  g1367(.din(new_new_n1719__), .dout(n4832));
  not1  g1368(.din(new_new_n467__), .dout(n4835));
  not1  g1369(.din(new_new_n469__), .dout(n4838));
  not1  g1370(.din(new_new_n471__), .dout(n4841));
  not1  g1371(.din(new_new_n473__), .dout(n4844));
  not1  g1372(.din(new_new_n475__), .dout(n4847));
  not1  g1373(.din(new_new_n477__), .dout(n4850));
  not1  g1374(.din(new_new_n479__), .dout(n4853));
  not1  g1375(.din(new_new_n481__), .dout(n4856));
  not1  g1376(.din(new_new_n483__), .dout(n4859));
  not1  g1377(.din(new_new_n485__), .dout(n4862));
  not1  g1378(.din(new_new_n487__), .dout(n4865));
  not1  g1379(.din(new_new_n489__), .dout(n4868));
  not1  g1380(.din(new_new_n491__), .dout(n4871));
  not1  g1381(.din(new_new_n493__), .dout(n4874));
  not1  g1382(.din(new_new_n495__), .dout(n4877));
  not1  g1383(.din(new_new_n497__), .dout(n4880));
  not1  g1384(.din(new_new_n499__), .dout(n4883));
  not1  g1385(.din(new_new_n501__), .dout(n4886));
  not1  g1386(.din(new_new_n503__), .dout(n4889));
  not1  g1387(.din(new_new_n505__), .dout(n4892));
  not1  g1388(.din(new_new_n507__), .dout(n4895));
  not1  g1389(.din(new_new_n509__), .dout(n4898));
  not1  g1390(.din(new_new_n511__), .dout(n4901));
  not1  g1391(.din(new_new_n513__), .dout(n4904));
  not1  g1392(.din(new_new_n515__), .dout(n4907));
  not1  g1393(.din(new_new_n517__), .dout(n4910));
  not1  g1394(.din(new_new_n519__), .dout(n4913));
  not1  g1395(.din(new_new_n521__), .dout(n4916));
  not1  g1396(.din(new_new_n523__), .dout(n4919));
  not1  g1397(.din(new_new_n525__), .dout(n4922));
  not1  g1398(.din(new_new_n527__), .dout(n4925));
  not1  g1399(.din(new_new_n529__), .dout(n4928));
  buf1  g1400(.din(new_new_n720__), .dout(new_new_n1948__));
  buf1  g1401(.din(new_new_n1948__), .dout(new_new_n1949__));
  buf1  g1402(.din(new_new_n1949__), .dout(new_new_n1950__));
  buf1  g1403(.din(new_new_n1949__), .dout(new_new_n1951__));
  buf1  g1404(.din(new_new_n1948__), .dout(new_new_n1952__));
  buf1  g1405(.din(new_new_n721__), .dout(new_new_n1953__));
  buf1  g1406(.din(new_new_n1953__), .dout(new_new_n1954__));
  buf1  g1407(.din(new_new_n1954__), .dout(new_new_n1955__));
  buf1  g1408(.din(new_new_n1954__), .dout(new_new_n1956__));
  buf1  g1409(.din(new_new_n1953__), .dout(new_new_n1957__));
  buf1  g1410(.din(new_new_n724__), .dout(new_new_n1958__));
  buf1  g1411(.din(new_new_n1958__), .dout(new_new_n1959__));
  buf1  g1412(.din(new_new_n1959__), .dout(new_new_n1960__));
  buf1  g1413(.din(new_new_n1959__), .dout(new_new_n1961__));
  buf1  g1414(.din(new_new_n1958__), .dout(new_new_n1962__));
  buf1  g1415(.din(new_new_n725__), .dout(new_new_n1963__));
  buf1  g1416(.din(new_new_n1963__), .dout(new_new_n1964__));
  buf1  g1417(.din(new_new_n1964__), .dout(new_new_n1965__));
  buf1  g1418(.din(new_new_n1964__), .dout(new_new_n1966__));
  buf1  g1419(.din(new_new_n1963__), .dout(new_new_n1967__));
  buf1  g1420(.din(new_new_n824__), .dout(new_new_n1968__));
  buf1  g1421(.din(new_new_n1968__), .dout(new_new_n1969__));
  buf1  g1422(.din(new_new_n1968__), .dout(new_new_n1970__));
  buf1  g1423(.din(new_new_n825__), .dout(new_new_n1971__));
  buf1  g1424(.din(new_new_n1971__), .dout(new_new_n1972__));
  buf1  g1425(.din(new_new_n1971__), .dout(new_new_n1973__));
  buf1  g1426(.din(new_new_n946__), .dout(new_new_n1974__));
  buf1  g1427(.din(new_new_n1974__), .dout(new_new_n1975__));
  buf1  g1428(.din(new_new_n1974__), .dout(new_new_n1976__));
  buf1  g1429(.din(new_new_n712__), .dout(new_new_n1977__));
  buf1  g1430(.din(new_new_n1977__), .dout(new_new_n1978__));
  buf1  g1431(.din(new_new_n1978__), .dout(new_new_n1979__));
  buf1  g1432(.din(new_new_n1978__), .dout(new_new_n1980__));
  buf1  g1433(.din(new_new_n1977__), .dout(new_new_n1981__));
  buf1  g1434(.din(new_new_n947__), .dout(new_new_n1982__));
  buf1  g1435(.din(new_new_n1982__), .dout(new_new_n1983__));
  buf1  g1436(.din(new_new_n1982__), .dout(new_new_n1984__));
  buf1  g1437(.din(new_new_n713__), .dout(new_new_n1985__));
  buf1  g1438(.din(new_new_n1985__), .dout(new_new_n1986__));
  buf1  g1439(.din(new_new_n1986__), .dout(new_new_n1987__));
  buf1  g1440(.din(new_new_n1986__), .dout(new_new_n1988__));
  buf1  g1441(.din(new_new_n1985__), .dout(new_new_n1989__));
  buf1  g1442(.din(new_new_n950__), .dout(new_new_n1990__));
  buf1  g1443(.din(new_new_n714__), .dout(new_new_n1991__));
  buf1  g1444(.din(new_new_n1991__), .dout(new_new_n1992__));
  buf1  g1445(.din(new_new_n1992__), .dout(new_new_n1993__));
  buf1  g1446(.din(new_new_n1992__), .dout(new_new_n1994__));
  buf1  g1447(.din(new_new_n1991__), .dout(new_new_n1995__));
  buf1  g1448(.din(new_new_n715__), .dout(new_new_n1996__));
  buf1  g1449(.din(new_new_n1996__), .dout(new_new_n1997__));
  buf1  g1450(.din(new_new_n1997__), .dout(new_new_n1998__));
  buf1  g1451(.din(new_new_n1997__), .dout(new_new_n1999__));
  buf1  g1452(.din(new_new_n1996__), .dout(new_new_n2000__));
  buf1  g1453(.din(new_new_n956__), .dout(new_new_n2001__));
  buf1  g1454(.din(new_new_n716__), .dout(new_new_n2002__));
  buf1  g1455(.din(new_new_n2002__), .dout(new_new_n2003__));
  buf1  g1456(.din(new_new_n2003__), .dout(new_new_n2004__));
  buf1  g1457(.din(new_new_n2003__), .dout(new_new_n2005__));
  buf1  g1458(.din(new_new_n2002__), .dout(new_new_n2006__));
  buf1  g1459(.din(new_new_n717__), .dout(new_new_n2007__));
  buf1  g1460(.din(new_new_n2007__), .dout(new_new_n2008__));
  buf1  g1461(.din(new_new_n2008__), .dout(new_new_n2009__));
  buf1  g1462(.din(new_new_n2008__), .dout(new_new_n2010__));
  buf1  g1463(.din(new_new_n2007__), .dout(new_new_n2011__));
  buf1  g1464(.din(new_new_n962__), .dout(new_new_n2012__));
  buf1  g1465(.din(new_new_n718__), .dout(new_new_n2013__));
  buf1  g1466(.din(new_new_n2013__), .dout(new_new_n2014__));
  buf1  g1467(.din(new_new_n2014__), .dout(new_new_n2015__));
  buf1  g1468(.din(new_new_n2014__), .dout(new_new_n2016__));
  buf1  g1469(.din(new_new_n2013__), .dout(new_new_n2017__));
  buf1  g1470(.din(new_new_n719__), .dout(new_new_n2018__));
  buf1  g1471(.din(new_new_n2018__), .dout(new_new_n2019__));
  buf1  g1472(.din(new_new_n2019__), .dout(new_new_n2020__));
  buf1  g1473(.din(new_new_n2019__), .dout(new_new_n2021__));
  buf1  g1474(.din(new_new_n2018__), .dout(new_new_n2022__));
  buf1  g1475(.din(new_new_n968__), .dout(new_new_n2023__));
  buf1  g1476(.din(new_new_n726__), .dout(new_new_n2024__));
  buf1  g1477(.din(new_new_n2024__), .dout(new_new_n2025__));
  buf1  g1478(.din(new_new_n2025__), .dout(new_new_n2026__));
  buf1  g1479(.din(new_new_n2025__), .dout(new_new_n2027__));
  buf1  g1480(.din(new_new_n2024__), .dout(new_new_n2028__));
  buf1  g1481(.din(new_new_n727__), .dout(new_new_n2029__));
  buf1  g1482(.din(new_new_n2029__), .dout(new_new_n2030__));
  buf1  g1483(.din(new_new_n2030__), .dout(new_new_n2031__));
  buf1  g1484(.din(new_new_n2030__), .dout(new_new_n2032__));
  buf1  g1485(.din(new_new_n2029__), .dout(new_new_n2033__));
  buf1  g1486(.din(new_new_n978__), .dout(new_new_n2034__));
  buf1  g1487(.din(new_new_n2034__), .dout(new_new_n2035__));
  buf1  g1488(.din(new_new_n2034__), .dout(new_new_n2036__));
  buf1  g1489(.din(new_new_n979__), .dout(new_new_n2037__));
  buf1  g1490(.din(new_new_n2037__), .dout(new_new_n2038__));
  buf1  g1491(.din(new_new_n2037__), .dout(new_new_n2039__));
  buf1  g1492(.din(new_new_n982__), .dout(new_new_n2040__));
  buf1  g1493(.din(new_new_n988__), .dout(new_new_n2041__));
  buf1  g1494(.din(new_new_n994__), .dout(new_new_n2042__));
  buf1  g1495(.din(new_new_n1000__), .dout(new_new_n2043__));
  buf1  g1496(.din(new_new_n722__), .dout(new_new_n2044__));
  buf1  g1497(.din(new_new_n2044__), .dout(new_new_n2045__));
  buf1  g1498(.din(new_new_n2045__), .dout(new_new_n2046__));
  buf1  g1499(.din(new_new_n2045__), .dout(new_new_n2047__));
  buf1  g1500(.din(new_new_n2044__), .dout(new_new_n2048__));
  buf1  g1501(.din(new_new_n723__), .dout(new_new_n2049__));
  buf1  g1502(.din(new_new_n2049__), .dout(new_new_n2050__));
  buf1  g1503(.din(new_new_n2050__), .dout(new_new_n2051__));
  buf1  g1504(.din(new_new_n2050__), .dout(new_new_n2052__));
  buf1  g1505(.din(new_new_n2049__), .dout(new_new_n2053__));
  buf1  g1506(.din(new_new_n1010__), .dout(new_new_n2054__));
  buf1  g1507(.din(new_new_n2054__), .dout(new_new_n2055__));
  buf1  g1508(.din(new_new_n2054__), .dout(new_new_n2056__));
  buf1  g1509(.din(new_new_n1011__), .dout(new_new_n2057__));
  buf1  g1510(.din(new_new_n2057__), .dout(new_new_n2058__));
  buf1  g1511(.din(new_new_n2057__), .dout(new_new_n2059__));
  buf1  g1512(.din(new_new_n1014__), .dout(new_new_n2060__));
  buf1  g1513(.din(new_new_n1020__), .dout(new_new_n2061__));
  buf1  g1514(.din(new_new_n1026__), .dout(new_new_n2062__));
  buf1  g1515(.din(new_new_n1032__), .dout(new_new_n2063__));
  buf1  g1516(.din(new_new_n1042__), .dout(new_new_n2064__));
  buf1  g1517(.din(new_new_n2064__), .dout(new_new_n2065__));
  buf1  g1518(.din(new_new_n2064__), .dout(new_new_n2066__));
  buf1  g1519(.din(new_new_n1043__), .dout(new_new_n2067__));
  buf1  g1520(.din(new_new_n2067__), .dout(new_new_n2068__));
  buf1  g1521(.din(new_new_n2067__), .dout(new_new_n2069__));
  buf1  g1522(.din(new_new_n1046__), .dout(new_new_n2070__));
  buf1  g1523(.din(new_new_n1052__), .dout(new_new_n2071__));
  buf1  g1524(.din(new_new_n1058__), .dout(new_new_n2072__));
  buf1  g1525(.din(new_new_n1064__), .dout(new_new_n2073__));
  buf1  g1526(.din(new_new_n826__), .dout(new_new_n2074__));
  buf1  g1527(.din(new_new_n2074__), .dout(new_new_n2075__));
  buf1  g1528(.din(new_new_n2074__), .dout(new_new_n2076__));
  buf1  g1529(.din(new_new_n827__), .dout(new_new_n2077__));
  buf1  g1530(.din(new_new_n2077__), .dout(new_new_n2078__));
  buf1  g1531(.din(new_new_n2077__), .dout(new_new_n2079__));
  buf1  g1532(.din(new_new_n1074__), .dout(new_new_n2080__));
  buf1  g1533(.din(new_new_n2080__), .dout(new_new_n2081__));
  buf1  g1534(.din(new_new_n2080__), .dout(new_new_n2082__));
  buf1  g1535(.din(new_new_n1075__), .dout(new_new_n2083__));
  buf1  g1536(.din(new_new_n2083__), .dout(new_new_n2084__));
  buf1  g1537(.din(new_new_n2083__), .dout(new_new_n2085__));
  buf1  g1538(.din(new_new_n1078__), .dout(new_new_n2086__));
  buf1  g1539(.din(new_new_n1084__), .dout(new_new_n2087__));
  buf1  g1540(.din(new_new_n1090__), .dout(new_new_n2088__));
  buf1  g1541(.din(new_new_n1096__), .dout(new_new_n2089__));
  buf1  g1542(.din(new_new_n1106__), .dout(new_new_n2090__));
  buf1  g1543(.din(new_new_n2090__), .dout(new_new_n2091__));
  buf1  g1544(.din(new_new_n2090__), .dout(new_new_n2092__));
  buf1  g1545(.din(new_new_n1107__), .dout(new_new_n2093__));
  buf1  g1546(.din(new_new_n2093__), .dout(new_new_n2094__));
  buf1  g1547(.din(new_new_n2093__), .dout(new_new_n2095__));
  buf1  g1548(.din(new_new_n1110__), .dout(new_new_n2096__));
  buf1  g1549(.din(new_new_n1116__), .dout(new_new_n2097__));
  buf1  g1550(.din(new_new_n1122__), .dout(new_new_n2098__));
  buf1  g1551(.din(new_new_n1128__), .dout(new_new_n2099__));
  buf1  g1552(.din(new_new_n1138__), .dout(new_new_n2100__));
  buf1  g1553(.din(new_new_n2100__), .dout(new_new_n2101__));
  buf1  g1554(.din(new_new_n2100__), .dout(new_new_n2102__));
  buf1  g1555(.din(new_new_n1139__), .dout(new_new_n2103__));
  buf1  g1556(.din(new_new_n2103__), .dout(new_new_n2104__));
  buf1  g1557(.din(new_new_n2103__), .dout(new_new_n2105__));
  buf1  g1558(.din(new_new_n1142__), .dout(new_new_n2106__));
  buf1  g1559(.din(new_new_n1148__), .dout(new_new_n2107__));
  buf1  g1560(.din(new_new_n1154__), .dout(new_new_n2108__));
  buf1  g1561(.din(new_new_n1160__), .dout(new_new_n2109__));
  buf1  g1562(.din(new_new_n1170__), .dout(new_new_n2110__));
  buf1  g1563(.din(new_new_n2110__), .dout(new_new_n2111__));
  buf1  g1564(.din(new_new_n2110__), .dout(new_new_n2112__));
  buf1  g1565(.din(new_new_n1171__), .dout(new_new_n2113__));
  buf1  g1566(.din(new_new_n2113__), .dout(new_new_n2114__));
  buf1  g1567(.din(new_new_n2113__), .dout(new_new_n2115__));
  buf1  g1568(.din(new_new_n1174__), .dout(new_new_n2116__));
  buf1  g1569(.din(new_new_n1180__), .dout(new_new_n2117__));
  buf1  g1570(.din(new_new_n1186__), .dout(new_new_n2118__));
  buf1  g1571(.din(new_new_n1192__), .dout(new_new_n2119__));
  buf1  g1572(.din(new_new_n844__), .dout(new_new_n2120__));
  buf1  g1573(.din(new_new_n828__), .dout(new_new_n2121__));
  buf1  g1574(.din(new_new_n845__), .dout(new_new_n2122__));
  buf1  g1575(.din(new_new_n829__), .dout(new_new_n2123__));
  buf1  g1576(.din(new_new_n1197__), .dout(new_new_n2124__));
  buf1  g1577(.din(new_new_n1196__), .dout(new_new_n2125__));
  buf1  g1578(.din(new_new_n846__), .dout(new_new_n2126__));
  buf1  g1579(.din(new_new_n830__), .dout(new_new_n2127__));
  buf1  g1580(.din(new_new_n847__), .dout(new_new_n2128__));
  buf1  g1581(.din(new_new_n831__), .dout(new_new_n2129__));
  buf1  g1582(.din(new_new_n1205__), .dout(new_new_n2130__));
  buf1  g1583(.din(new_new_n1204__), .dout(new_new_n2131__));
  buf1  g1584(.din(new_new_n848__), .dout(new_new_n2132__));
  buf1  g1585(.din(new_new_n832__), .dout(new_new_n2133__));
  buf1  g1586(.din(new_new_n849__), .dout(new_new_n2134__));
  buf1  g1587(.din(new_new_n833__), .dout(new_new_n2135__));
  buf1  g1588(.din(new_new_n1213__), .dout(new_new_n2136__));
  buf1  g1589(.din(new_new_n1212__), .dout(new_new_n2137__));
  buf1  g1590(.din(new_new_n850__), .dout(new_new_n2138__));
  buf1  g1591(.din(new_new_n834__), .dout(new_new_n2139__));
  buf1  g1592(.din(new_new_n851__), .dout(new_new_n2140__));
  buf1  g1593(.din(new_new_n835__), .dout(new_new_n2141__));
  buf1  g1594(.din(new_new_n1221__), .dout(new_new_n2142__));
  buf1  g1595(.din(new_new_n1220__), .dout(new_new_n2143__));
  buf1  g1596(.din(new_new_n852__), .dout(new_new_n2144__));
  buf1  g1597(.din(new_new_n836__), .dout(new_new_n2145__));
  buf1  g1598(.din(new_new_n853__), .dout(new_new_n2146__));
  buf1  g1599(.din(new_new_n837__), .dout(new_new_n2147__));
  buf1  g1600(.din(new_new_n1229__), .dout(new_new_n2148__));
  buf1  g1601(.din(new_new_n1228__), .dout(new_new_n2149__));
  buf1  g1602(.din(new_new_n854__), .dout(new_new_n2150__));
  buf1  g1603(.din(new_new_n838__), .dout(new_new_n2151__));
  buf1  g1604(.din(new_new_n855__), .dout(new_new_n2152__));
  buf1  g1605(.din(new_new_n839__), .dout(new_new_n2153__));
  buf1  g1606(.din(new_new_n1237__), .dout(new_new_n2154__));
  buf1  g1607(.din(new_new_n1236__), .dout(new_new_n2155__));
  buf1  g1608(.din(new_new_n856__), .dout(new_new_n2156__));
  buf1  g1609(.din(new_new_n840__), .dout(new_new_n2157__));
  buf1  g1610(.din(new_new_n857__), .dout(new_new_n2158__));
  buf1  g1611(.din(new_new_n841__), .dout(new_new_n2159__));
  buf1  g1612(.din(new_new_n1245__), .dout(new_new_n2160__));
  buf1  g1613(.din(new_new_n1244__), .dout(new_new_n2161__));
  buf1  g1614(.din(new_new_n858__), .dout(new_new_n2162__));
  buf1  g1615(.din(new_new_n842__), .dout(new_new_n2163__));
  buf1  g1616(.din(new_new_n859__), .dout(new_new_n2164__));
  buf1  g1617(.din(new_new_n843__), .dout(new_new_n2165__));
  buf1  g1618(.din(new_new_n1253__), .dout(new_new_n2166__));
  buf1  g1619(.din(new_new_n1252__), .dout(new_new_n2167__));
  buf1  g1620(.din(new_new_n1211__), .dout(new_new_n2168__));
  buf1  g1621(.din(new_new_n1203__), .dout(new_new_n2169__));
  buf1  g1622(.din(new_new_n1260__), .dout(new_new_n2170__));
  buf1  g1623(.din(new_new_n1219__), .dout(new_new_n2171__));
  buf1  g1624(.din(new_new_n2171__), .dout(new_new_n2172__));
  buf1  g1625(.din(new_new_n1226__), .dout(new_new_n2173__));
  buf1  g1626(.din(new_new_n2173__), .dout(new_new_n2174__));
  buf1  g1627(.din(new_new_n2173__), .dout(new_new_n2175__));
  buf1  g1628(.din(new_new_n1218__), .dout(new_new_n2176__));
  buf1  g1629(.din(new_new_n2176__), .dout(new_new_n2177__));
  buf1  g1630(.din(new_new_n2176__), .dout(new_new_n2178__));
  buf1  g1631(.din(new_new_n1227__), .dout(new_new_n2179__));
  buf1  g1632(.din(new_new_n2179__), .dout(new_new_n2180__));
  buf1  g1633(.din(new_new_n1210__), .dout(new_new_n2181__));
  buf1  g1634(.din(new_new_n2181__), .dout(new_new_n2182__));
  buf1  g1635(.din(new_new_n2181__), .dout(new_new_n2183__));
  buf1  g1636(.din(new_new_n1202__), .dout(new_new_n2184__));
  buf1  g1637(.din(new_new_n2184__), .dout(new_new_n2185__));
  buf1  g1638(.din(new_new_n2184__), .dout(new_new_n2186__));
  buf1  g1639(.din(new_new_n1243__), .dout(new_new_n2187__));
  buf1  g1640(.din(new_new_n1235__), .dout(new_new_n2188__));
  buf1  g1641(.din(new_new_n1274__), .dout(new_new_n2189__));
  buf1  g1642(.din(new_new_n1251__), .dout(new_new_n2190__));
  buf1  g1643(.din(new_new_n2190__), .dout(new_new_n2191__));
  buf1  g1644(.din(new_new_n1258__), .dout(new_new_n2192__));
  buf1  g1645(.din(new_new_n2192__), .dout(new_new_n2193__));
  buf1  g1646(.din(new_new_n2192__), .dout(new_new_n2194__));
  buf1  g1647(.din(new_new_n1250__), .dout(new_new_n2195__));
  buf1  g1648(.din(new_new_n2195__), .dout(new_new_n2196__));
  buf1  g1649(.din(new_new_n2195__), .dout(new_new_n2197__));
  buf1  g1650(.din(new_new_n1259__), .dout(new_new_n2198__));
  buf1  g1651(.din(new_new_n2198__), .dout(new_new_n2199__));
  buf1  g1652(.din(new_new_n1242__), .dout(new_new_n2200__));
  buf1  g1653(.din(new_new_n2200__), .dout(new_new_n2201__));
  buf1  g1654(.din(new_new_n2200__), .dout(new_new_n2202__));
  buf1  g1655(.din(new_new_n1234__), .dout(new_new_n2203__));
  buf1  g1656(.din(new_new_n2203__), .dout(new_new_n2204__));
  buf1  g1657(.din(new_new_n2203__), .dout(new_new_n2205__));
  buf1  g1658(.din(new_new_n646__), .dout(new_new_n2206__));
  buf1  g1659(.din(new_new_n2206__), .dout(new_new_n2207__));
  buf1  g1660(.din(new_new_n2207__), .dout(new_new_n2208__));
  buf1  g1661(.din(new_new_n2207__), .dout(new_new_n2209__));
  buf1  g1662(.din(new_new_n2206__), .dout(new_new_n2210__));
  buf1  g1663(.din(new_new_n2210__), .dout(new_new_n2211__));
  buf1  g1664(.din(new_new_n2210__), .dout(new_new_n2212__));
  buf1  g1665(.din(new_new_n647__), .dout(new_new_n2213__));
  buf1  g1666(.din(new_new_n2213__), .dout(new_new_n2214__));
  buf1  g1667(.din(new_new_n2214__), .dout(new_new_n2215__));
  buf1  g1668(.din(new_new_n2214__), .dout(new_new_n2216__));
  buf1  g1669(.din(new_new_n2213__), .dout(new_new_n2217__));
  buf1  g1670(.din(new_new_n2217__), .dout(new_new_n2218__));
  buf1  g1671(.din(new_new_n2217__), .dout(new_new_n2219__));
  buf1  g1672(.din(new_new_n870__), .dout(new_new_n2220__));
  buf1  g1673(.din(new_new_n2220__), .dout(new_new_n2221__));
  buf1  g1674(.din(new_new_n2220__), .dout(new_new_n2222__));
  buf1  g1675(.din(new_new_n868__), .dout(new_new_n2223__));
  buf1  g1676(.din(new_new_n2223__), .dout(new_new_n2224__));
  buf1  g1677(.din(new_new_n2223__), .dout(new_new_n2225__));
  buf1  g1678(.din(new_new_n871__), .dout(new_new_n2226__));
  buf1  g1679(.din(new_new_n2226__), .dout(new_new_n2227__));
  buf1  g1680(.din(new_new_n2226__), .dout(new_new_n2228__));
  buf1  g1681(.din(new_new_n869__), .dout(new_new_n2229__));
  buf1  g1682(.din(new_new_n2229__), .dout(new_new_n2230__));
  buf1  g1683(.din(new_new_n2229__), .dout(new_new_n2231__));
  buf1  g1684(.din(new_new_n1291__), .dout(new_new_n2232__));
  buf1  g1685(.din(new_new_n1290__), .dout(new_new_n2233__));
  buf1  g1686(.din(new_new_n1298__), .dout(new_new_n2234__));
  buf1  g1687(.din(new_new_n874__), .dout(new_new_n2235__));
  buf1  g1688(.din(new_new_n2235__), .dout(new_new_n2236__));
  buf1  g1689(.din(new_new_n2235__), .dout(new_new_n2237__));
  buf1  g1690(.din(new_new_n872__), .dout(new_new_n2238__));
  buf1  g1691(.din(new_new_n2238__), .dout(new_new_n2239__));
  buf1  g1692(.din(new_new_n2238__), .dout(new_new_n2240__));
  buf1  g1693(.din(new_new_n875__), .dout(new_new_n2241__));
  buf1  g1694(.din(new_new_n2241__), .dout(new_new_n2242__));
  buf1  g1695(.din(new_new_n2241__), .dout(new_new_n2243__));
  buf1  g1696(.din(new_new_n873__), .dout(new_new_n2244__));
  buf1  g1697(.din(new_new_n2244__), .dout(new_new_n2245__));
  buf1  g1698(.din(new_new_n2244__), .dout(new_new_n2246__));
  buf1  g1699(.din(new_new_n1305__), .dout(new_new_n2247__));
  buf1  g1700(.din(new_new_n1304__), .dout(new_new_n2248__));
  buf1  g1701(.din(new_new_n1312__), .dout(new_new_n2249__));
  buf1  g1702(.din(new_new_n1319__), .dout(new_new_n2250__));
  buf1  g1703(.din(new_new_n1318__), .dout(new_new_n2251__));
  buf1  g1704(.din(new_new_n1326__), .dout(new_new_n2252__));
  buf1  g1705(.din(new_new_n1333__), .dout(new_new_n2253__));
  buf1  g1706(.din(new_new_n1332__), .dout(new_new_n2254__));
  buf1  g1707(.din(new_new_n1340__), .dout(new_new_n2255__));
  buf1  g1708(.din(new_new_n862__), .dout(new_new_n2256__));
  buf1  g1709(.din(new_new_n2256__), .dout(new_new_n2257__));
  buf1  g1710(.din(new_new_n2256__), .dout(new_new_n2258__));
  buf1  g1711(.din(new_new_n860__), .dout(new_new_n2259__));
  buf1  g1712(.din(new_new_n2259__), .dout(new_new_n2260__));
  buf1  g1713(.din(new_new_n2259__), .dout(new_new_n2261__));
  buf1  g1714(.din(new_new_n863__), .dout(new_new_n2262__));
  buf1  g1715(.din(new_new_n2262__), .dout(new_new_n2263__));
  buf1  g1716(.din(new_new_n2262__), .dout(new_new_n2264__));
  buf1  g1717(.din(new_new_n861__), .dout(new_new_n2265__));
  buf1  g1718(.din(new_new_n2265__), .dout(new_new_n2266__));
  buf1  g1719(.din(new_new_n2265__), .dout(new_new_n2267__));
  buf1  g1720(.din(new_new_n1347__), .dout(new_new_n2268__));
  buf1  g1721(.din(new_new_n1346__), .dout(new_new_n2269__));
  buf1  g1722(.din(new_new_n1354__), .dout(new_new_n2270__));
  buf1  g1723(.din(new_new_n866__), .dout(new_new_n2271__));
  buf1  g1724(.din(new_new_n2271__), .dout(new_new_n2272__));
  buf1  g1725(.din(new_new_n2271__), .dout(new_new_n2273__));
  buf1  g1726(.din(new_new_n864__), .dout(new_new_n2274__));
  buf1  g1727(.din(new_new_n2274__), .dout(new_new_n2275__));
  buf1  g1728(.din(new_new_n2274__), .dout(new_new_n2276__));
  buf1  g1729(.din(new_new_n867__), .dout(new_new_n2277__));
  buf1  g1730(.din(new_new_n2277__), .dout(new_new_n2278__));
  buf1  g1731(.din(new_new_n2277__), .dout(new_new_n2279__));
  buf1  g1732(.din(new_new_n865__), .dout(new_new_n2280__));
  buf1  g1733(.din(new_new_n2280__), .dout(new_new_n2281__));
  buf1  g1734(.din(new_new_n2280__), .dout(new_new_n2282__));
  buf1  g1735(.din(new_new_n1361__), .dout(new_new_n2283__));
  buf1  g1736(.din(new_new_n1360__), .dout(new_new_n2284__));
  buf1  g1737(.din(new_new_n1368__), .dout(new_new_n2285__));
  buf1  g1738(.din(new_new_n1375__), .dout(new_new_n2286__));
  buf1  g1739(.din(new_new_n1374__), .dout(new_new_n2287__));
  buf1  g1740(.din(new_new_n1382__), .dout(new_new_n2288__));
  buf1  g1741(.din(new_new_n1389__), .dout(new_new_n2289__));
  buf1  g1742(.din(new_new_n1388__), .dout(new_new_n2290__));
  buf1  g1743(.din(new_new_n1396__), .dout(new_new_n2291__));
  buf1  g1744(.din(new_new_n736__), .dout(new_new_n2292__));
  buf1  g1745(.din(new_new_n728__), .dout(new_new_n2293__));
  buf1  g1746(.din(new_new_n737__), .dout(new_new_n2294__));
  buf1  g1747(.din(new_new_n2294__), .dout(new_new_n2295__));
  buf1  g1748(.din(new_new_n729__), .dout(new_new_n2296__));
  buf1  g1749(.din(new_new_n2296__), .dout(new_new_n2297__));
  buf1  g1750(.din(new_new_n1401__), .dout(new_new_n2298__));
  buf1  g1751(.din(new_new_n1400__), .dout(new_new_n2299__));
  buf1  g1752(.din(new_new_n752__), .dout(new_new_n2300__));
  buf1  g1753(.din(new_new_n744__), .dout(new_new_n2301__));
  buf1  g1754(.din(new_new_n753__), .dout(new_new_n2302__));
  buf1  g1755(.din(new_new_n2302__), .dout(new_new_n2303__));
  buf1  g1756(.din(new_new_n745__), .dout(new_new_n2304__));
  buf1  g1757(.din(new_new_n2304__), .dout(new_new_n2305__));
  buf1  g1758(.din(new_new_n1409__), .dout(new_new_n2306__));
  buf1  g1759(.din(new_new_n1408__), .dout(new_new_n2307__));
  buf1  g1760(.din(new_new_n1416__), .dout(new_new_n2308__));
  buf1  g1761(.din(new_new_n738__), .dout(new_new_n2309__));
  buf1  g1762(.din(new_new_n730__), .dout(new_new_n2310__));
  buf1  g1763(.din(new_new_n739__), .dout(new_new_n2311__));
  buf1  g1764(.din(new_new_n2311__), .dout(new_new_n2312__));
  buf1  g1765(.din(new_new_n731__), .dout(new_new_n2313__));
  buf1  g1766(.din(new_new_n2313__), .dout(new_new_n2314__));
  buf1  g1767(.din(new_new_n1421__), .dout(new_new_n2315__));
  buf1  g1768(.din(new_new_n1420__), .dout(new_new_n2316__));
  buf1  g1769(.din(new_new_n754__), .dout(new_new_n2317__));
  buf1  g1770(.din(new_new_n746__), .dout(new_new_n2318__));
  buf1  g1771(.din(new_new_n755__), .dout(new_new_n2319__));
  buf1  g1772(.din(new_new_n2319__), .dout(new_new_n2320__));
  buf1  g1773(.din(new_new_n747__), .dout(new_new_n2321__));
  buf1  g1774(.din(new_new_n2321__), .dout(new_new_n2322__));
  buf1  g1775(.din(new_new_n1429__), .dout(new_new_n2323__));
  buf1  g1776(.din(new_new_n1428__), .dout(new_new_n2324__));
  buf1  g1777(.din(new_new_n1436__), .dout(new_new_n2325__));
  buf1  g1778(.din(new_new_n740__), .dout(new_new_n2326__));
  buf1  g1779(.din(new_new_n732__), .dout(new_new_n2327__));
  buf1  g1780(.din(new_new_n741__), .dout(new_new_n2328__));
  buf1  g1781(.din(new_new_n2328__), .dout(new_new_n2329__));
  buf1  g1782(.din(new_new_n733__), .dout(new_new_n2330__));
  buf1  g1783(.din(new_new_n2330__), .dout(new_new_n2331__));
  buf1  g1784(.din(new_new_n1441__), .dout(new_new_n2332__));
  buf1  g1785(.din(new_new_n1440__), .dout(new_new_n2333__));
  buf1  g1786(.din(new_new_n756__), .dout(new_new_n2334__));
  buf1  g1787(.din(new_new_n748__), .dout(new_new_n2335__));
  buf1  g1788(.din(new_new_n757__), .dout(new_new_n2336__));
  buf1  g1789(.din(new_new_n2336__), .dout(new_new_n2337__));
  buf1  g1790(.din(new_new_n749__), .dout(new_new_n2338__));
  buf1  g1791(.din(new_new_n2338__), .dout(new_new_n2339__));
  buf1  g1792(.din(new_new_n1449__), .dout(new_new_n2340__));
  buf1  g1793(.din(new_new_n1448__), .dout(new_new_n2341__));
  buf1  g1794(.din(new_new_n1456__), .dout(new_new_n2342__));
  buf1  g1795(.din(new_new_n742__), .dout(new_new_n2343__));
  buf1  g1796(.din(new_new_n734__), .dout(new_new_n2344__));
  buf1  g1797(.din(new_new_n743__), .dout(new_new_n2345__));
  buf1  g1798(.din(new_new_n2345__), .dout(new_new_n2346__));
  buf1  g1799(.din(new_new_n735__), .dout(new_new_n2347__));
  buf1  g1800(.din(new_new_n2347__), .dout(new_new_n2348__));
  buf1  g1801(.din(new_new_n1461__), .dout(new_new_n2349__));
  buf1  g1802(.din(new_new_n1460__), .dout(new_new_n2350__));
  buf1  g1803(.din(new_new_n758__), .dout(new_new_n2351__));
  buf1  g1804(.din(new_new_n750__), .dout(new_new_n2352__));
  buf1  g1805(.din(new_new_n759__), .dout(new_new_n2353__));
  buf1  g1806(.din(new_new_n2353__), .dout(new_new_n2354__));
  buf1  g1807(.din(new_new_n751__), .dout(new_new_n2355__));
  buf1  g1808(.din(new_new_n2355__), .dout(new_new_n2356__));
  buf1  g1809(.din(new_new_n1469__), .dout(new_new_n2357__));
  buf1  g1810(.din(new_new_n1468__), .dout(new_new_n2358__));
  buf1  g1811(.din(new_new_n1476__), .dout(new_new_n2359__));
  buf1  g1812(.din(new_new_n768__), .dout(new_new_n2360__));
  buf1  g1813(.din(new_new_n760__), .dout(new_new_n2361__));
  buf1  g1814(.din(new_new_n769__), .dout(new_new_n2362__));
  buf1  g1815(.din(new_new_n2362__), .dout(new_new_n2363__));
  buf1  g1816(.din(new_new_n761__), .dout(new_new_n2364__));
  buf1  g1817(.din(new_new_n2364__), .dout(new_new_n2365__));
  buf1  g1818(.din(new_new_n1481__), .dout(new_new_n2366__));
  buf1  g1819(.din(new_new_n1480__), .dout(new_new_n2367__));
  buf1  g1820(.din(new_new_n784__), .dout(new_new_n2368__));
  buf1  g1821(.din(new_new_n776__), .dout(new_new_n2369__));
  buf1  g1822(.din(new_new_n785__), .dout(new_new_n2370__));
  buf1  g1823(.din(new_new_n2370__), .dout(new_new_n2371__));
  buf1  g1824(.din(new_new_n777__), .dout(new_new_n2372__));
  buf1  g1825(.din(new_new_n2372__), .dout(new_new_n2373__));
  buf1  g1826(.din(new_new_n1489__), .dout(new_new_n2374__));
  buf1  g1827(.din(new_new_n1488__), .dout(new_new_n2375__));
  buf1  g1828(.din(new_new_n1496__), .dout(new_new_n2376__));
  buf1  g1829(.din(new_new_n770__), .dout(new_new_n2377__));
  buf1  g1830(.din(new_new_n762__), .dout(new_new_n2378__));
  buf1  g1831(.din(new_new_n771__), .dout(new_new_n2379__));
  buf1  g1832(.din(new_new_n2379__), .dout(new_new_n2380__));
  buf1  g1833(.din(new_new_n763__), .dout(new_new_n2381__));
  buf1  g1834(.din(new_new_n2381__), .dout(new_new_n2382__));
  buf1  g1835(.din(new_new_n1501__), .dout(new_new_n2383__));
  buf1  g1836(.din(new_new_n1500__), .dout(new_new_n2384__));
  buf1  g1837(.din(new_new_n786__), .dout(new_new_n2385__));
  buf1  g1838(.din(new_new_n778__), .dout(new_new_n2386__));
  buf1  g1839(.din(new_new_n787__), .dout(new_new_n2387__));
  buf1  g1840(.din(new_new_n2387__), .dout(new_new_n2388__));
  buf1  g1841(.din(new_new_n779__), .dout(new_new_n2389__));
  buf1  g1842(.din(new_new_n2389__), .dout(new_new_n2390__));
  buf1  g1843(.din(new_new_n1509__), .dout(new_new_n2391__));
  buf1  g1844(.din(new_new_n1508__), .dout(new_new_n2392__));
  buf1  g1845(.din(new_new_n1516__), .dout(new_new_n2393__));
  buf1  g1846(.din(new_new_n772__), .dout(new_new_n2394__));
  buf1  g1847(.din(new_new_n764__), .dout(new_new_n2395__));
  buf1  g1848(.din(new_new_n773__), .dout(new_new_n2396__));
  buf1  g1849(.din(new_new_n2396__), .dout(new_new_n2397__));
  buf1  g1850(.din(new_new_n765__), .dout(new_new_n2398__));
  buf1  g1851(.din(new_new_n2398__), .dout(new_new_n2399__));
  buf1  g1852(.din(new_new_n1521__), .dout(new_new_n2400__));
  buf1  g1853(.din(new_new_n1520__), .dout(new_new_n2401__));
  buf1  g1854(.din(new_new_n788__), .dout(new_new_n2402__));
  buf1  g1855(.din(new_new_n780__), .dout(new_new_n2403__));
  buf1  g1856(.din(new_new_n789__), .dout(new_new_n2404__));
  buf1  g1857(.din(new_new_n2404__), .dout(new_new_n2405__));
  buf1  g1858(.din(new_new_n781__), .dout(new_new_n2406__));
  buf1  g1859(.din(new_new_n2406__), .dout(new_new_n2407__));
  buf1  g1860(.din(new_new_n1529__), .dout(new_new_n2408__));
  buf1  g1861(.din(new_new_n1528__), .dout(new_new_n2409__));
  buf1  g1862(.din(new_new_n1536__), .dout(new_new_n2410__));
  buf1  g1863(.din(new_new_n774__), .dout(new_new_n2411__));
  buf1  g1864(.din(new_new_n766__), .dout(new_new_n2412__));
  buf1  g1865(.din(new_new_n775__), .dout(new_new_n2413__));
  buf1  g1866(.din(new_new_n2413__), .dout(new_new_n2414__));
  buf1  g1867(.din(new_new_n767__), .dout(new_new_n2415__));
  buf1  g1868(.din(new_new_n2415__), .dout(new_new_n2416__));
  buf1  g1869(.din(new_new_n1541__), .dout(new_new_n2417__));
  buf1  g1870(.din(new_new_n1540__), .dout(new_new_n2418__));
  buf1  g1871(.din(new_new_n790__), .dout(new_new_n2419__));
  buf1  g1872(.din(new_new_n782__), .dout(new_new_n2420__));
  buf1  g1873(.din(new_new_n791__), .dout(new_new_n2421__));
  buf1  g1874(.din(new_new_n2421__), .dout(new_new_n2422__));
  buf1  g1875(.din(new_new_n783__), .dout(new_new_n2423__));
  buf1  g1876(.din(new_new_n2423__), .dout(new_new_n2424__));
  buf1  g1877(.din(new_new_n1549__), .dout(new_new_n2425__));
  buf1  g1878(.din(new_new_n1548__), .dout(new_new_n2426__));
  buf1  g1879(.din(new_new_n1556__), .dout(new_new_n2427__));
  buf1  g1880(.din(new_new_n878__), .dout(new_new_n2428__));
  buf1  g1881(.din(new_new_n876__), .dout(new_new_n2429__));
  buf1  g1882(.din(new_new_n879__), .dout(new_new_n2430__));
  buf1  g1883(.din(new_new_n2430__), .dout(new_new_n2431__));
  buf1  g1884(.din(new_new_n877__), .dout(new_new_n2432__));
  buf1  g1885(.din(new_new_n2432__), .dout(new_new_n2433__));
  buf1  g1886(.din(new_new_n1561__), .dout(new_new_n2434__));
  buf1  g1887(.din(new_new_n1560__), .dout(new_new_n2435__));
  buf1  g1888(.din(new_new_n882__), .dout(new_new_n2436__));
  buf1  g1889(.din(new_new_n880__), .dout(new_new_n2437__));
  buf1  g1890(.din(new_new_n883__), .dout(new_new_n2438__));
  buf1  g1891(.din(new_new_n2438__), .dout(new_new_n2439__));
  buf1  g1892(.din(new_new_n881__), .dout(new_new_n2440__));
  buf1  g1893(.din(new_new_n2440__), .dout(new_new_n2441__));
  buf1  g1894(.din(new_new_n1569__), .dout(new_new_n2442__));
  buf1  g1895(.din(new_new_n1568__), .dout(new_new_n2443__));
  buf1  g1896(.din(new_new_n1576__), .dout(new_new_n2444__));
  buf1  g1897(.din(new_new_n886__), .dout(new_new_n2445__));
  buf1  g1898(.din(new_new_n884__), .dout(new_new_n2446__));
  buf1  g1899(.din(new_new_n887__), .dout(new_new_n2447__));
  buf1  g1900(.din(new_new_n2447__), .dout(new_new_n2448__));
  buf1  g1901(.din(new_new_n885__), .dout(new_new_n2449__));
  buf1  g1902(.din(new_new_n2449__), .dout(new_new_n2450__));
  buf1  g1903(.din(new_new_n1581__), .dout(new_new_n2451__));
  buf1  g1904(.din(new_new_n1580__), .dout(new_new_n2452__));
  buf1  g1905(.din(new_new_n890__), .dout(new_new_n2453__));
  buf1  g1906(.din(new_new_n888__), .dout(new_new_n2454__));
  buf1  g1907(.din(new_new_n891__), .dout(new_new_n2455__));
  buf1  g1908(.din(new_new_n2455__), .dout(new_new_n2456__));
  buf1  g1909(.din(new_new_n889__), .dout(new_new_n2457__));
  buf1  g1910(.din(new_new_n2457__), .dout(new_new_n2458__));
  buf1  g1911(.din(new_new_n1589__), .dout(new_new_n2459__));
  buf1  g1912(.din(new_new_n1588__), .dout(new_new_n2460__));
  buf1  g1913(.din(new_new_n1596__), .dout(new_new_n2461__));
  buf1  g1914(.din(new_new_n894__), .dout(new_new_n2462__));
  buf1  g1915(.din(new_new_n892__), .dout(new_new_n2463__));
  buf1  g1916(.din(new_new_n895__), .dout(new_new_n2464__));
  buf1  g1917(.din(new_new_n2464__), .dout(new_new_n2465__));
  buf1  g1918(.din(new_new_n893__), .dout(new_new_n2466__));
  buf1  g1919(.din(new_new_n2466__), .dout(new_new_n2467__));
  buf1  g1920(.din(new_new_n1601__), .dout(new_new_n2468__));
  buf1  g1921(.din(new_new_n1600__), .dout(new_new_n2469__));
  buf1  g1922(.din(new_new_n898__), .dout(new_new_n2470__));
  buf1  g1923(.din(new_new_n896__), .dout(new_new_n2471__));
  buf1  g1924(.din(new_new_n899__), .dout(new_new_n2472__));
  buf1  g1925(.din(new_new_n2472__), .dout(new_new_n2473__));
  buf1  g1926(.din(new_new_n897__), .dout(new_new_n2474__));
  buf1  g1927(.din(new_new_n2474__), .dout(new_new_n2475__));
  buf1  g1928(.din(new_new_n1609__), .dout(new_new_n2476__));
  buf1  g1929(.din(new_new_n1608__), .dout(new_new_n2477__));
  buf1  g1930(.din(new_new_n1616__), .dout(new_new_n2478__));
  buf1  g1931(.din(new_new_n902__), .dout(new_new_n2479__));
  buf1  g1932(.din(new_new_n900__), .dout(new_new_n2480__));
  buf1  g1933(.din(new_new_n903__), .dout(new_new_n2481__));
  buf1  g1934(.din(new_new_n2481__), .dout(new_new_n2482__));
  buf1  g1935(.din(new_new_n901__), .dout(new_new_n2483__));
  buf1  g1936(.din(new_new_n2483__), .dout(new_new_n2484__));
  buf1  g1937(.din(new_new_n1621__), .dout(new_new_n2485__));
  buf1  g1938(.din(new_new_n1620__), .dout(new_new_n2486__));
  buf1  g1939(.din(new_new_n906__), .dout(new_new_n2487__));
  buf1  g1940(.din(new_new_n904__), .dout(new_new_n2488__));
  buf1  g1941(.din(new_new_n907__), .dout(new_new_n2489__));
  buf1  g1942(.din(new_new_n2489__), .dout(new_new_n2490__));
  buf1  g1943(.din(new_new_n905__), .dout(new_new_n2491__));
  buf1  g1944(.din(new_new_n2491__), .dout(new_new_n2492__));
  buf1  g1945(.din(new_new_n1629__), .dout(new_new_n2493__));
  buf1  g1946(.din(new_new_n1628__), .dout(new_new_n2494__));
  buf1  g1947(.din(new_new_n1636__), .dout(new_new_n2495__));
  buf1  g1948(.din(new_new_n910__), .dout(new_new_n2496__));
  buf1  g1949(.din(new_new_n908__), .dout(new_new_n2497__));
  buf1  g1950(.din(new_new_n911__), .dout(new_new_n2498__));
  buf1  g1951(.din(new_new_n2498__), .dout(new_new_n2499__));
  buf1  g1952(.din(new_new_n909__), .dout(new_new_n2500__));
  buf1  g1953(.din(new_new_n2500__), .dout(new_new_n2501__));
  buf1  g1954(.din(new_new_n1641__), .dout(new_new_n2502__));
  buf1  g1955(.din(new_new_n1640__), .dout(new_new_n2503__));
  buf1  g1956(.din(new_new_n914__), .dout(new_new_n2504__));
  buf1  g1957(.din(new_new_n912__), .dout(new_new_n2505__));
  buf1  g1958(.din(new_new_n915__), .dout(new_new_n2506__));
  buf1  g1959(.din(new_new_n2506__), .dout(new_new_n2507__));
  buf1  g1960(.din(new_new_n913__), .dout(new_new_n2508__));
  buf1  g1961(.din(new_new_n2508__), .dout(new_new_n2509__));
  buf1  g1962(.din(new_new_n1649__), .dout(new_new_n2510__));
  buf1  g1963(.din(new_new_n1648__), .dout(new_new_n2511__));
  buf1  g1964(.din(new_new_n1656__), .dout(new_new_n2512__));
  buf1  g1965(.din(new_new_n918__), .dout(new_new_n2513__));
  buf1  g1966(.din(new_new_n916__), .dout(new_new_n2514__));
  buf1  g1967(.din(new_new_n919__), .dout(new_new_n2515__));
  buf1  g1968(.din(new_new_n2515__), .dout(new_new_n2516__));
  buf1  g1969(.din(new_new_n917__), .dout(new_new_n2517__));
  buf1  g1970(.din(new_new_n2517__), .dout(new_new_n2518__));
  buf1  g1971(.din(new_new_n1661__), .dout(new_new_n2519__));
  buf1  g1972(.din(new_new_n1660__), .dout(new_new_n2520__));
  buf1  g1973(.din(new_new_n922__), .dout(new_new_n2521__));
  buf1  g1974(.din(new_new_n920__), .dout(new_new_n2522__));
  buf1  g1975(.din(new_new_n923__), .dout(new_new_n2523__));
  buf1  g1976(.din(new_new_n2523__), .dout(new_new_n2524__));
  buf1  g1977(.din(new_new_n921__), .dout(new_new_n2525__));
  buf1  g1978(.din(new_new_n2525__), .dout(new_new_n2526__));
  buf1  g1979(.din(new_new_n1669__), .dout(new_new_n2527__));
  buf1  g1980(.din(new_new_n1668__), .dout(new_new_n2528__));
  buf1  g1981(.din(new_new_n1676__), .dout(new_new_n2529__));
  buf1  g1982(.din(new_new_n926__), .dout(new_new_n2530__));
  buf1  g1983(.din(new_new_n924__), .dout(new_new_n2531__));
  buf1  g1984(.din(new_new_n927__), .dout(new_new_n2532__));
  buf1  g1985(.din(new_new_n2532__), .dout(new_new_n2533__));
  buf1  g1986(.din(new_new_n925__), .dout(new_new_n2534__));
  buf1  g1987(.din(new_new_n2534__), .dout(new_new_n2535__));
  buf1  g1988(.din(new_new_n1681__), .dout(new_new_n2536__));
  buf1  g1989(.din(new_new_n1680__), .dout(new_new_n2537__));
  buf1  g1990(.din(new_new_n930__), .dout(new_new_n2538__));
  buf1  g1991(.din(new_new_n928__), .dout(new_new_n2539__));
  buf1  g1992(.din(new_new_n931__), .dout(new_new_n2540__));
  buf1  g1993(.din(new_new_n2540__), .dout(new_new_n2541__));
  buf1  g1994(.din(new_new_n929__), .dout(new_new_n2542__));
  buf1  g1995(.din(new_new_n2542__), .dout(new_new_n2543__));
  buf1  g1996(.din(new_new_n1689__), .dout(new_new_n2544__));
  buf1  g1997(.din(new_new_n1688__), .dout(new_new_n2545__));
  buf1  g1998(.din(new_new_n1696__), .dout(new_new_n2546__));
  buf1  g1999(.din(new_new_n934__), .dout(new_new_n2547__));
  buf1  g2000(.din(new_new_n932__), .dout(new_new_n2548__));
  buf1  g2001(.din(new_new_n935__), .dout(new_new_n2549__));
  buf1  g2002(.din(new_new_n2549__), .dout(new_new_n2550__));
  buf1  g2003(.din(new_new_n933__), .dout(new_new_n2551__));
  buf1  g2004(.din(new_new_n2551__), .dout(new_new_n2552__));
  buf1  g2005(.din(new_new_n1701__), .dout(new_new_n2553__));
  buf1  g2006(.din(new_new_n1700__), .dout(new_new_n2554__));
  buf1  g2007(.din(new_new_n938__), .dout(new_new_n2555__));
  buf1  g2008(.din(new_new_n936__), .dout(new_new_n2556__));
  buf1  g2009(.din(new_new_n939__), .dout(new_new_n2557__));
  buf1  g2010(.din(new_new_n2557__), .dout(new_new_n2558__));
  buf1  g2011(.din(new_new_n937__), .dout(new_new_n2559__));
  buf1  g2012(.din(new_new_n2559__), .dout(new_new_n2560__));
  buf1  g2013(.din(new_new_n1709__), .dout(new_new_n2561__));
  buf1  g2014(.din(new_new_n1708__), .dout(new_new_n2562__));
  buf1  g2015(.din(new_new_n1716__), .dout(new_new_n2563__));
  always @ (posedge clock) begin
    n630_lo <= n4343;
    n642_lo <= n4346;
    n654_lo <= n4349;
    n666_lo <= n4352;
    n678_lo <= n4355;
    n690_lo <= n4358;
    n702_lo <= n4361;
    n714_lo <= n4364;
    n726_lo <= n4367;
    n738_lo <= n4370;
    n750_lo <= n4373;
    n762_lo <= n4376;
    n774_lo <= n4379;
    n786_lo <= n4382;
    n798_lo <= n4385;
    n810_lo <= n4388;
    n822_lo <= n4391;
    n834_lo <= n4394;
    n846_lo <= n4397;
    n858_lo <= n4400;
    n870_lo <= n4403;
    n882_lo <= n4406;
    n894_lo <= n4409;
    n906_lo <= n4412;
    n918_lo <= n4415;
    n930_lo <= n4418;
    n942_lo <= n4421;
    n954_lo <= n4424;
    n966_lo <= n4427;
    n978_lo <= n4430;
    n990_lo <= n4433;
    n1002_lo <= n4436;
    n1005_lo <= n4439;
    n1008_lo <= n4442;
    n1017_lo <= n4445;
    n1020_lo <= n4448;
    n1029_lo <= n4451;
    n1032_lo <= n4454;
    n1041_lo <= n4457;
    n1044_lo <= n4460;
    n1053_lo <= n4463;
    n1056_lo <= n4466;
    n1065_lo <= n4469;
    n1068_lo <= n4472;
    n1077_lo <= n4475;
    n1080_lo <= n4478;
    n1089_lo <= n4481;
    n1092_lo <= n4484;
    n1101_lo <= n4487;
    n1104_lo <= n4490;
    n1837_o2 <= n4493;
    n1838_o2 <= n4496;
    n1839_o2 <= n4499;
    n1840_o2 <= n4502;
    n1841_o2 <= n4505;
    n1842_o2 <= n4508;
    n1843_o2 <= n4511;
    n1844_o2 <= n4514;
    n1845_o2 <= n4517;
    n1846_o2 <= n4520;
    n1847_o2 <= n4523;
    n1848_o2 <= n4526;
    n1849_o2 <= n4529;
    n1850_o2 <= n4532;
    n1851_o2 <= n4535;
    n1852_o2 <= n4538;
    n1853_o2 <= n4541;
    n1854_o2 <= n4544;
    n1855_o2 <= n4547;
    n1856_o2 <= n4550;
    n1857_o2 <= n4553;
    n1858_o2 <= n4556;
    n1859_o2 <= n4559;
    n1860_o2 <= n4562;
    n1861_o2 <= n4565;
    n1862_o2 <= n4568;
    n1863_o2 <= n4571;
    n1864_o2 <= n4574;
    n1865_o2 <= n4577;
    n1866_o2 <= n4580;
    n1867_o2 <= n4583;
    n1868_o2 <= n4586;
    G834_o2 <= n4589;
    G847_o2 <= n4592;
    G860_o2 <= n4595;
    G873_o2 <= n4598;
    G925_o2 <= n4601;
    G886_o2 <= n4604;
    G912_o2 <= n4607;
    G899_o2 <= n4610;
    n2151_o2 <= n4613;
    n2152_o2 <= n4616;
    n2153_o2 <= n4619;
    n2154_o2 <= n4622;
    n2155_o2 <= n4625;
    n2156_o2 <= n4628;
    n2157_o2 <= n4631;
    n2158_o2 <= n4634;
    n2159_o2 <= n4637;
    n2160_o2 <= n4640;
    n2161_o2 <= n4643;
    n2162_o2 <= n4646;
    n2163_o2 <= n4649;
    n2164_o2 <= n4652;
    n2165_o2 <= n4655;
    n2166_o2 <= n4658;
    n2167_o2 <= n4661;
    n2168_o2 <= n4664;
    n2169_o2 <= n4667;
    n2170_o2 <= n4670;
    n2171_o2 <= n4673;
    n2172_o2 <= n4676;
    n2173_o2 <= n4679;
    n2174_o2 <= n4682;
    n2175_o2 <= n4685;
    n2176_o2 <= n4688;
    n2177_o2 <= n4691;
    n2178_o2 <= n4694;
    n2179_o2 <= n4697;
    n2180_o2 <= n4700;
    n2181_o2 <= n4703;
    n2182_o2 <= n4706;
    G974_o2 <= n4709;
    G976_o2 <= n4712;
    G970_o2 <= n4715;
    G972_o2 <= n4718;
    G973_o2 <= n4721;
    G977_o2 <= n4724;
    G971_o2 <= n4727;
    G975_o2 <= n4730;
    G954_o2 <= n4733;
    G956_o2 <= n4736;
    G950_o2 <= n4739;
    G952_o2 <= n4742;
    G953_o2 <= n4745;
    G957_o2 <= n4748;
    G951_o2 <= n4751;
    G955_o2 <= n4754;
    G986_o2 <= n4757;
    G991_o2 <= n4760;
    G770_o2 <= n4763;
    G773_o2 <= n4766;
    G776_o2 <= n4769;
    G779_o2 <= n4772;
    G782_o2 <= n4775;
    G785_o2 <= n4778;
    G788_o2 <= n4781;
    G791_o2 <= n4784;
    G642_o2 <= n4787;
    G645_o2 <= n4790;
    G648_o2 <= n4793;
    G651_o2 <= n4796;
    G654_o2 <= n4799;
    G657_o2 <= n4802;
    G660_o2 <= n4805;
    G663_o2 <= n4808;
    G602_o2 <= n4811;
    G607_o2 <= n4814;
    G612_o2 <= n4817;
    G617_o2 <= n4820;
    G622_o2 <= n4823;
    G627_o2 <= n4826;
    G632_o2 <= n4829;
    G637_o2 <= n4832;
    n627_lo_buf_o2 <= n4835;
    n639_lo_buf_o2 <= n4838;
    n651_lo_buf_o2 <= n4841;
    n663_lo_buf_o2 <= n4844;
    n675_lo_buf_o2 <= n4847;
    n687_lo_buf_o2 <= n4850;
    n699_lo_buf_o2 <= n4853;
    n711_lo_buf_o2 <= n4856;
    n723_lo_buf_o2 <= n4859;
    n735_lo_buf_o2 <= n4862;
    n747_lo_buf_o2 <= n4865;
    n759_lo_buf_o2 <= n4868;
    n771_lo_buf_o2 <= n4871;
    n783_lo_buf_o2 <= n4874;
    n795_lo_buf_o2 <= n4877;
    n807_lo_buf_o2 <= n4880;
    n819_lo_buf_o2 <= n4883;
    n831_lo_buf_o2 <= n4886;
    n843_lo_buf_o2 <= n4889;
    n855_lo_buf_o2 <= n4892;
    n867_lo_buf_o2 <= n4895;
    n879_lo_buf_o2 <= n4898;
    n891_lo_buf_o2 <= n4901;
    n903_lo_buf_o2 <= n4904;
    n915_lo_buf_o2 <= n4907;
    n927_lo_buf_o2 <= n4910;
    n939_lo_buf_o2 <= n4913;
    n951_lo_buf_o2 <= n4916;
    n963_lo_buf_o2 <= n4919;
    n975_lo_buf_o2 <= n4922;
    n987_lo_buf_o2 <= n4925;
    n999_lo_buf_o2 <= n4928;
  end
  initial begin
    n630_lo <= 1'b0;
    n642_lo <= 1'b0;
    n654_lo <= 1'b0;
    n666_lo <= 1'b0;
    n678_lo <= 1'b0;
    n690_lo <= 1'b0;
    n702_lo <= 1'b0;
    n714_lo <= 1'b0;
    n726_lo <= 1'b0;
    n738_lo <= 1'b0;
    n750_lo <= 1'b0;
    n762_lo <= 1'b0;
    n774_lo <= 1'b0;
    n786_lo <= 1'b0;
    n798_lo <= 1'b0;
    n810_lo <= 1'b0;
    n822_lo <= 1'b0;
    n834_lo <= 1'b0;
    n846_lo <= 1'b0;
    n858_lo <= 1'b0;
    n870_lo <= 1'b0;
    n882_lo <= 1'b0;
    n894_lo <= 1'b0;
    n906_lo <= 1'b0;
    n918_lo <= 1'b0;
    n930_lo <= 1'b0;
    n942_lo <= 1'b0;
    n954_lo <= 1'b0;
    n966_lo <= 1'b0;
    n978_lo <= 1'b0;
    n990_lo <= 1'b0;
    n1002_lo <= 1'b0;
    n1005_lo <= 1'b0;
    n1008_lo <= 1'b0;
    n1017_lo <= 1'b0;
    n1020_lo <= 1'b0;
    n1029_lo <= 1'b0;
    n1032_lo <= 1'b0;
    n1041_lo <= 1'b0;
    n1044_lo <= 1'b0;
    n1053_lo <= 1'b0;
    n1056_lo <= 1'b0;
    n1065_lo <= 1'b0;
    n1068_lo <= 1'b0;
    n1077_lo <= 1'b0;
    n1080_lo <= 1'b0;
    n1089_lo <= 1'b0;
    n1092_lo <= 1'b0;
    n1101_lo <= 1'b0;
    n1104_lo <= 1'b0;
    n1837_o2 <= 1'b0;
    n1838_o2 <= 1'b0;
    n1839_o2 <= 1'b0;
    n1840_o2 <= 1'b0;
    n1841_o2 <= 1'b0;
    n1842_o2 <= 1'b0;
    n1843_o2 <= 1'b0;
    n1844_o2 <= 1'b0;
    n1845_o2 <= 1'b0;
    n1846_o2 <= 1'b0;
    n1847_o2 <= 1'b0;
    n1848_o2 <= 1'b0;
    n1849_o2 <= 1'b0;
    n1850_o2 <= 1'b0;
    n1851_o2 <= 1'b0;
    n1852_o2 <= 1'b0;
    n1853_o2 <= 1'b0;
    n1854_o2 <= 1'b0;
    n1855_o2 <= 1'b0;
    n1856_o2 <= 1'b0;
    n1857_o2 <= 1'b0;
    n1858_o2 <= 1'b0;
    n1859_o2 <= 1'b0;
    n1860_o2 <= 1'b0;
    n1861_o2 <= 1'b0;
    n1862_o2 <= 1'b0;
    n1863_o2 <= 1'b0;
    n1864_o2 <= 1'b0;
    n1865_o2 <= 1'b0;
    n1866_o2 <= 1'b0;
    n1867_o2 <= 1'b0;
    n1868_o2 <= 1'b0;
    G834_o2 <= 1'b0;
    G847_o2 <= 1'b0;
    G860_o2 <= 1'b0;
    G873_o2 <= 1'b0;
    G925_o2 <= 1'b0;
    G886_o2 <= 1'b0;
    G912_o2 <= 1'b0;
    G899_o2 <= 1'b0;
    n2151_o2 <= 1'b0;
    n2152_o2 <= 1'b0;
    n2153_o2 <= 1'b0;
    n2154_o2 <= 1'b0;
    n2155_o2 <= 1'b0;
    n2156_o2 <= 1'b0;
    n2157_o2 <= 1'b0;
    n2158_o2 <= 1'b0;
    n2159_o2 <= 1'b0;
    n2160_o2 <= 1'b0;
    n2161_o2 <= 1'b0;
    n2162_o2 <= 1'b0;
    n2163_o2 <= 1'b0;
    n2164_o2 <= 1'b0;
    n2165_o2 <= 1'b0;
    n2166_o2 <= 1'b0;
    n2167_o2 <= 1'b0;
    n2168_o2 <= 1'b0;
    n2169_o2 <= 1'b0;
    n2170_o2 <= 1'b0;
    n2171_o2 <= 1'b0;
    n2172_o2 <= 1'b0;
    n2173_o2 <= 1'b0;
    n2174_o2 <= 1'b0;
    n2175_o2 <= 1'b0;
    n2176_o2 <= 1'b0;
    n2177_o2 <= 1'b0;
    n2178_o2 <= 1'b0;
    n2179_o2 <= 1'b0;
    n2180_o2 <= 1'b0;
    n2181_o2 <= 1'b0;
    n2182_o2 <= 1'b0;
    G974_o2 <= 1'b0;
    G976_o2 <= 1'b0;
    G970_o2 <= 1'b0;
    G972_o2 <= 1'b0;
    G973_o2 <= 1'b0;
    G977_o2 <= 1'b0;
    G971_o2 <= 1'b0;
    G975_o2 <= 1'b0;
    G954_o2 <= 1'b0;
    G956_o2 <= 1'b0;
    G950_o2 <= 1'b0;
    G952_o2 <= 1'b0;
    G953_o2 <= 1'b0;
    G957_o2 <= 1'b0;
    G951_o2 <= 1'b0;
    G955_o2 <= 1'b0;
    G986_o2 <= 1'b0;
    G991_o2 <= 1'b0;
    G770_o2 <= 1'b0;
    G773_o2 <= 1'b0;
    G776_o2 <= 1'b0;
    G779_o2 <= 1'b0;
    G782_o2 <= 1'b0;
    G785_o2 <= 1'b0;
    G788_o2 <= 1'b0;
    G791_o2 <= 1'b0;
    G642_o2 <= 1'b0;
    G645_o2 <= 1'b0;
    G648_o2 <= 1'b0;
    G651_o2 <= 1'b0;
    G654_o2 <= 1'b0;
    G657_o2 <= 1'b0;
    G660_o2 <= 1'b0;
    G663_o2 <= 1'b0;
    G602_o2 <= 1'b0;
    G607_o2 <= 1'b0;
    G612_o2 <= 1'b0;
    G617_o2 <= 1'b0;
    G622_o2 <= 1'b0;
    G627_o2 <= 1'b0;
    G632_o2 <= 1'b0;
    G637_o2 <= 1'b0;
    n627_lo_buf_o2 <= 1'b0;
    n639_lo_buf_o2 <= 1'b0;
    n651_lo_buf_o2 <= 1'b0;
    n663_lo_buf_o2 <= 1'b0;
    n675_lo_buf_o2 <= 1'b0;
    n687_lo_buf_o2 <= 1'b0;
    n699_lo_buf_o2 <= 1'b0;
    n711_lo_buf_o2 <= 1'b0;
    n723_lo_buf_o2 <= 1'b0;
    n735_lo_buf_o2 <= 1'b0;
    n747_lo_buf_o2 <= 1'b0;
    n759_lo_buf_o2 <= 1'b0;
    n771_lo_buf_o2 <= 1'b0;
    n783_lo_buf_o2 <= 1'b0;
    n795_lo_buf_o2 <= 1'b0;
    n807_lo_buf_o2 <= 1'b0;
    n819_lo_buf_o2 <= 1'b0;
    n831_lo_buf_o2 <= 1'b0;
    n843_lo_buf_o2 <= 1'b0;
    n855_lo_buf_o2 <= 1'b0;
    n867_lo_buf_o2 <= 1'b0;
    n879_lo_buf_o2 <= 1'b0;
    n891_lo_buf_o2 <= 1'b0;
    n903_lo_buf_o2 <= 1'b0;
    n915_lo_buf_o2 <= 1'b0;
    n927_lo_buf_o2 <= 1'b0;
    n939_lo_buf_o2 <= 1'b0;
    n951_lo_buf_o2 <= 1'b0;
    n963_lo_buf_o2 <= 1'b0;
    n975_lo_buf_o2 <= 1'b0;
    n987_lo_buf_o2 <= 1'b0;
    n999_lo_buf_o2 <= 1'b0;
  end
endmodule


