
module mymod
(
  G1_p,
  G1_n,
  G2_p,
  G2_n,
  G3_p,
  G3_n,
  G4_p,
  G4_n,
  G5_p,
  G5_n,
  G6_p,
  G6_n,
  G7_p,
  G7_n,
  G8_p,
  G8_n,
  G9_p,
  G9_n,
  G10_p,
  G10_n,
  G11_p,
  G11_n,
  G12_p,
  G12_n,
  G13_p,
  G13_n,
  G14_p,
  G14_n,
  G15_p,
  G15_n,
  G16_p,
  G16_n,
  G17_p,
  G17_n,
  G18_p,
  G18_n,
  G19_p,
  G19_n,
  G20_p,
  G20_n,
  G21_p,
  G21_n,
  G22_p,
  G22_n,
  G23_p,
  G23_n,
  G24_p,
  G24_n,
  G25_p,
  G25_n,
  G26_p,
  G26_n,
  G27_p,
  G27_n,
  G28_p,
  G28_n,
  G29_p,
  G29_n,
  G30_p,
  G30_n,
  G31_p,
  G31_n,
  G32_p,
  G32_n,
  G33_p,
  G33_n,
  G34_p,
  G34_n,
  G35_p,
  G35_n,
  G36_p,
  G36_n,
  G37_p,
  G37_n,
  G38_p,
  G38_n,
  G39_p,
  G39_n,
  G40_p,
  G40_n,
  G41_p,
  G41_n,
  G42_p,
  G42_n,
  G43_p,
  G43_n,
  G44_p,
  G44_n,
  G45_p,
  G45_n,
  G46_p,
  G46_n,
  G47_p,
  G47_n,
  G48_p,
  G48_n,
  G49_p,
  G49_n,
  G50_p,
  G50_n,
  G51_p,
  G51_n,
  G52_p,
  G52_n,
  G53_p,
  G53_n,
  G54_p,
  G54_n,
  G55_p,
  G55_n,
  G56_p,
  G56_n,
  G57_p,
  G57_n,
  G58_p,
  G58_n,
  G59_p,
  G59_n,
  G60_p,
  G60_n,
  G61_p,
  G61_n,
  G62_p,
  G62_n,
  G63_p,
  G63_n,
  G64_p,
  G64_n,
  G65_p,
  G65_n,
  G66_p,
  G66_n,
  G67_p,
  G67_n,
  G68_p,
  G68_n,
  G69_p,
  G69_n,
  G70_p,
  G70_n,
  G71_p,
  G71_n,
  G72_p,
  G72_n,
  G73_p,
  G73_n,
  G74_p,
  G74_n,
  G75_p,
  G75_n,
  G76_p,
  G76_n,
  G77_p,
  G77_n,
  G78_p,
  G78_n,
  G79_p,
  G79_n,
  G80_p,
  G80_n,
  G81_p,
  G81_n,
  G82_p,
  G82_n,
  G83_p,
  G83_n,
  G84_p,
  G84_n,
  G85_p,
  G85_n,
  G86_p,
  G86_n,
  G87_p,
  G87_n,
  G88_p,
  G88_n,
  G89_p,
  G89_n,
  G90_p,
  G90_n,
  G91_p,
  G91_n,
  G92_p,
  G92_n,
  G93_p,
  G93_n,
  G94_p,
  G94_n,
  G95_p,
  G95_n,
  G96_p,
  G96_n,
  G97_p,
  G97_n,
  G98_p,
  G98_n,
  G99_p,
  G99_n,
  G100_p,
  G100_n,
  G101_p,
  G101_n,
  G102_p,
  G102_n,
  G103_p,
  G103_n,
  G104_p,
  G104_n,
  G105_p,
  G105_n,
  G106_p,
  G106_n,
  G107_p,
  G107_n,
  G108_p,
  G108_n,
  G109_p,
  G109_n,
  G110_p,
  G110_n,
  G111_p,
  G111_n,
  G112_p,
  G112_n,
  G113_p,
  G113_n,
  G114_p,
  G114_n,
  G115_p,
  G115_n,
  G116_p,
  G116_n,
  G117_p,
  G117_n,
  G118_p,
  G118_n,
  G119_p,
  G119_n,
  G120_p,
  G120_n,
  G121_p,
  G121_n,
  G122_p,
  G122_n,
  G123_p,
  G123_n,
  G124_p,
  G124_n,
  G125_p,
  G125_n,
  G126_p,
  G126_n,
  G127_p,
  G127_n,
  G128_p,
  G128_n,
  G129_p,
  G129_n,
  G130_p,
  G130_n,
  G131_p,
  G131_n,
  G132_p,
  G132_n,
  G133_p,
  G133_n,
  G134_p,
  G134_n,
  G135_p,
  G135_n,
  G136_p,
  G136_n,
  G137_p,
  G137_n,
  G138_p,
  G138_n,
  G139_p,
  G139_n,
  G140_p,
  G140_n,
  G141_p,
  G141_n,
  G142_p,
  G142_n,
  G143_p,
  G143_n,
  G144_p,
  G144_n,
  G145_p,
  G145_n,
  G146_p,
  G146_n,
  G147_p,
  G147_n,
  G148_p,
  G148_n,
  G149_p,
  G149_n,
  G150_p,
  G150_n,
  G151_p,
  G151_n,
  G152_p,
  G152_n,
  G153_p,
  G153_n,
  G154_p,
  G154_n,
  G155_p,
  G155_n,
  G156_p,
  G156_n,
  G157_p,
  G157_n,
  G2531_p,
  G2532_p,
  G2533_p,
  G2534_p,
  G2535_p,
  G2536_p,
  G2537_p,
  G2538_p,
  G2539_p,
  G2540_p,
  G2541_p,
  G2542_p,
  G2543_p,
  G2544_p,
  G2545_p,
  G2546_p,
  G2547_p,
  G2548_p,
  G2549_p,
  G2550_p,
  G2551_p,
  G2552_p,
  G2553_p,
  G2554_p,
  G2555_p,
  G2556_p,
  G2557_p,
  G2558_p,
  G2559_p,
  G2560_p,
  G2561_n,
  G2562_p,
  G2563_p,
  G2564_p,
  G2565_p,
  G2566_p,
  G2567_p,
  G2568_p,
  G2569_p,
  G2570_p,
  G2571_p,
  G2572_p,
  G2573_p,
  G2574_p,
  G2575_n,
  G2576_n,
  G2577_p,
  G2578_p,
  G2579_p,
  G2580_p,
  G2581_n,
  G2582_p,
  G2583_p,
  G2584_p,
  G2585_p,
  G2586_p,
  G2587_n,
  G2588_p,
  G2589_p,
  G2590_n,
  G2591_p,
  G2592_p,
  G2593_p,
  G2594_p
);

  input G1_p;input G1_n;input G2_p;input G2_n;input G3_p;input G3_n;input G4_p;input G4_n;input G5_p;input G5_n;input G6_p;input G6_n;input G7_p;input G7_n;input G8_p;input G8_n;input G9_p;input G9_n;input G10_p;input G10_n;input G11_p;input G11_n;input G12_p;input G12_n;input G13_p;input G13_n;input G14_p;input G14_n;input G15_p;input G15_n;input G16_p;input G16_n;input G17_p;input G17_n;input G18_p;input G18_n;input G19_p;input G19_n;input G20_p;input G20_n;input G21_p;input G21_n;input G22_p;input G22_n;input G23_p;input G23_n;input G24_p;input G24_n;input G25_p;input G25_n;input G26_p;input G26_n;input G27_p;input G27_n;input G28_p;input G28_n;input G29_p;input G29_n;input G30_p;input G30_n;input G31_p;input G31_n;input G32_p;input G32_n;input G33_p;input G33_n;input G34_p;input G34_n;input G35_p;input G35_n;input G36_p;input G36_n;input G37_p;input G37_n;input G38_p;input G38_n;input G39_p;input G39_n;input G40_p;input G40_n;input G41_p;input G41_n;input G42_p;input G42_n;input G43_p;input G43_n;input G44_p;input G44_n;input G45_p;input G45_n;input G46_p;input G46_n;input G47_p;input G47_n;input G48_p;input G48_n;input G49_p;input G49_n;input G50_p;input G50_n;input G51_p;input G51_n;input G52_p;input G52_n;input G53_p;input G53_n;input G54_p;input G54_n;input G55_p;input G55_n;input G56_p;input G56_n;input G57_p;input G57_n;input G58_p;input G58_n;input G59_p;input G59_n;input G60_p;input G60_n;input G61_p;input G61_n;input G62_p;input G62_n;input G63_p;input G63_n;input G64_p;input G64_n;input G65_p;input G65_n;input G66_p;input G66_n;input G67_p;input G67_n;input G68_p;input G68_n;input G69_p;input G69_n;input G70_p;input G70_n;input G71_p;input G71_n;input G72_p;input G72_n;input G73_p;input G73_n;input G74_p;input G74_n;input G75_p;input G75_n;input G76_p;input G76_n;input G77_p;input G77_n;input G78_p;input G78_n;input G79_p;input G79_n;input G80_p;input G80_n;input G81_p;input G81_n;input G82_p;input G82_n;input G83_p;input G83_n;input G84_p;input G84_n;input G85_p;input G85_n;input G86_p;input G86_n;input G87_p;input G87_n;input G88_p;input G88_n;input G89_p;input G89_n;input G90_p;input G90_n;input G91_p;input G91_n;input G92_p;input G92_n;input G93_p;input G93_n;input G94_p;input G94_n;input G95_p;input G95_n;input G96_p;input G96_n;input G97_p;input G97_n;input G98_p;input G98_n;input G99_p;input G99_n;input G100_p;input G100_n;input G101_p;input G101_n;input G102_p;input G102_n;input G103_p;input G103_n;input G104_p;input G104_n;input G105_p;input G105_n;input G106_p;input G106_n;input G107_p;input G107_n;input G108_p;input G108_n;input G109_p;input G109_n;input G110_p;input G110_n;input G111_p;input G111_n;input G112_p;input G112_n;input G113_p;input G113_n;input G114_p;input G114_n;input G115_p;input G115_n;input G116_p;input G116_n;input G117_p;input G117_n;input G118_p;input G118_n;input G119_p;input G119_n;input G120_p;input G120_n;input G121_p;input G121_n;input G122_p;input G122_n;input G123_p;input G123_n;input G124_p;input G124_n;input G125_p;input G125_n;input G126_p;input G126_n;input G127_p;input G127_n;input G128_p;input G128_n;input G129_p;input G129_n;input G130_p;input G130_n;input G131_p;input G131_n;input G132_p;input G132_n;input G133_p;input G133_n;input G134_p;input G134_n;input G135_p;input G135_n;input G136_p;input G136_n;input G137_p;input G137_n;input G138_p;input G138_n;input G139_p;input G139_n;input G140_p;input G140_n;input G141_p;input G141_n;input G142_p;input G142_n;input G143_p;input G143_n;input G144_p;input G144_n;input G145_p;input G145_n;input G146_p;input G146_n;input G147_p;input G147_n;input G148_p;input G148_n;input G149_p;input G149_n;input G150_p;input G150_n;input G151_p;input G151_n;input G152_p;input G152_n;input G153_p;input G153_n;input G154_p;input G154_n;input G155_p;input G155_n;input G156_p;input G156_n;input G157_p;input G157_n;
  output G2531_p;output G2532_p;output G2533_p;output G2534_p;output G2535_p;output G2536_p;output G2537_p;output G2538_p;output G2539_p;output G2540_p;output G2541_p;output G2542_p;output G2543_p;output G2544_p;output G2545_p;output G2546_p;output G2547_p;output G2548_p;output G2549_p;output G2550_p;output G2551_p;output G2552_p;output G2553_p;output G2554_p;output G2555_p;output G2556_p;output G2557_p;output G2558_p;output G2559_p;output G2560_p;output G2561_n;output G2562_p;output G2563_p;output G2564_p;output G2565_p;output G2566_p;output G2567_p;output G2568_p;output G2569_p;output G2570_p;output G2571_p;output G2572_p;output G2573_p;output G2574_p;output G2575_n;output G2576_n;output G2577_p;output G2578_p;output G2579_p;output G2580_p;output G2581_n;output G2582_p;output G2583_p;output G2584_p;output G2585_p;output G2586_p;output G2587_n;output G2588_p;output G2589_p;output G2590_n;output G2591_p;output G2592_p;output G2593_p;output G2594_p;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire G51_p;
  wire G51_n;
  wire G52_p;
  wire G52_n;
  wire G53_p;
  wire G53_n;
  wire G54_p;
  wire G54_n;
  wire G55_p;
  wire G55_n;
  wire G56_p;
  wire G56_n;
  wire G57_p;
  wire G57_n;
  wire G58_p;
  wire G58_n;
  wire G59_p;
  wire G59_n;
  wire G60_p;
  wire G60_n;
  wire G61_p;
  wire G61_n;
  wire G62_p;
  wire G62_n;
  wire G63_p;
  wire G63_n;
  wire G64_p;
  wire G64_n;
  wire G65_p;
  wire G65_n;
  wire G66_p;
  wire G66_n;
  wire G67_p;
  wire G67_n;
  wire G68_p;
  wire G68_n;
  wire G69_p;
  wire G69_n;
  wire G70_p;
  wire G70_n;
  wire G71_p;
  wire G71_n;
  wire G72_p;
  wire G72_n;
  wire G73_p;
  wire G73_n;
  wire G74_p;
  wire G74_n;
  wire G75_p;
  wire G75_n;
  wire G76_p;
  wire G76_n;
  wire G77_p;
  wire G77_n;
  wire G78_p;
  wire G78_n;
  wire G79_p;
  wire G79_n;
  wire G80_p;
  wire G80_n;
  wire G81_p;
  wire G81_n;
  wire G82_p;
  wire G82_n;
  wire G83_p;
  wire G83_n;
  wire G84_p;
  wire G84_n;
  wire G85_p;
  wire G85_n;
  wire G86_p;
  wire G86_n;
  wire G87_p;
  wire G87_n;
  wire G88_p;
  wire G88_n;
  wire G89_p;
  wire G89_n;
  wire G90_p;
  wire G90_n;
  wire G91_p;
  wire G91_n;
  wire G92_p;
  wire G92_n;
  wire G93_p;
  wire G93_n;
  wire G94_p;
  wire G94_n;
  wire G95_p;
  wire G95_n;
  wire G96_p;
  wire G96_n;
  wire G97_p;
  wire G97_n;
  wire G98_p;
  wire G98_n;
  wire G99_p;
  wire G99_n;
  wire G100_p;
  wire G100_n;
  wire G101_p;
  wire G101_n;
  wire G102_p;
  wire G102_n;
  wire G103_p;
  wire G103_n;
  wire G104_p;
  wire G104_n;
  wire G105_p;
  wire G105_n;
  wire G106_p;
  wire G106_n;
  wire G107_p;
  wire G107_n;
  wire G108_p;
  wire G108_n;
  wire G109_p;
  wire G109_n;
  wire G110_p;
  wire G110_n;
  wire G111_p;
  wire G111_n;
  wire G112_p;
  wire G112_n;
  wire G113_p;
  wire G113_n;
  wire G114_p;
  wire G114_n;
  wire G115_p;
  wire G115_n;
  wire G116_p;
  wire G116_n;
  wire G117_p;
  wire G117_n;
  wire G118_p;
  wire G118_n;
  wire G119_p;
  wire G119_n;
  wire G120_p;
  wire G120_n;
  wire G121_p;
  wire G121_n;
  wire G122_p;
  wire G122_n;
  wire G123_p;
  wire G123_n;
  wire G124_p;
  wire G124_n;
  wire G125_p;
  wire G125_n;
  wire G126_p;
  wire G126_n;
  wire G127_p;
  wire G127_n;
  wire G128_p;
  wire G128_n;
  wire G129_p;
  wire G129_n;
  wire G130_p;
  wire G130_n;
  wire G131_p;
  wire G131_n;
  wire G132_p;
  wire G132_n;
  wire G133_p;
  wire G133_n;
  wire G134_p;
  wire G134_n;
  wire G135_p;
  wire G135_n;
  wire G136_p;
  wire G136_n;
  wire G137_p;
  wire G137_n;
  wire G138_p;
  wire G138_n;
  wire G139_p;
  wire G139_n;
  wire G140_p;
  wire G140_n;
  wire G141_p;
  wire G141_n;
  wire G142_p;
  wire G142_n;
  wire G143_p;
  wire G143_n;
  wire G144_p;
  wire G144_n;
  wire G145_p;
  wire G145_n;
  wire G146_p;
  wire G146_n;
  wire G147_p;
  wire G147_n;
  wire G148_p;
  wire G148_n;
  wire G149_p;
  wire G149_n;
  wire G150_p;
  wire G150_n;
  wire G151_p;
  wire G151_n;
  wire G152_p;
  wire G152_n;
  wire G153_p;
  wire G153_n;
  wire G154_p;
  wire G154_n;
  wire G155_p;
  wire G155_n;
  wire G156_p;
  wire G156_n;
  wire G157_p;
  wire G157_n;
  wire ffc_0_p;
  wire ffc_0_n;
  wire ffc_1_p;
  wire ffc_1_n;
  wire ffc_2_p;
  wire ffc_2_n;
  wire ffc_3_p;
  wire ffc_3_n;
  wire ffc_4_p;
  wire ffc_4_n;
  wire ffc_5_p;
  wire ffc_5_n;
  wire ffc_6_p;
  wire ffc_6_n;
  wire ffc_7_p;
  wire ffc_7_n;
  wire ffc_8_p;
  wire ffc_8_n;
  wire ffc_9_p;
  wire ffc_9_n;
  wire ffc_10_p;
  wire ffc_10_n;
  wire ffc_11_p;
  wire ffc_11_n;
  wire ffc_12_p;
  wire ffc_12_n;
  wire ffc_13_p;
  wire ffc_13_n;
  wire ffc_14_p;
  wire ffc_14_n;
  wire ffc_15_p;
  wire ffc_15_n;
  wire ffc_16_p;
  wire ffc_16_n;
  wire ffc_17_p;
  wire ffc_17_n;
  wire ffc_18_p;
  wire ffc_18_n;
  wire ffc_19_p;
  wire ffc_19_n;
  wire ffc_20_p;
  wire ffc_20_n;
  wire ffc_21_p;
  wire ffc_21_n;
  wire ffc_22_p;
  wire ffc_22_n;
  wire ffc_23_p;
  wire ffc_23_n;
  wire ffc_24_p;
  wire ffc_24_n;
  wire ffc_25_p;
  wire ffc_25_n;
  wire ffc_26_p;
  wire ffc_26_n;
  wire ffc_27_p;
  wire ffc_27_n;
  wire ffc_28_p;
  wire ffc_28_n;
  wire ffc_29_p;
  wire ffc_29_n;
  wire ffc_30_p;
  wire ffc_30_n;
  wire ffc_31_p;
  wire ffc_31_n;
  wire ffc_32_p;
  wire ffc_32_n;
  wire ffc_33_p;
  wire ffc_33_n;
  wire ffc_34_p;
  wire ffc_34_n;
  wire ffc_35_p;
  wire ffc_35_n;
  wire ffc_36_p;
  wire ffc_36_n;
  wire ffc_37_p;
  wire ffc_37_n;
  wire ffc_38_p;
  wire ffc_38_n;
  wire ffc_39_p;
  wire ffc_39_n;
  wire ffc_40_p;
  wire ffc_40_n;
  wire ffc_41_p;
  wire ffc_41_n;
  wire ffc_42_p;
  wire ffc_42_n;
  wire ffc_43_p;
  wire ffc_43_n;
  wire ffc_44_p;
  wire ffc_44_n;
  wire ffc_45_p;
  wire ffc_45_n;
  wire ffc_46_p;
  wire ffc_46_n;
  wire ffc_47_p;
  wire ffc_47_n;
  wire ffc_48_p;
  wire ffc_48_n;
  wire ffc_49_p;
  wire ffc_49_n;
  wire ffc_50_p;
  wire ffc_50_n;
  wire ffc_51_p;
  wire ffc_51_n;
  wire ffc_52_p;
  wire ffc_52_n;
  wire ffc_53_p;
  wire ffc_53_n;
  wire ffc_54_p;
  wire ffc_54_n;
  wire ffc_55_p;
  wire ffc_55_n;
  wire ffc_56_p;
  wire ffc_56_n;
  wire ffc_57_p;
  wire ffc_57_n;
  wire ffc_58_p;
  wire ffc_58_n;
  wire ffc_59_p;
  wire ffc_59_n;
  wire ffc_60_p;
  wire ffc_60_n;
  wire ffc_61_p;
  wire ffc_61_n;
  wire ffc_62_p;
  wire ffc_62_n;
  wire ffc_63_p;
  wire ffc_63_n;
  wire ffc_64_p;
  wire ffc_64_n;
  wire ffc_65_p;
  wire ffc_65_n;
  wire ffc_66_p;
  wire ffc_66_n;
  wire ffc_67_p;
  wire ffc_67_n;
  wire ffc_68_p;
  wire ffc_68_n;
  wire ffc_69_p;
  wire ffc_69_n;
  wire ffc_70_p;
  wire ffc_70_n;
  wire ffc_71_p;
  wire ffc_71_n;
  wire ffc_72_p;
  wire ffc_72_n;
  wire ffc_73_p;
  wire ffc_73_n;
  wire ffc_74_p;
  wire ffc_74_n;
  wire ffc_75_p;
  wire ffc_75_n;
  wire ffc_76_p;
  wire ffc_76_n;
  wire ffc_77_p;
  wire ffc_77_n;
  wire ffc_78_p;
  wire ffc_78_n;
  wire ffc_79_p;
  wire ffc_79_n;
  wire ffc_80_p;
  wire ffc_80_n;
  wire ffc_81_p;
  wire ffc_81_n;
  wire ffc_82_p;
  wire ffc_82_n;
  wire ffc_83_p;
  wire ffc_83_n;
  wire ffc_84_p;
  wire ffc_84_n;
  wire ffc_85_p;
  wire ffc_85_n;
  wire ffc_86_p;
  wire ffc_86_n;
  wire ffc_87_p;
  wire ffc_87_n;
  wire ffc_88_p;
  wire ffc_88_n;
  wire ffc_89_p;
  wire ffc_89_n;
  wire ffc_90_p;
  wire ffc_90_n;
  wire ffc_91_p;
  wire ffc_91_n;
  wire ffc_92_p;
  wire ffc_92_n;
  wire ffc_93_p;
  wire ffc_93_n;
  wire ffc_94_p;
  wire ffc_94_n;
  wire ffc_95_p;
  wire ffc_95_n;
  wire ffc_96_p;
  wire ffc_96_n;
  wire ffc_97_p;
  wire ffc_97_n;
  wire ffc_98_p;
  wire ffc_98_n;
  wire ffc_99_p;
  wire ffc_99_n;
  wire ffc_100_p;
  wire ffc_100_n;
  wire ffc_101_p;
  wire ffc_101_n;
  wire ffc_102_p;
  wire ffc_102_n;
  wire ffc_103_p;
  wire ffc_103_n;
  wire ffc_104_p;
  wire ffc_104_n;
  wire ffc_105_p;
  wire ffc_105_n;
  wire ffc_106_p;
  wire ffc_106_n;
  wire ffc_107_p;
  wire ffc_107_n;
  wire ffc_108_p;
  wire ffc_108_n;
  wire ffc_109_p;
  wire ffc_109_n;
  wire ffc_110_p;
  wire ffc_110_n;
  wire ffc_111_p;
  wire ffc_111_n;
  wire ffc_112_p;
  wire ffc_112_n;
  wire ffc_113_p;
  wire ffc_113_n;
  wire ffc_114_p;
  wire ffc_114_n;
  wire ffc_115_p;
  wire ffc_115_n;
  wire ffc_116_p;
  wire ffc_116_n;
  wire ffc_117_p;
  wire ffc_117_n;
  wire ffc_118_p;
  wire ffc_118_n;
  wire ffc_119_p;
  wire ffc_119_n;
  wire ffc_120_p;
  wire ffc_120_n;
  wire ffc_121_p;
  wire ffc_121_n;
  wire ffc_122_p;
  wire ffc_122_n;
  wire ffc_123_p;
  wire ffc_123_n;
  wire ffc_124_p;
  wire ffc_124_n;
  wire ffc_125_p;
  wire ffc_125_n;
  wire ffc_126_p;
  wire ffc_126_n;
  wire ffc_127_p;
  wire ffc_127_n;
  wire ffc_128_p;
  wire ffc_128_n;
  wire ffc_129_p;
  wire ffc_129_n;
  wire ffc_130_p;
  wire ffc_130_n;
  wire ffc_131_p;
  wire ffc_131_n;
  wire ffc_132_p;
  wire ffc_132_n;
  wire ffc_133_p;
  wire ffc_133_n;
  wire ffc_134_p;
  wire ffc_134_n;
  wire ffc_135_p;
  wire ffc_135_n;
  wire ffc_136_p;
  wire ffc_136_n;
  wire ffc_137_p;
  wire ffc_137_n;
  wire ffc_138_p;
  wire ffc_138_n;
  wire ffc_139_p;
  wire ffc_139_n;
  wire ffc_140_p;
  wire ffc_140_n;
  wire ffc_141_p;
  wire ffc_141_n;
  wire ffc_142_p;
  wire ffc_142_n;
  wire ffc_143_p;
  wire ffc_143_n;
  wire ffc_144_p;
  wire ffc_144_n;
  wire ffc_145_p;
  wire ffc_145_n;
  wire ffc_146_p;
  wire ffc_146_n;
  wire ffc_147_p;
  wire ffc_147_n;
  wire ffc_148_p;
  wire ffc_148_n;
  wire ffc_149_p;
  wire ffc_149_n;
  wire ffc_150_p;
  wire ffc_150_n;
  wire ffc_151_p;
  wire ffc_151_n;
  wire ffc_152_p;
  wire ffc_152_n;
  wire ffc_153_p;
  wire ffc_153_n;
  wire ffc_154_p;
  wire ffc_154_n;
  wire ffc_155_p;
  wire ffc_155_n;
  wire ffc_156_p;
  wire ffc_156_n;
  wire ffc_157_p;
  wire ffc_157_n;
  wire ffc_158_p;
  wire ffc_158_n;
  wire ffc_159_p;
  wire ffc_159_n;
  wire ffc_160_p;
  wire ffc_160_n;
  wire ffc_161_p;
  wire ffc_161_n;
  wire ffc_162_p;
  wire ffc_162_n;
  wire ffc_163_p;
  wire ffc_163_n;
  wire ffc_164_p;
  wire ffc_164_n;
  wire ffc_165_p;
  wire ffc_165_n;
  wire ffc_166_p;
  wire ffc_166_n;
  wire ffc_167_p;
  wire ffc_167_n;
  wire ffc_168_p;
  wire ffc_168_n;
  wire ffc_169_p;
  wire ffc_169_n;
  wire ffc_170_p;
  wire ffc_170_n;
  wire ffc_171_p;
  wire ffc_171_n;
  wire ffc_172_p;
  wire ffc_172_n;
  wire ffc_173_p;
  wire ffc_173_n;
  wire ffc_174_p;
  wire ffc_174_n;
  wire ffc_175_p;
  wire ffc_175_n;
  wire ffc_176_p;
  wire ffc_176_n;
  wire ffc_177_p;
  wire ffc_177_n;
  wire ffc_178_p;
  wire ffc_178_n;
  wire ffc_179_p;
  wire ffc_179_n;
  wire ffc_180_p;
  wire ffc_180_n;
  wire ffc_181_p;
  wire ffc_181_n;
  wire ffc_182_p;
  wire ffc_182_n;
  wire ffc_183_p;
  wire ffc_183_n;
  wire ffc_184_p;
  wire ffc_184_n;
  wire ffc_185_p;
  wire ffc_185_n;
  wire ffc_186_p;
  wire ffc_186_n;
  wire ffc_187_p;
  wire ffc_187_n;
  wire ffc_188_p;
  wire ffc_188_n;
  wire ffc_189_p;
  wire ffc_189_n;
  wire ffc_190_p;
  wire ffc_190_n;
  wire ffc_191_p;
  wire ffc_191_n;
  wire ffc_192_p;
  wire ffc_192_n;
  wire ffc_193_p;
  wire ffc_193_n;
  wire ffc_194_p;
  wire ffc_194_n;
  wire ffc_195_p;
  wire ffc_195_n;
  wire ffc_196_p;
  wire ffc_196_n;
  wire ffc_197_p;
  wire ffc_197_n;
  wire ffc_198_p;
  wire ffc_198_n;
  wire ffc_199_p;
  wire ffc_199_n;
  wire ffc_200_p;
  wire ffc_200_n;
  wire ffc_201_p;
  wire ffc_201_n;
  wire ffc_202_p;
  wire ffc_202_n;
  wire ffc_203_p;
  wire ffc_203_n;
  wire ffc_204_p;
  wire ffc_204_n;
  wire ffc_205_p;
  wire ffc_205_n;
  wire ffc_206_p;
  wire ffc_206_n;
  wire ffc_207_p;
  wire ffc_207_n;
  wire ffc_208_p;
  wire ffc_208_n;
  wire ffc_209_p;
  wire ffc_209_n;
  wire ffc_210_p;
  wire ffc_210_n;
  wire ffc_211_p;
  wire ffc_211_n;
  wire ffc_212_p;
  wire ffc_212_n;
  wire ffc_213_p;
  wire ffc_213_n;
  wire ffc_214_p;
  wire ffc_214_n;
  wire ffc_215_p;
  wire ffc_215_n;
  wire ffc_216_p;
  wire ffc_216_n;
  wire ffc_217_p;
  wire ffc_217_n;
  wire ffc_218_p;
  wire ffc_218_n;
  wire ffc_219_p;
  wire ffc_219_n;
  wire ffc_220_p;
  wire ffc_220_n;
  wire ffc_221_p;
  wire ffc_221_n;
  wire ffc_222_p;
  wire ffc_222_n;
  wire ffc_223_p;
  wire ffc_223_n;
  wire ffc_224_p;
  wire ffc_224_n;
  wire ffc_225_p;
  wire ffc_225_n;
  wire ffc_226_p;
  wire ffc_226_n;
  wire ffc_227_p;
  wire ffc_227_n;
  wire ffc_228_p;
  wire ffc_228_n;
  wire ffc_229_p;
  wire ffc_229_n;
  wire ffc_230_p;
  wire ffc_230_n;
  wire ffc_231_p;
  wire ffc_231_n;
  wire ffc_232_p;
  wire ffc_232_n;
  wire ffc_233_p;
  wire ffc_233_n;
  wire ffc_234_p;
  wire ffc_234_n;
  wire ffc_235_p;
  wire ffc_235_n;
  wire ffc_236_p;
  wire ffc_236_n;
  wire ffc_237_p;
  wire ffc_237_n;
  wire ffc_238_p;
  wire ffc_238_n;
  wire ffc_239_p;
  wire ffc_239_n;
  wire ffc_240_p;
  wire ffc_240_n;
  wire ffc_241_p;
  wire ffc_241_n;
  wire ffc_242_p;
  wire ffc_242_n;
  wire ffc_243_p;
  wire ffc_243_n;
  wire ffc_244_p;
  wire ffc_244_n;
  wire ffc_245_p;
  wire ffc_245_n;
  wire ffc_246_p;
  wire ffc_246_n;
  wire ffc_247_p;
  wire ffc_247_n;
  wire ffc_248_p;
  wire ffc_248_n;
  wire ffc_249_p;
  wire ffc_249_n;
  wire ffc_250_p;
  wire ffc_250_n;
  wire ffc_251_p;
  wire ffc_251_n;
  wire ffc_252_p;
  wire ffc_252_n;
  wire ffc_253_p;
  wire ffc_253_n;
  wire ffc_254_p;
  wire ffc_254_n;
  wire ffc_255_p;
  wire ffc_255_n;
  wire ffc_256_p;
  wire ffc_256_n;
  wire ffc_257_p;
  wire ffc_257_n;
  wire ffc_258_p;
  wire ffc_258_n;
  wire ffc_259_p;
  wire ffc_259_n;
  wire ffc_260_p;
  wire ffc_260_n;
  wire ffc_261_p;
  wire ffc_261_n;
  wire ffc_262_p;
  wire ffc_262_n;
  wire ffc_263_p;
  wire ffc_263_n;
  wire ffc_264_p;
  wire ffc_264_n;
  wire ffc_265_p;
  wire ffc_265_n;
  wire ffc_266_p;
  wire ffc_266_n;
  wire ffc_267_p;
  wire ffc_267_n;
  wire ffc_268_p;
  wire ffc_268_n;
  wire ffc_269_p;
  wire ffc_269_n;
  wire ffc_270_p;
  wire ffc_270_n;
  wire ffc_271_p;
  wire ffc_271_n;
  wire ffc_272_p;
  wire ffc_272_n;
  wire ffc_273_p;
  wire ffc_273_n;
  wire ffc_274_p;
  wire ffc_274_n;
  wire ffc_275_p;
  wire ffc_275_n;
  wire ffc_276_p;
  wire ffc_276_n;
  wire ffc_277_p;
  wire ffc_277_n;
  wire ffc_278_p;
  wire ffc_278_n;
  wire ffc_279_p;
  wire ffc_279_n;
  wire ffc_280_p;
  wire ffc_280_n;
  wire ffc_281_p;
  wire ffc_281_n;
  wire ffc_282_p;
  wire ffc_282_n;
  wire ffc_283_p;
  wire ffc_283_n;
  wire ffc_284_p;
  wire ffc_284_n;
  wire ffc_285_p;
  wire ffc_285_n;
  wire ffc_286_p;
  wire ffc_286_n;
  wire ffc_287_p;
  wire ffc_287_n;
  wire ffc_288_p;
  wire ffc_288_n;
  wire ffc_289_p;
  wire ffc_289_n;
  wire ffc_290_p;
  wire ffc_290_n;
  wire ffc_291_p;
  wire ffc_291_n;
  wire ffc_292_p;
  wire ffc_292_n;
  wire ffc_293_p;
  wire ffc_293_n;
  wire ffc_294_p;
  wire ffc_294_n;
  wire ffc_295_p;
  wire ffc_295_n;
  wire ffc_296_p;
  wire ffc_296_n;
  wire ffc_297_p;
  wire ffc_297_n;
  wire ffc_298_p;
  wire ffc_298_n;
  wire ffc_299_p;
  wire ffc_299_n;
  wire ffc_300_p;
  wire ffc_300_n;
  wire ffc_301_p;
  wire ffc_301_n;
  wire ffc_302_p;
  wire ffc_302_n;
  wire ffc_303_p;
  wire ffc_303_n;
  wire ffc_304_p;
  wire ffc_304_n;
  wire ffc_305_p;
  wire ffc_305_n;
  wire ffc_306_p;
  wire ffc_306_n;
  wire ffc_307_p;
  wire ffc_307_n;
  wire ffc_308_p;
  wire ffc_308_n;
  wire ffc_309_p;
  wire ffc_309_n;
  wire ffc_310_p;
  wire ffc_310_n;
  wire ffc_311_p;
  wire ffc_311_n;
  wire ffc_312_p;
  wire ffc_312_n;
  wire ffc_313_p;
  wire ffc_313_n;
  wire ffc_314_p;
  wire ffc_314_n;
  wire ffc_315_p;
  wire ffc_315_n;
  wire ffc_316_p;
  wire ffc_316_n;
  wire ffc_317_p;
  wire ffc_317_n;
  wire ffc_318_p;
  wire ffc_318_n;
  wire ffc_319_p;
  wire ffc_319_n;
  wire ffc_320_p;
  wire ffc_320_n;
  wire ffc_321_p;
  wire ffc_321_n;
  wire ffc_322_p;
  wire ffc_322_n;
  wire ffc_323_p;
  wire ffc_323_n;
  wire ffc_324_p;
  wire ffc_324_n;
  wire ffc_325_p;
  wire ffc_325_n;
  wire ffc_326_p;
  wire ffc_326_n;
  wire ffc_327_p;
  wire ffc_327_n;
  wire ffc_328_p;
  wire ffc_328_n;
  wire ffc_329_p;
  wire ffc_329_n;
  wire ffc_330_p;
  wire ffc_330_n;
  wire ffc_331_p;
  wire ffc_331_n;
  wire ffc_332_p;
  wire ffc_332_n;
  wire ffc_333_p;
  wire ffc_333_n;
  wire ffc_334_p;
  wire ffc_334_n;
  wire ffc_335_p;
  wire ffc_335_n;
  wire ffc_336_p;
  wire ffc_336_n;
  wire ffc_337_p;
  wire ffc_337_n;
  wire ffc_338_p;
  wire ffc_338_n;
  wire ffc_339_p;
  wire ffc_339_n;
  wire ffc_340_p;
  wire ffc_340_n;
  wire ffc_341_p;
  wire ffc_341_n;
  wire ffc_342_p;
  wire ffc_342_n;
  wire ffc_343_p;
  wire ffc_343_n;
  wire ffc_344_p;
  wire ffc_344_n;
  wire ffc_345_p;
  wire ffc_345_n;
  wire ffc_346_p;
  wire ffc_346_n;
  wire ffc_347_p;
  wire ffc_347_n;
  wire ffc_348_p;
  wire ffc_348_n;
  wire ffc_349_p;
  wire ffc_349_n;
  wire ffc_350_p;
  wire ffc_350_n;
  wire ffc_351_p;
  wire ffc_351_n;
  wire ffc_352_p;
  wire ffc_352_n;
  wire ffc_353_p;
  wire ffc_353_n;
  wire ffc_354_p;
  wire ffc_354_n;
  wire ffc_355_p;
  wire ffc_355_n;
  wire ffc_356_p;
  wire ffc_356_n;
  wire ffc_357_p;
  wire ffc_357_n;
  wire ffc_358_p;
  wire ffc_358_n;
  wire ffc_359_p;
  wire ffc_359_n;
  wire ffc_360_p;
  wire ffc_360_n;
  wire ffc_361_p;
  wire ffc_361_n;
  wire ffc_362_p;
  wire ffc_362_n;
  wire ffc_363_p;
  wire ffc_363_n;
  wire ffc_364_p;
  wire ffc_364_n;
  wire ffc_365_p;
  wire ffc_365_n;
  wire ffc_366_p;
  wire ffc_366_n;
  wire ffc_367_p;
  wire ffc_367_n;
  wire ffc_368_p;
  wire ffc_368_n;
  wire ffc_369_p;
  wire ffc_369_n;
  wire ffc_370_p;
  wire ffc_370_n;
  wire ffc_371_p;
  wire ffc_371_n;
  wire ffc_372_p;
  wire ffc_372_n;
  wire ffc_373_p;
  wire ffc_373_n;
  wire ffc_374_p;
  wire ffc_374_n;
  wire ffc_375_p;
  wire ffc_375_n;
  wire ffc_376_p;
  wire ffc_376_n;
  wire ffc_377_p;
  wire ffc_377_n;
  wire ffc_378_p;
  wire ffc_378_n;
  wire ffc_379_p;
  wire ffc_379_n;
  wire ffc_380_p;
  wire ffc_380_n;
  wire ffc_381_p;
  wire ffc_381_n;
  wire ffc_382_p;
  wire ffc_382_n;
  wire ffc_383_p;
  wire ffc_383_n;
  wire ffc_384_p;
  wire ffc_384_n;
  wire ffc_385_p;
  wire ffc_385_n;
  wire ffc_386_p;
  wire ffc_386_n;
  wire ffc_387_p;
  wire ffc_387_n;
  wire ffc_388_p;
  wire ffc_388_n;
  wire ffc_389_p;
  wire ffc_389_n;
  wire ffc_390_p;
  wire ffc_390_n;
  wire ffc_391_p;
  wire ffc_391_n;
  wire ffc_392_p;
  wire ffc_392_n;
  wire ffc_393_p;
  wire ffc_393_n;
  wire ffc_394_p;
  wire ffc_394_n;
  wire ffc_395_p;
  wire ffc_395_n;
  wire ffc_396_p;
  wire ffc_396_n;
  wire ffc_397_p;
  wire ffc_397_n;
  wire ffc_398_p;
  wire ffc_398_n;
  wire ffc_399_p;
  wire ffc_399_n;
  wire ffc_400_p;
  wire ffc_400_n;
  wire ffc_401_p;
  wire ffc_401_n;
  wire ffc_402_p;
  wire ffc_402_n;
  wire ffc_403_p;
  wire ffc_403_n;
  wire ffc_404_p;
  wire ffc_404_n;
  wire ffc_405_p;
  wire ffc_405_n;
  wire ffc_406_p;
  wire ffc_406_n;
  wire ffc_407_p;
  wire ffc_407_n;
  wire ffc_408_p;
  wire ffc_408_n;
  wire ffc_409_p;
  wire ffc_409_n;
  wire ffc_410_p;
  wire ffc_410_n;
  wire ffc_411_p;
  wire ffc_411_n;
  wire ffc_412_p;
  wire ffc_412_n;
  wire ffc_413_p;
  wire ffc_413_n;
  wire ffc_414_p;
  wire ffc_414_n;
  wire ffc_415_p;
  wire ffc_415_n;
  wire ffc_416_p;
  wire ffc_416_n;
  wire ffc_417_p;
  wire ffc_417_n;
  wire ffc_418_p;
  wire ffc_418_n;
  wire ffc_419_p;
  wire ffc_419_n;
  wire ffc_420_p;
  wire ffc_420_n;
  wire ffc_421_p;
  wire ffc_421_n;
  wire ffc_422_p;
  wire ffc_422_n;
  wire ffc_423_p;
  wire ffc_423_n;
  wire ffc_424_p;
  wire ffc_424_n;
  wire ffc_425_p;
  wire ffc_425_n;
  wire ffc_426_p;
  wire ffc_426_n;
  wire ffc_427_p;
  wire ffc_427_n;
  wire ffc_428_p;
  wire ffc_428_n;
  wire ffc_429_p;
  wire ffc_429_n;
  wire ffc_430_p;
  wire ffc_430_n;
  wire ffc_431_p;
  wire ffc_431_n;
  wire ffc_432_p;
  wire ffc_432_n;
  wire ffc_433_p;
  wire ffc_433_n;
  wire ffc_434_p;
  wire ffc_434_n;
  wire ffc_435_p;
  wire ffc_435_n;
  wire ffc_436_p;
  wire ffc_436_n;
  wire ffc_437_p;
  wire ffc_437_n;
  wire ffc_438_p;
  wire ffc_438_n;
  wire ffc_439_p;
  wire ffc_439_n;
  wire ffc_440_p;
  wire ffc_440_n;
  wire ffc_441_p;
  wire ffc_441_n;
  wire ffc_442_p;
  wire ffc_442_n;
  wire ffc_443_p;
  wire ffc_443_n;
  wire ffc_444_p;
  wire ffc_444_n;
  wire ffc_445_p;
  wire ffc_445_n;
  wire ffc_446_p;
  wire ffc_446_n;
  wire ffc_447_p;
  wire ffc_447_n;
  wire ffc_448_p;
  wire ffc_448_n;
  wire ffc_449_p;
  wire ffc_449_n;
  wire ffc_450_p;
  wire ffc_450_n;
  wire ffc_451_p;
  wire ffc_451_n;
  wire ffc_452_p;
  wire ffc_452_n;
  wire ffc_453_p;
  wire ffc_453_n;
  wire ffc_454_p;
  wire ffc_454_n;
  wire ffc_455_p;
  wire ffc_455_n;
  wire ffc_456_p;
  wire ffc_456_n;
  wire ffc_457_p;
  wire ffc_457_n;
  wire ffc_458_p;
  wire ffc_458_n;
  wire ffc_459_p;
  wire ffc_459_n;
  wire ffc_460_p;
  wire ffc_460_n;
  wire ffc_461_p;
  wire ffc_461_n;
  wire ffc_462_p;
  wire ffc_462_n;
  wire ffc_463_p;
  wire ffc_463_n;
  wire ffc_464_p;
  wire ffc_464_n;
  wire ffc_465_p;
  wire ffc_465_n;
  wire ffc_466_p;
  wire ffc_466_n;
  wire ffc_467_p;
  wire ffc_467_n;
  wire ffc_468_p;
  wire ffc_468_n;
  wire ffc_469_p;
  wire ffc_469_n;
  wire ffc_470_p;
  wire ffc_470_n;
  wire ffc_471_p;
  wire ffc_471_n;
  wire ffc_472_p;
  wire ffc_472_n;
  wire ffc_473_p;
  wire ffc_473_n;
  wire ffc_474_p;
  wire ffc_474_n;
  wire ffc_475_p;
  wire ffc_475_n;
  wire ffc_476_p;
  wire ffc_476_n;
  wire ffc_477_p;
  wire ffc_477_n;
  wire ffc_478_p;
  wire ffc_478_n;
  wire ffc_479_p;
  wire ffc_479_n;
  wire ffc_480_p;
  wire ffc_480_n;
  wire ffc_481_p;
  wire ffc_481_n;
  wire ffc_482_p;
  wire ffc_482_n;
  wire ffc_483_p;
  wire ffc_483_n;
  wire ffc_484_p;
  wire ffc_484_n;
  wire ffc_485_p;
  wire ffc_485_n;
  wire ffc_486_p;
  wire ffc_486_n;
  wire ffc_487_p;
  wire ffc_487_n;
  wire ffc_488_p;
  wire ffc_488_n;
  wire ffc_489_p;
  wire ffc_489_n;
  wire ffc_490_p;
  wire ffc_490_n;
  wire ffc_491_p;
  wire ffc_491_n;
  wire ffc_492_p;
  wire ffc_492_n;
  wire ffc_493_p;
  wire ffc_493_n;
  wire ffc_494_p;
  wire ffc_494_n;
  wire ffc_495_p;
  wire ffc_495_n;
  wire ffc_496_p;
  wire ffc_496_n;
  wire ffc_497_p;
  wire ffc_497_n;
  wire ffc_498_p;
  wire ffc_498_n;
  wire ffc_499_p;
  wire ffc_499_n;
  wire ffc_500_p;
  wire ffc_500_n;
  wire ffc_501_p;
  wire ffc_501_n;
  wire ffc_502_p;
  wire ffc_502_n;
  wire ffc_503_p;
  wire ffc_503_n;
  wire ffc_504_p;
  wire ffc_504_n;
  wire ffc_505_p;
  wire ffc_505_n;
  wire ffc_506_p;
  wire ffc_506_n;
  wire ffc_507_p;
  wire ffc_507_n;
  wire ffc_508_p;
  wire ffc_508_n;
  wire ffc_509_p;
  wire ffc_509_n;
  wire ffc_510_p;
  wire ffc_510_n;
  wire ffc_511_p;
  wire ffc_511_n;
  wire ffc_512_p;
  wire ffc_512_n;
  wire ffc_513_p;
  wire ffc_513_n;
  wire ffc_514_p;
  wire ffc_514_n;
  wire ffc_515_p;
  wire ffc_515_n;
  wire ffc_516_p;
  wire ffc_516_n;
  wire ffc_517_p;
  wire ffc_517_n;
  wire ffc_518_p;
  wire ffc_518_n;
  wire ffc_519_p;
  wire ffc_519_n;
  wire ffc_520_p;
  wire ffc_520_n;
  wire ffc_521_p;
  wire ffc_521_n;
  wire ffc_522_p;
  wire ffc_522_n;
  wire ffc_523_p;
  wire ffc_523_n;
  wire ffc_524_p;
  wire ffc_524_n;
  wire ffc_525_p;
  wire ffc_525_n;
  wire ffc_526_p;
  wire ffc_526_n;
  wire ffc_527_p;
  wire ffc_527_n;
  wire ffc_528_p;
  wire ffc_528_n;
  wire ffc_529_p;
  wire ffc_529_n;
  wire ffc_530_p;
  wire ffc_530_n;
  wire ffc_531_p;
  wire ffc_531_n;
  wire ffc_532_p;
  wire ffc_532_n;
  wire ffc_533_p;
  wire ffc_533_n;
  wire ffc_534_p;
  wire ffc_534_n;
  wire ffc_535_p;
  wire ffc_535_n;
  wire ffc_536_p;
  wire ffc_536_n;
  wire ffc_537_p;
  wire ffc_537_n;
  wire ffc_538_p;
  wire ffc_538_n;
  wire ffc_539_p;
  wire ffc_539_n;
  wire ffc_540_p;
  wire ffc_540_n;
  wire ffc_541_p;
  wire ffc_541_n;
  wire ffc_542_p;
  wire ffc_542_n;
  wire ffc_543_p;
  wire ffc_543_n;
  wire ffc_544_p;
  wire ffc_544_n;
  wire ffc_545_p;
  wire ffc_545_n;
  wire ffc_546_p;
  wire ffc_546_n;
  wire ffc_547_p;
  wire ffc_547_n;
  wire ffc_548_p;
  wire ffc_548_n;
  wire ffc_549_p;
  wire ffc_549_n;
  wire ffc_550_p;
  wire ffc_550_n;
  wire ffc_551_p;
  wire ffc_551_n;
  wire ffc_552_p;
  wire ffc_552_n;
  wire ffc_553_p;
  wire ffc_553_n;
  wire ffc_554_p;
  wire ffc_554_n;
  wire ffc_555_p;
  wire ffc_555_n;
  wire ffc_556_p;
  wire ffc_556_n;
  wire ffc_557_p;
  wire ffc_557_n;
  wire ffc_558_p;
  wire ffc_558_n;
  wire ffc_559_p;
  wire ffc_559_n;
  wire ffc_560_p;
  wire ffc_560_n;
  wire ffc_561_p;
  wire ffc_561_n;
  wire ffc_562_p;
  wire ffc_562_n;
  wire ffc_563_p;
  wire ffc_563_n;
  wire ffc_564_p;
  wire ffc_564_n;
  wire ffc_565_p;
  wire ffc_565_n;
  wire ffc_566_p;
  wire ffc_566_n;
  wire ffc_567_p;
  wire ffc_567_n;
  wire ffc_568_p;
  wire ffc_568_n;
  wire ffc_569_p;
  wire ffc_569_n;
  wire ffc_570_p;
  wire ffc_570_n;
  wire ffc_571_p;
  wire ffc_571_n;
  wire ffc_572_p;
  wire ffc_572_n;
  wire ffc_573_p;
  wire ffc_573_n;
  wire ffc_574_p;
  wire ffc_574_n;
  wire g733_p;
  wire g733_n;
  wire g734_p;
  wire g734_n;
  wire g735_p;
  wire g735_n;
  wire g736_p;
  wire g736_n;
  wire g737_p;
  wire g737_n;
  wire g738_p;
  wire g738_n;
  wire g739_p;
  wire g739_n;
  wire g740_p;
  wire g740_n;
  wire g741_p;
  wire g741_n;
  wire g742_p;
  wire g742_n;
  wire g743_p;
  wire g743_n;
  wire g744_p;
  wire g744_n;
  wire g745_p;
  wire g745_n;
  wire g746_p;
  wire g746_n;
  wire g747_p;
  wire g747_n;
  wire g748_p;
  wire g748_n;
  wire g749_p;
  wire g749_n;
  wire g750_p;
  wire g750_n;
  wire g751_p;
  wire g751_n;
  wire g752_p;
  wire g752_n;
  wire g753_p;
  wire g753_n;
  wire g754_p;
  wire g754_n;
  wire g755_p;
  wire g755_n;
  wire g756_p;
  wire g756_n;
  wire g757_p;
  wire g757_n;
  wire g758_p;
  wire g758_n;
  wire g759_p;
  wire g759_n;
  wire g760_p;
  wire g760_n;
  wire g761_p;
  wire g761_n;
  wire g762_p;
  wire g762_n;
  wire g763_p;
  wire g763_n;
  wire g764_p;
  wire g764_n;
  wire g765_p;
  wire g765_n;
  wire g766_p;
  wire g766_n;
  wire g767_p;
  wire g767_n;
  wire g768_p;
  wire g768_n;
  wire g769_p;
  wire g769_n;
  wire g770_p;
  wire g770_n;
  wire g771_p;
  wire g771_n;
  wire g772_p;
  wire g772_n;
  wire g773_p;
  wire g773_n;
  wire g774_p;
  wire g774_n;
  wire g775_p;
  wire g775_n;
  wire g776_p;
  wire g776_n;
  wire g777_p;
  wire g777_n;
  wire g778_p;
  wire g778_n;
  wire g779_p;
  wire g779_n;
  wire g780_p;
  wire g780_n;
  wire g781_p;
  wire g781_n;
  wire g782_p;
  wire g782_n;
  wire g783_p;
  wire g783_n;
  wire g784_p;
  wire g784_n;
  wire g785_p;
  wire g785_n;
  wire g786_p;
  wire g786_n;
  wire g787_p;
  wire g787_n;
  wire g788_p;
  wire g788_n;
  wire g789_p;
  wire g789_n;
  wire g790_p;
  wire g790_n;
  wire g791_p;
  wire g791_n;
  wire g792_p;
  wire g792_n;
  wire g793_p;
  wire g793_n;
  wire g794_p;
  wire g794_n;
  wire g795_p;
  wire g795_n;
  wire g796_p;
  wire g796_n;
  wire g797_p;
  wire g797_n;
  wire g798_p;
  wire g798_n;
  wire g799_p;
  wire g799_n;
  wire g800_p;
  wire g800_n;
  wire g801_p;
  wire g801_n;
  wire g802_p;
  wire g802_n;
  wire g803_p;
  wire g803_n;
  wire g804_p;
  wire g804_n;
  wire g805_p;
  wire g805_n;
  wire g806_p;
  wire g806_n;
  wire g807_p;
  wire g807_n;
  wire g808_p;
  wire g808_n;
  wire g809_p;
  wire g809_n;
  wire g810_p;
  wire g810_n;
  wire g811_p;
  wire g811_n;
  wire g812_p;
  wire g812_n;
  wire g813_p;
  wire g813_n;
  wire g814_p;
  wire g814_n;
  wire g815_p;
  wire g815_n;
  wire g816_p;
  wire g816_n;
  wire g817_p;
  wire g817_n;
  wire g818_p;
  wire g818_n;
  wire g819_p;
  wire g819_n;
  wire g820_p;
  wire g820_n;
  wire g821_p;
  wire g821_n;
  wire g822_p;
  wire g822_n;
  wire g823_p;
  wire g823_n;
  wire g824_p;
  wire g824_n;
  wire g825_p;
  wire g825_n;
  wire g826_p;
  wire g826_n;
  wire g827_p;
  wire g827_n;
  wire g828_p;
  wire g828_n;
  wire g829_p;
  wire g829_n;
  wire g830_p;
  wire g830_n;
  wire g831_p;
  wire g831_n;
  wire g832_p;
  wire g832_n;
  wire g833_p;
  wire g833_n;
  wire g834_p;
  wire g834_n;
  wire g835_p;
  wire g835_n;
  wire g836_p;
  wire g836_n;
  wire g837_p;
  wire g837_n;
  wire g838_p;
  wire g838_n;
  wire g839_p;
  wire g839_n;
  wire g840_p;
  wire g840_n;
  wire g841_p;
  wire g841_n;
  wire g842_p;
  wire g842_n;
  wire g843_p;
  wire g843_n;
  wire g844_p;
  wire g844_n;
  wire g845_p;
  wire g845_n;
  wire g846_p;
  wire g846_n;
  wire g847_p;
  wire g847_n;
  wire g848_p;
  wire g848_n;
  wire g849_p;
  wire g849_n;
  wire g850_p;
  wire g850_n;
  wire g851_p;
  wire g851_n;
  wire g852_p;
  wire g852_n;
  wire g853_p;
  wire g853_n;
  wire g854_p;
  wire g854_n;
  wire g855_p;
  wire g855_n;
  wire g856_p;
  wire g856_n;
  wire g857_p;
  wire g857_n;
  wire g858_p;
  wire g858_n;
  wire g859_p;
  wire g859_n;
  wire g860_p;
  wire g860_n;
  wire g861_p;
  wire g861_n;
  wire g862_p;
  wire g862_n;
  wire g863_p;
  wire g863_n;
  wire g864_p;
  wire g864_n;
  wire g865_p;
  wire g865_n;
  wire g866_p;
  wire g866_n;
  wire g867_p;
  wire g867_n;
  wire g868_p;
  wire g868_n;
  wire g869_p;
  wire g869_n;
  wire g870_p;
  wire g870_n;
  wire g871_p;
  wire g871_n;
  wire g872_p;
  wire g872_n;
  wire g873_p;
  wire g873_n;
  wire g874_p;
  wire g874_n;
  wire g875_p;
  wire g875_n;
  wire g876_p;
  wire g876_n;
  wire g877_p;
  wire g877_n;
  wire g878_p;
  wire g878_n;
  wire g879_p;
  wire g879_n;
  wire g880_p;
  wire g880_n;
  wire g881_p;
  wire g881_n;
  wire g882_p;
  wire g882_n;
  wire g883_p;
  wire g883_n;
  wire g884_p;
  wire g884_n;
  wire g885_p;
  wire g885_n;
  wire g886_p;
  wire g886_n;
  wire g887_p;
  wire g887_n;
  wire g888_p;
  wire g888_n;
  wire g889_p;
  wire g889_n;
  wire g890_p;
  wire g890_n;
  wire g891_p;
  wire g891_n;
  wire g892_p;
  wire g892_n;
  wire g893_p;
  wire g893_n;
  wire g894_p;
  wire g894_n;
  wire g895_p;
  wire g895_n;
  wire g896_p;
  wire g896_n;
  wire g897_p;
  wire g897_n;
  wire g898_p;
  wire g898_n;
  wire g899_p;
  wire g899_n;
  wire g900_p;
  wire g900_n;
  wire g901_p;
  wire g901_n;
  wire g902_p;
  wire g902_n;
  wire g903_p;
  wire g903_n;
  wire g904_p;
  wire g904_n;
  wire g905_p;
  wire g905_n;
  wire g906_p;
  wire g906_n;
  wire g907_p;
  wire g907_n;
  wire g908_p;
  wire g908_n;
  wire g909_p;
  wire g909_n;
  wire g910_p;
  wire g910_n;
  wire g911_p;
  wire g911_n;
  wire g912_p;
  wire g912_n;
  wire g913_p;
  wire g913_n;
  wire g914_p;
  wire g914_n;
  wire g915_p;
  wire g915_n;
  wire g916_p;
  wire g916_n;
  wire g917_p;
  wire g917_n;
  wire g918_p;
  wire g918_n;
  wire g919_p;
  wire g919_n;
  wire g920_p;
  wire g920_n;
  wire g921_p;
  wire g921_n;
  wire g922_p;
  wire g922_n;
  wire g923_p;
  wire g923_n;
  wire g924_p;
  wire g924_n;
  wire g925_p;
  wire g925_n;
  wire g926_p;
  wire g926_n;
  wire g927_p;
  wire g927_n;
  wire g928_p;
  wire g928_n;
  wire g929_p;
  wire g929_n;
  wire g930_p;
  wire g930_n;
  wire g931_p;
  wire g931_n;
  wire g932_p;
  wire g932_n;
  wire g933_p;
  wire g933_n;
  wire g934_p;
  wire g934_n;
  wire g935_p;
  wire g935_n;
  wire g936_p;
  wire g936_n;
  wire g937_p;
  wire g937_n;
  wire g938_p;
  wire g938_n;
  wire g939_p;
  wire g939_n;
  wire g940_p;
  wire g940_n;
  wire g941_p;
  wire g941_n;
  wire g942_p;
  wire g942_n;
  wire g943_p;
  wire g943_n;
  wire g944_p;
  wire g944_n;
  wire g945_p;
  wire g945_n;
  wire g946_p;
  wire g946_n;
  wire g947_p;
  wire g947_n;
  wire g948_p;
  wire g948_n;
  wire g949_p;
  wire g949_n;
  wire g950_p;
  wire g950_n;
  wire g951_p;
  wire g951_n;
  wire g952_p;
  wire g952_n;
  wire g953_p;
  wire g953_n;
  wire g954_p;
  wire g954_n;
  wire g955_p;
  wire g955_n;
  wire g956_p;
  wire g956_n;
  wire g957_p;
  wire g957_n;
  wire g958_p;
  wire g958_n;
  wire g959_p;
  wire g959_n;
  wire g960_p;
  wire g960_n;
  wire g961_p;
  wire g961_n;
  wire g962_p;
  wire g962_n;
  wire g963_p;
  wire g963_n;
  wire g964_p;
  wire g964_n;
  wire g965_p;
  wire g965_n;
  wire g966_p;
  wire g966_n;
  wire g967_p;
  wire g967_n;
  wire g968_p;
  wire g968_n;
  wire g969_p;
  wire g969_n;
  wire g970_p;
  wire g970_n;
  wire g971_p;
  wire g971_n;
  wire g972_p;
  wire g972_n;
  wire g973_p;
  wire g973_n;
  wire g974_p;
  wire g974_n;
  wire g975_p;
  wire g975_n;
  wire g976_p;
  wire g976_n;
  wire g977_p;
  wire g977_n;
  wire g978_p;
  wire g978_n;
  wire g979_p;
  wire g979_n;
  wire g980_p;
  wire g980_n;
  wire g981_p;
  wire g981_n;
  wire g982_p;
  wire g982_n;
  wire g983_p;
  wire g983_n;
  wire g984_p;
  wire g984_n;
  wire g985_p;
  wire g985_n;
  wire g986_p;
  wire g986_n;
  wire g987_p;
  wire g987_n;
  wire g988_p;
  wire g988_n;
  wire g989_p;
  wire g989_n;
  wire g990_p;
  wire g990_n;
  wire g991_p;
  wire g991_n;
  wire g992_p;
  wire g992_n;
  wire g993_p;
  wire g993_n;
  wire g994_p;
  wire g994_n;
  wire g995_p;
  wire g995_n;
  wire g996_p;
  wire g996_n;
  wire g997_p;
  wire g997_n;
  wire g998_p;
  wire g998_n;
  wire g999_p;
  wire g999_n;
  wire g1000_p;
  wire g1000_n;
  wire g1001_p;
  wire g1001_n;
  wire g1002_p;
  wire g1002_n;
  wire g1003_p;
  wire g1003_n;
  wire g1004_p;
  wire g1004_n;
  wire g1005_p;
  wire g1005_n;
  wire g1006_p;
  wire g1006_n;
  wire g1007_p;
  wire g1007_n;
  wire g1008_p;
  wire g1008_n;
  wire g1009_p;
  wire g1009_n;
  wire g1010_p;
  wire g1010_n;
  wire g1011_p;
  wire g1011_n;
  wire g1012_p;
  wire g1012_n;
  wire g1013_p;
  wire g1013_n;
  wire g1014_p;
  wire g1014_n;
  wire g1015_p;
  wire g1015_n;
  wire g1016_p;
  wire g1016_n;
  wire g1017_p;
  wire g1017_n;
  wire g1018_p;
  wire g1018_n;
  wire g1019_p;
  wire g1019_n;
  wire g1020_p;
  wire g1020_n;
  wire g1021_p;
  wire g1021_n;
  wire g1022_p;
  wire g1022_n;
  wire g1023_p;
  wire g1023_n;
  wire g1024_p;
  wire g1024_n;
  wire g1025_p;
  wire g1025_n;
  wire g1026_p;
  wire g1026_n;
  wire g1027_p;
  wire g1027_n;
  wire g1028_p;
  wire g1028_n;
  wire g1029_p;
  wire g1029_n;
  wire g1030_p;
  wire g1030_n;
  wire g1031_p;
  wire g1031_n;
  wire g1032_p;
  wire g1032_n;
  wire g1033_p;
  wire g1033_n;
  wire g1034_p;
  wire g1034_n;
  wire g1035_p;
  wire g1035_n;
  wire g1036_p;
  wire g1036_n;
  wire g1037_p;
  wire g1037_n;
  wire g1038_p;
  wire g1038_n;
  wire g1039_p;
  wire g1039_n;
  wire g1040_p;
  wire g1040_n;
  wire g1041_p;
  wire g1041_n;
  wire g1042_p;
  wire g1042_n;
  wire g1043_p;
  wire g1043_n;
  wire g1044_p;
  wire g1044_n;
  wire g1045_p;
  wire g1045_n;
  wire g1046_p;
  wire g1046_n;
  wire g1047_p;
  wire g1047_n;
  wire g1048_p;
  wire g1048_n;
  wire g1049_p;
  wire g1049_n;
  wire g1050_p;
  wire g1050_n;
  wire g1051_p;
  wire g1051_n;
  wire g1052_p;
  wire g1052_n;
  wire g1053_p;
  wire g1053_n;
  wire g1054_p;
  wire g1054_n;
  wire g1055_p;
  wire g1055_n;
  wire g1056_p;
  wire g1056_n;
  wire g1057_p;
  wire g1057_n;
  wire g1058_p;
  wire g1058_n;
  wire g1059_p;
  wire g1059_n;
  wire g1060_p;
  wire g1060_n;
  wire g1061_p;
  wire g1061_n;
  wire g1062_p;
  wire g1062_n;
  wire g1063_p;
  wire g1063_n;
  wire g1064_p;
  wire g1064_n;
  wire g1065_p;
  wire g1065_n;
  wire g1066_p;
  wire g1066_n;
  wire g1067_p;
  wire g1067_n;
  wire g1068_p;
  wire g1068_n;
  wire g1069_p;
  wire g1069_n;
  wire g1070_p;
  wire g1070_n;
  wire g1071_p;
  wire g1071_n;
  wire g1072_p;
  wire g1072_n;
  wire g1073_p;
  wire g1073_n;
  wire g1074_p;
  wire g1074_n;
  wire g1075_p;
  wire g1075_n;
  wire g1076_p;
  wire g1076_n;
  wire g1077_p;
  wire g1077_n;
  wire g1078_p;
  wire g1078_n;
  wire g1079_p;
  wire g1079_n;
  wire g1080_p;
  wire g1080_n;
  wire g1081_p;
  wire g1081_n;
  wire g1082_p;
  wire g1082_n;
  wire g1083_p;
  wire g1083_n;
  wire g1084_p;
  wire g1084_n;
  wire g1085_p;
  wire g1085_n;
  wire g1086_p;
  wire g1086_n;
  wire g1087_p;
  wire g1087_n;
  wire g1088_p;
  wire g1088_n;
  wire g1089_p;
  wire g1089_n;
  wire g1090_p;
  wire g1090_n;
  wire g1091_p;
  wire g1091_n;
  wire g1092_p;
  wire g1092_n;
  wire g1093_p;
  wire g1093_n;
  wire g1094_p;
  wire g1094_n;
  wire g1095_p;
  wire g1095_n;
  wire g1096_p;
  wire g1096_n;
  wire g1097_p;
  wire g1097_n;
  wire g1098_p;
  wire g1098_n;
  wire g1099_p;
  wire g1099_n;
  wire g1100_p;
  wire g1100_n;
  wire g1101_p;
  wire g1101_n;
  wire g1102_p;
  wire g1102_n;
  wire g1103_p;
  wire g1103_n;
  wire g1104_p;
  wire g1104_n;
  wire g1105_p;
  wire g1105_n;
  wire g1106_p;
  wire g1106_n;
  wire g1107_p;
  wire g1107_n;
  wire g1108_p;
  wire g1108_n;
  wire g1109_p;
  wire g1109_n;
  wire g1110_p;
  wire g1110_n;
  wire g1111_p;
  wire g1111_n;
  wire g1112_p;
  wire g1112_n;
  wire g1113_p;
  wire g1113_n;
  wire g1114_p;
  wire g1114_n;
  wire g1115_p;
  wire g1115_n;
  wire g1116_p;
  wire g1116_n;
  wire g1117_p;
  wire g1117_n;
  wire g1118_p;
  wire g1118_n;
  wire g1119_p;
  wire g1119_n;
  wire g1120_p;
  wire g1120_n;
  wire g1121_p;
  wire g1121_n;
  wire g1122_p;
  wire g1122_n;
  wire g1123_p;
  wire g1123_n;
  wire g1124_p;
  wire g1124_n;
  wire g1125_p;
  wire g1125_n;
  wire g1126_p;
  wire g1126_n;
  wire g1127_p;
  wire g1127_n;
  wire g1128_p;
  wire g1128_n;
  wire g1129_p;
  wire g1129_n;
  wire g1130_p;
  wire g1130_n;
  wire g1131_p;
  wire g1131_n;
  wire g1132_p;
  wire g1132_n;
  wire g1133_p;
  wire g1133_n;
  wire g1134_p;
  wire g1134_n;
  wire g1135_p;
  wire g1135_n;
  wire g1136_p;
  wire g1136_n;
  wire g1137_p;
  wire g1137_n;
  wire g1138_p;
  wire g1138_n;
  wire g1139_p;
  wire g1139_n;
  wire g1140_p;
  wire g1140_n;
  wire g1141_p;
  wire g1141_n;
  wire g1142_p;
  wire g1142_n;
  wire g1143_p;
  wire g1143_n;
  wire g1144_p;
  wire g1144_n;
  wire g1145_p;
  wire g1145_n;
  wire g1146_p;
  wire g1146_n;
  wire g1147_p;
  wire g1147_n;
  wire g1148_p;
  wire g1148_n;
  wire g1149_p;
  wire g1149_n;
  wire g1150_p;
  wire g1150_n;
  wire g1151_p;
  wire g1151_n;
  wire g1152_p;
  wire g1152_n;
  wire g1153_p;
  wire g1153_n;
  wire g1154_p;
  wire g1154_n;
  wire g1155_p;
  wire g1155_n;
  wire g1156_p;
  wire g1156_n;
  wire g1157_p;
  wire g1157_n;
  wire g1158_p;
  wire g1158_n;
  wire g1159_p;
  wire g1159_n;
  wire g1160_p;
  wire g1160_n;
  wire g1161_p;
  wire g1161_n;
  wire g1162_p;
  wire g1162_n;
  wire g1163_p;
  wire g1163_n;
  wire g1164_p;
  wire g1164_n;
  wire g1165_p;
  wire g1165_n;
  wire g1166_p;
  wire g1166_n;
  wire g1167_p;
  wire g1167_n;
  wire g1168_p;
  wire g1168_n;
  wire g1169_p;
  wire g1169_n;
  wire g1170_p;
  wire g1170_n;
  wire g1171_p;
  wire g1171_n;
  wire g1172_p;
  wire g1172_n;
  wire g1173_p;
  wire g1173_n;
  wire g1174_p;
  wire g1174_n;
  wire g1175_p;
  wire g1175_n;
  wire g1176_p;
  wire g1176_n;
  wire g1177_p;
  wire g1177_n;
  wire g1178_p;
  wire g1178_n;
  wire g1179_p;
  wire g1179_n;
  wire g1180_p;
  wire g1180_n;
  wire g1181_p;
  wire g1181_n;
  wire g1182_p;
  wire g1182_n;
  wire g1183_p;
  wire g1183_n;
  wire g1184_p;
  wire g1184_n;
  wire g1185_p;
  wire g1185_n;
  wire g1186_p;
  wire g1186_n;
  wire g1187_p;
  wire g1187_n;
  wire g1188_p;
  wire g1188_n;
  wire g1189_p;
  wire g1189_n;
  wire g1190_p;
  wire g1190_n;
  wire g1191_p;
  wire g1191_n;
  wire g1192_p;
  wire g1192_n;
  wire g1193_p;
  wire g1193_n;
  wire g1194_p;
  wire g1194_n;
  wire g1195_p;
  wire g1195_n;
  wire g1196_p;
  wire g1196_n;
  wire g1197_p;
  wire g1197_n;
  wire g1198_p;
  wire g1198_n;
  wire g1199_p;
  wire g1199_n;
  wire g1200_p;
  wire g1200_n;
  wire g1201_p;
  wire g1201_n;
  wire g1202_p;
  wire g1202_n;
  wire g1203_p;
  wire g1203_n;
  wire g1204_p;
  wire g1204_n;
  wire g1205_p;
  wire g1205_n;
  wire g1206_p;
  wire g1206_n;
  wire g1207_p;
  wire g1207_n;
  wire g1208_p;
  wire g1208_n;
  wire g1209_p;
  wire g1209_n;
  wire g1210_p;
  wire g1210_n;
  wire g1211_p;
  wire g1211_n;
  wire g1212_p;
  wire g1212_n;
  wire g1213_p;
  wire g1213_n;
  wire g1214_p;
  wire g1214_n;
  wire g1215_p;
  wire g1215_n;
  wire g1216_p;
  wire g1216_n;
  wire g1217_p;
  wire g1217_n;
  wire g1218_p;
  wire g1218_n;
  wire g1219_p;
  wire g1219_n;
  wire g1220_p;
  wire g1220_n;
  wire g1221_p;
  wire g1221_n;
  wire g1222_p;
  wire g1222_n;
  wire g1223_p;
  wire g1223_n;
  wire g1224_p;
  wire g1224_n;
  wire g1225_p;
  wire g1225_n;
  wire g1226_p;
  wire g1226_n;
  wire g1227_p;
  wire g1227_n;
  wire g1228_p;
  wire g1228_n;
  wire g1229_p;
  wire g1229_n;
  wire g1230_p;
  wire g1230_n;
  wire g1231_p;
  wire g1231_n;
  wire g1232_p;
  wire g1232_n;
  wire g1233_p;
  wire g1233_n;
  wire g1234_p;
  wire g1234_n;
  wire g1235_p;
  wire g1235_n;
  wire g1236_p;
  wire g1236_n;
  wire g1237_p;
  wire g1237_n;
  wire g1238_p;
  wire g1238_n;
  wire g1239_p;
  wire g1239_n;
  wire g1240_p;
  wire g1240_n;
  wire g1241_p;
  wire g1241_n;
  wire g1242_p;
  wire g1242_n;
  wire g1243_p;
  wire g1243_n;
  wire g1244_p;
  wire g1244_n;
  wire g1245_p;
  wire g1245_n;
  wire g1246_p;
  wire g1246_n;
  wire g1247_p;
  wire g1247_n;
  wire g1248_p;
  wire g1248_n;
  wire g1249_p;
  wire g1249_n;
  wire g1250_p;
  wire g1250_n;
  wire g1251_p;
  wire g1251_n;
  wire g1252_p;
  wire g1252_n;
  wire g1253_p;
  wire g1253_n;
  wire g1254_p;
  wire g1254_n;
  wire g1255_p;
  wire g1255_n;
  wire g1256_p;
  wire g1256_n;
  wire g1257_p;
  wire g1257_n;
  wire g1258_p;
  wire g1258_n;
  wire g1259_p;
  wire g1259_n;
  wire g1260_p;
  wire g1260_n;
  wire g1261_p;
  wire g1261_n;
  wire g1262_p;
  wire g1262_n;
  wire g1263_p;
  wire g1263_n;
  wire g1264_p;
  wire g1264_n;
  wire g1265_p;
  wire g1265_n;
  wire g1266_p;
  wire g1266_n;
  wire g1267_p;
  wire g1267_n;
  wire g1268_p;
  wire g1268_n;
  wire g1269_p;
  wire g1269_n;
  wire g1270_p;
  wire g1270_n;
  wire g1271_p;
  wire g1271_n;
  wire g1272_p;
  wire g1272_n;
  wire g1273_p;
  wire g1273_n;
  wire g1274_p;
  wire g1274_n;
  wire g1275_p;
  wire g1275_n;
  wire g1276_p;
  wire g1276_n;
  wire g1277_p;
  wire g1277_n;
  wire g1278_p;
  wire g1278_n;
  wire g1279_p;
  wire g1279_n;
  wire g1280_p;
  wire g1280_n;
  wire g1281_p;
  wire g1281_n;
  wire g1282_p;
  wire g1282_n;
  wire g1283_p;
  wire g1283_n;
  wire g1284_p;
  wire g1284_n;
  wire g1285_p;
  wire g1285_n;
  wire g1286_p;
  wire g1286_n;
  wire g1287_p;
  wire g1287_n;
  wire g1288_p;
  wire g1288_n;
  wire g1289_p;
  wire g1289_n;
  wire g1290_p;
  wire g1290_n;
  wire g1291_p;
  wire g1291_n;
  wire g1292_p;
  wire g1292_n;
  wire g1293_p;
  wire g1293_n;
  wire g1294_p;
  wire g1294_n;
  wire g1295_p;
  wire g1295_n;
  wire g1296_p;
  wire g1296_n;
  wire g1297_p;
  wire g1297_n;
  wire g1298_p;
  wire g1298_n;
  wire g1299_p;
  wire g1299_n;
  wire g1300_p;
  wire g1300_n;
  wire g1301_p;
  wire g1301_n;
  wire g1302_p;
  wire g1302_n;
  wire ffc_279_n_spl_;
  wire ffc_261_n_spl_;
  wire ffc_261_n_spl_0;
  wire ffc_261_n_spl_1;
  wire g737_n_spl_;
  wire g737_n_spl_0;
  wire g740_n_spl_;
  wire g741_n_spl_;
  wire ffc_283_n_spl_;
  wire ffc_283_n_spl_0;
  wire g745_n_spl_;
  wire g745_n_spl_0;
  wire g752_n_spl_;
  wire ffc_287_p_spl_;
  wire ffc_287_p_spl_0;
  wire ffc_287_p_spl_1;
  wire ffc_391_n_spl_;
  wire ffc_287_n_spl_;
  wire ffc_287_n_spl_0;
  wire ffc_287_n_spl_1;
  wire ffc_392_p_spl_;
  wire g749_n_spl_;
  wire ffc_270_p_spl_;
  wire ffc_391_p_spl_;
  wire ffc_452_n_spl_;
  wire ffc_452_n_spl_0;
  wire ffc_483_p_spl_;
  wire ffc_485_n_spl_;
  wire ffc_483_n_spl_;
  wire ffc_485_p_spl_;
  wire ffc_482_n_spl_;
  wire ffc_497_p_spl_;
  wire ffc_482_p_spl_;
  wire ffc_497_n_spl_;
  wire ffc_398_p_spl_;
  wire ffc_94_n_spl_;
  wire ffc_438_n_spl_;
  wire ffc_452_p_spl_;
  wire ffc_438_p_spl_;
  wire g851_p_spl_;
  wire g851_n_spl_;
  wire g868_n_spl_;
  wire ffc_491_p_spl_;
  wire g875_n_spl_;
  wire g877_n_spl_;
  wire g876_n_spl_;
  wire g774_p_spl_;
  wire g779_p_spl_;
  wire g788_p_spl_;
  wire g849_p_spl_;
  wire g864_p_spl_;
  wire ffc_415_p_spl_;
  wire ffc_415_p_spl_0;
  wire ffc_415_p_spl_1;
  wire ffc_415_n_spl_;
  wire ffc_415_n_spl_0;
  wire ffc_415_n_spl_1;
  wire ffc_404_p_spl_;
  wire ffc_404_p_spl_0;
  wire ffc_404_p_spl_00;
  wire ffc_404_p_spl_01;
  wire ffc_404_p_spl_1;
  wire ffc_404_p_spl_10;
  wire ffc_404_p_spl_11;
  wire ffc_404_n_spl_;
  wire ffc_404_n_spl_0;
  wire ffc_404_n_spl_00;
  wire ffc_404_n_spl_01;
  wire ffc_404_n_spl_1;
  wire ffc_404_n_spl_10;
  wire ffc_404_n_spl_11;
  wire ffc_442_p_spl_;
  wire ffc_442_p_spl_0;
  wire ffc_443_p_spl_;
  wire ffc_443_p_spl_0;
  wire ffc_442_n_spl_;
  wire ffc_442_n_spl_0;
  wire ffc_443_n_spl_;
  wire ffc_443_n_spl_0;
  wire g896_p_spl_;
  wire g899_p_spl_;
  wire ffc_406_n_spl_;
  wire ffc_406_n_spl_0;
  wire ffc_406_n_spl_00;
  wire ffc_406_n_spl_01;
  wire ffc_406_n_spl_1;
  wire ffc_406_p_spl_;
  wire ffc_406_p_spl_0;
  wire ffc_406_p_spl_00;
  wire ffc_406_p_spl_01;
  wire ffc_406_p_spl_1;
  wire g901_p_spl_;
  wire g906_p_spl_;
  wire ffc_405_n_spl_;
  wire ffc_405_p_spl_;
  wire ffc_439_n_spl_;
  wire g900_n_spl_;
  wire g900_n_spl_0;
  wire ffc_439_p_spl_;
  wire ffc_439_p_spl_0;
  wire ffc_439_p_spl_1;
  wire g900_p_spl_;
  wire ffc_342_n_spl_;
  wire ffc_342_n_spl_0;
  wire ffc_346_n_spl_;
  wire ffc_399_n_spl_;
  wire ffc_399_n_spl_0;
  wire ffc_399_n_spl_1;
  wire ffc_399_p_spl_;
  wire ffc_399_p_spl_0;
  wire ffc_399_p_spl_1;
  wire ffc_564_p_spl_;
  wire ffc_565_p_spl_;
  wire g939_p_spl_;
  wire g940_p_spl_;
  wire ffc_505_n_spl_;
  wire g908_n_spl_;
  wire g908_n_spl_0;
  wire g908_n_spl_1;
  wire ffc_318_p_spl_;
  wire ffc_318_p_spl_0;
  wire g943_n_spl_;
  wire g943_n_spl_0;
  wire g943_n_spl_00;
  wire g943_n_spl_1;
  wire g925_p_spl_;
  wire g943_p_spl_;
  wire g943_p_spl_0;
  wire g943_p_spl_00;
  wire g943_p_spl_1;
  wire ffc_41_p_spl_;
  wire ffc_41_p_spl_0;
  wire ffc_41_p_spl_00;
  wire ffc_41_p_spl_000;
  wire ffc_41_p_spl_01;
  wire ffc_41_p_spl_1;
  wire ffc_41_p_spl_10;
  wire ffc_41_p_spl_11;
  wire ffc_41_n_spl_;
  wire ffc_41_n_spl_0;
  wire ffc_41_n_spl_00;
  wire ffc_41_n_spl_000;
  wire ffc_41_n_spl_01;
  wire ffc_41_n_spl_1;
  wire ffc_41_n_spl_10;
  wire ffc_41_n_spl_11;
  wire ffc_445_p_spl_;
  wire ffc_445_p_spl_0;
  wire ffc_445_p_spl_00;
  wire ffc_445_p_spl_1;
  wire g925_n_spl_;
  wire g925_n_spl_0;
  wire g913_p_spl_;
  wire g913_p_spl_0;
  wire ffc_74_p_spl_;
  wire ffc_74_p_spl_0;
  wire ffc_74_p_spl_00;
  wire ffc_74_p_spl_01;
  wire ffc_74_p_spl_1;
  wire ffc_74_p_spl_10;
  wire ffc_74_p_spl_11;
  wire ffc_74_n_spl_;
  wire ffc_74_n_spl_0;
  wire ffc_74_n_spl_00;
  wire ffc_74_n_spl_01;
  wire ffc_74_n_spl_1;
  wire ffc_74_n_spl_10;
  wire ffc_74_n_spl_11;
  wire ffc_417_p_spl_;
  wire ffc_417_p_spl_0;
  wire ffc_417_p_spl_1;
  wire ffc_540_p_spl_;
  wire ffc_540_p_spl_0;
  wire ffc_416_p_spl_;
  wire ffc_416_p_spl_0;
  wire ffc_505_p_spl_;
  wire ffc_308_n_spl_;
  wire ffc_308_n_spl_0;
  wire ffc_308_n_spl_00;
  wire ffc_308_n_spl_1;
  wire g964_p_spl_;
  wire g964_p_spl_0;
  wire g964_p_spl_1;
  wire g966_p_spl_;
  wire g966_p_spl_0;
  wire g966_p_spl_1;
  wire g971_n_spl_;
  wire g971_n_spl_0;
  wire g971_n_spl_1;
  wire g971_p_spl_;
  wire g971_p_spl_0;
  wire ffc_428_n_spl_;
  wire ffc_428_p_spl_;
  wire ffc_428_p_spl_0;
  wire ffc_544_p_spl_;
  wire ffc_544_p_spl_0;
  wire ffc_544_p_spl_00;
  wire ffc_544_p_spl_01;
  wire ffc_544_p_spl_1;
  wire ffc_445_n_spl_;
  wire ffc_544_n_spl_;
  wire g928_n_spl_;
  wire ffc_533_p_spl_;
  wire ffc_533_p_spl_0;
  wire ffc_533_p_spl_00;
  wire ffc_533_p_spl_000;
  wire ffc_533_p_spl_001;
  wire ffc_533_p_spl_01;
  wire ffc_533_p_spl_010;
  wire ffc_533_p_spl_1;
  wire ffc_533_p_spl_10;
  wire ffc_533_p_spl_11;
  wire ffc_563_p_spl_;
  wire ffc_563_p_spl_0;
  wire ffc_563_p_spl_00;
  wire ffc_563_p_spl_1;
  wire ffc_533_n_spl_;
  wire ffc_533_n_spl_0;
  wire ffc_533_n_spl_00;
  wire ffc_533_n_spl_1;
  wire ffc_532_p_spl_;
  wire ffc_532_p_spl_0;
  wire ffc_532_p_spl_00;
  wire ffc_532_p_spl_000;
  wire ffc_532_p_spl_001;
  wire ffc_532_p_spl_01;
  wire ffc_532_p_spl_1;
  wire ffc_532_p_spl_10;
  wire ffc_532_p_spl_11;
  wire ffc_532_n_spl_;
  wire ffc_532_n_spl_0;
  wire ffc_532_n_spl_00;
  wire ffc_532_n_spl_000;
  wire ffc_532_n_spl_001;
  wire ffc_532_n_spl_01;
  wire ffc_532_n_spl_010;
  wire ffc_532_n_spl_011;
  wire ffc_532_n_spl_1;
  wire ffc_532_n_spl_10;
  wire ffc_532_n_spl_100;
  wire ffc_532_n_spl_101;
  wire ffc_532_n_spl_11;
  wire ffc_532_n_spl_110;
  wire g938_n_spl_;
  wire g938_n_spl_0;
  wire ffc_99_p_spl_;
  wire ffc_163_p_spl_;
  wire ffc_120_p_spl_;
  wire ffc_141_p_spl_;
  wire ffc_190_p_spl_;
  wire ffc_244_p_spl_;
  wire ffc_208_p_spl_;
  wire ffc_226_p_spl_;
  wire ffc_269_p_spl_;
  wire ffc_422_n_spl_;
  wire ffc_422_n_spl_0;
  wire ffc_422_n_spl_1;
  wire g1005_n_spl_;
  wire ffc_423_n_spl_;
  wire ffc_423_n_spl_0;
  wire g948_n_spl_;
  wire ffc_440_n_spl_;
  wire ffc_440_n_spl_0;
  wire ffc_440_n_spl_1;
  wire g1011_n_spl_;
  wire g903_n_spl_;
  wire g903_n_spl_0;
  wire g903_n_spl_1;
  wire ffc_305_n_spl_;
  wire ffc_305_n_spl_0;
  wire ffc_305_n_spl_1;
  wire g1016_n_spl_;
  wire g1021_n_spl_;
  wire ffc_311_n_spl_;
  wire ffc_311_n_spl_0;
  wire ffc_311_n_spl_1;
  wire g954_n_spl_;
  wire g919_n_spl_;
  wire g919_n_spl_0;
  wire ffc_315_n_spl_;
  wire ffc_315_n_spl_0;
  wire ffc_315_n_spl_1;
  wire g1028_n_spl_;
  wire ffc_318_n_spl_;
  wire g951_n_spl_;
  wire g960_n_spl_;
  wire g957_n_spl_;
  wire g963_n_spl_;
  wire ffc_350_p_spl_;
  wire ffc_354_p_spl_;
  wire g919_p_spl_;
  wire g913_n_spl_;
  wire ffc_546_p_spl_;
  wire ffc_546_p_spl_0;
  wire ffc_546_p_spl_1;
  wire g942_n_spl_;
  wire g968_n_spl_;
  wire ffc_541_p_spl_;
  wire ffc_541_p_spl_0;
  wire g1051_n_spl_;
  wire g1051_n_spl_0;
  wire g1051_n_spl_1;
  wire g897_p_spl_;
  wire g898_p_spl_;
  wire g1055_n_spl_;
  wire g1055_n_spl_0;
  wire ffc_441_p_spl_;
  wire g944_n_spl_;
  wire g945_p_spl_;
  wire ffc_322_p_spl_;
  wire ffc_322_n_spl_;
  wire ffc_541_n_spl_;
  wire ffc_541_n_spl_0;
  wire g1071_n_spl_;
  wire g1072_p_spl_;
  wire ffc_424_n_spl_;
  wire ffc_424_n_spl_0;
  wire g1075_n_spl_;
  wire g1076_p_spl_;
  wire g1079_n_spl_;
  wire g1082_n_spl_;
  wire ffc_548_n_spl_;
  wire ffc_547_n_spl_;
  wire g974_n_spl_;
  wire ffc_342_p_spl_;
  wire ffc_346_p_spl_;
  wire g929_n_spl_;
  wire g902_p_spl_;
  wire ffc_386_n_spl_;
  wire ffc_386_p_spl_;
  wire ffc_424_p_spl_;
  wire ffc_424_p_spl_0;
  wire g1099_p_spl_;
  wire g1107_p_spl_;
  wire g907_n_spl_;
  wire g980_n_spl_;
  wire g980_n_spl_0;
  wire g1112_n_spl_;
  wire ffc_377_p_spl_;
  wire ffc_380_n_spl_;
  wire ffc_377_n_spl_;
  wire ffc_380_p_spl_;
  wire ffc_422_p_spl_;
  wire ffc_423_p_spl_;
  wire ffc_423_p_spl_0;
  wire ffc_308_p_spl_;
  wire ffc_311_p_spl_;
  wire ffc_311_p_spl_0;
  wire ffc_383_n_spl_;
  wire ffc_383_p_spl_;
  wire ffc_440_p_spl_;
  wire ffc_416_n_spl_;
  wire g1055_p_spl_;
  wire ffc_516_p_spl_;
  wire ffc_517_n_spl_;
  wire ffc_516_n_spl_;
  wire ffc_517_p_spl_;
  wire ffc_514_p_spl_;
  wire ffc_515_n_spl_;
  wire ffc_514_n_spl_;
  wire ffc_515_p_spl_;
  wire g1141_p_spl_;
  wire g1144_p_spl_;
  wire g1141_n_spl_;
  wire g1144_n_spl_;
  wire ffc_367_p_spl_;
  wire ffc_370_n_spl_;
  wire ffc_367_n_spl_;
  wire ffc_370_p_spl_;
  wire g1156_n_spl_;
  wire g1159_p_spl_;
  wire ffc_542_p_spl_;
  wire ffc_542_n_spl_;
  wire ffc_417_n_spl_;
  wire ffc_540_n_spl_;
  wire g1164_p_spl_;
  wire g1167_p_spl_;
  wire g1164_n_spl_;
  wire g1167_n_spl_;
  wire g1051_p_spl_;
  wire ffc_332_p_spl_;
  wire g941_n_spl_;
  wire g941_n_spl_0;
  wire g941_n_spl_1;
  wire ffc_295_p_spl_;
  wire g941_p_spl_;
  wire g941_p_spl_0;
  wire g941_p_spl_00;
  wire g941_p_spl_1;
  wire g995_n_spl_;
  wire g995_n_spl_0;
  wire g1204_p_spl_;
  wire ffc_444_n_spl_;
  wire ffc_444_n_spl_0;
  wire ffc_444_n_spl_00;
  wire ffc_444_n_spl_000;
  wire ffc_444_n_spl_001;
  wire ffc_444_n_spl_01;
  wire ffc_444_n_spl_010;
  wire ffc_444_n_spl_011;
  wire ffc_444_n_spl_1;
  wire ffc_444_n_spl_10;
  wire ffc_444_n_spl_11;
  wire ffc_444_p_spl_;
  wire ffc_444_p_spl_0;
  wire ffc_444_p_spl_00;
  wire ffc_444_p_spl_000;
  wire ffc_444_p_spl_001;
  wire ffc_444_p_spl_01;
  wire ffc_444_p_spl_010;
  wire ffc_444_p_spl_011;
  wire ffc_444_p_spl_1;
  wire ffc_444_p_spl_10;
  wire ffc_444_p_spl_100;
  wire ffc_444_p_spl_11;
  wire ffc_504_p_spl_;
  wire ffc_504_p_spl_0;
  wire ffc_504_p_spl_1;
  wire ffc_504_n_spl_;
  wire ffc_504_n_spl_0;
  wire g1040_n_spl_;
  wire g1183_n_spl_;
  wire ffc_335_p_spl_;
  wire ffc_299_p_spl_;
  wire ffc_338_p_spl_;
  wire ffc_301_p_spl_;
  wire ffc_325_p_spl_;
  wire ffc_293_p_spl_;
  wire g986_n_spl_;
  wire ffc_574_p_spl_;
  wire ffc_574_p_spl_0;
  wire ffc_574_p_spl_00;
  wire ffc_574_p_spl_1;
  wire ffc_574_n_spl_;
  wire ffc_574_n_spl_0;
  wire ffc_574_n_spl_1;
  wire ffc_356_n_spl_;
  wire ffc_356_p_spl_;
  wire ffc_356_p_spl_0;
  wire ffc_266_n_spl_;
  wire ffc_266_p_spl_;
  wire ffc_266_p_spl_0;
  wire g1284_n_spl_;
  wire g1288_n_spl_;
  wire ffc_291_n_spl_;
  wire ffc_330_n_spl_;
  wire ffc_330_n_spl_0;
  wire g742_n_spl_;
  wire g758_p_spl_;
  wire g761_n_spl_;
  wire g766_p_spl_;
  wire g838_n_spl_;
  wire g859_p_spl_;
  wire g895_n_spl_;

  orX
  g_g733_n
  (
    .dout(g733_n),
    .din1(ffc_401_n),
    .din2(ffc_418_n)
  );


  orX
  g_g734_n
  (
    .dout(g734_n),
    .din1(ffc_7_n),
    .din2(ffc_38_n)
  );


  orX
  g_g735_n
  (
    .dout(g735_n),
    .din1(ffc_279_n_spl_),
    .din2(g734_n)
  );


  andX
  g_g736_p
  (
    .dout(g736_p),
    .din1(ffc_185_p),
    .din2(ffc_261_n_spl_0)
  );


  orX
  g_g737_n
  (
    .dout(g737_n),
    .din1(ffc_24_n),
    .din2(ffc_279_n_spl_)
  );


  orX
  g_g738_n
  (
    .dout(g738_n),
    .din1(ffc_274_n),
    .din2(g737_n_spl_0)
  );


  orX
  g_g739_n
  (
    .dout(g739_n),
    .din1(ffc_360_n),
    .din2(g737_n_spl_0)
  );


  orX
  g_g740_n
  (
    .dout(g740_n),
    .din1(ffc_449_n),
    .din2(ffc_451_n)
  );


  orX
  g_g741_n
  (
    .dout(g741_n),
    .din1(ffc_448_n),
    .din2(ffc_450_n)
  );


  orX
  g_g742_n
  (
    .dout(g742_n),
    .din1(g740_n_spl_),
    .din2(g741_n_spl_)
  );


  andX
  g_g743_p
  (
    .dout(g743_p),
    .din1(ffc_360_p),
    .din2(g741_n_spl_)
  );


  andX
  g_g744_p
  (
    .dout(g744_p),
    .din1(ffc_274_p),
    .din2(g740_n_spl_)
  );


  orX
  g_g745_n
  (
    .dout(g745_n),
    .din1(g743_p),
    .din2(g744_p)
  );


  andX
  g_g746_p
  (
    .dout(g746_p),
    .din1(ffc_387_n),
    .din2(ffc_388_n)
  );


  andX
  g_g747_p
  (
    .dout(g747_p),
    .din1(ffc_395_n),
    .din2(ffc_396_n)
  );


  andX
  g_g748_p
  (
    .dout(g748_p),
    .din1(ffc_400_n),
    .din2(ffc_403_n)
  );


  orX
  g_g749_n
  (
    .dout(g749_n),
    .din1(ffc_394_p),
    .din2(ffc_397_p)
  );


  orX
  g_g750_n
  (
    .dout(g750_n),
    .din1(ffc_283_n_spl_0),
    .din2(ffc_390_p)
  );


  orX
  g_g751_n
  (
    .dout(g751_n),
    .din1(ffc_265_n),
    .din2(ffc_279_p)
  );


  orX
  g_g752_n
  (
    .dout(g752_n),
    .din1(g745_n_spl_0),
    .din2(g751_n)
  );


  orX
  g_g753_n
  (
    .dout(g753_n),
    .din1(ffc_90_n),
    .din2(g752_n_spl_)
  );


  andX
  g_g754_p
  (
    .dout(g754_p),
    .din1(ffc_3_p),
    .din2(ffc_11_p)
  );


  orX
  g_g755_n
  (
    .dout(g755_n),
    .din1(g752_n_spl_),
    .din2(g754_p)
  );


  orX
  g_g756_n
  (
    .dout(g756_n),
    .din1(ffc_287_p_spl_0),
    .din2(ffc_391_n_spl_)
  );


  orX
  g_g757_n
  (
    .dout(g757_n),
    .din1(ffc_287_n_spl_0),
    .din2(ffc_392_p_spl_)
  );


  andX
  g_g758_p
  (
    .dout(g758_p),
    .din1(g756_n),
    .din2(g757_n)
  );


  andX
  g_g759_p
  (
    .dout(g759_p),
    .din1(ffc_287_n_spl_0),
    .din2(ffc_393_n)
  );


  andX
  g_g760_p
  (
    .dout(g760_p),
    .din1(ffc_287_p_spl_0),
    .din2(g749_n_spl_)
  );


  orX
  g_g761_n
  (
    .dout(g761_n),
    .din1(g759_p),
    .din2(g760_p)
  );


  andX
  g_g762_p
  (
    .dout(g762_p),
    .din1(ffc_270_p_spl_),
    .din2(ffc_283_n_spl_0)
  );


  orX
  g_g763_n
  (
    .dout(g763_n),
    .din1(ffc_391_p_spl_),
    .din2(g762_p)
  );


  orX
  g_g764_n
  (
    .dout(g764_n),
    .din1(ffc_287_p_spl_1),
    .din2(ffc_390_n)
  );


  orX
  g_g765_n
  (
    .dout(g765_n),
    .din1(ffc_287_n_spl_1),
    .din2(ffc_452_n_spl_0)
  );


  andX
  g_g766_p
  (
    .dout(g766_p),
    .din1(g764_n),
    .din2(g765_n)
  );


  orX
  g_g767_n
  (
    .dout(g767_n),
    .din1(ffc_351_p),
    .din2(ffc_419_n)
  );


  orX
  g_g768_n
  (
    .dout(g768_n),
    .din1(ffc_351_n),
    .din2(ffc_419_p)
  );


  andX
  g_g769_p
  (
    .dout(g769_p),
    .din1(g767_n),
    .din2(g768_n)
  );


  orX
  g_g770_n
  (
    .dout(g770_n),
    .din1(ffc_355_p),
    .din2(g769_p)
  );


  orX
  g_g771_n
  (
    .dout(g771_n),
    .din1(ffc_496_n),
    .din2(ffc_499_n)
  );


  orX
  g_g772_n
  (
    .dout(g772_n),
    .din1(ffc_496_p),
    .din2(ffc_499_p)
  );


  andX
  g_g773_p
  (
    .dout(g773_p),
    .din1(ffc_34_p),
    .din2(g772_n)
  );


  andX
  g_g774_p
  (
    .dout(g774_p),
    .din1(g771_n),
    .din2(g773_p)
  );


  andX
  g_g775_p
  (
    .dout(g775_p),
    .din1(ffc_492_n),
    .din2(ffc_493_n)
  );


  orX
  g_g775_n
  (
    .dout(g775_n),
    .din1(ffc_492_p),
    .din2(ffc_493_p)
  );


  andX
  g_g776_p
  (
    .dout(g776_p),
    .din1(ffc_471_n),
    .din2(ffc_472_n)
  );


  orX
  g_g776_n
  (
    .dout(g776_n),
    .din1(ffc_471_p),
    .din2(ffc_472_p)
  );


  orX
  g_g777_n
  (
    .dout(g777_n),
    .din1(g775_n),
    .din2(g776_p)
  );


  orX
  g_g778_n
  (
    .dout(g778_n),
    .din1(g775_p),
    .din2(g776_n)
  );


  andX
  g_g779_p
  (
    .dout(g779_p),
    .din1(g777_n),
    .din2(g778_n)
  );


  andX
  g_g780_p
  (
    .dout(g780_p),
    .din1(ffc_483_p_spl_),
    .din2(ffc_485_n_spl_)
  );


  orX
  g_g780_n
  (
    .dout(g780_n),
    .din1(ffc_483_n_spl_),
    .din2(ffc_485_p_spl_)
  );


  andX
  g_g781_p
  (
    .dout(g781_p),
    .din1(ffc_483_n_spl_),
    .din2(ffc_485_p_spl_)
  );


  orX
  g_g781_n
  (
    .dout(g781_n),
    .din1(ffc_483_p_spl_),
    .din2(ffc_485_n_spl_)
  );


  andX
  g_g782_p
  (
    .dout(g782_p),
    .din1(g780_n),
    .din2(g781_n)
  );


  orX
  g_g782_n
  (
    .dout(g782_n),
    .din1(g780_p),
    .din2(g781_p)
  );


  andX
  g_g783_p
  (
    .dout(g783_p),
    .din1(ffc_482_n_spl_),
    .din2(ffc_497_p_spl_)
  );


  orX
  g_g783_n
  (
    .dout(g783_n),
    .din1(ffc_482_p_spl_),
    .din2(ffc_497_n_spl_)
  );


  andX
  g_g784_p
  (
    .dout(g784_p),
    .din1(ffc_482_p_spl_),
    .din2(ffc_497_n_spl_)
  );


  orX
  g_g784_n
  (
    .dout(g784_n),
    .din1(ffc_482_n_spl_),
    .din2(ffc_497_p_spl_)
  );


  andX
  g_g785_p
  (
    .dout(g785_p),
    .din1(g783_n),
    .din2(g784_n)
  );


  orX
  g_g785_n
  (
    .dout(g785_n),
    .din1(g783_p),
    .din2(g784_p)
  );


  orX
  g_g786_n
  (
    .dout(g786_n),
    .din1(g782_p),
    .din2(g785_n)
  );


  orX
  g_g787_n
  (
    .dout(g787_n),
    .din1(g782_n),
    .din2(g785_p)
  );


  andX
  g_g788_p
  (
    .dout(g788_p),
    .din1(g786_n),
    .din2(g787_n)
  );


  andX
  g_g789_p
  (
    .dout(g789_p),
    .din1(ffc_347_n),
    .din2(ffc_480_p)
  );


  andX
  g_g790_p
  (
    .dout(g790_p),
    .din1(ffc_336_p),
    .din2(ffc_434_n)
  );


  andX
  g_g791_p
  (
    .dout(g791_p),
    .din1(ffc_302_n),
    .din2(ffc_476_p)
  );


  orX
  g_g792_n
  (
    .dout(g792_n),
    .din1(g790_p),
    .din2(g791_p)
  );


  orX
  g_g793_n
  (
    .dout(g793_n),
    .din1(g789_p),
    .din2(g792_n)
  );


  andX
  g_g794_p
  (
    .dout(g794_p),
    .din1(ffc_323_p),
    .din2(ffc_478_n)
  );


  andX
  g_g795_p
  (
    .dout(g795_p),
    .din1(ffc_339_n),
    .din2(ffc_433_p)
  );


  orX
  g_g796_n
  (
    .dout(g796_n),
    .din1(g794_p),
    .din2(g795_p)
  );


  andX
  g_g797_p
  (
    .dout(g797_p),
    .din1(ffc_343_p),
    .din2(ffc_435_n)
  );


  andX
  g_g798_p
  (
    .dout(g798_p),
    .din1(ffc_323_n),
    .din2(ffc_478_p)
  );


  orX
  g_g799_n
  (
    .dout(g799_n),
    .din1(g797_p),
    .din2(g798_p)
  );


  orX
  g_g800_n
  (
    .dout(g800_n),
    .din1(g796_n),
    .din2(g799_n)
  );


  andX
  g_g801_p
  (
    .dout(g801_p),
    .din1(ffc_296_n),
    .din2(ffc_430_p)
  );


  andX
  g_g802_p
  (
    .dout(g802_p),
    .din1(ffc_302_p),
    .din2(ffc_476_n)
  );


  orX
  g_g803_n
  (
    .dout(g803_n),
    .din1(g801_p),
    .din2(g802_p)
  );


  andX
  g_g804_p
  (
    .dout(g804_p),
    .din1(ffc_319_n),
    .din2(ffc_431_p)
  );


  andX
  g_g805_p
  (
    .dout(g805_p),
    .din1(ffc_347_p),
    .din2(ffc_480_n)
  );


  orX
  g_g806_n
  (
    .dout(g806_n),
    .din1(g804_p),
    .din2(g805_p)
  );


  orX
  g_g807_n
  (
    .dout(g807_n),
    .din1(g803_n),
    .din2(g806_n)
  );


  orX
  g_g808_n
  (
    .dout(g808_n),
    .din1(g800_n),
    .din2(g807_n)
  );


  orX
  g_g809_n
  (
    .dout(g809_n),
    .din1(g793_n),
    .din2(g808_n)
  );


  andX
  g_g810_p
  (
    .dout(g810_p),
    .din1(ffc_312_p),
    .din2(ffc_432_n)
  );


  andX
  g_g811_p
  (
    .dout(g811_p),
    .din1(ffc_446_n),
    .din2(ffc_447_n)
  );


  orX
  g_g812_n
  (
    .dout(g812_n),
    .din1(ffc_30_n),
    .din2(g811_p)
  );


  orX
  g_g813_n
  (
    .dout(g813_n),
    .din1(g810_p),
    .din2(g812_n)
  );


  andX
  g_g814_p
  (
    .dout(g814_p),
    .din1(ffc_333_n),
    .din2(ffc_479_p)
  );


  andX
  g_g815_p
  (
    .dout(g815_p),
    .din1(ffc_333_p),
    .din2(ffc_479_n)
  );


  orX
  g_g816_n
  (
    .dout(g816_n),
    .din1(g814_p),
    .din2(g815_p)
  );


  andX
  g_g817_p
  (
    .dout(g817_p),
    .din1(ffc_326_p),
    .din2(ffc_481_n)
  );


  andX
  g_g818_p
  (
    .dout(g818_p),
    .din1(ffc_326_n),
    .din2(ffc_481_p)
  );


  orX
  g_g819_n
  (
    .dout(g819_n),
    .din1(g817_p),
    .din2(g818_p)
  );


  orX
  g_g820_n
  (
    .dout(g820_n),
    .din1(g816_n),
    .din2(g819_n)
  );


  orX
  g_g821_n
  (
    .dout(g821_n),
    .din1(g813_n),
    .din2(g820_n)
  );


  orX
  g_g822_n
  (
    .dout(g822_n),
    .din1(ffc_462_p),
    .din2(ffc_464_p)
  );


  orX
  g_g823_n
  (
    .dout(g823_n),
    .din1(ffc_453_p),
    .din2(ffc_465_p)
  );


  orX
  g_g824_n
  (
    .dout(g824_n),
    .din1(g822_n),
    .din2(g823_n)
  );


  orX
  g_g825_n
  (
    .dout(g825_n),
    .din1(ffc_454_p),
    .din2(ffc_468_p)
  );


  orX
  g_g826_n
  (
    .dout(g826_n),
    .din1(ffc_456_p),
    .din2(ffc_469_p)
  );


  orX
  g_g827_n
  (
    .dout(g827_n),
    .din1(g825_n),
    .din2(g826_n)
  );


  orX
  g_g828_n
  (
    .dout(g828_n),
    .din1(g824_n),
    .din2(g827_n)
  );


  orX
  g_g829_n
  (
    .dout(g829_n),
    .din1(ffc_457_p),
    .din2(ffc_458_p)
  );


  orX
  g_g830_n
  (
    .dout(g830_n),
    .din1(ffc_455_p),
    .din2(ffc_470_p)
  );


  orX
  g_g831_n
  (
    .dout(g831_n),
    .din1(g829_n),
    .din2(g830_n)
  );


  orX
  g_g832_n
  (
    .dout(g832_n),
    .din1(ffc_460_p),
    .din2(ffc_461_p)
  );


  orX
  g_g833_n
  (
    .dout(g833_n),
    .din1(ffc_459_p),
    .din2(ffc_467_p)
  );


  orX
  g_g834_n
  (
    .dout(g834_n),
    .din1(g832_n),
    .din2(g833_n)
  );


  orX
  g_g835_n
  (
    .dout(g835_n),
    .din1(g831_n),
    .din2(g834_n)
  );


  orX
  g_g836_n
  (
    .dout(g836_n),
    .din1(g828_n),
    .din2(g835_n)
  );


  orX
  g_g837_n
  (
    .dout(g837_n),
    .din1(g821_n),
    .din2(g836_n)
  );


  orX
  g_g838_n
  (
    .dout(g838_n),
    .din1(g809_n),
    .din2(g837_n)
  );


  andX
  g_g839_p
  (
    .dout(g839_p),
    .din1(ffc_270_p_spl_),
    .din2(ffc_391_n_spl_)
  );


  orX
  g_g839_n
  (
    .dout(g839_n),
    .din1(ffc_270_n),
    .din2(ffc_391_p_spl_)
  );


  andX
  g_g840_p
  (
    .dout(g840_p),
    .din1(ffc_412_n),
    .din2(g839_p)
  );


  andX
  g_g841_p
  (
    .dout(g841_p),
    .din1(ffc_412_p),
    .din2(g839_n)
  );


  orX
  g_g842_n
  (
    .dout(g842_n),
    .din1(g840_p),
    .din2(g841_p)
  );


  andX
  g_g843_p
  (
    .dout(g843_p),
    .din1(ffc_283_n_spl_),
    .din2(g842_n)
  );


  andX
  g_g844_p
  (
    .dout(g844_p),
    .din1(ffc_283_p),
    .din2(ffc_398_p_spl_)
  );


  orX
  g_g845_n
  (
    .dout(g845_n),
    .din1(g843_p),
    .din2(g844_p)
  );


  orX
  g_g846_n
  (
    .dout(g846_n),
    .din1(ffc_498_p),
    .din2(ffc_502_p)
  );


  orX
  g_g847_n
  (
    .dout(g847_n),
    .din1(ffc_498_n),
    .din2(ffc_502_n)
  );


  andX
  g_g848_p
  (
    .dout(g848_p),
    .din1(ffc_94_n_spl_),
    .din2(g847_n)
  );


  andX
  g_g849_p
  (
    .dout(g849_p),
    .din1(g846_n),
    .din2(g848_p)
  );


  orX
  g_g850_n
  (
    .dout(g850_n),
    .din1(ffc_287_p_spl_1),
    .din2(ffc_398_p_spl_)
  );


  andX
  g_g851_p
  (
    .dout(g851_p),
    .din1(ffc_500_n),
    .din2(ffc_501_n)
  );


  orX
  g_g851_n
  (
    .dout(g851_n),
    .din1(ffc_500_p),
    .din2(ffc_501_p)
  );


  andX
  g_g852_p
  (
    .dout(g852_p),
    .din1(ffc_438_n_spl_),
    .din2(ffc_452_p_spl_)
  );


  orX
  g_g852_n
  (
    .dout(g852_n),
    .din1(ffc_438_p_spl_),
    .din2(ffc_452_n_spl_0)
  );


  andX
  g_g853_p
  (
    .dout(g853_p),
    .din1(ffc_438_p_spl_),
    .din2(ffc_452_n_spl_)
  );


  orX
  g_g853_n
  (
    .dout(g853_n),
    .din1(ffc_438_n_spl_),
    .din2(ffc_452_p_spl_)
  );


  andX
  g_g854_p
  (
    .dout(g854_p),
    .din1(g852_n),
    .din2(g853_n)
  );


  orX
  g_g854_n
  (
    .dout(g854_n),
    .din1(g852_p),
    .din2(g853_p)
  );


  orX
  g_g855_n
  (
    .dout(g855_n),
    .din1(g851_p_spl_),
    .din2(g854_p)
  );


  orX
  g_g856_n
  (
    .dout(g856_n),
    .din1(g851_n_spl_),
    .din2(g854_n)
  );


  andX
  g_g857_p
  (
    .dout(g857_p),
    .din1(g855_n),
    .din2(g856_n)
  );


  orX
  g_g858_n
  (
    .dout(g858_n),
    .din1(ffc_287_n_spl_1),
    .din2(g857_p)
  );


  andX
  g_g859_p
  (
    .dout(g859_p),
    .din1(g850_n),
    .din2(g858_n)
  );


  andX
  g_g860_p
  (
    .dout(g860_p),
    .din1(ffc_494_p),
    .din2(ffc_495_n)
  );


  orX
  g_g860_n
  (
    .dout(g860_n),
    .din1(ffc_494_n),
    .din2(ffc_495_p)
  );


  orX
  g_g861_n
  (
    .dout(g861_n),
    .din1(g851_p_spl_),
    .din2(g860_n)
  );


  orX
  g_g862_n
  (
    .dout(g862_n),
    .din1(g851_n_spl_),
    .din2(g860_p)
  );


  andX
  g_g863_p
  (
    .dout(g863_p),
    .din1(ffc_94_n_spl_),
    .din2(g862_n)
  );


  andX
  g_g864_p
  (
    .dout(g864_p),
    .din1(g861_n),
    .din2(g863_p)
  );


  orX
  g_g865_n
  (
    .dout(g865_n),
    .din1(ffc_426_p),
    .din2(ffc_436_n)
  );


  orX
  g_g866_n
  (
    .dout(g866_n),
    .din1(ffc_477_p),
    .din2(ffc_490_p)
  );


  andX
  g_g867_p
  (
    .dout(g867_p),
    .din1(g865_n),
    .din2(g866_n)
  );


  orX
  g_g868_n
  (
    .dout(g868_n),
    .din1(ffc_466_p),
    .din2(ffc_473_p)
  );


  orX
  g_g869_n
  (
    .dout(g869_n),
    .din1(ffc_463_p),
    .din2(ffc_474_p)
  );


  orX
  g_g870_n
  (
    .dout(g870_n),
    .din1(g868_n_spl_),
    .din2(g869_n)
  );


  orX
  g_g871_n
  (
    .dout(g871_n),
    .din1(g867_p),
    .din2(g870_n)
  );


  orX
  g_g872_n
  (
    .dout(g872_n),
    .din1(ffc_463_n),
    .din2(g868_n_spl_)
  );


  andX
  g_g873_p
  (
    .dout(g873_p),
    .din1(ffc_466_n),
    .din2(g872_n)
  );


  andX
  g_g874_p
  (
    .dout(g874_p),
    .din1(g871_n),
    .din2(g873_p)
  );


  orX
  g_g875_n
  (
    .dout(g875_n),
    .din1(ffc_488_p),
    .din2(ffc_489_p)
  );


  orX
  g_g876_n
  (
    .dout(g876_n),
    .din1(ffc_491_p_spl_),
    .din2(g875_n_spl_)
  );


  orX
  g_g877_n
  (
    .dout(g877_n),
    .din1(ffc_486_p),
    .din2(ffc_487_p)
  );


  andX
  g_g878_p
  (
    .dout(g878_p),
    .din1(ffc_427_n),
    .din2(ffc_429_p)
  );


  orX
  g_g879_n
  (
    .dout(g879_n),
    .din1(ffc_484_p),
    .din2(g878_p)
  );


  orX
  g_g880_n
  (
    .dout(g880_n),
    .din1(g877_n_spl_),
    .din2(g879_n)
  );


  orX
  g_g881_n
  (
    .dout(g881_n),
    .din1(g876_n_spl_),
    .din2(g880_n)
  );


  orX
  g_g882_n
  (
    .dout(g882_n),
    .din1(g874_p),
    .din2(g881_n)
  );


  orX
  g_g883_n
  (
    .dout(g883_n),
    .din1(ffc_484_n),
    .din2(ffc_491_p_spl_)
  );


  orX
  g_g884_n
  (
    .dout(g884_n),
    .din1(g877_n_spl_),
    .din2(g883_n)
  );


  andX
  g_g885_p
  (
    .dout(g885_p),
    .din1(ffc_437_n),
    .din2(g884_n)
  );


  orX
  g_g886_n
  (
    .dout(g886_n),
    .din1(g875_n_spl_),
    .din2(g885_p)
  );


  orX
  g_g887_n
  (
    .dout(g887_n),
    .din1(ffc_486_n),
    .din2(g876_n_spl_)
  );


  andX
  g_g888_p
  (
    .dout(g888_p),
    .din1(ffc_488_n),
    .din2(g887_n)
  );


  andX
  g_g889_p
  (
    .dout(g889_p),
    .din1(g886_n),
    .din2(g888_p)
  );


  andX
  g_g890_p
  (
    .dout(g890_p),
    .din1(g882_n),
    .din2(g889_p)
  );


  orX
  g_g891_n
  (
    .dout(g891_n),
    .din1(g774_p_spl_),
    .din2(g779_p_spl_)
  );


  orX
  g_g892_n
  (
    .dout(g892_n),
    .din1(g788_p_spl_),
    .din2(g891_n)
  );


  orX
  g_g893_n
  (
    .dout(g893_n),
    .din1(g745_n_spl_0),
    .din2(g849_p_spl_)
  );


  orX
  g_g894_n
  (
    .dout(g894_n),
    .din1(g864_p_spl_),
    .din2(g893_n)
  );


  orX
  g_g895_n
  (
    .dout(g895_n),
    .din1(g892_n),
    .din2(g894_n)
  );


  andX
  g_g896_p
  (
    .dout(g896_p),
    .din1(ffc_415_p_spl_0),
    .din2(ffc_508_p)
  );


  orX
  g_g896_n
  (
    .dout(g896_n),
    .din1(ffc_415_n_spl_0),
    .din2(ffc_508_n)
  );


  andX
  g_g897_p
  (
    .dout(g897_p),
    .din1(ffc_404_p_spl_00),
    .din2(ffc_534_p)
  );


  orX
  g_g897_n
  (
    .dout(g897_n),
    .din1(ffc_404_n_spl_00),
    .din2(ffc_534_n)
  );


  andX
  g_g898_p
  (
    .dout(g898_p),
    .din1(ffc_404_n_spl_00),
    .din2(ffc_537_p)
  );


  orX
  g_g898_n
  (
    .dout(g898_n),
    .din1(ffc_404_p_spl_00),
    .din2(ffc_537_n)
  );


  andX
  g_g899_p
  (
    .dout(g899_p),
    .din1(ffc_529_p),
    .din2(ffc_543_n)
  );


  orX
  g_g899_n
  (
    .dout(g899_n),
    .din1(ffc_529_n),
    .din2(ffc_543_p)
  );


  andX
  g_g900_p
  (
    .dout(g900_p),
    .din1(ffc_530_n),
    .din2(ffc_545_n)
  );


  orX
  g_g900_n
  (
    .dout(g900_n),
    .din1(ffc_530_p),
    .din2(ffc_545_p)
  );


  andX
  g_g901_p
  (
    .dout(g901_p),
    .din1(ffc_128_p),
    .din2(ffc_415_p_spl_0)
  );


  orX
  g_g901_n
  (
    .dout(g901_n),
    .din1(ffc_128_n),
    .din2(ffc_415_n_spl_0)
  );


  andX
  g_g902_p
  (
    .dout(g902_p),
    .din1(ffc_442_p_spl_0),
    .din2(ffc_443_p_spl_0)
  );


  orX
  g_g902_n
  (
    .dout(g902_n),
    .din1(ffc_442_n_spl_0),
    .din2(ffc_443_n_spl_0)
  );


  andX
  g_g903_p
  (
    .dout(g903_p),
    .din1(g896_n),
    .din2(g899_n)
  );


  orX
  g_g903_n
  (
    .dout(g903_n),
    .din1(g896_p_spl_),
    .din2(g899_p_spl_)
  );


  andX
  g_g904_p
  (
    .dout(g904_p),
    .din1(ffc_406_n_spl_00),
    .din2(ffc_522_n)
  );


  orX
  g_g904_n
  (
    .dout(g904_n),
    .din1(ffc_406_p_spl_00),
    .din2(ffc_522_p)
  );


  andX
  g_g905_p
  (
    .dout(g905_p),
    .din1(ffc_525_n),
    .din2(ffc_528_n)
  );


  orX
  g_g905_n
  (
    .dout(g905_n),
    .din1(ffc_525_p),
    .din2(ffc_528_p)
  );


  andX
  g_g906_p
  (
    .dout(g906_p),
    .din1(g904_n),
    .din2(g905_p)
  );


  orX
  g_g906_n
  (
    .dout(g906_n),
    .din1(g904_p),
    .din2(g905_n)
  );


  andX
  g_g907_p
  (
    .dout(g907_p),
    .din1(ffc_475_n),
    .din2(ffc_503_n)
  );


  orX
  g_g907_n
  (
    .dout(g907_n),
    .din1(ffc_475_p),
    .din2(ffc_503_p)
  );


  andX
  g_g908_p
  (
    .dout(g908_p),
    .din1(g901_n),
    .din2(g906_n)
  );


  orX
  g_g908_n
  (
    .dout(g908_n),
    .din1(g901_p_spl_),
    .din2(g906_p_spl_)
  );


  andX
  g_g909_p
  (
    .dout(g909_p),
    .din1(ffc_526_n),
    .din2(ffc_527_p)
  );


  orX
  g_g909_n
  (
    .dout(g909_n),
    .din1(ffc_526_p),
    .din2(ffc_527_n)
  );


  andX
  g_g910_p
  (
    .dout(g910_p),
    .din1(ffc_405_n_spl_),
    .din2(g909_n)
  );


  orX
  g_g910_n
  (
    .dout(g910_n),
    .din1(ffc_405_p_spl_),
    .din2(g909_p)
  );


  andX
  g_g911_p
  (
    .dout(g911_p),
    .din1(ffc_406_p_spl_00),
    .din2(ffc_509_n)
  );


  orX
  g_g911_n
  (
    .dout(g911_n),
    .din1(ffc_406_n_spl_00),
    .din2(ffc_509_p)
  );


  andX
  g_g912_p
  (
    .dout(g912_p),
    .din1(ffc_405_p_spl_),
    .din2(g911_p)
  );


  orX
  g_g912_n
  (
    .dout(g912_n),
    .din1(ffc_405_n_spl_),
    .din2(g911_n)
  );


  andX
  g_g913_p
  (
    .dout(g913_p),
    .din1(g910_n),
    .din2(g912_n)
  );


  orX
  g_g913_n
  (
    .dout(g913_n),
    .din1(g910_p),
    .din2(g912_p)
  );


  andX
  g_g914_p
  (
    .dout(g914_p),
    .din1(ffc_519_n),
    .din2(ffc_524_n)
  );


  orX
  g_g914_n
  (
    .dout(g914_n),
    .din1(ffc_519_p),
    .din2(ffc_524_p)
  );


  andX
  g_g915_p
  (
    .dout(g915_p),
    .din1(ffc_406_p_spl_01),
    .din2(g914_n)
  );


  orX
  g_g915_n
  (
    .dout(g915_n),
    .din1(ffc_406_n_spl_01),
    .din2(g914_p)
  );


  andX
  g_g916_p
  (
    .dout(g916_p),
    .din1(ffc_415_p_spl_1),
    .din2(ffc_507_p)
  );


  orX
  g_g916_n
  (
    .dout(g916_n),
    .din1(ffc_415_n_spl_1),
    .din2(ffc_507_n)
  );


  andX
  g_g917_p
  (
    .dout(g917_p),
    .din1(ffc_406_n_spl_01),
    .din2(ffc_521_p)
  );


  orX
  g_g917_n
  (
    .dout(g917_n),
    .din1(ffc_406_p_spl_01),
    .din2(ffc_521_n)
  );


  andX
  g_g918_p
  (
    .dout(g918_p),
    .din1(g916_n),
    .din2(g917_n)
  );


  orX
  g_g918_n
  (
    .dout(g918_n),
    .din1(g916_p),
    .din2(g917_p)
  );


  andX
  g_g919_p
  (
    .dout(g919_p),
    .din1(g915_n),
    .din2(g918_p)
  );


  orX
  g_g919_n
  (
    .dout(g919_n),
    .din1(g915_p),
    .din2(g918_n)
  );


  andX
  g_g920_p
  (
    .dout(g920_p),
    .din1(ffc_518_n),
    .din2(ffc_523_n)
  );


  orX
  g_g920_n
  (
    .dout(g920_n),
    .din1(ffc_518_p),
    .din2(ffc_523_p)
  );


  andX
  g_g921_p
  (
    .dout(g921_p),
    .din1(ffc_406_p_spl_1),
    .din2(g920_n)
  );


  orX
  g_g921_n
  (
    .dout(g921_n),
    .din1(ffc_406_n_spl_1),
    .din2(g920_p)
  );


  andX
  g_g922_p
  (
    .dout(g922_p),
    .din1(ffc_415_p_spl_1),
    .din2(ffc_506_p)
  );


  orX
  g_g922_n
  (
    .dout(g922_n),
    .din1(ffc_415_n_spl_1),
    .din2(ffc_506_n)
  );


  andX
  g_g923_p
  (
    .dout(g923_p),
    .din1(ffc_406_n_spl_1),
    .din2(ffc_520_p)
  );


  orX
  g_g923_n
  (
    .dout(g923_n),
    .din1(ffc_406_p_spl_1),
    .din2(ffc_520_n)
  );


  andX
  g_g924_p
  (
    .dout(g924_p),
    .din1(g922_n),
    .din2(g923_n)
  );


  orX
  g_g924_n
  (
    .dout(g924_n),
    .din1(g922_p),
    .din2(g923_p)
  );


  andX
  g_g925_p
  (
    .dout(g925_p),
    .din1(g921_n),
    .din2(g924_p)
  );


  orX
  g_g925_n
  (
    .dout(g925_n),
    .din1(g921_p),
    .din2(g924_n)
  );


  andX
  g_g926_p
  (
    .dout(g926_p),
    .din1(ffc_439_n_spl_),
    .din2(g900_n_spl_0)
  );


  orX
  g_g926_n
  (
    .dout(g926_n),
    .din1(ffc_439_p_spl_0),
    .din2(g900_p_spl_)
  );


  andX
  g_g927_p
  (
    .dout(g927_p),
    .din1(ffc_439_p_spl_0),
    .din2(g900_p_spl_)
  );


  orX
  g_g927_n
  (
    .dout(g927_n),
    .din1(ffc_439_n_spl_),
    .din2(g900_n_spl_0)
  );


  andX
  g_g928_p
  (
    .dout(g928_p),
    .din1(g926_n),
    .din2(g927_n)
  );


  orX
  g_g928_n
  (
    .dout(g928_n),
    .din1(g926_p),
    .din2(g927_p)
  );


  orX
  g_g929_n
  (
    .dout(g929_n),
    .din1(ffc_342_n_spl_0),
    .din2(ffc_346_n_spl_)
  );


  andX
  g_g930_p
  (
    .dout(g930_p),
    .din1(ffc_399_n_spl_0),
    .din2(ffc_510_p)
  );


  orX
  g_g930_n
  (
    .dout(g930_n),
    .din1(ffc_399_p_spl_0),
    .din2(ffc_510_n)
  );


  andX
  g_g931_p
  (
    .dout(g931_p),
    .din1(ffc_399_p_spl_0),
    .din2(ffc_513_p)
  );


  orX
  g_g931_n
  (
    .dout(g931_n),
    .din1(ffc_399_n_spl_0),
    .din2(ffc_513_n)
  );


  andX
  g_g932_p
  (
    .dout(g932_p),
    .din1(g930_n),
    .din2(g931_n)
  );


  orX
  g_g932_n
  (
    .dout(g932_n),
    .din1(g930_p),
    .din2(g931_p)
  );


  andX
  g_g933_p
  (
    .dout(g933_p),
    .din1(ffc_404_p_spl_01),
    .din2(g932_n)
  );


  orX
  g_g933_n
  (
    .dout(g933_n),
    .din1(ffc_404_n_spl_01),
    .din2(g932_p)
  );


  andX
  g_g934_p
  (
    .dout(g934_p),
    .din1(ffc_399_n_spl_1),
    .din2(ffc_511_p)
  );


  orX
  g_g934_n
  (
    .dout(g934_n),
    .din1(ffc_399_p_spl_1),
    .din2(ffc_511_n)
  );


  andX
  g_g935_p
  (
    .dout(g935_p),
    .din1(ffc_399_p_spl_1),
    .din2(ffc_512_p)
  );


  orX
  g_g935_n
  (
    .dout(g935_n),
    .din1(ffc_399_n_spl_1),
    .din2(ffc_512_n)
  );


  andX
  g_g936_p
  (
    .dout(g936_p),
    .din1(g934_n),
    .din2(g935_n)
  );


  orX
  g_g936_n
  (
    .dout(g936_n),
    .din1(g934_p),
    .din2(g935_p)
  );


  andX
  g_g937_p
  (
    .dout(g937_p),
    .din1(ffc_404_n_spl_01),
    .din2(g936_n)
  );


  orX
  g_g937_n
  (
    .dout(g937_n),
    .din1(ffc_404_p_spl_01),
    .din2(g936_p)
  );


  andX
  g_g938_p
  (
    .dout(g938_p),
    .din1(g933_n),
    .din2(g937_n)
  );


  orX
  g_g938_n
  (
    .dout(g938_n),
    .din1(g933_p),
    .din2(g937_p)
  );


  andX
  g_g939_p
  (
    .dout(g939_p),
    .din1(ffc_554_p),
    .din2(ffc_564_n)
  );


  orX
  g_g939_n
  (
    .dout(g939_n),
    .din1(ffc_554_n),
    .din2(ffc_564_p_spl_)
  );


  andX
  g_g940_p
  (
    .dout(g940_p),
    .din1(ffc_559_n),
    .din2(ffc_565_p_spl_)
  );


  orX
  g_g940_n
  (
    .dout(g940_n),
    .din1(ffc_559_p),
    .din2(ffc_565_n)
  );


  andX
  g_g941_p
  (
    .dout(g941_p),
    .din1(g939_p_spl_),
    .din2(g940_p_spl_)
  );


  orX
  g_g941_n
  (
    .dout(g941_n),
    .din1(g939_n),
    .din2(g940_n)
  );


  orX
  g_g942_n
  (
    .dout(g942_n),
    .din1(ffc_505_n_spl_),
    .din2(g908_n_spl_0)
  );


  andX
  g_g943_p
  (
    .dout(g943_p),
    .din1(ffc_420_p),
    .din2(ffc_421_n)
  );


  orX
  g_g943_n
  (
    .dout(g943_n),
    .din1(ffc_420_n),
    .din2(ffc_421_p)
  );


  orX
  g_g944_n
  (
    .dout(g944_n),
    .din1(ffc_318_p_spl_0),
    .din2(g943_n_spl_00)
  );


  andX
  g_g945_p
  (
    .dout(g945_p),
    .din1(g925_p_spl_),
    .din2(g943_p_spl_00)
  );


  andX
  g_g946_p
  (
    .dout(g946_p),
    .din1(ffc_14_p),
    .din2(ffc_41_p_spl_000)
  );


  andX
  g_g947_p
  (
    .dout(g947_p),
    .din1(ffc_41_n_spl_000),
    .din2(ffc_445_p_spl_00)
  );


  orX
  g_g948_n
  (
    .dout(g948_n),
    .din1(g946_p),
    .din2(g947_p)
  );


  andX
  g_g949_p
  (
    .dout(g949_p),
    .din1(ffc_41_p_spl_000),
    .din2(ffc_59_p)
  );


  andX
  g_g950_p
  (
    .dout(g950_p),
    .din1(ffc_41_n_spl_000),
    .din2(g925_n_spl_0)
  );


  orX
  g_g951_n
  (
    .dout(g951_n),
    .din1(g949_p),
    .din2(g950_p)
  );


  andX
  g_g952_p
  (
    .dout(g952_p),
    .din1(ffc_41_p_spl_00),
    .din2(ffc_56_p)
  );


  andX
  g_g953_p
  (
    .dout(g953_p),
    .din1(ffc_41_n_spl_00),
    .din2(g913_p_spl_0)
  );


  orX
  g_g954_n
  (
    .dout(g954_n),
    .din1(g952_p),
    .din2(g953_p)
  );


  andX
  g_g955_p
  (
    .dout(g955_p),
    .din1(ffc_68_p),
    .din2(ffc_74_p_spl_00)
  );


  andX
  g_g956_p
  (
    .dout(g956_p),
    .din1(ffc_74_n_spl_00),
    .din2(ffc_417_p_spl_0)
  );


  orX
  g_g957_n
  (
    .dout(g957_n),
    .din1(g955_p),
    .din2(g956_p)
  );


  andX
  g_g958_p
  (
    .dout(g958_p),
    .din1(ffc_74_p_spl_00),
    .din2(ffc_80_p)
  );


  andX
  g_g959_p
  (
    .dout(g959_p),
    .din1(ffc_74_n_spl_00),
    .din2(ffc_540_p_spl_0)
  );


  orX
  g_g960_n
  (
    .dout(g960_n),
    .din1(g958_p),
    .din2(g959_p)
  );


  andX
  g_g961_p
  (
    .dout(g961_p),
    .din1(ffc_74_p_spl_01),
    .din2(ffc_83_p)
  );


  andX
  g_g962_p
  (
    .dout(g962_p),
    .din1(ffc_74_n_spl_01),
    .din2(ffc_416_p_spl_0)
  );


  orX
  g_g963_n
  (
    .dout(g963_n),
    .din1(g961_p),
    .din2(g962_p)
  );


  andX
  g_g964_p
  (
    .dout(g964_p),
    .din1(ffc_425_n),
    .din2(ffc_505_p_spl_)
  );


  andX
  g_g965_p
  (
    .dout(g965_p),
    .din1(ffc_308_n_spl_00),
    .din2(g964_p_spl_0)
  );


  andX
  g_g966_p
  (
    .dout(g966_p),
    .din1(ffc_425_p),
    .din2(ffc_505_p_spl_)
  );


  andX
  g_g967_p
  (
    .dout(g967_p),
    .din1(ffc_346_n_spl_),
    .din2(g966_p_spl_0)
  );


  orX
  g_g968_n
  (
    .dout(g968_n),
    .din1(g965_p),
    .din2(g967_p)
  );


  andX
  g_g969_p
  (
    .dout(g969_p),
    .din1(ffc_404_p_spl_10),
    .din2(ffc_536_p)
  );


  orX
  g_g969_n
  (
    .dout(g969_n),
    .din1(ffc_404_n_spl_10),
    .din2(ffc_536_n)
  );


  andX
  g_g970_p
  (
    .dout(g970_p),
    .din1(ffc_404_n_spl_10),
    .din2(ffc_539_p)
  );


  orX
  g_g970_n
  (
    .dout(g970_n),
    .din1(ffc_404_p_spl_10),
    .din2(ffc_539_n)
  );


  andX
  g_g971_p
  (
    .dout(g971_p),
    .din1(g969_n),
    .din2(g970_n)
  );


  orX
  g_g971_n
  (
    .dout(g971_n),
    .din1(g969_p),
    .din2(g970_p)
  );


  andX
  g_g972_p
  (
    .dout(g972_p),
    .din1(g943_p_spl_00),
    .din2(g971_n_spl_0)
  );


  orX
  g_g972_n
  (
    .dout(g972_n),
    .din1(g943_n_spl_00),
    .din2(g971_p_spl_0)
  );


  andX
  g_g973_p
  (
    .dout(g973_p),
    .din1(ffc_428_n_spl_),
    .din2(g943_p_spl_0)
  );


  orX
  g_g973_n
  (
    .dout(g973_n),
    .din1(ffc_428_p_spl_0),
    .din2(g943_n_spl_0)
  );


  orX
  g_g974_n
  (
    .dout(g974_n),
    .din1(g972_p),
    .din2(g973_n)
  );


  andX
  g_g975_p
  (
    .dout(g975_p),
    .din1(ffc_445_p_spl_00),
    .din2(ffc_544_p_spl_00)
  );


  orX
  g_g975_n
  (
    .dout(g975_n),
    .din1(ffc_445_n_spl_),
    .din2(ffc_544_n_spl_)
  );


  andX
  g_g976_p
  (
    .dout(g976_p),
    .din1(ffc_445_n_spl_),
    .din2(ffc_544_n_spl_)
  );


  orX
  g_g976_n
  (
    .dout(g976_n),
    .din1(ffc_445_p_spl_0),
    .din2(ffc_544_p_spl_00)
  );


  andX
  g_g977_p
  (
    .dout(g977_p),
    .din1(g975_n),
    .din2(g976_n)
  );


  orX
  g_g977_n
  (
    .dout(g977_n),
    .din1(g975_p),
    .din2(g976_p)
  );


  andX
  g_g978_p
  (
    .dout(g978_p),
    .din1(g928_n_spl_),
    .din2(g977_p)
  );


  andX
  g_g979_p
  (
    .dout(g979_p),
    .din1(g928_p),
    .din2(g977_n)
  );


  orX
  g_g980_n
  (
    .dout(g980_n),
    .din1(g978_p),
    .din2(g979_p)
  );


  orX
  g_g981_n
  (
    .dout(g981_n),
    .din1(ffc_560_p),
    .din2(ffc_562_p)
  );


  andX
  g_g982_p
  (
    .dout(g982_p),
    .din1(ffc_533_p_spl_000),
    .din2(g981_n)
  );


  andX
  g_g983_p
  (
    .dout(g983_p),
    .din1(ffc_556_p),
    .din2(ffc_563_p_spl_00)
  );


  andX
  g_g984_p
  (
    .dout(g984_p),
    .din1(ffc_533_n_spl_00),
    .din2(ffc_561_p)
  );


  orX
  g_g985_n
  (
    .dout(g985_n),
    .din1(g983_p),
    .din2(g984_p)
  );


  orX
  g_g986_n
  (
    .dout(g986_n),
    .din1(g982_p),
    .din2(g985_n)
  );


  andX
  g_g987_p
  (
    .dout(g987_p),
    .din1(ffc_532_p_spl_000),
    .din2(ffc_558_p)
  );


  andX
  g_g988_p
  (
    .dout(g988_p),
    .din1(ffc_532_n_spl_000),
    .din2(ffc_555_p)
  );


  orX
  g_g989_n
  (
    .dout(g989_n),
    .din1(g987_p),
    .din2(g988_p)
  );


  andX
  g_g990_p
  (
    .dout(g990_p),
    .din1(ffc_533_p_spl_000),
    .din2(g989_n)
  );


  andX
  g_g991_p
  (
    .dout(g991_p),
    .din1(ffc_553_p),
    .din2(ffc_563_p_spl_00)
  );


  andX
  g_g992_p
  (
    .dout(g992_p),
    .din1(ffc_532_n_spl_000),
    .din2(ffc_557_p)
  );


  andX
  g_g993_p
  (
    .dout(g993_p),
    .din1(ffc_533_n_spl_00),
    .din2(g992_p)
  );


  orX
  g_g994_n
  (
    .dout(g994_n),
    .din1(g991_p),
    .din2(g993_p)
  );


  orX
  g_g995_n
  (
    .dout(g995_n),
    .din1(g990_p),
    .din2(g994_n)
  );


  andX
  g_g996_p
  (
    .dout(g996_p),
    .din1(ffc_71_p),
    .din2(ffc_74_p_spl_01)
  );


  andX
  g_g997_p
  (
    .dout(g997_p),
    .din1(ffc_74_n_spl_01),
    .din2(g938_n_spl_0)
  );


  andX
  g_g998_p
  (
    .dout(g998_p),
    .din1(ffc_99_p_spl_),
    .din2(ffc_163_p_spl_)
  );


  andX
  g_g999_p
  (
    .dout(g999_p),
    .din1(ffc_120_p_spl_),
    .din2(ffc_141_p_spl_)
  );


  andX
  g_g1000_p
  (
    .dout(g1000_p),
    .din1(ffc_190_p_spl_),
    .din2(ffc_244_p_spl_)
  );


  andX
  g_g1001_p
  (
    .dout(g1001_p),
    .din1(ffc_208_p_spl_),
    .din2(ffc_226_p_spl_)
  );


  orX
  g_g1002_n
  (
    .dout(g1002_n),
    .din1(ffc_269_p_spl_),
    .din2(ffc_445_p_spl_1)
  );


  andX
  g_g1003_p
  (
    .dout(g1003_p),
    .din1(ffc_41_p_spl_01),
    .din2(ffc_44_p)
  );


  andX
  g_g1004_p
  (
    .dout(g1004_p),
    .din1(ffc_41_n_spl_01),
    .din2(ffc_439_p_spl_1)
  );


  orX
  g_g1005_n
  (
    .dout(g1005_n),
    .din1(g1003_p),
    .din2(g1004_p)
  );


  orX
  g_g1006_n
  (
    .dout(g1006_n),
    .din1(ffc_422_n_spl_0),
    .din2(g1005_n_spl_)
  );


  andX
  g_g1007_p
  (
    .dout(g1007_p),
    .din1(ffc_422_n_spl_0),
    .din2(g1005_n_spl_)
  );


  orX
  g_g1008_n
  (
    .dout(g1008_n),
    .din1(ffc_423_n_spl_0),
    .din2(g948_n_spl_)
  );


  andX
  g_g1009_p
  (
    .dout(g1009_p),
    .din1(ffc_41_p_spl_01),
    .din2(ffc_47_p)
  );


  andX
  g_g1010_p
  (
    .dout(g1010_p),
    .din1(ffc_41_n_spl_01),
    .din2(ffc_544_p_spl_01)
  );


  orX
  g_g1011_n
  (
    .dout(g1011_n),
    .din1(g1009_p),
    .din2(g1010_p)
  );


  orX
  g_g1012_n
  (
    .dout(g1012_n),
    .din1(ffc_440_n_spl_0),
    .din2(g1011_n_spl_)
  );


  andX
  g_g1013_p
  (
    .dout(g1013_p),
    .din1(ffc_440_n_spl_0),
    .din2(g1011_n_spl_)
  );


  andX
  g_g1014_p
  (
    .dout(g1014_p),
    .din1(ffc_41_p_spl_10),
    .din2(ffc_50_p)
  );


  andX
  g_g1015_p
  (
    .dout(g1015_p),
    .din1(ffc_41_n_spl_10),
    .din2(g903_n_spl_0)
  );


  orX
  g_g1016_n
  (
    .dout(g1016_n),
    .din1(g1014_p),
    .din2(g1015_p)
  );


  andX
  g_g1017_p
  (
    .dout(g1017_p),
    .din1(ffc_305_n_spl_0),
    .din2(g1016_n_spl_)
  );


  orX
  g_g1018_n
  (
    .dout(g1018_n),
    .din1(ffc_305_n_spl_0),
    .din2(g1016_n_spl_)
  );


  andX
  g_g1019_p
  (
    .dout(g1019_p),
    .din1(ffc_41_p_spl_10),
    .din2(ffc_53_p)
  );


  andX
  g_g1020_p
  (
    .dout(g1020_p),
    .din1(ffc_41_n_spl_10),
    .din2(g908_n_spl_0)
  );


  orX
  g_g1021_n
  (
    .dout(g1021_n),
    .din1(g1019_p),
    .din2(g1020_p)
  );


  andX
  g_g1022_p
  (
    .dout(g1022_p),
    .din1(ffc_308_n_spl_00),
    .din2(g1021_n_spl_)
  );


  orX
  g_g1023_n
  (
    .dout(g1023_n),
    .din1(ffc_308_n_spl_0),
    .din2(g1021_n_spl_)
  );


  andX
  g_g1024_p
  (
    .dout(g1024_p),
    .din1(ffc_311_n_spl_0),
    .din2(g954_n_spl_)
  );


  andX
  g_g1025_p
  (
    .dout(g1025_p),
    .din1(ffc_311_n_spl_0),
    .din2(g964_p_spl_0)
  );


  andX
  g_g1026_p
  (
    .dout(g1026_p),
    .din1(ffc_20_p),
    .din2(ffc_41_p_spl_11)
  );


  andX
  g_g1027_p
  (
    .dout(g1027_p),
    .din1(ffc_41_n_spl_11),
    .din2(g919_n_spl_0)
  );


  orX
  g_g1028_n
  (
    .dout(g1028_n),
    .din1(g1026_p),
    .din2(g1027_p)
  );


  andX
  g_g1029_p
  (
    .dout(g1029_p),
    .din1(ffc_315_n_spl_0),
    .din2(g1028_n_spl_)
  );


  orX
  g_g1030_n
  (
    .dout(g1030_n),
    .din1(ffc_315_n_spl_0),
    .din2(g1028_n_spl_)
  );


  andX
  g_g1031_p
  (
    .dout(g1031_p),
    .din1(ffc_315_n_spl_1),
    .din2(g964_p_spl_1)
  );


  orX
  g_g1032_n
  (
    .dout(g1032_n),
    .din1(ffc_318_n_spl_),
    .din2(g951_n_spl_)
  );


  andX
  g_g1033_p
  (
    .dout(g1033_p),
    .din1(ffc_442_n_spl_0),
    .din2(g960_n_spl_)
  );


  orX
  g_g1034_n
  (
    .dout(g1034_n),
    .din1(ffc_443_n_spl_0),
    .din2(g957_n_spl_)
  );


  andX
  g_g1035_p
  (
    .dout(g1035_p),
    .din1(ffc_342_n_spl_0),
    .din2(g963_n_spl_)
  );


  andX
  g_g1036_p
  (
    .dout(g1036_p),
    .din1(ffc_350_p_spl_),
    .din2(ffc_354_n)
  );


  andX
  g_g1037_p
  (
    .dout(g1037_p),
    .din1(ffc_350_n),
    .din2(ffc_354_p_spl_)
  );


  andX
  g_g1038_p
  (
    .dout(g1038_p),
    .din1(g919_p_spl_),
    .din2(g966_p_spl_0)
  );


  andX
  g_g1039_p
  (
    .dout(g1039_p),
    .din1(g913_n_spl_),
    .din2(g966_p_spl_1)
  );


  orX
  g_g1040_n
  (
    .dout(g1040_n),
    .din1(ffc_132_n),
    .din2(ffc_563_n)
  );


  andX
  g_g1041_p
  (
    .dout(g1041_p),
    .din1(ffc_17_p),
    .din2(ffc_41_p_spl_11)
  );


  andX
  g_g1042_p
  (
    .dout(g1042_p),
    .din1(ffc_41_n_spl_11),
    .din2(ffc_546_p_spl_0)
  );


  orX
  g_g1043_n
  (
    .dout(g1043_n),
    .din1(g1041_p),
    .din2(g1042_p)
  );


  orX
  g_g1044_n
  (
    .dout(g1044_n),
    .din1(g942_n_spl_),
    .din2(g968_n_spl_)
  );


  andX
  g_g1045_p
  (
    .dout(g1045_p),
    .din1(ffc_62_p),
    .din2(ffc_74_p_spl_10)
  );


  andX
  g_g1046_p
  (
    .dout(g1046_p),
    .din1(ffc_74_n_spl_10),
    .din2(ffc_541_p_spl_0)
  );


  orX
  g_g1047_n
  (
    .dout(g1047_n),
    .din1(g1045_p),
    .din2(g1046_p)
  );


  andX
  g_g1048_p
  (
    .dout(g1048_p),
    .din1(ffc_65_p),
    .din2(ffc_74_p_spl_10)
  );


  andX
  g_g1049_p
  (
    .dout(g1049_p),
    .din1(ffc_404_p_spl_11),
    .din2(ffc_535_p)
  );


  orX
  g_g1049_n
  (
    .dout(g1049_n),
    .din1(ffc_404_n_spl_11),
    .din2(ffc_535_n)
  );


  andX
  g_g1050_p
  (
    .dout(g1050_p),
    .din1(ffc_404_n_spl_11),
    .din2(ffc_538_p)
  );


  orX
  g_g1050_n
  (
    .dout(g1050_n),
    .din1(ffc_404_p_spl_11),
    .din2(ffc_538_n)
  );


  andX
  g_g1051_p
  (
    .dout(g1051_p),
    .din1(g1049_n),
    .din2(g1050_n)
  );


  orX
  g_g1051_n
  (
    .dout(g1051_n),
    .din1(g1049_p),
    .din2(g1050_p)
  );


  andX
  g_g1052_p
  (
    .dout(g1052_p),
    .din1(ffc_74_n_spl_10),
    .din2(g1051_n_spl_0)
  );


  orX
  g_g1053_n
  (
    .dout(g1053_n),
    .din1(g1048_p),
    .din2(g1052_p)
  );


  andX
  g_g1054_p
  (
    .dout(g1054_p),
    .din1(ffc_74_p_spl_11),
    .din2(ffc_86_p)
  );


  andX
  g_g1055_p
  (
    .dout(g1055_p),
    .din1(g897_n),
    .din2(g898_n)
  );


  orX
  g_g1055_n
  (
    .dout(g1055_n),
    .din1(g897_p_spl_),
    .din2(g898_p_spl_)
  );


  andX
  g_g1056_p
  (
    .dout(g1056_p),
    .din1(ffc_74_n_spl_11),
    .din2(g1055_n_spl_0)
  );


  orX
  g_g1057_n
  (
    .dout(g1057_n),
    .din1(g1054_p),
    .din2(g1056_p)
  );


  andX
  g_g1058_p
  (
    .dout(g1058_p),
    .din1(ffc_74_p_spl_11),
    .din2(ffc_77_p)
  );


  andX
  g_g1059_p
  (
    .dout(g1059_p),
    .din1(ffc_74_n_spl_11),
    .din2(g971_n_spl_0)
  );


  orX
  g_g1060_n
  (
    .dout(g1060_n),
    .din1(g1058_p),
    .din2(g1059_p)
  );


  andX
  g_g1061_p
  (
    .dout(g1061_p),
    .din1(ffc_305_n_spl_1),
    .din2(ffc_441_p_spl_)
  );


  andX
  g_g1062_p
  (
    .dout(g1062_p),
    .din1(ffc_305_p),
    .din2(ffc_441_n)
  );


  orX
  g_g1063_n
  (
    .dout(g1063_n),
    .din1(g1061_p),
    .din2(g1062_p)
  );


  andX
  g_g1064_p
  (
    .dout(g1064_p),
    .din1(ffc_315_p),
    .din2(ffc_318_n_spl_)
  );


  andX
  g_g1065_p
  (
    .dout(g1065_p),
    .din1(ffc_315_n_spl_1),
    .din2(ffc_318_p_spl_0)
  );


  orX
  g_g1066_n
  (
    .dout(g1066_n),
    .din1(g1064_p),
    .din2(g1065_p)
  );


  orX
  g_g1067_n
  (
    .dout(g1067_n),
    .din1(g944_n_spl_),
    .din2(g945_p_spl_)
  );


  andX
  g_g1068_p
  (
    .dout(g1068_p),
    .din1(ffc_322_p_spl_),
    .din2(ffc_428_n_spl_)
  );


  andX
  g_g1069_p
  (
    .dout(g1069_p),
    .din1(ffc_322_n_spl_),
    .din2(ffc_428_p_spl_0)
  );


  orX
  g_g1070_n
  (
    .dout(g1070_n),
    .din1(g1068_p),
    .din2(g1069_p)
  );


  orX
  g_g1071_n
  (
    .dout(g1071_n),
    .din1(ffc_541_n_spl_0),
    .din2(g943_n_spl_1)
  );


  andX
  g_g1072_p
  (
    .dout(g1072_p),
    .din1(ffc_322_n_spl_),
    .din2(g943_p_spl_1)
  );


  andX
  g_g1073_p
  (
    .dout(g1073_p),
    .din1(g1071_n_spl_),
    .din2(g1072_p_spl_)
  );


  orX
  g_g1074_n
  (
    .dout(g1074_n),
    .din1(g1071_n_spl_),
    .din2(g1072_p_spl_)
  );


  orX
  g_g1075_n
  (
    .dout(g1075_n),
    .din1(g943_n_spl_1),
    .din2(g1051_n_spl_0)
  );


  andX
  g_g1076_p
  (
    .dout(g1076_p),
    .din1(ffc_424_n_spl_0),
    .din2(g943_p_spl_1)
  );


  andX
  g_g1077_p
  (
    .dout(g1077_p),
    .din1(g1075_n_spl_),
    .din2(g1076_p_spl_)
  );


  orX
  g_g1078_n
  (
    .dout(g1078_n),
    .din1(g1075_n_spl_),
    .din2(g1076_p_spl_)
  );


  orX
  g_g1079_n
  (
    .dout(g1079_n),
    .din1(ffc_505_n_spl_),
    .din2(g903_n_spl_0)
  );


  andX
  g_g1080_p
  (
    .dout(g1080_p),
    .din1(ffc_305_n_spl_1),
    .din2(g964_p_spl_1)
  );


  andX
  g_g1081_p
  (
    .dout(g1081_p),
    .din1(ffc_342_n_spl_),
    .din2(g966_p_spl_1)
  );


  orX
  g_g1082_n
  (
    .dout(g1082_n),
    .din1(g1080_p),
    .din2(g1081_p)
  );


  andX
  g_g1083_p
  (
    .dout(g1083_p),
    .din1(g1079_n_spl_),
    .din2(g1082_n_spl_)
  );


  orX
  g_g1084_n
  (
    .dout(g1084_n),
    .din1(g1079_n_spl_),
    .din2(g1082_n_spl_)
  );


  andX
  g_g1085_p
  (
    .dout(g1085_p),
    .din1(ffc_546_p_spl_0),
    .din2(ffc_548_n_spl_)
  );


  andX
  g_g1086_p
  (
    .dout(g1086_p),
    .din1(ffc_544_p_spl_01),
    .din2(ffc_547_n_spl_)
  );


  andX
  g_g1087_p
  (
    .dout(g1087_p),
    .din1(ffc_531_n),
    .din2(ffc_549_n)
  );


  orX
  g_g1088_n
  (
    .dout(g1088_n),
    .din1(g1086_p),
    .din2(g1087_p)
  );


  orX
  g_g1089_n
  (
    .dout(g1089_n),
    .din1(ffc_546_p_spl_1),
    .din2(ffc_548_n_spl_)
  );


  orX
  g_g1090_n
  (
    .dout(g1090_n),
    .din1(ffc_544_p_spl_1),
    .din2(ffc_547_n_spl_)
  );


  andX
  g_g1091_p
  (
    .dout(g1091_p),
    .din1(g1089_n),
    .din2(g1090_n)
  );


  andX
  g_g1092_p
  (
    .dout(g1092_p),
    .din1(g1088_n),
    .din2(g1091_p)
  );


  orX
  g_g1093_n
  (
    .dout(g1093_n),
    .din1(g1085_p),
    .din2(g1092_p)
  );


  andX
  g_g1094_p
  (
    .dout(g1094_p),
    .din1(g1084_n),
    .din2(g1093_n)
  );


  orX
  g_g1095_n
  (
    .dout(g1095_n),
    .din1(g1083_p),
    .din2(g1094_p)
  );


  orX
  g_g1096_n
  (
    .dout(g1096_n),
    .din1(g972_n),
    .din2(g973_p)
  );


  andX
  g_g1097_p
  (
    .dout(g1097_p),
    .din1(g974_n_spl_),
    .din2(g1096_n)
  );


  orX
  g_g1098_n
  (
    .dout(g1098_n),
    .din1(ffc_342_p_spl_),
    .din2(ffc_346_p_spl_)
  );


  andX
  g_g1099_p
  (
    .dout(g1099_p),
    .din1(g929_n_spl_),
    .din2(g1098_n)
  );


  andX
  g_g1100_p
  (
    .dout(g1100_p),
    .din1(ffc_442_n_spl_),
    .din2(ffc_443_n_spl_)
  );


  orX
  g_g1100_n
  (
    .dout(g1100_n),
    .din1(ffc_442_p_spl_0),
    .din2(ffc_443_p_spl_0)
  );


  andX
  g_g1101_p
  (
    .dout(g1101_p),
    .din1(g902_n),
    .din2(g1100_n)
  );


  orX
  g_g1101_n
  (
    .dout(g1101_n),
    .din1(g902_p_spl_),
    .din2(g1100_p)
  );


  andX
  g_g1102_p
  (
    .dout(g1102_p),
    .din1(ffc_386_n_spl_),
    .din2(ffc_424_n_spl_0)
  );


  orX
  g_g1102_n
  (
    .dout(g1102_n),
    .din1(ffc_386_p_spl_),
    .din2(ffc_424_p_spl_0)
  );


  andX
  g_g1103_p
  (
    .dout(g1103_p),
    .din1(ffc_386_p_spl_),
    .din2(ffc_424_p_spl_0)
  );


  orX
  g_g1103_n
  (
    .dout(g1103_n),
    .din1(ffc_386_n_spl_),
    .din2(ffc_424_n_spl_)
  );


  andX
  g_g1104_p
  (
    .dout(g1104_p),
    .din1(g1102_n),
    .din2(g1103_n)
  );


  orX
  g_g1104_n
  (
    .dout(g1104_n),
    .din1(g1102_p),
    .din2(g1103_p)
  );


  orX
  g_g1105_n
  (
    .dout(g1105_n),
    .din1(g1101_p),
    .din2(g1104_n)
  );


  orX
  g_g1106_n
  (
    .dout(g1106_n),
    .din1(g1101_n),
    .din2(g1104_p)
  );


  andX
  g_g1107_p
  (
    .dout(g1107_p),
    .din1(g1105_n),
    .din2(g1106_n)
  );


  orX
  g_g1108_n
  (
    .dout(g1108_n),
    .din1(g1099_p_spl_),
    .din2(g1107_p_spl_)
  );


  andX
  g_g1109_p
  (
    .dout(g1109_p),
    .din1(g1099_p_spl_),
    .din2(g1107_p_spl_)
  );


  andX
  g_g1110_p
  (
    .dout(g1110_p),
    .din1(g903_n_spl_1),
    .din2(g907_n_spl_)
  );


  andX
  g_g1111_p
  (
    .dout(g1111_p),
    .din1(g903_p),
    .din2(g907_p)
  );


  orX
  g_g1112_n
  (
    .dout(g1112_n),
    .din1(g1110_p),
    .din2(g1111_p)
  );


  andX
  g_g1113_p
  (
    .dout(g1113_p),
    .din1(g980_n_spl_0),
    .din2(g1112_n_spl_)
  );


  orX
  g_g1114_n
  (
    .dout(g1114_n),
    .din1(g980_n_spl_0),
    .din2(g1112_n_spl_)
  );


  andX
  g_g1115_p
  (
    .dout(g1115_p),
    .din1(ffc_377_p_spl_),
    .din2(ffc_380_n_spl_)
  );


  orX
  g_g1115_n
  (
    .dout(g1115_n),
    .din1(ffc_377_n_spl_),
    .din2(ffc_380_p_spl_)
  );


  andX
  g_g1116_p
  (
    .dout(g1116_p),
    .din1(ffc_377_n_spl_),
    .din2(ffc_380_p_spl_)
  );


  orX
  g_g1116_n
  (
    .dout(g1116_n),
    .din1(ffc_377_p_spl_),
    .din2(ffc_380_n_spl_)
  );


  andX
  g_g1117_p
  (
    .dout(g1117_p),
    .din1(g1115_n),
    .din2(g1116_n)
  );


  orX
  g_g1117_n
  (
    .dout(g1117_n),
    .din1(g1115_p),
    .din2(g1116_p)
  );


  andX
  g_g1118_p
  (
    .dout(g1118_p),
    .din1(ffc_422_p_spl_),
    .din2(ffc_423_n_spl_0)
  );


  orX
  g_g1118_n
  (
    .dout(g1118_n),
    .din1(ffc_422_n_spl_1),
    .din2(ffc_423_p_spl_0)
  );


  andX
  g_g1119_p
  (
    .dout(g1119_p),
    .din1(ffc_422_n_spl_1),
    .din2(ffc_423_p_spl_0)
  );


  orX
  g_g1119_n
  (
    .dout(g1119_n),
    .din1(ffc_422_p_spl_),
    .din2(ffc_423_n_spl_)
  );


  andX
  g_g1120_p
  (
    .dout(g1120_p),
    .din1(g1118_n),
    .din2(g1119_n)
  );


  orX
  g_g1120_n
  (
    .dout(g1120_n),
    .din1(g1118_p),
    .din2(g1119_p)
  );


  andX
  g_g1121_p
  (
    .dout(g1121_p),
    .din1(g1117_n),
    .din2(g1120_p)
  );


  andX
  g_g1122_p
  (
    .dout(g1122_p),
    .din1(g1117_p),
    .din2(g1120_n)
  );


  orX
  g_g1123_n
  (
    .dout(g1123_n),
    .din1(g1121_p),
    .din2(g1122_p)
  );


  andX
  g_g1124_p
  (
    .dout(g1124_p),
    .din1(ffc_308_p_spl_),
    .din2(ffc_311_n_spl_1)
  );


  orX
  g_g1124_n
  (
    .dout(g1124_n),
    .din1(ffc_308_n_spl_1),
    .din2(ffc_311_p_spl_0)
  );


  andX
  g_g1125_p
  (
    .dout(g1125_p),
    .din1(ffc_308_n_spl_1),
    .din2(ffc_311_p_spl_0)
  );


  orX
  g_g1125_n
  (
    .dout(g1125_n),
    .din1(ffc_308_p_spl_),
    .din2(ffc_311_n_spl_1)
  );


  andX
  g_g1126_p
  (
    .dout(g1126_p),
    .din1(g1124_n),
    .din2(g1125_n)
  );


  orX
  g_g1126_n
  (
    .dout(g1126_n),
    .din1(g1124_p),
    .din2(g1125_p)
  );


  andX
  g_g1127_p
  (
    .dout(g1127_p),
    .din1(ffc_383_n_spl_),
    .din2(ffc_440_n_spl_1)
  );


  orX
  g_g1127_n
  (
    .dout(g1127_n),
    .din1(ffc_383_p_spl_),
    .din2(ffc_440_p_spl_)
  );


  andX
  g_g1128_p
  (
    .dout(g1128_p),
    .din1(ffc_383_p_spl_),
    .din2(ffc_440_p_spl_)
  );


  orX
  g_g1128_n
  (
    .dout(g1128_n),
    .din1(ffc_383_n_spl_),
    .din2(ffc_440_n_spl_1)
  );


  andX
  g_g1129_p
  (
    .dout(g1129_p),
    .din1(g1127_n),
    .din2(g1128_n)
  );


  orX
  g_g1129_n
  (
    .dout(g1129_n),
    .din1(g1127_p),
    .din2(g1128_p)
  );


  andX
  g_g1130_p
  (
    .dout(g1130_p),
    .din1(g1126_p),
    .din2(g1129_p)
  );


  andX
  g_g1131_p
  (
    .dout(g1131_p),
    .din1(g1126_n),
    .din2(g1129_n)
  );


  orX
  g_g1132_n
  (
    .dout(g1132_n),
    .din1(g1130_p),
    .din2(g1131_p)
  );


  andX
  g_g1133_p
  (
    .dout(g1133_p),
    .din1(ffc_416_n_spl_),
    .din2(g1055_n_spl_0)
  );


  orX
  g_g1133_n
  (
    .dout(g1133_n),
    .din1(ffc_416_p_spl_0),
    .din2(g1055_p_spl_)
  );


  andX
  g_g1134_p
  (
    .dout(g1134_p),
    .din1(ffc_416_p_spl_),
    .din2(g1055_p_spl_)
  );


  orX
  g_g1134_n
  (
    .dout(g1134_n),
    .din1(ffc_416_n_spl_),
    .din2(g1055_n_spl_)
  );


  andX
  g_g1135_p
  (
    .dout(g1135_p),
    .din1(g1133_n),
    .din2(g1134_n)
  );


  orX
  g_g1135_n
  (
    .dout(g1135_n),
    .din1(g1133_p),
    .din2(g1134_p)
  );


  orX
  g_g1136_n
  (
    .dout(g1136_n),
    .din1(g938_p),
    .din2(g1135_p)
  );


  orX
  g_g1137_n
  (
    .dout(g1137_n),
    .din1(g938_n_spl_0),
    .din2(g1135_n)
  );


  andX
  g_g1138_p
  (
    .dout(g1138_p),
    .din1(g1136_n),
    .din2(g1137_n)
  );


  andX
  g_g1139_p
  (
    .dout(g1139_p),
    .din1(ffc_516_p_spl_),
    .din2(ffc_517_n_spl_)
  );


  orX
  g_g1139_n
  (
    .dout(g1139_n),
    .din1(ffc_516_n_spl_),
    .din2(ffc_517_p_spl_)
  );


  andX
  g_g1140_p
  (
    .dout(g1140_p),
    .din1(ffc_516_n_spl_),
    .din2(ffc_517_p_spl_)
  );


  orX
  g_g1140_n
  (
    .dout(g1140_n),
    .din1(ffc_516_p_spl_),
    .din2(ffc_517_n_spl_)
  );


  andX
  g_g1141_p
  (
    .dout(g1141_p),
    .din1(g1139_n),
    .din2(g1140_n)
  );


  orX
  g_g1141_n
  (
    .dout(g1141_n),
    .din1(g1139_p),
    .din2(g1140_p)
  );


  andX
  g_g1142_p
  (
    .dout(g1142_p),
    .din1(ffc_514_p_spl_),
    .din2(ffc_515_n_spl_)
  );


  orX
  g_g1142_n
  (
    .dout(g1142_n),
    .din1(ffc_514_n_spl_),
    .din2(ffc_515_p_spl_)
  );


  andX
  g_g1143_p
  (
    .dout(g1143_p),
    .din1(ffc_514_n_spl_),
    .din2(ffc_515_p_spl_)
  );


  orX
  g_g1143_n
  (
    .dout(g1143_n),
    .din1(ffc_514_p_spl_),
    .din2(ffc_515_n_spl_)
  );


  andX
  g_g1144_p
  (
    .dout(g1144_p),
    .din1(g1142_n),
    .din2(g1143_n)
  );


  orX
  g_g1144_n
  (
    .dout(g1144_n),
    .din1(g1142_p),
    .din2(g1143_p)
  );


  andX
  g_g1145_p
  (
    .dout(g1145_p),
    .din1(g1141_p_spl_),
    .din2(g1144_p_spl_)
  );


  orX
  g_g1145_n
  (
    .dout(g1145_n),
    .din1(g1141_n_spl_),
    .din2(g1144_n_spl_)
  );


  andX
  g_g1146_p
  (
    .dout(g1146_p),
    .din1(g1141_n_spl_),
    .din2(g1144_n_spl_)
  );


  orX
  g_g1146_n
  (
    .dout(g1146_n),
    .din1(g1141_p_spl_),
    .din2(g1144_p_spl_)
  );


  andX
  g_g1147_p
  (
    .dout(g1147_p),
    .din1(g1145_n),
    .din2(g1146_n)
  );


  orX
  g_g1147_n
  (
    .dout(g1147_n),
    .din1(g1145_p),
    .din2(g1146_p)
  );


  andX
  g_g1148_p
  (
    .dout(g1148_p),
    .din1(ffc_367_p_spl_),
    .din2(ffc_370_n_spl_)
  );


  orX
  g_g1148_n
  (
    .dout(g1148_n),
    .din1(ffc_367_n_spl_),
    .din2(ffc_370_p_spl_)
  );


  andX
  g_g1149_p
  (
    .dout(g1149_p),
    .din1(ffc_367_n_spl_),
    .din2(ffc_370_p_spl_)
  );


  orX
  g_g1149_n
  (
    .dout(g1149_n),
    .din1(ffc_367_p_spl_),
    .din2(ffc_370_n_spl_)
  );


  andX
  g_g1150_p
  (
    .dout(g1150_p),
    .din1(g1148_n),
    .din2(g1149_n)
  );


  orX
  g_g1150_n
  (
    .dout(g1150_n),
    .din1(g1148_p),
    .din2(g1149_p)
  );


  orX
  g_g1151_n
  (
    .dout(g1151_n),
    .din1(g1147_p),
    .din2(g1150_n)
  );


  orX
  g_g1152_n
  (
    .dout(g1152_n),
    .din1(g1147_n),
    .din2(g1150_p)
  );


  andX
  g_g1153_p
  (
    .dout(g1153_p),
    .din1(g1151_n),
    .din2(g1152_n)
  );


  andX
  g_g1154_p
  (
    .dout(g1154_p),
    .din1(g908_p),
    .din2(g913_p_spl_0)
  );


  andX
  g_g1155_p
  (
    .dout(g1155_p),
    .din1(g908_n_spl_1),
    .din2(g913_n_spl_)
  );


  orX
  g_g1156_n
  (
    .dout(g1156_n),
    .din1(g1154_p),
    .din2(g1155_p)
  );


  orX
  g_g1157_n
  (
    .dout(g1157_n),
    .din1(g919_n_spl_0),
    .din2(g925_p_spl_)
  );


  orX
  g_g1158_n
  (
    .dout(g1158_n),
    .din1(g919_p_spl_),
    .din2(g925_n_spl_0)
  );


  andX
  g_g1159_p
  (
    .dout(g1159_p),
    .din1(g1157_n),
    .din2(g1158_n)
  );


  andX
  g_g1160_p
  (
    .dout(g1160_p),
    .din1(g1156_n_spl_),
    .din2(g1159_p_spl_)
  );


  orX
  g_g1161_n
  (
    .dout(g1161_n),
    .din1(g1156_n_spl_),
    .din2(g1159_p_spl_)
  );


  andX
  g_g1162_p
  (
    .dout(g1162_p),
    .din1(ffc_541_p_spl_0),
    .din2(ffc_542_p_spl_)
  );


  orX
  g_g1162_n
  (
    .dout(g1162_n),
    .din1(ffc_541_n_spl_0),
    .din2(ffc_542_n_spl_)
  );


  andX
  g_g1163_p
  (
    .dout(g1163_p),
    .din1(ffc_541_n_spl_),
    .din2(ffc_542_n_spl_)
  );


  orX
  g_g1163_n
  (
    .dout(g1163_n),
    .din1(ffc_541_p_spl_),
    .din2(ffc_542_p_spl_)
  );


  andX
  g_g1164_p
  (
    .dout(g1164_p),
    .din1(g1162_n),
    .din2(g1163_n)
  );


  orX
  g_g1164_n
  (
    .dout(g1164_n),
    .din1(g1162_p),
    .din2(g1163_p)
  );


  andX
  g_g1165_p
  (
    .dout(g1165_p),
    .din1(ffc_417_n_spl_),
    .din2(ffc_540_p_spl_0)
  );


  orX
  g_g1165_n
  (
    .dout(g1165_n),
    .din1(ffc_417_p_spl_0),
    .din2(ffc_540_n_spl_)
  );


  andX
  g_g1166_p
  (
    .dout(g1166_p),
    .din1(ffc_417_p_spl_1),
    .din2(ffc_540_n_spl_)
  );


  orX
  g_g1166_n
  (
    .dout(g1166_n),
    .din1(ffc_417_n_spl_),
    .din2(ffc_540_p_spl_)
  );


  andX
  g_g1167_p
  (
    .dout(g1167_p),
    .din1(g1165_n),
    .din2(g1166_n)
  );


  orX
  g_g1167_n
  (
    .dout(g1167_n),
    .din1(g1165_p),
    .din2(g1166_p)
  );


  andX
  g_g1168_p
  (
    .dout(g1168_p),
    .din1(g1164_p_spl_),
    .din2(g1167_p_spl_)
  );


  orX
  g_g1168_n
  (
    .dout(g1168_n),
    .din1(g1164_n_spl_),
    .din2(g1167_n_spl_)
  );


  andX
  g_g1169_p
  (
    .dout(g1169_p),
    .din1(g1164_n_spl_),
    .din2(g1167_n_spl_)
  );


  orX
  g_g1169_n
  (
    .dout(g1169_n),
    .din1(g1164_p_spl_),
    .din2(g1167_p_spl_)
  );


  andX
  g_g1170_p
  (
    .dout(g1170_p),
    .din1(g1168_n),
    .din2(g1169_n)
  );


  orX
  g_g1170_n
  (
    .dout(g1170_n),
    .din1(g1168_p),
    .din2(g1169_p)
  );


  andX
  g_g1171_p
  (
    .dout(g1171_p),
    .din1(g971_n_spl_1),
    .din2(g1051_p_spl_)
  );


  orX
  g_g1171_n
  (
    .dout(g1171_n),
    .din1(g971_p_spl_0),
    .din2(g1051_n_spl_1)
  );


  andX
  g_g1172_p
  (
    .dout(g1172_p),
    .din1(g971_p_spl_),
    .din2(g1051_n_spl_1)
  );


  orX
  g_g1172_n
  (
    .dout(g1172_n),
    .din1(g971_n_spl_1),
    .din2(g1051_p_spl_)
  );


  andX
  g_g1173_p
  (
    .dout(g1173_p),
    .din1(g1171_n),
    .din2(g1172_n)
  );


  orX
  g_g1173_n
  (
    .dout(g1173_n),
    .din1(g1171_p),
    .din2(g1172_p)
  );


  andX
  g_g1174_p
  (
    .dout(g1174_p),
    .din1(g1170_n),
    .din2(g1173_p)
  );


  andX
  g_g1175_p
  (
    .dout(g1175_p),
    .din1(g1170_p),
    .din2(g1173_n)
  );


  orX
  g_g1176_n
  (
    .dout(g1176_n),
    .din1(g1174_p),
    .din2(g1175_p)
  );


  orX
  g_g1177_n
  (
    .dout(g1177_n),
    .din1(ffc_154_n),
    .din2(ffc_532_p_spl_000)
  );


  andX
  g_g1178_p
  (
    .dout(g1178_p),
    .din1(ffc_533_n_spl_0),
    .din2(g1177_n)
  );


  andX
  g_g1179_p
  (
    .dout(g1179_p),
    .din1(ffc_532_n_spl_001),
    .din2(ffc_552_n)
  );


  andX
  g_g1180_p
  (
    .dout(g1180_p),
    .din1(ffc_533_p_spl_001),
    .din2(g1179_p)
  );


  andX
  g_g1181_p
  (
    .dout(g1181_p),
    .din1(ffc_176_n),
    .din2(ffc_532_p_spl_001)
  );


  orX
  g_g1182_n
  (
    .dout(g1182_n),
    .din1(g1180_p),
    .din2(g1181_p)
  );


  orX
  g_g1183_n
  (
    .dout(g1183_n),
    .din1(g1178_p),
    .din2(g1182_n)
  );


  andX
  g_g1184_p
  (
    .dout(g1184_p),
    .din1(ffc_102_p),
    .din2(ffc_532_n_spl_001)
  );


  andX
  g_g1185_p
  (
    .dout(g1185_p),
    .din1(ffc_104_p),
    .din2(ffc_532_n_spl_010)
  );


  andX
  g_g1186_p
  (
    .dout(g1186_p),
    .din1(ffc_144_p),
    .din2(ffc_532_n_spl_010)
  );


  andX
  g_g1187_p
  (
    .dout(g1187_p),
    .din1(ffc_146_p),
    .din2(ffc_532_n_spl_011)
  );


  andX
  g_g1188_p
  (
    .dout(g1188_p),
    .din1(ffc_150_p),
    .din2(ffc_532_n_spl_011)
  );


  andX
  g_g1189_p
  (
    .dout(g1189_p),
    .din1(ffc_166_p),
    .din2(ffc_532_p_spl_001)
  );


  andX
  g_g1190_p
  (
    .dout(g1190_p),
    .din1(ffc_168_p),
    .din2(ffc_532_p_spl_01)
  );


  andX
  g_g1191_p
  (
    .dout(g1191_p),
    .din1(ffc_172_n),
    .din2(ffc_532_p_spl_01)
  );


  andX
  g_g1192_p
  (
    .dout(g1192_p),
    .din1(ffc_106_n),
    .din2(ffc_533_p_spl_001)
  );


  orX
  g_g1193_n
  (
    .dout(g1193_n),
    .din1(ffc_148_p),
    .din2(ffc_533_p_spl_010)
  );


  andX
  g_g1194_p
  (
    .dout(g1194_p),
    .din1(ffc_108_n),
    .din2(ffc_532_n_spl_100)
  );


  andX
  g_g1195_p
  (
    .dout(g1195_p),
    .din1(ffc_533_p_spl_010),
    .din2(g1194_p)
  );


  andX
  g_g1196_p
  (
    .dout(g1196_p),
    .din1(ffc_152_p),
    .din2(ffc_532_n_spl_100)
  );


  orX
  g_g1197_n
  (
    .dout(g1197_n),
    .din1(ffc_533_p_spl_01),
    .din2(g1196_p)
  );


  andX
  g_g1198_p
  (
    .dout(g1198_p),
    .din1(ffc_181_p),
    .din2(ffc_532_p_spl_10)
  );


  andX
  g_g1199_p
  (
    .dout(g1199_p),
    .din1(ffc_116_p),
    .din2(ffc_532_n_spl_101)
  );


  orX
  g_g1200_n
  (
    .dout(g1200_n),
    .din1(g1198_p),
    .din2(g1199_p)
  );


  andX
  g_g1201_p
  (
    .dout(g1201_p),
    .din1(ffc_533_p_spl_10),
    .din2(g1200_n)
  );


  orX
  g_g1202_n
  (
    .dout(g1202_n),
    .din1(ffc_332_p_spl_),
    .din2(g941_n_spl_0)
  );


  orX
  g_g1203_n
  (
    .dout(g1203_n),
    .din1(ffc_295_p_spl_),
    .din2(g941_p_spl_00)
  );


  andX
  g_g1204_p
  (
    .dout(g1204_p),
    .din1(g1202_n),
    .din2(g1203_n)
  );


  andX
  g_g1205_p
  (
    .dout(g1205_p),
    .din1(g995_n_spl_0),
    .din2(g1204_p_spl_)
  );


  andX
  g_g1206_p
  (
    .dout(g1206_p),
    .din1(ffc_195_p),
    .din2(ffc_444_n_spl_000)
  );


  andX
  g_g1207_p
  (
    .dout(g1207_p),
    .din1(ffc_249_p),
    .din2(ffc_444_p_spl_000)
  );


  orX
  g_g1208_n
  (
    .dout(g1208_n),
    .din1(g1206_p),
    .din2(g1207_p)
  );


  andX
  g_g1209_p
  (
    .dout(g1209_p),
    .din1(ffc_199_p),
    .din2(ffc_444_n_spl_000)
  );


  andX
  g_g1210_p
  (
    .dout(g1210_p),
    .din1(ffc_253_p),
    .din2(ffc_444_p_spl_000)
  );


  orX
  g_g1211_n
  (
    .dout(g1211_n),
    .din1(g1209_p),
    .din2(g1210_p)
  );


  andX
  g_g1212_p
  (
    .dout(g1212_p),
    .din1(ffc_201_p),
    .din2(ffc_444_n_spl_001)
  );


  andX
  g_g1213_p
  (
    .dout(g1213_p),
    .din1(ffc_255_p),
    .din2(ffc_444_p_spl_001)
  );


  orX
  g_g1214_n
  (
    .dout(g1214_n),
    .din1(g1212_p),
    .din2(g1213_p)
  );


  andX
  g_g1215_p
  (
    .dout(g1215_p),
    .din1(ffc_213_p),
    .din2(ffc_444_n_spl_001)
  );


  andX
  g_g1216_p
  (
    .dout(g1216_p),
    .din1(ffc_231_p),
    .din2(ffc_444_p_spl_001)
  );


  orX
  g_g1217_n
  (
    .dout(g1217_n),
    .din1(g1215_p),
    .din2(g1216_p)
  );


  andX
  g_g1218_p
  (
    .dout(g1218_p),
    .din1(ffc_217_p),
    .din2(ffc_444_n_spl_010)
  );


  andX
  g_g1219_p
  (
    .dout(g1219_p),
    .din1(ffc_235_p),
    .din2(ffc_444_p_spl_010)
  );


  orX
  g_g1220_n
  (
    .dout(g1220_n),
    .din1(g1218_p),
    .din2(g1219_p)
  );


  andX
  g_g1221_p
  (
    .dout(g1221_p),
    .din1(ffc_219_p),
    .din2(ffc_444_n_spl_010)
  );


  andX
  g_g1222_p
  (
    .dout(g1222_p),
    .din1(ffc_237_p),
    .din2(ffc_444_p_spl_010)
  );


  orX
  g_g1223_n
  (
    .dout(g1223_n),
    .din1(g1221_p),
    .din2(g1222_p)
  );


  andX
  g_g1224_p
  (
    .dout(g1224_p),
    .din1(ffc_197_p),
    .din2(ffc_444_n_spl_011)
  );


  andX
  g_g1225_p
  (
    .dout(g1225_p),
    .din1(ffc_251_p),
    .din2(ffc_444_p_spl_011)
  );


  orX
  g_g1226_n
  (
    .dout(g1226_n),
    .din1(g1224_p),
    .din2(g1225_p)
  );


  andX
  g_g1227_p
  (
    .dout(g1227_p),
    .din1(ffc_504_p_spl_0),
    .din2(g1226_n)
  );


  andX
  g_g1228_p
  (
    .dout(g1228_p),
    .din1(ffc_215_p),
    .din2(ffc_444_n_spl_011)
  );


  andX
  g_g1229_p
  (
    .dout(g1229_p),
    .din1(ffc_233_p),
    .din2(ffc_444_p_spl_011)
  );


  orX
  g_g1230_n
  (
    .dout(g1230_n),
    .din1(g1228_p),
    .din2(g1229_p)
  );


  andX
  g_g1231_p
  (
    .dout(g1231_p),
    .din1(ffc_504_n_spl_0),
    .din2(g1230_n)
  );


  orX
  g_g1232_n
  (
    .dout(g1232_n),
    .din1(g1227_p),
    .din2(g1231_p)
  );


  andX
  g_g1233_p
  (
    .dout(g1233_p),
    .din1(ffc_187_p),
    .din2(ffc_444_n_spl_10)
  );


  andX
  g_g1234_p
  (
    .dout(g1234_p),
    .din1(ffc_241_p),
    .din2(ffc_444_p_spl_100)
  );


  orX
  g_g1235_n
  (
    .dout(g1235_n),
    .din1(g1233_p),
    .din2(g1234_p)
  );


  andX
  g_g1236_p
  (
    .dout(g1236_p),
    .din1(ffc_504_p_spl_0),
    .din2(g1235_n)
  );


  andX
  g_g1237_p
  (
    .dout(g1237_p),
    .din1(ffc_205_p),
    .din2(ffc_444_n_spl_10)
  );


  andX
  g_g1238_p
  (
    .dout(g1238_p),
    .din1(ffc_223_p),
    .din2(ffc_444_p_spl_100)
  );


  orX
  g_g1239_n
  (
    .dout(g1239_n),
    .din1(g1237_p),
    .din2(g1238_p)
  );


  andX
  g_g1240_p
  (
    .dout(g1240_p),
    .din1(ffc_504_n_spl_0),
    .din2(g1239_n)
  );


  orX
  g_g1241_n
  (
    .dout(g1241_n),
    .din1(g1236_p),
    .din2(g1240_p)
  );


  andX
  g_g1242_p
  (
    .dout(g1242_p),
    .din1(ffc_203_p),
    .din2(ffc_444_n_spl_11)
  );


  andX
  g_g1243_p
  (
    .dout(g1243_p),
    .din1(ffc_257_p),
    .din2(ffc_444_p_spl_10)
  );


  orX
  g_g1244_n
  (
    .dout(g1244_n),
    .din1(g1242_p),
    .din2(g1243_p)
  );


  andX
  g_g1245_p
  (
    .dout(g1245_p),
    .din1(ffc_504_p_spl_1),
    .din2(g1244_n)
  );


  andX
  g_g1246_p
  (
    .dout(g1246_p),
    .din1(ffc_221_p),
    .din2(ffc_444_n_spl_11)
  );


  andX
  g_g1247_p
  (
    .dout(g1247_p),
    .din1(ffc_239_p),
    .din2(ffc_444_p_spl_11)
  );


  orX
  g_g1248_n
  (
    .dout(g1248_n),
    .din1(g1246_p),
    .din2(g1247_p)
  );


  andX
  g_g1249_p
  (
    .dout(g1249_p),
    .din1(ffc_504_n_spl_),
    .din2(g1248_n)
  );


  orX
  g_g1250_n
  (
    .dout(g1250_n),
    .din1(g1245_p),
    .din2(g1249_p)
  );


  andX
  g_g1251_p
  (
    .dout(g1251_p),
    .din1(ffc_110_n),
    .din2(ffc_532_n_spl_101)
  );


  andX
  g_g1252_p
  (
    .dout(g1252_p),
    .din1(ffc_533_p_spl_10),
    .din2(g1251_p)
  );


  andX
  g_g1253_p
  (
    .dout(g1253_p),
    .din1(ffc_174_n),
    .din2(ffc_532_p_spl_10)
  );


  orX
  g_g1254_n
  (
    .dout(g1254_n),
    .din1(g1252_p),
    .din2(g1253_p)
  );


  andX
  g_g1255_p
  (
    .dout(g1255_p),
    .din1(ffc_178_p),
    .din2(ffc_532_p_spl_11)
  );


  andX
  g_g1256_p
  (
    .dout(g1256_p),
    .din1(ffc_113_p),
    .din2(ffc_532_n_spl_110)
  );


  orX
  g_g1257_n
  (
    .dout(g1257_n),
    .din1(g1255_p),
    .din2(g1256_p)
  );


  andX
  g_g1258_p
  (
    .dout(g1258_p),
    .din1(ffc_533_p_spl_11),
    .din2(g1257_n)
  );


  andX
  g_g1259_p
  (
    .dout(g1259_p),
    .din1(ffc_134_p),
    .din2(ffc_563_p_spl_0)
  );


  andX
  g_g1260_p
  (
    .dout(g1260_p),
    .din1(ffc_156_p),
    .din2(ffc_532_n_spl_110)
  );


  andX
  g_g1261_p
  (
    .dout(g1261_p),
    .din1(ffc_533_n_spl_1),
    .din2(g1260_p)
  );


  orX
  g_g1262_n
  (
    .dout(g1262_n),
    .din1(g1259_p),
    .din2(g1261_p)
  );


  orX
  g_g1263_n
  (
    .dout(g1263_n),
    .din1(g1258_p),
    .din2(g1262_n)
  );


  andX
  g_g1264_p
  (
    .dout(g1264_p),
    .din1(ffc_137_p),
    .din2(ffc_563_p_spl_1)
  );


  andX
  g_g1265_p
  (
    .dout(g1265_p),
    .din1(ffc_159_p),
    .din2(ffc_532_n_spl_11)
  );


  andX
  g_g1266_p
  (
    .dout(g1266_p),
    .din1(ffc_533_n_spl_1),
    .din2(g1265_p)
  );


  orX
  g_g1267_n
  (
    .dout(g1267_n),
    .din1(g1264_p),
    .din2(g1266_p)
  );


  andX
  g_g1268_p
  (
    .dout(g1268_p),
    .din1(g1040_n_spl_),
    .din2(g1183_n_spl_)
  );


  orX
  g_g1269_n
  (
    .dout(g1269_n),
    .din1(ffc_335_p_spl_),
    .din2(g941_n_spl_0)
  );


  orX
  g_g1270_n
  (
    .dout(g1270_n),
    .din1(ffc_299_p_spl_),
    .din2(g941_p_spl_00)
  );


  andX
  g_g1271_p
  (
    .dout(g1271_p),
    .din1(g1269_n),
    .din2(g1270_n)
  );


  orX
  g_g1272_n
  (
    .dout(g1272_n),
    .din1(ffc_338_p_spl_),
    .din2(g941_n_spl_1)
  );


  orX
  g_g1273_n
  (
    .dout(g1273_n),
    .din1(ffc_301_p_spl_),
    .din2(g941_p_spl_0)
  );


  andX
  g_g1274_p
  (
    .dout(g1274_p),
    .din1(g1272_n),
    .din2(g1273_n)
  );


  orX
  g_g1275_n
  (
    .dout(g1275_n),
    .din1(g995_n_spl_0),
    .din2(g1204_p_spl_)
  );


  andX
  g_g1276_p
  (
    .dout(g1276_p),
    .din1(ffc_325_p_spl_),
    .din2(g941_p_spl_1)
  );


  andX
  g_g1277_p
  (
    .dout(g1277_p),
    .din1(ffc_293_p_spl_),
    .din2(g941_n_spl_1)
  );


  orX
  g_g1278_n
  (
    .dout(g1278_n),
    .din1(g986_n_spl_),
    .din2(g1277_p)
  );


  orX
  g_g1279_n
  (
    .dout(g1279_n),
    .din1(g1276_p),
    .din2(g1278_n)
  );


  andX
  g_g1280_p
  (
    .dout(g1280_p),
    .din1(g1275_n),
    .din2(g1279_n)
  );


  orX
  g_g1281_n
  (
    .dout(g1281_n),
    .din1(ffc_566_n),
    .din2(ffc_574_p_spl_00)
  );


  orX
  g_g1282_n
  (
    .dout(g1282_n),
    .din1(ffc_572_n),
    .din2(ffc_574_n_spl_0)
  );


  andX
  g_g1283_p
  (
    .dout(g1283_p),
    .din1(g1281_n),
    .din2(g1282_n)
  );


  orX
  g_g1284_n
  (
    .dout(g1284_n),
    .din1(ffc_356_n_spl_),
    .din2(g1283_p)
  );


  orX
  g_g1285_n
  (
    .dout(g1285_n),
    .din1(ffc_568_n),
    .din2(ffc_574_p_spl_00)
  );


  orX
  g_g1286_n
  (
    .dout(g1286_n),
    .din1(ffc_570_n),
    .din2(ffc_574_n_spl_0)
  );


  andX
  g_g1287_p
  (
    .dout(g1287_p),
    .din1(g1285_n),
    .din2(g1286_n)
  );


  orX
  g_g1288_n
  (
    .dout(g1288_n),
    .din1(ffc_356_p_spl_0),
    .din2(g1287_p)
  );


  andX
  g_g1289_p
  (
    .dout(g1289_p),
    .din1(ffc_96_p),
    .din2(ffc_266_n_spl_)
  );


  andX
  g_g1290_p
  (
    .dout(g1290_p),
    .din1(ffc_138_p),
    .din2(ffc_266_n_spl_)
  );


  andX
  g_g1291_p
  (
    .dout(g1291_p),
    .din1(ffc_160_p),
    .din2(ffc_266_p_spl_0)
  );


  andX
  g_g1292_p
  (
    .dout(g1292_p),
    .din1(ffc_266_p_spl_0),
    .din2(ffc_275_n)
  );


  andX
  g_g1293_p
  (
    .dout(g1293_p),
    .din1(g1284_n_spl_),
    .din2(g1288_n_spl_)
  );


  andX
  g_g1294_p
  (
    .dout(g1294_p),
    .din1(ffc_567_p),
    .din2(ffc_574_n_spl_1)
  );


  andX
  g_g1295_p
  (
    .dout(g1295_p),
    .din1(ffc_573_p),
    .din2(ffc_574_p_spl_0)
  );


  orX
  g_g1296_n
  (
    .dout(g1296_n),
    .din1(g1294_p),
    .din2(g1295_p)
  );


  andX
  g_g1297_p
  (
    .dout(g1297_p),
    .din1(ffc_356_p_spl_0),
    .din2(g1296_n)
  );


  andX
  g_g1298_p
  (
    .dout(g1298_p),
    .din1(ffc_569_p),
    .din2(ffc_574_n_spl_1)
  );


  andX
  g_g1299_p
  (
    .dout(g1299_p),
    .din1(ffc_571_p),
    .din2(ffc_574_p_spl_1)
  );


  orX
  g_g1300_n
  (
    .dout(g1300_n),
    .din1(g1298_p),
    .din2(g1299_p)
  );


  andX
  g_g1301_p
  (
    .dout(g1301_p),
    .din1(ffc_356_n_spl_),
    .din2(g1300_n)
  );


  orX
  g_g1302_n
  (
    .dout(g1302_n),
    .din1(g1297_p),
    .din2(g1301_p)
  );


  buf

  (
    G2531_p,
    ffc_261_n_spl_0
  );


  buf

  (
    G2532_p,
    ffc_261_n_spl_1
  );


  buf

  (
    G2533_p,
    ffc_261_n_spl_1
  );


  buf

  (
    G2534_p,
    ffc_291_n_spl_
  );


  buf

  (
    G2535_p,
    ffc_291_n_spl_
  );


  buf

  (
    G2536_p,
    ffc_330_n_spl_0
  );


  buf

  (
    G2537_p,
    ffc_330_n_spl_0
  );


  buf

  (
    G2538_p,
    ffc_330_n_spl_
  );


  buf

  (
    G2539_p,
    ffc_100_n
  );


  buf

  (
    G2540_p,
    ffc_245_n
  );


  buf

  (
    G2541_p,
    ffc_164_n
  );


  buf

  (
    G2542_p,
    ffc_191_n
  );


  buf

  (
    G2543_p,
    ffc_142_n
  );


  buf

  (
    G2544_p,
    ffc_227_n
  );


  buf

  (
    G2545_p,
    ffc_121_n
  );


  buf

  (
    G2546_p,
    ffc_209_n
  );


  buf

  (
    G2547_p,
    g733_n
  );


  buf

  (
    G2548_p,
    g735_n
  );


  buf

  (
    G2549_p,
    ffc_261_p
  );


  buf

  (
    G2550_p,
    g736_p
  );


  buf

  (
    G2551_p,
    g737_n_spl_
  );


  buf

  (
    G2552_p,
    g738_n
  );


  buf

  (
    G2553_p,
    g739_n
  );


  buf

  (
    G2554_p,
    g742_n_spl_
  );


  buf

  (
    G2555_p,
    g742_n_spl_
  );


  buf

  (
    G2556_p,
    g745_n_spl_
  );


  buf

  (
    G2557_p,
    g746_p
  );


  buf

  (
    G2558_p,
    g747_p
  );


  buf

  (
    G2559_p,
    ffc_389_n
  );


  buf

  (
    G2560_p,
    g748_p
  );


  buf

  (
    G2561_n,
    g749_n_spl_
  );


  buf

  (
    G2562_p,
    ffc_407_n
  );


  buf

  (
    G2563_p,
    g750_n
  );


  buf

  (
    G2564_p,
    g753_n
  );


  buf

  (
    G2565_p,
    g755_n
  );


  buf

  (
    G2566_p,
    ffc_393_p
  );


  buf

  (
    G2567_p,
    ffc_392_p_spl_
  );


  buf

  (
    G2568_p,
    ffc_402_p
  );


  buf

  (
    G2569_p,
    ffc_408_p
  );


  buf

  (
    G2570_p,
    ffc_409_p
  );


  buf

  (
    G2571_p,
    ffc_410_p
  );


  buf

  (
    G2572_p,
    ffc_411_p
  );


  buf

  (
    G2573_p,
    g758_p_spl_
  );


  buf

  (
    G2574_p,
    g758_p_spl_
  );


  buf

  (
    G2575_n,
    g761_n_spl_
  );


  buf

  (
    G2576_n,
    g761_n_spl_
  );


  buf

  (
    G2577_p,
    g763_n
  );


  buf

  (
    G2578_p,
    g766_p_spl_
  );


  buf

  (
    G2579_p,
    g766_p_spl_
  );


  buf

  (
    G2580_p,
    g770_n
  );


  buf

  (
    G2581_n,
    g774_p_spl_
  );


  buf

  (
    G2582_p,
    g779_p_spl_
  );


  buf

  (
    G2583_p,
    g788_p_spl_
  );


  buf

  (
    G2584_p,
    g838_n_spl_
  );


  buf

  (
    G2585_p,
    g838_n_spl_
  );


  buf

  (
    G2586_p,
    g845_n
  );


  buf

  (
    G2587_n,
    g849_p_spl_
  );


  buf

  (
    G2588_p,
    g859_p_spl_
  );


  buf

  (
    G2589_p,
    g859_p_spl_
  );


  buf

  (
    G2590_n,
    g864_p_spl_
  );


  buf

  (
    G2591_p,
    g890_p
  );


  buf

  (
    G2592_p,
    1'b0
  );


  buf

  (
    G2593_p,
    g895_n_spl_
  );


  buf

  (
    G2594_p,
    g895_n_spl_
  );


  DROC
  ffc_0
  (
    .doutp(ffc_0_p),
    .doutn(ffc_0_n),
    .din(G1_p)
  );


  DROC
  ffc_1
  (
    .doutp(ffc_1_p),
    .doutn(ffc_1_n),
    .din(ffc_0_p)
  );


  DROC
  ffc_2
  (
    .doutp(ffc_2_p),
    .doutn(ffc_2_n),
    .din(ffc_1_p)
  );


  DROC
  ffc_3
  (
    .doutp(ffc_3_p),
    .doutn(ffc_3_n),
    .din(ffc_2_p)
  );


  DROC
  ffc_4
  (
    .doutp(ffc_4_p),
    .doutn(ffc_4_n),
    .din(G2_p)
  );


  DROC
  ffc_5
  (
    .doutp(ffc_5_p),
    .doutn(ffc_5_n),
    .din(ffc_4_p)
  );


  DROC
  ffc_6
  (
    .doutp(ffc_6_p),
    .doutn(ffc_6_n),
    .din(ffc_5_p)
  );


  DROC
  ffc_7
  (
    .doutp(ffc_7_p),
    .doutn(ffc_7_n),
    .din(ffc_6_p)
  );


  DROC
  ffc_8
  (
    .doutp(ffc_8_p),
    .doutn(ffc_8_n),
    .din(G3_p)
  );


  DROC
  ffc_9
  (
    .doutp(ffc_9_p),
    .doutn(ffc_9_n),
    .din(ffc_8_p)
  );


  DROC
  ffc_10
  (
    .doutp(ffc_10_p),
    .doutn(ffc_10_n),
    .din(ffc_9_p)
  );


  DROC
  ffc_11
  (
    .doutp(ffc_11_p),
    .doutn(ffc_11_n),
    .din(ffc_10_p)
  );


  DROC
  ffc_12
  (
    .doutp(ffc_12_p),
    .doutn(ffc_12_n),
    .din(G4_p)
  );


  DROC
  ffc_13
  (
    .doutp(ffc_13_p),
    .doutn(ffc_13_n),
    .din(ffc_12_p)
  );


  DROC
  ffc_14
  (
    .doutp(ffc_14_p),
    .doutn(ffc_14_n),
    .din(ffc_13_p)
  );


  DROC
  ffc_15
  (
    .doutp(ffc_15_p),
    .doutn(ffc_15_n),
    .din(G5_p)
  );


  DROC
  ffc_16
  (
    .doutp(ffc_16_p),
    .doutn(ffc_16_n),
    .din(ffc_15_p)
  );


  DROC
  ffc_17
  (
    .doutp(ffc_17_p),
    .doutn(ffc_17_n),
    .din(ffc_16_p)
  );


  DROC
  ffc_18
  (
    .doutp(ffc_18_p),
    .doutn(ffc_18_n),
    .din(G6_p)
  );


  DROC
  ffc_19
  (
    .doutp(ffc_19_p),
    .doutn(ffc_19_n),
    .din(ffc_18_p)
  );


  DROC
  ffc_20
  (
    .doutp(ffc_20_p),
    .doutn(ffc_20_n),
    .din(ffc_19_p)
  );


  DROC
  ffc_21
  (
    .doutp(ffc_21_p),
    .doutn(ffc_21_n),
    .din(G7_p)
  );


  DROC
  ffc_22
  (
    .doutp(ffc_22_p),
    .doutn(ffc_22_n),
    .din(ffc_21_p)
  );


  DROC
  ffc_23
  (
    .doutp(ffc_23_p),
    .doutn(ffc_23_n),
    .din(ffc_22_p)
  );


  DROC
  ffc_24
  (
    .doutp(ffc_24_p),
    .doutn(ffc_24_n),
    .din(ffc_23_p)
  );


  DROC
  ffc_25
  (
    .doutp(ffc_25_p),
    .doutn(ffc_25_n),
    .din(G8_p)
  );


  DROC
  ffc_26
  (
    .doutp(ffc_26_p),
    .doutn(ffc_26_n),
    .din(ffc_25_p)
  );


  DROC
  ffc_27
  (
    .doutp(ffc_27_p),
    .doutn(ffc_27_n),
    .din(G9_p)
  );


  DROC
  ffc_28
  (
    .doutp(ffc_28_p),
    .doutn(ffc_28_n),
    .din(ffc_27_p)
  );


  DROC
  ffc_29
  (
    .doutp(ffc_29_p),
    .doutn(ffc_29_n),
    .din(ffc_28_p)
  );


  DROC
  ffc_30
  (
    .doutp(ffc_30_p),
    .doutn(ffc_30_n),
    .din(ffc_29_p)
  );


  DROC
  ffc_31
  (
    .doutp(ffc_31_p),
    .doutn(ffc_31_n),
    .din(G10_p)
  );


  DROC
  ffc_32
  (
    .doutp(ffc_32_p),
    .doutn(ffc_32_n),
    .din(ffc_31_p)
  );


  DROC
  ffc_33
  (
    .doutp(ffc_33_p),
    .doutn(ffc_33_n),
    .din(ffc_32_p)
  );


  DROC
  ffc_34
  (
    .doutp(ffc_34_p),
    .doutn(ffc_34_n),
    .din(ffc_33_p)
  );


  DROC
  ffc_35
  (
    .doutp(ffc_35_p),
    .doutn(ffc_35_n),
    .din(G11_p)
  );


  DROC
  ffc_36
  (
    .doutp(ffc_36_p),
    .doutn(ffc_36_n),
    .din(ffc_35_p)
  );


  DROC
  ffc_37
  (
    .doutp(ffc_37_p),
    .doutn(ffc_37_n),
    .din(ffc_36_p)
  );


  DROC
  ffc_38
  (
    .doutp(ffc_38_p),
    .doutn(ffc_38_n),
    .din(ffc_37_p)
  );


  DROC
  ffc_39
  (
    .doutp(ffc_39_p),
    .doutn(ffc_39_n),
    .din(G12_p)
  );


  DROC
  ffc_40
  (
    .doutp(ffc_40_p),
    .doutn(ffc_40_n),
    .din(ffc_39_p)
  );


  DROC
  ffc_41
  (
    .doutp(ffc_41_p),
    .doutn(ffc_41_n),
    .din(ffc_40_p)
  );


  DROC
  ffc_42
  (
    .doutp(ffc_42_p),
    .doutn(ffc_42_n),
    .din(G13_p)
  );


  DROC
  ffc_43
  (
    .doutp(ffc_43_p),
    .doutn(ffc_43_n),
    .din(ffc_42_p)
  );


  DROC
  ffc_44
  (
    .doutp(ffc_44_p),
    .doutn(ffc_44_n),
    .din(ffc_43_p)
  );


  DROC
  ffc_45
  (
    .doutp(ffc_45_p),
    .doutn(ffc_45_n),
    .din(G14_p)
  );


  DROC
  ffc_46
  (
    .doutp(ffc_46_p),
    .doutn(ffc_46_n),
    .din(ffc_45_p)
  );


  DROC
  ffc_47
  (
    .doutp(ffc_47_p),
    .doutn(ffc_47_n),
    .din(ffc_46_p)
  );


  DROC
  ffc_48
  (
    .doutp(ffc_48_p),
    .doutn(ffc_48_n),
    .din(G15_p)
  );


  DROC
  ffc_49
  (
    .doutp(ffc_49_p),
    .doutn(ffc_49_n),
    .din(ffc_48_p)
  );


  DROC
  ffc_50
  (
    .doutp(ffc_50_p),
    .doutn(ffc_50_n),
    .din(ffc_49_p)
  );


  DROC
  ffc_51
  (
    .doutp(ffc_51_p),
    .doutn(ffc_51_n),
    .din(G16_p)
  );


  DROC
  ffc_52
  (
    .doutp(ffc_52_p),
    .doutn(ffc_52_n),
    .din(ffc_51_p)
  );


  DROC
  ffc_53
  (
    .doutp(ffc_53_p),
    .doutn(ffc_53_n),
    .din(ffc_52_p)
  );


  DROC
  ffc_54
  (
    .doutp(ffc_54_p),
    .doutn(ffc_54_n),
    .din(G17_p)
  );


  DROC
  ffc_55
  (
    .doutp(ffc_55_p),
    .doutn(ffc_55_n),
    .din(ffc_54_p)
  );


  DROC
  ffc_56
  (
    .doutp(ffc_56_p),
    .doutn(ffc_56_n),
    .din(ffc_55_p)
  );


  DROC
  ffc_57
  (
    .doutp(ffc_57_p),
    .doutn(ffc_57_n),
    .din(G18_p)
  );


  DROC
  ffc_58
  (
    .doutp(ffc_58_p),
    .doutn(ffc_58_n),
    .din(ffc_57_p)
  );


  DROC
  ffc_59
  (
    .doutp(ffc_59_p),
    .doutn(ffc_59_n),
    .din(ffc_58_p)
  );


  DROC
  ffc_60
  (
    .doutp(ffc_60_p),
    .doutn(ffc_60_n),
    .din(G19_p)
  );


  DROC
  ffc_61
  (
    .doutp(ffc_61_p),
    .doutn(ffc_61_n),
    .din(ffc_60_p)
  );


  DROC
  ffc_62
  (
    .doutp(ffc_62_p),
    .doutn(ffc_62_n),
    .din(ffc_61_p)
  );


  DROC
  ffc_63
  (
    .doutp(ffc_63_p),
    .doutn(ffc_63_n),
    .din(G20_p)
  );


  DROC
  ffc_64
  (
    .doutp(ffc_64_p),
    .doutn(ffc_64_n),
    .din(ffc_63_p)
  );


  DROC
  ffc_65
  (
    .doutp(ffc_65_p),
    .doutn(ffc_65_n),
    .din(ffc_64_p)
  );


  DROC
  ffc_66
  (
    .doutp(ffc_66_p),
    .doutn(ffc_66_n),
    .din(G21_p)
  );


  DROC
  ffc_67
  (
    .doutp(ffc_67_p),
    .doutn(ffc_67_n),
    .din(ffc_66_p)
  );


  DROC
  ffc_68
  (
    .doutp(ffc_68_p),
    .doutn(ffc_68_n),
    .din(ffc_67_p)
  );


  DROC
  ffc_69
  (
    .doutp(ffc_69_p),
    .doutn(ffc_69_n),
    .din(G22_p)
  );


  DROC
  ffc_70
  (
    .doutp(ffc_70_p),
    .doutn(ffc_70_n),
    .din(ffc_69_p)
  );


  DROC
  ffc_71
  (
    .doutp(ffc_71_p),
    .doutn(ffc_71_n),
    .din(ffc_70_p)
  );


  DROC
  ffc_72
  (
    .doutp(ffc_72_p),
    .doutn(ffc_72_n),
    .din(G23_p)
  );


  DROC
  ffc_73
  (
    .doutp(ffc_73_p),
    .doutn(ffc_73_n),
    .din(ffc_72_p)
  );


  DROC
  ffc_74
  (
    .doutp(ffc_74_p),
    .doutn(ffc_74_n),
    .din(ffc_73_p)
  );


  DROC
  ffc_75
  (
    .doutp(ffc_75_p),
    .doutn(ffc_75_n),
    .din(G24_p)
  );


  DROC
  ffc_76
  (
    .doutp(ffc_76_p),
    .doutn(ffc_76_n),
    .din(ffc_75_p)
  );


  DROC
  ffc_77
  (
    .doutp(ffc_77_p),
    .doutn(ffc_77_n),
    .din(ffc_76_p)
  );


  DROC
  ffc_78
  (
    .doutp(ffc_78_p),
    .doutn(ffc_78_n),
    .din(G25_p)
  );


  DROC
  ffc_79
  (
    .doutp(ffc_79_p),
    .doutn(ffc_79_n),
    .din(ffc_78_p)
  );


  DROC
  ffc_80
  (
    .doutp(ffc_80_p),
    .doutn(ffc_80_n),
    .din(ffc_79_p)
  );


  DROC
  ffc_81
  (
    .doutp(ffc_81_p),
    .doutn(ffc_81_n),
    .din(G26_p)
  );


  DROC
  ffc_82
  (
    .doutp(ffc_82_p),
    .doutn(ffc_82_n),
    .din(ffc_81_p)
  );


  DROC
  ffc_83
  (
    .doutp(ffc_83_p),
    .doutn(ffc_83_n),
    .din(ffc_82_p)
  );


  DROC
  ffc_84
  (
    .doutp(ffc_84_p),
    .doutn(ffc_84_n),
    .din(G27_p)
  );


  DROC
  ffc_85
  (
    .doutp(ffc_85_p),
    .doutn(ffc_85_n),
    .din(ffc_84_p)
  );


  DROC
  ffc_86
  (
    .doutp(ffc_86_p),
    .doutn(ffc_86_n),
    .din(ffc_85_p)
  );


  DROC
  ffc_87
  (
    .doutp(ffc_87_p),
    .doutn(ffc_87_n),
    .din(G28_p)
  );


  DROC
  ffc_88
  (
    .doutp(ffc_88_p),
    .doutn(ffc_88_n),
    .din(ffc_87_p)
  );


  DROC
  ffc_89
  (
    .doutp(ffc_89_p),
    .doutn(ffc_89_n),
    .din(ffc_88_p)
  );


  DROC
  ffc_90
  (
    .doutp(ffc_90_p),
    .doutn(ffc_90_n),
    .din(ffc_89_p)
  );


  DROC
  ffc_91
  (
    .doutp(ffc_91_p),
    .doutn(ffc_91_n),
    .din(G29_p)
  );


  DROC
  ffc_92
  (
    .doutp(ffc_92_p),
    .doutn(ffc_92_n),
    .din(ffc_91_p)
  );


  DROC
  ffc_93
  (
    .doutp(ffc_93_p),
    .doutn(ffc_93_n),
    .din(ffc_92_p)
  );


  DROC
  ffc_94
  (
    .doutp(ffc_94_p),
    .doutn(ffc_94_n),
    .din(ffc_93_p)
  );


  DROC
  ffc_95
  (
    .doutp(ffc_95_p),
    .doutn(ffc_95_n),
    .din(G30_p)
  );


  DROC
  ffc_96
  (
    .doutp(ffc_96_p),
    .doutn(ffc_96_n),
    .din(G31_p)
  );


  DROC
  ffc_97
  (
    .doutp(ffc_97_p),
    .doutn(ffc_97_n),
    .din(G32_p)
  );


  DROC
  ffc_98
  (
    .doutp(ffc_98_p),
    .doutn(ffc_98_n),
    .din(ffc_97_p)
  );


  DROC
  ffc_99
  (
    .doutp(ffc_99_p),
    .doutn(ffc_99_n),
    .din(ffc_98_p)
  );


  DROC
  ffc_100
  (
    .doutp(ffc_100_p),
    .doutn(ffc_100_n),
    .din(ffc_99_p_spl_)
  );


  DROC
  ffc_101
  (
    .doutp(ffc_101_p),
    .doutn(ffc_101_n),
    .din(G33_p)
  );


  DROC
  ffc_102
  (
    .doutp(ffc_102_p),
    .doutn(ffc_102_n),
    .din(ffc_101_p)
  );


  DROC
  ffc_103
  (
    .doutp(ffc_103_p),
    .doutn(ffc_103_n),
    .din(G34_p)
  );


  DROC
  ffc_104
  (
    .doutp(ffc_104_p),
    .doutn(ffc_104_n),
    .din(ffc_103_p)
  );


  DROC
  ffc_105
  (
    .doutp(ffc_105_p),
    .doutn(ffc_105_n),
    .din(G35_p)
  );


  DROC
  ffc_106
  (
    .doutp(ffc_106_p),
    .doutn(ffc_106_n),
    .din(ffc_105_p)
  );


  DROC
  ffc_107
  (
    .doutp(ffc_107_p),
    .doutn(ffc_107_n),
    .din(G36_p)
  );


  DROC
  ffc_108
  (
    .doutp(ffc_108_p),
    .doutn(ffc_108_n),
    .din(ffc_107_p)
  );


  DROC
  ffc_109
  (
    .doutp(ffc_109_p),
    .doutn(ffc_109_n),
    .din(G37_p)
  );


  DROC
  ffc_110
  (
    .doutp(ffc_110_p),
    .doutn(ffc_110_n),
    .din(ffc_109_p)
  );


  DROC
  ffc_111
  (
    .doutp(ffc_111_p),
    .doutn(ffc_111_n),
    .din(G38_p)
  );


  DROC
  ffc_112
  (
    .doutp(ffc_112_p),
    .doutn(ffc_112_n),
    .din(G39_p)
  );


  DROC
  ffc_113
  (
    .doutp(ffc_113_p),
    .doutn(ffc_113_n),
    .din(ffc_112_p)
  );


  DROC
  ffc_114
  (
    .doutp(ffc_114_p),
    .doutn(ffc_114_n),
    .din(G40_p)
  );


  DROC
  ffc_115
  (
    .doutp(ffc_115_p),
    .doutn(ffc_115_n),
    .din(G41_p)
  );


  DROC
  ffc_116
  (
    .doutp(ffc_116_p),
    .doutn(ffc_116_n),
    .din(ffc_115_p)
  );


  DROC
  ffc_117
  (
    .doutp(ffc_117_p),
    .doutn(ffc_117_n),
    .din(G42_p)
  );


  DROC
  ffc_118
  (
    .doutp(ffc_118_p),
    .doutn(ffc_118_n),
    .din(G43_p)
  );


  DROC
  ffc_119
  (
    .doutp(ffc_119_p),
    .doutn(ffc_119_n),
    .din(ffc_118_p)
  );


  DROC
  ffc_120
  (
    .doutp(ffc_120_p),
    .doutn(ffc_120_n),
    .din(ffc_119_p)
  );


  DROC
  ffc_121
  (
    .doutp(ffc_121_p),
    .doutn(ffc_121_n),
    .din(ffc_120_p_spl_)
  );


  DROC
  ffc_122
  (
    .doutp(ffc_122_p),
    .doutn(ffc_122_n),
    .din(G44_p)
  );


  DROC
  ffc_123
  (
    .doutp(ffc_123_p),
    .doutn(ffc_123_n),
    .din(ffc_122_p)
  );


  DROC
  ffc_124
  (
    .doutp(ffc_124_p),
    .doutn(ffc_124_n),
    .din(G45_p)
  );


  DROC
  ffc_125
  (
    .doutp(ffc_125_p),
    .doutn(ffc_125_n),
    .din(ffc_124_p)
  );


  DROC
  ffc_126
  (
    .doutp(ffc_126_p),
    .doutn(ffc_126_n),
    .din(G46_p)
  );


  DROC
  ffc_127
  (
    .doutp(ffc_127_p),
    .doutn(ffc_127_n),
    .din(ffc_126_p)
  );


  DROC
  ffc_128
  (
    .doutp(ffc_128_p),
    .doutn(ffc_128_n),
    .din(ffc_127_p)
  );


  DROC
  ffc_129
  (
    .doutp(ffc_129_p),
    .doutn(ffc_129_n),
    .din(G47_p)
  );


  DROC
  ffc_130
  (
    .doutp(ffc_130_p),
    .doutn(ffc_130_n),
    .din(ffc_129_p)
  );


  DROC
  ffc_131
  (
    .doutp(ffc_131_p),
    .doutn(ffc_131_n),
    .din(G48_p)
  );


  DROC
  ffc_132
  (
    .doutp(ffc_132_p),
    .doutn(ffc_132_n),
    .din(ffc_131_p)
  );


  DROC
  ffc_133
  (
    .doutp(ffc_133_p),
    .doutn(ffc_133_n),
    .din(G49_p)
  );


  DROC
  ffc_134
  (
    .doutp(ffc_134_p),
    .doutn(ffc_134_n),
    .din(ffc_133_p)
  );


  DROC
  ffc_135
  (
    .doutp(ffc_135_p),
    .doutn(ffc_135_n),
    .din(G50_p)
  );


  DROC
  ffc_136
  (
    .doutp(ffc_136_p),
    .doutn(ffc_136_n),
    .din(G51_p)
  );


  DROC
  ffc_137
  (
    .doutp(ffc_137_p),
    .doutn(ffc_137_n),
    .din(ffc_136_p)
  );


  DROC
  ffc_138
  (
    .doutp(ffc_138_p),
    .doutn(ffc_138_n),
    .din(G52_p)
  );


  DROC
  ffc_139
  (
    .doutp(ffc_139_p),
    .doutn(ffc_139_n),
    .din(G53_p)
  );


  DROC
  ffc_140
  (
    .doutp(ffc_140_p),
    .doutn(ffc_140_n),
    .din(ffc_139_p)
  );


  DROC
  ffc_141
  (
    .doutp(ffc_141_p),
    .doutn(ffc_141_n),
    .din(ffc_140_p)
  );


  DROC
  ffc_142
  (
    .doutp(ffc_142_p),
    .doutn(ffc_142_n),
    .din(ffc_141_p_spl_)
  );


  DROC
  ffc_143
  (
    .doutp(ffc_143_p),
    .doutn(ffc_143_n),
    .din(G54_p)
  );


  DROC
  ffc_144
  (
    .doutp(ffc_144_p),
    .doutn(ffc_144_n),
    .din(ffc_143_p)
  );


  DROC
  ffc_145
  (
    .doutp(ffc_145_p),
    .doutn(ffc_145_n),
    .din(G55_p)
  );


  DROC
  ffc_146
  (
    .doutp(ffc_146_p),
    .doutn(ffc_146_n),
    .din(ffc_145_p)
  );


  DROC
  ffc_147
  (
    .doutp(ffc_147_p),
    .doutn(ffc_147_n),
    .din(G56_p)
  );


  DROC
  ffc_148
  (
    .doutp(ffc_148_p),
    .doutn(ffc_148_n),
    .din(ffc_147_p)
  );


  DROC
  ffc_149
  (
    .doutp(ffc_149_p),
    .doutn(ffc_149_n),
    .din(G57_p)
  );


  DROC
  ffc_150
  (
    .doutp(ffc_150_p),
    .doutn(ffc_150_n),
    .din(ffc_149_p)
  );


  DROC
  ffc_151
  (
    .doutp(ffc_151_p),
    .doutn(ffc_151_n),
    .din(G58_p)
  );


  DROC
  ffc_152
  (
    .doutp(ffc_152_p),
    .doutn(ffc_152_n),
    .din(ffc_151_p)
  );


  DROC
  ffc_153
  (
    .doutp(ffc_153_p),
    .doutn(ffc_153_n),
    .din(G59_p)
  );


  DROC
  ffc_154
  (
    .doutp(ffc_154_p),
    .doutn(ffc_154_n),
    .din(ffc_153_p)
  );


  DROC
  ffc_155
  (
    .doutp(ffc_155_p),
    .doutn(ffc_155_n),
    .din(G60_p)
  );


  DROC
  ffc_156
  (
    .doutp(ffc_156_p),
    .doutn(ffc_156_n),
    .din(ffc_155_p)
  );


  DROC
  ffc_157
  (
    .doutp(ffc_157_p),
    .doutn(ffc_157_n),
    .din(G61_p)
  );


  DROC
  ffc_158
  (
    .doutp(ffc_158_p),
    .doutn(ffc_158_n),
    .din(G62_p)
  );


  DROC
  ffc_159
  (
    .doutp(ffc_159_p),
    .doutn(ffc_159_n),
    .din(ffc_158_p)
  );


  DROC
  ffc_160
  (
    .doutp(ffc_160_p),
    .doutn(ffc_160_n),
    .din(G63_p)
  );


  DROC
  ffc_161
  (
    .doutp(ffc_161_p),
    .doutn(ffc_161_n),
    .din(G64_p)
  );


  DROC
  ffc_162
  (
    .doutp(ffc_162_p),
    .doutn(ffc_162_n),
    .din(ffc_161_p)
  );


  DROC
  ffc_163
  (
    .doutp(ffc_163_p),
    .doutn(ffc_163_n),
    .din(ffc_162_p)
  );


  DROC
  ffc_164
  (
    .doutp(ffc_164_p),
    .doutn(ffc_164_n),
    .din(ffc_163_p_spl_)
  );


  DROC
  ffc_165
  (
    .doutp(ffc_165_p),
    .doutn(ffc_165_n),
    .din(G65_p)
  );


  DROC
  ffc_166
  (
    .doutp(ffc_166_p),
    .doutn(ffc_166_n),
    .din(ffc_165_p)
  );


  DROC
  ffc_167
  (
    .doutp(ffc_167_p),
    .doutn(ffc_167_n),
    .din(G66_p)
  );


  DROC
  ffc_168
  (
    .doutp(ffc_168_p),
    .doutn(ffc_168_n),
    .din(ffc_167_p)
  );


  DROC
  ffc_169
  (
    .doutp(ffc_169_p),
    .doutn(ffc_169_n),
    .din(G67_p)
  );


  DROC
  ffc_170
  (
    .doutp(ffc_170_p),
    .doutn(ffc_170_n),
    .din(ffc_169_p)
  );


  DROC
  ffc_171
  (
    .doutp(ffc_171_p),
    .doutn(ffc_171_n),
    .din(G68_p)
  );


  DROC
  ffc_172
  (
    .doutp(ffc_172_p),
    .doutn(ffc_172_n),
    .din(ffc_171_p)
  );


  DROC
  ffc_173
  (
    .doutp(ffc_173_p),
    .doutn(ffc_173_n),
    .din(G69_p)
  );


  DROC
  ffc_174
  (
    .doutp(ffc_174_p),
    .doutn(ffc_174_n),
    .din(ffc_173_p)
  );


  DROC
  ffc_175
  (
    .doutp(ffc_175_p),
    .doutn(ffc_175_n),
    .din(G70_p)
  );


  DROC
  ffc_176
  (
    .doutp(ffc_176_p),
    .doutn(ffc_176_n),
    .din(ffc_175_p)
  );


  DROC
  ffc_177
  (
    .doutp(ffc_177_p),
    .doutn(ffc_177_n),
    .din(G71_p)
  );


  DROC
  ffc_178
  (
    .doutp(ffc_178_p),
    .doutn(ffc_178_n),
    .din(ffc_177_p)
  );


  DROC
  ffc_179
  (
    .doutp(ffc_179_p),
    .doutn(ffc_179_n),
    .din(G72_p)
  );


  DROC
  ffc_180
  (
    .doutp(ffc_180_p),
    .doutn(ffc_180_n),
    .din(G73_p)
  );


  DROC
  ffc_181
  (
    .doutp(ffc_181_p),
    .doutn(ffc_181_n),
    .din(ffc_180_p)
  );


  DROC
  ffc_182
  (
    .doutp(ffc_182_p),
    .doutn(ffc_182_n),
    .din(G74_p)
  );


  DROC
  ffc_183
  (
    .doutp(ffc_183_p),
    .doutn(ffc_183_n),
    .din(ffc_182_p)
  );


  DROC
  ffc_184
  (
    .doutp(ffc_184_p),
    .doutn(ffc_184_n),
    .din(ffc_183_p)
  );


  DROC
  ffc_185
  (
    .doutp(ffc_185_p),
    .doutn(ffc_185_n),
    .din(ffc_184_p)
  );


  DROC
  ffc_186
  (
    .doutp(ffc_186_p),
    .doutn(ffc_186_n),
    .din(G75_p)
  );


  DROC
  ffc_187
  (
    .doutp(ffc_187_p),
    .doutn(ffc_187_n),
    .din(ffc_186_p)
  );


  DROC
  ffc_188
  (
    .doutp(ffc_188_p),
    .doutn(ffc_188_n),
    .din(G76_p)
  );


  DROC
  ffc_189
  (
    .doutp(ffc_189_p),
    .doutn(ffc_189_n),
    .din(ffc_188_p)
  );


  DROC
  ffc_190
  (
    .doutp(ffc_190_p),
    .doutn(ffc_190_n),
    .din(ffc_189_p)
  );


  DROC
  ffc_191
  (
    .doutp(ffc_191_p),
    .doutn(ffc_191_n),
    .din(ffc_190_p_spl_)
  );


  DROC
  ffc_192
  (
    .doutp(ffc_192_p),
    .doutn(ffc_192_n),
    .din(G77_p)
  );


  DROC
  ffc_193
  (
    .doutp(ffc_193_p),
    .doutn(ffc_193_n),
    .din(ffc_192_p)
  );


  DROC
  ffc_194
  (
    .doutp(ffc_194_p),
    .doutn(ffc_194_n),
    .din(G78_p)
  );


  DROC
  ffc_195
  (
    .doutp(ffc_195_p),
    .doutn(ffc_195_n),
    .din(ffc_194_p)
  );


  DROC
  ffc_196
  (
    .doutp(ffc_196_p),
    .doutn(ffc_196_n),
    .din(G81_p)
  );


  DROC
  ffc_197
  (
    .doutp(ffc_197_p),
    .doutn(ffc_197_n),
    .din(ffc_196_p)
  );


  DROC
  ffc_198
  (
    .doutp(ffc_198_p),
    .doutn(ffc_198_n),
    .din(G82_p)
  );


  DROC
  ffc_199
  (
    .doutp(ffc_199_p),
    .doutn(ffc_199_n),
    .din(ffc_198_p)
  );


  DROC
  ffc_200
  (
    .doutp(ffc_200_p),
    .doutn(ffc_200_n),
    .din(G83_p)
  );


  DROC
  ffc_201
  (
    .doutp(ffc_201_p),
    .doutn(ffc_201_n),
    .din(ffc_200_p)
  );


  DROC
  ffc_202
  (
    .doutp(ffc_202_p),
    .doutn(ffc_202_n),
    .din(G84_p)
  );


  DROC
  ffc_203
  (
    .doutp(ffc_203_p),
    .doutn(ffc_203_n),
    .din(ffc_202_p)
  );


  DROC
  ffc_204
  (
    .doutp(ffc_204_p),
    .doutn(ffc_204_n),
    .din(G85_p)
  );


  DROC
  ffc_205
  (
    .doutp(ffc_205_p),
    .doutn(ffc_205_n),
    .din(ffc_204_p)
  );


  DROC
  ffc_206
  (
    .doutp(ffc_206_p),
    .doutn(ffc_206_n),
    .din(G86_p)
  );


  DROC
  ffc_207
  (
    .doutp(ffc_207_p),
    .doutn(ffc_207_n),
    .din(ffc_206_p)
  );


  DROC
  ffc_208
  (
    .doutp(ffc_208_p),
    .doutn(ffc_208_n),
    .din(ffc_207_p)
  );


  DROC
  ffc_209
  (
    .doutp(ffc_209_p),
    .doutn(ffc_209_n),
    .din(ffc_208_p_spl_)
  );


  DROC
  ffc_210
  (
    .doutp(ffc_210_p),
    .doutn(ffc_210_n),
    .din(G87_p)
  );


  DROC
  ffc_211
  (
    .doutp(ffc_211_p),
    .doutn(ffc_211_n),
    .din(ffc_210_p)
  );


  DROC
  ffc_212
  (
    .doutp(ffc_212_p),
    .doutn(ffc_212_n),
    .din(G88_p)
  );


  DROC
  ffc_213
  (
    .doutp(ffc_213_p),
    .doutn(ffc_213_n),
    .din(ffc_212_p)
  );


  DROC
  ffc_214
  (
    .doutp(ffc_214_p),
    .doutn(ffc_214_n),
    .din(G91_p)
  );


  DROC
  ffc_215
  (
    .doutp(ffc_215_p),
    .doutn(ffc_215_n),
    .din(ffc_214_p)
  );


  DROC
  ffc_216
  (
    .doutp(ffc_216_p),
    .doutn(ffc_216_n),
    .din(G92_p)
  );


  DROC
  ffc_217
  (
    .doutp(ffc_217_p),
    .doutn(ffc_217_n),
    .din(ffc_216_p)
  );


  DROC
  ffc_218
  (
    .doutp(ffc_218_p),
    .doutn(ffc_218_n),
    .din(G93_p)
  );


  DROC
  ffc_219
  (
    .doutp(ffc_219_p),
    .doutn(ffc_219_n),
    .din(ffc_218_p)
  );


  DROC
  ffc_220
  (
    .doutp(ffc_220_p),
    .doutn(ffc_220_n),
    .din(G94_p)
  );


  DROC
  ffc_221
  (
    .doutp(ffc_221_p),
    .doutn(ffc_221_n),
    .din(ffc_220_p)
  );


  DROC
  ffc_222
  (
    .doutp(ffc_222_p),
    .doutn(ffc_222_n),
    .din(G95_p)
  );


  DROC
  ffc_223
  (
    .doutp(ffc_223_p),
    .doutn(ffc_223_n),
    .din(ffc_222_p)
  );


  DROC
  ffc_224
  (
    .doutp(ffc_224_p),
    .doutn(ffc_224_n),
    .din(G96_p)
  );


  DROC
  ffc_225
  (
    .doutp(ffc_225_p),
    .doutn(ffc_225_n),
    .din(ffc_224_p)
  );


  DROC
  ffc_226
  (
    .doutp(ffc_226_p),
    .doutn(ffc_226_n),
    .din(ffc_225_p)
  );


  DROC
  ffc_227
  (
    .doutp(ffc_227_p),
    .doutn(ffc_227_n),
    .din(ffc_226_p_spl_)
  );


  DROC
  ffc_228
  (
    .doutp(ffc_228_p),
    .doutn(ffc_228_n),
    .din(G97_p)
  );


  DROC
  ffc_229
  (
    .doutp(ffc_229_p),
    .doutn(ffc_229_n),
    .din(ffc_228_p)
  );


  DROC
  ffc_230
  (
    .doutp(ffc_230_p),
    .doutn(ffc_230_n),
    .din(G98_p)
  );


  DROC
  ffc_231
  (
    .doutp(ffc_231_p),
    .doutn(ffc_231_n),
    .din(ffc_230_p)
  );


  DROC
  ffc_232
  (
    .doutp(ffc_232_p),
    .doutn(ffc_232_n),
    .din(G101_p)
  );


  DROC
  ffc_233
  (
    .doutp(ffc_233_p),
    .doutn(ffc_233_n),
    .din(ffc_232_p)
  );


  DROC
  ffc_234
  (
    .doutp(ffc_234_p),
    .doutn(ffc_234_n),
    .din(G102_p)
  );


  DROC
  ffc_235
  (
    .doutp(ffc_235_p),
    .doutn(ffc_235_n),
    .din(ffc_234_p)
  );


  DROC
  ffc_236
  (
    .doutp(ffc_236_p),
    .doutn(ffc_236_n),
    .din(G103_p)
  );


  DROC
  ffc_237
  (
    .doutp(ffc_237_p),
    .doutn(ffc_237_n),
    .din(ffc_236_p)
  );


  DROC
  ffc_238
  (
    .doutp(ffc_238_p),
    .doutn(ffc_238_n),
    .din(G104_p)
  );


  DROC
  ffc_239
  (
    .doutp(ffc_239_p),
    .doutn(ffc_239_n),
    .din(ffc_238_p)
  );


  DROC
  ffc_240
  (
    .doutp(ffc_240_p),
    .doutn(ffc_240_n),
    .din(G105_p)
  );


  DROC
  ffc_241
  (
    .doutp(ffc_241_p),
    .doutn(ffc_241_n),
    .din(ffc_240_p)
  );


  DROC
  ffc_242
  (
    .doutp(ffc_242_p),
    .doutn(ffc_242_n),
    .din(G106_p)
  );


  DROC
  ffc_243
  (
    .doutp(ffc_243_p),
    .doutn(ffc_243_n),
    .din(ffc_242_p)
  );


  DROC
  ffc_244
  (
    .doutp(ffc_244_p),
    .doutn(ffc_244_n),
    .din(ffc_243_p)
  );


  DROC
  ffc_245
  (
    .doutp(ffc_245_p),
    .doutn(ffc_245_n),
    .din(ffc_244_p_spl_)
  );


  DROC
  ffc_246
  (
    .doutp(ffc_246_p),
    .doutn(ffc_246_n),
    .din(G107_p)
  );


  DROC
  ffc_247
  (
    .doutp(ffc_247_p),
    .doutn(ffc_247_n),
    .din(ffc_246_p)
  );


  DROC
  ffc_248
  (
    .doutp(ffc_248_p),
    .doutn(ffc_248_n),
    .din(G108_p)
  );


  DROC
  ffc_249
  (
    .doutp(ffc_249_p),
    .doutn(ffc_249_n),
    .din(ffc_248_p)
  );


  DROC
  ffc_250
  (
    .doutp(ffc_250_p),
    .doutn(ffc_250_n),
    .din(G111_p)
  );


  DROC
  ffc_251
  (
    .doutp(ffc_251_p),
    .doutn(ffc_251_n),
    .din(ffc_250_p)
  );


  DROC
  ffc_252
  (
    .doutp(ffc_252_p),
    .doutn(ffc_252_n),
    .din(G112_p)
  );


  DROC
  ffc_253
  (
    .doutp(ffc_253_p),
    .doutn(ffc_253_n),
    .din(ffc_252_p)
  );


  DROC
  ffc_254
  (
    .doutp(ffc_254_p),
    .doutn(ffc_254_n),
    .din(G113_p)
  );


  DROC
  ffc_255
  (
    .doutp(ffc_255_p),
    .doutn(ffc_255_n),
    .din(ffc_254_p)
  );


  DROC
  ffc_256
  (
    .doutp(ffc_256_p),
    .doutn(ffc_256_n),
    .din(G114_p)
  );


  DROC
  ffc_257
  (
    .doutp(ffc_257_p),
    .doutn(ffc_257_n),
    .din(ffc_256_p)
  );


  DROC
  ffc_258
  (
    .doutp(ffc_258_p),
    .doutn(ffc_258_n),
    .din(G115_p)
  );


  DROC
  ffc_259
  (
    .doutp(ffc_259_p),
    .doutn(ffc_259_n),
    .din(ffc_258_p)
  );


  DROC
  ffc_260
  (
    .doutp(ffc_260_p),
    .doutn(ffc_260_n),
    .din(ffc_259_p)
  );


  DROC
  ffc_261
  (
    .doutp(ffc_261_p),
    .doutn(ffc_261_n),
    .din(ffc_260_p)
  );


  DROC
  ffc_262
  (
    .doutp(ffc_262_p),
    .doutn(ffc_262_n),
    .din(G116_p)
  );


  DROC
  ffc_263
  (
    .doutp(ffc_263_p),
    .doutn(ffc_263_n),
    .din(ffc_262_p)
  );


  DROC
  ffc_264
  (
    .doutp(ffc_264_p),
    .doutn(ffc_264_n),
    .din(ffc_263_p)
  );


  DROC
  ffc_265
  (
    .doutp(ffc_265_p),
    .doutn(ffc_265_n),
    .din(ffc_264_p)
  );


  DROC
  ffc_266
  (
    .doutp(ffc_266_p),
    .doutn(ffc_266_n),
    .din(G117_p)
  );


  DROC
  ffc_267
  (
    .doutp(ffc_267_p),
    .doutn(ffc_267_n),
    .din(G118_p)
  );


  DROC
  ffc_268
  (
    .doutp(ffc_268_p),
    .doutn(ffc_268_n),
    .din(ffc_267_p)
  );


  DROC
  ffc_269
  (
    .doutp(ffc_269_p),
    .doutn(ffc_269_n),
    .din(ffc_268_p)
  );


  DROC
  ffc_270
  (
    .doutp(ffc_270_p),
    .doutn(ffc_270_n),
    .din(ffc_269_p_spl_)
  );


  DROC
  ffc_271
  (
    .doutp(ffc_271_p),
    .doutn(ffc_271_n),
    .din(G119_p)
  );


  DROC
  ffc_272
  (
    .doutp(ffc_272_p),
    .doutn(ffc_272_n),
    .din(ffc_271_p)
  );


  DROC
  ffc_273
  (
    .doutp(ffc_273_p),
    .doutn(ffc_273_n),
    .din(ffc_272_p)
  );


  DROC
  ffc_274
  (
    .doutp(ffc_274_p),
    .doutn(ffc_274_n),
    .din(ffc_273_p)
  );


  DROC
  ffc_275
  (
    .doutp(ffc_275_p),
    .doutn(ffc_275_n),
    .din(G120_p)
  );


  DROC
  ffc_276
  (
    .doutp(ffc_276_p),
    .doutn(ffc_276_n),
    .din(G121_p)
  );


  DROC
  ffc_277
  (
    .doutp(ffc_277_p),
    .doutn(ffc_277_n),
    .din(ffc_276_p)
  );


  DROC
  ffc_278
  (
    .doutp(ffc_278_p),
    .doutn(ffc_278_n),
    .din(ffc_277_p)
  );


  DROC
  ffc_279
  (
    .doutp(ffc_279_p),
    .doutn(ffc_279_n),
    .din(ffc_278_p)
  );


  DROC
  ffc_280
  (
    .doutp(ffc_280_p),
    .doutn(ffc_280_n),
    .din(G122_p)
  );


  DROC
  ffc_281
  (
    .doutp(ffc_281_p),
    .doutn(ffc_281_n),
    .din(ffc_280_p)
  );


  DROC
  ffc_282
  (
    .doutp(ffc_282_p),
    .doutn(ffc_282_n),
    .din(ffc_281_p)
  );


  DROC
  ffc_283
  (
    .doutp(ffc_283_p),
    .doutn(ffc_283_n),
    .din(ffc_282_p)
  );


  DROC
  ffc_284
  (
    .doutp(ffc_284_p),
    .doutn(ffc_284_n),
    .din(G123_p)
  );


  DROC
  ffc_285
  (
    .doutp(ffc_285_p),
    .doutn(ffc_285_n),
    .din(ffc_284_p)
  );


  DROC
  ffc_286
  (
    .doutp(ffc_286_p),
    .doutn(ffc_286_n),
    .din(ffc_285_p)
  );


  DROC
  ffc_287
  (
    .doutp(ffc_287_p),
    .doutn(ffc_287_n),
    .din(ffc_286_p)
  );


  DROC
  ffc_288
  (
    .doutp(ffc_288_p),
    .doutn(ffc_288_n),
    .din(G124_p)
  );


  DROC
  ffc_289
  (
    .doutp(ffc_289_p),
    .doutn(ffc_289_n),
    .din(ffc_288_p)
  );


  DROC
  ffc_290
  (
    .doutp(ffc_290_p),
    .doutn(ffc_290_n),
    .din(ffc_289_p)
  );


  DROC
  ffc_291
  (
    .doutp(ffc_291_p),
    .doutn(ffc_291_n),
    .din(ffc_290_p)
  );


  DROC
  ffc_292
  (
    .doutp(ffc_292_p),
    .doutn(ffc_292_n),
    .din(G125_p)
  );


  DROC
  ffc_293
  (
    .doutp(ffc_293_p),
    .doutn(ffc_293_n),
    .din(ffc_292_p)
  );


  DROC
  ffc_294
  (
    .doutp(ffc_294_p),
    .doutn(ffc_294_n),
    .din(G126_p)
  );


  DROC
  ffc_295
  (
    .doutp(ffc_295_p),
    .doutn(ffc_295_n),
    .din(ffc_294_p)
  );


  DROC
  ffc_296
  (
    .doutp(ffc_296_p),
    .doutn(ffc_296_n),
    .din(ffc_423_p_spl_)
  );


  DROC
  ffc_297
  (
    .doutp(ffc_297_p),
    .doutn(ffc_297_n),
    .din(G127_p)
  );


  DROC
  ffc_298
  (
    .doutp(ffc_298_p),
    .doutn(ffc_298_n),
    .din(G128_p)
  );


  DROC
  ffc_299
  (
    .doutp(ffc_299_p),
    .doutn(ffc_299_n),
    .din(ffc_298_p)
  );


  DROC
  ffc_300
  (
    .doutp(ffc_300_p),
    .doutn(ffc_300_n),
    .din(G129_p)
  );


  DROC
  ffc_301
  (
    .doutp(ffc_301_p),
    .doutn(ffc_301_n),
    .din(ffc_300_p)
  );


  DROC
  ffc_302
  (
    .doutp(ffc_302_p),
    .doutn(ffc_302_n),
    .din(ffc_441_p_spl_)
  );


  DROC
  ffc_303
  (
    .doutp(ffc_303_p),
    .doutn(ffc_303_n),
    .din(G130_p)
  );


  DROC
  ffc_304
  (
    .doutp(ffc_304_p),
    .doutn(ffc_304_n),
    .din(ffc_303_p)
  );


  DROC
  ffc_305
  (
    .doutp(ffc_305_p),
    .doutn(ffc_305_n),
    .din(ffc_304_p)
  );


  DROC
  ffc_306
  (
    .doutp(ffc_306_p),
    .doutn(ffc_306_n),
    .din(G131_p)
  );


  DROC
  ffc_307
  (
    .doutp(ffc_307_p),
    .doutn(ffc_307_n),
    .din(ffc_306_p)
  );


  DROC
  ffc_308
  (
    .doutp(ffc_308_p),
    .doutn(ffc_308_n),
    .din(ffc_307_p)
  );


  DROC
  ffc_309
  (
    .doutp(ffc_309_p),
    .doutn(ffc_309_n),
    .din(G132_p)
  );


  DROC
  ffc_310
  (
    .doutp(ffc_310_p),
    .doutn(ffc_310_n),
    .din(ffc_309_p)
  );


  DROC
  ffc_311
  (
    .doutp(ffc_311_p),
    .doutn(ffc_311_n),
    .din(ffc_310_p)
  );


  DROC
  ffc_312
  (
    .doutp(ffc_312_p),
    .doutn(ffc_312_n),
    .din(ffc_311_p_spl_)
  );


  DROC
  ffc_313
  (
    .doutp(ffc_313_p),
    .doutn(ffc_313_n),
    .din(G133_p)
  );


  DROC
  ffc_314
  (
    .doutp(ffc_314_p),
    .doutn(ffc_314_n),
    .din(ffc_313_p)
  );


  DROC
  ffc_315
  (
    .doutp(ffc_315_p),
    .doutn(ffc_315_n),
    .din(ffc_314_p)
  );


  DROC
  ffc_316
  (
    .doutp(ffc_316_p),
    .doutn(ffc_316_n),
    .din(G134_p)
  );


  DROC
  ffc_317
  (
    .doutp(ffc_317_p),
    .doutn(ffc_317_n),
    .din(ffc_316_p)
  );


  DROC
  ffc_318
  (
    .doutp(ffc_318_p),
    .doutn(ffc_318_n),
    .din(ffc_317_p)
  );


  DROC
  ffc_319
  (
    .doutp(ffc_319_p),
    .doutn(ffc_319_n),
    .din(ffc_318_p_spl_)
  );


  DROC
  ffc_320
  (
    .doutp(ffc_320_p),
    .doutn(ffc_320_n),
    .din(G135_p)
  );


  DROC
  ffc_321
  (
    .doutp(ffc_321_p),
    .doutn(ffc_321_n),
    .din(ffc_320_p)
  );


  DROC
  ffc_322
  (
    .doutp(ffc_322_p),
    .doutn(ffc_322_n),
    .din(ffc_321_p)
  );


  DROC
  ffc_323
  (
    .doutp(ffc_323_p),
    .doutn(ffc_323_n),
    .din(ffc_322_p_spl_)
  );


  DROC
  ffc_324
  (
    .doutp(ffc_324_p),
    .doutn(ffc_324_n),
    .din(G136_p)
  );


  DROC
  ffc_325
  (
    .doutp(ffc_325_p),
    .doutn(ffc_325_n),
    .din(ffc_324_p)
  );


  DROC
  ffc_326
  (
    .doutp(ffc_326_p),
    .doutn(ffc_326_n),
    .din(ffc_428_p_spl_)
  );


  DROC
  ffc_327
  (
    .doutp(ffc_327_p),
    .doutn(ffc_327_n),
    .din(G137_p)
  );


  DROC
  ffc_328
  (
    .doutp(ffc_328_p),
    .doutn(ffc_328_n),
    .din(ffc_327_p)
  );


  DROC
  ffc_329
  (
    .doutp(ffc_329_p),
    .doutn(ffc_329_n),
    .din(ffc_328_p)
  );


  DROC
  ffc_330
  (
    .doutp(ffc_330_p),
    .doutn(ffc_330_n),
    .din(ffc_329_p)
  );


  DROC
  ffc_331
  (
    .doutp(ffc_331_p),
    .doutn(ffc_331_n),
    .din(G138_p)
  );


  DROC
  ffc_332
  (
    .doutp(ffc_332_p),
    .doutn(ffc_332_n),
    .din(ffc_331_p)
  );


  DROC
  ffc_333
  (
    .doutp(ffc_333_p),
    .doutn(ffc_333_n),
    .din(ffc_424_p_spl_)
  );


  DROC
  ffc_334
  (
    .doutp(ffc_334_p),
    .doutn(ffc_334_n),
    .din(G139_p)
  );


  DROC
  ffc_335
  (
    .doutp(ffc_335_p),
    .doutn(ffc_335_n),
    .din(ffc_334_p)
  );


  DROC
  ffc_336
  (
    .doutp(ffc_336_p),
    .doutn(ffc_336_n),
    .din(ffc_442_p_spl_)
  );


  DROC
  ffc_337
  (
    .doutp(ffc_337_p),
    .doutn(ffc_337_n),
    .din(G140_p)
  );


  DROC
  ffc_338
  (
    .doutp(ffc_338_p),
    .doutn(ffc_338_n),
    .din(ffc_337_p)
  );


  DROC
  ffc_339
  (
    .doutp(ffc_339_p),
    .doutn(ffc_339_n),
    .din(ffc_443_p_spl_)
  );


  DROC
  ffc_340
  (
    .doutp(ffc_340_p),
    .doutn(ffc_340_n),
    .din(G141_p)
  );


  DROC
  ffc_341
  (
    .doutp(ffc_341_p),
    .doutn(ffc_341_n),
    .din(ffc_340_p)
  );


  DROC
  ffc_342
  (
    .doutp(ffc_342_p),
    .doutn(ffc_342_n),
    .din(ffc_341_p)
  );


  DROC
  ffc_343
  (
    .doutp(ffc_343_p),
    .doutn(ffc_343_n),
    .din(ffc_342_p_spl_)
  );


  DROC
  ffc_344
  (
    .doutp(ffc_344_p),
    .doutn(ffc_344_n),
    .din(G142_p)
  );


  DROC
  ffc_345
  (
    .doutp(ffc_345_p),
    .doutn(ffc_345_n),
    .din(ffc_344_p)
  );


  DROC
  ffc_346
  (
    .doutp(ffc_346_p),
    .doutn(ffc_346_n),
    .din(ffc_345_p)
  );


  DROC
  ffc_347
  (
    .doutp(ffc_347_p),
    .doutn(ffc_347_n),
    .din(ffc_346_p_spl_)
  );


  DROC
  ffc_348
  (
    .doutp(ffc_348_p),
    .doutn(ffc_348_n),
    .din(G143_p)
  );


  DROC
  ffc_349
  (
    .doutp(ffc_349_p),
    .doutn(ffc_349_n),
    .din(ffc_348_p)
  );


  DROC
  ffc_350
  (
    .doutp(ffc_350_p),
    .doutn(ffc_350_n),
    .din(ffc_349_p)
  );


  DROC
  ffc_351
  (
    .doutp(ffc_351_p),
    .doutn(ffc_351_n),
    .din(ffc_350_p_spl_)
  );


  DROC
  ffc_352
  (
    .doutp(ffc_352_p),
    .doutn(ffc_352_n),
    .din(G144_p)
  );


  DROC
  ffc_353
  (
    .doutp(ffc_353_p),
    .doutn(ffc_353_n),
    .din(ffc_352_p)
  );


  DROC
  ffc_354
  (
    .doutp(ffc_354_p),
    .doutn(ffc_354_n),
    .din(ffc_353_p)
  );


  DROC
  ffc_355
  (
    .doutp(ffc_355_p),
    .doutn(ffc_355_n),
    .din(ffc_354_p_spl_)
  );


  DROC
  ffc_356
  (
    .doutp(ffc_356_p),
    .doutn(ffc_356_n),
    .din(G146_p)
  );


  DROC
  ffc_357
  (
    .doutp(ffc_357_p),
    .doutn(ffc_357_n),
    .din(G147_p)
  );


  DROC
  ffc_358
  (
    .doutp(ffc_358_p),
    .doutn(ffc_358_n),
    .din(ffc_357_p)
  );


  DROC
  ffc_359
  (
    .doutp(ffc_359_p),
    .doutn(ffc_359_n),
    .din(ffc_358_p)
  );


  DROC
  ffc_360
  (
    .doutp(ffc_360_p),
    .doutn(ffc_360_n),
    .din(ffc_359_p)
  );


  DROC
  ffc_361
  (
    .doutp(ffc_361_p),
    .doutn(ffc_361_n),
    .din(G148_p)
  );


  DROC
  ffc_362
  (
    .doutp(ffc_362_p),
    .doutn(ffc_362_n),
    .din(ffc_361_p)
  );


  DROC
  ffc_363
  (
    .doutp(ffc_363_p),
    .doutn(ffc_363_n),
    .din(G149_p)
  );


  DROC
  ffc_364
  (
    .doutp(ffc_364_p),
    .doutn(ffc_364_n),
    .din(ffc_363_p)
  );


  DROC
  ffc_365
  (
    .doutp(ffc_365_p),
    .doutn(ffc_365_n),
    .din(G150_p)
  );


  DROC
  ffc_366
  (
    .doutp(ffc_366_p),
    .doutn(ffc_366_n),
    .din(ffc_365_p)
  );


  DROC
  ffc_367
  (
    .doutp(ffc_367_p),
    .doutn(ffc_367_n),
    .din(ffc_366_p)
  );


  DROC
  ffc_368
  (
    .doutp(ffc_368_p),
    .doutn(ffc_368_n),
    .din(G151_p)
  );


  DROC
  ffc_369
  (
    .doutp(ffc_369_p),
    .doutn(ffc_369_n),
    .din(ffc_368_p)
  );


  DROC
  ffc_370
  (
    .doutp(ffc_370_p),
    .doutn(ffc_370_n),
    .din(ffc_369_p)
  );


  DROC
  ffc_371
  (
    .doutp(ffc_371_p),
    .doutn(ffc_371_n),
    .din(G152_p)
  );


  DROC
  ffc_372
  (
    .doutp(ffc_372_p),
    .doutn(ffc_372_n),
    .din(ffc_371_p)
  );


  DROC
  ffc_373
  (
    .doutp(ffc_373_p),
    .doutn(ffc_373_n),
    .din(G153_p)
  );


  DROC
  ffc_374
  (
    .doutp(ffc_374_p),
    .doutn(ffc_374_n),
    .din(ffc_373_p)
  );


  DROC
  ffc_375
  (
    .doutp(ffc_375_p),
    .doutn(ffc_375_n),
    .din(G154_p)
  );


  DROC
  ffc_376
  (
    .doutp(ffc_376_p),
    .doutn(ffc_376_n),
    .din(ffc_375_p)
  );


  DROC
  ffc_377
  (
    .doutp(ffc_377_p),
    .doutn(ffc_377_n),
    .din(ffc_376_p)
  );


  DROC
  ffc_378
  (
    .doutp(ffc_378_p),
    .doutn(ffc_378_n),
    .din(G155_p)
  );


  DROC
  ffc_379
  (
    .doutp(ffc_379_p),
    .doutn(ffc_379_n),
    .din(ffc_378_p)
  );


  DROC
  ffc_380
  (
    .doutp(ffc_380_p),
    .doutn(ffc_380_n),
    .din(ffc_379_p)
  );


  DROC
  ffc_381
  (
    .doutp(ffc_381_p),
    .doutn(ffc_381_n),
    .din(G156_p)
  );


  DROC
  ffc_382
  (
    .doutp(ffc_382_p),
    .doutn(ffc_382_n),
    .din(ffc_381_p)
  );


  DROC
  ffc_383
  (
    .doutp(ffc_383_p),
    .doutn(ffc_383_n),
    .din(ffc_382_p)
  );


  DROC
  ffc_384
  (
    .doutp(ffc_384_p),
    .doutn(ffc_384_n),
    .din(G157_p)
  );


  DROC
  ffc_385
  (
    .doutp(ffc_385_p),
    .doutn(ffc_385_n),
    .din(ffc_384_p)
  );


  DROC
  ffc_386
  (
    .doutp(ffc_386_p),
    .doutn(ffc_386_n),
    .din(ffc_385_p)
  );


  DROC
  ffc_387
  (
    .doutp(ffc_387_p),
    .doutn(ffc_387_n),
    .din(ffc_413_p)
  );


  DROC
  ffc_388
  (
    .doutp(ffc_388_p),
    .doutn(ffc_388_n),
    .din(ffc_414_p)
  );


  DROC
  ffc_389
  (
    .doutp(ffc_389_p),
    .doutn(ffc_389_n),
    .din(ffc_417_p_spl_1)
  );


  DROC
  ffc_390
  (
    .doutp(ffc_390_p),
    .doutn(ffc_390_n),
    .din(ffc_439_p_spl_1)
  );


  DROC
  ffc_391
  (
    .doutp(ffc_391_p),
    .doutn(ffc_391_n),
    .din(ffc_445_p_spl_1)
  );


  DROC
  ffc_392
  (
    .doutp(ffc_392_p),
    .doutn(ffc_392_n),
    .din(ffc_546_p_spl_1)
  );


  DROC
  ffc_393
  (
    .doutp(ffc_393_p),
    .doutn(ffc_393_n),
    .din(ffc_544_p_spl_1)
  );


  DROC
  ffc_394
  (
    .doutp(ffc_394_p),
    .doutn(ffc_394_n),
    .din(g896_p_spl_)
  );


  DROC
  ffc_395
  (
    .doutp(ffc_395_p),
    .doutn(ffc_395_n),
    .din(g897_p_spl_)
  );


  DROC
  ffc_396
  (
    .doutp(ffc_396_p),
    .doutn(ffc_396_n),
    .din(g898_p_spl_)
  );


  DROC
  ffc_397
  (
    .doutp(ffc_397_p),
    .doutn(ffc_397_n),
    .din(g899_p_spl_)
  );


  DROC
  ffc_398
  (
    .doutp(ffc_398_p),
    .doutn(ffc_398_n),
    .din(g900_n_spl_)
  );


  DROC
  ffc_399
  (
    .doutp(ffc_399_p),
    .doutn(ffc_399_n),
    .din(ffc_444_p_spl_11)
  );


  DROC
  ffc_400
  (
    .doutp(ffc_400_p),
    .doutn(ffc_400_n),
    .din(g901_p_spl_)
  );


  DROC
  ffc_401
  (
    .doutp(ffc_401_p),
    .doutn(ffc_401_n),
    .din(g902_p_spl_)
  );


  DROC
  ffc_402
  (
    .doutp(ffc_402_p),
    .doutn(ffc_402_n),
    .din(g903_n_spl_1)
  );


  DROC
  ffc_403
  (
    .doutp(ffc_403_p),
    .doutn(ffc_403_n),
    .din(g906_p_spl_)
  );


  DROC
  ffc_404
  (
    .doutp(ffc_404_p),
    .doutn(ffc_404_n),
    .din(ffc_504_p_spl_1)
  );


  DROC
  ffc_405
  (
    .doutp(ffc_405_p),
    .doutn(ffc_405_n),
    .din(ffc_532_p_spl_11)
  );


  DROC
  ffc_406
  (
    .doutp(ffc_406_p),
    .doutn(ffc_406_n),
    .din(ffc_533_p_spl_11)
  );


  DROC
  ffc_407
  (
    .doutp(ffc_407_p),
    .doutn(ffc_407_n),
    .din(g907_n_spl_)
  );


  DROC
  ffc_408
  (
    .doutp(ffc_408_p),
    .doutn(ffc_408_n),
    .din(g908_n_spl_1)
  );


  DROC
  ffc_409
  (
    .doutp(ffc_409_p),
    .doutn(ffc_409_n),
    .din(g913_p_spl_)
  );


  DROC
  ffc_410
  (
    .doutp(ffc_410_p),
    .doutn(ffc_410_n),
    .din(g919_n_spl_)
  );


  DROC
  ffc_411
  (
    .doutp(ffc_411_p),
    .doutn(ffc_411_n),
    .din(g925_n_spl_)
  );


  DROC
  ffc_412
  (
    .doutp(ffc_412_p),
    .doutn(ffc_412_n),
    .din(g928_n_spl_)
  );


  DROC
  ffc_413
  (
    .doutp(ffc_413_p),
    .doutn(ffc_413_n),
    .din(ffc_550_p)
  );


  DROC
  ffc_414
  (
    .doutp(ffc_414_p),
    .doutn(ffc_414_n),
    .din(ffc_551_p)
  );


  DROC
  ffc_415
  (
    .doutp(ffc_415_p),
    .doutn(ffc_415_n),
    .din(ffc_563_p_spl_1)
  );


  DROC
  ffc_416
  (
    .doutp(ffc_416_p),
    .doutn(ffc_416_n),
    .din(ffc_564_p_spl_)
  );


  DROC
  ffc_417
  (
    .doutp(ffc_417_p),
    .doutn(ffc_417_n),
    .din(ffc_565_p_spl_)
  );


  DROC
  ffc_418
  (
    .doutp(ffc_418_n),
    .doutn(ffc_418_p),
    .din(g929_n_spl_)
  );


  DROC
  ffc_419
  (
    .doutp(ffc_419_p),
    .doutn(ffc_419_n),
    .din(g938_n_spl_)
  );


  DROC
  ffc_420
  (
    .doutp(ffc_420_p),
    .doutn(ffc_420_n),
    .din(g939_p_spl_)
  );


  DROC
  ffc_421
  (
    .doutp(ffc_421_p),
    .doutn(ffc_421_n),
    .din(g940_p_spl_)
  );


  DROC
  ffc_422
  (
    .doutp(ffc_422_p),
    .doutn(ffc_422_n),
    .din(ffc_293_p_spl_)
  );


  DROC
  ffc_423
  (
    .doutp(ffc_423_p),
    .doutn(ffc_423_n),
    .din(ffc_295_p_spl_)
  );


  DROC
  ffc_424
  (
    .doutp(ffc_424_p),
    .doutn(ffc_424_n),
    .din(ffc_332_p_spl_)
  );


  DROC
  ffc_425
  (
    .doutp(ffc_425_p),
    .doutn(ffc_425_n),
    .din(g941_p_spl_1)
  );


  DROC
  ffc_426
  (
    .doutp(ffc_426_n),
    .doutn(ffc_426_p),
    .din(g942_n_spl_)
  );


  DROC
  ffc_427
  (
    .doutp(ffc_427_n),
    .doutn(ffc_427_p),
    .din(g944_n_spl_)
  );


  DROC
  ffc_428
  (
    .doutp(ffc_428_p),
    .doutn(ffc_428_n),
    .din(ffc_325_p_spl_)
  );


  DROC
  ffc_429
  (
    .doutp(ffc_429_p),
    .doutn(ffc_429_n),
    .din(g945_p_spl_)
  );


  DROC
  ffc_430
  (
    .doutp(ffc_430_p),
    .doutn(ffc_430_n),
    .din(g948_n_spl_)
  );


  DROC
  ffc_431
  (
    .doutp(ffc_431_p),
    .doutn(ffc_431_n),
    .din(g951_n_spl_)
  );


  DROC
  ffc_432
  (
    .doutp(ffc_432_p),
    .doutn(ffc_432_n),
    .din(g954_n_spl_)
  );


  DROC
  ffc_433
  (
    .doutp(ffc_433_p),
    .doutn(ffc_433_n),
    .din(g957_n_spl_)
  );


  DROC
  ffc_434
  (
    .doutp(ffc_434_p),
    .doutn(ffc_434_n),
    .din(g960_n_spl_)
  );


  DROC
  ffc_435
  (
    .doutp(ffc_435_p),
    .doutn(ffc_435_n),
    .din(g963_n_spl_)
  );


  DROC
  ffc_436
  (
    .doutp(ffc_436_p),
    .doutn(ffc_436_n),
    .din(g968_n_spl_)
  );


  DROC
  ffc_437
  (
    .doutp(ffc_437_n),
    .doutn(ffc_437_p),
    .din(g974_n_spl_)
  );


  DROC
  ffc_438
  (
    .doutp(ffc_438_n),
    .doutn(ffc_438_p),
    .din(g980_n_spl_)
  );


  DROC
  ffc_439
  (
    .doutp(ffc_439_p),
    .doutn(ffc_439_n),
    .din(g986_n_spl_)
  );


  DROC
  ffc_440
  (
    .doutp(ffc_440_p),
    .doutn(ffc_440_n),
    .din(ffc_299_p_spl_)
  );


  DROC
  ffc_441
  (
    .doutp(ffc_441_p),
    .doutn(ffc_441_n),
    .din(ffc_301_p_spl_)
  );


  DROC
  ffc_442
  (
    .doutp(ffc_442_p),
    .doutn(ffc_442_n),
    .din(ffc_335_p_spl_)
  );


  DROC
  ffc_443
  (
    .doutp(ffc_443_p),
    .doutn(ffc_443_n),
    .din(ffc_338_p_spl_)
  );


  DROC
  ffc_444
  (
    .doutp(ffc_444_p),
    .doutn(ffc_444_n),
    .din(ffc_574_p_spl_1)
  );


  DROC
  ffc_445
  (
    .doutp(ffc_445_p),
    .doutn(ffc_445_n),
    .din(g995_n_spl_)
  );


  DROC
  ffc_446
  (
    .doutp(ffc_446_p),
    .doutn(ffc_446_n),
    .din(g996_p)
  );


  DROC
  ffc_447
  (
    .doutp(ffc_447_p),
    .doutn(ffc_447_n),
    .din(g997_p)
  );


  DROC
  ffc_448
  (
    .doutp(ffc_448_p),
    .doutn(ffc_448_n),
    .din(g998_p)
  );


  DROC
  ffc_449
  (
    .doutp(ffc_449_p),
    .doutn(ffc_449_n),
    .din(g999_p)
  );


  DROC
  ffc_450
  (
    .doutp(ffc_450_p),
    .doutn(ffc_450_n),
    .din(g1000_p)
  );


  DROC
  ffc_451
  (
    .doutp(ffc_451_p),
    .doutn(ffc_451_n),
    .din(g1001_p)
  );


  DROC
  ffc_452
  (
    .doutp(ffc_452_p),
    .doutn(ffc_452_n),
    .din(g1002_n)
  );


  DROC
  ffc_453
  (
    .doutp(ffc_453_n),
    .doutn(ffc_453_p),
    .din(g1006_n)
  );


  DROC
  ffc_454
  (
    .doutp(ffc_454_p),
    .doutn(ffc_454_n),
    .din(g1007_p)
  );


  DROC
  ffc_455
  (
    .doutp(ffc_455_n),
    .doutn(ffc_455_p),
    .din(g1008_n)
  );


  DROC
  ffc_456
  (
    .doutp(ffc_456_n),
    .doutn(ffc_456_p),
    .din(g1012_n)
  );


  DROC
  ffc_457
  (
    .doutp(ffc_457_p),
    .doutn(ffc_457_n),
    .din(g1013_p)
  );


  DROC
  ffc_458
  (
    .doutp(ffc_458_p),
    .doutn(ffc_458_n),
    .din(g1017_p)
  );


  DROC
  ffc_459
  (
    .doutp(ffc_459_n),
    .doutn(ffc_459_p),
    .din(g1018_n)
  );


  DROC
  ffc_460
  (
    .doutp(ffc_460_p),
    .doutn(ffc_460_n),
    .din(g1022_p)
  );


  DROC
  ffc_461
  (
    .doutp(ffc_461_n),
    .doutn(ffc_461_p),
    .din(g1023_n)
  );


  DROC
  ffc_462
  (
    .doutp(ffc_462_p),
    .doutn(ffc_462_n),
    .din(g1024_p)
  );


  DROC
  ffc_463
  (
    .doutp(ffc_463_p),
    .doutn(ffc_463_n),
    .din(g1025_p)
  );


  DROC
  ffc_464
  (
    .doutp(ffc_464_p),
    .doutn(ffc_464_n),
    .din(g1029_p)
  );


  DROC
  ffc_465
  (
    .doutp(ffc_465_n),
    .doutn(ffc_465_p),
    .din(g1030_n)
  );


  DROC
  ffc_466
  (
    .doutp(ffc_466_p),
    .doutn(ffc_466_n),
    .din(g1031_p)
  );


  DROC
  ffc_467
  (
    .doutp(ffc_467_n),
    .doutn(ffc_467_p),
    .din(g1032_n)
  );


  DROC
  ffc_468
  (
    .doutp(ffc_468_p),
    .doutn(ffc_468_n),
    .din(g1033_p)
  );


  DROC
  ffc_469
  (
    .doutp(ffc_469_n),
    .doutn(ffc_469_p),
    .din(g1034_n)
  );


  DROC
  ffc_470
  (
    .doutp(ffc_470_p),
    .doutn(ffc_470_n),
    .din(g1035_p)
  );


  DROC
  ffc_471
  (
    .doutp(ffc_471_p),
    .doutn(ffc_471_n),
    .din(g1036_p)
  );


  DROC
  ffc_472
  (
    .doutp(ffc_472_p),
    .doutn(ffc_472_n),
    .din(g1037_p)
  );


  DROC
  ffc_473
  (
    .doutp(ffc_473_p),
    .doutn(ffc_473_n),
    .din(g1038_p)
  );


  DROC
  ffc_474
  (
    .doutp(ffc_474_p),
    .doutn(ffc_474_n),
    .din(g1039_p)
  );


  DROC
  ffc_475
  (
    .doutp(ffc_475_n),
    .doutn(ffc_475_p),
    .din(g1040_n_spl_)
  );


  DROC
  ffc_476
  (
    .doutp(ffc_476_p),
    .doutn(ffc_476_n),
    .din(g1043_n)
  );


  DROC
  ffc_477
  (
    .doutp(ffc_477_n),
    .doutn(ffc_477_p),
    .din(g1044_n)
  );


  DROC
  ffc_478
  (
    .doutp(ffc_478_p),
    .doutn(ffc_478_n),
    .din(g1047_n)
  );


  DROC
  ffc_479
  (
    .doutp(ffc_479_p),
    .doutn(ffc_479_n),
    .din(g1053_n)
  );


  DROC
  ffc_480
  (
    .doutp(ffc_480_p),
    .doutn(ffc_480_n),
    .din(g1057_n)
  );


  DROC
  ffc_481
  (
    .doutp(ffc_481_p),
    .doutn(ffc_481_n),
    .din(g1060_n)
  );


  DROC
  ffc_482
  (
    .doutp(ffc_482_p),
    .doutn(ffc_482_n),
    .din(g1063_n)
  );


  DROC
  ffc_483
  (
    .doutp(ffc_483_p),
    .doutn(ffc_483_n),
    .din(g1066_n)
  );


  DROC
  ffc_484
  (
    .doutp(ffc_484_n),
    .doutn(ffc_484_p),
    .din(g1067_n)
  );


  DROC
  ffc_485
  (
    .doutp(ffc_485_p),
    .doutn(ffc_485_n),
    .din(g1070_n)
  );


  DROC
  ffc_486
  (
    .doutp(ffc_486_p),
    .doutn(ffc_486_n),
    .din(g1073_p)
  );


  DROC
  ffc_487
  (
    .doutp(ffc_487_n),
    .doutn(ffc_487_p),
    .din(g1074_n)
  );


  DROC
  ffc_488
  (
    .doutp(ffc_488_p),
    .doutn(ffc_488_n),
    .din(g1077_p)
  );


  DROC
  ffc_489
  (
    .doutp(ffc_489_n),
    .doutn(ffc_489_p),
    .din(g1078_n)
  );


  DROC
  ffc_490
  (
    .doutp(ffc_490_n),
    .doutn(ffc_490_p),
    .din(g1095_n)
  );


  DROC
  ffc_491
  (
    .doutp(ffc_491_n),
    .doutn(ffc_491_p),
    .din(g1097_p)
  );


  DROC
  ffc_492
  (
    .doutp(ffc_492_n),
    .doutn(ffc_492_p),
    .din(g1108_n)
  );


  DROC
  ffc_493
  (
    .doutp(ffc_493_p),
    .doutn(ffc_493_n),
    .din(g1109_p)
  );


  DROC
  ffc_494
  (
    .doutp(ffc_494_n),
    .doutn(ffc_494_p),
    .din(g1113_p)
  );


  DROC
  ffc_495
  (
    .doutp(ffc_495_n),
    .doutn(ffc_495_p),
    .din(g1114_n)
  );


  DROC
  ffc_496
  (
    .doutp(ffc_496_p),
    .doutn(ffc_496_n),
    .din(g1123_n)
  );


  DROC
  ffc_497
  (
    .doutp(ffc_497_p),
    .doutn(ffc_497_n),
    .din(g1132_n)
  );


  DROC
  ffc_498
  (
    .doutp(ffc_498_p),
    .doutn(ffc_498_n),
    .din(g1138_p)
  );


  DROC
  ffc_499
  (
    .doutp(ffc_499_p),
    .doutn(ffc_499_n),
    .din(g1153_p)
  );


  DROC
  ffc_500
  (
    .doutp(ffc_500_p),
    .doutn(ffc_500_n),
    .din(g1160_p)
  );


  DROC
  ffc_501
  (
    .doutp(ffc_501_n),
    .doutn(ffc_501_p),
    .din(g1161_n)
  );


  DROC
  ffc_502
  (
    .doutp(ffc_502_p),
    .doutn(ffc_502_n),
    .din(g1176_n)
  );


  DROC
  ffc_503
  (
    .doutp(ffc_503_n),
    .doutn(ffc_503_p),
    .din(g1183_n_spl_)
  );


  DROC
  ffc_504
  (
    .doutp(ffc_504_p),
    .doutn(ffc_504_n),
    .din(ffc_356_p_spl_)
  );


  DROC
  ffc_505
  (
    .doutp(ffc_505_p),
    .doutn(ffc_505_n),
    .din(ffc_26_p)
  );


  DROC
  ffc_506
  (
    .doutp(ffc_506_p),
    .doutn(ffc_506_n),
    .din(ffc_123_p)
  );


  DROC
  ffc_507
  (
    .doutp(ffc_507_p),
    .doutn(ffc_507_n),
    .din(ffc_125_p)
  );


  DROC
  ffc_508
  (
    .doutp(ffc_508_p),
    .doutn(ffc_508_n),
    .din(ffc_130_p)
  );


  DROC
  ffc_509
  (
    .doutp(ffc_509_p),
    .doutn(ffc_509_n),
    .din(ffc_170_p)
  );


  DROC
  ffc_510
  (
    .doutp(ffc_510_p),
    .doutn(ffc_510_n),
    .din(ffc_193_p)
  );


  DROC
  ffc_511
  (
    .doutp(ffc_511_p),
    .doutn(ffc_511_n),
    .din(ffc_211_p)
  );


  DROC
  ffc_512
  (
    .doutp(ffc_512_p),
    .doutn(ffc_512_n),
    .din(ffc_229_p)
  );


  DROC
  ffc_513
  (
    .doutp(ffc_513_p),
    .doutn(ffc_513_n),
    .din(ffc_247_p)
  );


  DROC
  ffc_514
  (
    .doutp(ffc_514_p),
    .doutn(ffc_514_n),
    .din(ffc_362_p)
  );


  DROC
  ffc_515
  (
    .doutp(ffc_515_p),
    .doutn(ffc_515_n),
    .din(ffc_364_p)
  );


  DROC
  ffc_516
  (
    .doutp(ffc_516_p),
    .doutn(ffc_516_n),
    .din(ffc_372_p)
  );


  DROC
  ffc_517
  (
    .doutp(ffc_517_p),
    .doutn(ffc_517_n),
    .din(ffc_374_p)
  );


  DROC
  ffc_518
  (
    .doutp(ffc_518_p),
    .doutn(ffc_518_n),
    .din(g1184_p)
  );


  DROC
  ffc_519
  (
    .doutp(ffc_519_p),
    .doutn(ffc_519_n),
    .din(g1185_p)
  );


  DROC
  ffc_520
  (
    .doutp(ffc_520_p),
    .doutn(ffc_520_n),
    .din(g1186_p)
  );


  DROC
  ffc_521
  (
    .doutp(ffc_521_p),
    .doutn(ffc_521_n),
    .din(g1187_p)
  );


  DROC
  ffc_522
  (
    .doutp(ffc_522_p),
    .doutn(ffc_522_n),
    .din(g1188_p)
  );


  DROC
  ffc_523
  (
    .doutp(ffc_523_p),
    .doutn(ffc_523_n),
    .din(g1189_p)
  );


  DROC
  ffc_524
  (
    .doutp(ffc_524_p),
    .doutn(ffc_524_n),
    .din(g1190_p)
  );


  DROC
  ffc_525
  (
    .doutp(ffc_525_p),
    .doutn(ffc_525_n),
    .din(g1191_p)
  );


  DROC
  ffc_526
  (
    .doutp(ffc_526_p),
    .doutn(ffc_526_n),
    .din(g1192_p)
  );


  DROC
  ffc_527
  (
    .doutp(ffc_527_p),
    .doutn(ffc_527_n),
    .din(g1193_n)
  );


  DROC
  ffc_528
  (
    .doutp(ffc_528_p),
    .doutn(ffc_528_n),
    .din(g1195_p)
  );


  DROC
  ffc_529
  (
    .doutp(ffc_529_p),
    .doutn(ffc_529_n),
    .din(g1197_n)
  );


  DROC
  ffc_530
  (
    .doutp(ffc_530_p),
    .doutn(ffc_530_n),
    .din(g1201_p)
  );


  DROC
  ffc_531
  (
    .doutp(ffc_531_p),
    .doutn(ffc_531_n),
    .din(g1205_p)
  );


  DROC
  ffc_532
  (
    .doutp(ffc_532_p),
    .doutn(ffc_532_n),
    .din(ffc_266_p_spl_)
  );


  DROC
  ffc_533
  (
    .doutp(ffc_533_p),
    .doutn(ffc_533_n),
    .din(ffc_275_p)
  );


  DROC
  ffc_534
  (
    .doutp(ffc_534_p),
    .doutn(ffc_534_n),
    .din(g1208_n)
  );


  DROC
  ffc_535
  (
    .doutp(ffc_535_p),
    .doutn(ffc_535_n),
    .din(g1211_n)
  );


  DROC
  ffc_536
  (
    .doutp(ffc_536_p),
    .doutn(ffc_536_n),
    .din(g1214_n)
  );


  DROC
  ffc_537
  (
    .doutp(ffc_537_p),
    .doutn(ffc_537_n),
    .din(g1217_n)
  );


  DROC
  ffc_538
  (
    .doutp(ffc_538_p),
    .doutn(ffc_538_n),
    .din(g1220_n)
  );


  DROC
  ffc_539
  (
    .doutp(ffc_539_p),
    .doutn(ffc_539_n),
    .din(g1223_n)
  );


  DROC
  ffc_540
  (
    .doutp(ffc_540_p),
    .doutn(ffc_540_n),
    .din(g1232_n)
  );


  DROC
  ffc_541
  (
    .doutp(ffc_541_p),
    .doutn(ffc_541_n),
    .din(g1241_n)
  );


  DROC
  ffc_542
  (
    .doutp(ffc_542_p),
    .doutn(ffc_542_n),
    .din(g1250_n)
  );


  DROC
  ffc_543
  (
    .doutp(ffc_543_p),
    .doutn(ffc_543_n),
    .din(g1254_n)
  );


  DROC
  ffc_544
  (
    .doutp(ffc_544_p),
    .doutn(ffc_544_n),
    .din(g1263_n)
  );


  DROC
  ffc_545
  (
    .doutp(ffc_545_p),
    .doutn(ffc_545_n),
    .din(g1267_n)
  );


  DROC
  ffc_546
  (
    .doutp(ffc_546_n),
    .doutn(ffc_546_p),
    .din(g1268_p)
  );


  DROC
  ffc_547
  (
    .doutp(ffc_547_p),
    .doutn(ffc_547_n),
    .din(g1271_p)
  );


  DROC
  ffc_548
  (
    .doutp(ffc_548_p),
    .doutn(ffc_548_n),
    .din(g1274_p)
  );


  DROC
  ffc_549
  (
    .doutp(ffc_549_p),
    .doutn(ffc_549_n),
    .din(g1280_p)
  );


  DROC
  ffc_550
  (
    .doutp(ffc_550_n),
    .doutn(ffc_550_p),
    .din(g1284_n_spl_)
  );


  DROC
  ffc_551
  (
    .doutp(ffc_551_n),
    .doutn(ffc_551_p),
    .din(g1288_n_spl_)
  );


  DROC
  ffc_552
  (
    .doutp(ffc_552_p),
    .doutn(ffc_552_n),
    .din(ffc_111_p)
  );


  DROC
  ffc_553
  (
    .doutp(ffc_553_p),
    .doutn(ffc_553_n),
    .din(ffc_135_p)
  );


  DROC
  ffc_554
  (
    .doutp(ffc_554_p),
    .doutn(ffc_554_n),
    .din(ffc_95_p)
  );


  DROC
  ffc_555
  (
    .doutp(ffc_555_p),
    .doutn(ffc_555_n),
    .din(ffc_114_p)
  );


  DROC
  ffc_556
  (
    .doutp(ffc_556_p),
    .doutn(ffc_556_n),
    .din(ffc_117_p)
  );


  DROC
  ffc_557
  (
    .doutp(ffc_557_p),
    .doutn(ffc_557_n),
    .din(ffc_157_p)
  );


  DROC
  ffc_558
  (
    .doutp(ffc_558_p),
    .doutn(ffc_558_n),
    .din(ffc_179_p)
  );


  DROC
  ffc_559
  (
    .doutp(ffc_559_p),
    .doutn(ffc_559_n),
    .din(ffc_297_p)
  );


  DROC
  ffc_560
  (
    .doutp(ffc_560_p),
    .doutn(ffc_560_n),
    .din(g1289_p)
  );


  DROC
  ffc_561
  (
    .doutp(ffc_561_p),
    .doutn(ffc_561_n),
    .din(g1290_p)
  );


  DROC
  ffc_562
  (
    .doutp(ffc_562_p),
    .doutn(ffc_562_n),
    .din(g1291_p)
  );


  DROC
  ffc_563
  (
    .doutp(ffc_563_p),
    .doutn(ffc_563_n),
    .din(g1292_p)
  );


  DROC
  ffc_564
  (
    .doutp(ffc_564_n),
    .doutn(ffc_564_p),
    .din(g1293_p)
  );


  DROC
  ffc_565
  (
    .doutp(ffc_565_p),
    .doutn(ffc_565_n),
    .din(g1302_n)
  );


  DROC
  ffc_566
  (
    .doutp(ffc_566_p),
    .doutn(ffc_566_n),
    .din(G79_p)
  );


  DROC
  ffc_567
  (
    .doutp(ffc_567_p),
    .doutn(ffc_567_n),
    .din(G80_p)
  );


  DROC
  ffc_568
  (
    .doutp(ffc_568_p),
    .doutn(ffc_568_n),
    .din(G89_p)
  );


  DROC
  ffc_569
  (
    .doutp(ffc_569_p),
    .doutn(ffc_569_n),
    .din(G90_p)
  );


  DROC
  ffc_570
  (
    .doutp(ffc_570_p),
    .doutn(ffc_570_n),
    .din(G99_p)
  );


  DROC
  ffc_571
  (
    .doutp(ffc_571_p),
    .doutn(ffc_571_n),
    .din(G100_p)
  );


  DROC
  ffc_572
  (
    .doutp(ffc_572_p),
    .doutn(ffc_572_n),
    .din(G109_p)
  );


  DROC
  ffc_573
  (
    .doutp(ffc_573_p),
    .doutn(ffc_573_n),
    .din(G110_p)
  );


  DROC
  ffc_574
  (
    .doutp(ffc_574_p),
    .doutn(ffc_574_n),
    .din(G145_p)
  );


  buf

  (
    ffc_279_n_spl_,
    ffc_279_n
  );


  buf

  (
    ffc_261_n_spl_,
    ffc_261_n
  );


  buf

  (
    ffc_261_n_spl_0,
    ffc_261_n_spl_
  );


  buf

  (
    ffc_261_n_spl_1,
    ffc_261_n_spl_
  );


  buf

  (
    g737_n_spl_,
    g737_n
  );


  buf

  (
    g737_n_spl_0,
    g737_n_spl_
  );


  buf

  (
    g740_n_spl_,
    g740_n
  );


  buf

  (
    g741_n_spl_,
    g741_n
  );


  buf

  (
    ffc_283_n_spl_,
    ffc_283_n
  );


  buf

  (
    ffc_283_n_spl_0,
    ffc_283_n_spl_
  );


  buf

  (
    g745_n_spl_,
    g745_n
  );


  buf

  (
    g745_n_spl_0,
    g745_n_spl_
  );


  buf

  (
    g752_n_spl_,
    g752_n
  );


  buf

  (
    ffc_287_p_spl_,
    ffc_287_p
  );


  buf

  (
    ffc_287_p_spl_0,
    ffc_287_p_spl_
  );


  buf

  (
    ffc_287_p_spl_1,
    ffc_287_p_spl_
  );


  buf

  (
    ffc_391_n_spl_,
    ffc_391_n
  );


  buf

  (
    ffc_287_n_spl_,
    ffc_287_n
  );


  buf

  (
    ffc_287_n_spl_0,
    ffc_287_n_spl_
  );


  buf

  (
    ffc_287_n_spl_1,
    ffc_287_n_spl_
  );


  buf

  (
    ffc_392_p_spl_,
    ffc_392_p
  );


  buf

  (
    g749_n_spl_,
    g749_n
  );


  buf

  (
    ffc_270_p_spl_,
    ffc_270_p
  );


  buf

  (
    ffc_391_p_spl_,
    ffc_391_p
  );


  buf

  (
    ffc_452_n_spl_,
    ffc_452_n
  );


  buf

  (
    ffc_452_n_spl_0,
    ffc_452_n_spl_
  );


  buf

  (
    ffc_483_p_spl_,
    ffc_483_p
  );


  buf

  (
    ffc_485_n_spl_,
    ffc_485_n
  );


  buf

  (
    ffc_483_n_spl_,
    ffc_483_n
  );


  buf

  (
    ffc_485_p_spl_,
    ffc_485_p
  );


  buf

  (
    ffc_482_n_spl_,
    ffc_482_n
  );


  buf

  (
    ffc_497_p_spl_,
    ffc_497_p
  );


  buf

  (
    ffc_482_p_spl_,
    ffc_482_p
  );


  buf

  (
    ffc_497_n_spl_,
    ffc_497_n
  );


  buf

  (
    ffc_398_p_spl_,
    ffc_398_p
  );


  buf

  (
    ffc_94_n_spl_,
    ffc_94_n
  );


  buf

  (
    ffc_438_n_spl_,
    ffc_438_n
  );


  buf

  (
    ffc_452_p_spl_,
    ffc_452_p
  );


  buf

  (
    ffc_438_p_spl_,
    ffc_438_p
  );


  buf

  (
    g851_p_spl_,
    g851_p
  );


  buf

  (
    g851_n_spl_,
    g851_n
  );


  buf

  (
    g868_n_spl_,
    g868_n
  );


  buf

  (
    ffc_491_p_spl_,
    ffc_491_p
  );


  buf

  (
    g875_n_spl_,
    g875_n
  );


  buf

  (
    g877_n_spl_,
    g877_n
  );


  buf

  (
    g876_n_spl_,
    g876_n
  );


  buf

  (
    g774_p_spl_,
    g774_p
  );


  buf

  (
    g779_p_spl_,
    g779_p
  );


  buf

  (
    g788_p_spl_,
    g788_p
  );


  buf

  (
    g849_p_spl_,
    g849_p
  );


  buf

  (
    g864_p_spl_,
    g864_p
  );


  buf

  (
    ffc_415_p_spl_,
    ffc_415_p
  );


  buf

  (
    ffc_415_p_spl_0,
    ffc_415_p_spl_
  );


  buf

  (
    ffc_415_p_spl_1,
    ffc_415_p_spl_
  );


  buf

  (
    ffc_415_n_spl_,
    ffc_415_n
  );


  buf

  (
    ffc_415_n_spl_0,
    ffc_415_n_spl_
  );


  buf

  (
    ffc_415_n_spl_1,
    ffc_415_n_spl_
  );


  buf

  (
    ffc_404_p_spl_,
    ffc_404_p
  );


  buf

  (
    ffc_404_p_spl_0,
    ffc_404_p_spl_
  );


  buf

  (
    ffc_404_p_spl_00,
    ffc_404_p_spl_0
  );


  buf

  (
    ffc_404_p_spl_01,
    ffc_404_p_spl_0
  );


  buf

  (
    ffc_404_p_spl_1,
    ffc_404_p_spl_
  );


  buf

  (
    ffc_404_p_spl_10,
    ffc_404_p_spl_1
  );


  buf

  (
    ffc_404_p_spl_11,
    ffc_404_p_spl_1
  );


  buf

  (
    ffc_404_n_spl_,
    ffc_404_n
  );


  buf

  (
    ffc_404_n_spl_0,
    ffc_404_n_spl_
  );


  buf

  (
    ffc_404_n_spl_00,
    ffc_404_n_spl_0
  );


  buf

  (
    ffc_404_n_spl_01,
    ffc_404_n_spl_0
  );


  buf

  (
    ffc_404_n_spl_1,
    ffc_404_n_spl_
  );


  buf

  (
    ffc_404_n_spl_10,
    ffc_404_n_spl_1
  );


  buf

  (
    ffc_404_n_spl_11,
    ffc_404_n_spl_1
  );


  buf

  (
    ffc_442_p_spl_,
    ffc_442_p
  );


  buf

  (
    ffc_442_p_spl_0,
    ffc_442_p_spl_
  );


  buf

  (
    ffc_443_p_spl_,
    ffc_443_p
  );


  buf

  (
    ffc_443_p_spl_0,
    ffc_443_p_spl_
  );


  buf

  (
    ffc_442_n_spl_,
    ffc_442_n
  );


  buf

  (
    ffc_442_n_spl_0,
    ffc_442_n_spl_
  );


  buf

  (
    ffc_443_n_spl_,
    ffc_443_n
  );


  buf

  (
    ffc_443_n_spl_0,
    ffc_443_n_spl_
  );


  buf

  (
    g896_p_spl_,
    g896_p
  );


  buf

  (
    g899_p_spl_,
    g899_p
  );


  buf

  (
    ffc_406_n_spl_,
    ffc_406_n
  );


  buf

  (
    ffc_406_n_spl_0,
    ffc_406_n_spl_
  );


  buf

  (
    ffc_406_n_spl_00,
    ffc_406_n_spl_0
  );


  buf

  (
    ffc_406_n_spl_01,
    ffc_406_n_spl_0
  );


  buf

  (
    ffc_406_n_spl_1,
    ffc_406_n_spl_
  );


  buf

  (
    ffc_406_p_spl_,
    ffc_406_p
  );


  buf

  (
    ffc_406_p_spl_0,
    ffc_406_p_spl_
  );


  buf

  (
    ffc_406_p_spl_00,
    ffc_406_p_spl_0
  );


  buf

  (
    ffc_406_p_spl_01,
    ffc_406_p_spl_0
  );


  buf

  (
    ffc_406_p_spl_1,
    ffc_406_p_spl_
  );


  buf

  (
    g901_p_spl_,
    g901_p
  );


  buf

  (
    g906_p_spl_,
    g906_p
  );


  buf

  (
    ffc_405_n_spl_,
    ffc_405_n
  );


  buf

  (
    ffc_405_p_spl_,
    ffc_405_p
  );


  buf

  (
    ffc_439_n_spl_,
    ffc_439_n
  );


  buf

  (
    g900_n_spl_,
    g900_n
  );


  buf

  (
    g900_n_spl_0,
    g900_n_spl_
  );


  buf

  (
    ffc_439_p_spl_,
    ffc_439_p
  );


  buf

  (
    ffc_439_p_spl_0,
    ffc_439_p_spl_
  );


  buf

  (
    ffc_439_p_spl_1,
    ffc_439_p_spl_
  );


  buf

  (
    g900_p_spl_,
    g900_p
  );


  buf

  (
    ffc_342_n_spl_,
    ffc_342_n
  );


  buf

  (
    ffc_342_n_spl_0,
    ffc_342_n_spl_
  );


  buf

  (
    ffc_346_n_spl_,
    ffc_346_n
  );


  buf

  (
    ffc_399_n_spl_,
    ffc_399_n
  );


  buf

  (
    ffc_399_n_spl_0,
    ffc_399_n_spl_
  );


  buf

  (
    ffc_399_n_spl_1,
    ffc_399_n_spl_
  );


  buf

  (
    ffc_399_p_spl_,
    ffc_399_p
  );


  buf

  (
    ffc_399_p_spl_0,
    ffc_399_p_spl_
  );


  buf

  (
    ffc_399_p_spl_1,
    ffc_399_p_spl_
  );


  buf

  (
    ffc_564_p_spl_,
    ffc_564_p
  );


  buf

  (
    ffc_565_p_spl_,
    ffc_565_p
  );


  buf

  (
    g939_p_spl_,
    g939_p
  );


  buf

  (
    g940_p_spl_,
    g940_p
  );


  buf

  (
    ffc_505_n_spl_,
    ffc_505_n
  );


  buf

  (
    g908_n_spl_,
    g908_n
  );


  buf

  (
    g908_n_spl_0,
    g908_n_spl_
  );


  buf

  (
    g908_n_spl_1,
    g908_n_spl_
  );


  buf

  (
    ffc_318_p_spl_,
    ffc_318_p
  );


  buf

  (
    ffc_318_p_spl_0,
    ffc_318_p_spl_
  );


  buf

  (
    g943_n_spl_,
    g943_n
  );


  buf

  (
    g943_n_spl_0,
    g943_n_spl_
  );


  buf

  (
    g943_n_spl_00,
    g943_n_spl_0
  );


  buf

  (
    g943_n_spl_1,
    g943_n_spl_
  );


  buf

  (
    g925_p_spl_,
    g925_p
  );


  buf

  (
    g943_p_spl_,
    g943_p
  );


  buf

  (
    g943_p_spl_0,
    g943_p_spl_
  );


  buf

  (
    g943_p_spl_00,
    g943_p_spl_0
  );


  buf

  (
    g943_p_spl_1,
    g943_p_spl_
  );


  buf

  (
    ffc_41_p_spl_,
    ffc_41_p
  );


  buf

  (
    ffc_41_p_spl_0,
    ffc_41_p_spl_
  );


  buf

  (
    ffc_41_p_spl_00,
    ffc_41_p_spl_0
  );


  buf

  (
    ffc_41_p_spl_000,
    ffc_41_p_spl_00
  );


  buf

  (
    ffc_41_p_spl_01,
    ffc_41_p_spl_0
  );


  buf

  (
    ffc_41_p_spl_1,
    ffc_41_p_spl_
  );


  buf

  (
    ffc_41_p_spl_10,
    ffc_41_p_spl_1
  );


  buf

  (
    ffc_41_p_spl_11,
    ffc_41_p_spl_1
  );


  buf

  (
    ffc_41_n_spl_,
    ffc_41_n
  );


  buf

  (
    ffc_41_n_spl_0,
    ffc_41_n_spl_
  );


  buf

  (
    ffc_41_n_spl_00,
    ffc_41_n_spl_0
  );


  buf

  (
    ffc_41_n_spl_000,
    ffc_41_n_spl_00
  );


  buf

  (
    ffc_41_n_spl_01,
    ffc_41_n_spl_0
  );


  buf

  (
    ffc_41_n_spl_1,
    ffc_41_n_spl_
  );


  buf

  (
    ffc_41_n_spl_10,
    ffc_41_n_spl_1
  );


  buf

  (
    ffc_41_n_spl_11,
    ffc_41_n_spl_1
  );


  buf

  (
    ffc_445_p_spl_,
    ffc_445_p
  );


  buf

  (
    ffc_445_p_spl_0,
    ffc_445_p_spl_
  );


  buf

  (
    ffc_445_p_spl_00,
    ffc_445_p_spl_0
  );


  buf

  (
    ffc_445_p_spl_1,
    ffc_445_p_spl_
  );


  buf

  (
    g925_n_spl_,
    g925_n
  );


  buf

  (
    g925_n_spl_0,
    g925_n_spl_
  );


  buf

  (
    g913_p_spl_,
    g913_p
  );


  buf

  (
    g913_p_spl_0,
    g913_p_spl_
  );


  buf

  (
    ffc_74_p_spl_,
    ffc_74_p
  );


  buf

  (
    ffc_74_p_spl_0,
    ffc_74_p_spl_
  );


  buf

  (
    ffc_74_p_spl_00,
    ffc_74_p_spl_0
  );


  buf

  (
    ffc_74_p_spl_01,
    ffc_74_p_spl_0
  );


  buf

  (
    ffc_74_p_spl_1,
    ffc_74_p_spl_
  );


  buf

  (
    ffc_74_p_spl_10,
    ffc_74_p_spl_1
  );


  buf

  (
    ffc_74_p_spl_11,
    ffc_74_p_spl_1
  );


  buf

  (
    ffc_74_n_spl_,
    ffc_74_n
  );


  buf

  (
    ffc_74_n_spl_0,
    ffc_74_n_spl_
  );


  buf

  (
    ffc_74_n_spl_00,
    ffc_74_n_spl_0
  );


  buf

  (
    ffc_74_n_spl_01,
    ffc_74_n_spl_0
  );


  buf

  (
    ffc_74_n_spl_1,
    ffc_74_n_spl_
  );


  buf

  (
    ffc_74_n_spl_10,
    ffc_74_n_spl_1
  );


  buf

  (
    ffc_74_n_spl_11,
    ffc_74_n_spl_1
  );


  buf

  (
    ffc_417_p_spl_,
    ffc_417_p
  );


  buf

  (
    ffc_417_p_spl_0,
    ffc_417_p_spl_
  );


  buf

  (
    ffc_417_p_spl_1,
    ffc_417_p_spl_
  );


  buf

  (
    ffc_540_p_spl_,
    ffc_540_p
  );


  buf

  (
    ffc_540_p_spl_0,
    ffc_540_p_spl_
  );


  buf

  (
    ffc_416_p_spl_,
    ffc_416_p
  );


  buf

  (
    ffc_416_p_spl_0,
    ffc_416_p_spl_
  );


  buf

  (
    ffc_505_p_spl_,
    ffc_505_p
  );


  buf

  (
    ffc_308_n_spl_,
    ffc_308_n
  );


  buf

  (
    ffc_308_n_spl_0,
    ffc_308_n_spl_
  );


  buf

  (
    ffc_308_n_spl_00,
    ffc_308_n_spl_0
  );


  buf

  (
    ffc_308_n_spl_1,
    ffc_308_n_spl_
  );


  buf

  (
    g964_p_spl_,
    g964_p
  );


  buf

  (
    g964_p_spl_0,
    g964_p_spl_
  );


  buf

  (
    g964_p_spl_1,
    g964_p_spl_
  );


  buf

  (
    g966_p_spl_,
    g966_p
  );


  buf

  (
    g966_p_spl_0,
    g966_p_spl_
  );


  buf

  (
    g966_p_spl_1,
    g966_p_spl_
  );


  buf

  (
    g971_n_spl_,
    g971_n
  );


  buf

  (
    g971_n_spl_0,
    g971_n_spl_
  );


  buf

  (
    g971_n_spl_1,
    g971_n_spl_
  );


  buf

  (
    g971_p_spl_,
    g971_p
  );


  buf

  (
    g971_p_spl_0,
    g971_p_spl_
  );


  buf

  (
    ffc_428_n_spl_,
    ffc_428_n
  );


  buf

  (
    ffc_428_p_spl_,
    ffc_428_p
  );


  buf

  (
    ffc_428_p_spl_0,
    ffc_428_p_spl_
  );


  buf

  (
    ffc_544_p_spl_,
    ffc_544_p
  );


  buf

  (
    ffc_544_p_spl_0,
    ffc_544_p_spl_
  );


  buf

  (
    ffc_544_p_spl_00,
    ffc_544_p_spl_0
  );


  buf

  (
    ffc_544_p_spl_01,
    ffc_544_p_spl_0
  );


  buf

  (
    ffc_544_p_spl_1,
    ffc_544_p_spl_
  );


  buf

  (
    ffc_445_n_spl_,
    ffc_445_n
  );


  buf

  (
    ffc_544_n_spl_,
    ffc_544_n
  );


  buf

  (
    g928_n_spl_,
    g928_n
  );


  buf

  (
    ffc_533_p_spl_,
    ffc_533_p
  );


  buf

  (
    ffc_533_p_spl_0,
    ffc_533_p_spl_
  );


  buf

  (
    ffc_533_p_spl_00,
    ffc_533_p_spl_0
  );


  buf

  (
    ffc_533_p_spl_000,
    ffc_533_p_spl_00
  );


  buf

  (
    ffc_533_p_spl_001,
    ffc_533_p_spl_00
  );


  buf

  (
    ffc_533_p_spl_01,
    ffc_533_p_spl_0
  );


  buf

  (
    ffc_533_p_spl_010,
    ffc_533_p_spl_01
  );


  buf

  (
    ffc_533_p_spl_1,
    ffc_533_p_spl_
  );


  buf

  (
    ffc_533_p_spl_10,
    ffc_533_p_spl_1
  );


  buf

  (
    ffc_533_p_spl_11,
    ffc_533_p_spl_1
  );


  buf

  (
    ffc_563_p_spl_,
    ffc_563_p
  );


  buf

  (
    ffc_563_p_spl_0,
    ffc_563_p_spl_
  );


  buf

  (
    ffc_563_p_spl_00,
    ffc_563_p_spl_0
  );


  buf

  (
    ffc_563_p_spl_1,
    ffc_563_p_spl_
  );


  buf

  (
    ffc_533_n_spl_,
    ffc_533_n
  );


  buf

  (
    ffc_533_n_spl_0,
    ffc_533_n_spl_
  );


  buf

  (
    ffc_533_n_spl_00,
    ffc_533_n_spl_0
  );


  buf

  (
    ffc_533_n_spl_1,
    ffc_533_n_spl_
  );


  buf

  (
    ffc_532_p_spl_,
    ffc_532_p
  );


  buf

  (
    ffc_532_p_spl_0,
    ffc_532_p_spl_
  );


  buf

  (
    ffc_532_p_spl_00,
    ffc_532_p_spl_0
  );


  buf

  (
    ffc_532_p_spl_000,
    ffc_532_p_spl_00
  );


  buf

  (
    ffc_532_p_spl_001,
    ffc_532_p_spl_00
  );


  buf

  (
    ffc_532_p_spl_01,
    ffc_532_p_spl_0
  );


  buf

  (
    ffc_532_p_spl_1,
    ffc_532_p_spl_
  );


  buf

  (
    ffc_532_p_spl_10,
    ffc_532_p_spl_1
  );


  buf

  (
    ffc_532_p_spl_11,
    ffc_532_p_spl_1
  );


  buf

  (
    ffc_532_n_spl_,
    ffc_532_n
  );


  buf

  (
    ffc_532_n_spl_0,
    ffc_532_n_spl_
  );


  buf

  (
    ffc_532_n_spl_00,
    ffc_532_n_spl_0
  );


  buf

  (
    ffc_532_n_spl_000,
    ffc_532_n_spl_00
  );


  buf

  (
    ffc_532_n_spl_001,
    ffc_532_n_spl_00
  );


  buf

  (
    ffc_532_n_spl_01,
    ffc_532_n_spl_0
  );


  buf

  (
    ffc_532_n_spl_010,
    ffc_532_n_spl_01
  );


  buf

  (
    ffc_532_n_spl_011,
    ffc_532_n_spl_01
  );


  buf

  (
    ffc_532_n_spl_1,
    ffc_532_n_spl_
  );


  buf

  (
    ffc_532_n_spl_10,
    ffc_532_n_spl_1
  );


  buf

  (
    ffc_532_n_spl_100,
    ffc_532_n_spl_10
  );


  buf

  (
    ffc_532_n_spl_101,
    ffc_532_n_spl_10
  );


  buf

  (
    ffc_532_n_spl_11,
    ffc_532_n_spl_1
  );


  buf

  (
    ffc_532_n_spl_110,
    ffc_532_n_spl_11
  );


  buf

  (
    g938_n_spl_,
    g938_n
  );


  buf

  (
    g938_n_spl_0,
    g938_n_spl_
  );


  buf

  (
    ffc_99_p_spl_,
    ffc_99_p
  );


  buf

  (
    ffc_163_p_spl_,
    ffc_163_p
  );


  buf

  (
    ffc_120_p_spl_,
    ffc_120_p
  );


  buf

  (
    ffc_141_p_spl_,
    ffc_141_p
  );


  buf

  (
    ffc_190_p_spl_,
    ffc_190_p
  );


  buf

  (
    ffc_244_p_spl_,
    ffc_244_p
  );


  buf

  (
    ffc_208_p_spl_,
    ffc_208_p
  );


  buf

  (
    ffc_226_p_spl_,
    ffc_226_p
  );


  buf

  (
    ffc_269_p_spl_,
    ffc_269_p
  );


  buf

  (
    ffc_422_n_spl_,
    ffc_422_n
  );


  buf

  (
    ffc_422_n_spl_0,
    ffc_422_n_spl_
  );


  buf

  (
    ffc_422_n_spl_1,
    ffc_422_n_spl_
  );


  buf

  (
    g1005_n_spl_,
    g1005_n
  );


  buf

  (
    ffc_423_n_spl_,
    ffc_423_n
  );


  buf

  (
    ffc_423_n_spl_0,
    ffc_423_n_spl_
  );


  buf

  (
    g948_n_spl_,
    g948_n
  );


  buf

  (
    ffc_440_n_spl_,
    ffc_440_n
  );


  buf

  (
    ffc_440_n_spl_0,
    ffc_440_n_spl_
  );


  buf

  (
    ffc_440_n_spl_1,
    ffc_440_n_spl_
  );


  buf

  (
    g1011_n_spl_,
    g1011_n
  );


  buf

  (
    g903_n_spl_,
    g903_n
  );


  buf

  (
    g903_n_spl_0,
    g903_n_spl_
  );


  buf

  (
    g903_n_spl_1,
    g903_n_spl_
  );


  buf

  (
    ffc_305_n_spl_,
    ffc_305_n
  );


  buf

  (
    ffc_305_n_spl_0,
    ffc_305_n_spl_
  );


  buf

  (
    ffc_305_n_spl_1,
    ffc_305_n_spl_
  );


  buf

  (
    g1016_n_spl_,
    g1016_n
  );


  buf

  (
    g1021_n_spl_,
    g1021_n
  );


  buf

  (
    ffc_311_n_spl_,
    ffc_311_n
  );


  buf

  (
    ffc_311_n_spl_0,
    ffc_311_n_spl_
  );


  buf

  (
    ffc_311_n_spl_1,
    ffc_311_n_spl_
  );


  buf

  (
    g954_n_spl_,
    g954_n
  );


  buf

  (
    g919_n_spl_,
    g919_n
  );


  buf

  (
    g919_n_spl_0,
    g919_n_spl_
  );


  buf

  (
    ffc_315_n_spl_,
    ffc_315_n
  );


  buf

  (
    ffc_315_n_spl_0,
    ffc_315_n_spl_
  );


  buf

  (
    ffc_315_n_spl_1,
    ffc_315_n_spl_
  );


  buf

  (
    g1028_n_spl_,
    g1028_n
  );


  buf

  (
    ffc_318_n_spl_,
    ffc_318_n
  );


  buf

  (
    g951_n_spl_,
    g951_n
  );


  buf

  (
    g960_n_spl_,
    g960_n
  );


  buf

  (
    g957_n_spl_,
    g957_n
  );


  buf

  (
    g963_n_spl_,
    g963_n
  );


  buf

  (
    ffc_350_p_spl_,
    ffc_350_p
  );


  buf

  (
    ffc_354_p_spl_,
    ffc_354_p
  );


  buf

  (
    g919_p_spl_,
    g919_p
  );


  buf

  (
    g913_n_spl_,
    g913_n
  );


  buf

  (
    ffc_546_p_spl_,
    ffc_546_p
  );


  buf

  (
    ffc_546_p_spl_0,
    ffc_546_p_spl_
  );


  buf

  (
    ffc_546_p_spl_1,
    ffc_546_p_spl_
  );


  buf

  (
    g942_n_spl_,
    g942_n
  );


  buf

  (
    g968_n_spl_,
    g968_n
  );


  buf

  (
    ffc_541_p_spl_,
    ffc_541_p
  );


  buf

  (
    ffc_541_p_spl_0,
    ffc_541_p_spl_
  );


  buf

  (
    g1051_n_spl_,
    g1051_n
  );


  buf

  (
    g1051_n_spl_0,
    g1051_n_spl_
  );


  buf

  (
    g1051_n_spl_1,
    g1051_n_spl_
  );


  buf

  (
    g897_p_spl_,
    g897_p
  );


  buf

  (
    g898_p_spl_,
    g898_p
  );


  buf

  (
    g1055_n_spl_,
    g1055_n
  );


  buf

  (
    g1055_n_spl_0,
    g1055_n_spl_
  );


  buf

  (
    ffc_441_p_spl_,
    ffc_441_p
  );


  buf

  (
    g944_n_spl_,
    g944_n
  );


  buf

  (
    g945_p_spl_,
    g945_p
  );


  buf

  (
    ffc_322_p_spl_,
    ffc_322_p
  );


  buf

  (
    ffc_322_n_spl_,
    ffc_322_n
  );


  buf

  (
    ffc_541_n_spl_,
    ffc_541_n
  );


  buf

  (
    ffc_541_n_spl_0,
    ffc_541_n_spl_
  );


  buf

  (
    g1071_n_spl_,
    g1071_n
  );


  buf

  (
    g1072_p_spl_,
    g1072_p
  );


  buf

  (
    ffc_424_n_spl_,
    ffc_424_n
  );


  buf

  (
    ffc_424_n_spl_0,
    ffc_424_n_spl_
  );


  buf

  (
    g1075_n_spl_,
    g1075_n
  );


  buf

  (
    g1076_p_spl_,
    g1076_p
  );


  buf

  (
    g1079_n_spl_,
    g1079_n
  );


  buf

  (
    g1082_n_spl_,
    g1082_n
  );


  buf

  (
    ffc_548_n_spl_,
    ffc_548_n
  );


  buf

  (
    ffc_547_n_spl_,
    ffc_547_n
  );


  buf

  (
    g974_n_spl_,
    g974_n
  );


  buf

  (
    ffc_342_p_spl_,
    ffc_342_p
  );


  buf

  (
    ffc_346_p_spl_,
    ffc_346_p
  );


  buf

  (
    g929_n_spl_,
    g929_n
  );


  buf

  (
    g902_p_spl_,
    g902_p
  );


  buf

  (
    ffc_386_n_spl_,
    ffc_386_n
  );


  buf

  (
    ffc_386_p_spl_,
    ffc_386_p
  );


  buf

  (
    ffc_424_p_spl_,
    ffc_424_p
  );


  buf

  (
    ffc_424_p_spl_0,
    ffc_424_p_spl_
  );


  buf

  (
    g1099_p_spl_,
    g1099_p
  );


  buf

  (
    g1107_p_spl_,
    g1107_p
  );


  buf

  (
    g907_n_spl_,
    g907_n
  );


  buf

  (
    g980_n_spl_,
    g980_n
  );


  buf

  (
    g980_n_spl_0,
    g980_n_spl_
  );


  buf

  (
    g1112_n_spl_,
    g1112_n
  );


  buf

  (
    ffc_377_p_spl_,
    ffc_377_p
  );


  buf

  (
    ffc_380_n_spl_,
    ffc_380_n
  );


  buf

  (
    ffc_377_n_spl_,
    ffc_377_n
  );


  buf

  (
    ffc_380_p_spl_,
    ffc_380_p
  );


  buf

  (
    ffc_422_p_spl_,
    ffc_422_p
  );


  buf

  (
    ffc_423_p_spl_,
    ffc_423_p
  );


  buf

  (
    ffc_423_p_spl_0,
    ffc_423_p_spl_
  );


  buf

  (
    ffc_308_p_spl_,
    ffc_308_p
  );


  buf

  (
    ffc_311_p_spl_,
    ffc_311_p
  );


  buf

  (
    ffc_311_p_spl_0,
    ffc_311_p_spl_
  );


  buf

  (
    ffc_383_n_spl_,
    ffc_383_n
  );


  buf

  (
    ffc_383_p_spl_,
    ffc_383_p
  );


  buf

  (
    ffc_440_p_spl_,
    ffc_440_p
  );


  buf

  (
    ffc_416_n_spl_,
    ffc_416_n
  );


  buf

  (
    g1055_p_spl_,
    g1055_p
  );


  buf

  (
    ffc_516_p_spl_,
    ffc_516_p
  );


  buf

  (
    ffc_517_n_spl_,
    ffc_517_n
  );


  buf

  (
    ffc_516_n_spl_,
    ffc_516_n
  );


  buf

  (
    ffc_517_p_spl_,
    ffc_517_p
  );


  buf

  (
    ffc_514_p_spl_,
    ffc_514_p
  );


  buf

  (
    ffc_515_n_spl_,
    ffc_515_n
  );


  buf

  (
    ffc_514_n_spl_,
    ffc_514_n
  );


  buf

  (
    ffc_515_p_spl_,
    ffc_515_p
  );


  buf

  (
    g1141_p_spl_,
    g1141_p
  );


  buf

  (
    g1144_p_spl_,
    g1144_p
  );


  buf

  (
    g1141_n_spl_,
    g1141_n
  );


  buf

  (
    g1144_n_spl_,
    g1144_n
  );


  buf

  (
    ffc_367_p_spl_,
    ffc_367_p
  );


  buf

  (
    ffc_370_n_spl_,
    ffc_370_n
  );


  buf

  (
    ffc_367_n_spl_,
    ffc_367_n
  );


  buf

  (
    ffc_370_p_spl_,
    ffc_370_p
  );


  buf

  (
    g1156_n_spl_,
    g1156_n
  );


  buf

  (
    g1159_p_spl_,
    g1159_p
  );


  buf

  (
    ffc_542_p_spl_,
    ffc_542_p
  );


  buf

  (
    ffc_542_n_spl_,
    ffc_542_n
  );


  buf

  (
    ffc_417_n_spl_,
    ffc_417_n
  );


  buf

  (
    ffc_540_n_spl_,
    ffc_540_n
  );


  buf

  (
    g1164_p_spl_,
    g1164_p
  );


  buf

  (
    g1167_p_spl_,
    g1167_p
  );


  buf

  (
    g1164_n_spl_,
    g1164_n
  );


  buf

  (
    g1167_n_spl_,
    g1167_n
  );


  buf

  (
    g1051_p_spl_,
    g1051_p
  );


  buf

  (
    ffc_332_p_spl_,
    ffc_332_p
  );


  buf

  (
    g941_n_spl_,
    g941_n
  );


  buf

  (
    g941_n_spl_0,
    g941_n_spl_
  );


  buf

  (
    g941_n_spl_1,
    g941_n_spl_
  );


  buf

  (
    ffc_295_p_spl_,
    ffc_295_p
  );


  buf

  (
    g941_p_spl_,
    g941_p
  );


  buf

  (
    g941_p_spl_0,
    g941_p_spl_
  );


  buf

  (
    g941_p_spl_00,
    g941_p_spl_0
  );


  buf

  (
    g941_p_spl_1,
    g941_p_spl_
  );


  buf

  (
    g995_n_spl_,
    g995_n
  );


  buf

  (
    g995_n_spl_0,
    g995_n_spl_
  );


  buf

  (
    g1204_p_spl_,
    g1204_p
  );


  buf

  (
    ffc_444_n_spl_,
    ffc_444_n
  );


  buf

  (
    ffc_444_n_spl_0,
    ffc_444_n_spl_
  );


  buf

  (
    ffc_444_n_spl_00,
    ffc_444_n_spl_0
  );


  buf

  (
    ffc_444_n_spl_000,
    ffc_444_n_spl_00
  );


  buf

  (
    ffc_444_n_spl_001,
    ffc_444_n_spl_00
  );


  buf

  (
    ffc_444_n_spl_01,
    ffc_444_n_spl_0
  );


  buf

  (
    ffc_444_n_spl_010,
    ffc_444_n_spl_01
  );


  buf

  (
    ffc_444_n_spl_011,
    ffc_444_n_spl_01
  );


  buf

  (
    ffc_444_n_spl_1,
    ffc_444_n_spl_
  );


  buf

  (
    ffc_444_n_spl_10,
    ffc_444_n_spl_1
  );


  buf

  (
    ffc_444_n_spl_11,
    ffc_444_n_spl_1
  );


  buf

  (
    ffc_444_p_spl_,
    ffc_444_p
  );


  buf

  (
    ffc_444_p_spl_0,
    ffc_444_p_spl_
  );


  buf

  (
    ffc_444_p_spl_00,
    ffc_444_p_spl_0
  );


  buf

  (
    ffc_444_p_spl_000,
    ffc_444_p_spl_00
  );


  buf

  (
    ffc_444_p_spl_001,
    ffc_444_p_spl_00
  );


  buf

  (
    ffc_444_p_spl_01,
    ffc_444_p_spl_0
  );


  buf

  (
    ffc_444_p_spl_010,
    ffc_444_p_spl_01
  );


  buf

  (
    ffc_444_p_spl_011,
    ffc_444_p_spl_01
  );


  buf

  (
    ffc_444_p_spl_1,
    ffc_444_p_spl_
  );


  buf

  (
    ffc_444_p_spl_10,
    ffc_444_p_spl_1
  );


  buf

  (
    ffc_444_p_spl_100,
    ffc_444_p_spl_10
  );


  buf

  (
    ffc_444_p_spl_11,
    ffc_444_p_spl_1
  );


  buf

  (
    ffc_504_p_spl_,
    ffc_504_p
  );


  buf

  (
    ffc_504_p_spl_0,
    ffc_504_p_spl_
  );


  buf

  (
    ffc_504_p_spl_1,
    ffc_504_p_spl_
  );


  buf

  (
    ffc_504_n_spl_,
    ffc_504_n
  );


  buf

  (
    ffc_504_n_spl_0,
    ffc_504_n_spl_
  );


  buf

  (
    g1040_n_spl_,
    g1040_n
  );


  buf

  (
    g1183_n_spl_,
    g1183_n
  );


  buf

  (
    ffc_335_p_spl_,
    ffc_335_p
  );


  buf

  (
    ffc_299_p_spl_,
    ffc_299_p
  );


  buf

  (
    ffc_338_p_spl_,
    ffc_338_p
  );


  buf

  (
    ffc_301_p_spl_,
    ffc_301_p
  );


  buf

  (
    ffc_325_p_spl_,
    ffc_325_p
  );


  buf

  (
    ffc_293_p_spl_,
    ffc_293_p
  );


  buf

  (
    g986_n_spl_,
    g986_n
  );


  buf

  (
    ffc_574_p_spl_,
    ffc_574_p
  );


  buf

  (
    ffc_574_p_spl_0,
    ffc_574_p_spl_
  );


  buf

  (
    ffc_574_p_spl_00,
    ffc_574_p_spl_0
  );


  buf

  (
    ffc_574_p_spl_1,
    ffc_574_p_spl_
  );


  buf

  (
    ffc_574_n_spl_,
    ffc_574_n
  );


  buf

  (
    ffc_574_n_spl_0,
    ffc_574_n_spl_
  );


  buf

  (
    ffc_574_n_spl_1,
    ffc_574_n_spl_
  );


  buf

  (
    ffc_356_n_spl_,
    ffc_356_n
  );


  buf

  (
    ffc_356_p_spl_,
    ffc_356_p
  );


  buf

  (
    ffc_356_p_spl_0,
    ffc_356_p_spl_
  );


  buf

  (
    ffc_266_n_spl_,
    ffc_266_n
  );


  buf

  (
    ffc_266_p_spl_,
    ffc_266_p
  );


  buf

  (
    ffc_266_p_spl_0,
    ffc_266_p_spl_
  );


  buf

  (
    g1284_n_spl_,
    g1284_n
  );


  buf

  (
    g1288_n_spl_,
    g1288_n
  );


  buf

  (
    ffc_291_n_spl_,
    ffc_291_n
  );


  buf

  (
    ffc_330_n_spl_,
    ffc_330_n
  );


  buf

  (
    ffc_330_n_spl_0,
    ffc_330_n_spl_
  );


  buf

  (
    g742_n_spl_,
    g742_n
  );


  buf

  (
    g758_p_spl_,
    g758_p
  );


  buf

  (
    g761_n_spl_,
    g761_n
  );


  buf

  (
    g766_p_spl_,
    g766_p
  );


  buf

  (
    g838_n_spl_,
    g838_n
  );


  buf

  (
    g859_p_spl_,
    g859_p
  );


  buf

  (
    g895_n_spl_,
    g895_n
  );


endmodule
