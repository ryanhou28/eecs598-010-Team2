module tb();

reg [0:177] in_ram [0:9];
reg [0:177] inz;
wire [0:122] outz;
reg clk=0;
c5315_clk dup(clk,
inz[0],
inz[1],
inz[2],
inz[3],
inz[4],
inz[5],
inz[6],
inz[7],
inz[8],
inz[9],
inz[10],
inz[11],
inz[12],
inz[13],
inz[14],
inz[15],
inz[16],
inz[17],
inz[18],
inz[19],
inz[20],
inz[21],
inz[22],
inz[23],
inz[24],
inz[25],
inz[26],
inz[27],
inz[28],
inz[29],
inz[30],
inz[31],
inz[32],
inz[33],
inz[34],
inz[35],
inz[36],
inz[37],
inz[38],
inz[39],
inz[40],
inz[41],
inz[42],
inz[43],
inz[44],
inz[45],
inz[46],
inz[47],
inz[48],
inz[49],
inz[50],
inz[51],
inz[52],
inz[53],
inz[54],
inz[55],
inz[56],
inz[57],
inz[58],
inz[59],
inz[60],
inz[61],
inz[62],
inz[63],
inz[64],
inz[65],
inz[66],
inz[67],
inz[68],
inz[69],
inz[70],
inz[71],
inz[72],
inz[73],
inz[74],
inz[75],
inz[76],
inz[77],
inz[78],
inz[79],
inz[80],
inz[81],
inz[82],
inz[83],
inz[84],
inz[85],
inz[86],
inz[87],
inz[88],
inz[89],
inz[90],
inz[91],
inz[92],
inz[93],
inz[94],
inz[95],
inz[96],
inz[97],
inz[98],
inz[99],
inz[100],
inz[101],
inz[102],
inz[103],
inz[104],
inz[105],
inz[106],
inz[107],
inz[108],
inz[109],
inz[110],
inz[111],
inz[112],
inz[113],
inz[114],
inz[115],
inz[116],
inz[117],
inz[118],
inz[119],
inz[120],
inz[121],
inz[122],
inz[123],
inz[124],
inz[125],
inz[126],
inz[127],
inz[128],
inz[129],
inz[130],
inz[131],
inz[132],
inz[133],
inz[134],
inz[135],
inz[136],
inz[137],
inz[138],
inz[139],
inz[140],
inz[141],
inz[142],
inz[143],
inz[144],
inz[145],
inz[146],
inz[147],
inz[148],
inz[149],
inz[150],
inz[151],
inz[152],
inz[153],
inz[154],
inz[155],
inz[156],
inz[157],
inz[158],
inz[159],
inz[160],
inz[161],
inz[162],
inz[163],
inz[164],
inz[165],
inz[166],
inz[167],
inz[168],
inz[169],
inz[170],
inz[171],
inz[172],
inz[173],
inz[174],
inz[175],
inz[176],
inz[177],
outz[0],
outz[1],
outz[2],
outz[3],
outz[4],
outz[5],
outz[6],
outz[7],
outz[8],
outz[9],
outz[10],
outz[11],
outz[12],
outz[13],
outz[14],
outz[15],
outz[16],
outz[17],
outz[18],
outz[19],
outz[20],
outz[21],
outz[22],
outz[23],
outz[24],
outz[25],
outz[26],
outz[27],
outz[28],
outz[29],
outz[30],
outz[31],
outz[32],
outz[33],
outz[34],
outz[35],
outz[36],
outz[37],
outz[38],
outz[39],
outz[40],
outz[41],
outz[42],
outz[43],
outz[44],
outz[45],
outz[46],
outz[47],
outz[48],
outz[49],
outz[50],
outz[51],
outz[52],
outz[53],
outz[54],
outz[55],
outz[56],
outz[57],
outz[58],
outz[59],
outz[60],
outz[61],
outz[62],
outz[63],
outz[64],
outz[65],
outz[66],
outz[67],
outz[68],
outz[69],
outz[70],
outz[71],
outz[72],
outz[73],
outz[74],
outz[75],
outz[76],
outz[77],
outz[78],
outz[79],
outz[80],
outz[81],
outz[82],
outz[83],
outz[84],
outz[85],
outz[86],
outz[87],
outz[88],
outz[89],
outz[90],
outz[91],
outz[92],
outz[93],
outz[94],
outz[95],
outz[96],
outz[97],
outz[98],
outz[99],
outz[100],
outz[101],
outz[102],
outz[103],
outz[104],
outz[105],
outz[106],
outz[107],
outz[108],
outz[109],
outz[110],
outz[111],
outz[112],
outz[113],
outz[114],
outz[115],
outz[116],
outz[117],
outz[118],
outz[119],
outz[120],
outz[121],
outz[122]
);

initial begin 
  $readmemb("l5315.txt", in_ram);
  for (integer i = 0; i < 13; i=i+1) begin
  inz <= in_ram[i];
  #10 clk<=~clk;
  #10 clk<=~clk;
  $displayb(outz);
  end
end

endmodule
