
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  G42,
  G43,
  G44,
  G45,
  G46,
  G47,
  G48,
  G49,
  G50,
  G51,
  G52,
  G53,
  G54,
  G55,
  G56,
  G57,
  G58,
  G59,
  G60,
  G61,
  G62,
  G63,
  G64,
  G65,
  G66,
  G67,
  G68,
  G69,
  G70,
  G71,
  G72,
  G73,
  G74,
  G75,
  G76,
  G77,
  G78,
  G79,
  G80,
  G81,
  G82,
  G83,
  G84,
  G85,
  G86,
  G87,
  G88,
  G89,
  G90,
  G91,
  G92,
  G93,
  G94,
  G95,
  G96,
  G97,
  G98,
  G99,
  G100,
  G101,
  G102,
  G103,
  G104,
  G105,
  G106,
  G107,
  G108,
  G109,
  G110,
  G111,
  G112,
  G113,
  G114,
  G115,
  G116,
  G117,
  G118,
  G119,
  G120,
  G121,
  G122,
  G123,
  G124,
  G125,
  G126,
  G127,
  G128,
  G129,
  G130,
  G131,
  G132,
  G133,
  G134,
  G135,
  G136,
  G137,
  G138,
  G139,
  G140,
  G141,
  G142,
  G143,
  G144,
  G145,
  G146,
  G147,
  G148,
  G149,
  G150,
  G151,
  G152,
  G153,
  G154,
  G155,
  G156,
  G157,
  G2531,
  G2532,
  G2533,
  G2534,
  G2535,
  G2536,
  G2537,
  G2538,
  G2539,
  G2540,
  G2541,
  G2542,
  G2543,
  G2544,
  G2545,
  G2546,
  G2547,
  G2548,
  G2549,
  G2550,
  G2551,
  G2552,
  G2553,
  G2554,
  G2555,
  G2556,
  G2557,
  G2558,
  G2559,
  G2560,
  G2561,
  G2562,
  G2563,
  G2564,
  G2565,
  G2566,
  G2567,
  G2568,
  G2569,
  G2570,
  G2571,
  G2572,
  G2573,
  G2574,
  G2575,
  G2576,
  G2577,
  G2578,
  G2579,
  G2580,
  G2581,
  G2582,
  G2583,
  G2584,
  G2585,
  G2586,
  G2587,
  G2588,
  G2589,
  G2590,
  G2591,
  G2592,
  G2593,
  G2594
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input G42;input G43;input G44;input G45;input G46;input G47;input G48;input G49;input G50;input G51;input G52;input G53;input G54;input G55;input G56;input G57;input G58;input G59;input G60;input G61;input G62;input G63;input G64;input G65;input G66;input G67;input G68;input G69;input G70;input G71;input G72;input G73;input G74;input G75;input G76;input G77;input G78;input G79;input G80;input G81;input G82;input G83;input G84;input G85;input G86;input G87;input G88;input G89;input G90;input G91;input G92;input G93;input G94;input G95;input G96;input G97;input G98;input G99;input G100;input G101;input G102;input G103;input G104;input G105;input G106;input G107;input G108;input G109;input G110;input G111;input G112;input G113;input G114;input G115;input G116;input G117;input G118;input G119;input G120;input G121;input G122;input G123;input G124;input G125;input G126;input G127;input G128;input G129;input G130;input G131;input G132;input G133;input G134;input G135;input G136;input G137;input G138;input G139;input G140;input G141;input G142;input G143;input G144;input G145;input G146;input G147;input G148;input G149;input G150;input G151;input G152;input G153;input G154;input G155;input G156;input G157;
  output G2531;output G2532;output G2533;output G2534;output G2535;output G2536;output G2537;output G2538;output G2539;output G2540;output G2541;output G2542;output G2543;output G2544;output G2545;output G2546;output G2547;output G2548;output G2549;output G2550;output G2551;output G2552;output G2553;output G2554;output G2555;output G2556;output G2557;output G2558;output G2559;output G2560;output G2561;output G2562;output G2563;output G2564;output G2565;output G2566;output G2567;output G2568;output G2569;output G2570;output G2571;output G2572;output G2573;output G2574;output G2575;output G2576;output G2577;output G2578;output G2579;output G2580;output G2581;output G2582;output G2583;output G2584;output G2585;output G2586;output G2587;output G2588;output G2589;output G2590;output G2591;output G2592;output G2593;output G2594;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire G51_p;
  wire G51_n;
  wire G52_p;
  wire G52_n;
  wire G53_p;
  wire G53_n;
  wire G54_p;
  wire G54_n;
  wire G55_p;
  wire G55_n;
  wire G56_p;
  wire G56_n;
  wire G57_p;
  wire G57_n;
  wire G58_p;
  wire G58_n;
  wire G59_p;
  wire G59_n;
  wire G60_p;
  wire G60_n;
  wire G61_p;
  wire G61_n;
  wire G62_p;
  wire G62_n;
  wire G63_p;
  wire G63_n;
  wire G64_p;
  wire G64_n;
  wire G65_p;
  wire G65_n;
  wire G66_p;
  wire G66_n;
  wire G67_p;
  wire G67_n;
  wire G68_p;
  wire G68_n;
  wire G69_p;
  wire G69_n;
  wire G70_p;
  wire G70_n;
  wire G71_p;
  wire G71_n;
  wire G72_p;
  wire G72_n;
  wire G73_p;
  wire G73_n;
  wire G74_p;
  wire G74_n;
  wire G75_p;
  wire G75_n;
  wire G76_p;
  wire G76_n;
  wire G77_p;
  wire G77_n;
  wire G78_p;
  wire G78_n;
  wire G79_p;
  wire G79_n;
  wire G80_p;
  wire G80_n;
  wire G81_p;
  wire G81_n;
  wire G82_p;
  wire G82_n;
  wire G83_p;
  wire G83_n;
  wire G84_p;
  wire G84_n;
  wire G85_p;
  wire G85_n;
  wire G86_p;
  wire G86_n;
  wire G87_p;
  wire G87_n;
  wire G88_p;
  wire G88_n;
  wire G89_p;
  wire G89_n;
  wire G90_p;
  wire G90_n;
  wire G91_p;
  wire G91_n;
  wire G92_p;
  wire G92_n;
  wire G93_p;
  wire G93_n;
  wire G94_p;
  wire G94_n;
  wire G95_p;
  wire G95_n;
  wire G96_p;
  wire G96_n;
  wire G97_p;
  wire G97_n;
  wire G98_p;
  wire G98_n;
  wire G99_p;
  wire G99_n;
  wire G100_p;
  wire G100_n;
  wire G101_p;
  wire G101_n;
  wire G102_p;
  wire G102_n;
  wire G103_p;
  wire G103_n;
  wire G104_p;
  wire G104_n;
  wire G105_p;
  wire G105_n;
  wire G106_p;
  wire G106_n;
  wire G107_p;
  wire G107_n;
  wire G108_p;
  wire G108_n;
  wire G109_p;
  wire G109_n;
  wire G110_p;
  wire G110_n;
  wire G111_p;
  wire G111_n;
  wire G112_p;
  wire G112_n;
  wire G113_p;
  wire G113_n;
  wire G114_p;
  wire G114_n;
  wire G115_p;
  wire G115_n;
  wire G116_p;
  wire G116_n;
  wire G117_p;
  wire G117_n;
  wire G118_p;
  wire G118_n;
  wire G119_p;
  wire G119_n;
  wire G120_p;
  wire G120_n;
  wire G121_p;
  wire G121_n;
  wire G122_p;
  wire G122_n;
  wire G123_p;
  wire G123_n;
  wire G124_p;
  wire G124_n;
  wire G125_p;
  wire G125_n;
  wire G126_p;
  wire G126_n;
  wire G127_p;
  wire G127_n;
  wire G128_p;
  wire G128_n;
  wire G129_p;
  wire G129_n;
  wire G130_p;
  wire G130_n;
  wire G131_p;
  wire G131_n;
  wire G132_p;
  wire G132_n;
  wire G133_p;
  wire G133_n;
  wire G134_p;
  wire G134_n;
  wire G135_p;
  wire G135_n;
  wire G136_p;
  wire G136_n;
  wire G137_p;
  wire G137_n;
  wire G138_p;
  wire G138_n;
  wire G139_p;
  wire G139_n;
  wire G140_p;
  wire G140_n;
  wire G141_p;
  wire G141_n;
  wire G142_p;
  wire G142_n;
  wire G143_p;
  wire G143_n;
  wire G144_p;
  wire G144_n;
  wire G145_p;
  wire G145_n;
  wire G146_p;
  wire G146_n;
  wire G147_p;
  wire G147_n;
  wire G148_p;
  wire G148_n;
  wire G149_p;
  wire G149_n;
  wire G150_p;
  wire G150_n;
  wire G151_p;
  wire G151_n;
  wire G152_p;
  wire G152_n;
  wire G153_p;
  wire G153_n;
  wire G154_p;
  wire G154_n;
  wire G155_p;
  wire G155_n;
  wire G156_p;
  wire G156_n;
  wire G157_p;
  wire G157_n;
  wire g158_p;
  wire g158_n;
  wire g159_p;
  wire g159_n;
  wire g160_p;
  wire g160_n;
  wire g161_p;
  wire g161_n;
  wire g162_p;
  wire g162_n;
  wire g163_p;
  wire g163_n;
  wire g164_p;
  wire g164_n;
  wire g165_p;
  wire g165_n;
  wire g166_p;
  wire g166_n;
  wire g167_p;
  wire g167_n;
  wire g168_p;
  wire g168_n;
  wire g169_p;
  wire g169_n;
  wire g170_p;
  wire g170_n;
  wire g171_p;
  wire g171_n;
  wire g172_p;
  wire g172_n;
  wire g173_p;
  wire g173_n;
  wire g174_p;
  wire g174_n;
  wire g175_p;
  wire g175_n;
  wire g176_p;
  wire g176_n;
  wire g177_p;
  wire g177_n;
  wire g178_p;
  wire g178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire g686_p;
  wire g686_n;
  wire g687_p;
  wire g687_n;
  wire g688_p;
  wire g688_n;
  wire g689_p;
  wire g689_n;
  wire g690_p;
  wire g690_n;
  wire g691_p;
  wire g691_n;
  wire g692_p;
  wire g692_n;
  wire g693_p;
  wire g693_n;
  wire g694_p;
  wire g694_n;
  wire g695_p;
  wire g695_n;
  wire g696_p;
  wire g696_n;
  wire g697_p;
  wire g697_n;
  wire g698_p;
  wire g698_n;
  wire g699_p;
  wire g699_n;
  wire g700_p;
  wire g700_n;
  wire g701_p;
  wire g701_n;
  wire g702_p;
  wire g702_n;
  wire g703_p;
  wire g703_n;
  wire g704_p;
  wire g704_n;
  wire g705_p;
  wire g705_n;
  wire g706_p;
  wire g706_n;
  wire g707_p;
  wire g707_n;
  wire g708_p;
  wire g708_n;
  wire g709_p;
  wire g709_n;
  wire g710_p;
  wire g710_n;
  wire g711_p;
  wire g711_n;
  wire g712_p;
  wire g712_n;
  wire g713_p;
  wire g713_n;
  wire g714_p;
  wire g714_n;
  wire g715_p;
  wire g715_n;
  wire g716_p;
  wire g716_n;
  wire g717_p;
  wire g717_n;
  wire g718_p;
  wire g718_n;
  wire G142_p_spl_;
  wire G142_p_spl_0;
  wire G142_p_spl_1;
  wire G141_p_spl_;
  wire G141_p_spl_0;
  wire G141_p_spl_1;
  wire G142_n_spl_;
  wire G142_n_spl_0;
  wire G141_n_spl_;
  wire G141_n_spl_0;
  wire G140_p_spl_;
  wire G140_p_spl_0;
  wire G140_p_spl_1;
  wire G139_p_spl_;
  wire G139_p_spl_0;
  wire G139_p_spl_1;
  wire G140_n_spl_;
  wire G140_n_spl_0;
  wire G139_n_spl_;
  wire G139_n_spl_0;
  wire g159_n_spl_;
  wire g158_n_spl_;
  wire G121_n_spl_;
  wire G115_n_spl_;
  wire G115_n_spl_0;
  wire G115_n_spl_1;
  wire g164_n_spl_;
  wire g164_n_spl_0;
  wire G53_n_spl_;
  wire G43_n_spl_;
  wire G96_n_spl_;
  wire G86_n_spl_;
  wire G64_n_spl_;
  wire G32_n_spl_;
  wire G106_n_spl_;
  wire G76_n_spl_;
  wire g172_n_spl_;
  wire g169_n_spl_;
  wire G145_n_spl_;
  wire G145_n_spl_0;
  wire G145_n_spl_00;
  wire G145_n_spl_000;
  wire G145_n_spl_0000;
  wire G145_n_spl_00000;
  wire G145_n_spl_00001;
  wire G145_n_spl_0001;
  wire G145_n_spl_00010;
  wire G145_n_spl_00011;
  wire G145_n_spl_001;
  wire G145_n_spl_0010;
  wire G145_n_spl_0011;
  wire G145_n_spl_01;
  wire G145_n_spl_010;
  wire G145_n_spl_0100;
  wire G145_n_spl_0101;
  wire G145_n_spl_011;
  wire G145_n_spl_0110;
  wire G145_n_spl_0111;
  wire G145_n_spl_1;
  wire G145_n_spl_10;
  wire G145_n_spl_100;
  wire G145_n_spl_1000;
  wire G145_n_spl_1001;
  wire G145_n_spl_101;
  wire G145_n_spl_1010;
  wire G145_n_spl_1011;
  wire G145_n_spl_11;
  wire G145_n_spl_110;
  wire G145_n_spl_1100;
  wire G145_n_spl_1101;
  wire G145_n_spl_111;
  wire G145_n_spl_1110;
  wire G145_n_spl_1111;
  wire G145_p_spl_;
  wire G145_p_spl_0;
  wire G145_p_spl_00;
  wire G145_p_spl_000;
  wire G145_p_spl_0000;
  wire G145_p_spl_00000;
  wire G145_p_spl_00001;
  wire G145_p_spl_0001;
  wire G145_p_spl_00010;
  wire G145_p_spl_00011;
  wire G145_p_spl_001;
  wire G145_p_spl_0010;
  wire G145_p_spl_0011;
  wire G145_p_spl_01;
  wire G145_p_spl_010;
  wire G145_p_spl_0100;
  wire G145_p_spl_0101;
  wire G145_p_spl_011;
  wire G145_p_spl_0110;
  wire G145_p_spl_0111;
  wire G145_p_spl_1;
  wire G145_p_spl_10;
  wire G145_p_spl_100;
  wire G145_p_spl_1000;
  wire G145_p_spl_1001;
  wire G145_p_spl_101;
  wire G145_p_spl_1010;
  wire G145_p_spl_1011;
  wire G145_p_spl_11;
  wire G145_p_spl_110;
  wire G145_p_spl_1100;
  wire G145_p_spl_1101;
  wire G145_p_spl_111;
  wire G145_p_spl_1110;
  wire G145_p_spl_1111;
  wire G146_p_spl_;
  wire G146_p_spl_0;
  wire G146_p_spl_00;
  wire G146_p_spl_000;
  wire G146_p_spl_0000;
  wire G146_p_spl_0001;
  wire G146_p_spl_001;
  wire G146_p_spl_01;
  wire G146_p_spl_010;
  wire G146_p_spl_011;
  wire G146_p_spl_1;
  wire G146_p_spl_10;
  wire G146_p_spl_100;
  wire G146_p_spl_101;
  wire G146_p_spl_11;
  wire G146_p_spl_110;
  wire G146_p_spl_111;
  wire G146_n_spl_;
  wire G146_n_spl_0;
  wire G146_n_spl_00;
  wire G146_n_spl_000;
  wire G146_n_spl_0000;
  wire G146_n_spl_0001;
  wire G146_n_spl_001;
  wire G146_n_spl_01;
  wire G146_n_spl_010;
  wire G146_n_spl_011;
  wire G146_n_spl_1;
  wire G146_n_spl_10;
  wire G146_n_spl_100;
  wire G146_n_spl_101;
  wire G146_n_spl_11;
  wire G146_n_spl_110;
  wire G146_n_spl_111;
  wire G120_n_spl_;
  wire G120_n_spl_0;
  wire G120_n_spl_00;
  wire G120_n_spl_000;
  wire G120_n_spl_0000;
  wire G120_n_spl_0001;
  wire G120_n_spl_001;
  wire G120_n_spl_0010;
  wire G120_n_spl_0011;
  wire G120_n_spl_01;
  wire G120_n_spl_010;
  wire G120_n_spl_0100;
  wire G120_n_spl_011;
  wire G120_n_spl_1;
  wire G120_n_spl_10;
  wire G120_n_spl_100;
  wire G120_n_spl_101;
  wire G120_n_spl_11;
  wire G120_n_spl_110;
  wire G120_n_spl_111;
  wire G117_p_spl_;
  wire G117_p_spl_0;
  wire G117_p_spl_00;
  wire G117_p_spl_000;
  wire G117_p_spl_0000;
  wire G117_p_spl_0001;
  wire G117_p_spl_001;
  wire G117_p_spl_0010;
  wire G117_p_spl_0011;
  wire G117_p_spl_01;
  wire G117_p_spl_010;
  wire G117_p_spl_0100;
  wire G117_p_spl_0101;
  wire G117_p_spl_011;
  wire G117_p_spl_0110;
  wire G117_p_spl_0111;
  wire G117_p_spl_1;
  wire G117_p_spl_10;
  wire G117_p_spl_100;
  wire G117_p_spl_1000;
  wire G117_p_spl_1001;
  wire G117_p_spl_101;
  wire G117_p_spl_1010;
  wire G117_p_spl_1011;
  wire G117_p_spl_11;
  wire G117_p_spl_110;
  wire G117_p_spl_1100;
  wire G117_p_spl_1101;
  wire G117_p_spl_111;
  wire G117_p_spl_1110;
  wire G120_p_spl_;
  wire G120_p_spl_0;
  wire G120_p_spl_00;
  wire G120_p_spl_000;
  wire G120_p_spl_0000;
  wire G120_p_spl_0001;
  wire G120_p_spl_001;
  wire G120_p_spl_0010;
  wire G120_p_spl_0011;
  wire G120_p_spl_01;
  wire G120_p_spl_010;
  wire G120_p_spl_0100;
  wire G120_p_spl_011;
  wire G120_p_spl_1;
  wire G120_p_spl_10;
  wire G120_p_spl_100;
  wire G120_p_spl_101;
  wire G120_p_spl_11;
  wire G120_p_spl_110;
  wire G120_p_spl_111;
  wire G117_n_spl_;
  wire G117_n_spl_0;
  wire G117_n_spl_00;
  wire G117_n_spl_000;
  wire G117_n_spl_0000;
  wire G117_n_spl_0001;
  wire G117_n_spl_001;
  wire G117_n_spl_0010;
  wire G117_n_spl_0011;
  wire G117_n_spl_01;
  wire G117_n_spl_010;
  wire G117_n_spl_0100;
  wire G117_n_spl_0101;
  wire G117_n_spl_011;
  wire G117_n_spl_0110;
  wire G117_n_spl_0111;
  wire G117_n_spl_1;
  wire G117_n_spl_10;
  wire G117_n_spl_100;
  wire G117_n_spl_1000;
  wire G117_n_spl_1001;
  wire G117_n_spl_101;
  wire G117_n_spl_1010;
  wire G117_n_spl_1011;
  wire G117_n_spl_11;
  wire G117_n_spl_110;
  wire G117_n_spl_1100;
  wire G117_n_spl_1101;
  wire G117_n_spl_111;
  wire G117_n_spl_1110;
  wire g204_p_spl_;
  wire g204_p_spl_0;
  wire g204_p_spl_00;
  wire g204_p_spl_000;
  wire g204_p_spl_01;
  wire g204_p_spl_1;
  wire g204_p_spl_10;
  wire g204_p_spl_11;
  wire g204_n_spl_;
  wire g204_n_spl_0;
  wire g204_n_spl_00;
  wire g204_n_spl_000;
  wire g204_n_spl_01;
  wire g204_n_spl_1;
  wire g204_n_spl_10;
  wire g204_n_spl_11;
  wire g240_n_spl_;
  wire g240_n_spl_0;
  wire g240_n_spl_00;
  wire g240_n_spl_1;
  wire G122_n_spl_;
  wire G122_n_spl_0;
  wire g176_n_spl_;
  wire g176_n_spl_0;
  wire g243_n_spl_;
  wire g231_n_spl_;
  wire g231_n_spl_0;
  wire g231_n_spl_00;
  wire g231_n_spl_1;
  wire G123_p_spl_;
  wire G123_p_spl_0;
  wire G123_p_spl_1;
  wire g290_p_spl_;
  wire g290_p_spl_0;
  wire g290_p_spl_00;
  wire g290_p_spl_01;
  wire g290_p_spl_1;
  wire G123_n_spl_;
  wire G123_n_spl_0;
  wire G123_n_spl_1;
  wire g222_p_spl_;
  wire g222_p_spl_0;
  wire g222_p_spl_00;
  wire g222_p_spl_01;
  wire g222_p_spl_1;
  wire g255_n_spl_;
  wire g255_n_spl_0;
  wire g255_n_spl_00;
  wire g255_n_spl_1;
  wire G118_p_spl_;
  wire G118_p_spl_0;
  wire g290_n_spl_;
  wire g290_n_spl_0;
  wire g290_n_spl_00;
  wire g290_n_spl_01;
  wire g290_n_spl_1;
  wire g290_n_spl_10;
  wire g290_n_spl_11;
  wire G118_n_spl_;
  wire g298_p_spl_;
  wire g298_p_spl_0;
  wire g240_p_spl_;
  wire g240_p_spl_0;
  wire g240_p_spl_1;
  wire g310_p_spl_;
  wire g310_p_spl_0;
  wire G143_n_spl_;
  wire G143_n_spl_0;
  wire g310_n_spl_;
  wire g310_n_spl_0;
  wire g310_n_spl_1;
  wire G143_p_spl_;
  wire G143_p_spl_0;
  wire G144_p_spl_;
  wire G144_p_spl_0;
  wire G155_n_spl_;
  wire G154_n_spl_;
  wire G155_p_spl_;
  wire G154_p_spl_;
  wire G126_n_spl_;
  wire G126_n_spl_0;
  wire G125_n_spl_;
  wire G125_n_spl_0;
  wire G126_p_spl_;
  wire G126_p_spl_0;
  wire G126_p_spl_1;
  wire G125_p_spl_;
  wire G125_p_spl_0;
  wire G125_p_spl_1;
  wire g320_n_spl_;
  wire g317_p_spl_;
  wire g320_p_spl_;
  wire g317_n_spl_;
  wire G153_n_spl_;
  wire G152_n_spl_;
  wire G153_p_spl_;
  wire G152_p_spl_;
  wire G149_n_spl_;
  wire G148_n_spl_;
  wire G149_p_spl_;
  wire G148_p_spl_;
  wire g329_n_spl_;
  wire g326_n_spl_;
  wire g329_p_spl_;
  wire g326_p_spl_;
  wire G151_n_spl_;
  wire G150_n_spl_;
  wire G151_p_spl_;
  wire G150_p_spl_;
  wire g335_n_spl_;
  wire g332_n_spl_;
  wire g335_p_spl_;
  wire g332_p_spl_;
  wire G157_n_spl_;
  wire G138_p_spl_;
  wire G138_p_spl_0;
  wire G138_p_spl_00;
  wire G138_p_spl_1;
  wire G157_p_spl_;
  wire G138_n_spl_;
  wire G138_n_spl_0;
  wire G138_n_spl_1;
  wire g349_n_spl_;
  wire g346_n_spl_;
  wire g349_p_spl_;
  wire g346_p_spl_;
  wire g352_n_spl_;
  wire g344_n_spl_;
  wire g352_p_spl_;
  wire g344_p_spl_;
  wire G144_n_spl_;
  wire G134_n_spl_;
  wire G134_n_spl_0;
  wire G134_n_spl_1;
  wire G133_n_spl_;
  wire G133_n_spl_0;
  wire G134_p_spl_;
  wire G134_p_spl_0;
  wire G134_p_spl_1;
  wire G133_p_spl_;
  wire G133_p_spl_0;
  wire G133_p_spl_1;
  wire G136_n_spl_;
  wire G136_n_spl_0;
  wire G136_n_spl_1;
  wire G135_n_spl_;
  wire G135_n_spl_0;
  wire G135_n_spl_1;
  wire G136_p_spl_;
  wire G136_p_spl_0;
  wire G136_p_spl_00;
  wire G136_p_spl_1;
  wire G135_p_spl_;
  wire G135_p_spl_0;
  wire G135_p_spl_1;
  wire g367_n_spl_;
  wire g364_p_spl_;
  wire g367_p_spl_;
  wire g364_n_spl_;
  wire G132_n_spl_;
  wire G132_n_spl_0;
  wire G131_n_spl_;
  wire G131_n_spl_0;
  wire G132_p_spl_;
  wire G132_p_spl_0;
  wire G132_p_spl_1;
  wire G131_p_spl_;
  wire G131_p_spl_0;
  wire G131_p_spl_1;
  wire G156_n_spl_;
  wire G128_p_spl_;
  wire G128_p_spl_0;
  wire G128_p_spl_1;
  wire G156_p_spl_;
  wire G128_n_spl_;
  wire G128_n_spl_0;
  wire g376_n_spl_;
  wire g373_n_spl_;
  wire g376_p_spl_;
  wire g373_p_spl_;
  wire G130_n_spl_;
  wire G130_n_spl_0;
  wire G129_n_spl_;
  wire G129_n_spl_0;
  wire G130_p_spl_;
  wire G130_p_spl_0;
  wire G130_p_spl_1;
  wire G129_p_spl_;
  wire G129_p_spl_0;
  wire G129_p_spl_1;
  wire g382_n_spl_;
  wire g379_n_spl_;
  wire g382_p_spl_;
  wire g379_p_spl_;
  wire G12_n_spl_;
  wire G12_n_spl_0;
  wire G12_n_spl_00;
  wire G12_n_spl_000;
  wire G12_n_spl_0000;
  wire G12_n_spl_0001;
  wire G12_n_spl_001;
  wire G12_n_spl_01;
  wire G12_n_spl_010;
  wire G12_n_spl_011;
  wire G12_n_spl_1;
  wire G12_n_spl_10;
  wire G12_n_spl_100;
  wire G12_n_spl_101;
  wire G12_n_spl_11;
  wire G12_n_spl_110;
  wire G12_n_spl_111;
  wire g222_n_spl_;
  wire g222_n_spl_0;
  wire g222_n_spl_1;
  wire G12_p_spl_;
  wire G12_p_spl_0;
  wire G12_p_spl_00;
  wire G12_p_spl_000;
  wire G12_p_spl_0000;
  wire G12_p_spl_0001;
  wire G12_p_spl_001;
  wire G12_p_spl_01;
  wire G12_p_spl_010;
  wire G12_p_spl_011;
  wire G12_p_spl_1;
  wire G12_p_spl_10;
  wire G12_p_spl_100;
  wire G12_p_spl_101;
  wire G12_p_spl_11;
  wire G12_p_spl_110;
  wire G12_p_spl_111;
  wire g231_p_spl_;
  wire g231_p_spl_0;
  wire g231_p_spl_00;
  wire g231_p_spl_01;
  wire g231_p_spl_1;
  wire g213_p_spl_;
  wire g213_p_spl_0;
  wire g213_p_spl_00;
  wire g213_p_spl_1;
  wire g213_n_spl_;
  wire g213_n_spl_0;
  wire g213_n_spl_1;
  wire G23_n_spl_;
  wire G23_n_spl_0;
  wire G23_n_spl_00;
  wire G23_n_spl_000;
  wire G23_n_spl_001;
  wire G23_n_spl_01;
  wire G23_n_spl_010;
  wire G23_n_spl_011;
  wire G23_n_spl_1;
  wire G23_n_spl_10;
  wire G23_n_spl_100;
  wire G23_n_spl_101;
  wire G23_n_spl_11;
  wire G23_n_spl_110;
  wire G23_p_spl_;
  wire G23_p_spl_0;
  wire G23_p_spl_00;
  wire G23_p_spl_000;
  wire G23_p_spl_001;
  wire G23_p_spl_01;
  wire G23_p_spl_010;
  wire G23_p_spl_011;
  wire G23_p_spl_1;
  wire G23_p_spl_10;
  wire G23_p_spl_100;
  wire G23_p_spl_101;
  wire G23_p_spl_11;
  wire G23_p_spl_110;
  wire g185_n_spl_;
  wire g185_n_spl_0;
  wire g185_n_spl_00;
  wire g185_n_spl_1;
  wire g185_p_spl_;
  wire g185_p_spl_0;
  wire g185_p_spl_1;
  wire g203_n_spl_;
  wire g203_n_spl_0;
  wire g203_n_spl_00;
  wire g203_n_spl_1;
  wire g203_p_spl_;
  wire g203_p_spl_0;
  wire g203_p_spl_1;
  wire g427_n_spl_;
  wire g427_n_spl_0;
  wire g427_n_spl_1;
  wire g427_p_spl_;
  wire g427_p_spl_0;
  wire g427_p_spl_1;
  wire g255_p_spl_;
  wire g255_p_spl_0;
  wire g255_p_spl_00;
  wire g255_p_spl_1;
  wire g262_n_spl_;
  wire g262_n_spl_0;
  wire g262_n_spl_1;
  wire g262_p_spl_;
  wire g262_p_spl_0;
  wire g262_p_spl_1;
  wire g271_p_spl_;
  wire g271_p_spl_0;
  wire g271_p_spl_1;
  wire g271_n_spl_;
  wire g271_n_spl_0;
  wire g271_n_spl_1;
  wire g280_p_spl_;
  wire g280_p_spl_0;
  wire g280_p_spl_1;
  wire g280_n_spl_;
  wire g280_n_spl_0;
  wire g280_n_spl_00;
  wire g280_n_spl_1;
  wire g484_n_spl_;
  wire g484_n_spl_0;
  wire g484_n_spl_1;
  wire g484_p_spl_;
  wire g484_p_spl_0;
  wire g484_p_spl_1;
  wire g503_n_spl_;
  wire g503_n_spl_0;
  wire g503_p_spl_;
  wire g503_p_spl_0;
  wire g194_n_spl_;
  wire g194_n_spl_0;
  wire g194_n_spl_1;
  wire g194_p_spl_;
  wire g194_p_spl_0;
  wire g522_n_spl_;
  wire g522_n_spl_0;
  wire g522_n_spl_1;
  wire g522_p_spl_;
  wire g522_p_spl_0;
  wire g522_p_spl_1;
  wire g550_n_spl_;
  wire g550_n_spl_0;
  wire g550_n_spl_1;
  wire g550_p_spl_;
  wire g553_n_spl_;
  wire g553_n_spl_0;
  wire g553_p_spl_;
  wire g553_p_spl_0;
  wire g562_p_spl_;
  wire g562_n_spl_;
  wire g574_p_spl_;
  wire g574_n_spl_;
  wire g580_n_spl_;
  wire g577_p_spl_;
  wire g580_p_spl_;
  wire g577_n_spl_;
  wire g586_n_spl_;
  wire g583_n_spl_;
  wire g586_p_spl_;
  wire g583_p_spl_;
  wire G29_n_spl_;
  wire g600_n_spl_;
  wire g597_p_spl_;
  wire g600_p_spl_;
  wire g597_n_spl_;
  wire g606_n_spl_;
  wire g606_p_spl_;
  wire g609_n_spl_;
  wire g609_n_spl_0;
  wire g609_n_spl_1;
  wire g609_p_spl_;
  wire g609_p_spl_0;
  wire g609_p_spl_1;
  wire g298_n_spl_;
  wire g603_p_spl_;
  wire g603_n_spl_;
  wire g620_p_spl_;
  wire g620_n_spl_;
  wire g629_p_spl_;
  wire g628_p_spl_;
  wire g629_n_spl_;
  wire g628_n_spl_;
  wire g630_p_spl_;
  wire g630_p_spl_0;
  wire g630_p_spl_00;
  wire g630_p_spl_01;
  wire g630_p_spl_1;
  wire G8_n_spl_;
  wire g631_n_spl_;
  wire g631_n_spl_0;
  wire g631_n_spl_1;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire g630_n_spl_;
  wire g630_n_spl_0;
  wire g630_n_spl_00;
  wire g630_n_spl_1;
  wire g633_p_spl_;
  wire g633_n_spl_;
  wire g640_p_spl_;
  wire g637_p_spl_;
  wire g646_p_spl_;
  wire g643_p_spl_;
  wire g651_n_spl_;
  wire g656_n_spl_;
  wire g661_n_spl_;
  wire g682_p_spl_;
  wire g682_p_spl_0;
  wire g682_p_spl_00;
  wire g682_p_spl_01;
  wire g682_p_spl_1;
  wire g682_p_spl_10;
  wire g682_p_spl_11;
  wire g682_n_spl_;
  wire g682_n_spl_0;
  wire g682_n_spl_00;
  wire g682_n_spl_01;
  wire g682_n_spl_1;
  wire g682_n_spl_10;
  wire g682_n_spl_11;
  wire g684_p_spl_;
  wire g683_n_spl_;
  wire g687_p_spl_;
  wire g686_n_spl_;
  wire g690_n_spl_;
  wire g695_p_spl_;
  wire g694_n_spl_;
  wire g700_n_spl_;
  wire g699_p_spl_;
  wire g698_n_spl_;
  wire g693_n_spl_;
  wire g361_p_spl_;
  wire g342_p_spl_;
  wire g388_p_spl_;
  wire g593_p_spl_;
  wire g627_p_spl_;
  wire G124_n_spl_;
  wire G137_n_spl_;
  wire G137_n_spl_0;
  wire g173_n_spl_;
  wire g292_n_spl_;
  wire g295_n_spl_;
  wire g301_n_spl_;
  wire g540_n_spl_;
  wire g617_p_spl_;
  wire g718_n_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    G37_p,
    G37
  );


  not

  (
    G37_n,
    G37
  );


  buf

  (
    G38_p,
    G38
  );


  not

  (
    G38_n,
    G38
  );


  buf

  (
    G39_p,
    G39
  );


  not

  (
    G39_n,
    G39
  );


  buf

  (
    G40_p,
    G40
  );


  not

  (
    G40_n,
    G40
  );


  buf

  (
    G41_p,
    G41
  );


  not

  (
    G41_n,
    G41
  );


  buf

  (
    G42_p,
    G42
  );


  not

  (
    G42_n,
    G42
  );


  buf

  (
    G43_p,
    G43
  );


  not

  (
    G43_n,
    G43
  );


  buf

  (
    G44_p,
    G44
  );


  not

  (
    G44_n,
    G44
  );


  buf

  (
    G45_p,
    G45
  );


  not

  (
    G45_n,
    G45
  );


  buf

  (
    G46_p,
    G46
  );


  not

  (
    G46_n,
    G46
  );


  buf

  (
    G47_p,
    G47
  );


  not

  (
    G47_n,
    G47
  );


  buf

  (
    G48_p,
    G48
  );


  not

  (
    G48_n,
    G48
  );


  buf

  (
    G49_p,
    G49
  );


  not

  (
    G49_n,
    G49
  );


  buf

  (
    G50_p,
    G50
  );


  not

  (
    G50_n,
    G50
  );


  buf

  (
    G51_p,
    G51
  );


  not

  (
    G51_n,
    G51
  );


  buf

  (
    G52_p,
    G52
  );


  not

  (
    G52_n,
    G52
  );


  buf

  (
    G53_p,
    G53
  );


  not

  (
    G53_n,
    G53
  );


  buf

  (
    G54_p,
    G54
  );


  not

  (
    G54_n,
    G54
  );


  buf

  (
    G55_p,
    G55
  );


  not

  (
    G55_n,
    G55
  );


  buf

  (
    G56_p,
    G56
  );


  not

  (
    G56_n,
    G56
  );


  buf

  (
    G57_p,
    G57
  );


  not

  (
    G57_n,
    G57
  );


  buf

  (
    G58_p,
    G58
  );


  not

  (
    G58_n,
    G58
  );


  buf

  (
    G59_p,
    G59
  );


  not

  (
    G59_n,
    G59
  );


  buf

  (
    G60_p,
    G60
  );


  not

  (
    G60_n,
    G60
  );


  buf

  (
    G61_p,
    G61
  );


  not

  (
    G61_n,
    G61
  );


  buf

  (
    G62_p,
    G62
  );


  not

  (
    G62_n,
    G62
  );


  buf

  (
    G63_p,
    G63
  );


  not

  (
    G63_n,
    G63
  );


  buf

  (
    G64_p,
    G64
  );


  not

  (
    G64_n,
    G64
  );


  buf

  (
    G65_p,
    G65
  );


  not

  (
    G65_n,
    G65
  );


  buf

  (
    G66_p,
    G66
  );


  not

  (
    G66_n,
    G66
  );


  buf

  (
    G67_p,
    G67
  );


  not

  (
    G67_n,
    G67
  );


  buf

  (
    G68_p,
    G68
  );


  not

  (
    G68_n,
    G68
  );


  buf

  (
    G69_p,
    G69
  );


  not

  (
    G69_n,
    G69
  );


  buf

  (
    G70_p,
    G70
  );


  not

  (
    G70_n,
    G70
  );


  buf

  (
    G71_p,
    G71
  );


  not

  (
    G71_n,
    G71
  );


  buf

  (
    G72_p,
    G72
  );


  not

  (
    G72_n,
    G72
  );


  buf

  (
    G73_p,
    G73
  );


  not

  (
    G73_n,
    G73
  );


  buf

  (
    G74_p,
    G74
  );


  not

  (
    G74_n,
    G74
  );


  buf

  (
    G75_p,
    G75
  );


  not

  (
    G75_n,
    G75
  );


  buf

  (
    G76_p,
    G76
  );


  not

  (
    G76_n,
    G76
  );


  buf

  (
    G77_p,
    G77
  );


  not

  (
    G77_n,
    G77
  );


  buf

  (
    G78_p,
    G78
  );


  not

  (
    G78_n,
    G78
  );


  buf

  (
    G79_p,
    G79
  );


  not

  (
    G79_n,
    G79
  );


  buf

  (
    G80_p,
    G80
  );


  not

  (
    G80_n,
    G80
  );


  buf

  (
    G81_p,
    G81
  );


  not

  (
    G81_n,
    G81
  );


  buf

  (
    G82_p,
    G82
  );


  not

  (
    G82_n,
    G82
  );


  buf

  (
    G83_p,
    G83
  );


  not

  (
    G83_n,
    G83
  );


  buf

  (
    G84_p,
    G84
  );


  not

  (
    G84_n,
    G84
  );


  buf

  (
    G85_p,
    G85
  );


  not

  (
    G85_n,
    G85
  );


  buf

  (
    G86_p,
    G86
  );


  not

  (
    G86_n,
    G86
  );


  buf

  (
    G87_p,
    G87
  );


  not

  (
    G87_n,
    G87
  );


  buf

  (
    G88_p,
    G88
  );


  not

  (
    G88_n,
    G88
  );


  buf

  (
    G89_p,
    G89
  );


  not

  (
    G89_n,
    G89
  );


  buf

  (
    G90_p,
    G90
  );


  not

  (
    G90_n,
    G90
  );


  buf

  (
    G91_p,
    G91
  );


  not

  (
    G91_n,
    G91
  );


  buf

  (
    G92_p,
    G92
  );


  not

  (
    G92_n,
    G92
  );


  buf

  (
    G93_p,
    G93
  );


  not

  (
    G93_n,
    G93
  );


  buf

  (
    G94_p,
    G94
  );


  not

  (
    G94_n,
    G94
  );


  buf

  (
    G95_p,
    G95
  );


  not

  (
    G95_n,
    G95
  );


  buf

  (
    G96_p,
    G96
  );


  not

  (
    G96_n,
    G96
  );


  buf

  (
    G97_p,
    G97
  );


  not

  (
    G97_n,
    G97
  );


  buf

  (
    G98_p,
    G98
  );


  not

  (
    G98_n,
    G98
  );


  buf

  (
    G99_p,
    G99
  );


  not

  (
    G99_n,
    G99
  );


  buf

  (
    G100_p,
    G100
  );


  not

  (
    G100_n,
    G100
  );


  buf

  (
    G101_p,
    G101
  );


  not

  (
    G101_n,
    G101
  );


  buf

  (
    G102_p,
    G102
  );


  not

  (
    G102_n,
    G102
  );


  buf

  (
    G103_p,
    G103
  );


  not

  (
    G103_n,
    G103
  );


  buf

  (
    G104_p,
    G104
  );


  not

  (
    G104_n,
    G104
  );


  buf

  (
    G105_p,
    G105
  );


  not

  (
    G105_n,
    G105
  );


  buf

  (
    G106_p,
    G106
  );


  not

  (
    G106_n,
    G106
  );


  buf

  (
    G107_p,
    G107
  );


  not

  (
    G107_n,
    G107
  );


  buf

  (
    G108_p,
    G108
  );


  not

  (
    G108_n,
    G108
  );


  buf

  (
    G109_p,
    G109
  );


  not

  (
    G109_n,
    G109
  );


  buf

  (
    G110_p,
    G110
  );


  not

  (
    G110_n,
    G110
  );


  buf

  (
    G111_p,
    G111
  );


  not

  (
    G111_n,
    G111
  );


  buf

  (
    G112_p,
    G112
  );


  not

  (
    G112_n,
    G112
  );


  buf

  (
    G113_p,
    G113
  );


  not

  (
    G113_n,
    G113
  );


  buf

  (
    G114_p,
    G114
  );


  not

  (
    G114_n,
    G114
  );


  buf

  (
    G115_p,
    G115
  );


  not

  (
    G115_n,
    G115
  );


  buf

  (
    G116_p,
    G116
  );


  not

  (
    G116_n,
    G116
  );


  buf

  (
    G117_p,
    G117
  );


  not

  (
    G117_n,
    G117
  );


  buf

  (
    G118_p,
    G118
  );


  not

  (
    G118_n,
    G118
  );


  buf

  (
    G119_p,
    G119
  );


  not

  (
    G119_n,
    G119
  );


  buf

  (
    G120_p,
    G120
  );


  not

  (
    G120_n,
    G120
  );


  buf

  (
    G121_p,
    G121
  );


  not

  (
    G121_n,
    G121
  );


  buf

  (
    G122_p,
    G122
  );


  not

  (
    G122_n,
    G122
  );


  buf

  (
    G123_p,
    G123
  );


  not

  (
    G123_n,
    G123
  );


  buf

  (
    G124_p,
    G124
  );


  not

  (
    G124_n,
    G124
  );


  buf

  (
    G125_p,
    G125
  );


  not

  (
    G125_n,
    G125
  );


  buf

  (
    G126_p,
    G126
  );


  not

  (
    G126_n,
    G126
  );


  buf

  (
    G127_p,
    G127
  );


  not

  (
    G127_n,
    G127
  );


  buf

  (
    G128_p,
    G128
  );


  not

  (
    G128_n,
    G128
  );


  buf

  (
    G129_p,
    G129
  );


  not

  (
    G129_n,
    G129
  );


  buf

  (
    G130_p,
    G130
  );


  not

  (
    G130_n,
    G130
  );


  buf

  (
    G131_p,
    G131
  );


  not

  (
    G131_n,
    G131
  );


  buf

  (
    G132_p,
    G132
  );


  not

  (
    G132_n,
    G132
  );


  buf

  (
    G133_p,
    G133
  );


  not

  (
    G133_n,
    G133
  );


  buf

  (
    G134_p,
    G134
  );


  not

  (
    G134_n,
    G134
  );


  buf

  (
    G135_p,
    G135
  );


  not

  (
    G135_n,
    G135
  );


  buf

  (
    G136_p,
    G136
  );


  not

  (
    G136_n,
    G136
  );


  buf

  (
    G137_p,
    G137
  );


  not

  (
    G137_n,
    G137
  );


  buf

  (
    G138_p,
    G138
  );


  not

  (
    G138_n,
    G138
  );


  buf

  (
    G139_p,
    G139
  );


  not

  (
    G139_n,
    G139
  );


  buf

  (
    G140_p,
    G140
  );


  not

  (
    G140_n,
    G140
  );


  buf

  (
    G141_p,
    G141
  );


  not

  (
    G141_n,
    G141
  );


  buf

  (
    G142_p,
    G142
  );


  not

  (
    G142_n,
    G142
  );


  buf

  (
    G143_p,
    G143
  );


  not

  (
    G143_n,
    G143
  );


  buf

  (
    G144_p,
    G144
  );


  not

  (
    G144_n,
    G144
  );


  buf

  (
    G145_p,
    G145
  );


  not

  (
    G145_n,
    G145
  );


  buf

  (
    G146_p,
    G146
  );


  not

  (
    G146_n,
    G146
  );


  buf

  (
    G147_p,
    G147
  );


  not

  (
    G147_n,
    G147
  );


  buf

  (
    G148_p,
    G148
  );


  not

  (
    G148_n,
    G148
  );


  buf

  (
    G149_p,
    G149
  );


  not

  (
    G149_n,
    G149
  );


  buf

  (
    G150_p,
    G150
  );


  not

  (
    G150_n,
    G150
  );


  buf

  (
    G151_p,
    G151
  );


  not

  (
    G151_n,
    G151
  );


  buf

  (
    G152_p,
    G152
  );


  not

  (
    G152_n,
    G152
  );


  buf

  (
    G153_p,
    G153
  );


  not

  (
    G153_n,
    G153
  );


  buf

  (
    G154_p,
    G154
  );


  not

  (
    G154_n,
    G154
  );


  buf

  (
    G155_p,
    G155
  );


  not

  (
    G155_n,
    G155
  );


  buf

  (
    G156_p,
    G156
  );


  not

  (
    G156_n,
    G156
  );


  buf

  (
    G157_p,
    G157
  );


  not

  (
    G157_n,
    G157
  );


  and

  (
    g158_p,
    G142_p_spl_0,
    G141_p_spl_0
  );


  or

  (
    g158_n,
    G142_n_spl_0,
    G141_n_spl_0
  );


  and

  (
    g159_p,
    G140_p_spl_0,
    G139_p_spl_0
  );


  or

  (
    g159_n,
    G140_n_spl_0,
    G139_n_spl_0
  );


  or

  (
    g160_n,
    g159_n_spl_,
    g158_n_spl_
  );


  or

  (
    g161_n,
    G121_n_spl_,
    G2_n
  );


  or

  (
    g162_n,
    g161_n,
    G11_n
  );


  and

  (
    g163_p,
    G115_n_spl_0,
    G74_p
  );


  or

  (
    g164_n,
    G121_n_spl_,
    G7_n
  );


  or

  (
    g165_n,
    g164_n_spl_0,
    G119_n
  );


  or

  (
    g166_n,
    g164_n_spl_0,
    G147_n
  );


  or

  (
    g167_n,
    G53_n_spl_,
    G43_n_spl_
  );


  or

  (
    g168_n,
    G96_n_spl_,
    G86_n_spl_
  );


  or

  (
    g169_n,
    g168_n,
    g167_n
  );


  or

  (
    g170_n,
    G64_n_spl_,
    G32_n_spl_
  );


  or

  (
    g171_n,
    G106_n_spl_,
    G76_n_spl_
  );


  or

  (
    g172_n,
    g171_n,
    g170_n
  );


  or

  (
    g173_n,
    g172_n_spl_,
    g169_n_spl_
  );


  and

  (
    g174_p,
    g172_n_spl_,
    G147_p
  );


  and

  (
    g175_p,
    g169_n_spl_,
    G119_p
  );


  or

  (
    g176_n,
    g175_p,
    g174_p
  );


  and

  (
    g177_p,
    G145_n_spl_00000,
    G79_n
  );


  or

  (
    g177_n,
    G145_p_spl_00000,
    G79_p
  );


  and

  (
    g178_p,
    G145_p_spl_00000,
    G109_n
  );


  or

  (
    g178_n,
    G145_n_spl_00000,
    G109_p
  );


  and

  (
    g179_p,
    g178_n,
    g177_n
  );


  or

  (
    g179_n,
    g178_p,
    g177_p
  );


  and

  (
    g180_p,
    g179_n,
    G146_p_spl_0000
  );


  or

  (
    g180_n,
    g179_p,
    G146_n_spl_0000
  );


  and

  (
    g181_p,
    G145_p_spl_00001,
    G99_n
  );


  or

  (
    g181_n,
    G145_n_spl_00001,
    G99_p
  );


  and

  (
    g182_p,
    G145_n_spl_00001,
    G89_n
  );


  or

  (
    g182_n,
    G145_p_spl_00001,
    G89_p
  );


  and

  (
    g183_p,
    g182_n,
    g181_n
  );


  or

  (
    g183_n,
    g182_p,
    g181_p
  );


  and

  (
    g184_p,
    g183_n,
    G146_n_spl_0000
  );


  or

  (
    g184_n,
    g183_p,
    G146_p_spl_0000
  );


  and

  (
    g185_p,
    g184_n,
    g180_n
  );


  or

  (
    g185_n,
    g184_p,
    g180_p
  );


  and

  (
    g186_p,
    G145_n_spl_00010,
    G78_n
  );


  or

  (
    g186_n,
    G145_p_spl_00010,
    G78_p
  );


  and

  (
    g187_p,
    G145_p_spl_00010,
    G108_n
  );


  or

  (
    g187_n,
    G145_n_spl_00010,
    G108_p
  );


  and

  (
    g188_p,
    g187_n,
    g186_n
  );


  or

  (
    g188_n,
    g187_p,
    g186_p
  );


  and

  (
    g189_p,
    g188_n,
    G146_p_spl_0001
  );


  or

  (
    g189_n,
    g188_p,
    G146_n_spl_0001
  );


  and

  (
    g190_p,
    G145_p_spl_00011,
    G98_n
  );


  or

  (
    g190_n,
    G145_n_spl_00011,
    G98_p
  );


  and

  (
    g191_p,
    G145_n_spl_00011,
    G88_n
  );


  or

  (
    g191_n,
    G145_p_spl_00011,
    G88_p
  );


  and

  (
    g192_p,
    g191_n,
    g190_n
  );


  or

  (
    g192_n,
    g191_p,
    g190_p
  );


  and

  (
    g193_p,
    g192_n,
    G146_n_spl_0001
  );


  or

  (
    g193_n,
    g192_p,
    G146_p_spl_0001
  );


  and

  (
    g194_p,
    g193_n,
    g189_n
  );


  or

  (
    g194_n,
    g193_p,
    g189_p
  );


  and

  (
    g195_p,
    G145_n_spl_0010,
    G80_n
  );


  or

  (
    g195_n,
    G145_p_spl_0010,
    G80_p
  );


  and

  (
    g196_p,
    G145_p_spl_0010,
    G110_n
  );


  or

  (
    g196_n,
    G145_n_spl_0010,
    G110_p
  );


  and

  (
    g197_p,
    g196_n,
    g195_n
  );


  or

  (
    g197_n,
    g196_p,
    g195_p
  );


  and

  (
    g198_p,
    g197_n,
    G146_p_spl_001
  );


  or

  (
    g198_n,
    g197_p,
    G146_n_spl_001
  );


  and

  (
    g199_p,
    G145_p_spl_0011,
    G100_n
  );


  or

  (
    g199_n,
    G145_n_spl_0011,
    G100_p
  );


  and

  (
    g200_p,
    G145_n_spl_0011,
    G90_n
  );


  or

  (
    g200_n,
    G145_p_spl_0011,
    G90_p
  );


  and

  (
    g201_p,
    g200_n,
    g199_n
  );


  or

  (
    g201_n,
    g200_p,
    g199_p
  );


  and

  (
    g202_p,
    g201_n,
    G146_n_spl_001
  );


  or

  (
    g202_n,
    g201_p,
    G146_p_spl_001
  );


  and

  (
    g203_p,
    g202_n,
    g198_n
  );


  or

  (
    g203_n,
    g202_p,
    g198_p
  );


  and

  (
    g204_p,
    G120_n_spl_0000,
    G117_p_spl_0000
  );


  or

  (
    g204_n,
    G120_p_spl_0000,
    G117_n_spl_0000
  );


  and

  (
    g205_p,
    g204_p_spl_000,
    G46_p
  );


  or

  (
    g205_n,
    g204_n_spl_000,
    G46_n
  );


  and

  (
    g206_p,
    G117_n_spl_0000,
    G57_p
  );


  or

  (
    g206_n,
    G117_p_spl_0000,
    G57_n
  );


  and

  (
    g207_p,
    g206_n,
    G120_n_spl_0000
  );


  or

  (
    g207_n,
    g206_p,
    G120_p_spl_0000
  );


  and

  (
    g208_p,
    G117_n_spl_0001,
    G36_n
  );


  or

  (
    g208_n,
    G117_p_spl_0001,
    G36_p
  );


  and

  (
    g209_p,
    g208_p,
    G120_p_spl_0001
  );


  or

  (
    g209_n,
    g208_n,
    G120_n_spl_0001
  );


  and

  (
    g210_p,
    G117_p_spl_0001,
    G68_n
  );


  or

  (
    g210_n,
    G117_n_spl_0001,
    G68_p
  );


  and

  (
    g211_p,
    g210_n,
    g209_n
  );


  or

  (
    g211_n,
    g210_p,
    g209_p
  );


  and

  (
    g212_p,
    g211_p,
    g207_n
  );


  or

  (
    g212_n,
    g211_n,
    g207_p
  );


  and

  (
    g213_p,
    g212_n,
    g205_n
  );


  or

  (
    g213_n,
    g212_p,
    g205_p
  );


  and

  (
    g214_p,
    g204_p_spl_000,
    G47_p
  );


  or

  (
    g214_n,
    g204_n_spl_000,
    G47_n
  );


  and

  (
    g215_p,
    G117_n_spl_0010,
    G58_p
  );


  or

  (
    g215_n,
    G117_p_spl_0010,
    G58_n
  );


  and

  (
    g216_p,
    g215_n,
    G120_n_spl_0001
  );


  or

  (
    g216_n,
    g215_p,
    G120_p_spl_0001
  );


  and

  (
    g217_p,
    G117_n_spl_0010,
    G37_n
  );


  or

  (
    g217_n,
    G117_p_spl_0010,
    G37_p
  );


  and

  (
    g218_p,
    g217_p,
    G120_p_spl_0010
  );


  or

  (
    g218_n,
    g217_n,
    G120_n_spl_0010
  );


  and

  (
    g219_p,
    G117_p_spl_0011,
    G69_n
  );


  or

  (
    g219_n,
    G117_n_spl_0011,
    G69_p
  );


  and

  (
    g220_p,
    g219_n,
    g218_n
  );


  or

  (
    g220_n,
    g219_p,
    g218_p
  );


  and

  (
    g221_p,
    g220_p,
    g216_n
  );


  or

  (
    g221_n,
    g220_n,
    g216_p
  );


  and

  (
    g222_p,
    g221_n,
    g214_n
  );


  or

  (
    g222_n,
    g221_p,
    g214_p
  );


  and

  (
    g223_p,
    g204_p_spl_00,
    G48_p
  );


  or

  (
    g223_n,
    g204_n_spl_00,
    G48_n
  );


  and

  (
    g224_p,
    G117_n_spl_0011,
    G59_p
  );


  or

  (
    g224_n,
    G117_p_spl_0011,
    G59_n
  );


  and

  (
    g225_p,
    g224_n,
    G120_n_spl_0010
  );


  or

  (
    g225_n,
    g224_p,
    G120_p_spl_0010
  );


  and

  (
    g226_p,
    G117_n_spl_0100,
    G38_n
  );


  or

  (
    g226_n,
    G117_p_spl_0100,
    G38_p
  );


  and

  (
    g227_p,
    g226_p,
    G120_p_spl_0011
  );


  or

  (
    g227_n,
    g226_n,
    G120_n_spl_0011
  );


  and

  (
    g228_p,
    G117_p_spl_0100,
    G70_n
  );


  or

  (
    g228_n,
    G117_n_spl_0100,
    G70_p
  );


  and

  (
    g229_p,
    g228_n,
    g227_n
  );


  or

  (
    g229_n,
    g228_p,
    g227_p
  );


  and

  (
    g230_p,
    g229_p,
    g225_n
  );


  or

  (
    g230_n,
    g229_n,
    g225_p
  );


  and

  (
    g231_p,
    g230_n,
    g223_n
  );


  or

  (
    g231_n,
    g230_p,
    g223_p
  );


  and

  (
    g232_p,
    g204_p_spl_01,
    G42_p
  );


  or

  (
    g232_n,
    g204_n_spl_01,
    G42_n
  );


  and

  (
    g233_p,
    G117_n_spl_0101,
    G52_p
  );


  or

  (
    g233_n,
    G117_p_spl_0101,
    G52_n
  );


  and

  (
    g234_p,
    g233_n,
    G120_n_spl_0011
  );


  or

  (
    g234_n,
    g233_p,
    G120_p_spl_0011
  );


  and

  (
    g235_p,
    G117_n_spl_0101,
    G31_n
  );


  or

  (
    g235_n,
    G117_p_spl_0101,
    G31_p
  );


  and

  (
    g236_p,
    g235_p,
    G120_p_spl_0100
  );


  or

  (
    g236_n,
    g235_n,
    G120_n_spl_0100
  );


  and

  (
    g237_p,
    G117_p_spl_0110,
    G63_n
  );


  or

  (
    g237_n,
    G117_n_spl_0110,
    G63_p
  );


  and

  (
    g238_p,
    g237_n,
    g236_n
  );


  or

  (
    g238_n,
    g237_p,
    g236_p
  );


  and

  (
    g239_p,
    g238_p,
    g234_n
  );


  or

  (
    g239_n,
    g238_n,
    g234_p
  );


  and

  (
    g240_p,
    g239_n,
    g232_n
  );


  or

  (
    g240_n,
    g239_p,
    g232_p
  );


  or

  (
    g241_n,
    g240_n_spl_00,
    G122_n_spl_0
  );


  or

  (
    g242_n,
    g176_n_spl_0,
    G116_n
  );


  or

  (
    g243_n,
    g242_n,
    G121_p
  );


  or

  (
    g244_n,
    g243_n_spl_,
    G28_n
  );


  and

  (
    g245_p,
    G3_p,
    G1_p
  );


  or

  (
    g246_n,
    g245_p,
    g243_n_spl_
  );


  and

  (
    g247_p,
    g204_p_spl_01,
    G49_p
  );


  or

  (
    g247_n,
    g204_n_spl_01,
    G49_n
  );


  and

  (
    g248_p,
    G117_n_spl_0110,
    G60_p
  );


  or

  (
    g248_n,
    G117_p_spl_0110,
    G60_n
  );


  and

  (
    g249_p,
    g248_n,
    G120_n_spl_0100
  );


  or

  (
    g249_n,
    g248_p,
    G120_p_spl_0100
  );


  and

  (
    g250_p,
    G117_n_spl_0111,
    G39_n
  );


  or

  (
    g250_n,
    G117_p_spl_0111,
    G39_p
  );


  and

  (
    g251_p,
    g250_p,
    G120_p_spl_010
  );


  or

  (
    g251_n,
    g250_n,
    G120_n_spl_010
  );


  and

  (
    g252_p,
    G117_p_spl_0111,
    G71_n
  );


  or

  (
    g252_n,
    G117_n_spl_0111,
    G71_p
  );


  and

  (
    g253_p,
    g252_n,
    g251_n
  );


  or

  (
    g253_n,
    g252_p,
    g251_p
  );


  and

  (
    g254_p,
    g253_p,
    g249_n
  );


  or

  (
    g254_n,
    g253_n,
    g249_p
  );


  and

  (
    g255_p,
    g254_n,
    g247_n
  );


  or

  (
    g255_n,
    g254_p,
    g247_p
  );


  and

  (
    g256_p,
    G117_n_spl_1000,
    G35_n
  );


  or

  (
    g256_n,
    G117_p_spl_1000,
    G35_p
  );


  and

  (
    g257_p,
    G117_p_spl_1000,
    G67_n
  );


  or

  (
    g257_n,
    G117_n_spl_1000,
    G67_p
  );


  and

  (
    g258_p,
    g257_n,
    g256_n
  );


  or

  (
    g258_n,
    g257_p,
    g256_p
  );


  and

  (
    g259_p,
    g258_n,
    G120_p_spl_011
  );


  or

  (
    g259_n,
    g258_p,
    G120_n_spl_011
  );


  and

  (
    g260_p,
    G117_n_spl_1001,
    G56_n
  );


  or

  (
    g260_n,
    G117_p_spl_1001,
    G56_p
  );


  and

  (
    g261_p,
    g260_p,
    G120_n_spl_011
  );


  or

  (
    g261_n,
    g260_n,
    G120_p_spl_011
  );


  and

  (
    g262_p,
    g261_n,
    g259_n
  );


  or

  (
    g262_n,
    g261_p,
    g259_p
  );


  and

  (
    g263_p,
    g204_p_spl_10,
    G45_p
  );


  or

  (
    g263_n,
    g204_n_spl_10,
    G45_n
  );


  and

  (
    g264_p,
    G117_n_spl_1001,
    G55_p
  );


  or

  (
    g264_n,
    G117_p_spl_1001,
    G55_n
  );


  and

  (
    g265_p,
    g264_n,
    G120_n_spl_100
  );


  or

  (
    g265_n,
    g264_p,
    G120_p_spl_100
  );


  and

  (
    g266_p,
    G117_n_spl_1010,
    G34_n
  );


  or

  (
    g266_n,
    G117_p_spl_1010,
    G34_p
  );


  and

  (
    g267_p,
    g266_p,
    G120_p_spl_100
  );


  or

  (
    g267_n,
    g266_n,
    G120_n_spl_100
  );


  and

  (
    g268_p,
    G117_p_spl_1010,
    G66_n
  );


  or

  (
    g268_n,
    G117_n_spl_1010,
    G66_p
  );


  and

  (
    g269_p,
    g268_n,
    g267_n
  );


  or

  (
    g269_n,
    g268_p,
    g267_p
  );


  and

  (
    g270_p,
    g269_p,
    g265_n
  );


  or

  (
    g270_n,
    g269_n,
    g265_p
  );


  and

  (
    g271_p,
    g270_n,
    g263_n
  );


  or

  (
    g271_n,
    g270_p,
    g263_p
  );


  and

  (
    g272_p,
    g204_p_spl_10,
    G44_p
  );


  or

  (
    g272_n,
    g204_n_spl_10,
    G44_n
  );


  and

  (
    g273_p,
    G117_n_spl_1011,
    G54_p
  );


  or

  (
    g273_n,
    G117_p_spl_1011,
    G54_n
  );


  and

  (
    g274_p,
    g273_n,
    G120_n_spl_101
  );


  or

  (
    g274_n,
    g273_p,
    G120_p_spl_101
  );


  and

  (
    g275_p,
    G117_n_spl_1011,
    G33_n
  );


  or

  (
    g275_n,
    G117_p_spl_1011,
    G33_p
  );


  and

  (
    g276_p,
    g275_p,
    G120_p_spl_101
  );


  or

  (
    g276_n,
    g275_n,
    G120_n_spl_101
  );


  and

  (
    g277_p,
    G117_p_spl_1100,
    G65_n
  );


  or

  (
    g277_n,
    G117_n_spl_1100,
    G65_p
  );


  and

  (
    g278_p,
    g277_n,
    g276_n
  );


  or

  (
    g278_n,
    g277_p,
    g276_p
  );


  and

  (
    g279_p,
    g278_p,
    g274_n
  );


  or

  (
    g279_n,
    g278_n,
    g274_p
  );


  and

  (
    g280_p,
    g279_n,
    g272_n
  );


  or

  (
    g280_n,
    g279_p,
    g272_p
  );


  and

  (
    g281_p,
    g231_n_spl_00,
    G123_p_spl_0
  );


  and

  (
    g282_p,
    g204_p_spl_11,
    G50_p
  );


  or

  (
    g282_n,
    g204_n_spl_11,
    G50_n
  );


  and

  (
    g283_p,
    G117_n_spl_1100,
    G61_p
  );


  or

  (
    g283_n,
    G117_p_spl_1100,
    G61_n
  );


  and

  (
    g284_p,
    g283_n,
    G120_n_spl_110
  );


  or

  (
    g284_n,
    g283_p,
    G120_p_spl_110
  );


  and

  (
    g285_p,
    G117_n_spl_1101,
    G40_n
  );


  or

  (
    g285_n,
    G117_p_spl_1101,
    G40_p
  );


  and

  (
    g286_p,
    g285_p,
    G120_p_spl_110
  );


  or

  (
    g286_n,
    g285_n,
    G120_n_spl_110
  );


  and

  (
    g287_p,
    G117_p_spl_1101,
    G72_n
  );


  or

  (
    g287_n,
    G117_n_spl_1101,
    G72_p
  );


  and

  (
    g288_p,
    g287_n,
    g286_n
  );


  or

  (
    g288_n,
    g287_p,
    g286_p
  );


  and

  (
    g289_p,
    g288_p,
    g284_n
  );


  or

  (
    g289_n,
    g288_n,
    g284_p
  );


  and

  (
    g290_p,
    g289_n,
    g282_n
  );


  or

  (
    g290_n,
    g289_p,
    g282_p
  );


  and

  (
    g291_p,
    g290_p_spl_00,
    G123_n_spl_0
  );


  or

  (
    g292_n,
    g291_p,
    g281_p
  );


  and

  (
    g293_p,
    g222_p_spl_00,
    G123_p_spl_0
  );


  and

  (
    g294_p,
    g255_n_spl_00,
    G123_n_spl_0
  );


  or

  (
    g295_n,
    g294_p,
    g293_p
  );


  and

  (
    g296_p,
    G122_n_spl_0,
    G118_p_spl_0
  );


  or

  (
    g297_n,
    g296_p,
    g290_n_spl_00
  );


  and

  (
    g298_p,
    g290_p_spl_00,
    G118_n_spl_
  );


  or

  (
    g298_n,
    g290_n_spl_00,
    G118_p_spl_0
  );


  and

  (
    g299_p,
    g298_p_spl_0,
    G123_p_spl_1
  );


  and

  (
    g300_p,
    g240_p_spl_0,
    G123_n_spl_1
  );


  or

  (
    g301_n,
    g300_p,
    g299_p
  );


  and

  (
    g302_p,
    G145_n_spl_0100,
    G77_n
  );


  or

  (
    g302_n,
    G145_p_spl_0100,
    G77_p
  );


  and

  (
    g303_p,
    G145_p_spl_0100,
    G107_n
  );


  or

  (
    g303_n,
    G145_n_spl_0100,
    G107_p
  );


  and

  (
    g304_p,
    g303_n,
    g302_n
  );


  or

  (
    g304_n,
    g303_p,
    g302_p
  );


  and

  (
    g305_p,
    g304_n,
    G146_p_spl_010
  );


  or

  (
    g305_n,
    g304_p,
    G146_n_spl_010
  );


  and

  (
    g306_p,
    G145_p_spl_0101,
    G97_n
  );


  or

  (
    g306_n,
    G145_n_spl_0101,
    G97_p
  );


  and

  (
    g307_p,
    G145_n_spl_0101,
    G87_n
  );


  or

  (
    g307_n,
    G145_p_spl_0101,
    G87_p
  );


  and

  (
    g308_p,
    g307_n,
    g306_n
  );


  or

  (
    g308_n,
    g307_p,
    g306_p
  );


  and

  (
    g309_p,
    g308_n,
    G146_n_spl_010
  );


  or

  (
    g309_n,
    g308_p,
    G146_p_spl_010
  );


  and

  (
    g310_p,
    g309_n,
    g305_n
  );


  or

  (
    g310_n,
    g309_p,
    g305_p
  );


  or

  (
    g311_n,
    g310_p_spl_0,
    G143_n_spl_0
  );


  or

  (
    g312_n,
    g310_n_spl_0,
    G143_p_spl_0
  );


  and

  (
    g313_p,
    g312_n,
    g311_n
  );


  or

  (
    g314_n,
    g313_p,
    G144_p_spl_0
  );


  and

  (
    g315_p,
    G155_n_spl_,
    G154_n_spl_
  );


  or

  (
    g315_n,
    G155_p_spl_,
    G154_p_spl_
  );


  and

  (
    g316_p,
    G155_p_spl_,
    G154_p_spl_
  );


  or

  (
    g316_n,
    G155_n_spl_,
    G154_n_spl_
  );


  and

  (
    g317_p,
    g316_n,
    g315_n
  );


  or

  (
    g317_n,
    g316_p,
    g315_p
  );


  and

  (
    g318_p,
    G126_n_spl_0,
    G125_n_spl_0
  );


  or

  (
    g318_n,
    G126_p_spl_0,
    G125_p_spl_0
  );


  and

  (
    g319_p,
    G126_p_spl_0,
    G125_p_spl_0
  );


  or

  (
    g319_n,
    G126_n_spl_0,
    G125_n_spl_0
  );


  and

  (
    g320_p,
    g319_n,
    g318_n
  );


  or

  (
    g320_n,
    g319_p,
    g318_p
  );


  and

  (
    g321_p,
    g320_n_spl_,
    g317_p_spl_
  );


  or

  (
    g321_n,
    g320_p_spl_,
    g317_n_spl_
  );


  and

  (
    g322_p,
    g320_p_spl_,
    g317_n_spl_
  );


  or

  (
    g322_n,
    g320_n_spl_,
    g317_p_spl_
  );


  and

  (
    g323_p,
    g322_n,
    g321_n
  );


  or

  (
    g323_n,
    g322_p,
    g321_p
  );


  and

  (
    g324_p,
    G153_n_spl_,
    G152_n_spl_
  );


  or

  (
    g324_n,
    G153_p_spl_,
    G152_p_spl_
  );


  and

  (
    g325_p,
    G153_p_spl_,
    G152_p_spl_
  );


  or

  (
    g325_n,
    G153_n_spl_,
    G152_n_spl_
  );


  and

  (
    g326_p,
    g325_n,
    g324_n
  );


  or

  (
    g326_n,
    g325_p,
    g324_p
  );


  and

  (
    g327_p,
    G149_n_spl_,
    G148_n_spl_
  );


  or

  (
    g327_n,
    G149_p_spl_,
    G148_p_spl_
  );


  and

  (
    g328_p,
    G149_p_spl_,
    G148_p_spl_
  );


  or

  (
    g328_n,
    G149_n_spl_,
    G148_n_spl_
  );


  and

  (
    g329_p,
    g328_n,
    g327_n
  );


  or

  (
    g329_n,
    g328_p,
    g327_p
  );


  and

  (
    g330_p,
    g329_n_spl_,
    g326_n_spl_
  );


  or

  (
    g330_n,
    g329_p_spl_,
    g326_p_spl_
  );


  and

  (
    g331_p,
    g329_p_spl_,
    g326_p_spl_
  );


  or

  (
    g331_n,
    g329_n_spl_,
    g326_n_spl_
  );


  and

  (
    g332_p,
    g331_n,
    g330_n
  );


  or

  (
    g332_n,
    g331_p,
    g330_p
  );


  and

  (
    g333_p,
    G151_n_spl_,
    G150_n_spl_
  );


  or

  (
    g333_n,
    G151_p_spl_,
    G150_p_spl_
  );


  and

  (
    g334_p,
    G151_p_spl_,
    G150_p_spl_
  );


  or

  (
    g334_n,
    G151_n_spl_,
    G150_n_spl_
  );


  and

  (
    g335_p,
    g334_n,
    g333_n
  );


  or

  (
    g335_n,
    g334_p,
    g333_p
  );


  and

  (
    g336_p,
    g335_n_spl_,
    g332_n_spl_
  );


  or

  (
    g336_n,
    g335_p_spl_,
    g332_p_spl_
  );


  and

  (
    g337_p,
    g335_p_spl_,
    g332_p_spl_
  );


  or

  (
    g337_n,
    g335_n_spl_,
    g332_n_spl_
  );


  and

  (
    g338_p,
    g337_n,
    g336_n
  );


  or

  (
    g338_n,
    g337_p,
    g336_p
  );


  or

  (
    g339_n,
    g338_p,
    g323_n
  );


  or

  (
    g340_n,
    g338_n,
    g323_p
  );


  and

  (
    g341_p,
    g340_n,
    G10_p
  );


  and

  (
    g342_p,
    g341_p,
    g339_n
  );


  and

  (
    g343_p,
    G142_n_spl_0,
    G141_n_spl_0
  );


  or

  (
    g343_n,
    G142_p_spl_0,
    G141_p_spl_0
  );


  and

  (
    g344_p,
    g343_n,
    g158_n_spl_
  );


  or

  (
    g344_n,
    g343_p,
    g158_p
  );


  and

  (
    g345_p,
    G140_n_spl_0,
    G139_n_spl_0
  );


  or

  (
    g345_n,
    G140_p_spl_0,
    G139_p_spl_0
  );


  and

  (
    g346_p,
    g345_n,
    g159_n_spl_
  );


  or

  (
    g346_n,
    g345_p,
    g159_p
  );


  and

  (
    g347_p,
    G157_n_spl_,
    G138_p_spl_00
  );


  or

  (
    g347_n,
    G157_p_spl_,
    G138_n_spl_0
  );


  and

  (
    g348_p,
    G157_p_spl_,
    G138_n_spl_0
  );


  or

  (
    g348_n,
    G157_n_spl_,
    G138_p_spl_00
  );


  and

  (
    g349_p,
    g348_n,
    g347_n
  );


  or

  (
    g349_n,
    g348_p,
    g347_p
  );


  and

  (
    g350_p,
    g349_n_spl_,
    g346_n_spl_
  );


  or

  (
    g350_n,
    g349_p_spl_,
    g346_p_spl_
  );


  and

  (
    g351_p,
    g349_p_spl_,
    g346_p_spl_
  );


  or

  (
    g351_n,
    g349_n_spl_,
    g346_n_spl_
  );


  and

  (
    g352_p,
    g351_n,
    g350_n
  );


  or

  (
    g352_n,
    g351_p,
    g350_p
  );


  and

  (
    g353_p,
    g352_n_spl_,
    g344_n_spl_
  );


  or

  (
    g353_n,
    g352_p_spl_,
    g344_p_spl_
  );


  and

  (
    g354_p,
    g352_p_spl_,
    g344_p_spl_
  );


  or

  (
    g354_n,
    g352_n_spl_,
    g344_n_spl_
  );


  and

  (
    g355_p,
    g354_n,
    g353_n
  );


  or

  (
    g355_n,
    g354_p,
    g353_p
  );


  and

  (
    g356_p,
    G144_n_spl_,
    G143_n_spl_0
  );


  or

  (
    g356_n,
    G144_p_spl_0,
    G143_p_spl_0
  );


  and

  (
    g357_p,
    G144_p_spl_,
    G143_p_spl_
  );


  or

  (
    g357_n,
    G144_n_spl_,
    G143_n_spl_
  );


  and

  (
    g358_p,
    g357_n,
    g356_n
  );


  or

  (
    g358_n,
    g357_p,
    g356_p
  );


  or

  (
    g359_n,
    g358_n,
    g355_n
  );


  or

  (
    g360_n,
    g358_p,
    g355_p
  );


  and

  (
    g361_p,
    g360_n,
    g359_n
  );


  and

  (
    g362_p,
    G134_n_spl_0,
    G133_n_spl_0
  );


  or

  (
    g362_n,
    G134_p_spl_0,
    G133_p_spl_0
  );


  and

  (
    g363_p,
    G134_p_spl_0,
    G133_p_spl_0
  );


  or

  (
    g363_n,
    G134_n_spl_0,
    G133_n_spl_0
  );


  and

  (
    g364_p,
    g363_n,
    g362_n
  );


  or

  (
    g364_n,
    g363_p,
    g362_p
  );


  and

  (
    g365_p,
    G136_n_spl_0,
    G135_n_spl_0
  );


  or

  (
    g365_n,
    G136_p_spl_00,
    G135_p_spl_0
  );


  and

  (
    g366_p,
    G136_p_spl_00,
    G135_p_spl_0
  );


  or

  (
    g366_n,
    G136_n_spl_0,
    G135_n_spl_0
  );


  and

  (
    g367_p,
    g366_n,
    g365_n
  );


  or

  (
    g367_n,
    g366_p,
    g365_p
  );


  and

  (
    g368_p,
    g367_n_spl_,
    g364_p_spl_
  );


  or

  (
    g368_n,
    g367_p_spl_,
    g364_n_spl_
  );


  and

  (
    g369_p,
    g367_p_spl_,
    g364_n_spl_
  );


  or

  (
    g369_n,
    g367_n_spl_,
    g364_p_spl_
  );


  and

  (
    g370_p,
    g369_n,
    g368_n
  );


  or

  (
    g370_n,
    g369_p,
    g368_p
  );


  and

  (
    g371_p,
    G132_n_spl_0,
    G131_n_spl_0
  );


  or

  (
    g371_n,
    G132_p_spl_0,
    G131_p_spl_0
  );


  and

  (
    g372_p,
    G132_p_spl_0,
    G131_p_spl_0
  );


  or

  (
    g372_n,
    G132_n_spl_0,
    G131_n_spl_0
  );


  and

  (
    g373_p,
    g372_n,
    g371_n
  );


  or

  (
    g373_n,
    g372_p,
    g371_p
  );


  and

  (
    g374_p,
    G156_n_spl_,
    G128_p_spl_0
  );


  or

  (
    g374_n,
    G156_p_spl_,
    G128_n_spl_0
  );


  and

  (
    g375_p,
    G156_p_spl_,
    G128_n_spl_0
  );


  or

  (
    g375_n,
    G156_n_spl_,
    G128_p_spl_0
  );


  and

  (
    g376_p,
    g375_n,
    g374_n
  );


  or

  (
    g376_n,
    g375_p,
    g374_p
  );


  and

  (
    g377_p,
    g376_n_spl_,
    g373_n_spl_
  );


  or

  (
    g377_n,
    g376_p_spl_,
    g373_p_spl_
  );


  and

  (
    g378_p,
    g376_p_spl_,
    g373_p_spl_
  );


  or

  (
    g378_n,
    g376_n_spl_,
    g373_n_spl_
  );


  and

  (
    g379_p,
    g378_n,
    g377_n
  );


  or

  (
    g379_n,
    g378_p,
    g377_p
  );


  and

  (
    g380_p,
    G130_n_spl_0,
    G129_n_spl_0
  );


  or

  (
    g380_n,
    G130_p_spl_0,
    G129_p_spl_0
  );


  and

  (
    g381_p,
    G130_p_spl_0,
    G129_p_spl_0
  );


  or

  (
    g381_n,
    G130_n_spl_0,
    G129_n_spl_0
  );


  and

  (
    g382_p,
    g381_n,
    g380_n
  );


  or

  (
    g382_n,
    g381_p,
    g380_p
  );


  and

  (
    g383_p,
    g382_n_spl_,
    g379_n_spl_
  );


  or

  (
    g383_n,
    g382_p_spl_,
    g379_p_spl_
  );


  and

  (
    g384_p,
    g382_p_spl_,
    g379_p_spl_
  );


  or

  (
    g384_n,
    g382_n_spl_,
    g379_n_spl_
  );


  and

  (
    g385_p,
    g384_n,
    g383_n
  );


  or

  (
    g385_n,
    g384_p,
    g383_p
  );


  or

  (
    g386_n,
    g385_n,
    g370_p
  );


  or

  (
    g387_n,
    g385_p,
    g370_n
  );


  and

  (
    g388_p,
    g387_n,
    g386_n
  );


  and

  (
    g389_p,
    g222_p_spl_00,
    G12_n_spl_0000
  );


  or

  (
    g389_n,
    g222_n_spl_0,
    G12_p_spl_0000
  );


  and

  (
    g390_p,
    G15_n,
    G12_p_spl_0000
  );


  or

  (
    g390_n,
    G15_p,
    G12_n_spl_0000
  );


  and

  (
    g391_p,
    g390_n,
    g389_n
  );


  or

  (
    g391_n,
    g390_p,
    g389_p
  );


  and

  (
    g392_p,
    g391_n,
    G130_p_spl_1
  );


  and

  (
    g393_p,
    g231_p_spl_00,
    G12_n_spl_0001
  );


  or

  (
    g393_n,
    g231_n_spl_00,
    G12_p_spl_0001
  );


  and

  (
    g394_p,
    G12_p_spl_0001,
    G5_n
  );


  or

  (
    g394_n,
    G12_n_spl_0001,
    G5_p
  );


  and

  (
    g395_p,
    g394_n,
    g393_n
  );


  or

  (
    g395_n,
    g394_p,
    g393_p
  );


  and

  (
    g396_p,
    g395_p,
    G129_n_spl_
  );


  or

  (
    g397_n,
    g396_p,
    g392_p
  );


  and

  (
    g398_p,
    g213_p_spl_00,
    G12_n_spl_001
  );


  or

  (
    g398_n,
    g213_n_spl_0,
    G12_p_spl_001
  );


  and

  (
    g399_p,
    G16_n,
    G12_p_spl_001
  );


  or

  (
    g399_n,
    G16_p,
    G12_n_spl_001
  );


  and

  (
    g400_p,
    g399_n,
    g398_n
  );


  or

  (
    g400_n,
    g399_p,
    g398_p
  );


  and

  (
    g401_p,
    g400_p,
    G131_n_spl_
  );


  or

  (
    g402_n,
    G23_n_spl_000,
    G22_n
  );


  or

  (
    g403_n,
    g310_n_spl_0,
    G23_p_spl_000
  );


  and

  (
    g404_p,
    g403_n,
    g402_n
  );


  or

  (
    g405_n,
    g404_p,
    g401_p
  );


  or

  (
    g406_n,
    g405_n,
    G9_n
  );


  and

  (
    g407_p,
    g185_n_spl_00,
    G23_n_spl_000
  );


  or

  (
    g407_n,
    g185_p_spl_0,
    G23_p_spl_000
  );


  and

  (
    g408_p,
    G26_n,
    G23_p_spl_001
  );


  or

  (
    g408_n,
    G26_p,
    G23_n_spl_001
  );


  and

  (
    g409_p,
    g408_n,
    g407_n
  );


  or

  (
    g409_n,
    g408_p,
    g407_p
  );


  and

  (
    g410_p,
    g409_n,
    G141_p_spl_1
  );


  and

  (
    g411_p,
    g203_n_spl_00,
    G23_n_spl_001
  );


  or

  (
    g411_n,
    g203_p_spl_0,
    G23_p_spl_001
  );


  and

  (
    g412_p,
    G23_p_spl_010,
    G21_n
  );


  or

  (
    g412_n,
    G23_n_spl_010,
    G21_p
  );


  and

  (
    g413_p,
    g412_n,
    g411_n
  );


  or

  (
    g413_n,
    g412_p,
    g411_p
  );


  and

  (
    g414_p,
    g413_n,
    G140_p_spl_1
  );


  and

  (
    g415_p,
    g409_p,
    G141_n_spl_
  );


  or

  (
    g416_n,
    g415_p,
    g414_p
  );


  or

  (
    g417_n,
    g416_n,
    g410_p
  );


  and

  (
    g418_p,
    g413_p,
    G140_n_spl_
  );


  and

  (
    g419_p,
    G145_n_spl_0110,
    G83_n
  );


  or

  (
    g419_n,
    G145_p_spl_0110,
    G83_p
  );


  and

  (
    g420_p,
    G145_p_spl_0110,
    G113_n
  );


  or

  (
    g420_n,
    G145_n_spl_0110,
    G113_p
  );


  and

  (
    g421_p,
    g420_n,
    g419_n
  );


  or

  (
    g421_n,
    g420_p,
    g419_p
  );


  and

  (
    g422_p,
    g421_n,
    G146_p_spl_011
  );


  or

  (
    g422_n,
    g421_p,
    G146_n_spl_011
  );


  and

  (
    g423_p,
    G145_p_spl_0111,
    G103_n
  );


  or

  (
    g423_n,
    G145_n_spl_0111,
    G103_p
  );


  and

  (
    g424_p,
    G145_n_spl_0111,
    G93_n
  );


  or

  (
    g424_n,
    G145_p_spl_0111,
    G93_p
  );


  and

  (
    g425_p,
    g424_n,
    g423_n
  );


  or

  (
    g425_n,
    g424_p,
    g423_p
  );


  and

  (
    g426_p,
    g425_n,
    G146_n_spl_011
  );


  or

  (
    g426_n,
    g425_p,
    G146_p_spl_011
  );


  and

  (
    g427_p,
    g426_n,
    g422_n
  );


  or

  (
    g427_n,
    g426_p,
    g422_p
  );


  and

  (
    g428_p,
    g427_n_spl_0,
    G23_n_spl_010
  );


  or

  (
    g428_n,
    g427_p_spl_0,
    G23_p_spl_010
  );


  and

  (
    g429_p,
    G24_n,
    G23_p_spl_011
  );


  or

  (
    g429_n,
    G24_p,
    G23_n_spl_011
  );


  and

  (
    g430_p,
    g429_n,
    g428_n
  );


  or

  (
    g430_n,
    g429_p,
    g428_p
  );


  and

  (
    g431_p,
    g430_p,
    G136_n_spl_1
  );


  and

  (
    g432_p,
    g430_n,
    G136_p_spl_0
  );


  or

  (
    g433_n,
    g432_p,
    g431_p
  );


  or

  (
    g434_n,
    g433_n,
    g418_p
  );


  or

  (
    g435_n,
    g434_n,
    g417_n
  );


  or

  (
    g436_n,
    g435_n,
    g406_n
  );


  or

  (
    g437_n,
    g436_n,
    g397_n
  );


  and

  (
    g438_p,
    g255_p_spl_00,
    G12_n_spl_010
  );


  or

  (
    g438_n,
    g255_n_spl_00,
    G12_p_spl_010
  );


  and

  (
    g439_p,
    G14_n,
    G12_p_spl_010
  );


  or

  (
    g439_n,
    G14_p,
    G12_n_spl_010
  );


  and

  (
    g440_p,
    g439_n,
    g438_n
  );


  or

  (
    g440_n,
    g439_p,
    g438_p
  );


  and

  (
    g441_p,
    g440_n,
    G128_p_spl_1
  );


  and

  (
    g442_p,
    g391_p,
    G130_n_spl_
  );


  or

  (
    g443_n,
    g442_p,
    g441_p
  );


  and

  (
    g444_p,
    g400_n,
    G131_p_spl_1
  );


  and

  (
    g445_p,
    g262_n_spl_0,
    G12_n_spl_011
  );


  or

  (
    g445_n,
    g262_p_spl_0,
    G12_p_spl_011
  );


  and

  (
    g446_p,
    G17_n,
    G12_p_spl_011
  );


  or

  (
    g446_n,
    G17_p,
    G12_n_spl_011
  );


  and

  (
    g447_p,
    g446_n,
    g445_n
  );


  or

  (
    g447_n,
    g446_p,
    g445_p
  );


  and

  (
    g448_p,
    g447_p,
    G132_n_spl_
  );


  or

  (
    g449_n,
    g448_p,
    g444_p
  );


  and

  (
    g450_p,
    g447_n,
    G132_p_spl_1
  );


  and

  (
    g451_p,
    g271_p_spl_0,
    G12_n_spl_100
  );


  or

  (
    g451_n,
    g271_n_spl_0,
    G12_p_spl_100
  );


  and

  (
    g452_p,
    G12_p_spl_100,
    G6_n
  );


  or

  (
    g452_n,
    G12_n_spl_100,
    G6_p
  );


  and

  (
    g453_p,
    g452_n,
    g451_n
  );


  or

  (
    g453_n,
    g452_p,
    g451_p
  );


  and

  (
    g454_p,
    g453_p,
    G133_n_spl_
  );


  or

  (
    g455_n,
    g454_p,
    g450_p
  );


  and

  (
    g456_p,
    g240_p_spl_0,
    G12_n_spl_101
  );


  or

  (
    g456_n,
    g240_n_spl_00,
    G12_p_spl_101
  );


  and

  (
    g457_p,
    G13_n,
    G12_p_spl_101
  );


  or

  (
    g457_n,
    G13_p,
    G12_n_spl_101
  );


  and

  (
    g458_p,
    g457_n,
    g456_n
  );


  or

  (
    g458_n,
    g457_p,
    g456_p
  );


  and

  (
    g459_p,
    g458_n,
    G125_p_spl_1
  );


  or

  (
    g460_n,
    g459_p,
    g455_n
  );


  or

  (
    g461_n,
    g460_n,
    g449_n
  );


  or

  (
    g462_n,
    g461_n,
    g443_n
  );


  or

  (
    g463_n,
    g462_n,
    g437_n
  );


  and

  (
    g464_p,
    g290_p_spl_01,
    G12_n_spl_110
  );


  or

  (
    g464_n,
    g290_n_spl_01,
    G12_p_spl_110
  );


  and

  (
    g465_p,
    G12_p_spl_110,
    G4_n
  );


  or

  (
    g465_n,
    G12_n_spl_110,
    G4_p
  );


  and

  (
    g466_p,
    g465_n,
    g464_n
  );


  or

  (
    g466_n,
    g465_p,
    g464_p
  );


  and

  (
    g467_p,
    g466_p,
    G126_n_spl_
  );


  and

  (
    g468_p,
    g453_n,
    G133_p_spl_1
  );


  or

  (
    g469_n,
    g468_p,
    g467_p
  );


  and

  (
    g470_p,
    g280_p_spl_0,
    G12_n_spl_111
  );


  or

  (
    g470_n,
    g280_n_spl_00,
    G12_p_spl_111
  );


  and

  (
    g471_p,
    G18_n,
    G12_p_spl_111
  );


  or

  (
    g471_n,
    G18_p,
    G12_n_spl_111
  );


  and

  (
    g472_p,
    g471_n,
    g470_n
  );


  or

  (
    g472_n,
    g471_p,
    g470_p
  );


  and

  (
    g473_p,
    g472_n,
    G134_p_spl_1
  );


  and

  (
    g474_p,
    g458_p,
    G125_n_spl_
  );


  or

  (
    g475_n,
    g474_p,
    g473_p
  );


  and

  (
    g476_p,
    G145_n_spl_1000,
    G75_n
  );


  or

  (
    g476_n,
    G145_p_spl_1000,
    G75_p
  );


  and

  (
    g477_p,
    G145_p_spl_1000,
    G105_n
  );


  or

  (
    g477_n,
    G145_n_spl_1000,
    G105_p
  );


  and

  (
    g478_p,
    g477_n,
    g476_n
  );


  or

  (
    g478_n,
    g477_p,
    g476_p
  );


  and

  (
    g479_p,
    g478_n,
    G146_p_spl_100
  );


  or

  (
    g479_n,
    g478_p,
    G146_n_spl_100
  );


  and

  (
    g480_p,
    G145_p_spl_1001,
    G95_n
  );


  or

  (
    g480_n,
    G145_n_spl_1001,
    G95_p
  );


  and

  (
    g481_p,
    G145_n_spl_1001,
    G85_n
  );


  or

  (
    g481_n,
    G145_p_spl_1001,
    G85_p
  );


  and

  (
    g482_p,
    g481_n,
    g480_n
  );


  or

  (
    g482_n,
    g481_p,
    g480_p
  );


  and

  (
    g483_p,
    g482_n,
    G146_n_spl_100
  );


  or

  (
    g483_n,
    g482_p,
    G146_p_spl_100
  );


  and

  (
    g484_p,
    g483_n,
    g479_n
  );


  or

  (
    g484_n,
    g483_p,
    g479_p
  );


  and

  (
    g485_p,
    g484_n_spl_0,
    G23_n_spl_011
  );


  or

  (
    g485_n,
    g484_p_spl_0,
    G23_p_spl_011
  );


  and

  (
    g486_p,
    G23_p_spl_100,
    G19_n
  );


  or

  (
    g486_n,
    G23_n_spl_100,
    G19_p
  );


  and

  (
    g487_p,
    g486_n,
    g485_n
  );


  or

  (
    g487_n,
    g486_p,
    g485_p
  );


  and

  (
    g488_p,
    g487_p,
    G135_n_spl_1
  );


  and

  (
    g489_p,
    g487_n,
    G135_p_spl_1
  );


  and

  (
    g490_p,
    g472_p,
    G134_n_spl_1
  );


  or

  (
    g491_n,
    g490_p,
    g489_p
  );


  or

  (
    g492_n,
    g491_n,
    g488_p
  );


  or

  (
    g493_n,
    g492_n,
    g475_n
  );


  or

  (
    g494_n,
    g493_n,
    g469_n
  );


  and

  (
    g495_p,
    G145_n_spl_1010,
    G81_n
  );


  or

  (
    g495_n,
    G145_p_spl_1010,
    G81_p
  );


  and

  (
    g496_p,
    G145_p_spl_1010,
    G111_n
  );


  or

  (
    g496_n,
    G145_n_spl_1010,
    G111_p
  );


  and

  (
    g497_p,
    g496_n,
    g495_n
  );


  or

  (
    g497_n,
    g496_p,
    g495_p
  );


  and

  (
    g498_p,
    g497_n,
    G146_p_spl_101
  );


  or

  (
    g498_n,
    g497_p,
    G146_n_spl_101
  );


  and

  (
    g499_p,
    G145_p_spl_1011,
    G101_n
  );


  or

  (
    g499_n,
    G145_n_spl_1011,
    G101_p
  );


  and

  (
    g500_p,
    G145_n_spl_1011,
    G91_n
  );


  or

  (
    g500_n,
    G145_p_spl_1011,
    G91_p
  );


  and

  (
    g501_p,
    g500_n,
    g499_n
  );


  or

  (
    g501_n,
    g500_p,
    g499_p
  );


  and

  (
    g502_p,
    g501_n,
    G146_n_spl_101
  );


  or

  (
    g502_n,
    g501_p,
    G146_p_spl_101
  );


  and

  (
    g503_p,
    g502_n,
    g498_n
  );


  or

  (
    g503_n,
    g502_p,
    g498_p
  );


  and

  (
    g504_p,
    g503_n_spl_0,
    G23_n_spl_100
  );


  or

  (
    g504_n,
    g503_p_spl_0,
    G23_p_spl_100
  );


  and

  (
    g505_p,
    G25_n,
    G23_p_spl_101
  );


  or

  (
    g505_n,
    G25_p,
    G23_n_spl_101
  );


  and

  (
    g506_p,
    g505_n,
    g504_n
  );


  or

  (
    g506_n,
    g505_p,
    g504_p
  );


  and

  (
    g507_p,
    g506_n,
    G139_p_spl_1
  );


  and

  (
    g508_p,
    g194_n_spl_0,
    G23_n_spl_101
  );


  or

  (
    g508_n,
    g194_p_spl_0,
    G23_p_spl_101
  );


  and

  (
    g509_p,
    G27_n,
    G23_p_spl_110
  );


  or

  (
    g509_n,
    G27_p,
    G23_n_spl_110
  );


  and

  (
    g510_p,
    g509_n,
    g508_n
  );


  or

  (
    g510_n,
    g509_p,
    g508_p
  );


  and

  (
    g511_p,
    g510_n,
    G142_p_spl_1
  );


  or

  (
    g512_n,
    g511_p,
    g507_p
  );


  and

  (
    g513_p,
    g506_p,
    G139_n_spl_
  );


  and

  (
    g514_p,
    G145_n_spl_1100,
    G82_n
  );


  or

  (
    g514_n,
    G145_p_spl_1100,
    G82_p
  );


  and

  (
    g515_p,
    G145_p_spl_1100,
    G112_n
  );


  or

  (
    g515_n,
    G145_n_spl_1100,
    G112_p
  );


  and

  (
    g516_p,
    g515_n,
    g514_n
  );


  or

  (
    g516_n,
    g515_p,
    g514_p
  );


  and

  (
    g517_p,
    g516_n,
    G146_p_spl_110
  );


  or

  (
    g517_n,
    g516_p,
    G146_n_spl_110
  );


  and

  (
    g518_p,
    G145_p_spl_1101,
    G102_n
  );


  or

  (
    g518_n,
    G145_n_spl_1101,
    G102_p
  );


  and

  (
    g519_p,
    G145_n_spl_1101,
    G92_n
  );


  or

  (
    g519_n,
    G145_p_spl_1101,
    G92_p
  );


  and

  (
    g520_p,
    g519_n,
    g518_n
  );


  or

  (
    g520_n,
    g519_p,
    g518_p
  );


  and

  (
    g521_p,
    g520_n,
    G146_n_spl_110
  );


  or

  (
    g521_n,
    g520_p,
    G146_p_spl_110
  );


  and

  (
    g522_p,
    g521_n,
    g517_n
  );


  or

  (
    g522_n,
    g521_p,
    g517_p
  );


  and

  (
    g523_p,
    g522_n_spl_0,
    G23_n_spl_110
  );


  or

  (
    g523_n,
    g522_p_spl_0,
    G23_p_spl_110
  );


  and

  (
    g524_p,
    G23_p_spl_11,
    G20_n
  );


  or

  (
    g524_n,
    G23_n_spl_11,
    G20_p
  );


  and

  (
    g525_p,
    g524_n,
    g523_n
  );


  or

  (
    g525_n,
    g524_p,
    g523_p
  );


  and

  (
    g526_p,
    g525_n,
    G138_p_spl_0
  );


  and

  (
    g527_p,
    g525_p,
    G138_n_spl_1
  );


  or

  (
    g528_n,
    g527_p,
    g526_p
  );


  or

  (
    g529_n,
    g528_n,
    g513_p
  );


  or

  (
    g530_n,
    g529_n,
    g512_n
  );


  and

  (
    g531_p,
    g395_n,
    G129_p_spl_1
  );


  and

  (
    g532_p,
    g510_p,
    G142_n_spl_
  );


  or

  (
    g533_n,
    g532_p,
    g531_p
  );


  and

  (
    g534_p,
    g466_n,
    G126_p_spl_1
  );


  and

  (
    g535_p,
    g440_p,
    G128_n_spl_
  );


  or

  (
    g536_n,
    g535_p,
    g534_p
  );


  or

  (
    g537_n,
    g536_n,
    g533_n
  );


  or

  (
    g538_n,
    g537_n,
    g530_n
  );


  or

  (
    g539_n,
    g538_n,
    g494_n
  );


  or

  (
    g540_n,
    g539_n,
    g463_n
  );


  and

  (
    g541_p,
    g290_p_spl_01,
    G118_p_spl_
  );


  or

  (
    g541_n,
    g290_n_spl_01,
    G118_n_spl_
  );


  and

  (
    g542_p,
    g204_p_spl_11,
    G51_p
  );


  or

  (
    g542_n,
    g204_n_spl_11,
    G51_n
  );


  and

  (
    g543_p,
    G117_n_spl_1110,
    G62_p
  );


  or

  (
    g543_n,
    G117_p_spl_1110,
    G62_n
  );


  and

  (
    g544_p,
    g543_n,
    G120_n_spl_111
  );


  or

  (
    g544_n,
    g543_p,
    G120_p_spl_111
  );


  and

  (
    g545_p,
    G117_n_spl_1110,
    G41_n
  );


  or

  (
    g545_n,
    G117_p_spl_1110,
    G41_p
  );


  and

  (
    g546_p,
    g545_p,
    G120_p_spl_111
  );


  or

  (
    g546_n,
    g545_n,
    G120_n_spl_111
  );


  and

  (
    g547_p,
    G117_p_spl_111,
    G73_n
  );


  or

  (
    g547_n,
    G117_n_spl_111,
    G73_p
  );


  and

  (
    g548_p,
    g547_n,
    g546_n
  );


  or

  (
    g548_n,
    g547_p,
    g546_p
  );


  and

  (
    g549_p,
    g548_p,
    g544_n
  );


  or

  (
    g549_n,
    g548_n,
    g544_p
  );


  and

  (
    g550_p,
    g549_n,
    g542_n
  );


  or

  (
    g550_n,
    g549_p,
    g542_p
  );


  and

  (
    g551_p,
    g550_n_spl_0,
    g240_n_spl_0
  );


  or

  (
    g551_n,
    g550_p_spl_,
    g240_p_spl_1
  );


  and

  (
    g552_p,
    g550_p_spl_,
    g240_p_spl_1
  );


  or

  (
    g552_n,
    g550_n_spl_0,
    g240_n_spl_1
  );


  and

  (
    g553_p,
    g552_n,
    g551_n
  );


  or

  (
    g553_n,
    g552_p,
    g551_p
  );


  and

  (
    g554_p,
    g553_n_spl_0,
    g541_p
  );


  and

  (
    g555_p,
    g553_p_spl_0,
    g541_n
  );


  or

  (
    g556_n,
    g555_p,
    g554_p
  );


  and

  (
    g557_p,
    g556_n,
    G122_n_spl_
  );


  and

  (
    g558_p,
    g550_n_spl_1,
    G122_p
  );


  or

  (
    g559_n,
    g558_p,
    g557_p
  );


  and

  (
    g560_p,
    g194_n_spl_0,
    g185_n_spl_00
  );


  or

  (
    g560_n,
    g194_p_spl_0,
    g185_p_spl_0
  );


  and

  (
    g561_p,
    g194_p_spl_,
    g185_p_spl_1
  );


  or

  (
    g561_n,
    g194_n_spl_1,
    g185_n_spl_0
  );


  and

  (
    g562_p,
    g561_n,
    g560_n
  );


  or

  (
    g562_n,
    g561_p,
    g560_p
  );


  and

  (
    g563_p,
    g562_p_spl_,
    g310_p_spl_0
  );


  or

  (
    g563_n,
    g562_n_spl_,
    g310_n_spl_1
  );


  and

  (
    g564_p,
    g562_n_spl_,
    g310_n_spl_1
  );


  or

  (
    g564_n,
    g562_p_spl_,
    g310_p_spl_
  );


  and

  (
    g565_p,
    g564_n,
    g563_n
  );


  or

  (
    g565_n,
    g564_p,
    g563_p
  );


  and

  (
    g566_p,
    G145_n_spl_1110,
    G84_n
  );


  or

  (
    g566_n,
    G145_p_spl_1110,
    G84_p
  );


  and

  (
    g567_p,
    G145_p_spl_1110,
    G114_n
  );


  or

  (
    g567_n,
    G145_n_spl_1110,
    G114_p
  );


  and

  (
    g568_p,
    g567_n,
    g566_n
  );


  or

  (
    g568_n,
    g567_p,
    g566_p
  );


  and

  (
    g569_p,
    g568_n,
    G146_p_spl_111
  );


  or

  (
    g569_n,
    g568_p,
    G146_n_spl_111
  );


  and

  (
    g570_p,
    G145_p_spl_1111,
    G104_n
  );


  or

  (
    g570_n,
    G145_n_spl_1111,
    G104_p
  );


  and

  (
    g571_p,
    G145_n_spl_1111,
    G94_n
  );


  or

  (
    g571_n,
    G145_p_spl_1111,
    G94_p
  );


  and

  (
    g572_p,
    g571_n,
    g570_n
  );


  or

  (
    g572_n,
    g571_p,
    g570_p
  );


  and

  (
    g573_p,
    g572_n,
    G146_n_spl_111
  );


  or

  (
    g573_n,
    g572_p,
    G146_p_spl_111
  );


  and

  (
    g574_p,
    g573_n,
    g569_n
  );


  or

  (
    g574_n,
    g573_p,
    g569_p
  );


  and

  (
    g575_p,
    g574_p_spl_,
    g484_p_spl_0
  );


  or

  (
    g575_n,
    g574_n_spl_,
    g484_n_spl_0
  );


  and

  (
    g576_p,
    g574_n_spl_,
    g484_n_spl_1
  );


  or

  (
    g576_n,
    g574_p_spl_,
    g484_p_spl_1
  );


  and

  (
    g577_p,
    g576_n,
    g575_n
  );


  or

  (
    g577_n,
    g576_p,
    g575_p
  );


  and

  (
    g578_p,
    g503_n_spl_0,
    g203_n_spl_00
  );


  or

  (
    g578_n,
    g503_p_spl_0,
    g203_p_spl_0
  );


  and

  (
    g579_p,
    g503_p_spl_,
    g203_p_spl_1
  );


  or

  (
    g579_n,
    g503_n_spl_,
    g203_n_spl_0
  );


  and

  (
    g580_p,
    g579_n,
    g578_n
  );


  or

  (
    g580_n,
    g579_p,
    g578_p
  );


  and

  (
    g581_p,
    g580_n_spl_,
    g577_p_spl_
  );


  or

  (
    g581_n,
    g580_p_spl_,
    g577_n_spl_
  );


  and

  (
    g582_p,
    g580_p_spl_,
    g577_n_spl_
  );


  or

  (
    g582_n,
    g580_n_spl_,
    g577_p_spl_
  );


  and

  (
    g583_p,
    g582_n,
    g581_n
  );


  or

  (
    g583_n,
    g582_p,
    g581_p
  );


  and

  (
    g584_p,
    g522_n_spl_0,
    g427_n_spl_0
  );


  or

  (
    g584_n,
    g522_p_spl_0,
    g427_p_spl_0
  );


  and

  (
    g585_p,
    g522_p_spl_1,
    g427_p_spl_1
  );


  or

  (
    g585_n,
    g522_n_spl_1,
    g427_n_spl_1
  );


  and

  (
    g586_p,
    g585_n,
    g584_n
  );


  or

  (
    g586_n,
    g585_p,
    g584_p
  );


  and

  (
    g587_p,
    g586_n_spl_,
    g583_n_spl_
  );


  or

  (
    g587_n,
    g586_p_spl_,
    g583_p_spl_
  );


  and

  (
    g588_p,
    g586_p_spl_,
    g583_p_spl_
  );


  or

  (
    g588_n,
    g586_n_spl_,
    g583_n_spl_
  );


  and

  (
    g589_p,
    g588_n,
    g587_n
  );


  or

  (
    g589_n,
    g588_p,
    g587_p
  );


  or

  (
    g590_n,
    g589_p,
    g565_n
  );


  or

  (
    g591_n,
    g589_n,
    g565_p
  );


  and

  (
    g592_p,
    g591_n,
    G29_n_spl_
  );


  and

  (
    g593_p,
    g592_p,
    g590_n
  );


  or

  (
    g594_n,
    g550_n_spl_1,
    G123_p_spl_1
  );


  and

  (
    g595_p,
    g262_n_spl_0,
    g213_p_spl_00
  );


  or

  (
    g595_n,
    g262_p_spl_0,
    g213_n_spl_0
  );


  and

  (
    g596_p,
    g262_p_spl_1,
    g213_n_spl_1
  );


  or

  (
    g596_n,
    g262_n_spl_1,
    g213_p_spl_0
  );


  and

  (
    g597_p,
    g596_n,
    g595_n
  );


  or

  (
    g597_n,
    g596_p,
    g595_p
  );


  and

  (
    g598_p,
    g280_n_spl_00,
    g271_n_spl_0
  );


  or

  (
    g598_n,
    g280_p_spl_0,
    g271_p_spl_0
  );


  and

  (
    g599_p,
    g280_p_spl_1,
    g271_p_spl_1
  );


  or

  (
    g599_n,
    g280_n_spl_0,
    g271_n_spl_1
  );


  and

  (
    g600_p,
    g599_n,
    g598_n
  );


  or

  (
    g600_n,
    g599_p,
    g598_p
  );


  and

  (
    g601_p,
    g600_n_spl_,
    g597_p_spl_
  );


  or

  (
    g601_n,
    g600_p_spl_,
    g597_n_spl_
  );


  and

  (
    g602_p,
    g600_p_spl_,
    g597_n_spl_
  );


  or

  (
    g602_n,
    g600_n_spl_,
    g597_p_spl_
  );


  and

  (
    g603_p,
    g602_n,
    g601_n
  );


  or

  (
    g603_n,
    g602_p,
    g601_p
  );


  and

  (
    g604_p,
    g290_n_spl_10,
    g255_p_spl_00
  );


  or

  (
    g604_n,
    g290_p_spl_1,
    g255_n_spl_0
  );


  and

  (
    g605_p,
    g290_p_spl_1,
    g255_n_spl_1
  );


  or

  (
    g605_n,
    g290_n_spl_10,
    g255_p_spl_0
  );


  and

  (
    g606_p,
    g605_n,
    g604_n
  );


  or

  (
    g606_n,
    g605_p,
    g604_p
  );


  and

  (
    g607_p,
    g606_n_spl_,
    g553_p_spl_0
  );


  or

  (
    g607_n,
    g606_p_spl_,
    g553_n_spl_0
  );


  and

  (
    g608_p,
    g606_p_spl_,
    g553_n_spl_
  );


  or

  (
    g608_n,
    g606_n_spl_,
    g553_p_spl_
  );


  and

  (
    g609_p,
    g608_n,
    g607_n
  );


  or

  (
    g609_n,
    g608_p,
    g607_p
  );


  and

  (
    g610_p,
    g609_n_spl_0,
    g298_p_spl_0
  );


  or

  (
    g610_n,
    g609_p_spl_0,
    g298_n_spl_
  );


  and

  (
    g611_p,
    g609_p_spl_0,
    g298_n_spl_
  );


  or

  (
    g611_n,
    g609_n_spl_0,
    g298_p_spl_
  );


  and

  (
    g612_p,
    g611_n,
    g610_n
  );


  or

  (
    g612_n,
    g611_p,
    g610_p
  );


  or

  (
    g613_n,
    g612_n,
    g603_p_spl_
  );


  or

  (
    g614_n,
    g612_p,
    g603_n_spl_
  );


  and

  (
    g615_p,
    g614_n,
    g613_n
  );


  or

  (
    g616_n,
    g615_p,
    G123_n_spl_1
  );


  and

  (
    g617_p,
    g616_n,
    g594_n
  );


  and

  (
    g618_p,
    g231_n_spl_0,
    g222_p_spl_01
  );


  or

  (
    g618_n,
    g231_p_spl_00,
    g222_n_spl_0
  );


  and

  (
    g619_p,
    g231_p_spl_01,
    g222_n_spl_1
  );


  or

  (
    g619_n,
    g231_n_spl_1,
    g222_p_spl_01
  );


  and

  (
    g620_p,
    g619_n,
    g618_n
  );


  or

  (
    g620_n,
    g619_p,
    g618_p
  );


  and

  (
    g621_p,
    g620_p_spl_,
    g609_n_spl_1
  );


  or

  (
    g621_n,
    g620_n_spl_,
    g609_p_spl_1
  );


  and

  (
    g622_p,
    g620_n_spl_,
    g609_p_spl_1
  );


  or

  (
    g622_n,
    g620_p_spl_,
    g609_n_spl_1
  );


  and

  (
    g623_p,
    g622_n,
    g621_n
  );


  or

  (
    g623_n,
    g622_p,
    g621_p
  );


  or

  (
    g624_n,
    g623_p,
    g603_n_spl_
  );


  or

  (
    g625_n,
    g623_n,
    g603_p_spl_
  );


  and

  (
    g626_p,
    g625_n,
    G29_n_spl_
  );


  and

  (
    g627_p,
    g626_p,
    g624_n
  );


  and

  (
    g628_p,
    g203_p_spl_1,
    G127_n
  );


  or

  (
    g628_n,
    g203_n_spl_1,
    G127_p
  );


  and

  (
    g629_p,
    g185_n_spl_1,
    G30_p
  );


  or

  (
    g629_n,
    g185_p_spl_1,
    G30_n
  );


  and

  (
    g630_p,
    g629_p_spl_,
    g628_p_spl_
  );


  or

  (
    g630_n,
    g629_n_spl_,
    g628_n_spl_
  );


  or

  (
    g631_n,
    g630_p_spl_00,
    G8_n_spl_
  );


  or

  (
    g632_n,
    g631_n_spl_0,
    G133_p_spl_1
  );


  and

  (
    g633_p,
    g630_p_spl_00,
    G8_p_spl_0
  );


  or

  (
    g633_n,
    g630_n_spl_00,
    G8_n_spl_
  );


  and

  (
    g634_p,
    g633_p_spl_,
    g271_p_spl_1
  );


  or

  (
    g635_n,
    g631_n_spl_0,
    G132_p_spl_1
  );


  and

  (
    g636_p,
    g633_p_spl_,
    g262_n_spl_1
  );


  and

  (
    g637_p,
    g213_p_spl_1,
    G8_p_spl_0
  );


  or

  (
    g638_n,
    g631_n_spl_1,
    G131_p_spl_1
  );


  or

  (
    g639_n,
    g633_n_spl_,
    G142_p_spl_1
  );


  and

  (
    g640_p,
    g639_n,
    g638_n
  );


  or

  (
    g641_n,
    g640_p_spl_,
    g637_p_spl_
  );


  and

  (
    g642_p,
    g640_p_spl_,
    g637_p_spl_
  );


  and

  (
    g643_p,
    g222_p_spl_1,
    G8_p_spl_
  );


  or

  (
    g644_n,
    g631_n_spl_1,
    G130_p_spl_1
  );


  or

  (
    g645_n,
    g633_n_spl_,
    G141_p_spl_1
  );


  and

  (
    g646_p,
    g645_n,
    g644_n
  );


  or

  (
    g647_n,
    g646_p_spl_,
    g643_p_spl_
  );


  and

  (
    g648_p,
    g646_p_spl_,
    g643_p_spl_
  );


  and

  (
    g649_p,
    g630_n_spl_00,
    G129_p_spl_1
  );


  and

  (
    g650_p,
    g630_p_spl_01,
    G140_p_spl_1
  );


  or

  (
    g651_n,
    g650_p,
    g649_p
  );


  or

  (
    g652_n,
    g651_n_spl_,
    g231_p_spl_01
  );


  and

  (
    g653_p,
    g651_n_spl_,
    g231_p_spl_1
  );


  and

  (
    g654_p,
    g630_n_spl_0,
    G128_p_spl_1
  );


  and

  (
    g655_p,
    g630_p_spl_01,
    G139_p_spl_1
  );


  or

  (
    g656_n,
    g655_p,
    g654_p
  );


  and

  (
    g657_p,
    g656_n_spl_,
    g255_p_spl_1
  );


  or

  (
    g658_n,
    g657_p,
    g653_p
  );


  and

  (
    g659_p,
    g630_n_spl_1,
    G126_p_spl_1
  );


  and

  (
    g660_p,
    g630_p_spl_1,
    G138_p_spl_1
  );


  or

  (
    g661_n,
    g660_p,
    g659_p
  );


  and

  (
    g662_p,
    g661_n_spl_,
    g290_n_spl_11
  );


  or

  (
    g663_n,
    g630_n_spl_1,
    G136_p_spl_1
  );


  or

  (
    g664_n,
    g630_p_spl_1,
    G125_p_spl_1
  );


  and

  (
    g665_p,
    g664_n,
    g663_n
  );


  or

  (
    g666_n,
    g665_p,
    g662_p
  );


  or

  (
    g667_n,
    g666_n,
    g240_n_spl_1
  );


  or

  (
    g668_n,
    g661_n_spl_,
    g290_n_spl_11
  );


  or

  (
    g669_n,
    g656_n_spl_,
    g255_p_spl_1
  );


  and

  (
    g670_p,
    g669_n,
    g668_n
  );


  and

  (
    g671_p,
    g670_p,
    g667_n
  );


  or

  (
    g672_n,
    g671_p,
    g658_n
  );


  and

  (
    g673_p,
    g672_n,
    g652_n
  );


  or

  (
    g674_n,
    g673_p,
    g648_p
  );


  and

  (
    g675_p,
    g674_n,
    g647_n
  );


  or

  (
    g676_n,
    g675_p,
    g642_p
  );


  and

  (
    g677_p,
    g676_n,
    g641_n
  );


  or

  (
    g678_n,
    g677_p,
    g636_p
  );


  and

  (
    g679_p,
    g678_n,
    g635_n
  );


  or

  (
    g680_n,
    g679_p,
    g634_p
  );


  and

  (
    g681_p,
    g680_n,
    g632_n
  );


  and

  (
    g682_p,
    g629_p_spl_,
    g628_n_spl_
  );


  or

  (
    g682_n,
    g629_n_spl_,
    g628_p_spl_
  );


  and

  (
    g683_p,
    g682_p_spl_00,
    G136_n_spl_1
  );


  or

  (
    g683_n,
    g682_n_spl_00,
    G136_p_spl_1
  );


  and

  (
    g684_p,
    g682_p_spl_00,
    g427_p_spl_1
  );


  or

  (
    g684_n,
    g682_n_spl_00,
    g427_n_spl_1
  );


  and

  (
    g685_p,
    g684_p_spl_,
    g683_n_spl_
  );


  and

  (
    g686_p,
    g682_p_spl_01,
    G138_n_spl_1
  );


  or

  (
    g686_n,
    g682_n_spl_01,
    G138_p_spl_1
  );


  and

  (
    g687_p,
    g682_p_spl_01,
    g522_n_spl_1
  );


  or

  (
    g687_n,
    g682_n_spl_01,
    g522_p_spl_1
  );


  and

  (
    g688_p,
    g687_n,
    g686_p
  );


  or

  (
    g688_n,
    g687_p_spl_,
    g686_n_spl_
  );


  and

  (
    g689_p,
    g687_p_spl_,
    g686_n_spl_
  );


  or

  (
    g690_n,
    g689_p,
    g688_p
  );


  and

  (
    g691_p,
    g684_n,
    g683_p
  );


  or

  (
    g691_n,
    g684_p_spl_,
    g683_n_spl_
  );


  or

  (
    g692_n,
    g691_p,
    g690_n_spl_
  );


  or

  (
    g693_n,
    g692_n,
    g685_p
  );


  and

  (
    g694_p,
    g682_p_spl_10,
    G135_n_spl_1
  );


  or

  (
    g694_n,
    g682_n_spl_10,
    G135_p_spl_1
  );


  and

  (
    g695_p,
    g682_p_spl_10,
    g484_p_spl_1
  );


  or

  (
    g695_n,
    g682_n_spl_10,
    g484_n_spl_1
  );


  and

  (
    g696_p,
    g695_n,
    g694_p
  );


  or

  (
    g696_n,
    g695_p_spl_,
    g694_n_spl_
  );


  and

  (
    g697_p,
    g695_p_spl_,
    g694_n_spl_
  );


  or

  (
    g698_n,
    g697_p,
    g696_p
  );


  and

  (
    g699_p,
    g682_p_spl_11,
    g280_p_spl_1
  );


  or

  (
    g699_n,
    g682_n_spl_11,
    g280_n_spl_1
  );


  and

  (
    g700_p,
    g682_p_spl_11,
    G134_n_spl_1
  );


  or

  (
    g700_n,
    g682_n_spl_11,
    G134_p_spl_1
  );


  and

  (
    g701_p,
    g700_p,
    g699_n
  );


  or

  (
    g701_n,
    g700_n_spl_,
    g699_p_spl_
  );


  and

  (
    g702_p,
    g700_n_spl_,
    g699_p_spl_
  );


  or

  (
    g703_n,
    g702_p,
    g701_p
  );


  or

  (
    g704_n,
    g703_n,
    g698_n_spl_
  );


  or

  (
    g705_n,
    g704_n,
    g693_n_spl_
  );


  or

  (
    g706_n,
    g705_n,
    g681_p
  );


  or

  (
    g707_n,
    g701_n,
    g698_n_spl_
  );


  and

  (
    g708_p,
    g707_n,
    g696_n
  );


  or

  (
    g709_n,
    g708_p,
    g693_n_spl_
  );


  or

  (
    g710_n,
    g691_n,
    g690_n_spl_
  );


  and

  (
    g711_p,
    g710_n,
    g709_n
  );


  and

  (
    g712_p,
    g711_p,
    g688_n
  );


  and

  (
    g713_p,
    g712_p,
    g706_n
  );


  or

  (
    g714_n,
    g361_p_spl_,
    g342_p_spl_
  );


  or

  (
    g715_n,
    g714_n,
    g388_p_spl_
  );


  or

  (
    g716_n,
    g593_p_spl_,
    g176_n_spl_0
  );


  or

  (
    g717_n,
    g716_n,
    g627_p_spl_
  );


  or

  (
    g718_n,
    g717_n,
    g715_n
  );


  buf

  (
    G2531,
    G115_n_spl_0
  );


  buf

  (
    G2532,
    G115_n_spl_1
  );


  buf

  (
    G2533,
    G115_n_spl_1
  );


  buf

  (
    G2534,
    G124_n_spl_
  );


  buf

  (
    G2535,
    G124_n_spl_
  );


  buf

  (
    G2536,
    G137_n_spl_0
  );


  buf

  (
    G2537,
    G137_n_spl_0
  );


  buf

  (
    G2538,
    G137_n_spl_
  );


  buf

  (
    G2539,
    G32_n_spl_
  );


  buf

  (
    G2540,
    G106_n_spl_
  );


  buf

  (
    G2541,
    G64_n_spl_
  );


  buf

  (
    G2542,
    G76_n_spl_
  );


  buf

  (
    G2543,
    G53_n_spl_
  );


  buf

  (
    G2544,
    G96_n_spl_
  );


  buf

  (
    G2545,
    G43_n_spl_
  );


  buf

  (
    G2546,
    G86_n_spl_
  );


  buf

  (
    G2547,
    g160_n
  );


  buf

  (
    G2548,
    g162_n
  );


  buf

  (
    G2549,
    G115_p
  );


  buf

  (
    G2550,
    g163_p
  );


  buf

  (
    G2551,
    g164_n_spl_
  );


  buf

  (
    G2552,
    g165_n
  );


  buf

  (
    G2553,
    g166_n
  );


  buf

  (
    G2554,
    g173_n_spl_
  );


  buf

  (
    G2555,
    g173_n_spl_
  );


  buf

  (
    G2556,
    g176_n_spl_
  );


  buf

  (
    G2557,
    g185_n_spl_1
  );


  buf

  (
    G2558,
    g194_n_spl_1
  );


  buf

  (
    G2559,
    g203_n_spl_1
  );


  buf

  (
    G2560,
    g213_p_spl_1
  );


  buf

  (
    G2561,
    g222_p_spl_1
  );


  buf

  (
    G2562,
    g231_p_spl_1
  );


  buf

  (
    G2563,
    g241_n
  );


  buf

  (
    G2564,
    g244_n
  );


  buf

  (
    G2565,
    g246_n
  );


  buf

  (
    G2566,
    g255_n_spl_1
  );


  buf

  (
    G2567,
    g231_n_spl_1
  );


  buf

  (
    G2568,
    g222_n_spl_1
  );


  buf

  (
    G2569,
    g213_n_spl_1
  );


  buf

  (
    G2570,
    g262_p_spl_1
  );


  buf

  (
    G2571,
    g271_n_spl_1
  );


  buf

  (
    G2572,
    g280_n_spl_1
  );


  buf

  (
    G2573,
    g292_n_spl_
  );


  buf

  (
    G2574,
    g292_n_spl_
  );


  buf

  (
    G2575,
    g295_n_spl_
  );


  buf

  (
    G2576,
    g295_n_spl_
  );


  buf

  (
    G2577,
    g297_n
  );


  buf

  (
    G2578,
    g301_n_spl_
  );


  buf

  (
    G2579,
    g301_n_spl_
  );


  buf

  (
    G2580,
    g314_n
  );


  not

  (
    G2581,
    g342_p_spl_
  );


  buf

  (
    G2582,
    g361_p_spl_
  );


  buf

  (
    G2583,
    g388_p_spl_
  );


  buf

  (
    G2584,
    g540_n_spl_
  );


  buf

  (
    G2585,
    g540_n_spl_
  );


  buf

  (
    G2586,
    g559_n
  );


  not

  (
    G2587,
    g593_p_spl_
  );


  buf

  (
    G2588,
    g617_p_spl_
  );


  buf

  (
    G2589,
    g617_p_spl_
  );


  not

  (
    G2590,
    g627_p_spl_
  );


  buf

  (
    G2591,
    g713_p
  );


  buf

  (
    G2592,
    1'b0
  );


  buf

  (
    G2593,
    g718_n_spl_
  );


  buf

  (
    G2594,
    g718_n_spl_
  );


  buf

  (
    G142_p_spl_,
    G142_p
  );


  buf

  (
    G142_p_spl_0,
    G142_p_spl_
  );


  buf

  (
    G142_p_spl_1,
    G142_p_spl_
  );


  buf

  (
    G141_p_spl_,
    G141_p
  );


  buf

  (
    G141_p_spl_0,
    G141_p_spl_
  );


  buf

  (
    G141_p_spl_1,
    G141_p_spl_
  );


  buf

  (
    G142_n_spl_,
    G142_n
  );


  buf

  (
    G142_n_spl_0,
    G142_n_spl_
  );


  buf

  (
    G141_n_spl_,
    G141_n
  );


  buf

  (
    G141_n_spl_0,
    G141_n_spl_
  );


  buf

  (
    G140_p_spl_,
    G140_p
  );


  buf

  (
    G140_p_spl_0,
    G140_p_spl_
  );


  buf

  (
    G140_p_spl_1,
    G140_p_spl_
  );


  buf

  (
    G139_p_spl_,
    G139_p
  );


  buf

  (
    G139_p_spl_0,
    G139_p_spl_
  );


  buf

  (
    G139_p_spl_1,
    G139_p_spl_
  );


  buf

  (
    G140_n_spl_,
    G140_n
  );


  buf

  (
    G140_n_spl_0,
    G140_n_spl_
  );


  buf

  (
    G139_n_spl_,
    G139_n
  );


  buf

  (
    G139_n_spl_0,
    G139_n_spl_
  );


  buf

  (
    g159_n_spl_,
    g159_n
  );


  buf

  (
    g158_n_spl_,
    g158_n
  );


  buf

  (
    G121_n_spl_,
    G121_n
  );


  buf

  (
    G115_n_spl_,
    G115_n
  );


  buf

  (
    G115_n_spl_0,
    G115_n_spl_
  );


  buf

  (
    G115_n_spl_1,
    G115_n_spl_
  );


  buf

  (
    g164_n_spl_,
    g164_n
  );


  buf

  (
    g164_n_spl_0,
    g164_n_spl_
  );


  buf

  (
    G53_n_spl_,
    G53_n
  );


  buf

  (
    G43_n_spl_,
    G43_n
  );


  buf

  (
    G96_n_spl_,
    G96_n
  );


  buf

  (
    G86_n_spl_,
    G86_n
  );


  buf

  (
    G64_n_spl_,
    G64_n
  );


  buf

  (
    G32_n_spl_,
    G32_n
  );


  buf

  (
    G106_n_spl_,
    G106_n
  );


  buf

  (
    G76_n_spl_,
    G76_n
  );


  buf

  (
    g172_n_spl_,
    g172_n
  );


  buf

  (
    g169_n_spl_,
    g169_n
  );


  buf

  (
    G145_n_spl_,
    G145_n
  );


  buf

  (
    G145_n_spl_0,
    G145_n_spl_
  );


  buf

  (
    G145_n_spl_00,
    G145_n_spl_0
  );


  buf

  (
    G145_n_spl_000,
    G145_n_spl_00
  );


  buf

  (
    G145_n_spl_0000,
    G145_n_spl_000
  );


  buf

  (
    G145_n_spl_00000,
    G145_n_spl_0000
  );


  buf

  (
    G145_n_spl_00001,
    G145_n_spl_0000
  );


  buf

  (
    G145_n_spl_0001,
    G145_n_spl_000
  );


  buf

  (
    G145_n_spl_00010,
    G145_n_spl_0001
  );


  buf

  (
    G145_n_spl_00011,
    G145_n_spl_0001
  );


  buf

  (
    G145_n_spl_001,
    G145_n_spl_00
  );


  buf

  (
    G145_n_spl_0010,
    G145_n_spl_001
  );


  buf

  (
    G145_n_spl_0011,
    G145_n_spl_001
  );


  buf

  (
    G145_n_spl_01,
    G145_n_spl_0
  );


  buf

  (
    G145_n_spl_010,
    G145_n_spl_01
  );


  buf

  (
    G145_n_spl_0100,
    G145_n_spl_010
  );


  buf

  (
    G145_n_spl_0101,
    G145_n_spl_010
  );


  buf

  (
    G145_n_spl_011,
    G145_n_spl_01
  );


  buf

  (
    G145_n_spl_0110,
    G145_n_spl_011
  );


  buf

  (
    G145_n_spl_0111,
    G145_n_spl_011
  );


  buf

  (
    G145_n_spl_1,
    G145_n_spl_
  );


  buf

  (
    G145_n_spl_10,
    G145_n_spl_1
  );


  buf

  (
    G145_n_spl_100,
    G145_n_spl_10
  );


  buf

  (
    G145_n_spl_1000,
    G145_n_spl_100
  );


  buf

  (
    G145_n_spl_1001,
    G145_n_spl_100
  );


  buf

  (
    G145_n_spl_101,
    G145_n_spl_10
  );


  buf

  (
    G145_n_spl_1010,
    G145_n_spl_101
  );


  buf

  (
    G145_n_spl_1011,
    G145_n_spl_101
  );


  buf

  (
    G145_n_spl_11,
    G145_n_spl_1
  );


  buf

  (
    G145_n_spl_110,
    G145_n_spl_11
  );


  buf

  (
    G145_n_spl_1100,
    G145_n_spl_110
  );


  buf

  (
    G145_n_spl_1101,
    G145_n_spl_110
  );


  buf

  (
    G145_n_spl_111,
    G145_n_spl_11
  );


  buf

  (
    G145_n_spl_1110,
    G145_n_spl_111
  );


  buf

  (
    G145_n_spl_1111,
    G145_n_spl_111
  );


  buf

  (
    G145_p_spl_,
    G145_p
  );


  buf

  (
    G145_p_spl_0,
    G145_p_spl_
  );


  buf

  (
    G145_p_spl_00,
    G145_p_spl_0
  );


  buf

  (
    G145_p_spl_000,
    G145_p_spl_00
  );


  buf

  (
    G145_p_spl_0000,
    G145_p_spl_000
  );


  buf

  (
    G145_p_spl_00000,
    G145_p_spl_0000
  );


  buf

  (
    G145_p_spl_00001,
    G145_p_spl_0000
  );


  buf

  (
    G145_p_spl_0001,
    G145_p_spl_000
  );


  buf

  (
    G145_p_spl_00010,
    G145_p_spl_0001
  );


  buf

  (
    G145_p_spl_00011,
    G145_p_spl_0001
  );


  buf

  (
    G145_p_spl_001,
    G145_p_spl_00
  );


  buf

  (
    G145_p_spl_0010,
    G145_p_spl_001
  );


  buf

  (
    G145_p_spl_0011,
    G145_p_spl_001
  );


  buf

  (
    G145_p_spl_01,
    G145_p_spl_0
  );


  buf

  (
    G145_p_spl_010,
    G145_p_spl_01
  );


  buf

  (
    G145_p_spl_0100,
    G145_p_spl_010
  );


  buf

  (
    G145_p_spl_0101,
    G145_p_spl_010
  );


  buf

  (
    G145_p_spl_011,
    G145_p_spl_01
  );


  buf

  (
    G145_p_spl_0110,
    G145_p_spl_011
  );


  buf

  (
    G145_p_spl_0111,
    G145_p_spl_011
  );


  buf

  (
    G145_p_spl_1,
    G145_p_spl_
  );


  buf

  (
    G145_p_spl_10,
    G145_p_spl_1
  );


  buf

  (
    G145_p_spl_100,
    G145_p_spl_10
  );


  buf

  (
    G145_p_spl_1000,
    G145_p_spl_100
  );


  buf

  (
    G145_p_spl_1001,
    G145_p_spl_100
  );


  buf

  (
    G145_p_spl_101,
    G145_p_spl_10
  );


  buf

  (
    G145_p_spl_1010,
    G145_p_spl_101
  );


  buf

  (
    G145_p_spl_1011,
    G145_p_spl_101
  );


  buf

  (
    G145_p_spl_11,
    G145_p_spl_1
  );


  buf

  (
    G145_p_spl_110,
    G145_p_spl_11
  );


  buf

  (
    G145_p_spl_1100,
    G145_p_spl_110
  );


  buf

  (
    G145_p_spl_1101,
    G145_p_spl_110
  );


  buf

  (
    G145_p_spl_111,
    G145_p_spl_11
  );


  buf

  (
    G145_p_spl_1110,
    G145_p_spl_111
  );


  buf

  (
    G145_p_spl_1111,
    G145_p_spl_111
  );


  buf

  (
    G146_p_spl_,
    G146_p
  );


  buf

  (
    G146_p_spl_0,
    G146_p_spl_
  );


  buf

  (
    G146_p_spl_00,
    G146_p_spl_0
  );


  buf

  (
    G146_p_spl_000,
    G146_p_spl_00
  );


  buf

  (
    G146_p_spl_0000,
    G146_p_spl_000
  );


  buf

  (
    G146_p_spl_0001,
    G146_p_spl_000
  );


  buf

  (
    G146_p_spl_001,
    G146_p_spl_00
  );


  buf

  (
    G146_p_spl_01,
    G146_p_spl_0
  );


  buf

  (
    G146_p_spl_010,
    G146_p_spl_01
  );


  buf

  (
    G146_p_spl_011,
    G146_p_spl_01
  );


  buf

  (
    G146_p_spl_1,
    G146_p_spl_
  );


  buf

  (
    G146_p_spl_10,
    G146_p_spl_1
  );


  buf

  (
    G146_p_spl_100,
    G146_p_spl_10
  );


  buf

  (
    G146_p_spl_101,
    G146_p_spl_10
  );


  buf

  (
    G146_p_spl_11,
    G146_p_spl_1
  );


  buf

  (
    G146_p_spl_110,
    G146_p_spl_11
  );


  buf

  (
    G146_p_spl_111,
    G146_p_spl_11
  );


  buf

  (
    G146_n_spl_,
    G146_n
  );


  buf

  (
    G146_n_spl_0,
    G146_n_spl_
  );


  buf

  (
    G146_n_spl_00,
    G146_n_spl_0
  );


  buf

  (
    G146_n_spl_000,
    G146_n_spl_00
  );


  buf

  (
    G146_n_spl_0000,
    G146_n_spl_000
  );


  buf

  (
    G146_n_spl_0001,
    G146_n_spl_000
  );


  buf

  (
    G146_n_spl_001,
    G146_n_spl_00
  );


  buf

  (
    G146_n_spl_01,
    G146_n_spl_0
  );


  buf

  (
    G146_n_spl_010,
    G146_n_spl_01
  );


  buf

  (
    G146_n_spl_011,
    G146_n_spl_01
  );


  buf

  (
    G146_n_spl_1,
    G146_n_spl_
  );


  buf

  (
    G146_n_spl_10,
    G146_n_spl_1
  );


  buf

  (
    G146_n_spl_100,
    G146_n_spl_10
  );


  buf

  (
    G146_n_spl_101,
    G146_n_spl_10
  );


  buf

  (
    G146_n_spl_11,
    G146_n_spl_1
  );


  buf

  (
    G146_n_spl_110,
    G146_n_spl_11
  );


  buf

  (
    G146_n_spl_111,
    G146_n_spl_11
  );


  buf

  (
    G120_n_spl_,
    G120_n
  );


  buf

  (
    G120_n_spl_0,
    G120_n_spl_
  );


  buf

  (
    G120_n_spl_00,
    G120_n_spl_0
  );


  buf

  (
    G120_n_spl_000,
    G120_n_spl_00
  );


  buf

  (
    G120_n_spl_0000,
    G120_n_spl_000
  );


  buf

  (
    G120_n_spl_0001,
    G120_n_spl_000
  );


  buf

  (
    G120_n_spl_001,
    G120_n_spl_00
  );


  buf

  (
    G120_n_spl_0010,
    G120_n_spl_001
  );


  buf

  (
    G120_n_spl_0011,
    G120_n_spl_001
  );


  buf

  (
    G120_n_spl_01,
    G120_n_spl_0
  );


  buf

  (
    G120_n_spl_010,
    G120_n_spl_01
  );


  buf

  (
    G120_n_spl_0100,
    G120_n_spl_010
  );


  buf

  (
    G120_n_spl_011,
    G120_n_spl_01
  );


  buf

  (
    G120_n_spl_1,
    G120_n_spl_
  );


  buf

  (
    G120_n_spl_10,
    G120_n_spl_1
  );


  buf

  (
    G120_n_spl_100,
    G120_n_spl_10
  );


  buf

  (
    G120_n_spl_101,
    G120_n_spl_10
  );


  buf

  (
    G120_n_spl_11,
    G120_n_spl_1
  );


  buf

  (
    G120_n_spl_110,
    G120_n_spl_11
  );


  buf

  (
    G120_n_spl_111,
    G120_n_spl_11
  );


  buf

  (
    G117_p_spl_,
    G117_p
  );


  buf

  (
    G117_p_spl_0,
    G117_p_spl_
  );


  buf

  (
    G117_p_spl_00,
    G117_p_spl_0
  );


  buf

  (
    G117_p_spl_000,
    G117_p_spl_00
  );


  buf

  (
    G117_p_spl_0000,
    G117_p_spl_000
  );


  buf

  (
    G117_p_spl_0001,
    G117_p_spl_000
  );


  buf

  (
    G117_p_spl_001,
    G117_p_spl_00
  );


  buf

  (
    G117_p_spl_0010,
    G117_p_spl_001
  );


  buf

  (
    G117_p_spl_0011,
    G117_p_spl_001
  );


  buf

  (
    G117_p_spl_01,
    G117_p_spl_0
  );


  buf

  (
    G117_p_spl_010,
    G117_p_spl_01
  );


  buf

  (
    G117_p_spl_0100,
    G117_p_spl_010
  );


  buf

  (
    G117_p_spl_0101,
    G117_p_spl_010
  );


  buf

  (
    G117_p_spl_011,
    G117_p_spl_01
  );


  buf

  (
    G117_p_spl_0110,
    G117_p_spl_011
  );


  buf

  (
    G117_p_spl_0111,
    G117_p_spl_011
  );


  buf

  (
    G117_p_spl_1,
    G117_p_spl_
  );


  buf

  (
    G117_p_spl_10,
    G117_p_spl_1
  );


  buf

  (
    G117_p_spl_100,
    G117_p_spl_10
  );


  buf

  (
    G117_p_spl_1000,
    G117_p_spl_100
  );


  buf

  (
    G117_p_spl_1001,
    G117_p_spl_100
  );


  buf

  (
    G117_p_spl_101,
    G117_p_spl_10
  );


  buf

  (
    G117_p_spl_1010,
    G117_p_spl_101
  );


  buf

  (
    G117_p_spl_1011,
    G117_p_spl_101
  );


  buf

  (
    G117_p_spl_11,
    G117_p_spl_1
  );


  buf

  (
    G117_p_spl_110,
    G117_p_spl_11
  );


  buf

  (
    G117_p_spl_1100,
    G117_p_spl_110
  );


  buf

  (
    G117_p_spl_1101,
    G117_p_spl_110
  );


  buf

  (
    G117_p_spl_111,
    G117_p_spl_11
  );


  buf

  (
    G117_p_spl_1110,
    G117_p_spl_111
  );


  buf

  (
    G120_p_spl_,
    G120_p
  );


  buf

  (
    G120_p_spl_0,
    G120_p_spl_
  );


  buf

  (
    G120_p_spl_00,
    G120_p_spl_0
  );


  buf

  (
    G120_p_spl_000,
    G120_p_spl_00
  );


  buf

  (
    G120_p_spl_0000,
    G120_p_spl_000
  );


  buf

  (
    G120_p_spl_0001,
    G120_p_spl_000
  );


  buf

  (
    G120_p_spl_001,
    G120_p_spl_00
  );


  buf

  (
    G120_p_spl_0010,
    G120_p_spl_001
  );


  buf

  (
    G120_p_spl_0011,
    G120_p_spl_001
  );


  buf

  (
    G120_p_spl_01,
    G120_p_spl_0
  );


  buf

  (
    G120_p_spl_010,
    G120_p_spl_01
  );


  buf

  (
    G120_p_spl_0100,
    G120_p_spl_010
  );


  buf

  (
    G120_p_spl_011,
    G120_p_spl_01
  );


  buf

  (
    G120_p_spl_1,
    G120_p_spl_
  );


  buf

  (
    G120_p_spl_10,
    G120_p_spl_1
  );


  buf

  (
    G120_p_spl_100,
    G120_p_spl_10
  );


  buf

  (
    G120_p_spl_101,
    G120_p_spl_10
  );


  buf

  (
    G120_p_spl_11,
    G120_p_spl_1
  );


  buf

  (
    G120_p_spl_110,
    G120_p_spl_11
  );


  buf

  (
    G120_p_spl_111,
    G120_p_spl_11
  );


  buf

  (
    G117_n_spl_,
    G117_n
  );


  buf

  (
    G117_n_spl_0,
    G117_n_spl_
  );


  buf

  (
    G117_n_spl_00,
    G117_n_spl_0
  );


  buf

  (
    G117_n_spl_000,
    G117_n_spl_00
  );


  buf

  (
    G117_n_spl_0000,
    G117_n_spl_000
  );


  buf

  (
    G117_n_spl_0001,
    G117_n_spl_000
  );


  buf

  (
    G117_n_spl_001,
    G117_n_spl_00
  );


  buf

  (
    G117_n_spl_0010,
    G117_n_spl_001
  );


  buf

  (
    G117_n_spl_0011,
    G117_n_spl_001
  );


  buf

  (
    G117_n_spl_01,
    G117_n_spl_0
  );


  buf

  (
    G117_n_spl_010,
    G117_n_spl_01
  );


  buf

  (
    G117_n_spl_0100,
    G117_n_spl_010
  );


  buf

  (
    G117_n_spl_0101,
    G117_n_spl_010
  );


  buf

  (
    G117_n_spl_011,
    G117_n_spl_01
  );


  buf

  (
    G117_n_spl_0110,
    G117_n_spl_011
  );


  buf

  (
    G117_n_spl_0111,
    G117_n_spl_011
  );


  buf

  (
    G117_n_spl_1,
    G117_n_spl_
  );


  buf

  (
    G117_n_spl_10,
    G117_n_spl_1
  );


  buf

  (
    G117_n_spl_100,
    G117_n_spl_10
  );


  buf

  (
    G117_n_spl_1000,
    G117_n_spl_100
  );


  buf

  (
    G117_n_spl_1001,
    G117_n_spl_100
  );


  buf

  (
    G117_n_spl_101,
    G117_n_spl_10
  );


  buf

  (
    G117_n_spl_1010,
    G117_n_spl_101
  );


  buf

  (
    G117_n_spl_1011,
    G117_n_spl_101
  );


  buf

  (
    G117_n_spl_11,
    G117_n_spl_1
  );


  buf

  (
    G117_n_spl_110,
    G117_n_spl_11
  );


  buf

  (
    G117_n_spl_1100,
    G117_n_spl_110
  );


  buf

  (
    G117_n_spl_1101,
    G117_n_spl_110
  );


  buf

  (
    G117_n_spl_111,
    G117_n_spl_11
  );


  buf

  (
    G117_n_spl_1110,
    G117_n_spl_111
  );


  buf

  (
    g204_p_spl_,
    g204_p
  );


  buf

  (
    g204_p_spl_0,
    g204_p_spl_
  );


  buf

  (
    g204_p_spl_00,
    g204_p_spl_0
  );


  buf

  (
    g204_p_spl_000,
    g204_p_spl_00
  );


  buf

  (
    g204_p_spl_01,
    g204_p_spl_0
  );


  buf

  (
    g204_p_spl_1,
    g204_p_spl_
  );


  buf

  (
    g204_p_spl_10,
    g204_p_spl_1
  );


  buf

  (
    g204_p_spl_11,
    g204_p_spl_1
  );


  buf

  (
    g204_n_spl_,
    g204_n
  );


  buf

  (
    g204_n_spl_0,
    g204_n_spl_
  );


  buf

  (
    g204_n_spl_00,
    g204_n_spl_0
  );


  buf

  (
    g204_n_spl_000,
    g204_n_spl_00
  );


  buf

  (
    g204_n_spl_01,
    g204_n_spl_0
  );


  buf

  (
    g204_n_spl_1,
    g204_n_spl_
  );


  buf

  (
    g204_n_spl_10,
    g204_n_spl_1
  );


  buf

  (
    g204_n_spl_11,
    g204_n_spl_1
  );


  buf

  (
    g240_n_spl_,
    g240_n
  );


  buf

  (
    g240_n_spl_0,
    g240_n_spl_
  );


  buf

  (
    g240_n_spl_00,
    g240_n_spl_0
  );


  buf

  (
    g240_n_spl_1,
    g240_n_spl_
  );


  buf

  (
    G122_n_spl_,
    G122_n
  );


  buf

  (
    G122_n_spl_0,
    G122_n_spl_
  );


  buf

  (
    g176_n_spl_,
    g176_n
  );


  buf

  (
    g176_n_spl_0,
    g176_n_spl_
  );


  buf

  (
    g243_n_spl_,
    g243_n
  );


  buf

  (
    g231_n_spl_,
    g231_n
  );


  buf

  (
    g231_n_spl_0,
    g231_n_spl_
  );


  buf

  (
    g231_n_spl_00,
    g231_n_spl_0
  );


  buf

  (
    g231_n_spl_1,
    g231_n_spl_
  );


  buf

  (
    G123_p_spl_,
    G123_p
  );


  buf

  (
    G123_p_spl_0,
    G123_p_spl_
  );


  buf

  (
    G123_p_spl_1,
    G123_p_spl_
  );


  buf

  (
    g290_p_spl_,
    g290_p
  );


  buf

  (
    g290_p_spl_0,
    g290_p_spl_
  );


  buf

  (
    g290_p_spl_00,
    g290_p_spl_0
  );


  buf

  (
    g290_p_spl_01,
    g290_p_spl_0
  );


  buf

  (
    g290_p_spl_1,
    g290_p_spl_
  );


  buf

  (
    G123_n_spl_,
    G123_n
  );


  buf

  (
    G123_n_spl_0,
    G123_n_spl_
  );


  buf

  (
    G123_n_spl_1,
    G123_n_spl_
  );


  buf

  (
    g222_p_spl_,
    g222_p
  );


  buf

  (
    g222_p_spl_0,
    g222_p_spl_
  );


  buf

  (
    g222_p_spl_00,
    g222_p_spl_0
  );


  buf

  (
    g222_p_spl_01,
    g222_p_spl_0
  );


  buf

  (
    g222_p_spl_1,
    g222_p_spl_
  );


  buf

  (
    g255_n_spl_,
    g255_n
  );


  buf

  (
    g255_n_spl_0,
    g255_n_spl_
  );


  buf

  (
    g255_n_spl_00,
    g255_n_spl_0
  );


  buf

  (
    g255_n_spl_1,
    g255_n_spl_
  );


  buf

  (
    G118_p_spl_,
    G118_p
  );


  buf

  (
    G118_p_spl_0,
    G118_p_spl_
  );


  buf

  (
    g290_n_spl_,
    g290_n
  );


  buf

  (
    g290_n_spl_0,
    g290_n_spl_
  );


  buf

  (
    g290_n_spl_00,
    g290_n_spl_0
  );


  buf

  (
    g290_n_spl_01,
    g290_n_spl_0
  );


  buf

  (
    g290_n_spl_1,
    g290_n_spl_
  );


  buf

  (
    g290_n_spl_10,
    g290_n_spl_1
  );


  buf

  (
    g290_n_spl_11,
    g290_n_spl_1
  );


  buf

  (
    G118_n_spl_,
    G118_n
  );


  buf

  (
    g298_p_spl_,
    g298_p
  );


  buf

  (
    g298_p_spl_0,
    g298_p_spl_
  );


  buf

  (
    g240_p_spl_,
    g240_p
  );


  buf

  (
    g240_p_spl_0,
    g240_p_spl_
  );


  buf

  (
    g240_p_spl_1,
    g240_p_spl_
  );


  buf

  (
    g310_p_spl_,
    g310_p
  );


  buf

  (
    g310_p_spl_0,
    g310_p_spl_
  );


  buf

  (
    G143_n_spl_,
    G143_n
  );


  buf

  (
    G143_n_spl_0,
    G143_n_spl_
  );


  buf

  (
    g310_n_spl_,
    g310_n
  );


  buf

  (
    g310_n_spl_0,
    g310_n_spl_
  );


  buf

  (
    g310_n_spl_1,
    g310_n_spl_
  );


  buf

  (
    G143_p_spl_,
    G143_p
  );


  buf

  (
    G143_p_spl_0,
    G143_p_spl_
  );


  buf

  (
    G144_p_spl_,
    G144_p
  );


  buf

  (
    G144_p_spl_0,
    G144_p_spl_
  );


  buf

  (
    G155_n_spl_,
    G155_n
  );


  buf

  (
    G154_n_spl_,
    G154_n
  );


  buf

  (
    G155_p_spl_,
    G155_p
  );


  buf

  (
    G154_p_spl_,
    G154_p
  );


  buf

  (
    G126_n_spl_,
    G126_n
  );


  buf

  (
    G126_n_spl_0,
    G126_n_spl_
  );


  buf

  (
    G125_n_spl_,
    G125_n
  );


  buf

  (
    G125_n_spl_0,
    G125_n_spl_
  );


  buf

  (
    G126_p_spl_,
    G126_p
  );


  buf

  (
    G126_p_spl_0,
    G126_p_spl_
  );


  buf

  (
    G126_p_spl_1,
    G126_p_spl_
  );


  buf

  (
    G125_p_spl_,
    G125_p
  );


  buf

  (
    G125_p_spl_0,
    G125_p_spl_
  );


  buf

  (
    G125_p_spl_1,
    G125_p_spl_
  );


  buf

  (
    g320_n_spl_,
    g320_n
  );


  buf

  (
    g317_p_spl_,
    g317_p
  );


  buf

  (
    g320_p_spl_,
    g320_p
  );


  buf

  (
    g317_n_spl_,
    g317_n
  );


  buf

  (
    G153_n_spl_,
    G153_n
  );


  buf

  (
    G152_n_spl_,
    G152_n
  );


  buf

  (
    G153_p_spl_,
    G153_p
  );


  buf

  (
    G152_p_spl_,
    G152_p
  );


  buf

  (
    G149_n_spl_,
    G149_n
  );


  buf

  (
    G148_n_spl_,
    G148_n
  );


  buf

  (
    G149_p_spl_,
    G149_p
  );


  buf

  (
    G148_p_spl_,
    G148_p
  );


  buf

  (
    g329_n_spl_,
    g329_n
  );


  buf

  (
    g326_n_spl_,
    g326_n
  );


  buf

  (
    g329_p_spl_,
    g329_p
  );


  buf

  (
    g326_p_spl_,
    g326_p
  );


  buf

  (
    G151_n_spl_,
    G151_n
  );


  buf

  (
    G150_n_spl_,
    G150_n
  );


  buf

  (
    G151_p_spl_,
    G151_p
  );


  buf

  (
    G150_p_spl_,
    G150_p
  );


  buf

  (
    g335_n_spl_,
    g335_n
  );


  buf

  (
    g332_n_spl_,
    g332_n
  );


  buf

  (
    g335_p_spl_,
    g335_p
  );


  buf

  (
    g332_p_spl_,
    g332_p
  );


  buf

  (
    G157_n_spl_,
    G157_n
  );


  buf

  (
    G138_p_spl_,
    G138_p
  );


  buf

  (
    G138_p_spl_0,
    G138_p_spl_
  );


  buf

  (
    G138_p_spl_00,
    G138_p_spl_0
  );


  buf

  (
    G138_p_spl_1,
    G138_p_spl_
  );


  buf

  (
    G157_p_spl_,
    G157_p
  );


  buf

  (
    G138_n_spl_,
    G138_n
  );


  buf

  (
    G138_n_spl_0,
    G138_n_spl_
  );


  buf

  (
    G138_n_spl_1,
    G138_n_spl_
  );


  buf

  (
    g349_n_spl_,
    g349_n
  );


  buf

  (
    g346_n_spl_,
    g346_n
  );


  buf

  (
    g349_p_spl_,
    g349_p
  );


  buf

  (
    g346_p_spl_,
    g346_p
  );


  buf

  (
    g352_n_spl_,
    g352_n
  );


  buf

  (
    g344_n_spl_,
    g344_n
  );


  buf

  (
    g352_p_spl_,
    g352_p
  );


  buf

  (
    g344_p_spl_,
    g344_p
  );


  buf

  (
    G144_n_spl_,
    G144_n
  );


  buf

  (
    G134_n_spl_,
    G134_n
  );


  buf

  (
    G134_n_spl_0,
    G134_n_spl_
  );


  buf

  (
    G134_n_spl_1,
    G134_n_spl_
  );


  buf

  (
    G133_n_spl_,
    G133_n
  );


  buf

  (
    G133_n_spl_0,
    G133_n_spl_
  );


  buf

  (
    G134_p_spl_,
    G134_p
  );


  buf

  (
    G134_p_spl_0,
    G134_p_spl_
  );


  buf

  (
    G134_p_spl_1,
    G134_p_spl_
  );


  buf

  (
    G133_p_spl_,
    G133_p
  );


  buf

  (
    G133_p_spl_0,
    G133_p_spl_
  );


  buf

  (
    G133_p_spl_1,
    G133_p_spl_
  );


  buf

  (
    G136_n_spl_,
    G136_n
  );


  buf

  (
    G136_n_spl_0,
    G136_n_spl_
  );


  buf

  (
    G136_n_spl_1,
    G136_n_spl_
  );


  buf

  (
    G135_n_spl_,
    G135_n
  );


  buf

  (
    G135_n_spl_0,
    G135_n_spl_
  );


  buf

  (
    G135_n_spl_1,
    G135_n_spl_
  );


  buf

  (
    G136_p_spl_,
    G136_p
  );


  buf

  (
    G136_p_spl_0,
    G136_p_spl_
  );


  buf

  (
    G136_p_spl_00,
    G136_p_spl_0
  );


  buf

  (
    G136_p_spl_1,
    G136_p_spl_
  );


  buf

  (
    G135_p_spl_,
    G135_p
  );


  buf

  (
    G135_p_spl_0,
    G135_p_spl_
  );


  buf

  (
    G135_p_spl_1,
    G135_p_spl_
  );


  buf

  (
    g367_n_spl_,
    g367_n
  );


  buf

  (
    g364_p_spl_,
    g364_p
  );


  buf

  (
    g367_p_spl_,
    g367_p
  );


  buf

  (
    g364_n_spl_,
    g364_n
  );


  buf

  (
    G132_n_spl_,
    G132_n
  );


  buf

  (
    G132_n_spl_0,
    G132_n_spl_
  );


  buf

  (
    G131_n_spl_,
    G131_n
  );


  buf

  (
    G131_n_spl_0,
    G131_n_spl_
  );


  buf

  (
    G132_p_spl_,
    G132_p
  );


  buf

  (
    G132_p_spl_0,
    G132_p_spl_
  );


  buf

  (
    G132_p_spl_1,
    G132_p_spl_
  );


  buf

  (
    G131_p_spl_,
    G131_p
  );


  buf

  (
    G131_p_spl_0,
    G131_p_spl_
  );


  buf

  (
    G131_p_spl_1,
    G131_p_spl_
  );


  buf

  (
    G156_n_spl_,
    G156_n
  );


  buf

  (
    G128_p_spl_,
    G128_p
  );


  buf

  (
    G128_p_spl_0,
    G128_p_spl_
  );


  buf

  (
    G128_p_spl_1,
    G128_p_spl_
  );


  buf

  (
    G156_p_spl_,
    G156_p
  );


  buf

  (
    G128_n_spl_,
    G128_n
  );


  buf

  (
    G128_n_spl_0,
    G128_n_spl_
  );


  buf

  (
    g376_n_spl_,
    g376_n
  );


  buf

  (
    g373_n_spl_,
    g373_n
  );


  buf

  (
    g376_p_spl_,
    g376_p
  );


  buf

  (
    g373_p_spl_,
    g373_p
  );


  buf

  (
    G130_n_spl_,
    G130_n
  );


  buf

  (
    G130_n_spl_0,
    G130_n_spl_
  );


  buf

  (
    G129_n_spl_,
    G129_n
  );


  buf

  (
    G129_n_spl_0,
    G129_n_spl_
  );


  buf

  (
    G130_p_spl_,
    G130_p
  );


  buf

  (
    G130_p_spl_0,
    G130_p_spl_
  );


  buf

  (
    G130_p_spl_1,
    G130_p_spl_
  );


  buf

  (
    G129_p_spl_,
    G129_p
  );


  buf

  (
    G129_p_spl_0,
    G129_p_spl_
  );


  buf

  (
    G129_p_spl_1,
    G129_p_spl_
  );


  buf

  (
    g382_n_spl_,
    g382_n
  );


  buf

  (
    g379_n_spl_,
    g379_n
  );


  buf

  (
    g382_p_spl_,
    g382_p
  );


  buf

  (
    g379_p_spl_,
    g379_p
  );


  buf

  (
    G12_n_spl_,
    G12_n
  );


  buf

  (
    G12_n_spl_0,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_00,
    G12_n_spl_0
  );


  buf

  (
    G12_n_spl_000,
    G12_n_spl_00
  );


  buf

  (
    G12_n_spl_0000,
    G12_n_spl_000
  );


  buf

  (
    G12_n_spl_0001,
    G12_n_spl_000
  );


  buf

  (
    G12_n_spl_001,
    G12_n_spl_00
  );


  buf

  (
    G12_n_spl_01,
    G12_n_spl_0
  );


  buf

  (
    G12_n_spl_010,
    G12_n_spl_01
  );


  buf

  (
    G12_n_spl_011,
    G12_n_spl_01
  );


  buf

  (
    G12_n_spl_1,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_10,
    G12_n_spl_1
  );


  buf

  (
    G12_n_spl_100,
    G12_n_spl_10
  );


  buf

  (
    G12_n_spl_101,
    G12_n_spl_10
  );


  buf

  (
    G12_n_spl_11,
    G12_n_spl_1
  );


  buf

  (
    G12_n_spl_110,
    G12_n_spl_11
  );


  buf

  (
    G12_n_spl_111,
    G12_n_spl_11
  );


  buf

  (
    g222_n_spl_,
    g222_n
  );


  buf

  (
    g222_n_spl_0,
    g222_n_spl_
  );


  buf

  (
    g222_n_spl_1,
    g222_n_spl_
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G12_p_spl_0,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_00,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_000,
    G12_p_spl_00
  );


  buf

  (
    G12_p_spl_0000,
    G12_p_spl_000
  );


  buf

  (
    G12_p_spl_0001,
    G12_p_spl_000
  );


  buf

  (
    G12_p_spl_001,
    G12_p_spl_00
  );


  buf

  (
    G12_p_spl_01,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_010,
    G12_p_spl_01
  );


  buf

  (
    G12_p_spl_011,
    G12_p_spl_01
  );


  buf

  (
    G12_p_spl_1,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_10,
    G12_p_spl_1
  );


  buf

  (
    G12_p_spl_100,
    G12_p_spl_10
  );


  buf

  (
    G12_p_spl_101,
    G12_p_spl_10
  );


  buf

  (
    G12_p_spl_11,
    G12_p_spl_1
  );


  buf

  (
    G12_p_spl_110,
    G12_p_spl_11
  );


  buf

  (
    G12_p_spl_111,
    G12_p_spl_11
  );


  buf

  (
    g231_p_spl_,
    g231_p
  );


  buf

  (
    g231_p_spl_0,
    g231_p_spl_
  );


  buf

  (
    g231_p_spl_00,
    g231_p_spl_0
  );


  buf

  (
    g231_p_spl_01,
    g231_p_spl_0
  );


  buf

  (
    g231_p_spl_1,
    g231_p_spl_
  );


  buf

  (
    g213_p_spl_,
    g213_p
  );


  buf

  (
    g213_p_spl_0,
    g213_p_spl_
  );


  buf

  (
    g213_p_spl_00,
    g213_p_spl_0
  );


  buf

  (
    g213_p_spl_1,
    g213_p_spl_
  );


  buf

  (
    g213_n_spl_,
    g213_n
  );


  buf

  (
    g213_n_spl_0,
    g213_n_spl_
  );


  buf

  (
    g213_n_spl_1,
    g213_n_spl_
  );


  buf

  (
    G23_n_spl_,
    G23_n
  );


  buf

  (
    G23_n_spl_0,
    G23_n_spl_
  );


  buf

  (
    G23_n_spl_00,
    G23_n_spl_0
  );


  buf

  (
    G23_n_spl_000,
    G23_n_spl_00
  );


  buf

  (
    G23_n_spl_001,
    G23_n_spl_00
  );


  buf

  (
    G23_n_spl_01,
    G23_n_spl_0
  );


  buf

  (
    G23_n_spl_010,
    G23_n_spl_01
  );


  buf

  (
    G23_n_spl_011,
    G23_n_spl_01
  );


  buf

  (
    G23_n_spl_1,
    G23_n_spl_
  );


  buf

  (
    G23_n_spl_10,
    G23_n_spl_1
  );


  buf

  (
    G23_n_spl_100,
    G23_n_spl_10
  );


  buf

  (
    G23_n_spl_101,
    G23_n_spl_10
  );


  buf

  (
    G23_n_spl_11,
    G23_n_spl_1
  );


  buf

  (
    G23_n_spl_110,
    G23_n_spl_11
  );


  buf

  (
    G23_p_spl_,
    G23_p
  );


  buf

  (
    G23_p_spl_0,
    G23_p_spl_
  );


  buf

  (
    G23_p_spl_00,
    G23_p_spl_0
  );


  buf

  (
    G23_p_spl_000,
    G23_p_spl_00
  );


  buf

  (
    G23_p_spl_001,
    G23_p_spl_00
  );


  buf

  (
    G23_p_spl_01,
    G23_p_spl_0
  );


  buf

  (
    G23_p_spl_010,
    G23_p_spl_01
  );


  buf

  (
    G23_p_spl_011,
    G23_p_spl_01
  );


  buf

  (
    G23_p_spl_1,
    G23_p_spl_
  );


  buf

  (
    G23_p_spl_10,
    G23_p_spl_1
  );


  buf

  (
    G23_p_spl_100,
    G23_p_spl_10
  );


  buf

  (
    G23_p_spl_101,
    G23_p_spl_10
  );


  buf

  (
    G23_p_spl_11,
    G23_p_spl_1
  );


  buf

  (
    G23_p_spl_110,
    G23_p_spl_11
  );


  buf

  (
    g185_n_spl_,
    g185_n
  );


  buf

  (
    g185_n_spl_0,
    g185_n_spl_
  );


  buf

  (
    g185_n_spl_00,
    g185_n_spl_0
  );


  buf

  (
    g185_n_spl_1,
    g185_n_spl_
  );


  buf

  (
    g185_p_spl_,
    g185_p
  );


  buf

  (
    g185_p_spl_0,
    g185_p_spl_
  );


  buf

  (
    g185_p_spl_1,
    g185_p_spl_
  );


  buf

  (
    g203_n_spl_,
    g203_n
  );


  buf

  (
    g203_n_spl_0,
    g203_n_spl_
  );


  buf

  (
    g203_n_spl_00,
    g203_n_spl_0
  );


  buf

  (
    g203_n_spl_1,
    g203_n_spl_
  );


  buf

  (
    g203_p_spl_,
    g203_p
  );


  buf

  (
    g203_p_spl_0,
    g203_p_spl_
  );


  buf

  (
    g203_p_spl_1,
    g203_p_spl_
  );


  buf

  (
    g427_n_spl_,
    g427_n
  );


  buf

  (
    g427_n_spl_0,
    g427_n_spl_
  );


  buf

  (
    g427_n_spl_1,
    g427_n_spl_
  );


  buf

  (
    g427_p_spl_,
    g427_p
  );


  buf

  (
    g427_p_spl_0,
    g427_p_spl_
  );


  buf

  (
    g427_p_spl_1,
    g427_p_spl_
  );


  buf

  (
    g255_p_spl_,
    g255_p
  );


  buf

  (
    g255_p_spl_0,
    g255_p_spl_
  );


  buf

  (
    g255_p_spl_00,
    g255_p_spl_0
  );


  buf

  (
    g255_p_spl_1,
    g255_p_spl_
  );


  buf

  (
    g262_n_spl_,
    g262_n
  );


  buf

  (
    g262_n_spl_0,
    g262_n_spl_
  );


  buf

  (
    g262_n_spl_1,
    g262_n_spl_
  );


  buf

  (
    g262_p_spl_,
    g262_p
  );


  buf

  (
    g262_p_spl_0,
    g262_p_spl_
  );


  buf

  (
    g262_p_spl_1,
    g262_p_spl_
  );


  buf

  (
    g271_p_spl_,
    g271_p
  );


  buf

  (
    g271_p_spl_0,
    g271_p_spl_
  );


  buf

  (
    g271_p_spl_1,
    g271_p_spl_
  );


  buf

  (
    g271_n_spl_,
    g271_n
  );


  buf

  (
    g271_n_spl_0,
    g271_n_spl_
  );


  buf

  (
    g271_n_spl_1,
    g271_n_spl_
  );


  buf

  (
    g280_p_spl_,
    g280_p
  );


  buf

  (
    g280_p_spl_0,
    g280_p_spl_
  );


  buf

  (
    g280_p_spl_1,
    g280_p_spl_
  );


  buf

  (
    g280_n_spl_,
    g280_n
  );


  buf

  (
    g280_n_spl_0,
    g280_n_spl_
  );


  buf

  (
    g280_n_spl_00,
    g280_n_spl_0
  );


  buf

  (
    g280_n_spl_1,
    g280_n_spl_
  );


  buf

  (
    g484_n_spl_,
    g484_n
  );


  buf

  (
    g484_n_spl_0,
    g484_n_spl_
  );


  buf

  (
    g484_n_spl_1,
    g484_n_spl_
  );


  buf

  (
    g484_p_spl_,
    g484_p
  );


  buf

  (
    g484_p_spl_0,
    g484_p_spl_
  );


  buf

  (
    g484_p_spl_1,
    g484_p_spl_
  );


  buf

  (
    g503_n_spl_,
    g503_n
  );


  buf

  (
    g503_n_spl_0,
    g503_n_spl_
  );


  buf

  (
    g503_p_spl_,
    g503_p
  );


  buf

  (
    g503_p_spl_0,
    g503_p_spl_
  );


  buf

  (
    g194_n_spl_,
    g194_n
  );


  buf

  (
    g194_n_spl_0,
    g194_n_spl_
  );


  buf

  (
    g194_n_spl_1,
    g194_n_spl_
  );


  buf

  (
    g194_p_spl_,
    g194_p
  );


  buf

  (
    g194_p_spl_0,
    g194_p_spl_
  );


  buf

  (
    g522_n_spl_,
    g522_n
  );


  buf

  (
    g522_n_spl_0,
    g522_n_spl_
  );


  buf

  (
    g522_n_spl_1,
    g522_n_spl_
  );


  buf

  (
    g522_p_spl_,
    g522_p
  );


  buf

  (
    g522_p_spl_0,
    g522_p_spl_
  );


  buf

  (
    g522_p_spl_1,
    g522_p_spl_
  );


  buf

  (
    g550_n_spl_,
    g550_n
  );


  buf

  (
    g550_n_spl_0,
    g550_n_spl_
  );


  buf

  (
    g550_n_spl_1,
    g550_n_spl_
  );


  buf

  (
    g550_p_spl_,
    g550_p
  );


  buf

  (
    g553_n_spl_,
    g553_n
  );


  buf

  (
    g553_n_spl_0,
    g553_n_spl_
  );


  buf

  (
    g553_p_spl_,
    g553_p
  );


  buf

  (
    g553_p_spl_0,
    g553_p_spl_
  );


  buf

  (
    g562_p_spl_,
    g562_p
  );


  buf

  (
    g562_n_spl_,
    g562_n
  );


  buf

  (
    g574_p_spl_,
    g574_p
  );


  buf

  (
    g574_n_spl_,
    g574_n
  );


  buf

  (
    g580_n_spl_,
    g580_n
  );


  buf

  (
    g577_p_spl_,
    g577_p
  );


  buf

  (
    g580_p_spl_,
    g580_p
  );


  buf

  (
    g577_n_spl_,
    g577_n
  );


  buf

  (
    g586_n_spl_,
    g586_n
  );


  buf

  (
    g583_n_spl_,
    g583_n
  );


  buf

  (
    g586_p_spl_,
    g586_p
  );


  buf

  (
    g583_p_spl_,
    g583_p
  );


  buf

  (
    G29_n_spl_,
    G29_n
  );


  buf

  (
    g600_n_spl_,
    g600_n
  );


  buf

  (
    g597_p_spl_,
    g597_p
  );


  buf

  (
    g600_p_spl_,
    g600_p
  );


  buf

  (
    g597_n_spl_,
    g597_n
  );


  buf

  (
    g606_n_spl_,
    g606_n
  );


  buf

  (
    g606_p_spl_,
    g606_p
  );


  buf

  (
    g609_n_spl_,
    g609_n
  );


  buf

  (
    g609_n_spl_0,
    g609_n_spl_
  );


  buf

  (
    g609_n_spl_1,
    g609_n_spl_
  );


  buf

  (
    g609_p_spl_,
    g609_p
  );


  buf

  (
    g609_p_spl_0,
    g609_p_spl_
  );


  buf

  (
    g609_p_spl_1,
    g609_p_spl_
  );


  buf

  (
    g298_n_spl_,
    g298_n
  );


  buf

  (
    g603_p_spl_,
    g603_p
  );


  buf

  (
    g603_n_spl_,
    g603_n
  );


  buf

  (
    g620_p_spl_,
    g620_p
  );


  buf

  (
    g620_n_spl_,
    g620_n
  );


  buf

  (
    g629_p_spl_,
    g629_p
  );


  buf

  (
    g628_p_spl_,
    g628_p
  );


  buf

  (
    g629_n_spl_,
    g629_n
  );


  buf

  (
    g628_n_spl_,
    g628_n
  );


  buf

  (
    g630_p_spl_,
    g630_p
  );


  buf

  (
    g630_p_spl_0,
    g630_p_spl_
  );


  buf

  (
    g630_p_spl_00,
    g630_p_spl_0
  );


  buf

  (
    g630_p_spl_01,
    g630_p_spl_0
  );


  buf

  (
    g630_p_spl_1,
    g630_p_spl_
  );


  buf

  (
    G8_n_spl_,
    G8_n
  );


  buf

  (
    g631_n_spl_,
    g631_n
  );


  buf

  (
    g631_n_spl_0,
    g631_n_spl_
  );


  buf

  (
    g631_n_spl_1,
    g631_n_spl_
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    g630_n_spl_,
    g630_n
  );


  buf

  (
    g630_n_spl_0,
    g630_n_spl_
  );


  buf

  (
    g630_n_spl_00,
    g630_n_spl_0
  );


  buf

  (
    g630_n_spl_1,
    g630_n_spl_
  );


  buf

  (
    g633_p_spl_,
    g633_p
  );


  buf

  (
    g633_n_spl_,
    g633_n
  );


  buf

  (
    g640_p_spl_,
    g640_p
  );


  buf

  (
    g637_p_spl_,
    g637_p
  );


  buf

  (
    g646_p_spl_,
    g646_p
  );


  buf

  (
    g643_p_spl_,
    g643_p
  );


  buf

  (
    g651_n_spl_,
    g651_n
  );


  buf

  (
    g656_n_spl_,
    g656_n
  );


  buf

  (
    g661_n_spl_,
    g661_n
  );


  buf

  (
    g682_p_spl_,
    g682_p
  );


  buf

  (
    g682_p_spl_0,
    g682_p_spl_
  );


  buf

  (
    g682_p_spl_00,
    g682_p_spl_0
  );


  buf

  (
    g682_p_spl_01,
    g682_p_spl_0
  );


  buf

  (
    g682_p_spl_1,
    g682_p_spl_
  );


  buf

  (
    g682_p_spl_10,
    g682_p_spl_1
  );


  buf

  (
    g682_p_spl_11,
    g682_p_spl_1
  );


  buf

  (
    g682_n_spl_,
    g682_n
  );


  buf

  (
    g682_n_spl_0,
    g682_n_spl_
  );


  buf

  (
    g682_n_spl_00,
    g682_n_spl_0
  );


  buf

  (
    g682_n_spl_01,
    g682_n_spl_0
  );


  buf

  (
    g682_n_spl_1,
    g682_n_spl_
  );


  buf

  (
    g682_n_spl_10,
    g682_n_spl_1
  );


  buf

  (
    g682_n_spl_11,
    g682_n_spl_1
  );


  buf

  (
    g684_p_spl_,
    g684_p
  );


  buf

  (
    g683_n_spl_,
    g683_n
  );


  buf

  (
    g687_p_spl_,
    g687_p
  );


  buf

  (
    g686_n_spl_,
    g686_n
  );


  buf

  (
    g690_n_spl_,
    g690_n
  );


  buf

  (
    g695_p_spl_,
    g695_p
  );


  buf

  (
    g694_n_spl_,
    g694_n
  );


  buf

  (
    g700_n_spl_,
    g700_n
  );


  buf

  (
    g699_p_spl_,
    g699_p
  );


  buf

  (
    g698_n_spl_,
    g698_n
  );


  buf

  (
    g693_n_spl_,
    g693_n
  );


  buf

  (
    g361_p_spl_,
    g361_p
  );


  buf

  (
    g342_p_spl_,
    g342_p
  );


  buf

  (
    g388_p_spl_,
    g388_p
  );


  buf

  (
    g593_p_spl_,
    g593_p
  );


  buf

  (
    g627_p_spl_,
    g627_p
  );


  buf

  (
    G124_n_spl_,
    G124_n
  );


  buf

  (
    G137_n_spl_,
    G137_n
  );


  buf

  (
    G137_n_spl_0,
    G137_n_spl_
  );


  buf

  (
    g173_n_spl_,
    g173_n
  );


  buf

  (
    g292_n_spl_,
    g292_n
  );


  buf

  (
    g295_n_spl_,
    g295_n
  );


  buf

  (
    g301_n_spl_,
    g301_n
  );


  buf

  (
    g540_n_spl_,
    g540_n
  );


  buf

  (
    g617_p_spl_,
    g617_p
  );


  buf

  (
    g718_n_spl_,
    g718_n
  );


endmodule
