// Benchmark "mymod" written by ABC on Sun Oct 29 19:31:47 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36,
    G426, G427, G428, G429, G430, G431, G432  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36;
  output G426, G427, G428, G429, G430, G431, G432;
  reg n205_lo, n214_lo, n217_lo, n226_lo, n229_lo, n232_lo, n238_lo,
    n241_lo, n250_lo, n253_lo, n256_lo, n262_lo, n265_lo, n274_lo, n277_lo,
    n280_lo, n286_lo, n289_lo, n298_lo, n301_lo, n304_lo, n310_lo, n313_lo,
    n322_lo, n325_lo, n328_lo, n334_lo, n337_lo, n346_lo, n349_lo, n352_lo,
    n358_lo, n361_lo, n370_lo, n373_lo, n376_lo, n382_lo, n385_lo, n394_lo,
    n397_lo, n400_lo, n406_lo, n409_lo, n418_lo, n421_lo, n424_lo, n430_lo,
    n433_lo, n442_lo, n445_lo, n448_lo, n454_lo, n457_lo, n466_lo, n469_lo,
    n472_lo, n478_lo, n481_lo, n490_lo, n493_lo, n496_lo, n502_lo, n505_lo,
    n514_lo, n517_lo, n520_lo, n526_lo, n529_lo, n538_lo, n541_lo, n544_lo,
    n550_lo, n553_lo, n562_lo, n565_lo, n568_lo, n574_lo, n577_lo, n586_lo,
    n589_lo, n592_lo, n598_lo, n601_lo, n610_lo, n613_lo, n616_lo, n622_lo,
    n625_lo, n628_lo, n634_lo, n316_inv, n319_inv, n997_o2, n998_o2,
    n999_o2, n1000_o2, n1001_o2, n1002_o2, n1003_o2, n1004_o2, n1005_o2,
    n1015_o2, n1016_o2, n1017_o2, n1018_o2, n1019_o2, n1020_o2, n1021_o2,
    n1022_o2, n1023_o2, n376_1_inv, n235_lo_buf_o2, n283_lo_buf_o2,
    n331_lo_buf_o2, n379_lo_buf_o2, n427_lo_buf_o2, n475_lo_buf_o2,
    n523_lo_buf_o2, n571_lo_buf_o2, n619_lo_buf_o2, n406_1_inv, G223_o2,
    G226_o2, G229_o2, G232_o2, G235_o2, G238_o2, G242_o2, G246_o2, G250_o2,
    n259_lo_buf_o2, n307_lo_buf_o2, n355_lo_buf_o2, n403_lo_buf_o2,
    n451_lo_buf_o2, n499_lo_buf_o2, n547_lo_buf_o2, n595_lo_buf_o2,
    n631_lo_buf_o2, G213_o2, G318_o2, G358_o2, G259_o2, G263_o2, G266_o2,
    G269_o2, G272_o2, G275_o2, G278_o2, G281_o2, G284_o2, n211_lo_buf_o2,
    n247_lo_buf_o2, n295_lo_buf_o2, n343_lo_buf_o2, n391_lo_buf_o2,
    n439_lo_buf_o2, n487_lo_buf_o2, n535_lo_buf_o2, n583_lo_buf_o2,
    G158_o2, G184_o2, G186_o2, G188_o2, G190_o2, G192_o2, G194_o2, G196_o2,
    G198_o2, n223_lo_buf_o2, n271_lo_buf_o2, n319_lo_buf_o2,
    n367_lo_buf_o2, n415_lo_buf_o2, n463_lo_buf_o2, n511_lo_buf_o2,
    n559_lo_buf_o2, n607_lo_buf_o2, n580_inv, G154_o2, G159_o2, G162_o2,
    G165_o2, G168_o2, G171_o2, G174_o2, G177_o2, G180_o2;
  wire new_n420_, new_n422_, new_n424_, new_n426_, new_n428_, new_n430_,
    new_n432_, new_n434_, new_n436_, new_n438_, new_n440_, new_n442_,
    new_n444_, new_n446_, new_n448_, new_n450_, new_n452_, new_n454_,
    new_n456_, new_n458_, new_n460_, new_n462_, new_n464_, new_n466_,
    new_n468_, new_n470_, new_n472_, new_n474_, new_n476_, new_n478_,
    new_n480_, new_n482_, new_n484_, new_n486_, new_n488_, new_n490_,
    new_n492_, new_n493_, new_n495_, new_n496_, new_n498_, new_n500_,
    new_n502_, new_n503_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n510_, new_n512_, new_n513_, new_n515_, new_n516_, new_n519_,
    new_n520_, new_n522_, new_n523_, new_n524_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n532_, new_n533_, new_n534_,
    new_n536_, new_n538_, new_n539_, new_n540_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n558_, new_n559_, new_n560_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n578_,
    new_n579_, new_n580_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n590_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n599_, new_n600_, new_n602_,
    new_n603_, new_n604_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n616_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n630_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n650_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n674_, new_n676_, new_n678_, new_n680_,
    new_n682_, new_n684_, new_n686_, new_n688_, new_n690_, new_n692_,
    new_n694_, new_n696_, new_n698_, new_n700_, new_n702_, new_n704_,
    new_n706_, new_n708_, new_n710_, new_n712_, new_n714_, new_n716_,
    new_n718_, new_n720_, new_n722_, new_n724_, new_n726_, new_n728_,
    new_n730_, new_n732_, new_n735_, new_n737_, new_n739_, new_n741_,
    new_n743_, new_n745_, new_n747_, new_n749_, new_n751_, new_n752_,
    new_n754_, new_n756_, new_n758_, new_n760_, new_n762_, new_n764_,
    new_n766_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n798_, new_n800_,
    new_n802_, new_n804_, new_n806_, new_n808_, new_n810_, new_n812_,
    new_n814_, new_n816_, new_n818_, new_n820_, new_n822_, new_n824_,
    new_n826_, new_n828_, new_n830_, new_n832_, new_n834_, new_n836_,
    new_n838_, new_n840_, new_n842_, new_n844_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1304_, new_n1305_, new_n1306_, new_n1307_,
    new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_,
    new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_,
    new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_,
    new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_,
    new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_,
    new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_,
    new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_,
    new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_,
    new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_,
    new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_,
    new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_,
    new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_,
    new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_,
    new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_,
    new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, n205_li,
    n214_li, n217_li, n226_li, n229_li, n232_li, n238_li, n241_li, n250_li,
    n253_li, n256_li, n262_li, n265_li, n274_li, n277_li, n280_li, n286_li,
    n289_li, n298_li, n301_li, n304_li, n310_li, n313_li, n322_li, n325_li,
    n328_li, n334_li, n337_li, n346_li, n349_li, n352_li, n358_li, n361_li,
    n370_li, n373_li, n376_li, n382_li, n385_li, n394_li, n397_li, n400_li,
    n406_li, n409_li, n418_li, n421_li, n424_li, n430_li, n433_li, n442_li,
    n445_li, n448_li, n454_li, n457_li, n466_li, n469_li, n472_li, n478_li,
    n481_li, n490_li, n493_li, n496_li, n502_li, n505_li, n514_li, n517_li,
    n520_li, n526_li, n529_li, n538_li, n541_li, n544_li, n550_li, n553_li,
    n562_li, n565_li, n568_li, n574_li, n577_li, n586_li, n589_li, n592_li,
    n598_li, n601_li, n610_li, n613_li, n616_li, n622_li, n625_li, n628_li,
    n634_li, n919_i2, n1024_i2, n997_i2, n998_i2, n999_i2, n1000_i2,
    n1001_i2, n1002_i2, n1003_i2, n1004_i2, n1005_i2, n1015_i2, n1016_i2,
    n1017_i2, n1018_i2, n1019_i2, n1020_i2, n1021_i2, n1022_i2, n1023_i2,
    G199_i2, n235_lo_buf_i2, n283_lo_buf_i2, n331_lo_buf_i2,
    n379_lo_buf_i2, n427_lo_buf_i2, n475_lo_buf_i2, n523_lo_buf_i2,
    n571_lo_buf_i2, n619_lo_buf_i2, G355_i2, G223_i2, G226_i2, G229_i2,
    G232_i2, G235_i2, G238_i2, G242_i2, G246_i2, G250_i2, n259_lo_buf_i2,
    n307_lo_buf_i2, n355_lo_buf_i2, n403_lo_buf_i2, n451_lo_buf_i2,
    n499_lo_buf_i2, n547_lo_buf_i2, n595_lo_buf_i2, n631_lo_buf_i2,
    G213_i2, G318_i2, G358_i2, G259_i2, G263_i2, G266_i2, G269_i2, G272_i2,
    G275_i2, G278_i2, G281_i2, G284_i2, n211_lo_buf_i2, n247_lo_buf_i2,
    n295_lo_buf_i2, n343_lo_buf_i2, n391_lo_buf_i2, n439_lo_buf_i2,
    n487_lo_buf_i2, n535_lo_buf_i2, n583_lo_buf_i2, G158_i2, G184_i2,
    G186_i2, G188_i2, G190_i2, G192_i2, G194_i2, G196_i2, G198_i2,
    n223_lo_buf_i2, n271_lo_buf_i2, n319_lo_buf_i2, n367_lo_buf_i2,
    n415_lo_buf_i2, n463_lo_buf_i2, n511_lo_buf_i2, n559_lo_buf_i2,
    n607_lo_buf_i2, G295_i2, G154_i2, G159_i2, G162_i2, G165_i2, G168_i2,
    G171_i2, G174_i2, G177_i2, G180_i2;
  assign new_n420_ = G1;
  assign new_n422_ = G2;
  assign new_n424_ = G3;
  assign new_n426_ = G4;
  assign new_n428_ = G5;
  assign new_n430_ = G6;
  assign new_n432_ = G7;
  assign new_n434_ = G8;
  assign new_n436_ = G9;
  assign new_n438_ = G10;
  assign new_n440_ = G11;
  assign new_n442_ = G12;
  assign new_n444_ = G13;
  assign new_n446_ = G14;
  assign new_n448_ = G15;
  assign new_n450_ = G16;
  assign new_n452_ = G17;
  assign new_n454_ = G18;
  assign new_n456_ = G19;
  assign new_n458_ = G20;
  assign new_n460_ = G21;
  assign new_n462_ = G22;
  assign new_n464_ = G23;
  assign new_n466_ = G24;
  assign new_n468_ = G25;
  assign new_n470_ = G26;
  assign new_n472_ = G27;
  assign new_n474_ = G28;
  assign new_n476_ = G29;
  assign new_n478_ = G30;
  assign new_n480_ = G31;
  assign new_n482_ = G32;
  assign new_n484_ = G33;
  assign new_n486_ = G34;
  assign new_n488_ = G35;
  assign new_n490_ = G36;
  assign new_n492_ = n205_lo;
  assign new_n493_ = ~n205_lo;
  assign new_n495_ = ~n214_lo;
  assign new_n496_ = n217_lo;
  assign new_n498_ = n226_lo;
  assign new_n500_ = n229_lo;
  assign new_n502_ = n232_lo;
  assign new_n503_ = ~n232_lo;
  assign new_n505_ = ~n238_lo;
  assign new_n506_ = n241_lo;
  assign new_n507_ = ~n241_lo;
  assign new_n508_ = n250_lo;
  assign new_n510_ = n253_lo;
  assign new_n512_ = n256_lo;
  assign new_n513_ = ~n256_lo;
  assign new_n515_ = ~n262_lo;
  assign new_n516_ = n265_lo;
  assign new_n519_ = ~n274_lo;
  assign new_n520_ = n277_lo;
  assign new_n522_ = n280_lo;
  assign new_n523_ = ~n280_lo;
  assign new_n524_ = n286_lo;
  assign new_n526_ = n289_lo;
  assign new_n527_ = ~n289_lo;
  assign new_n528_ = n298_lo;
  assign new_n529_ = ~n298_lo;
  assign new_n530_ = n301_lo;
  assign new_n532_ = n304_lo;
  assign new_n533_ = ~n304_lo;
  assign new_n534_ = n310_lo;
  assign new_n536_ = n313_lo;
  assign new_n538_ = n322_lo;
  assign new_n539_ = ~n322_lo;
  assign new_n540_ = n325_lo;
  assign new_n542_ = n328_lo;
  assign new_n543_ = ~n328_lo;
  assign new_n544_ = n334_lo;
  assign new_n545_ = ~n334_lo;
  assign new_n546_ = n337_lo;
  assign new_n547_ = ~n337_lo;
  assign new_n548_ = n346_lo;
  assign new_n549_ = ~n346_lo;
  assign new_n550_ = n349_lo;
  assign new_n552_ = n352_lo;
  assign new_n553_ = ~n352_lo;
  assign new_n554_ = n358_lo;
  assign new_n555_ = ~n358_lo;
  assign new_n556_ = n361_lo;
  assign new_n558_ = n370_lo;
  assign new_n559_ = ~n370_lo;
  assign new_n560_ = n373_lo;
  assign new_n562_ = n376_lo;
  assign new_n563_ = ~n376_lo;
  assign new_n564_ = n382_lo;
  assign new_n565_ = ~n382_lo;
  assign new_n566_ = n385_lo;
  assign new_n567_ = ~n385_lo;
  assign new_n568_ = n394_lo;
  assign new_n569_ = ~n394_lo;
  assign new_n570_ = n397_lo;
  assign new_n572_ = n400_lo;
  assign new_n573_ = ~n400_lo;
  assign new_n574_ = n406_lo;
  assign new_n575_ = ~n406_lo;
  assign new_n576_ = n409_lo;
  assign new_n578_ = n418_lo;
  assign new_n579_ = ~n418_lo;
  assign new_n580_ = n421_lo;
  assign new_n582_ = n424_lo;
  assign new_n583_ = ~n424_lo;
  assign new_n584_ = n430_lo;
  assign new_n585_ = ~n430_lo;
  assign new_n586_ = n433_lo;
  assign new_n587_ = ~n433_lo;
  assign new_n588_ = n442_lo;
  assign new_n590_ = n445_lo;
  assign new_n592_ = n448_lo;
  assign new_n593_ = ~n448_lo;
  assign new_n594_ = n454_lo;
  assign new_n595_ = ~n454_lo;
  assign new_n596_ = n457_lo;
  assign new_n599_ = ~n466_lo;
  assign new_n600_ = n469_lo;
  assign new_n602_ = n472_lo;
  assign new_n603_ = ~n472_lo;
  assign new_n604_ = n478_lo;
  assign new_n606_ = n481_lo;
  assign new_n607_ = ~n481_lo;
  assign new_n608_ = n490_lo;
  assign new_n609_ = ~n490_lo;
  assign new_n610_ = n493_lo;
  assign new_n612_ = n496_lo;
  assign new_n613_ = ~n496_lo;
  assign new_n614_ = n502_lo;
  assign new_n616_ = n505_lo;
  assign new_n618_ = n514_lo;
  assign new_n619_ = ~n514_lo;
  assign new_n620_ = n517_lo;
  assign new_n622_ = n520_lo;
  assign new_n623_ = ~n520_lo;
  assign new_n624_ = n526_lo;
  assign new_n625_ = ~n526_lo;
  assign new_n626_ = n529_lo;
  assign new_n627_ = ~n529_lo;
  assign new_n628_ = n538_lo;
  assign new_n630_ = n541_lo;
  assign new_n632_ = n544_lo;
  assign new_n633_ = ~n544_lo;
  assign new_n634_ = n550_lo;
  assign new_n635_ = ~n550_lo;
  assign new_n636_ = n553_lo;
  assign new_n639_ = ~n562_lo;
  assign new_n640_ = n565_lo;
  assign new_n642_ = n568_lo;
  assign new_n643_ = ~n568_lo;
  assign new_n644_ = n574_lo;
  assign new_n646_ = n577_lo;
  assign new_n647_ = ~n577_lo;
  assign new_n648_ = n586_lo;
  assign new_n650_ = n589_lo;
  assign new_n652_ = n592_lo;
  assign new_n653_ = ~n592_lo;
  assign new_n654_ = n598_lo;
  assign new_n656_ = n601_lo;
  assign new_n659_ = ~n610_lo;
  assign new_n660_ = n613_lo;
  assign new_n662_ = n616_lo;
  assign new_n663_ = ~n616_lo;
  assign new_n664_ = n622_lo;
  assign new_n666_ = n625_lo;
  assign new_n668_ = n628_lo;
  assign new_n669_ = ~n628_lo;
  assign new_n670_ = n634_lo;
  assign new_n672_ = n316_inv;
  assign new_n674_ = n319_inv;
  assign new_n676_ = n997_o2;
  assign new_n678_ = n998_o2;
  assign new_n680_ = n999_o2;
  assign new_n682_ = n1000_o2;
  assign new_n684_ = n1001_o2;
  assign new_n686_ = n1002_o2;
  assign new_n688_ = n1003_o2;
  assign new_n690_ = n1004_o2;
  assign new_n692_ = n1005_o2;
  assign new_n694_ = n1015_o2;
  assign new_n696_ = n1016_o2;
  assign new_n698_ = n1017_o2;
  assign new_n700_ = n1018_o2;
  assign new_n702_ = n1019_o2;
  assign new_n704_ = n1020_o2;
  assign new_n706_ = n1021_o2;
  assign new_n708_ = n1022_o2;
  assign new_n710_ = n1023_o2;
  assign new_n712_ = n376_1_inv;
  assign new_n714_ = n235_lo_buf_o2;
  assign new_n716_ = n283_lo_buf_o2;
  assign new_n718_ = n331_lo_buf_o2;
  assign new_n720_ = n379_lo_buf_o2;
  assign new_n722_ = n427_lo_buf_o2;
  assign new_n724_ = n475_lo_buf_o2;
  assign new_n726_ = n523_lo_buf_o2;
  assign new_n728_ = n571_lo_buf_o2;
  assign new_n730_ = n619_lo_buf_o2;
  assign new_n732_ = n406_1_inv;
  assign new_n735_ = ~G223_o2;
  assign new_n737_ = ~G226_o2;
  assign new_n739_ = ~G229_o2;
  assign new_n741_ = ~G232_o2;
  assign new_n743_ = ~G235_o2;
  assign new_n745_ = ~G238_o2;
  assign new_n747_ = ~G242_o2;
  assign new_n749_ = ~G246_o2;
  assign new_n751_ = ~G250_o2;
  assign new_n752_ = n259_lo_buf_o2;
  assign new_n754_ = n307_lo_buf_o2;
  assign new_n756_ = n355_lo_buf_o2;
  assign new_n758_ = n403_lo_buf_o2;
  assign new_n760_ = n451_lo_buf_o2;
  assign new_n762_ = n499_lo_buf_o2;
  assign new_n764_ = n547_lo_buf_o2;
  assign new_n766_ = n595_lo_buf_o2;
  assign new_n768_ = n631_lo_buf_o2;
  assign new_n770_ = G213_o2;
  assign new_n771_ = ~G213_o2;
  assign new_n772_ = G318_o2;
  assign new_n773_ = ~G318_o2;
  assign new_n774_ = G358_o2;
  assign new_n775_ = ~G358_o2;
  assign new_n776_ = G259_o2;
  assign new_n777_ = ~G259_o2;
  assign new_n778_ = G263_o2;
  assign new_n779_ = ~G263_o2;
  assign new_n780_ = G266_o2;
  assign new_n781_ = ~G266_o2;
  assign new_n782_ = G269_o2;
  assign new_n783_ = ~G269_o2;
  assign new_n784_ = G272_o2;
  assign new_n785_ = ~G272_o2;
  assign new_n786_ = G275_o2;
  assign new_n787_ = ~G275_o2;
  assign new_n788_ = G278_o2;
  assign new_n789_ = ~G278_o2;
  assign new_n790_ = G281_o2;
  assign new_n791_ = ~G281_o2;
  assign new_n792_ = G284_o2;
  assign new_n793_ = ~G284_o2;
  assign new_n794_ = n211_lo_buf_o2;
  assign new_n796_ = n247_lo_buf_o2;
  assign new_n798_ = n295_lo_buf_o2;
  assign new_n800_ = n343_lo_buf_o2;
  assign new_n802_ = n391_lo_buf_o2;
  assign new_n804_ = n439_lo_buf_o2;
  assign new_n806_ = n487_lo_buf_o2;
  assign new_n808_ = n535_lo_buf_o2;
  assign new_n810_ = n583_lo_buf_o2;
  assign new_n812_ = G158_o2;
  assign new_n814_ = G184_o2;
  assign new_n816_ = G186_o2;
  assign new_n818_ = G188_o2;
  assign new_n820_ = G190_o2;
  assign new_n822_ = G192_o2;
  assign new_n824_ = G194_o2;
  assign new_n826_ = G196_o2;
  assign new_n828_ = G198_o2;
  assign new_n830_ = n223_lo_buf_o2;
  assign new_n832_ = n271_lo_buf_o2;
  assign new_n834_ = n319_lo_buf_o2;
  assign new_n836_ = n367_lo_buf_o2;
  assign new_n838_ = n415_lo_buf_o2;
  assign new_n840_ = n463_lo_buf_o2;
  assign new_n842_ = n511_lo_buf_o2;
  assign new_n844_ = n559_lo_buf_o2;
  assign new_n846_ = n607_lo_buf_o2;
  assign new_n848_ = n580_inv;
  assign new_n849_ = ~n580_inv;
  assign new_n850_ = G154_o2;
  assign new_n851_ = ~G154_o2;
  assign new_n852_ = G159_o2;
  assign new_n853_ = ~G159_o2;
  assign new_n854_ = G162_o2;
  assign new_n855_ = ~G162_o2;
  assign new_n856_ = G165_o2;
  assign new_n857_ = ~G165_o2;
  assign new_n858_ = G168_o2;
  assign new_n859_ = ~G168_o2;
  assign new_n860_ = G171_o2;
  assign new_n861_ = ~G171_o2;
  assign new_n862_ = G174_o2;
  assign new_n863_ = ~G174_o2;
  assign new_n864_ = G177_o2;
  assign new_n865_ = ~G177_o2;
  assign new_n866_ = G180_o2;
  assign new_n867_ = ~G180_o2;
  assign new_n868_ = new_n1306_ | new_n495_;
  assign new_n869_ = new_n1310_ | new_n505_;
  assign new_n870_ = new_n1314_ | new_n515_;
  assign new_n871_ = new_n868_ & new_n498_;
  assign new_n872_ = new_n871_ & new_n869_;
  assign new_n873_ = new_n872_ & new_n870_;
  assign new_n874_ = new_n1318_ & new_n508_;
  assign new_n875_ = new_n1325_ & new_n524_;
  assign new_n876_ = new_n1332_ & new_n534_;
  assign new_n877_ = new_n875_ | new_n874_;
  assign new_n878_ = new_n877_ | new_n876_;
  assign new_n879_ = new_n878_ | new_n519_;
  assign new_n880_ = new_n1318_ & new_n528_;
  assign new_n881_ = new_n1306_ | new_n529_;
  assign new_n882_ = new_n1325_ & new_n544_;
  assign new_n883_ = new_n1310_ | new_n545_;
  assign new_n884_ = new_n1332_ & new_n554_;
  assign new_n885_ = new_n1314_ | new_n555_;
  assign new_n886_ = new_n883_ & new_n881_;
  assign new_n887_ = new_n882_ | new_n880_;
  assign new_n888_ = new_n886_ & new_n885_;
  assign new_n889_ = new_n887_ | new_n884_;
  assign new_n890_ = new_n888_ & new_n538_;
  assign new_n891_ = new_n889_ | new_n539_;
  assign new_n892_ = new_n1319_ & new_n548_;
  assign new_n893_ = new_n1305_ | new_n549_;
  assign new_n894_ = new_n1326_ & new_n564_;
  assign new_n895_ = new_n1309_ | new_n565_;
  assign new_n896_ = new_n1333_ & new_n574_;
  assign new_n897_ = new_n1313_ | new_n575_;
  assign new_n898_ = new_n895_ & new_n893_;
  assign new_n899_ = new_n894_ | new_n892_;
  assign new_n900_ = new_n898_ & new_n897_;
  assign new_n901_ = new_n899_ | new_n896_;
  assign new_n902_ = new_n900_ & new_n558_;
  assign new_n903_ = new_n901_ | new_n559_;
  assign new_n904_ = new_n1319_ & new_n568_;
  assign new_n905_ = new_n1307_ | new_n569_;
  assign new_n906_ = new_n1326_ & new_n584_;
  assign new_n907_ = new_n1311_ | new_n585_;
  assign new_n908_ = new_n1333_ & new_n594_;
  assign new_n909_ = new_n1315_ | new_n595_;
  assign new_n910_ = new_n907_ & new_n905_;
  assign new_n911_ = new_n906_ | new_n904_;
  assign new_n912_ = new_n910_ & new_n909_;
  assign new_n913_ = new_n911_ | new_n908_;
  assign new_n914_ = new_n912_ & new_n578_;
  assign new_n915_ = new_n913_ | new_n579_;
  assign new_n916_ = new_n1321_ & new_n588_;
  assign new_n917_ = new_n1328_ & new_n604_;
  assign new_n918_ = new_n1335_ & new_n614_;
  assign new_n919_ = new_n917_ | new_n916_;
  assign new_n920_ = new_n919_ | new_n918_;
  assign new_n921_ = new_n920_ | new_n599_;
  assign new_n922_ = new_n1321_ & new_n608_;
  assign new_n923_ = new_n1307_ | new_n609_;
  assign new_n924_ = new_n1328_ & new_n624_;
  assign new_n925_ = new_n1311_ | new_n625_;
  assign new_n926_ = new_n1335_ & new_n634_;
  assign new_n927_ = new_n1315_ | new_n635_;
  assign new_n928_ = new_n925_ & new_n923_;
  assign new_n929_ = new_n924_ | new_n922_;
  assign new_n930_ = new_n928_ & new_n927_;
  assign new_n931_ = new_n929_ | new_n926_;
  assign new_n932_ = new_n930_ & new_n618_;
  assign new_n933_ = new_n931_ | new_n619_;
  assign new_n934_ = new_n1322_ & new_n628_;
  assign new_n935_ = new_n1329_ & new_n644_;
  assign new_n936_ = new_n1336_ & new_n654_;
  assign new_n937_ = new_n935_ | new_n934_;
  assign new_n938_ = new_n937_ | new_n936_;
  assign new_n939_ = new_n938_ | new_n639_;
  assign new_n940_ = new_n1322_ & new_n648_;
  assign new_n941_ = new_n1329_ & new_n664_;
  assign new_n942_ = new_n1336_ & new_n670_;
  assign new_n943_ = new_n941_ | new_n940_;
  assign new_n944_ = new_n943_ | new_n942_;
  assign new_n945_ = new_n944_ | new_n659_;
  assign new_n946_ = new_n891_ & new_n1337_;
  assign new_n947_ = new_n1339_ & new_n1340_;
  assign new_n948_ = new_n947_ & new_n1341_;
  assign new_n949_ = new_n948_ & new_n1342_;
  assign new_n950_ = new_n949_ & new_n1343_;
  assign new_n951_ = new_n950_ & new_n1344_;
  assign new_n952_ = new_n951_ & new_n945_;
  assign new_n953_ = new_n952_ | new_n873_;
  assign new_n954_ = new_n1340_ | new_n1345_;
  assign new_n955_ = new_n1346_ & new_n1339_;
  assign new_n956_ = new_n955_ & new_n1341_;
  assign new_n957_ = new_n1347_ | new_n1345_;
  assign new_n958_ = new_n1348_ | new_n1342_;
  assign new_n959_ = new_n958_ | new_n1349_;
  assign new_n960_ = new_n1349_ | new_n1347_;
  assign new_n961_ = new_n960_ | new_n1343_;
  assign new_n962_ = new_n1350_ & new_n1338_;
  assign new_n963_ = new_n962_ & new_n961_;
  assign new_n964_ = new_n1348_ | new_n932_;
  assign new_n965_ = new_n964_ | new_n1344_;
  assign new_n966_ = new_n1346_ & new_n1337_;
  assign new_n967_ = new_n966_ & new_n1350_;
  assign new_n968_ = new_n967_ & new_n965_;
  assign new_n969_ = new_n1351_ & new_n1352_;
  assign new_n970_ = new_n1353_ | new_n1354_;
  assign new_n971_ = new_n969_ & new_n1355_;
  assign new_n972_ = new_n970_ | new_n1356_;
  assign new_n973_ = new_n971_ & new_n1357_;
  assign new_n974_ = new_n972_ | new_n1358_;
  assign new_n975_ = new_n973_ & new_n1359_;
  assign new_n976_ = new_n974_ | new_n1360_;
  assign new_n977_ = new_n975_ & new_n1361_;
  assign new_n978_ = new_n976_ | new_n1362_;
  assign new_n979_ = new_n977_ & new_n1363_;
  assign new_n980_ = new_n978_ | new_n1364_;
  assign new_n981_ = new_n979_ & new_n1365_;
  assign new_n982_ = new_n980_ | new_n1366_;
  assign new_n983_ = new_n981_ & new_n1367_;
  assign new_n984_ = new_n982_ | new_n1368_;
  assign new_n985_ = new_n1372_ & new_n777_;
  assign new_n986_ = new_n1380_ & new_n776_;
  assign new_n987_ = new_n986_ | new_n985_;
  assign new_n988_ = new_n812_ & new_n735_;
  assign new_n989_ = new_n988_ & new_n987_;
  assign new_n990_ = new_n1372_ & new_n779_;
  assign new_n991_ = new_n1380_ & new_n778_;
  assign new_n992_ = new_n991_ | new_n990_;
  assign new_n993_ = new_n814_ & new_n737_;
  assign new_n994_ = new_n993_ & new_n992_;
  assign new_n995_ = new_n1371_ & new_n781_;
  assign new_n996_ = new_n1381_ & new_n780_;
  assign new_n997_ = new_n996_ | new_n995_;
  assign new_n998_ = new_n816_ & new_n739_;
  assign new_n999_ = new_n998_ & new_n997_;
  assign new_n1000_ = new_n1373_ & new_n783_;
  assign new_n1001_ = new_n1381_ & new_n782_;
  assign new_n1002_ = new_n1001_ | new_n1000_;
  assign new_n1003_ = new_n818_ & new_n741_;
  assign new_n1004_ = new_n1003_ & new_n1002_;
  assign new_n1005_ = new_n1373_ & new_n785_;
  assign new_n1006_ = new_n1383_ & new_n784_;
  assign new_n1007_ = new_n1006_ | new_n1005_;
  assign new_n1008_ = new_n820_ & new_n743_;
  assign new_n1009_ = new_n1008_ & new_n1007_;
  assign new_n1010_ = new_n1375_ & new_n787_;
  assign new_n1011_ = new_n1383_ & new_n786_;
  assign new_n1012_ = new_n1011_ | new_n1010_;
  assign new_n1013_ = new_n822_ & new_n745_;
  assign new_n1014_ = new_n1013_ & new_n1012_;
  assign new_n1015_ = new_n1375_ & new_n789_;
  assign new_n1016_ = new_n1382_ & new_n788_;
  assign new_n1017_ = new_n1016_ | new_n1015_;
  assign new_n1018_ = new_n824_ & new_n747_;
  assign new_n1019_ = new_n1018_ & new_n1017_;
  assign new_n1020_ = new_n1376_ & new_n791_;
  assign new_n1021_ = new_n1385_ & new_n790_;
  assign new_n1022_ = new_n1021_ | new_n1020_;
  assign new_n1023_ = new_n826_ & new_n749_;
  assign new_n1024_ = new_n1023_ & new_n1022_;
  assign new_n1025_ = new_n1376_ & new_n793_;
  assign new_n1026_ = new_n1385_ & new_n792_;
  assign new_n1027_ = new_n1026_ | new_n1025_;
  assign new_n1028_ = new_n828_ & new_n751_;
  assign new_n1029_ = new_n1028_ & new_n1027_;
  assign new_n1030_ = new_n994_ | new_n989_;
  assign new_n1031_ = new_n1030_ | new_n999_;
  assign new_n1032_ = new_n1031_ | new_n1004_;
  assign new_n1033_ = new_n1032_ | new_n1009_;
  assign new_n1034_ = new_n1033_ | new_n1014_;
  assign new_n1035_ = new_n1034_ | new_n1019_;
  assign new_n1036_ = new_n1035_ | new_n1024_;
  assign new_n1037_ = new_n1036_ | new_n1029_;
  assign new_n1038_ = new_n1390_ & new_n1352_;
  assign new_n1039_ = new_n1398_ & new_n1354_;
  assign new_n1040_ = new_n1039_ | new_n1038_;
  assign new_n1041_ = new_n1390_ & new_n1351_;
  assign new_n1042_ = new_n1398_ & new_n1353_;
  assign new_n1043_ = new_n1042_ | new_n1041_;
  assign new_n1044_ = new_n1389_ & new_n1355_;
  assign new_n1045_ = new_n1399_ & new_n1356_;
  assign new_n1046_ = new_n1045_ | new_n1044_;
  assign new_n1047_ = new_n1391_ & new_n1357_;
  assign new_n1048_ = new_n1399_ & new_n1358_;
  assign new_n1049_ = new_n1048_ | new_n1047_;
  assign new_n1050_ = new_n1391_ & new_n1359_;
  assign new_n1051_ = new_n1400_ & new_n1360_;
  assign new_n1052_ = new_n1051_ | new_n1050_;
  assign new_n1053_ = new_n1393_ & new_n1361_;
  assign new_n1054_ = new_n1400_ & new_n1362_;
  assign new_n1055_ = new_n1054_ | new_n1053_;
  assign new_n1056_ = new_n1393_ & new_n1363_;
  assign new_n1057_ = new_n1402_ & new_n1364_;
  assign new_n1058_ = new_n1057_ | new_n1056_;
  assign new_n1059_ = new_n1394_ & new_n1365_;
  assign new_n1060_ = new_n1402_ & new_n1366_;
  assign new_n1061_ = new_n1060_ | new_n1059_;
  assign new_n1062_ = new_n1394_ & new_n1367_;
  assign new_n1063_ = new_n1403_ & new_n1368_;
  assign new_n1064_ = new_n1063_ | new_n1062_;
  assign new_n1065_ = new_n1405_ & new_n503_;
  assign new_n1066_ = new_n1065_ & new_n1406_;
  assign new_n1067_ = new_n1408_ & new_n523_;
  assign new_n1068_ = new_n1067_ & new_n1409_;
  assign new_n1069_ = new_n1411_ & new_n543_;
  assign new_n1070_ = new_n1069_ & new_n1412_;
  assign new_n1071_ = new_n1414_ & new_n563_;
  assign new_n1072_ = new_n1071_ & new_n1415_;
  assign new_n1073_ = new_n1417_ & new_n583_;
  assign new_n1074_ = new_n1073_ & new_n1418_;
  assign new_n1075_ = new_n1420_ & new_n603_;
  assign new_n1076_ = new_n1075_ & new_n1421_;
  assign new_n1077_ = new_n1423_ & new_n623_;
  assign new_n1078_ = new_n1077_ & new_n1424_;
  assign new_n1079_ = new_n1426_ & new_n643_;
  assign new_n1080_ = new_n1079_ & new_n1427_;
  assign new_n1081_ = new_n1429_ & new_n663_;
  assign new_n1082_ = new_n1081_ & new_n1430_;
  assign new_n1083_ = new_n1405_ & new_n513_;
  assign new_n1084_ = new_n1408_ & new_n533_;
  assign new_n1085_ = new_n1411_ & new_n553_;
  assign new_n1086_ = new_n1414_ & new_n573_;
  assign new_n1087_ = new_n1417_ & new_n593_;
  assign new_n1088_ = new_n1420_ & new_n613_;
  assign new_n1089_ = new_n1423_ & new_n633_;
  assign new_n1090_ = new_n1426_ & new_n653_;
  assign new_n1091_ = new_n1429_ & new_n669_;
  assign new_n1092_ = new_n1431_ | new_n1432_;
  assign new_n1093_ = new_n1092_ | new_n1433_;
  assign new_n1094_ = new_n1093_ | new_n1434_;
  assign new_n1095_ = new_n1094_ | new_n1435_;
  assign new_n1096_ = new_n1095_ | new_n1436_;
  assign new_n1097_ = new_n1096_ | new_n1437_;
  assign new_n1098_ = new_n1097_ | new_n1438_;
  assign new_n1099_ = new_n1098_ | new_n1439_;
  assign new_n1100_ = new_n1440_ & new_n493_;
  assign new_n1101_ = new_n1441_ & new_n507_;
  assign new_n1102_ = new_n1442_ & new_n527_;
  assign new_n1103_ = new_n1443_ & new_n547_;
  assign new_n1104_ = new_n1444_ & new_n567_;
  assign new_n1105_ = new_n1445_ & new_n587_;
  assign new_n1106_ = new_n1446_ & new_n607_;
  assign new_n1107_ = new_n1447_ & new_n627_;
  assign new_n1108_ = new_n1448_ & new_n647_;
  assign G426 = new_n672_;
  assign G427 = new_n674_;
  assign G428 = new_n732_;
  assign G429 = ~new_n953_;
  assign G430 = ~new_n956_;
  assign G431 = ~new_n963_;
  assign G432 = ~new_n968_;
  assign n205_li = new_n420_;
  assign n214_li = new_n676_;
  assign n217_li = new_n422_;
  assign n226_li = new_n694_;
  assign n229_li = new_n424_;
  assign n232_li = new_n500_;
  assign n238_li = new_n714_;
  assign n241_li = new_n426_;
  assign n250_li = new_n678_;
  assign n253_li = new_n428_;
  assign n256_li = new_n510_;
  assign n262_li = new_n752_;
  assign n265_li = new_n430_;
  assign n274_li = new_n696_;
  assign n277_li = new_n432_;
  assign n280_li = new_n520_;
  assign n286_li = new_n716_;
  assign n289_li = new_n434_;
  assign n298_li = new_n680_;
  assign n301_li = new_n436_;
  assign n304_li = new_n530_;
  assign n310_li = new_n754_;
  assign n313_li = new_n438_;
  assign n322_li = new_n698_;
  assign n325_li = new_n440_;
  assign n328_li = new_n540_;
  assign n334_li = new_n718_;
  assign n337_li = new_n442_;
  assign n346_li = new_n682_;
  assign n349_li = new_n444_;
  assign n352_li = new_n550_;
  assign n358_li = new_n756_;
  assign n361_li = new_n446_;
  assign n370_li = new_n700_;
  assign n373_li = new_n448_;
  assign n376_li = new_n560_;
  assign n382_li = new_n720_;
  assign n385_li = new_n450_;
  assign n394_li = new_n684_;
  assign n397_li = new_n452_;
  assign n400_li = new_n570_;
  assign n406_li = new_n758_;
  assign n409_li = new_n454_;
  assign n418_li = new_n702_;
  assign n421_li = new_n456_;
  assign n424_li = new_n580_;
  assign n430_li = new_n722_;
  assign n433_li = new_n458_;
  assign n442_li = new_n686_;
  assign n445_li = new_n460_;
  assign n448_li = new_n590_;
  assign n454_li = new_n760_;
  assign n457_li = new_n462_;
  assign n466_li = new_n704_;
  assign n469_li = new_n464_;
  assign n472_li = new_n600_;
  assign n478_li = new_n724_;
  assign n481_li = new_n466_;
  assign n490_li = new_n688_;
  assign n493_li = new_n468_;
  assign n496_li = new_n610_;
  assign n502_li = new_n762_;
  assign n505_li = new_n470_;
  assign n514_li = new_n706_;
  assign n517_li = new_n472_;
  assign n520_li = new_n620_;
  assign n526_li = new_n726_;
  assign n529_li = new_n474_;
  assign n538_li = new_n690_;
  assign n541_li = new_n476_;
  assign n544_li = new_n630_;
  assign n550_li = new_n764_;
  assign n553_li = new_n478_;
  assign n562_li = new_n708_;
  assign n565_li = new_n480_;
  assign n568_li = new_n640_;
  assign n574_li = new_n728_;
  assign n577_li = new_n482_;
  assign n586_li = new_n692_;
  assign n589_li = new_n484_;
  assign n592_li = new_n650_;
  assign n598_li = new_n766_;
  assign n601_li = new_n486_;
  assign n610_li = new_n710_;
  assign n613_li = new_n488_;
  assign n616_li = new_n660_;
  assign n622_li = new_n730_;
  assign n625_li = new_n490_;
  assign n628_li = new_n666_;
  assign n634_li = new_n768_;
  assign n919_i2 = new_n1449_;
  assign n1024_i2 = new_n1386_;
  assign n997_i2 = new_n794_;
  assign n998_i2 = new_n796_;
  assign n999_i2 = new_n798_;
  assign n1000_i2 = new_n800_;
  assign n1001_i2 = new_n802_;
  assign n1002_i2 = new_n804_;
  assign n1003_i2 = new_n806_;
  assign n1004_i2 = new_n808_;
  assign n1005_i2 = new_n810_;
  assign n1015_i2 = new_n1404_;
  assign n1016_i2 = new_n1407_;
  assign n1017_i2 = new_n1410_;
  assign n1018_i2 = new_n1413_;
  assign n1019_i2 = new_n1416_;
  assign n1020_i2 = new_n1419_;
  assign n1021_i2 = new_n1422_;
  assign n1022_i2 = new_n1425_;
  assign n1023_i2 = new_n1428_;
  assign G199_i2 = new_n1403_;
  assign n235_lo_buf_i2 = new_n502_;
  assign n283_lo_buf_i2 = new_n522_;
  assign n331_lo_buf_i2 = new_n542_;
  assign n379_lo_buf_i2 = new_n562_;
  assign n427_lo_buf_i2 = new_n582_;
  assign n475_lo_buf_i2 = new_n602_;
  assign n523_lo_buf_i2 = new_n622_;
  assign n571_lo_buf_i2 = new_n642_;
  assign n619_lo_buf_i2 = new_n662_;
  assign G355_i2 = new_n1450_;
  assign G223_i2 = ~new_n1406_;
  assign G226_i2 = ~new_n1409_;
  assign G229_i2 = ~new_n1412_;
  assign G232_i2 = ~new_n1415_;
  assign G235_i2 = ~new_n1418_;
  assign G238_i2 = ~new_n1421_;
  assign G242_i2 = ~new_n1424_;
  assign G246_i2 = ~new_n1427_;
  assign G250_i2 = ~new_n1430_;
  assign n259_lo_buf_i2 = new_n512_;
  assign n307_lo_buf_i2 = new_n532_;
  assign n355_lo_buf_i2 = new_n552_;
  assign n403_lo_buf_i2 = new_n572_;
  assign n451_lo_buf_i2 = new_n592_;
  assign n499_lo_buf_i2 = new_n612_;
  assign n547_lo_buf_i2 = new_n632_;
  assign n595_lo_buf_i2 = new_n652_;
  assign n631_lo_buf_i2 = new_n668_;
  assign G213_i2 = n919_i2;
  assign G318_i2 = n1024_i2;
  assign G358_i2 = G355_i2;
  assign G259_i2 = new_n1432_;
  assign G263_i2 = new_n1431_;
  assign G266_i2 = new_n1433_;
  assign G269_i2 = new_n1434_;
  assign G272_i2 = new_n1435_;
  assign G275_i2 = new_n1436_;
  assign G278_i2 = new_n1437_;
  assign G281_i2 = new_n1438_;
  assign G284_i2 = new_n1439_;
  assign n211_lo_buf_i2 = new_n492_;
  assign n247_lo_buf_i2 = new_n506_;
  assign n295_lo_buf_i2 = new_n526_;
  assign n343_lo_buf_i2 = new_n546_;
  assign n391_lo_buf_i2 = new_n566_;
  assign n439_lo_buf_i2 = new_n586_;
  assign n487_lo_buf_i2 = new_n606_;
  assign n535_lo_buf_i2 = new_n626_;
  assign n583_lo_buf_i2 = new_n646_;
  assign G158_i2 = new_n1083_;
  assign G184_i2 = new_n1084_;
  assign G186_i2 = new_n1085_;
  assign G188_i2 = new_n1086_;
  assign G190_i2 = new_n1087_;
  assign G192_i2 = new_n1088_;
  assign G194_i2 = new_n1089_;
  assign G196_i2 = new_n1090_;
  assign G198_i2 = new_n1091_;
  assign n223_lo_buf_i2 = new_n1440_;
  assign n271_lo_buf_i2 = new_n1441_;
  assign n319_lo_buf_i2 = new_n1442_;
  assign n367_lo_buf_i2 = new_n1443_;
  assign n415_lo_buf_i2 = new_n1444_;
  assign n463_lo_buf_i2 = new_n1445_;
  assign n511_lo_buf_i2 = new_n1446_;
  assign n559_lo_buf_i2 = new_n1447_;
  assign n607_lo_buf_i2 = new_n1448_;
  assign G295_i2 = new_n1099_;
  assign G154_i2 = new_n1100_;
  assign G159_i2 = new_n1101_;
  assign G162_i2 = new_n1102_;
  assign G165_i2 = new_n1103_;
  assign G168_i2 = new_n1104_;
  assign G171_i2 = new_n1105_;
  assign G174_i2 = new_n1106_;
  assign G177_i2 = new_n1107_;
  assign G180_i2 = new_n1108_;
  assign new_n1304_ = new_n771_;
  assign new_n1305_ = new_n1304_;
  assign new_n1306_ = new_n1305_;
  assign new_n1307_ = new_n1304_;
  assign new_n1308_ = new_n773_;
  assign new_n1309_ = new_n1308_;
  assign new_n1310_ = new_n1309_;
  assign new_n1311_ = new_n1308_;
  assign new_n1312_ = new_n775_;
  assign new_n1313_ = new_n1312_;
  assign new_n1314_ = new_n1313_;
  assign new_n1315_ = new_n1312_;
  assign new_n1316_ = new_n770_;
  assign new_n1317_ = new_n1316_;
  assign new_n1318_ = new_n1317_;
  assign new_n1319_ = new_n1317_;
  assign new_n1320_ = new_n1316_;
  assign new_n1321_ = new_n1320_;
  assign new_n1322_ = new_n1320_;
  assign new_n1323_ = new_n772_;
  assign new_n1324_ = new_n1323_;
  assign new_n1325_ = new_n1324_;
  assign new_n1326_ = new_n1324_;
  assign new_n1327_ = new_n1323_;
  assign new_n1328_ = new_n1327_;
  assign new_n1329_ = new_n1327_;
  assign new_n1330_ = new_n774_;
  assign new_n1331_ = new_n1330_;
  assign new_n1332_ = new_n1331_;
  assign new_n1333_ = new_n1331_;
  assign new_n1334_ = new_n1330_;
  assign new_n1335_ = new_n1334_;
  assign new_n1336_ = new_n1334_;
  assign new_n1337_ = new_n879_;
  assign new_n1338_ = new_n946_;
  assign new_n1339_ = new_n1338_;
  assign new_n1340_ = new_n903_;
  assign new_n1341_ = new_n915_;
  assign new_n1342_ = new_n921_;
  assign new_n1343_ = new_n933_;
  assign new_n1344_ = new_n939_;
  assign new_n1345_ = new_n890_;
  assign new_n1346_ = new_n954_;
  assign new_n1347_ = new_n902_;
  assign new_n1348_ = new_n957_;
  assign new_n1349_ = new_n914_;
  assign new_n1350_ = new_n959_;
  assign new_n1351_ = new_n853_;
  assign new_n1352_ = new_n851_;
  assign new_n1353_ = new_n852_;
  assign new_n1354_ = new_n850_;
  assign new_n1355_ = new_n855_;
  assign new_n1356_ = new_n854_;
  assign new_n1357_ = new_n857_;
  assign new_n1358_ = new_n856_;
  assign new_n1359_ = new_n859_;
  assign new_n1360_ = new_n858_;
  assign new_n1361_ = new_n861_;
  assign new_n1362_ = new_n860_;
  assign new_n1363_ = new_n863_;
  assign new_n1364_ = new_n862_;
  assign new_n1365_ = new_n865_;
  assign new_n1366_ = new_n864_;
  assign new_n1367_ = new_n867_;
  assign new_n1368_ = new_n866_;
  assign new_n1369_ = new_n849_;
  assign new_n1370_ = new_n1369_;
  assign new_n1371_ = new_n1370_;
  assign new_n1372_ = new_n1371_;
  assign new_n1373_ = new_n1370_;
  assign new_n1374_ = new_n1369_;
  assign new_n1375_ = new_n1374_;
  assign new_n1376_ = new_n1374_;
  assign new_n1377_ = new_n848_;
  assign new_n1378_ = new_n1377_;
  assign new_n1379_ = new_n1378_;
  assign new_n1380_ = new_n1379_;
  assign new_n1381_ = new_n1379_;
  assign new_n1382_ = new_n1378_;
  assign new_n1383_ = new_n1382_;
  assign new_n1384_ = new_n1377_;
  assign new_n1385_ = new_n1384_;
  assign new_n1386_ = new_n1384_;
  assign new_n1387_ = new_n983_;
  assign new_n1388_ = new_n1387_;
  assign new_n1389_ = new_n1388_;
  assign new_n1390_ = new_n1389_;
  assign new_n1391_ = new_n1388_;
  assign new_n1392_ = new_n1387_;
  assign new_n1393_ = new_n1392_;
  assign new_n1394_ = new_n1392_;
  assign new_n1395_ = new_n984_;
  assign new_n1396_ = new_n1395_;
  assign new_n1397_ = new_n1396_;
  assign new_n1398_ = new_n1397_;
  assign new_n1399_ = new_n1397_;
  assign new_n1400_ = new_n1396_;
  assign new_n1401_ = new_n1395_;
  assign new_n1402_ = new_n1401_;
  assign new_n1403_ = new_n1401_;
  assign new_n1404_ = new_n830_;
  assign new_n1405_ = new_n1404_;
  assign new_n1406_ = new_n1040_;
  assign new_n1407_ = new_n832_;
  assign new_n1408_ = new_n1407_;
  assign new_n1409_ = new_n1043_;
  assign new_n1410_ = new_n834_;
  assign new_n1411_ = new_n1410_;
  assign new_n1412_ = new_n1046_;
  assign new_n1413_ = new_n836_;
  assign new_n1414_ = new_n1413_;
  assign new_n1415_ = new_n1049_;
  assign new_n1416_ = new_n838_;
  assign new_n1417_ = new_n1416_;
  assign new_n1418_ = new_n1052_;
  assign new_n1419_ = new_n840_;
  assign new_n1420_ = new_n1419_;
  assign new_n1421_ = new_n1055_;
  assign new_n1422_ = new_n842_;
  assign new_n1423_ = new_n1422_;
  assign new_n1424_ = new_n1058_;
  assign new_n1425_ = new_n844_;
  assign new_n1426_ = new_n1425_;
  assign new_n1427_ = new_n1061_;
  assign new_n1428_ = new_n846_;
  assign new_n1429_ = new_n1428_;
  assign new_n1430_ = new_n1064_;
  assign new_n1431_ = new_n1068_;
  assign new_n1432_ = new_n1066_;
  assign new_n1433_ = new_n1070_;
  assign new_n1434_ = new_n1072_;
  assign new_n1435_ = new_n1074_;
  assign new_n1436_ = new_n1076_;
  assign new_n1437_ = new_n1078_;
  assign new_n1438_ = new_n1080_;
  assign new_n1439_ = new_n1082_;
  assign new_n1440_ = new_n496_;
  assign new_n1441_ = new_n516_;
  assign new_n1442_ = new_n536_;
  assign new_n1443_ = new_n556_;
  assign new_n1444_ = new_n576_;
  assign new_n1445_ = new_n596_;
  assign new_n1446_ = new_n616_;
  assign new_n1447_ = new_n636_;
  assign new_n1448_ = new_n656_;
  assign new_n1449_ = new_n712_;
  assign new_n1450_ = new_n1037_;
  always @ (posedge clock) begin
    n205_lo <= n205_li;
    n214_lo <= n214_li;
    n217_lo <= n217_li;
    n226_lo <= n226_li;
    n229_lo <= n229_li;
    n232_lo <= n232_li;
    n238_lo <= n238_li;
    n241_lo <= n241_li;
    n250_lo <= n250_li;
    n253_lo <= n253_li;
    n256_lo <= n256_li;
    n262_lo <= n262_li;
    n265_lo <= n265_li;
    n274_lo <= n274_li;
    n277_lo <= n277_li;
    n280_lo <= n280_li;
    n286_lo <= n286_li;
    n289_lo <= n289_li;
    n298_lo <= n298_li;
    n301_lo <= n301_li;
    n304_lo <= n304_li;
    n310_lo <= n310_li;
    n313_lo <= n313_li;
    n322_lo <= n322_li;
    n325_lo <= n325_li;
    n328_lo <= n328_li;
    n334_lo <= n334_li;
    n337_lo <= n337_li;
    n346_lo <= n346_li;
    n349_lo <= n349_li;
    n352_lo <= n352_li;
    n358_lo <= n358_li;
    n361_lo <= n361_li;
    n370_lo <= n370_li;
    n373_lo <= n373_li;
    n376_lo <= n376_li;
    n382_lo <= n382_li;
    n385_lo <= n385_li;
    n394_lo <= n394_li;
    n397_lo <= n397_li;
    n400_lo <= n400_li;
    n406_lo <= n406_li;
    n409_lo <= n409_li;
    n418_lo <= n418_li;
    n421_lo <= n421_li;
    n424_lo <= n424_li;
    n430_lo <= n430_li;
    n433_lo <= n433_li;
    n442_lo <= n442_li;
    n445_lo <= n445_li;
    n448_lo <= n448_li;
    n454_lo <= n454_li;
    n457_lo <= n457_li;
    n466_lo <= n466_li;
    n469_lo <= n469_li;
    n472_lo <= n472_li;
    n478_lo <= n478_li;
    n481_lo <= n481_li;
    n490_lo <= n490_li;
    n493_lo <= n493_li;
    n496_lo <= n496_li;
    n502_lo <= n502_li;
    n505_lo <= n505_li;
    n514_lo <= n514_li;
    n517_lo <= n517_li;
    n520_lo <= n520_li;
    n526_lo <= n526_li;
    n529_lo <= n529_li;
    n538_lo <= n538_li;
    n541_lo <= n541_li;
    n544_lo <= n544_li;
    n550_lo <= n550_li;
    n553_lo <= n553_li;
    n562_lo <= n562_li;
    n565_lo <= n565_li;
    n568_lo <= n568_li;
    n574_lo <= n574_li;
    n577_lo <= n577_li;
    n586_lo <= n586_li;
    n589_lo <= n589_li;
    n592_lo <= n592_li;
    n598_lo <= n598_li;
    n601_lo <= n601_li;
    n610_lo <= n610_li;
    n613_lo <= n613_li;
    n616_lo <= n616_li;
    n622_lo <= n622_li;
    n625_lo <= n625_li;
    n628_lo <= n628_li;
    n634_lo <= n634_li;
    n316_inv <= n919_i2;
    n319_inv <= n1024_i2;
    n997_o2 <= n997_i2;
    n998_o2 <= n998_i2;
    n999_o2 <= n999_i2;
    n1000_o2 <= n1000_i2;
    n1001_o2 <= n1001_i2;
    n1002_o2 <= n1002_i2;
    n1003_o2 <= n1003_i2;
    n1004_o2 <= n1004_i2;
    n1005_o2 <= n1005_i2;
    n1015_o2 <= n1015_i2;
    n1016_o2 <= n1016_i2;
    n1017_o2 <= n1017_i2;
    n1018_o2 <= n1018_i2;
    n1019_o2 <= n1019_i2;
    n1020_o2 <= n1020_i2;
    n1021_o2 <= n1021_i2;
    n1022_o2 <= n1022_i2;
    n1023_o2 <= n1023_i2;
    n376_1_inv <= G199_i2;
    n235_lo_buf_o2 <= n235_lo_buf_i2;
    n283_lo_buf_o2 <= n283_lo_buf_i2;
    n331_lo_buf_o2 <= n331_lo_buf_i2;
    n379_lo_buf_o2 <= n379_lo_buf_i2;
    n427_lo_buf_o2 <= n427_lo_buf_i2;
    n475_lo_buf_o2 <= n475_lo_buf_i2;
    n523_lo_buf_o2 <= n523_lo_buf_i2;
    n571_lo_buf_o2 <= n571_lo_buf_i2;
    n619_lo_buf_o2 <= n619_lo_buf_i2;
    n406_1_inv <= G355_i2;
    G223_o2 <= G223_i2;
    G226_o2 <= G226_i2;
    G229_o2 <= G229_i2;
    G232_o2 <= G232_i2;
    G235_o2 <= G235_i2;
    G238_o2 <= G238_i2;
    G242_o2 <= G242_i2;
    G246_o2 <= G246_i2;
    G250_o2 <= G250_i2;
    n259_lo_buf_o2 <= n259_lo_buf_i2;
    n307_lo_buf_o2 <= n307_lo_buf_i2;
    n355_lo_buf_o2 <= n355_lo_buf_i2;
    n403_lo_buf_o2 <= n403_lo_buf_i2;
    n451_lo_buf_o2 <= n451_lo_buf_i2;
    n499_lo_buf_o2 <= n499_lo_buf_i2;
    n547_lo_buf_o2 <= n547_lo_buf_i2;
    n595_lo_buf_o2 <= n595_lo_buf_i2;
    n631_lo_buf_o2 <= n631_lo_buf_i2;
    G213_o2 <= G213_i2;
    G318_o2 <= G318_i2;
    G358_o2 <= G358_i2;
    G259_o2 <= G259_i2;
    G263_o2 <= G263_i2;
    G266_o2 <= G266_i2;
    G269_o2 <= G269_i2;
    G272_o2 <= G272_i2;
    G275_o2 <= G275_i2;
    G278_o2 <= G278_i2;
    G281_o2 <= G281_i2;
    G284_o2 <= G284_i2;
    n211_lo_buf_o2 <= n211_lo_buf_i2;
    n247_lo_buf_o2 <= n247_lo_buf_i2;
    n295_lo_buf_o2 <= n295_lo_buf_i2;
    n343_lo_buf_o2 <= n343_lo_buf_i2;
    n391_lo_buf_o2 <= n391_lo_buf_i2;
    n439_lo_buf_o2 <= n439_lo_buf_i2;
    n487_lo_buf_o2 <= n487_lo_buf_i2;
    n535_lo_buf_o2 <= n535_lo_buf_i2;
    n583_lo_buf_o2 <= n583_lo_buf_i2;
    G158_o2 <= G158_i2;
    G184_o2 <= G184_i2;
    G186_o2 <= G186_i2;
    G188_o2 <= G188_i2;
    G190_o2 <= G190_i2;
    G192_o2 <= G192_i2;
    G194_o2 <= G194_i2;
    G196_o2 <= G196_i2;
    G198_o2 <= G198_i2;
    n223_lo_buf_o2 <= n223_lo_buf_i2;
    n271_lo_buf_o2 <= n271_lo_buf_i2;
    n319_lo_buf_o2 <= n319_lo_buf_i2;
    n367_lo_buf_o2 <= n367_lo_buf_i2;
    n415_lo_buf_o2 <= n415_lo_buf_i2;
    n463_lo_buf_o2 <= n463_lo_buf_i2;
    n511_lo_buf_o2 <= n511_lo_buf_i2;
    n559_lo_buf_o2 <= n559_lo_buf_i2;
    n607_lo_buf_o2 <= n607_lo_buf_i2;
    n580_inv <= G295_i2;
    G154_o2 <= G154_i2;
    G159_o2 <= G159_i2;
    G162_o2 <= G162_i2;
    G165_o2 <= G165_i2;
    G168_o2 <= G168_i2;
    G171_o2 <= G171_i2;
    G174_o2 <= G174_i2;
    G177_o2 <= G177_i2;
    G180_o2 <= G180_i2;
  end
  initial begin
    n205_lo <= 1'b0;
    n214_lo <= 1'b0;
    n217_lo <= 1'b0;
    n226_lo <= 1'b0;
    n229_lo <= 1'b0;
    n232_lo <= 1'b0;
    n238_lo <= 1'b0;
    n241_lo <= 1'b0;
    n250_lo <= 1'b0;
    n253_lo <= 1'b0;
    n256_lo <= 1'b0;
    n262_lo <= 1'b0;
    n265_lo <= 1'b0;
    n274_lo <= 1'b0;
    n277_lo <= 1'b0;
    n280_lo <= 1'b0;
    n286_lo <= 1'b0;
    n289_lo <= 1'b0;
    n298_lo <= 1'b0;
    n301_lo <= 1'b0;
    n304_lo <= 1'b0;
    n310_lo <= 1'b0;
    n313_lo <= 1'b0;
    n322_lo <= 1'b0;
    n325_lo <= 1'b0;
    n328_lo <= 1'b0;
    n334_lo <= 1'b0;
    n337_lo <= 1'b0;
    n346_lo <= 1'b0;
    n349_lo <= 1'b0;
    n352_lo <= 1'b0;
    n358_lo <= 1'b0;
    n361_lo <= 1'b0;
    n370_lo <= 1'b0;
    n373_lo <= 1'b0;
    n376_lo <= 1'b0;
    n382_lo <= 1'b0;
    n385_lo <= 1'b0;
    n394_lo <= 1'b0;
    n397_lo <= 1'b0;
    n400_lo <= 1'b0;
    n406_lo <= 1'b0;
    n409_lo <= 1'b0;
    n418_lo <= 1'b0;
    n421_lo <= 1'b0;
    n424_lo <= 1'b0;
    n430_lo <= 1'b0;
    n433_lo <= 1'b0;
    n442_lo <= 1'b0;
    n445_lo <= 1'b0;
    n448_lo <= 1'b0;
    n454_lo <= 1'b0;
    n457_lo <= 1'b0;
    n466_lo <= 1'b0;
    n469_lo <= 1'b0;
    n472_lo <= 1'b0;
    n478_lo <= 1'b0;
    n481_lo <= 1'b0;
    n490_lo <= 1'b0;
    n493_lo <= 1'b0;
    n496_lo <= 1'b0;
    n502_lo <= 1'b0;
    n505_lo <= 1'b0;
    n514_lo <= 1'b0;
    n517_lo <= 1'b0;
    n520_lo <= 1'b0;
    n526_lo <= 1'b0;
    n529_lo <= 1'b0;
    n538_lo <= 1'b0;
    n541_lo <= 1'b0;
    n544_lo <= 1'b0;
    n550_lo <= 1'b0;
    n553_lo <= 1'b0;
    n562_lo <= 1'b0;
    n565_lo <= 1'b0;
    n568_lo <= 1'b0;
    n574_lo <= 1'b0;
    n577_lo <= 1'b0;
    n586_lo <= 1'b0;
    n589_lo <= 1'b0;
    n592_lo <= 1'b0;
    n598_lo <= 1'b0;
    n601_lo <= 1'b0;
    n610_lo <= 1'b0;
    n613_lo <= 1'b0;
    n616_lo <= 1'b0;
    n622_lo <= 1'b0;
    n625_lo <= 1'b0;
    n628_lo <= 1'b0;
    n634_lo <= 1'b0;
    n316_inv <= 1'b0;
    n319_inv <= 1'b0;
    n997_o2 <= 1'b0;
    n998_o2 <= 1'b0;
    n999_o2 <= 1'b0;
    n1000_o2 <= 1'b0;
    n1001_o2 <= 1'b0;
    n1002_o2 <= 1'b0;
    n1003_o2 <= 1'b0;
    n1004_o2 <= 1'b0;
    n1005_o2 <= 1'b0;
    n1015_o2 <= 1'b0;
    n1016_o2 <= 1'b0;
    n1017_o2 <= 1'b0;
    n1018_o2 <= 1'b0;
    n1019_o2 <= 1'b0;
    n1020_o2 <= 1'b0;
    n1021_o2 <= 1'b0;
    n1022_o2 <= 1'b0;
    n1023_o2 <= 1'b0;
    n376_1_inv <= 1'b0;
    n235_lo_buf_o2 <= 1'b0;
    n283_lo_buf_o2 <= 1'b0;
    n331_lo_buf_o2 <= 1'b0;
    n379_lo_buf_o2 <= 1'b0;
    n427_lo_buf_o2 <= 1'b0;
    n475_lo_buf_o2 <= 1'b0;
    n523_lo_buf_o2 <= 1'b0;
    n571_lo_buf_o2 <= 1'b0;
    n619_lo_buf_o2 <= 1'b0;
    n406_1_inv <= 1'b0;
    G223_o2 <= 1'b0;
    G226_o2 <= 1'b0;
    G229_o2 <= 1'b0;
    G232_o2 <= 1'b0;
    G235_o2 <= 1'b0;
    G238_o2 <= 1'b0;
    G242_o2 <= 1'b0;
    G246_o2 <= 1'b0;
    G250_o2 <= 1'b0;
    n259_lo_buf_o2 <= 1'b0;
    n307_lo_buf_o2 <= 1'b0;
    n355_lo_buf_o2 <= 1'b0;
    n403_lo_buf_o2 <= 1'b0;
    n451_lo_buf_o2 <= 1'b0;
    n499_lo_buf_o2 <= 1'b0;
    n547_lo_buf_o2 <= 1'b0;
    n595_lo_buf_o2 <= 1'b0;
    n631_lo_buf_o2 <= 1'b0;
    G213_o2 <= 1'b0;
    G318_o2 <= 1'b0;
    G358_o2 <= 1'b0;
    G259_o2 <= 1'b0;
    G263_o2 <= 1'b0;
    G266_o2 <= 1'b0;
    G269_o2 <= 1'b0;
    G272_o2 <= 1'b0;
    G275_o2 <= 1'b0;
    G278_o2 <= 1'b0;
    G281_o2 <= 1'b0;
    G284_o2 <= 1'b0;
    n211_lo_buf_o2 <= 1'b0;
    n247_lo_buf_o2 <= 1'b0;
    n295_lo_buf_o2 <= 1'b0;
    n343_lo_buf_o2 <= 1'b0;
    n391_lo_buf_o2 <= 1'b0;
    n439_lo_buf_o2 <= 1'b0;
    n487_lo_buf_o2 <= 1'b0;
    n535_lo_buf_o2 <= 1'b0;
    n583_lo_buf_o2 <= 1'b0;
    G158_o2 <= 1'b0;
    G184_o2 <= 1'b0;
    G186_o2 <= 1'b0;
    G188_o2 <= 1'b0;
    G190_o2 <= 1'b0;
    G192_o2 <= 1'b0;
    G194_o2 <= 1'b0;
    G196_o2 <= 1'b0;
    G198_o2 <= 1'b0;
    n223_lo_buf_o2 <= 1'b0;
    n271_lo_buf_o2 <= 1'b0;
    n319_lo_buf_o2 <= 1'b0;
    n367_lo_buf_o2 <= 1'b0;
    n415_lo_buf_o2 <= 1'b0;
    n463_lo_buf_o2 <= 1'b0;
    n511_lo_buf_o2 <= 1'b0;
    n559_lo_buf_o2 <= 1'b0;
    n607_lo_buf_o2 <= 1'b0;
    n580_inv <= 1'b0;
    G154_o2 <= 1'b0;
    G159_o2 <= 1'b0;
    G162_o2 <= 1'b0;
    G165_o2 <= 1'b0;
    G168_o2 <= 1'b0;
    G171_o2 <= 1'b0;
    G174_o2 <= 1'b0;
    G177_o2 <= 1'b0;
    G180_o2 <= 1'b0;
  end
endmodule


