
module mymod
(
  G1_p,
  G1_n,
  G2_p,
  G2_n,
  G3_p,
  G3_n,
  G4_p,
  G4_n,
  G5_p,
  G5_n,
  G6_p,
  G6_n,
  G7_p,
  G7_n,
  G8_p,
  G8_n,
  G9_p,
  G9_n,
  G10_p,
  G10_n,
  G11_p,
  G11_n,
  G12_p,
  G12_n,
  G13_p,
  G13_n,
  G14_p,
  G14_n,
  G15_p,
  G15_n,
  G16_p,
  G16_n,
  G17_p,
  G17_n,
  G18_p,
  G18_n,
  G19_p,
  G19_n,
  G20_p,
  G20_n,
  G21_p,
  G21_n,
  G22_p,
  G22_n,
  G23_p,
  G23_n,
  G24_p,
  G24_n,
  G25_p,
  G25_n,
  G26_p,
  G26_n,
  G27_p,
  G27_n,
  G28_p,
  G28_n,
  G29_p,
  G29_n,
  G30_p,
  G30_n,
  G31_p,
  G31_n,
  G32_p,
  G32_n,
  G33_p,
  G33_n,
  G1884_n,
  G1885_n,
  G1886_n,
  G1887_n,
  G1888_n,
  G1889_n,
  G1890_n,
  G1891_n,
  G1892_n,
  G1893_n,
  G1894_n,
  G1895_n,
  G1896_n,
  G1897_n,
  G1898_n,
  G1899_n,
  G1900_n,
  G1901_n,
  G1902_n,
  G1903_n,
  G1904_n,
  G1905_n,
  G1906_n,
  G1907_n,
  G1908_n
);

  input G1_p;input G1_n;input G2_p;input G2_n;input G3_p;input G3_n;input G4_p;input G4_n;input G5_p;input G5_n;input G6_p;input G6_n;input G7_p;input G7_n;input G8_p;input G8_n;input G9_p;input G9_n;input G10_p;input G10_n;input G11_p;input G11_n;input G12_p;input G12_n;input G13_p;input G13_n;input G14_p;input G14_n;input G15_p;input G15_n;input G16_p;input G16_n;input G17_p;input G17_n;input G18_p;input G18_n;input G19_p;input G19_n;input G20_p;input G20_n;input G21_p;input G21_n;input G22_p;input G22_n;input G23_p;input G23_n;input G24_p;input G24_n;input G25_p;input G25_n;input G26_p;input G26_n;input G27_p;input G27_n;input G28_p;input G28_n;input G29_p;input G29_n;input G30_p;input G30_n;input G31_p;input G31_n;input G32_p;input G32_n;input G33_p;input G33_n;
  output G1884_n;output G1885_n;output G1886_n;output G1887_n;output G1888_n;output G1889_n;output G1890_n;output G1891_n;output G1892_n;output G1893_n;output G1894_n;output G1895_n;output G1896_n;output G1897_n;output G1898_n;output G1899_n;output G1900_n;output G1901_n;output G1902_n;output G1903_n;output G1904_n;output G1905_n;output G1906_n;output G1907_n;output G1908_n;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire g34_p;
  wire g34_n;
  wire g35_p;
  wire g35_n;
  wire g36_p;
  wire g36_n;
  wire g37_p;
  wire g37_n;
  wire g38_p;
  wire g38_n;
  wire g39_p;
  wire g39_n;
  wire g40_p;
  wire g40_n;
  wire g41_p;
  wire g41_n;
  wire g42_p;
  wire g42_n;
  wire g43_p;
  wire g43_n;
  wire g44_p;
  wire g44_n;
  wire g45_p;
  wire g45_n;
  wire g46_p;
  wire g46_n;
  wire g47_p;
  wire g47_n;
  wire g48_p;
  wire g48_n;
  wire g49_p;
  wire g49_n;
  wire g50_p;
  wire g50_n;
  wire g51_p;
  wire g51_n;
  wire g52_p;
  wire g52_n;
  wire g53_p;
  wire g53_n;
  wire g54_p;
  wire g54_n;
  wire g55_p;
  wire g55_n;
  wire g56_p;
  wire g56_n;
  wire g57_p;
  wire g57_n;
  wire g58_p;
  wire g58_n;
  wire g59_p;
  wire g59_n;
  wire g60_p;
  wire g60_n;
  wire g61_p;
  wire g61_n;
  wire g62_p;
  wire g62_n;
  wire g63_p;
  wire g63_n;
  wire g64_p;
  wire g64_n;
  wire g65_p;
  wire g65_n;
  wire g66_p;
  wire g66_n;
  wire g67_p;
  wire g67_n;
  wire g68_p;
  wire g68_n;
  wire g69_p;
  wire g69_n;
  wire g70_p;
  wire g70_n;
  wire g71_p;
  wire g71_n;
  wire g72_p;
  wire g72_n;
  wire g73_p;
  wire g73_n;
  wire g74_p;
  wire g74_n;
  wire g75_p;
  wire g75_n;
  wire g76_p;
  wire g76_n;
  wire g77_p;
  wire g77_n;
  wire g78_p;
  wire g78_n;
  wire g79_p;
  wire g79_n;
  wire g80_p;
  wire g80_n;
  wire g81_p;
  wire g81_n;
  wire g82_p;
  wire g82_n;
  wire g83_p;
  wire g83_n;
  wire g84_p;
  wire g84_n;
  wire g85_p;
  wire g85_n;
  wire g86_p;
  wire g86_n;
  wire g87_p;
  wire g87_n;
  wire g88_p;
  wire g88_n;
  wire g89_p;
  wire g89_n;
  wire g90_p;
  wire g90_n;
  wire g91_p;
  wire g91_n;
  wire g92_p;
  wire g92_n;
  wire g93_p;
  wire g93_n;
  wire g94_p;
  wire g94_n;
  wire g95_p;
  wire g95_n;
  wire g96_p;
  wire g96_n;
  wire g97_p;
  wire g97_n;
  wire g98_p;
  wire g98_n;
  wire g99_p;
  wire g99_n;
  wire g100_p;
  wire g100_n;
  wire g101_p;
  wire g101_n;
  wire g102_p;
  wire g102_n;
  wire g103_p;
  wire g103_n;
  wire g104_p;
  wire g104_n;
  wire g105_p;
  wire g105_n;
  wire g106_p;
  wire g106_n;
  wire g107_p;
  wire g107_n;
  wire g108_p;
  wire g108_n;
  wire g109_p;
  wire g109_n;
  wire g110_p;
  wire g110_n;
  wire g111_p;
  wire g111_n;
  wire g112_p;
  wire g112_n;
  wire g113_p;
  wire g113_n;
  wire g114_p;
  wire g114_n;
  wire g115_p;
  wire g115_n;
  wire g116_p;
  wire g116_n;
  wire g117_p;
  wire g117_n;
  wire g118_p;
  wire g118_n;
  wire g119_p;
  wire g119_n;
  wire g120_p;
  wire g120_n;
  wire g121_p;
  wire g121_n;
  wire g122_p;
  wire g122_n;
  wire g123_p;
  wire g123_n;
  wire g124_p;
  wire g124_n;
  wire g125_p;
  wire g125_n;
  wire g126_p;
  wire g126_n;
  wire g127_p;
  wire g127_n;
  wire g128_p;
  wire g128_n;
  wire g129_p;
  wire g129_n;
  wire g130_p;
  wire g130_n;
  wire g131_p;
  wire g131_n;
  wire g132_p;
  wire g132_n;
  wire g133_p;
  wire g133_n;
  wire g134_p;
  wire g134_n;
  wire g135_p;
  wire g135_n;
  wire g136_p;
  wire g136_n;
  wire g137_p;
  wire g137_n;
  wire g138_p;
  wire g138_n;
  wire g139_p;
  wire g139_n;
  wire g140_p;
  wire g140_n;
  wire g141_p;
  wire g141_n;
  wire g142_p;
  wire g142_n;
  wire g143_p;
  wire g143_n;
  wire g144_p;
  wire g144_n;
  wire g145_p;
  wire g145_n;
  wire g146_p;
  wire g146_n;
  wire g147_p;
  wire g147_n;
  wire g148_p;
  wire g148_n;
  wire g149_p;
  wire g149_n;
  wire g150_p;
  wire g150_n;
  wire g151_p;
  wire g151_n;
  wire g152_p;
  wire g152_n;
  wire g153_p;
  wire g153_n;
  wire g154_p;
  wire g154_n;
  wire g155_p;
  wire g155_n;
  wire g156_p;
  wire g156_n;
  wire g157_p;
  wire g157_n;
  wire g158_p;
  wire g158_n;
  wire g159_p;
  wire g159_n;
  wire g160_p;
  wire g160_n;
  wire g161_p;
  wire g161_n;
  wire g162_p;
  wire g162_n;
  wire g163_p;
  wire g163_n;
  wire g164_p;
  wire g164_n;
  wire g165_p;
  wire g165_n;
  wire g166_p;
  wire g166_n;
  wire g167_p;
  wire g167_n;
  wire g168_p;
  wire g168_n;
  wire g169_p;
  wire g169_n;
  wire g170_p;
  wire g170_n;
  wire g171_p;
  wire g171_n;
  wire g172_p;
  wire g172_n;
  wire g173_p;
  wire g173_n;
  wire g174_p;
  wire g174_n;
  wire g175_p;
  wire g175_n;
  wire g176_p;
  wire g176_n;
  wire g177_p;
  wire g177_n;
  wire g178_p;
  wire g178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire G29_n_spl_;
  wire G33_n_spl_;
  wire G33_n_spl_0;
  wire G33_n_spl_00;
  wire G33_n_spl_000;
  wire G33_n_spl_001;
  wire G33_n_spl_01;
  wire G33_n_spl_010;
  wire G33_n_spl_011;
  wire G33_n_spl_1;
  wire G33_n_spl_10;
  wire G33_n_spl_11;
  wire G29_p_spl_;
  wire G33_p_spl_;
  wire G33_p_spl_0;
  wire G33_p_spl_00;
  wire G33_p_spl_000;
  wire G33_p_spl_001;
  wire G33_p_spl_01;
  wire G33_p_spl_010;
  wire G33_p_spl_1;
  wire G33_p_spl_10;
  wire G33_p_spl_11;
  wire G23_n_spl_;
  wire G23_n_spl_0;
  wire G23_n_spl_1;
  wire G24_p_spl_;
  wire G24_p_spl_0;
  wire G24_p_spl_1;
  wire G23_p_spl_;
  wire G23_p_spl_0;
  wire G23_p_spl_1;
  wire G24_n_spl_;
  wire G24_n_spl_0;
  wire G24_n_spl_1;
  wire G31_n_spl_;
  wire G31_n_spl_0;
  wire G31_n_spl_00;
  wire G31_n_spl_000;
  wire G31_n_spl_001;
  wire G31_n_spl_01;
  wire G31_n_spl_010;
  wire G31_n_spl_011;
  wire G31_n_spl_1;
  wire G31_n_spl_10;
  wire G31_n_spl_11;
  wire g35_n_spl_;
  wire G31_p_spl_;
  wire G31_p_spl_0;
  wire G31_p_spl_00;
  wire G31_p_spl_000;
  wire G31_p_spl_001;
  wire G31_p_spl_01;
  wire G31_p_spl_010;
  wire G31_p_spl_011;
  wire G31_p_spl_1;
  wire G31_p_spl_10;
  wire G31_p_spl_100;
  wire G31_p_spl_101;
  wire G31_p_spl_11;
  wire G31_p_spl_110;
  wire g35_p_spl_;
  wire g34_p_spl_;
  wire g36_p_spl_;
  wire g34_n_spl_;
  wire g36_n_spl_;
  wire G32_n_spl_;
  wire g38_p_spl_;
  wire g38_p_spl_0;
  wire g38_p_spl_00;
  wire g38_p_spl_01;
  wire g38_p_spl_1;
  wire g38_p_spl_10;
  wire g39_n_spl_;
  wire g39_p_spl_;
  wire G20_p_spl_;
  wire g41_n_spl_;
  wire G20_n_spl_;
  wire g41_p_spl_;
  wire G22_p_spl_;
  wire G22_n_spl_;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_00;
  wire G4_p_spl_01;
  wire G4_p_spl_1;
  wire G4_p_spl_10;
  wire G14_n_spl_;
  wire G14_n_spl_0;
  wire G14_n_spl_00;
  wire G14_n_spl_1;
  wire G4_n_spl_;
  wire G4_n_spl_0;
  wire G4_n_spl_00;
  wire G4_n_spl_01;
  wire G4_n_spl_1;
  wire G4_n_spl_10;
  wire G14_p_spl_;
  wire G14_p_spl_0;
  wire G14_p_spl_00;
  wire G14_p_spl_1;
  wire g43_p_spl_;
  wire g46_p_spl_;
  wire g43_n_spl_;
  wire g46_n_spl_;
  wire G12_p_spl_;
  wire G12_p_spl_0;
  wire G12_p_spl_00;
  wire G12_p_spl_1;
  wire G13_n_spl_;
  wire G13_n_spl_0;
  wire G13_n_spl_00;
  wire G13_n_spl_1;
  wire G12_n_spl_;
  wire G12_n_spl_0;
  wire G12_n_spl_00;
  wire G12_n_spl_1;
  wire G13_p_spl_;
  wire G13_p_spl_0;
  wire G13_p_spl_00;
  wire G13_p_spl_1;
  wire G11_p_spl_;
  wire G11_p_spl_0;
  wire G11_p_spl_00;
  wire G11_p_spl_1;
  wire g52_p_spl_;
  wire G11_n_spl_;
  wire G11_n_spl_0;
  wire G11_n_spl_00;
  wire G11_n_spl_1;
  wire g52_n_spl_;
  wire G10_n_spl_;
  wire G10_n_spl_0;
  wire G10_n_spl_00;
  wire G10_n_spl_1;
  wire G15_n_spl_;
  wire G15_n_spl_0;
  wire G15_n_spl_00;
  wire G15_n_spl_1;
  wire G10_p_spl_;
  wire G10_p_spl_0;
  wire G10_p_spl_00;
  wire G10_p_spl_1;
  wire G15_p_spl_;
  wire G15_p_spl_0;
  wire G15_p_spl_00;
  wire G15_p_spl_1;
  wire G16_p_spl_;
  wire G16_p_spl_0;
  wire G16_p_spl_00;
  wire G16_p_spl_1;
  wire g58_n_spl_;
  wire g58_n_spl_0;
  wire g58_n_spl_1;
  wire G16_n_spl_;
  wire G16_n_spl_0;
  wire G16_n_spl_00;
  wire G16_n_spl_1;
  wire g58_p_spl_;
  wire g58_p_spl_0;
  wire g58_p_spl_1;
  wire g55_n_spl_;
  wire g61_p_spl_;
  wire g61_p_spl_0;
  wire g61_p_spl_1;
  wire g55_p_spl_;
  wire g61_n_spl_;
  wire g61_n_spl_0;
  wire g61_n_spl_1;
  wire G2_p_spl_;
  wire G2_p_spl_0;
  wire G2_p_spl_00;
  wire G2_p_spl_1;
  wire G3_n_spl_;
  wire G3_n_spl_0;
  wire G3_n_spl_00;
  wire G3_n_spl_1;
  wire G2_n_spl_;
  wire G2_n_spl_0;
  wire G2_n_spl_00;
  wire G2_n_spl_1;
  wire G3_p_spl_;
  wire G3_p_spl_0;
  wire G3_p_spl_00;
  wire G3_p_spl_1;
  wire G1_p_spl_;
  wire G1_p_spl_0;
  wire G1_p_spl_00;
  wire G1_p_spl_1;
  wire g67_p_spl_;
  wire G1_n_spl_;
  wire G1_n_spl_0;
  wire G1_n_spl_00;
  wire G1_n_spl_1;
  wire g67_n_spl_;
  wire g64_n_spl_;
  wire g64_n_spl_0;
  wire g64_n_spl_00;
  wire g64_n_spl_01;
  wire g64_n_spl_1;
  wire g70_n_spl_;
  wire g70_n_spl_0;
  wire g70_n_spl_1;
  wire g64_p_spl_;
  wire g64_p_spl_0;
  wire g64_p_spl_00;
  wire g64_p_spl_01;
  wire g64_p_spl_1;
  wire g70_p_spl_;
  wire g70_p_spl_0;
  wire g70_p_spl_1;
  wire g49_n_spl_;
  wire g73_n_spl_;
  wire g49_p_spl_;
  wire g73_p_spl_;
  wire g76_n_spl_;
  wire g76_p_spl_;
  wire G25_n_spl_;
  wire G25_n_spl_0;
  wire g77_p_spl_;
  wire G25_p_spl_;
  wire G25_p_spl_0;
  wire g77_n_spl_;
  wire g42_p_spl_;
  wire g42_p_spl_0;
  wire g80_n_spl_;
  wire g80_n_spl_0;
  wire g42_n_spl_;
  wire g80_p_spl_;
  wire G18_p_spl_;
  wire G18_n_spl_;
  wire g83_n_spl_;
  wire g83_p_spl_;
  wire g86_n_spl_;
  wire g86_p_spl_;
  wire G9_p_spl_;
  wire G9_p_spl_0;
  wire G9_p_spl_00;
  wire G9_p_spl_1;
  wire G9_n_spl_;
  wire G9_n_spl_0;
  wire G9_n_spl_00;
  wire G9_n_spl_1;
  wire g92_n_spl_;
  wire g92_n_spl_0;
  wire g92_n_spl_1;
  wire g92_p_spl_;
  wire g92_p_spl_0;
  wire g92_p_spl_1;
  wire g89_p_spl_;
  wire g95_p_spl_;
  wire g95_p_spl_0;
  wire g95_p_spl_1;
  wire g89_n_spl_;
  wire g95_n_spl_;
  wire g95_n_spl_0;
  wire g95_n_spl_1;
  wire G5_n_spl_;
  wire G5_n_spl_0;
  wire G5_n_spl_00;
  wire G5_n_spl_1;
  wire G8_n_spl_;
  wire G8_n_spl_0;
  wire G8_n_spl_00;
  wire G8_n_spl_01;
  wire G8_n_spl_1;
  wire G8_n_spl_10;
  wire G5_p_spl_;
  wire G5_p_spl_0;
  wire G5_p_spl_00;
  wire G5_p_spl_1;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire G8_p_spl_00;
  wire G8_p_spl_01;
  wire G8_p_spl_1;
  wire G8_p_spl_10;
  wire g101_p_spl_;
  wire g101_n_spl_;
  wire g98_n_spl_;
  wire g104_p_spl_;
  wire g98_p_spl_;
  wire g104_n_spl_;
  wire g107_n_spl_;
  wire G27_n_spl_;
  wire G27_n_spl_0;
  wire g108_p_spl_;
  wire G27_p_spl_;
  wire g108_n_spl_;
  wire G6_n_spl_;
  wire G6_n_spl_0;
  wire G6_n_spl_00;
  wire G6_n_spl_1;
  wire G6_p_spl_;
  wire G6_p_spl_0;
  wire G6_p_spl_00;
  wire G6_p_spl_1;
  wire g112_p_spl_;
  wire g112_n_spl_;
  wire g115_n_spl_;
  wire g118_n_spl_;
  wire g115_p_spl_;
  wire g118_p_spl_;
  wire G19_p_spl_;
  wire G19_n_spl_;
  wire g121_n_spl_;
  wire g123_n_spl_;
  wire g121_p_spl_;
  wire g123_p_spl_;
  wire g126_n_spl_;
  wire G28_n_spl_;
  wire G28_n_spl_0;
  wire g127_p_spl_;
  wire G28_p_spl_;
  wire g127_n_spl_;
  wire G7_n_spl_;
  wire G7_n_spl_0;
  wire G7_n_spl_00;
  wire G7_n_spl_1;
  wire G7_p_spl_;
  wire G7_p_spl_0;
  wire G7_p_spl_00;
  wire G7_p_spl_1;
  wire g133_p_spl_;
  wire g133_n_spl_;
  wire g136_n_spl_;
  wire g136_p_spl_;
  wire g141_p_spl_;
  wire g141_n_spl_;
  wire g139_n_spl_;
  wire g144_n_spl_;
  wire g139_p_spl_;
  wire g144_p_spl_;
  wire g147_n_spl_;
  wire g148_p_spl_;
  wire g149_n_spl_;
  wire g149_n_spl_0;
  wire g148_n_spl_;
  wire g149_p_spl_;
  wire G17_p_spl_;
  wire G17_n_spl_;
  wire g156_p_spl_;
  wire g156_n_spl_;
  wire g162_p_spl_;
  wire g162_n_spl_;
  wire g165_n_spl_;
  wire g165_n_spl_0;
  wire g165_n_spl_1;
  wire g165_p_spl_;
  wire g165_p_spl_0;
  wire g165_p_spl_1;
  wire g159_p_spl_;
  wire g168_p_spl_;
  wire g159_n_spl_;
  wire g168_n_spl_;
  wire g171_n_spl_;
  wire g171_p_spl_;
  wire G26_p_spl_;
  wire G26_p_spl_0;
  wire g172_n_spl_;
  wire G26_n_spl_;
  wire G26_n_spl_0;
  wire g172_p_spl_;
  wire g179_n_spl_;
  wire g179_p_spl_;
  wire G21_p_spl_;
  wire G21_n_spl_;
  wire g181_p_spl_;
  wire g184_p_spl_;
  wire g181_n_spl_;
  wire g184_n_spl_;
  wire g190_p_spl_;
  wire g193_n_spl_;
  wire g190_n_spl_;
  wire g193_p_spl_;
  wire g187_p_spl_;
  wire g196_n_spl_;
  wire g196_n_spl_0;
  wire g187_n_spl_;
  wire g196_p_spl_;
  wire g196_p_spl_0;
  wire g199_p_spl_;
  wire g199_n_spl_;
  wire g200_p_spl_;
  wire g201_n_spl_;
  wire g201_n_spl_0;
  wire g200_n_spl_;
  wire g201_p_spl_;
  wire g201_p_spl_0;
  wire g180_p_spl_;
  wire g180_p_spl_0;
  wire g204_n_spl_;
  wire g204_n_spl_0;
  wire g180_n_spl_;
  wire g204_p_spl_;
  wire g178_p_spl_;
  wire g178_n_spl_;
  wire g178_n_spl_0;
  wire g81_n_spl_;
  wire g206_p_spl_;
  wire g81_p_spl_;
  wire g206_n_spl_;
  wire g40_n_spl_;
  wire g207_p_spl_;
  wire g40_p_spl_;
  wire g207_n_spl_;
  wire g208_n_spl_;
  wire g208_n_spl_0;
  wire g208_n_spl_00;
  wire g208_n_spl_01;
  wire g208_n_spl_1;
  wire g208_n_spl_10;
  wire g208_p_spl_;
  wire g208_p_spl_0;
  wire g208_p_spl_00;
  wire g208_p_spl_01;
  wire g208_p_spl_1;
  wire g208_p_spl_10;
  wire G30_n_spl_;
  wire G30_p_spl_;
  wire g221_p_spl_;
  wire g221_n_spl_;
  wire g223_n_spl_;
  wire g223_n_spl_0;
  wire g223_p_spl_;
  wire g223_p_spl_0;
  wire g224_n_spl_;
  wire g224_n_spl_0;
  wire g224_n_spl_00;
  wire g224_n_spl_01;
  wire g224_n_spl_1;
  wire g224_p_spl_;
  wire g224_p_spl_0;
  wire g224_p_spl_00;
  wire g224_p_spl_01;
  wire g224_p_spl_1;
  wire g235_p_spl_;
  wire g235_n_spl_;
  wire g236_n_spl_;
  wire g236_n_spl_0;
  wire g236_n_spl_1;
  wire g236_p_spl_;
  wire g236_p_spl_0;
  wire g236_p_spl_1;
  wire g256_n_spl_;
  wire g256_n_spl_0;
  wire g256_n_spl_1;
  wire g256_p_spl_;
  wire g256_p_spl_0;
  wire g256_p_spl_1;
  wire g269_p_spl_;
  wire g269_p_spl_0;
  wire g269_p_spl_00;
  wire g269_p_spl_01;
  wire g269_p_spl_1;
  wire g269_p_spl_10;
  wire g269_n_spl_;
  wire g269_n_spl_0;
  wire g303_n_spl_;
  wire g303_p_spl_;
  wire g315_n_spl_;
  wire g315_p_spl_;

  LA
  g_g34_p
  (
    .dout(g34_p),
    .din1(G29_n_spl_),
    .din2(G33_n_spl_000)
  );


  FA
  g_g34_n
  (
    .dout(g34_n),
    .din1(G29_p_spl_),
    .din2(G33_p_spl_000)
  );


  LA
  g_g35_p
  (
    .dout(g35_p),
    .din1(G23_n_spl_0),
    .din2(G24_p_spl_0)
  );


  FA
  g_g35_n
  (
    .dout(g35_n),
    .din1(G23_p_spl_0),
    .din2(G24_n_spl_0)
  );


  LA
  g_g36_p
  (
    .dout(g36_p),
    .din1(G31_n_spl_000),
    .din2(g35_n_spl_)
  );


  FA
  g_g36_n
  (
    .dout(g36_n),
    .din1(G31_p_spl_000),
    .din2(g35_p_spl_)
  );


  LA
  g_g37_p
  (
    .dout(g37_p),
    .din1(g34_p_spl_),
    .din2(g36_p_spl_)
  );


  FA
  g_g37_n
  (
    .dout(g37_n),
    .din1(g34_n_spl_),
    .din2(g36_n_spl_)
  );


  LA
  g_g38_p
  (
    .dout(g38_p),
    .din1(G32_n_spl_),
    .din2(G33_n_spl_000)
  );


  FA
  g_g38_n
  (
    .dout(g38_n),
    .din1(G32_p),
    .din2(G33_p_spl_000)
  );


  LA
  g_g39_p
  (
    .dout(g39_p),
    .din1(g35_n_spl_),
    .din2(g38_p_spl_00)
  );


  FA
  g_g39_n
  (
    .dout(g39_n),
    .din1(g35_p_spl_),
    .din2(g38_n)
  );


  LA
  g_g40_p
  (
    .dout(g40_p),
    .din1(g37_n),
    .din2(g39_n_spl_)
  );


  FA
  g_g40_n
  (
    .dout(g40_n),
    .din1(g37_p),
    .din2(g39_p_spl_)
  );


  LA
  g_g41_p
  (
    .dout(g41_p),
    .din1(G23_n_spl_0),
    .din2(G31_n_spl_000)
  );


  FA
  g_g41_n
  (
    .dout(g41_n),
    .din1(G23_p_spl_0),
    .din2(G31_p_spl_000)
  );


  LA
  g_g42_p
  (
    .dout(g42_p),
    .din1(G20_p_spl_),
    .din2(g41_n_spl_)
  );


  FA
  g_g42_n
  (
    .dout(g42_n),
    .din1(G20_n_spl_),
    .din2(g41_p_spl_)
  );


  LA
  g_g43_p
  (
    .dout(g43_p),
    .din1(G22_p_spl_),
    .din2(G33_n_spl_001)
  );


  FA
  g_g43_n
  (
    .dout(g43_n),
    .din1(G22_n_spl_),
    .din2(G33_p_spl_001)
  );


  LA
  g_g44_p
  (
    .dout(g44_p),
    .din1(G4_p_spl_00),
    .din2(G14_n_spl_00)
  );


  FA
  g_g44_n
  (
    .dout(g44_n),
    .din1(G4_n_spl_00),
    .din2(G14_p_spl_00)
  );


  LA
  g_g45_p
  (
    .dout(g45_p),
    .din1(G4_n_spl_00),
    .din2(G14_p_spl_00)
  );


  FA
  g_g45_n
  (
    .dout(g45_n),
    .din1(G4_p_spl_00),
    .din2(G14_n_spl_00)
  );


  LA
  g_g46_p
  (
    .dout(g46_p),
    .din1(g44_n),
    .din2(g45_n)
  );


  FA
  g_g46_n
  (
    .dout(g46_n),
    .din1(g44_p),
    .din2(g45_p)
  );


  LA
  g_g47_p
  (
    .dout(g47_p),
    .din1(g43_p_spl_),
    .din2(g46_p_spl_)
  );


  FA
  g_g47_n
  (
    .dout(g47_n),
    .din1(g43_n_spl_),
    .din2(g46_n_spl_)
  );


  LA
  g_g48_p
  (
    .dout(g48_p),
    .din1(g43_n_spl_),
    .din2(g46_n_spl_)
  );


  FA
  g_g48_n
  (
    .dout(g48_n),
    .din1(g43_p_spl_),
    .din2(g46_p_spl_)
  );


  LA
  g_g49_p
  (
    .dout(g49_p),
    .din1(g47_n),
    .din2(g48_n)
  );


  FA
  g_g49_n
  (
    .dout(g49_n),
    .din1(g47_p),
    .din2(g48_p)
  );


  LA
  g_g50_p
  (
    .dout(g50_p),
    .din1(G12_p_spl_00),
    .din2(G13_n_spl_00)
  );


  FA
  g_g50_n
  (
    .dout(g50_n),
    .din1(G12_n_spl_00),
    .din2(G13_p_spl_00)
  );


  LA
  g_g51_p
  (
    .dout(g51_p),
    .din1(G12_n_spl_00),
    .din2(G13_p_spl_00)
  );


  FA
  g_g51_n
  (
    .dout(g51_n),
    .din1(G12_p_spl_00),
    .din2(G13_n_spl_00)
  );


  LA
  g_g52_p
  (
    .dout(g52_p),
    .din1(g50_n),
    .din2(g51_n)
  );


  FA
  g_g52_n
  (
    .dout(g52_n),
    .din1(g50_p),
    .din2(g51_p)
  );


  LA
  g_g53_p
  (
    .dout(g53_p),
    .din1(G11_p_spl_00),
    .din2(g52_p_spl_)
  );


  FA
  g_g53_n
  (
    .dout(g53_n),
    .din1(G11_n_spl_00),
    .din2(g52_n_spl_)
  );


  LA
  g_g54_p
  (
    .dout(g54_p),
    .din1(G11_n_spl_00),
    .din2(g52_n_spl_)
  );


  FA
  g_g54_n
  (
    .dout(g54_n),
    .din1(G11_p_spl_00),
    .din2(g52_p_spl_)
  );


  LA
  g_g55_p
  (
    .dout(g55_p),
    .din1(g53_n),
    .din2(g54_n)
  );


  FA
  g_g55_n
  (
    .dout(g55_n),
    .din1(g53_p),
    .din2(g54_p)
  );


  LA
  g_g56_p
  (
    .dout(g56_p),
    .din1(G10_n_spl_00),
    .din2(G15_n_spl_00)
  );


  FA
  g_g56_n
  (
    .dout(g56_n),
    .din1(G10_p_spl_00),
    .din2(G15_p_spl_00)
  );


  LA
  g_g57_p
  (
    .dout(g57_p),
    .din1(G10_p_spl_00),
    .din2(G15_p_spl_00)
  );


  FA
  g_g57_n
  (
    .dout(g57_n),
    .din1(G10_n_spl_00),
    .din2(G15_n_spl_00)
  );


  LA
  g_g58_p
  (
    .dout(g58_p),
    .din1(g56_n),
    .din2(g57_n)
  );


  FA
  g_g58_n
  (
    .dout(g58_n),
    .din1(g56_p),
    .din2(g57_p)
  );


  LA
  g_g59_p
  (
    .dout(g59_p),
    .din1(G16_p_spl_00),
    .din2(g58_n_spl_0)
  );


  FA
  g_g59_n
  (
    .dout(g59_n),
    .din1(G16_n_spl_00),
    .din2(g58_p_spl_0)
  );


  LA
  g_g60_p
  (
    .dout(g60_p),
    .din1(G16_n_spl_00),
    .din2(g58_p_spl_0)
  );


  FA
  g_g60_n
  (
    .dout(g60_n),
    .din1(G16_p_spl_00),
    .din2(g58_n_spl_0)
  );


  LA
  g_g61_p
  (
    .dout(g61_p),
    .din1(g59_n),
    .din2(g60_n)
  );


  FA
  g_g61_n
  (
    .dout(g61_n),
    .din1(g59_p),
    .din2(g60_p)
  );


  LA
  g_g62_p
  (
    .dout(g62_p),
    .din1(g55_n_spl_),
    .din2(g61_p_spl_0)
  );


  FA
  g_g62_n
  (
    .dout(g62_n),
    .din1(g55_p_spl_),
    .din2(g61_n_spl_0)
  );


  LA
  g_g63_p
  (
    .dout(g63_p),
    .din1(g55_p_spl_),
    .din2(g61_n_spl_0)
  );


  FA
  g_g63_n
  (
    .dout(g63_n),
    .din1(g55_n_spl_),
    .din2(g61_p_spl_0)
  );


  LA
  g_g64_p
  (
    .dout(g64_p),
    .din1(g62_n),
    .din2(g63_n)
  );


  FA
  g_g64_n
  (
    .dout(g64_n),
    .din1(g62_p),
    .din2(g63_p)
  );


  LA
  g_g65_p
  (
    .dout(g65_p),
    .din1(G2_p_spl_00),
    .din2(G3_n_spl_00)
  );


  FA
  g_g65_n
  (
    .dout(g65_n),
    .din1(G2_n_spl_00),
    .din2(G3_p_spl_00)
  );


  LA
  g_g66_p
  (
    .dout(g66_p),
    .din1(G2_n_spl_00),
    .din2(G3_p_spl_00)
  );


  FA
  g_g66_n
  (
    .dout(g66_n),
    .din1(G2_p_spl_00),
    .din2(G3_n_spl_00)
  );


  LA
  g_g67_p
  (
    .dout(g67_p),
    .din1(g65_n),
    .din2(g66_n)
  );


  FA
  g_g67_n
  (
    .dout(g67_n),
    .din1(g65_p),
    .din2(g66_p)
  );


  LA
  g_g68_p
  (
    .dout(g68_p),
    .din1(G1_p_spl_00),
    .din2(g67_p_spl_)
  );


  FA
  g_g68_n
  (
    .dout(g68_n),
    .din1(G1_n_spl_00),
    .din2(g67_n_spl_)
  );


  LA
  g_g69_p
  (
    .dout(g69_p),
    .din1(G1_n_spl_00),
    .din2(g67_n_spl_)
  );


  FA
  g_g69_n
  (
    .dout(g69_n),
    .din1(G1_p_spl_00),
    .din2(g67_p_spl_)
  );


  LA
  g_g70_p
  (
    .dout(g70_p),
    .din1(g68_n),
    .din2(g69_n)
  );


  FA
  g_g70_n
  (
    .dout(g70_n),
    .din1(g68_p),
    .din2(g69_p)
  );


  LA
  g_g71_p
  (
    .dout(g71_p),
    .din1(g64_n_spl_00),
    .din2(g70_n_spl_0)
  );


  FA
  g_g71_n
  (
    .dout(g71_n),
    .din1(g64_p_spl_00),
    .din2(g70_p_spl_0)
  );


  LA
  g_g72_p
  (
    .dout(g72_p),
    .din1(g64_p_spl_00),
    .din2(g70_p_spl_0)
  );


  FA
  g_g72_n
  (
    .dout(g72_n),
    .din1(g64_n_spl_00),
    .din2(g70_n_spl_0)
  );


  LA
  g_g73_p
  (
    .dout(g73_p),
    .din1(g71_n),
    .din2(g72_n)
  );


  FA
  g_g73_n
  (
    .dout(g73_n),
    .din1(g71_p),
    .din2(g72_p)
  );


  LA
  g_g74_p
  (
    .dout(g74_p),
    .din1(g49_n_spl_),
    .din2(g73_n_spl_)
  );


  FA
  g_g74_n
  (
    .dout(g74_n),
    .din1(g49_p_spl_),
    .din2(g73_p_spl_)
  );


  LA
  g_g75_p
  (
    .dout(g75_p),
    .din1(g49_p_spl_),
    .din2(g73_p_spl_)
  );


  FA
  g_g75_n
  (
    .dout(g75_n),
    .din1(g49_n_spl_),
    .din2(g73_n_spl_)
  );


  LA
  g_g76_p
  (
    .dout(g76_p),
    .din1(g74_n),
    .din2(g75_n)
  );


  FA
  g_g76_n
  (
    .dout(g76_n),
    .din1(g74_p),
    .din2(g75_p)
  );


  LA
  g_g77_p
  (
    .dout(g77_p),
    .din1(G31_n_spl_001),
    .din2(g76_n_spl_)
  );


  FA
  g_g77_n
  (
    .dout(g77_n),
    .din1(G31_p_spl_001),
    .din2(g76_p_spl_)
  );


  LA
  g_g78_p
  (
    .dout(g78_p),
    .din1(G25_n_spl_0),
    .din2(g77_p_spl_)
  );


  FA
  g_g78_n
  (
    .dout(g78_n),
    .din1(G25_p_spl_0),
    .din2(g77_n_spl_)
  );


  LA
  g_g79_p
  (
    .dout(g79_p),
    .din1(G25_p_spl_0),
    .din2(g77_n_spl_)
  );


  FA
  g_g79_n
  (
    .dout(g79_n),
    .din1(G25_n_spl_0),
    .din2(g77_p_spl_)
  );


  LA
  g_g80_p
  (
    .dout(g80_p),
    .din1(g78_n),
    .din2(g79_n)
  );


  FA
  g_g80_n
  (
    .dout(g80_n),
    .din1(g78_p),
    .din2(g79_p)
  );


  LA
  g_g81_p
  (
    .dout(g81_p),
    .din1(g42_p_spl_0),
    .din2(g80_n_spl_0)
  );


  FA
  g_g81_n
  (
    .dout(g81_n),
    .din1(g42_n_spl_),
    .din2(g80_p_spl_)
  );


  LA
  g_g82_p
  (
    .dout(g82_p),
    .din1(G18_p_spl_),
    .din2(G33_n_spl_001)
  );


  FA
  g_g82_n
  (
    .dout(g82_n),
    .din1(G18_n_spl_),
    .din2(G33_p_spl_001)
  );


  LA
  g_g83_p
  (
    .dout(g83_p),
    .din1(G24_n_spl_0),
    .din2(g82_p)
  );


  FA
  g_g83_n
  (
    .dout(g83_n),
    .din1(G24_p_spl_0),
    .din2(g82_n)
  );


  LA
  g_g84_p
  (
    .dout(g84_p),
    .din1(G15_p_spl_0),
    .din2(g83_n_spl_)
  );


  FA
  g_g84_n
  (
    .dout(g84_n),
    .din1(G15_n_spl_0),
    .din2(g83_p_spl_)
  );


  LA
  g_g85_p
  (
    .dout(g85_p),
    .din1(G15_n_spl_1),
    .din2(g83_p_spl_)
  );


  FA
  g_g85_n
  (
    .dout(g85_n),
    .din1(G15_p_spl_1),
    .din2(g83_n_spl_)
  );


  LA
  g_g86_p
  (
    .dout(g86_p),
    .din1(g84_n),
    .din2(g85_n)
  );


  FA
  g_g86_n
  (
    .dout(g86_n),
    .din1(g84_p),
    .din2(g85_p)
  );


  LA
  g_g87_p
  (
    .dout(g87_p),
    .din1(G11_n_spl_0),
    .din2(g86_n_spl_)
  );


  FA
  g_g87_n
  (
    .dout(g87_n),
    .din1(G11_p_spl_0),
    .din2(g86_p_spl_)
  );


  LA
  g_g88_p
  (
    .dout(g88_p),
    .din1(G11_p_spl_1),
    .din2(g86_p_spl_)
  );


  FA
  g_g88_n
  (
    .dout(g88_n),
    .din1(G11_n_spl_1),
    .din2(g86_n_spl_)
  );


  LA
  g_g89_p
  (
    .dout(g89_p),
    .din1(g87_n),
    .din2(g88_n)
  );


  FA
  g_g89_n
  (
    .dout(g89_n),
    .din1(g87_p),
    .din2(g88_p)
  );


  LA
  g_g90_p
  (
    .dout(g90_p),
    .din1(G9_p_spl_00),
    .din2(G14_n_spl_0)
  );


  FA
  g_g90_n
  (
    .dout(g90_n),
    .din1(G9_n_spl_00),
    .din2(G14_p_spl_0)
  );


  LA
  g_g91_p
  (
    .dout(g91_p),
    .din1(G9_n_spl_00),
    .din2(G14_p_spl_1)
  );


  FA
  g_g91_n
  (
    .dout(g91_n),
    .din1(G9_p_spl_00),
    .din2(G14_n_spl_1)
  );


  LA
  g_g92_p
  (
    .dout(g92_p),
    .din1(g90_n),
    .din2(g91_n)
  );


  FA
  g_g92_n
  (
    .dout(g92_n),
    .din1(g90_p),
    .din2(g91_p)
  );


  LA
  g_g93_p
  (
    .dout(g93_p),
    .din1(G16_p_spl_0),
    .din2(g92_n_spl_0)
  );


  FA
  g_g93_n
  (
    .dout(g93_n),
    .din1(G16_n_spl_0),
    .din2(g92_p_spl_0)
  );


  LA
  g_g94_p
  (
    .dout(g94_p),
    .din1(G16_n_spl_1),
    .din2(g92_p_spl_0)
  );


  FA
  g_g94_n
  (
    .dout(g94_n),
    .din1(G16_p_spl_1),
    .din2(g92_n_spl_0)
  );


  LA
  g_g95_p
  (
    .dout(g95_p),
    .din1(g93_n),
    .din2(g94_n)
  );


  FA
  g_g95_n
  (
    .dout(g95_n),
    .din1(g93_p),
    .din2(g94_p)
  );


  LA
  g_g96_p
  (
    .dout(g96_p),
    .din1(g89_p_spl_),
    .din2(g95_p_spl_0)
  );


  FA
  g_g96_n
  (
    .dout(g96_n),
    .din1(g89_n_spl_),
    .din2(g95_n_spl_0)
  );


  LA
  g_g97_p
  (
    .dout(g97_p),
    .din1(g89_n_spl_),
    .din2(g95_n_spl_0)
  );


  FA
  g_g97_n
  (
    .dout(g97_n),
    .din1(g89_p_spl_),
    .din2(g95_p_spl_0)
  );


  LA
  g_g98_p
  (
    .dout(g98_p),
    .din1(g96_n),
    .din2(g97_n)
  );


  FA
  g_g98_n
  (
    .dout(g98_n),
    .din1(g96_p),
    .din2(g97_p)
  );


  LA
  g_g99_p
  (
    .dout(g99_p),
    .din1(G5_n_spl_00),
    .din2(G8_n_spl_00)
  );


  FA
  g_g99_n
  (
    .dout(g99_n),
    .din1(G5_p_spl_00),
    .din2(G8_p_spl_00)
  );


  LA
  g_g100_p
  (
    .dout(g100_p),
    .din1(G5_p_spl_00),
    .din2(G8_p_spl_00)
  );


  FA
  g_g100_n
  (
    .dout(g100_n),
    .din1(G5_n_spl_00),
    .din2(G8_n_spl_00)
  );


  LA
  g_g101_p
  (
    .dout(g101_p),
    .din1(g99_n),
    .din2(g100_n)
  );


  FA
  g_g101_n
  (
    .dout(g101_n),
    .din1(g99_p),
    .din2(g100_p)
  );


  LA
  g_g102_p
  (
    .dout(g102_p),
    .din1(G2_n_spl_0),
    .din2(g101_p_spl_)
  );


  FA
  g_g102_n
  (
    .dout(g102_n),
    .din1(G2_p_spl_0),
    .din2(g101_n_spl_)
  );


  LA
  g_g103_p
  (
    .dout(g103_p),
    .din1(G2_p_spl_1),
    .din2(g101_n_spl_)
  );


  FA
  g_g103_n
  (
    .dout(g103_n),
    .din1(G2_n_spl_1),
    .din2(g101_p_spl_)
  );


  LA
  g_g104_p
  (
    .dout(g104_p),
    .din1(g102_n),
    .din2(g103_n)
  );


  FA
  g_g104_n
  (
    .dout(g104_n),
    .din1(g102_p),
    .din2(g103_p)
  );


  LA
  g_g105_p
  (
    .dout(g105_p),
    .din1(g98_n_spl_),
    .din2(g104_p_spl_)
  );


  FA
  g_g105_n
  (
    .dout(g105_n),
    .din1(g98_p_spl_),
    .din2(g104_n_spl_)
  );


  LA
  g_g106_p
  (
    .dout(g106_p),
    .din1(g98_p_spl_),
    .din2(g104_n_spl_)
  );


  FA
  g_g106_n
  (
    .dout(g106_n),
    .din1(g98_n_spl_),
    .din2(g104_p_spl_)
  );


  LA
  g_g107_p
  (
    .dout(g107_p),
    .din1(g105_n),
    .din2(g106_n)
  );


  FA
  g_g107_n
  (
    .dout(g107_n),
    .din1(g105_p),
    .din2(g106_p)
  );


  LA
  g_g108_p
  (
    .dout(g108_p),
    .din1(G31_n_spl_001),
    .din2(g107_n_spl_)
  );


  FA
  g_g108_n
  (
    .dout(g108_n),
    .din1(G31_p_spl_001),
    .din2(g107_p)
  );


  LA
  g_g109_p
  (
    .dout(g109_p),
    .din1(G27_n_spl_0),
    .din2(g108_p_spl_)
  );


  FA
  g_g109_n
  (
    .dout(g109_n),
    .din1(G27_p_spl_),
    .din2(g108_n_spl_)
  );


  LA
  g_g110_p
  (
    .dout(g110_p),
    .din1(G6_n_spl_00),
    .din2(G8_n_spl_01)
  );


  FA
  g_g110_n
  (
    .dout(g110_n),
    .din1(G6_p_spl_00),
    .din2(G8_p_spl_01)
  );


  LA
  g_g111_p
  (
    .dout(g111_p),
    .din1(G6_p_spl_00),
    .din2(G8_p_spl_01)
  );


  FA
  g_g111_n
  (
    .dout(g111_n),
    .din1(G6_n_spl_00),
    .din2(G8_n_spl_01)
  );


  LA
  g_g112_p
  (
    .dout(g112_p),
    .din1(g110_n),
    .din2(g111_n)
  );


  FA
  g_g112_n
  (
    .dout(g112_n),
    .din1(g110_p),
    .din2(g111_p)
  );


  LA
  g_g113_p
  (
    .dout(g113_p),
    .din1(G3_n_spl_0),
    .din2(g112_p_spl_)
  );


  FA
  g_g113_n
  (
    .dout(g113_n),
    .din1(G3_p_spl_0),
    .din2(g112_n_spl_)
  );


  LA
  g_g114_p
  (
    .dout(g114_p),
    .din1(G3_p_spl_1),
    .din2(g112_n_spl_)
  );


  FA
  g_g114_n
  (
    .dout(g114_n),
    .din1(G3_n_spl_1),
    .din2(g112_p_spl_)
  );


  LA
  g_g115_p
  (
    .dout(g115_p),
    .din1(g113_n),
    .din2(g114_n)
  );


  FA
  g_g115_n
  (
    .dout(g115_n),
    .din1(g113_p),
    .din2(g114_p)
  );


  LA
  g_g116_p
  (
    .dout(g116_p),
    .din1(G12_n_spl_0),
    .din2(g58_n_spl_1)
  );


  FA
  g_g116_n
  (
    .dout(g116_n),
    .din1(G12_p_spl_0),
    .din2(g58_p_spl_1)
  );


  LA
  g_g117_p
  (
    .dout(g117_p),
    .din1(G12_p_spl_1),
    .din2(g58_p_spl_1)
  );


  FA
  g_g117_n
  (
    .dout(g117_n),
    .din1(G12_n_spl_1),
    .din2(g58_n_spl_1)
  );


  LA
  g_g118_p
  (
    .dout(g118_p),
    .din1(g116_n),
    .din2(g117_n)
  );


  FA
  g_g118_n
  (
    .dout(g118_n),
    .din1(g116_p),
    .din2(g117_p)
  );


  LA
  g_g119_p
  (
    .dout(g119_p),
    .din1(g115_n_spl_),
    .din2(g118_n_spl_)
  );


  FA
  g_g119_n
  (
    .dout(g119_n),
    .din1(g115_p_spl_),
    .din2(g118_p_spl_)
  );


  LA
  g_g120_p
  (
    .dout(g120_p),
    .din1(g115_p_spl_),
    .din2(g118_p_spl_)
  );


  FA
  g_g120_n
  (
    .dout(g120_n),
    .din1(g115_n_spl_),
    .din2(g118_n_spl_)
  );


  LA
  g_g121_p
  (
    .dout(g121_p),
    .din1(g119_n),
    .din2(g120_n)
  );


  FA
  g_g121_n
  (
    .dout(g121_n),
    .din1(g119_p),
    .din2(g120_p)
  );


  LA
  g_g122_p
  (
    .dout(g122_p),
    .din1(G19_p_spl_),
    .din2(G33_n_spl_010)
  );


  FA
  g_g122_n
  (
    .dout(g122_n),
    .din1(G19_n_spl_),
    .din2(G33_p_spl_010)
  );


  LA
  g_g123_p
  (
    .dout(g123_p),
    .din1(G23_n_spl_1),
    .din2(g122_p)
  );


  FA
  g_g123_n
  (
    .dout(g123_n),
    .din1(G23_p_spl_1),
    .din2(g122_n)
  );


  LA
  g_g124_p
  (
    .dout(g124_p),
    .din1(g121_n_spl_),
    .din2(g123_n_spl_)
  );


  FA
  g_g124_n
  (
    .dout(g124_n),
    .din1(g121_p_spl_),
    .din2(g123_p_spl_)
  );


  LA
  g_g125_p
  (
    .dout(g125_p),
    .din1(g121_p_spl_),
    .din2(g123_p_spl_)
  );


  FA
  g_g125_n
  (
    .dout(g125_n),
    .din1(g121_n_spl_),
    .din2(g123_n_spl_)
  );


  LA
  g_g126_p
  (
    .dout(g126_p),
    .din1(g124_n),
    .din2(g125_n)
  );


  FA
  g_g126_n
  (
    .dout(g126_n),
    .din1(g124_p),
    .din2(g125_p)
  );


  LA
  g_g127_p
  (
    .dout(g127_p),
    .din1(G31_n_spl_010),
    .din2(g126_n_spl_)
  );


  FA
  g_g127_n
  (
    .dout(g127_n),
    .din1(G31_p_spl_010),
    .din2(g126_p)
  );


  LA
  g_g128_p
  (
    .dout(g128_p),
    .din1(G28_n_spl_0),
    .din2(g127_p_spl_)
  );


  FA
  g_g128_n
  (
    .dout(g128_n),
    .din1(G28_p_spl_),
    .din2(g127_n_spl_)
  );


  LA
  g_g129_p
  (
    .dout(g129_p),
    .din1(G28_p_spl_),
    .din2(g127_n_spl_)
  );


  FA
  g_g129_n
  (
    .dout(g129_n),
    .din1(G28_n_spl_0),
    .din2(g127_p_spl_)
  );


  LA
  g_g130_p
  (
    .dout(g130_p),
    .din1(g128_n),
    .din2(g129_n)
  );


  FA
  g_g130_n
  (
    .dout(g130_n),
    .din1(g128_p),
    .din2(g129_p)
  );


  LA
  g_g131_p
  (
    .dout(g131_p),
    .din1(G7_n_spl_00),
    .din2(G10_n_spl_0)
  );


  FA
  g_g131_n
  (
    .dout(g131_n),
    .din1(G7_p_spl_00),
    .din2(G10_p_spl_0)
  );


  LA
  g_g132_p
  (
    .dout(g132_p),
    .din1(G7_p_spl_00),
    .din2(G10_p_spl_1)
  );


  FA
  g_g132_n
  (
    .dout(g132_n),
    .din1(G7_n_spl_00),
    .din2(G10_n_spl_1)
  );


  LA
  g_g133_p
  (
    .dout(g133_p),
    .din1(g131_n),
    .din2(g132_n)
  );


  FA
  g_g133_n
  (
    .dout(g133_n),
    .din1(g131_p),
    .din2(g132_p)
  );


  LA
  g_g134_p
  (
    .dout(g134_p),
    .din1(G4_n_spl_01),
    .din2(g133_p_spl_)
  );


  FA
  g_g134_n
  (
    .dout(g134_n),
    .din1(G4_p_spl_01),
    .din2(g133_n_spl_)
  );


  LA
  g_g135_p
  (
    .dout(g135_p),
    .din1(G4_p_spl_01),
    .din2(g133_n_spl_)
  );


  FA
  g_g135_n
  (
    .dout(g135_n),
    .din1(G4_n_spl_01),
    .din2(g133_p_spl_)
  );


  LA
  g_g136_p
  (
    .dout(g136_p),
    .din1(g134_n),
    .din2(g135_n)
  );


  FA
  g_g136_n
  (
    .dout(g136_n),
    .din1(g134_p),
    .din2(g135_p)
  );


  LA
  g_g137_p
  (
    .dout(g137_p),
    .din1(g95_n_spl_1),
    .din2(g136_n_spl_)
  );


  FA
  g_g137_n
  (
    .dout(g137_n),
    .din1(g95_p_spl_1),
    .din2(g136_p_spl_)
  );


  LA
  g_g138_p
  (
    .dout(g138_p),
    .din1(g95_p_spl_1),
    .din2(g136_p_spl_)
  );


  FA
  g_g138_n
  (
    .dout(g138_n),
    .din1(g95_n_spl_1),
    .din2(g136_n_spl_)
  );


  LA
  g_g139_p
  (
    .dout(g139_p),
    .din1(g137_n),
    .din2(g138_n)
  );


  FA
  g_g139_n
  (
    .dout(g139_n),
    .din1(g137_p),
    .din2(g138_p)
  );


  LA
  g_g140_p
  (
    .dout(g140_p),
    .din1(G20_p_spl_),
    .din2(G33_n_spl_010)
  );


  FA
  g_g140_n
  (
    .dout(g140_n),
    .din1(G20_n_spl_),
    .din2(G33_p_spl_010)
  );


  LA
  g_g141_p
  (
    .dout(g141_p),
    .din1(G23_n_spl_1),
    .din2(g140_p)
  );


  FA
  g_g141_n
  (
    .dout(g141_n),
    .din1(G23_p_spl_1),
    .din2(g140_n)
  );


  LA
  g_g142_p
  (
    .dout(g142_p),
    .din1(G13_n_spl_0),
    .din2(g141_p_spl_)
  );


  FA
  g_g142_n
  (
    .dout(g142_n),
    .din1(G13_p_spl_0),
    .din2(g141_n_spl_)
  );


  LA
  g_g143_p
  (
    .dout(g143_p),
    .din1(G13_p_spl_1),
    .din2(g141_n_spl_)
  );


  FA
  g_g143_n
  (
    .dout(g143_n),
    .din1(G13_n_spl_1),
    .din2(g141_p_spl_)
  );


  LA
  g_g144_p
  (
    .dout(g144_p),
    .din1(g142_n),
    .din2(g143_n)
  );


  FA
  g_g144_n
  (
    .dout(g144_n),
    .din1(g142_p),
    .din2(g143_p)
  );


  LA
  g_g145_p
  (
    .dout(g145_p),
    .din1(g139_n_spl_),
    .din2(g144_n_spl_)
  );


  FA
  g_g145_n
  (
    .dout(g145_n),
    .din1(g139_p_spl_),
    .din2(g144_p_spl_)
  );


  LA
  g_g146_p
  (
    .dout(g146_p),
    .din1(g139_p_spl_),
    .din2(g144_p_spl_)
  );


  FA
  g_g146_n
  (
    .dout(g146_n),
    .din1(g139_n_spl_),
    .din2(g144_n_spl_)
  );


  LA
  g_g147_p
  (
    .dout(g147_p),
    .din1(g145_n),
    .din2(g146_n)
  );


  FA
  g_g147_n
  (
    .dout(g147_n),
    .din1(g145_p),
    .din2(g146_p)
  );


  LA
  g_g148_p
  (
    .dout(g148_p),
    .din1(G31_n_spl_010),
    .din2(g147_n_spl_)
  );


  FA
  g_g148_n
  (
    .dout(g148_n),
    .din1(G31_p_spl_010),
    .din2(g147_p)
  );


  LA
  g_g149_p
  (
    .dout(g149_p),
    .din1(G19_p_spl_),
    .din2(g41_n_spl_)
  );


  FA
  g_g149_n
  (
    .dout(g149_n),
    .din1(G19_n_spl_),
    .din2(g41_p_spl_)
  );


  LA
  g_g150_p
  (
    .dout(g150_p),
    .din1(g148_p_spl_),
    .din2(g149_n_spl_0)
  );


  FA
  g_g150_n
  (
    .dout(g150_n),
    .din1(g148_n_spl_),
    .din2(g149_p_spl_)
  );


  LA
  g_g151_p
  (
    .dout(g151_p),
    .din1(g148_n_spl_),
    .din2(g149_p_spl_)
  );


  FA
  g_g151_n
  (
    .dout(g151_n),
    .din1(g148_p_spl_),
    .din2(g149_n_spl_0)
  );


  LA
  g_g152_p
  (
    .dout(g152_p),
    .din1(g150_n),
    .din2(g151_n)
  );


  FA
  g_g152_n
  (
    .dout(g152_n),
    .din1(g150_p),
    .din2(g151_p)
  );


  LA
  g_g153_p
  (
    .dout(g153_p),
    .din1(g130_p),
    .din2(g152_p)
  );


  FA
  g_g153_n
  (
    .dout(g153_n),
    .din1(g130_n),
    .din2(g152_n)
  );


  LA
  g_g154_p
  (
    .dout(g154_p),
    .din1(g109_n),
    .din2(g153_p)
  );


  FA
  g_g154_n
  (
    .dout(g154_n),
    .din1(g109_p),
    .din2(g153_n)
  );


  LA
  g_g155_p
  (
    .dout(g155_p),
    .din1(G17_p_spl_),
    .din2(G33_n_spl_011)
  );


  FA
  g_g155_n
  (
    .dout(g155_n),
    .din1(G17_n_spl_),
    .din2(G33_p_spl_01)
  );


  LA
  g_g156_p
  (
    .dout(g156_p),
    .din1(G24_n_spl_1),
    .din2(g155_p)
  );


  FA
  g_g156_n
  (
    .dout(g156_n),
    .din1(G24_p_spl_1),
    .din2(g155_n)
  );


  LA
  g_g157_p
  (
    .dout(g157_p),
    .din1(G1_p_spl_0),
    .din2(g156_p_spl_)
  );


  FA
  g_g157_n
  (
    .dout(g157_n),
    .din1(G1_n_spl_0),
    .din2(g156_n_spl_)
  );


  LA
  g_g158_p
  (
    .dout(g158_p),
    .din1(G1_n_spl_1),
    .din2(g156_n_spl_)
  );


  FA
  g_g158_n
  (
    .dout(g158_n),
    .din1(G1_p_spl_1),
    .din2(g156_p_spl_)
  );


  LA
  g_g159_p
  (
    .dout(g159_p),
    .din1(g157_n),
    .din2(g158_n)
  );


  FA
  g_g159_n
  (
    .dout(g159_n),
    .din1(g157_p),
    .din2(g158_p)
  );


  LA
  g_g160_p
  (
    .dout(g160_p),
    .din1(G6_p_spl_0),
    .din2(G7_n_spl_0)
  );


  FA
  g_g160_n
  (
    .dout(g160_n),
    .din1(G6_n_spl_0),
    .din2(G7_p_spl_0)
  );


  LA
  g_g161_p
  (
    .dout(g161_p),
    .din1(G6_n_spl_1),
    .din2(G7_p_spl_1)
  );


  FA
  g_g161_n
  (
    .dout(g161_n),
    .din1(G6_p_spl_1),
    .din2(G7_n_spl_1)
  );


  LA
  g_g162_p
  (
    .dout(g162_p),
    .din1(g160_n),
    .din2(g161_n)
  );


  FA
  g_g162_n
  (
    .dout(g162_n),
    .din1(g160_p),
    .din2(g161_p)
  );


  LA
  g_g163_p
  (
    .dout(g163_p),
    .din1(G5_p_spl_0),
    .din2(g162_p_spl_)
  );


  FA
  g_g163_n
  (
    .dout(g163_n),
    .din1(G5_n_spl_0),
    .din2(g162_n_spl_)
  );


  LA
  g_g164_p
  (
    .dout(g164_p),
    .din1(G5_n_spl_1),
    .din2(g162_n_spl_)
  );


  FA
  g_g164_n
  (
    .dout(g164_n),
    .din1(G5_p_spl_1),
    .din2(g162_p_spl_)
  );


  LA
  g_g165_p
  (
    .dout(g165_p),
    .din1(g163_n),
    .din2(g164_n)
  );


  FA
  g_g165_n
  (
    .dout(g165_n),
    .din1(g163_p),
    .din2(g164_p)
  );


  LA
  g_g166_p
  (
    .dout(g166_p),
    .din1(g64_n_spl_01),
    .din2(g165_n_spl_0)
  );


  FA
  g_g166_n
  (
    .dout(g166_n),
    .din1(g64_p_spl_01),
    .din2(g165_p_spl_0)
  );


  LA
  g_g167_p
  (
    .dout(g167_p),
    .din1(g64_p_spl_01),
    .din2(g165_p_spl_0)
  );


  FA
  g_g167_n
  (
    .dout(g167_n),
    .din1(g64_n_spl_01),
    .din2(g165_n_spl_0)
  );


  LA
  g_g168_p
  (
    .dout(g168_p),
    .din1(g166_n),
    .din2(g167_n)
  );


  FA
  g_g168_n
  (
    .dout(g168_n),
    .din1(g166_p),
    .din2(g167_p)
  );


  LA
  g_g169_p
  (
    .dout(g169_p),
    .din1(g159_p_spl_),
    .din2(g168_p_spl_)
  );


  FA
  g_g169_n
  (
    .dout(g169_n),
    .din1(g159_n_spl_),
    .din2(g168_n_spl_)
  );


  LA
  g_g170_p
  (
    .dout(g170_p),
    .din1(g159_n_spl_),
    .din2(g168_n_spl_)
  );


  FA
  g_g170_n
  (
    .dout(g170_n),
    .din1(g159_p_spl_),
    .din2(g168_p_spl_)
  );


  LA
  g_g171_p
  (
    .dout(g171_p),
    .din1(g169_n),
    .din2(g170_n)
  );


  FA
  g_g171_n
  (
    .dout(g171_n),
    .din1(g169_p),
    .din2(g170_p)
  );


  LA
  g_g172_p
  (
    .dout(g172_p),
    .din1(G31_n_spl_011),
    .din2(g171_n_spl_)
  );


  FA
  g_g172_n
  (
    .dout(g172_n),
    .din1(G31_p_spl_011),
    .din2(g171_p_spl_)
  );


  LA
  g_g173_p
  (
    .dout(g173_p),
    .din1(G26_p_spl_0),
    .din2(g172_n_spl_)
  );


  FA
  g_g173_n
  (
    .dout(g173_n),
    .din1(G26_n_spl_0),
    .din2(g172_p_spl_)
  );


  LA
  g_g174_p
  (
    .dout(g174_p),
    .din1(G27_p_spl_),
    .din2(g108_n_spl_)
  );


  FA
  g_g174_n
  (
    .dout(g174_n),
    .din1(G27_n_spl_0),
    .din2(g108_p_spl_)
  );


  LA
  g_g175_p
  (
    .dout(g175_p),
    .din1(G26_n_spl_0),
    .din2(g172_p_spl_)
  );


  FA
  g_g175_n
  (
    .dout(g175_n),
    .din1(G26_p_spl_0),
    .din2(g172_n_spl_)
  );


  LA
  g_g176_p
  (
    .dout(g176_p),
    .din1(g174_n),
    .din2(g175_n)
  );


  FA
  g_g176_n
  (
    .dout(g176_n),
    .din1(g174_p),
    .din2(g175_p)
  );


  LA
  g_g177_p
  (
    .dout(g177_p),
    .din1(g173_n),
    .din2(g176_p)
  );


  FA
  g_g177_n
  (
    .dout(g177_n),
    .din1(g173_p),
    .din2(g176_n)
  );


  LA
  g_g178_p
  (
    .dout(g178_p),
    .din1(g154_p),
    .din2(g177_p)
  );


  FA
  g_g178_n
  (
    .dout(g178_n),
    .din1(g154_n),
    .din2(g177_n)
  );


  LA
  g_g179_p
  (
    .dout(g179_p),
    .din1(G24_n_spl_1),
    .din2(G31_n_spl_011)
  );


  FA
  g_g179_n
  (
    .dout(g179_n),
    .din1(G24_p_spl_1),
    .din2(G31_p_spl_011)
  );


  LA
  g_g180_p
  (
    .dout(g180_p),
    .din1(G18_p_spl_),
    .din2(g179_n_spl_)
  );


  FA
  g_g180_n
  (
    .dout(g180_n),
    .din1(G18_n_spl_),
    .din2(g179_p_spl_)
  );


  LA
  g_g181_p
  (
    .dout(g181_p),
    .din1(G21_p_spl_),
    .din2(G33_n_spl_011)
  );


  FA
  g_g181_n
  (
    .dout(g181_n),
    .din1(G21_n_spl_),
    .din2(G33_p_spl_10)
  );


  LA
  g_g182_p
  (
    .dout(g182_p),
    .din1(G9_p_spl_0),
    .din2(g61_n_spl_1)
  );


  FA
  g_g182_n
  (
    .dout(g182_n),
    .din1(G9_n_spl_0),
    .din2(g61_p_spl_1)
  );


  LA
  g_g183_p
  (
    .dout(g183_p),
    .din1(G9_n_spl_1),
    .din2(g61_p_spl_1)
  );


  FA
  g_g183_n
  (
    .dout(g183_n),
    .din1(G9_p_spl_1),
    .din2(g61_n_spl_1)
  );


  LA
  g_g184_p
  (
    .dout(g184_p),
    .din1(g182_n),
    .din2(g183_n)
  );


  FA
  g_g184_n
  (
    .dout(g184_n),
    .din1(g182_p),
    .din2(g183_p)
  );


  LA
  g_g185_p
  (
    .dout(g185_p),
    .din1(g181_p_spl_),
    .din2(g184_p_spl_)
  );


  FA
  g_g185_n
  (
    .dout(g185_n),
    .din1(g181_n_spl_),
    .din2(g184_n_spl_)
  );


  LA
  g_g186_p
  (
    .dout(g186_p),
    .din1(g181_n_spl_),
    .din2(g184_n_spl_)
  );


  FA
  g_g186_n
  (
    .dout(g186_n),
    .din1(g181_p_spl_),
    .din2(g184_p_spl_)
  );


  LA
  g_g187_p
  (
    .dout(g187_p),
    .din1(g185_n),
    .din2(g186_n)
  );


  FA
  g_g187_n
  (
    .dout(g187_n),
    .din1(g185_p),
    .din2(g186_p)
  );


  LA
  g_g188_p
  (
    .dout(g188_p),
    .din1(g70_n_spl_1),
    .din2(g165_p_spl_1)
  );


  FA
  g_g188_n
  (
    .dout(g188_n),
    .din1(g70_p_spl_1),
    .din2(g165_n_spl_1)
  );


  LA
  g_g189_p
  (
    .dout(g189_p),
    .din1(g70_p_spl_1),
    .din2(g165_n_spl_1)
  );


  FA
  g_g189_n
  (
    .dout(g189_n),
    .din1(g70_n_spl_1),
    .din2(g165_p_spl_1)
  );


  LA
  g_g190_p
  (
    .dout(g190_p),
    .din1(g188_n),
    .din2(g189_n)
  );


  FA
  g_g190_n
  (
    .dout(g190_n),
    .din1(g188_p),
    .din2(g189_p)
  );


  LA
  g_g191_p
  (
    .dout(g191_p),
    .din1(G4_n_spl_10),
    .din2(G8_n_spl_10)
  );


  FA
  g_g191_n
  (
    .dout(g191_n),
    .din1(G4_p_spl_10),
    .din2(G8_p_spl_10)
  );


  LA
  g_g192_p
  (
    .dout(g192_p),
    .din1(G4_p_spl_10),
    .din2(G8_p_spl_10)
  );


  FA
  g_g192_n
  (
    .dout(g192_n),
    .din1(G4_n_spl_10),
    .din2(G8_n_spl_10)
  );


  LA
  g_g193_p
  (
    .dout(g193_p),
    .din1(g191_n),
    .din2(g192_n)
  );


  FA
  g_g193_n
  (
    .dout(g193_n),
    .din1(g191_p),
    .din2(g192_p)
  );


  LA
  g_g194_p
  (
    .dout(g194_p),
    .din1(g190_p_spl_),
    .din2(g193_n_spl_)
  );


  FA
  g_g194_n
  (
    .dout(g194_n),
    .din1(g190_n_spl_),
    .din2(g193_p_spl_)
  );


  LA
  g_g195_p
  (
    .dout(g195_p),
    .din1(g190_n_spl_),
    .din2(g193_p_spl_)
  );


  FA
  g_g195_n
  (
    .dout(g195_n),
    .din1(g190_p_spl_),
    .din2(g193_n_spl_)
  );


  LA
  g_g196_p
  (
    .dout(g196_p),
    .din1(g194_n),
    .din2(g195_n)
  );


  FA
  g_g196_n
  (
    .dout(g196_n),
    .din1(g194_p),
    .din2(g195_p)
  );


  LA
  g_g197_p
  (
    .dout(g197_p),
    .din1(g187_p_spl_),
    .din2(g196_n_spl_0)
  );


  FA
  g_g197_n
  (
    .dout(g197_n),
    .din1(g187_n_spl_),
    .din2(g196_p_spl_0)
  );


  LA
  g_g198_p
  (
    .dout(g198_p),
    .din1(g187_n_spl_),
    .din2(g196_p_spl_0)
  );


  FA
  g_g198_n
  (
    .dout(g198_n),
    .din1(g187_p_spl_),
    .din2(g196_n_spl_0)
  );


  LA
  g_g199_p
  (
    .dout(g199_p),
    .din1(g197_n),
    .din2(g198_n)
  );


  FA
  g_g199_n
  (
    .dout(g199_n),
    .din1(g197_p),
    .din2(g198_p)
  );


  LA
  g_g200_p
  (
    .dout(g200_p),
    .din1(G31_n_spl_10),
    .din2(g199_p_spl_)
  );


  FA
  g_g200_n
  (
    .dout(g200_n),
    .din1(G31_p_spl_100),
    .din2(g199_n_spl_)
  );


  LA
  g_g201_p
  (
    .dout(g201_p),
    .din1(G17_p_spl_),
    .din2(g179_n_spl_)
  );


  FA
  g_g201_n
  (
    .dout(g201_n),
    .din1(G17_n_spl_),
    .din2(g179_p_spl_)
  );


  LA
  g_g202_p
  (
    .dout(g202_p),
    .din1(g200_p_spl_),
    .din2(g201_n_spl_0)
  );


  FA
  g_g202_n
  (
    .dout(g202_n),
    .din1(g200_n_spl_),
    .din2(g201_p_spl_0)
  );


  LA
  g_g203_p
  (
    .dout(g203_p),
    .din1(g200_n_spl_),
    .din2(g201_p_spl_0)
  );


  FA
  g_g203_n
  (
    .dout(g203_n),
    .din1(g200_p_spl_),
    .din2(g201_n_spl_0)
  );


  LA
  g_g204_p
  (
    .dout(g204_p),
    .din1(g202_n),
    .din2(g203_n)
  );


  FA
  g_g204_n
  (
    .dout(g204_n),
    .din1(g202_p),
    .din2(g203_p)
  );


  LA
  g_g205_p
  (
    .dout(g205_p),
    .din1(g180_p_spl_0),
    .din2(g204_n_spl_0)
  );


  FA
  g_g205_n
  (
    .dout(g205_n),
    .din1(g180_n_spl_),
    .din2(g204_p_spl_)
  );


  LA
  g_g206_p
  (
    .dout(g206_p),
    .din1(g178_p_spl_),
    .din2(g205_n)
  );


  FA
  g_g206_n
  (
    .dout(g206_n),
    .din1(g178_n_spl_0),
    .din2(g205_p)
  );


  LA
  g_g207_p
  (
    .dout(g207_p),
    .din1(g81_n_spl_),
    .din2(g206_p_spl_)
  );


  FA
  g_g207_n
  (
    .dout(g207_n),
    .din1(g81_p_spl_),
    .din2(g206_n_spl_)
  );


  LA
  g_g208_p
  (
    .dout(g208_p),
    .din1(g40_n_spl_),
    .din2(g207_p_spl_)
  );


  FA
  g_g208_n
  (
    .dout(g208_n),
    .din1(g40_p_spl_),
    .din2(g207_n_spl_)
  );


  LA
  g_g209_p
  (
    .dout(g209_p),
    .din1(G1_p_spl_1),
    .din2(g208_n_spl_00)
  );


  LA
  g_g210_p
  (
    .dout(g210_p),
    .din1(G1_n_spl_1),
    .din2(g208_p_spl_00)
  );


  FA
  g_g211_n
  (
    .dout(g211_n),
    .din1(g209_p),
    .din2(g210_p)
  );


  LA
  g_g212_p
  (
    .dout(g212_p),
    .din1(G2_p_spl_1),
    .din2(g208_n_spl_00)
  );


  LA
  g_g213_p
  (
    .dout(g213_p),
    .din1(G2_n_spl_1),
    .din2(g208_p_spl_00)
  );


  FA
  g_g214_n
  (
    .dout(g214_n),
    .din1(g212_p),
    .din2(g213_p)
  );


  LA
  g_g215_p
  (
    .dout(g215_p),
    .din1(G3_p_spl_1),
    .din2(g208_n_spl_01)
  );


  LA
  g_g216_p
  (
    .dout(g216_p),
    .din1(G3_n_spl_1),
    .din2(g208_p_spl_01)
  );


  FA
  g_g217_n
  (
    .dout(g217_n),
    .din1(g215_p),
    .din2(g216_p)
  );


  LA
  g_g218_p
  (
    .dout(g218_p),
    .din1(G4_p_spl_1),
    .din2(g208_n_spl_01)
  );


  LA
  g_g219_p
  (
    .dout(g219_p),
    .din1(G4_n_spl_1),
    .din2(g208_p_spl_01)
  );


  FA
  g_g220_n
  (
    .dout(g220_n),
    .din1(g218_p),
    .din2(g219_p)
  );


  LA
  g_g221_p
  (
    .dout(g221_p),
    .din1(G30_n_spl_),
    .din2(G33_n_spl_10)
  );


  FA
  g_g221_n
  (
    .dout(g221_n),
    .din1(G30_p_spl_),
    .din2(G33_p_spl_10)
  );


  LA
  g_g222_p
  (
    .dout(g222_p),
    .din1(g36_p_spl_),
    .din2(g221_p_spl_)
  );


  FA
  g_g222_n
  (
    .dout(g222_n),
    .din1(g36_n_spl_),
    .din2(g221_n_spl_)
  );


  LA
  g_g223_p
  (
    .dout(g223_p),
    .din1(g39_n_spl_),
    .din2(g222_n)
  );


  FA
  g_g223_n
  (
    .dout(g223_n),
    .din1(g39_p_spl_),
    .din2(g222_p)
  );


  LA
  g_g224_p
  (
    .dout(g224_p),
    .din1(g207_p_spl_),
    .din2(g223_n_spl_0)
  );


  FA
  g_g224_n
  (
    .dout(g224_n),
    .din1(g207_n_spl_),
    .din2(g223_p_spl_0)
  );


  LA
  g_g225_p
  (
    .dout(g225_p),
    .din1(G10_p_spl_1),
    .din2(g224_n_spl_00)
  );


  LA
  g_g226_p
  (
    .dout(g226_p),
    .din1(G10_n_spl_1),
    .din2(g224_p_spl_00)
  );


  FA
  g_g227_n
  (
    .dout(g227_n),
    .din1(g225_p),
    .din2(g226_p)
  );


  LA
  g_g228_p
  (
    .dout(g228_p),
    .din1(G15_p_spl_1),
    .din2(g224_n_spl_00)
  );


  LA
  g_g229_p
  (
    .dout(g229_p),
    .din1(G15_n_spl_1),
    .din2(g224_p_spl_00)
  );


  FA
  g_g230_n
  (
    .dout(g230_n),
    .din1(g228_p),
    .din2(g229_p)
  );


  LA
  g_g231_p
  (
    .dout(g231_p),
    .din1(G16_p_spl_1),
    .din2(g224_n_spl_01)
  );


  LA
  g_g232_p
  (
    .dout(g232_p),
    .din1(G16_n_spl_1),
    .din2(g224_p_spl_01)
  );


  FA
  g_g233_n
  (
    .dout(g233_n),
    .din1(g231_p),
    .din2(g232_p)
  );


  LA
  g_g234_p
  (
    .dout(g234_p),
    .din1(g42_p_spl_0),
    .din2(g80_p_spl_)
  );


  FA
  g_g234_n
  (
    .dout(g234_n),
    .din1(g42_n_spl_),
    .din2(g80_n_spl_0)
  );


  LA
  g_g235_p
  (
    .dout(g235_p),
    .din1(g206_p_spl_),
    .din2(g234_p)
  );


  FA
  g_g235_n
  (
    .dout(g235_n),
    .din1(g206_n_spl_),
    .din2(g234_n)
  );


  LA
  g_g236_p
  (
    .dout(g236_p),
    .din1(g40_n_spl_),
    .din2(g235_p_spl_)
  );


  FA
  g_g236_n
  (
    .dout(g236_n),
    .din1(g40_p_spl_),
    .din2(g235_n_spl_)
  );


  LA
  g_g237_p
  (
    .dout(g237_p),
    .din1(G5_p_spl_1),
    .din2(g236_n_spl_0)
  );


  LA
  g_g238_p
  (
    .dout(g238_p),
    .din1(G5_n_spl_1),
    .din2(g236_p_spl_0)
  );


  FA
  g_g239_n
  (
    .dout(g239_n),
    .din1(g237_p),
    .din2(g238_p)
  );


  LA
  g_g240_p
  (
    .dout(g240_p),
    .din1(G6_p_spl_1),
    .din2(g236_n_spl_0)
  );


  LA
  g_g241_p
  (
    .dout(g241_p),
    .din1(G6_n_spl_1),
    .din2(g236_p_spl_0)
  );


  FA
  g_g242_n
  (
    .dout(g242_n),
    .din1(g240_p),
    .din2(g241_p)
  );


  LA
  g_g243_p
  (
    .dout(g243_p),
    .din1(G7_p_spl_1),
    .din2(g236_n_spl_1)
  );


  LA
  g_g244_p
  (
    .dout(g244_p),
    .din1(G7_n_spl_1),
    .din2(g236_p_spl_1)
  );


  FA
  g_g245_n
  (
    .dout(g245_n),
    .din1(g243_p),
    .din2(g244_p)
  );


  LA
  g_g246_p
  (
    .dout(g246_p),
    .din1(G8_p_spl_1),
    .din2(g236_n_spl_1)
  );


  LA
  g_g247_p
  (
    .dout(g247_p),
    .din1(G8_n_spl_1),
    .din2(g236_p_spl_1)
  );


  FA
  g_g248_n
  (
    .dout(g248_n),
    .din1(g246_p),
    .din2(g247_p)
  );


  LA
  g_g249_p
  (
    .dout(g249_p),
    .din1(g223_n_spl_0),
    .din2(g235_p_spl_)
  );


  FA
  g_g249_n
  (
    .dout(g249_n),
    .din1(g223_p_spl_0),
    .din2(g235_n_spl_)
  );


  FA
  g_g250_n
  (
    .dout(g250_n),
    .din1(G9_n_spl_1),
    .din2(g249_n)
  );


  FA
  g_g251_n
  (
    .dout(g251_n),
    .din1(G9_p_spl_1),
    .din2(g249_p)
  );


  LA
  g_g252_p
  (
    .dout(g252_p),
    .din1(g250_n),
    .din2(g251_n)
  );


  LA
  g_g253_p
  (
    .dout(g253_p),
    .din1(g178_p_spl_),
    .din2(g180_p_spl_0)
  );


  FA
  g_g253_n
  (
    .dout(g253_n),
    .din1(g178_n_spl_0),
    .din2(g180_n_spl_)
  );


  LA
  g_g254_p
  (
    .dout(g254_p),
    .din1(g81_n_spl_),
    .din2(g223_n_spl_)
  );


  FA
  g_g254_n
  (
    .dout(g254_n),
    .din1(g81_p_spl_),
    .din2(g223_p_spl_)
  );


  LA
  g_g255_p
  (
    .dout(g255_p),
    .din1(g204_p_spl_),
    .din2(g254_p)
  );


  FA
  g_g255_n
  (
    .dout(g255_n),
    .din1(g204_n_spl_0),
    .din2(g254_n)
  );


  LA
  g_g256_p
  (
    .dout(g256_p),
    .din1(g253_p),
    .din2(g255_p)
  );


  FA
  g_g256_n
  (
    .dout(g256_n),
    .din1(g253_n),
    .din2(g255_n)
  );


  LA
  g_g257_p
  (
    .dout(g257_p),
    .din1(G11_p_spl_1),
    .din2(g256_n_spl_0)
  );


  LA
  g_g258_p
  (
    .dout(g258_p),
    .din1(G11_n_spl_1),
    .din2(g256_p_spl_0)
  );


  FA
  g_g259_n
  (
    .dout(g259_n),
    .din1(g257_p),
    .din2(g258_p)
  );


  LA
  g_g260_p
  (
    .dout(g260_p),
    .din1(G12_p_spl_1),
    .din2(g256_n_spl_0)
  );


  LA
  g_g261_p
  (
    .dout(g261_p),
    .din1(G12_n_spl_1),
    .din2(g256_p_spl_0)
  );


  FA
  g_g262_n
  (
    .dout(g262_n),
    .din1(g260_p),
    .din2(g261_p)
  );


  LA
  g_g263_p
  (
    .dout(g263_p),
    .din1(G13_p_spl_1),
    .din2(g256_n_spl_1)
  );


  LA
  g_g264_p
  (
    .dout(g264_p),
    .din1(G13_n_spl_1),
    .din2(g256_p_spl_1)
  );


  FA
  g_g265_n
  (
    .dout(g265_n),
    .din1(g263_p),
    .din2(g264_p)
  );


  LA
  g_g266_p
  (
    .dout(g266_p),
    .din1(G14_p_spl_1),
    .din2(g256_n_spl_1)
  );


  LA
  g_g267_p
  (
    .dout(g267_p),
    .din1(G14_n_spl_1),
    .din2(g256_p_spl_1)
  );


  FA
  g_g268_n
  (
    .dout(g268_n),
    .din1(g266_p),
    .din2(g267_p)
  );


  LA
  g_g269_p
  (
    .dout(g269_p),
    .din1(g208_n_spl_10),
    .din2(g224_n_spl_01)
  );


  FA
  g_g269_n
  (
    .dout(g269_n),
    .din1(g208_p_spl_10),
    .din2(g224_p_spl_01)
  );


  FA
  g_g270_n
  (
    .dout(g270_n),
    .din1(G32_n_spl_),
    .din2(g269_p_spl_00)
  );


  FA
  g_g271_n
  (
    .dout(g271_n),
    .din1(g80_n_spl_),
    .din2(g204_n_spl_)
  );


  FA
  g_g272_n
  (
    .dout(g272_n),
    .din1(g42_p_spl_),
    .din2(g180_p_spl_)
  );


  FA
  g_g273_n
  (
    .dout(g273_n),
    .din1(g178_n_spl_),
    .din2(g272_n)
  );


  FA
  g_g274_n
  (
    .dout(g274_n),
    .din1(g271_n),
    .din2(g273_n)
  );


  LA
  g_g275_p
  (
    .dout(g275_p),
    .din1(g270_n),
    .din2(g274_n)
  );


  LA
  g_g276_p
  (
    .dout(g276_p),
    .din1(G33_n_spl_10),
    .din2(g275_p)
  );


  LA
  g_g277_p
  (
    .dout(g277_p),
    .din1(G31_n_spl_10),
    .din2(g201_p_spl_)
  );


  FA
  g_g277_n
  (
    .dout(g277_n),
    .din1(G31_p_spl_100),
    .din2(g201_n_spl_)
  );


  LA
  g_g278_p
  (
    .dout(g278_p),
    .din1(g269_n_spl_0),
    .din2(g277_p)
  );


  FA
  g_g278_n
  (
    .dout(g278_n),
    .din1(g269_p_spl_00),
    .din2(g277_n)
  );


  FA
  g_g279_n
  (
    .dout(g279_n),
    .din1(g199_n_spl_),
    .din2(g278_p)
  );


  FA
  g_g280_n
  (
    .dout(g280_n),
    .din1(g199_p_spl_),
    .din2(g278_n)
  );


  LA
  g_g281_p
  (
    .dout(g281_p),
    .din1(g279_n),
    .din2(g280_n)
  );


  FA
  g_g282_n
  (
    .dout(g282_n),
    .din1(g38_p_spl_00),
    .din2(g281_p)
  );


  LA
  g_g283_p
  (
    .dout(g283_p),
    .din1(G25_p_spl_),
    .din2(G31_n_spl_11)
  );


  FA
  g_g283_n
  (
    .dout(g283_n),
    .din1(G25_n_spl_),
    .din2(G31_p_spl_101)
  );


  LA
  g_g284_p
  (
    .dout(g284_p),
    .din1(g269_n_spl_0),
    .din2(g283_p)
  );


  FA
  g_g284_n
  (
    .dout(g284_n),
    .din1(g269_p_spl_01),
    .din2(g283_n)
  );


  FA
  g_g285_n
  (
    .dout(g285_n),
    .din1(g76_p_spl_),
    .din2(g284_p)
  );


  FA
  g_g286_n
  (
    .dout(g286_n),
    .din1(g76_n_spl_),
    .din2(g284_n)
  );


  LA
  g_g287_p
  (
    .dout(g287_p),
    .din1(g285_n),
    .din2(g286_n)
  );


  FA
  g_g288_n
  (
    .dout(g288_n),
    .din1(g38_p_spl_01),
    .din2(g287_p)
  );


  FA
  g_g289_n
  (
    .dout(g289_n),
    .din1(G27_n_spl_),
    .din2(G31_p_spl_101)
  );


  FA
  g_g290_n
  (
    .dout(g290_n),
    .din1(g269_p_spl_01),
    .din2(g289_n)
  );


  LA
  g_g291_p
  (
    .dout(g291_p),
    .din1(g107_n_spl_),
    .din2(g290_n)
  );


  FA
  g_g292_n
  (
    .dout(g292_n),
    .din1(g38_p_spl_01),
    .din2(g291_p)
  );


  FA
  g_g293_n
  (
    .dout(g293_n),
    .din1(G28_n_spl_),
    .din2(G31_p_spl_110)
  );


  FA
  g_g294_n
  (
    .dout(g294_n),
    .din1(g269_p_spl_10),
    .din2(g293_n)
  );


  LA
  g_g295_p
  (
    .dout(g295_p),
    .din1(g126_n_spl_),
    .din2(g294_n)
  );


  FA
  g_g296_n
  (
    .dout(g296_n),
    .din1(g38_p_spl_10),
    .din2(g295_p)
  );


  FA
  g_g297_n
  (
    .dout(g297_n),
    .din1(G31_p_spl_110),
    .din2(g149_n_spl_)
  );


  FA
  g_g298_n
  (
    .dout(g298_n),
    .din1(g269_p_spl_10),
    .din2(g297_n)
  );


  LA
  g_g299_p
  (
    .dout(g299_p),
    .din1(g147_n_spl_),
    .din2(g298_n)
  );


  FA
  g_g300_n
  (
    .dout(g300_n),
    .din1(g38_p_spl_10),
    .din2(g299_p)
  );


  LA
  g_g301_p
  (
    .dout(g301_p),
    .din1(G21_p_spl_),
    .din2(G29_p_spl_)
  );


  FA
  g_g301_n
  (
    .dout(g301_n),
    .din1(G21_n_spl_),
    .din2(G29_n_spl_)
  );


  LA
  g_g302_p
  (
    .dout(g302_p),
    .din1(G33_n_spl_11),
    .din2(g301_n)
  );


  FA
  g_g302_n
  (
    .dout(g302_n),
    .din1(G33_p_spl_11),
    .din2(g301_p)
  );


  LA
  g_g303_p
  (
    .dout(g303_p),
    .din1(g34_n_spl_),
    .din2(g196_p_spl_)
  );


  FA
  g_g303_n
  (
    .dout(g303_n),
    .din1(g34_p_spl_),
    .din2(g196_n_spl_)
  );


  LA
  g_g304_p
  (
    .dout(g304_p),
    .din1(g208_n_spl_10),
    .din2(g303_n_spl_)
  );


  FA
  g_g304_n
  (
    .dout(g304_n),
    .din1(g208_p_spl_10),
    .din2(g303_p_spl_)
  );


  LA
  g_g305_p
  (
    .dout(g305_p),
    .din1(g208_p_spl_1),
    .din2(g303_p_spl_)
  );


  FA
  g_g305_n
  (
    .dout(g305_n),
    .din1(g208_n_spl_1),
    .din2(g303_n_spl_)
  );


  LA
  g_g306_p
  (
    .dout(g306_p),
    .din1(g304_n),
    .din2(g305_n)
  );


  FA
  g_g306_n
  (
    .dout(g306_n),
    .din1(g304_p),
    .din2(g305_p)
  );


  FA
  g_g307_n
  (
    .dout(g307_n),
    .din1(g302_p),
    .din2(g306_n)
  );


  FA
  g_g308_n
  (
    .dout(g308_n),
    .din1(g302_n),
    .din2(g306_p)
  );


  LA
  g_g309_p
  (
    .dout(g309_p),
    .din1(g307_n),
    .din2(g308_n)
  );


  LA
  g_g310_p
  (
    .dout(g310_p),
    .din1(G22_p_spl_),
    .din2(G30_p_spl_)
  );


  FA
  g_g310_n
  (
    .dout(g310_n),
    .din1(G22_n_spl_),
    .din2(G30_n_spl_)
  );


  LA
  g_g311_p
  (
    .dout(g311_p),
    .din1(G33_n_spl_11),
    .din2(g310_n)
  );


  FA
  g_g311_n
  (
    .dout(g311_n),
    .din1(G33_p_spl_11),
    .din2(g310_p)
  );


  LA
  g_g312_p
  (
    .dout(g312_p),
    .din1(g64_p_spl_1),
    .din2(g92_n_spl_1)
  );


  FA
  g_g312_n
  (
    .dout(g312_n),
    .din1(g64_n_spl_1),
    .din2(g92_p_spl_1)
  );


  LA
  g_g313_p
  (
    .dout(g313_p),
    .din1(g64_n_spl_1),
    .din2(g92_p_spl_1)
  );


  FA
  g_g313_n
  (
    .dout(g313_n),
    .din1(g64_p_spl_1),
    .din2(g92_n_spl_1)
  );


  LA
  g_g314_p
  (
    .dout(g314_p),
    .din1(g312_n),
    .din2(g313_n)
  );


  FA
  g_g314_n
  (
    .dout(g314_n),
    .din1(g312_p),
    .din2(g313_p)
  );


  LA
  g_g315_p
  (
    .dout(g315_p),
    .din1(g221_n_spl_),
    .din2(g314_n)
  );


  FA
  g_g315_n
  (
    .dout(g315_n),
    .din1(g221_p_spl_),
    .din2(g314_p)
  );


  LA
  g_g316_p
  (
    .dout(g316_p),
    .din1(g224_n_spl_1),
    .din2(g315_n_spl_)
  );


  FA
  g_g316_n
  (
    .dout(g316_n),
    .din1(g224_p_spl_1),
    .din2(g315_p_spl_)
  );


  LA
  g_g317_p
  (
    .dout(g317_p),
    .din1(g224_p_spl_1),
    .din2(g315_p_spl_)
  );


  FA
  g_g317_n
  (
    .dout(g317_n),
    .din1(g224_n_spl_1),
    .din2(g315_n_spl_)
  );


  LA
  g_g318_p
  (
    .dout(g318_p),
    .din1(g316_n),
    .din2(g317_n)
  );


  FA
  g_g318_n
  (
    .dout(g318_n),
    .din1(g316_p),
    .din2(g317_p)
  );


  FA
  g_g319_n
  (
    .dout(g319_n),
    .din1(g311_p),
    .din2(g318_n)
  );


  FA
  g_g320_n
  (
    .dout(g320_n),
    .din1(g311_n),
    .din2(g318_p)
  );


  LA
  g_g321_p
  (
    .dout(g321_p),
    .din1(g319_n),
    .din2(g320_n)
  );


  LA
  g_g322_p
  (
    .dout(g322_p),
    .din1(G26_p_spl_),
    .din2(G31_n_spl_11)
  );


  FA
  g_g322_n
  (
    .dout(g322_n),
    .din1(G26_n_spl_),
    .din2(G31_p_spl_11)
  );


  LA
  g_g323_p
  (
    .dout(g323_p),
    .din1(g269_n_spl_),
    .din2(g322_p)
  );


  FA
  g_g323_n
  (
    .dout(g323_n),
    .din1(g269_p_spl_1),
    .din2(g322_n)
  );


  FA
  g_g324_n
  (
    .dout(g324_n),
    .din1(g171_p_spl_),
    .din2(g323_p)
  );


  FA
  g_g325_n
  (
    .dout(g325_n),
    .din1(g171_n_spl_),
    .din2(g323_n)
  );


  LA
  g_g326_p
  (
    .dout(g326_p),
    .din1(g324_n),
    .din2(g325_n)
  );


  FA
  g_g327_n
  (
    .dout(g327_n),
    .din1(g38_p_spl_1),
    .din2(g326_p)
  );


  buf

  (
    G1884_n,
    g211_n
  );


  buf

  (
    G1885_n,
    g214_n
  );


  buf

  (
    G1886_n,
    g217_n
  );


  buf

  (
    G1887_n,
    g220_n
  );


  buf

  (
    G1888_n,
    g227_n
  );


  buf

  (
    G1889_n,
    g230_n
  );


  buf

  (
    G1890_n,
    g233_n
  );


  buf

  (
    G1891_n,
    g239_n
  );


  buf

  (
    G1892_n,
    g242_n
  );


  buf

  (
    G1893_n,
    g245_n
  );


  buf

  (
    G1894_n,
    g248_n
  );


  buf

  (
    G1895_n,
    g252_p
  );


  buf

  (
    G1896_n,
    g259_n
  );


  buf

  (
    G1897_n,
    g262_n
  );


  buf

  (
    G1898_n,
    g265_n
  );


  buf

  (
    G1899_n,
    g268_n
  );


  buf

  (
    G1900_n,
    g276_p
  );


  buf

  (
    G1901_n,
    g282_n
  );


  buf

  (
    G1902_n,
    g288_n
  );


  buf

  (
    G1903_n,
    g292_n
  );


  buf

  (
    G1904_n,
    g296_n
  );


  buf

  (
    G1905_n,
    g300_n
  );


  buf

  (
    G1906_n,
    g309_p
  );


  buf

  (
    G1907_n,
    g321_p
  );


  buf

  (
    G1908_n,
    g327_n
  );


  buf

  (
    G29_n_spl_,
    G29_n
  );


  buf

  (
    G33_n_spl_,
    G33_n
  );


  buf

  (
    G33_n_spl_0,
    G33_n_spl_
  );


  buf

  (
    G33_n_spl_00,
    G33_n_spl_0
  );


  buf

  (
    G33_n_spl_000,
    G33_n_spl_00
  );


  buf

  (
    G33_n_spl_001,
    G33_n_spl_00
  );


  buf

  (
    G33_n_spl_01,
    G33_n_spl_0
  );


  buf

  (
    G33_n_spl_010,
    G33_n_spl_01
  );


  buf

  (
    G33_n_spl_011,
    G33_n_spl_01
  );


  buf

  (
    G33_n_spl_1,
    G33_n_spl_
  );


  buf

  (
    G33_n_spl_10,
    G33_n_spl_1
  );


  buf

  (
    G33_n_spl_11,
    G33_n_spl_1
  );


  buf

  (
    G29_p_spl_,
    G29_p
  );


  buf

  (
    G33_p_spl_,
    G33_p
  );


  buf

  (
    G33_p_spl_0,
    G33_p_spl_
  );


  buf

  (
    G33_p_spl_00,
    G33_p_spl_0
  );


  buf

  (
    G33_p_spl_000,
    G33_p_spl_00
  );


  buf

  (
    G33_p_spl_001,
    G33_p_spl_00
  );


  buf

  (
    G33_p_spl_01,
    G33_p_spl_0
  );


  buf

  (
    G33_p_spl_010,
    G33_p_spl_01
  );


  buf

  (
    G33_p_spl_1,
    G33_p_spl_
  );


  buf

  (
    G33_p_spl_10,
    G33_p_spl_1
  );


  buf

  (
    G33_p_spl_11,
    G33_p_spl_1
  );


  buf

  (
    G23_n_spl_,
    G23_n
  );


  buf

  (
    G23_n_spl_0,
    G23_n_spl_
  );


  buf

  (
    G23_n_spl_1,
    G23_n_spl_
  );


  buf

  (
    G24_p_spl_,
    G24_p
  );


  buf

  (
    G24_p_spl_0,
    G24_p_spl_
  );


  buf

  (
    G24_p_spl_1,
    G24_p_spl_
  );


  buf

  (
    G23_p_spl_,
    G23_p
  );


  buf

  (
    G23_p_spl_0,
    G23_p_spl_
  );


  buf

  (
    G23_p_spl_1,
    G23_p_spl_
  );


  buf

  (
    G24_n_spl_,
    G24_n
  );


  buf

  (
    G24_n_spl_0,
    G24_n_spl_
  );


  buf

  (
    G24_n_spl_1,
    G24_n_spl_
  );


  buf

  (
    G31_n_spl_,
    G31_n
  );


  buf

  (
    G31_n_spl_0,
    G31_n_spl_
  );


  buf

  (
    G31_n_spl_00,
    G31_n_spl_0
  );


  buf

  (
    G31_n_spl_000,
    G31_n_spl_00
  );


  buf

  (
    G31_n_spl_001,
    G31_n_spl_00
  );


  buf

  (
    G31_n_spl_01,
    G31_n_spl_0
  );


  buf

  (
    G31_n_spl_010,
    G31_n_spl_01
  );


  buf

  (
    G31_n_spl_011,
    G31_n_spl_01
  );


  buf

  (
    G31_n_spl_1,
    G31_n_spl_
  );


  buf

  (
    G31_n_spl_10,
    G31_n_spl_1
  );


  buf

  (
    G31_n_spl_11,
    G31_n_spl_1
  );


  buf

  (
    g35_n_spl_,
    g35_n
  );


  buf

  (
    G31_p_spl_,
    G31_p
  );


  buf

  (
    G31_p_spl_0,
    G31_p_spl_
  );


  buf

  (
    G31_p_spl_00,
    G31_p_spl_0
  );


  buf

  (
    G31_p_spl_000,
    G31_p_spl_00
  );


  buf

  (
    G31_p_spl_001,
    G31_p_spl_00
  );


  buf

  (
    G31_p_spl_01,
    G31_p_spl_0
  );


  buf

  (
    G31_p_spl_010,
    G31_p_spl_01
  );


  buf

  (
    G31_p_spl_011,
    G31_p_spl_01
  );


  buf

  (
    G31_p_spl_1,
    G31_p_spl_
  );


  buf

  (
    G31_p_spl_10,
    G31_p_spl_1
  );


  buf

  (
    G31_p_spl_100,
    G31_p_spl_10
  );


  buf

  (
    G31_p_spl_101,
    G31_p_spl_10
  );


  buf

  (
    G31_p_spl_11,
    G31_p_spl_1
  );


  buf

  (
    G31_p_spl_110,
    G31_p_spl_11
  );


  buf

  (
    g35_p_spl_,
    g35_p
  );


  buf

  (
    g34_p_spl_,
    g34_p
  );


  buf

  (
    g36_p_spl_,
    g36_p
  );


  buf

  (
    g34_n_spl_,
    g34_n
  );


  buf

  (
    g36_n_spl_,
    g36_n
  );


  buf

  (
    G32_n_spl_,
    G32_n
  );


  buf

  (
    g38_p_spl_,
    g38_p
  );


  buf

  (
    g38_p_spl_0,
    g38_p_spl_
  );


  buf

  (
    g38_p_spl_00,
    g38_p_spl_0
  );


  buf

  (
    g38_p_spl_01,
    g38_p_spl_0
  );


  buf

  (
    g38_p_spl_1,
    g38_p_spl_
  );


  buf

  (
    g38_p_spl_10,
    g38_p_spl_1
  );


  buf

  (
    g39_n_spl_,
    g39_n
  );


  buf

  (
    g39_p_spl_,
    g39_p
  );


  buf

  (
    G20_p_spl_,
    G20_p
  );


  buf

  (
    g41_n_spl_,
    g41_n
  );


  buf

  (
    G20_n_spl_,
    G20_n
  );


  buf

  (
    g41_p_spl_,
    g41_p
  );


  buf

  (
    G22_p_spl_,
    G22_p
  );


  buf

  (
    G22_n_spl_,
    G22_n
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_00,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_01,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_10,
    G4_p_spl_1
  );


  buf

  (
    G14_n_spl_,
    G14_n
  );


  buf

  (
    G14_n_spl_0,
    G14_n_spl_
  );


  buf

  (
    G14_n_spl_00,
    G14_n_spl_0
  );


  buf

  (
    G14_n_spl_1,
    G14_n_spl_
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    G4_n_spl_0,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_00,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_01,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_1,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_10,
    G4_n_spl_1
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G14_p_spl_0,
    G14_p_spl_
  );


  buf

  (
    G14_p_spl_00,
    G14_p_spl_0
  );


  buf

  (
    G14_p_spl_1,
    G14_p_spl_
  );


  buf

  (
    g43_p_spl_,
    g43_p
  );


  buf

  (
    g46_p_spl_,
    g46_p
  );


  buf

  (
    g43_n_spl_,
    g43_n
  );


  buf

  (
    g46_n_spl_,
    g46_n
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G12_p_spl_0,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_00,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_1,
    G12_p_spl_
  );


  buf

  (
    G13_n_spl_,
    G13_n
  );


  buf

  (
    G13_n_spl_0,
    G13_n_spl_
  );


  buf

  (
    G13_n_spl_00,
    G13_n_spl_0
  );


  buf

  (
    G13_n_spl_1,
    G13_n_spl_
  );


  buf

  (
    G12_n_spl_,
    G12_n
  );


  buf

  (
    G12_n_spl_0,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_00,
    G12_n_spl_0
  );


  buf

  (
    G12_n_spl_1,
    G12_n_spl_
  );


  buf

  (
    G13_p_spl_,
    G13_p
  );


  buf

  (
    G13_p_spl_0,
    G13_p_spl_
  );


  buf

  (
    G13_p_spl_00,
    G13_p_spl_0
  );


  buf

  (
    G13_p_spl_1,
    G13_p_spl_
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    G11_p_spl_0,
    G11_p_spl_
  );


  buf

  (
    G11_p_spl_00,
    G11_p_spl_0
  );


  buf

  (
    G11_p_spl_1,
    G11_p_spl_
  );


  buf

  (
    g52_p_spl_,
    g52_p
  );


  buf

  (
    G11_n_spl_,
    G11_n
  );


  buf

  (
    G11_n_spl_0,
    G11_n_spl_
  );


  buf

  (
    G11_n_spl_00,
    G11_n_spl_0
  );


  buf

  (
    G11_n_spl_1,
    G11_n_spl_
  );


  buf

  (
    g52_n_spl_,
    g52_n
  );


  buf

  (
    G10_n_spl_,
    G10_n
  );


  buf

  (
    G10_n_spl_0,
    G10_n_spl_
  );


  buf

  (
    G10_n_spl_00,
    G10_n_spl_0
  );


  buf

  (
    G10_n_spl_1,
    G10_n_spl_
  );


  buf

  (
    G15_n_spl_,
    G15_n
  );


  buf

  (
    G15_n_spl_0,
    G15_n_spl_
  );


  buf

  (
    G15_n_spl_00,
    G15_n_spl_0
  );


  buf

  (
    G15_n_spl_1,
    G15_n_spl_
  );


  buf

  (
    G10_p_spl_,
    G10_p
  );


  buf

  (
    G10_p_spl_0,
    G10_p_spl_
  );


  buf

  (
    G10_p_spl_00,
    G10_p_spl_0
  );


  buf

  (
    G10_p_spl_1,
    G10_p_spl_
  );


  buf

  (
    G15_p_spl_,
    G15_p
  );


  buf

  (
    G15_p_spl_0,
    G15_p_spl_
  );


  buf

  (
    G15_p_spl_00,
    G15_p_spl_0
  );


  buf

  (
    G15_p_spl_1,
    G15_p_spl_
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    G16_p_spl_0,
    G16_p_spl_
  );


  buf

  (
    G16_p_spl_00,
    G16_p_spl_0
  );


  buf

  (
    G16_p_spl_1,
    G16_p_spl_
  );


  buf

  (
    g58_n_spl_,
    g58_n
  );


  buf

  (
    g58_n_spl_0,
    g58_n_spl_
  );


  buf

  (
    g58_n_spl_1,
    g58_n_spl_
  );


  buf

  (
    G16_n_spl_,
    G16_n
  );


  buf

  (
    G16_n_spl_0,
    G16_n_spl_
  );


  buf

  (
    G16_n_spl_00,
    G16_n_spl_0
  );


  buf

  (
    G16_n_spl_1,
    G16_n_spl_
  );


  buf

  (
    g58_p_spl_,
    g58_p
  );


  buf

  (
    g58_p_spl_0,
    g58_p_spl_
  );


  buf

  (
    g58_p_spl_1,
    g58_p_spl_
  );


  buf

  (
    g55_n_spl_,
    g55_n
  );


  buf

  (
    g61_p_spl_,
    g61_p
  );


  buf

  (
    g61_p_spl_0,
    g61_p_spl_
  );


  buf

  (
    g61_p_spl_1,
    g61_p_spl_
  );


  buf

  (
    g55_p_spl_,
    g55_p
  );


  buf

  (
    g61_n_spl_,
    g61_n
  );


  buf

  (
    g61_n_spl_0,
    g61_n_spl_
  );


  buf

  (
    g61_n_spl_1,
    g61_n_spl_
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G2_p_spl_0,
    G2_p_spl_
  );


  buf

  (
    G2_p_spl_00,
    G2_p_spl_0
  );


  buf

  (
    G2_p_spl_1,
    G2_p_spl_
  );


  buf

  (
    G3_n_spl_,
    G3_n
  );


  buf

  (
    G3_n_spl_0,
    G3_n_spl_
  );


  buf

  (
    G3_n_spl_00,
    G3_n_spl_0
  );


  buf

  (
    G3_n_spl_1,
    G3_n_spl_
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G2_n_spl_0,
    G2_n_spl_
  );


  buf

  (
    G2_n_spl_00,
    G2_n_spl_0
  );


  buf

  (
    G2_n_spl_1,
    G2_n_spl_
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G3_p_spl_0,
    G3_p_spl_
  );


  buf

  (
    G3_p_spl_00,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_1,
    G3_p_spl_
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G1_p_spl_0,
    G1_p_spl_
  );


  buf

  (
    G1_p_spl_00,
    G1_p_spl_0
  );


  buf

  (
    G1_p_spl_1,
    G1_p_spl_
  );


  buf

  (
    g67_p_spl_,
    g67_p
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G1_n_spl_0,
    G1_n_spl_
  );


  buf

  (
    G1_n_spl_00,
    G1_n_spl_0
  );


  buf

  (
    G1_n_spl_1,
    G1_n_spl_
  );


  buf

  (
    g67_n_spl_,
    g67_n
  );


  buf

  (
    g64_n_spl_,
    g64_n
  );


  buf

  (
    g64_n_spl_0,
    g64_n_spl_
  );


  buf

  (
    g64_n_spl_00,
    g64_n_spl_0
  );


  buf

  (
    g64_n_spl_01,
    g64_n_spl_0
  );


  buf

  (
    g64_n_spl_1,
    g64_n_spl_
  );


  buf

  (
    g70_n_spl_,
    g70_n
  );


  buf

  (
    g70_n_spl_0,
    g70_n_spl_
  );


  buf

  (
    g70_n_spl_1,
    g70_n_spl_
  );


  buf

  (
    g64_p_spl_,
    g64_p
  );


  buf

  (
    g64_p_spl_0,
    g64_p_spl_
  );


  buf

  (
    g64_p_spl_00,
    g64_p_spl_0
  );


  buf

  (
    g64_p_spl_01,
    g64_p_spl_0
  );


  buf

  (
    g64_p_spl_1,
    g64_p_spl_
  );


  buf

  (
    g70_p_spl_,
    g70_p
  );


  buf

  (
    g70_p_spl_0,
    g70_p_spl_
  );


  buf

  (
    g70_p_spl_1,
    g70_p_spl_
  );


  buf

  (
    g49_n_spl_,
    g49_n
  );


  buf

  (
    g73_n_spl_,
    g73_n
  );


  buf

  (
    g49_p_spl_,
    g49_p
  );


  buf

  (
    g73_p_spl_,
    g73_p
  );


  buf

  (
    g76_n_spl_,
    g76_n
  );


  buf

  (
    g76_p_spl_,
    g76_p
  );


  buf

  (
    G25_n_spl_,
    G25_n
  );


  buf

  (
    G25_n_spl_0,
    G25_n_spl_
  );


  buf

  (
    g77_p_spl_,
    g77_p
  );


  buf

  (
    G25_p_spl_,
    G25_p
  );


  buf

  (
    G25_p_spl_0,
    G25_p_spl_
  );


  buf

  (
    g77_n_spl_,
    g77_n
  );


  buf

  (
    g42_p_spl_,
    g42_p
  );


  buf

  (
    g42_p_spl_0,
    g42_p_spl_
  );


  buf

  (
    g80_n_spl_,
    g80_n
  );


  buf

  (
    g80_n_spl_0,
    g80_n_spl_
  );


  buf

  (
    g42_n_spl_,
    g42_n
  );


  buf

  (
    g80_p_spl_,
    g80_p
  );


  buf

  (
    G18_p_spl_,
    G18_p
  );


  buf

  (
    G18_n_spl_,
    G18_n
  );


  buf

  (
    g83_n_spl_,
    g83_n
  );


  buf

  (
    g83_p_spl_,
    g83_p
  );


  buf

  (
    g86_n_spl_,
    g86_n
  );


  buf

  (
    g86_p_spl_,
    g86_p
  );


  buf

  (
    G9_p_spl_,
    G9_p
  );


  buf

  (
    G9_p_spl_0,
    G9_p_spl_
  );


  buf

  (
    G9_p_spl_00,
    G9_p_spl_0
  );


  buf

  (
    G9_p_spl_1,
    G9_p_spl_
  );


  buf

  (
    G9_n_spl_,
    G9_n
  );


  buf

  (
    G9_n_spl_0,
    G9_n_spl_
  );


  buf

  (
    G9_n_spl_00,
    G9_n_spl_0
  );


  buf

  (
    G9_n_spl_1,
    G9_n_spl_
  );


  buf

  (
    g92_n_spl_,
    g92_n
  );


  buf

  (
    g92_n_spl_0,
    g92_n_spl_
  );


  buf

  (
    g92_n_spl_1,
    g92_n_spl_
  );


  buf

  (
    g92_p_spl_,
    g92_p
  );


  buf

  (
    g92_p_spl_0,
    g92_p_spl_
  );


  buf

  (
    g92_p_spl_1,
    g92_p_spl_
  );


  buf

  (
    g89_p_spl_,
    g89_p
  );


  buf

  (
    g95_p_spl_,
    g95_p
  );


  buf

  (
    g95_p_spl_0,
    g95_p_spl_
  );


  buf

  (
    g95_p_spl_1,
    g95_p_spl_
  );


  buf

  (
    g89_n_spl_,
    g89_n
  );


  buf

  (
    g95_n_spl_,
    g95_n
  );


  buf

  (
    g95_n_spl_0,
    g95_n_spl_
  );


  buf

  (
    g95_n_spl_1,
    g95_n_spl_
  );


  buf

  (
    G5_n_spl_,
    G5_n
  );


  buf

  (
    G5_n_spl_0,
    G5_n_spl_
  );


  buf

  (
    G5_n_spl_00,
    G5_n_spl_0
  );


  buf

  (
    G5_n_spl_1,
    G5_n_spl_
  );


  buf

  (
    G8_n_spl_,
    G8_n
  );


  buf

  (
    G8_n_spl_0,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_00,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_01,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_1,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_10,
    G8_n_spl_1
  );


  buf

  (
    G5_p_spl_,
    G5_p
  );


  buf

  (
    G5_p_spl_0,
    G5_p_spl_
  );


  buf

  (
    G5_p_spl_00,
    G5_p_spl_0
  );


  buf

  (
    G5_p_spl_1,
    G5_p_spl_
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_00,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_01,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_1,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_10,
    G8_p_spl_1
  );


  buf

  (
    g101_p_spl_,
    g101_p
  );


  buf

  (
    g101_n_spl_,
    g101_n
  );


  buf

  (
    g98_n_spl_,
    g98_n
  );


  buf

  (
    g104_p_spl_,
    g104_p
  );


  buf

  (
    g98_p_spl_,
    g98_p
  );


  buf

  (
    g104_n_spl_,
    g104_n
  );


  buf

  (
    g107_n_spl_,
    g107_n
  );


  buf

  (
    G27_n_spl_,
    G27_n
  );


  buf

  (
    G27_n_spl_0,
    G27_n_spl_
  );


  buf

  (
    g108_p_spl_,
    g108_p
  );


  buf

  (
    G27_p_spl_,
    G27_p
  );


  buf

  (
    g108_n_spl_,
    g108_n
  );


  buf

  (
    G6_n_spl_,
    G6_n
  );


  buf

  (
    G6_n_spl_0,
    G6_n_spl_
  );


  buf

  (
    G6_n_spl_00,
    G6_n_spl_0
  );


  buf

  (
    G6_n_spl_1,
    G6_n_spl_
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G6_p_spl_0,
    G6_p_spl_
  );


  buf

  (
    G6_p_spl_00,
    G6_p_spl_0
  );


  buf

  (
    G6_p_spl_1,
    G6_p_spl_
  );


  buf

  (
    g112_p_spl_,
    g112_p
  );


  buf

  (
    g112_n_spl_,
    g112_n
  );


  buf

  (
    g115_n_spl_,
    g115_n
  );


  buf

  (
    g118_n_spl_,
    g118_n
  );


  buf

  (
    g115_p_spl_,
    g115_p
  );


  buf

  (
    g118_p_spl_,
    g118_p
  );


  buf

  (
    G19_p_spl_,
    G19_p
  );


  buf

  (
    G19_n_spl_,
    G19_n
  );


  buf

  (
    g121_n_spl_,
    g121_n
  );


  buf

  (
    g123_n_spl_,
    g123_n
  );


  buf

  (
    g121_p_spl_,
    g121_p
  );


  buf

  (
    g123_p_spl_,
    g123_p
  );


  buf

  (
    g126_n_spl_,
    g126_n
  );


  buf

  (
    G28_n_spl_,
    G28_n
  );


  buf

  (
    G28_n_spl_0,
    G28_n_spl_
  );


  buf

  (
    g127_p_spl_,
    g127_p
  );


  buf

  (
    G28_p_spl_,
    G28_p
  );


  buf

  (
    g127_n_spl_,
    g127_n
  );


  buf

  (
    G7_n_spl_,
    G7_n
  );


  buf

  (
    G7_n_spl_0,
    G7_n_spl_
  );


  buf

  (
    G7_n_spl_00,
    G7_n_spl_0
  );


  buf

  (
    G7_n_spl_1,
    G7_n_spl_
  );


  buf

  (
    G7_p_spl_,
    G7_p
  );


  buf

  (
    G7_p_spl_0,
    G7_p_spl_
  );


  buf

  (
    G7_p_spl_00,
    G7_p_spl_0
  );


  buf

  (
    G7_p_spl_1,
    G7_p_spl_
  );


  buf

  (
    g133_p_spl_,
    g133_p
  );


  buf

  (
    g133_n_spl_,
    g133_n
  );


  buf

  (
    g136_n_spl_,
    g136_n
  );


  buf

  (
    g136_p_spl_,
    g136_p
  );


  buf

  (
    g141_p_spl_,
    g141_p
  );


  buf

  (
    g141_n_spl_,
    g141_n
  );


  buf

  (
    g139_n_spl_,
    g139_n
  );


  buf

  (
    g144_n_spl_,
    g144_n
  );


  buf

  (
    g139_p_spl_,
    g139_p
  );


  buf

  (
    g144_p_spl_,
    g144_p
  );


  buf

  (
    g147_n_spl_,
    g147_n
  );


  buf

  (
    g148_p_spl_,
    g148_p
  );


  buf

  (
    g149_n_spl_,
    g149_n
  );


  buf

  (
    g149_n_spl_0,
    g149_n_spl_
  );


  buf

  (
    g148_n_spl_,
    g148_n
  );


  buf

  (
    g149_p_spl_,
    g149_p
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


  buf

  (
    G17_n_spl_,
    G17_n
  );


  buf

  (
    g156_p_spl_,
    g156_p
  );


  buf

  (
    g156_n_spl_,
    g156_n
  );


  buf

  (
    g162_p_spl_,
    g162_p
  );


  buf

  (
    g162_n_spl_,
    g162_n
  );


  buf

  (
    g165_n_spl_,
    g165_n
  );


  buf

  (
    g165_n_spl_0,
    g165_n_spl_
  );


  buf

  (
    g165_n_spl_1,
    g165_n_spl_
  );


  buf

  (
    g165_p_spl_,
    g165_p
  );


  buf

  (
    g165_p_spl_0,
    g165_p_spl_
  );


  buf

  (
    g165_p_spl_1,
    g165_p_spl_
  );


  buf

  (
    g159_p_spl_,
    g159_p
  );


  buf

  (
    g168_p_spl_,
    g168_p
  );


  buf

  (
    g159_n_spl_,
    g159_n
  );


  buf

  (
    g168_n_spl_,
    g168_n
  );


  buf

  (
    g171_n_spl_,
    g171_n
  );


  buf

  (
    g171_p_spl_,
    g171_p
  );


  buf

  (
    G26_p_spl_,
    G26_p
  );


  buf

  (
    G26_p_spl_0,
    G26_p_spl_
  );


  buf

  (
    g172_n_spl_,
    g172_n
  );


  buf

  (
    G26_n_spl_,
    G26_n
  );


  buf

  (
    G26_n_spl_0,
    G26_n_spl_
  );


  buf

  (
    g172_p_spl_,
    g172_p
  );


  buf

  (
    g179_n_spl_,
    g179_n
  );


  buf

  (
    g179_p_spl_,
    g179_p
  );


  buf

  (
    G21_p_spl_,
    G21_p
  );


  buf

  (
    G21_n_spl_,
    G21_n
  );


  buf

  (
    g181_p_spl_,
    g181_p
  );


  buf

  (
    g184_p_spl_,
    g184_p
  );


  buf

  (
    g181_n_spl_,
    g181_n
  );


  buf

  (
    g184_n_spl_,
    g184_n
  );


  buf

  (
    g190_p_spl_,
    g190_p
  );


  buf

  (
    g193_n_spl_,
    g193_n
  );


  buf

  (
    g190_n_spl_,
    g190_n
  );


  buf

  (
    g193_p_spl_,
    g193_p
  );


  buf

  (
    g187_p_spl_,
    g187_p
  );


  buf

  (
    g196_n_spl_,
    g196_n
  );


  buf

  (
    g196_n_spl_0,
    g196_n_spl_
  );


  buf

  (
    g187_n_spl_,
    g187_n
  );


  buf

  (
    g196_p_spl_,
    g196_p
  );


  buf

  (
    g196_p_spl_0,
    g196_p_spl_
  );


  buf

  (
    g199_p_spl_,
    g199_p
  );


  buf

  (
    g199_n_spl_,
    g199_n
  );


  buf

  (
    g200_p_spl_,
    g200_p
  );


  buf

  (
    g201_n_spl_,
    g201_n
  );


  buf

  (
    g201_n_spl_0,
    g201_n_spl_
  );


  buf

  (
    g200_n_spl_,
    g200_n
  );


  buf

  (
    g201_p_spl_,
    g201_p
  );


  buf

  (
    g201_p_spl_0,
    g201_p_spl_
  );


  buf

  (
    g180_p_spl_,
    g180_p
  );


  buf

  (
    g180_p_spl_0,
    g180_p_spl_
  );


  buf

  (
    g204_n_spl_,
    g204_n
  );


  buf

  (
    g204_n_spl_0,
    g204_n_spl_
  );


  buf

  (
    g180_n_spl_,
    g180_n
  );


  buf

  (
    g204_p_spl_,
    g204_p
  );


  buf

  (
    g178_p_spl_,
    g178_p
  );


  buf

  (
    g178_n_spl_,
    g178_n
  );


  buf

  (
    g178_n_spl_0,
    g178_n_spl_
  );


  buf

  (
    g81_n_spl_,
    g81_n
  );


  buf

  (
    g206_p_spl_,
    g206_p
  );


  buf

  (
    g81_p_spl_,
    g81_p
  );


  buf

  (
    g206_n_spl_,
    g206_n
  );


  buf

  (
    g40_n_spl_,
    g40_n
  );


  buf

  (
    g207_p_spl_,
    g207_p
  );


  buf

  (
    g40_p_spl_,
    g40_p
  );


  buf

  (
    g207_n_spl_,
    g207_n
  );


  buf

  (
    g208_n_spl_,
    g208_n
  );


  buf

  (
    g208_n_spl_0,
    g208_n_spl_
  );


  buf

  (
    g208_n_spl_00,
    g208_n_spl_0
  );


  buf

  (
    g208_n_spl_01,
    g208_n_spl_0
  );


  buf

  (
    g208_n_spl_1,
    g208_n_spl_
  );


  buf

  (
    g208_n_spl_10,
    g208_n_spl_1
  );


  buf

  (
    g208_p_spl_,
    g208_p
  );


  buf

  (
    g208_p_spl_0,
    g208_p_spl_
  );


  buf

  (
    g208_p_spl_00,
    g208_p_spl_0
  );


  buf

  (
    g208_p_spl_01,
    g208_p_spl_0
  );


  buf

  (
    g208_p_spl_1,
    g208_p_spl_
  );


  buf

  (
    g208_p_spl_10,
    g208_p_spl_1
  );


  buf

  (
    G30_n_spl_,
    G30_n
  );


  buf

  (
    G30_p_spl_,
    G30_p
  );


  buf

  (
    g221_p_spl_,
    g221_p
  );


  buf

  (
    g221_n_spl_,
    g221_n
  );


  buf

  (
    g223_n_spl_,
    g223_n
  );


  buf

  (
    g223_n_spl_0,
    g223_n_spl_
  );


  buf

  (
    g223_p_spl_,
    g223_p
  );


  buf

  (
    g223_p_spl_0,
    g223_p_spl_
  );


  buf

  (
    g224_n_spl_,
    g224_n
  );


  buf

  (
    g224_n_spl_0,
    g224_n_spl_
  );


  buf

  (
    g224_n_spl_00,
    g224_n_spl_0
  );


  buf

  (
    g224_n_spl_01,
    g224_n_spl_0
  );


  buf

  (
    g224_n_spl_1,
    g224_n_spl_
  );


  buf

  (
    g224_p_spl_,
    g224_p
  );


  buf

  (
    g224_p_spl_0,
    g224_p_spl_
  );


  buf

  (
    g224_p_spl_00,
    g224_p_spl_0
  );


  buf

  (
    g224_p_spl_01,
    g224_p_spl_0
  );


  buf

  (
    g224_p_spl_1,
    g224_p_spl_
  );


  buf

  (
    g235_p_spl_,
    g235_p
  );


  buf

  (
    g235_n_spl_,
    g235_n
  );


  buf

  (
    g236_n_spl_,
    g236_n
  );


  buf

  (
    g236_n_spl_0,
    g236_n_spl_
  );


  buf

  (
    g236_n_spl_1,
    g236_n_spl_
  );


  buf

  (
    g236_p_spl_,
    g236_p
  );


  buf

  (
    g236_p_spl_0,
    g236_p_spl_
  );


  buf

  (
    g236_p_spl_1,
    g236_p_spl_
  );


  buf

  (
    g256_n_spl_,
    g256_n
  );


  buf

  (
    g256_n_spl_0,
    g256_n_spl_
  );


  buf

  (
    g256_n_spl_1,
    g256_n_spl_
  );


  buf

  (
    g256_p_spl_,
    g256_p
  );


  buf

  (
    g256_p_spl_0,
    g256_p_spl_
  );


  buf

  (
    g256_p_spl_1,
    g256_p_spl_
  );


  buf

  (
    g269_p_spl_,
    g269_p
  );


  buf

  (
    g269_p_spl_0,
    g269_p_spl_
  );


  buf

  (
    g269_p_spl_00,
    g269_p_spl_0
  );


  buf

  (
    g269_p_spl_01,
    g269_p_spl_0
  );


  buf

  (
    g269_p_spl_1,
    g269_p_spl_
  );


  buf

  (
    g269_p_spl_10,
    g269_p_spl_1
  );


  buf

  (
    g269_n_spl_,
    g269_n
  );


  buf

  (
    g269_n_spl_0,
    g269_n_spl_
  );


  buf

  (
    g303_n_spl_,
    g303_n
  );


  buf

  (
    g303_p_spl_,
    g303_p
  );


  buf

  (
    g315_n_spl_,
    g315_n
  );


  buf

  (
    g315_p_spl_,
    g315_p
  );


endmodule
