
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  G42,
  G43,
  G44,
  G45,
  G46,
  G47,
  G48,
  G49,
  G50,
  G51,
  G52,
  G53,
  G54,
  G55,
  G56,
  G57,
  G58,
  G59,
  G60,
  G855,
  G856,
  G857,
  G858,
  G859,
  G860,
  G861,
  G862,
  G863,
  G864,
  G865,
  G866,
  G867,
  G868,
  G869,
  G870,
  G871,
  G872,
  G873,
  G874,
  G875,
  G876,
  G877,
  G878,
  G879,
  G880
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input G42;input G43;input G44;input G45;input G46;input G47;input G48;input G49;input G50;input G51;input G52;input G53;input G54;input G55;input G56;input G57;input G58;input G59;input G60;
  output G855;output G856;output G857;output G858;output G859;output G860;output G861;output G862;output G863;output G864;output G865;output G866;output G867;output G868;output G869;output G870;output G871;output G872;output G873;output G874;output G875;output G876;output G877;output G878;output G879;output G880;
  wire new_n87_;wire new_n89_;wire new_n93_;wire new_n94_;wire new_n96_;wire new_n97_;wire new_n98_;wire new_n100_;wire new_n102_;wire new_n105_;wire new_n109_;wire new_n110_;wire new_n112_;wire new_n113_;wire new_n116_;wire new_n117_;wire new_n118_;wire new_n119_;wire new_n120_;wire new_n121_;wire new_n122_;wire new_n123_;wire new_n124_;wire new_n125_;wire new_n126_;wire new_n127_;wire new_n128_;wire new_n129_;wire new_n130_;wire new_n131_;wire new_n132_;wire new_n133_;wire new_n134_;wire new_n135_;wire new_n136_;wire new_n137_;wire new_n138_;wire new_n139_;wire new_n140_;wire new_n141_;wire new_n143_;wire new_n144_;wire new_n145_;wire new_n146_;wire new_n147_;wire new_n148_;wire new_n149_;wire new_n150_;wire new_n151_;wire new_n152_;wire new_n153_;wire new_n154_;wire new_n155_;wire new_n156_;wire new_n157_;wire new_n158_;wire new_n159_;wire new_n160_;wire new_n161_;wire new_n162_;wire new_n163_;wire new_n164_;wire new_n165_;wire new_n166_;wire new_n167_;wire new_n168_;wire new_n170_;wire new_n171_;wire new_n172_;wire new_n173_;wire new_n174_;wire new_n175_;wire new_n176_;wire new_n177_;wire new_n178_;wire new_n179_;wire new_n180_;wire new_n181_;wire new_n182_;wire new_n183_;wire new_n184_;wire new_n185_;wire new_n186_;wire new_n187_;wire new_n188_;wire new_n189_;wire new_n190_;wire new_n191_;wire new_n192_;wire new_n193_;wire new_n194_;wire new_n195_;wire new_n196_;wire new_n197_;wire new_n198_;wire new_n199_;wire new_n200_;wire new_n201_;wire new_n202_;wire new_n203_;wire new_n204_;wire new_n205_;wire new_n206_;wire new_n207_;wire new_n208_;wire new_n209_;wire new_n210_;wire new_n211_;wire new_n212_;wire new_n213_;wire new_n215_;wire new_n216_;wire new_n217_;wire new_n218_;wire new_n219_;wire new_n220_;wire new_n221_;wire new_n222_;wire new_n223_;wire new_n224_;wire new_n225_;wire new_n226_;wire new_n227_;wire new_n228_;wire new_n229_;wire new_n230_;wire new_n231_;wire new_n232_;wire new_n233_;wire new_n234_;wire new_n235_;wire new_n236_;wire new_n237_;wire new_n238_;wire new_n239_;wire new_n240_;wire new_n241_;wire new_n242_;wire new_n243_;wire new_n244_;wire new_n245_;wire new_n246_;wire new_n247_;wire new_n248_;wire new_n249_;wire new_n250_;wire new_n251_;wire new_n253_;wire new_n254_;wire new_n255_;wire new_n256_;wire new_n257_;wire new_n258_;wire new_n259_;wire new_n260_;wire new_n261_;wire new_n262_;wire new_n263_;wire new_n264_;wire new_n265_;wire new_n266_;wire new_n267_;wire new_n269_;wire new_n270_;wire new_n271_;wire new_n272_;wire new_n273_;wire new_n274_;wire new_n275_;wire new_n276_;wire new_n277_;wire new_n278_;wire new_n279_;wire new_n280_;wire new_n281_;wire new_n282_;wire new_n283_;wire new_n285_;wire new_n286_;wire new_n287_;wire new_n288_;wire new_n289_;wire new_n290_;wire new_n291_;wire new_n292_;wire new_n293_;wire new_n294_;wire new_n295_;wire new_n296_;wire new_n297_;wire new_n298_;wire new_n299_;wire new_n300_;wire new_n301_;wire new_n302_;wire new_n303_;wire new_n304_;wire new_n305_;wire new_n306_;wire new_n307_;wire new_n308_;wire new_n309_;wire new_n310_;wire new_n311_;wire new_n312_;wire new_n313_;wire new_n314_;wire new_n315_;wire new_n316_;wire new_n317_;wire new_n318_;wire new_n319_;wire new_n320_;wire new_n321_;wire new_n322_;wire new_n323_;wire new_n324_;wire new_n325_;wire new_n326_;wire new_n327_;wire new_n329_;wire new_n330_;wire new_n331_;wire new_n332_;wire new_n333_;wire new_n334_;wire new_n335_;wire new_n336_;wire new_n337_;wire new_n338_;wire new_n339_;wire new_n340_;wire new_n341_;wire new_n342_;wire new_n344_;wire new_n345_;wire new_n346_;wire new_n347_;wire new_n348_;wire new_n349_;wire new_n350_;wire new_n351_;wire new_n352_;wire new_n353_;wire new_n354_;wire new_n355_;wire new_n356_;wire new_n357_;wire new_n359_;wire new_n360_;wire new_n361_;wire new_n362_;wire new_n363_;wire new_n364_;wire new_n365_;wire new_n366_;wire new_n367_;wire new_n368_;wire new_n369_;wire new_n370_;wire new_n371_;wire new_n372_;wire new_n374_;wire new_n375_;wire new_n376_;wire new_n377_;wire new_n378_;wire new_n379_;wire new_n380_;wire new_n381_;wire new_n382_;wire new_n383_;wire new_n384_;wire new_n385_;wire new_n386_;wire new_n387_;
  wire G6_spl_;
  wire G6_spl_0;
  wire G16_spl_;
  wire G8_spl_;
  wire G8_spl_0;
  wire G8_spl_00;
  wire G8_spl_01;
  wire G8_spl_1;
  wire G8_spl_10;
  wire new_n87__spl_;
  wire G7_spl_;
  wire G17_spl_;
  wire G17_spl_0;
  wire G17_spl_1;
  wire new_n89__spl_;
  wire G1_spl_;
  wire G1_spl_0;
  wire G2_spl_;
  wire G3_spl_;
  wire new_n93__spl_;
  wire G4_spl_;
  wire G4_spl_0;
  wire G4_spl_00;
  wire G4_spl_01;
  wire G4_spl_1;
  wire G4_spl_10;
  wire G4_spl_11;
  wire new_n94__spl_;
  wire new_n96__spl_;
  wire G857_spl_;
  wire new_n98__spl_;
  wire G11_spl_;
  wire G11_spl_0;
  wire G11_spl_1;
  wire new_n100__spl_;
  wire new_n102__spl_;
  wire new_n105__spl_;
  wire G9_spl_;
  wire G9_spl_0;
  wire G10_spl_;
  wire G10_spl_0;
  wire G12_spl_;
  wire new_n109__spl_;
  wire new_n109__spl_0;
  wire new_n112__spl_;
  wire G24_spl_;
  wire G24_spl_0;
  wire G24_spl_1;
  wire G25_spl_;
  wire G25_spl_0;
  wire G25_spl_1;
  wire G26_spl_;
  wire G26_spl_0;
  wire G26_spl_1;
  wire G27_spl_;
  wire G27_spl_0;
  wire G27_spl_1;
  wire new_n118__spl_;
  wire new_n121__spl_;
  wire G32_spl_;
  wire G32_spl_0;
  wire G32_spl_1;
  wire new_n124__spl_;
  wire G28_spl_;
  wire G28_spl_0;
  wire G28_spl_1;
  wire G29_spl_;
  wire G29_spl_0;
  wire G29_spl_1;
  wire G30_spl_;
  wire G30_spl_0;
  wire G30_spl_1;
  wire G31_spl_;
  wire G31_spl_0;
  wire new_n130__spl_;
  wire new_n133__spl_;
  wire G33_spl_;
  wire new_n136__spl_;
  wire new_n127__spl_;
  wire new_n139__spl_;
  wire G41_spl_;
  wire G41_spl_0;
  wire G41_spl_00;
  wire G41_spl_1;
  wire G42_spl_;
  wire G42_spl_0;
  wire G42_spl_00;
  wire G42_spl_1;
  wire G43_spl_;
  wire G43_spl_0;
  wire G43_spl_00;
  wire G43_spl_1;
  wire G44_spl_;
  wire G44_spl_0;
  wire G44_spl_00;
  wire G44_spl_1;
  wire new_n145__spl_;
  wire new_n148__spl_;
  wire new_n151__spl_;
  wire G45_spl_;
  wire G45_spl_0;
  wire G45_spl_00;
  wire G45_spl_1;
  wire G46_spl_;
  wire G46_spl_0;
  wire G46_spl_00;
  wire G46_spl_1;
  wire G47_spl_;
  wire G47_spl_0;
  wire G47_spl_00;
  wire G47_spl_1;
  wire G48_spl_;
  wire G48_spl_0;
  wire G48_spl_00;
  wire G48_spl_1;
  wire new_n157__spl_;
  wire new_n160__spl_;
  wire G49_spl_;
  wire new_n163__spl_;
  wire new_n154__spl_;
  wire new_n166__spl_;
  wire G866_spl_;
  wire G866_spl_0;
  wire new_n170__spl_;
  wire new_n171__spl_;
  wire G39_spl_;
  wire new_n173__spl_;
  wire new_n173__spl_0;
  wire new_n173__spl_1;
  wire G60_spl_;
  wire G60_spl_0;
  wire new_n176__spl_;
  wire new_n188__spl_;
  wire new_n188__spl_0;
  wire new_n188__spl_00;
  wire new_n188__spl_01;
  wire new_n188__spl_1;
  wire new_n188__spl_10;
  wire new_n188__spl_11;
  wire new_n178__spl_;
  wire new_n178__spl_0;
  wire new_n178__spl_1;
  wire new_n191__spl_;
  wire new_n191__spl_0;
  wire G53_spl_;
  wire G53_spl_0;
  wire G53_spl_00;
  wire G53_spl_01;
  wire G53_spl_1;
  wire G53_spl_10;
  wire G53_spl_11;
  wire new_n192__spl_;
  wire new_n192__spl_0;
  wire new_n194__spl_;
  wire G51_spl_;
  wire G51_spl_0;
  wire G51_spl_00;
  wire G51_spl_000;
  wire G51_spl_001;
  wire G51_spl_01;
  wire G51_spl_010;
  wire G51_spl_011;
  wire G51_spl_1;
  wire G51_spl_10;
  wire G51_spl_11;
  wire G58_spl_;
  wire new_n198__spl_;
  wire G52_spl_;
  wire G52_spl_0;
  wire G52_spl_00;
  wire G52_spl_01;
  wire G52_spl_1;
  wire G52_spl_10;
  wire G52_spl_11;
  wire G54_spl_;
  wire G54_spl_0;
  wire G54_spl_00;
  wire G54_spl_01;
  wire G54_spl_1;
  wire G54_spl_10;
  wire G54_spl_11;
  wire new_n207__spl_;
  wire new_n207__spl_0;
  wire new_n207__spl_00;
  wire new_n207__spl_01;
  wire new_n207__spl_1;
  wire new_n207__spl_10;
  wire new_n207__spl_11;
  wire G55_spl_;
  wire G55_spl_0;
  wire G50_spl_;
  wire G50_spl_0;
  wire G50_spl_00;
  wire G50_spl_01;
  wire G50_spl_1;
  wire G50_spl_10;
  wire G50_spl_11;
  wire G36_spl_;
  wire new_n218__spl_;
  wire new_n218__spl_0;
  wire G37_spl_;
  wire new_n224__spl_;
  wire new_n224__spl_0;
  wire new_n226__spl_;
  wire new_n227__spl_;
  wire new_n225__spl_;
  wire new_n225__spl_0;
  wire new_n228__spl_;
  wire new_n220__spl_;
  wire new_n229__spl_;
  wire new_n219__spl_;
  wire new_n219__spl_0;
  wire new_n230__spl_;
  wire new_n231__spl_;
  wire G35_spl_;
  wire new_n236__spl_;
  wire new_n236__spl_0;
  wire new_n237__spl_;
  wire new_n237__spl_0;
  wire new_n239__spl_;
  wire new_n242__spl_;
  wire new_n286__spl_;
  wire new_n286__spl_0;
  wire new_n286__spl_1;
  wire G34_spl_;
  wire G34_spl_0;
  wire G34_spl_1;
  wire new_n290__spl_;
  wire new_n290__spl_0;
  wire new_n290__spl_1;
  wire new_n293__spl_;
  wire new_n293__spl_0;
  wire new_n300__spl_;
  wire new_n300__spl_0;
  wire new_n308__spl_;
  wire new_n308__spl_0;
  wire new_n317__spl_;
  wire new_n317__spl_0;
  wire new_n311__spl_;
  wire new_n311__spl_0;
  wire new_n318__spl_;
  wire new_n320__spl_;
  wire new_n320__spl_0;
  wire new_n310__spl_;
  wire new_n321__spl_;
  wire new_n321__spl_0;
  wire new_n309__spl_;
  wire new_n309__spl_0;
  wire new_n302__spl_;
  wire new_n323__spl_;
  wire new_n323__spl_0;
  wire new_n301__spl_;
  wire new_n301__spl_0;
  wire new_n325__spl_;
  wire new_n325__spl_0;
  wire new_n326__spl_;
  wire new_n294__spl_;
  wire new_n294__spl_0;
  wire new_n329__spl_;
  wire new_n329__spl_0;
  wire new_n344__spl_;
  wire new_n344__spl_0;
  wire new_n359__spl_;
  wire new_n359__spl_0;
  wire new_n374__spl_;
  wire new_n374__spl_0;

  nor2
  g000
  (
    .dina(G6_spl_0),
    .dinb(G16_spl_),
    .dout(new_n87_)
  );


  nab2
  g001
  (
    .dina(G8_spl_00),
    .dinb(new_n87__spl_),
    .dout(G855)
  );


  nor2
  g002
  (
    .dina(G6_spl_0),
    .dinb(G7_spl_),
    .dout(new_n89_)
  );


  nab2
  g003
  (
    .dina(G17_spl_0),
    .dinb(new_n89__spl_),
    .dout(G856)
  );


  nab2
  g004
  (
    .dina(G8_spl_00),
    .dinb(new_n89__spl_),
    .dout(G857)
  );


  nor2
  g005
  (
    .dina(G18),
    .dinb(G19),
    .dout(G858)
  );


  nor2
  g006
  (
    .dina(G1_spl_0),
    .dinb(G2_spl_),
    .dout(new_n93_)
  );


  nab2
  g007
  (
    .dina(G3_spl_),
    .dinb(new_n93__spl_),
    .dout(new_n94_)
  );


  nab2
  g008
  (
    .dina(G4_spl_00),
    .dinb(new_n94__spl_),
    .dout(G859)
  );


  nor2
  g009
  (
    .dina(G1_spl_0),
    .dinb(G5),
    .dout(new_n96_)
  );


  and1
  g010
  (
    .dina(G3_spl_),
    .dinb(G4_spl_00),
    .dout(new_n97_)
  );


  anb2
  g011
  (
    .dina(new_n96__spl_),
    .dinb(new_n97_),
    .dout(new_n98_)
  );


  anb1
  g012
  (
    .dina(G857_spl_),
    .dinb(new_n98__spl_),
    .dout(G860)
  );


  nor2
  g013
  (
    .dina(G11_spl_0),
    .dinb(G16_spl_),
    .dout(new_n100_)
  );


  anb1
  g014
  (
    .dina(G17_spl_0),
    .dinb(new_n100__spl_),
    .dout(G861)
  );


  nor2
  g015
  (
    .dina(G7_spl_),
    .dinb(G11_spl_0),
    .dout(new_n102_)
  );


  anb1
  g016
  (
    .dina(G17_spl_1),
    .dinb(new_n102__spl_),
    .dout(G862)
  );


  anb1
  g017
  (
    .dina(G8_spl_01),
    .dinb(new_n102__spl_),
    .dout(G863)
  );


  nor1
  g018
  (
    .dina(G20),
    .dinb(G21),
    .dout(new_n105_)
  );


  anb2
  g019
  (
    .dina(new_n105__spl_),
    .dinb(G23),
    .dout(G864)
  );


  nor1
  g020
  (
    .dina(G857_spl_),
    .dinb(new_n98__spl_),
    .dout(G865)
  );


  nab2
  g021
  (
    .dina(G9_spl_0),
    .dinb(new_n96__spl_),
    .dout(G866)
  );


  nab2
  g022
  (
    .dina(G10_spl_0),
    .dinb(new_n94__spl_),
    .dout(new_n109_)
  );


  and1
  g023
  (
    .dina(G6_spl_),
    .dinb(G12_spl_),
    .dout(new_n110_)
  );


  anb2
  g024
  (
    .dina(new_n109__spl_0),
    .dinb(new_n110_),
    .dout(G867)
  );


  nor2
  g025
  (
    .dina(G11_spl_1),
    .dinb(G12_spl_),
    .dout(new_n112_)
  );


  anb1
  g026
  (
    .dina(G15),
    .dinb(new_n112__spl_),
    .dout(new_n113_)
  );


  anb2
  g027
  (
    .dina(new_n109__spl_0),
    .dinb(new_n113_),
    .dout(G868)
  );


  anb2
  g028
  (
    .dina(new_n105__spl_),
    .dinb(G22),
    .dout(G869)
  );


  nor1
  g029
  (
    .dina(G24_spl_0),
    .dinb(G25_spl_0),
    .dout(new_n116_)
  );


  nor2
  g030
  (
    .dina(G24_spl_0),
    .dinb(G25_spl_0),
    .dout(new_n117_)
  );


  anb2
  g031
  (
    .dina(new_n116_),
    .dinb(new_n117_),
    .dout(new_n118_)
  );


  and2
  g032
  (
    .dina(G26_spl_0),
    .dinb(G27_spl_0),
    .dout(new_n119_)
  );


  and1
  g033
  (
    .dina(G26_spl_0),
    .dinb(G27_spl_0),
    .dout(new_n120_)
  );


  anb1
  g034
  (
    .dina(new_n119_),
    .dinb(new_n120_),
    .dout(new_n121_)
  );


  anb1
  g035
  (
    .dina(new_n118__spl_),
    .dinb(new_n121__spl_),
    .dout(new_n122_)
  );


  anb2
  g036
  (
    .dina(new_n118__spl_),
    .dinb(new_n121__spl_),
    .dout(new_n123_)
  );


  anb2
  g037
  (
    .dina(new_n122_),
    .dinb(new_n123_),
    .dout(new_n124_)
  );


  anb1
  g038
  (
    .dina(G32_spl_0),
    .dinb(new_n124__spl_),
    .dout(new_n125_)
  );


  anb2
  g039
  (
    .dina(G32_spl_0),
    .dinb(new_n124__spl_),
    .dout(new_n126_)
  );


  anb2
  g040
  (
    .dina(new_n125_),
    .dinb(new_n126_),
    .dout(new_n127_)
  );


  nor1
  g041
  (
    .dina(G28_spl_0),
    .dinb(G29_spl_0),
    .dout(new_n128_)
  );


  nor2
  g042
  (
    .dina(G28_spl_0),
    .dinb(G29_spl_0),
    .dout(new_n129_)
  );


  anb2
  g043
  (
    .dina(new_n128_),
    .dinb(new_n129_),
    .dout(new_n130_)
  );


  and2
  g044
  (
    .dina(G30_spl_0),
    .dinb(G31_spl_0),
    .dout(new_n131_)
  );


  and1
  g045
  (
    .dina(G30_spl_0),
    .dinb(G31_spl_0),
    .dout(new_n132_)
  );


  anb1
  g046
  (
    .dina(new_n131_),
    .dinb(new_n132_),
    .dout(new_n133_)
  );


  anb1
  g047
  (
    .dina(new_n130__spl_),
    .dinb(new_n133__spl_),
    .dout(new_n134_)
  );


  anb2
  g048
  (
    .dina(new_n130__spl_),
    .dinb(new_n133__spl_),
    .dout(new_n135_)
  );


  anb2
  g049
  (
    .dina(new_n134_),
    .dinb(new_n135_),
    .dout(new_n136_)
  );


  nab2
  g050
  (
    .dina(G33_spl_),
    .dinb(new_n136__spl_),
    .dout(new_n137_)
  );


  nab1
  g051
  (
    .dina(G33_spl_),
    .dinb(new_n136__spl_),
    .dout(new_n138_)
  );


  anb1
  g052
  (
    .dina(new_n137_),
    .dinb(new_n138_),
    .dout(new_n139_)
  );


  anb1
  g053
  (
    .dina(new_n127__spl_),
    .dinb(new_n139__spl_),
    .dout(new_n140_)
  );


  anb2
  g054
  (
    .dina(new_n127__spl_),
    .dinb(new_n139__spl_),
    .dout(new_n141_)
  );


  anb2
  g055
  (
    .dina(new_n140_),
    .dinb(new_n141_),
    .dout(G870)
  );


  nor1
  g056
  (
    .dina(G41_spl_00),
    .dinb(G42_spl_00),
    .dout(new_n143_)
  );


  nor2
  g057
  (
    .dina(G41_spl_00),
    .dinb(G42_spl_00),
    .dout(new_n144_)
  );


  anb2
  g058
  (
    .dina(new_n143_),
    .dinb(new_n144_),
    .dout(new_n145_)
  );


  and2
  g059
  (
    .dina(G43_spl_00),
    .dinb(G44_spl_00),
    .dout(new_n146_)
  );


  and1
  g060
  (
    .dina(G43_spl_00),
    .dinb(G44_spl_00),
    .dout(new_n147_)
  );


  anb1
  g061
  (
    .dina(new_n146_),
    .dinb(new_n147_),
    .dout(new_n148_)
  );


  anb1
  g062
  (
    .dina(new_n145__spl_),
    .dinb(new_n148__spl_),
    .dout(new_n149_)
  );


  anb2
  g063
  (
    .dina(new_n145__spl_),
    .dinb(new_n148__spl_),
    .dout(new_n150_)
  );


  anb2
  g064
  (
    .dina(new_n149_),
    .dinb(new_n150_),
    .dout(new_n151_)
  );


  anb1
  g065
  (
    .dina(G32_spl_1),
    .dinb(new_n151__spl_),
    .dout(new_n152_)
  );


  anb2
  g066
  (
    .dina(G32_spl_1),
    .dinb(new_n151__spl_),
    .dout(new_n153_)
  );


  anb2
  g067
  (
    .dina(new_n152_),
    .dinb(new_n153_),
    .dout(new_n154_)
  );


  nor1
  g068
  (
    .dina(G45_spl_00),
    .dinb(G46_spl_00),
    .dout(new_n155_)
  );


  nor2
  g069
  (
    .dina(G45_spl_00),
    .dinb(G46_spl_00),
    .dout(new_n156_)
  );


  anb2
  g070
  (
    .dina(new_n155_),
    .dinb(new_n156_),
    .dout(new_n157_)
  );


  and2
  g071
  (
    .dina(G47_spl_00),
    .dinb(G48_spl_00),
    .dout(new_n158_)
  );


  and1
  g072
  (
    .dina(G47_spl_00),
    .dinb(G48_spl_00),
    .dout(new_n159_)
  );


  anb1
  g073
  (
    .dina(new_n158_),
    .dinb(new_n159_),
    .dout(new_n160_)
  );


  anb1
  g074
  (
    .dina(new_n157__spl_),
    .dinb(new_n160__spl_),
    .dout(new_n161_)
  );


  anb2
  g075
  (
    .dina(new_n157__spl_),
    .dinb(new_n160__spl_),
    .dout(new_n162_)
  );


  anb2
  g076
  (
    .dina(new_n161_),
    .dinb(new_n162_),
    .dout(new_n163_)
  );


  nab2
  g077
  (
    .dina(G49_spl_),
    .dinb(new_n163__spl_),
    .dout(new_n164_)
  );


  nab1
  g078
  (
    .dina(G49_spl_),
    .dinb(new_n163__spl_),
    .dout(new_n165_)
  );


  anb1
  g079
  (
    .dina(new_n164_),
    .dinb(new_n165_),
    .dout(new_n166_)
  );


  anb1
  g080
  (
    .dina(new_n154__spl_),
    .dinb(new_n166__spl_),
    .dout(new_n167_)
  );


  anb2
  g081
  (
    .dina(new_n154__spl_),
    .dinb(new_n166__spl_),
    .dout(new_n168_)
  );


  anb2
  g082
  (
    .dina(new_n167_),
    .dinb(new_n168_),
    .dout(G871)
  );


  nor2
  g083
  (
    .dina(G11_spl_1),
    .dinb(G40),
    .dout(new_n170_)
  );


  anb2
  g084
  (
    .dina(G866_spl_0),
    .dinb(new_n170__spl_),
    .dout(new_n171_)
  );


  anb1
  g085
  (
    .dina(G4_spl_01),
    .dinb(new_n171__spl_),
    .dout(new_n172_)
  );


  anb1
  g086
  (
    .dina(G1_spl_),
    .dinb(new_n172_),
    .dout(new_n173_)
  );


  anb1
  g087
  (
    .dina(G39_spl_),
    .dinb(new_n173__spl_0),
    .dout(new_n174_)
  );


  anb1
  g088
  (
    .dina(G17_spl_1),
    .dinb(new_n87__spl_),
    .dout(new_n175_)
  );


  anb2
  g089
  (
    .dina(G866_spl_0),
    .dinb(new_n175_),
    .dout(new_n176_)
  );


  anb1
  g090
  (
    .dina(G10_spl_0),
    .dinb(G60_spl_0),
    .dout(new_n177_)
  );


  anb2
  g091
  (
    .dina(new_n176__spl_),
    .dinb(new_n177_),
    .dout(new_n178_)
  );


  and2
  g092
  (
    .dina(G4_spl_01),
    .dinb(G8_spl_01),
    .dout(new_n179_)
  );


  and1
  g093
  (
    .dina(G4_spl_10),
    .dinb(G8_spl_10),
    .dout(new_n180_)
  );


  anb1
  g094
  (
    .dina(new_n179_),
    .dinb(new_n180_),
    .dout(new_n181_)
  );


  anb2
  g095
  (
    .dina(new_n170__spl_),
    .dinb(new_n181_),
    .dout(new_n182_)
  );


  and2
  g096
  (
    .dina(G866_spl_),
    .dinb(new_n182_),
    .dout(new_n183_)
  );


  nab2
  g097
  (
    .dina(G8_spl_10),
    .dinb(new_n100__spl_),
    .dout(new_n184_)
  );


  and1
  g098
  (
    .dina(G4_spl_10),
    .dinb(G9_spl_0),
    .dout(new_n185_)
  );


  anb2
  g099
  (
    .dina(new_n93__spl_),
    .dinb(new_n185_),
    .dout(new_n186_)
  );


  anb1
  g100
  (
    .dina(new_n184_),
    .dinb(new_n186_),
    .dout(new_n187_)
  );


  anb1
  g101
  (
    .dina(new_n183_),
    .dinb(new_n187_),
    .dout(new_n188_)
  );


  anb2
  g102
  (
    .dina(new_n188__spl_00),
    .dinb(G31_spl_),
    .dout(new_n189_)
  );


  anb2
  g103
  (
    .dina(new_n174_),
    .dinb(new_n189_),
    .dout(new_n190_)
  );


  anb1
  g104
  (
    .dina(new_n178__spl_0),
    .dinb(new_n190_),
    .dout(new_n191_)
  );


  anb2
  g105
  (
    .dina(new_n191__spl_0),
    .dinb(G48_spl_0),
    .dout(new_n192_)
  );


  nor1
  g106
  (
    .dina(G53_spl_00),
    .dinb(new_n192__spl_0),
    .dout(new_n193_)
  );


  anb1
  g107
  (
    .dina(new_n191__spl_0),
    .dinb(G48_spl_1),
    .dout(new_n194_)
  );


  and2
  g108
  (
    .dina(new_n193_),
    .dinb(new_n194__spl_),
    .dout(new_n195_)
  );


  and1
  g109
  (
    .dina(G51_spl_000),
    .dinb(G58_spl_),
    .dout(new_n196_)
  );


  anb1
  g110
  (
    .dina(new_n195_),
    .dinb(new_n196_),
    .dout(new_n197_)
  );


  anb1
  g111
  (
    .dina(G58_spl_),
    .dinb(new_n194__spl_),
    .dout(new_n198_)
  );


  anb1
  g112
  (
    .dina(G51_spl_000),
    .dinb(new_n198__spl_),
    .dout(new_n199_)
  );


  nab1
  g113
  (
    .dina(G52_spl_00),
    .dinb(new_n192__spl_0),
    .dout(new_n200_)
  );


  anb2
  g114
  (
    .dina(new_n199_),
    .dinb(new_n200_),
    .dout(new_n201_)
  );


  anb2
  g115
  (
    .dina(new_n197_),
    .dinb(new_n201_),
    .dout(new_n202_)
  );


  anb1
  g116
  (
    .dina(G54_spl_00),
    .dinb(new_n191__spl_),
    .dout(new_n203_)
  );


  nor2
  g117
  (
    .dina(G8_spl_1),
    .dinb(G13),
    .dout(new_n204_)
  );


  anb1
  g118
  (
    .dina(G14),
    .dinb(new_n204_),
    .dout(new_n205_)
  );


  nab1
  g119
  (
    .dina(new_n112__spl_),
    .dinb(new_n205_),
    .dout(new_n206_)
  );


  anb2
  g120
  (
    .dina(new_n109__spl_),
    .dinb(new_n206_),
    .dout(new_n207_)
  );


  nab2
  g121
  (
    .dina(G48_spl_1),
    .dinb(new_n207__spl_00),
    .dout(new_n208_)
  );


  and1
  g122
  (
    .dina(G55_spl_0),
    .dinb(G59),
    .dout(new_n209_)
  );


  nor2
  g123
  (
    .dina(G30_spl_1),
    .dinb(G50_spl_00),
    .dout(new_n210_)
  );


  anb2
  g124
  (
    .dina(new_n209_),
    .dinb(new_n210_),
    .dout(new_n211_)
  );


  anb1
  g125
  (
    .dina(new_n208_),
    .dinb(new_n211_),
    .dout(new_n212_)
  );


  anb2
  g126
  (
    .dina(new_n203_),
    .dinb(new_n212_),
    .dout(new_n213_)
  );


  anb1
  g127
  (
    .dina(new_n202_),
    .dinb(new_n213_),
    .dout(G872)
  );


  anb1
  g128
  (
    .dina(G36_spl_),
    .dinb(new_n173__spl_0),
    .dout(new_n215_)
  );


  anb2
  g129
  (
    .dina(new_n188__spl_00),
    .dinb(G29_spl_1),
    .dout(new_n216_)
  );


  anb2
  g130
  (
    .dina(new_n215_),
    .dinb(new_n216_),
    .dout(new_n217_)
  );


  anb1
  g131
  (
    .dina(new_n178__spl_0),
    .dinb(new_n217_),
    .dout(new_n218_)
  );


  anb2
  g132
  (
    .dina(new_n218__spl_0),
    .dinb(G46_spl_0),
    .dout(new_n219_)
  );


  anb2
  g133
  (
    .dina(G46_spl_1),
    .dinb(new_n218__spl_0),
    .dout(new_n220_)
  );


  anb1
  g134
  (
    .dina(G37_spl_),
    .dinb(new_n173__spl_1),
    .dout(new_n221_)
  );


  anb2
  g135
  (
    .dina(new_n188__spl_01),
    .dinb(G30_spl_1),
    .dout(new_n222_)
  );


  anb2
  g136
  (
    .dina(new_n221_),
    .dinb(new_n222_),
    .dout(new_n223_)
  );


  anb1
  g137
  (
    .dina(new_n178__spl_1),
    .dinb(new_n223_),
    .dout(new_n224_)
  );


  anb2
  g138
  (
    .dina(new_n224__spl_0),
    .dinb(G47_spl_0),
    .dout(new_n225_)
  );


  anb2
  g139
  (
    .dina(G47_spl_1),
    .dinb(new_n224__spl_0),
    .dout(new_n226_)
  );


  anb1
  g140
  (
    .dina(new_n192__spl_),
    .dinb(new_n198__spl_),
    .dout(new_n227_)
  );


  anb1
  g141
  (
    .dina(new_n226__spl_),
    .dinb(new_n227__spl_),
    .dout(new_n228_)
  );


  anb1
  g142
  (
    .dina(new_n225__spl_0),
    .dinb(new_n228__spl_),
    .dout(new_n229_)
  );


  anb1
  g143
  (
    .dina(new_n220__spl_),
    .dinb(new_n229__spl_),
    .dout(new_n230_)
  );


  anb1
  g144
  (
    .dina(new_n219__spl_0),
    .dinb(new_n230__spl_),
    .dout(new_n231_)
  );


  anb2
  g145
  (
    .dina(new_n231__spl_),
    .dinb(G51_spl_001),
    .dout(new_n232_)
  );


  anb1
  g146
  (
    .dina(G35_spl_),
    .dinb(new_n173__spl_1),
    .dout(new_n233_)
  );


  anb2
  g147
  (
    .dina(new_n188__spl_01),
    .dinb(G28_spl_1),
    .dout(new_n234_)
  );


  anb2
  g148
  (
    .dina(new_n233_),
    .dinb(new_n234_),
    .dout(new_n235_)
  );


  anb1
  g149
  (
    .dina(new_n178__spl_1),
    .dinb(new_n235_),
    .dout(new_n236_)
  );


  anb1
  g150
  (
    .dina(G45_spl_0),
    .dinb(new_n236__spl_0),
    .dout(new_n237_)
  );


  anb2
  g151
  (
    .dina(G53_spl_00),
    .dinb(new_n237__spl_0),
    .dout(new_n238_)
  );


  anb1
  g152
  (
    .dina(new_n236__spl_0),
    .dinb(G45_spl_1),
    .dout(new_n239_)
  );


  anb1
  g153
  (
    .dina(new_n238_),
    .dinb(new_n239__spl_),
    .dout(new_n240_)
  );


  anb1
  g154
  (
    .dina(new_n232_),
    .dinb(new_n240_),
    .dout(new_n241_)
  );


  nor1
  g155
  (
    .dina(new_n231__spl_),
    .dinb(new_n239__spl_),
    .dout(new_n242_)
  );


  anb1
  g156
  (
    .dina(G51_spl_001),
    .dinb(new_n242__spl_),
    .dout(new_n243_)
  );


  nor1
  g157
  (
    .dina(G52_spl_00),
    .dinb(new_n237__spl_0),
    .dout(new_n244_)
  );


  anb2
  g158
  (
    .dina(new_n243_),
    .dinb(new_n244_),
    .dout(new_n245_)
  );


  anb2
  g159
  (
    .dina(new_n241_),
    .dinb(new_n245_),
    .dout(new_n246_)
  );


  anb1
  g160
  (
    .dina(G54_spl_00),
    .dinb(new_n236__spl_),
    .dout(new_n247_)
  );


  nor2
  g161
  (
    .dina(G27_spl_1),
    .dinb(G50_spl_00),
    .dout(new_n248_)
  );


  anb1
  g162
  (
    .dina(G45_spl_1),
    .dinb(new_n207__spl_00),
    .dout(new_n249_)
  );


  anb1
  g163
  (
    .dina(new_n248_),
    .dinb(new_n249_),
    .dout(new_n250_)
  );


  anb2
  g164
  (
    .dina(new_n247_),
    .dinb(new_n250_),
    .dout(new_n251_)
  );


  anb1
  g165
  (
    .dina(new_n246_),
    .dinb(new_n251_),
    .dout(G873)
  );


  nor1
  g166
  (
    .dina(G53_spl_01),
    .dinb(new_n219__spl_0),
    .dout(new_n253_)
  );


  nab2
  g167
  (
    .dina(new_n220__spl_),
    .dinb(new_n253_),
    .dout(new_n254_)
  );


  anb1
  g168
  (
    .dina(G51_spl_010),
    .dinb(new_n229__spl_),
    .dout(new_n255_)
  );


  anb1
  g169
  (
    .dina(new_n254_),
    .dinb(new_n255_),
    .dout(new_n256_)
  );


  anb1
  g170
  (
    .dina(G51_spl_010),
    .dinb(new_n230__spl_),
    .dout(new_n257_)
  );


  nab1
  g171
  (
    .dina(G52_spl_01),
    .dinb(new_n219__spl_),
    .dout(new_n258_)
  );


  anb2
  g172
  (
    .dina(new_n257_),
    .dinb(new_n258_),
    .dout(new_n259_)
  );


  anb2
  g173
  (
    .dina(new_n256_),
    .dinb(new_n259_),
    .dout(new_n260_)
  );


  anb1
  g174
  (
    .dina(G54_spl_01),
    .dinb(new_n218__spl_),
    .dout(new_n261_)
  );


  nab2
  g175
  (
    .dina(G46_spl_1),
    .dinb(new_n207__spl_01),
    .dout(new_n262_)
  );


  and1
  g176
  (
    .dina(G55_spl_0),
    .dinb(G56),
    .dout(new_n263_)
  );


  nor2
  g177
  (
    .dina(G28_spl_1),
    .dinb(G50_spl_01),
    .dout(new_n264_)
  );


  anb2
  g178
  (
    .dina(new_n263_),
    .dinb(new_n264_),
    .dout(new_n265_)
  );


  anb1
  g179
  (
    .dina(new_n262_),
    .dinb(new_n265_),
    .dout(new_n266_)
  );


  anb2
  g180
  (
    .dina(new_n261_),
    .dinb(new_n266_),
    .dout(new_n267_)
  );


  anb1
  g181
  (
    .dina(new_n260_),
    .dinb(new_n267_),
    .dout(G874)
  );


  nor1
  g182
  (
    .dina(G53_spl_01),
    .dinb(new_n225__spl_0),
    .dout(new_n269_)
  );


  nab2
  g183
  (
    .dina(new_n226__spl_),
    .dinb(new_n269_),
    .dout(new_n270_)
  );


  anb1
  g184
  (
    .dina(G51_spl_011),
    .dinb(new_n227__spl_),
    .dout(new_n271_)
  );


  anb1
  g185
  (
    .dina(new_n270_),
    .dinb(new_n271_),
    .dout(new_n272_)
  );


  anb1
  g186
  (
    .dina(G51_spl_011),
    .dinb(new_n228__spl_),
    .dout(new_n273_)
  );


  nab1
  g187
  (
    .dina(G52_spl_01),
    .dinb(new_n225__spl_),
    .dout(new_n274_)
  );


  anb2
  g188
  (
    .dina(new_n273_),
    .dinb(new_n274_),
    .dout(new_n275_)
  );


  anb2
  g189
  (
    .dina(new_n272_),
    .dinb(new_n275_),
    .dout(new_n276_)
  );


  anb1
  g190
  (
    .dina(G54_spl_01),
    .dinb(new_n224__spl_),
    .dout(new_n277_)
  );


  nab2
  g191
  (
    .dina(G47_spl_1),
    .dinb(new_n207__spl_01),
    .dout(new_n278_)
  );


  and1
  g192
  (
    .dina(G55_spl_),
    .dinb(G57),
    .dout(new_n279_)
  );


  nor2
  g193
  (
    .dina(G29_spl_1),
    .dinb(G50_spl_01),
    .dout(new_n280_)
  );


  anb2
  g194
  (
    .dina(new_n279_),
    .dinb(new_n280_),
    .dout(new_n281_)
  );


  anb1
  g195
  (
    .dina(new_n278_),
    .dinb(new_n281_),
    .dout(new_n282_)
  );


  anb2
  g196
  (
    .dina(new_n277_),
    .dinb(new_n282_),
    .dout(new_n283_)
  );


  anb1
  g197
  (
    .dina(new_n276_),
    .dinb(new_n283_),
    .dout(G875)
  );


  anb2
  g198
  (
    .dina(new_n188__spl_10),
    .dinb(G24_spl_1),
    .dout(new_n285_)
  );


  nab2
  g199
  (
    .dina(G10_spl_),
    .dinb(new_n171__spl_),
    .dout(new_n286_)
  );


  anb1
  g200
  (
    .dina(G35_spl_),
    .dinb(new_n286__spl_0),
    .dout(new_n287_)
  );


  nor2
  g201
  (
    .dina(G2_spl_),
    .dinb(G34_spl_0),
    .dout(new_n288_)
  );


  anb1
  g202
  (
    .dina(G4_spl_11),
    .dinb(G60_spl_0),
    .dout(new_n289_)
  );


  anb2
  g203
  (
    .dina(new_n176__spl_),
    .dinb(new_n289_),
    .dout(new_n290_)
  );


  and1
  g204
  (
    .dina(new_n288_),
    .dinb(new_n290__spl_0),
    .dout(new_n291_)
  );


  anb2
  g205
  (
    .dina(new_n287_),
    .dinb(new_n291_),
    .dout(new_n292_)
  );


  anb1
  g206
  (
    .dina(new_n285_),
    .dinb(new_n292_),
    .dout(new_n293_)
  );


  anb2
  g207
  (
    .dina(new_n293__spl_0),
    .dinb(G41_spl_0),
    .dout(new_n294_)
  );


  anb2
  g208
  (
    .dina(new_n188__spl_10),
    .dinb(G25_spl_1),
    .dout(new_n295_)
  );


  anb1
  g209
  (
    .dina(G36_spl_),
    .dinb(new_n286__spl_0),
    .dout(new_n296_)
  );


  and1
  g210
  (
    .dina(G9_spl_),
    .dinb(G34_spl_0),
    .dout(new_n297_)
  );


  anb1
  g211
  (
    .dina(new_n290__spl_0),
    .dinb(new_n297_),
    .dout(new_n298_)
  );


  anb2
  g212
  (
    .dina(new_n296_),
    .dinb(new_n298_),
    .dout(new_n299_)
  );


  anb1
  g213
  (
    .dina(new_n295_),
    .dinb(new_n299_),
    .dout(new_n300_)
  );


  anb2
  g214
  (
    .dina(new_n300__spl_0),
    .dinb(G42_spl_0),
    .dout(new_n301_)
  );


  anb2
  g215
  (
    .dina(G42_spl_1),
    .dinb(new_n300__spl_0),
    .dout(new_n302_)
  );


  anb2
  g216
  (
    .dina(new_n188__spl_11),
    .dinb(G26_spl_1),
    .dout(new_n303_)
  );


  anb1
  g217
  (
    .dina(G37_spl_),
    .dinb(new_n286__spl_1),
    .dout(new_n304_)
  );


  and1
  g218
  (
    .dina(G4_spl_11),
    .dinb(G34_spl_1),
    .dout(new_n305_)
  );


  anb1
  g219
  (
    .dina(new_n290__spl_1),
    .dinb(new_n305_),
    .dout(new_n306_)
  );


  anb2
  g220
  (
    .dina(new_n304_),
    .dinb(new_n306_),
    .dout(new_n307_)
  );


  anb1
  g221
  (
    .dina(new_n303_),
    .dinb(new_n307_),
    .dout(new_n308_)
  );


  anb2
  g222
  (
    .dina(new_n308__spl_0),
    .dinb(G43_spl_0),
    .dout(new_n309_)
  );


  anb2
  g223
  (
    .dina(G43_spl_1),
    .dinb(new_n308__spl_0),
    .dout(new_n310_)
  );


  nor1
  g224
  (
    .dina(new_n237__spl_),
    .dinb(new_n242__spl_),
    .dout(new_n311_)
  );


  anb2
  g225
  (
    .dina(new_n188__spl_11),
    .dinb(G27_spl_1),
    .dout(new_n312_)
  );


  anb1
  g226
  (
    .dina(G39_spl_),
    .dinb(new_n286__spl_1),
    .dout(new_n313_)
  );


  and1
  g227
  (
    .dina(G34_spl_1),
    .dinb(G38),
    .dout(new_n314_)
  );


  anb1
  g228
  (
    .dina(new_n290__spl_1),
    .dinb(new_n314_),
    .dout(new_n315_)
  );


  anb2
  g229
  (
    .dina(new_n313_),
    .dinb(new_n315_),
    .dout(new_n316_)
  );


  anb1
  g230
  (
    .dina(new_n312_),
    .dinb(new_n316_),
    .dout(new_n317_)
  );


  anb1
  g231
  (
    .dina(new_n317__spl_0),
    .dinb(G44_spl_0),
    .dout(new_n318_)
  );


  nor1
  g232
  (
    .dina(new_n311__spl_0),
    .dinb(new_n318__spl_),
    .dout(new_n319_)
  );


  anb2
  g233
  (
    .dina(new_n317__spl_0),
    .dinb(G44_spl_1),
    .dout(new_n320_)
  );


  anb2
  g234
  (
    .dina(new_n319_),
    .dinb(new_n320__spl_0),
    .dout(new_n321_)
  );


  and1
  g235
  (
    .dina(new_n310__spl_),
    .dinb(new_n321__spl_0),
    .dout(new_n322_)
  );


  nab2
  g236
  (
    .dina(new_n309__spl_0),
    .dinb(new_n322_),
    .dout(new_n323_)
  );


  and1
  g237
  (
    .dina(new_n302__spl_),
    .dinb(new_n323__spl_0),
    .dout(new_n324_)
  );


  nab2
  g238
  (
    .dina(new_n301__spl_0),
    .dinb(new_n324_),
    .dout(new_n325_)
  );


  anb1
  g239
  (
    .dina(new_n293__spl_0),
    .dinb(G41_spl_1),
    .dout(new_n326_)
  );


  anb1
  g240
  (
    .dina(new_n325__spl_0),
    .dinb(new_n326__spl_),
    .dout(new_n327_)
  );


  anb1
  g241
  (
    .dina(new_n294__spl_0),
    .dinb(new_n327_),
    .dout(G876)
  );


  anb2
  g242
  (
    .dina(new_n318__spl_),
    .dinb(new_n320__spl_0),
    .dout(new_n329_)
  );


  anb2
  g243
  (
    .dina(new_n311__spl_0),
    .dinb(new_n329__spl_0),
    .dout(new_n330_)
  );


  anb1
  g244
  (
    .dina(new_n311__spl_),
    .dinb(new_n329__spl_0),
    .dout(new_n331_)
  );


  anb1
  g245
  (
    .dina(new_n330_),
    .dinb(new_n331_),
    .dout(new_n332_)
  );


  anb2
  g246
  (
    .dina(new_n332_),
    .dinb(G51_spl_10),
    .dout(new_n333_)
  );


  anb1
  g247
  (
    .dina(G52_spl_10),
    .dinb(new_n329__spl_),
    .dout(new_n334_)
  );


  nab2
  g248
  (
    .dina(G53_spl_10),
    .dinb(new_n320__spl_),
    .dout(new_n335_)
  );


  anb1
  g249
  (
    .dina(G54_spl_10),
    .dinb(new_n317__spl_),
    .dout(new_n336_)
  );


  nor2
  g250
  (
    .dina(G26_spl_1),
    .dinb(G50_spl_10),
    .dout(new_n337_)
  );


  anb1
  g251
  (
    .dina(G44_spl_1),
    .dinb(new_n207__spl_10),
    .dout(new_n338_)
  );


  anb1
  g252
  (
    .dina(new_n337_),
    .dinb(new_n338_),
    .dout(new_n339_)
  );


  anb2
  g253
  (
    .dina(new_n336_),
    .dinb(new_n339_),
    .dout(new_n340_)
  );


  anb1
  g254
  (
    .dina(new_n335_),
    .dinb(new_n340_),
    .dout(new_n341_)
  );


  anb2
  g255
  (
    .dina(new_n334_),
    .dinb(new_n341_),
    .dout(new_n342_)
  );


  anb1
  g256
  (
    .dina(new_n333_),
    .dinb(new_n342_),
    .dout(G877)
  );


  nab2
  g257
  (
    .dina(new_n294__spl_0),
    .dinb(new_n326__spl_),
    .dout(new_n344_)
  );


  anb1
  g258
  (
    .dina(new_n325__spl_0),
    .dinb(new_n344__spl_0),
    .dout(new_n345_)
  );


  anb1
  g259
  (
    .dina(new_n344__spl_0),
    .dinb(new_n325__spl_),
    .dout(new_n346_)
  );


  anb1
  g260
  (
    .dina(G51_spl_10),
    .dinb(new_n346_),
    .dout(new_n347_)
  );


  anb2
  g261
  (
    .dina(new_n345_),
    .dinb(new_n347_),
    .dout(new_n348_)
  );


  anb1
  g262
  (
    .dina(G52_spl_10),
    .dinb(new_n344__spl_),
    .dout(new_n349_)
  );


  nab2
  g263
  (
    .dina(G53_spl_10),
    .dinb(new_n294__spl_),
    .dout(new_n350_)
  );


  anb1
  g264
  (
    .dina(G54_spl_10),
    .dinb(new_n293__spl_),
    .dout(new_n351_)
  );


  nor2
  g265
  (
    .dina(G50_spl_10),
    .dinb(G60_spl_),
    .dout(new_n352_)
  );


  anb1
  g266
  (
    .dina(G41_spl_1),
    .dinb(new_n207__spl_10),
    .dout(new_n353_)
  );


  anb1
  g267
  (
    .dina(new_n352_),
    .dinb(new_n353_),
    .dout(new_n354_)
  );


  anb2
  g268
  (
    .dina(new_n351_),
    .dinb(new_n354_),
    .dout(new_n355_)
  );


  anb1
  g269
  (
    .dina(new_n350_),
    .dinb(new_n355_),
    .dout(new_n356_)
  );


  anb2
  g270
  (
    .dina(new_n349_),
    .dinb(new_n356_),
    .dout(new_n357_)
  );


  anb1
  g271
  (
    .dina(new_n348_),
    .dinb(new_n357_),
    .dout(G878)
  );


  nor2
  g272
  (
    .dina(new_n301__spl_0),
    .dinb(new_n302__spl_),
    .dout(new_n359_)
  );


  anb1
  g273
  (
    .dina(new_n323__spl_0),
    .dinb(new_n359__spl_0),
    .dout(new_n360_)
  );


  anb1
  g274
  (
    .dina(new_n359__spl_0),
    .dinb(new_n323__spl_),
    .dout(new_n361_)
  );


  anb1
  g275
  (
    .dina(G51_spl_11),
    .dinb(new_n361_),
    .dout(new_n362_)
  );


  anb2
  g276
  (
    .dina(new_n360_),
    .dinb(new_n362_),
    .dout(new_n363_)
  );


  anb1
  g277
  (
    .dina(G52_spl_11),
    .dinb(new_n359__spl_),
    .dout(new_n364_)
  );


  nab2
  g278
  (
    .dina(G53_spl_11),
    .dinb(new_n301__spl_),
    .dout(new_n365_)
  );


  anb1
  g279
  (
    .dina(G54_spl_11),
    .dinb(new_n300__spl_),
    .dout(new_n366_)
  );


  nor2
  g280
  (
    .dina(G24_spl_1),
    .dinb(G50_spl_11),
    .dout(new_n367_)
  );


  anb1
  g281
  (
    .dina(G42_spl_1),
    .dinb(new_n207__spl_11),
    .dout(new_n368_)
  );


  anb1
  g282
  (
    .dina(new_n367_),
    .dinb(new_n368_),
    .dout(new_n369_)
  );


  anb2
  g283
  (
    .dina(new_n366_),
    .dinb(new_n369_),
    .dout(new_n370_)
  );


  anb1
  g284
  (
    .dina(new_n365_),
    .dinb(new_n370_),
    .dout(new_n371_)
  );


  anb2
  g285
  (
    .dina(new_n364_),
    .dinb(new_n371_),
    .dout(new_n372_)
  );


  anb1
  g286
  (
    .dina(new_n363_),
    .dinb(new_n372_),
    .dout(G879)
  );


  nor2
  g287
  (
    .dina(new_n309__spl_0),
    .dinb(new_n310__spl_),
    .dout(new_n374_)
  );


  anb1
  g288
  (
    .dina(new_n321__spl_0),
    .dinb(new_n374__spl_0),
    .dout(new_n375_)
  );


  anb1
  g289
  (
    .dina(new_n374__spl_0),
    .dinb(new_n321__spl_),
    .dout(new_n376_)
  );


  anb1
  g290
  (
    .dina(G51_spl_11),
    .dinb(new_n376_),
    .dout(new_n377_)
  );


  anb2
  g291
  (
    .dina(new_n375_),
    .dinb(new_n377_),
    .dout(new_n378_)
  );


  anb1
  g292
  (
    .dina(G52_spl_11),
    .dinb(new_n374__spl_),
    .dout(new_n379_)
  );


  nab2
  g293
  (
    .dina(G53_spl_11),
    .dinb(new_n309__spl_),
    .dout(new_n380_)
  );


  anb1
  g294
  (
    .dina(G54_spl_11),
    .dinb(new_n308__spl_),
    .dout(new_n381_)
  );


  nor2
  g295
  (
    .dina(G25_spl_1),
    .dinb(G50_spl_11),
    .dout(new_n382_)
  );


  anb1
  g296
  (
    .dina(G43_spl_1),
    .dinb(new_n207__spl_11),
    .dout(new_n383_)
  );


  anb1
  g297
  (
    .dina(new_n382_),
    .dinb(new_n383_),
    .dout(new_n384_)
  );


  anb2
  g298
  (
    .dina(new_n381_),
    .dinb(new_n384_),
    .dout(new_n385_)
  );


  anb1
  g299
  (
    .dina(new_n380_),
    .dinb(new_n385_),
    .dout(new_n386_)
  );


  anb2
  g300
  (
    .dina(new_n379_),
    .dinb(new_n386_),
    .dout(new_n387_)
  );


  anb1
  g301
  (
    .dina(new_n378_),
    .dinb(new_n387_),
    .dout(G880)
  );


  splt
  gG6
  (
    .dout(G6_spl_),
    .din(G6)
  );


  splt
  gG6_spl_
  (
    .dout(G6_spl_0),
    .din(G6_spl_)
  );


  splt
  gG16
  (
    .dout(G16_spl_),
    .din(G16)
  );


  splt
  gG8
  (
    .dout(G8_spl_),
    .din(G8)
  );


  splt
  gG8_spl_
  (
    .dout(G8_spl_0),
    .din(G8_spl_)
  );


  splt
  gG8_spl_0
  (
    .dout(G8_spl_00),
    .din(G8_spl_0)
  );


  splt
  gG8_spl_0
  (
    .dout(G8_spl_01),
    .din(G8_spl_0)
  );


  splt
  gG8_spl_
  (
    .dout(G8_spl_1),
    .din(G8_spl_)
  );


  splt
  gG8_spl_1
  (
    .dout(G8_spl_10),
    .din(G8_spl_1)
  );


  splt
  gnew_n87_
  (
    .dout(new_n87__spl_),
    .din(new_n87_)
  );


  splt
  gG7
  (
    .dout(G7_spl_),
    .din(G7)
  );


  splt
  gG17
  (
    .dout(G17_spl_),
    .din(G17)
  );


  splt
  gG17_spl_
  (
    .dout(G17_spl_0),
    .din(G17_spl_)
  );


  splt
  gG17_spl_
  (
    .dout(G17_spl_1),
    .din(G17_spl_)
  );


  splt
  gnew_n89_
  (
    .dout(new_n89__spl_),
    .din(new_n89_)
  );


  splt
  gG1
  (
    .dout(G1_spl_),
    .din(G1)
  );


  splt
  gG1_spl_
  (
    .dout(G1_spl_0),
    .din(G1_spl_)
  );


  splt
  gG2
  (
    .dout(G2_spl_),
    .din(G2)
  );


  splt
  gG3
  (
    .dout(G3_spl_),
    .din(G3)
  );


  splt
  gnew_n93_
  (
    .dout(new_n93__spl_),
    .din(new_n93_)
  );


  splt
  gG4
  (
    .dout(G4_spl_),
    .din(G4)
  );


  splt
  gG4_spl_
  (
    .dout(G4_spl_0),
    .din(G4_spl_)
  );


  splt
  gG4_spl_0
  (
    .dout(G4_spl_00),
    .din(G4_spl_0)
  );


  splt
  gG4_spl_0
  (
    .dout(G4_spl_01),
    .din(G4_spl_0)
  );


  splt
  gG4_spl_
  (
    .dout(G4_spl_1),
    .din(G4_spl_)
  );


  splt
  gG4_spl_1
  (
    .dout(G4_spl_10),
    .din(G4_spl_1)
  );


  splt
  gG4_spl_1
  (
    .dout(G4_spl_11),
    .din(G4_spl_1)
  );


  splt
  gnew_n94_
  (
    .dout(new_n94__spl_),
    .din(new_n94_)
  );


  splt
  gnew_n96_
  (
    .dout(new_n96__spl_),
    .din(new_n96_)
  );


  splt
  gG857
  (
    .dout(G857_spl_),
    .din(G857)
  );


  splt
  gnew_n98_
  (
    .dout(new_n98__spl_),
    .din(new_n98_)
  );


  splt
  gG11
  (
    .dout(G11_spl_),
    .din(G11)
  );


  splt
  gG11_spl_
  (
    .dout(G11_spl_0),
    .din(G11_spl_)
  );


  splt
  gG11_spl_
  (
    .dout(G11_spl_1),
    .din(G11_spl_)
  );


  splt
  gnew_n100_
  (
    .dout(new_n100__spl_),
    .din(new_n100_)
  );


  splt
  gnew_n102_
  (
    .dout(new_n102__spl_),
    .din(new_n102_)
  );


  splt
  gnew_n105_
  (
    .dout(new_n105__spl_),
    .din(new_n105_)
  );


  splt
  gG9
  (
    .dout(G9_spl_),
    .din(G9)
  );


  splt
  gG9_spl_
  (
    .dout(G9_spl_0),
    .din(G9_spl_)
  );


  splt
  gG10
  (
    .dout(G10_spl_),
    .din(G10)
  );


  splt
  gG10_spl_
  (
    .dout(G10_spl_0),
    .din(G10_spl_)
  );


  splt
  gG12
  (
    .dout(G12_spl_),
    .din(G12)
  );


  splt
  gnew_n109_
  (
    .dout(new_n109__spl_),
    .din(new_n109_)
  );


  splt
  gnew_n109__spl_
  (
    .dout(new_n109__spl_0),
    .din(new_n109__spl_)
  );


  splt
  gnew_n112_
  (
    .dout(new_n112__spl_),
    .din(new_n112_)
  );


  splt
  gG24
  (
    .dout(G24_spl_),
    .din(G24)
  );


  splt
  gG24_spl_
  (
    .dout(G24_spl_0),
    .din(G24_spl_)
  );


  splt
  gG24_spl_
  (
    .dout(G24_spl_1),
    .din(G24_spl_)
  );


  splt
  gG25
  (
    .dout(G25_spl_),
    .din(G25)
  );


  splt
  gG25_spl_
  (
    .dout(G25_spl_0),
    .din(G25_spl_)
  );


  splt
  gG25_spl_
  (
    .dout(G25_spl_1),
    .din(G25_spl_)
  );


  splt
  gG26
  (
    .dout(G26_spl_),
    .din(G26)
  );


  splt
  gG26_spl_
  (
    .dout(G26_spl_0),
    .din(G26_spl_)
  );


  splt
  gG26_spl_
  (
    .dout(G26_spl_1),
    .din(G26_spl_)
  );


  splt
  gG27
  (
    .dout(G27_spl_),
    .din(G27)
  );


  splt
  gG27_spl_
  (
    .dout(G27_spl_0),
    .din(G27_spl_)
  );


  splt
  gG27_spl_
  (
    .dout(G27_spl_1),
    .din(G27_spl_)
  );


  splt
  gnew_n118_
  (
    .dout(new_n118__spl_),
    .din(new_n118_)
  );


  splt
  gnew_n121_
  (
    .dout(new_n121__spl_),
    .din(new_n121_)
  );


  splt
  gG32
  (
    .dout(G32_spl_),
    .din(G32)
  );


  splt
  gG32_spl_
  (
    .dout(G32_spl_0),
    .din(G32_spl_)
  );


  splt
  gG32_spl_
  (
    .dout(G32_spl_1),
    .din(G32_spl_)
  );


  splt
  gnew_n124_
  (
    .dout(new_n124__spl_),
    .din(new_n124_)
  );


  splt
  gG28
  (
    .dout(G28_spl_),
    .din(G28)
  );


  splt
  gG28_spl_
  (
    .dout(G28_spl_0),
    .din(G28_spl_)
  );


  splt
  gG28_spl_
  (
    .dout(G28_spl_1),
    .din(G28_spl_)
  );


  splt
  gG29
  (
    .dout(G29_spl_),
    .din(G29)
  );


  splt
  gG29_spl_
  (
    .dout(G29_spl_0),
    .din(G29_spl_)
  );


  splt
  gG29_spl_
  (
    .dout(G29_spl_1),
    .din(G29_spl_)
  );


  splt
  gG30
  (
    .dout(G30_spl_),
    .din(G30)
  );


  splt
  gG30_spl_
  (
    .dout(G30_spl_0),
    .din(G30_spl_)
  );


  splt
  gG30_spl_
  (
    .dout(G30_spl_1),
    .din(G30_spl_)
  );


  splt
  gG31
  (
    .dout(G31_spl_),
    .din(G31)
  );


  splt
  gG31_spl_
  (
    .dout(G31_spl_0),
    .din(G31_spl_)
  );


  splt
  gnew_n130_
  (
    .dout(new_n130__spl_),
    .din(new_n130_)
  );


  splt
  gnew_n133_
  (
    .dout(new_n133__spl_),
    .din(new_n133_)
  );


  splt
  gG33
  (
    .dout(G33_spl_),
    .din(G33)
  );


  splt
  gnew_n136_
  (
    .dout(new_n136__spl_),
    .din(new_n136_)
  );


  splt
  gnew_n127_
  (
    .dout(new_n127__spl_),
    .din(new_n127_)
  );


  splt
  gnew_n139_
  (
    .dout(new_n139__spl_),
    .din(new_n139_)
  );


  splt
  gG41
  (
    .dout(G41_spl_),
    .din(G41)
  );


  splt
  gG41_spl_
  (
    .dout(G41_spl_0),
    .din(G41_spl_)
  );


  splt
  gG41_spl_0
  (
    .dout(G41_spl_00),
    .din(G41_spl_0)
  );


  splt
  gG41_spl_
  (
    .dout(G41_spl_1),
    .din(G41_spl_)
  );


  splt
  gG42
  (
    .dout(G42_spl_),
    .din(G42)
  );


  splt
  gG42_spl_
  (
    .dout(G42_spl_0),
    .din(G42_spl_)
  );


  splt
  gG42_spl_0
  (
    .dout(G42_spl_00),
    .din(G42_spl_0)
  );


  splt
  gG42_spl_
  (
    .dout(G42_spl_1),
    .din(G42_spl_)
  );


  splt
  gG43
  (
    .dout(G43_spl_),
    .din(G43)
  );


  splt
  gG43_spl_
  (
    .dout(G43_spl_0),
    .din(G43_spl_)
  );


  splt
  gG43_spl_0
  (
    .dout(G43_spl_00),
    .din(G43_spl_0)
  );


  splt
  gG43_spl_
  (
    .dout(G43_spl_1),
    .din(G43_spl_)
  );


  splt
  gG44
  (
    .dout(G44_spl_),
    .din(G44)
  );


  splt
  gG44_spl_
  (
    .dout(G44_spl_0),
    .din(G44_spl_)
  );


  splt
  gG44_spl_0
  (
    .dout(G44_spl_00),
    .din(G44_spl_0)
  );


  splt
  gG44_spl_
  (
    .dout(G44_spl_1),
    .din(G44_spl_)
  );


  splt
  gnew_n145_
  (
    .dout(new_n145__spl_),
    .din(new_n145_)
  );


  splt
  gnew_n148_
  (
    .dout(new_n148__spl_),
    .din(new_n148_)
  );


  splt
  gnew_n151_
  (
    .dout(new_n151__spl_),
    .din(new_n151_)
  );


  splt
  gG45
  (
    .dout(G45_spl_),
    .din(G45)
  );


  splt
  gG45_spl_
  (
    .dout(G45_spl_0),
    .din(G45_spl_)
  );


  splt
  gG45_spl_0
  (
    .dout(G45_spl_00),
    .din(G45_spl_0)
  );


  splt
  gG45_spl_
  (
    .dout(G45_spl_1),
    .din(G45_spl_)
  );


  splt
  gG46
  (
    .dout(G46_spl_),
    .din(G46)
  );


  splt
  gG46_spl_
  (
    .dout(G46_spl_0),
    .din(G46_spl_)
  );


  splt
  gG46_spl_0
  (
    .dout(G46_spl_00),
    .din(G46_spl_0)
  );


  splt
  gG46_spl_
  (
    .dout(G46_spl_1),
    .din(G46_spl_)
  );


  splt
  gG47
  (
    .dout(G47_spl_),
    .din(G47)
  );


  splt
  gG47_spl_
  (
    .dout(G47_spl_0),
    .din(G47_spl_)
  );


  splt
  gG47_spl_0
  (
    .dout(G47_spl_00),
    .din(G47_spl_0)
  );


  splt
  gG47_spl_
  (
    .dout(G47_spl_1),
    .din(G47_spl_)
  );


  splt
  gG48
  (
    .dout(G48_spl_),
    .din(G48)
  );


  splt
  gG48_spl_
  (
    .dout(G48_spl_0),
    .din(G48_spl_)
  );


  splt
  gG48_spl_0
  (
    .dout(G48_spl_00),
    .din(G48_spl_0)
  );


  splt
  gG48_spl_
  (
    .dout(G48_spl_1),
    .din(G48_spl_)
  );


  splt
  gnew_n157_
  (
    .dout(new_n157__spl_),
    .din(new_n157_)
  );


  splt
  gnew_n160_
  (
    .dout(new_n160__spl_),
    .din(new_n160_)
  );


  splt
  gG49
  (
    .dout(G49_spl_),
    .din(G49)
  );


  splt
  gnew_n163_
  (
    .dout(new_n163__spl_),
    .din(new_n163_)
  );


  splt
  gnew_n154_
  (
    .dout(new_n154__spl_),
    .din(new_n154_)
  );


  splt
  gnew_n166_
  (
    .dout(new_n166__spl_),
    .din(new_n166_)
  );


  splt
  gG866
  (
    .dout(G866_spl_),
    .din(G866)
  );


  splt
  gG866_spl_
  (
    .dout(G866_spl_0),
    .din(G866_spl_)
  );


  splt
  gnew_n170_
  (
    .dout(new_n170__spl_),
    .din(new_n170_)
  );


  splt
  gnew_n171_
  (
    .dout(new_n171__spl_),
    .din(new_n171_)
  );


  splt
  gG39
  (
    .dout(G39_spl_),
    .din(G39)
  );


  splt
  gnew_n173_
  (
    .dout(new_n173__spl_),
    .din(new_n173_)
  );


  splt
  gnew_n173__spl_
  (
    .dout(new_n173__spl_0),
    .din(new_n173__spl_)
  );


  splt
  gnew_n173__spl_
  (
    .dout(new_n173__spl_1),
    .din(new_n173__spl_)
  );


  splt
  gG60
  (
    .dout(G60_spl_),
    .din(G60)
  );


  splt
  gG60_spl_
  (
    .dout(G60_spl_0),
    .din(G60_spl_)
  );


  splt
  gnew_n176_
  (
    .dout(new_n176__spl_),
    .din(new_n176_)
  );


  splt
  gnew_n188_
  (
    .dout(new_n188__spl_),
    .din(new_n188_)
  );


  splt
  gnew_n188__spl_
  (
    .dout(new_n188__spl_0),
    .din(new_n188__spl_)
  );


  splt
  gnew_n188__spl_0
  (
    .dout(new_n188__spl_00),
    .din(new_n188__spl_0)
  );


  splt
  gnew_n188__spl_0
  (
    .dout(new_n188__spl_01),
    .din(new_n188__spl_0)
  );


  splt
  gnew_n188__spl_
  (
    .dout(new_n188__spl_1),
    .din(new_n188__spl_)
  );


  splt
  gnew_n188__spl_1
  (
    .dout(new_n188__spl_10),
    .din(new_n188__spl_1)
  );


  splt
  gnew_n188__spl_1
  (
    .dout(new_n188__spl_11),
    .din(new_n188__spl_1)
  );


  splt
  gnew_n178_
  (
    .dout(new_n178__spl_),
    .din(new_n178_)
  );


  splt
  gnew_n178__spl_
  (
    .dout(new_n178__spl_0),
    .din(new_n178__spl_)
  );


  splt
  gnew_n178__spl_
  (
    .dout(new_n178__spl_1),
    .din(new_n178__spl_)
  );


  splt
  gnew_n191_
  (
    .dout(new_n191__spl_),
    .din(new_n191_)
  );


  splt
  gnew_n191__spl_
  (
    .dout(new_n191__spl_0),
    .din(new_n191__spl_)
  );


  splt
  gG53
  (
    .dout(G53_spl_),
    .din(G53)
  );


  splt
  gG53_spl_
  (
    .dout(G53_spl_0),
    .din(G53_spl_)
  );


  splt
  gG53_spl_0
  (
    .dout(G53_spl_00),
    .din(G53_spl_0)
  );


  splt
  gG53_spl_0
  (
    .dout(G53_spl_01),
    .din(G53_spl_0)
  );


  splt
  gG53_spl_
  (
    .dout(G53_spl_1),
    .din(G53_spl_)
  );


  splt
  gG53_spl_1
  (
    .dout(G53_spl_10),
    .din(G53_spl_1)
  );


  splt
  gG53_spl_1
  (
    .dout(G53_spl_11),
    .din(G53_spl_1)
  );


  splt
  gnew_n192_
  (
    .dout(new_n192__spl_),
    .din(new_n192_)
  );


  splt
  gnew_n192__spl_
  (
    .dout(new_n192__spl_0),
    .din(new_n192__spl_)
  );


  splt
  gnew_n194_
  (
    .dout(new_n194__spl_),
    .din(new_n194_)
  );


  splt
  gG51
  (
    .dout(G51_spl_),
    .din(G51)
  );


  splt
  gG51_spl_
  (
    .dout(G51_spl_0),
    .din(G51_spl_)
  );


  splt
  gG51_spl_0
  (
    .dout(G51_spl_00),
    .din(G51_spl_0)
  );


  splt
  gG51_spl_00
  (
    .dout(G51_spl_000),
    .din(G51_spl_00)
  );


  splt
  gG51_spl_00
  (
    .dout(G51_spl_001),
    .din(G51_spl_00)
  );


  splt
  gG51_spl_0
  (
    .dout(G51_spl_01),
    .din(G51_spl_0)
  );


  splt
  gG51_spl_01
  (
    .dout(G51_spl_010),
    .din(G51_spl_01)
  );


  splt
  gG51_spl_01
  (
    .dout(G51_spl_011),
    .din(G51_spl_01)
  );


  splt
  gG51_spl_
  (
    .dout(G51_spl_1),
    .din(G51_spl_)
  );


  splt
  gG51_spl_1
  (
    .dout(G51_spl_10),
    .din(G51_spl_1)
  );


  splt
  gG51_spl_1
  (
    .dout(G51_spl_11),
    .din(G51_spl_1)
  );


  splt
  gG58
  (
    .dout(G58_spl_),
    .din(G58)
  );


  splt
  gnew_n198_
  (
    .dout(new_n198__spl_),
    .din(new_n198_)
  );


  splt
  gG52
  (
    .dout(G52_spl_),
    .din(G52)
  );


  splt
  gG52_spl_
  (
    .dout(G52_spl_0),
    .din(G52_spl_)
  );


  splt
  gG52_spl_0
  (
    .dout(G52_spl_00),
    .din(G52_spl_0)
  );


  splt
  gG52_spl_0
  (
    .dout(G52_spl_01),
    .din(G52_spl_0)
  );


  splt
  gG52_spl_
  (
    .dout(G52_spl_1),
    .din(G52_spl_)
  );


  splt
  gG52_spl_1
  (
    .dout(G52_spl_10),
    .din(G52_spl_1)
  );


  splt
  gG52_spl_1
  (
    .dout(G52_spl_11),
    .din(G52_spl_1)
  );


  splt
  gG54
  (
    .dout(G54_spl_),
    .din(G54)
  );


  splt
  gG54_spl_
  (
    .dout(G54_spl_0),
    .din(G54_spl_)
  );


  splt
  gG54_spl_0
  (
    .dout(G54_spl_00),
    .din(G54_spl_0)
  );


  splt
  gG54_spl_0
  (
    .dout(G54_spl_01),
    .din(G54_spl_0)
  );


  splt
  gG54_spl_
  (
    .dout(G54_spl_1),
    .din(G54_spl_)
  );


  splt
  gG54_spl_1
  (
    .dout(G54_spl_10),
    .din(G54_spl_1)
  );


  splt
  gG54_spl_1
  (
    .dout(G54_spl_11),
    .din(G54_spl_1)
  );


  splt
  gnew_n207_
  (
    .dout(new_n207__spl_),
    .din(new_n207_)
  );


  splt
  gnew_n207__spl_
  (
    .dout(new_n207__spl_0),
    .din(new_n207__spl_)
  );


  splt
  gnew_n207__spl_0
  (
    .dout(new_n207__spl_00),
    .din(new_n207__spl_0)
  );


  splt
  gnew_n207__spl_0
  (
    .dout(new_n207__spl_01),
    .din(new_n207__spl_0)
  );


  splt
  gnew_n207__spl_
  (
    .dout(new_n207__spl_1),
    .din(new_n207__spl_)
  );


  splt
  gnew_n207__spl_1
  (
    .dout(new_n207__spl_10),
    .din(new_n207__spl_1)
  );


  splt
  gnew_n207__spl_1
  (
    .dout(new_n207__spl_11),
    .din(new_n207__spl_1)
  );


  splt
  gG55
  (
    .dout(G55_spl_),
    .din(G55)
  );


  splt
  gG55_spl_
  (
    .dout(G55_spl_0),
    .din(G55_spl_)
  );


  splt
  gG50
  (
    .dout(G50_spl_),
    .din(G50)
  );


  splt
  gG50_spl_
  (
    .dout(G50_spl_0),
    .din(G50_spl_)
  );


  splt
  gG50_spl_0
  (
    .dout(G50_spl_00),
    .din(G50_spl_0)
  );


  splt
  gG50_spl_0
  (
    .dout(G50_spl_01),
    .din(G50_spl_0)
  );


  splt
  gG50_spl_
  (
    .dout(G50_spl_1),
    .din(G50_spl_)
  );


  splt
  gG50_spl_1
  (
    .dout(G50_spl_10),
    .din(G50_spl_1)
  );


  splt
  gG50_spl_1
  (
    .dout(G50_spl_11),
    .din(G50_spl_1)
  );


  splt
  gG36
  (
    .dout(G36_spl_),
    .din(G36)
  );


  splt
  gnew_n218_
  (
    .dout(new_n218__spl_),
    .din(new_n218_)
  );


  splt
  gnew_n218__spl_
  (
    .dout(new_n218__spl_0),
    .din(new_n218__spl_)
  );


  splt
  gG37
  (
    .dout(G37_spl_),
    .din(G37)
  );


  splt
  gnew_n224_
  (
    .dout(new_n224__spl_),
    .din(new_n224_)
  );


  splt
  gnew_n224__spl_
  (
    .dout(new_n224__spl_0),
    .din(new_n224__spl_)
  );


  splt
  gnew_n226_
  (
    .dout(new_n226__spl_),
    .din(new_n226_)
  );


  splt
  gnew_n227_
  (
    .dout(new_n227__spl_),
    .din(new_n227_)
  );


  splt
  gnew_n225_
  (
    .dout(new_n225__spl_),
    .din(new_n225_)
  );


  splt
  gnew_n225__spl_
  (
    .dout(new_n225__spl_0),
    .din(new_n225__spl_)
  );


  splt
  gnew_n228_
  (
    .dout(new_n228__spl_),
    .din(new_n228_)
  );


  splt
  gnew_n220_
  (
    .dout(new_n220__spl_),
    .din(new_n220_)
  );


  splt
  gnew_n229_
  (
    .dout(new_n229__spl_),
    .din(new_n229_)
  );


  splt
  gnew_n219_
  (
    .dout(new_n219__spl_),
    .din(new_n219_)
  );


  splt
  gnew_n219__spl_
  (
    .dout(new_n219__spl_0),
    .din(new_n219__spl_)
  );


  splt
  gnew_n230_
  (
    .dout(new_n230__spl_),
    .din(new_n230_)
  );


  splt
  gnew_n231_
  (
    .dout(new_n231__spl_),
    .din(new_n231_)
  );


  splt
  gG35
  (
    .dout(G35_spl_),
    .din(G35)
  );


  splt
  gnew_n236_
  (
    .dout(new_n236__spl_),
    .din(new_n236_)
  );


  splt
  gnew_n236__spl_
  (
    .dout(new_n236__spl_0),
    .din(new_n236__spl_)
  );


  splt
  gnew_n237_
  (
    .dout(new_n237__spl_),
    .din(new_n237_)
  );


  splt
  gnew_n237__spl_
  (
    .dout(new_n237__spl_0),
    .din(new_n237__spl_)
  );


  splt
  gnew_n239_
  (
    .dout(new_n239__spl_),
    .din(new_n239_)
  );


  splt
  gnew_n242_
  (
    .dout(new_n242__spl_),
    .din(new_n242_)
  );


  splt
  gnew_n286_
  (
    .dout(new_n286__spl_),
    .din(new_n286_)
  );


  splt
  gnew_n286__spl_
  (
    .dout(new_n286__spl_0),
    .din(new_n286__spl_)
  );


  splt
  gnew_n286__spl_
  (
    .dout(new_n286__spl_1),
    .din(new_n286__spl_)
  );


  splt
  gG34
  (
    .dout(G34_spl_),
    .din(G34)
  );


  splt
  gG34_spl_
  (
    .dout(G34_spl_0),
    .din(G34_spl_)
  );


  splt
  gG34_spl_
  (
    .dout(G34_spl_1),
    .din(G34_spl_)
  );


  splt
  gnew_n290_
  (
    .dout(new_n290__spl_),
    .din(new_n290_)
  );


  splt
  gnew_n290__spl_
  (
    .dout(new_n290__spl_0),
    .din(new_n290__spl_)
  );


  splt
  gnew_n290__spl_
  (
    .dout(new_n290__spl_1),
    .din(new_n290__spl_)
  );


  splt
  gnew_n293_
  (
    .dout(new_n293__spl_),
    .din(new_n293_)
  );


  splt
  gnew_n293__spl_
  (
    .dout(new_n293__spl_0),
    .din(new_n293__spl_)
  );


  splt
  gnew_n300_
  (
    .dout(new_n300__spl_),
    .din(new_n300_)
  );


  splt
  gnew_n300__spl_
  (
    .dout(new_n300__spl_0),
    .din(new_n300__spl_)
  );


  splt
  gnew_n308_
  (
    .dout(new_n308__spl_),
    .din(new_n308_)
  );


  splt
  gnew_n308__spl_
  (
    .dout(new_n308__spl_0),
    .din(new_n308__spl_)
  );


  splt
  gnew_n317_
  (
    .dout(new_n317__spl_),
    .din(new_n317_)
  );


  splt
  gnew_n317__spl_
  (
    .dout(new_n317__spl_0),
    .din(new_n317__spl_)
  );


  splt
  gnew_n311_
  (
    .dout(new_n311__spl_),
    .din(new_n311_)
  );


  splt
  gnew_n311__spl_
  (
    .dout(new_n311__spl_0),
    .din(new_n311__spl_)
  );


  splt
  gnew_n318_
  (
    .dout(new_n318__spl_),
    .din(new_n318_)
  );


  splt
  gnew_n320_
  (
    .dout(new_n320__spl_),
    .din(new_n320_)
  );


  splt
  gnew_n320__spl_
  (
    .dout(new_n320__spl_0),
    .din(new_n320__spl_)
  );


  splt
  gnew_n310_
  (
    .dout(new_n310__spl_),
    .din(new_n310_)
  );


  splt
  gnew_n321_
  (
    .dout(new_n321__spl_),
    .din(new_n321_)
  );


  splt
  gnew_n321__spl_
  (
    .dout(new_n321__spl_0),
    .din(new_n321__spl_)
  );


  splt
  gnew_n309_
  (
    .dout(new_n309__spl_),
    .din(new_n309_)
  );


  splt
  gnew_n309__spl_
  (
    .dout(new_n309__spl_0),
    .din(new_n309__spl_)
  );


  splt
  gnew_n302_
  (
    .dout(new_n302__spl_),
    .din(new_n302_)
  );


  splt
  gnew_n323_
  (
    .dout(new_n323__spl_),
    .din(new_n323_)
  );


  splt
  gnew_n323__spl_
  (
    .dout(new_n323__spl_0),
    .din(new_n323__spl_)
  );


  splt
  gnew_n301_
  (
    .dout(new_n301__spl_),
    .din(new_n301_)
  );


  splt
  gnew_n301__spl_
  (
    .dout(new_n301__spl_0),
    .din(new_n301__spl_)
  );


  splt
  gnew_n325_
  (
    .dout(new_n325__spl_),
    .din(new_n325_)
  );


  splt
  gnew_n325__spl_
  (
    .dout(new_n325__spl_0),
    .din(new_n325__spl_)
  );


  splt
  gnew_n326_
  (
    .dout(new_n326__spl_),
    .din(new_n326_)
  );


  splt
  gnew_n294_
  (
    .dout(new_n294__spl_),
    .din(new_n294_)
  );


  splt
  gnew_n294__spl_
  (
    .dout(new_n294__spl_0),
    .din(new_n294__spl_)
  );


  splt
  gnew_n329_
  (
    .dout(new_n329__spl_),
    .din(new_n329_)
  );


  splt
  gnew_n329__spl_
  (
    .dout(new_n329__spl_0),
    .din(new_n329__spl_)
  );


  splt
  gnew_n344_
  (
    .dout(new_n344__spl_),
    .din(new_n344_)
  );


  splt
  gnew_n344__spl_
  (
    .dout(new_n344__spl_0),
    .din(new_n344__spl_)
  );


  splt
  gnew_n359_
  (
    .dout(new_n359__spl_),
    .din(new_n359_)
  );


  splt
  gnew_n359__spl_
  (
    .dout(new_n359__spl_0),
    .din(new_n359__spl_)
  );


  splt
  gnew_n374_
  (
    .dout(new_n374__spl_),
    .din(new_n374_)
  );


  splt
  gnew_n374__spl_
  (
    .dout(new_n374__spl_0),
    .din(new_n374__spl_)
  );


endmodule
