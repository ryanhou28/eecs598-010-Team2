module rrr(clk, X_0, Y_0, X_1, Y_1, X_2, Y_2, X_3, Y_3, S_0, S_1, S_2, S_3, Co);
input clk;
 input X_0, Y_0, X_1, Y_1, X_2, Y_2, X_3, Y_3;
 output S_0, S_1, S_2, S_3;
 output Co;
 wire w1, w2, w3;
 reg xw1, xw2, xw3;
 reg XX_1, XX_2, XX_3, XXX_2, XXX_3, XXXX_3;
 reg YY_1, YY_2, YY_3, YYY_2, YYY_3, YYYY_3;
 // reg SS_2, SS_1, SS_0, SSS_1, SSS_0, SSSS_0;
 reg SS_1, SS_0, SSS_0;
 reg sS_0, sS_1, sS_2;
 assign S_0 = sS_0;
 assign S_1 = sS_1;
 assign S_2 = sS_2;
 // instantiating 4 1-bit full adders in Verilog
 fulladder u1(X_0, Y_0, 1'b0, SSSS_0, w1);
 fulladder u2(XX_1, YY_1, xw1, SSS_1, w2);
 fulladder u3(XXX_2, YYY_2, xw2, SS_2, w3);
 fulladder u4(XXXX_3, YYYY_3, xw3, S_3, Co);
 always @ (posedge clk) begin
   XX_1 <= X_1;
   XX_2 <= X_2;
   XXX_2 <= XX_2;
   XX_3 <= X_3;
   XXX_3 <= XX_3;
   XXXX_3 <= XXX_3;
   YY_1 <= Y_1;
   YY_2 <= Y_2;
   YYY_2 <= YY_2;
   YY_3 <= Y_3;
   YYY_3 <= YY_3;
   YYYY_3 <= YYY_3;
   sS_0 <= SS_0;
   SS_0 <= SSS_0;
   SSS_0 <= SSSS_0;
   sS_1 <= SS_1;
   SS_1 <= SSS_1;
   sS_2 <= SS_2;
   xw1 <= w1;
   xw2 <= w2;
   xw3 <= w3;
 end
 initial begin
   XX_1 <= 1'b0;
   XX_2 <= 1'b0;
   XXX_2 <= 1'b0;
   XX_3 <= 1'b0;
   XXX_3 <= 1'b0;
   XXXX_3 <= 1'b0;
   YY_1 <= 1'b0;
   YY_2 <= 1'b0;
   YYY_2 <= 1'b0;
   YY_3 <= 1'b0;
   YYY_3 <= 1'b0;
   YYYY_3 <= 1'b0;
   sS_0 <= 1'b0;
   SS_0 <= 1'b0;
   SSS_0 <= 1'b0;
   sS_1 <= 1'b0;
   SS_1 <= 1'b0;
   sS_2 <= 1'b0;
   xw1 <= 1'b0;
   xw2 <= 1'b0;
   xw3 <= 1'b0;
 end
endmodule

module fulladder(X, Y, Ci, S, Co);
  input X, Y, Ci;
  output S, Co;
  wire w1,w2,w3;
  //Structural code for one bit full adder
  xor (w1, X, Y);
  xor (S, w1, Ci);
  and (w2, w1, Ci);
  and (w3, X, Y);
  or (Co, w2, w3);
endmodule
