
module mymod
(
  G1_p,
  G1_n,
  G2_p,
  G2_n,
  G3_p,
  G3_n,
  G4_p,
  G4_n,
  G5_p,
  G5_n,
  G6_p,
  G6_n,
  G7_p,
  G7_n,
  G8_p,
  G8_n,
  G9_p,
  G9_n,
  G10_p,
  G10_n,
  G11_p,
  G11_n,
  G12_p,
  G12_n,
  G13_p,
  G13_n,
  G14_p,
  G14_n,
  G15_p,
  G15_n,
  G16_p,
  G16_n,
  G17_p,
  G17_n,
  G18_p,
  G18_n,
  G19_p,
  G19_n,
  G20_p,
  G20_n,
  G21_p,
  G21_n,
  G22_p,
  G22_n,
  G23_p,
  G23_n,
  G24_p,
  G24_n,
  G25_p,
  G25_n,
  G26_p,
  G26_n,
  G27_p,
  G27_n,
  G28_p,
  G28_n,
  G29_p,
  G29_n,
  G30_p,
  G30_n,
  G31_p,
  G31_n,
  G32_p,
  G32_n,
  G33_p,
  G33_n,
  G34_p,
  G34_n,
  G35_p,
  G35_n,
  G36_p,
  G36_n,
  G37_p,
  G37_n,
  G38_p,
  G38_n,
  G39_p,
  G39_n,
  G40_p,
  G40_n,
  G41_p,
  G41_n,
  G42_p,
  G42_n,
  G43_p,
  G43_n,
  G44_p,
  G44_n,
  G45_p,
  G45_n,
  G46_p,
  G46_n,
  G47_p,
  G47_n,
  G48_p,
  G48_n,
  G49_p,
  G49_n,
  G50_p,
  G50_n,
  G51_p,
  G51_n,
  G52_p,
  G52_n,
  G53_p,
  G53_n,
  G54_p,
  G54_n,
  G55_p,
  G55_n,
  G56_p,
  G56_n,
  G57_p,
  G57_n,
  G58_p,
  G58_n,
  G59_p,
  G59_n,
  G60_p,
  G60_n,
  G855_p,
  G856_p,
  G857_p,
  G858_p,
  G859_p,
  G860_p,
  G861_p,
  G862_n,
  G863_n,
  G864_n,
  G865_n,
  G866_p,
  G867_p,
  G868_p,
  G869_n,
  G870_p,
  G871_p,
  G872_p,
  G873_p,
  G874_p,
  G875_p,
  G876_p,
  G877_p,
  G878_p,
  G879_p,
  G880_p
);

  input G1_p;input G1_n;input G2_p;input G2_n;input G3_p;input G3_n;input G4_p;input G4_n;input G5_p;input G5_n;input G6_p;input G6_n;input G7_p;input G7_n;input G8_p;input G8_n;input G9_p;input G9_n;input G10_p;input G10_n;input G11_p;input G11_n;input G12_p;input G12_n;input G13_p;input G13_n;input G14_p;input G14_n;input G15_p;input G15_n;input G16_p;input G16_n;input G17_p;input G17_n;input G18_p;input G18_n;input G19_p;input G19_n;input G20_p;input G20_n;input G21_p;input G21_n;input G22_p;input G22_n;input G23_p;input G23_n;input G24_p;input G24_n;input G25_p;input G25_n;input G26_p;input G26_n;input G27_p;input G27_n;input G28_p;input G28_n;input G29_p;input G29_n;input G30_p;input G30_n;input G31_p;input G31_n;input G32_p;input G32_n;input G33_p;input G33_n;input G34_p;input G34_n;input G35_p;input G35_n;input G36_p;input G36_n;input G37_p;input G37_n;input G38_p;input G38_n;input G39_p;input G39_n;input G40_p;input G40_n;input G41_p;input G41_n;input G42_p;input G42_n;input G43_p;input G43_n;input G44_p;input G44_n;input G45_p;input G45_n;input G46_p;input G46_n;input G47_p;input G47_n;input G48_p;input G48_n;input G49_p;input G49_n;input G50_p;input G50_n;input G51_p;input G51_n;input G52_p;input G52_n;input G53_p;input G53_n;input G54_p;input G54_n;input G55_p;input G55_n;input G56_p;input G56_n;input G57_p;input G57_n;input G58_p;input G58_n;input G59_p;input G59_n;input G60_p;input G60_n;
  output G855_p;output G856_p;output G857_p;output G858_p;output G859_p;output G860_p;output G861_p;output G862_n;output G863_n;output G864_n;output G865_n;output G866_p;output G867_p;output G868_p;output G869_n;output G870_p;output G871_p;output G872_p;output G873_p;output G874_p;output G875_p;output G876_p;output G877_p;output G878_p;output G879_p;output G880_p;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire G51_p;
  wire G51_n;
  wire G52_p;
  wire G52_n;
  wire G53_p;
  wire G53_n;
  wire G54_p;
  wire G54_n;
  wire G55_p;
  wire G55_n;
  wire G56_p;
  wire G56_n;
  wire G57_p;
  wire G57_n;
  wire G58_p;
  wire G58_n;
  wire G59_p;
  wire G59_n;
  wire G60_p;
  wire G60_n;
  wire g61_p;
  wire g61_n;
  wire g62_p;
  wire g62_n;
  wire g63_p;
  wire g63_n;
  wire g64_p;
  wire g64_n;
  wire g65_p;
  wire g65_n;
  wire g66_p;
  wire g66_n;
  wire g67_p;
  wire g67_n;
  wire g68_p;
  wire g68_n;
  wire g69_p;
  wire g69_n;
  wire g70_p;
  wire g70_n;
  wire g71_p;
  wire g71_n;
  wire g72_p;
  wire g72_n;
  wire g73_p;
  wire g73_n;
  wire g74_p;
  wire g74_n;
  wire g75_p;
  wire g75_n;
  wire g76_p;
  wire g76_n;
  wire g77_p;
  wire g77_n;
  wire g78_p;
  wire g78_n;
  wire g79_p;
  wire g79_n;
  wire g80_p;
  wire g80_n;
  wire g81_p;
  wire g81_n;
  wire g82_p;
  wire g82_n;
  wire g83_p;
  wire g83_n;
  wire g84_p;
  wire g84_n;
  wire g85_p;
  wire g85_n;
  wire g86_p;
  wire g86_n;
  wire g87_p;
  wire g87_n;
  wire g88_p;
  wire g88_n;
  wire g89_p;
  wire g89_n;
  wire g90_p;
  wire g90_n;
  wire g91_p;
  wire g91_n;
  wire g92_p;
  wire g92_n;
  wire g93_p;
  wire g93_n;
  wire g94_p;
  wire g94_n;
  wire g95_p;
  wire g95_n;
  wire g96_p;
  wire g96_n;
  wire g97_p;
  wire g97_n;
  wire g98_p;
  wire g98_n;
  wire g99_p;
  wire g99_n;
  wire g100_p;
  wire g100_n;
  wire g101_p;
  wire g101_n;
  wire g102_p;
  wire g102_n;
  wire g103_p;
  wire g103_n;
  wire g104_p;
  wire g104_n;
  wire g105_p;
  wire g105_n;
  wire g106_p;
  wire g106_n;
  wire g107_p;
  wire g107_n;
  wire g108_p;
  wire g108_n;
  wire g109_p;
  wire g109_n;
  wire g110_p;
  wire g110_n;
  wire g111_p;
  wire g111_n;
  wire g112_p;
  wire g112_n;
  wire g113_p;
  wire g113_n;
  wire g114_p;
  wire g114_n;
  wire g115_p;
  wire g115_n;
  wire g116_p;
  wire g116_n;
  wire g117_p;
  wire g117_n;
  wire g118_p;
  wire g118_n;
  wire g119_p;
  wire g119_n;
  wire g120_p;
  wire g120_n;
  wire g121_p;
  wire g121_n;
  wire g122_p;
  wire g122_n;
  wire g123_p;
  wire g123_n;
  wire g124_p;
  wire g124_n;
  wire g125_p;
  wire g125_n;
  wire g126_p;
  wire g126_n;
  wire g127_p;
  wire g127_n;
  wire g128_p;
  wire g128_n;
  wire g129_p;
  wire g129_n;
  wire g130_p;
  wire g130_n;
  wire g131_p;
  wire g131_n;
  wire g132_p;
  wire g132_n;
  wire g133_p;
  wire g133_n;
  wire g134_p;
  wire g134_n;
  wire g135_p;
  wire g135_n;
  wire g136_p;
  wire g136_n;
  wire g137_p;
  wire g137_n;
  wire g138_p;
  wire g138_n;
  wire g139_p;
  wire g139_n;
  wire g140_p;
  wire g140_n;
  wire g141_p;
  wire g141_n;
  wire g142_p;
  wire g142_n;
  wire g143_p;
  wire g143_n;
  wire g144_p;
  wire g144_n;
  wire g145_p;
  wire g145_n;
  wire g146_p;
  wire g146_n;
  wire g147_p;
  wire g147_n;
  wire g148_p;
  wire g148_n;
  wire g149_p;
  wire g149_n;
  wire g150_p;
  wire g150_n;
  wire g151_p;
  wire g151_n;
  wire g152_p;
  wire g152_n;
  wire g153_p;
  wire g153_n;
  wire g154_p;
  wire g154_n;
  wire g155_p;
  wire g155_n;
  wire g156_p;
  wire g156_n;
  wire g157_p;
  wire g157_n;
  wire g158_p;
  wire g158_n;
  wire g159_p;
  wire g159_n;
  wire g160_p;
  wire g160_n;
  wire g161_p;
  wire g161_n;
  wire g162_p;
  wire g162_n;
  wire g163_p;
  wire g163_n;
  wire g164_p;
  wire g164_n;
  wire g165_p;
  wire g165_n;
  wire g166_p;
  wire g166_n;
  wire g167_p;
  wire g167_n;
  wire g168_p;
  wire g168_n;
  wire g169_p;
  wire g169_n;
  wire g170_p;
  wire g170_n;
  wire g171_p;
  wire g171_n;
  wire g172_p;
  wire g172_n;
  wire g173_p;
  wire g173_n;
  wire g174_p;
  wire g174_n;
  wire g175_p;
  wire g175_n;
  wire g176_p;
  wire g176_n;
  wire g177_p;
  wire g177_n;
  wire g178_p;
  wire g178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire G16_p_spl_;
  wire G6_n_spl_;
  wire G6_n_spl_0;
  wire G16_n_spl_;
  wire G8_n_spl_;
  wire G8_n_spl_0;
  wire G8_n_spl_00;
  wire G8_n_spl_01;
  wire G8_n_spl_1;
  wire G8_n_spl_10;
  wire g61_n_spl_;
  wire G7_n_spl_;
  wire G17_n_spl_;
  wire G17_n_spl_0;
  wire g63_n_spl_;
  wire G1_p_spl_;
  wire G1_p_spl_0;
  wire G2_p_spl_;
  wire G1_n_spl_;
  wire G1_n_spl_0;
  wire G2_n_spl_;
  wire G3_n_spl_;
  wire g67_n_spl_;
  wire G4_n_spl_;
  wire G4_n_spl_0;
  wire G4_n_spl_00;
  wire G4_n_spl_01;
  wire G4_n_spl_1;
  wire G4_n_spl_10;
  wire G4_n_spl_11;
  wire g68_n_spl_;
  wire g70_p_spl_;
  wire g70_n_spl_;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_00;
  wire G4_p_spl_01;
  wire G4_p_spl_1;
  wire G4_p_spl_10;
  wire g65_n_spl_;
  wire g65_n_spl_0;
  wire G11_p_spl_;
  wire G11_n_spl_;
  wire G11_n_spl_0;
  wire G11_n_spl_1;
  wire G17_p_spl_;
  wire g74_p_spl_;
  wire g76_n_spl_;
  wire g79_n_spl_;
  wire G9_p_spl_;
  wire G9_p_spl_0;
  wire G9_n_spl_;
  wire G9_n_spl_0;
  wire G10_n_spl_;
  wire G10_n_spl_0;
  wire g83_n_spl_;
  wire g83_n_spl_0;
  wire G12_n_spl_;
  wire g86_n_spl_;
  wire G24_p_spl_;
  wire G24_p_spl_0;
  wire G25_n_spl_;
  wire G25_n_spl_0;
  wire G25_n_spl_1;
  wire G24_n_spl_;
  wire G24_n_spl_0;
  wire G24_n_spl_1;
  wire G25_p_spl_;
  wire G25_p_spl_0;
  wire G26_p_spl_;
  wire G26_p_spl_0;
  wire G27_n_spl_;
  wire G27_n_spl_0;
  wire G27_n_spl_1;
  wire G26_n_spl_;
  wire G26_n_spl_0;
  wire G26_n_spl_1;
  wire G27_p_spl_;
  wire G27_p_spl_0;
  wire g92_p_spl_;
  wire g95_p_spl_;
  wire g92_n_spl_;
  wire g95_n_spl_;
  wire G32_p_spl_;
  wire G32_p_spl_0;
  wire G32_p_spl_1;
  wire g98_p_spl_;
  wire G32_n_spl_;
  wire G32_n_spl_0;
  wire G32_n_spl_1;
  wire g98_n_spl_;
  wire G28_p_spl_;
  wire G28_p_spl_0;
  wire G29_n_spl_;
  wire G29_n_spl_0;
  wire G29_n_spl_1;
  wire G28_n_spl_;
  wire G28_n_spl_0;
  wire G28_n_spl_1;
  wire G29_p_spl_;
  wire G29_p_spl_0;
  wire G30_p_spl_;
  wire G30_p_spl_0;
  wire G31_n_spl_;
  wire G31_n_spl_0;
  wire G30_n_spl_;
  wire G30_n_spl_0;
  wire G30_n_spl_1;
  wire G31_p_spl_;
  wire G31_p_spl_0;
  wire g104_p_spl_;
  wire g107_p_spl_;
  wire g104_n_spl_;
  wire g107_n_spl_;
  wire G33_p_spl_;
  wire g110_p_spl_;
  wire G33_n_spl_;
  wire g110_n_spl_;
  wire G41_p_spl_;
  wire G41_p_spl_0;
  wire G41_p_spl_1;
  wire G42_n_spl_;
  wire G42_n_spl_0;
  wire G42_n_spl_00;
  wire G42_n_spl_1;
  wire G41_n_spl_;
  wire G41_n_spl_0;
  wire G41_n_spl_00;
  wire G41_n_spl_1;
  wire G42_p_spl_;
  wire G42_p_spl_0;
  wire G42_p_spl_1;
  wire G43_p_spl_;
  wire G43_p_spl_0;
  wire G43_p_spl_1;
  wire G44_n_spl_;
  wire G44_n_spl_0;
  wire G44_n_spl_00;
  wire G44_n_spl_1;
  wire G43_n_spl_;
  wire G43_n_spl_0;
  wire G43_n_spl_00;
  wire G43_n_spl_1;
  wire G44_p_spl_;
  wire G44_p_spl_0;
  wire G44_p_spl_1;
  wire g119_p_spl_;
  wire g122_p_spl_;
  wire g119_n_spl_;
  wire g122_n_spl_;
  wire g125_p_spl_;
  wire g125_n_spl_;
  wire G45_p_spl_;
  wire G45_p_spl_0;
  wire G45_p_spl_1;
  wire G46_n_spl_;
  wire G46_n_spl_0;
  wire G46_n_spl_00;
  wire G46_n_spl_1;
  wire G45_n_spl_;
  wire G45_n_spl_0;
  wire G45_n_spl_00;
  wire G45_n_spl_1;
  wire G46_p_spl_;
  wire G46_p_spl_0;
  wire G46_p_spl_1;
  wire G47_p_spl_;
  wire G47_p_spl_0;
  wire G47_p_spl_1;
  wire G48_n_spl_;
  wire G48_n_spl_0;
  wire G48_n_spl_00;
  wire G48_n_spl_1;
  wire G47_n_spl_;
  wire G47_n_spl_0;
  wire G47_n_spl_00;
  wire G47_n_spl_1;
  wire G48_p_spl_;
  wire G48_p_spl_0;
  wire G48_p_spl_1;
  wire g131_p_spl_;
  wire g134_p_spl_;
  wire g131_n_spl_;
  wire g134_n_spl_;
  wire G49_p_spl_;
  wire g137_p_spl_;
  wire G49_n_spl_;
  wire g137_n_spl_;
  wire G55_n_spl_;
  wire G55_n_spl_0;
  wire G50_n_spl_;
  wire G50_n_spl_0;
  wire G50_n_spl_00;
  wire G50_n_spl_01;
  wire G50_n_spl_1;
  wire G50_n_spl_10;
  wire G50_n_spl_11;
  wire g82_p_spl_;
  wire g82_p_spl_0;
  wire g82_n_spl_;
  wire g82_n_spl_0;
  wire g82_n_spl_1;
  wire G10_p_spl_;
  wire g147_p_spl_;
  wire g147_n_spl_;
  wire G60_n_spl_;
  wire G60_n_spl_0;
  wire G60_p_spl_;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire g153_p_spl_;
  wire g153_n_spl_;
  wire g160_n_spl_;
  wire g160_n_spl_0;
  wire g160_n_spl_00;
  wire g160_n_spl_01;
  wire g160_n_spl_1;
  wire g160_n_spl_10;
  wire g160_n_spl_11;
  wire g160_p_spl_;
  wire g160_p_spl_0;
  wire g160_p_spl_00;
  wire g160_p_spl_01;
  wire g160_p_spl_1;
  wire g160_p_spl_10;
  wire g160_p_spl_11;
  wire g162_p_spl_;
  wire g162_n_spl_;
  wire G39_p_spl_;
  wire g164_n_spl_;
  wire g164_n_spl_0;
  wire g164_n_spl_1;
  wire G39_n_spl_;
  wire g164_p_spl_;
  wire g164_p_spl_0;
  wire g164_p_spl_1;
  wire g149_n_spl_;
  wire g149_n_spl_0;
  wire g149_n_spl_1;
  wire g149_p_spl_;
  wire g149_p_spl_0;
  wire g149_p_spl_1;
  wire G54_n_spl_;
  wire G54_n_spl_0;
  wire G54_n_spl_00;
  wire G54_n_spl_01;
  wire G54_n_spl_1;
  wire G54_n_spl_10;
  wire G54_n_spl_11;
  wire g167_p_spl_;
  wire g167_p_spl_0;
  wire g172_n_spl_;
  wire g172_n_spl_0;
  wire g172_n_spl_00;
  wire g172_n_spl_01;
  wire g172_n_spl_1;
  wire g172_n_spl_10;
  wire g172_n_spl_11;
  wire g167_n_spl_;
  wire G53_n_spl_;
  wire G53_n_spl_0;
  wire G53_n_spl_00;
  wire G53_n_spl_01;
  wire G53_n_spl_1;
  wire G53_n_spl_10;
  wire G53_n_spl_11;
  wire g174_p_spl_;
  wire g176_p_spl_;
  wire G51_n_spl_;
  wire G51_n_spl_0;
  wire G51_n_spl_00;
  wire G51_n_spl_000;
  wire G51_n_spl_001;
  wire G51_n_spl_01;
  wire G51_n_spl_010;
  wire G51_n_spl_011;
  wire G51_n_spl_1;
  wire G51_n_spl_10;
  wire G51_n_spl_11;
  wire G58_n_spl_;
  wire g180_p_spl_;
  wire G52_n_spl_;
  wire G52_n_spl_0;
  wire G52_n_spl_00;
  wire G52_n_spl_01;
  wire G52_n_spl_1;
  wire G52_n_spl_10;
  wire G52_n_spl_11;
  wire g174_n_spl_;
  wire G35_p_spl_;
  wire G35_n_spl_;
  wire g194_p_spl_;
  wire g194_p_spl_0;
  wire G36_p_spl_;
  wire G36_n_spl_;
  wire g199_n_spl_;
  wire g199_p_spl_;
  wire g199_p_spl_0;
  wire G37_p_spl_;
  wire G37_n_spl_;
  wire g205_n_spl_;
  wire g205_p_spl_;
  wire g205_p_spl_0;
  wire g207_p_spl_;
  wire g208_p_spl_;
  wire g206_n_spl_;
  wire g206_p_spl_;
  wire g209_p_spl_;
  wire g201_p_spl_;
  wire g210_p_spl_;
  wire g200_n_spl_;
  wire g200_p_spl_;
  wire g211_p_spl_;
  wire g212_p_spl_;
  wire g194_n_spl_;
  wire g214_p_spl_;
  wire g216_p_spl_;
  wire g219_p_spl_;
  wire g214_n_spl_;
  wire g259_p_spl_;
  wire g259_p_spl_0;
  wire g259_p_spl_1;
  wire g259_n_spl_;
  wire g259_n_spl_0;
  wire g259_n_spl_1;
  wire G34_p_spl_;
  wire G34_p_spl_0;
  wire G34_p_spl_1;
  wire G34_n_spl_;
  wire G34_n_spl_0;
  wire G34_n_spl_1;
  wire g265_n_spl_;
  wire g265_n_spl_0;
  wire g265_n_spl_1;
  wire g265_p_spl_;
  wire g265_p_spl_0;
  wire g265_p_spl_1;
  wire g267_n_spl_;
  wire g267_p_spl_;
  wire g267_p_spl_0;
  wire g274_n_spl_;
  wire g274_p_spl_;
  wire g274_p_spl_0;
  wire g282_n_spl_;
  wire g282_p_spl_;
  wire g282_p_spl_0;
  wire g291_p_spl_;
  wire g291_p_spl_0;
  wire g291_n_spl_;
  wire g285_n_spl_;
  wire g292_n_spl_;
  wire g285_p_spl_;
  wire g292_p_spl_;
  wire g294_n_spl_;
  wire g294_n_spl_0;
  wire g294_p_spl_;
  wire g284_n_spl_;
  wire g295_n_spl_;
  wire g284_p_spl_;
  wire g295_p_spl_;
  wire g283_n_spl_;
  wire g283_n_spl_0;
  wire g283_p_spl_;
  wire g276_n_spl_;
  wire g297_n_spl_;
  wire g276_p_spl_;
  wire g297_p_spl_;
  wire g275_n_spl_;
  wire g275_n_spl_0;
  wire g275_p_spl_;
  wire g299_p_spl_;
  wire g300_p_spl_;
  wire g268_n_spl_;
  wire g268_n_spl_0;
  wire g303_n_spl_;
  wire g322_n_spl_;
  wire g337_n_spl_;
  wire g352_n_spl_;

  LA
  g_g61_p
  (
    .dout(g61_p),
    .din1(G6_p),
    .din2(G16_p_spl_)
  );


  FA
  g_g61_n
  (
    .dout(g61_n),
    .din1(G6_n_spl_0),
    .din2(G16_n_spl_)
  );


  FA
  g_g62_n
  (
    .dout(g62_n),
    .din1(G8_n_spl_00),
    .din2(g61_n_spl_)
  );


  FA
  g_g63_n
  (
    .dout(g63_n),
    .din1(G6_n_spl_0),
    .din2(G7_n_spl_)
  );


  FA
  g_g64_n
  (
    .dout(g64_n),
    .din1(G17_n_spl_0),
    .din2(g63_n_spl_)
  );


  FA
  g_g65_n
  (
    .dout(g65_n),
    .din1(G8_n_spl_00),
    .din2(g63_n_spl_)
  );


  FA
  g_g66_n
  (
    .dout(g66_n),
    .din1(G18_n),
    .din2(G19_n)
  );


  LA
  g_g67_p
  (
    .dout(g67_p),
    .din1(G1_p_spl_0),
    .din2(G2_p_spl_)
  );


  FA
  g_g67_n
  (
    .dout(g67_n),
    .din1(G1_n_spl_0),
    .din2(G2_n_spl_)
  );


  FA
  g_g68_n
  (
    .dout(g68_n),
    .din1(G3_n_spl_),
    .din2(g67_n_spl_)
  );


  FA
  g_g69_n
  (
    .dout(g69_n),
    .din1(G4_n_spl_00),
    .din2(g68_n_spl_)
  );


  LA
  g_g70_p
  (
    .dout(g70_p),
    .din1(G1_p_spl_0),
    .din2(G5_p)
  );


  FA
  g_g70_n
  (
    .dout(g70_n),
    .din1(G1_n_spl_0),
    .din2(G5_n)
  );


  LA
  g_g71_p
  (
    .dout(g71_p),
    .din1(G3_p),
    .din2(g70_p_spl_)
  );


  FA
  g_g71_n
  (
    .dout(g71_n),
    .din1(G3_n_spl_),
    .din2(g70_n_spl_)
  );


  LA
  g_g72_p
  (
    .dout(g72_p),
    .din1(G4_p_spl_00),
    .din2(g71_p)
  );


  FA
  g_g72_n
  (
    .dout(g72_n),
    .din1(G4_n_spl_00),
    .din2(g71_n)
  );


  LA
  g_g73_p
  (
    .dout(g73_p),
    .din1(g65_n_spl_0),
    .din2(g72_p)
  );


  LA
  g_g74_p
  (
    .dout(g74_p),
    .din1(G11_p_spl_),
    .din2(G16_p_spl_)
  );


  FA
  g_g74_n
  (
    .dout(g74_n),
    .din1(G11_n_spl_0),
    .din2(G16_n_spl_)
  );


  LA
  g_g75_p
  (
    .dout(g75_p),
    .din1(G17_p_spl_),
    .din2(g74_p_spl_)
  );


  FA
  g_g76_n
  (
    .dout(g76_n),
    .din1(G7_n_spl_),
    .din2(G11_n_spl_0)
  );


  FA
  g_g77_n
  (
    .dout(g77_n),
    .din1(G17_n_spl_0),
    .din2(g76_n_spl_)
  );


  FA
  g_g78_n
  (
    .dout(g78_n),
    .din1(G8_n_spl_01),
    .din2(g76_n_spl_)
  );


  FA
  g_g79_n
  (
    .dout(g79_n),
    .din1(G20_p),
    .din2(G21_p)
  );


  LA
  g_g80_p
  (
    .dout(g80_p),
    .din1(G23_p),
    .din2(g79_n_spl_)
  );


  FA
  g_g81_n
  (
    .dout(g81_n),
    .din1(g65_n_spl_0),
    .din2(g72_n)
  );


  LA
  g_g82_p
  (
    .dout(g82_p),
    .din1(G9_p_spl_0),
    .din2(g70_p_spl_)
  );


  FA
  g_g82_n
  (
    .dout(g82_n),
    .din1(G9_n_spl_0),
    .din2(g70_n_spl_)
  );


  FA
  g_g83_n
  (
    .dout(g83_n),
    .din1(G10_n_spl_0),
    .din2(g68_n_spl_)
  );


  FA
  g_g84_n
  (
    .dout(g84_n),
    .din1(G6_n_spl_),
    .din2(g83_n_spl_0)
  );


  FA
  g_g85_n
  (
    .dout(g85_n),
    .din1(G12_n_spl_),
    .din2(g84_n)
  );


  FA
  g_g86_n
  (
    .dout(g86_n),
    .din1(G11_n_spl_1),
    .din2(G12_n_spl_)
  );


  FA
  g_g87_n
  (
    .dout(g87_n),
    .din1(G15_n),
    .din2(g83_n_spl_0)
  );


  FA
  g_g88_n
  (
    .dout(g88_n),
    .din1(g86_n_spl_),
    .din2(g87_n)
  );


  LA
  g_g89_p
  (
    .dout(g89_p),
    .din1(G22_p),
    .din2(g79_n_spl_)
  );


  LA
  g_g90_p
  (
    .dout(g90_p),
    .din1(G24_p_spl_0),
    .din2(G25_n_spl_0)
  );


  FA
  g_g90_n
  (
    .dout(g90_n),
    .din1(G24_n_spl_0),
    .din2(G25_p_spl_0)
  );


  LA
  g_g91_p
  (
    .dout(g91_p),
    .din1(G24_n_spl_0),
    .din2(G25_p_spl_0)
  );


  FA
  g_g91_n
  (
    .dout(g91_n),
    .din1(G24_p_spl_0),
    .din2(G25_n_spl_0)
  );


  LA
  g_g92_p
  (
    .dout(g92_p),
    .din1(g90_n),
    .din2(g91_n)
  );


  FA
  g_g92_n
  (
    .dout(g92_n),
    .din1(g90_p),
    .din2(g91_p)
  );


  LA
  g_g93_p
  (
    .dout(g93_p),
    .din1(G26_p_spl_0),
    .din2(G27_n_spl_0)
  );


  FA
  g_g93_n
  (
    .dout(g93_n),
    .din1(G26_n_spl_0),
    .din2(G27_p_spl_0)
  );


  LA
  g_g94_p
  (
    .dout(g94_p),
    .din1(G26_n_spl_0),
    .din2(G27_p_spl_0)
  );


  FA
  g_g94_n
  (
    .dout(g94_n),
    .din1(G26_p_spl_0),
    .din2(G27_n_spl_0)
  );


  LA
  g_g95_p
  (
    .dout(g95_p),
    .din1(g93_n),
    .din2(g94_n)
  );


  FA
  g_g95_n
  (
    .dout(g95_n),
    .din1(g93_p),
    .din2(g94_p)
  );


  LA
  g_g96_p
  (
    .dout(g96_p),
    .din1(g92_p_spl_),
    .din2(g95_p_spl_)
  );


  FA
  g_g96_n
  (
    .dout(g96_n),
    .din1(g92_n_spl_),
    .din2(g95_n_spl_)
  );


  LA
  g_g97_p
  (
    .dout(g97_p),
    .din1(g92_n_spl_),
    .din2(g95_n_spl_)
  );


  FA
  g_g97_n
  (
    .dout(g97_n),
    .din1(g92_p_spl_),
    .din2(g95_p_spl_)
  );


  LA
  g_g98_p
  (
    .dout(g98_p),
    .din1(g96_n),
    .din2(g97_n)
  );


  FA
  g_g98_n
  (
    .dout(g98_n),
    .din1(g96_p),
    .din2(g97_p)
  );


  LA
  g_g99_p
  (
    .dout(g99_p),
    .din1(G32_p_spl_0),
    .din2(g98_p_spl_)
  );


  FA
  g_g99_n
  (
    .dout(g99_n),
    .din1(G32_n_spl_0),
    .din2(g98_n_spl_)
  );


  LA
  g_g100_p
  (
    .dout(g100_p),
    .din1(G32_n_spl_0),
    .din2(g98_n_spl_)
  );


  FA
  g_g100_n
  (
    .dout(g100_n),
    .din1(G32_p_spl_0),
    .din2(g98_p_spl_)
  );


  LA
  g_g101_p
  (
    .dout(g101_p),
    .din1(g99_n),
    .din2(g100_n)
  );


  FA
  g_g101_n
  (
    .dout(g101_n),
    .din1(g99_p),
    .din2(g100_p)
  );


  LA
  g_g102_p
  (
    .dout(g102_p),
    .din1(G28_p_spl_0),
    .din2(G29_n_spl_0)
  );


  FA
  g_g102_n
  (
    .dout(g102_n),
    .din1(G28_n_spl_0),
    .din2(G29_p_spl_0)
  );


  LA
  g_g103_p
  (
    .dout(g103_p),
    .din1(G28_n_spl_0),
    .din2(G29_p_spl_0)
  );


  FA
  g_g103_n
  (
    .dout(g103_n),
    .din1(G28_p_spl_0),
    .din2(G29_n_spl_0)
  );


  LA
  g_g104_p
  (
    .dout(g104_p),
    .din1(g102_n),
    .din2(g103_n)
  );


  FA
  g_g104_n
  (
    .dout(g104_n),
    .din1(g102_p),
    .din2(g103_p)
  );


  LA
  g_g105_p
  (
    .dout(g105_p),
    .din1(G30_p_spl_0),
    .din2(G31_n_spl_0)
  );


  FA
  g_g105_n
  (
    .dout(g105_n),
    .din1(G30_n_spl_0),
    .din2(G31_p_spl_0)
  );


  LA
  g_g106_p
  (
    .dout(g106_p),
    .din1(G30_n_spl_0),
    .din2(G31_p_spl_0)
  );


  FA
  g_g106_n
  (
    .dout(g106_n),
    .din1(G30_p_spl_0),
    .din2(G31_n_spl_0)
  );


  LA
  g_g107_p
  (
    .dout(g107_p),
    .din1(g105_n),
    .din2(g106_n)
  );


  FA
  g_g107_n
  (
    .dout(g107_n),
    .din1(g105_p),
    .din2(g106_p)
  );


  LA
  g_g108_p
  (
    .dout(g108_p),
    .din1(g104_p_spl_),
    .din2(g107_p_spl_)
  );


  FA
  g_g108_n
  (
    .dout(g108_n),
    .din1(g104_n_spl_),
    .din2(g107_n_spl_)
  );


  LA
  g_g109_p
  (
    .dout(g109_p),
    .din1(g104_n_spl_),
    .din2(g107_n_spl_)
  );


  FA
  g_g109_n
  (
    .dout(g109_n),
    .din1(g104_p_spl_),
    .din2(g107_p_spl_)
  );


  LA
  g_g110_p
  (
    .dout(g110_p),
    .din1(g108_n),
    .din2(g109_n)
  );


  FA
  g_g110_n
  (
    .dout(g110_n),
    .din1(g108_p),
    .din2(g109_p)
  );


  LA
  g_g111_p
  (
    .dout(g111_p),
    .din1(G33_p_spl_),
    .din2(g110_p_spl_)
  );


  FA
  g_g111_n
  (
    .dout(g111_n),
    .din1(G33_n_spl_),
    .din2(g110_n_spl_)
  );


  LA
  g_g112_p
  (
    .dout(g112_p),
    .din1(G33_n_spl_),
    .din2(g110_n_spl_)
  );


  FA
  g_g112_n
  (
    .dout(g112_n),
    .din1(G33_p_spl_),
    .din2(g110_p_spl_)
  );


  LA
  g_g113_p
  (
    .dout(g113_p),
    .din1(g111_n),
    .din2(g112_n)
  );


  FA
  g_g113_n
  (
    .dout(g113_n),
    .din1(g111_p),
    .din2(g112_p)
  );


  LA
  g_g114_p
  (
    .dout(g114_p),
    .din1(g101_n),
    .din2(g113_n)
  );


  LA
  g_g115_p
  (
    .dout(g115_p),
    .din1(g101_p),
    .din2(g113_p)
  );


  FA
  g_g116_n
  (
    .dout(g116_n),
    .din1(g114_p),
    .din2(g115_p)
  );


  LA
  g_g117_p
  (
    .dout(g117_p),
    .din1(G41_p_spl_0),
    .din2(G42_n_spl_00)
  );


  FA
  g_g117_n
  (
    .dout(g117_n),
    .din1(G41_n_spl_00),
    .din2(G42_p_spl_0)
  );


  LA
  g_g118_p
  (
    .dout(g118_p),
    .din1(G41_n_spl_00),
    .din2(G42_p_spl_0)
  );


  FA
  g_g118_n
  (
    .dout(g118_n),
    .din1(G41_p_spl_0),
    .din2(G42_n_spl_00)
  );


  LA
  g_g119_p
  (
    .dout(g119_p),
    .din1(g117_n),
    .din2(g118_n)
  );


  FA
  g_g119_n
  (
    .dout(g119_n),
    .din1(g117_p),
    .din2(g118_p)
  );


  LA
  g_g120_p
  (
    .dout(g120_p),
    .din1(G43_p_spl_0),
    .din2(G44_n_spl_00)
  );


  FA
  g_g120_n
  (
    .dout(g120_n),
    .din1(G43_n_spl_00),
    .din2(G44_p_spl_0)
  );


  LA
  g_g121_p
  (
    .dout(g121_p),
    .din1(G43_n_spl_00),
    .din2(G44_p_spl_0)
  );


  FA
  g_g121_n
  (
    .dout(g121_n),
    .din1(G43_p_spl_0),
    .din2(G44_n_spl_00)
  );


  LA
  g_g122_p
  (
    .dout(g122_p),
    .din1(g120_n),
    .din2(g121_n)
  );


  FA
  g_g122_n
  (
    .dout(g122_n),
    .din1(g120_p),
    .din2(g121_p)
  );


  LA
  g_g123_p
  (
    .dout(g123_p),
    .din1(g119_p_spl_),
    .din2(g122_p_spl_)
  );


  FA
  g_g123_n
  (
    .dout(g123_n),
    .din1(g119_n_spl_),
    .din2(g122_n_spl_)
  );


  LA
  g_g124_p
  (
    .dout(g124_p),
    .din1(g119_n_spl_),
    .din2(g122_n_spl_)
  );


  FA
  g_g124_n
  (
    .dout(g124_n),
    .din1(g119_p_spl_),
    .din2(g122_p_spl_)
  );


  LA
  g_g125_p
  (
    .dout(g125_p),
    .din1(g123_n),
    .din2(g124_n)
  );


  FA
  g_g125_n
  (
    .dout(g125_n),
    .din1(g123_p),
    .din2(g124_p)
  );


  LA
  g_g126_p
  (
    .dout(g126_p),
    .din1(G32_p_spl_1),
    .din2(g125_p_spl_)
  );


  FA
  g_g126_n
  (
    .dout(g126_n),
    .din1(G32_n_spl_1),
    .din2(g125_n_spl_)
  );


  LA
  g_g127_p
  (
    .dout(g127_p),
    .din1(G32_n_spl_1),
    .din2(g125_n_spl_)
  );


  FA
  g_g127_n
  (
    .dout(g127_n),
    .din1(G32_p_spl_1),
    .din2(g125_p_spl_)
  );


  LA
  g_g128_p
  (
    .dout(g128_p),
    .din1(g126_n),
    .din2(g127_n)
  );


  FA
  g_g128_n
  (
    .dout(g128_n),
    .din1(g126_p),
    .din2(g127_p)
  );


  LA
  g_g129_p
  (
    .dout(g129_p),
    .din1(G45_p_spl_0),
    .din2(G46_n_spl_00)
  );


  FA
  g_g129_n
  (
    .dout(g129_n),
    .din1(G45_n_spl_00),
    .din2(G46_p_spl_0)
  );


  LA
  g_g130_p
  (
    .dout(g130_p),
    .din1(G45_n_spl_00),
    .din2(G46_p_spl_0)
  );


  FA
  g_g130_n
  (
    .dout(g130_n),
    .din1(G45_p_spl_0),
    .din2(G46_n_spl_00)
  );


  LA
  g_g131_p
  (
    .dout(g131_p),
    .din1(g129_n),
    .din2(g130_n)
  );


  FA
  g_g131_n
  (
    .dout(g131_n),
    .din1(g129_p),
    .din2(g130_p)
  );


  LA
  g_g132_p
  (
    .dout(g132_p),
    .din1(G47_p_spl_0),
    .din2(G48_n_spl_00)
  );


  FA
  g_g132_n
  (
    .dout(g132_n),
    .din1(G47_n_spl_00),
    .din2(G48_p_spl_0)
  );


  LA
  g_g133_p
  (
    .dout(g133_p),
    .din1(G47_n_spl_00),
    .din2(G48_p_spl_0)
  );


  FA
  g_g133_n
  (
    .dout(g133_n),
    .din1(G47_p_spl_0),
    .din2(G48_n_spl_00)
  );


  LA
  g_g134_p
  (
    .dout(g134_p),
    .din1(g132_n),
    .din2(g133_n)
  );


  FA
  g_g134_n
  (
    .dout(g134_n),
    .din1(g132_p),
    .din2(g133_p)
  );


  LA
  g_g135_p
  (
    .dout(g135_p),
    .din1(g131_p_spl_),
    .din2(g134_p_spl_)
  );


  FA
  g_g135_n
  (
    .dout(g135_n),
    .din1(g131_n_spl_),
    .din2(g134_n_spl_)
  );


  LA
  g_g136_p
  (
    .dout(g136_p),
    .din1(g131_n_spl_),
    .din2(g134_n_spl_)
  );


  FA
  g_g136_n
  (
    .dout(g136_n),
    .din1(g131_p_spl_),
    .din2(g134_p_spl_)
  );


  LA
  g_g137_p
  (
    .dout(g137_p),
    .din1(g135_n),
    .din2(g136_n)
  );


  FA
  g_g137_n
  (
    .dout(g137_n),
    .din1(g135_p),
    .din2(g136_p)
  );


  LA
  g_g138_p
  (
    .dout(g138_p),
    .din1(G49_p_spl_),
    .din2(g137_p_spl_)
  );


  FA
  g_g138_n
  (
    .dout(g138_n),
    .din1(G49_n_spl_),
    .din2(g137_n_spl_)
  );


  LA
  g_g139_p
  (
    .dout(g139_p),
    .din1(G49_n_spl_),
    .din2(g137_n_spl_)
  );


  FA
  g_g139_n
  (
    .dout(g139_n),
    .din1(G49_p_spl_),
    .din2(g137_p_spl_)
  );


  LA
  g_g140_p
  (
    .dout(g140_p),
    .din1(g138_n),
    .din2(g139_n)
  );


  FA
  g_g140_n
  (
    .dout(g140_n),
    .din1(g138_p),
    .din2(g139_p)
  );


  LA
  g_g141_p
  (
    .dout(g141_p),
    .din1(g128_n),
    .din2(g140_n)
  );


  LA
  g_g142_p
  (
    .dout(g142_p),
    .din1(g128_p),
    .din2(g140_p)
  );


  FA
  g_g143_n
  (
    .dout(g143_n),
    .din1(g141_p),
    .din2(g142_p)
  );


  FA
  g_g144_n
  (
    .dout(g144_n),
    .din1(G55_n_spl_0),
    .din2(G59_n)
  );


  FA
  g_g145_n
  (
    .dout(g145_n),
    .din1(G30_n_spl_1),
    .din2(G50_n_spl_00)
  );


  LA
  g_g146_p
  (
    .dout(g146_p),
    .din1(G17_p_spl_),
    .din2(g82_p_spl_0)
  );


  FA
  g_g146_n
  (
    .dout(g146_n),
    .din1(G17_n_spl_),
    .din2(g82_n_spl_0)
  );


  LA
  g_g147_p
  (
    .dout(g147_p),
    .din1(g61_p),
    .din2(g146_p)
  );


  FA
  g_g147_n
  (
    .dout(g147_n),
    .din1(g61_n_spl_),
    .din2(g146_n)
  );


  LA
  g_g148_p
  (
    .dout(g148_p),
    .din1(G10_p_spl_),
    .din2(g147_p_spl_)
  );


  FA
  g_g148_n
  (
    .dout(g148_n),
    .din1(G10_n_spl_0),
    .din2(g147_n_spl_)
  );


  LA
  g_g149_p
  (
    .dout(g149_p),
    .din1(G60_n_spl_0),
    .din2(g148_p)
  );


  FA
  g_g149_n
  (
    .dout(g149_n),
    .din1(G60_p_spl_),
    .din2(g148_n)
  );


  LA
  g_g150_p
  (
    .dout(g150_p),
    .din1(G4_n_spl_01),
    .din2(G8_n_spl_01)
  );


  FA
  g_g150_n
  (
    .dout(g150_n),
    .din1(G4_p_spl_00),
    .din2(G8_p_spl_0)
  );


  LA
  g_g151_p
  (
    .dout(g151_p),
    .din1(G4_p_spl_01),
    .din2(G8_p_spl_0)
  );


  FA
  g_g151_n
  (
    .dout(g151_n),
    .din1(G4_n_spl_01),
    .din2(G8_n_spl_10)
  );


  LA
  g_g152_p
  (
    .dout(g152_p),
    .din1(g150_n),
    .din2(g151_n)
  );


  FA
  g_g152_n
  (
    .dout(g152_n),
    .din1(g150_p),
    .din2(g151_p)
  );


  LA
  g_g153_p
  (
    .dout(g153_p),
    .din1(G11_p_spl_),
    .din2(G40_p)
  );


  FA
  g_g153_n
  (
    .dout(g153_n),
    .din1(G11_n_spl_1),
    .din2(G40_n)
  );


  LA
  g_g154_p
  (
    .dout(g154_p),
    .din1(g82_p_spl_0),
    .din2(g153_p_spl_)
  );


  FA
  g_g154_n
  (
    .dout(g154_n),
    .din1(g82_n_spl_0),
    .din2(g153_n_spl_)
  );


  LA
  g_g155_p
  (
    .dout(g155_p),
    .din1(g152_p),
    .din2(g154_p)
  );


  FA
  g_g155_n
  (
    .dout(g155_n),
    .din1(g152_n),
    .din2(g154_n)
  );


  LA
  g_g156_p
  (
    .dout(g156_p),
    .din1(G4_p_spl_01),
    .din2(g67_p)
  );


  FA
  g_g156_n
  (
    .dout(g156_n),
    .din1(G4_n_spl_10),
    .din2(g67_n_spl_)
  );


  LA
  g_g157_p
  (
    .dout(g157_p),
    .din1(G8_p_spl_),
    .din2(g74_p_spl_)
  );


  FA
  g_g157_n
  (
    .dout(g157_n),
    .din1(G8_n_spl_10),
    .din2(g74_n)
  );


  LA
  g_g158_p
  (
    .dout(g158_p),
    .din1(G9_p_spl_0),
    .din2(g157_n)
  );


  FA
  g_g158_n
  (
    .dout(g158_n),
    .din1(G9_n_spl_0),
    .din2(g157_p)
  );


  LA
  g_g159_p
  (
    .dout(g159_p),
    .din1(g156_p),
    .din2(g158_p)
  );


  FA
  g_g159_n
  (
    .dout(g159_n),
    .din1(g156_n),
    .din2(g158_n)
  );


  LA
  g_g160_p
  (
    .dout(g160_p),
    .din1(g155_n),
    .din2(g159_n)
  );


  FA
  g_g160_n
  (
    .dout(g160_n),
    .din1(g155_p),
    .din2(g159_p)
  );


  LA
  g_g161_p
  (
    .dout(g161_p),
    .din1(G31_p_spl_),
    .din2(g160_n_spl_00)
  );


  FA
  g_g161_n
  (
    .dout(g161_n),
    .din1(G31_n_spl_),
    .din2(g160_p_spl_00)
  );


  LA
  g_g162_p
  (
    .dout(g162_p),
    .din1(g82_p_spl_),
    .din2(g153_n_spl_)
  );


  FA
  g_g162_n
  (
    .dout(g162_n),
    .din1(g82_n_spl_1),
    .din2(g153_p_spl_)
  );


  LA
  g_g163_p
  (
    .dout(g163_p),
    .din1(G4_p_spl_10),
    .din2(g162_p_spl_)
  );


  FA
  g_g163_n
  (
    .dout(g163_n),
    .din1(G4_n_spl_10),
    .din2(g162_n_spl_)
  );


  LA
  g_g164_p
  (
    .dout(g164_p),
    .din1(G1_p_spl_),
    .din2(g163_n)
  );


  FA
  g_g164_n
  (
    .dout(g164_n),
    .din1(G1_n_spl_),
    .din2(g163_p)
  );


  LA
  g_g165_p
  (
    .dout(g165_p),
    .din1(G39_p_spl_),
    .din2(g164_n_spl_0)
  );


  FA
  g_g165_n
  (
    .dout(g165_n),
    .din1(G39_n_spl_),
    .din2(g164_p_spl_0)
  );


  LA
  g_g166_p
  (
    .dout(g166_p),
    .din1(g161_n),
    .din2(g165_n)
  );


  FA
  g_g166_n
  (
    .dout(g166_n),
    .din1(g161_p),
    .din2(g165_p)
  );


  LA
  g_g167_p
  (
    .dout(g167_p),
    .din1(g149_n_spl_0),
    .din2(g166_p)
  );


  FA
  g_g167_n
  (
    .dout(g167_n),
    .din1(g149_p_spl_0),
    .din2(g166_n)
  );


  FA
  g_g168_n
  (
    .dout(g168_n),
    .din1(G54_n_spl_00),
    .din2(g167_p_spl_0)
  );


  FA
  g_g169_n
  (
    .dout(g169_n),
    .din1(G8_n_spl_1),
    .din2(g83_n_spl_)
  );


  FA
  g_g170_n
  (
    .dout(g170_n),
    .din1(G13_n),
    .din2(g86_n_spl_)
  );


  FA
  g_g171_n
  (
    .dout(g171_n),
    .din1(G14_n),
    .din2(g170_n)
  );


  FA
  g_g172_n
  (
    .dout(g172_n),
    .din1(g169_n),
    .din2(g171_n)
  );


  FA
  g_g173_n
  (
    .dout(g173_n),
    .din1(G48_n_spl_0),
    .din2(g172_n_spl_00)
  );


  LA
  g_g174_p
  (
    .dout(g174_p),
    .din1(G48_p_spl_1),
    .din2(g167_n_spl_)
  );


  FA
  g_g174_n
  (
    .dout(g174_n),
    .din1(G48_n_spl_1),
    .din2(g167_p_spl_0)
  );


  LA
  g_g175_p
  (
    .dout(g175_p),
    .din1(G53_n_spl_00),
    .din2(g174_p_spl_)
  );


  LA
  g_g176_p
  (
    .dout(g176_p),
    .din1(G48_n_spl_1),
    .din2(g167_p_spl_)
  );


  FA
  g_g176_n
  (
    .dout(g176_n),
    .din1(G48_p_spl_1),
    .din2(g167_n_spl_)
  );


  FA
  g_g177_n
  (
    .dout(g177_n),
    .din1(g175_p),
    .din2(g176_p_spl_)
  );


  FA
  g_g178_n
  (
    .dout(g178_n),
    .din1(G51_n_spl_000),
    .din2(G58_n_spl_)
  );


  LA
  g_g179_p
  (
    .dout(g179_p),
    .din1(g177_n),
    .din2(g178_n)
  );


  LA
  g_g180_p
  (
    .dout(g180_p),
    .din1(G58_p),
    .din2(g176_n)
  );


  FA
  g_g180_n
  (
    .dout(g180_n),
    .din1(G58_n_spl_),
    .din2(g176_p_spl_)
  );


  FA
  g_g181_n
  (
    .dout(g181_n),
    .din1(G51_n_spl_000),
    .din2(g180_p_spl_)
  );


  LA
  g_g182_p
  (
    .dout(g182_p),
    .din1(G52_n_spl_00),
    .din2(g181_n)
  );


  LA
  g_g183_p
  (
    .dout(g183_p),
    .din1(g174_n_spl_),
    .din2(g182_p)
  );


  FA
  g_g184_n
  (
    .dout(g184_n),
    .din1(g179_p),
    .din2(g183_p)
  );


  LA
  g_g185_p
  (
    .dout(g185_p),
    .din1(g173_n),
    .din2(g184_n)
  );


  LA
  g_g186_p
  (
    .dout(g186_p),
    .din1(g168_n),
    .din2(g185_p)
  );


  LA
  g_g187_p
  (
    .dout(g187_p),
    .din1(g145_n),
    .din2(g186_p)
  );


  LA
  g_g188_p
  (
    .dout(g188_p),
    .din1(g144_n),
    .din2(g187_p)
  );


  FA
  g_g189_n
  (
    .dout(g189_n),
    .din1(G27_n_spl_1),
    .din2(G50_n_spl_00)
  );


  FA
  g_g190_n
  (
    .dout(g190_n),
    .din1(G45_n_spl_0),
    .din2(g172_n_spl_00)
  );


  LA
  g_g191_p
  (
    .dout(g191_p),
    .din1(G28_p_spl_),
    .din2(g160_n_spl_00)
  );


  FA
  g_g191_n
  (
    .dout(g191_n),
    .din1(G28_n_spl_1),
    .din2(g160_p_spl_00)
  );


  LA
  g_g192_p
  (
    .dout(g192_p),
    .din1(G35_p_spl_),
    .din2(g164_n_spl_0)
  );


  FA
  g_g192_n
  (
    .dout(g192_n),
    .din1(G35_n_spl_),
    .din2(g164_p_spl_0)
  );


  LA
  g_g193_p
  (
    .dout(g193_p),
    .din1(g191_n),
    .din2(g192_n)
  );


  FA
  g_g193_n
  (
    .dout(g193_n),
    .din1(g191_p),
    .din2(g192_p)
  );


  LA
  g_g194_p
  (
    .dout(g194_p),
    .din1(g149_n_spl_0),
    .din2(g193_p)
  );


  FA
  g_g194_n
  (
    .dout(g194_n),
    .din1(g149_p_spl_0),
    .din2(g193_n)
  );


  FA
  g_g195_n
  (
    .dout(g195_n),
    .din1(G54_n_spl_00),
    .din2(g194_p_spl_0)
  );


  LA
  g_g196_p
  (
    .dout(g196_p),
    .din1(G29_p_spl_),
    .din2(g160_n_spl_01)
  );


  FA
  g_g196_n
  (
    .dout(g196_n),
    .din1(G29_n_spl_1),
    .din2(g160_p_spl_01)
  );


  LA
  g_g197_p
  (
    .dout(g197_p),
    .din1(G36_p_spl_),
    .din2(g164_n_spl_1)
  );


  FA
  g_g197_n
  (
    .dout(g197_n),
    .din1(G36_n_spl_),
    .din2(g164_p_spl_1)
  );


  LA
  g_g198_p
  (
    .dout(g198_p),
    .din1(g196_n),
    .din2(g197_n)
  );


  FA
  g_g198_n
  (
    .dout(g198_n),
    .din1(g196_p),
    .din2(g197_p)
  );


  LA
  g_g199_p
  (
    .dout(g199_p),
    .din1(g149_n_spl_1),
    .din2(g198_p)
  );


  FA
  g_g199_n
  (
    .dout(g199_n),
    .din1(g149_p_spl_1),
    .din2(g198_n)
  );


  LA
  g_g200_p
  (
    .dout(g200_p),
    .din1(G46_p_spl_1),
    .din2(g199_n_spl_)
  );


  FA
  g_g200_n
  (
    .dout(g200_n),
    .din1(G46_n_spl_0),
    .din2(g199_p_spl_0)
  );


  LA
  g_g201_p
  (
    .dout(g201_p),
    .din1(G46_n_spl_1),
    .din2(g199_p_spl_0)
  );


  FA
  g_g201_n
  (
    .dout(g201_n),
    .din1(G46_p_spl_1),
    .din2(g199_n_spl_)
  );


  LA
  g_g202_p
  (
    .dout(g202_p),
    .din1(G30_p_spl_),
    .din2(g160_n_spl_01)
  );


  FA
  g_g202_n
  (
    .dout(g202_n),
    .din1(G30_n_spl_1),
    .din2(g160_p_spl_01)
  );


  LA
  g_g203_p
  (
    .dout(g203_p),
    .din1(G37_p_spl_),
    .din2(g164_n_spl_1)
  );


  FA
  g_g203_n
  (
    .dout(g203_n),
    .din1(G37_n_spl_),
    .din2(g164_p_spl_1)
  );


  LA
  g_g204_p
  (
    .dout(g204_p),
    .din1(g202_n),
    .din2(g203_n)
  );


  FA
  g_g204_n
  (
    .dout(g204_n),
    .din1(g202_p),
    .din2(g203_p)
  );


  LA
  g_g205_p
  (
    .dout(g205_p),
    .din1(g149_n_spl_1),
    .din2(g204_p)
  );


  FA
  g_g205_n
  (
    .dout(g205_n),
    .din1(g149_p_spl_1),
    .din2(g204_n)
  );


  LA
  g_g206_p
  (
    .dout(g206_p),
    .din1(G47_p_spl_1),
    .din2(g205_n_spl_)
  );


  FA
  g_g206_n
  (
    .dout(g206_n),
    .din1(G47_n_spl_0),
    .din2(g205_p_spl_0)
  );


  LA
  g_g207_p
  (
    .dout(g207_p),
    .din1(G47_n_spl_1),
    .din2(g205_p_spl_0)
  );


  FA
  g_g207_n
  (
    .dout(g207_n),
    .din1(G47_p_spl_1),
    .din2(g205_n_spl_)
  );


  LA
  g_g208_p
  (
    .dout(g208_p),
    .din1(g174_n_spl_),
    .din2(g180_n)
  );


  FA
  g_g208_n
  (
    .dout(g208_n),
    .din1(g174_p_spl_),
    .din2(g180_p_spl_)
  );


  LA
  g_g209_p
  (
    .dout(g209_p),
    .din1(g207_n),
    .din2(g208_n)
  );


  FA
  g_g209_n
  (
    .dout(g209_n),
    .din1(g207_p_spl_),
    .din2(g208_p_spl_)
  );


  LA
  g_g210_p
  (
    .dout(g210_p),
    .din1(g206_n_spl_),
    .din2(g209_n)
  );


  FA
  g_g210_n
  (
    .dout(g210_n),
    .din1(g206_p_spl_),
    .din2(g209_p_spl_)
  );


  LA
  g_g211_p
  (
    .dout(g211_p),
    .din1(g201_n),
    .din2(g210_n)
  );


  FA
  g_g211_n
  (
    .dout(g211_n),
    .din1(g201_p_spl_),
    .din2(g210_p_spl_)
  );


  LA
  g_g212_p
  (
    .dout(g212_p),
    .din1(g200_n_spl_),
    .din2(g211_n)
  );


  FA
  g_g212_n
  (
    .dout(g212_n),
    .din1(g200_p_spl_),
    .din2(g211_p_spl_)
  );


  FA
  g_g213_n
  (
    .dout(g213_n),
    .din1(G51_n_spl_001),
    .din2(g212_p_spl_)
  );


  LA
  g_g214_p
  (
    .dout(g214_p),
    .din1(G45_p_spl_1),
    .din2(g194_n_spl_)
  );


  FA
  g_g214_n
  (
    .dout(g214_n),
    .din1(G45_n_spl_1),
    .din2(g194_p_spl_0)
  );


  LA
  g_g215_p
  (
    .dout(g215_p),
    .din1(G53_n_spl_00),
    .din2(g214_p_spl_)
  );


  LA
  g_g216_p
  (
    .dout(g216_p),
    .din1(G45_n_spl_1),
    .din2(g194_p_spl_)
  );


  FA
  g_g216_n
  (
    .dout(g216_n),
    .din1(G45_p_spl_1),
    .din2(g194_n_spl_)
  );


  FA
  g_g217_n
  (
    .dout(g217_n),
    .din1(g215_p),
    .din2(g216_p_spl_)
  );


  LA
  g_g218_p
  (
    .dout(g218_p),
    .din1(g213_n),
    .din2(g217_n)
  );


  LA
  g_g219_p
  (
    .dout(g219_p),
    .din1(g212_n),
    .din2(g216_n)
  );


  FA
  g_g219_n
  (
    .dout(g219_n),
    .din1(g212_p_spl_),
    .din2(g216_p_spl_)
  );


  FA
  g_g220_n
  (
    .dout(g220_n),
    .din1(G51_n_spl_001),
    .din2(g219_p_spl_)
  );


  LA
  g_g221_p
  (
    .dout(g221_p),
    .din1(G52_n_spl_00),
    .din2(g220_n)
  );


  LA
  g_g222_p
  (
    .dout(g222_p),
    .din1(g214_n_spl_),
    .din2(g221_p)
  );


  FA
  g_g223_n
  (
    .dout(g223_n),
    .din1(g218_p),
    .din2(g222_p)
  );


  LA
  g_g224_p
  (
    .dout(g224_p),
    .din1(g195_n),
    .din2(g223_n)
  );


  LA
  g_g225_p
  (
    .dout(g225_p),
    .din1(g190_n),
    .din2(g224_p)
  );


  LA
  g_g226_p
  (
    .dout(g226_p),
    .din1(g189_n),
    .din2(g225_p)
  );


  FA
  g_g227_n
  (
    .dout(g227_n),
    .din1(G46_n_spl_1),
    .din2(g172_n_spl_01)
  );


  FA
  g_g228_n
  (
    .dout(g228_n),
    .din1(G55_n_spl_0),
    .din2(G56_n)
  );


  FA
  g_g229_n
  (
    .dout(g229_n),
    .din1(G28_n_spl_1),
    .din2(G50_n_spl_01)
  );


  FA
  g_g230_n
  (
    .dout(g230_n),
    .din1(G54_n_spl_01),
    .din2(g199_p_spl_)
  );


  LA
  g_g231_p
  (
    .dout(g231_p),
    .din1(G53_n_spl_01),
    .din2(g200_p_spl_)
  );


  FA
  g_g232_n
  (
    .dout(g232_n),
    .din1(g201_p_spl_),
    .din2(g231_p)
  );


  FA
  g_g233_n
  (
    .dout(g233_n),
    .din1(G51_n_spl_010),
    .din2(g210_p_spl_)
  );


  LA
  g_g234_p
  (
    .dout(g234_p),
    .din1(g232_n),
    .din2(g233_n)
  );


  FA
  g_g235_n
  (
    .dout(g235_n),
    .din1(G51_n_spl_010),
    .din2(g211_p_spl_)
  );


  LA
  g_g236_p
  (
    .dout(g236_p),
    .din1(G52_n_spl_01),
    .din2(g235_n)
  );


  LA
  g_g237_p
  (
    .dout(g237_p),
    .din1(g200_n_spl_),
    .din2(g236_p)
  );


  FA
  g_g238_n
  (
    .dout(g238_n),
    .din1(g234_p),
    .din2(g237_p)
  );


  LA
  g_g239_p
  (
    .dout(g239_p),
    .din1(g230_n),
    .din2(g238_n)
  );


  LA
  g_g240_p
  (
    .dout(g240_p),
    .din1(g229_n),
    .din2(g239_p)
  );


  LA
  g_g241_p
  (
    .dout(g241_p),
    .din1(g228_n),
    .din2(g240_p)
  );


  LA
  g_g242_p
  (
    .dout(g242_p),
    .din1(g227_n),
    .din2(g241_p)
  );


  FA
  g_g243_n
  (
    .dout(g243_n),
    .din1(G55_n_spl_),
    .din2(G57_n)
  );


  FA
  g_g244_n
  (
    .dout(g244_n),
    .din1(G29_n_spl_1),
    .din2(G50_n_spl_01)
  );


  FA
  g_g245_n
  (
    .dout(g245_n),
    .din1(G54_n_spl_01),
    .din2(g205_p_spl_)
  );


  FA
  g_g246_n
  (
    .dout(g246_n),
    .din1(G47_n_spl_1),
    .din2(g172_n_spl_01)
  );


  LA
  g_g247_p
  (
    .dout(g247_p),
    .din1(G53_n_spl_01),
    .din2(g206_p_spl_)
  );


  FA
  g_g248_n
  (
    .dout(g248_n),
    .din1(g207_p_spl_),
    .din2(g247_p)
  );


  FA
  g_g249_n
  (
    .dout(g249_n),
    .din1(G51_n_spl_011),
    .din2(g208_p_spl_)
  );


  LA
  g_g250_p
  (
    .dout(g250_p),
    .din1(g248_n),
    .din2(g249_n)
  );


  FA
  g_g251_n
  (
    .dout(g251_n),
    .din1(G51_n_spl_011),
    .din2(g209_p_spl_)
  );


  LA
  g_g252_p
  (
    .dout(g252_p),
    .din1(G52_n_spl_01),
    .din2(g251_n)
  );


  LA
  g_g253_p
  (
    .dout(g253_p),
    .din1(g206_n_spl_),
    .din2(g252_p)
  );


  FA
  g_g254_n
  (
    .dout(g254_n),
    .din1(g250_p),
    .din2(g253_p)
  );


  LA
  g_g255_p
  (
    .dout(g255_p),
    .din1(g246_n),
    .din2(g254_n)
  );


  LA
  g_g256_p
  (
    .dout(g256_p),
    .din1(g245_n),
    .din2(g255_p)
  );


  LA
  g_g257_p
  (
    .dout(g257_p),
    .din1(g244_n),
    .din2(g256_p)
  );


  LA
  g_g258_p
  (
    .dout(g258_p),
    .din1(g243_n),
    .din2(g257_p)
  );


  LA
  g_g259_p
  (
    .dout(g259_p),
    .din1(G10_p_spl_),
    .din2(g162_p_spl_)
  );


  FA
  g_g259_n
  (
    .dout(g259_n),
    .din1(G10_n_spl_),
    .din2(g162_n_spl_)
  );


  LA
  g_g260_p
  (
    .dout(g260_p),
    .din1(G35_p_spl_),
    .din2(g259_p_spl_0)
  );


  FA
  g_g260_n
  (
    .dout(g260_n),
    .din1(G35_n_spl_),
    .din2(g259_n_spl_0)
  );


  LA
  g_g261_p
  (
    .dout(g261_p),
    .din1(G2_p_spl_),
    .din2(G34_p_spl_0)
  );


  FA
  g_g261_n
  (
    .dout(g261_n),
    .din1(G2_n_spl_),
    .din2(G34_n_spl_0)
  );


  LA
  g_g262_p
  (
    .dout(g262_p),
    .din1(g260_n),
    .din2(g261_n)
  );


  FA
  g_g262_n
  (
    .dout(g262_n),
    .din1(g260_p),
    .din2(g261_p)
  );


  LA
  g_g263_p
  (
    .dout(g263_p),
    .din1(G24_p_spl_),
    .din2(g160_n_spl_10)
  );


  FA
  g_g263_n
  (
    .dout(g263_n),
    .din1(G24_n_spl_1),
    .din2(g160_p_spl_10)
  );


  LA
  g_g264_p
  (
    .dout(g264_p),
    .din1(G4_p_spl_10),
    .din2(g147_p_spl_)
  );


  FA
  g_g264_n
  (
    .dout(g264_n),
    .din1(G4_n_spl_11),
    .din2(g147_n_spl_)
  );


  LA
  g_g265_p
  (
    .dout(g265_p),
    .din1(G60_n_spl_0),
    .din2(g264_p)
  );


  FA
  g_g265_n
  (
    .dout(g265_n),
    .din1(G60_p_spl_),
    .din2(g264_n)
  );


  LA
  g_g266_p
  (
    .dout(g266_p),
    .din1(g263_n),
    .din2(g265_n_spl_0)
  );


  FA
  g_g266_n
  (
    .dout(g266_n),
    .din1(g263_p),
    .din2(g265_p_spl_0)
  );


  LA
  g_g267_p
  (
    .dout(g267_p),
    .din1(g262_p),
    .din2(g266_p)
  );


  FA
  g_g267_n
  (
    .dout(g267_n),
    .din1(g262_n),
    .din2(g266_n)
  );


  LA
  g_g268_p
  (
    .dout(g268_p),
    .din1(G41_p_spl_1),
    .din2(g267_n_spl_)
  );


  FA
  g_g268_n
  (
    .dout(g268_n),
    .din1(G41_n_spl_0),
    .din2(g267_p_spl_0)
  );


  LA
  g_g269_p
  (
    .dout(g269_p),
    .din1(G36_p_spl_),
    .din2(g259_p_spl_0)
  );


  FA
  g_g269_n
  (
    .dout(g269_n),
    .din1(G36_n_spl_),
    .din2(g259_n_spl_0)
  );


  LA
  g_g270_p
  (
    .dout(g270_p),
    .din1(G9_p_spl_),
    .din2(G34_p_spl_0)
  );


  FA
  g_g270_n
  (
    .dout(g270_n),
    .din1(G9_n_spl_),
    .din2(G34_n_spl_0)
  );


  LA
  g_g271_p
  (
    .dout(g271_p),
    .din1(g269_n),
    .din2(g270_n)
  );


  FA
  g_g271_n
  (
    .dout(g271_n),
    .din1(g269_p),
    .din2(g270_p)
  );


  LA
  g_g272_p
  (
    .dout(g272_p),
    .din1(G25_p_spl_),
    .din2(g160_n_spl_10)
  );


  FA
  g_g272_n
  (
    .dout(g272_n),
    .din1(G25_n_spl_1),
    .din2(g160_p_spl_10)
  );


  LA
  g_g273_p
  (
    .dout(g273_p),
    .din1(g265_n_spl_0),
    .din2(g272_n)
  );


  FA
  g_g273_n
  (
    .dout(g273_n),
    .din1(g265_p_spl_0),
    .din2(g272_p)
  );


  LA
  g_g274_p
  (
    .dout(g274_p),
    .din1(g271_p),
    .din2(g273_p)
  );


  FA
  g_g274_n
  (
    .dout(g274_n),
    .din1(g271_n),
    .din2(g273_n)
  );


  LA
  g_g275_p
  (
    .dout(g275_p),
    .din1(G42_p_spl_1),
    .din2(g274_n_spl_)
  );


  FA
  g_g275_n
  (
    .dout(g275_n),
    .din1(G42_n_spl_0),
    .din2(g274_p_spl_0)
  );


  LA
  g_g276_p
  (
    .dout(g276_p),
    .din1(G42_n_spl_1),
    .din2(g274_p_spl_0)
  );


  FA
  g_g276_n
  (
    .dout(g276_n),
    .din1(G42_p_spl_1),
    .din2(g274_n_spl_)
  );


  LA
  g_g277_p
  (
    .dout(g277_p),
    .din1(G37_p_spl_),
    .din2(g259_p_spl_1)
  );


  FA
  g_g277_n
  (
    .dout(g277_n),
    .din1(G37_n_spl_),
    .din2(g259_n_spl_1)
  );


  LA
  g_g278_p
  (
    .dout(g278_p),
    .din1(G4_p_spl_1),
    .din2(G34_p_spl_1)
  );


  FA
  g_g278_n
  (
    .dout(g278_n),
    .din1(G4_n_spl_11),
    .din2(G34_n_spl_1)
  );


  LA
  g_g279_p
  (
    .dout(g279_p),
    .din1(g277_n),
    .din2(g278_n)
  );


  FA
  g_g279_n
  (
    .dout(g279_n),
    .din1(g277_p),
    .din2(g278_p)
  );


  LA
  g_g280_p
  (
    .dout(g280_p),
    .din1(G26_p_spl_),
    .din2(g160_n_spl_11)
  );


  FA
  g_g280_n
  (
    .dout(g280_n),
    .din1(G26_n_spl_1),
    .din2(g160_p_spl_11)
  );


  LA
  g_g281_p
  (
    .dout(g281_p),
    .din1(g265_n_spl_1),
    .din2(g280_n)
  );


  FA
  g_g281_n
  (
    .dout(g281_n),
    .din1(g265_p_spl_1),
    .din2(g280_p)
  );


  LA
  g_g282_p
  (
    .dout(g282_p),
    .din1(g279_p),
    .din2(g281_p)
  );


  FA
  g_g282_n
  (
    .dout(g282_n),
    .din1(g279_n),
    .din2(g281_n)
  );


  LA
  g_g283_p
  (
    .dout(g283_p),
    .din1(G43_p_spl_1),
    .din2(g282_n_spl_)
  );


  FA
  g_g283_n
  (
    .dout(g283_n),
    .din1(G43_n_spl_0),
    .din2(g282_p_spl_0)
  );


  LA
  g_g284_p
  (
    .dout(g284_p),
    .din1(G43_n_spl_1),
    .din2(g282_p_spl_0)
  );


  FA
  g_g284_n
  (
    .dout(g284_n),
    .din1(G43_p_spl_1),
    .din2(g282_n_spl_)
  );


  LA
  g_g285_p
  (
    .dout(g285_p),
    .din1(g214_n_spl_),
    .din2(g219_n)
  );


  FA
  g_g285_n
  (
    .dout(g285_n),
    .din1(g214_p_spl_),
    .din2(g219_p_spl_)
  );


  LA
  g_g286_p
  (
    .dout(g286_p),
    .din1(G39_p_spl_),
    .din2(g259_p_spl_1)
  );


  FA
  g_g286_n
  (
    .dout(g286_n),
    .din1(G39_n_spl_),
    .din2(g259_n_spl_1)
  );


  LA
  g_g287_p
  (
    .dout(g287_p),
    .din1(G34_p_spl_1),
    .din2(G38_p)
  );


  FA
  g_g287_n
  (
    .dout(g287_n),
    .din1(G34_n_spl_1),
    .din2(G38_n)
  );


  LA
  g_g288_p
  (
    .dout(g288_p),
    .din1(g286_n),
    .din2(g287_n)
  );


  FA
  g_g288_n
  (
    .dout(g288_n),
    .din1(g286_p),
    .din2(g287_p)
  );


  LA
  g_g289_p
  (
    .dout(g289_p),
    .din1(G27_p_spl_),
    .din2(g160_n_spl_11)
  );


  FA
  g_g289_n
  (
    .dout(g289_n),
    .din1(G27_n_spl_1),
    .din2(g160_p_spl_11)
  );


  LA
  g_g290_p
  (
    .dout(g290_p),
    .din1(g265_n_spl_1),
    .din2(g289_n)
  );


  FA
  g_g290_n
  (
    .dout(g290_n),
    .din1(g265_p_spl_1),
    .din2(g289_p)
  );


  LA
  g_g291_p
  (
    .dout(g291_p),
    .din1(g288_p),
    .din2(g290_p)
  );


  FA
  g_g291_n
  (
    .dout(g291_n),
    .din1(g288_n),
    .din2(g290_n)
  );


  LA
  g_g292_p
  (
    .dout(g292_p),
    .din1(G44_n_spl_0),
    .din2(g291_p_spl_0)
  );


  FA
  g_g292_n
  (
    .dout(g292_n),
    .din1(G44_p_spl_1),
    .din2(g291_n_spl_)
  );


  LA
  g_g293_p
  (
    .dout(g293_p),
    .din1(g285_n_spl_),
    .din2(g292_n_spl_)
  );


  FA
  g_g293_n
  (
    .dout(g293_n),
    .din1(g285_p_spl_),
    .din2(g292_p_spl_)
  );


  LA
  g_g294_p
  (
    .dout(g294_p),
    .din1(G44_p_spl_1),
    .din2(g291_n_spl_)
  );


  FA
  g_g294_n
  (
    .dout(g294_n),
    .din1(G44_n_spl_1),
    .din2(g291_p_spl_0)
  );


  LA
  g_g295_p
  (
    .dout(g295_p),
    .din1(g293_n),
    .din2(g294_n_spl_0)
  );


  FA
  g_g295_n
  (
    .dout(g295_n),
    .din1(g293_p),
    .din2(g294_p_spl_)
  );


  LA
  g_g296_p
  (
    .dout(g296_p),
    .din1(g284_n_spl_),
    .din2(g295_n_spl_)
  );


  FA
  g_g296_n
  (
    .dout(g296_n),
    .din1(g284_p_spl_),
    .din2(g295_p_spl_)
  );


  LA
  g_g297_p
  (
    .dout(g297_p),
    .din1(g283_n_spl_0),
    .din2(g296_n)
  );


  FA
  g_g297_n
  (
    .dout(g297_n),
    .din1(g283_p_spl_),
    .din2(g296_p)
  );


  LA
  g_g298_p
  (
    .dout(g298_p),
    .din1(g276_n_spl_),
    .din2(g297_n_spl_)
  );


  FA
  g_g298_n
  (
    .dout(g298_n),
    .din1(g276_p_spl_),
    .din2(g297_p_spl_)
  );


  LA
  g_g299_p
  (
    .dout(g299_p),
    .din1(g275_n_spl_0),
    .din2(g298_n)
  );


  FA
  g_g299_n
  (
    .dout(g299_n),
    .din1(g275_p_spl_),
    .din2(g298_p)
  );


  LA
  g_g300_p
  (
    .dout(g300_p),
    .din1(G41_n_spl_1),
    .din2(g267_p_spl_0)
  );


  FA
  g_g300_n
  (
    .dout(g300_n),
    .din1(G41_p_spl_1),
    .din2(g267_n_spl_)
  );


  FA
  g_g301_n
  (
    .dout(g301_n),
    .din1(g299_p_spl_),
    .din2(g300_p_spl_)
  );


  LA
  g_g302_p
  (
    .dout(g302_p),
    .din1(g268_n_spl_0),
    .din2(g301_n)
  );


  LA
  g_g303_p
  (
    .dout(g303_p),
    .din1(g292_n_spl_),
    .din2(g294_n_spl_0)
  );


  FA
  g_g303_n
  (
    .dout(g303_n),
    .din1(g292_p_spl_),
    .din2(g294_p_spl_)
  );


  FA
  g_g304_n
  (
    .dout(g304_n),
    .din1(g285_p_spl_),
    .din2(g303_p)
  );


  FA
  g_g305_n
  (
    .dout(g305_n),
    .din1(g285_n_spl_),
    .din2(g303_n_spl_)
  );


  LA
  g_g306_p
  (
    .dout(g306_p),
    .din1(g304_n),
    .din2(g305_n)
  );


  FA
  g_g307_n
  (
    .dout(g307_n),
    .din1(G51_n_spl_10),
    .din2(g306_p)
  );


  FA
  g_g308_n
  (
    .dout(g308_n),
    .din1(G52_n_spl_10),
    .din2(g303_n_spl_)
  );


  FA
  g_g309_n
  (
    .dout(g309_n),
    .din1(G54_n_spl_10),
    .din2(g291_p_spl_)
  );


  LA
  g_g310_p
  (
    .dout(g310_p),
    .din1(g308_n),
    .din2(g309_n)
  );


  FA
  g_g311_n
  (
    .dout(g311_n),
    .din1(G44_n_spl_1),
    .din2(g172_n_spl_10)
  );


  FA
  g_g312_n
  (
    .dout(g312_n),
    .din1(G53_n_spl_10),
    .din2(g294_n_spl_)
  );


  FA
  g_g313_n
  (
    .dout(g313_n),
    .din1(G26_n_spl_1),
    .din2(G50_n_spl_10)
  );


  LA
  g_g314_p
  (
    .dout(g314_p),
    .din1(g312_n),
    .din2(g313_n)
  );


  LA
  g_g315_p
  (
    .dout(g315_p),
    .din1(g311_n),
    .din2(g314_p)
  );


  LA
  g_g316_p
  (
    .dout(g316_p),
    .din1(g310_p),
    .din2(g315_p)
  );


  LA
  g_g317_p
  (
    .dout(g317_p),
    .din1(g307_n),
    .din2(g316_p)
  );


  FA
  g_g318_n
  (
    .dout(g318_n),
    .din1(G53_n_spl_10),
    .din2(g268_n_spl_0)
  );


  FA
  g_g319_n
  (
    .dout(g319_n),
    .din1(G50_n_spl_10),
    .din2(G60_n_spl_)
  );


  LA
  g_g320_p
  (
    .dout(g320_p),
    .din1(g318_n),
    .din2(g319_n)
  );


  FA
  g_g321_n
  (
    .dout(g321_n),
    .din1(G41_n_spl_1),
    .din2(g172_n_spl_10)
  );


  LA
  g_g322_p
  (
    .dout(g322_p),
    .din1(g268_n_spl_),
    .din2(g300_n)
  );


  FA
  g_g322_n
  (
    .dout(g322_n),
    .din1(g268_p),
    .din2(g300_p_spl_)
  );


  FA
  g_g323_n
  (
    .dout(g323_n),
    .din1(G52_n_spl_10),
    .din2(g322_n_spl_)
  );


  FA
  g_g324_n
  (
    .dout(g324_n),
    .din1(G54_n_spl_10),
    .din2(g267_p_spl_)
  );


  LA
  g_g325_p
  (
    .dout(g325_p),
    .din1(g323_n),
    .din2(g324_n)
  );


  LA
  g_g326_p
  (
    .dout(g326_p),
    .din1(g321_n),
    .din2(g325_p)
  );


  LA
  g_g327_p
  (
    .dout(g327_p),
    .din1(g320_p),
    .din2(g326_p)
  );


  LA
  g_g328_p
  (
    .dout(g328_p),
    .din1(g299_p_spl_),
    .din2(g322_n_spl_)
  );


  LA
  g_g329_p
  (
    .dout(g329_p),
    .din1(g299_n),
    .din2(g322_p)
  );


  FA
  g_g330_n
  (
    .dout(g330_n),
    .din1(G51_n_spl_10),
    .din2(g329_p)
  );


  FA
  g_g331_n
  (
    .dout(g331_n),
    .din1(g328_p),
    .din2(g330_n)
  );


  LA
  g_g332_p
  (
    .dout(g332_p),
    .din1(g327_p),
    .din2(g331_n)
  );


  FA
  g_g333_n
  (
    .dout(g333_n),
    .din1(G53_n_spl_11),
    .din2(g275_n_spl_0)
  );


  FA
  g_g334_n
  (
    .dout(g334_n),
    .din1(G24_n_spl_1),
    .din2(G50_n_spl_11)
  );


  LA
  g_g335_p
  (
    .dout(g335_p),
    .din1(g333_n),
    .din2(g334_n)
  );


  FA
  g_g336_n
  (
    .dout(g336_n),
    .din1(G42_n_spl_1),
    .din2(g172_n_spl_11)
  );


  LA
  g_g337_p
  (
    .dout(g337_p),
    .din1(g275_n_spl_),
    .din2(g276_n_spl_)
  );


  FA
  g_g337_n
  (
    .dout(g337_n),
    .din1(g275_p_spl_),
    .din2(g276_p_spl_)
  );


  FA
  g_g338_n
  (
    .dout(g338_n),
    .din1(G52_n_spl_11),
    .din2(g337_n_spl_)
  );


  FA
  g_g339_n
  (
    .dout(g339_n),
    .din1(G54_n_spl_11),
    .din2(g274_p_spl_)
  );


  LA
  g_g340_p
  (
    .dout(g340_p),
    .din1(g338_n),
    .din2(g339_n)
  );


  LA
  g_g341_p
  (
    .dout(g341_p),
    .din1(g336_n),
    .din2(g340_p)
  );


  LA
  g_g342_p
  (
    .dout(g342_p),
    .din1(g335_p),
    .din2(g341_p)
  );


  LA
  g_g343_p
  (
    .dout(g343_p),
    .din1(g297_p_spl_),
    .din2(g337_n_spl_)
  );


  LA
  g_g344_p
  (
    .dout(g344_p),
    .din1(g297_n_spl_),
    .din2(g337_p)
  );


  FA
  g_g345_n
  (
    .dout(g345_n),
    .din1(G51_n_spl_11),
    .din2(g344_p)
  );


  FA
  g_g346_n
  (
    .dout(g346_n),
    .din1(g343_p),
    .din2(g345_n)
  );


  LA
  g_g347_p
  (
    .dout(g347_p),
    .din1(g342_p),
    .din2(g346_n)
  );


  FA
  g_g348_n
  (
    .dout(g348_n),
    .din1(G53_n_spl_11),
    .din2(g283_n_spl_0)
  );


  FA
  g_g349_n
  (
    .dout(g349_n),
    .din1(G25_n_spl_1),
    .din2(G50_n_spl_11)
  );


  LA
  g_g350_p
  (
    .dout(g350_p),
    .din1(g348_n),
    .din2(g349_n)
  );


  FA
  g_g351_n
  (
    .dout(g351_n),
    .din1(G43_n_spl_1),
    .din2(g172_n_spl_11)
  );


  LA
  g_g352_p
  (
    .dout(g352_p),
    .din1(g283_n_spl_),
    .din2(g284_n_spl_)
  );


  FA
  g_g352_n
  (
    .dout(g352_n),
    .din1(g283_p_spl_),
    .din2(g284_p_spl_)
  );


  FA
  g_g353_n
  (
    .dout(g353_n),
    .din1(G52_n_spl_11),
    .din2(g352_n_spl_)
  );


  FA
  g_g354_n
  (
    .dout(g354_n),
    .din1(G54_n_spl_11),
    .din2(g282_p_spl_)
  );


  LA
  g_g355_p
  (
    .dout(g355_p),
    .din1(g353_n),
    .din2(g354_n)
  );


  LA
  g_g356_p
  (
    .dout(g356_p),
    .din1(g351_n),
    .din2(g355_p)
  );


  LA
  g_g357_p
  (
    .dout(g357_p),
    .din1(g295_p_spl_),
    .din2(g352_n_spl_)
  );


  LA
  g_g358_p
  (
    .dout(g358_p),
    .din1(g295_n_spl_),
    .din2(g352_p)
  );


  FA
  g_g359_n
  (
    .dout(g359_n),
    .din1(G51_n_spl_11),
    .din2(g358_p)
  );


  FA
  g_g360_n
  (
    .dout(g360_n),
    .din1(g357_p),
    .din2(g359_n)
  );


  LA
  g_g361_p
  (
    .dout(g361_p),
    .din1(g356_p),
    .din2(g360_n)
  );


  LA
  g_g362_p
  (
    .dout(g362_p),
    .din1(g350_p),
    .din2(g361_p)
  );


  buf

  (
    G855_p,
    g62_n
  );


  buf

  (
    G856_p,
    g64_n
  );


  buf

  (
    G857_p,
    g65_n_spl_
  );


  buf

  (
    G858_p,
    g66_n
  );


  buf

  (
    G859_p,
    g69_n
  );


  buf

  (
    G860_p,
    g73_p
  );


  buf

  (
    G861_p,
    g75_p
  );


  buf

  (
    G862_n,
    g77_n
  );


  buf

  (
    G863_n,
    g78_n
  );


  buf

  (
    G864_n,
    g80_p
  );


  buf

  (
    G865_n,
    g81_n
  );


  buf

  (
    G866_p,
    g82_n_spl_1
  );


  buf

  (
    G867_p,
    g85_n
  );


  buf

  (
    G868_p,
    g88_n
  );


  buf

  (
    G869_n,
    g89_p
  );


  buf

  (
    G870_p,
    g116_n
  );


  buf

  (
    G871_p,
    g143_n
  );


  buf

  (
    G872_p,
    g188_p
  );


  buf

  (
    G873_p,
    g226_p
  );


  buf

  (
    G874_p,
    g242_p
  );


  buf

  (
    G875_p,
    g258_p
  );


  buf

  (
    G876_p,
    g302_p
  );


  buf

  (
    G877_p,
    g317_p
  );


  buf

  (
    G878_p,
    g332_p
  );


  buf

  (
    G879_p,
    g347_p
  );


  buf

  (
    G880_p,
    g362_p
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    G6_n_spl_,
    G6_n
  );


  buf

  (
    G6_n_spl_0,
    G6_n_spl_
  );


  buf

  (
    G16_n_spl_,
    G16_n
  );


  buf

  (
    G8_n_spl_,
    G8_n
  );


  buf

  (
    G8_n_spl_0,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_00,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_01,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_1,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_10,
    G8_n_spl_1
  );


  buf

  (
    g61_n_spl_,
    g61_n
  );


  buf

  (
    G7_n_spl_,
    G7_n
  );


  buf

  (
    G17_n_spl_,
    G17_n
  );


  buf

  (
    G17_n_spl_0,
    G17_n_spl_
  );


  buf

  (
    g63_n_spl_,
    g63_n
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G1_p_spl_0,
    G1_p_spl_
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G1_n_spl_0,
    G1_n_spl_
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G3_n_spl_,
    G3_n
  );


  buf

  (
    g67_n_spl_,
    g67_n
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    G4_n_spl_0,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_00,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_01,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_1,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_10,
    G4_n_spl_1
  );


  buf

  (
    G4_n_spl_11,
    G4_n_spl_1
  );


  buf

  (
    g68_n_spl_,
    g68_n
  );


  buf

  (
    g70_p_spl_,
    g70_p
  );


  buf

  (
    g70_n_spl_,
    g70_n
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_00,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_01,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_10,
    G4_p_spl_1
  );


  buf

  (
    g65_n_spl_,
    g65_n
  );


  buf

  (
    g65_n_spl_0,
    g65_n_spl_
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    G11_n_spl_,
    G11_n
  );


  buf

  (
    G11_n_spl_0,
    G11_n_spl_
  );


  buf

  (
    G11_n_spl_1,
    G11_n_spl_
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


  buf

  (
    g74_p_spl_,
    g74_p
  );


  buf

  (
    g76_n_spl_,
    g76_n
  );


  buf

  (
    g79_n_spl_,
    g79_n
  );


  buf

  (
    G9_p_spl_,
    G9_p
  );


  buf

  (
    G9_p_spl_0,
    G9_p_spl_
  );


  buf

  (
    G9_n_spl_,
    G9_n
  );


  buf

  (
    G9_n_spl_0,
    G9_n_spl_
  );


  buf

  (
    G10_n_spl_,
    G10_n
  );


  buf

  (
    G10_n_spl_0,
    G10_n_spl_
  );


  buf

  (
    g83_n_spl_,
    g83_n
  );


  buf

  (
    g83_n_spl_0,
    g83_n_spl_
  );


  buf

  (
    G12_n_spl_,
    G12_n
  );


  buf

  (
    g86_n_spl_,
    g86_n
  );


  buf

  (
    G24_p_spl_,
    G24_p
  );


  buf

  (
    G24_p_spl_0,
    G24_p_spl_
  );


  buf

  (
    G25_n_spl_,
    G25_n
  );


  buf

  (
    G25_n_spl_0,
    G25_n_spl_
  );


  buf

  (
    G25_n_spl_1,
    G25_n_spl_
  );


  buf

  (
    G24_n_spl_,
    G24_n
  );


  buf

  (
    G24_n_spl_0,
    G24_n_spl_
  );


  buf

  (
    G24_n_spl_1,
    G24_n_spl_
  );


  buf

  (
    G25_p_spl_,
    G25_p
  );


  buf

  (
    G25_p_spl_0,
    G25_p_spl_
  );


  buf

  (
    G26_p_spl_,
    G26_p
  );


  buf

  (
    G26_p_spl_0,
    G26_p_spl_
  );


  buf

  (
    G27_n_spl_,
    G27_n
  );


  buf

  (
    G27_n_spl_0,
    G27_n_spl_
  );


  buf

  (
    G27_n_spl_1,
    G27_n_spl_
  );


  buf

  (
    G26_n_spl_,
    G26_n
  );


  buf

  (
    G26_n_spl_0,
    G26_n_spl_
  );


  buf

  (
    G26_n_spl_1,
    G26_n_spl_
  );


  buf

  (
    G27_p_spl_,
    G27_p
  );


  buf

  (
    G27_p_spl_0,
    G27_p_spl_
  );


  buf

  (
    g92_p_spl_,
    g92_p
  );


  buf

  (
    g95_p_spl_,
    g95_p
  );


  buf

  (
    g92_n_spl_,
    g92_n
  );


  buf

  (
    g95_n_spl_,
    g95_n
  );


  buf

  (
    G32_p_spl_,
    G32_p
  );


  buf

  (
    G32_p_spl_0,
    G32_p_spl_
  );


  buf

  (
    G32_p_spl_1,
    G32_p_spl_
  );


  buf

  (
    g98_p_spl_,
    g98_p
  );


  buf

  (
    G32_n_spl_,
    G32_n
  );


  buf

  (
    G32_n_spl_0,
    G32_n_spl_
  );


  buf

  (
    G32_n_spl_1,
    G32_n_spl_
  );


  buf

  (
    g98_n_spl_,
    g98_n
  );


  buf

  (
    G28_p_spl_,
    G28_p
  );


  buf

  (
    G28_p_spl_0,
    G28_p_spl_
  );


  buf

  (
    G29_n_spl_,
    G29_n
  );


  buf

  (
    G29_n_spl_0,
    G29_n_spl_
  );


  buf

  (
    G29_n_spl_1,
    G29_n_spl_
  );


  buf

  (
    G28_n_spl_,
    G28_n
  );


  buf

  (
    G28_n_spl_0,
    G28_n_spl_
  );


  buf

  (
    G28_n_spl_1,
    G28_n_spl_
  );


  buf

  (
    G29_p_spl_,
    G29_p
  );


  buf

  (
    G29_p_spl_0,
    G29_p_spl_
  );


  buf

  (
    G30_p_spl_,
    G30_p
  );


  buf

  (
    G30_p_spl_0,
    G30_p_spl_
  );


  buf

  (
    G31_n_spl_,
    G31_n
  );


  buf

  (
    G31_n_spl_0,
    G31_n_spl_
  );


  buf

  (
    G30_n_spl_,
    G30_n
  );


  buf

  (
    G30_n_spl_0,
    G30_n_spl_
  );


  buf

  (
    G30_n_spl_1,
    G30_n_spl_
  );


  buf

  (
    G31_p_spl_,
    G31_p
  );


  buf

  (
    G31_p_spl_0,
    G31_p_spl_
  );


  buf

  (
    g104_p_spl_,
    g104_p
  );


  buf

  (
    g107_p_spl_,
    g107_p
  );


  buf

  (
    g104_n_spl_,
    g104_n
  );


  buf

  (
    g107_n_spl_,
    g107_n
  );


  buf

  (
    G33_p_spl_,
    G33_p
  );


  buf

  (
    g110_p_spl_,
    g110_p
  );


  buf

  (
    G33_n_spl_,
    G33_n
  );


  buf

  (
    g110_n_spl_,
    g110_n
  );


  buf

  (
    G41_p_spl_,
    G41_p
  );


  buf

  (
    G41_p_spl_0,
    G41_p_spl_
  );


  buf

  (
    G41_p_spl_1,
    G41_p_spl_
  );


  buf

  (
    G42_n_spl_,
    G42_n
  );


  buf

  (
    G42_n_spl_0,
    G42_n_spl_
  );


  buf

  (
    G42_n_spl_00,
    G42_n_spl_0
  );


  buf

  (
    G42_n_spl_1,
    G42_n_spl_
  );


  buf

  (
    G41_n_spl_,
    G41_n
  );


  buf

  (
    G41_n_spl_0,
    G41_n_spl_
  );


  buf

  (
    G41_n_spl_00,
    G41_n_spl_0
  );


  buf

  (
    G41_n_spl_1,
    G41_n_spl_
  );


  buf

  (
    G42_p_spl_,
    G42_p
  );


  buf

  (
    G42_p_spl_0,
    G42_p_spl_
  );


  buf

  (
    G42_p_spl_1,
    G42_p_spl_
  );


  buf

  (
    G43_p_spl_,
    G43_p
  );


  buf

  (
    G43_p_spl_0,
    G43_p_spl_
  );


  buf

  (
    G43_p_spl_1,
    G43_p_spl_
  );


  buf

  (
    G44_n_spl_,
    G44_n
  );


  buf

  (
    G44_n_spl_0,
    G44_n_spl_
  );


  buf

  (
    G44_n_spl_00,
    G44_n_spl_0
  );


  buf

  (
    G44_n_spl_1,
    G44_n_spl_
  );


  buf

  (
    G43_n_spl_,
    G43_n
  );


  buf

  (
    G43_n_spl_0,
    G43_n_spl_
  );


  buf

  (
    G43_n_spl_00,
    G43_n_spl_0
  );


  buf

  (
    G43_n_spl_1,
    G43_n_spl_
  );


  buf

  (
    G44_p_spl_,
    G44_p
  );


  buf

  (
    G44_p_spl_0,
    G44_p_spl_
  );


  buf

  (
    G44_p_spl_1,
    G44_p_spl_
  );


  buf

  (
    g119_p_spl_,
    g119_p
  );


  buf

  (
    g122_p_spl_,
    g122_p
  );


  buf

  (
    g119_n_spl_,
    g119_n
  );


  buf

  (
    g122_n_spl_,
    g122_n
  );


  buf

  (
    g125_p_spl_,
    g125_p
  );


  buf

  (
    g125_n_spl_,
    g125_n
  );


  buf

  (
    G45_p_spl_,
    G45_p
  );


  buf

  (
    G45_p_spl_0,
    G45_p_spl_
  );


  buf

  (
    G45_p_spl_1,
    G45_p_spl_
  );


  buf

  (
    G46_n_spl_,
    G46_n
  );


  buf

  (
    G46_n_spl_0,
    G46_n_spl_
  );


  buf

  (
    G46_n_spl_00,
    G46_n_spl_0
  );


  buf

  (
    G46_n_spl_1,
    G46_n_spl_
  );


  buf

  (
    G45_n_spl_,
    G45_n
  );


  buf

  (
    G45_n_spl_0,
    G45_n_spl_
  );


  buf

  (
    G45_n_spl_00,
    G45_n_spl_0
  );


  buf

  (
    G45_n_spl_1,
    G45_n_spl_
  );


  buf

  (
    G46_p_spl_,
    G46_p
  );


  buf

  (
    G46_p_spl_0,
    G46_p_spl_
  );


  buf

  (
    G46_p_spl_1,
    G46_p_spl_
  );


  buf

  (
    G47_p_spl_,
    G47_p
  );


  buf

  (
    G47_p_spl_0,
    G47_p_spl_
  );


  buf

  (
    G47_p_spl_1,
    G47_p_spl_
  );


  buf

  (
    G48_n_spl_,
    G48_n
  );


  buf

  (
    G48_n_spl_0,
    G48_n_spl_
  );


  buf

  (
    G48_n_spl_00,
    G48_n_spl_0
  );


  buf

  (
    G48_n_spl_1,
    G48_n_spl_
  );


  buf

  (
    G47_n_spl_,
    G47_n
  );


  buf

  (
    G47_n_spl_0,
    G47_n_spl_
  );


  buf

  (
    G47_n_spl_00,
    G47_n_spl_0
  );


  buf

  (
    G47_n_spl_1,
    G47_n_spl_
  );


  buf

  (
    G48_p_spl_,
    G48_p
  );


  buf

  (
    G48_p_spl_0,
    G48_p_spl_
  );


  buf

  (
    G48_p_spl_1,
    G48_p_spl_
  );


  buf

  (
    g131_p_spl_,
    g131_p
  );


  buf

  (
    g134_p_spl_,
    g134_p
  );


  buf

  (
    g131_n_spl_,
    g131_n
  );


  buf

  (
    g134_n_spl_,
    g134_n
  );


  buf

  (
    G49_p_spl_,
    G49_p
  );


  buf

  (
    g137_p_spl_,
    g137_p
  );


  buf

  (
    G49_n_spl_,
    G49_n
  );


  buf

  (
    g137_n_spl_,
    g137_n
  );


  buf

  (
    G55_n_spl_,
    G55_n
  );


  buf

  (
    G55_n_spl_0,
    G55_n_spl_
  );


  buf

  (
    G50_n_spl_,
    G50_n
  );


  buf

  (
    G50_n_spl_0,
    G50_n_spl_
  );


  buf

  (
    G50_n_spl_00,
    G50_n_spl_0
  );


  buf

  (
    G50_n_spl_01,
    G50_n_spl_0
  );


  buf

  (
    G50_n_spl_1,
    G50_n_spl_
  );


  buf

  (
    G50_n_spl_10,
    G50_n_spl_1
  );


  buf

  (
    G50_n_spl_11,
    G50_n_spl_1
  );


  buf

  (
    g82_p_spl_,
    g82_p
  );


  buf

  (
    g82_p_spl_0,
    g82_p_spl_
  );


  buf

  (
    g82_n_spl_,
    g82_n
  );


  buf

  (
    g82_n_spl_0,
    g82_n_spl_
  );


  buf

  (
    g82_n_spl_1,
    g82_n_spl_
  );


  buf

  (
    G10_p_spl_,
    G10_p
  );


  buf

  (
    g147_p_spl_,
    g147_p
  );


  buf

  (
    g147_n_spl_,
    g147_n
  );


  buf

  (
    G60_n_spl_,
    G60_n
  );


  buf

  (
    G60_n_spl_0,
    G60_n_spl_
  );


  buf

  (
    G60_p_spl_,
    G60_p
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    g153_p_spl_,
    g153_p
  );


  buf

  (
    g153_n_spl_,
    g153_n
  );


  buf

  (
    g160_n_spl_,
    g160_n
  );


  buf

  (
    g160_n_spl_0,
    g160_n_spl_
  );


  buf

  (
    g160_n_spl_00,
    g160_n_spl_0
  );


  buf

  (
    g160_n_spl_01,
    g160_n_spl_0
  );


  buf

  (
    g160_n_spl_1,
    g160_n_spl_
  );


  buf

  (
    g160_n_spl_10,
    g160_n_spl_1
  );


  buf

  (
    g160_n_spl_11,
    g160_n_spl_1
  );


  buf

  (
    g160_p_spl_,
    g160_p
  );


  buf

  (
    g160_p_spl_0,
    g160_p_spl_
  );


  buf

  (
    g160_p_spl_00,
    g160_p_spl_0
  );


  buf

  (
    g160_p_spl_01,
    g160_p_spl_0
  );


  buf

  (
    g160_p_spl_1,
    g160_p_spl_
  );


  buf

  (
    g160_p_spl_10,
    g160_p_spl_1
  );


  buf

  (
    g160_p_spl_11,
    g160_p_spl_1
  );


  buf

  (
    g162_p_spl_,
    g162_p
  );


  buf

  (
    g162_n_spl_,
    g162_n
  );


  buf

  (
    G39_p_spl_,
    G39_p
  );


  buf

  (
    g164_n_spl_,
    g164_n
  );


  buf

  (
    g164_n_spl_0,
    g164_n_spl_
  );


  buf

  (
    g164_n_spl_1,
    g164_n_spl_
  );


  buf

  (
    G39_n_spl_,
    G39_n
  );


  buf

  (
    g164_p_spl_,
    g164_p
  );


  buf

  (
    g164_p_spl_0,
    g164_p_spl_
  );


  buf

  (
    g164_p_spl_1,
    g164_p_spl_
  );


  buf

  (
    g149_n_spl_,
    g149_n
  );


  buf

  (
    g149_n_spl_0,
    g149_n_spl_
  );


  buf

  (
    g149_n_spl_1,
    g149_n_spl_
  );


  buf

  (
    g149_p_spl_,
    g149_p
  );


  buf

  (
    g149_p_spl_0,
    g149_p_spl_
  );


  buf

  (
    g149_p_spl_1,
    g149_p_spl_
  );


  buf

  (
    G54_n_spl_,
    G54_n
  );


  buf

  (
    G54_n_spl_0,
    G54_n_spl_
  );


  buf

  (
    G54_n_spl_00,
    G54_n_spl_0
  );


  buf

  (
    G54_n_spl_01,
    G54_n_spl_0
  );


  buf

  (
    G54_n_spl_1,
    G54_n_spl_
  );


  buf

  (
    G54_n_spl_10,
    G54_n_spl_1
  );


  buf

  (
    G54_n_spl_11,
    G54_n_spl_1
  );


  buf

  (
    g167_p_spl_,
    g167_p
  );


  buf

  (
    g167_p_spl_0,
    g167_p_spl_
  );


  buf

  (
    g172_n_spl_,
    g172_n
  );


  buf

  (
    g172_n_spl_0,
    g172_n_spl_
  );


  buf

  (
    g172_n_spl_00,
    g172_n_spl_0
  );


  buf

  (
    g172_n_spl_01,
    g172_n_spl_0
  );


  buf

  (
    g172_n_spl_1,
    g172_n_spl_
  );


  buf

  (
    g172_n_spl_10,
    g172_n_spl_1
  );


  buf

  (
    g172_n_spl_11,
    g172_n_spl_1
  );


  buf

  (
    g167_n_spl_,
    g167_n
  );


  buf

  (
    G53_n_spl_,
    G53_n
  );


  buf

  (
    G53_n_spl_0,
    G53_n_spl_
  );


  buf

  (
    G53_n_spl_00,
    G53_n_spl_0
  );


  buf

  (
    G53_n_spl_01,
    G53_n_spl_0
  );


  buf

  (
    G53_n_spl_1,
    G53_n_spl_
  );


  buf

  (
    G53_n_spl_10,
    G53_n_spl_1
  );


  buf

  (
    G53_n_spl_11,
    G53_n_spl_1
  );


  buf

  (
    g174_p_spl_,
    g174_p
  );


  buf

  (
    g176_p_spl_,
    g176_p
  );


  buf

  (
    G51_n_spl_,
    G51_n
  );


  buf

  (
    G51_n_spl_0,
    G51_n_spl_
  );


  buf

  (
    G51_n_spl_00,
    G51_n_spl_0
  );


  buf

  (
    G51_n_spl_000,
    G51_n_spl_00
  );


  buf

  (
    G51_n_spl_001,
    G51_n_spl_00
  );


  buf

  (
    G51_n_spl_01,
    G51_n_spl_0
  );


  buf

  (
    G51_n_spl_010,
    G51_n_spl_01
  );


  buf

  (
    G51_n_spl_011,
    G51_n_spl_01
  );


  buf

  (
    G51_n_spl_1,
    G51_n_spl_
  );


  buf

  (
    G51_n_spl_10,
    G51_n_spl_1
  );


  buf

  (
    G51_n_spl_11,
    G51_n_spl_1
  );


  buf

  (
    G58_n_spl_,
    G58_n
  );


  buf

  (
    g180_p_spl_,
    g180_p
  );


  buf

  (
    G52_n_spl_,
    G52_n
  );


  buf

  (
    G52_n_spl_0,
    G52_n_spl_
  );


  buf

  (
    G52_n_spl_00,
    G52_n_spl_0
  );


  buf

  (
    G52_n_spl_01,
    G52_n_spl_0
  );


  buf

  (
    G52_n_spl_1,
    G52_n_spl_
  );


  buf

  (
    G52_n_spl_10,
    G52_n_spl_1
  );


  buf

  (
    G52_n_spl_11,
    G52_n_spl_1
  );


  buf

  (
    g174_n_spl_,
    g174_n
  );


  buf

  (
    G35_p_spl_,
    G35_p
  );


  buf

  (
    G35_n_spl_,
    G35_n
  );


  buf

  (
    g194_p_spl_,
    g194_p
  );


  buf

  (
    g194_p_spl_0,
    g194_p_spl_
  );


  buf

  (
    G36_p_spl_,
    G36_p
  );


  buf

  (
    G36_n_spl_,
    G36_n
  );


  buf

  (
    g199_n_spl_,
    g199_n
  );


  buf

  (
    g199_p_spl_,
    g199_p
  );


  buf

  (
    g199_p_spl_0,
    g199_p_spl_
  );


  buf

  (
    G37_p_spl_,
    G37_p
  );


  buf

  (
    G37_n_spl_,
    G37_n
  );


  buf

  (
    g205_n_spl_,
    g205_n
  );


  buf

  (
    g205_p_spl_,
    g205_p
  );


  buf

  (
    g205_p_spl_0,
    g205_p_spl_
  );


  buf

  (
    g207_p_spl_,
    g207_p
  );


  buf

  (
    g208_p_spl_,
    g208_p
  );


  buf

  (
    g206_n_spl_,
    g206_n
  );


  buf

  (
    g206_p_spl_,
    g206_p
  );


  buf

  (
    g209_p_spl_,
    g209_p
  );


  buf

  (
    g201_p_spl_,
    g201_p
  );


  buf

  (
    g210_p_spl_,
    g210_p
  );


  buf

  (
    g200_n_spl_,
    g200_n
  );


  buf

  (
    g200_p_spl_,
    g200_p
  );


  buf

  (
    g211_p_spl_,
    g211_p
  );


  buf

  (
    g212_p_spl_,
    g212_p
  );


  buf

  (
    g194_n_spl_,
    g194_n
  );


  buf

  (
    g214_p_spl_,
    g214_p
  );


  buf

  (
    g216_p_spl_,
    g216_p
  );


  buf

  (
    g219_p_spl_,
    g219_p
  );


  buf

  (
    g214_n_spl_,
    g214_n
  );


  buf

  (
    g259_p_spl_,
    g259_p
  );


  buf

  (
    g259_p_spl_0,
    g259_p_spl_
  );


  buf

  (
    g259_p_spl_1,
    g259_p_spl_
  );


  buf

  (
    g259_n_spl_,
    g259_n
  );


  buf

  (
    g259_n_spl_0,
    g259_n_spl_
  );


  buf

  (
    g259_n_spl_1,
    g259_n_spl_
  );


  buf

  (
    G34_p_spl_,
    G34_p
  );


  buf

  (
    G34_p_spl_0,
    G34_p_spl_
  );


  buf

  (
    G34_p_spl_1,
    G34_p_spl_
  );


  buf

  (
    G34_n_spl_,
    G34_n
  );


  buf

  (
    G34_n_spl_0,
    G34_n_spl_
  );


  buf

  (
    G34_n_spl_1,
    G34_n_spl_
  );


  buf

  (
    g265_n_spl_,
    g265_n
  );


  buf

  (
    g265_n_spl_0,
    g265_n_spl_
  );


  buf

  (
    g265_n_spl_1,
    g265_n_spl_
  );


  buf

  (
    g265_p_spl_,
    g265_p
  );


  buf

  (
    g265_p_spl_0,
    g265_p_spl_
  );


  buf

  (
    g265_p_spl_1,
    g265_p_spl_
  );


  buf

  (
    g267_n_spl_,
    g267_n
  );


  buf

  (
    g267_p_spl_,
    g267_p
  );


  buf

  (
    g267_p_spl_0,
    g267_p_spl_
  );


  buf

  (
    g274_n_spl_,
    g274_n
  );


  buf

  (
    g274_p_spl_,
    g274_p
  );


  buf

  (
    g274_p_spl_0,
    g274_p_spl_
  );


  buf

  (
    g282_n_spl_,
    g282_n
  );


  buf

  (
    g282_p_spl_,
    g282_p
  );


  buf

  (
    g282_p_spl_0,
    g282_p_spl_
  );


  buf

  (
    g291_p_spl_,
    g291_p
  );


  buf

  (
    g291_p_spl_0,
    g291_p_spl_
  );


  buf

  (
    g291_n_spl_,
    g291_n
  );


  buf

  (
    g285_n_spl_,
    g285_n
  );


  buf

  (
    g292_n_spl_,
    g292_n
  );


  buf

  (
    g285_p_spl_,
    g285_p
  );


  buf

  (
    g292_p_spl_,
    g292_p
  );


  buf

  (
    g294_n_spl_,
    g294_n
  );


  buf

  (
    g294_n_spl_0,
    g294_n_spl_
  );


  buf

  (
    g294_p_spl_,
    g294_p
  );


  buf

  (
    g284_n_spl_,
    g284_n
  );


  buf

  (
    g295_n_spl_,
    g295_n
  );


  buf

  (
    g284_p_spl_,
    g284_p
  );


  buf

  (
    g295_p_spl_,
    g295_p
  );


  buf

  (
    g283_n_spl_,
    g283_n
  );


  buf

  (
    g283_n_spl_0,
    g283_n_spl_
  );


  buf

  (
    g283_p_spl_,
    g283_p
  );


  buf

  (
    g276_n_spl_,
    g276_n
  );


  buf

  (
    g297_n_spl_,
    g297_n
  );


  buf

  (
    g276_p_spl_,
    g276_p
  );


  buf

  (
    g297_p_spl_,
    g297_p
  );


  buf

  (
    g275_n_spl_,
    g275_n
  );


  buf

  (
    g275_n_spl_0,
    g275_n_spl_
  );


  buf

  (
    g275_p_spl_,
    g275_p
  );


  buf

  (
    g299_p_spl_,
    g299_p
  );


  buf

  (
    g300_p_spl_,
    g300_p
  );


  buf

  (
    g268_n_spl_,
    g268_n
  );


  buf

  (
    g268_n_spl_0,
    g268_n_spl_
  );


  buf

  (
    g303_n_spl_,
    g303_n
  );


  buf

  (
    g322_n_spl_,
    g322_n
  );


  buf

  (
    g337_n_spl_,
    g337_n
  );


  buf

  (
    g352_n_spl_,
    g352_n
  );


endmodule
