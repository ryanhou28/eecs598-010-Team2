// Benchmark "mymod" written by ABC on Sun Oct 29 19:32:01 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32,
    G6257, G6258, G6259, G6260, G6261, G6262, G6263, G6264, G6265, G6266,
    G6267, G6268, G6269, G6270, G6271, G6272, G6273, G6274, G6275, G6276,
    G6277, G6278, G6279, G6280, G6281, G6282, G6283, G6284, G6285, G6286,
    G6287, G6288  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32;
  output G6257, G6258, G6259, G6260, G6261, G6262, G6263, G6264, G6265, G6266,
    G6267, G6268, G6269, G6270, G6271, G6272, G6273, G6274, G6275, G6276,
    G6277, G6278, G6279, G6280, G6281, G6282, G6283, G6284, G6285, G6286,
    G6287, G6288;
  reg n2491_lo, n2575_lo, n2587_lo, n2599_lo, n2611_lo, n2623_lo, n2635_lo,
    n2647_lo, n2659_lo, n2671_lo, n2683_lo, n2734_lo, n2746_lo, n2758_lo,
    n2770_lo, n2782_lo, n2785_lo, n2794_lo, n2797_lo, n2806_lo, n2809_lo,
    n2818_lo, n2821_lo, n2830_lo, n2833_lo, n2836_lo, n2839_lo, n2842_lo,
    n2845_lo, n2848_lo, n2851_lo, n2854_lo, n2857_lo, n2860_lo, n2863_lo,
    n4871_o2, n4893_o2, n4938_o2, n5056_o2, n5100_o2, n5122_o2, n5254_o2,
    n5276_o2, n5316_o2, n5434_o2, n5473_o2, n5494_o2, n5620_o2, n5643_o2,
    n5682_o2, n5798_o2, n5839_o2, n5867_o2, n6052_o2, n6087_o2, n6153_o2,
    n6408_o2, n6454_o2, n6509_o2, n6775_o2, n6818_o2, n6892_o2, n5779_o2,
    n5780_o2, n7156_o2, n5792_o2, n7205_o2, n5842_o2, n5863_o2, n7263_o2,
    n5881_o2, n5930_o2, n5959_o2, n5981_o2, n6042_o2, n6075_o2, n6103_o2,
    n7610_o2, n6169_o2, n7665_o2, n6205_o2, n6239_o2, n7788_o2, n6309_o2,
    n6461_o2, n6476_o2, n325_inv, n6545_o2, G578_o2, G5106_o2, n6713_o2,
    G5164_o2, n343_inv, n6810_o2, n6973_o2, n352_inv, n7053_o2, G581_o2,
    G5467_o2, n7231_o2, G5527_o2, n370_inv, n7304_o2, n7530_o2, n379_inv,
    n7653_o2, G584_o2, G5820_o2, n7148_o2, n7149_o2, n7224_o2, n7916_o2,
    G5868_o2, n406_inv, n7280_o2, n7313_o2, n8056_o2, n7323_o2, n7398_o2,
    n7459_o2, n7501_o2, n7518_o2, G563_o2, n7606_o2, n439_inv, n7675_o2,
    G3410_o2, n7722_o2, n7747_o2, n7835_o2, G587_o2, G6046_o2, n7909_o2,
    G566_o2, G6070_o2, n472_inv, n8086_o2, n8093_o2, G3752_o2, n484_inv,
    n8199_o2, n2800_lo_buf_o2, G548_o2, n496_inv, G569_o2, G1761_o2,
    n505_inv, G4101_o2, G551_o2, n514_inv, G4743_o2, G5271_o2, G5790_o2,
    G6122_o2, G2082_o2, n2812_lo_buf_o2, n2668_lo_buf_o2, n2680_lo_buf_o2,
    G572_o2, G6125_o2, n547_inv, n2656_lo_buf_o2, G554_o2, G4452_o2,
    n559_inv, n2644_lo_buf_o2, G2410_o2, n2632_lo_buf_o2, n2620_lo_buf_o2,
    G6131_o2, G4693_o2, G5209_o2, G5741_o2, G6082_o2, G6119_o2,
    n2608_lo_buf_o2, n2596_lo_buf_o2, n2584_lo_buf_o2, n2572_lo_buf_o2,
    n2704_lo_buf_o2, G557_o2, G5936_o2, G5442_o2, G4926_o2, G6134_o2,
    G3929_o2, G4425_o2, G4947_o2, n2764_lo_buf_o2, n634_inv,
    n2560_lo_buf_o2, n2824_lo_buf_o2, G575_o2, G2740_o2, n649_inv,
    n2548_lo_buf_o2, n2536_lo_buf_o2, n2524_lo_buf_o2, G875_o2, G1064_o2,
    G1253_o2, G6140_o2, G5151_o2, G5686_o2, G6061_o2, G4803_o2, G5332_o2,
    G5844_o2, G6114_o2, G4806_o2, G3881_o2, G4370_o2, G4896_o2, G5001_o2,
    G3121_o2, n2512_lo_buf_o2, G4085_o2, G4605_o2, G5118_o2, G4997_o2,
    n2500_lo_buf_o2, n2716_lo_buf_o2, G560_o2, G1895_o2, G3064_o2,
    G3269_o2, G3569_o2, n748_inv, G1196_o2, G1007_o2, G818_o2, G674_o2,
    G5041_o2, G5562_o2, G6005_o2, G5214_o2, G5746_o2, G6087_o2, G6086_o2,
    G5745_o2, G5213_o2, G5893_o2, G5391_o2, G4864_o2, G6143_o2, G6008_o2,
    G5565_o2, G5044_o2, G3813_o2, G4325_o2, G4834_o2, G4993_o2, G3989_o2,
    G4490_o2, G5011_o2, G5112_o2, n2776_lo_buf_o2, G3298_o2, G3073_o2,
    G3265_o2, G3624_o2, G1642_o2, G1980_o2, n2488_lo_buf_o2, G626_o2,
    G1139_o2, G950_o2, G707_o2, G545_o2, G4217_o2, G4716_o2, G5244_o2,
    G3136_o2, G3499_o2, G3885_o2, G5243_o2, G3886_o2, G4375_o2, G4901_o2,
    G5054_o2, G4374_o2, G4900_o2, G5053_o2, G5242_o2, G4034_o2, G4556_o2,
    G5064_o2, G5172_o2, G2030_o2, G3016_o2, G3520_o2, G3261_o2, G3620_o2,
    G4220_o2, G4719_o2, G5247_o2, G5109_o2, G1638_o2, G1976_o2, G3560_o2,
    G3205_o2, G3193_o2, G3367_o2, G3670_o2, n979_inv, G1280_o2, G902_o2,
    G659_o2, G983_o2, G740_o2, G2917_o2, G3391_o2, G3494_o2, G1512_o2,
    G1854_o2, G2203_o2, G3493_o2, G3069_o2, G3574_o2, G3319_o2, G3667_o2,
    G3068_o2, G3573_o2, G3666_o2, G3318_o2, G3492_o2, G3241_o2, G3722_o2,
    G3422_o2, G1445_o2, G3257_o2, G3616_o2, G1634_o2, G1972_o2, G2256_o2,
    G3394_o2, G3557_o2, G3364_o2, G3719_o2, G2253_o2, G1583_o2, G1917_o2,
    G1727_o2, G2061_o2, G935_o2, G692_o2, G2136_o2, G1507_o2, G1849_o2,
    G2198_o2, G2197_o2, G1848_o2, G1689_o2, G2016_o2, G2314_o2, G2313_o2,
    G1688_o2, G2015_o2, G1847_o2, G2196_o2, G2118_o2, G1777_o2, G1630_o2,
    G1968_o2, G2309_o2, G2139_o2, G1580_o2, G2250_o2, G1914_o2, G1724_o2,
    G2058_o2, n2728_lo_buf_o2;
  wire new_new_n809__, new_new_n810__, new_new_n811__, new_new_n812__,
    new_new_n813__, new_new_n814__, new_new_n815__, new_new_n816__,
    new_new_n817__, new_new_n818__, new_new_n819__, new_new_n820__,
    new_new_n821__, new_new_n822__, new_new_n823__, new_new_n824__,
    new_new_n825__, new_new_n826__, new_new_n827__, new_new_n828__,
    new_new_n829__, new_new_n830__, new_new_n831__, new_new_n832__,
    new_new_n833__, new_new_n834__, new_new_n835__, new_new_n836__,
    new_new_n837__, new_new_n838__, new_new_n839__, new_new_n840__,
    new_new_n841__, new_new_n842__, new_new_n843__, new_new_n844__,
    new_new_n845__, new_new_n846__, new_new_n847__, new_new_n848__,
    new_new_n849__, new_new_n851__, new_new_n853__, new_new_n855__,
    new_new_n857__, new_new_n859__, new_new_n861__, new_new_n863__,
    new_new_n865__, new_new_n867__, new_new_n869__, new_new_n871__,
    new_new_n873__, new_new_n875__, new_new_n876__, new_new_n877__,
    new_new_n878__, new_new_n879__, new_new_n880__, new_new_n881__,
    new_new_n882__, new_new_n883__, new_new_n884__, new_new_n885__,
    new_new_n886__, new_new_n887__, new_new_n888__, new_new_n889__,
    new_new_n890__, new_new_n891__, new_new_n892__, new_new_n893__,
    new_new_n895__, new_new_n896__, new_new_n897__, new_new_n898__,
    new_new_n899__, new_new_n900__, new_new_n901__, new_new_n902__,
    new_new_n903__, new_new_n905__, new_new_n906__, new_new_n907__,
    new_new_n909__, new_new_n910__, new_new_n911__, new_new_n913__,
    new_new_n914__, new_new_n915__, new_new_n917__, new_new_n918__,
    new_new_n919__, new_new_n921__, new_new_n923__, new_new_n924__,
    new_new_n925__, new_new_n926__, new_new_n927__, new_new_n929__,
    new_new_n931__, new_new_n932__, new_new_n933__, new_new_n934__,
    new_new_n935__, new_new_n937__, new_new_n939__, new_new_n940__,
    new_new_n941__, new_new_n942__, new_new_n943__, new_new_n946__,
    new_new_n947__, new_new_n949__, new_new_n952__, new_new_n953__,
    new_new_n955__, new_new_n958__, new_new_n959__, new_new_n961__,
    new_new_n964__, new_new_n965__, new_new_n967__, new_new_n970__,
    new_new_n971__, new_new_n973__, new_new_n976__, new_new_n977__,
    new_new_n979__, new_new_n982__, new_new_n983__, new_new_n985__,
    new_new_n988__, new_new_n989__, new_new_n991__, new_new_n994__,
    new_new_n995__, new_new_n997__, new_new_n998__, new_new_n999__,
    new_new_n1001__, new_new_n1003__, new_new_n1004__, new_new_n1006__,
    new_new_n1007__, new_new_n1008__, new_new_n1009__, new_new_n1010__,
    new_new_n1011__, new_new_n1013__, new_new_n1014__, new_new_n1015__,
    new_new_n1016__, new_new_n1017__, new_new_n1018__, new_new_n1019__,
    new_new_n1020__, new_new_n1021__, new_new_n1022__, new_new_n1023__,
    new_new_n1024__, new_new_n1025__, new_new_n1026__, new_new_n1027__,
    new_new_n1029__, new_new_n1030__, new_new_n1032__, new_new_n1033__,
    new_new_n1034__, new_new_n1035__, new_new_n1036__, new_new_n1037__,
    new_new_n1039__, new_new_n1040__, new_new_n1041__, new_new_n1042__,
    new_new_n1043__, new_new_n1045__, new_new_n1047__, new_new_n1049__,
    new_new_n1052__, new_new_n1053__, new_new_n1055__, new_new_n1057__,
    new_new_n1059__, new_new_n1061__, new_new_n1063__, new_new_n1065__,
    new_new_n1067__, new_new_n1070__, new_new_n1071__, new_new_n1073__,
    new_new_n1075__, new_new_n1077__, new_new_n1079__, new_new_n1081__,
    new_new_n1083__, new_new_n1085__, new_new_n1088__, new_new_n1089__,
    new_new_n1090__, new_new_n1091__, new_new_n1093__, new_new_n1094__,
    new_new_n1095__, new_new_n1097__, new_new_n1099__, new_new_n1101__,
    new_new_n1102__, new_new_n1103__, new_new_n1104__, new_new_n1105__,
    new_new_n1107__, new_new_n1108__, new_new_n1109__, new_new_n1110__,
    new_new_n1111__, new_new_n1112__, new_new_n1113__, new_new_n1114__,
    new_new_n1115__, new_new_n1116__, new_new_n1117__, new_new_n1119__,
    new_new_n1120__, new_new_n1121__, new_new_n1123__, new_new_n1124__,
    new_new_n1125__, new_new_n1127__, new_new_n1128__, new_new_n1129__,
    new_new_n1130__, new_new_n1131__, new_new_n1132__, new_new_n1133__,
    new_new_n1136__, new_new_n1137__, new_new_n1138__, new_new_n1139__,
    new_new_n1141__, new_new_n1143__, new_new_n1145__, new_new_n1146__,
    new_new_n1147__, new_new_n1149__, new_new_n1151__, new_new_n1153__,
    new_new_n1155__, new_new_n1156__, new_new_n1157__, new_new_n1159__,
    new_new_n1161__, new_new_n1163__, new_new_n1165__, new_new_n1167__,
    new_new_n1169__, new_new_n1171__, new_new_n1173__, new_new_n1174__,
    new_new_n1175__, new_new_n1176__, new_new_n1177__, new_new_n1178__,
    new_new_n1180__, new_new_n1181__, new_new_n1183__, new_new_n1184__,
    new_new_n1185__, new_new_n1186__, new_new_n1187__, new_new_n1189__,
    new_new_n1191__, new_new_n1193__, new_new_n1195__, new_new_n1196__,
    new_new_n1197__, new_new_n1199__, new_new_n1201__, new_new_n1203__,
    new_new_n1204__, new_new_n1205__, new_new_n1207__, new_new_n1208__,
    new_new_n1209__, new_new_n1210__, new_new_n1211__, new_new_n1213__,
    new_new_n1214__, new_new_n1215__, new_new_n1216__, new_new_n1217__,
    new_new_n1218__, new_new_n1219__, new_new_n1220__, new_new_n1222__,
    new_new_n1223__, new_new_n1224__, new_new_n1225__, new_new_n1226__,
    new_new_n1227__, new_new_n1228__, new_new_n1229__, new_new_n1230__,
    new_new_n1231__, new_new_n1232__, new_new_n1233__, new_new_n1235__,
    new_new_n1236__, new_new_n1237__, new_new_n1238__, new_new_n1239__,
    new_new_n1240__, new_new_n1241__, new_new_n1243__, new_new_n1244__,
    new_new_n1245__, new_new_n1246__, new_new_n1247__, new_new_n1248__,
    new_new_n1249__, new_new_n1250__, new_new_n1251__, new_new_n1253__,
    new_new_n1254__, new_new_n1255__, new_new_n1256__, new_new_n1257__,
    new_new_n1259__, new_new_n1261__, new_new_n1263__, new_new_n1264__,
    new_new_n1265__, new_new_n1266__, new_new_n1267__, new_new_n1268__,
    new_new_n1269__, new_new_n1270__, new_new_n1271__, new_new_n1272__,
    new_new_n1273__, new_new_n1274__, new_new_n1275__, new_new_n1277__,
    new_new_n1278__, new_new_n1279__, new_new_n1280__, new_new_n1281__,
    new_new_n1282__, new_new_n1283__, new_new_n1284__, new_new_n1285__,
    new_new_n1286__, new_new_n1287__, new_new_n1288__, new_new_n1290__,
    new_new_n1291__, new_new_n1293__, new_new_n1294__, new_new_n1295__,
    new_new_n1296__, new_new_n1297__, new_new_n1298__, new_new_n1299__,
    new_new_n1300__, new_new_n1301__, new_new_n1302__, new_new_n1303__,
    new_new_n1304__, new_new_n1305__, new_new_n1306__, new_new_n1307__,
    new_new_n1308__, new_new_n1309__, new_new_n1310__, new_new_n1311__,
    new_new_n1312__, new_new_n1313__, new_new_n1314__, new_new_n1315__,
    new_new_n1316__, new_new_n1317__, new_new_n1319__, new_new_n1320__,
    new_new_n1321__, new_new_n1322__, new_new_n1323__, new_new_n1324__,
    new_new_n1325__, new_new_n1326__, new_new_n1327__, new_new_n1329__,
    new_new_n1330__, new_new_n1331__, new_new_n1332__, new_new_n1333__,
    new_new_n1334__, new_new_n1335__, new_new_n1336__, new_new_n1337__,
    new_new_n1338__, new_new_n1339__, new_new_n1340__, new_new_n1341__,
    new_new_n1342__, new_new_n1343__, new_new_n1344__, new_new_n1345__,
    new_new_n1346__, new_new_n1347__, new_new_n1348__, new_new_n1349__,
    new_new_n1350__, new_new_n1351__, new_new_n1352__, new_new_n1353__,
    new_new_n1354__, new_new_n1355__, new_new_n1356__, new_new_n1357__,
    new_new_n1358__, new_new_n1359__, new_new_n1360__, new_new_n1361__,
    new_new_n1362__, new_new_n1363__, new_new_n1364__, new_new_n1365__,
    new_new_n1366__, new_new_n1367__, new_new_n1368__, new_new_n1369__,
    new_new_n1370__, new_new_n1371__, new_new_n1372__, new_new_n1373__,
    new_new_n1374__, new_new_n1375__, new_new_n1376__, new_new_n1377__,
    new_new_n1378__, new_new_n1379__, new_new_n1380__, new_new_n1381__,
    new_new_n1382__, new_new_n1383__, new_new_n1384__, new_new_n1385__,
    new_new_n1386__, new_new_n1387__, new_new_n1388__, new_new_n1389__,
    new_new_n1391__, new_new_n1392__, new_new_n1393__, new_new_n1394__,
    new_new_n1395__, new_new_n1396__, new_new_n1397__, new_new_n1398__,
    new_new_n1399__, new_new_n1400__, new_new_n1401__, new_new_n1402__,
    new_new_n1403__, new_new_n1404__, new_new_n1405__, new_new_n1406__,
    new_new_n1407__, new_new_n1408__, new_new_n1409__, new_new_n1411__,
    new_new_n1412__, new_new_n1413__, new_new_n1414__, new_new_n1415__,
    new_new_n1416__, new_new_n1417__, new_new_n1418__, new_new_n1419__,
    new_new_n1420__, new_new_n1421__, new_new_n1422__, new_new_n1423__,
    new_new_n1424__, new_new_n1425__, new_new_n1426__, new_new_n1427__,
    new_new_n1428__, new_new_n1429__, new_new_n1430__, new_new_n1431__,
    new_new_n1432__, new_new_n1433__, new_new_n1434__, new_new_n1435__,
    new_new_n1436__, new_new_n1437__, new_new_n1438__, new_new_n1439__,
    new_new_n1440__, new_new_n1441__, new_new_n1442__, new_new_n1443__,
    new_new_n1444__, new_new_n1445__, new_new_n1446__, new_new_n1447__,
    new_new_n1448__, new_new_n1449__, new_new_n1450__, new_new_n1451__,
    new_new_n1452__, new_new_n1453__, new_new_n1454__, new_new_n1455__,
    new_new_n1456__, new_new_n1457__, new_new_n1458__, new_new_n1459__,
    new_new_n1460__, new_new_n1461__, new_new_n1462__, new_new_n1463__,
    new_new_n1464__, new_new_n1465__, new_new_n1466__, new_new_n1467__,
    new_new_n1468__, new_new_n1469__, new_new_n1470__, new_new_n1471__,
    new_new_n1472__, new_new_n1473__, new_new_n1474__, new_new_n1475__,
    new_new_n1476__, new_new_n1477__, new_new_n1478__, new_new_n1479__,
    new_new_n1480__, new_new_n1481__, new_new_n1483__, new_new_n1484__,
    new_new_n1485__, new_new_n1486__, new_new_n1487__, new_new_n1488__,
    new_new_n1489__, new_new_n1490__, new_new_n1491__, new_new_n1492__,
    new_new_n1493__, new_new_n1494__, new_new_n1495__, new_new_n1496__,
    new_new_n1497__, new_new_n1498__, new_new_n1499__, new_new_n1500__,
    new_new_n1501__, new_new_n1502__, new_new_n1503__, new_new_n1504__,
    new_new_n1505__, new_new_n1506__, new_new_n1507__, new_new_n1508__,
    new_new_n1509__, new_new_n1510__, new_new_n1511__, new_new_n1512__,
    new_new_n1513__, new_new_n1514__, new_new_n1515__, new_new_n1516__,
    new_new_n1517__, new_new_n1518__, new_new_n1519__, new_new_n1520__,
    new_new_n1521__, new_new_n1522__, new_new_n1523__, new_new_n1524__,
    new_new_n1525__, new_new_n1526__, new_new_n1527__, new_new_n1528__,
    new_new_n1529__, new_new_n1530__, new_new_n1531__, new_new_n1533__,
    new_new_n1534__, new_new_n1535__, new_new_n1536__, new_new_n1537__,
    new_new_n1538__, new_new_n1539__, new_new_n1540__, new_new_n1541__,
    new_new_n1542__, new_new_n1543__, new_new_n1544__, new_new_n1545__,
    new_new_n1546__, new_new_n1547__, new_new_n1548__, new_new_n1549__,
    new_new_n1550__, new_new_n1551__, new_new_n1552__, new_new_n1553__,
    new_new_n1554__, new_new_n1555__, new_new_n1556__, new_new_n1557__,
    new_new_n1558__, new_new_n1559__, new_new_n1560__, new_new_n1561__,
    new_new_n1562__, new_new_n1563__, new_new_n1564__, new_new_n1565__,
    new_new_n1566__, new_new_n1567__, new_new_n1568__, new_new_n1569__,
    new_new_n1570__, new_new_n1571__, new_new_n1572__, new_new_n1573__,
    new_new_n1574__, new_new_n1575__, new_new_n1576__, new_new_n1577__,
    new_new_n1578__, new_new_n1579__, new_new_n1580__, new_new_n1581__,
    new_new_n1582__, new_new_n1583__, new_new_n1584__, new_new_n1585__,
    new_new_n1586__, new_new_n1587__, new_new_n1588__, new_new_n1589__,
    new_new_n1590__, new_new_n1591__, new_new_n1592__, new_new_n1593__,
    new_new_n1594__, new_new_n1595__, new_new_n1596__, new_new_n1597__,
    new_new_n1598__, new_new_n1599__, new_new_n1600__, new_new_n1601__,
    new_new_n1602__, new_new_n1603__, new_new_n1604__, new_new_n1605__,
    new_new_n1606__, new_new_n1607__, new_new_n1608__, new_new_n1609__,
    new_new_n1610__, new_new_n1611__, new_new_n1612__, new_new_n1613__,
    new_new_n1614__, new_new_n1615__, new_new_n1616__, new_new_n1617__,
    new_new_n1618__, new_new_n1619__, new_new_n1620__, new_new_n1621__,
    new_new_n1622__, new_new_n1623__, new_new_n1624__, new_new_n1625__,
    new_new_n1626__, new_new_n1627__, new_new_n1628__, new_new_n1629__,
    new_new_n1630__, new_new_n1631__, new_new_n1632__, new_new_n1633__,
    new_new_n1634__, new_new_n1635__, new_new_n1636__, new_new_n1637__,
    new_new_n1638__, new_new_n1639__, new_new_n1640__, new_new_n1641__,
    new_new_n1642__, new_new_n1643__, new_new_n1644__, new_new_n1645__,
    new_new_n1646__, new_new_n1647__, new_new_n1648__, new_new_n1649__,
    new_new_n1650__, new_new_n1651__, new_new_n1652__, new_new_n1653__,
    new_new_n1654__, new_new_n1655__, new_new_n1656__, new_new_n1657__,
    new_new_n1658__, new_new_n1659__, new_new_n1660__, new_new_n1661__,
    new_new_n1662__, new_new_n1663__, new_new_n1664__, new_new_n1665__,
    new_new_n1666__, new_new_n1667__, new_new_n1668__, new_new_n1669__,
    new_new_n1670__, new_new_n1671__, new_new_n1672__, new_new_n1673__,
    new_new_n1674__, new_new_n1675__, new_new_n1676__, new_new_n1677__,
    new_new_n1678__, new_new_n1679__, new_new_n1680__, new_new_n1681__,
    new_new_n1682__, new_new_n1683__, new_new_n1684__, new_new_n1685__,
    new_new_n1686__, new_new_n1687__, new_new_n1688__, new_new_n1689__,
    new_new_n1690__, new_new_n1691__, new_new_n1692__, new_new_n1693__,
    new_new_n1694__, new_new_n1695__, new_new_n1696__, new_new_n1697__,
    new_new_n1698__, new_new_n1699__, new_new_n1700__, new_new_n1701__,
    new_new_n1702__, new_new_n1703__, new_new_n1704__, new_new_n1705__,
    new_new_n1706__, new_new_n1707__, new_new_n1708__, new_new_n1709__,
    new_new_n1710__, new_new_n1711__, new_new_n1712__, new_new_n1713__,
    new_new_n1714__, new_new_n1715__, new_new_n1716__, new_new_n1717__,
    new_new_n1718__, new_new_n1719__, new_new_n1720__, new_new_n1721__,
    new_new_n1722__, new_new_n1723__, new_new_n1724__, new_new_n1725__,
    new_new_n1726__, new_new_n1727__, new_new_n1728__, new_new_n1729__,
    new_new_n1730__, new_new_n1731__, new_new_n1732__, new_new_n1733__,
    new_new_n1734__, new_new_n1735__, new_new_n1736__, new_new_n1737__,
    new_new_n1738__, new_new_n1739__, new_new_n1740__, new_new_n1741__,
    new_new_n1742__, new_new_n1743__, new_new_n1744__, new_new_n1745__,
    new_new_n1746__, new_new_n1747__, new_new_n1748__, new_new_n1749__,
    new_new_n1750__, new_new_n1751__, new_new_n1752__, new_new_n1753__,
    new_new_n1754__, new_new_n1755__, new_new_n1756__, new_new_n1757__,
    new_new_n1758__, new_new_n1759__, new_new_n1760__, new_new_n1761__,
    new_new_n1762__, new_new_n1763__, new_new_n1764__, new_new_n1765__,
    new_new_n1766__, new_new_n1767__, new_new_n1768__, new_new_n1769__,
    new_new_n1770__, new_new_n1771__, new_new_n1772__, new_new_n1773__,
    new_new_n1774__, new_new_n1775__, new_new_n1776__, new_new_n1777__,
    new_new_n1778__, new_new_n1779__, new_new_n1780__, new_new_n1781__,
    new_new_n1782__, new_new_n1783__, new_new_n1784__, new_new_n1785__,
    new_new_n1786__, new_new_n1787__, new_new_n1788__, new_new_n1789__,
    new_new_n1790__, new_new_n1791__, new_new_n1792__, new_new_n1793__,
    new_new_n1794__, new_new_n1795__, new_new_n1796__, new_new_n1797__,
    new_new_n1798__, new_new_n1799__, new_new_n1800__, new_new_n1801__,
    new_new_n1802__, new_new_n1803__, new_new_n1804__, new_new_n1805__,
    new_new_n1806__, new_new_n1807__, new_new_n1808__, new_new_n1809__,
    new_new_n1810__, new_new_n1811__, new_new_n1812__, new_new_n1813__,
    new_new_n1814__, new_new_n1815__, new_new_n1816__, new_new_n1817__,
    new_new_n1818__, new_new_n1819__, new_new_n1820__, new_new_n1821__,
    new_new_n1822__, new_new_n1823__, new_new_n1824__, new_new_n1825__,
    new_new_n1826__, new_new_n1827__, new_new_n1828__, new_new_n1829__,
    new_new_n1830__, new_new_n1831__, new_new_n1832__, new_new_n1833__,
    new_new_n1834__, new_new_n1835__, new_new_n1836__, new_new_n1837__,
    new_new_n1838__, new_new_n1839__, new_new_n1840__, new_new_n1841__,
    new_new_n1842__, new_new_n1843__, new_new_n1844__, new_new_n1845__,
    new_new_n1846__, new_new_n1847__, new_new_n1848__, new_new_n1849__,
    new_new_n1850__, new_new_n1851__, new_new_n1852__, new_new_n1853__,
    new_new_n1854__, new_new_n1855__, new_new_n1856__, new_new_n1857__,
    new_new_n1858__, new_new_n1859__, new_new_n1860__, new_new_n1861__,
    new_new_n1862__, new_new_n1863__, new_new_n1864__, new_new_n1865__,
    new_new_n1866__, new_new_n1867__, new_new_n1868__, new_new_n1869__,
    new_new_n1870__, new_new_n1871__, new_new_n1872__, new_new_n1873__,
    new_new_n1874__, new_new_n1875__, new_new_n1876__, new_new_n1877__,
    new_new_n1878__, new_new_n1879__, new_new_n1880__, new_new_n1881__,
    new_new_n1882__, new_new_n1883__, new_new_n1884__, new_new_n1885__,
    new_new_n1886__, new_new_n1887__, new_new_n1888__, new_new_n1889__,
    new_new_n1890__, new_new_n1891__, new_new_n1892__, new_new_n1893__,
    new_new_n1894__, new_new_n1895__, new_new_n1896__, new_new_n1897__,
    new_new_n1898__, new_new_n1899__, new_new_n1900__, new_new_n1901__,
    new_new_n1902__, new_new_n1903__, new_new_n1904__, new_new_n1905__,
    new_new_n1906__, new_new_n1907__, new_new_n1908__, new_new_n1909__,
    new_new_n1910__, new_new_n1911__, new_new_n1912__, new_new_n1913__,
    new_new_n1914__, new_new_n1915__, new_new_n1916__, new_new_n1917__,
    new_new_n1918__, new_new_n1919__, new_new_n1920__, new_new_n1921__,
    new_new_n1922__, new_new_n1923__, new_new_n1924__, new_new_n1925__,
    new_new_n1926__, new_new_n1927__, new_new_n1928__, new_new_n1929__,
    new_new_n1930__, new_new_n1931__, new_new_n1932__, new_new_n1933__,
    new_new_n1934__, new_new_n1935__, new_new_n1936__, new_new_n1937__,
    new_new_n1938__, new_new_n1939__, new_new_n1940__, new_new_n1941__,
    new_new_n1942__, new_new_n1943__, new_new_n1944__, new_new_n1945__,
    new_new_n1946__, new_new_n1947__, new_new_n1948__, new_new_n1949__,
    new_new_n1950__, new_new_n1951__, new_new_n1952__, new_new_n1953__,
    new_new_n1954__, new_new_n1955__, new_new_n1956__, new_new_n1957__,
    new_new_n1958__, new_new_n1959__, new_new_n1960__, new_new_n1961__,
    new_new_n1962__, new_new_n1963__, new_new_n1964__, new_new_n1965__,
    new_new_n1966__, new_new_n1967__, new_new_n1968__, new_new_n1969__,
    new_new_n1970__, new_new_n1971__, new_new_n1972__, new_new_n1973__,
    new_new_n1974__, new_new_n1975__, new_new_n1976__, new_new_n1977__,
    new_new_n1978__, new_new_n1979__, new_new_n1980__, new_new_n1981__,
    new_new_n1982__, new_new_n1983__, new_new_n1984__, new_new_n1985__,
    new_new_n1986__, new_new_n1987__, new_new_n1988__, new_new_n1989__,
    new_new_n1990__, new_new_n1991__, new_new_n1992__, new_new_n1993__,
    new_new_n1994__, new_new_n1995__, new_new_n1996__, new_new_n1997__,
    new_new_n1998__, new_new_n1999__, new_new_n2000__, new_new_n2001__,
    new_new_n2002__, new_new_n2003__, new_new_n2004__, new_new_n2005__,
    new_new_n2006__, new_new_n2007__, new_new_n2008__, new_new_n2009__,
    new_new_n2010__, new_new_n2011__, new_new_n2012__, new_new_n2013__,
    new_new_n2014__, new_new_n2015__, new_new_n2016__, new_new_n2017__,
    new_new_n2018__, new_new_n2019__, new_new_n2020__, new_new_n2021__,
    new_new_n2022__, new_new_n2023__, new_new_n2024__, new_new_n2025__,
    new_new_n2026__, new_new_n2027__, new_new_n2028__, new_new_n2029__,
    new_new_n2030__, new_new_n2031__, new_new_n2032__, new_new_n2033__,
    new_new_n2034__, new_new_n2035__, new_new_n2036__, new_new_n2037__,
    new_new_n2038__, new_new_n2039__, new_new_n2040__, new_new_n2041__,
    new_new_n2042__, new_new_n2043__, new_new_n2044__, new_new_n2045__,
    new_new_n2046__, new_new_n2047__, new_new_n2048__, new_new_n2049__,
    new_new_n2050__, new_new_n2051__, new_new_n2052__, new_new_n2053__,
    new_new_n2054__, new_new_n2055__, new_new_n2056__, new_new_n2057__,
    new_new_n2058__, new_new_n2059__, new_new_n2060__, new_new_n2061__,
    new_new_n2062__, new_new_n2063__, new_new_n2064__, new_new_n2065__,
    new_new_n2066__, new_new_n2067__, new_new_n2068__, new_new_n2069__,
    new_new_n2070__, new_new_n2071__, new_new_n2072__, new_new_n2073__,
    new_new_n2074__, new_new_n2075__, new_new_n2076__, new_new_n2077__,
    new_new_n2078__, new_new_n2079__, new_new_n2080__, new_new_n2081__,
    new_new_n2082__, new_new_n2083__, new_new_n2084__, new_new_n2085__,
    new_new_n2086__, new_new_n2087__, new_new_n2088__, new_new_n2089__,
    new_new_n2090__, new_new_n2091__, new_new_n2092__, new_new_n2093__,
    new_new_n2094__, new_new_n2095__, new_new_n2096__, new_new_n2097__,
    new_new_n2098__, new_new_n2099__, new_new_n2100__, new_new_n2101__,
    new_new_n2102__, new_new_n2103__, new_new_n2104__, new_new_n2105__,
    new_new_n2106__, new_new_n2107__, new_new_n2108__, new_new_n2109__,
    new_new_n2110__, new_new_n2111__, new_new_n2112__, new_new_n2113__,
    new_new_n2114__, new_new_n2115__, new_new_n2116__, new_new_n2117__,
    new_new_n2118__, new_new_n2119__, new_new_n2120__, new_new_n2121__,
    new_new_n2122__, new_new_n2123__, new_new_n2124__, new_new_n2125__,
    new_new_n2126__, new_new_n2127__, new_new_n2128__, new_new_n2129__,
    new_new_n2130__, new_new_n2131__, new_new_n2132__, new_new_n2133__,
    new_new_n2134__, new_new_n2135__, new_new_n2136__, new_new_n2137__,
    new_new_n2138__, new_new_n2139__, new_new_n2140__, new_new_n2141__,
    new_new_n2142__, new_new_n2143__, new_new_n2144__, new_new_n2145__,
    new_new_n2146__, new_new_n2147__, new_new_n2148__, new_new_n2149__,
    new_new_n2150__, new_new_n2151__, new_new_n2152__, new_new_n2153__,
    new_new_n2154__, new_new_n2155__, new_new_n2156__, new_new_n2157__,
    new_new_n2158__, new_new_n2159__, new_new_n2160__, new_new_n2161__,
    new_new_n2162__, new_new_n2163__, new_new_n2164__, new_new_n2165__,
    new_new_n2166__, new_new_n2167__, new_new_n2168__, new_new_n2169__,
    new_new_n2170__, new_new_n2171__, new_new_n2172__, new_new_n2173__,
    new_new_n2174__, new_new_n2175__, new_new_n2176__, new_new_n2177__,
    new_new_n2178__, new_new_n2179__, new_new_n2180__, new_new_n2181__,
    new_new_n2182__, new_new_n2183__, new_new_n2184__, new_new_n2185__,
    new_new_n2186__, new_new_n2187__, new_new_n2188__, new_new_n2189__,
    new_new_n2190__, new_new_n2191__, new_new_n2192__, new_new_n2193__,
    new_new_n2194__, new_new_n2195__, new_new_n2196__, new_new_n2197__,
    new_new_n2198__, new_new_n2199__, new_new_n2200__, new_new_n2201__,
    new_new_n2202__, new_new_n2203__, new_new_n2204__, new_new_n2205__,
    new_new_n2206__, new_new_n2207__, new_new_n2208__, new_new_n2209__,
    new_new_n2210__, new_new_n2211__, new_new_n2212__, new_new_n2213__,
    new_new_n2214__, new_new_n2215__, new_new_n2216__, new_new_n2217__,
    new_new_n2218__, new_new_n2219__, new_new_n2220__, new_new_n2221__,
    new_new_n2222__, new_new_n2223__, new_new_n2224__, new_new_n2225__,
    new_new_n2226__, new_new_n2227__, new_new_n2228__, new_new_n2229__,
    new_new_n2230__, new_new_n2231__, new_new_n2232__, new_new_n2233__,
    new_new_n2234__, new_new_n2235__, new_new_n2236__, new_new_n2237__,
    new_new_n2238__, new_new_n2239__, new_new_n2240__, new_new_n2241__,
    new_new_n2242__, new_new_n2243__, new_new_n2244__, new_new_n2245__,
    new_new_n2246__, new_new_n2247__, new_new_n2248__, new_new_n2249__,
    new_new_n2250__, new_new_n2251__, new_new_n2252__, new_new_n2253__,
    new_new_n2254__, new_new_n2255__, new_new_n2256__, new_new_n2257__,
    new_new_n2258__, new_new_n2259__, new_new_n2260__, new_new_n2261__,
    new_new_n2262__, new_new_n2263__, new_new_n2264__, new_new_n2265__,
    new_new_n2266__, new_new_n2267__, new_new_n2268__, new_new_n2269__,
    new_new_n2270__, new_new_n2271__, new_new_n2272__, new_new_n2273__,
    new_new_n2274__, new_new_n2275__, new_new_n2276__, new_new_n2277__,
    new_new_n2278__, new_new_n2279__, new_new_n2280__, new_new_n2281__,
    new_new_n2282__, new_new_n2283__, new_new_n2284__, new_new_n2285__,
    new_new_n2286__, new_new_n2287__, new_new_n2288__, new_new_n2289__,
    new_new_n2290__, new_new_n2291__, new_new_n2292__, new_new_n2293__,
    new_new_n2294__, new_new_n2295__, new_new_n2296__, new_new_n2297__,
    new_new_n2298__, new_new_n2299__, new_new_n2300__, new_new_n2301__,
    new_new_n2302__, new_new_n2303__, new_new_n2304__, new_new_n2305__,
    new_new_n2306__, new_new_n2307__, new_new_n2308__, new_new_n2309__,
    new_new_n2310__, new_new_n2311__, new_new_n2312__, new_new_n2313__,
    new_new_n2314__, new_new_n2315__, new_new_n2316__, new_new_n2317__,
    new_new_n2318__, new_new_n2319__, new_new_n2320__, new_new_n2321__,
    new_new_n2322__, new_new_n2323__, new_new_n2324__, new_new_n2325__,
    new_new_n2326__, new_new_n2327__, new_new_n2328__, new_new_n2329__,
    new_new_n2330__, new_new_n2331__, new_new_n2332__, new_new_n2333__,
    new_new_n2334__, new_new_n2335__, new_new_n2336__, new_new_n2337__,
    new_new_n2338__, new_new_n2339__, new_new_n2340__, new_new_n2341__,
    new_new_n2342__, new_new_n2343__, new_new_n2344__, new_new_n2345__,
    new_new_n2346__, new_new_n2347__, new_new_n2348__, new_new_n2349__,
    new_new_n2350__, new_new_n2351__, new_new_n2352__, new_new_n2353__,
    new_new_n2354__, new_new_n2355__, new_new_n2356__, new_new_n2357__,
    new_new_n2358__, new_new_n2359__, new_new_n2360__, new_new_n2361__,
    new_new_n2362__, new_new_n2363__, new_new_n2364__, new_new_n2365__,
    new_new_n2366__, new_new_n2367__, new_new_n2368__, new_new_n2369__,
    new_new_n2370__, new_new_n2371__, new_new_n2372__, new_new_n2373__,
    new_new_n2374__, new_new_n2375__, new_new_n2376__, new_new_n2377__,
    new_new_n2378__, new_new_n2379__, new_new_n2380__, new_new_n2381__,
    new_new_n2382__, new_new_n2383__, new_new_n2384__, new_new_n2385__,
    new_new_n2386__, new_new_n2387__, new_new_n2388__, new_new_n2389__,
    new_new_n2390__, new_new_n2391__, new_new_n2392__, new_new_n2393__,
    new_new_n2394__, new_new_n2395__, new_new_n2396__, new_new_n2397__,
    new_new_n2398__, new_new_n2399__, new_new_n2400__, new_new_n2401__,
    new_new_n2402__, new_new_n2403__, new_new_n2404__, new_new_n2405__,
    new_new_n2406__, new_new_n2407__, new_new_n2408__, new_new_n2409__,
    new_new_n2410__, new_new_n2411__, new_new_n2412__, new_new_n2413__,
    new_new_n2414__, new_new_n2415__, new_new_n2416__, new_new_n2417__,
    new_new_n2418__, new_new_n2419__, new_new_n2420__, new_new_n2421__,
    new_new_n2422__, new_new_n2423__, new_new_n2424__, new_new_n2425__,
    new_new_n2426__, new_new_n2427__, new_new_n2428__, new_new_n2429__,
    new_new_n2430__, new_new_n2431__, new_new_n2432__, new_new_n2433__,
    new_new_n2434__, new_new_n2435__, new_new_n2436__, new_new_n2437__,
    new_new_n2438__, new_new_n2439__, new_new_n2440__, new_new_n2441__,
    new_new_n2442__, new_new_n2443__, new_new_n2444__, new_new_n2445__,
    new_new_n2446__, new_new_n2447__, new_new_n2448__, new_new_n2449__,
    new_new_n2450__, new_new_n2451__, new_new_n2452__, new_new_n2453__,
    new_new_n2454__, new_new_n2455__, new_new_n2456__, new_new_n2457__,
    new_new_n2458__, new_new_n2459__, new_new_n2460__, new_new_n2461__,
    new_new_n2462__, new_new_n2463__, new_new_n2464__, new_new_n2465__,
    new_new_n2466__, new_new_n2467__, new_new_n2468__, new_new_n2469__,
    new_new_n2470__, new_new_n2471__, new_new_n2472__, new_new_n2473__,
    new_new_n2474__, new_new_n2475__, new_new_n2476__, new_new_n2477__,
    new_new_n2478__, new_new_n2479__, new_new_n2480__, new_new_n2481__,
    new_new_n2482__, new_new_n2483__, new_new_n2484__, new_new_n2485__,
    new_new_n2486__, new_new_n2487__, new_new_n2488__, new_new_n2489__,
    new_new_n2490__, new_new_n2491__, new_new_n2492__, new_new_n2493__,
    new_new_n2494__, new_new_n2495__, new_new_n2496__, new_new_n2497__,
    new_new_n2498__, new_new_n2499__, new_new_n2500__, new_new_n2501__,
    new_new_n2502__, new_new_n2503__, new_new_n2504__, new_new_n2505__,
    new_new_n2506__, new_new_n2507__, new_new_n2508__, new_new_n2509__,
    new_new_n2510__, new_new_n2511__, new_new_n2512__, new_new_n2513__,
    new_new_n2514__, new_new_n2515__, new_new_n2516__, new_new_n2517__,
    new_new_n2518__, new_new_n2519__, new_new_n2520__, new_new_n2521__,
    new_new_n2522__, new_new_n2523__, new_new_n2524__, new_new_n2525__,
    new_new_n2526__, new_new_n2527__, new_new_n2528__, new_new_n2529__,
    new_new_n2530__, new_new_n2531__, new_new_n2532__, new_new_n2533__,
    new_new_n2534__, new_new_n2535__, new_new_n2536__, new_new_n2537__,
    new_new_n2538__, new_new_n2539__, new_new_n2540__, new_new_n2541__,
    new_new_n2542__, new_new_n2543__, new_new_n2544__, new_new_n2545__,
    new_new_n2546__, new_new_n2547__, new_new_n2548__, new_new_n2549__,
    new_new_n2550__, new_new_n2551__, new_new_n2552__, new_new_n2553__,
    new_new_n2554__, new_new_n2555__, new_new_n2556__, new_new_n2557__,
    new_new_n2558__, new_new_n2559__, new_new_n2560__, new_new_n2561__,
    new_new_n2562__, new_new_n2563__, new_new_n2564__, new_new_n2565__,
    new_new_n2566__, new_new_n2567__, new_new_n2568__, new_new_n2569__,
    new_new_n2570__, new_new_n2571__, new_new_n2572__, new_new_n2573__,
    new_new_n2574__, new_new_n2575__, new_new_n2576__, new_new_n2577__,
    new_new_n2578__, new_new_n2579__, new_new_n2580__, new_new_n2581__,
    new_new_n2582__, new_new_n2583__, new_new_n2584__, new_new_n2585__,
    new_new_n2586__, new_new_n2587__, new_new_n2588__, new_new_n2589__,
    new_new_n2590__, new_new_n2591__, new_new_n2592__, new_new_n2593__,
    new_new_n2594__, new_new_n2595__, new_new_n2596__, new_new_n2597__,
    new_new_n2598__, new_new_n2599__, new_new_n2600__, new_new_n2601__,
    new_new_n2602__, new_new_n2603__, new_new_n2604__, new_new_n2605__,
    new_new_n2606__, new_new_n2607__, new_new_n2608__, new_new_n2609__,
    new_new_n2610__, new_new_n2611__, new_new_n2612__, new_new_n2613__,
    new_new_n2614__, new_new_n2615__, new_new_n2616__, new_new_n2617__,
    new_new_n2618__, new_new_n2619__, new_new_n2620__, new_new_n2621__,
    new_new_n2622__, new_new_n2623__, new_new_n2624__, new_new_n2625__,
    new_new_n2626__, new_new_n2627__, new_new_n2628__, new_new_n2629__,
    new_new_n2630__, new_new_n2631__, new_new_n2632__, new_new_n2633__,
    new_new_n2634__, new_new_n2635__, new_new_n2636__, new_new_n2637__,
    new_new_n2638__, new_new_n2639__, new_new_n2640__, new_new_n2641__,
    new_new_n2642__, new_new_n2643__, new_new_n2644__, new_new_n2645__,
    new_new_n2646__, new_new_n2647__, new_new_n2648__, new_new_n2649__,
    new_new_n2650__, new_new_n2651__, new_new_n2652__, new_new_n2653__,
    new_new_n2654__, new_new_n2655__, new_new_n2656__, new_new_n2657__,
    new_new_n2658__, new_new_n2659__, new_new_n2660__, new_new_n2661__,
    new_new_n2662__, new_new_n2663__, new_new_n2664__, new_new_n2665__,
    new_new_n2666__, new_new_n2667__, new_new_n2668__, new_new_n2669__,
    new_new_n2670__, new_new_n2671__, new_new_n2672__, new_new_n2673__,
    new_new_n2674__, new_new_n2675__, new_new_n2676__, new_new_n2677__,
    new_new_n2678__, new_new_n2679__, new_new_n2680__, new_new_n2681__,
    new_new_n2682__, new_new_n2683__, new_new_n2684__, new_new_n2685__,
    new_new_n2686__, new_new_n2687__, new_new_n2688__, new_new_n2689__,
    new_new_n2690__, new_new_n2691__, new_new_n2692__, new_new_n2693__,
    new_new_n2694__, new_new_n2695__, new_new_n2696__, new_new_n2697__,
    new_new_n2698__, new_new_n2699__, new_new_n2700__, new_new_n2701__,
    new_new_n2702__, new_new_n2703__, new_new_n2704__, new_new_n2705__,
    new_new_n2706__, new_new_n2707__, new_new_n2708__, new_new_n2709__,
    new_new_n2710__, new_new_n2711__, new_new_n2712__, new_new_n2713__,
    new_new_n2714__, new_new_n2715__, new_new_n2716__, new_new_n2717__,
    new_new_n2718__, new_new_n2719__, new_new_n2720__, new_new_n2721__,
    new_new_n2722__, new_new_n2723__, new_new_n2724__, new_new_n2725__,
    new_new_n2726__, new_new_n2727__, new_new_n2728__, new_new_n2729__,
    new_new_n2730__, new_new_n2731__, new_new_n2732__, new_new_n2733__,
    new_new_n2734__, new_new_n2735__, new_new_n2736__, new_new_n2737__,
    new_new_n2738__, new_new_n2739__, new_new_n2740__, new_new_n2741__,
    new_new_n2742__, new_new_n2743__, new_new_n2744__, new_new_n2745__,
    new_new_n2746__, new_new_n2747__, new_new_n2748__, new_new_n2749__,
    new_new_n2750__, new_new_n2751__, new_new_n2752__, new_new_n2753__,
    new_new_n2754__, new_new_n2755__, new_new_n2756__, new_new_n2757__,
    new_new_n2758__, new_new_n2759__, new_new_n2760__, new_new_n2761__,
    new_new_n2762__, new_new_n2763__, new_new_n2764__, new_new_n2765__,
    new_new_n2766__, new_new_n2767__, new_new_n2768__, new_new_n2769__,
    new_new_n2770__, new_new_n2771__, new_new_n2772__, new_new_n2773__,
    new_new_n2774__, new_new_n2775__, new_new_n2776__, new_new_n2777__,
    new_new_n2778__, new_new_n2779__, new_new_n2780__, new_new_n2781__,
    new_new_n2782__, new_new_n2783__, new_new_n2784__, new_new_n2785__,
    new_new_n2786__, new_new_n2787__, new_new_n2788__, new_new_n2789__,
    new_new_n2790__, new_new_n2791__, new_new_n2792__, new_new_n2793__,
    new_new_n2794__, new_new_n2795__, new_new_n2796__, new_new_n2797__,
    new_new_n2798__, new_new_n2799__, new_new_n2800__, new_new_n2801__,
    new_new_n2802__, new_new_n2803__, new_new_n2804__, new_new_n2805__,
    new_new_n2806__, new_new_n2807__, new_new_n2808__, new_new_n2809__,
    new_new_n2810__, new_new_n2811__, new_new_n2812__, new_new_n2813__,
    new_new_n2814__, new_new_n2815__, new_new_n2816__, new_new_n2817__,
    new_new_n2818__, new_new_n2819__, new_new_n2820__, new_new_n2821__,
    new_new_n2822__, new_new_n2823__, new_new_n2824__, new_new_n2825__,
    new_new_n2826__, new_new_n2827__, new_new_n2828__, new_new_n2829__,
    new_new_n2830__, new_new_n2831__, new_new_n2832__, new_new_n2833__,
    new_new_n2834__, new_new_n2835__, new_new_n2836__, new_new_n2837__,
    new_new_n2838__, new_new_n2839__, new_new_n2840__, new_new_n2841__,
    new_new_n2842__, new_new_n2843__, new_new_n2844__, new_new_n2845__,
    new_new_n2846__, new_new_n2847__, new_new_n2848__, new_new_n2849__,
    new_new_n2850__, new_new_n2851__, new_new_n2852__, new_new_n2853__,
    new_new_n2854__, new_new_n2855__, new_new_n2856__, new_new_n2857__,
    new_new_n2858__, new_new_n2859__, new_new_n2860__, new_new_n2861__,
    new_new_n2862__, new_new_n2863__, new_new_n2864__, new_new_n2865__,
    new_new_n2866__, new_new_n2867__, new_new_n2868__, new_new_n2869__,
    new_new_n2870__, new_new_n2871__, new_new_n2872__, new_new_n2873__,
    new_new_n2874__, new_new_n2875__, new_new_n2876__, new_new_n2877__,
    new_new_n2878__, new_new_n2879__, new_new_n2880__, new_new_n2881__,
    new_new_n2882__, new_new_n2883__, new_new_n2884__, new_new_n2885__,
    new_new_n2886__, new_new_n2887__, new_new_n2888__, new_new_n2889__,
    new_new_n2890__, new_new_n2891__, new_new_n2892__, new_new_n2893__,
    new_new_n2894__, new_new_n2895__, new_new_n2896__, new_new_n2897__,
    new_new_n2898__, new_new_n2899__, new_new_n2900__, new_new_n2901__,
    new_new_n2902__, new_new_n2903__, new_new_n2904__, new_new_n2905__,
    new_new_n2906__, new_new_n2907__, new_new_n2908__, new_new_n2909__,
    new_new_n2910__, new_new_n2911__, new_new_n2912__, new_new_n2913__,
    new_new_n2914__, new_new_n2915__, new_new_n2916__, new_new_n2917__,
    new_new_n2918__, new_new_n2919__, new_new_n2920__, new_new_n2921__,
    new_new_n2922__, new_new_n2923__, new_new_n2924__, new_new_n2925__,
    new_new_n2926__, new_new_n2927__, new_new_n2928__, new_new_n2929__,
    new_new_n2930__, new_new_n2931__, new_new_n2932__, new_new_n2933__,
    new_new_n2934__, new_new_n2935__, new_new_n2936__, new_new_n2937__,
    new_new_n2938__, new_new_n2939__, new_new_n2940__, new_new_n2941__,
    new_new_n2942__, new_new_n2943__, new_new_n2944__, new_new_n2945__,
    new_new_n2946__, new_new_n2947__, new_new_n2948__, new_new_n2949__,
    new_new_n2950__, new_new_n2951__, new_new_n2952__, new_new_n2953__,
    new_new_n2954__, new_new_n2955__, new_new_n2956__, new_new_n2957__,
    new_new_n2958__, new_new_n2959__, new_new_n2960__, new_new_n2961__,
    new_new_n2962__, new_new_n2963__, new_new_n2964__, new_new_n2965__,
    new_new_n2966__, new_new_n2967__, new_new_n2968__, new_new_n2969__,
    new_new_n2970__, new_new_n2971__, new_new_n2972__, new_new_n2973__,
    new_new_n2974__, new_new_n2975__, new_new_n2976__, new_new_n2977__,
    new_new_n2978__, new_new_n2979__, new_new_n2980__, new_new_n2981__,
    new_new_n2982__, new_new_n2983__, new_new_n2984__, new_new_n2985__,
    new_new_n2986__, new_new_n2987__, new_new_n2988__, new_new_n2989__,
    new_new_n2990__, new_new_n2991__, new_new_n2992__, new_new_n2993__,
    new_new_n2994__, new_new_n2995__, new_new_n2996__, new_new_n2997__,
    new_new_n2998__, new_new_n2999__, new_new_n3000__, new_new_n3001__,
    new_new_n3002__, new_new_n3003__, new_new_n3004__, new_new_n3005__,
    new_new_n3006__, new_new_n3007__, new_new_n3008__, new_new_n3009__,
    new_new_n3010__, new_new_n3011__, new_new_n3012__, new_new_n3013__,
    new_new_n3014__, new_new_n3015__, new_new_n3016__, new_new_n3017__,
    new_new_n3018__, new_new_n3019__, new_new_n3020__, new_new_n3021__,
    new_new_n3022__, new_new_n3023__, new_new_n3024__, new_new_n3025__,
    new_new_n3026__, new_new_n3027__, new_new_n3028__, new_new_n3029__,
    new_new_n3030__, new_new_n3031__, new_new_n3032__, new_new_n3033__,
    new_new_n3034__, new_new_n3035__, new_new_n3036__, new_new_n3037__,
    new_new_n3038__, new_new_n3039__, new_new_n3040__, new_new_n3041__,
    new_new_n3042__, new_new_n3043__, new_new_n3044__, new_new_n3045__,
    new_new_n3046__, new_new_n3047__, new_new_n3048__, new_new_n3049__,
    new_new_n3050__, new_new_n3051__, new_new_n3052__, new_new_n3053__,
    new_new_n3054__, new_new_n3055__, new_new_n3056__, new_new_n3057__,
    new_new_n3058__, new_new_n3059__, new_new_n3060__, new_new_n3061__,
    new_new_n3062__, new_new_n3063__, new_new_n3064__, new_new_n3065__,
    new_new_n3066__, new_new_n3067__, new_new_n3068__, new_new_n3069__,
    new_new_n3070__, new_new_n3071__, new_new_n3072__, new_new_n3073__,
    new_new_n3074__, new_new_n3075__, new_new_n3076__, new_new_n3077__,
    new_new_n3078__, new_new_n3079__, new_new_n3080__, new_new_n3081__,
    new_new_n3082__, new_new_n3083__, new_new_n3084__, new_new_n3085__,
    new_new_n3086__, new_new_n3087__, new_new_n3088__, new_new_n3089__,
    new_new_n3090__, new_new_n3091__, new_new_n3092__, new_new_n3093__,
    new_new_n3094__, new_new_n3095__, new_new_n3096__, new_new_n3097__,
    new_new_n3098__, new_new_n3099__, new_new_n3100__, new_new_n3101__,
    new_new_n3102__, new_new_n3103__, new_new_n3104__, new_new_n3105__,
    new_new_n3106__, new_new_n3107__, new_new_n3108__, new_new_n3109__,
    new_new_n3110__, new_new_n3111__, new_new_n3112__, new_new_n3113__,
    new_new_n3114__, new_new_n3115__, new_new_n3116__, new_new_n3117__,
    new_new_n3118__, new_new_n3119__, new_new_n3120__, new_new_n3121__,
    new_new_n3122__, new_new_n3123__, new_new_n3124__, new_new_n3125__,
    new_new_n3126__, new_new_n3127__, new_new_n3128__, new_new_n3129__,
    new_new_n3130__, new_new_n3131__, new_new_n3132__, new_new_n3133__,
    new_new_n3134__, new_new_n3135__, new_new_n3136__, new_new_n3137__,
    new_new_n3138__, new_new_n3139__, new_new_n3140__, new_new_n3141__,
    new_new_n3142__, new_new_n3143__, new_new_n3144__, new_new_n3145__,
    new_new_n3146__, new_new_n3147__, new_new_n3148__, new_new_n3149__,
    new_new_n3150__, new_new_n3151__, new_new_n3152__, new_new_n3153__,
    new_new_n3154__, new_new_n3155__, new_new_n3156__, new_new_n3157__,
    new_new_n3158__, new_new_n3159__, new_new_n3160__, new_new_n3161__,
    new_new_n3162__, new_new_n3163__, new_new_n3164__, new_new_n3165__,
    new_new_n3166__, new_new_n3167__, new_new_n3168__, new_new_n3169__,
    new_new_n3170__, new_new_n3171__, new_new_n3172__, new_new_n3173__,
    new_new_n3174__, new_new_n3175__, new_new_n3176__, new_new_n3177__,
    new_new_n3178__, new_new_n3179__, new_new_n3180__, new_new_n3181__,
    new_new_n3182__, new_new_n3183__, new_new_n3184__, new_new_n3185__,
    new_new_n3186__, new_new_n3187__, new_new_n3188__, new_new_n3189__,
    new_new_n3190__, new_new_n3191__, new_new_n3192__, new_new_n3193__,
    new_new_n3194__, new_new_n3195__, new_new_n3196__, new_new_n3197__,
    new_new_n3198__, new_new_n3199__, new_new_n3200__, new_new_n3201__,
    new_new_n3202__, new_new_n3203__, new_new_n3204__, new_new_n3205__,
    new_new_n3206__, new_new_n3207__, new_new_n3208__, new_new_n3209__,
    new_new_n3210__, new_new_n3211__, new_new_n3212__, new_new_n3213__,
    new_new_n3214__, new_new_n3215__, new_new_n3216__, new_new_n3217__,
    new_new_n3218__, new_new_n3219__, new_new_n3220__, new_new_n3221__,
    new_new_n3222__, new_new_n3223__, new_new_n3224__, new_new_n3225__,
    new_new_n3226__, new_new_n3227__, new_new_n3228__, new_new_n3229__,
    new_new_n3230__, new_new_n3231__, new_new_n3232__, new_new_n3233__,
    new_new_n3234__, new_new_n3235__, new_new_n3236__, new_new_n3237__,
    new_new_n3238__, new_new_n3239__, new_new_n3240__, new_new_n3241__,
    new_new_n3242__, new_new_n3243__, new_new_n3244__, new_new_n3245__,
    new_new_n3246__, new_new_n3247__, new_new_n3248__, new_new_n3249__,
    new_new_n3250__, new_new_n3251__, new_new_n3252__, new_new_n3253__,
    new_new_n3254__, new_new_n3255__, new_new_n3256__, new_new_n3257__,
    new_new_n3258__, new_new_n3259__, new_new_n3260__, new_new_n3261__,
    new_new_n3262__, new_new_n3263__, new_new_n3264__, new_new_n3265__,
    new_new_n3266__, new_new_n3267__, new_new_n3268__, new_new_n3269__,
    new_new_n3270__, new_new_n3271__, new_new_n3272__, new_new_n3273__,
    new_new_n3274__, new_new_n3275__, new_new_n3276__, new_new_n3277__,
    new_new_n3278__, new_new_n3279__, new_new_n3280__, new_new_n3281__,
    new_new_n3282__, new_new_n3283__, new_new_n3284__, new_new_n3285__,
    new_new_n3286__, new_new_n3287__, new_new_n3288__, new_new_n3289__,
    new_new_n3290__, new_new_n3291__, new_new_n3292__, new_new_n3293__,
    new_new_n3294__, new_new_n3295__, new_new_n3296__, new_new_n3297__,
    new_new_n3298__, new_new_n3299__, new_new_n3300__, new_new_n3301__,
    new_new_n3302__, new_new_n3303__, new_new_n3304__, new_new_n3305__,
    new_new_n3306__, new_new_n3307__, new_new_n3308__, new_new_n3309__,
    new_new_n3310__, new_new_n3311__, new_new_n3312__, new_new_n3313__,
    new_new_n3314__, new_new_n3315__, new_new_n3316__, new_new_n3317__,
    new_new_n3318__, new_new_n3319__, new_new_n3320__, new_new_n3321__,
    new_new_n3322__, new_new_n3323__, new_new_n3324__, new_new_n3325__,
    new_new_n3326__, new_new_n3327__, new_new_n3328__, new_new_n3329__,
    new_new_n3330__, new_new_n3331__, new_new_n3332__, new_new_n3333__,
    new_new_n3334__, new_new_n3335__, new_new_n3336__, new_new_n3337__,
    new_new_n3338__, new_new_n3339__, new_new_n3340__, new_new_n3341__,
    new_new_n3342__, new_new_n3343__, new_new_n3344__, new_new_n3345__,
    new_new_n3346__, new_new_n3347__, new_new_n3348__, new_new_n3349__,
    new_new_n3350__, new_new_n3351__, new_new_n3352__, new_new_n3353__,
    new_new_n3354__, new_new_n3355__, new_new_n3356__, new_new_n3357__,
    new_new_n3358__, new_new_n3359__, new_new_n3360__, new_new_n3361__,
    new_new_n3362__, new_new_n3363__, new_new_n3364__, new_new_n3365__,
    new_new_n3366__, new_new_n3367__, new_new_n3368__, new_new_n3369__,
    new_new_n3370__, new_new_n3371__, new_new_n3372__, new_new_n3373__,
    new_new_n3374__, new_new_n3375__, new_new_n3376__, new_new_n3377__,
    new_new_n3378__, new_new_n3379__, new_new_n3380__, new_new_n3381__,
    new_new_n3382__, new_new_n3383__, new_new_n3384__, new_new_n3385__,
    new_new_n3386__, new_new_n3387__, new_new_n3388__, new_new_n3389__,
    new_new_n3390__, new_new_n3391__, new_new_n3392__, new_new_n3393__,
    new_new_n3394__, new_new_n3395__, new_new_n3396__, new_new_n3397__,
    new_new_n3398__, new_new_n3399__, new_new_n3400__, new_new_n3401__,
    new_new_n3402__, new_new_n3403__, new_new_n3404__, new_new_n3405__,
    new_new_n3406__, new_new_n3407__, new_new_n3408__, new_new_n3409__,
    new_new_n3410__, new_new_n3411__, new_new_n3412__, new_new_n3413__,
    new_new_n3414__, new_new_n3415__, new_new_n3416__, new_new_n3417__,
    new_new_n3418__, new_new_n3419__, new_new_n3420__, new_new_n3421__,
    new_new_n3422__, new_new_n3423__, new_new_n3424__, new_new_n3425__,
    new_new_n3426__, new_new_n3427__, new_new_n3428__, new_new_n3429__,
    new_new_n3430__, new_new_n3431__, new_new_n3432__, new_new_n3433__,
    new_new_n3434__, new_new_n3435__, new_new_n3436__, new_new_n3437__,
    new_new_n3438__, new_new_n3439__, new_new_n3440__, new_new_n3441__,
    new_new_n3442__, new_new_n3443__, new_new_n3444__, new_new_n3445__,
    new_new_n3446__, new_new_n3447__, new_new_n3448__, new_new_n3449__,
    new_new_n3450__, new_new_n3451__, new_new_n3452__, new_new_n3453__,
    new_new_n3454__, new_new_n3455__, new_new_n3456__, new_new_n3457__,
    new_new_n3458__, new_new_n3459__, new_new_n3460__, new_new_n3461__,
    new_new_n3462__, new_new_n3463__, new_new_n3464__, new_new_n3465__,
    new_new_n3466__, new_new_n3467__, new_new_n3468__, new_new_n3469__,
    new_new_n3470__, new_new_n3471__, new_new_n3472__, new_new_n3473__,
    new_new_n3474__, new_new_n3475__, new_new_n3476__, new_new_n3477__,
    new_new_n3478__, new_new_n3479__, new_new_n3480__, new_new_n3481__,
    new_new_n3482__, new_new_n3483__, new_new_n3484__, new_new_n3485__,
    new_new_n3486__, new_new_n3487__, new_new_n3488__, new_new_n3489__,
    new_new_n3490__, new_new_n3491__, new_new_n3492__, new_new_n3493__,
    new_new_n3494__, new_new_n3495__, new_new_n3496__, new_new_n3497__,
    new_new_n3498__, new_new_n3499__, new_new_n3500__, new_new_n3501__,
    new_new_n3502__, new_new_n3503__, new_new_n3504__, new_new_n3505__,
    new_new_n3506__, new_new_n3507__, new_new_n3508__, new_new_n3509__,
    new_new_n3510__, new_new_n3511__, new_new_n3512__, new_new_n3513__,
    new_new_n3514__, new_new_n3515__, new_new_n3516__, new_new_n3517__,
    new_new_n3518__, new_new_n3519__, new_new_n3520__, new_new_n3521__,
    new_new_n3522__, new_new_n3523__, new_new_n3524__, new_new_n3525__,
    new_new_n3526__, new_new_n3527__, new_new_n3528__, new_new_n3529__,
    new_new_n3530__, new_new_n3531__, new_new_n3532__, new_new_n3533__,
    new_new_n3534__, new_new_n3535__, new_new_n3536__, new_new_n3537__,
    new_new_n3538__, new_new_n3539__, new_new_n3540__, new_new_n3541__,
    new_new_n3542__, new_new_n3543__, new_new_n3544__, new_new_n3545__,
    new_new_n3546__, new_new_n3547__, new_new_n3548__, new_new_n3549__,
    new_new_n3550__, new_new_n3551__, new_new_n3552__, new_new_n3553__,
    new_new_n3554__, new_new_n3555__, new_new_n3556__, new_new_n3557__,
    new_new_n3558__, new_new_n3559__, new_new_n3560__, new_new_n3561__,
    new_new_n3562__, new_new_n3563__, new_new_n3564__, new_new_n3565__,
    new_new_n3566__, new_new_n3567__, new_new_n3568__, new_new_n3569__,
    new_new_n3570__, new_new_n3571__, new_new_n3572__, new_new_n3573__,
    new_new_n3574__, new_new_n3575__, new_new_n3576__, new_new_n3577__,
    new_new_n3578__, new_new_n3579__, new_new_n3580__, new_new_n3581__,
    new_new_n3582__, new_new_n3583__, new_new_n3584__, new_new_n3585__,
    new_new_n3586__, new_new_n3587__, new_new_n3588__, new_new_n3589__,
    new_new_n3590__, new_new_n3591__, new_new_n3592__, new_new_n3593__,
    new_new_n3594__, new_new_n3595__, new_new_n3596__, new_new_n3597__,
    new_new_n3598__, new_new_n3599__, new_new_n3600__, new_new_n3601__,
    new_new_n3602__, new_new_n3603__, new_new_n3604__, new_new_n3605__,
    new_new_n3606__, new_new_n3607__, new_new_n3608__, new_new_n3609__,
    new_new_n3610__, new_new_n3611__, new_new_n3612__, new_new_n3613__,
    new_new_n3614__, new_new_n3615__, new_new_n3616__, new_new_n3617__,
    new_new_n3618__, new_new_n3619__, new_new_n3620__, new_new_n3621__,
    new_new_n3622__, new_new_n3623__, new_new_n3624__, new_new_n3625__,
    new_new_n3626__, new_new_n3627__, new_new_n3628__, new_new_n3629__,
    new_new_n3630__, new_new_n3631__, new_new_n3632__, new_new_n3633__,
    new_new_n3634__, new_new_n3635__, new_new_n3636__, new_new_n3637__,
    new_new_n3638__, new_new_n3639__, new_new_n3640__, new_new_n3641__,
    new_new_n3642__, new_new_n3643__, new_new_n3644__, new_new_n3645__,
    new_new_n3646__, new_new_n3647__, new_new_n3648__, new_new_n3649__,
    new_new_n3650__, new_new_n3651__, new_new_n3652__, new_new_n3653__,
    new_new_n3654__, new_new_n3655__, new_new_n3656__, new_new_n3657__,
    new_new_n3658__, new_new_n3659__, new_new_n3660__, new_new_n3661__,
    new_new_n3662__, new_new_n3663__, new_new_n3664__, new_new_n3665__,
    new_new_n3666__, new_new_n3667__, new_new_n3668__, new_new_n3669__,
    new_new_n3670__, new_new_n3671__, new_new_n3672__, new_new_n3673__,
    new_new_n3674__, new_new_n3675__, new_new_n3676__, new_new_n3677__,
    new_new_n3678__, new_new_n3679__, new_new_n3680__, new_new_n3681__,
    new_new_n3682__, new_new_n3683__, new_new_n3684__, new_new_n3685__,
    new_new_n3686__, new_new_n3687__, new_new_n3688__, new_new_n3689__,
    new_new_n3690__, new_new_n3691__, new_new_n3692__, new_new_n3693__,
    new_new_n3694__, new_new_n3695__, new_new_n3696__, new_new_n3697__,
    new_new_n3698__, new_new_n3699__, new_new_n3700__, new_new_n3701__,
    new_new_n3702__, new_new_n3703__, new_new_n3704__, new_new_n3705__,
    new_new_n3706__, new_new_n3707__, new_new_n3708__, new_new_n3709__,
    new_new_n3710__, new_new_n3711__, new_new_n3712__, new_new_n3713__,
    new_new_n3714__, new_new_n3715__, new_new_n3716__, new_new_n3717__,
    new_new_n3718__, new_new_n3719__, new_new_n3720__, new_new_n3721__,
    new_new_n3722__, new_new_n3723__, new_new_n3724__, new_new_n3725__,
    new_new_n3726__, new_new_n3727__, new_new_n3728__, new_new_n3729__,
    new_new_n3730__, new_new_n3731__, new_new_n3732__, new_new_n3733__,
    new_new_n3734__, new_new_n3735__, new_new_n3736__, new_new_n3737__,
    new_new_n3738__, new_new_n3739__, new_new_n3740__, new_new_n3741__,
    new_new_n3742__, new_new_n3743__, new_new_n3744__, new_new_n3745__,
    new_new_n3746__, new_new_n3747__, new_new_n3748__, new_new_n3749__,
    new_new_n3750__, new_new_n3751__, new_new_n3752__, new_new_n3753__,
    new_new_n3754__, new_new_n3755__, new_new_n3756__, new_new_n3757__,
    new_new_n3758__, new_new_n3759__, new_new_n3760__, new_new_n3761__,
    new_new_n3762__, new_new_n3763__, new_new_n3764__, new_new_n3765__,
    new_new_n3766__, new_new_n3767__, new_new_n3768__, new_new_n3769__,
    new_new_n3770__, new_new_n3771__, new_new_n3772__, new_new_n3773__,
    new_new_n3774__, new_new_n3775__, new_new_n3776__, new_new_n3777__,
    new_new_n3778__, new_new_n3779__, new_new_n3780__, new_new_n3781__,
    new_new_n3782__, new_new_n3783__, new_new_n3784__, new_new_n3785__,
    new_new_n3786__, new_new_n3787__, new_new_n3788__, new_new_n3789__,
    new_new_n3790__, new_new_n3791__, new_new_n3792__, new_new_n3793__,
    new_new_n3794__, new_new_n3795__, new_new_n3796__, new_new_n3797__,
    new_new_n3798__, new_new_n3799__, new_new_n3800__, new_new_n3801__,
    new_new_n3802__, new_new_n3803__, new_new_n3804__, new_new_n3805__,
    new_new_n3806__, new_new_n3807__, new_new_n3808__, new_new_n3809__,
    new_new_n3810__, new_new_n3811__, new_new_n3812__, new_new_n3813__,
    new_new_n3814__, new_new_n3815__, new_new_n3816__, new_new_n3817__,
    new_new_n3818__, new_new_n3819__, new_new_n3820__, new_new_n3821__,
    new_new_n3822__, new_new_n3823__, new_new_n3824__, new_new_n3825__,
    new_new_n3826__, new_new_n3827__, new_new_n3828__, new_new_n3829__,
    new_new_n3830__, new_new_n3831__, new_new_n3832__, new_new_n3833__,
    new_new_n3834__, new_new_n3835__, new_new_n3836__, new_new_n3837__,
    new_new_n3838__, new_new_n3839__, new_new_n3840__, new_new_n3841__,
    new_new_n3842__, new_new_n3843__, new_new_n3844__, new_new_n3845__,
    new_new_n3846__, new_new_n3847__, new_new_n3848__, new_new_n3849__,
    new_new_n3850__, new_new_n3851__, new_new_n3852__, new_new_n3853__,
    new_new_n3854__, new_new_n3855__, new_new_n3856__, new_new_n3857__,
    new_new_n3858__, new_new_n3859__, new_new_n3860__, new_new_n3861__,
    new_new_n3862__, new_new_n3863__, new_new_n3864__, new_new_n3865__,
    new_new_n3866__, new_new_n3867__, new_new_n3868__, new_new_n3869__,
    new_new_n3870__, new_new_n3871__, new_new_n3872__, new_new_n3873__,
    new_new_n3874__, new_new_n3875__, new_new_n3876__, new_new_n3877__,
    new_new_n3878__, new_new_n3879__, new_new_n3880__, new_new_n3881__,
    new_new_n3882__, new_new_n3883__, new_new_n3884__, new_new_n3885__,
    new_new_n3886__, new_new_n3887__, new_new_n3888__, new_new_n3889__,
    new_new_n3890__, new_new_n3891__, new_new_n3892__, new_new_n3893__,
    new_new_n3894__, new_new_n3895__, new_new_n3896__, new_new_n3897__,
    new_new_n3898__, new_new_n3899__, new_new_n3900__, new_new_n3901__,
    new_new_n3902__, new_new_n3903__, new_new_n3904__, new_new_n3905__,
    new_new_n3906__, new_new_n3907__, new_new_n3908__, new_new_n3909__,
    new_new_n3910__, new_new_n3911__, new_new_n3912__, new_new_n3913__,
    new_new_n3914__, new_new_n3915__, new_new_n3916__, new_new_n3917__,
    new_new_n3918__, new_new_n3919__, new_new_n3920__, new_new_n3921__,
    new_new_n3922__, new_new_n3923__, new_new_n3924__, new_new_n3925__,
    new_new_n3926__, new_new_n3927__, new_new_n3928__, new_new_n3929__,
    new_new_n3930__, new_new_n3931__, new_new_n3932__, new_new_n3933__,
    new_new_n3934__, new_new_n3935__, new_new_n3936__, new_new_n3937__,
    new_new_n3938__, new_new_n3939__, new_new_n3940__, new_new_n3941__,
    new_new_n3942__, new_new_n3943__, new_new_n3944__, new_new_n3945__,
    new_new_n3946__, new_new_n3947__, new_new_n3948__, new_new_n3949__,
    new_new_n3950__, new_new_n3951__, new_new_n3952__, new_new_n3953__,
    new_new_n3954__, new_new_n3955__, new_new_n3956__, new_new_n3957__,
    new_new_n3958__, new_new_n3959__, new_new_n3960__, new_new_n3961__,
    new_new_n3962__, new_new_n3963__, new_new_n3964__, new_new_n3965__,
    new_new_n3966__, new_new_n3967__, new_new_n3968__, new_new_n3969__,
    new_new_n3970__, new_new_n3971__, new_new_n3972__, new_new_n3973__,
    new_new_n3974__, new_new_n3975__, new_new_n3976__, new_new_n3977__,
    new_new_n3978__, new_new_n3979__, new_new_n3980__, new_new_n3981__,
    new_new_n3982__, new_new_n3983__, new_new_n3984__, new_new_n3985__,
    new_new_n3986__, new_new_n3987__, new_new_n3988__, new_new_n3989__,
    new_new_n3990__, new_new_n3991__, new_new_n3992__, new_new_n3993__,
    new_new_n3994__, new_new_n3995__, new_new_n3996__, new_new_n3997__,
    new_new_n3998__, new_new_n3999__, new_new_n4000__, new_new_n4001__,
    new_new_n4002__, new_new_n4003__, new_new_n4004__, new_new_n4005__,
    new_new_n4006__, new_new_n4007__, new_new_n4008__, new_new_n4009__,
    new_new_n4010__, new_new_n4011__, new_new_n4012__, new_new_n4013__,
    new_new_n4014__, new_new_n4015__, new_new_n4016__, new_new_n4017__,
    new_new_n4018__, new_new_n4019__, new_new_n4020__, new_new_n4021__,
    new_new_n4022__, new_new_n4023__, new_new_n4024__, new_new_n4025__,
    new_new_n4026__, new_new_n4027__, new_new_n4028__, new_new_n4029__,
    new_new_n4030__, new_new_n4031__, new_new_n4032__, new_new_n4033__,
    new_new_n4034__, new_new_n4035__, new_new_n4036__, new_new_n4037__,
    new_new_n4038__, new_new_n4039__, new_new_n4040__, new_new_n4041__,
    new_new_n4042__, new_new_n4043__, new_new_n4044__, new_new_n4045__,
    new_new_n4046__, new_new_n4047__, new_new_n4048__, new_new_n4049__,
    new_new_n4050__, new_new_n4051__, new_new_n4052__, new_new_n4053__,
    new_new_n4054__, new_new_n4055__, new_new_n4056__, new_new_n4057__,
    new_new_n4058__, new_new_n4059__, new_new_n4060__, new_new_n4061__,
    new_new_n4062__, new_new_n4063__, new_new_n4064__, new_new_n4065__,
    new_new_n4066__, new_new_n4067__, new_new_n4068__, new_new_n4069__,
    new_new_n4070__, new_new_n4071__, new_new_n4072__, new_new_n4073__,
    new_new_n4074__, new_new_n4075__, new_new_n4076__, new_new_n4077__,
    new_new_n4078__, new_new_n4079__, new_new_n4080__, new_new_n4081__,
    new_new_n4082__, new_new_n4083__, new_new_n4084__, new_new_n4085__,
    new_new_n4086__, new_new_n4087__, new_new_n4088__, new_new_n4089__,
    new_new_n4090__, new_new_n4091__, new_new_n4092__, new_new_n4093__,
    new_new_n4094__, new_new_n4095__, new_new_n4096__, new_new_n4097__,
    new_new_n4098__, new_new_n4099__, new_new_n4100__, new_new_n4101__,
    new_new_n4102__, new_new_n4103__, new_new_n4104__, new_new_n4105__,
    new_new_n4106__, new_new_n4107__, new_new_n4108__, new_new_n4109__,
    new_new_n4110__, new_new_n4111__, new_new_n4112__, new_new_n4113__,
    new_new_n4114__, new_new_n4115__, new_new_n4116__, new_new_n4117__,
    new_new_n4118__, new_new_n4119__, new_new_n4120__, new_new_n4121__,
    new_new_n4122__, new_new_n4123__, new_new_n4124__, new_new_n4125__,
    new_new_n4126__, new_new_n4127__, new_new_n4128__, new_new_n4129__,
    new_new_n4130__, new_new_n4131__, new_new_n4132__, new_new_n4133__,
    new_new_n4134__, new_new_n4135__, new_new_n4136__, new_new_n4137__,
    new_new_n4138__, new_new_n4139__, new_new_n4140__, new_new_n4141__,
    new_new_n4142__, new_new_n4143__, new_new_n4144__, new_new_n4145__,
    new_new_n4146__, new_new_n4147__, new_new_n4148__, new_new_n4149__,
    new_new_n4150__, new_new_n4151__, new_new_n4152__, new_new_n4153__,
    new_new_n4154__, new_new_n4155__, new_new_n4156__, new_new_n4157__,
    new_new_n4158__, new_new_n4159__, new_new_n4160__, new_new_n4161__,
    new_new_n4162__, new_new_n4163__, new_new_n4164__, new_new_n4165__,
    new_new_n4166__, new_new_n4167__, new_new_n4168__, new_new_n4169__,
    new_new_n4170__, new_new_n4171__, new_new_n4172__, new_new_n4173__,
    new_new_n4174__, new_new_n4175__, new_new_n4176__, new_new_n4177__,
    new_new_n4178__, new_new_n4179__, new_new_n4180__, new_new_n4181__,
    new_new_n4182__, new_new_n4183__, new_new_n4184__, new_new_n4185__,
    new_new_n4186__, new_new_n4187__, new_new_n4188__, new_new_n4189__,
    new_new_n4190__, new_new_n4191__, new_new_n4192__, new_new_n4193__,
    new_new_n4194__, new_new_n4195__, new_new_n4196__, new_new_n4197__,
    new_new_n4198__, new_new_n4199__, new_new_n4200__, new_new_n4201__,
    new_new_n4202__, new_new_n4203__, new_new_n4204__, new_new_n4205__,
    new_new_n4206__, new_new_n4207__, new_new_n4208__, new_new_n4209__,
    new_new_n4210__, new_new_n4211__, new_new_n4212__, new_new_n4213__,
    new_new_n4214__, new_new_n4215__, new_new_n4216__, new_new_n4217__,
    new_new_n4218__, new_new_n4219__, new_new_n4220__, new_new_n4221__,
    new_new_n4222__, new_new_n4223__, new_new_n4224__, new_new_n4225__,
    new_new_n4226__, new_new_n4227__, new_new_n4228__, new_new_n4229__,
    new_new_n4230__, new_new_n4231__, new_new_n4232__, new_new_n4233__,
    new_new_n4234__, new_new_n4235__, new_new_n4236__, new_new_n4237__,
    new_new_n4238__, new_new_n4239__, new_new_n4240__, new_new_n4241__,
    new_new_n4242__, new_new_n4243__, new_new_n4244__, new_new_n4245__,
    new_new_n4246__, new_new_n4247__, new_new_n4248__, new_new_n4249__,
    new_new_n4250__, new_new_n4251__, new_new_n4252__, new_new_n4253__,
    new_new_n4254__, new_new_n4255__, new_new_n4256__, new_new_n4257__,
    new_new_n4258__, new_new_n4259__, new_new_n4260__, new_new_n4261__,
    new_new_n4262__, new_new_n4263__, new_new_n4264__, new_new_n4265__,
    new_new_n4266__, new_new_n4267__, new_new_n4268__, new_new_n4269__,
    new_new_n4270__, new_new_n4271__, new_new_n4272__, new_new_n4273__,
    new_new_n4274__, new_new_n4275__, new_new_n4276__, new_new_n4277__,
    new_new_n4278__, new_new_n4279__, new_new_n4280__, new_new_n4281__,
    new_new_n4282__, new_new_n4283__, new_new_n4284__, new_new_n4285__,
    new_new_n4286__, new_new_n4287__, new_new_n4288__, new_new_n4289__,
    new_new_n4290__, new_new_n4291__, new_new_n4292__, new_new_n4293__,
    new_new_n4294__, new_new_n4295__, new_new_n4296__, new_new_n4297__,
    new_new_n4298__, new_new_n4299__, new_new_n4300__, new_new_n4301__,
    new_new_n4302__, new_new_n4303__, new_new_n4304__, new_new_n4305__,
    new_new_n4306__, new_new_n4307__, new_new_n4308__, new_new_n4309__,
    new_new_n4310__, new_new_n4311__, new_new_n4312__, new_new_n4313__,
    new_new_n4314__, new_new_n4315__, new_new_n4316__, new_new_n4317__,
    new_new_n4318__, new_new_n4319__, new_new_n4320__, new_new_n4321__,
    new_new_n4322__, new_new_n4323__, new_new_n4324__, new_new_n4325__,
    new_new_n4326__, new_new_n4327__, new_new_n4328__, new_new_n4329__,
    new_new_n4330__, new_new_n4331__, new_new_n4332__, new_new_n4333__,
    new_new_n4334__, new_new_n4335__, new_new_n4336__, new_new_n4337__,
    new_new_n4338__, new_new_n4339__, new_new_n4340__, new_new_n4341__,
    new_new_n4342__, new_new_n4343__, new_new_n4344__, new_new_n4345__,
    new_new_n4346__, new_new_n4347__, new_new_n4348__, new_new_n4349__,
    new_new_n4350__, new_new_n4351__, new_new_n4352__, new_new_n4353__,
    new_new_n4354__, new_new_n4355__, new_new_n4356__, new_new_n4357__,
    new_new_n4358__, new_new_n4359__, new_new_n4360__, new_new_n4361__,
    new_new_n4362__, new_new_n4363__, new_new_n4364__, new_new_n4365__,
    new_new_n4366__, new_new_n4367__, new_new_n4368__, new_new_n4369__,
    new_new_n4370__, new_new_n4371__, new_new_n4372__, new_new_n4373__,
    new_new_n4374__, new_new_n4375__, new_new_n4376__, new_new_n4377__,
    new_new_n4378__, new_new_n4379__, new_new_n4380__, new_new_n4381__,
    new_new_n4382__, new_new_n4383__, new_new_n4384__, new_new_n4385__,
    new_new_n4386__, new_new_n4387__, new_new_n4388__, new_new_n4389__,
    new_new_n4390__, new_new_n4391__, new_new_n4392__, new_new_n4393__,
    new_new_n4394__, new_new_n4395__, new_new_n4396__, new_new_n4397__,
    new_new_n4398__, new_new_n4399__, new_new_n4400__, new_new_n4401__,
    new_new_n4402__, new_new_n4403__, new_new_n4404__, new_new_n4405__,
    new_new_n4406__, new_new_n4407__, new_new_n4408__, new_new_n4409__,
    new_new_n4410__, new_new_n4411__, new_new_n4412__, new_new_n4413__,
    new_new_n4414__, new_new_n4415__, new_new_n4416__, new_new_n4417__,
    new_new_n4418__, new_new_n4419__, new_new_n4420__, new_new_n4421__,
    new_new_n4422__, new_new_n4423__, new_new_n4424__, new_new_n4425__,
    new_new_n4426__, new_new_n4427__, new_new_n4428__, new_new_n4429__,
    new_new_n4430__, new_new_n4431__, new_new_n4432__, new_new_n4433__,
    new_new_n4434__, new_new_n4435__, new_new_n4436__, new_new_n4437__,
    new_new_n4438__, new_new_n4439__, new_new_n4440__, new_new_n4441__,
    new_new_n4442__, new_new_n4443__, new_new_n4444__, new_new_n4445__,
    new_new_n4446__, new_new_n4447__, new_new_n4448__, new_new_n4449__,
    new_new_n4450__, new_new_n4451__, new_new_n4452__, new_new_n4453__,
    new_new_n4454__, new_new_n4455__, new_new_n4456__, new_new_n4457__,
    new_new_n4458__, new_new_n4459__, new_new_n4460__, new_new_n4461__,
    new_new_n4462__, new_new_n4463__, new_new_n4464__, new_new_n4465__,
    new_new_n4466__, new_new_n4467__, new_new_n4468__, new_new_n4469__,
    new_new_n4470__, new_new_n4471__, new_new_n4472__, new_new_n4473__,
    new_new_n4474__, new_new_n4475__, new_new_n4476__, new_new_n4477__,
    new_new_n4478__, new_new_n4479__, new_new_n4480__, new_new_n4481__,
    new_new_n4482__, new_new_n4483__, new_new_n4484__, new_new_n4485__,
    new_new_n4486__, new_new_n4487__, new_new_n4488__, new_new_n4489__,
    new_new_n4490__, new_new_n4491__, new_new_n4492__, new_new_n4493__,
    new_new_n4494__, new_new_n4495__, new_new_n4496__, new_new_n4497__,
    new_new_n4498__, new_new_n4499__, new_new_n4500__, new_new_n4501__,
    new_new_n4502__, new_new_n4503__, new_new_n4504__, new_new_n4505__,
    new_new_n4506__, new_new_n4507__, new_new_n4508__, new_new_n4509__,
    new_new_n4510__, new_new_n4511__, new_new_n4512__, new_new_n4513__,
    new_new_n4514__, new_new_n4515__, new_new_n4516__, new_new_n4517__,
    new_new_n4518__, new_new_n4519__, new_new_n4520__, new_new_n4521__,
    new_new_n4522__, new_new_n4523__, new_new_n4524__, new_new_n4525__,
    new_new_n4526__, new_new_n4527__, new_new_n4528__, new_new_n4529__,
    new_new_n4530__, new_new_n4531__, new_new_n4532__, new_new_n4533__,
    new_new_n4534__, new_new_n4535__, new_new_n4536__, new_new_n4537__,
    new_new_n4538__, new_new_n4539__, new_new_n4540__, new_new_n4541__,
    new_new_n4542__, new_new_n4543__, new_new_n4544__, new_new_n4545__,
    new_new_n4546__, new_new_n4547__, new_new_n4548__, new_new_n4549__,
    new_new_n4550__, new_new_n4551__, new_new_n4552__, new_new_n4553__,
    new_new_n4554__, new_new_n4555__, new_new_n4556__, new_new_n4557__,
    new_new_n4558__, new_new_n4559__, new_new_n4560__, new_new_n4561__,
    new_new_n4562__, new_new_n4563__, new_new_n4564__, new_new_n4565__,
    new_new_n4566__, new_new_n4567__, new_new_n4568__, new_new_n4569__,
    new_new_n4570__, new_new_n4571__, new_new_n4572__, new_new_n4573__,
    new_new_n4574__, new_new_n4575__, new_new_n4576__, new_new_n4577__,
    new_new_n4578__, new_new_n4579__, new_new_n4580__, new_new_n4581__,
    new_new_n4582__, new_new_n4583__, new_new_n4584__, new_new_n4585__,
    new_new_n4586__, new_new_n4587__, new_new_n4588__, new_new_n4589__,
    new_new_n4590__, new_new_n4591__, new_new_n4592__, new_new_n4593__,
    new_new_n4594__, new_new_n4595__, new_new_n4596__, new_new_n4597__,
    new_new_n4598__, new_new_n4599__, new_new_n4600__, new_new_n4601__,
    new_new_n4602__, new_new_n4603__, new_new_n4604__, new_new_n4605__,
    new_new_n4606__, new_new_n4607__, new_new_n4608__, new_new_n4609__,
    new_new_n4610__, new_new_n4611__, new_new_n4612__, new_new_n4613__,
    new_new_n4614__, new_new_n4615__, new_new_n4616__, new_new_n4617__,
    new_new_n4618__, new_new_n4619__, new_new_n4620__, new_new_n4621__,
    new_new_n4622__, new_new_n4623__, new_new_n4624__, new_new_n4625__,
    new_new_n4626__, new_new_n4627__, new_new_n4628__, new_new_n4629__,
    new_new_n4630__, new_new_n4631__, new_new_n4632__, new_new_n4633__,
    new_new_n4634__, new_new_n4635__, new_new_n4636__, new_new_n4637__,
    new_new_n4638__, new_new_n4639__, new_new_n4640__, new_new_n4641__,
    new_new_n4642__, new_new_n4643__, new_new_n4644__, new_new_n4645__,
    new_new_n4646__, new_new_n4647__, new_new_n4648__, new_new_n4649__,
    new_new_n4650__, new_new_n4651__, new_new_n4652__, new_new_n4653__,
    new_new_n4654__, new_new_n4655__, new_new_n4656__, new_new_n4657__,
    new_new_n4658__, new_new_n4659__, new_new_n4660__, new_new_n4661__,
    new_new_n4662__, new_new_n4663__, new_new_n4664__, new_new_n4665__,
    new_new_n4666__, new_new_n4667__, new_new_n4668__, new_new_n4669__,
    new_new_n4670__, new_new_n4671__, new_new_n4672__, new_new_n4673__,
    new_new_n4674__, new_new_n4675__, new_new_n4676__, new_new_n4677__,
    new_new_n4678__, new_new_n4679__, new_new_n4680__, new_new_n4681__,
    new_new_n4682__, new_new_n4683__, new_new_n4684__, new_new_n4685__,
    new_new_n4686__, new_new_n4687__, new_new_n4688__, new_new_n4689__,
    new_new_n4690__, new_new_n4691__, new_new_n4692__, new_new_n4693__,
    new_new_n4694__, new_new_n4695__, new_new_n4696__, new_new_n4697__,
    new_new_n4698__, new_new_n4699__, new_new_n4700__, new_new_n4701__,
    new_new_n4702__, new_new_n4703__, new_new_n4704__, new_new_n4705__,
    new_new_n4706__, new_new_n4707__, new_new_n4708__, new_new_n4709__,
    new_new_n4710__, new_new_n4711__, new_new_n4712__, new_new_n4713__,
    new_new_n4714__, new_new_n4715__, new_new_n4716__, new_new_n4717__,
    new_new_n4718__, new_new_n4719__, new_new_n4720__, new_new_n4721__,
    new_new_n4722__, new_new_n4723__, new_new_n4724__, new_new_n4725__,
    new_new_n4726__, new_new_n4727__, new_new_n4728__, new_new_n4729__,
    new_new_n4730__, new_new_n4731__, new_new_n4732__, new_new_n4733__,
    new_new_n4734__, new_new_n4735__, new_new_n4736__, new_new_n4737__,
    new_new_n4738__, new_new_n4739__, new_new_n4740__, new_new_n4741__,
    new_new_n4742__, new_new_n4743__, new_new_n4744__, new_new_n4745__,
    new_new_n4746__, new_new_n4747__, new_new_n4748__, new_new_n4749__,
    new_new_n4750__, new_new_n4751__, new_new_n4752__, new_new_n4753__,
    new_new_n4754__, new_new_n4755__, new_new_n4756__, new_new_n4757__,
    new_new_n4758__, new_new_n4759__, new_new_n4760__, new_new_n4761__,
    new_new_n4762__, new_new_n4763__, new_new_n4764__, new_new_n4765__,
    new_new_n4766__, new_new_n4767__, new_new_n4768__, new_new_n4769__,
    new_new_n4770__, new_new_n4771__, new_new_n4772__, new_new_n4773__,
    new_new_n4774__, new_new_n4775__, new_new_n4776__, new_new_n4777__,
    new_new_n4778__, new_new_n4779__, new_new_n4780__, new_new_n4781__,
    new_new_n4782__, new_new_n4783__, new_new_n4784__, new_new_n4785__,
    new_new_n4786__, new_new_n4787__, new_new_n4788__, new_new_n4789__,
    new_new_n4790__, new_new_n4791__, new_new_n4792__, new_new_n4793__,
    new_new_n4794__, new_new_n4795__, new_new_n4796__, new_new_n4797__,
    new_new_n4798__, new_new_n4799__, new_new_n4800__, new_new_n4801__,
    new_new_n4802__, new_new_n4803__, new_new_n4804__, new_new_n4805__,
    new_new_n4806__, new_new_n4807__, new_new_n4808__, new_new_n4809__,
    new_new_n4810__, new_new_n4811__, new_new_n4812__, new_new_n4813__,
    new_new_n4814__, new_new_n4815__, new_new_n4816__, new_new_n4817__,
    new_new_n4818__, new_new_n4819__, new_new_n4820__, new_new_n4821__,
    new_new_n4822__, new_new_n4823__, new_new_n4824__, new_new_n4825__,
    new_new_n4826__, new_new_n4827__, new_new_n4828__, new_new_n4829__,
    new_new_n4830__, new_new_n4831__, new_new_n4832__, new_new_n4833__,
    new_new_n4834__, new_new_n4835__, new_new_n4836__, new_new_n4837__,
    new_new_n4838__, new_new_n4839__, new_new_n4840__, new_new_n4841__,
    new_new_n4842__, new_new_n4843__, new_new_n4844__, new_new_n4845__,
    new_new_n4846__, new_new_n4847__, new_new_n4848__, new_new_n4849__,
    new_new_n4850__, new_new_n4851__, new_new_n4852__, new_new_n4853__,
    new_new_n4854__, new_new_n4855__, new_new_n4856__, new_new_n4857__,
    new_new_n4858__, new_new_n4859__, new_new_n4860__, new_new_n4861__,
    new_new_n4862__, new_new_n4863__, new_new_n4864__, new_new_n4865__,
    new_new_n4866__, new_new_n4867__, new_new_n4868__, new_new_n4869__,
    new_new_n4870__, new_new_n4871__, new_new_n4872__, new_new_n4873__,
    new_new_n4874__, new_new_n4875__, new_new_n4876__, new_new_n4877__,
    new_new_n4878__, new_new_n4879__, new_new_n4880__, new_new_n4881__,
    new_new_n4882__, new_new_n4883__, new_new_n4884__, new_new_n4885__,
    new_new_n4886__, new_new_n4887__, new_new_n4888__, new_new_n4889__,
    new_new_n4890__, new_new_n4891__, new_new_n4892__, new_new_n4893__,
    new_new_n4894__, new_new_n4895__, new_new_n4896__, new_new_n4897__,
    new_new_n4898__, new_new_n4899__, new_new_n4900__, new_new_n4901__,
    new_new_n4902__, new_new_n4903__, new_new_n4904__, new_new_n4905__,
    new_new_n4906__, new_new_n4907__, new_new_n4908__, new_new_n4909__,
    new_new_n4910__, new_new_n4911__, new_new_n4912__, new_new_n4913__,
    new_new_n4914__, new_new_n4915__, new_new_n4916__, new_new_n4917__,
    new_new_n4918__, new_new_n4919__, new_new_n4920__, new_new_n4921__,
    new_new_n4922__, new_new_n4923__, new_new_n4924__, new_new_n4925__,
    new_new_n4926__, new_new_n4927__, new_new_n4928__, new_new_n4929__,
    new_new_n4930__, new_new_n4931__, new_new_n4932__, new_new_n4933__,
    new_new_n4934__, new_new_n4935__, new_new_n4936__, new_new_n4937__,
    new_new_n4938__, new_new_n4939__, new_new_n4940__, new_new_n4941__,
    new_new_n4942__, new_new_n4943__, new_new_n4944__, new_new_n4945__,
    new_new_n4946__, new_new_n4947__, new_new_n4948__, new_new_n4949__,
    new_new_n4950__, new_new_n4951__, new_new_n4952__, new_new_n4953__,
    new_new_n4954__, new_new_n4955__, new_new_n4956__, new_new_n4957__,
    new_new_n4958__, new_new_n4959__, new_new_n4960__, new_new_n4961__,
    new_new_n4962__, new_new_n4963__, new_new_n4964__, new_new_n4965__,
    new_new_n4966__, new_new_n4967__, new_new_n4968__, new_new_n4969__,
    new_new_n4970__, new_new_n4971__, new_new_n4972__, new_new_n4973__,
    new_new_n4974__, new_new_n4975__, new_new_n4976__, new_new_n4977__,
    new_new_n4978__, new_new_n4979__, new_new_n4980__, new_new_n4981__,
    new_new_n4982__, new_new_n4983__, new_new_n4984__, new_new_n4985__,
    new_new_n4986__, new_new_n4987__, new_new_n4988__, new_new_n4989__,
    new_new_n4990__, new_new_n4991__, new_new_n4992__, new_new_n4993__,
    new_new_n4994__, new_new_n4995__, new_new_n4996__, new_new_n4997__,
    new_new_n4998__, new_new_n4999__, new_new_n5000__, new_new_n5001__,
    new_new_n5002__, new_new_n5003__, new_new_n5004__, new_new_n5005__,
    new_new_n5006__, new_new_n5007__, new_new_n5008__, new_new_n5009__,
    new_new_n5010__, new_new_n5011__, new_new_n5012__, new_new_n5013__,
    new_new_n5014__, new_new_n5015__, new_new_n5016__, new_new_n5017__,
    new_new_n5018__, new_new_n5019__, new_new_n5020__, new_new_n5021__,
    new_new_n5022__, new_new_n5023__, new_new_n5024__, new_new_n5025__,
    new_new_n5026__, new_new_n5027__, new_new_n5028__, new_new_n5029__,
    new_new_n5030__, new_new_n5031__, new_new_n5032__, new_new_n5033__,
    new_new_n5034__, new_new_n5035__, new_new_n5036__, new_new_n5037__,
    new_new_n5038__, new_new_n5039__, new_new_n5040__, new_new_n5041__,
    new_new_n5042__, new_new_n5043__, new_new_n5044__, new_new_n5045__,
    new_new_n5046__, new_new_n5047__, new_new_n5048__, new_new_n5049__,
    new_new_n5050__, new_new_n5051__, new_new_n5052__, new_new_n5053__,
    new_new_n5054__, new_new_n5055__, new_new_n5056__, new_new_n5057__,
    new_new_n5058__, new_new_n5059__, new_new_n5060__, new_new_n5061__,
    new_new_n5062__, new_new_n5063__, new_new_n5064__, new_new_n5065__,
    new_new_n5066__, new_new_n5067__, new_new_n5068__, new_new_n5069__,
    new_new_n5070__, new_new_n5071__, new_new_n5072__, new_new_n5073__,
    new_new_n5074__, new_new_n5075__, new_new_n5076__, new_new_n5077__,
    new_new_n5078__, new_new_n5079__, new_new_n5080__, new_new_n5081__,
    new_new_n5082__, new_new_n5083__, new_new_n5084__, new_new_n5085__,
    new_new_n5086__, new_new_n5087__, new_new_n5088__, new_new_n5089__,
    new_new_n5090__, new_new_n5091__, new_new_n5092__, new_new_n5093__,
    new_new_n5094__, new_new_n5095__, new_new_n5096__, new_new_n5097__,
    new_new_n5098__, new_new_n5099__, new_new_n5100__, new_new_n5101__,
    new_new_n5102__, new_new_n5103__, new_new_n5104__, new_new_n5105__,
    new_new_n5106__, new_new_n5107__, new_new_n5108__, new_new_n5109__,
    new_new_n5110__, new_new_n5111__, new_new_n5112__, new_new_n5113__,
    new_new_n5114__, new_new_n5115__, new_new_n5116__, new_new_n5117__,
    new_new_n5118__, new_new_n5119__, new_new_n5120__, new_new_n5121__,
    new_new_n5122__, new_new_n5123__, new_new_n5124__, new_new_n5125__,
    new_new_n5126__, new_new_n5127__, new_new_n5128__, new_new_n5129__,
    new_new_n5130__, new_new_n5131__, new_new_n5132__, new_new_n5133__,
    new_new_n5134__, new_new_n5135__, new_new_n5136__, new_new_n5137__,
    new_new_n5138__, new_new_n5139__, new_new_n5140__, new_new_n5141__,
    new_new_n5142__, new_new_n5143__, new_new_n5144__, new_new_n5145__,
    new_new_n5146__, new_new_n5147__, new_new_n5148__, new_new_n5149__,
    new_new_n5150__, new_new_n5151__, new_new_n5152__, new_new_n5153__,
    new_new_n5154__, new_new_n5155__, new_new_n5156__, new_new_n5157__,
    new_new_n5158__, new_new_n5159__, new_new_n5160__, new_new_n5161__,
    new_new_n5162__, new_new_n5163__, new_new_n5164__, new_new_n5165__,
    new_new_n5166__, new_new_n5167__, new_new_n5168__, new_new_n5169__,
    new_new_n5170__, new_new_n5171__, new_new_n5172__, new_new_n5173__,
    new_new_n5174__, new_new_n5175__, new_new_n5176__, new_new_n5177__,
    new_new_n5178__, new_new_n5179__, new_new_n5180__, new_new_n5181__,
    new_new_n5182__, new_new_n5183__, new_new_n5184__, new_new_n5185__,
    new_new_n5186__, new_new_n5187__, new_new_n5188__, new_new_n5189__,
    new_new_n5190__, new_new_n5191__, new_new_n5192__, new_new_n5193__,
    new_new_n5194__, new_new_n5195__, new_new_n5196__, new_new_n5197__,
    new_new_n5198__, new_new_n5199__, new_new_n5200__, new_new_n5201__,
    new_new_n5202__, new_new_n5203__, new_new_n5204__, new_new_n5205__,
    new_new_n5206__, new_new_n5207__, new_new_n5208__, new_new_n5209__,
    new_new_n5210__, new_new_n5211__, new_new_n5212__, new_new_n5213__,
    new_new_n5214__, new_new_n5215__, new_new_n5216__, new_new_n5217__,
    new_new_n5218__, new_new_n5219__, new_new_n5220__, new_new_n5221__,
    new_new_n5222__, new_new_n5223__, new_new_n5224__, new_new_n5225__,
    new_new_n5226__, new_new_n5227__, new_new_n5228__, new_new_n5229__,
    new_new_n5230__, new_new_n5231__, new_new_n5232__, new_new_n5233__,
    new_new_n5234__, new_new_n5235__, new_new_n5236__, new_new_n5237__,
    new_new_n5238__, new_new_n5239__, new_new_n5240__, new_new_n5241__,
    new_new_n5242__, new_new_n5243__, new_new_n5244__, new_new_n5245__,
    new_new_n5246__, new_new_n5247__, new_new_n5248__, new_new_n5249__,
    new_new_n5250__, new_new_n5251__, new_new_n5252__, new_new_n5253__,
    new_new_n5254__, new_new_n5255__, new_new_n5256__, new_new_n5257__,
    new_new_n5258__, new_new_n5259__, new_new_n5260__, new_new_n5261__,
    new_new_n5262__, new_new_n5263__, new_new_n5264__, new_new_n5265__,
    new_new_n5266__, new_new_n5267__, new_new_n5268__, new_new_n5269__,
    new_new_n5270__, new_new_n5271__, new_new_n5272__, new_new_n5273__,
    new_new_n5274__, new_new_n5275__, new_new_n5276__, new_new_n5277__,
    new_new_n5278__, new_new_n5279__, new_new_n5280__, new_new_n5281__,
    new_new_n5282__, new_new_n5283__, new_new_n5284__, new_new_n5285__,
    new_new_n5286__, new_new_n5287__, new_new_n5288__, new_new_n5289__,
    new_new_n5290__, new_new_n5291__, new_new_n5292__, new_new_n5293__,
    new_new_n5294__, new_new_n5295__, new_new_n5296__, new_new_n5297__,
    new_new_n5298__, new_new_n5299__, new_new_n5300__, new_new_n5301__,
    new_new_n5302__, new_new_n5303__, new_new_n5304__, new_new_n5305__,
    new_new_n5306__, new_new_n5307__, new_new_n5308__, new_new_n5309__,
    new_new_n5310__, new_new_n5311__, new_new_n5312__, new_new_n5313__,
    new_new_n5314__, new_new_n5315__, new_new_n5316__, new_new_n5317__,
    new_new_n5318__, new_new_n5319__, new_new_n5320__, new_new_n5321__,
    new_new_n5322__, new_new_n5323__, new_new_n5324__, new_new_n5325__,
    new_new_n5326__, new_new_n5327__, new_new_n5328__, new_new_n5329__,
    new_new_n5330__, new_new_n5331__, new_new_n5332__, new_new_n5333__,
    new_new_n5334__, new_new_n5335__, new_new_n5336__, new_new_n5337__,
    new_new_n5338__, new_new_n5339__, new_new_n5340__, new_new_n5341__,
    new_new_n5342__, new_new_n5343__, new_new_n5344__, new_new_n5345__,
    new_new_n5346__, new_new_n5347__, new_new_n5348__, new_new_n5349__,
    new_new_n5350__, new_new_n5351__, new_new_n5352__, new_new_n5353__,
    new_new_n5354__, new_new_n5355__, new_new_n5356__, new_new_n5357__,
    new_new_n5358__, new_new_n5359__, new_new_n5360__, new_new_n5361__,
    new_new_n5362__, new_new_n5363__, new_new_n5364__, new_new_n5365__,
    new_new_n5366__, new_new_n5367__, new_new_n5368__, new_new_n5369__,
    new_new_n5370__, new_new_n5371__, new_new_n5372__, new_new_n5373__,
    new_new_n5374__, new_new_n5375__, new_new_n5376__, new_new_n5377__,
    new_new_n5378__, new_new_n5379__, new_new_n5380__, new_new_n5381__,
    new_new_n5382__, new_new_n5383__, new_new_n5384__, new_new_n5385__,
    new_new_n5386__, new_new_n5387__, new_new_n5388__, new_new_n5389__,
    new_new_n5390__, new_new_n5391__, new_new_n5392__, new_new_n5393__,
    new_new_n5394__, new_new_n5395__, new_new_n5396__, new_new_n5397__,
    new_new_n5398__, new_new_n5399__, new_new_n5400__, new_new_n5401__,
    new_new_n5402__, new_new_n5403__, new_new_n5404__, new_new_n5405__,
    new_new_n5406__, new_new_n5407__, new_new_n5408__, new_new_n5409__,
    new_new_n5410__, new_new_n5411__, new_new_n5412__, new_new_n5413__,
    new_new_n5414__, new_new_n5415__, new_new_n5416__, new_new_n5417__,
    new_new_n5418__, new_new_n5419__, new_new_n5420__, new_new_n5421__,
    new_new_n5422__, new_new_n5423__, new_new_n5424__, new_new_n5425__,
    new_new_n5426__, new_new_n5427__, new_new_n5428__, new_new_n5429__,
    new_new_n5430__, new_new_n5431__, new_new_n5432__, new_new_n5433__,
    new_new_n5434__, new_new_n5435__, new_new_n5436__, new_new_n5437__,
    new_new_n5438__, new_new_n5439__, new_new_n5440__, new_new_n5441__,
    new_new_n5442__, new_new_n5443__, new_new_n5444__, new_new_n5445__,
    new_new_n5446__, new_new_n5447__, new_new_n5448__, new_new_n5449__,
    new_new_n5450__, new_new_n5451__, new_new_n5452__, new_new_n5453__,
    new_new_n5454__, new_new_n5455__, new_new_n5456__, new_new_n5457__,
    new_new_n5458__, new_new_n5459__, new_new_n5460__, new_new_n5461__,
    new_new_n5462__, new_new_n5463__, new_new_n5464__, new_new_n5465__,
    new_new_n5466__, new_new_n5467__, new_new_n5468__, new_new_n5469__,
    new_new_n5470__, new_new_n5471__, new_new_n5472__, new_new_n5473__,
    new_new_n5474__, new_new_n5475__, new_new_n5476__, new_new_n5477__,
    new_new_n5478__, new_new_n5479__, new_new_n5480__, new_new_n5481__,
    new_new_n5482__, new_new_n5483__, new_new_n5484__, new_new_n5485__,
    new_new_n5486__, new_new_n5487__, new_new_n5488__, new_new_n5489__,
    new_new_n5490__, new_new_n5491__, new_new_n5492__, new_new_n5493__,
    new_new_n5494__, new_new_n5495__, new_new_n5496__, new_new_n5497__,
    new_new_n5498__, new_new_n5499__, new_new_n5500__, new_new_n5501__,
    new_new_n5502__, new_new_n5503__, new_new_n5504__, new_new_n5505__,
    new_new_n5506__, new_new_n5507__, new_new_n5508__, new_new_n5509__,
    new_new_n5510__, new_new_n5511__, new_new_n5512__, new_new_n5513__,
    new_new_n5514__, new_new_n5515__, new_new_n5516__, new_new_n5517__,
    new_new_n5518__, new_new_n5519__, new_new_n5520__, new_new_n5521__,
    new_new_n5522__, new_new_n5523__, new_new_n5524__, new_new_n5525__,
    new_new_n5526__, new_new_n5527__, new_new_n5528__, new_new_n5529__,
    new_new_n5530__, new_new_n5531__, new_new_n5532__, new_new_n5533__,
    new_new_n5534__, new_new_n5535__, new_new_n5536__, new_new_n5537__,
    new_new_n5538__, new_new_n5539__, new_new_n5540__, new_new_n5541__,
    new_new_n5542__, new_new_n5543__, new_new_n5544__, new_new_n5545__,
    new_new_n5546__, new_new_n5547__, new_new_n5548__, new_new_n5549__,
    new_new_n5550__, new_new_n5551__, new_new_n5552__, new_new_n5553__,
    new_new_n5554__, new_new_n5555__, new_new_n5556__, new_new_n5557__,
    new_new_n5558__, new_new_n5559__, new_new_n5560__, new_new_n5561__,
    new_new_n5562__, new_new_n5563__, new_new_n5564__, new_new_n5565__,
    new_new_n5566__, new_new_n5567__, new_new_n5568__, new_new_n5569__,
    new_new_n5570__, new_new_n5571__, new_new_n5572__, new_new_n5573__,
    new_new_n5574__, new_new_n5575__, new_new_n5576__, new_new_n5577__,
    new_new_n5578__, new_new_n5579__, new_new_n5580__, new_new_n5581__,
    new_new_n5582__, new_new_n5583__, new_new_n5584__, new_new_n5585__,
    new_new_n5586__, new_new_n5587__, new_new_n5588__, new_new_n5589__,
    new_new_n5590__, new_new_n5591__, new_new_n5592__, new_new_n5593__,
    new_new_n5594__, new_new_n5595__, new_new_n5596__, new_new_n5597__,
    new_new_n5598__, new_new_n5599__, new_new_n5600__, new_new_n5601__,
    new_new_n5602__, new_new_n5603__, new_new_n5604__, new_new_n5605__,
    new_new_n5606__, new_new_n5607__, new_new_n5608__, new_new_n5609__,
    new_new_n5610__, new_new_n5611__, new_new_n5612__, new_new_n5613__,
    new_new_n5614__, new_new_n5615__, new_new_n5616__, new_new_n5617__,
    new_new_n5618__, new_new_n5619__, new_new_n5620__, new_new_n5621__,
    new_new_n5622__, new_new_n5623__, new_new_n5624__, new_new_n5625__,
    new_new_n5626__, new_new_n5627__, new_new_n5628__, new_new_n5629__,
    new_new_n5630__, new_new_n5631__, new_new_n5632__, new_new_n5633__,
    new_new_n5634__, new_new_n5635__, new_new_n5636__, new_new_n5637__,
    new_new_n5638__, new_new_n5639__, new_new_n5640__, new_new_n5641__,
    new_new_n5642__, new_new_n5643__, new_new_n5644__, new_new_n5645__,
    new_new_n5646__, new_new_n5647__, new_new_n5648__, new_new_n5649__,
    new_new_n5650__, new_new_n5651__, new_new_n5652__, new_new_n5653__,
    new_new_n5654__, new_new_n5655__, new_new_n5656__, new_new_n5657__,
    new_new_n5658__, new_new_n5659__, new_new_n5660__, new_new_n5661__,
    new_new_n5662__, new_new_n5663__, new_new_n5664__, new_new_n5665__,
    new_new_n5666__, new_new_n5667__, new_new_n5668__, new_new_n5669__,
    new_new_n5670__, new_new_n5671__, new_new_n5672__, new_new_n5673__,
    new_new_n5674__, new_new_n5675__, new_new_n5676__, new_new_n5677__,
    new_new_n5678__, new_new_n5679__, new_new_n5680__, new_new_n5681__,
    new_new_n5682__, new_new_n5683__, new_new_n5684__, new_new_n5685__,
    new_new_n5686__, new_new_n5687__, new_new_n5688__, new_new_n5689__,
    new_new_n5690__, new_new_n5691__, new_new_n5692__, new_new_n5693__,
    new_new_n5694__, new_new_n5695__, new_new_n5696__, new_new_n5697__,
    new_new_n5698__, new_new_n5699__, new_new_n5700__, new_new_n5701__,
    new_new_n5702__, new_new_n5703__, new_new_n5704__, new_new_n5705__,
    new_new_n5706__, new_new_n5707__, new_new_n5708__, new_new_n5709__,
    new_new_n5710__, new_new_n5711__, new_new_n5712__, new_new_n5713__,
    new_new_n5714__, new_new_n5715__, new_new_n5716__, new_new_n5717__,
    new_new_n5718__, new_new_n5719__, new_new_n5720__, new_new_n5721__,
    new_new_n5722__, new_new_n5723__, new_new_n5724__, new_new_n5725__,
    new_new_n5726__, new_new_n5727__, new_new_n5728__, new_new_n5729__,
    new_new_n5730__, new_new_n5731__, new_new_n5732__, new_new_n5733__,
    new_new_n5734__, new_new_n5735__, new_new_n5736__, new_new_n5737__,
    new_new_n5738__, new_new_n5739__, new_new_n5740__, new_new_n5741__,
    new_new_n5742__, new_new_n5743__, new_new_n5744__, new_new_n5745__,
    new_new_n5746__, new_new_n5747__, new_new_n5748__, new_new_n5749__,
    new_new_n5750__, new_new_n5751__, new_new_n5752__, new_new_n5753__,
    new_new_n5754__, new_new_n5755__, new_new_n5756__, new_new_n5757__,
    new_new_n5758__, new_new_n5759__, new_new_n5760__, new_new_n5761__,
    new_new_n5762__, new_new_n5763__, new_new_n5764__, new_new_n5765__,
    new_new_n5766__, new_new_n5767__, new_new_n5768__, new_new_n5769__,
    new_new_n5770__, new_new_n5771__, new_new_n5772__, new_new_n5773__,
    new_new_n5774__, new_new_n5775__, new_new_n5776__, new_new_n5777__,
    new_new_n5778__, new_new_n5779__, new_new_n5780__, new_new_n5781__,
    new_new_n5782__, new_new_n5783__, new_new_n5784__, new_new_n5785__,
    new_new_n5786__, new_new_n5787__, new_new_n5788__, new_new_n5789__,
    new_new_n5790__, new_new_n5791__, new_new_n5792__, new_new_n5793__,
    new_new_n5794__, new_new_n5795__, new_new_n5796__, new_new_n5797__,
    new_new_n5798__, new_new_n5799__, new_new_n5800__, new_new_n5801__,
    new_new_n5802__, new_new_n5803__, new_new_n5804__, new_new_n5805__,
    new_new_n5806__, new_new_n5807__, new_new_n5808__, new_new_n5809__,
    new_new_n5810__, new_new_n5811__, new_new_n5812__, new_new_n5813__,
    new_new_n5814__, new_new_n5815__, new_new_n5816__, new_new_n5817__,
    new_new_n5818__, new_new_n5819__, new_new_n5820__, new_new_n5821__,
    new_new_n5822__, new_new_n5823__, new_new_n5824__, new_new_n5825__,
    new_new_n5826__, new_new_n5827__, new_new_n5828__, new_new_n5829__,
    new_new_n5830__, new_new_n5831__, new_new_n5832__, new_new_n5833__,
    new_new_n5834__, new_new_n5835__, new_new_n5836__, new_new_n5837__,
    new_new_n5838__, new_new_n5839__, new_new_n5840__, new_new_n5841__,
    new_new_n5842__, new_new_n5843__, new_new_n5844__, new_new_n5845__,
    new_new_n5846__, new_new_n5847__, new_new_n5848__, new_new_n5849__,
    new_new_n5850__, new_new_n5851__, new_new_n5852__, new_new_n5853__,
    new_new_n5854__, new_new_n5855__, new_new_n5856__, new_new_n5857__,
    new_new_n5858__, new_new_n5859__, new_new_n5860__, new_new_n5861__,
    new_new_n5862__, new_new_n5863__, new_new_n5864__, new_new_n5865__,
    new_new_n5866__, new_new_n5867__, new_new_n5868__, new_new_n5869__,
    new_new_n5870__, new_new_n5871__, new_new_n5872__, new_new_n5873__,
    new_new_n5874__, new_new_n5875__, new_new_n5876__, new_new_n5877__,
    new_new_n5878__, new_new_n5879__, new_new_n5880__, new_new_n5881__,
    new_new_n5882__, new_new_n5883__, new_new_n5884__, new_new_n5885__,
    new_new_n5886__, new_new_n5887__, new_new_n5888__, new_new_n5889__,
    new_new_n5890__, new_new_n5891__, new_new_n5892__, new_new_n5893__,
    new_new_n5894__, new_new_n5895__, new_new_n5896__, new_new_n5897__,
    new_new_n5898__, new_new_n5899__, new_new_n5900__, new_new_n5901__,
    new_new_n5902__, new_new_n5903__, new_new_n5904__, new_new_n5905__,
    new_new_n5906__, new_new_n5907__, new_new_n5908__, new_new_n5909__,
    new_new_n5910__, new_new_n5911__, new_new_n5912__, new_new_n5913__,
    new_new_n5914__, new_new_n5915__, new_new_n5916__, new_new_n5917__,
    new_new_n5918__, new_new_n5919__, new_new_n5920__, new_new_n5921__,
    new_new_n5922__, new_new_n5923__, new_new_n5924__, new_new_n5925__,
    new_new_n5926__, new_new_n5927__, new_new_n5928__, new_new_n5929__,
    new_new_n5930__, new_new_n5931__, new_new_n5932__, new_new_n5933__,
    new_new_n5934__, new_new_n5935__, new_new_n5936__, new_new_n5937__,
    new_new_n5938__, new_new_n5939__, new_new_n5940__, new_new_n5941__,
    new_new_n5942__, new_new_n5943__, new_new_n5944__, new_new_n5945__,
    new_new_n5946__, new_new_n5947__, new_new_n6352__, new_new_n6353__,
    new_new_n6354__, new_new_n6355__, new_new_n6356__, new_new_n6357__,
    new_new_n6358__, new_new_n6359__, new_new_n6360__, new_new_n6361__,
    new_new_n6362__, new_new_n6363__, new_new_n6364__, new_new_n6365__,
    new_new_n6366__, new_new_n6367__, new_new_n6368__, new_new_n6369__,
    new_new_n6370__, new_new_n6371__, new_new_n6372__, new_new_n6373__,
    new_new_n6374__, new_new_n6375__, new_new_n6376__, new_new_n6377__,
    new_new_n6378__, new_new_n6379__, new_new_n6380__, new_new_n6381__,
    new_new_n6382__, new_new_n6383__, new_new_n6384__, new_new_n6385__,
    new_new_n6386__, new_new_n6387__, new_new_n6388__, new_new_n6389__,
    new_new_n6390__, new_new_n6391__, new_new_n6392__, new_new_n6393__,
    new_new_n6394__, new_new_n6395__, new_new_n6396__, new_new_n6397__,
    new_new_n6398__, new_new_n6399__, new_new_n6400__, new_new_n6401__,
    new_new_n6402__, new_new_n6403__, new_new_n6404__, new_new_n6405__,
    new_new_n6406__, new_new_n6407__, new_new_n6408__, new_new_n6409__,
    new_new_n6410__, new_new_n6411__, new_new_n6412__, new_new_n6413__,
    new_new_n6414__, new_new_n6415__, new_new_n6416__, new_new_n6417__,
    new_new_n6418__, new_new_n6419__, new_new_n6420__, new_new_n6421__,
    new_new_n6422__, new_new_n6423__, new_new_n6424__, new_new_n6425__,
    new_new_n6426__, new_new_n6427__, new_new_n6428__, new_new_n6429__,
    new_new_n6430__, new_new_n6431__, new_new_n6432__, new_new_n6433__,
    new_new_n6434__, new_new_n6435__, new_new_n6436__, new_new_n6437__,
    new_new_n6438__, new_new_n6439__, new_new_n6440__, new_new_n6441__,
    new_new_n6442__, new_new_n6443__, new_new_n6444__, new_new_n6445__,
    new_new_n6446__, new_new_n6447__, new_new_n6448__, new_new_n6449__,
    new_new_n6450__, new_new_n6451__, new_new_n6452__, new_new_n6453__,
    new_new_n6454__, new_new_n6455__, new_new_n6456__, new_new_n6457__,
    new_new_n6458__, new_new_n6459__, new_new_n6460__, new_new_n6461__,
    new_new_n6462__, new_new_n6463__, new_new_n6464__, new_new_n6465__,
    new_new_n6466__, new_new_n6467__, new_new_n6468__, new_new_n6469__,
    new_new_n6470__, new_new_n6471__, new_new_n6472__, new_new_n6473__,
    new_new_n6474__, new_new_n6475__, new_new_n6476__, new_new_n6477__,
    new_new_n6478__, new_new_n6479__, new_new_n6480__, new_new_n6481__,
    new_new_n6482__, new_new_n6483__, new_new_n6484__, new_new_n6485__,
    new_new_n6486__, new_new_n6487__, new_new_n6488__, new_new_n6489__,
    new_new_n6490__, new_new_n6491__, new_new_n6492__, new_new_n6493__,
    new_new_n6494__, new_new_n6495__, new_new_n6496__, new_new_n6497__,
    new_new_n6498__, new_new_n6499__, new_new_n6500__, new_new_n6501__,
    new_new_n6502__, new_new_n6503__, new_new_n6504__, new_new_n6505__,
    new_new_n6506__, new_new_n6507__, new_new_n6508__, new_new_n6509__,
    new_new_n6510__, new_new_n6511__, new_new_n6512__, new_new_n6513__,
    new_new_n6514__, new_new_n6515__, new_new_n6516__, new_new_n6517__,
    new_new_n6518__, new_new_n6519__, new_new_n6520__, new_new_n6521__,
    new_new_n6522__, new_new_n6523__, new_new_n6524__, new_new_n6525__,
    new_new_n6526__, new_new_n6527__, new_new_n6528__, new_new_n6529__,
    new_new_n6530__, new_new_n6531__, new_new_n6532__, new_new_n6533__,
    new_new_n6534__, new_new_n6535__, new_new_n6536__, new_new_n6537__,
    new_new_n6538__, new_new_n6539__, new_new_n6540__, new_new_n6541__,
    new_new_n6542__, new_new_n6543__, new_new_n6544__, new_new_n6545__,
    new_new_n6546__, new_new_n6547__, new_new_n6548__, new_new_n6549__,
    new_new_n6550__, new_new_n6551__, new_new_n6552__, new_new_n6553__,
    new_new_n6554__, new_new_n6555__, new_new_n6556__, new_new_n6557__,
    new_new_n6558__, new_new_n6559__, new_new_n6560__, new_new_n6561__,
    new_new_n6562__, new_new_n6563__, new_new_n6564__, new_new_n6565__,
    new_new_n6566__, new_new_n6567__, new_new_n6568__, new_new_n6569__,
    new_new_n6570__, new_new_n6571__, new_new_n6572__, new_new_n6573__,
    new_new_n6574__, new_new_n6575__, new_new_n6576__, new_new_n6577__,
    new_new_n6578__, new_new_n6579__, new_new_n6580__, new_new_n6581__,
    new_new_n6582__, new_new_n6583__, new_new_n6584__, new_new_n6585__,
    new_new_n6586__, new_new_n6587__, new_new_n6588__, new_new_n6589__,
    new_new_n6590__, new_new_n6591__, new_new_n6592__, new_new_n6593__,
    new_new_n6594__, new_new_n6595__, new_new_n6596__, new_new_n6597__,
    new_new_n6598__, new_new_n6599__, new_new_n6600__, new_new_n6601__,
    new_new_n6602__, new_new_n6603__, new_new_n6604__, new_new_n6605__,
    new_new_n6606__, new_new_n6607__, new_new_n6608__, new_new_n6609__,
    new_new_n6610__, new_new_n6611__, new_new_n6612__, new_new_n6613__,
    new_new_n6614__, new_new_n6615__, new_new_n6616__, new_new_n6617__,
    new_new_n6618__, new_new_n6619__, new_new_n6620__, new_new_n6621__,
    new_new_n6622__, new_new_n6623__, new_new_n6624__, new_new_n6625__,
    new_new_n6626__, new_new_n6627__, new_new_n6628__, new_new_n6629__,
    new_new_n6630__, new_new_n6631__, new_new_n6632__, new_new_n6633__,
    new_new_n6634__, new_new_n6635__, new_new_n6636__, new_new_n6637__,
    new_new_n6638__, new_new_n6639__, new_new_n6640__, new_new_n6641__,
    new_new_n6642__, new_new_n6643__, new_new_n6644__, new_new_n6645__,
    new_new_n6646__, new_new_n6647__, new_new_n6648__, new_new_n6649__,
    new_new_n6650__, new_new_n6651__, new_new_n6652__, new_new_n6653__,
    new_new_n6654__, new_new_n6655__, new_new_n6656__, new_new_n6657__,
    new_new_n6658__, new_new_n6659__, new_new_n6660__, new_new_n6661__,
    new_new_n6662__, new_new_n6663__, new_new_n6664__, new_new_n6665__,
    new_new_n6666__, new_new_n6667__, new_new_n6668__, new_new_n6669__,
    new_new_n6670__, new_new_n6671__, new_new_n6672__, new_new_n6673__,
    new_new_n6674__, new_new_n6675__, new_new_n6676__, new_new_n6677__,
    new_new_n6678__, new_new_n6679__, new_new_n6680__, new_new_n6681__,
    new_new_n6682__, new_new_n6683__, new_new_n6684__, new_new_n6685__,
    new_new_n6686__, new_new_n6687__, new_new_n6688__, new_new_n6689__,
    new_new_n6690__, new_new_n6691__, new_new_n6692__, new_new_n6693__,
    new_new_n6694__, new_new_n6695__, new_new_n6696__, new_new_n6697__,
    new_new_n6698__, new_new_n6699__, new_new_n6700__, new_new_n6701__,
    new_new_n6702__, new_new_n6703__, new_new_n6704__, new_new_n6705__,
    new_new_n6706__, new_new_n6707__, new_new_n6708__, new_new_n6709__,
    new_new_n6710__, new_new_n6711__, new_new_n6712__, new_new_n6713__,
    new_new_n6714__, new_new_n6715__, new_new_n6716__, new_new_n6717__,
    new_new_n6718__, new_new_n6719__, new_new_n6720__, new_new_n6721__,
    new_new_n6722__, new_new_n6723__, new_new_n6724__, new_new_n6725__,
    new_new_n6726__, new_new_n6727__, new_new_n6728__, new_new_n6729__,
    new_new_n6730__, new_new_n6731__, new_new_n6732__, new_new_n6733__,
    new_new_n6734__, new_new_n6735__, new_new_n6736__, new_new_n6737__,
    new_new_n6738__, new_new_n6739__, new_new_n6740__, new_new_n6741__,
    new_new_n6742__, new_new_n6743__, new_new_n6744__, new_new_n6745__,
    new_new_n6746__, new_new_n6747__, new_new_n6748__, new_new_n6749__,
    new_new_n6750__, new_new_n6751__, new_new_n6752__, new_new_n6753__,
    new_new_n6754__, new_new_n6755__, new_new_n6756__, new_new_n6757__,
    new_new_n6758__, new_new_n6759__, new_new_n6760__, new_new_n6761__,
    new_new_n6762__, new_new_n6763__, new_new_n6764__, new_new_n6765__,
    new_new_n6766__, new_new_n6767__, new_new_n6768__, new_new_n6769__,
    new_new_n6770__, new_new_n6771__, new_new_n6772__, new_new_n6773__,
    new_new_n6774__, new_new_n6775__, new_new_n6776__, new_new_n6777__,
    new_new_n6778__, new_new_n6779__, new_new_n6780__, new_new_n6781__,
    new_new_n6782__, new_new_n6783__, new_new_n6784__, new_new_n6785__,
    new_new_n6786__, new_new_n6787__, new_new_n6788__, new_new_n6789__,
    new_new_n6790__, new_new_n6791__, new_new_n6792__, new_new_n6793__,
    new_new_n6794__, new_new_n6795__, new_new_n6796__, new_new_n6797__,
    new_new_n6798__, new_new_n6799__, new_new_n6800__, new_new_n6801__,
    new_new_n6802__, new_new_n6803__, new_new_n6804__, new_new_n6805__,
    new_new_n6806__, new_new_n6807__, new_new_n6808__, new_new_n6809__,
    new_new_n6810__, new_new_n6811__, new_new_n6812__, new_new_n6813__,
    new_new_n6814__, new_new_n6815__, new_new_n6816__, new_new_n6817__,
    new_new_n6818__, new_new_n6819__, new_new_n6820__, new_new_n6821__,
    new_new_n6822__, new_new_n6823__, new_new_n6824__, new_new_n6825__,
    new_new_n6826__, new_new_n6827__, new_new_n6828__, new_new_n6829__,
    new_new_n6830__, new_new_n6831__, new_new_n6832__, new_new_n6833__,
    new_new_n6834__, new_new_n6835__, new_new_n6836__, new_new_n6837__,
    new_new_n6838__, new_new_n6839__, new_new_n6840__, new_new_n6841__,
    new_new_n6842__, new_new_n6843__, new_new_n6844__, new_new_n6845__,
    new_new_n6846__, new_new_n6847__, new_new_n6848__, new_new_n6849__,
    new_new_n6850__, new_new_n6851__, new_new_n6852__, new_new_n6853__,
    new_new_n6854__, new_new_n6855__, new_new_n6856__, new_new_n6857__,
    new_new_n6858__, new_new_n6859__, new_new_n6860__, new_new_n6861__,
    new_new_n6862__, new_new_n6863__, new_new_n6864__, new_new_n6865__,
    new_new_n6866__, new_new_n6867__, new_new_n6868__, new_new_n6869__,
    new_new_n6870__, new_new_n6871__, new_new_n6872__, new_new_n6873__,
    new_new_n6874__, new_new_n6875__, new_new_n6876__, new_new_n6877__,
    new_new_n6878__, new_new_n6879__, new_new_n6880__, new_new_n6881__,
    new_new_n6882__, new_new_n6883__, new_new_n6884__, new_new_n6885__,
    new_new_n6886__, new_new_n6887__, new_new_n6888__, new_new_n6889__,
    new_new_n6890__, new_new_n6891__, new_new_n6892__, new_new_n6893__,
    new_new_n6894__, new_new_n6895__, new_new_n6896__, new_new_n6897__,
    new_new_n6898__, new_new_n6899__, new_new_n6900__, new_new_n6901__,
    new_new_n6902__, new_new_n6903__, new_new_n6904__, new_new_n6905__,
    new_new_n6906__, new_new_n6907__, new_new_n6908__, new_new_n6909__,
    new_new_n6910__, new_new_n6911__, new_new_n6912__, new_new_n6913__,
    new_new_n6914__, new_new_n6915__, new_new_n6916__, new_new_n6917__,
    new_new_n6918__, new_new_n6919__, new_new_n6920__, new_new_n6921__,
    new_new_n6922__, new_new_n6923__, new_new_n6924__, new_new_n6925__,
    new_new_n6926__, new_new_n6927__, new_new_n6928__, new_new_n6929__,
    new_new_n6930__, new_new_n6931__, new_new_n6932__, new_new_n6933__,
    new_new_n6934__, new_new_n6935__, new_new_n6936__, new_new_n6937__,
    new_new_n6938__, new_new_n6939__, new_new_n6940__, new_new_n6941__,
    new_new_n6942__, new_new_n6943__, new_new_n6944__, new_new_n6945__,
    new_new_n6946__, new_new_n6947__, new_new_n6948__, new_new_n6949__,
    new_new_n6950__, new_new_n6951__, new_new_n6952__, new_new_n6953__,
    new_new_n6954__, new_new_n6955__, new_new_n6956__, new_new_n6957__,
    new_new_n6958__, new_new_n6959__, new_new_n6960__, new_new_n6961__,
    new_new_n6962__, new_new_n6963__, new_new_n6964__, new_new_n6965__,
    new_new_n6966__, new_new_n6967__, new_new_n6968__, new_new_n6969__,
    new_new_n6970__, new_new_n6971__, new_new_n6972__, new_new_n6973__,
    new_new_n6974__, new_new_n6975__, new_new_n6976__, new_new_n6977__,
    new_new_n6978__, new_new_n6979__, new_new_n6980__, new_new_n6981__,
    new_new_n6982__, new_new_n6983__, new_new_n6984__, new_new_n6985__,
    new_new_n6986__, new_new_n6987__, new_new_n6988__, new_new_n6989__,
    new_new_n6990__, new_new_n6991__, new_new_n6992__, new_new_n6993__,
    new_new_n6994__, new_new_n6995__, new_new_n6996__, new_new_n6997__,
    new_new_n6998__, new_new_n6999__, new_new_n7000__, new_new_n7001__,
    new_new_n7002__, new_new_n7003__, new_new_n7004__, new_new_n7005__,
    new_new_n7006__, new_new_n7007__, new_new_n7008__, new_new_n7009__,
    new_new_n7010__, new_new_n7011__, new_new_n7012__, new_new_n7013__,
    new_new_n7014__, new_new_n7015__, new_new_n7016__, new_new_n7017__,
    new_new_n7018__, new_new_n7019__, new_new_n7020__, new_new_n7021__,
    new_new_n7022__, new_new_n7023__, new_new_n7024__, new_new_n7025__,
    new_new_n7026__, new_new_n7027__, new_new_n7028__, new_new_n7029__,
    new_new_n7030__, new_new_n7031__, new_new_n7032__, new_new_n7033__,
    new_new_n7034__, new_new_n7035__, new_new_n7036__, new_new_n7037__,
    new_new_n7038__, new_new_n7039__, new_new_n7040__, new_new_n7041__,
    new_new_n7042__, new_new_n7043__, new_new_n7044__, new_new_n7045__,
    new_new_n7046__, new_new_n7047__, new_new_n7048__, new_new_n7049__,
    new_new_n7050__, new_new_n7051__, new_new_n7052__, new_new_n7053__,
    new_new_n7054__, new_new_n7055__, new_new_n7056__, new_new_n7057__,
    new_new_n7058__, new_new_n7059__, new_new_n7060__, new_new_n7061__,
    new_new_n7062__, new_new_n7063__, new_new_n7064__, new_new_n7065__,
    new_new_n7066__, new_new_n7067__, new_new_n7068__, new_new_n7069__,
    new_new_n7070__, new_new_n7071__, new_new_n7072__, new_new_n7073__,
    new_new_n7074__, new_new_n7075__, new_new_n7076__, new_new_n7077__,
    new_new_n7078__, new_new_n7079__, new_new_n7080__, new_new_n7081__,
    new_new_n7082__, new_new_n7083__, new_new_n7084__, new_new_n7085__,
    new_new_n7086__, new_new_n7087__, new_new_n7088__, new_new_n7089__,
    new_new_n7090__, new_new_n7091__, new_new_n7092__, new_new_n7093__,
    new_new_n7094__, new_new_n7095__, new_new_n7096__, new_new_n7097__,
    new_new_n7098__, new_new_n7099__, new_new_n7100__, new_new_n7101__,
    new_new_n7102__, new_new_n7103__, new_new_n7104__, new_new_n7105__,
    new_new_n7106__, new_new_n7107__, new_new_n7108__, new_new_n7109__,
    new_new_n7110__, new_new_n7111__, new_new_n7112__, new_new_n7113__,
    new_new_n7114__, new_new_n7115__, new_new_n7116__, new_new_n7117__,
    new_new_n7118__, new_new_n7119__, new_new_n7120__, new_new_n7121__,
    new_new_n7122__, new_new_n7123__, new_new_n7124__, new_new_n7125__,
    new_new_n7126__, new_new_n7127__, new_new_n7128__, new_new_n7129__,
    new_new_n7130__, new_new_n7131__, new_new_n7132__, new_new_n7133__,
    new_new_n7134__, new_new_n7135__, new_new_n7136__, new_new_n7137__,
    new_new_n7138__, new_new_n7139__, new_new_n7140__, new_new_n7141__,
    new_new_n7142__, new_new_n7143__, new_new_n7144__, new_new_n7145__,
    new_new_n7146__, new_new_n7147__, new_new_n7148__, new_new_n7149__,
    new_new_n7150__, new_new_n7151__, new_new_n7152__, new_new_n7153__,
    new_new_n7154__, new_new_n7155__, new_new_n7156__, new_new_n7157__,
    new_new_n7158__, new_new_n7159__, new_new_n7160__, new_new_n7161__,
    new_new_n7162__, new_new_n7163__, new_new_n7164__, new_new_n7165__,
    new_new_n7166__, new_new_n7167__, new_new_n7168__, new_new_n7169__,
    new_new_n7170__, new_new_n7171__, new_new_n7172__, new_new_n7173__,
    new_new_n7174__, new_new_n7175__, new_new_n7176__, new_new_n7177__,
    new_new_n7178__, new_new_n7179__, new_new_n7180__, new_new_n7181__,
    new_new_n7182__, new_new_n7183__, new_new_n7184__, new_new_n7185__,
    new_new_n7186__, new_new_n7187__, new_new_n7188__, new_new_n7189__,
    new_new_n7190__, new_new_n7191__, new_new_n7192__, new_new_n7193__,
    new_new_n7194__, new_new_n7195__, new_new_n7196__, new_new_n7197__,
    new_new_n7198__, new_new_n7199__, new_new_n7200__, new_new_n7201__,
    new_new_n7202__, new_new_n7203__, new_new_n7204__, new_new_n7205__,
    new_new_n7206__, new_new_n7207__, new_new_n7208__, new_new_n7209__,
    new_new_n7210__, new_new_n7211__, new_new_n7212__, new_new_n7213__,
    new_new_n7214__, new_new_n7215__, new_new_n7216__, new_new_n7217__,
    new_new_n7218__, new_new_n7219__, new_new_n7220__, new_new_n7221__,
    new_new_n7222__, new_new_n7223__, new_new_n7224__, new_new_n7225__,
    new_new_n7226__, new_new_n7227__, new_new_n7228__, new_new_n7229__,
    new_new_n7230__, new_new_n7231__, new_new_n7232__, new_new_n7233__,
    new_new_n7234__, new_new_n7235__, new_new_n7236__, new_new_n7237__,
    new_new_n7238__, new_new_n7239__, new_new_n7240__, new_new_n7241__,
    new_new_n7242__, new_new_n7243__, new_new_n7244__, new_new_n7245__,
    new_new_n7246__, new_new_n7247__, new_new_n7248__, new_new_n7249__,
    new_new_n7250__, new_new_n7251__, new_new_n7252__, new_new_n7253__,
    new_new_n7254__, new_new_n7255__, new_new_n7256__, new_new_n7257__,
    new_new_n7258__, new_new_n7259__, new_new_n7260__, new_new_n7261__,
    new_new_n7262__, new_new_n7263__, new_new_n7264__, new_new_n7265__,
    new_new_n7266__, new_new_n7267__, new_new_n7268__, new_new_n7269__,
    new_new_n7270__, new_new_n7271__, new_new_n7272__, new_new_n7273__,
    new_new_n7274__, new_new_n7275__, new_new_n7276__, new_new_n7277__,
    new_new_n7278__, new_new_n7279__, new_new_n7280__, new_new_n7281__,
    new_new_n7282__, new_new_n7283__, new_new_n7284__, new_new_n7285__,
    new_new_n7286__, new_new_n7287__, new_new_n7288__, new_new_n7289__,
    new_new_n7290__, new_new_n7291__, new_new_n7292__, new_new_n7293__,
    new_new_n7294__, new_new_n7295__, new_new_n7296__, new_new_n7297__,
    new_new_n7298__, new_new_n7299__, new_new_n7300__, new_new_n7301__,
    new_new_n7302__, new_new_n7303__, new_new_n7304__, new_new_n7305__,
    new_new_n7306__, new_new_n7307__, new_new_n7308__, new_new_n7309__,
    new_new_n7310__, new_new_n7311__, new_new_n7312__, new_new_n7313__,
    new_new_n7314__, new_new_n7315__, new_new_n7316__, new_new_n7317__,
    new_new_n7318__, new_new_n7319__, new_new_n7320__, new_new_n7321__,
    new_new_n7322__, new_new_n7323__, new_new_n7324__, new_new_n7325__,
    new_new_n7326__, new_new_n7327__, new_new_n7328__, new_new_n7329__,
    new_new_n7330__, new_new_n7331__, new_new_n7332__, new_new_n7333__,
    new_new_n7334__, new_new_n7335__, new_new_n7336__, new_new_n7337__,
    new_new_n7338__, new_new_n7339__, new_new_n7340__, new_new_n7341__,
    new_new_n7342__, new_new_n7343__, new_new_n7344__, new_new_n7345__,
    new_new_n7346__, new_new_n7347__, new_new_n7348__, new_new_n7349__,
    new_new_n7350__, new_new_n7351__, new_new_n7352__, new_new_n7353__,
    new_new_n7354__, new_new_n7355__, new_new_n7356__, new_new_n7357__,
    new_new_n7358__, new_new_n7359__, new_new_n7360__, new_new_n7361__,
    new_new_n7362__, new_new_n7363__, new_new_n7364__, new_new_n7365__,
    new_new_n7366__, new_new_n7367__, new_new_n7368__, new_new_n7369__,
    new_new_n7370__, new_new_n7371__, new_new_n7372__, new_new_n7373__,
    new_new_n7374__, new_new_n7375__, new_new_n7376__, new_new_n7377__,
    new_new_n7378__, new_new_n7379__, new_new_n7380__, new_new_n7381__,
    new_new_n7382__, new_new_n7383__, new_new_n7384__, new_new_n7385__,
    new_new_n7386__, new_new_n7387__, new_new_n7388__, new_new_n7389__,
    new_new_n7390__, new_new_n7391__, new_new_n7392__, new_new_n7393__,
    new_new_n7394__, new_new_n7395__, new_new_n7396__, new_new_n7397__,
    new_new_n7398__, new_new_n7399__, new_new_n7400__, new_new_n7401__,
    new_new_n7402__, new_new_n7403__, new_new_n7404__, new_new_n7405__,
    new_new_n7406__, new_new_n7407__, new_new_n7408__, new_new_n7409__,
    new_new_n7410__, new_new_n7411__, new_new_n7412__, new_new_n7413__,
    new_new_n7414__, new_new_n7415__, new_new_n7416__, new_new_n7417__,
    new_new_n7418__, new_new_n7419__, new_new_n7420__, new_new_n7421__,
    new_new_n7422__, new_new_n7423__, new_new_n7424__, new_new_n7425__,
    new_new_n7426__, new_new_n7427__, new_new_n7428__, new_new_n7429__,
    new_new_n7430__, new_new_n7431__, new_new_n7432__, new_new_n7433__,
    new_new_n7434__, new_new_n7435__, new_new_n7436__, new_new_n7437__,
    new_new_n7438__, new_new_n7439__, new_new_n7440__, new_new_n7441__,
    new_new_n7442__, new_new_n7443__, new_new_n7444__, new_new_n7445__,
    new_new_n7446__, new_new_n7447__, new_new_n7448__, new_new_n7449__,
    new_new_n7450__, new_new_n7451__, new_new_n7452__, new_new_n7453__,
    new_new_n7454__, new_new_n7455__, new_new_n7456__, new_new_n7457__,
    new_new_n7458__, new_new_n7459__, new_new_n7460__, new_new_n7461__,
    new_new_n7462__, new_new_n7463__, new_new_n7464__, new_new_n7465__,
    new_new_n7466__, new_new_n7467__, new_new_n7468__, new_new_n7469__,
    new_new_n7470__, new_new_n7471__, new_new_n7472__, new_new_n7473__,
    new_new_n7474__, new_new_n7475__, new_new_n7476__, new_new_n7477__,
    new_new_n7478__, new_new_n7479__, new_new_n7480__, new_new_n7481__,
    new_new_n7482__, new_new_n7483__, new_new_n7484__, new_new_n7485__,
    new_new_n7486__, new_new_n7487__, new_new_n7488__, new_new_n7489__,
    new_new_n7490__, new_new_n7491__, new_new_n7492__, new_new_n7493__,
    new_new_n7494__, new_new_n7495__, new_new_n7496__, new_new_n7497__,
    new_new_n7498__, new_new_n7499__, new_new_n7500__, new_new_n7501__,
    new_new_n7502__, new_new_n7503__, new_new_n7504__, new_new_n7505__,
    new_new_n7506__, new_new_n7507__, new_new_n7508__, new_new_n7509__,
    new_new_n7510__, new_new_n7511__, new_new_n7512__, new_new_n7513__,
    new_new_n7514__, new_new_n7515__, new_new_n7516__, new_new_n7517__,
    new_new_n7518__, new_new_n7519__, new_new_n7520__, new_new_n7521__,
    new_new_n7522__, new_new_n7523__, new_new_n7524__, new_new_n7525__,
    new_new_n7526__, new_new_n7527__, new_new_n7528__, new_new_n7529__,
    new_new_n7530__, new_new_n7531__, new_new_n7532__, new_new_n7533__,
    new_new_n7534__, new_new_n7535__, new_new_n7536__, new_new_n7537__,
    new_new_n7538__, new_new_n7539__, new_new_n7540__, new_new_n7541__,
    new_new_n7542__, new_new_n7543__, new_new_n7544__, new_new_n7545__,
    new_new_n7546__, new_new_n7547__, new_new_n7548__, new_new_n7549__,
    new_new_n7550__, new_new_n7551__, new_new_n7552__, new_new_n7553__,
    new_new_n7554__, new_new_n7555__, new_new_n7556__, new_new_n7557__,
    new_new_n7558__, new_new_n7559__, new_new_n7560__, new_new_n7561__,
    new_new_n7562__, new_new_n7563__, new_new_n7564__, new_new_n7565__,
    new_new_n7566__, new_new_n7567__, new_new_n7568__, new_new_n7569__,
    new_new_n7570__, new_new_n7571__, new_new_n7572__, new_new_n7573__,
    new_new_n7574__, new_new_n7575__, new_new_n7576__, new_new_n7577__,
    new_new_n7578__, new_new_n7579__, new_new_n7580__, new_new_n7581__,
    new_new_n7582__, new_new_n7583__, new_new_n7584__, new_new_n7585__,
    new_new_n7586__, new_new_n7587__, new_new_n7588__, new_new_n7589__,
    new_new_n7590__, new_new_n7591__, new_new_n7592__, new_new_n7593__,
    new_new_n7594__, new_new_n7595__, new_new_n7596__, new_new_n7597__,
    new_new_n7598__, new_new_n7599__, new_new_n7600__, new_new_n7601__,
    new_new_n7602__, new_new_n7603__, new_new_n7604__, new_new_n7605__,
    new_new_n7606__, new_new_n7607__, new_new_n7608__, new_new_n7609__,
    new_new_n7610__, new_new_n7611__, new_new_n7612__, new_new_n7613__,
    new_new_n7614__, new_new_n7615__, new_new_n7616__, new_new_n7617__,
    new_new_n7618__, new_new_n7619__, new_new_n7620__, new_new_n7621__,
    new_new_n7622__, new_new_n7623__, new_new_n7624__, new_new_n7625__,
    new_new_n7626__, new_new_n7627__, new_new_n7628__, new_new_n7629__,
    new_new_n7630__, new_new_n7631__, new_new_n7632__, new_new_n7633__,
    new_new_n7634__, new_new_n7635__, new_new_n7636__, new_new_n7637__,
    new_new_n7638__, new_new_n7639__, new_new_n7640__, new_new_n7641__,
    new_new_n7642__, new_new_n7643__, new_new_n7644__, new_new_n7645__,
    new_new_n7646__, new_new_n7647__, new_new_n7648__, new_new_n7649__,
    new_new_n7650__, new_new_n7651__, new_new_n7652__, new_new_n7653__,
    new_new_n7654__, new_new_n7655__, new_new_n7656__, new_new_n7657__,
    new_new_n7658__, new_new_n7659__, new_new_n7660__, new_new_n7661__,
    new_new_n7662__, new_new_n7663__, new_new_n7664__, new_new_n7665__,
    new_new_n7666__, new_new_n7667__, new_new_n7668__, new_new_n7669__,
    new_new_n7670__, new_new_n7671__, new_new_n7672__, new_new_n7673__,
    new_new_n7674__, new_new_n7675__, new_new_n7676__, new_new_n7677__,
    new_new_n7678__, new_new_n7679__, new_new_n7680__, new_new_n7681__,
    new_new_n7682__, new_new_n7683__, new_new_n7684__, new_new_n7685__,
    new_new_n7686__, new_new_n7687__, new_new_n7688__, new_new_n7689__,
    new_new_n7690__, new_new_n7691__, new_new_n7692__, new_new_n7693__,
    new_new_n7694__, new_new_n7695__, new_new_n7696__, new_new_n7697__,
    new_new_n7698__, new_new_n7699__, new_new_n7700__, new_new_n7701__,
    new_new_n7702__, new_new_n7703__, new_new_n7704__, new_new_n7705__,
    new_new_n7706__, new_new_n7707__, new_new_n7708__, new_new_n7709__,
    new_new_n7710__, new_new_n7711__, new_new_n7712__, new_new_n7713__,
    new_new_n7714__, new_new_n7715__, new_new_n7716__, new_new_n7717__,
    new_new_n7718__, new_new_n7719__, new_new_n7720__, new_new_n7721__,
    new_new_n7722__, new_new_n7723__, new_new_n7724__, new_new_n7725__,
    new_new_n7726__, new_new_n7727__, new_new_n7728__, new_new_n7729__,
    new_new_n7730__, new_new_n7731__, new_new_n7732__, new_new_n7733__,
    new_new_n7734__, new_new_n7735__, new_new_n7736__, new_new_n7737__,
    new_new_n7738__, new_new_n7739__, new_new_n7740__, new_new_n7741__,
    new_new_n7742__, new_new_n7743__, new_new_n7744__, new_new_n7745__,
    new_new_n7746__, new_new_n7747__, new_new_n7748__, new_new_n7749__,
    new_new_n7750__, new_new_n7751__, new_new_n7752__, new_new_n7753__,
    new_new_n7754__, new_new_n7755__, new_new_n7756__, new_new_n7757__,
    new_new_n7758__, new_new_n7759__, new_new_n7760__, new_new_n7761__,
    new_new_n7762__, new_new_n7763__, new_new_n7764__, new_new_n7765__,
    new_new_n7766__, new_new_n7767__, new_new_n7768__, new_new_n7769__,
    new_new_n7770__, new_new_n7771__, new_new_n7772__, new_new_n7773__,
    new_new_n7774__, new_new_n7775__, new_new_n7776__, new_new_n7777__,
    new_new_n7778__, new_new_n7779__, new_new_n7780__, new_new_n7781__,
    new_new_n7782__, new_new_n7783__, new_new_n7784__, new_new_n7785__,
    new_new_n7786__, new_new_n7787__, new_new_n7788__, new_new_n7789__,
    new_new_n7790__, new_new_n7791__, new_new_n7792__, new_new_n7793__,
    new_new_n7794__, new_new_n7795__, new_new_n7796__, new_new_n7797__,
    new_new_n7798__, new_new_n7799__, new_new_n7800__, new_new_n7801__,
    new_new_n7802__, new_new_n7803__, new_new_n7804__, new_new_n7805__,
    new_new_n7806__, new_new_n7807__, new_new_n7808__, new_new_n7809__,
    new_new_n7810__, new_new_n7811__, new_new_n7812__, new_new_n7813__,
    new_new_n7814__, new_new_n7815__, new_new_n7816__, new_new_n7817__,
    new_new_n7818__, new_new_n7819__, new_new_n7820__, new_new_n7821__,
    new_new_n7822__, new_new_n7823__, new_new_n7824__, new_new_n7825__,
    new_new_n7826__, new_new_n7827__, new_new_n7828__, new_new_n7829__,
    new_new_n7830__, new_new_n7831__, new_new_n7832__, new_new_n7833__,
    new_new_n7834__, new_new_n7835__, new_new_n7836__, new_new_n7837__,
    new_new_n7838__, new_new_n7839__, new_new_n7840__, new_new_n7841__,
    new_new_n7842__, new_new_n7843__, new_new_n7844__, new_new_n7845__,
    new_new_n7846__, new_new_n7847__, new_new_n7848__, new_new_n7849__,
    new_new_n7850__, new_new_n7851__, new_new_n7852__, new_new_n7853__,
    new_new_n7854__, new_new_n7855__, new_new_n7856__, new_new_n7857__,
    new_new_n7858__, new_new_n7859__, new_new_n7860__, new_new_n7861__,
    new_new_n7862__, new_new_n7863__, new_new_n7864__, new_new_n7865__,
    new_new_n7866__, new_new_n7867__, new_new_n7868__, new_new_n7869__,
    new_new_n7870__, new_new_n7871__, new_new_n7872__, new_new_n7873__,
    new_new_n7874__, new_new_n7875__, new_new_n7876__, new_new_n7877__,
    new_new_n7878__, new_new_n7879__, new_new_n7880__, new_new_n7881__,
    new_new_n7882__, new_new_n7883__, new_new_n7884__, new_new_n7885__,
    new_new_n7886__, new_new_n7887__, new_new_n7888__, new_new_n7889__,
    new_new_n7890__, new_new_n7891__, new_new_n7892__, new_new_n7893__,
    new_new_n7894__, new_new_n7895__, new_new_n7896__, new_new_n7897__,
    new_new_n7898__, new_new_n7899__, new_new_n7900__, new_new_n7901__,
    new_new_n7902__, new_new_n7903__, new_new_n7904__, new_new_n7905__,
    new_new_n7906__, new_new_n7907__, new_new_n7908__, new_new_n7909__,
    new_new_n7910__, new_new_n7911__, new_new_n7912__, new_new_n7913__,
    new_new_n7914__, new_new_n7915__, new_new_n7916__, new_new_n7917__,
    new_new_n7918__, new_new_n7919__, new_new_n7920__, new_new_n7921__,
    new_new_n7922__, new_new_n7923__, new_new_n7924__, new_new_n7925__,
    new_new_n7926__, new_new_n7927__, new_new_n7928__, new_new_n7929__,
    new_new_n7930__, new_new_n7931__, new_new_n7932__, new_new_n7933__,
    new_new_n7934__, new_new_n7935__, new_new_n7936__, new_new_n7937__,
    new_new_n7938__, new_new_n7939__, new_new_n7940__, new_new_n7941__,
    new_new_n7942__, new_new_n7943__, new_new_n7944__, new_new_n7945__,
    new_new_n7946__, new_new_n7947__, new_new_n7948__, new_new_n7949__,
    new_new_n7950__, new_new_n7951__, new_new_n7952__, new_new_n7953__,
    new_new_n7954__, new_new_n7955__, new_new_n7956__, new_new_n7957__,
    new_new_n7958__, new_new_n7959__, new_new_n7960__, new_new_n7961__,
    new_new_n7962__, new_new_n7963__, new_new_n7964__, new_new_n7965__,
    new_new_n7966__, new_new_n7967__, new_new_n7968__, new_new_n7969__,
    new_new_n7970__, new_new_n7971__, new_new_n7972__, new_new_n7973__,
    new_new_n7974__, new_new_n7975__, new_new_n7976__, new_new_n7977__,
    new_new_n7978__, new_new_n7979__, new_new_n7980__, new_new_n7981__,
    new_new_n7982__, new_new_n7983__, new_new_n7984__, new_new_n7985__,
    new_new_n7986__, new_new_n7987__, new_new_n7988__, new_new_n7989__,
    new_new_n7990__, new_new_n7991__, new_new_n7992__, new_new_n7993__,
    new_new_n7994__, new_new_n7995__, new_new_n7996__, new_new_n7997__,
    new_new_n7998__, new_new_n7999__, new_new_n8000__, new_new_n8001__,
    new_new_n8002__, new_new_n8003__, new_new_n8004__, new_new_n8005__,
    new_new_n8006__, new_new_n8007__, new_new_n8008__, new_new_n8009__,
    new_new_n8010__, new_new_n8011__, new_new_n8012__, new_new_n8013__,
    new_new_n8014__, new_new_n8015__, new_new_n8016__, new_new_n8017__,
    new_new_n8018__, new_new_n8019__, new_new_n8020__, new_new_n8021__,
    new_new_n8022__, new_new_n8023__, new_new_n8024__, new_new_n8025__,
    new_new_n8026__, new_new_n8027__, new_new_n8028__, new_new_n8029__,
    new_new_n8030__, new_new_n8031__, new_new_n8032__, new_new_n8033__,
    new_new_n8034__, new_new_n8035__, new_new_n8036__, new_new_n8037__,
    new_new_n8038__, new_new_n8039__, new_new_n8040__, new_new_n8041__,
    new_new_n8042__, new_new_n8043__, new_new_n8044__, new_new_n8045__,
    new_new_n8046__, new_new_n8047__, new_new_n8048__, new_new_n8049__,
    new_new_n8050__, new_new_n8051__, new_new_n8052__, new_new_n8053__,
    new_new_n8054__, new_new_n8055__, new_new_n8056__, new_new_n8057__,
    new_new_n8058__, new_new_n8059__, new_new_n8060__, new_new_n8061__,
    new_new_n8062__, new_new_n8063__, new_new_n8064__, new_new_n8065__,
    new_new_n8066__, new_new_n8067__, new_new_n8068__, new_new_n8069__,
    new_new_n8070__, new_new_n8071__, new_new_n8072__, new_new_n8073__,
    new_new_n8074__, new_new_n8075__, new_new_n8076__, new_new_n8077__,
    new_new_n8078__, new_new_n8079__, new_new_n8080__, new_new_n8081__,
    new_new_n8082__, new_new_n8083__, new_new_n8084__, new_new_n8085__,
    new_new_n8086__, new_new_n8087__, new_new_n8088__, new_new_n8089__,
    new_new_n8090__, new_new_n8091__, new_new_n8092__, new_new_n8093__,
    new_new_n8094__, new_new_n8095__, new_new_n8096__, new_new_n8097__,
    new_new_n8098__, new_new_n8099__, new_new_n8100__, new_new_n8101__,
    new_new_n8102__, new_new_n8103__, new_new_n8104__, new_new_n8105__,
    new_new_n8106__, new_new_n8107__, new_new_n8108__, new_new_n8109__,
    new_new_n8110__, new_new_n8111__, new_new_n8112__, new_new_n8113__,
    new_new_n8114__, new_new_n8115__, new_new_n8116__, new_new_n8117__,
    new_new_n8118__, new_new_n8119__, new_new_n8120__, new_new_n8121__,
    new_new_n8122__, new_new_n8123__, new_new_n8124__, new_new_n8125__,
    new_new_n8126__, new_new_n8127__, new_new_n8128__, new_new_n8129__,
    new_new_n8130__, new_new_n8131__, new_new_n8132__, new_new_n8133__,
    new_new_n8134__, new_new_n8135__, new_new_n8136__, new_new_n8137__,
    new_new_n8138__, new_new_n8139__, new_new_n8140__, new_new_n8141__,
    new_new_n8142__, new_new_n8143__, new_new_n8144__, new_new_n8145__,
    new_new_n8146__, new_new_n8147__, new_new_n8148__, new_new_n8149__,
    new_new_n8150__, new_new_n8151__, new_new_n8152__, new_new_n8153__,
    new_new_n8154__, new_new_n8155__, new_new_n8156__, new_new_n8157__,
    new_new_n8158__, new_new_n8159__, new_new_n8160__, new_new_n8161__,
    new_new_n8162__, new_new_n8163__, new_new_n8164__, new_new_n8165__,
    new_new_n8166__, new_new_n8167__, new_new_n8168__, new_new_n8169__,
    new_new_n8170__, new_new_n8171__, new_new_n8172__, new_new_n8173__,
    new_new_n8174__, new_new_n8175__, new_new_n8176__, new_new_n8177__,
    new_new_n8178__, new_new_n8179__, new_new_n8180__, new_new_n8181__,
    new_new_n8182__, new_new_n8183__, new_new_n8184__, new_new_n8185__,
    new_new_n8186__, new_new_n8187__, new_new_n8188__, new_new_n8189__,
    new_new_n8190__, new_new_n8191__, new_new_n8192__, new_new_n8193__,
    new_new_n8194__, new_new_n8195__, new_new_n8196__, new_new_n8197__,
    new_new_n8198__, new_new_n8199__, new_new_n8200__, new_new_n8201__,
    new_new_n8202__, new_new_n8203__, new_new_n8204__, new_new_n8205__,
    new_new_n8206__, new_new_n8207__, new_new_n8208__, new_new_n8209__,
    new_new_n8210__, new_new_n8211__, new_new_n8212__, new_new_n8213__,
    new_new_n8214__, new_new_n8215__, new_new_n8216__, new_new_n8217__,
    new_new_n8218__, new_new_n8219__, new_new_n8220__, new_new_n8221__,
    new_new_n8222__, new_new_n8223__, new_new_n8224__, new_new_n8225__,
    new_new_n8226__, new_new_n8227__, new_new_n8228__, new_new_n8229__,
    new_new_n8230__, new_new_n8231__, new_new_n8232__, new_new_n8233__,
    new_new_n8234__, new_new_n8235__, new_new_n8236__, new_new_n8237__,
    new_new_n8238__, new_new_n8239__, new_new_n8240__, new_new_n8241__,
    new_new_n8242__, new_new_n8243__, new_new_n8244__, new_new_n8245__,
    new_new_n8246__, new_new_n8247__, new_new_n8248__, new_new_n8249__,
    new_new_n8250__, new_new_n8251__, new_new_n8252__, new_new_n8253__,
    new_new_n8254__, new_new_n8255__, new_new_n8256__, new_new_n8257__,
    new_new_n8258__, new_new_n8259__, new_new_n8260__, new_new_n8261__,
    new_new_n8262__, new_new_n8263__, new_new_n8264__, new_new_n8265__,
    new_new_n8266__, new_new_n8267__, new_new_n8268__, new_new_n8269__,
    new_new_n8270__, new_new_n8271__, new_new_n8272__, new_new_n8273__,
    new_new_n8274__, new_new_n8275__, new_new_n8276__, new_new_n8277__,
    new_new_n8278__, new_new_n8279__, new_new_n8280__, new_new_n8281__,
    new_new_n8282__, new_new_n8283__, new_new_n8284__, new_new_n8285__,
    new_new_n8286__, new_new_n8287__, new_new_n8288__, new_new_n8289__,
    new_new_n8290__, new_new_n8291__, new_new_n8292__, new_new_n8293__,
    new_new_n8294__, new_new_n8295__, new_new_n8296__, new_new_n8297__,
    new_new_n8298__, new_new_n8299__, new_new_n8300__, new_new_n8301__,
    new_new_n8302__, new_new_n8303__, new_new_n8304__, new_new_n8305__,
    new_new_n8306__, new_new_n8307__, new_new_n8308__, new_new_n8309__,
    new_new_n8310__, new_new_n8311__, new_new_n8312__, new_new_n8313__,
    new_new_n8314__, new_new_n8315__, new_new_n8316__, new_new_n8317__,
    new_new_n8318__, new_new_n8319__, new_new_n8320__, new_new_n8321__,
    new_new_n8322__, new_new_n8323__, new_new_n8324__, new_new_n8325__,
    new_new_n8326__, new_new_n8327__, new_new_n8328__, new_new_n8329__,
    new_new_n8330__, new_new_n8331__, new_new_n8332__, new_new_n8333__,
    new_new_n8334__, new_new_n8335__, new_new_n8336__, new_new_n8337__,
    new_new_n8338__, new_new_n8339__, new_new_n8340__, new_new_n8341__,
    new_new_n8342__, new_new_n8343__, new_new_n8344__, new_new_n8345__,
    new_new_n8346__, new_new_n8347__, new_new_n8348__, new_new_n8349__,
    new_new_n8350__, new_new_n8351__, new_new_n8352__, new_new_n8353__,
    new_new_n8354__, new_new_n8355__, new_new_n8356__, new_new_n8357__,
    new_new_n8358__, new_new_n8359__, new_new_n8360__, new_new_n8361__,
    new_new_n8362__, new_new_n8363__, new_new_n8364__, new_new_n8365__,
    new_new_n8366__, new_new_n8367__, new_new_n8368__, new_new_n8369__,
    new_new_n8370__, new_new_n8371__, new_new_n8372__, new_new_n8373__,
    new_new_n8374__, new_new_n8375__, new_new_n8376__, new_new_n8377__,
    new_new_n8378__, new_new_n8379__, new_new_n8380__, new_new_n8381__,
    new_new_n8382__, new_new_n8383__, new_new_n8384__, new_new_n8385__,
    new_new_n8386__, new_new_n8387__, new_new_n8388__, new_new_n8389__,
    new_new_n8390__, new_new_n8391__, new_new_n8392__, new_new_n8393__,
    new_new_n8394__, new_new_n8395__, new_new_n8396__, new_new_n8397__,
    new_new_n8398__, new_new_n8399__, new_new_n8400__, new_new_n8401__,
    new_new_n8402__, new_new_n8403__, new_new_n8404__, new_new_n8405__,
    new_new_n8406__, new_new_n8407__, new_new_n8408__, new_new_n8409__,
    new_new_n8410__, new_new_n8411__, new_new_n8412__, new_new_n8413__,
    new_new_n8414__, new_new_n8415__, new_new_n8416__, new_new_n8417__,
    new_new_n8418__, new_new_n8419__, new_new_n8420__, new_new_n8421__,
    new_new_n8422__, new_new_n8423__, new_new_n8424__, new_new_n8425__,
    new_new_n8426__, new_new_n8427__, new_new_n8428__, new_new_n8429__,
    new_new_n8430__, new_new_n8431__, new_new_n8432__, new_new_n8433__,
    new_new_n8434__, new_new_n8435__, new_new_n8436__, new_new_n8437__,
    new_new_n8438__, new_new_n8439__, new_new_n8440__, new_new_n8441__,
    new_new_n8442__, new_new_n8443__, new_new_n8444__, new_new_n8445__,
    new_new_n8446__, new_new_n8447__, new_new_n8448__, new_new_n8449__,
    new_new_n8450__, new_new_n8451__, new_new_n8452__, new_new_n8453__,
    new_new_n8454__, new_new_n8455__, new_new_n8456__, new_new_n8457__,
    new_new_n8458__, new_new_n8459__, new_new_n8460__, new_new_n8461__,
    new_new_n8462__, new_new_n8463__, new_new_n8464__, new_new_n8465__,
    new_new_n8466__, new_new_n8467__, new_new_n8468__, new_new_n8469__,
    new_new_n8470__, new_new_n8471__, new_new_n8472__, new_new_n8473__,
    new_new_n8474__, new_new_n8475__, new_new_n8476__, new_new_n8477__,
    new_new_n8478__, new_new_n8479__, new_new_n8480__, new_new_n8481__,
    new_new_n8482__, new_new_n8483__, new_new_n8484__, new_new_n8485__,
    new_new_n8486__, new_new_n8487__, new_new_n8488__, new_new_n8489__,
    new_new_n8490__, new_new_n8491__, new_new_n8492__, new_new_n8493__,
    new_new_n8494__, new_new_n8495__, new_new_n8496__, new_new_n8497__,
    new_new_n8498__, new_new_n8499__, new_new_n8500__, new_new_n8501__,
    new_new_n8502__, new_new_n8503__, new_new_n8504__, new_new_n8505__,
    new_new_n8506__, new_new_n8507__, new_new_n8508__, new_new_n8509__,
    new_new_n8510__, new_new_n8511__, new_new_n8512__, new_new_n8513__,
    new_new_n8514__, new_new_n8515__, new_new_n8516__, new_new_n8517__,
    new_new_n8518__, new_new_n8519__, new_new_n8520__, new_new_n8521__,
    new_new_n8522__, new_new_n8523__, new_new_n8524__, new_new_n8525__,
    new_new_n8526__, new_new_n8527__, new_new_n8528__, new_new_n8529__,
    new_new_n8530__, new_new_n8531__, new_new_n8532__, new_new_n8533__,
    new_new_n8534__, new_new_n8535__, new_new_n8536__, new_new_n8537__,
    new_new_n8538__, new_new_n8539__, new_new_n8540__, new_new_n8541__,
    new_new_n8542__, new_new_n8543__, new_new_n8544__, new_new_n8545__,
    new_new_n8546__, new_new_n8547__, new_new_n8548__, new_new_n8549__,
    new_new_n8550__, new_new_n8551__, new_new_n8552__, new_new_n8553__,
    new_new_n8554__, new_new_n8555__, new_new_n8556__, new_new_n8557__,
    new_new_n8558__, new_new_n8559__, new_new_n8560__, new_new_n8561__,
    new_new_n8562__, new_new_n8563__, new_new_n8564__, new_new_n8565__,
    new_new_n8566__, new_new_n8567__, new_new_n8568__, new_new_n8569__,
    new_new_n8570__, new_new_n8571__, new_new_n8572__, new_new_n8573__,
    new_new_n8574__, new_new_n8575__, new_new_n8576__, new_new_n8577__,
    new_new_n8578__, new_new_n8579__, new_new_n8580__, new_new_n8581__,
    new_new_n8582__, new_new_n8583__, new_new_n8584__, new_new_n8585__,
    new_new_n8586__, new_new_n8587__, new_new_n8588__, new_new_n8589__,
    new_new_n8590__, new_new_n8591__, new_new_n8592__, new_new_n8593__,
    new_new_n8594__, new_new_n8595__, new_new_n8596__, new_new_n8597__,
    new_new_n8598__, new_new_n8599__, new_new_n8600__, new_new_n8601__,
    new_new_n8602__, new_new_n8603__, new_new_n8604__, new_new_n8605__,
    new_new_n8606__, new_new_n8607__, new_new_n8608__, new_new_n8609__,
    new_new_n8610__, new_new_n8611__, new_new_n8612__, new_new_n8613__,
    new_new_n8614__, new_new_n8615__, new_new_n8616__, new_new_n8617__,
    new_new_n8618__, new_new_n8619__, new_new_n8620__, new_new_n8621__,
    new_new_n8622__, new_new_n8623__, new_new_n8624__, new_new_n8625__,
    new_new_n8626__, new_new_n8627__, new_new_n8628__, new_new_n8629__,
    new_new_n8630__, new_new_n8631__, new_new_n8632__, new_new_n8633__,
    new_new_n8634__, new_new_n8635__, new_new_n8636__, new_new_n8637__,
    new_new_n8638__, new_new_n8639__, new_new_n8640__, new_new_n8641__,
    new_new_n8642__, new_new_n8643__, new_new_n8644__, new_new_n8645__,
    new_new_n8646__, new_new_n8647__, new_new_n8648__, new_new_n8649__,
    new_new_n8650__, new_new_n8651__, new_new_n8652__, new_new_n8653__,
    new_new_n8654__, new_new_n8655__, new_new_n8656__, new_new_n8657__,
    new_new_n8658__, new_new_n8659__, new_new_n8660__, new_new_n8661__,
    new_new_n8662__, new_new_n8663__, new_new_n8664__, new_new_n8665__,
    new_new_n8666__, new_new_n8667__, new_new_n8668__, new_new_n8669__,
    new_new_n8670__, new_new_n8671__, new_new_n8672__, new_new_n8673__,
    new_new_n8674__, new_new_n8675__, new_new_n8676__, new_new_n8677__,
    new_new_n8678__, new_new_n8679__, new_new_n8680__, new_new_n8681__,
    new_new_n8682__, new_new_n8683__, new_new_n8684__, new_new_n8685__,
    new_new_n8686__, new_new_n8687__, new_new_n8688__, new_new_n8689__,
    new_new_n8690__, new_new_n8691__, new_new_n8692__, new_new_n8693__,
    new_new_n8694__, new_new_n8695__, new_new_n8696__, new_new_n8697__,
    new_new_n8698__, new_new_n8699__, new_new_n8700__, new_new_n8701__,
    new_new_n8702__, new_new_n8703__, new_new_n8704__, new_new_n8705__,
    new_new_n8706__, new_new_n8707__, new_new_n8708__, new_new_n8709__,
    new_new_n8710__, new_new_n8711__, new_new_n8712__, new_new_n8713__,
    new_new_n8714__, new_new_n8715__, new_new_n8716__, new_new_n8717__,
    new_new_n8718__, new_new_n8719__, new_new_n8720__, new_new_n8721__,
    new_new_n8722__, new_new_n8723__, new_new_n8724__, new_new_n8725__,
    new_new_n8726__, new_new_n8727__, new_new_n8728__, new_new_n8729__,
    new_new_n8730__, new_new_n8731__, new_new_n8732__, new_new_n8733__,
    new_new_n8734__, new_new_n8735__, new_new_n8736__, new_new_n8737__,
    new_new_n8738__, new_new_n8739__, new_new_n8740__, new_new_n8741__,
    new_new_n8742__, new_new_n8743__, new_new_n8744__, new_new_n8745__,
    new_new_n8746__, new_new_n8747__, new_new_n8748__, new_new_n8749__,
    new_new_n8750__, new_new_n8751__, new_new_n8752__, new_new_n8753__,
    new_new_n8754__, new_new_n8755__, new_new_n8756__, new_new_n8757__,
    new_new_n8758__, new_new_n8759__, new_new_n8760__, new_new_n8761__,
    new_new_n8762__, new_new_n8763__, new_new_n8764__, new_new_n8765__,
    new_new_n8766__, new_new_n8767__, new_new_n8768__, new_new_n8769__,
    new_new_n8770__, new_new_n8771__, new_new_n8772__, new_new_n8773__,
    new_new_n8774__, new_new_n8775__, new_new_n8776__, new_new_n8777__,
    new_new_n8778__, new_new_n8779__, new_new_n8780__, new_new_n8781__,
    new_new_n8782__, new_new_n8783__, new_new_n8784__, new_new_n8785__,
    new_new_n8786__, new_new_n8787__, new_new_n8788__, new_new_n8789__,
    new_new_n8790__, new_new_n8791__, new_new_n8792__, new_new_n8793__,
    new_new_n8794__, new_new_n8795__, new_new_n8796__, new_new_n8797__,
    new_new_n8798__, new_new_n8799__, new_new_n8800__, new_new_n8801__,
    new_new_n8802__, new_new_n8803__, new_new_n8804__, new_new_n8805__,
    new_new_n8806__, new_new_n8807__, new_new_n8808__, new_new_n8809__,
    new_new_n8810__, new_new_n8811__, new_new_n8812__, new_new_n8813__,
    new_new_n8814__, new_new_n8815__, new_new_n8816__, new_new_n8817__,
    new_new_n8818__, new_new_n8819__, new_new_n8820__, new_new_n8821__,
    new_new_n8822__, new_new_n8823__, new_new_n8824__, new_new_n8825__,
    new_new_n8826__, new_new_n8827__, new_new_n8828__, new_new_n8829__,
    new_new_n8830__, new_new_n8831__, new_new_n8832__, new_new_n8833__,
    new_new_n8834__, new_new_n8835__, new_new_n8836__, new_new_n8837__,
    new_new_n8838__, new_new_n8839__, new_new_n8840__, new_new_n8841__,
    new_new_n8842__, new_new_n8843__, new_new_n8844__, new_new_n8845__,
    new_new_n8846__, new_new_n8847__, new_new_n8848__, new_new_n8849__,
    new_new_n8850__, new_new_n8851__, new_new_n8852__, new_new_n8853__,
    new_new_n8854__, new_new_n8855__, new_new_n8856__, new_new_n8857__,
    new_new_n8858__, new_new_n8859__, new_new_n8860__, new_new_n8861__,
    new_new_n8862__, new_new_n8863__, new_new_n8864__, new_new_n8865__,
    new_new_n8866__, new_new_n8867__, new_new_n8868__, new_new_n8869__,
    new_new_n8870__, new_new_n8871__, new_new_n8872__, new_new_n8873__,
    new_new_n8874__, new_new_n8875__, new_new_n8876__, new_new_n8877__,
    new_new_n8878__, new_new_n8879__, new_new_n8880__, new_new_n8881__,
    new_new_n8882__, new_new_n8883__, new_new_n8884__, new_new_n8885__,
    new_new_n8886__, new_new_n8887__, new_new_n8888__, new_new_n8889__,
    new_new_n8890__, new_new_n8891__, new_new_n8892__, new_new_n8893__,
    new_new_n8894__, new_new_n8895__, new_new_n8896__, new_new_n8897__,
    new_new_n8898__, new_new_n8899__, new_new_n8900__, new_new_n8901__,
    new_new_n8902__, new_new_n8903__, new_new_n8904__, new_new_n8905__,
    new_new_n8906__, new_new_n8907__, new_new_n8908__, new_new_n8909__,
    new_new_n8910__, new_new_n8911__, new_new_n8912__, new_new_n8913__,
    new_new_n8914__, new_new_n8915__, new_new_n8916__, new_new_n8917__,
    new_new_n8918__, new_new_n8919__, new_new_n8920__, new_new_n8921__,
    new_new_n8922__, new_new_n8923__, new_new_n8924__, new_new_n8925__,
    new_new_n8926__, new_new_n8927__, new_new_n8928__, new_new_n8929__,
    new_new_n8930__, new_new_n8931__, new_new_n8932__, new_new_n8933__,
    new_new_n8934__, new_new_n8935__, new_new_n8936__, new_new_n8937__,
    new_new_n8938__, new_new_n8939__, new_new_n8940__, new_new_n8941__,
    new_new_n8942__, new_new_n8943__, new_new_n8944__, new_new_n8945__,
    new_new_n8946__, new_new_n8947__, new_new_n8948__, new_new_n8949__,
    new_new_n8950__, new_new_n8951__, new_new_n8952__, new_new_n8953__,
    new_new_n8954__, new_new_n8955__, new_new_n8956__, new_new_n8957__,
    new_new_n8958__, new_new_n8959__, new_new_n8960__, new_new_n8961__,
    new_new_n8962__, new_new_n8963__, new_new_n8964__, new_new_n8965__,
    new_new_n8966__, new_new_n8967__, new_new_n8968__, new_new_n8969__,
    new_new_n8970__, new_new_n8971__, new_new_n8972__, new_new_n8973__,
    new_new_n8974__, new_new_n8975__, new_new_n8976__, new_new_n8977__,
    new_new_n8978__, new_new_n8979__, new_new_n8980__, new_new_n8981__,
    new_new_n8982__, new_new_n8983__, new_new_n8984__, new_new_n8985__,
    new_new_n8986__, new_new_n8987__, new_new_n8988__, new_new_n8989__,
    new_new_n8990__, new_new_n8991__, new_new_n8992__, new_new_n8993__,
    new_new_n8994__, new_new_n8995__, new_new_n8996__, new_new_n8997__,
    new_new_n8998__, new_new_n8999__, new_new_n9000__, new_new_n9001__,
    new_new_n9002__, new_new_n9003__, new_new_n9004__, new_new_n9005__,
    new_new_n9006__, new_new_n9007__, new_new_n9008__, new_new_n9009__,
    new_new_n9010__, new_new_n9011__, new_new_n9012__, new_new_n9013__,
    new_new_n9014__, new_new_n9015__, new_new_n9016__, new_new_n9017__,
    new_new_n9018__, new_new_n9019__, new_new_n9020__, new_new_n9021__,
    new_new_n9022__, new_new_n9023__, new_new_n9024__, new_new_n9025__,
    new_new_n9026__, new_new_n9027__, new_new_n9028__, new_new_n9029__,
    new_new_n9030__, new_new_n9031__, new_new_n9032__, new_new_n9033__,
    new_new_n9034__, new_new_n9035__, new_new_n9036__, new_new_n9037__,
    new_new_n9038__, new_new_n9039__, new_new_n9040__, new_new_n9041__,
    new_new_n9042__, new_new_n9043__, new_new_n9044__, new_new_n9045__,
    new_new_n9046__, new_new_n9047__, new_new_n9048__, new_new_n9049__,
    new_new_n9050__, new_new_n9051__, new_new_n9052__, new_new_n9053__,
    new_new_n9054__, new_new_n9055__, new_new_n9056__, new_new_n9057__,
    new_new_n9058__, new_new_n9059__, new_new_n9060__, new_new_n9061__,
    new_new_n9062__, new_new_n9063__, new_new_n9064__, new_new_n9065__,
    new_new_n9066__, new_new_n9067__, new_new_n9068__, new_new_n9069__,
    new_new_n9070__, new_new_n9071__, new_new_n9072__, new_new_n9073__,
    new_new_n9074__, new_new_n9075__, new_new_n9076__, new_new_n9077__,
    new_new_n9078__, new_new_n9079__, new_new_n9080__, new_new_n9081__,
    new_new_n9082__, new_new_n9083__, new_new_n9084__, new_new_n9085__,
    new_new_n9086__, new_new_n9087__, new_new_n9088__, new_new_n9089__,
    new_new_n9090__, new_new_n9091__, new_new_n9092__, new_new_n9093__,
    new_new_n9094__, new_new_n9095__, new_new_n9096__, new_new_n9097__,
    new_new_n9098__, new_new_n9099__, new_new_n9100__, new_new_n9101__,
    new_new_n9102__, new_new_n9103__, new_new_n9104__, new_new_n9105__,
    new_new_n9106__, new_new_n9107__, new_new_n9108__, new_new_n9109__,
    new_new_n9110__, new_new_n9111__, new_new_n9112__, new_new_n9113__,
    new_new_n9114__, new_new_n9115__, new_new_n9116__, new_new_n9117__,
    new_new_n9118__, new_new_n9119__, new_new_n9120__, new_new_n9121__,
    new_new_n9122__, new_new_n9123__, new_new_n9124__, new_new_n9125__,
    new_new_n9126__, new_new_n9127__, new_new_n9128__, new_new_n9129__,
    new_new_n9130__, new_new_n9131__, new_new_n9132__, new_new_n9133__,
    new_new_n9134__, new_new_n9135__, new_new_n9136__, new_new_n9137__,
    new_new_n9138__, new_new_n9139__, new_new_n9140__, new_new_n9141__,
    new_new_n9142__, new_new_n9143__, new_new_n9144__, new_new_n9145__,
    new_new_n9146__, new_new_n9147__, new_new_n9148__, new_new_n9149__,
    new_new_n9150__, new_new_n9151__, new_new_n9152__, new_new_n9153__,
    new_new_n9154__, new_new_n9155__, new_new_n9156__, new_new_n9157__,
    new_new_n9158__, new_new_n9159__, new_new_n9160__, new_new_n9161__,
    new_new_n9162__, new_new_n9163__, new_new_n9164__, new_new_n9165__,
    new_new_n9166__, new_new_n9167__, new_new_n9168__, new_new_n9169__,
    new_new_n9170__, new_new_n9171__, new_new_n9172__, new_new_n9173__,
    new_new_n9174__, new_new_n9175__, new_new_n9176__, new_new_n9177__,
    new_new_n9178__, new_new_n9179__, new_new_n9180__, new_new_n9181__,
    new_new_n9182__, new_new_n9183__, new_new_n9184__, new_new_n9185__,
    new_new_n9186__, new_new_n9187__, new_new_n9188__, new_new_n9189__,
    new_new_n9190__, new_new_n9191__, new_new_n9192__, new_new_n9193__,
    new_new_n9194__, new_new_n9195__, new_new_n9196__, new_new_n9197__,
    new_new_n9198__, new_new_n9199__, new_new_n9200__, new_new_n9201__,
    new_new_n9202__, new_new_n9203__, new_new_n9204__, new_new_n9205__,
    new_new_n9206__, new_new_n9207__, new_new_n9208__, new_new_n9209__,
    new_new_n9210__, new_new_n9211__, new_new_n9212__, new_new_n9213__,
    new_new_n9214__, new_new_n9215__, new_new_n9216__, new_new_n9217__,
    new_new_n9218__, new_new_n9219__, new_new_n9220__, new_new_n9221__,
    new_new_n9222__, new_new_n9223__, new_new_n9224__, new_new_n9225__,
    new_new_n9226__, new_new_n9227__, new_new_n9228__, new_new_n9229__,
    new_new_n9230__, new_new_n9231__, new_new_n9232__, new_new_n9233__,
    new_new_n9234__, new_new_n9235__, new_new_n9236__, new_new_n9237__,
    new_new_n9238__, new_new_n9239__, new_new_n9240__, new_new_n9241__,
    new_new_n9242__, new_new_n9243__, new_new_n9244__, new_new_n9245__,
    new_new_n9246__, new_new_n9247__, new_new_n9248__, new_new_n9249__,
    new_new_n9250__, new_new_n9251__, new_new_n9252__, new_new_n9253__,
    new_new_n9254__, new_new_n9255__, new_new_n9256__, new_new_n9257__,
    new_new_n9258__, new_new_n9259__, new_new_n9260__, new_new_n9261__,
    new_new_n9262__, new_new_n9263__, new_new_n9264__, new_new_n9265__,
    new_new_n9266__, new_new_n9267__, new_new_n9268__, new_new_n9269__,
    new_new_n9270__, new_new_n9271__, new_new_n9272__, new_new_n9273__,
    new_new_n9274__, new_new_n9275__, new_new_n9276__, new_new_n9277__,
    new_new_n9278__, new_new_n9279__, new_new_n9280__, new_new_n9281__,
    new_new_n9282__, new_new_n9283__, new_new_n9284__, new_new_n9285__,
    new_new_n9286__, new_new_n9287__, new_new_n9288__, new_new_n9289__,
    new_new_n9290__, new_new_n9291__, new_new_n9292__, new_new_n9293__,
    new_new_n9294__, new_new_n9295__, new_new_n9296__, new_new_n9297__,
    new_new_n9298__, new_new_n9299__, new_new_n9300__, new_new_n9301__,
    new_new_n9302__, new_new_n9303__, new_new_n9304__, new_new_n9305__,
    new_new_n9306__, new_new_n9307__, new_new_n9308__, new_new_n9309__,
    new_new_n9310__, new_new_n9311__, new_new_n9312__, new_new_n9313__,
    new_new_n9314__, new_new_n9315__, new_new_n9316__, new_new_n9317__,
    new_new_n9318__, new_new_n9319__, new_new_n9320__, new_new_n9321__,
    new_new_n9322__, new_new_n9323__, new_new_n9324__, new_new_n9325__,
    new_new_n9326__, new_new_n9327__, new_new_n9328__, new_new_n9329__,
    new_new_n9330__, new_new_n9331__, new_new_n9332__, new_new_n9333__,
    new_new_n9334__, new_new_n9335__, new_new_n9336__, new_new_n9337__,
    new_new_n9338__, new_new_n9339__, new_new_n9340__, new_new_n9341__,
    new_new_n9342__, new_new_n9343__, new_new_n9344__, new_new_n9345__,
    new_new_n9346__, new_new_n9347__, new_new_n9348__, new_new_n9349__,
    new_new_n9350__, new_new_n9351__, new_new_n9352__, new_new_n9353__,
    new_new_n9354__, new_new_n9355__, new_new_n9356__, new_new_n9357__,
    new_new_n9358__, new_new_n9359__, new_new_n9360__, new_new_n9361__,
    new_new_n9362__, new_new_n9363__, new_new_n9364__, new_new_n9365__,
    new_new_n9366__, new_new_n9367__, new_new_n9368__, new_new_n9369__,
    new_new_n9370__, new_new_n9371__, new_new_n9372__, new_new_n9373__,
    new_new_n9374__, new_new_n9375__, new_new_n9376__, new_new_n9377__,
    new_new_n9378__, new_new_n9379__, new_new_n9380__, new_new_n9381__,
    new_new_n9382__, new_new_n9383__, new_new_n9384__, new_new_n9385__,
    new_new_n9386__, new_new_n9387__, new_new_n9388__, new_new_n9389__,
    new_new_n9390__, new_new_n9391__, new_new_n9392__, new_new_n9393__,
    new_new_n9394__, new_new_n9395__, new_new_n9396__, new_new_n9397__,
    new_new_n9398__, new_new_n9399__, new_new_n9400__, new_new_n9401__,
    new_new_n9402__, new_new_n9403__, new_new_n9404__, new_new_n9405__,
    new_new_n9406__, new_new_n9407__, new_new_n9408__, new_new_n9409__,
    new_new_n9410__, new_new_n9411__, new_new_n9412__, new_new_n9413__,
    new_new_n9414__, new_new_n9415__, new_new_n9416__, new_new_n9417__,
    new_new_n9418__, new_new_n9419__, new_new_n9420__, new_new_n9421__,
    new_new_n9422__, new_new_n9423__, new_new_n9424__, new_new_n9425__,
    new_new_n9426__, new_new_n9427__, new_new_n9428__, new_new_n9429__,
    new_new_n9430__, new_new_n9431__, new_new_n9432__, new_new_n9433__,
    new_new_n9434__, new_new_n9435__, new_new_n9436__, new_new_n9437__,
    new_new_n9438__, new_new_n9439__, new_new_n9440__, new_new_n9441__,
    new_new_n9442__, new_new_n9443__, new_new_n9444__, new_new_n9445__,
    new_new_n9446__, new_new_n9447__, new_new_n9448__, new_new_n9449__,
    new_new_n9450__, new_new_n9451__, new_new_n9452__, new_new_n9453__,
    new_new_n9454__, new_new_n9455__, new_new_n9456__, new_new_n9457__,
    new_new_n9458__, new_new_n9459__, new_new_n9460__, new_new_n9461__,
    new_new_n9462__, new_new_n9463__, new_new_n9464__, new_new_n9465__,
    new_new_n9466__, new_new_n9467__, new_new_n9468__, new_new_n9469__,
    new_new_n9470__, new_new_n9471__, new_new_n9472__, new_new_n9473__,
    new_new_n9474__, new_new_n9475__, new_new_n9476__, new_new_n9477__,
    new_new_n9478__, new_new_n9479__, new_new_n9480__, new_new_n9481__,
    new_new_n9482__, new_new_n9483__, new_new_n9484__, new_new_n9485__,
    new_new_n9486__, new_new_n9487__, new_new_n9488__, new_new_n9489__,
    new_new_n9490__, new_new_n9491__, new_new_n9492__, new_new_n9493__,
    new_new_n9494__, new_new_n9495__, new_new_n9496__, new_new_n9497__,
    new_new_n9498__, new_new_n9499__, new_new_n9500__, new_new_n9501__,
    new_new_n9502__, new_new_n9503__, new_new_n9504__, new_new_n9505__,
    new_new_n9506__, new_new_n9507__, new_new_n9508__, new_new_n9509__,
    new_new_n9510__, new_new_n9511__, new_new_n9512__, new_new_n9513__,
    new_new_n9514__, new_new_n9515__, new_new_n9516__, new_new_n9517__,
    new_new_n9518__, new_new_n9519__, new_new_n9520__, new_new_n9521__,
    new_new_n9522__, new_new_n9523__, new_new_n9524__, new_new_n9525__,
    new_new_n9526__, new_new_n9527__, new_new_n9528__, new_new_n9529__,
    new_new_n9530__, new_new_n9531__, new_new_n9532__, new_new_n9533__,
    new_new_n9534__, new_new_n9535__, new_new_n9536__, new_new_n9537__,
    new_new_n9538__, new_new_n9539__, new_new_n9540__, new_new_n9541__,
    new_new_n9542__, new_new_n9543__, new_new_n9544__, new_new_n9545__,
    new_new_n9546__, new_new_n9547__, new_new_n9548__, new_new_n9549__,
    new_new_n9550__, new_new_n9551__, new_new_n9552__, new_new_n9553__,
    new_new_n9554__, new_new_n9555__, new_new_n9556__, new_new_n9557__,
    new_new_n9558__, new_new_n9559__, new_new_n9560__, new_new_n9561__,
    new_new_n9562__, new_new_n9563__, new_new_n9564__, new_new_n9565__,
    new_new_n9566__, new_new_n9567__, new_new_n9568__, new_new_n9569__,
    new_new_n9570__, new_new_n9571__, new_new_n9572__, new_new_n9573__,
    new_new_n9574__, new_new_n9575__, new_new_n9576__, new_new_n9577__,
    new_new_n9578__, new_new_n9579__, new_new_n9580__, new_new_n9581__,
    new_new_n9582__, new_new_n9583__, new_new_n9584__, new_new_n9585__,
    new_new_n9586__, new_new_n9587__, new_new_n9588__, new_new_n9589__,
    new_new_n9590__, new_new_n9591__, new_new_n9592__, new_new_n9593__,
    new_new_n9594__, new_new_n9595__, new_new_n9596__, new_new_n9597__,
    new_new_n9598__, new_new_n9599__, new_new_n9600__, new_new_n9601__,
    new_new_n9602__, new_new_n9603__, new_new_n9604__, new_new_n9605__,
    new_new_n9606__, new_new_n9607__, new_new_n9608__, new_new_n9609__,
    new_new_n9610__, new_new_n9611__, new_new_n9612__, new_new_n9613__,
    new_new_n9614__, new_new_n9615__, new_new_n9616__, new_new_n9617__,
    new_new_n9618__, new_new_n9619__, new_new_n9620__, new_new_n9621__,
    new_new_n9622__, new_new_n9623__, new_new_n9624__, new_new_n9625__,
    new_new_n9626__, new_new_n9627__, new_new_n9628__, new_new_n9629__,
    new_new_n9630__, new_new_n9631__, new_new_n9632__, new_new_n9633__,
    new_new_n9634__, new_new_n9635__, new_new_n9636__, new_new_n9637__,
    new_new_n9638__, new_new_n9639__, new_new_n9640__, new_new_n9641__,
    new_new_n9642__, new_new_n9643__, new_new_n9644__, new_new_n9645__,
    new_new_n9646__, new_new_n9647__, new_new_n9648__, new_new_n9649__,
    new_new_n9650__, new_new_n9651__, new_new_n9652__, new_new_n9653__,
    new_new_n9654__, new_new_n9655__, new_new_n9656__, new_new_n9657__,
    new_new_n9658__, new_new_n9659__, new_new_n9660__, new_new_n9661__,
    new_new_n9662__, new_new_n9663__, new_new_n9664__, new_new_n9665__,
    new_new_n9666__, new_new_n9667__, new_new_n9668__, new_new_n9669__,
    new_new_n9670__, new_new_n9671__, new_new_n9672__, new_new_n9673__,
    new_new_n9674__, new_new_n9675__, new_new_n9676__, new_new_n9677__,
    new_new_n9678__, new_new_n9679__, new_new_n9680__, new_new_n9681__,
    new_new_n9682__, new_new_n9683__, new_new_n9684__, new_new_n9685__,
    new_new_n9686__, new_new_n9687__, new_new_n9688__, new_new_n9689__,
    new_new_n9690__, new_new_n9691__, new_new_n9692__, new_new_n9693__,
    new_new_n9694__, new_new_n9695__, new_new_n9696__, new_new_n9697__,
    new_new_n9698__, new_new_n9699__, new_new_n9700__, new_new_n9701__,
    new_new_n9702__, new_new_n9703__, new_new_n9704__, new_new_n9705__,
    new_new_n9706__, new_new_n9707__, new_new_n9708__, new_new_n9709__,
    new_new_n9710__, new_new_n9711__, new_new_n9712__, new_new_n9713__,
    new_new_n9714__, new_new_n9715__, new_new_n9716__, new_new_n9717__,
    new_new_n9718__, new_new_n9719__, new_new_n9720__, new_new_n9721__,
    new_new_n9722__, new_new_n9723__, new_new_n9724__, new_new_n9725__,
    new_new_n9726__, new_new_n9727__, new_new_n9728__, new_new_n9729__,
    new_new_n9730__, new_new_n9731__, new_new_n9732__, new_new_n9733__,
    new_new_n9734__, new_new_n9735__, new_new_n9736__, new_new_n9737__,
    new_new_n9738__, new_new_n9739__, new_new_n9740__, new_new_n9741__,
    new_new_n9742__, new_new_n9743__, new_new_n9744__, new_new_n9745__,
    new_new_n9746__, new_new_n9747__, new_new_n9748__, new_new_n9749__,
    new_new_n9750__, new_new_n9751__, new_new_n9752__, new_new_n9753__,
    new_new_n9754__, new_new_n9755__, new_new_n9756__, new_new_n9757__,
    new_new_n9758__, new_new_n9759__, new_new_n9760__, new_new_n9761__,
    new_new_n9762__, new_new_n9763__, new_new_n9764__, new_new_n9765__,
    new_new_n9766__, new_new_n9767__, new_new_n9768__, new_new_n9769__,
    new_new_n9770__, new_new_n9771__, new_new_n9772__, new_new_n9773__,
    new_new_n9774__, new_new_n9775__, new_new_n9776__, new_new_n9777__,
    new_new_n9778__, new_new_n9779__, new_new_n9780__, new_new_n9781__,
    new_new_n9782__, new_new_n9783__, new_new_n9784__, new_new_n9785__,
    new_new_n9786__, new_new_n9787__, new_new_n9788__, new_new_n9789__,
    new_new_n9790__, new_new_n9791__, new_new_n9792__, new_new_n9793__,
    new_new_n9794__, new_new_n9795__, new_new_n9796__, new_new_n9797__,
    new_new_n9798__, new_new_n9799__, new_new_n9800__, new_new_n9801__,
    new_new_n9802__, new_new_n9803__, new_new_n9804__, new_new_n9805__,
    new_new_n9806__, new_new_n9807__, new_new_n9808__, new_new_n9809__,
    new_new_n9810__, new_new_n9811__, new_new_n9812__, new_new_n9813__,
    new_new_n9814__, new_new_n9815__, new_new_n9816__, new_new_n9817__,
    new_new_n9818__, new_new_n9819__, new_new_n9820__, new_new_n9821__,
    new_new_n9822__, new_new_n9823__, new_new_n9824__, new_new_n9825__,
    new_new_n9826__, new_new_n9827__, new_new_n9828__, new_new_n9829__,
    new_new_n9830__, new_new_n9831__, new_new_n9832__, new_new_n9833__,
    new_new_n9834__, new_new_n9835__, new_new_n9836__, new_new_n9837__,
    new_new_n9838__, new_new_n9839__, new_new_n9840__, new_new_n9841__,
    new_new_n9842__, new_new_n9843__, new_new_n9844__, new_new_n9845__,
    new_new_n9846__, new_new_n9847__, new_new_n9848__, new_new_n9849__,
    new_new_n9850__, new_new_n9851__, new_new_n9852__, new_new_n9853__,
    new_new_n9854__, new_new_n9855__, new_new_n9856__, new_new_n9857__,
    new_new_n9858__, new_new_n9859__, new_new_n9860__, new_new_n9861__,
    new_new_n9862__, new_new_n9863__, new_new_n9864__, new_new_n9865__,
    new_new_n9866__, new_new_n9867__, new_new_n9868__, new_new_n9869__,
    new_new_n9870__, new_new_n9871__, new_new_n9872__, new_new_n9873__,
    new_new_n9874__, new_new_n9875__, new_new_n9876__, new_new_n9877__,
    new_new_n9878__, new_new_n9879__, new_new_n9880__, new_new_n9881__,
    new_new_n9882__, new_new_n9883__, new_new_n9884__, new_new_n9885__,
    new_new_n9886__, new_new_n9887__, new_new_n9888__, new_new_n9889__,
    new_new_n9890__, new_new_n9891__, new_new_n9892__, new_new_n9893__,
    new_new_n9894__, new_new_n9895__, new_new_n9896__, new_new_n9897__,
    new_new_n9898__, new_new_n9899__, new_new_n9900__, new_new_n9901__,
    new_new_n9902__, new_new_n9903__, new_new_n9904__, new_new_n9905__,
    new_new_n9906__, new_new_n9907__, new_new_n9908__, new_new_n9909__,
    new_new_n9910__, new_new_n9911__, new_new_n9912__, new_new_n9913__,
    new_new_n9914__, new_new_n9915__, new_new_n9916__, new_new_n9917__,
    new_new_n9918__, new_new_n9919__, new_new_n9920__, new_new_n9921__,
    new_new_n9922__, new_new_n9923__, new_new_n9924__, new_new_n9925__,
    new_new_n9926__, new_new_n9927__, new_new_n9928__, new_new_n9929__,
    new_new_n9930__, new_new_n9931__, new_new_n9932__, new_new_n9933__,
    new_new_n9934__, new_new_n9935__, new_new_n9936__, new_new_n9937__,
    new_new_n9938__, new_new_n9939__, new_new_n9940__, new_new_n9941__,
    new_new_n9942__, new_new_n9943__, new_new_n9944__, new_new_n9945__,
    new_new_n9946__, new_new_n9947__, new_new_n9948__, new_new_n9949__,
    new_new_n9950__, new_new_n9951__, new_new_n9952__, new_new_n9953__,
    new_new_n9954__, new_new_n9955__, new_new_n9956__, new_new_n9957__,
    new_new_n9958__, new_new_n9959__, new_new_n9960__, new_new_n9961__,
    new_new_n9962__, new_new_n9963__, new_new_n9964__, new_new_n9965__,
    new_new_n9966__, new_new_n9967__, new_new_n9968__, new_new_n9969__,
    new_new_n9970__, new_new_n9971__, new_new_n9972__, new_new_n9973__,
    new_new_n9974__, new_new_n9975__, new_new_n9976__, new_new_n9977__,
    new_new_n9978__, new_new_n9979__, new_new_n9980__, new_new_n9981__,
    new_new_n9982__, new_new_n9983__, new_new_n9984__, new_new_n9985__,
    new_new_n9986__, new_new_n9987__, new_new_n9988__, new_new_n9989__,
    new_new_n9990__, new_new_n9991__, new_new_n9992__, new_new_n9993__,
    new_new_n9994__, new_new_n9995__, new_new_n9996__, new_new_n9997__,
    new_new_n9998__, new_new_n9999__, new_new_n10000__, new_new_n10001__,
    new_new_n10002__, new_new_n10003__, new_new_n10004__, new_new_n10005__,
    new_new_n10006__, new_new_n10007__, new_new_n10008__, new_new_n10009__,
    new_new_n10010__, new_new_n10011__, new_new_n10012__, new_new_n10013__,
    new_new_n10014__, new_new_n10015__, new_new_n10016__, new_new_n10017__,
    new_new_n10018__, new_new_n10019__, new_new_n10020__, new_new_n10021__,
    new_new_n10022__, new_new_n10023__, new_new_n10024__, new_new_n10025__,
    new_new_n10026__, new_new_n10027__, new_new_n10028__, new_new_n10029__,
    new_new_n10030__, new_new_n10031__, new_new_n10032__, new_new_n10033__,
    new_new_n10034__, new_new_n10035__, new_new_n10036__, new_new_n10037__,
    new_new_n10038__, new_new_n10039__, new_new_n10040__, new_new_n10041__,
    new_new_n10042__, new_new_n10043__, new_new_n10044__, new_new_n10045__,
    new_new_n10046__, new_new_n10047__, new_new_n10048__, new_new_n10049__,
    new_new_n10050__, new_new_n10051__, new_new_n10052__, new_new_n10053__,
    new_new_n10054__, new_new_n10055__, new_new_n10056__, new_new_n10057__,
    new_new_n10058__, new_new_n10059__, new_new_n10060__, new_new_n10061__,
    new_new_n10062__, new_new_n10063__, new_new_n10064__, new_new_n10065__,
    new_new_n10066__, new_new_n10067__, new_new_n10068__, new_new_n10069__,
    new_new_n10070__, new_new_n10071__, new_new_n10072__, new_new_n10073__,
    new_new_n10074__, new_new_n10075__, new_new_n10076__, new_new_n10077__,
    new_new_n10078__, new_new_n10079__, new_new_n10080__, new_new_n10081__,
    new_new_n10082__, new_new_n10083__, new_new_n10084__, new_new_n10085__,
    new_new_n10086__, new_new_n10087__, new_new_n10088__, new_new_n10089__,
    new_new_n10090__, new_new_n10091__, new_new_n10092__, new_new_n10093__,
    new_new_n10094__, new_new_n10095__, new_new_n10096__, new_new_n10097__,
    new_new_n10098__, new_new_n10099__, new_new_n10100__, new_new_n10101__,
    new_new_n10102__, new_new_n10103__, new_new_n10104__, new_new_n10105__,
    new_new_n10106__, new_new_n10107__, new_new_n10108__, new_new_n10109__,
    new_new_n10110__, new_new_n10111__, new_new_n10112__, new_new_n10113__,
    new_new_n10114__, new_new_n10115__, new_new_n10116__, new_new_n10117__,
    new_new_n10118__, new_new_n10119__, new_new_n10120__, new_new_n10121__,
    new_new_n10122__, new_new_n10123__, new_new_n10124__, new_new_n10125__,
    new_new_n10126__, new_new_n10127__, new_new_n10128__, new_new_n10129__,
    new_new_n10130__, new_new_n10131__, new_new_n10132__, new_new_n10133__,
    new_new_n10134__, new_new_n10135__, new_new_n10136__, new_new_n10137__,
    new_new_n10138__, new_new_n10139__, new_new_n10140__, new_new_n10141__,
    new_new_n10142__, new_new_n10143__, new_new_n10144__, new_new_n10145__,
    new_new_n10146__, new_new_n10147__, new_new_n10148__, new_new_n10149__,
    new_new_n10150__, new_new_n10151__, new_new_n10152__, new_new_n10153__,
    new_new_n10154__, new_new_n10155__, new_new_n10156__, new_new_n10157__,
    new_new_n10158__, new_new_n10159__, new_new_n10160__, new_new_n10161__,
    new_new_n10162__, new_new_n10163__, new_new_n10164__, new_new_n10165__,
    new_new_n10166__, new_new_n10167__, new_new_n10168__, new_new_n10169__,
    new_new_n10170__, new_new_n10171__, new_new_n10172__, new_new_n10173__,
    new_new_n10174__, new_new_n10175__, new_new_n10176__, new_new_n10177__,
    new_new_n10178__, new_new_n10179__, new_new_n10180__, new_new_n10181__,
    new_new_n10182__, new_new_n10183__, new_new_n10184__, new_new_n10185__,
    new_new_n10186__, new_new_n10187__, new_new_n10188__, new_new_n10189__,
    new_new_n10190__, new_new_n10191__, new_new_n10192__, new_new_n10193__,
    new_new_n10194__, new_new_n10195__, new_new_n10196__, new_new_n10197__,
    new_new_n10198__, new_new_n10199__, new_new_n10200__, new_new_n10201__,
    new_new_n10202__, new_new_n10203__, new_new_n10204__, new_new_n10205__,
    new_new_n10206__, new_new_n10207__, new_new_n10208__, new_new_n10209__,
    new_new_n10210__, new_new_n10211__, new_new_n10212__, new_new_n10213__,
    new_new_n10214__, new_new_n10215__, new_new_n10216__, new_new_n10217__,
    new_new_n10218__, new_new_n10219__, new_new_n10220__, new_new_n10221__,
    new_new_n10222__, new_new_n10223__, new_new_n10224__, new_new_n10225__,
    new_new_n10226__, new_new_n10227__, new_new_n10228__, new_new_n10229__,
    new_new_n10230__, new_new_n10231__, new_new_n10232__, new_new_n10233__,
    new_new_n10234__, new_new_n10235__, new_new_n10236__, new_new_n10237__,
    new_new_n10238__, new_new_n10239__, new_new_n10240__, new_new_n10241__,
    new_new_n10242__, new_new_n10243__, new_new_n10244__, new_new_n10245__,
    new_new_n10246__, new_new_n10247__, new_new_n10248__, new_new_n10249__,
    new_new_n10250__, new_new_n10251__, new_new_n10252__, new_new_n10253__,
    new_new_n10254__, new_new_n10255__, new_new_n10256__, new_new_n10257__,
    new_new_n10258__, new_new_n10259__, new_new_n10260__, new_new_n10261__,
    new_new_n10262__, new_new_n10263__, new_new_n10264__, new_new_n10265__,
    new_new_n10266__, new_new_n10267__, new_new_n10268__, new_new_n10269__,
    new_new_n10270__, new_new_n10271__, new_new_n10272__, new_new_n10273__,
    new_new_n10274__, new_new_n10275__, new_new_n10276__, new_new_n10277__,
    new_new_n10278__, new_new_n10279__, new_new_n10280__, new_new_n10281__,
    new_new_n10282__, new_new_n10283__, new_new_n10284__, new_new_n10285__,
    new_new_n10286__, new_new_n10287__, new_new_n10288__, new_new_n10289__,
    new_new_n10290__, new_new_n10291__, new_new_n10292__, new_new_n10293__,
    new_new_n10294__, new_new_n10295__, new_new_n10296__, new_new_n10297__,
    new_new_n10298__, new_new_n10299__, new_new_n10300__, new_new_n10301__,
    new_new_n10302__, new_new_n10303__, new_new_n10304__, new_new_n10305__,
    new_new_n10306__, new_new_n10307__, new_new_n10308__, new_new_n10309__,
    new_new_n10310__, new_new_n10311__, new_new_n10312__, new_new_n10313__,
    new_new_n10314__, new_new_n10315__, new_new_n10316__, new_new_n10317__,
    new_new_n10318__, new_new_n10319__, new_new_n10320__, new_new_n10321__,
    new_new_n10322__, new_new_n10323__, new_new_n10324__, new_new_n10325__,
    new_new_n10326__, new_new_n10327__, new_new_n10328__, new_new_n10329__,
    new_new_n10330__, new_new_n10331__, new_new_n10332__, new_new_n10333__,
    new_new_n10334__, new_new_n10335__, new_new_n10336__, new_new_n10337__,
    new_new_n10338__, new_new_n10339__, new_new_n10340__, new_new_n10341__,
    new_new_n10342__, new_new_n10343__, new_new_n10344__, new_new_n10345__,
    new_new_n10346__, new_new_n10347__, new_new_n10348__, new_new_n10349__,
    new_new_n10350__, new_new_n10351__, new_new_n10352__, new_new_n10353__,
    new_new_n10354__, new_new_n10355__, new_new_n10356__, new_new_n10357__,
    new_new_n10358__, new_new_n10359__, new_new_n10360__, new_new_n10361__,
    new_new_n10362__, new_new_n10363__, new_new_n10364__, new_new_n10365__,
    new_new_n10366__, new_new_n10367__, new_new_n10368__, new_new_n10369__,
    new_new_n10370__, new_new_n10371__, new_new_n10372__, new_new_n10373__,
    new_new_n10374__, new_new_n10375__, new_new_n10376__, new_new_n10377__,
    new_new_n10378__, new_new_n10379__, new_new_n10380__, new_new_n10381__,
    new_new_n10382__, new_new_n10383__, new_new_n10384__, new_new_n10385__,
    new_new_n10386__, new_new_n10387__, new_new_n10388__, new_new_n10389__,
    new_new_n10390__, new_new_n10391__, new_new_n10392__, new_new_n10393__,
    new_new_n10394__, new_new_n10395__, new_new_n10396__, new_new_n10397__,
    new_new_n10398__, new_new_n10399__, new_new_n10400__, new_new_n10401__,
    new_new_n10402__, new_new_n10403__, new_new_n10404__, new_new_n10405__,
    new_new_n10406__, new_new_n10407__, new_new_n10408__, new_new_n10409__,
    new_new_n10410__, new_new_n10411__, n19409, n19412, n19415, n19418,
    n19421, n19424, n19427, n19430, n19433, n19436, n19439, n19442, n19445,
    n19448, n19451, n19454, n19457, n19460, n19463, n19466, n19469, n19472,
    n19475, n19478, n19481, n19484, n19487, n19490, n19493, n19496, n19499,
    n19502, n19505, n19508, n19511, n19514, n19517, n19520, n19523, n19526,
    n19529, n19532, n19535, n19538, n19541, n19544, n19547, n19550, n19553,
    n19556, n19559, n19562, n19565, n19568, n19571, n19574, n19577, n19580,
    n19583, n19586, n19589, n19592, n19595, n19598, n19601, n19604, n19607,
    n19610, n19613, n19616, n19619, n19622, n19625, n19628, n19631, n19634,
    n19637, n19640, n19643, n19646, n19649, n19652, n19655, n19658, n19661,
    n19664, n19667, n19670, n19673, n19676, n19679, n19682, n19685, n19688,
    n19691, n19694, n19697, n19700, n19703, n19706, n19709, n19712, n19715,
    n19718, n19721, n19724, n19727, n19730, n19733, n19736, n19739, n19742,
    n19745, n19748, n19751, n19754, n19757, n19760, n19763, n19766, n19769,
    n19772, n19775, n19778, n19781, n19784, n19787, n19790, n19793, n19796,
    n19799, n19802, n19805, n19808, n19811, n19814, n19817, n19820, n19823,
    n19826, n19829, n19832, n19835, n19838, n19841, n19844, n19847, n19850,
    n19853, n19856, n19859, n19862, n19865, n19868, n19871, n19874, n19877,
    n19880, n19883, n19886, n19889, n19892, n19895, n19898, n19901, n19904,
    n19907, n19910, n19913, n19916, n19919, n19922, n19925, n19928, n19931,
    n19934, n19937, n19940, n19943, n19946, n19949, n19952, n19955, n19958,
    n19961, n19964, n19967, n19970, n19973, n19976, n19979, n19982, n19985,
    n19988, n19991, n19994, n19997, n20000, n20003, n20006, n20009, n20012,
    n20015, n20018, n20021, n20024, n20027, n20030, n20033, n20036, n20039,
    n20042, n20045, n20048, n20051, n20054, n20057, n20060, n20063, n20066,
    n20069, n20072, n20075, n20078, n20081, n20084, n20087, n20090, n20093,
    n20096, n20099, n20102, n20105, n20108, n20111, n20114, n20117, n20120,
    n20123, n20126, n20129, n20132, n20135, n20138, n20141, n20144, n20147,
    n20150, n20153, n20156, n20159, n20162, n20165, n20168, n20171, n20174,
    n20177, n20180, n20183, n20186, n20189, n20192, n20195, n20198, n20201,
    n20204, n20207, n20210, n20213, n20216, n20219, n20222, n20225, n20228,
    n20231, n20234, n20237, n20240, n20243, n20246, n20249, n20252, n20255,
    n20258, n20261, n20264, n20267, n20270, n20273, n20276, n20279, n20282,
    n20285, n20288, n20291, n20294, n20297, n20300, n20303, n20306, n20309,
    n20312, n20315, n20318, n20321, n20324, n20327, n20330, n20333, n20336,
    n20339, n20342, n20345, n20348, n20351, n20354, n20357, n20360, n20363,
    n20366, n20369, n20372, n20375, n20378, n20381, n20384, n20387, n20390,
    n20393, n20396, n20399, n20402, n20405, n20408, n20411, n20414, n20417,
    n20420, n20423, n20426, n20429, n20432, n20435, n20438, n20441, n20444,
    n20447, n20450, n20453, n20456, n20459, n20462, n20465, n20468, n20471,
    n20474, n20477, n20480, n20483, n20486, n20489, n20492, n20495, n20498,
    n20501, n20504, n20507, n20510, n20513, n20516, n20519, n20522;
  buf1  g0000(.din(G1), .dout(new_new_n809__));
  not1  g0001(.din(G1), .dout(new_new_n810__));
  buf1  g0002(.din(G2), .dout(new_new_n811__));
  not1  g0003(.din(G2), .dout(new_new_n812__));
  buf1  g0004(.din(G3), .dout(new_new_n813__));
  not1  g0005(.din(G3), .dout(new_new_n814__));
  buf1  g0006(.din(G4), .dout(new_new_n815__));
  not1  g0007(.din(G4), .dout(new_new_n816__));
  buf1  g0008(.din(G5), .dout(new_new_n817__));
  not1  g0009(.din(G5), .dout(new_new_n818__));
  buf1  g0010(.din(G6), .dout(new_new_n819__));
  not1  g0011(.din(G6), .dout(new_new_n820__));
  buf1  g0012(.din(G7), .dout(new_new_n821__));
  not1  g0013(.din(G7), .dout(new_new_n822__));
  buf1  g0014(.din(G8), .dout(new_new_n823__));
  not1  g0015(.din(G8), .dout(new_new_n824__));
  buf1  g0016(.din(G9), .dout(new_new_n825__));
  not1  g0017(.din(G9), .dout(new_new_n826__));
  buf1  g0018(.din(G10), .dout(new_new_n827__));
  not1  g0019(.din(G10), .dout(new_new_n828__));
  buf1  g0020(.din(G11), .dout(new_new_n829__));
  not1  g0021(.din(G11), .dout(new_new_n830__));
  buf1  g0022(.din(G12), .dout(new_new_n831__));
  not1  g0023(.din(G12), .dout(new_new_n832__));
  buf1  g0024(.din(G13), .dout(new_new_n833__));
  not1  g0025(.din(G13), .dout(new_new_n834__));
  buf1  g0026(.din(G14), .dout(new_new_n835__));
  not1  g0027(.din(G14), .dout(new_new_n836__));
  buf1  g0028(.din(G15), .dout(new_new_n837__));
  not1  g0029(.din(G15), .dout(new_new_n838__));
  buf1  g0030(.din(G16), .dout(new_new_n839__));
  not1  g0031(.din(G16), .dout(new_new_n840__));
  buf1  g0032(.din(G17), .dout(new_new_n841__));
  not1  g0033(.din(G17), .dout(new_new_n842__));
  buf1  g0034(.din(G18), .dout(new_new_n843__));
  not1  g0035(.din(G18), .dout(new_new_n844__));
  buf1  g0036(.din(G19), .dout(new_new_n845__));
  not1  g0037(.din(G19), .dout(new_new_n846__));
  buf1  g0038(.din(G20), .dout(new_new_n847__));
  not1  g0039(.din(G20), .dout(new_new_n848__));
  buf1  g0040(.din(G21), .dout(new_new_n849__));
  buf1  g0041(.din(G22), .dout(new_new_n851__));
  buf1  g0042(.din(G23), .dout(new_new_n853__));
  buf1  g0043(.din(G24), .dout(new_new_n855__));
  buf1  g0044(.din(G25), .dout(new_new_n857__));
  buf1  g0045(.din(G26), .dout(new_new_n859__));
  buf1  g0046(.din(G27), .dout(new_new_n861__));
  buf1  g0047(.din(G28), .dout(new_new_n863__));
  buf1  g0048(.din(G29), .dout(new_new_n865__));
  buf1  g0049(.din(G30), .dout(new_new_n867__));
  buf1  g0050(.din(G31), .dout(new_new_n869__));
  buf1  g0051(.din(G32), .dout(new_new_n871__));
  buf1  g0052(.din(n2491_lo), .dout(new_new_n873__));
  buf1  g0053(.din(n2575_lo), .dout(new_new_n875__));
  not1  g0054(.din(n2575_lo), .dout(new_new_n876__));
  buf1  g0055(.din(n2587_lo), .dout(new_new_n877__));
  not1  g0056(.din(n2587_lo), .dout(new_new_n878__));
  buf1  g0057(.din(n2599_lo), .dout(new_new_n879__));
  not1  g0058(.din(n2599_lo), .dout(new_new_n880__));
  buf1  g0059(.din(n2611_lo), .dout(new_new_n881__));
  not1  g0060(.din(n2611_lo), .dout(new_new_n882__));
  buf1  g0061(.din(n2623_lo), .dout(new_new_n883__));
  not1  g0062(.din(n2623_lo), .dout(new_new_n884__));
  buf1  g0063(.din(n2635_lo), .dout(new_new_n885__));
  not1  g0064(.din(n2635_lo), .dout(new_new_n886__));
  buf1  g0065(.din(n2647_lo), .dout(new_new_n887__));
  not1  g0066(.din(n2647_lo), .dout(new_new_n888__));
  buf1  g0067(.din(n2659_lo), .dout(new_new_n889__));
  not1  g0068(.din(n2659_lo), .dout(new_new_n890__));
  buf1  g0069(.din(n2671_lo), .dout(new_new_n891__));
  not1  g0070(.din(n2671_lo), .dout(new_new_n892__));
  buf1  g0071(.din(n2683_lo), .dout(new_new_n893__));
  buf1  g0072(.din(n2734_lo), .dout(new_new_n895__));
  not1  g0073(.din(n2734_lo), .dout(new_new_n896__));
  buf1  g0074(.din(n2746_lo), .dout(new_new_n897__));
  not1  g0075(.din(n2746_lo), .dout(new_new_n898__));
  buf1  g0076(.din(n2758_lo), .dout(new_new_n899__));
  not1  g0077(.din(n2758_lo), .dout(new_new_n900__));
  buf1  g0078(.din(n2770_lo), .dout(new_new_n901__));
  not1  g0079(.din(n2770_lo), .dout(new_new_n902__));
  buf1  g0080(.din(n2782_lo), .dout(new_new_n903__));
  buf1  g0081(.din(n2785_lo), .dout(new_new_n905__));
  not1  g0082(.din(n2785_lo), .dout(new_new_n906__));
  buf1  g0083(.din(n2794_lo), .dout(new_new_n907__));
  buf1  g0084(.din(n2797_lo), .dout(new_new_n909__));
  not1  g0085(.din(n2797_lo), .dout(new_new_n910__));
  buf1  g0086(.din(n2806_lo), .dout(new_new_n911__));
  buf1  g0087(.din(n2809_lo), .dout(new_new_n913__));
  not1  g0088(.din(n2809_lo), .dout(new_new_n914__));
  buf1  g0089(.din(n2818_lo), .dout(new_new_n915__));
  buf1  g0090(.din(n2821_lo), .dout(new_new_n917__));
  not1  g0091(.din(n2821_lo), .dout(new_new_n918__));
  buf1  g0092(.din(n2830_lo), .dout(new_new_n919__));
  buf1  g0093(.din(n2833_lo), .dout(new_new_n921__));
  buf1  g0094(.din(n2836_lo), .dout(new_new_n923__));
  not1  g0095(.din(n2836_lo), .dout(new_new_n924__));
  buf1  g0096(.din(n2839_lo), .dout(new_new_n925__));
  not1  g0097(.din(n2839_lo), .dout(new_new_n926__));
  buf1  g0098(.din(n2842_lo), .dout(new_new_n927__));
  buf1  g0099(.din(n2845_lo), .dout(new_new_n929__));
  buf1  g0100(.din(n2848_lo), .dout(new_new_n931__));
  not1  g0101(.din(n2848_lo), .dout(new_new_n932__));
  buf1  g0102(.din(n2851_lo), .dout(new_new_n933__));
  not1  g0103(.din(n2851_lo), .dout(new_new_n934__));
  buf1  g0104(.din(n2854_lo), .dout(new_new_n935__));
  buf1  g0105(.din(n2857_lo), .dout(new_new_n937__));
  buf1  g0106(.din(n2860_lo), .dout(new_new_n939__));
  not1  g0107(.din(n2860_lo), .dout(new_new_n940__));
  buf1  g0108(.din(n2863_lo), .dout(new_new_n941__));
  not1  g0109(.din(n2863_lo), .dout(new_new_n942__));
  buf1  g0110(.din(n4871_o2), .dout(new_new_n943__));
  not1  g0111(.din(n4893_o2), .dout(new_new_n946__));
  buf1  g0112(.din(n4938_o2), .dout(new_new_n947__));
  buf1  g0113(.din(n5056_o2), .dout(new_new_n949__));
  not1  g0114(.din(n5100_o2), .dout(new_new_n952__));
  buf1  g0115(.din(n5122_o2), .dout(new_new_n953__));
  buf1  g0116(.din(n5254_o2), .dout(new_new_n955__));
  not1  g0117(.din(n5276_o2), .dout(new_new_n958__));
  buf1  g0118(.din(n5316_o2), .dout(new_new_n959__));
  buf1  g0119(.din(n5434_o2), .dout(new_new_n961__));
  not1  g0120(.din(n5473_o2), .dout(new_new_n964__));
  buf1  g0121(.din(n5494_o2), .dout(new_new_n965__));
  buf1  g0122(.din(n5620_o2), .dout(new_new_n967__));
  not1  g0123(.din(n5643_o2), .dout(new_new_n970__));
  buf1  g0124(.din(n5682_o2), .dout(new_new_n971__));
  buf1  g0125(.din(n5798_o2), .dout(new_new_n973__));
  not1  g0126(.din(n5839_o2), .dout(new_new_n976__));
  buf1  g0127(.din(n5867_o2), .dout(new_new_n977__));
  buf1  g0128(.din(n6052_o2), .dout(new_new_n979__));
  not1  g0129(.din(n6087_o2), .dout(new_new_n982__));
  buf1  g0130(.din(n6153_o2), .dout(new_new_n983__));
  buf1  g0131(.din(n6408_o2), .dout(new_new_n985__));
  not1  g0132(.din(n6454_o2), .dout(new_new_n988__));
  buf1  g0133(.din(n6509_o2), .dout(new_new_n989__));
  buf1  g0134(.din(n6775_o2), .dout(new_new_n991__));
  not1  g0135(.din(n6818_o2), .dout(new_new_n994__));
  buf1  g0136(.din(n6892_o2), .dout(new_new_n995__));
  buf1  g0137(.din(n5779_o2), .dout(new_new_n997__));
  not1  g0138(.din(n5779_o2), .dout(new_new_n998__));
  buf1  g0139(.din(n5780_o2), .dout(new_new_n999__));
  buf1  g0140(.din(n7156_o2), .dout(new_new_n1001__));
  buf1  g0141(.din(n5792_o2), .dout(new_new_n1003__));
  not1  g0142(.din(n5792_o2), .dout(new_new_n1004__));
  not1  g0143(.din(n7205_o2), .dout(new_new_n1006__));
  buf1  g0144(.din(n5842_o2), .dout(new_new_n1007__));
  not1  g0145(.din(n5842_o2), .dout(new_new_n1008__));
  buf1  g0146(.din(n5863_o2), .dout(new_new_n1009__));
  not1  g0147(.din(n5863_o2), .dout(new_new_n1010__));
  buf1  g0148(.din(n7263_o2), .dout(new_new_n1011__));
  buf1  g0149(.din(n5881_o2), .dout(new_new_n1013__));
  not1  g0150(.din(n5881_o2), .dout(new_new_n1014__));
  buf1  g0151(.din(n5930_o2), .dout(new_new_n1015__));
  not1  g0152(.din(n5930_o2), .dout(new_new_n1016__));
  buf1  g0153(.din(n5959_o2), .dout(new_new_n1017__));
  not1  g0154(.din(n5959_o2), .dout(new_new_n1018__));
  buf1  g0155(.din(n5981_o2), .dout(new_new_n1019__));
  not1  g0156(.din(n5981_o2), .dout(new_new_n1020__));
  buf1  g0157(.din(n6042_o2), .dout(new_new_n1021__));
  not1  g0158(.din(n6042_o2), .dout(new_new_n1022__));
  buf1  g0159(.din(n6075_o2), .dout(new_new_n1023__));
  not1  g0160(.din(n6075_o2), .dout(new_new_n1024__));
  buf1  g0161(.din(n6103_o2), .dout(new_new_n1025__));
  not1  g0162(.din(n6103_o2), .dout(new_new_n1026__));
  buf1  g0163(.din(n7610_o2), .dout(new_new_n1027__));
  buf1  g0164(.din(n6169_o2), .dout(new_new_n1029__));
  not1  g0165(.din(n6169_o2), .dout(new_new_n1030__));
  not1  g0166(.din(n7665_o2), .dout(new_new_n1032__));
  buf1  g0167(.din(n6205_o2), .dout(new_new_n1033__));
  not1  g0168(.din(n6205_o2), .dout(new_new_n1034__));
  buf1  g0169(.din(n6239_o2), .dout(new_new_n1035__));
  not1  g0170(.din(n6239_o2), .dout(new_new_n1036__));
  buf1  g0171(.din(n7788_o2), .dout(new_new_n1037__));
  buf1  g0172(.din(n6309_o2), .dout(new_new_n1039__));
  not1  g0173(.din(n6309_o2), .dout(new_new_n1040__));
  buf1  g0174(.din(n6461_o2), .dout(new_new_n1041__));
  not1  g0175(.din(n6461_o2), .dout(new_new_n1042__));
  buf1  g0176(.din(n6476_o2), .dout(new_new_n1043__));
  buf1  g0177(.din(n325_inv), .dout(new_new_n1045__));
  buf1  g0178(.din(n6545_o2), .dout(new_new_n1047__));
  buf1  g0179(.din(G578_o2), .dout(new_new_n1049__));
  not1  g0180(.din(G5106_o2), .dout(new_new_n1052__));
  buf1  g0181(.din(n6713_o2), .dout(new_new_n1053__));
  buf1  g0182(.din(G5164_o2), .dout(new_new_n1055__));
  buf1  g0183(.din(n343_inv), .dout(new_new_n1057__));
  buf1  g0184(.din(n6810_o2), .dout(new_new_n1059__));
  buf1  g0185(.din(n6973_o2), .dout(new_new_n1061__));
  buf1  g0186(.din(n352_inv), .dout(new_new_n1063__));
  buf1  g0187(.din(n7053_o2), .dout(new_new_n1065__));
  buf1  g0188(.din(G581_o2), .dout(new_new_n1067__));
  not1  g0189(.din(G5467_o2), .dout(new_new_n1070__));
  buf1  g0190(.din(n7231_o2), .dout(new_new_n1071__));
  buf1  g0191(.din(G5527_o2), .dout(new_new_n1073__));
  buf1  g0192(.din(n370_inv), .dout(new_new_n1075__));
  buf1  g0193(.din(n7304_o2), .dout(new_new_n1077__));
  buf1  g0194(.din(n7530_o2), .dout(new_new_n1079__));
  buf1  g0195(.din(n379_inv), .dout(new_new_n1081__));
  buf1  g0196(.din(n7653_o2), .dout(new_new_n1083__));
  buf1  g0197(.din(G584_o2), .dout(new_new_n1085__));
  not1  g0198(.din(G5820_o2), .dout(new_new_n1088__));
  buf1  g0199(.din(n7148_o2), .dout(new_new_n1089__));
  not1  g0200(.din(n7148_o2), .dout(new_new_n1090__));
  buf1  g0201(.din(n7149_o2), .dout(new_new_n1091__));
  buf1  g0202(.din(n7224_o2), .dout(new_new_n1093__));
  not1  g0203(.din(n7224_o2), .dout(new_new_n1094__));
  buf1  g0204(.din(n7916_o2), .dout(new_new_n1095__));
  buf1  g0205(.din(G5868_o2), .dout(new_new_n1097__));
  buf1  g0206(.din(n406_inv), .dout(new_new_n1099__));
  buf1  g0207(.din(n7280_o2), .dout(new_new_n1101__));
  not1  g0208(.din(n7280_o2), .dout(new_new_n1102__));
  buf1  g0209(.din(n7313_o2), .dout(new_new_n1103__));
  not1  g0210(.din(n7313_o2), .dout(new_new_n1104__));
  buf1  g0211(.din(n8056_o2), .dout(new_new_n1105__));
  buf1  g0212(.din(n7323_o2), .dout(new_new_n1107__));
  not1  g0213(.din(n7323_o2), .dout(new_new_n1108__));
  buf1  g0214(.din(n7398_o2), .dout(new_new_n1109__));
  not1  g0215(.din(n7398_o2), .dout(new_new_n1110__));
  buf1  g0216(.din(n7459_o2), .dout(new_new_n1111__));
  not1  g0217(.din(n7459_o2), .dout(new_new_n1112__));
  buf1  g0218(.din(n7501_o2), .dout(new_new_n1113__));
  not1  g0219(.din(n7501_o2), .dout(new_new_n1114__));
  buf1  g0220(.din(n7518_o2), .dout(new_new_n1115__));
  not1  g0221(.din(n7518_o2), .dout(new_new_n1116__));
  buf1  g0222(.din(G563_o2), .dout(new_new_n1117__));
  buf1  g0223(.din(n7606_o2), .dout(new_new_n1119__));
  not1  g0224(.din(n7606_o2), .dout(new_new_n1120__));
  buf1  g0225(.din(n439_inv), .dout(new_new_n1121__));
  buf1  g0226(.din(n7675_o2), .dout(new_new_n1123__));
  not1  g0227(.din(n7675_o2), .dout(new_new_n1124__));
  buf1  g0228(.din(G3410_o2), .dout(new_new_n1125__));
  buf1  g0229(.din(n7722_o2), .dout(new_new_n1127__));
  not1  g0230(.din(n7722_o2), .dout(new_new_n1128__));
  buf1  g0231(.din(n7747_o2), .dout(new_new_n1129__));
  not1  g0232(.din(n7747_o2), .dout(new_new_n1130__));
  buf1  g0233(.din(n7835_o2), .dout(new_new_n1131__));
  not1  g0234(.din(n7835_o2), .dout(new_new_n1132__));
  buf1  g0235(.din(G587_o2), .dout(new_new_n1133__));
  not1  g0236(.din(G6046_o2), .dout(new_new_n1136__));
  buf1  g0237(.din(n7909_o2), .dout(new_new_n1137__));
  not1  g0238(.din(n7909_o2), .dout(new_new_n1138__));
  buf1  g0239(.din(G566_o2), .dout(new_new_n1139__));
  buf1  g0240(.din(G6070_o2), .dout(new_new_n1141__));
  buf1  g0241(.din(n472_inv), .dout(new_new_n1143__));
  buf1  g0242(.din(n8086_o2), .dout(new_new_n1145__));
  not1  g0243(.din(n8086_o2), .dout(new_new_n1146__));
  buf1  g0244(.din(n8093_o2), .dout(new_new_n1147__));
  buf1  g0245(.din(G3752_o2), .dout(new_new_n1149__));
  buf1  g0246(.din(n484_inv), .dout(new_new_n1151__));
  buf1  g0247(.din(n8199_o2), .dout(new_new_n1153__));
  buf1  g0248(.din(n2800_lo_buf_o2), .dout(new_new_n1155__));
  not1  g0249(.din(n2800_lo_buf_o2), .dout(new_new_n1156__));
  buf1  g0250(.din(G548_o2), .dout(new_new_n1157__));
  buf1  g0251(.din(n496_inv), .dout(new_new_n1159__));
  buf1  g0252(.din(G569_o2), .dout(new_new_n1161__));
  buf1  g0253(.din(G1761_o2), .dout(new_new_n1163__));
  buf1  g0254(.din(n505_inv), .dout(new_new_n1165__));
  buf1  g0255(.din(G4101_o2), .dout(new_new_n1167__));
  buf1  g0256(.din(G551_o2), .dout(new_new_n1169__));
  buf1  g0257(.din(n514_inv), .dout(new_new_n1171__));
  buf1  g0258(.din(G4743_o2), .dout(new_new_n1173__));
  not1  g0259(.din(G4743_o2), .dout(new_new_n1174__));
  buf1  g0260(.din(G5271_o2), .dout(new_new_n1175__));
  not1  g0261(.din(G5271_o2), .dout(new_new_n1176__));
  buf1  g0262(.din(G5790_o2), .dout(new_new_n1177__));
  not1  g0263(.din(G5790_o2), .dout(new_new_n1178__));
  not1  g0264(.din(G6122_o2), .dout(new_new_n1180__));
  buf1  g0265(.din(G2082_o2), .dout(new_new_n1181__));
  buf1  g0266(.din(n2812_lo_buf_o2), .dout(new_new_n1183__));
  not1  g0267(.din(n2812_lo_buf_o2), .dout(new_new_n1184__));
  buf1  g0268(.din(n2668_lo_buf_o2), .dout(new_new_n1185__));
  not1  g0269(.din(n2668_lo_buf_o2), .dout(new_new_n1186__));
  buf1  g0270(.din(n2680_lo_buf_o2), .dout(new_new_n1187__));
  buf1  g0271(.din(G572_o2), .dout(new_new_n1189__));
  buf1  g0272(.din(G6125_o2), .dout(new_new_n1191__));
  buf1  g0273(.din(n547_inv), .dout(new_new_n1193__));
  buf1  g0274(.din(n2656_lo_buf_o2), .dout(new_new_n1195__));
  not1  g0275(.din(n2656_lo_buf_o2), .dout(new_new_n1196__));
  buf1  g0276(.din(G554_o2), .dout(new_new_n1197__));
  buf1  g0277(.din(G4452_o2), .dout(new_new_n1199__));
  buf1  g0278(.din(n559_inv), .dout(new_new_n1201__));
  buf1  g0279(.din(n2644_lo_buf_o2), .dout(new_new_n1203__));
  not1  g0280(.din(n2644_lo_buf_o2), .dout(new_new_n1204__));
  buf1  g0281(.din(G2410_o2), .dout(new_new_n1205__));
  buf1  g0282(.din(n2632_lo_buf_o2), .dout(new_new_n1207__));
  not1  g0283(.din(n2632_lo_buf_o2), .dout(new_new_n1208__));
  buf1  g0284(.din(n2620_lo_buf_o2), .dout(new_new_n1209__));
  not1  g0285(.din(n2620_lo_buf_o2), .dout(new_new_n1210__));
  buf1  g0286(.din(G6131_o2), .dout(new_new_n1211__));
  buf1  g0287(.din(G4693_o2), .dout(new_new_n1213__));
  not1  g0288(.din(G4693_o2), .dout(new_new_n1214__));
  buf1  g0289(.din(G5209_o2), .dout(new_new_n1215__));
  not1  g0290(.din(G5209_o2), .dout(new_new_n1216__));
  buf1  g0291(.din(G5741_o2), .dout(new_new_n1217__));
  not1  g0292(.din(G5741_o2), .dout(new_new_n1218__));
  buf1  g0293(.din(G6082_o2), .dout(new_new_n1219__));
  not1  g0294(.din(G6082_o2), .dout(new_new_n1220__));
  not1  g0295(.din(G6119_o2), .dout(new_new_n1222__));
  buf1  g0296(.din(n2608_lo_buf_o2), .dout(new_new_n1223__));
  not1  g0297(.din(n2608_lo_buf_o2), .dout(new_new_n1224__));
  buf1  g0298(.din(n2596_lo_buf_o2), .dout(new_new_n1225__));
  not1  g0299(.din(n2596_lo_buf_o2), .dout(new_new_n1226__));
  buf1  g0300(.din(n2584_lo_buf_o2), .dout(new_new_n1227__));
  not1  g0301(.din(n2584_lo_buf_o2), .dout(new_new_n1228__));
  buf1  g0302(.din(n2572_lo_buf_o2), .dout(new_new_n1229__));
  not1  g0303(.din(n2572_lo_buf_o2), .dout(new_new_n1230__));
  buf1  g0304(.din(n2704_lo_buf_o2), .dout(new_new_n1231__));
  not1  g0305(.din(n2704_lo_buf_o2), .dout(new_new_n1232__));
  buf1  g0306(.din(G557_o2), .dout(new_new_n1233__));
  buf1  g0307(.din(G5936_o2), .dout(new_new_n1235__));
  not1  g0308(.din(G5936_o2), .dout(new_new_n1236__));
  buf1  g0309(.din(G5442_o2), .dout(new_new_n1237__));
  not1  g0310(.din(G5442_o2), .dout(new_new_n1238__));
  buf1  g0311(.din(G4926_o2), .dout(new_new_n1239__));
  not1  g0312(.din(G4926_o2), .dout(new_new_n1240__));
  buf1  g0313(.din(G6134_o2), .dout(new_new_n1241__));
  buf1  g0314(.din(G3929_o2), .dout(new_new_n1243__));
  not1  g0315(.din(G3929_o2), .dout(new_new_n1244__));
  buf1  g0316(.din(G4425_o2), .dout(new_new_n1245__));
  not1  g0317(.din(G4425_o2), .dout(new_new_n1246__));
  buf1  g0318(.din(G4947_o2), .dout(new_new_n1247__));
  not1  g0319(.din(G4947_o2), .dout(new_new_n1248__));
  buf1  g0320(.din(n2764_lo_buf_o2), .dout(new_new_n1249__));
  not1  g0321(.din(n2764_lo_buf_o2), .dout(new_new_n1250__));
  buf1  g0322(.din(n634_inv), .dout(new_new_n1251__));
  buf1  g0323(.din(n2560_lo_buf_o2), .dout(new_new_n1253__));
  not1  g0324(.din(n2560_lo_buf_o2), .dout(new_new_n1254__));
  buf1  g0325(.din(n2824_lo_buf_o2), .dout(new_new_n1255__));
  not1  g0326(.din(n2824_lo_buf_o2), .dout(new_new_n1256__));
  buf1  g0327(.din(G575_o2), .dout(new_new_n1257__));
  buf1  g0328(.din(G2740_o2), .dout(new_new_n1259__));
  buf1  g0329(.din(n649_inv), .dout(new_new_n1261__));
  buf1  g0330(.din(n2548_lo_buf_o2), .dout(new_new_n1263__));
  not1  g0331(.din(n2548_lo_buf_o2), .dout(new_new_n1264__));
  buf1  g0332(.din(n2536_lo_buf_o2), .dout(new_new_n1265__));
  not1  g0333(.din(n2536_lo_buf_o2), .dout(new_new_n1266__));
  buf1  g0334(.din(n2524_lo_buf_o2), .dout(new_new_n1267__));
  not1  g0335(.din(n2524_lo_buf_o2), .dout(new_new_n1268__));
  buf1  g0336(.din(G875_o2), .dout(new_new_n1269__));
  not1  g0337(.din(G875_o2), .dout(new_new_n1270__));
  buf1  g0338(.din(G1064_o2), .dout(new_new_n1271__));
  not1  g0339(.din(G1064_o2), .dout(new_new_n1272__));
  buf1  g0340(.din(G1253_o2), .dout(new_new_n1273__));
  not1  g0341(.din(G1253_o2), .dout(new_new_n1274__));
  buf1  g0342(.din(G6140_o2), .dout(new_new_n1275__));
  buf1  g0343(.din(G5151_o2), .dout(new_new_n1277__));
  not1  g0344(.din(G5151_o2), .dout(new_new_n1278__));
  buf1  g0345(.din(G5686_o2), .dout(new_new_n1279__));
  not1  g0346(.din(G5686_o2), .dout(new_new_n1280__));
  buf1  g0347(.din(G6061_o2), .dout(new_new_n1281__));
  not1  g0348(.din(G6061_o2), .dout(new_new_n1282__));
  buf1  g0349(.din(G4803_o2), .dout(new_new_n1283__));
  not1  g0350(.din(G4803_o2), .dout(new_new_n1284__));
  buf1  g0351(.din(G5332_o2), .dout(new_new_n1285__));
  not1  g0352(.din(G5332_o2), .dout(new_new_n1286__));
  buf1  g0353(.din(G5844_o2), .dout(new_new_n1287__));
  not1  g0354(.din(G5844_o2), .dout(new_new_n1288__));
  not1  g0355(.din(G6114_o2), .dout(new_new_n1290__));
  buf1  g0356(.din(G4806_o2), .dout(new_new_n1291__));
  buf1  g0357(.din(G3881_o2), .dout(new_new_n1293__));
  not1  g0358(.din(G3881_o2), .dout(new_new_n1294__));
  buf1  g0359(.din(G4370_o2), .dout(new_new_n1295__));
  not1  g0360(.din(G4370_o2), .dout(new_new_n1296__));
  buf1  g0361(.din(G4896_o2), .dout(new_new_n1297__));
  not1  g0362(.din(G4896_o2), .dout(new_new_n1298__));
  buf1  g0363(.din(G5001_o2), .dout(new_new_n1299__));
  not1  g0364(.din(G5001_o2), .dout(new_new_n1300__));
  buf1  g0365(.din(G3121_o2), .dout(new_new_n1301__));
  not1  g0366(.din(G3121_o2), .dout(new_new_n1302__));
  buf1  g0367(.din(n2512_lo_buf_o2), .dout(new_new_n1303__));
  not1  g0368(.din(n2512_lo_buf_o2), .dout(new_new_n1304__));
  buf1  g0369(.din(G4085_o2), .dout(new_new_n1305__));
  not1  g0370(.din(G4085_o2), .dout(new_new_n1306__));
  buf1  g0371(.din(G4605_o2), .dout(new_new_n1307__));
  not1  g0372(.din(G4605_o2), .dout(new_new_n1308__));
  buf1  g0373(.din(G5118_o2), .dout(new_new_n1309__));
  not1  g0374(.din(G5118_o2), .dout(new_new_n1310__));
  buf1  g0375(.din(G4997_o2), .dout(new_new_n1311__));
  not1  g0376(.din(G4997_o2), .dout(new_new_n1312__));
  buf1  g0377(.din(n2500_lo_buf_o2), .dout(new_new_n1313__));
  not1  g0378(.din(n2500_lo_buf_o2), .dout(new_new_n1314__));
  buf1  g0379(.din(n2716_lo_buf_o2), .dout(new_new_n1315__));
  not1  g0380(.din(n2716_lo_buf_o2), .dout(new_new_n1316__));
  buf1  g0381(.din(G560_o2), .dout(new_new_n1317__));
  buf1  g0382(.din(G1895_o2), .dout(new_new_n1319__));
  not1  g0383(.din(G1895_o2), .dout(new_new_n1320__));
  buf1  g0384(.din(G3064_o2), .dout(new_new_n1321__));
  not1  g0385(.din(G3064_o2), .dout(new_new_n1322__));
  buf1  g0386(.din(G3269_o2), .dout(new_new_n1323__));
  not1  g0387(.din(G3269_o2), .dout(new_new_n1324__));
  buf1  g0388(.din(G3569_o2), .dout(new_new_n1325__));
  not1  g0389(.din(G3569_o2), .dout(new_new_n1326__));
  buf1  g0390(.din(n748_inv), .dout(new_new_n1327__));
  buf1  g0391(.din(G1196_o2), .dout(new_new_n1329__));
  not1  g0392(.din(G1196_o2), .dout(new_new_n1330__));
  buf1  g0393(.din(G1007_o2), .dout(new_new_n1331__));
  not1  g0394(.din(G1007_o2), .dout(new_new_n1332__));
  buf1  g0395(.din(G818_o2), .dout(new_new_n1333__));
  not1  g0396(.din(G818_o2), .dout(new_new_n1334__));
  buf1  g0397(.din(G674_o2), .dout(new_new_n1335__));
  not1  g0398(.din(G674_o2), .dout(new_new_n1336__));
  buf1  g0399(.din(G5041_o2), .dout(new_new_n1337__));
  not1  g0400(.din(G5041_o2), .dout(new_new_n1338__));
  buf1  g0401(.din(G5562_o2), .dout(new_new_n1339__));
  not1  g0402(.din(G5562_o2), .dout(new_new_n1340__));
  buf1  g0403(.din(G6005_o2), .dout(new_new_n1341__));
  not1  g0404(.din(G6005_o2), .dout(new_new_n1342__));
  buf1  g0405(.din(G5214_o2), .dout(new_new_n1343__));
  not1  g0406(.din(G5214_o2), .dout(new_new_n1344__));
  buf1  g0407(.din(G5746_o2), .dout(new_new_n1345__));
  not1  g0408(.din(G5746_o2), .dout(new_new_n1346__));
  buf1  g0409(.din(G6087_o2), .dout(new_new_n1347__));
  not1  g0410(.din(G6087_o2), .dout(new_new_n1348__));
  buf1  g0411(.din(G6086_o2), .dout(new_new_n1349__));
  not1  g0412(.din(G6086_o2), .dout(new_new_n1350__));
  buf1  g0413(.din(G5745_o2), .dout(new_new_n1351__));
  not1  g0414(.din(G5745_o2), .dout(new_new_n1352__));
  buf1  g0415(.din(G5213_o2), .dout(new_new_n1353__));
  not1  g0416(.din(G5213_o2), .dout(new_new_n1354__));
  buf1  g0417(.din(G5893_o2), .dout(new_new_n1355__));
  not1  g0418(.din(G5893_o2), .dout(new_new_n1356__));
  buf1  g0419(.din(G5391_o2), .dout(new_new_n1357__));
  not1  g0420(.din(G5391_o2), .dout(new_new_n1358__));
  buf1  g0421(.din(G4864_o2), .dout(new_new_n1359__));
  not1  g0422(.din(G4864_o2), .dout(new_new_n1360__));
  buf1  g0423(.din(G6143_o2), .dout(new_new_n1361__));
  not1  g0424(.din(G6143_o2), .dout(new_new_n1362__));
  buf1  g0425(.din(G6008_o2), .dout(new_new_n1363__));
  not1  g0426(.din(G6008_o2), .dout(new_new_n1364__));
  buf1  g0427(.din(G5565_o2), .dout(new_new_n1365__));
  not1  g0428(.din(G5565_o2), .dout(new_new_n1366__));
  buf1  g0429(.din(G5044_o2), .dout(new_new_n1367__));
  not1  g0430(.din(G5044_o2), .dout(new_new_n1368__));
  buf1  g0431(.din(G3813_o2), .dout(new_new_n1369__));
  not1  g0432(.din(G3813_o2), .dout(new_new_n1370__));
  buf1  g0433(.din(G4325_o2), .dout(new_new_n1371__));
  not1  g0434(.din(G4325_o2), .dout(new_new_n1372__));
  buf1  g0435(.din(G4834_o2), .dout(new_new_n1373__));
  not1  g0436(.din(G4834_o2), .dout(new_new_n1374__));
  buf1  g0437(.din(G4993_o2), .dout(new_new_n1375__));
  not1  g0438(.din(G4993_o2), .dout(new_new_n1376__));
  buf1  g0439(.din(G3989_o2), .dout(new_new_n1377__));
  not1  g0440(.din(G3989_o2), .dout(new_new_n1378__));
  buf1  g0441(.din(G4490_o2), .dout(new_new_n1379__));
  not1  g0442(.din(G4490_o2), .dout(new_new_n1380__));
  buf1  g0443(.din(G5011_o2), .dout(new_new_n1381__));
  not1  g0444(.din(G5011_o2), .dout(new_new_n1382__));
  buf1  g0445(.din(G5112_o2), .dout(new_new_n1383__));
  not1  g0446(.din(G5112_o2), .dout(new_new_n1384__));
  buf1  g0447(.din(n2776_lo_buf_o2), .dout(new_new_n1385__));
  not1  g0448(.din(n2776_lo_buf_o2), .dout(new_new_n1386__));
  buf1  g0449(.din(G3298_o2), .dout(new_new_n1387__));
  not1  g0450(.din(G3298_o2), .dout(new_new_n1388__));
  buf1  g0451(.din(G3073_o2), .dout(new_new_n1389__));
  buf1  g0452(.din(G3265_o2), .dout(new_new_n1391__));
  not1  g0453(.din(G3265_o2), .dout(new_new_n1392__));
  buf1  g0454(.din(G3624_o2), .dout(new_new_n1393__));
  not1  g0455(.din(G3624_o2), .dout(new_new_n1394__));
  buf1  g0456(.din(G1642_o2), .dout(new_new_n1395__));
  not1  g0457(.din(G1642_o2), .dout(new_new_n1396__));
  buf1  g0458(.din(G1980_o2), .dout(new_new_n1397__));
  not1  g0459(.din(G1980_o2), .dout(new_new_n1398__));
  buf1  g0460(.din(n2488_lo_buf_o2), .dout(new_new_n1399__));
  not1  g0461(.din(n2488_lo_buf_o2), .dout(new_new_n1400__));
  buf1  g0462(.din(G626_o2), .dout(new_new_n1401__));
  not1  g0463(.din(G626_o2), .dout(new_new_n1402__));
  buf1  g0464(.din(G1139_o2), .dout(new_new_n1403__));
  not1  g0465(.din(G1139_o2), .dout(new_new_n1404__));
  buf1  g0466(.din(G950_o2), .dout(new_new_n1405__));
  not1  g0467(.din(G950_o2), .dout(new_new_n1406__));
  buf1  g0468(.din(G707_o2), .dout(new_new_n1407__));
  not1  g0469(.din(G707_o2), .dout(new_new_n1408__));
  buf1  g0470(.din(G545_o2), .dout(new_new_n1409__));
  buf1  g0471(.din(G4217_o2), .dout(new_new_n1411__));
  not1  g0472(.din(G4217_o2), .dout(new_new_n1412__));
  buf1  g0473(.din(G4716_o2), .dout(new_new_n1413__));
  not1  g0474(.din(G4716_o2), .dout(new_new_n1414__));
  buf1  g0475(.din(G5244_o2), .dout(new_new_n1415__));
  not1  g0476(.din(G5244_o2), .dout(new_new_n1416__));
  buf1  g0477(.din(G3136_o2), .dout(new_new_n1417__));
  not1  g0478(.din(G3136_o2), .dout(new_new_n1418__));
  buf1  g0479(.din(G3499_o2), .dout(new_new_n1419__));
  not1  g0480(.din(G3499_o2), .dout(new_new_n1420__));
  buf1  g0481(.din(G3885_o2), .dout(new_new_n1421__));
  not1  g0482(.din(G3885_o2), .dout(new_new_n1422__));
  buf1  g0483(.din(G5243_o2), .dout(new_new_n1423__));
  not1  g0484(.din(G5243_o2), .dout(new_new_n1424__));
  buf1  g0485(.din(G3886_o2), .dout(new_new_n1425__));
  not1  g0486(.din(G3886_o2), .dout(new_new_n1426__));
  buf1  g0487(.din(G4375_o2), .dout(new_new_n1427__));
  not1  g0488(.din(G4375_o2), .dout(new_new_n1428__));
  buf1  g0489(.din(G4901_o2), .dout(new_new_n1429__));
  not1  g0490(.din(G4901_o2), .dout(new_new_n1430__));
  buf1  g0491(.din(G5054_o2), .dout(new_new_n1431__));
  not1  g0492(.din(G5054_o2), .dout(new_new_n1432__));
  buf1  g0493(.din(G4374_o2), .dout(new_new_n1433__));
  not1  g0494(.din(G4374_o2), .dout(new_new_n1434__));
  buf1  g0495(.din(G4900_o2), .dout(new_new_n1435__));
  not1  g0496(.din(G4900_o2), .dout(new_new_n1436__));
  buf1  g0497(.din(G5053_o2), .dout(new_new_n1437__));
  not1  g0498(.din(G5053_o2), .dout(new_new_n1438__));
  buf1  g0499(.din(G5242_o2), .dout(new_new_n1439__));
  not1  g0500(.din(G5242_o2), .dout(new_new_n1440__));
  buf1  g0501(.din(G4034_o2), .dout(new_new_n1441__));
  not1  g0502(.din(G4034_o2), .dout(new_new_n1442__));
  buf1  g0503(.din(G4556_o2), .dout(new_new_n1443__));
  not1  g0504(.din(G4556_o2), .dout(new_new_n1444__));
  buf1  g0505(.din(G5064_o2), .dout(new_new_n1445__));
  not1  g0506(.din(G5064_o2), .dout(new_new_n1446__));
  buf1  g0507(.din(G5172_o2), .dout(new_new_n1447__));
  not1  g0508(.din(G5172_o2), .dout(new_new_n1448__));
  buf1  g0509(.din(G2030_o2), .dout(new_new_n1449__));
  not1  g0510(.din(G2030_o2), .dout(new_new_n1450__));
  buf1  g0511(.din(G3016_o2), .dout(new_new_n1451__));
  not1  g0512(.din(G3016_o2), .dout(new_new_n1452__));
  buf1  g0513(.din(G3520_o2), .dout(new_new_n1453__));
  not1  g0514(.din(G3520_o2), .dout(new_new_n1454__));
  buf1  g0515(.din(G3261_o2), .dout(new_new_n1455__));
  not1  g0516(.din(G3261_o2), .dout(new_new_n1456__));
  buf1  g0517(.din(G3620_o2), .dout(new_new_n1457__));
  not1  g0518(.din(G3620_o2), .dout(new_new_n1458__));
  buf1  g0519(.din(G4220_o2), .dout(new_new_n1459__));
  not1  g0520(.din(G4220_o2), .dout(new_new_n1460__));
  buf1  g0521(.din(G4719_o2), .dout(new_new_n1461__));
  not1  g0522(.din(G4719_o2), .dout(new_new_n1462__));
  buf1  g0523(.din(G5247_o2), .dout(new_new_n1463__));
  not1  g0524(.din(G5247_o2), .dout(new_new_n1464__));
  buf1  g0525(.din(G5109_o2), .dout(new_new_n1465__));
  not1  g0526(.din(G5109_o2), .dout(new_new_n1466__));
  buf1  g0527(.din(G1638_o2), .dout(new_new_n1467__));
  not1  g0528(.din(G1638_o2), .dout(new_new_n1468__));
  buf1  g0529(.din(G1976_o2), .dout(new_new_n1469__));
  not1  g0530(.din(G1976_o2), .dout(new_new_n1470__));
  buf1  g0531(.din(G3560_o2), .dout(new_new_n1471__));
  not1  g0532(.din(G3560_o2), .dout(new_new_n1472__));
  buf1  g0533(.din(G3205_o2), .dout(new_new_n1473__));
  not1  g0534(.din(G3205_o2), .dout(new_new_n1474__));
  buf1  g0535(.din(G3193_o2), .dout(new_new_n1475__));
  not1  g0536(.din(G3193_o2), .dout(new_new_n1476__));
  buf1  g0537(.din(G3367_o2), .dout(new_new_n1477__));
  not1  g0538(.din(G3367_o2), .dout(new_new_n1478__));
  buf1  g0539(.din(G3670_o2), .dout(new_new_n1479__));
  not1  g0540(.din(G3670_o2), .dout(new_new_n1480__));
  buf1  g0541(.din(n979_inv), .dout(new_new_n1481__));
  buf1  g0542(.din(G1280_o2), .dout(new_new_n1483__));
  not1  g0543(.din(G1280_o2), .dout(new_new_n1484__));
  buf1  g0544(.din(G902_o2), .dout(new_new_n1485__));
  not1  g0545(.din(G902_o2), .dout(new_new_n1486__));
  buf1  g0546(.din(G659_o2), .dout(new_new_n1487__));
  not1  g0547(.din(G659_o2), .dout(new_new_n1488__));
  buf1  g0548(.din(G983_o2), .dout(new_new_n1489__));
  not1  g0549(.din(G983_o2), .dout(new_new_n1490__));
  buf1  g0550(.din(G740_o2), .dout(new_new_n1491__));
  not1  g0551(.din(G740_o2), .dout(new_new_n1492__));
  buf1  g0552(.din(G2917_o2), .dout(new_new_n1493__));
  not1  g0553(.din(G2917_o2), .dout(new_new_n1494__));
  buf1  g0554(.din(G3391_o2), .dout(new_new_n1495__));
  not1  g0555(.din(G3391_o2), .dout(new_new_n1496__));
  buf1  g0556(.din(G3494_o2), .dout(new_new_n1497__));
  not1  g0557(.din(G3494_o2), .dout(new_new_n1498__));
  buf1  g0558(.din(G1512_o2), .dout(new_new_n1499__));
  not1  g0559(.din(G1512_o2), .dout(new_new_n1500__));
  buf1  g0560(.din(G1854_o2), .dout(new_new_n1501__));
  not1  g0561(.din(G1854_o2), .dout(new_new_n1502__));
  buf1  g0562(.din(G2203_o2), .dout(new_new_n1503__));
  not1  g0563(.din(G2203_o2), .dout(new_new_n1504__));
  buf1  g0564(.din(G3493_o2), .dout(new_new_n1505__));
  not1  g0565(.din(G3493_o2), .dout(new_new_n1506__));
  buf1  g0566(.din(G3069_o2), .dout(new_new_n1507__));
  not1  g0567(.din(G3069_o2), .dout(new_new_n1508__));
  buf1  g0568(.din(G3574_o2), .dout(new_new_n1509__));
  not1  g0569(.din(G3574_o2), .dout(new_new_n1510__));
  buf1  g0570(.din(G3319_o2), .dout(new_new_n1511__));
  not1  g0571(.din(G3319_o2), .dout(new_new_n1512__));
  buf1  g0572(.din(G3667_o2), .dout(new_new_n1513__));
  not1  g0573(.din(G3667_o2), .dout(new_new_n1514__));
  buf1  g0574(.din(G3068_o2), .dout(new_new_n1515__));
  not1  g0575(.din(G3068_o2), .dout(new_new_n1516__));
  buf1  g0576(.din(G3573_o2), .dout(new_new_n1517__));
  not1  g0577(.din(G3573_o2), .dout(new_new_n1518__));
  buf1  g0578(.din(G3666_o2), .dout(new_new_n1519__));
  not1  g0579(.din(G3666_o2), .dout(new_new_n1520__));
  buf1  g0580(.din(G3318_o2), .dout(new_new_n1521__));
  not1  g0581(.din(G3318_o2), .dout(new_new_n1522__));
  buf1  g0582(.din(G3492_o2), .dout(new_new_n1523__));
  not1  g0583(.din(G3492_o2), .dout(new_new_n1524__));
  buf1  g0584(.din(G3241_o2), .dout(new_new_n1525__));
  not1  g0585(.din(G3241_o2), .dout(new_new_n1526__));
  buf1  g0586(.din(G3722_o2), .dout(new_new_n1527__));
  not1  g0587(.din(G3722_o2), .dout(new_new_n1528__));
  buf1  g0588(.din(G3422_o2), .dout(new_new_n1529__));
  not1  g0589(.din(G3422_o2), .dout(new_new_n1530__));
  buf1  g0590(.din(G1445_o2), .dout(new_new_n1531__));
  buf1  g0591(.din(G3257_o2), .dout(new_new_n1533__));
  not1  g0592(.din(G3257_o2), .dout(new_new_n1534__));
  buf1  g0593(.din(G3616_o2), .dout(new_new_n1535__));
  not1  g0594(.din(G3616_o2), .dout(new_new_n1536__));
  buf1  g0595(.din(G1634_o2), .dout(new_new_n1537__));
  not1  g0596(.din(G1634_o2), .dout(new_new_n1538__));
  buf1  g0597(.din(G1972_o2), .dout(new_new_n1539__));
  not1  g0598(.din(G1972_o2), .dout(new_new_n1540__));
  buf1  g0599(.din(G2256_o2), .dout(new_new_n1541__));
  not1  g0600(.din(G2256_o2), .dout(new_new_n1542__));
  buf1  g0601(.din(G3394_o2), .dout(new_new_n1543__));
  not1  g0602(.din(G3394_o2), .dout(new_new_n1544__));
  buf1  g0603(.din(G3557_o2), .dout(new_new_n1545__));
  not1  g0604(.din(G3557_o2), .dout(new_new_n1546__));
  buf1  g0605(.din(G3364_o2), .dout(new_new_n1547__));
  not1  g0606(.din(G3364_o2), .dout(new_new_n1548__));
  buf1  g0607(.din(G3719_o2), .dout(new_new_n1549__));
  not1  g0608(.din(G3719_o2), .dout(new_new_n1550__));
  buf1  g0609(.din(G2253_o2), .dout(new_new_n1551__));
  not1  g0610(.din(G2253_o2), .dout(new_new_n1552__));
  buf1  g0611(.din(G1583_o2), .dout(new_new_n1553__));
  not1  g0612(.din(G1583_o2), .dout(new_new_n1554__));
  buf1  g0613(.din(G1917_o2), .dout(new_new_n1555__));
  not1  g0614(.din(G1917_o2), .dout(new_new_n1556__));
  buf1  g0615(.din(G1727_o2), .dout(new_new_n1557__));
  not1  g0616(.din(G1727_o2), .dout(new_new_n1558__));
  buf1  g0617(.din(G2061_o2), .dout(new_new_n1559__));
  not1  g0618(.din(G2061_o2), .dout(new_new_n1560__));
  buf1  g0619(.din(G935_o2), .dout(new_new_n1561__));
  not1  g0620(.din(G935_o2), .dout(new_new_n1562__));
  buf1  g0621(.din(G692_o2), .dout(new_new_n1563__));
  not1  g0622(.din(G692_o2), .dout(new_new_n1564__));
  buf1  g0623(.din(G2136_o2), .dout(new_new_n1565__));
  not1  g0624(.din(G2136_o2), .dout(new_new_n1566__));
  buf1  g0625(.din(G1507_o2), .dout(new_new_n1567__));
  not1  g0626(.din(G1507_o2), .dout(new_new_n1568__));
  buf1  g0627(.din(G1849_o2), .dout(new_new_n1569__));
  not1  g0628(.din(G1849_o2), .dout(new_new_n1570__));
  buf1  g0629(.din(G2198_o2), .dout(new_new_n1571__));
  not1  g0630(.din(G2198_o2), .dout(new_new_n1572__));
  buf1  g0631(.din(G2197_o2), .dout(new_new_n1573__));
  not1  g0632(.din(G2197_o2), .dout(new_new_n1574__));
  buf1  g0633(.din(G1848_o2), .dout(new_new_n1575__));
  not1  g0634(.din(G1848_o2), .dout(new_new_n1576__));
  buf1  g0635(.din(G1689_o2), .dout(new_new_n1577__));
  not1  g0636(.din(G1689_o2), .dout(new_new_n1578__));
  buf1  g0637(.din(G2016_o2), .dout(new_new_n1579__));
  not1  g0638(.din(G2016_o2), .dout(new_new_n1580__));
  buf1  g0639(.din(G2314_o2), .dout(new_new_n1581__));
  not1  g0640(.din(G2314_o2), .dout(new_new_n1582__));
  buf1  g0641(.din(G2313_o2), .dout(new_new_n1583__));
  not1  g0642(.din(G2313_o2), .dout(new_new_n1584__));
  buf1  g0643(.din(G1688_o2), .dout(new_new_n1585__));
  not1  g0644(.din(G1688_o2), .dout(new_new_n1586__));
  buf1  g0645(.din(G2015_o2), .dout(new_new_n1587__));
  not1  g0646(.din(G2015_o2), .dout(new_new_n1588__));
  buf1  g0647(.din(G1847_o2), .dout(new_new_n1589__));
  not1  g0648(.din(G1847_o2), .dout(new_new_n1590__));
  buf1  g0649(.din(G2196_o2), .dout(new_new_n1591__));
  not1  g0650(.din(G2196_o2), .dout(new_new_n1592__));
  buf1  g0651(.din(G2118_o2), .dout(new_new_n1593__));
  not1  g0652(.din(G2118_o2), .dout(new_new_n1594__));
  buf1  g0653(.din(G1777_o2), .dout(new_new_n1595__));
  not1  g0654(.din(G1777_o2), .dout(new_new_n1596__));
  buf1  g0655(.din(G1630_o2), .dout(new_new_n1597__));
  not1  g0656(.din(G1630_o2), .dout(new_new_n1598__));
  buf1  g0657(.din(G1968_o2), .dout(new_new_n1599__));
  not1  g0658(.din(G1968_o2), .dout(new_new_n1600__));
  buf1  g0659(.din(G2309_o2), .dout(new_new_n1601__));
  not1  g0660(.din(G2309_o2), .dout(new_new_n1602__));
  buf1  g0661(.din(G2139_o2), .dout(new_new_n1603__));
  not1  g0662(.din(G2139_o2), .dout(new_new_n1604__));
  buf1  g0663(.din(G1580_o2), .dout(new_new_n1605__));
  not1  g0664(.din(G1580_o2), .dout(new_new_n1606__));
  buf1  g0665(.din(G2250_o2), .dout(new_new_n1607__));
  not1  g0666(.din(G2250_o2), .dout(new_new_n1608__));
  buf1  g0667(.din(G1914_o2), .dout(new_new_n1609__));
  not1  g0668(.din(G1914_o2), .dout(new_new_n1610__));
  buf1  g0669(.din(G1724_o2), .dout(new_new_n1611__));
  not1  g0670(.din(G1724_o2), .dout(new_new_n1612__));
  buf1  g0671(.din(G2058_o2), .dout(new_new_n1613__));
  not1  g0672(.din(G2058_o2), .dout(new_new_n1614__));
  buf1  g0673(.din(n2728_lo_buf_o2), .dout(new_new_n1615__));
  not1  g0674(.din(n2728_lo_buf_o2), .dout(new_new_n1616__));
  and1  g0675(.dina(new_new_n893__), .dinb(new_new_n873__), .dout(new_new_n1617__));
  or1   g0676(.dina(new_new_n6352__), .dinb(new_new_n946__), .dout(new_new_n1618__));
  or1   g0677(.dina(new_new_n6352__), .dinb(new_new_n943__), .dout(new_new_n1619__));
  and1  g0678(.dina(new_new_n1619__), .dinb(new_new_n1618__), .dout(new_new_n1620__));
  or1   g0679(.dina(new_new_n6353__), .dinb(new_new_n952__), .dout(new_new_n1621__));
  or1   g0680(.dina(new_new_n6353__), .dinb(new_new_n949__), .dout(new_new_n1622__));
  and1  g0681(.dina(new_new_n1622__), .dinb(new_new_n1621__), .dout(new_new_n1623__));
  or1   g0682(.dina(new_new_n6354__), .dinb(new_new_n958__), .dout(new_new_n1624__));
  or1   g0683(.dina(new_new_n6354__), .dinb(new_new_n955__), .dout(new_new_n1625__));
  and1  g0684(.dina(new_new_n1625__), .dinb(new_new_n1624__), .dout(new_new_n1626__));
  or1   g0685(.dina(new_new_n6355__), .dinb(new_new_n964__), .dout(new_new_n1627__));
  or1   g0686(.dina(new_new_n6355__), .dinb(new_new_n961__), .dout(new_new_n1628__));
  and1  g0687(.dina(new_new_n1628__), .dinb(new_new_n1627__), .dout(new_new_n1629__));
  or1   g0688(.dina(new_new_n6356__), .dinb(new_new_n970__), .dout(new_new_n1630__));
  or1   g0689(.dina(new_new_n6356__), .dinb(new_new_n967__), .dout(new_new_n1631__));
  and1  g0690(.dina(new_new_n1631__), .dinb(new_new_n1630__), .dout(new_new_n1632__));
  or1   g0691(.dina(new_new_n6357__), .dinb(new_new_n976__), .dout(new_new_n1633__));
  or1   g0692(.dina(new_new_n6357__), .dinb(new_new_n973__), .dout(new_new_n1634__));
  and1  g0693(.dina(new_new_n1634__), .dinb(new_new_n1633__), .dout(new_new_n1635__));
  or1   g0694(.dina(new_new_n6358__), .dinb(new_new_n982__), .dout(new_new_n1636__));
  or1   g0695(.dina(new_new_n6358__), .dinb(new_new_n979__), .dout(new_new_n1637__));
  and1  g0696(.dina(new_new_n1637__), .dinb(new_new_n1636__), .dout(new_new_n1638__));
  or1   g0697(.dina(new_new_n6359__), .dinb(new_new_n988__), .dout(new_new_n1639__));
  or1   g0698(.dina(new_new_n6359__), .dinb(new_new_n985__), .dout(new_new_n1640__));
  and1  g0699(.dina(new_new_n1640__), .dinb(new_new_n1639__), .dout(new_new_n1641__));
  or1   g0700(.dina(new_new_n6360__), .dinb(new_new_n994__), .dout(new_new_n1642__));
  or1   g0701(.dina(new_new_n6360__), .dinb(new_new_n991__), .dout(new_new_n1643__));
  and1  g0702(.dina(new_new_n1643__), .dinb(new_new_n1642__), .dout(new_new_n1644__));
  or1   g0703(.dina(new_new_n6361__), .dinb(new_new_n1006__), .dout(new_new_n1645__));
  or1   g0704(.dina(new_new_n6361__), .dinb(new_new_n1001__), .dout(new_new_n1646__));
  and1  g0705(.dina(new_new_n1646__), .dinb(new_new_n1645__), .dout(new_new_n1647__));
  or1   g0706(.dina(new_new_n6362__), .dinb(new_new_n1032__), .dout(new_new_n1648__));
  or1   g0707(.dina(new_new_n6362__), .dinb(new_new_n1027__), .dout(new_new_n1649__));
  and1  g0708(.dina(new_new_n1649__), .dinb(new_new_n1648__), .dout(new_new_n1650__));
  or1   g0709(.dina(new_new_n6363__), .dinb(new_new_n1052__), .dout(new_new_n1651__));
  or1   g0710(.dina(new_new_n6363__), .dinb(new_new_n1049__), .dout(new_new_n1652__));
  and1  g0711(.dina(new_new_n1652__), .dinb(new_new_n1651__), .dout(new_new_n1653__));
  or1   g0712(.dina(new_new_n6364__), .dinb(new_new_n1070__), .dout(new_new_n1654__));
  or1   g0713(.dina(new_new_n6364__), .dinb(new_new_n1067__), .dout(new_new_n1655__));
  and1  g0714(.dina(new_new_n1655__), .dinb(new_new_n1654__), .dout(new_new_n1656__));
  or1   g0715(.dina(new_new_n6365__), .dinb(new_new_n1088__), .dout(new_new_n1657__));
  or1   g0716(.dina(new_new_n6365__), .dinb(new_new_n1085__), .dout(new_new_n1658__));
  and1  g0717(.dina(new_new_n1658__), .dinb(new_new_n1657__), .dout(new_new_n1659__));
  or1   g0718(.dina(new_new_n6366__), .dinb(new_new_n1136__), .dout(new_new_n1660__));
  or1   g0719(.dina(new_new_n6366__), .dinb(new_new_n1133__), .dout(new_new_n1661__));
  and1  g0720(.dina(new_new_n1661__), .dinb(new_new_n1660__), .dout(new_new_n1662__));
  or1   g0721(.dina(new_new_n6367__), .dinb(new_new_n1180__), .dout(new_new_n1663__));
  and1  g0722(.dina(new_new_n1663__), .dinb(new_new_n6367__), .dout(new_new_n1664__));
  or1   g0723(.dina(new_new_n6368__), .dinb(new_new_n1222__), .dout(new_new_n1665__));
  or1   g0724(.dina(new_new_n6368__), .dinb(new_new_n1211__), .dout(new_new_n1666__));
  and1  g0725(.dina(new_new_n1666__), .dinb(new_new_n1665__), .dout(new_new_n1667__));
  or1   g0726(.dina(new_new_n6370__), .dinb(new_new_n1290__), .dout(new_new_n1668__));
  or1   g0727(.dina(new_new_n6370__), .dinb(new_new_n1275__), .dout(new_new_n1669__));
  and1  g0728(.dina(new_new_n1669__), .dinb(new_new_n1668__), .dout(new_new_n1670__));
  and1  g0729(.dina(new_new_n1350__), .dinb(new_new_n1348__), .dout(new_new_n1671__));
  or1   g0730(.dina(new_new_n1349__), .dinb(new_new_n1347__), .dout(new_new_n1672__));
  and1  g0731(.dina(new_new_n1362__), .dinb(new_new_n1219__), .dout(new_new_n1673__));
  or1   g0732(.dina(new_new_n6369__), .dinb(new_new_n1220__), .dout(new_new_n1674__));
  and1  g0733(.dina(new_new_n1674__), .dinb(new_new_n1672__), .dout(new_new_n1675__));
  or1   g0734(.dina(new_new_n6371__), .dinb(new_new_n6372__), .dout(new_new_n1676__));
  or1   g0735(.dina(new_new_n6374__), .dinb(new_new_n6372__), .dout(new_new_n1677__));
  or1   g0736(.dina(new_new_n6374__), .dinb(new_new_n6371__), .dout(new_new_n1678__));
  and1  g0737(.dina(new_new_n1678__), .dinb(new_new_n1677__), .dout(new_new_n1679__));
  and1  g0738(.dina(new_new_n6375__), .dinb(new_new_n6376__), .dout(new_new_n1680__));
  or1   g0739(.dina(new_new_n6377__), .dinb(new_new_n6378__), .dout(new_new_n1681__));
  and1  g0740(.dina(new_new_n6380__), .dinb(new_new_n6375__), .dout(new_new_n1682__));
  or1   g0741(.dina(new_new_n6382__), .dinb(new_new_n6377__), .dout(new_new_n1683__));
  and1  g0742(.dina(new_new_n6380__), .dinb(new_new_n6376__), .dout(new_new_n1684__));
  or1   g0743(.dina(new_new_n6382__), .dinb(new_new_n6378__), .dout(new_new_n1685__));
  and1  g0744(.dina(new_new_n1685__), .dinb(new_new_n1683__), .dout(new_new_n1686__));
  or1   g0745(.dina(new_new_n1684__), .dinb(new_new_n1682__), .dout(new_new_n1687__));
  and1  g0746(.dina(new_new_n1676__), .dinb(new_new_n1281__), .dout(new_new_n1688__));
  or1   g0747(.dina(new_new_n6373__), .dinb(new_new_n1282__), .dout(new_new_n1689__));
  and1  g0748(.dina(new_new_n1689__), .dinb(new_new_n1687__), .dout(new_new_n1690__));
  or1   g0749(.dina(new_new_n6383__), .dinb(new_new_n6384__), .dout(new_new_n1691__));
  or1   g0750(.dina(new_new_n6386__), .dinb(new_new_n6384__), .dout(new_new_n1692__));
  or1   g0751(.dina(new_new_n6386__), .dinb(new_new_n6383__), .dout(new_new_n1693__));
  and1  g0752(.dina(new_new_n1693__), .dinb(new_new_n1692__), .dout(new_new_n1694__));
  and1  g0753(.dina(new_new_n6388__), .dinb(new_new_n1287__), .dout(new_new_n1695__));
  or1   g0754(.dina(new_new_n6390__), .dinb(new_new_n1288__), .dout(new_new_n1696__));
  and1  g0755(.dina(new_new_n6388__), .dinb(new_new_n1270__), .dout(new_new_n1697__));
  or1   g0756(.dina(new_new_n6390__), .dinb(new_new_n1269__), .dout(new_new_n1698__));
  and1  g0757(.dina(new_new_n1698__), .dinb(new_new_n1696__), .dout(new_new_n1699__));
  or1   g0758(.dina(new_new_n1697__), .dinb(new_new_n1695__), .dout(new_new_n1700__));
  and1  g0759(.dina(new_new_n1236__), .dinb(new_new_n1177__), .dout(new_new_n1701__));
  or1   g0760(.dina(new_new_n1235__), .dinb(new_new_n1178__), .dout(new_new_n1702__));
  and1  g0761(.dina(new_new_n6391__), .dinb(new_new_n6392__), .dout(new_new_n1703__));
  or1   g0762(.dina(new_new_n6393__), .dinb(new_new_n6394__), .dout(new_new_n1704__));
  and1  g0763(.dina(new_new_n6396__), .dinb(new_new_n6392__), .dout(new_new_n1705__));
  or1   g0764(.dina(new_new_n6398__), .dinb(new_new_n6394__), .dout(new_new_n1706__));
  and1  g0765(.dina(new_new_n6396__), .dinb(new_new_n6391__), .dout(new_new_n1707__));
  or1   g0766(.dina(new_new_n6398__), .dinb(new_new_n6393__), .dout(new_new_n1708__));
  and1  g0767(.dina(new_new_n1708__), .dinb(new_new_n1706__), .dout(new_new_n1709__));
  or1   g0768(.dina(new_new_n1707__), .dinb(new_new_n1705__), .dout(new_new_n1710__));
  and1  g0769(.dina(new_new_n1691__), .dinb(new_new_n6379__), .dout(new_new_n1711__));
  or1   g0770(.dina(new_new_n6385__), .dinb(new_new_n6381__), .dout(new_new_n1712__));
  and1  g0771(.dina(new_new_n1712__), .dinb(new_new_n1710__), .dout(new_new_n1713__));
  or1   g0772(.dina(new_new_n6399__), .dinb(new_new_n6400__), .dout(new_new_n1714__));
  or1   g0773(.dina(new_new_n6402__), .dinb(new_new_n6400__), .dout(new_new_n1715__));
  or1   g0774(.dina(new_new_n6402__), .dinb(new_new_n6399__), .dout(new_new_n1716__));
  and1  g0775(.dina(new_new_n1716__), .dinb(new_new_n1715__), .dout(new_new_n1717__));
  and1  g0776(.dina(new_new_n1352__), .dinb(new_new_n1346__), .dout(new_new_n1718__));
  or1   g0777(.dina(new_new_n1351__), .dinb(new_new_n1345__), .dout(new_new_n1719__));
  and1  g0778(.dina(new_new_n6406__), .dinb(new_new_n875__), .dout(new_new_n1720__));
  or1   g0779(.dina(new_new_n6414__), .dinb(new_new_n876__), .dout(new_new_n1721__));
  and1  g0780(.dina(new_new_n6419__), .dinb(new_new_n6420__), .dout(new_new_n1722__));
  or1   g0781(.dina(new_new_n6421__), .dinb(new_new_n6422__), .dout(new_new_n1723__));
  and1  g0782(.dina(new_new_n6424__), .dinb(new_new_n6420__), .dout(new_new_n1724__));
  or1   g0783(.dina(new_new_n6426__), .dinb(new_new_n6422__), .dout(new_new_n1725__));
  and1  g0784(.dina(new_new_n6424__), .dinb(new_new_n6419__), .dout(new_new_n1726__));
  or1   g0785(.dina(new_new_n6426__), .dinb(new_new_n6421__), .dout(new_new_n1727__));
  and1  g0786(.dina(new_new_n1727__), .dinb(new_new_n1725__), .dout(new_new_n1728__));
  or1   g0787(.dina(new_new_n1726__), .dinb(new_new_n1724__), .dout(new_new_n1729__));
  and1  g0788(.dina(new_new_n6387__), .dinb(new_new_n1217__), .dout(new_new_n1730__));
  or1   g0789(.dina(new_new_n6389__), .dinb(new_new_n1218__), .dout(new_new_n1731__));
  and1  g0790(.dina(new_new_n6427__), .dinb(new_new_n6428__), .dout(new_new_n1732__));
  or1   g0791(.dina(new_new_n6429__), .dinb(new_new_n6430__), .dout(new_new_n1733__));
  and1  g0792(.dina(new_new_n6432__), .dinb(new_new_n6428__), .dout(new_new_n1734__));
  or1   g0793(.dina(new_new_n6434__), .dinb(new_new_n6430__), .dout(new_new_n1735__));
  and1  g0794(.dina(new_new_n6432__), .dinb(new_new_n6427__), .dout(new_new_n1736__));
  or1   g0795(.dina(new_new_n6434__), .dinb(new_new_n6429__), .dout(new_new_n1737__));
  and1  g0796(.dina(new_new_n1737__), .dinb(new_new_n1735__), .dout(new_new_n1738__));
  or1   g0797(.dina(new_new_n1736__), .dinb(new_new_n1734__), .dout(new_new_n1739__));
  and1  g0798(.dina(new_new_n1714__), .dinb(new_new_n6395__), .dout(new_new_n1740__));
  or1   g0799(.dina(new_new_n6401__), .dinb(new_new_n6397__), .dout(new_new_n1741__));
  and1  g0800(.dina(new_new_n1741__), .dinb(new_new_n1739__), .dout(new_new_n1742__));
  or1   g0801(.dina(new_new_n6435__), .dinb(new_new_n6436__), .dout(new_new_n1743__));
  or1   g0802(.dina(new_new_n6438__), .dinb(new_new_n6436__), .dout(new_new_n1744__));
  or1   g0803(.dina(new_new_n6438__), .dinb(new_new_n6435__), .dout(new_new_n1745__));
  and1  g0804(.dina(new_new_n1745__), .dinb(new_new_n1744__), .dout(new_new_n1746__));
  and1  g0805(.dina(new_new_n6439__), .dinb(new_new_n6440__), .dout(new_new_n1747__));
  or1   g0806(.dina(new_new_n6441__), .dinb(new_new_n6442__), .dout(new_new_n1748__));
  and1  g0807(.dina(new_new_n6444__), .dinb(new_new_n6439__), .dout(new_new_n1749__));
  or1   g0808(.dina(new_new_n6446__), .dinb(new_new_n6441__), .dout(new_new_n1750__));
  and1  g0809(.dina(new_new_n6444__), .dinb(new_new_n6440__), .dout(new_new_n1751__));
  or1   g0810(.dina(new_new_n6446__), .dinb(new_new_n6442__), .dout(new_new_n1752__));
  and1  g0811(.dina(new_new_n1752__), .dinb(new_new_n1750__), .dout(new_new_n1753__));
  or1   g0812(.dina(new_new_n1751__), .dinb(new_new_n1749__), .dout(new_new_n1754__));
  and1  g0813(.dina(new_new_n6406__), .dinb(new_new_n877__), .dout(new_new_n1755__));
  or1   g0814(.dina(new_new_n6414__), .dinb(new_new_n878__), .dout(new_new_n1756__));
  and1  g0815(.dina(new_new_n6447__), .dinb(new_new_n6448__), .dout(new_new_n1757__));
  or1   g0816(.dina(new_new_n6449__), .dinb(new_new_n6450__), .dout(new_new_n1758__));
  and1  g0817(.dina(new_new_n6452__), .dinb(new_new_n6448__), .dout(new_new_n1759__));
  or1   g0818(.dina(new_new_n6454__), .dinb(new_new_n6450__), .dout(new_new_n1760__));
  and1  g0819(.dina(new_new_n6452__), .dinb(new_new_n6447__), .dout(new_new_n1761__));
  or1   g0820(.dina(new_new_n6454__), .dinb(new_new_n6449__), .dout(new_new_n1762__));
  and1  g0821(.dina(new_new_n1762__), .dinb(new_new_n1760__), .dout(new_new_n1763__));
  or1   g0822(.dina(new_new_n1761__), .dinb(new_new_n1759__), .dout(new_new_n1764__));
  and1  g0823(.dina(new_new_n6423__), .dinb(new_new_n1279__), .dout(new_new_n1765__));
  or1   g0824(.dina(new_new_n6425__), .dinb(new_new_n1280__), .dout(new_new_n1766__));
  and1  g0825(.dina(new_new_n6455__), .dinb(new_new_n6456__), .dout(new_new_n1767__));
  or1   g0826(.dina(new_new_n6457__), .dinb(new_new_n6458__), .dout(new_new_n1768__));
  and1  g0827(.dina(new_new_n6460__), .dinb(new_new_n6456__), .dout(new_new_n1769__));
  or1   g0828(.dina(new_new_n6462__), .dinb(new_new_n6458__), .dout(new_new_n1770__));
  and1  g0829(.dina(new_new_n6460__), .dinb(new_new_n6455__), .dout(new_new_n1771__));
  or1   g0830(.dina(new_new_n6462__), .dinb(new_new_n6457__), .dout(new_new_n1772__));
  and1  g0831(.dina(new_new_n1772__), .dinb(new_new_n1770__), .dout(new_new_n1773__));
  or1   g0832(.dina(new_new_n1771__), .dinb(new_new_n1769__), .dout(new_new_n1774__));
  and1  g0833(.dina(new_new_n1743__), .dinb(new_new_n6431__), .dout(new_new_n1775__));
  or1   g0834(.dina(new_new_n6437__), .dinb(new_new_n6433__), .dout(new_new_n1776__));
  and1  g0835(.dina(new_new_n1776__), .dinb(new_new_n1774__), .dout(new_new_n1777__));
  or1   g0836(.dina(new_new_n6463__), .dinb(new_new_n6464__), .dout(new_new_n1778__));
  or1   g0837(.dina(new_new_n6466__), .dinb(new_new_n6464__), .dout(new_new_n1779__));
  or1   g0838(.dina(new_new_n6466__), .dinb(new_new_n6463__), .dout(new_new_n1780__));
  and1  g0839(.dina(new_new_n1780__), .dinb(new_new_n1779__), .dout(new_new_n1781__));
  and1  g0840(.dina(new_new_n6468__), .dinb(new_new_n1285__), .dout(new_new_n1782__));
  or1   g0841(.dina(new_new_n6470__), .dinb(new_new_n1286__), .dout(new_new_n1783__));
  and1  g0842(.dina(new_new_n6468__), .dinb(new_new_n1272__), .dout(new_new_n1784__));
  or1   g0843(.dina(new_new_n6470__), .dinb(new_new_n1271__), .dout(new_new_n1785__));
  and1  g0844(.dina(new_new_n1785__), .dinb(new_new_n1783__), .dout(new_new_n1786__));
  or1   g0845(.dina(new_new_n1784__), .dinb(new_new_n1782__), .dout(new_new_n1787__));
  and1  g0846(.dina(new_new_n1238__), .dinb(new_new_n1175__), .dout(new_new_n1788__));
  or1   g0847(.dina(new_new_n1237__), .dinb(new_new_n1176__), .dout(new_new_n1789__));
  and1  g0848(.dina(new_new_n6471__), .dinb(new_new_n6472__), .dout(new_new_n1790__));
  or1   g0849(.dina(new_new_n6473__), .dinb(new_new_n6474__), .dout(new_new_n1791__));
  and1  g0850(.dina(new_new_n6476__), .dinb(new_new_n6472__), .dout(new_new_n1792__));
  or1   g0851(.dina(new_new_n6478__), .dinb(new_new_n6474__), .dout(new_new_n1793__));
  and1  g0852(.dina(new_new_n6476__), .dinb(new_new_n6471__), .dout(new_new_n1794__));
  or1   g0853(.dina(new_new_n6478__), .dinb(new_new_n6473__), .dout(new_new_n1795__));
  and1  g0854(.dina(new_new_n1795__), .dinb(new_new_n1793__), .dout(new_new_n1796__));
  or1   g0855(.dina(new_new_n1794__), .dinb(new_new_n1792__), .dout(new_new_n1797__));
  and1  g0856(.dina(new_new_n6405__), .dinb(new_new_n879__), .dout(new_new_n1798__));
  or1   g0857(.dina(new_new_n6413__), .dinb(new_new_n880__), .dout(new_new_n1799__));
  and1  g0858(.dina(new_new_n6479__), .dinb(new_new_n6480__), .dout(new_new_n1800__));
  or1   g0859(.dina(new_new_n6481__), .dinb(new_new_n6482__), .dout(new_new_n1801__));
  and1  g0860(.dina(new_new_n6484__), .dinb(new_new_n6480__), .dout(new_new_n1802__));
  or1   g0861(.dina(new_new_n6486__), .dinb(new_new_n6482__), .dout(new_new_n1803__));
  and1  g0862(.dina(new_new_n6484__), .dinb(new_new_n6479__), .dout(new_new_n1804__));
  or1   g0863(.dina(new_new_n6486__), .dinb(new_new_n6481__), .dout(new_new_n1805__));
  and1  g0864(.dina(new_new_n1805__), .dinb(new_new_n1803__), .dout(new_new_n1806__));
  or1   g0865(.dina(new_new_n1804__), .dinb(new_new_n1802__), .dout(new_new_n1807__));
  and1  g0866(.dina(new_new_n6451__), .dinb(new_new_n6443__), .dout(new_new_n1808__));
  or1   g0867(.dina(new_new_n6453__), .dinb(new_new_n6445__), .dout(new_new_n1809__));
  and1  g0868(.dina(new_new_n6487__), .dinb(new_new_n6488__), .dout(new_new_n1810__));
  or1   g0869(.dina(new_new_n6489__), .dinb(new_new_n6490__), .dout(new_new_n1811__));
  and1  g0870(.dina(new_new_n6492__), .dinb(new_new_n6488__), .dout(new_new_n1812__));
  or1   g0871(.dina(new_new_n6494__), .dinb(new_new_n6490__), .dout(new_new_n1813__));
  and1  g0872(.dina(new_new_n6492__), .dinb(new_new_n6487__), .dout(new_new_n1814__));
  or1   g0873(.dina(new_new_n6494__), .dinb(new_new_n6489__), .dout(new_new_n1815__));
  and1  g0874(.dina(new_new_n1815__), .dinb(new_new_n1813__), .dout(new_new_n1816__));
  or1   g0875(.dina(new_new_n1814__), .dinb(new_new_n1812__), .dout(new_new_n1817__));
  and1  g0876(.dina(new_new_n1778__), .dinb(new_new_n6459__), .dout(new_new_n1818__));
  or1   g0877(.dina(new_new_n6465__), .dinb(new_new_n6461__), .dout(new_new_n1819__));
  and1  g0878(.dina(new_new_n1819__), .dinb(new_new_n1817__), .dout(new_new_n1820__));
  or1   g0879(.dina(new_new_n6495__), .dinb(new_new_n6496__), .dout(new_new_n1821__));
  or1   g0880(.dina(new_new_n6498__), .dinb(new_new_n6496__), .dout(new_new_n1822__));
  or1   g0881(.dina(new_new_n6498__), .dinb(new_new_n6495__), .dout(new_new_n1823__));
  and1  g0882(.dina(new_new_n1823__), .dinb(new_new_n1822__), .dout(new_new_n1824__));
  and1  g0883(.dina(new_new_n1354__), .dinb(new_new_n1344__), .dout(new_new_n1825__));
  or1   g0884(.dina(new_new_n1353__), .dinb(new_new_n1343__), .dout(new_new_n1826__));
  and1  g0885(.dina(new_new_n6501__), .dinb(new_new_n6503__), .dout(new_new_n1827__));
  or1   g0886(.dina(new_new_n6506__), .dinb(new_new_n6508__), .dout(new_new_n1828__));
  and1  g0887(.dina(new_new_n6509__), .dinb(new_new_n6510__), .dout(new_new_n1829__));
  or1   g0888(.dina(new_new_n6511__), .dinb(new_new_n6512__), .dout(new_new_n1830__));
  and1  g0889(.dina(new_new_n6514__), .dinb(new_new_n6510__), .dout(new_new_n1831__));
  or1   g0890(.dina(new_new_n6516__), .dinb(new_new_n6512__), .dout(new_new_n1832__));
  and1  g0891(.dina(new_new_n6514__), .dinb(new_new_n6509__), .dout(new_new_n1833__));
  or1   g0892(.dina(new_new_n6516__), .dinb(new_new_n6511__), .dout(new_new_n1834__));
  and1  g0893(.dina(new_new_n1834__), .dinb(new_new_n1832__), .dout(new_new_n1835__));
  or1   g0894(.dina(new_new_n1833__), .dinb(new_new_n1831__), .dout(new_new_n1836__));
  and1  g0895(.dina(new_new_n6467__), .dinb(new_new_n1215__), .dout(new_new_n1837__));
  or1   g0896(.dina(new_new_n6469__), .dinb(new_new_n1216__), .dout(new_new_n1838__));
  and1  g0897(.dina(new_new_n6517__), .dinb(new_new_n6518__), .dout(new_new_n1839__));
  or1   g0898(.dina(new_new_n6519__), .dinb(new_new_n6520__), .dout(new_new_n1840__));
  and1  g0899(.dina(new_new_n6522__), .dinb(new_new_n6518__), .dout(new_new_n1841__));
  or1   g0900(.dina(new_new_n6524__), .dinb(new_new_n6520__), .dout(new_new_n1842__));
  and1  g0901(.dina(new_new_n6522__), .dinb(new_new_n6517__), .dout(new_new_n1843__));
  or1   g0902(.dina(new_new_n6524__), .dinb(new_new_n6519__), .dout(new_new_n1844__));
  and1  g0903(.dina(new_new_n1844__), .dinb(new_new_n1842__), .dout(new_new_n1845__));
  or1   g0904(.dina(new_new_n1843__), .dinb(new_new_n1841__), .dout(new_new_n1846__));
  and1  g0905(.dina(new_new_n6407__), .dinb(new_new_n881__), .dout(new_new_n1847__));
  or1   g0906(.dina(new_new_n6415__), .dinb(new_new_n882__), .dout(new_new_n1848__));
  and1  g0907(.dina(new_new_n6525__), .dinb(new_new_n6526__), .dout(new_new_n1849__));
  or1   g0908(.dina(new_new_n6527__), .dinb(new_new_n6528__), .dout(new_new_n1850__));
  and1  g0909(.dina(new_new_n6530__), .dinb(new_new_n6526__), .dout(new_new_n1851__));
  or1   g0910(.dina(new_new_n6532__), .dinb(new_new_n6528__), .dout(new_new_n1852__));
  and1  g0911(.dina(new_new_n6530__), .dinb(new_new_n6525__), .dout(new_new_n1853__));
  or1   g0912(.dina(new_new_n6532__), .dinb(new_new_n6527__), .dout(new_new_n1854__));
  and1  g0913(.dina(new_new_n1854__), .dinb(new_new_n1852__), .dout(new_new_n1855__));
  or1   g0914(.dina(new_new_n1853__), .dinb(new_new_n1851__), .dout(new_new_n1856__));
  and1  g0915(.dina(new_new_n6483__), .dinb(new_new_n6475__), .dout(new_new_n1857__));
  or1   g0916(.dina(new_new_n6485__), .dinb(new_new_n6477__), .dout(new_new_n1858__));
  and1  g0917(.dina(new_new_n6533__), .dinb(new_new_n6534__), .dout(new_new_n1859__));
  or1   g0918(.dina(new_new_n6535__), .dinb(new_new_n6536__), .dout(new_new_n1860__));
  and1  g0919(.dina(new_new_n6538__), .dinb(new_new_n6534__), .dout(new_new_n1861__));
  or1   g0920(.dina(new_new_n6540__), .dinb(new_new_n6536__), .dout(new_new_n1862__));
  and1  g0921(.dina(new_new_n6538__), .dinb(new_new_n6533__), .dout(new_new_n1863__));
  or1   g0922(.dina(new_new_n6540__), .dinb(new_new_n6535__), .dout(new_new_n1864__));
  and1  g0923(.dina(new_new_n1864__), .dinb(new_new_n1862__), .dout(new_new_n1865__));
  or1   g0924(.dina(new_new_n1863__), .dinb(new_new_n1861__), .dout(new_new_n1866__));
  and1  g0925(.dina(new_new_n1821__), .dinb(new_new_n6491__), .dout(new_new_n1867__));
  or1   g0926(.dina(new_new_n6497__), .dinb(new_new_n6493__), .dout(new_new_n1868__));
  and1  g0927(.dina(new_new_n1868__), .dinb(new_new_n1866__), .dout(new_new_n1869__));
  or1   g0928(.dina(new_new_n6541__), .dinb(new_new_n6542__), .dout(new_new_n1870__));
  or1   g0929(.dina(new_new_n6544__), .dinb(new_new_n6542__), .dout(new_new_n1871__));
  or1   g0930(.dina(new_new_n6544__), .dinb(new_new_n6541__), .dout(new_new_n1872__));
  and1  g0931(.dina(new_new_n1872__), .dinb(new_new_n1871__), .dout(new_new_n1873__));
  and1  g0932(.dina(new_new_n6545__), .dinb(new_new_n6546__), .dout(new_new_n1874__));
  or1   g0933(.dina(new_new_n6547__), .dinb(new_new_n6548__), .dout(new_new_n1875__));
  and1  g0934(.dina(new_new_n6550__), .dinb(new_new_n6545__), .dout(new_new_n1876__));
  or1   g0935(.dina(new_new_n6552__), .dinb(new_new_n6547__), .dout(new_new_n1877__));
  and1  g0936(.dina(new_new_n6550__), .dinb(new_new_n6546__), .dout(new_new_n1878__));
  or1   g0937(.dina(new_new_n6552__), .dinb(new_new_n6548__), .dout(new_new_n1879__));
  and1  g0938(.dina(new_new_n1879__), .dinb(new_new_n1877__), .dout(new_new_n1880__));
  or1   g0939(.dina(new_new_n1878__), .dinb(new_new_n1876__), .dout(new_new_n1881__));
  and1  g0940(.dina(new_new_n6501__), .dinb(new_new_n6553__), .dout(new_new_n1882__));
  or1   g0941(.dina(new_new_n6506__), .dinb(new_new_n6554__), .dout(new_new_n1883__));
  and1  g0942(.dina(new_new_n6555__), .dinb(new_new_n6556__), .dout(new_new_n1884__));
  or1   g0943(.dina(new_new_n6557__), .dinb(new_new_n6558__), .dout(new_new_n1885__));
  and1  g0944(.dina(new_new_n6560__), .dinb(new_new_n6556__), .dout(new_new_n1886__));
  or1   g0945(.dina(new_new_n6562__), .dinb(new_new_n6558__), .dout(new_new_n1887__));
  and1  g0946(.dina(new_new_n6560__), .dinb(new_new_n6555__), .dout(new_new_n1888__));
  or1   g0947(.dina(new_new_n6562__), .dinb(new_new_n6557__), .dout(new_new_n1889__));
  and1  g0948(.dina(new_new_n1889__), .dinb(new_new_n1887__), .dout(new_new_n1890__));
  or1   g0949(.dina(new_new_n1888__), .dinb(new_new_n1886__), .dout(new_new_n1891__));
  and1  g0950(.dina(new_new_n6513__), .dinb(new_new_n1277__), .dout(new_new_n1892__));
  or1   g0951(.dina(new_new_n6515__), .dinb(new_new_n1278__), .dout(new_new_n1893__));
  and1  g0952(.dina(new_new_n6563__), .dinb(new_new_n6564__), .dout(new_new_n1894__));
  or1   g0953(.dina(new_new_n6565__), .dinb(new_new_n6566__), .dout(new_new_n1895__));
  and1  g0954(.dina(new_new_n6568__), .dinb(new_new_n6564__), .dout(new_new_n1896__));
  or1   g0955(.dina(new_new_n6570__), .dinb(new_new_n6566__), .dout(new_new_n1897__));
  and1  g0956(.dina(new_new_n6568__), .dinb(new_new_n6563__), .dout(new_new_n1898__));
  or1   g0957(.dina(new_new_n6570__), .dinb(new_new_n6565__), .dout(new_new_n1899__));
  and1  g0958(.dina(new_new_n1899__), .dinb(new_new_n1897__), .dout(new_new_n1900__));
  or1   g0959(.dina(new_new_n1898__), .dinb(new_new_n1896__), .dout(new_new_n1901__));
  and1  g0960(.dina(new_new_n6407__), .dinb(new_new_n6503__), .dout(new_new_n1902__));
  or1   g0961(.dina(new_new_n6415__), .dinb(new_new_n6508__), .dout(new_new_n1903__));
  and1  g0962(.dina(new_new_n6571__), .dinb(new_new_n6572__), .dout(new_new_n1904__));
  or1   g0963(.dina(new_new_n6573__), .dinb(new_new_n6574__), .dout(new_new_n1905__));
  and1  g0964(.dina(new_new_n6576__), .dinb(new_new_n6572__), .dout(new_new_n1906__));
  or1   g0965(.dina(new_new_n6578__), .dinb(new_new_n6574__), .dout(new_new_n1907__));
  and1  g0966(.dina(new_new_n6576__), .dinb(new_new_n6571__), .dout(new_new_n1908__));
  or1   g0967(.dina(new_new_n6578__), .dinb(new_new_n6573__), .dout(new_new_n1909__));
  and1  g0968(.dina(new_new_n1909__), .dinb(new_new_n1907__), .dout(new_new_n1910__));
  or1   g0969(.dina(new_new_n1908__), .dinb(new_new_n1906__), .dout(new_new_n1911__));
  and1  g0970(.dina(new_new_n6529__), .dinb(new_new_n6521__), .dout(new_new_n1912__));
  or1   g0971(.dina(new_new_n6531__), .dinb(new_new_n6523__), .dout(new_new_n1913__));
  and1  g0972(.dina(new_new_n6579__), .dinb(new_new_n6580__), .dout(new_new_n1914__));
  or1   g0973(.dina(new_new_n6581__), .dinb(new_new_n6582__), .dout(new_new_n1915__));
  and1  g0974(.dina(new_new_n6584__), .dinb(new_new_n6580__), .dout(new_new_n1916__));
  or1   g0975(.dina(new_new_n6586__), .dinb(new_new_n6582__), .dout(new_new_n1917__));
  and1  g0976(.dina(new_new_n6584__), .dinb(new_new_n6579__), .dout(new_new_n1918__));
  or1   g0977(.dina(new_new_n6586__), .dinb(new_new_n6581__), .dout(new_new_n1919__));
  and1  g0978(.dina(new_new_n1919__), .dinb(new_new_n1917__), .dout(new_new_n1920__));
  or1   g0979(.dina(new_new_n1918__), .dinb(new_new_n1916__), .dout(new_new_n1921__));
  and1  g0980(.dina(new_new_n1870__), .dinb(new_new_n6537__), .dout(new_new_n1922__));
  or1   g0981(.dina(new_new_n6543__), .dinb(new_new_n6539__), .dout(new_new_n1923__));
  and1  g0982(.dina(new_new_n1923__), .dinb(new_new_n1921__), .dout(new_new_n1924__));
  or1   g0983(.dina(new_new_n6587__), .dinb(new_new_n6588__), .dout(new_new_n1925__));
  or1   g0984(.dina(new_new_n6590__), .dinb(new_new_n6588__), .dout(new_new_n1926__));
  or1   g0985(.dina(new_new_n6590__), .dinb(new_new_n6587__), .dout(new_new_n1927__));
  and1  g0986(.dina(new_new_n1927__), .dinb(new_new_n1926__), .dout(new_new_n1928__));
  and1  g0987(.dina(new_new_n6592__), .dinb(new_new_n1283__), .dout(new_new_n1929__));
  or1   g0988(.dina(new_new_n6594__), .dinb(new_new_n1284__), .dout(new_new_n1930__));
  and1  g0989(.dina(new_new_n6592__), .dinb(new_new_n1274__), .dout(new_new_n1931__));
  or1   g0990(.dina(new_new_n6594__), .dinb(new_new_n1273__), .dout(new_new_n1932__));
  and1  g0991(.dina(new_new_n1932__), .dinb(new_new_n1930__), .dout(new_new_n1933__));
  or1   g0992(.dina(new_new_n1931__), .dinb(new_new_n1929__), .dout(new_new_n1934__));
  and1  g0993(.dina(new_new_n1240__), .dinb(new_new_n1173__), .dout(new_new_n1935__));
  or1   g0994(.dina(new_new_n1239__), .dinb(new_new_n1174__), .dout(new_new_n1936__));
  and1  g0995(.dina(new_new_n6595__), .dinb(new_new_n6596__), .dout(new_new_n1937__));
  or1   g0996(.dina(new_new_n6597__), .dinb(new_new_n6598__), .dout(new_new_n1938__));
  and1  g0997(.dina(new_new_n6600__), .dinb(new_new_n6596__), .dout(new_new_n1939__));
  or1   g0998(.dina(new_new_n6602__), .dinb(new_new_n6598__), .dout(new_new_n1940__));
  and1  g0999(.dina(new_new_n6600__), .dinb(new_new_n6595__), .dout(new_new_n1941__));
  or1   g1000(.dina(new_new_n6602__), .dinb(new_new_n6597__), .dout(new_new_n1942__));
  and1  g1001(.dina(new_new_n1942__), .dinb(new_new_n1940__), .dout(new_new_n1943__));
  or1   g1002(.dina(new_new_n1941__), .dinb(new_new_n1939__), .dout(new_new_n1944__));
  and1  g1003(.dina(new_new_n6500__), .dinb(new_new_n6603__), .dout(new_new_n1945__));
  or1   g1004(.dina(new_new_n6505__), .dinb(new_new_n6604__), .dout(new_new_n1946__));
  and1  g1005(.dina(new_new_n6605__), .dinb(new_new_n6606__), .dout(new_new_n1947__));
  or1   g1006(.dina(new_new_n6607__), .dinb(new_new_n6608__), .dout(new_new_n1948__));
  and1  g1007(.dina(new_new_n6610__), .dinb(new_new_n6606__), .dout(new_new_n1949__));
  or1   g1008(.dina(new_new_n6612__), .dinb(new_new_n6608__), .dout(new_new_n1950__));
  and1  g1009(.dina(new_new_n6610__), .dinb(new_new_n6605__), .dout(new_new_n1951__));
  or1   g1010(.dina(new_new_n6612__), .dinb(new_new_n6607__), .dout(new_new_n1952__));
  and1  g1011(.dina(new_new_n1952__), .dinb(new_new_n1950__), .dout(new_new_n1953__));
  or1   g1012(.dina(new_new_n1951__), .dinb(new_new_n1949__), .dout(new_new_n1954__));
  and1  g1013(.dina(new_new_n6559__), .dinb(new_new_n6549__), .dout(new_new_n1955__));
  or1   g1014(.dina(new_new_n6561__), .dinb(new_new_n6551__), .dout(new_new_n1956__));
  and1  g1015(.dina(new_new_n6613__), .dinb(new_new_n6614__), .dout(new_new_n1957__));
  or1   g1016(.dina(new_new_n6615__), .dinb(new_new_n6616__), .dout(new_new_n1958__));
  and1  g1017(.dina(new_new_n6618__), .dinb(new_new_n6614__), .dout(new_new_n1959__));
  or1   g1018(.dina(new_new_n6620__), .dinb(new_new_n6616__), .dout(new_new_n1960__));
  and1  g1019(.dina(new_new_n6618__), .dinb(new_new_n6613__), .dout(new_new_n1961__));
  or1   g1020(.dina(new_new_n6620__), .dinb(new_new_n6615__), .dout(new_new_n1962__));
  and1  g1021(.dina(new_new_n1962__), .dinb(new_new_n1960__), .dout(new_new_n1963__));
  or1   g1022(.dina(new_new_n1961__), .dinb(new_new_n1959__), .dout(new_new_n1964__));
  and1  g1023(.dina(new_new_n6409__), .dinb(new_new_n6553__), .dout(new_new_n1965__));
  or1   g1024(.dina(new_new_n6417__), .dinb(new_new_n6554__), .dout(new_new_n1966__));
  and1  g1025(.dina(new_new_n6621__), .dinb(new_new_n6622__), .dout(new_new_n1967__));
  or1   g1026(.dina(new_new_n6623__), .dinb(new_new_n6624__), .dout(new_new_n1968__));
  and1  g1027(.dina(new_new_n6626__), .dinb(new_new_n6622__), .dout(new_new_n1969__));
  or1   g1028(.dina(new_new_n6628__), .dinb(new_new_n6624__), .dout(new_new_n1970__));
  and1  g1029(.dina(new_new_n6626__), .dinb(new_new_n6621__), .dout(new_new_n1971__));
  or1   g1030(.dina(new_new_n6628__), .dinb(new_new_n6623__), .dout(new_new_n1972__));
  and1  g1031(.dina(new_new_n1972__), .dinb(new_new_n1970__), .dout(new_new_n1973__));
  or1   g1032(.dina(new_new_n1971__), .dinb(new_new_n1969__), .dout(new_new_n1974__));
  and1  g1033(.dina(new_new_n6575__), .dinb(new_new_n6567__), .dout(new_new_n1975__));
  or1   g1034(.dina(new_new_n6577__), .dinb(new_new_n6569__), .dout(new_new_n1976__));
  and1  g1035(.dina(new_new_n6629__), .dinb(new_new_n6630__), .dout(new_new_n1977__));
  or1   g1036(.dina(new_new_n6631__), .dinb(new_new_n6632__), .dout(new_new_n1978__));
  and1  g1037(.dina(new_new_n6634__), .dinb(new_new_n6630__), .dout(new_new_n1979__));
  or1   g1038(.dina(new_new_n6636__), .dinb(new_new_n6632__), .dout(new_new_n1980__));
  and1  g1039(.dina(new_new_n6634__), .dinb(new_new_n6629__), .dout(new_new_n1981__));
  or1   g1040(.dina(new_new_n6636__), .dinb(new_new_n6631__), .dout(new_new_n1982__));
  and1  g1041(.dina(new_new_n1982__), .dinb(new_new_n1980__), .dout(new_new_n1983__));
  or1   g1042(.dina(new_new_n1981__), .dinb(new_new_n1979__), .dout(new_new_n1984__));
  and1  g1043(.dina(new_new_n1925__), .dinb(new_new_n6583__), .dout(new_new_n1985__));
  or1   g1044(.dina(new_new_n6589__), .dinb(new_new_n6585__), .dout(new_new_n1986__));
  and1  g1045(.dina(new_new_n1986__), .dinb(new_new_n1984__), .dout(new_new_n1987__));
  or1   g1046(.dina(new_new_n6637__), .dinb(new_new_n6638__), .dout(new_new_n1988__));
  or1   g1047(.dina(new_new_n6640__), .dinb(new_new_n6638__), .dout(new_new_n1989__));
  or1   g1048(.dina(new_new_n6640__), .dinb(new_new_n6637__), .dout(new_new_n1990__));
  and1  g1049(.dina(new_new_n1990__), .dinb(new_new_n1989__), .dout(new_new_n1991__));
  and1  g1050(.dina(new_new_n925__), .dinb(new_new_n6642__), .dout(new_new_n1992__));
  or1   g1051(.dina(new_new_n926__), .dinb(new_new_n6644__), .dout(new_new_n1993__));
  and1  g1052(.dina(new_new_n6591__), .dinb(new_new_n1213__), .dout(new_new_n1994__));
  or1   g1053(.dina(new_new_n6593__), .dinb(new_new_n1214__), .dout(new_new_n1995__));
  and1  g1054(.dina(new_new_n6645__), .dinb(new_new_n6646__), .dout(new_new_n1996__));
  or1   g1055(.dina(new_new_n6647__), .dinb(new_new_n6648__), .dout(new_new_n1997__));
  and1  g1056(.dina(new_new_n6650__), .dinb(new_new_n6646__), .dout(new_new_n1998__));
  or1   g1057(.dina(new_new_n6652__), .dinb(new_new_n6648__), .dout(new_new_n1999__));
  and1  g1058(.dina(new_new_n6650__), .dinb(new_new_n6645__), .dout(new_new_n2000__));
  or1   g1059(.dina(new_new_n6652__), .dinb(new_new_n6647__), .dout(new_new_n2001__));
  and1  g1060(.dina(new_new_n2001__), .dinb(new_new_n1999__), .dout(new_new_n2002__));
  or1   g1061(.dina(new_new_n2000__), .dinb(new_new_n1998__), .dout(new_new_n2003__));
  and1  g1062(.dina(new_new_n6502__), .dinb(new_new_n6653__), .dout(new_new_n2004__));
  or1   g1063(.dina(new_new_n6507__), .dinb(new_new_n6654__), .dout(new_new_n2005__));
  and1  g1064(.dina(new_new_n6655__), .dinb(new_new_n6656__), .dout(new_new_n2006__));
  or1   g1065(.dina(new_new_n6657__), .dinb(new_new_n6658__), .dout(new_new_n2007__));
  and1  g1066(.dina(new_new_n6660__), .dinb(new_new_n6656__), .dout(new_new_n2008__));
  or1   g1067(.dina(new_new_n6662__), .dinb(new_new_n6658__), .dout(new_new_n2009__));
  and1  g1068(.dina(new_new_n6660__), .dinb(new_new_n6655__), .dout(new_new_n2010__));
  or1   g1069(.dina(new_new_n6662__), .dinb(new_new_n6657__), .dout(new_new_n2011__));
  and1  g1070(.dina(new_new_n2011__), .dinb(new_new_n2009__), .dout(new_new_n2012__));
  or1   g1071(.dina(new_new_n2010__), .dinb(new_new_n2008__), .dout(new_new_n2013__));
  and1  g1072(.dina(new_new_n6609__), .dinb(new_new_n6599__), .dout(new_new_n2014__));
  or1   g1073(.dina(new_new_n6611__), .dinb(new_new_n6601__), .dout(new_new_n2015__));
  and1  g1074(.dina(new_new_n6663__), .dinb(new_new_n6664__), .dout(new_new_n2016__));
  or1   g1075(.dina(new_new_n6665__), .dinb(new_new_n6666__), .dout(new_new_n2017__));
  and1  g1076(.dina(new_new_n6668__), .dinb(new_new_n6664__), .dout(new_new_n2018__));
  or1   g1077(.dina(new_new_n6670__), .dinb(new_new_n6666__), .dout(new_new_n2019__));
  and1  g1078(.dina(new_new_n6668__), .dinb(new_new_n6663__), .dout(new_new_n2020__));
  or1   g1079(.dina(new_new_n6670__), .dinb(new_new_n6665__), .dout(new_new_n2021__));
  and1  g1080(.dina(new_new_n2021__), .dinb(new_new_n2019__), .dout(new_new_n2022__));
  or1   g1081(.dina(new_new_n2020__), .dinb(new_new_n2018__), .dout(new_new_n2023__));
  and1  g1082(.dina(new_new_n6409__), .dinb(new_new_n6603__), .dout(new_new_n2024__));
  or1   g1083(.dina(new_new_n6417__), .dinb(new_new_n6604__), .dout(new_new_n2025__));
  and1  g1084(.dina(new_new_n6671__), .dinb(new_new_n6672__), .dout(new_new_n2026__));
  or1   g1085(.dina(new_new_n6673__), .dinb(new_new_n6674__), .dout(new_new_n2027__));
  and1  g1086(.dina(new_new_n6676__), .dinb(new_new_n6672__), .dout(new_new_n2028__));
  or1   g1087(.dina(new_new_n6678__), .dinb(new_new_n6674__), .dout(new_new_n2029__));
  and1  g1088(.dina(new_new_n6676__), .dinb(new_new_n6671__), .dout(new_new_n2030__));
  or1   g1089(.dina(new_new_n6678__), .dinb(new_new_n6673__), .dout(new_new_n2031__));
  and1  g1090(.dina(new_new_n2031__), .dinb(new_new_n2029__), .dout(new_new_n2032__));
  or1   g1091(.dina(new_new_n2030__), .dinb(new_new_n2028__), .dout(new_new_n2033__));
  and1  g1092(.dina(new_new_n6625__), .dinb(new_new_n6617__), .dout(new_new_n2034__));
  or1   g1093(.dina(new_new_n6627__), .dinb(new_new_n6619__), .dout(new_new_n2035__));
  and1  g1094(.dina(new_new_n6679__), .dinb(new_new_n6680__), .dout(new_new_n2036__));
  or1   g1095(.dina(new_new_n6681__), .dinb(new_new_n6682__), .dout(new_new_n2037__));
  and1  g1096(.dina(new_new_n6684__), .dinb(new_new_n6680__), .dout(new_new_n2038__));
  or1   g1097(.dina(new_new_n6686__), .dinb(new_new_n6682__), .dout(new_new_n2039__));
  and1  g1098(.dina(new_new_n6684__), .dinb(new_new_n6679__), .dout(new_new_n2040__));
  or1   g1099(.dina(new_new_n6686__), .dinb(new_new_n6681__), .dout(new_new_n2041__));
  and1  g1100(.dina(new_new_n2041__), .dinb(new_new_n2039__), .dout(new_new_n2042__));
  or1   g1101(.dina(new_new_n2040__), .dinb(new_new_n2038__), .dout(new_new_n2043__));
  and1  g1102(.dina(new_new_n1988__), .dinb(new_new_n6633__), .dout(new_new_n2044__));
  or1   g1103(.dina(new_new_n6639__), .dinb(new_new_n6635__), .dout(new_new_n2045__));
  and1  g1104(.dina(new_new_n2045__), .dinb(new_new_n2043__), .dout(new_new_n2046__));
  or1   g1105(.dina(new_new_n6687__), .dinb(new_new_n6688__), .dout(new_new_n2047__));
  or1   g1106(.dina(new_new_n6690__), .dinb(new_new_n6688__), .dout(new_new_n2048__));
  or1   g1107(.dina(new_new_n6690__), .dinb(new_new_n6687__), .dout(new_new_n2049__));
  and1  g1108(.dina(new_new_n2049__), .dinb(new_new_n2048__), .dout(new_new_n2050__));
  and1  g1109(.dina(new_new_n6502__), .dinb(new_new_n6642__), .dout(new_new_n2051__));
  or1   g1110(.dina(new_new_n6507__), .dinb(new_new_n6644__), .dout(new_new_n2052__));
  and1  g1111(.dina(new_new_n6659__), .dinb(new_new_n6649__), .dout(new_new_n2053__));
  or1   g1112(.dina(new_new_n6661__), .dinb(new_new_n6651__), .dout(new_new_n2054__));
  and1  g1113(.dina(new_new_n6691__), .dinb(new_new_n6692__), .dout(new_new_n2055__));
  or1   g1114(.dina(new_new_n6693__), .dinb(new_new_n6694__), .dout(new_new_n2056__));
  and1  g1115(.dina(new_new_n6696__), .dinb(new_new_n6692__), .dout(new_new_n2057__));
  or1   g1116(.dina(new_new_n6698__), .dinb(new_new_n6694__), .dout(new_new_n2058__));
  and1  g1117(.dina(new_new_n6696__), .dinb(new_new_n6691__), .dout(new_new_n2059__));
  or1   g1118(.dina(new_new_n6698__), .dinb(new_new_n6693__), .dout(new_new_n2060__));
  and1  g1119(.dina(new_new_n2060__), .dinb(new_new_n2058__), .dout(new_new_n2061__));
  or1   g1120(.dina(new_new_n2059__), .dinb(new_new_n2057__), .dout(new_new_n2062__));
  and1  g1121(.dina(new_new_n6410__), .dinb(new_new_n6653__), .dout(new_new_n2063__));
  or1   g1122(.dina(new_new_n6418__), .dinb(new_new_n6654__), .dout(new_new_n2064__));
  and1  g1123(.dina(new_new_n6699__), .dinb(new_new_n6700__), .dout(new_new_n2065__));
  or1   g1124(.dina(new_new_n6701__), .dinb(new_new_n6702__), .dout(new_new_n2066__));
  and1  g1125(.dina(new_new_n6704__), .dinb(new_new_n6700__), .dout(new_new_n2067__));
  or1   g1126(.dina(new_new_n6706__), .dinb(new_new_n6702__), .dout(new_new_n2068__));
  and1  g1127(.dina(new_new_n6704__), .dinb(new_new_n6699__), .dout(new_new_n2069__));
  or1   g1128(.dina(new_new_n6706__), .dinb(new_new_n6701__), .dout(new_new_n2070__));
  and1  g1129(.dina(new_new_n2070__), .dinb(new_new_n2068__), .dout(new_new_n2071__));
  or1   g1130(.dina(new_new_n2069__), .dinb(new_new_n2067__), .dout(new_new_n2072__));
  and1  g1131(.dina(new_new_n6675__), .dinb(new_new_n6667__), .dout(new_new_n2073__));
  or1   g1132(.dina(new_new_n6677__), .dinb(new_new_n6669__), .dout(new_new_n2074__));
  and1  g1133(.dina(new_new_n6707__), .dinb(new_new_n6708__), .dout(new_new_n2075__));
  or1   g1134(.dina(new_new_n6709__), .dinb(new_new_n6710__), .dout(new_new_n2076__));
  and1  g1135(.dina(new_new_n6712__), .dinb(new_new_n6708__), .dout(new_new_n2077__));
  or1   g1136(.dina(new_new_n6714__), .dinb(new_new_n6710__), .dout(new_new_n2078__));
  and1  g1137(.dina(new_new_n6712__), .dinb(new_new_n6707__), .dout(new_new_n2079__));
  or1   g1138(.dina(new_new_n6714__), .dinb(new_new_n6709__), .dout(new_new_n2080__));
  and1  g1139(.dina(new_new_n2080__), .dinb(new_new_n2078__), .dout(new_new_n2081__));
  or1   g1140(.dina(new_new_n2079__), .dinb(new_new_n2077__), .dout(new_new_n2082__));
  and1  g1141(.dina(new_new_n2047__), .dinb(new_new_n6683__), .dout(new_new_n2083__));
  or1   g1142(.dina(new_new_n6689__), .dinb(new_new_n6685__), .dout(new_new_n2084__));
  and1  g1143(.dina(new_new_n2084__), .dinb(new_new_n2082__), .dout(new_new_n2085__));
  or1   g1144(.dina(new_new_n6715__), .dinb(new_new_n6716__), .dout(new_new_n2086__));
  or1   g1145(.dina(new_new_n6718__), .dinb(new_new_n6716__), .dout(new_new_n2087__));
  or1   g1146(.dina(new_new_n6718__), .dinb(new_new_n6715__), .dout(new_new_n2088__));
  and1  g1147(.dina(new_new_n2088__), .dinb(new_new_n2087__), .dout(new_new_n2089__));
  and1  g1148(.dina(new_new_n6410__), .dinb(new_new_n6641__), .dout(new_new_n2090__));
  or1   g1149(.dina(new_new_n6418__), .dinb(new_new_n6643__), .dout(new_new_n2091__));
  and1  g1150(.dina(new_new_n6703__), .dinb(new_new_n6695__), .dout(new_new_n2092__));
  or1   g1151(.dina(new_new_n6705__), .dinb(new_new_n6697__), .dout(new_new_n2093__));
  and1  g1152(.dina(new_new_n6719__), .dinb(new_new_n6720__), .dout(new_new_n2094__));
  or1   g1153(.dina(new_new_n6721__), .dinb(new_new_n6722__), .dout(new_new_n2095__));
  and1  g1154(.dina(new_new_n6724__), .dinb(new_new_n6720__), .dout(new_new_n2096__));
  or1   g1155(.dina(new_new_n6725__), .dinb(new_new_n6722__), .dout(new_new_n2097__));
  and1  g1156(.dina(new_new_n6724__), .dinb(new_new_n6719__), .dout(new_new_n2098__));
  or1   g1157(.dina(new_new_n6725__), .dinb(new_new_n6721__), .dout(new_new_n2099__));
  and1  g1158(.dina(new_new_n2099__), .dinb(new_new_n2097__), .dout(new_new_n2100__));
  or1   g1159(.dina(new_new_n2098__), .dinb(new_new_n2096__), .dout(new_new_n2101__));
  and1  g1160(.dina(new_new_n2086__), .dinb(new_new_n6711__), .dout(new_new_n2102__));
  or1   g1161(.dina(new_new_n6717__), .dinb(new_new_n6713__), .dout(new_new_n2103__));
  or1   g1162(.dina(new_new_n2102__), .dinb(new_new_n2100__), .dout(new_new_n2104__));
  and1  g1163(.dina(new_new_n6727__), .dinb(new_new_n6723__), .dout(new_new_n2105__));
  and1  g1164(.dina(new_new_n6727__), .dinb(new_new_n2101__), .dout(new_new_n2106__));
  and1  g1165(.dina(new_new_n6726__), .dinb(new_new_n2103__), .dout(new_new_n2107__));
  or1   g1166(.dina(new_new_n2107__), .dinb(new_new_n2106__), .dout(new_new_n2108__));
  and1  g1167(.dina(new_new_n6731__), .dinb(new_new_n6740__), .dout(new_new_n2109__));
  or1   g1168(.dina(new_new_n6745__), .dinb(new_new_n6753__), .dout(new_new_n2110__));
  and1  g1169(.dina(new_new_n1438__), .dinb(new_new_n1432__), .dout(new_new_n2111__));
  or1   g1170(.dina(new_new_n1437__), .dinb(new_new_n1431__), .dout(new_new_n2112__));
  and1  g1171(.dina(new_new_n6755__), .dinb(new_new_n2110__), .dout(new_new_n2113__));
  or1   g1172(.dina(new_new_n2111__), .dinb(new_new_n6756__), .dout(new_new_n2114__));
  and1  g1173(.dina(new_new_n6740__), .dinb(new_new_n6760__), .dout(new_new_n2115__));
  or1   g1174(.dina(new_new_n6753__), .dinb(new_new_n6774__), .dout(new_new_n2116__));
  and1  g1175(.dina(new_new_n6785__), .dinb(new_new_n6786__), .dout(new_new_n2117__));
  or1   g1176(.dina(new_new_n6787__), .dinb(new_new_n6788__), .dout(new_new_n2118__));
  and1  g1177(.dina(new_new_n6790__), .dinb(new_new_n6785__), .dout(new_new_n2119__));
  or1   g1178(.dina(new_new_n6792__), .dinb(new_new_n6787__), .dout(new_new_n2120__));
  and1  g1179(.dina(new_new_n6790__), .dinb(new_new_n6786__), .dout(new_new_n2121__));
  or1   g1180(.dina(new_new_n6792__), .dinb(new_new_n6788__), .dout(new_new_n2122__));
  and1  g1181(.dina(new_new_n2122__), .dinb(new_new_n2120__), .dout(new_new_n2123__));
  or1   g1182(.dina(new_new_n2121__), .dinb(new_new_n2119__), .dout(new_new_n2124__));
  and1  g1183(.dina(new_new_n2114__), .dinb(new_new_n1375__), .dout(new_new_n2125__));
  or1   g1184(.dina(new_new_n6793__), .dinb(new_new_n1376__), .dout(new_new_n2126__));
  and1  g1185(.dina(new_new_n6794__), .dinb(new_new_n6795__), .dout(new_new_n2127__));
  or1   g1186(.dina(new_new_n6796__), .dinb(new_new_n6797__), .dout(new_new_n2128__));
  and1  g1187(.dina(new_new_n6799__), .dinb(new_new_n6795__), .dout(new_new_n2129__));
  or1   g1188(.dina(new_new_n6801__), .dinb(new_new_n6797__), .dout(new_new_n2130__));
  and1  g1189(.dina(new_new_n6799__), .dinb(new_new_n6794__), .dout(new_new_n2131__));
  or1   g1190(.dina(new_new_n6801__), .dinb(new_new_n6796__), .dout(new_new_n2132__));
  and1  g1191(.dina(new_new_n2132__), .dinb(new_new_n2130__), .dout(new_new_n2133__));
  or1   g1192(.dina(new_new_n2131__), .dinb(new_new_n2129__), .dout(new_new_n2134__));
  and1  g1193(.dina(new_new_n6802__), .dinb(new_new_n2116__), .dout(new_new_n2135__));
  or1   g1194(.dina(new_new_n2133__), .dinb(new_new_n6803__), .dout(new_new_n2136__));
  and1  g1195(.dina(new_new_n6739__), .dinb(new_new_n6807__), .dout(new_new_n2137__));
  or1   g1196(.dina(new_new_n6754__), .dinb(new_new_n6817__), .dout(new_new_n2138__));
  and1  g1197(.dina(new_new_n6825__), .dinb(new_new_n1383__), .dout(new_new_n2139__));
  or1   g1198(.dina(new_new_n6827__), .dinb(new_new_n1384__), .dout(new_new_n2140__));
  and1  g1199(.dina(new_new_n6825__), .dinb(new_new_n1336__), .dout(new_new_n2141__));
  or1   g1200(.dina(new_new_n6827__), .dinb(new_new_n1335__), .dout(new_new_n2142__));
  and1  g1201(.dina(new_new_n2142__), .dinb(new_new_n2140__), .dout(new_new_n2143__));
  or1   g1202(.dina(new_new_n2141__), .dinb(new_new_n2139__), .dout(new_new_n2144__));
  and1  g1203(.dina(new_new_n6789__), .dinb(new_new_n1311__), .dout(new_new_n2145__));
  or1   g1204(.dina(new_new_n6791__), .dinb(new_new_n1312__), .dout(new_new_n2146__));
  and1  g1205(.dina(new_new_n6828__), .dinb(new_new_n6829__), .dout(new_new_n2147__));
  or1   g1206(.dina(new_new_n6830__), .dinb(new_new_n6831__), .dout(new_new_n2148__));
  and1  g1207(.dina(new_new_n6833__), .dinb(new_new_n6829__), .dout(new_new_n2149__));
  or1   g1208(.dina(new_new_n6835__), .dinb(new_new_n6831__), .dout(new_new_n2150__));
  and1  g1209(.dina(new_new_n6833__), .dinb(new_new_n6828__), .dout(new_new_n2151__));
  or1   g1210(.dina(new_new_n6835__), .dinb(new_new_n6830__), .dout(new_new_n2152__));
  and1  g1211(.dina(new_new_n2152__), .dinb(new_new_n2150__), .dout(new_new_n2153__));
  or1   g1212(.dina(new_new_n2151__), .dinb(new_new_n2149__), .dout(new_new_n2154__));
  and1  g1213(.dina(new_new_n6837__), .dinb(new_new_n6760__), .dout(new_new_n2155__));
  or1   g1214(.dina(new_new_n6839__), .dinb(new_new_n6774__), .dout(new_new_n2156__));
  and1  g1215(.dina(new_new_n6840__), .dinb(new_new_n6841__), .dout(new_new_n2157__));
  or1   g1216(.dina(new_new_n6842__), .dinb(new_new_n6843__), .dout(new_new_n2158__));
  and1  g1217(.dina(new_new_n6845__), .dinb(new_new_n6841__), .dout(new_new_n2159__));
  or1   g1218(.dina(new_new_n6847__), .dinb(new_new_n6843__), .dout(new_new_n2160__));
  and1  g1219(.dina(new_new_n6845__), .dinb(new_new_n6840__), .dout(new_new_n2161__));
  or1   g1220(.dina(new_new_n6847__), .dinb(new_new_n6842__), .dout(new_new_n2162__));
  and1  g1221(.dina(new_new_n2162__), .dinb(new_new_n2160__), .dout(new_new_n2163__));
  or1   g1222(.dina(new_new_n2161__), .dinb(new_new_n2159__), .dout(new_new_n2164__));
  and1  g1223(.dina(new_new_n2136__), .dinb(new_new_n6798__), .dout(new_new_n2165__));
  or1   g1224(.dina(new_new_n6848__), .dinb(new_new_n6800__), .dout(new_new_n2166__));
  and1  g1225(.dina(new_new_n6849__), .dinb(new_new_n6850__), .dout(new_new_n2167__));
  or1   g1226(.dina(new_new_n6851__), .dinb(new_new_n6852__), .dout(new_new_n2168__));
  and1  g1227(.dina(new_new_n6854__), .dinb(new_new_n6850__), .dout(new_new_n2169__));
  or1   g1228(.dina(new_new_n6856__), .dinb(new_new_n6852__), .dout(new_new_n2170__));
  and1  g1229(.dina(new_new_n6854__), .dinb(new_new_n6849__), .dout(new_new_n2171__));
  or1   g1230(.dina(new_new_n6856__), .dinb(new_new_n6851__), .dout(new_new_n2172__));
  and1  g1231(.dina(new_new_n2172__), .dinb(new_new_n2170__), .dout(new_new_n2173__));
  or1   g1232(.dina(new_new_n2171__), .dinb(new_new_n2169__), .dout(new_new_n2174__));
  and1  g1233(.dina(new_new_n6857__), .dinb(new_new_n2138__), .dout(new_new_n2175__));
  or1   g1234(.dina(new_new_n2173__), .dinb(new_new_n6858__), .dout(new_new_n2176__));
  and1  g1235(.dina(new_new_n6861__), .dinb(new_new_n6865__), .dout(new_new_n2177__));
  or1   g1236(.dina(new_new_n6870__), .dinb(new_new_n6874__), .dout(new_new_n2178__));
  and1  g1237(.dina(new_new_n6877__), .dinb(new_new_n1474__), .dout(new_new_n2179__));
  or1   g1238(.dina(new_new_n6879__), .dinb(new_new_n1473__), .dout(new_new_n2180__));
  and1  g1239(.dina(new_new_n6877__), .dinb(new_new_n1418__), .dout(new_new_n2181__));
  or1   g1240(.dina(new_new_n6879__), .dinb(new_new_n1417__), .dout(new_new_n2182__));
  and1  g1241(.dina(new_new_n2182__), .dinb(new_new_n2180__), .dout(new_new_n2183__));
  or1   g1242(.dina(new_new_n2181__), .dinb(new_new_n2179__), .dout(new_new_n2184__));
  and1  g1243(.dina(new_new_n6880__), .dinb(new_new_n2178__), .dout(new_new_n2185__));
  or1   g1244(.dina(new_new_n2183__), .dinb(new_new_n6881__), .dout(new_new_n2186__));
  and1  g1245(.dina(new_new_n6741__), .dinb(new_new_n6884__), .dout(new_new_n2187__));
  or1   g1246(.dina(new_new_n6754__), .dinb(new_new_n6890__), .dout(new_new_n2188__));
  and1  g1247(.dina(new_new_n1440__), .dinb(new_new_n1423__), .dout(new_new_n2189__));
  or1   g1248(.dina(new_new_n1439__), .dinb(new_new_n1424__), .dout(new_new_n2190__));
  and1  g1249(.dina(new_new_n6824__), .dinb(new_new_n1299__), .dout(new_new_n2191__));
  or1   g1250(.dina(new_new_n6826__), .dinb(new_new_n1300__), .dout(new_new_n2192__));
  and1  g1251(.dina(new_new_n6894__), .dinb(new_new_n6895__), .dout(new_new_n2193__));
  or1   g1252(.dina(new_new_n6896__), .dinb(new_new_n6897__), .dout(new_new_n2194__));
  and1  g1253(.dina(new_new_n6899__), .dinb(new_new_n6895__), .dout(new_new_n2195__));
  or1   g1254(.dina(new_new_n6901__), .dinb(new_new_n6897__), .dout(new_new_n2196__));
  and1  g1255(.dina(new_new_n6899__), .dinb(new_new_n6894__), .dout(new_new_n2197__));
  or1   g1256(.dina(new_new_n6901__), .dinb(new_new_n6896__), .dout(new_new_n2198__));
  and1  g1257(.dina(new_new_n2198__), .dinb(new_new_n2196__), .dout(new_new_n2199__));
  or1   g1258(.dina(new_new_n2197__), .dinb(new_new_n2195__), .dout(new_new_n2200__));
  and1  g1259(.dina(new_new_n6903__), .dinb(new_new_n6761__), .dout(new_new_n2201__));
  or1   g1260(.dina(new_new_n6905__), .dinb(new_new_n6775__), .dout(new_new_n2202__));
  and1  g1261(.dina(new_new_n6906__), .dinb(new_new_n6907__), .dout(new_new_n2203__));
  or1   g1262(.dina(new_new_n6908__), .dinb(new_new_n6909__), .dout(new_new_n2204__));
  and1  g1263(.dina(new_new_n6911__), .dinb(new_new_n6907__), .dout(new_new_n2205__));
  or1   g1264(.dina(new_new_n6913__), .dinb(new_new_n6909__), .dout(new_new_n2206__));
  and1  g1265(.dina(new_new_n6911__), .dinb(new_new_n6906__), .dout(new_new_n2207__));
  or1   g1266(.dina(new_new_n6913__), .dinb(new_new_n6908__), .dout(new_new_n2208__));
  and1  g1267(.dina(new_new_n2208__), .dinb(new_new_n2206__), .dout(new_new_n2209__));
  or1   g1268(.dina(new_new_n2207__), .dinb(new_new_n2205__), .dout(new_new_n2210__));
  and1  g1269(.dina(new_new_n6844__), .dinb(new_new_n6832__), .dout(new_new_n2211__));
  or1   g1270(.dina(new_new_n6846__), .dinb(new_new_n6834__), .dout(new_new_n2212__));
  and1  g1271(.dina(new_new_n6914__), .dinb(new_new_n6915__), .dout(new_new_n2213__));
  or1   g1272(.dina(new_new_n6916__), .dinb(new_new_n6917__), .dout(new_new_n2214__));
  and1  g1273(.dina(new_new_n6919__), .dinb(new_new_n6915__), .dout(new_new_n2215__));
  or1   g1274(.dina(new_new_n6921__), .dinb(new_new_n6917__), .dout(new_new_n2216__));
  and1  g1275(.dina(new_new_n6919__), .dinb(new_new_n6914__), .dout(new_new_n2217__));
  or1   g1276(.dina(new_new_n6921__), .dinb(new_new_n6916__), .dout(new_new_n2218__));
  and1  g1277(.dina(new_new_n2218__), .dinb(new_new_n2216__), .dout(new_new_n2219__));
  or1   g1278(.dina(new_new_n2217__), .dinb(new_new_n2215__), .dout(new_new_n2220__));
  and1  g1279(.dina(new_new_n6837__), .dinb(new_new_n6807__), .dout(new_new_n2221__));
  or1   g1280(.dina(new_new_n6839__), .dinb(new_new_n6817__), .dout(new_new_n2222__));
  and1  g1281(.dina(new_new_n6922__), .dinb(new_new_n6923__), .dout(new_new_n2223__));
  or1   g1282(.dina(new_new_n6924__), .dinb(new_new_n6925__), .dout(new_new_n2224__));
  and1  g1283(.dina(new_new_n6927__), .dinb(new_new_n6923__), .dout(new_new_n2225__));
  or1   g1284(.dina(new_new_n6929__), .dinb(new_new_n6925__), .dout(new_new_n2226__));
  and1  g1285(.dina(new_new_n6927__), .dinb(new_new_n6922__), .dout(new_new_n2227__));
  or1   g1286(.dina(new_new_n6929__), .dinb(new_new_n6924__), .dout(new_new_n2228__));
  and1  g1287(.dina(new_new_n2228__), .dinb(new_new_n2226__), .dout(new_new_n2229__));
  or1   g1288(.dina(new_new_n2227__), .dinb(new_new_n2225__), .dout(new_new_n2230__));
  and1  g1289(.dina(new_new_n2176__), .dinb(new_new_n6853__), .dout(new_new_n2231__));
  or1   g1290(.dina(new_new_n6930__), .dinb(new_new_n6855__), .dout(new_new_n2232__));
  and1  g1291(.dina(new_new_n6931__), .dinb(new_new_n6932__), .dout(new_new_n2233__));
  or1   g1292(.dina(new_new_n6933__), .dinb(new_new_n6934__), .dout(new_new_n2234__));
  and1  g1293(.dina(new_new_n6936__), .dinb(new_new_n6932__), .dout(new_new_n2235__));
  or1   g1294(.dina(new_new_n6938__), .dinb(new_new_n6934__), .dout(new_new_n2236__));
  and1  g1295(.dina(new_new_n6936__), .dinb(new_new_n6931__), .dout(new_new_n2237__));
  or1   g1296(.dina(new_new_n6938__), .dinb(new_new_n6933__), .dout(new_new_n2238__));
  and1  g1297(.dina(new_new_n2238__), .dinb(new_new_n2236__), .dout(new_new_n2239__));
  or1   g1298(.dina(new_new_n2237__), .dinb(new_new_n2235__), .dout(new_new_n2240__));
  and1  g1299(.dina(new_new_n6942__), .dinb(new_new_n6865__), .dout(new_new_n2241__));
  or1   g1300(.dina(new_new_n6955__), .dinb(new_new_n6874__), .dout(new_new_n2242__));
  and1  g1301(.dina(new_new_n6965__), .dinb(new_new_n2188__), .dout(new_new_n2243__));
  or1   g1302(.dina(new_new_n2239__), .dinb(new_new_n6966__), .dout(new_new_n2244__));
  and1  g1303(.dina(new_new_n1522__), .dinb(new_new_n1512__), .dout(new_new_n2245__));
  or1   g1304(.dina(new_new_n1521__), .dinb(new_new_n1511__), .dout(new_new_n2246__));
  and1  g1305(.dina(new_new_n6861__), .dinb(new_new_n6969__), .dout(new_new_n2247__));
  or1   g1306(.dina(new_new_n6870__), .dinb(new_new_n6975__), .dout(new_new_n2248__));
  and1  g1307(.dina(new_new_n6977__), .dinb(new_new_n6978__), .dout(new_new_n2249__));
  or1   g1308(.dina(new_new_n6979__), .dinb(new_new_n6980__), .dout(new_new_n2250__));
  and1  g1309(.dina(new_new_n6982__), .dinb(new_new_n6978__), .dout(new_new_n2251__));
  or1   g1310(.dina(new_new_n6984__), .dinb(new_new_n6980__), .dout(new_new_n2252__));
  and1  g1311(.dina(new_new_n6982__), .dinb(new_new_n6977__), .dout(new_new_n2253__));
  or1   g1312(.dina(new_new_n6984__), .dinb(new_new_n6979__), .dout(new_new_n2254__));
  and1  g1313(.dina(new_new_n2254__), .dinb(new_new_n2252__), .dout(new_new_n2255__));
  or1   g1314(.dina(new_new_n2253__), .dinb(new_new_n2251__), .dout(new_new_n2256__));
  and1  g1315(.dina(new_new_n2186__), .dinb(new_new_n6876__), .dout(new_new_n2257__));
  or1   g1316(.dina(new_new_n6985__), .dinb(new_new_n6878__), .dout(new_new_n2258__));
  and1  g1317(.dina(new_new_n6986__), .dinb(new_new_n6987__), .dout(new_new_n2259__));
  or1   g1318(.dina(new_new_n6988__), .dinb(new_new_n6989__), .dout(new_new_n2260__));
  and1  g1319(.dina(new_new_n6991__), .dinb(new_new_n6987__), .dout(new_new_n2261__));
  or1   g1320(.dina(new_new_n6993__), .dinb(new_new_n6989__), .dout(new_new_n2262__));
  and1  g1321(.dina(new_new_n6991__), .dinb(new_new_n6986__), .dout(new_new_n2263__));
  or1   g1322(.dina(new_new_n6993__), .dinb(new_new_n6988__), .dout(new_new_n2264__));
  and1  g1323(.dina(new_new_n2264__), .dinb(new_new_n2262__), .dout(new_new_n2265__));
  or1   g1324(.dina(new_new_n2263__), .dinb(new_new_n2261__), .dout(new_new_n2266__));
  and1  g1325(.dina(new_new_n6994__), .dinb(new_new_n2242__), .dout(new_new_n2267__));
  or1   g1326(.dina(new_new_n2265__), .dinb(new_new_n6995__), .dout(new_new_n2268__));
  and1  g1327(.dina(new_new_n6998__), .dinb(new_new_n7001__), .dout(new_new_n2269__));
  or1   g1328(.dina(new_new_n7004__), .dinb(new_new_n7007__), .dout(new_new_n2270__));
  and1  g1329(.dina(new_new_n7008__), .dinb(new_new_n7009__), .dout(new_new_n2271__));
  or1   g1330(.dina(new_new_n7010__), .dinb(new_new_n7011__), .dout(new_new_n2272__));
  and1  g1331(.dina(new_new_n7013__), .dinb(new_new_n7008__), .dout(new_new_n2273__));
  or1   g1332(.dina(new_new_n7015__), .dinb(new_new_n7010__), .dout(new_new_n2274__));
  and1  g1333(.dina(new_new_n7013__), .dinb(new_new_n7009__), .dout(new_new_n2275__));
  or1   g1334(.dina(new_new_n7015__), .dinb(new_new_n7011__), .dout(new_new_n2276__));
  and1  g1335(.dina(new_new_n2276__), .dinb(new_new_n2274__), .dout(new_new_n2277__));
  or1   g1336(.dina(new_new_n2275__), .dinb(new_new_n2273__), .dout(new_new_n2278__));
  and1  g1337(.dina(new_new_n6866__), .dinb(new_new_n7019__), .dout(new_new_n2279__));
  or1   g1338(.dina(new_new_n6873__), .dinb(new_new_n7034__), .dout(new_new_n2280__));
  and1  g1339(.dina(new_new_n7046__), .dinb(new_new_n2270__), .dout(new_new_n2281__));
  or1   g1340(.dina(new_new_n2277__), .dinb(new_new_n7047__), .dout(new_new_n2282__));
  and1  g1341(.dina(new_new_n7048__), .dinb(new_new_n7049__), .dout(new_new_n2283__));
  or1   g1342(.dina(new_new_n7050__), .dinb(new_new_n7051__), .dout(new_new_n2284__));
  and1  g1343(.dina(new_new_n7053__), .dinb(new_new_n7048__), .dout(new_new_n2285__));
  or1   g1344(.dina(new_new_n7055__), .dinb(new_new_n7050__), .dout(new_new_n2286__));
  and1  g1345(.dina(new_new_n7053__), .dinb(new_new_n7049__), .dout(new_new_n2287__));
  or1   g1346(.dina(new_new_n7055__), .dinb(new_new_n7051__), .dout(new_new_n2288__));
  and1  g1347(.dina(new_new_n2288__), .dinb(new_new_n2286__), .dout(new_new_n2289__));
  or1   g1348(.dina(new_new_n2287__), .dinb(new_new_n2285__), .dout(new_new_n2290__));
  and1  g1349(.dina(new_new_n6981__), .dinb(new_new_n1455__), .dout(new_new_n2291__));
  or1   g1350(.dina(new_new_n6983__), .dinb(new_new_n1456__), .dout(new_new_n2292__));
  and1  g1351(.dina(new_new_n7056__), .dinb(new_new_n7057__), .dout(new_new_n2293__));
  or1   g1352(.dina(new_new_n7058__), .dinb(new_new_n7059__), .dout(new_new_n2294__));
  and1  g1353(.dina(new_new_n7061__), .dinb(new_new_n7057__), .dout(new_new_n2295__));
  or1   g1354(.dina(new_new_n7063__), .dinb(new_new_n7059__), .dout(new_new_n2296__));
  and1  g1355(.dina(new_new_n7061__), .dinb(new_new_n7056__), .dout(new_new_n2297__));
  or1   g1356(.dina(new_new_n7063__), .dinb(new_new_n7058__), .dout(new_new_n2298__));
  and1  g1357(.dina(new_new_n2298__), .dinb(new_new_n2296__), .dout(new_new_n2299__));
  or1   g1358(.dina(new_new_n2297__), .dinb(new_new_n2295__), .dout(new_new_n2300__));
  and1  g1359(.dina(new_new_n6942__), .dinb(new_new_n6969__), .dout(new_new_n2301__));
  or1   g1360(.dina(new_new_n6955__), .dinb(new_new_n6975__), .dout(new_new_n2302__));
  and1  g1361(.dina(new_new_n7064__), .dinb(new_new_n7065__), .dout(new_new_n2303__));
  or1   g1362(.dina(new_new_n7066__), .dinb(new_new_n7067__), .dout(new_new_n2304__));
  and1  g1363(.dina(new_new_n7069__), .dinb(new_new_n7065__), .dout(new_new_n2305__));
  or1   g1364(.dina(new_new_n7071__), .dinb(new_new_n7067__), .dout(new_new_n2306__));
  and1  g1365(.dina(new_new_n7069__), .dinb(new_new_n7064__), .dout(new_new_n2307__));
  or1   g1366(.dina(new_new_n7071__), .dinb(new_new_n7066__), .dout(new_new_n2308__));
  and1  g1367(.dina(new_new_n2308__), .dinb(new_new_n2306__), .dout(new_new_n2309__));
  or1   g1368(.dina(new_new_n2307__), .dinb(new_new_n2305__), .dout(new_new_n2310__));
  and1  g1369(.dina(new_new_n2268__), .dinb(new_new_n6990__), .dout(new_new_n2311__));
  or1   g1370(.dina(new_new_n7072__), .dinb(new_new_n6992__), .dout(new_new_n2312__));
  and1  g1371(.dina(new_new_n7073__), .dinb(new_new_n7074__), .dout(new_new_n2313__));
  or1   g1372(.dina(new_new_n7075__), .dinb(new_new_n7076__), .dout(new_new_n2314__));
  and1  g1373(.dina(new_new_n7078__), .dinb(new_new_n7074__), .dout(new_new_n2315__));
  or1   g1374(.dina(new_new_n7080__), .dinb(new_new_n7076__), .dout(new_new_n2316__));
  and1  g1375(.dina(new_new_n7078__), .dinb(new_new_n7073__), .dout(new_new_n2317__));
  or1   g1376(.dina(new_new_n7080__), .dinb(new_new_n7075__), .dout(new_new_n2318__));
  and1  g1377(.dina(new_new_n2318__), .dinb(new_new_n2316__), .dout(new_new_n2319__));
  or1   g1378(.dina(new_new_n2317__), .dinb(new_new_n2315__), .dout(new_new_n2320__));
  and1  g1379(.dina(new_new_n7081__), .dinb(new_new_n2280__), .dout(new_new_n2321__));
  or1   g1380(.dina(new_new_n2319__), .dinb(new_new_n7082__), .dout(new_new_n2322__));
  and1  g1381(.dina(new_new_n6998__), .dinb(new_new_n7086__), .dout(new_new_n2323__));
  or1   g1382(.dina(new_new_n7004__), .dinb(new_new_n7094__), .dout(new_new_n2324__));
  and1  g1383(.dina(new_new_n7100__), .dinb(new_new_n1554__), .dout(new_new_n2325__));
  or1   g1384(.dina(new_new_n7102__), .dinb(new_new_n1553__), .dout(new_new_n2326__));
  and1  g1385(.dina(new_new_n7100__), .dinb(new_new_n1500__), .dout(new_new_n2327__));
  or1   g1386(.dina(new_new_n7102__), .dinb(new_new_n1499__), .dout(new_new_n2328__));
  and1  g1387(.dina(new_new_n2328__), .dinb(new_new_n2326__), .dout(new_new_n2329__));
  or1   g1388(.dina(new_new_n2327__), .dinb(new_new_n2325__), .dout(new_new_n2330__));
  and1  g1389(.dina(new_new_n7105__), .dinb(new_new_n7001__), .dout(new_new_n2331__));
  or1   g1390(.dina(new_new_n7110__), .dinb(new_new_n7007__), .dout(new_new_n2332__));
  and1  g1391(.dina(new_new_n7112__), .dinb(new_new_n7113__), .dout(new_new_n2333__));
  or1   g1392(.dina(new_new_n7114__), .dinb(new_new_n7115__), .dout(new_new_n2334__));
  and1  g1393(.dina(new_new_n7117__), .dinb(new_new_n7113__), .dout(new_new_n2335__));
  or1   g1394(.dina(new_new_n7119__), .dinb(new_new_n7115__), .dout(new_new_n2336__));
  and1  g1395(.dina(new_new_n7117__), .dinb(new_new_n7112__), .dout(new_new_n2337__));
  or1   g1396(.dina(new_new_n7119__), .dinb(new_new_n7114__), .dout(new_new_n2338__));
  and1  g1397(.dina(new_new_n2338__), .dinb(new_new_n2336__), .dout(new_new_n2339__));
  or1   g1398(.dina(new_new_n2337__), .dinb(new_new_n2335__), .dout(new_new_n2340__));
  and1  g1399(.dina(new_new_n2282__), .dinb(new_new_n7012__), .dout(new_new_n2341__));
  or1   g1400(.dina(new_new_n7120__), .dinb(new_new_n7014__), .dout(new_new_n2342__));
  and1  g1401(.dina(new_new_n7121__), .dinb(new_new_n7122__), .dout(new_new_n2343__));
  or1   g1402(.dina(new_new_n7123__), .dinb(new_new_n7124__), .dout(new_new_n2344__));
  and1  g1403(.dina(new_new_n7126__), .dinb(new_new_n7122__), .dout(new_new_n2345__));
  or1   g1404(.dina(new_new_n7128__), .dinb(new_new_n7124__), .dout(new_new_n2346__));
  and1  g1405(.dina(new_new_n7126__), .dinb(new_new_n7121__), .dout(new_new_n2347__));
  or1   g1406(.dina(new_new_n7128__), .dinb(new_new_n7123__), .dout(new_new_n2348__));
  and1  g1407(.dina(new_new_n2348__), .dinb(new_new_n2346__), .dout(new_new_n2349__));
  or1   g1408(.dina(new_new_n2347__), .dinb(new_new_n2345__), .dout(new_new_n2350__));
  and1  g1409(.dina(new_new_n7131__), .dinb(new_new_n7135__), .dout(new_new_n2351__));
  or1   g1410(.dina(new_new_n7139__), .dinb(new_new_n7143__), .dout(new_new_n2352__));
  and1  g1411(.dina(new_new_n7144__), .dinb(new_new_n7135__), .dout(new_new_n2353__));
  or1   g1412(.dina(new_new_n7145__), .dinb(new_new_n7143__), .dout(new_new_n2354__));
  and1  g1413(.dina(new_new_n1426__), .dinb(new_new_n1422__), .dout(new_new_n2355__));
  or1   g1414(.dina(new_new_n1425__), .dinb(new_new_n1421__), .dout(new_new_n2356__));
  and1  g1415(.dina(new_new_n7144__), .dinb(new_new_n7147__), .dout(new_new_n2357__));
  or1   g1416(.dina(new_new_n7145__), .dinb(new_new_n7150__), .dout(new_new_n2358__));
  and1  g1417(.dina(new_new_n7152__), .dinb(new_new_n7153__), .dout(new_new_n2359__));
  or1   g1418(.dina(new_new_n7154__), .dinb(new_new_n7155__), .dout(new_new_n2360__));
  and1  g1419(.dina(new_new_n7157__), .dinb(new_new_n1369__), .dout(new_new_n2361__));
  or1   g1420(.dina(new_new_n7159__), .dinb(new_new_n1370__), .dout(new_new_n2362__));
  and1  g1421(.dina(new_new_n7160__), .dinb(new_new_n7161__), .dout(new_new_n2363__));
  or1   g1422(.dina(new_new_n7162__), .dinb(new_new_n7163__), .dout(new_new_n2364__));
  and1  g1423(.dina(new_new_n7165__), .dinb(new_new_n7161__), .dout(new_new_n2365__));
  or1   g1424(.dina(new_new_n7167__), .dinb(new_new_n7163__), .dout(new_new_n2366__));
  and1  g1425(.dina(new_new_n7165__), .dinb(new_new_n7160__), .dout(new_new_n2367__));
  or1   g1426(.dina(new_new_n7167__), .dinb(new_new_n7162__), .dout(new_new_n2368__));
  and1  g1427(.dina(new_new_n2368__), .dinb(new_new_n2366__), .dout(new_new_n2369__));
  or1   g1428(.dina(new_new_n2367__), .dinb(new_new_n2365__), .dout(new_new_n2370__));
  and1  g1429(.dina(new_new_n7131__), .dinb(new_new_n7147__), .dout(new_new_n2371__));
  or1   g1430(.dina(new_new_n7139__), .dinb(new_new_n7150__), .dout(new_new_n2372__));
  and1  g1431(.dina(new_new_n7168__), .dinb(new_new_n7169__), .dout(new_new_n2373__));
  or1   g1432(.dina(new_new_n7170__), .dinb(new_new_n7171__), .dout(new_new_n2374__));
  and1  g1433(.dina(new_new_n7173__), .dinb(new_new_n7164__), .dout(new_new_n2375__));
  or1   g1434(.dina(new_new_n7175__), .dinb(new_new_n7166__), .dout(new_new_n2376__));
  and1  g1435(.dina(new_new_n7176__), .dinb(new_new_n7177__), .dout(new_new_n2377__));
  or1   g1436(.dina(new_new_n7178__), .dinb(new_new_n7179__), .dout(new_new_n2378__));
  and1  g1437(.dina(new_new_n7181__), .dinb(new_new_n7177__), .dout(new_new_n2379__));
  or1   g1438(.dina(new_new_n7183__), .dinb(new_new_n7179__), .dout(new_new_n2380__));
  and1  g1439(.dina(new_new_n7181__), .dinb(new_new_n7176__), .dout(new_new_n2381__));
  or1   g1440(.dina(new_new_n7183__), .dinb(new_new_n7178__), .dout(new_new_n2382__));
  and1  g1441(.dina(new_new_n2382__), .dinb(new_new_n2380__), .dout(new_new_n2383__));
  or1   g1442(.dina(new_new_n2381__), .dinb(new_new_n2379__), .dout(new_new_n2384__));
  and1  g1443(.dina(new_new_n6731__), .dinb(new_new_n7148__), .dout(new_new_n2385__));
  or1   g1444(.dina(new_new_n6745__), .dinb(new_new_n7151__), .dout(new_new_n2386__));
  and1  g1445(.dina(new_new_n7184__), .dinb(new_new_n7185__), .dout(new_new_n2387__));
  or1   g1446(.dina(new_new_n7186__), .dinb(new_new_n7187__), .dout(new_new_n2388__));
  and1  g1447(.dina(new_new_n7189__), .dinb(new_new_n7185__), .dout(new_new_n2389__));
  or1   g1448(.dina(new_new_n7191__), .dinb(new_new_n7187__), .dout(new_new_n2390__));
  and1  g1449(.dina(new_new_n7189__), .dinb(new_new_n7184__), .dout(new_new_n2391__));
  or1   g1450(.dina(new_new_n7191__), .dinb(new_new_n7186__), .dout(new_new_n2392__));
  and1  g1451(.dina(new_new_n2392__), .dinb(new_new_n2390__), .dout(new_new_n2393__));
  or1   g1452(.dina(new_new_n2391__), .dinb(new_new_n2389__), .dout(new_new_n2394__));
  and1  g1453(.dina(new_new_n7173__), .dinb(new_new_n7169__), .dout(new_new_n2395__));
  or1   g1454(.dina(new_new_n7175__), .dinb(new_new_n7171__), .dout(new_new_n2396__));
  and1  g1455(.dina(new_new_n7172__), .dinb(new_new_n7168__), .dout(new_new_n2397__));
  or1   g1456(.dina(new_new_n7174__), .dinb(new_new_n7170__), .dout(new_new_n2398__));
  and1  g1457(.dina(new_new_n2398__), .dinb(new_new_n2396__), .dout(new_new_n2399__));
  or1   g1458(.dina(new_new_n2397__), .dinb(new_new_n2395__), .dout(new_new_n2400__));
  and1  g1459(.dina(new_new_n7157__), .dinb(new_new_n7153__), .dout(new_new_n2401__));
  or1   g1460(.dina(new_new_n7159__), .dinb(new_new_n7155__), .dout(new_new_n2402__));
  and1  g1461(.dina(new_new_n7156__), .dinb(new_new_n7152__), .dout(new_new_n2403__));
  or1   g1462(.dina(new_new_n7158__), .dinb(new_new_n7154__), .dout(new_new_n2404__));
  and1  g1463(.dina(new_new_n2404__), .dinb(new_new_n2402__), .dout(new_new_n2405__));
  or1   g1464(.dina(new_new_n2403__), .dinb(new_new_n2401__), .dout(new_new_n2406__));
  and1  g1465(.dina(new_new_n7193__), .dinb(new_new_n1293__), .dout(new_new_n2407__));
  or1   g1466(.dina(new_new_n7195__), .dinb(new_new_n1294__), .dout(new_new_n2408__));
  and1  g1467(.dina(new_new_n7196__), .dinb(new_new_n7197__), .dout(new_new_n2409__));
  or1   g1468(.dina(new_new_n7198__), .dinb(new_new_n7199__), .dout(new_new_n2410__));
  and1  g1469(.dina(new_new_n7201__), .dinb(new_new_n7197__), .dout(new_new_n2411__));
  or1   g1470(.dina(new_new_n7203__), .dinb(new_new_n7199__), .dout(new_new_n2412__));
  and1  g1471(.dina(new_new_n7201__), .dinb(new_new_n7196__), .dout(new_new_n2413__));
  or1   g1472(.dina(new_new_n7203__), .dinb(new_new_n7198__), .dout(new_new_n2414__));
  and1  g1473(.dina(new_new_n2414__), .dinb(new_new_n2412__), .dout(new_new_n2415__));
  or1   g1474(.dina(new_new_n2413__), .dinb(new_new_n2411__), .dout(new_new_n2416__));
  and1  g1475(.dina(new_new_n7132__), .dinb(new_new_n7205__), .dout(new_new_n2417__));
  or1   g1476(.dina(new_new_n7140__), .dinb(new_new_n7208__), .dout(new_new_n2418__));
  and1  g1477(.dina(new_new_n7209__), .dinb(new_new_n7210__), .dout(new_new_n2419__));
  or1   g1478(.dina(new_new_n7211__), .dinb(new_new_n7212__), .dout(new_new_n2420__));
  and1  g1479(.dina(new_new_n7214__), .dinb(new_new_n7200__), .dout(new_new_n2421__));
  or1   g1480(.dina(new_new_n7216__), .dinb(new_new_n7202__), .dout(new_new_n2422__));
  and1  g1481(.dina(new_new_n7217__), .dinb(new_new_n7218__), .dout(new_new_n2423__));
  or1   g1482(.dina(new_new_n7219__), .dinb(new_new_n7220__), .dout(new_new_n2424__));
  and1  g1483(.dina(new_new_n7222__), .dinb(new_new_n7218__), .dout(new_new_n2425__));
  or1   g1484(.dina(new_new_n7224__), .dinb(new_new_n7220__), .dout(new_new_n2426__));
  and1  g1485(.dina(new_new_n7222__), .dinb(new_new_n7217__), .dout(new_new_n2427__));
  or1   g1486(.dina(new_new_n7224__), .dinb(new_new_n7219__), .dout(new_new_n2428__));
  and1  g1487(.dina(new_new_n2428__), .dinb(new_new_n2426__), .dout(new_new_n2429__));
  or1   g1488(.dina(new_new_n2427__), .dinb(new_new_n2425__), .dout(new_new_n2430__));
  and1  g1489(.dina(new_new_n6732__), .dinb(new_new_n7205__), .dout(new_new_n2431__));
  or1   g1490(.dina(new_new_n6746__), .dinb(new_new_n7208__), .dout(new_new_n2432__));
  and1  g1491(.dina(new_new_n7225__), .dinb(new_new_n7226__), .dout(new_new_n2433__));
  or1   g1492(.dina(new_new_n7227__), .dinb(new_new_n7228__), .dout(new_new_n2434__));
  and1  g1493(.dina(new_new_n7230__), .dinb(new_new_n7221__), .dout(new_new_n2435__));
  or1   g1494(.dina(new_new_n7232__), .dinb(new_new_n7223__), .dout(new_new_n2436__));
  and1  g1495(.dina(new_new_n7233__), .dinb(new_new_n7234__), .dout(new_new_n2437__));
  or1   g1496(.dina(new_new_n7235__), .dinb(new_new_n7236__), .dout(new_new_n2438__));
  and1  g1497(.dina(new_new_n7193__), .dinb(new_new_n1377__), .dout(new_new_n2439__));
  or1   g1498(.dina(new_new_n7195__), .dinb(new_new_n1378__), .dout(new_new_n2440__));
  and1  g1499(.dina(new_new_n7192__), .dinb(new_new_n1330__), .dout(new_new_n2441__));
  or1   g1500(.dina(new_new_n7194__), .dinb(new_new_n1329__), .dout(new_new_n2442__));
  and1  g1501(.dina(new_new_n2442__), .dinb(new_new_n2440__), .dout(new_new_n2443__));
  or1   g1502(.dina(new_new_n2441__), .dinb(new_new_n2439__), .dout(new_new_n2444__));
  and1  g1503(.dina(new_new_n1306__), .dinb(new_new_n1243__), .dout(new_new_n2445__));
  or1   g1504(.dina(new_new_n1305__), .dinb(new_new_n1244__), .dout(new_new_n2446__));
  and1  g1505(.dina(new_new_n7237__), .dinb(new_new_n7238__), .dout(new_new_n2447__));
  or1   g1506(.dina(new_new_n7239__), .dinb(new_new_n7240__), .dout(new_new_n2448__));
  and1  g1507(.dina(new_new_n7242__), .dinb(new_new_n7238__), .dout(new_new_n2449__));
  or1   g1508(.dina(new_new_n7244__), .dinb(new_new_n7240__), .dout(new_new_n2450__));
  and1  g1509(.dina(new_new_n7242__), .dinb(new_new_n7237__), .dout(new_new_n2451__));
  or1   g1510(.dina(new_new_n7244__), .dinb(new_new_n7239__), .dout(new_new_n2452__));
  and1  g1511(.dina(new_new_n2452__), .dinb(new_new_n2450__), .dout(new_new_n2453__));
  or1   g1512(.dina(new_new_n2451__), .dinb(new_new_n2449__), .dout(new_new_n2454__));
  and1  g1513(.dina(new_new_n7132__), .dinb(new_new_n7246__), .dout(new_new_n2455__));
  or1   g1514(.dina(new_new_n7140__), .dinb(new_new_n7249__), .dout(new_new_n2456__));
  and1  g1515(.dina(new_new_n7250__), .dinb(new_new_n7251__), .dout(new_new_n2457__));
  or1   g1516(.dina(new_new_n7252__), .dinb(new_new_n7253__), .dout(new_new_n2458__));
  and1  g1517(.dina(new_new_n7255__), .dinb(new_new_n7251__), .dout(new_new_n2459__));
  or1   g1518(.dina(new_new_n7257__), .dinb(new_new_n7253__), .dout(new_new_n2460__));
  and1  g1519(.dina(new_new_n7255__), .dinb(new_new_n7250__), .dout(new_new_n2461__));
  or1   g1520(.dina(new_new_n7257__), .dinb(new_new_n7252__), .dout(new_new_n2462__));
  and1  g1521(.dina(new_new_n2462__), .dinb(new_new_n2460__), .dout(new_new_n2463__));
  or1   g1522(.dina(new_new_n2461__), .dinb(new_new_n2459__), .dout(new_new_n2464__));
  and1  g1523(.dina(new_new_n7258__), .dinb(new_new_n7259__), .dout(new_new_n2465__));
  or1   g1524(.dina(new_new_n7260__), .dinb(new_new_n7261__), .dout(new_new_n2466__));
  and1  g1525(.dina(new_new_n7263__), .dinb(new_new_n7258__), .dout(new_new_n2467__));
  or1   g1526(.dina(new_new_n7265__), .dinb(new_new_n7260__), .dout(new_new_n2468__));
  and1  g1527(.dina(new_new_n7263__), .dinb(new_new_n7259__), .dout(new_new_n2469__));
  or1   g1528(.dina(new_new_n7265__), .dinb(new_new_n7261__), .dout(new_new_n2470__));
  and1  g1529(.dina(new_new_n2470__), .dinb(new_new_n2468__), .dout(new_new_n2471__));
  or1   g1530(.dina(new_new_n2469__), .dinb(new_new_n2467__), .dout(new_new_n2472__));
  and1  g1531(.dina(new_new_n7133__), .dinb(new_new_n7267__), .dout(new_new_n2473__));
  or1   g1532(.dina(new_new_n7141__), .dinb(new_new_n7270__), .dout(new_new_n2474__));
  and1  g1533(.dina(new_new_n7271__), .dinb(new_new_n7272__), .dout(new_new_n2475__));
  or1   g1534(.dina(new_new_n7273__), .dinb(new_new_n7274__), .dout(new_new_n2476__));
  and1  g1535(.dina(new_new_n7276__), .dinb(new_new_n7262__), .dout(new_new_n2477__));
  or1   g1536(.dina(new_new_n7278__), .dinb(new_new_n7264__), .dout(new_new_n2478__));
  and1  g1537(.dina(new_new_n7279__), .dinb(new_new_n7280__), .dout(new_new_n2479__));
  or1   g1538(.dina(new_new_n7281__), .dinb(new_new_n7282__), .dout(new_new_n2480__));
  and1  g1539(.dina(new_new_n7284__), .dinb(new_new_n7280__), .dout(new_new_n2481__));
  or1   g1540(.dina(new_new_n7286__), .dinb(new_new_n7282__), .dout(new_new_n2482__));
  and1  g1541(.dina(new_new_n7284__), .dinb(new_new_n7279__), .dout(new_new_n2483__));
  or1   g1542(.dina(new_new_n7286__), .dinb(new_new_n7281__), .dout(new_new_n2484__));
  and1  g1543(.dina(new_new_n2484__), .dinb(new_new_n2482__), .dout(new_new_n2485__));
  or1   g1544(.dina(new_new_n2483__), .dinb(new_new_n2481__), .dout(new_new_n2486__));
  and1  g1545(.dina(new_new_n6732__), .dinb(new_new_n7267__), .dout(new_new_n2487__));
  or1   g1546(.dina(new_new_n6746__), .dinb(new_new_n7270__), .dout(new_new_n2488__));
  and1  g1547(.dina(new_new_n7287__), .dinb(new_new_n7288__), .dout(new_new_n2489__));
  or1   g1548(.dina(new_new_n7289__), .dinb(new_new_n7290__), .dout(new_new_n2490__));
  and1  g1549(.dina(new_new_n7292__), .dinb(new_new_n7288__), .dout(new_new_n2491__));
  or1   g1550(.dina(new_new_n7294__), .dinb(new_new_n7290__), .dout(new_new_n2492__));
  and1  g1551(.dina(new_new_n7292__), .dinb(new_new_n7287__), .dout(new_new_n2493__));
  or1   g1552(.dina(new_new_n7294__), .dinb(new_new_n7289__), .dout(new_new_n2494__));
  and1  g1553(.dina(new_new_n2494__), .dinb(new_new_n2492__), .dout(new_new_n2495__));
  or1   g1554(.dina(new_new_n2493__), .dinb(new_new_n2491__), .dout(new_new_n2496__));
  and1  g1555(.dina(new_new_n7276__), .dinb(new_new_n7272__), .dout(new_new_n2497__));
  or1   g1556(.dina(new_new_n7278__), .dinb(new_new_n7274__), .dout(new_new_n2498__));
  and1  g1557(.dina(new_new_n7275__), .dinb(new_new_n7271__), .dout(new_new_n2499__));
  or1   g1558(.dina(new_new_n7277__), .dinb(new_new_n7273__), .dout(new_new_n2500__));
  and1  g1559(.dina(new_new_n2500__), .dinb(new_new_n2498__), .dout(new_new_n2501__));
  or1   g1560(.dina(new_new_n2499__), .dinb(new_new_n2497__), .dout(new_new_n2502__));
  and1  g1561(.dina(new_new_n1434__), .dinb(new_new_n1428__), .dout(new_new_n2503__));
  or1   g1562(.dina(new_new_n1433__), .dinb(new_new_n1427__), .dout(new_new_n2504__));
  and1  g1563(.dina(new_new_n7133__), .dinb(new_new_n7296__), .dout(new_new_n2505__));
  or1   g1564(.dina(new_new_n7141__), .dinb(new_new_n7299__), .dout(new_new_n2506__));
  and1  g1565(.dina(new_new_n7301__), .dinb(new_new_n7302__), .dout(new_new_n2507__));
  or1   g1566(.dina(new_new_n7303__), .dinb(new_new_n7304__), .dout(new_new_n2508__));
  and1  g1567(.dina(new_new_n7306__), .dinb(new_new_n1371__), .dout(new_new_n2509__));
  or1   g1568(.dina(new_new_n7308__), .dinb(new_new_n1372__), .dout(new_new_n2510__));
  and1  g1569(.dina(new_new_n7309__), .dinb(new_new_n7310__), .dout(new_new_n2511__));
  or1   g1570(.dina(new_new_n7311__), .dinb(new_new_n7312__), .dout(new_new_n2512__));
  and1  g1571(.dina(new_new_n7314__), .dinb(new_new_n7310__), .dout(new_new_n2513__));
  or1   g1572(.dina(new_new_n7316__), .dinb(new_new_n7312__), .dout(new_new_n2514__));
  and1  g1573(.dina(new_new_n7314__), .dinb(new_new_n7309__), .dout(new_new_n2515__));
  or1   g1574(.dina(new_new_n7316__), .dinb(new_new_n7311__), .dout(new_new_n2516__));
  and1  g1575(.dina(new_new_n2516__), .dinb(new_new_n2514__), .dout(new_new_n2517__));
  or1   g1576(.dina(new_new_n2515__), .dinb(new_new_n2513__), .dout(new_new_n2518__));
  and1  g1577(.dina(new_new_n6734__), .dinb(new_new_n7296__), .dout(new_new_n2519__));
  or1   g1578(.dina(new_new_n6748__), .dinb(new_new_n7299__), .dout(new_new_n2520__));
  and1  g1579(.dina(new_new_n7317__), .dinb(new_new_n7318__), .dout(new_new_n2521__));
  or1   g1580(.dina(new_new_n7319__), .dinb(new_new_n7320__), .dout(new_new_n2522__));
  and1  g1581(.dina(new_new_n7322__), .dinb(new_new_n7313__), .dout(new_new_n2523__));
  or1   g1582(.dina(new_new_n7324__), .dinb(new_new_n7315__), .dout(new_new_n2524__));
  and1  g1583(.dina(new_new_n7325__), .dinb(new_new_n7326__), .dout(new_new_n2525__));
  or1   g1584(.dina(new_new_n7327__), .dinb(new_new_n7328__), .dout(new_new_n2526__));
  and1  g1585(.dina(new_new_n7330__), .dinb(new_new_n7326__), .dout(new_new_n2527__));
  or1   g1586(.dina(new_new_n7332__), .dinb(new_new_n7328__), .dout(new_new_n2528__));
  and1  g1587(.dina(new_new_n7330__), .dinb(new_new_n7325__), .dout(new_new_n2529__));
  or1   g1588(.dina(new_new_n7332__), .dinb(new_new_n7327__), .dout(new_new_n2530__));
  and1  g1589(.dina(new_new_n2530__), .dinb(new_new_n2528__), .dout(new_new_n2531__));
  or1   g1590(.dina(new_new_n2529__), .dinb(new_new_n2527__), .dout(new_new_n2532__));
  and1  g1591(.dina(new_new_n7297__), .dinb(new_new_n6761__), .dout(new_new_n2533__));
  or1   g1592(.dina(new_new_n7300__), .dinb(new_new_n6775__), .dout(new_new_n2534__));
  and1  g1593(.dina(new_new_n7333__), .dinb(new_new_n7334__), .dout(new_new_n2535__));
  or1   g1594(.dina(new_new_n7335__), .dinb(new_new_n7336__), .dout(new_new_n2536__));
  and1  g1595(.dina(new_new_n7338__), .dinb(new_new_n7334__), .dout(new_new_n2537__));
  or1   g1596(.dina(new_new_n7340__), .dinb(new_new_n7336__), .dout(new_new_n2538__));
  and1  g1597(.dina(new_new_n7338__), .dinb(new_new_n7333__), .dout(new_new_n2539__));
  or1   g1598(.dina(new_new_n7340__), .dinb(new_new_n7335__), .dout(new_new_n2540__));
  and1  g1599(.dina(new_new_n2540__), .dinb(new_new_n2538__), .dout(new_new_n2541__));
  or1   g1600(.dina(new_new_n2539__), .dinb(new_new_n2537__), .dout(new_new_n2542__));
  and1  g1601(.dina(new_new_n7322__), .dinb(new_new_n7318__), .dout(new_new_n2543__));
  or1   g1602(.dina(new_new_n7324__), .dinb(new_new_n7320__), .dout(new_new_n2544__));
  and1  g1603(.dina(new_new_n7321__), .dinb(new_new_n7317__), .dout(new_new_n2545__));
  or1   g1604(.dina(new_new_n7323__), .dinb(new_new_n7319__), .dout(new_new_n2546__));
  and1  g1605(.dina(new_new_n2546__), .dinb(new_new_n2544__), .dout(new_new_n2547__));
  or1   g1606(.dina(new_new_n2545__), .dinb(new_new_n2543__), .dout(new_new_n2548__));
  and1  g1607(.dina(new_new_n7306__), .dinb(new_new_n7302__), .dout(new_new_n2549__));
  or1   g1608(.dina(new_new_n7308__), .dinb(new_new_n7304__), .dout(new_new_n2550__));
  and1  g1609(.dina(new_new_n7305__), .dinb(new_new_n7301__), .dout(new_new_n2551__));
  or1   g1610(.dina(new_new_n7307__), .dinb(new_new_n7303__), .dout(new_new_n2552__));
  and1  g1611(.dina(new_new_n2552__), .dinb(new_new_n2550__), .dout(new_new_n2553__));
  or1   g1612(.dina(new_new_n2551__), .dinb(new_new_n2549__), .dout(new_new_n2554__));
  and1  g1613(.dina(new_new_n7342__), .dinb(new_new_n1295__), .dout(new_new_n2555__));
  or1   g1614(.dina(new_new_n7344__), .dinb(new_new_n1296__), .dout(new_new_n2556__));
  and1  g1615(.dina(new_new_n7345__), .dinb(new_new_n7346__), .dout(new_new_n2557__));
  or1   g1616(.dina(new_new_n7347__), .dinb(new_new_n7348__), .dout(new_new_n2558__));
  and1  g1617(.dina(new_new_n7350__), .dinb(new_new_n7346__), .dout(new_new_n2559__));
  or1   g1618(.dina(new_new_n7352__), .dinb(new_new_n7348__), .dout(new_new_n2560__));
  and1  g1619(.dina(new_new_n7350__), .dinb(new_new_n7345__), .dout(new_new_n2561__));
  or1   g1620(.dina(new_new_n7352__), .dinb(new_new_n7347__), .dout(new_new_n2562__));
  and1  g1621(.dina(new_new_n2562__), .dinb(new_new_n2560__), .dout(new_new_n2563__));
  or1   g1622(.dina(new_new_n2561__), .dinb(new_new_n2559__), .dout(new_new_n2564__));
  and1  g1623(.dina(new_new_n6734__), .dinb(new_new_n7354__), .dout(new_new_n2565__));
  or1   g1624(.dina(new_new_n6748__), .dinb(new_new_n7357__), .dout(new_new_n2566__));
  and1  g1625(.dina(new_new_n7358__), .dinb(new_new_n7359__), .dout(new_new_n2567__));
  or1   g1626(.dina(new_new_n7360__), .dinb(new_new_n7361__), .dout(new_new_n2568__));
  and1  g1627(.dina(new_new_n7363__), .dinb(new_new_n7349__), .dout(new_new_n2569__));
  or1   g1628(.dina(new_new_n7365__), .dinb(new_new_n7351__), .dout(new_new_n2570__));
  and1  g1629(.dina(new_new_n7366__), .dinb(new_new_n7367__), .dout(new_new_n2571__));
  or1   g1630(.dina(new_new_n7368__), .dinb(new_new_n7369__), .dout(new_new_n2572__));
  and1  g1631(.dina(new_new_n7371__), .dinb(new_new_n7367__), .dout(new_new_n2573__));
  or1   g1632(.dina(new_new_n7373__), .dinb(new_new_n7369__), .dout(new_new_n2574__));
  and1  g1633(.dina(new_new_n7371__), .dinb(new_new_n7366__), .dout(new_new_n2575__));
  or1   g1634(.dina(new_new_n7373__), .dinb(new_new_n7368__), .dout(new_new_n2576__));
  and1  g1635(.dina(new_new_n2576__), .dinb(new_new_n2574__), .dout(new_new_n2577__));
  or1   g1636(.dina(new_new_n2575__), .dinb(new_new_n2573__), .dout(new_new_n2578__));
  and1  g1637(.dina(new_new_n7354__), .dinb(new_new_n6763__), .dout(new_new_n2579__));
  or1   g1638(.dina(new_new_n7357__), .dinb(new_new_n6777__), .dout(new_new_n2580__));
  and1  g1639(.dina(new_new_n7374__), .dinb(new_new_n7375__), .dout(new_new_n2581__));
  or1   g1640(.dina(new_new_n7376__), .dinb(new_new_n7377__), .dout(new_new_n2582__));
  and1  g1641(.dina(new_new_n7379__), .dinb(new_new_n7370__), .dout(new_new_n2583__));
  or1   g1642(.dina(new_new_n7381__), .dinb(new_new_n7372__), .dout(new_new_n2584__));
  and1  g1643(.dina(new_new_n7382__), .dinb(new_new_n7383__), .dout(new_new_n2585__));
  or1   g1644(.dina(new_new_n7384__), .dinb(new_new_n7385__), .dout(new_new_n2586__));
  and1  g1645(.dina(new_new_n7342__), .dinb(new_new_n1379__), .dout(new_new_n2587__));
  or1   g1646(.dina(new_new_n7344__), .dinb(new_new_n1380__), .dout(new_new_n2588__));
  and1  g1647(.dina(new_new_n7341__), .dinb(new_new_n1332__), .dout(new_new_n2589__));
  or1   g1648(.dina(new_new_n7343__), .dinb(new_new_n1331__), .dout(new_new_n2590__));
  and1  g1649(.dina(new_new_n2590__), .dinb(new_new_n2588__), .dout(new_new_n2591__));
  or1   g1650(.dina(new_new_n2589__), .dinb(new_new_n2587__), .dout(new_new_n2592__));
  and1  g1651(.dina(new_new_n1308__), .dinb(new_new_n1245__), .dout(new_new_n2593__));
  or1   g1652(.dina(new_new_n1307__), .dinb(new_new_n1246__), .dout(new_new_n2594__));
  and1  g1653(.dina(new_new_n7386__), .dinb(new_new_n7387__), .dout(new_new_n2595__));
  or1   g1654(.dina(new_new_n7388__), .dinb(new_new_n7389__), .dout(new_new_n2596__));
  and1  g1655(.dina(new_new_n7391__), .dinb(new_new_n7387__), .dout(new_new_n2597__));
  or1   g1656(.dina(new_new_n7393__), .dinb(new_new_n7389__), .dout(new_new_n2598__));
  and1  g1657(.dina(new_new_n7391__), .dinb(new_new_n7386__), .dout(new_new_n2599__));
  or1   g1658(.dina(new_new_n7393__), .dinb(new_new_n7388__), .dout(new_new_n2600__));
  and1  g1659(.dina(new_new_n2600__), .dinb(new_new_n2598__), .dout(new_new_n2601__));
  or1   g1660(.dina(new_new_n2599__), .dinb(new_new_n2597__), .dout(new_new_n2602__));
  and1  g1661(.dina(new_new_n6733__), .dinb(new_new_n7395__), .dout(new_new_n2603__));
  or1   g1662(.dina(new_new_n6747__), .dinb(new_new_n7398__), .dout(new_new_n2604__));
  and1  g1663(.dina(new_new_n7399__), .dinb(new_new_n7400__), .dout(new_new_n2605__));
  or1   g1664(.dina(new_new_n7401__), .dinb(new_new_n7402__), .dout(new_new_n2606__));
  and1  g1665(.dina(new_new_n7404__), .dinb(new_new_n7400__), .dout(new_new_n2607__));
  or1   g1666(.dina(new_new_n7406__), .dinb(new_new_n7402__), .dout(new_new_n2608__));
  and1  g1667(.dina(new_new_n7404__), .dinb(new_new_n7399__), .dout(new_new_n2609__));
  or1   g1668(.dina(new_new_n7406__), .dinb(new_new_n7401__), .dout(new_new_n2610__));
  and1  g1669(.dina(new_new_n2610__), .dinb(new_new_n2608__), .dout(new_new_n2611__));
  or1   g1670(.dina(new_new_n2609__), .dinb(new_new_n2607__), .dout(new_new_n2612__));
  and1  g1671(.dina(new_new_n7407__), .dinb(new_new_n7408__), .dout(new_new_n2613__));
  or1   g1672(.dina(new_new_n7409__), .dinb(new_new_n7410__), .dout(new_new_n2614__));
  and1  g1673(.dina(new_new_n7412__), .dinb(new_new_n7407__), .dout(new_new_n2615__));
  or1   g1674(.dina(new_new_n7414__), .dinb(new_new_n7409__), .dout(new_new_n2616__));
  and1  g1675(.dina(new_new_n7412__), .dinb(new_new_n7408__), .dout(new_new_n2617__));
  or1   g1676(.dina(new_new_n7414__), .dinb(new_new_n7410__), .dout(new_new_n2618__));
  and1  g1677(.dina(new_new_n2618__), .dinb(new_new_n2616__), .dout(new_new_n2619__));
  or1   g1678(.dina(new_new_n2617__), .dinb(new_new_n2615__), .dout(new_new_n2620__));
  and1  g1679(.dina(new_new_n6736__), .dinb(new_new_n7416__), .dout(new_new_n2621__));
  or1   g1680(.dina(new_new_n6750__), .dinb(new_new_n7419__), .dout(new_new_n2622__));
  and1  g1681(.dina(new_new_n7420__), .dinb(new_new_n7421__), .dout(new_new_n2623__));
  or1   g1682(.dina(new_new_n7422__), .dinb(new_new_n7423__), .dout(new_new_n2624__));
  and1  g1683(.dina(new_new_n7425__), .dinb(new_new_n7411__), .dout(new_new_n2625__));
  or1   g1684(.dina(new_new_n7427__), .dinb(new_new_n7413__), .dout(new_new_n2626__));
  and1  g1685(.dina(new_new_n7428__), .dinb(new_new_n7429__), .dout(new_new_n2627__));
  or1   g1686(.dina(new_new_n7430__), .dinb(new_new_n7431__), .dout(new_new_n2628__));
  and1  g1687(.dina(new_new_n7433__), .dinb(new_new_n7429__), .dout(new_new_n2629__));
  or1   g1688(.dina(new_new_n7435__), .dinb(new_new_n7431__), .dout(new_new_n2630__));
  and1  g1689(.dina(new_new_n7433__), .dinb(new_new_n7428__), .dout(new_new_n2631__));
  or1   g1690(.dina(new_new_n7435__), .dinb(new_new_n7430__), .dout(new_new_n2632__));
  and1  g1691(.dina(new_new_n2632__), .dinb(new_new_n2630__), .dout(new_new_n2633__));
  or1   g1692(.dina(new_new_n2631__), .dinb(new_new_n2629__), .dout(new_new_n2634__));
  and1  g1693(.dina(new_new_n7416__), .dinb(new_new_n6763__), .dout(new_new_n2635__));
  or1   g1694(.dina(new_new_n7419__), .dinb(new_new_n6777__), .dout(new_new_n2636__));
  and1  g1695(.dina(new_new_n7436__), .dinb(new_new_n7437__), .dout(new_new_n2637__));
  or1   g1696(.dina(new_new_n7438__), .dinb(new_new_n7439__), .dout(new_new_n2638__));
  and1  g1697(.dina(new_new_n7441__), .dinb(new_new_n7437__), .dout(new_new_n2639__));
  or1   g1698(.dina(new_new_n7443__), .dinb(new_new_n7439__), .dout(new_new_n2640__));
  and1  g1699(.dina(new_new_n7441__), .dinb(new_new_n7436__), .dout(new_new_n2641__));
  or1   g1700(.dina(new_new_n7443__), .dinb(new_new_n7438__), .dout(new_new_n2642__));
  and1  g1701(.dina(new_new_n2642__), .dinb(new_new_n2640__), .dout(new_new_n2643__));
  or1   g1702(.dina(new_new_n2641__), .dinb(new_new_n2639__), .dout(new_new_n2644__));
  and1  g1703(.dina(new_new_n7425__), .dinb(new_new_n7421__), .dout(new_new_n2645__));
  or1   g1704(.dina(new_new_n7427__), .dinb(new_new_n7423__), .dout(new_new_n2646__));
  and1  g1705(.dina(new_new_n7424__), .dinb(new_new_n7420__), .dout(new_new_n2647__));
  or1   g1706(.dina(new_new_n7426__), .dinb(new_new_n7422__), .dout(new_new_n2648__));
  and1  g1707(.dina(new_new_n2648__), .dinb(new_new_n2646__), .dout(new_new_n2649__));
  or1   g1708(.dina(new_new_n2647__), .dinb(new_new_n2645__), .dout(new_new_n2650__));
  and1  g1709(.dina(new_new_n1436__), .dinb(new_new_n1430__), .dout(new_new_n2651__));
  or1   g1710(.dina(new_new_n1435__), .dinb(new_new_n1429__), .dout(new_new_n2652__));
  and1  g1711(.dina(new_new_n6736__), .dinb(new_new_n7445__), .dout(new_new_n2653__));
  or1   g1712(.dina(new_new_n6750__), .dinb(new_new_n7447__), .dout(new_new_n2654__));
  and1  g1713(.dina(new_new_n7449__), .dinb(new_new_n7450__), .dout(new_new_n2655__));
  or1   g1714(.dina(new_new_n7451__), .dinb(new_new_n7452__), .dout(new_new_n2656__));
  and1  g1715(.dina(new_new_n7454__), .dinb(new_new_n1373__), .dout(new_new_n2657__));
  or1   g1716(.dina(new_new_n7456__), .dinb(new_new_n1374__), .dout(new_new_n2658__));
  and1  g1717(.dina(new_new_n7457__), .dinb(new_new_n7458__), .dout(new_new_n2659__));
  or1   g1718(.dina(new_new_n7459__), .dinb(new_new_n7460__), .dout(new_new_n2660__));
  and1  g1719(.dina(new_new_n7462__), .dinb(new_new_n7458__), .dout(new_new_n2661__));
  or1   g1720(.dina(new_new_n7464__), .dinb(new_new_n7460__), .dout(new_new_n2662__));
  and1  g1721(.dina(new_new_n7462__), .dinb(new_new_n7457__), .dout(new_new_n2663__));
  or1   g1722(.dina(new_new_n7464__), .dinb(new_new_n7459__), .dout(new_new_n2664__));
  and1  g1723(.dina(new_new_n2664__), .dinb(new_new_n2662__), .dout(new_new_n2665__));
  or1   g1724(.dina(new_new_n2663__), .dinb(new_new_n2661__), .dout(new_new_n2666__));
  and1  g1725(.dina(new_new_n7445__), .dinb(new_new_n6764__), .dout(new_new_n2667__));
  or1   g1726(.dina(new_new_n7447__), .dinb(new_new_n6778__), .dout(new_new_n2668__));
  and1  g1727(.dina(new_new_n7465__), .dinb(new_new_n7466__), .dout(new_new_n2669__));
  or1   g1728(.dina(new_new_n7467__), .dinb(new_new_n7468__), .dout(new_new_n2670__));
  and1  g1729(.dina(new_new_n7470__), .dinb(new_new_n7461__), .dout(new_new_n2671__));
  or1   g1730(.dina(new_new_n7472__), .dinb(new_new_n7463__), .dout(new_new_n2672__));
  and1  g1731(.dina(new_new_n7473__), .dinb(new_new_n7474__), .dout(new_new_n2673__));
  or1   g1732(.dina(new_new_n7475__), .dinb(new_new_n7476__), .dout(new_new_n2674__));
  and1  g1733(.dina(new_new_n7478__), .dinb(new_new_n7474__), .dout(new_new_n2675__));
  or1   g1734(.dina(new_new_n7480__), .dinb(new_new_n7476__), .dout(new_new_n2676__));
  and1  g1735(.dina(new_new_n7478__), .dinb(new_new_n7473__), .dout(new_new_n2677__));
  or1   g1736(.dina(new_new_n7480__), .dinb(new_new_n7475__), .dout(new_new_n2678__));
  and1  g1737(.dina(new_new_n2678__), .dinb(new_new_n2676__), .dout(new_new_n2679__));
  or1   g1738(.dina(new_new_n2677__), .dinb(new_new_n2675__), .dout(new_new_n2680__));
  and1  g1739(.dina(new_new_n7444__), .dinb(new_new_n6808__), .dout(new_new_n2681__));
  or1   g1740(.dina(new_new_n7448__), .dinb(new_new_n6818__), .dout(new_new_n2682__));
  and1  g1741(.dina(new_new_n7481__), .dinb(new_new_n7482__), .dout(new_new_n2683__));
  or1   g1742(.dina(new_new_n7483__), .dinb(new_new_n7484__), .dout(new_new_n2684__));
  and1  g1743(.dina(new_new_n7486__), .dinb(new_new_n7482__), .dout(new_new_n2685__));
  or1   g1744(.dina(new_new_n7488__), .dinb(new_new_n7484__), .dout(new_new_n2686__));
  and1  g1745(.dina(new_new_n7486__), .dinb(new_new_n7481__), .dout(new_new_n2687__));
  or1   g1746(.dina(new_new_n7488__), .dinb(new_new_n7483__), .dout(new_new_n2688__));
  and1  g1747(.dina(new_new_n2688__), .dinb(new_new_n2686__), .dout(new_new_n2689__));
  or1   g1748(.dina(new_new_n2687__), .dinb(new_new_n2685__), .dout(new_new_n2690__));
  and1  g1749(.dina(new_new_n7470__), .dinb(new_new_n7466__), .dout(new_new_n2691__));
  or1   g1750(.dina(new_new_n7472__), .dinb(new_new_n7468__), .dout(new_new_n2692__));
  and1  g1751(.dina(new_new_n7469__), .dinb(new_new_n7465__), .dout(new_new_n2693__));
  or1   g1752(.dina(new_new_n7471__), .dinb(new_new_n7467__), .dout(new_new_n2694__));
  and1  g1753(.dina(new_new_n2694__), .dinb(new_new_n2692__), .dout(new_new_n2695__));
  or1   g1754(.dina(new_new_n2693__), .dinb(new_new_n2691__), .dout(new_new_n2696__));
  and1  g1755(.dina(new_new_n7454__), .dinb(new_new_n7450__), .dout(new_new_n2697__));
  or1   g1756(.dina(new_new_n7456__), .dinb(new_new_n7452__), .dout(new_new_n2698__));
  and1  g1757(.dina(new_new_n7453__), .dinb(new_new_n7449__), .dout(new_new_n2699__));
  or1   g1758(.dina(new_new_n7455__), .dinb(new_new_n7451__), .dout(new_new_n2700__));
  and1  g1759(.dina(new_new_n2700__), .dinb(new_new_n2698__), .dout(new_new_n2701__));
  or1   g1760(.dina(new_new_n2699__), .dinb(new_new_n2697__), .dout(new_new_n2702__));
  and1  g1761(.dina(new_new_n7490__), .dinb(new_new_n1297__), .dout(new_new_n2703__));
  or1   g1762(.dina(new_new_n7492__), .dinb(new_new_n1298__), .dout(new_new_n2704__));
  and1  g1763(.dina(new_new_n7493__), .dinb(new_new_n7494__), .dout(new_new_n2705__));
  or1   g1764(.dina(new_new_n7495__), .dinb(new_new_n7496__), .dout(new_new_n2706__));
  and1  g1765(.dina(new_new_n7498__), .dinb(new_new_n7494__), .dout(new_new_n2707__));
  or1   g1766(.dina(new_new_n7500__), .dinb(new_new_n7496__), .dout(new_new_n2708__));
  and1  g1767(.dina(new_new_n7498__), .dinb(new_new_n7493__), .dout(new_new_n2709__));
  or1   g1768(.dina(new_new_n7500__), .dinb(new_new_n7495__), .dout(new_new_n2710__));
  and1  g1769(.dina(new_new_n2710__), .dinb(new_new_n2708__), .dout(new_new_n2711__));
  or1   g1770(.dina(new_new_n2709__), .dinb(new_new_n2707__), .dout(new_new_n2712__));
  and1  g1771(.dina(new_new_n7502__), .dinb(new_new_n6764__), .dout(new_new_n2713__));
  or1   g1772(.dina(new_new_n7504__), .dinb(new_new_n6778__), .dout(new_new_n2714__));
  and1  g1773(.dina(new_new_n7505__), .dinb(new_new_n7506__), .dout(new_new_n2715__));
  or1   g1774(.dina(new_new_n7507__), .dinb(new_new_n7508__), .dout(new_new_n2716__));
  and1  g1775(.dina(new_new_n7510__), .dinb(new_new_n7497__), .dout(new_new_n2717__));
  or1   g1776(.dina(new_new_n7512__), .dinb(new_new_n7499__), .dout(new_new_n2718__));
  and1  g1777(.dina(new_new_n7513__), .dinb(new_new_n7514__), .dout(new_new_n2719__));
  or1   g1778(.dina(new_new_n7515__), .dinb(new_new_n7516__), .dout(new_new_n2720__));
  and1  g1779(.dina(new_new_n7518__), .dinb(new_new_n7514__), .dout(new_new_n2721__));
  or1   g1780(.dina(new_new_n7520__), .dinb(new_new_n7516__), .dout(new_new_n2722__));
  and1  g1781(.dina(new_new_n7518__), .dinb(new_new_n7513__), .dout(new_new_n2723__));
  or1   g1782(.dina(new_new_n7520__), .dinb(new_new_n7515__), .dout(new_new_n2724__));
  and1  g1783(.dina(new_new_n2724__), .dinb(new_new_n2722__), .dout(new_new_n2725__));
  or1   g1784(.dina(new_new_n2723__), .dinb(new_new_n2721__), .dout(new_new_n2726__));
  and1  g1785(.dina(new_new_n7502__), .dinb(new_new_n6808__), .dout(new_new_n2727__));
  or1   g1786(.dina(new_new_n7504__), .dinb(new_new_n6818__), .dout(new_new_n2728__));
  and1  g1787(.dina(new_new_n7521__), .dinb(new_new_n7522__), .dout(new_new_n2729__));
  or1   g1788(.dina(new_new_n7523__), .dinb(new_new_n7524__), .dout(new_new_n2730__));
  and1  g1789(.dina(new_new_n7526__), .dinb(new_new_n7517__), .dout(new_new_n2731__));
  or1   g1790(.dina(new_new_n7528__), .dinb(new_new_n7519__), .dout(new_new_n2732__));
  and1  g1791(.dina(new_new_n7529__), .dinb(new_new_n7530__), .dout(new_new_n2733__));
  or1   g1792(.dina(new_new_n7531__), .dinb(new_new_n7532__), .dout(new_new_n2734__));
  and1  g1793(.dina(new_new_n7533__), .dinb(new_new_n7534__), .dout(new_new_n2735__));
  or1   g1794(.dina(new_new_n7535__), .dinb(new_new_n7536__), .dout(new_new_n2736__));
  and1  g1795(.dina(new_new_n7538__), .dinb(new_new_n7533__), .dout(new_new_n2737__));
  or1   g1796(.dina(new_new_n7540__), .dinb(new_new_n7535__), .dout(new_new_n2738__));
  and1  g1797(.dina(new_new_n7538__), .dinb(new_new_n7534__), .dout(new_new_n2739__));
  or1   g1798(.dina(new_new_n7540__), .dinb(new_new_n7536__), .dout(new_new_n2740__));
  and1  g1799(.dina(new_new_n2740__), .dinb(new_new_n2738__), .dout(new_new_n2741__));
  or1   g1800(.dina(new_new_n2739__), .dinb(new_new_n2737__), .dout(new_new_n2742__));
  and1  g1801(.dina(new_new_n7542__), .dinb(new_new_n6767__), .dout(new_new_n2743__));
  or1   g1802(.dina(new_new_n7544__), .dinb(new_new_n6781__), .dout(new_new_n2744__));
  and1  g1803(.dina(new_new_n7545__), .dinb(new_new_n7546__), .dout(new_new_n2745__));
  or1   g1804(.dina(new_new_n7547__), .dinb(new_new_n7548__), .dout(new_new_n2746__));
  and1  g1805(.dina(new_new_n7550__), .dinb(new_new_n7546__), .dout(new_new_n2747__));
  or1   g1806(.dina(new_new_n7552__), .dinb(new_new_n7548__), .dout(new_new_n2748__));
  and1  g1807(.dina(new_new_n7550__), .dinb(new_new_n7545__), .dout(new_new_n2749__));
  or1   g1808(.dina(new_new_n7552__), .dinb(new_new_n7547__), .dout(new_new_n2750__));
  and1  g1809(.dina(new_new_n2750__), .dinb(new_new_n2748__), .dout(new_new_n2751__));
  or1   g1810(.dina(new_new_n2749__), .dinb(new_new_n2747__), .dout(new_new_n2752__));
  and1  g1811(.dina(new_new_n6910__), .dinb(new_new_n6898__), .dout(new_new_n2753__));
  or1   g1812(.dina(new_new_n6912__), .dinb(new_new_n6900__), .dout(new_new_n2754__));
  and1  g1813(.dina(new_new_n7553__), .dinb(new_new_n7554__), .dout(new_new_n2755__));
  or1   g1814(.dina(new_new_n7555__), .dinb(new_new_n7556__), .dout(new_new_n2756__));
  and1  g1815(.dina(new_new_n7558__), .dinb(new_new_n7554__), .dout(new_new_n2757__));
  or1   g1816(.dina(new_new_n7560__), .dinb(new_new_n7556__), .dout(new_new_n2758__));
  and1  g1817(.dina(new_new_n7558__), .dinb(new_new_n7553__), .dout(new_new_n2759__));
  or1   g1818(.dina(new_new_n7560__), .dinb(new_new_n7555__), .dout(new_new_n2760__));
  and1  g1819(.dina(new_new_n2760__), .dinb(new_new_n2758__), .dout(new_new_n2761__));
  or1   g1820(.dina(new_new_n2759__), .dinb(new_new_n2757__), .dout(new_new_n2762__));
  and1  g1821(.dina(new_new_n6903__), .dinb(new_new_n6810__), .dout(new_new_n2763__));
  or1   g1822(.dina(new_new_n6905__), .dinb(new_new_n6820__), .dout(new_new_n2764__));
  and1  g1823(.dina(new_new_n7561__), .dinb(new_new_n7562__), .dout(new_new_n2765__));
  or1   g1824(.dina(new_new_n7563__), .dinb(new_new_n7564__), .dout(new_new_n2766__));
  and1  g1825(.dina(new_new_n7566__), .dinb(new_new_n7562__), .dout(new_new_n2767__));
  or1   g1826(.dina(new_new_n7568__), .dinb(new_new_n7564__), .dout(new_new_n2768__));
  and1  g1827(.dina(new_new_n7566__), .dinb(new_new_n7561__), .dout(new_new_n2769__));
  or1   g1828(.dina(new_new_n7568__), .dinb(new_new_n7563__), .dout(new_new_n2770__));
  and1  g1829(.dina(new_new_n2770__), .dinb(new_new_n2768__), .dout(new_new_n2771__));
  or1   g1830(.dina(new_new_n2769__), .dinb(new_new_n2767__), .dout(new_new_n2772__));
  and1  g1831(.dina(new_new_n6926__), .dinb(new_new_n6918__), .dout(new_new_n2773__));
  or1   g1832(.dina(new_new_n6928__), .dinb(new_new_n6920__), .dout(new_new_n2774__));
  and1  g1833(.dina(new_new_n7569__), .dinb(new_new_n7570__), .dout(new_new_n2775__));
  or1   g1834(.dina(new_new_n7571__), .dinb(new_new_n7572__), .dout(new_new_n2776__));
  and1  g1835(.dina(new_new_n7574__), .dinb(new_new_n7570__), .dout(new_new_n2777__));
  or1   g1836(.dina(new_new_n7576__), .dinb(new_new_n7572__), .dout(new_new_n2778__));
  and1  g1837(.dina(new_new_n7574__), .dinb(new_new_n7569__), .dout(new_new_n2779__));
  or1   g1838(.dina(new_new_n7576__), .dinb(new_new_n7571__), .dout(new_new_n2780__));
  and1  g1839(.dina(new_new_n2780__), .dinb(new_new_n2778__), .dout(new_new_n2781__));
  or1   g1840(.dina(new_new_n2779__), .dinb(new_new_n2777__), .dout(new_new_n2782__));
  and1  g1841(.dina(new_new_n6836__), .dinb(new_new_n6884__), .dout(new_new_n2783__));
  or1   g1842(.dina(new_new_n6838__), .dinb(new_new_n6890__), .dout(new_new_n2784__));
  and1  g1843(.dina(new_new_n7577__), .dinb(new_new_n7578__), .dout(new_new_n2785__));
  or1   g1844(.dina(new_new_n7579__), .dinb(new_new_n7580__), .dout(new_new_n2786__));
  and1  g1845(.dina(new_new_n7582__), .dinb(new_new_n7578__), .dout(new_new_n2787__));
  or1   g1846(.dina(new_new_n7584__), .dinb(new_new_n7580__), .dout(new_new_n2788__));
  and1  g1847(.dina(new_new_n7582__), .dinb(new_new_n7577__), .dout(new_new_n2789__));
  or1   g1848(.dina(new_new_n7584__), .dinb(new_new_n7579__), .dout(new_new_n2790__));
  and1  g1849(.dina(new_new_n2790__), .dinb(new_new_n2788__), .dout(new_new_n2791__));
  or1   g1850(.dina(new_new_n2789__), .dinb(new_new_n2787__), .dout(new_new_n2792__));
  and1  g1851(.dina(new_new_n2244__), .dinb(new_new_n6935__), .dout(new_new_n2793__));
  or1   g1852(.dina(new_new_n7585__), .dinb(new_new_n6937__), .dout(new_new_n2794__));
  and1  g1853(.dina(new_new_n7586__), .dinb(new_new_n7587__), .dout(new_new_n2795__));
  or1   g1854(.dina(new_new_n2793__), .dinb(new_new_n2791__), .dout(new_new_n2796__));
  and1  g1855(.dina(new_new_n7588__), .dinb(new_new_n7587__), .dout(new_new_n2797__));
  and1  g1856(.dina(new_new_n7588__), .dinb(new_new_n7586__), .dout(new_new_n2798__));
  or1   g1857(.dina(new_new_n2798__), .dinb(new_new_n2797__), .dout(new_new_n2799__));
  and1  g1858(.dina(new_new_n7589__), .dinb(new_new_n2324__), .dout(new_new_n2800__));
  or1   g1859(.dina(new_new_n2349__), .dinb(new_new_n7590__), .dout(new_new_n2801__));
  and1  g1860(.dina(new_new_n6866__), .dinb(new_new_n7594__), .dout(new_new_n2802__));
  or1   g1861(.dina(new_new_n6875__), .dinb(new_new_n7607__), .dout(new_new_n2803__));
  and1  g1862(.dina(new_new_n7618__), .dinb(new_new_n1477__), .dout(new_new_n2804__));
  or1   g1863(.dina(new_new_n7620__), .dinb(new_new_n1478__), .dout(new_new_n2805__));
  and1  g1864(.dina(new_new_n7618__), .dinb(new_new_n1408__), .dout(new_new_n2806__));
  or1   g1865(.dina(new_new_n7620__), .dinb(new_new_n1407__), .dout(new_new_n2807__));
  and1  g1866(.dina(new_new_n2807__), .dinb(new_new_n2805__), .dout(new_new_n2808__));
  or1   g1867(.dina(new_new_n2806__), .dinb(new_new_n2804__), .dout(new_new_n2809__));
  and1  g1868(.dina(new_new_n7052__), .dinb(new_new_n1391__), .dout(new_new_n2810__));
  or1   g1869(.dina(new_new_n7054__), .dinb(new_new_n1392__), .dout(new_new_n2811__));
  and1  g1870(.dina(new_new_n7621__), .dinb(new_new_n7622__), .dout(new_new_n2812__));
  or1   g1871(.dina(new_new_n7623__), .dinb(new_new_n7624__), .dout(new_new_n2813__));
  and1  g1872(.dina(new_new_n7626__), .dinb(new_new_n7622__), .dout(new_new_n2814__));
  or1   g1873(.dina(new_new_n7628__), .dinb(new_new_n7624__), .dout(new_new_n2815__));
  and1  g1874(.dina(new_new_n7626__), .dinb(new_new_n7621__), .dout(new_new_n2816__));
  or1   g1875(.dina(new_new_n7628__), .dinb(new_new_n7623__), .dout(new_new_n2817__));
  and1  g1876(.dina(new_new_n2817__), .dinb(new_new_n2815__), .dout(new_new_n2818__));
  or1   g1877(.dina(new_new_n2816__), .dinb(new_new_n2814__), .dout(new_new_n2819__));
  and1  g1878(.dina(new_new_n6943__), .dinb(new_new_n7631__), .dout(new_new_n2820__));
  or1   g1879(.dina(new_new_n6956__), .dinb(new_new_n7635__), .dout(new_new_n2821__));
  and1  g1880(.dina(new_new_n7637__), .dinb(new_new_n7638__), .dout(new_new_n2822__));
  or1   g1881(.dina(new_new_n7639__), .dinb(new_new_n7640__), .dout(new_new_n2823__));
  and1  g1882(.dina(new_new_n7642__), .dinb(new_new_n7638__), .dout(new_new_n2824__));
  or1   g1883(.dina(new_new_n7644__), .dinb(new_new_n7640__), .dout(new_new_n2825__));
  and1  g1884(.dina(new_new_n7642__), .dinb(new_new_n7637__), .dout(new_new_n2826__));
  or1   g1885(.dina(new_new_n7644__), .dinb(new_new_n7639__), .dout(new_new_n2827__));
  and1  g1886(.dina(new_new_n2827__), .dinb(new_new_n2825__), .dout(new_new_n2828__));
  or1   g1887(.dina(new_new_n2826__), .dinb(new_new_n2824__), .dout(new_new_n2829__));
  and1  g1888(.dina(new_new_n7068__), .dinb(new_new_n7060__), .dout(new_new_n2830__));
  or1   g1889(.dina(new_new_n7070__), .dinb(new_new_n7062__), .dout(new_new_n2831__));
  and1  g1890(.dina(new_new_n7645__), .dinb(new_new_n7646__), .dout(new_new_n2832__));
  or1   g1891(.dina(new_new_n7647__), .dinb(new_new_n7648__), .dout(new_new_n2833__));
  and1  g1892(.dina(new_new_n7650__), .dinb(new_new_n7646__), .dout(new_new_n2834__));
  or1   g1893(.dina(new_new_n7652__), .dinb(new_new_n7648__), .dout(new_new_n2835__));
  and1  g1894(.dina(new_new_n7650__), .dinb(new_new_n7645__), .dout(new_new_n2836__));
  or1   g1895(.dina(new_new_n7652__), .dinb(new_new_n7647__), .dout(new_new_n2837__));
  and1  g1896(.dina(new_new_n2837__), .dinb(new_new_n2835__), .dout(new_new_n2838__));
  or1   g1897(.dina(new_new_n2836__), .dinb(new_new_n2834__), .dout(new_new_n2839__));
  and1  g1898(.dina(new_new_n6970__), .dinb(new_new_n7019__), .dout(new_new_n2840__));
  or1   g1899(.dina(new_new_n6974__), .dinb(new_new_n7034__), .dout(new_new_n2841__));
  and1  g1900(.dina(new_new_n7653__), .dinb(new_new_n7654__), .dout(new_new_n2842__));
  or1   g1901(.dina(new_new_n7655__), .dinb(new_new_n7656__), .dout(new_new_n2843__));
  and1  g1902(.dina(new_new_n7658__), .dinb(new_new_n7654__), .dout(new_new_n2844__));
  or1   g1903(.dina(new_new_n7660__), .dinb(new_new_n7656__), .dout(new_new_n2845__));
  and1  g1904(.dina(new_new_n7658__), .dinb(new_new_n7653__), .dout(new_new_n2846__));
  or1   g1905(.dina(new_new_n7660__), .dinb(new_new_n7655__), .dout(new_new_n2847__));
  and1  g1906(.dina(new_new_n2847__), .dinb(new_new_n2845__), .dout(new_new_n2848__));
  or1   g1907(.dina(new_new_n2846__), .dinb(new_new_n2844__), .dout(new_new_n2849__));
  and1  g1908(.dina(new_new_n2322__), .dinb(new_new_n7077__), .dout(new_new_n2850__));
  or1   g1909(.dina(new_new_n7661__), .dinb(new_new_n7079__), .dout(new_new_n2851__));
  and1  g1910(.dina(new_new_n7662__), .dinb(new_new_n7663__), .dout(new_new_n2852__));
  or1   g1911(.dina(new_new_n7664__), .dinb(new_new_n7665__), .dout(new_new_n2853__));
  and1  g1912(.dina(new_new_n7667__), .dinb(new_new_n7663__), .dout(new_new_n2854__));
  or1   g1913(.dina(new_new_n7669__), .dinb(new_new_n7665__), .dout(new_new_n2855__));
  and1  g1914(.dina(new_new_n7667__), .dinb(new_new_n7662__), .dout(new_new_n2856__));
  or1   g1915(.dina(new_new_n7669__), .dinb(new_new_n7664__), .dout(new_new_n2857__));
  and1  g1916(.dina(new_new_n2857__), .dinb(new_new_n2855__), .dout(new_new_n2858__));
  or1   g1917(.dina(new_new_n2856__), .dinb(new_new_n2854__), .dout(new_new_n2859__));
  and1  g1918(.dina(new_new_n7673__), .dinb(new_new_n6997__), .dout(new_new_n2860__));
  or1   g1919(.dina(new_new_n7688__), .dinb(new_new_n7003__), .dout(new_new_n2861__));
  and1  g1920(.dina(new_new_n7700__), .dinb(new_new_n2803__), .dout(new_new_n2862__));
  or1   g1921(.dina(new_new_n2858__), .dinb(new_new_n7701__), .dout(new_new_n2863__));
  and1  g1922(.dina(new_new_n1586__), .dinb(new_new_n1578__), .dout(new_new_n2864__));
  or1   g1923(.dina(new_new_n1585__), .dinb(new_new_n1577__), .dout(new_new_n2865__));
  and1  g1924(.dina(new_new_n7704__), .dinb(new_new_n7000__), .dout(new_new_n2866__));
  or1   g1925(.dina(new_new_n7710__), .dinb(new_new_n7006__), .dout(new_new_n2867__));
  and1  g1926(.dina(new_new_n7712__), .dinb(new_new_n7713__), .dout(new_new_n2868__));
  or1   g1927(.dina(new_new_n7714__), .dinb(new_new_n7715__), .dout(new_new_n2869__));
  and1  g1928(.dina(new_new_n7717__), .dinb(new_new_n7713__), .dout(new_new_n2870__));
  or1   g1929(.dina(new_new_n7719__), .dinb(new_new_n7715__), .dout(new_new_n2871__));
  and1  g1930(.dina(new_new_n7717__), .dinb(new_new_n7712__), .dout(new_new_n2872__));
  or1   g1931(.dina(new_new_n7719__), .dinb(new_new_n7714__), .dout(new_new_n2873__));
  and1  g1932(.dina(new_new_n2873__), .dinb(new_new_n2871__), .dout(new_new_n2874__));
  or1   g1933(.dina(new_new_n2872__), .dinb(new_new_n2870__), .dout(new_new_n2875__));
  and1  g1934(.dina(new_new_n7116__), .dinb(new_new_n7099__), .dout(new_new_n2876__));
  or1   g1935(.dina(new_new_n7118__), .dinb(new_new_n7101__), .dout(new_new_n2877__));
  and1  g1936(.dina(new_new_n7720__), .dinb(new_new_n7721__), .dout(new_new_n2878__));
  or1   g1937(.dina(new_new_n7722__), .dinb(new_new_n7723__), .dout(new_new_n2879__));
  and1  g1938(.dina(new_new_n7725__), .dinb(new_new_n7721__), .dout(new_new_n2880__));
  or1   g1939(.dina(new_new_n7727__), .dinb(new_new_n7723__), .dout(new_new_n2881__));
  and1  g1940(.dina(new_new_n7725__), .dinb(new_new_n7720__), .dout(new_new_n2882__));
  or1   g1941(.dina(new_new_n7727__), .dinb(new_new_n7722__), .dout(new_new_n2883__));
  and1  g1942(.dina(new_new_n2883__), .dinb(new_new_n2881__), .dout(new_new_n2884__));
  or1   g1943(.dina(new_new_n2882__), .dinb(new_new_n2880__), .dout(new_new_n2885__));
  and1  g1944(.dina(new_new_n7086__), .dinb(new_new_n7105__), .dout(new_new_n2886__));
  or1   g1945(.dina(new_new_n7094__), .dinb(new_new_n7110__), .dout(new_new_n2887__));
  and1  g1946(.dina(new_new_n7728__), .dinb(new_new_n7729__), .dout(new_new_n2888__));
  or1   g1947(.dina(new_new_n7730__), .dinb(new_new_n7731__), .dout(new_new_n2889__));
  and1  g1948(.dina(new_new_n7733__), .dinb(new_new_n7729__), .dout(new_new_n2890__));
  or1   g1949(.dina(new_new_n7735__), .dinb(new_new_n7731__), .dout(new_new_n2891__));
  and1  g1950(.dina(new_new_n7733__), .dinb(new_new_n7728__), .dout(new_new_n2892__));
  or1   g1951(.dina(new_new_n7735__), .dinb(new_new_n7730__), .dout(new_new_n2893__));
  and1  g1952(.dina(new_new_n2893__), .dinb(new_new_n2891__), .dout(new_new_n2894__));
  or1   g1953(.dina(new_new_n2892__), .dinb(new_new_n2890__), .dout(new_new_n2895__));
  and1  g1954(.dina(new_new_n2801__), .dinb(new_new_n7125__), .dout(new_new_n2896__));
  or1   g1955(.dina(new_new_n7736__), .dinb(new_new_n7127__), .dout(new_new_n2897__));
  and1  g1956(.dina(new_new_n7737__), .dinb(new_new_n7738__), .dout(new_new_n2898__));
  or1   g1957(.dina(new_new_n7739__), .dinb(new_new_n7740__), .dout(new_new_n2899__));
  and1  g1958(.dina(new_new_n7742__), .dinb(new_new_n7738__), .dout(new_new_n2900__));
  or1   g1959(.dina(new_new_n7744__), .dinb(new_new_n7740__), .dout(new_new_n2901__));
  and1  g1960(.dina(new_new_n7742__), .dinb(new_new_n7737__), .dout(new_new_n2902__));
  or1   g1961(.dina(new_new_n7744__), .dinb(new_new_n7739__), .dout(new_new_n2903__));
  and1  g1962(.dina(new_new_n2903__), .dinb(new_new_n2901__), .dout(new_new_n2904__));
  or1   g1963(.dina(new_new_n2902__), .dinb(new_new_n2900__), .dout(new_new_n2905__));
  and1  g1964(.dina(new_new_n7745__), .dinb(new_new_n2861__), .dout(new_new_n2906__));
  or1   g1965(.dina(new_new_n2904__), .dinb(new_new_n7746__), .dout(new_new_n2907__));
  or1   g1966(.dina(new_new_n7748__), .dinb(new_new_n2795__), .dout(new_new_n2908__));
  and1  g1967(.dina(new_new_n6737__), .dinb(new_new_n7136__), .dout(new_new_n2909__));
  or1   g1968(.dina(new_new_n6751__), .dinb(new_new_n7142__), .dout(new_new_n2910__));
  and1  g1969(.dina(new_new_n7188__), .dinb(new_new_n7180__), .dout(new_new_n2911__));
  or1   g1970(.dina(new_new_n7190__), .dinb(new_new_n7182__), .dout(new_new_n2912__));
  or1   g1971(.dina(new_new_n2911__), .dinb(new_new_n2909__), .dout(new_new_n2913__));
  and1  g1972(.dina(new_new_n7214__), .dinb(new_new_n7210__), .dout(new_new_n2914__));
  or1   g1973(.dina(new_new_n7216__), .dinb(new_new_n7212__), .dout(new_new_n2915__));
  and1  g1974(.dina(new_new_n7213__), .dinb(new_new_n7209__), .dout(new_new_n2916__));
  or1   g1975(.dina(new_new_n7215__), .dinb(new_new_n7211__), .dout(new_new_n2917__));
  and1  g1976(.dina(new_new_n2917__), .dinb(new_new_n2915__), .dout(new_new_n2918__));
  or1   g1977(.dina(new_new_n2916__), .dinb(new_new_n2914__), .dout(new_new_n2919__));
  and1  g1978(.dina(new_new_n7254__), .dinb(new_new_n7241__), .dout(new_new_n2920__));
  or1   g1979(.dina(new_new_n7256__), .dinb(new_new_n7243__), .dout(new_new_n2921__));
  and1  g1980(.dina(new_new_n7749__), .dinb(new_new_n7750__), .dout(new_new_n2922__));
  or1   g1981(.dina(new_new_n7751__), .dinb(new_new_n7752__), .dout(new_new_n2923__));
  and1  g1982(.dina(new_new_n7754__), .dinb(new_new_n7750__), .dout(new_new_n2924__));
  or1   g1983(.dina(new_new_n7756__), .dinb(new_new_n7752__), .dout(new_new_n2925__));
  and1  g1984(.dina(new_new_n7754__), .dinb(new_new_n7749__), .dout(new_new_n2926__));
  or1   g1985(.dina(new_new_n7756__), .dinb(new_new_n7751__), .dout(new_new_n2927__));
  and1  g1986(.dina(new_new_n2927__), .dinb(new_new_n2925__), .dout(new_new_n2928__));
  or1   g1987(.dina(new_new_n2926__), .dinb(new_new_n2924__), .dout(new_new_n2929__));
  and1  g1988(.dina(new_new_n6737__), .dinb(new_new_n7246__), .dout(new_new_n2930__));
  or1   g1989(.dina(new_new_n6751__), .dinb(new_new_n7249__), .dout(new_new_n2931__));
  and1  g1990(.dina(new_new_n7757__), .dinb(new_new_n7758__), .dout(new_new_n2932__));
  or1   g1991(.dina(new_new_n7759__), .dinb(new_new_n7760__), .dout(new_new_n2933__));
  and1  g1992(.dina(new_new_n7762__), .dinb(new_new_n7758__), .dout(new_new_n2934__));
  or1   g1993(.dina(new_new_n7764__), .dinb(new_new_n7760__), .dout(new_new_n2935__));
  and1  g1994(.dina(new_new_n7762__), .dinb(new_new_n7757__), .dout(new_new_n2936__));
  or1   g1995(.dina(new_new_n7764__), .dinb(new_new_n7759__), .dout(new_new_n2937__));
  and1  g1996(.dina(new_new_n2937__), .dinb(new_new_n2935__), .dout(new_new_n2938__));
  or1   g1997(.dina(new_new_n2936__), .dinb(new_new_n2934__), .dout(new_new_n2939__));
  and1  g1998(.dina(new_new_n7291__), .dinb(new_new_n7283__), .dout(new_new_n2940__));
  or1   g1999(.dina(new_new_n7293__), .dinb(new_new_n7285__), .dout(new_new_n2941__));
  and1  g2000(.dina(new_new_n7765__), .dinb(new_new_n7766__), .dout(new_new_n2942__));
  or1   g2001(.dina(new_new_n7767__), .dinb(new_new_n7768__), .dout(new_new_n2943__));
  and1  g2002(.dina(new_new_n7770__), .dinb(new_new_n7766__), .dout(new_new_n2944__));
  or1   g2003(.dina(new_new_n7772__), .dinb(new_new_n7768__), .dout(new_new_n2945__));
  and1  g2004(.dina(new_new_n7770__), .dinb(new_new_n7765__), .dout(new_new_n2946__));
  or1   g2005(.dina(new_new_n7772__), .dinb(new_new_n7767__), .dout(new_new_n2947__));
  and1  g2006(.dina(new_new_n2947__), .dinb(new_new_n2945__), .dout(new_new_n2948__));
  or1   g2007(.dina(new_new_n2946__), .dinb(new_new_n2944__), .dout(new_new_n2949__));
  and1  g2008(.dina(new_new_n7268__), .dinb(new_new_n6767__), .dout(new_new_n2950__));
  or1   g2009(.dina(new_new_n7269__), .dinb(new_new_n6781__), .dout(new_new_n2951__));
  and1  g2010(.dina(new_new_n7773__), .dinb(new_new_n7774__), .dout(new_new_n2952__));
  or1   g2011(.dina(new_new_n7775__), .dinb(new_new_n7776__), .dout(new_new_n2953__));
  and1  g2012(.dina(new_new_n7778__), .dinb(new_new_n7774__), .dout(new_new_n2954__));
  or1   g2013(.dina(new_new_n7780__), .dinb(new_new_n7776__), .dout(new_new_n2955__));
  and1  g2014(.dina(new_new_n7778__), .dinb(new_new_n7773__), .dout(new_new_n2956__));
  or1   g2015(.dina(new_new_n7780__), .dinb(new_new_n7775__), .dout(new_new_n2957__));
  and1  g2016(.dina(new_new_n2957__), .dinb(new_new_n2955__), .dout(new_new_n2958__));
  or1   g2017(.dina(new_new_n2956__), .dinb(new_new_n2954__), .dout(new_new_n2959__));
  and1  g2018(.dina(new_new_n7337__), .dinb(new_new_n7329__), .dout(new_new_n2960__));
  or1   g2019(.dina(new_new_n7339__), .dinb(new_new_n7331__), .dout(new_new_n2961__));
  or1   g2020(.dina(new_new_n2960__), .dinb(new_new_n2958__), .dout(new_new_n2962__));
  and1  g2021(.dina(new_new_n7363__), .dinb(new_new_n7359__), .dout(new_new_n2963__));
  or1   g2022(.dina(new_new_n7365__), .dinb(new_new_n7361__), .dout(new_new_n2964__));
  and1  g2023(.dina(new_new_n7362__), .dinb(new_new_n7358__), .dout(new_new_n2965__));
  or1   g2024(.dina(new_new_n7364__), .dinb(new_new_n7360__), .dout(new_new_n2966__));
  and1  g2025(.dina(new_new_n2966__), .dinb(new_new_n2964__), .dout(new_new_n2967__));
  or1   g2026(.dina(new_new_n2965__), .dinb(new_new_n2963__), .dout(new_new_n2968__));
  and1  g2027(.dina(new_new_n7403__), .dinb(new_new_n7390__), .dout(new_new_n2969__));
  or1   g2028(.dina(new_new_n7405__), .dinb(new_new_n7392__), .dout(new_new_n2970__));
  and1  g2029(.dina(new_new_n7781__), .dinb(new_new_n7782__), .dout(new_new_n2971__));
  or1   g2030(.dina(new_new_n7783__), .dinb(new_new_n7784__), .dout(new_new_n2972__));
  and1  g2031(.dina(new_new_n7786__), .dinb(new_new_n7782__), .dout(new_new_n2973__));
  or1   g2032(.dina(new_new_n7788__), .dinb(new_new_n7784__), .dout(new_new_n2974__));
  and1  g2033(.dina(new_new_n7786__), .dinb(new_new_n7781__), .dout(new_new_n2975__));
  or1   g2034(.dina(new_new_n7788__), .dinb(new_new_n7783__), .dout(new_new_n2976__));
  and1  g2035(.dina(new_new_n2976__), .dinb(new_new_n2974__), .dout(new_new_n2977__));
  or1   g2036(.dina(new_new_n2975__), .dinb(new_new_n2973__), .dout(new_new_n2978__));
  and1  g2037(.dina(new_new_n7395__), .dinb(new_new_n6768__), .dout(new_new_n2979__));
  or1   g2038(.dina(new_new_n7398__), .dinb(new_new_n6782__), .dout(new_new_n2980__));
  and1  g2039(.dina(new_new_n7789__), .dinb(new_new_n7790__), .dout(new_new_n2981__));
  or1   g2040(.dina(new_new_n7791__), .dinb(new_new_n7792__), .dout(new_new_n2982__));
  and1  g2041(.dina(new_new_n7794__), .dinb(new_new_n7790__), .dout(new_new_n2983__));
  or1   g2042(.dina(new_new_n7796__), .dinb(new_new_n7792__), .dout(new_new_n2984__));
  and1  g2043(.dina(new_new_n7794__), .dinb(new_new_n7789__), .dout(new_new_n2985__));
  or1   g2044(.dina(new_new_n7796__), .dinb(new_new_n7791__), .dout(new_new_n2986__));
  and1  g2045(.dina(new_new_n2986__), .dinb(new_new_n2984__), .dout(new_new_n2987__));
  or1   g2046(.dina(new_new_n2985__), .dinb(new_new_n2983__), .dout(new_new_n2988__));
  and1  g2047(.dina(new_new_n7440__), .dinb(new_new_n7432__), .dout(new_new_n2989__));
  or1   g2048(.dina(new_new_n7442__), .dinb(new_new_n7434__), .dout(new_new_n2990__));
  and1  g2049(.dina(new_new_n7797__), .dinb(new_new_n7798__), .dout(new_new_n2991__));
  or1   g2050(.dina(new_new_n7799__), .dinb(new_new_n7800__), .dout(new_new_n2992__));
  and1  g2051(.dina(new_new_n7802__), .dinb(new_new_n7798__), .dout(new_new_n2993__));
  or1   g2052(.dina(new_new_n7804__), .dinb(new_new_n7800__), .dout(new_new_n2994__));
  and1  g2053(.dina(new_new_n7802__), .dinb(new_new_n7797__), .dout(new_new_n2995__));
  or1   g2054(.dina(new_new_n7804__), .dinb(new_new_n7799__), .dout(new_new_n2996__));
  and1  g2055(.dina(new_new_n2996__), .dinb(new_new_n2994__), .dout(new_new_n2997__));
  or1   g2056(.dina(new_new_n2995__), .dinb(new_new_n2993__), .dout(new_new_n2998__));
  and1  g2057(.dina(new_new_n7417__), .dinb(new_new_n6810__), .dout(new_new_n2999__));
  or1   g2058(.dina(new_new_n7418__), .dinb(new_new_n6820__), .dout(new_new_n3000__));
  and1  g2059(.dina(new_new_n7805__), .dinb(new_new_n7806__), .dout(new_new_n3001__));
  or1   g2060(.dina(new_new_n7807__), .dinb(new_new_n7808__), .dout(new_new_n3002__));
  and1  g2061(.dina(new_new_n7810__), .dinb(new_new_n7806__), .dout(new_new_n3003__));
  or1   g2062(.dina(new_new_n7812__), .dinb(new_new_n7808__), .dout(new_new_n3004__));
  and1  g2063(.dina(new_new_n7810__), .dinb(new_new_n7805__), .dout(new_new_n3005__));
  or1   g2064(.dina(new_new_n7812__), .dinb(new_new_n7807__), .dout(new_new_n3006__));
  and1  g2065(.dina(new_new_n3006__), .dinb(new_new_n3004__), .dout(new_new_n3007__));
  or1   g2066(.dina(new_new_n3005__), .dinb(new_new_n3003__), .dout(new_new_n3008__));
  and1  g2067(.dina(new_new_n7485__), .dinb(new_new_n7477__), .dout(new_new_n3009__));
  or1   g2068(.dina(new_new_n7487__), .dinb(new_new_n7479__), .dout(new_new_n3010__));
  or1   g2069(.dina(new_new_n3009__), .dinb(new_new_n3007__), .dout(new_new_n3011__));
  and1  g2070(.dina(new_new_n7510__), .dinb(new_new_n7506__), .dout(new_new_n3012__));
  or1   g2071(.dina(new_new_n7512__), .dinb(new_new_n7508__), .dout(new_new_n3013__));
  and1  g2072(.dina(new_new_n7509__), .dinb(new_new_n7505__), .dout(new_new_n3014__));
  or1   g2073(.dina(new_new_n7511__), .dinb(new_new_n7507__), .dout(new_new_n3015__));
  and1  g2074(.dina(new_new_n3015__), .dinb(new_new_n3013__), .dout(new_new_n3016__));
  or1   g2075(.dina(new_new_n3014__), .dinb(new_new_n3012__), .dout(new_new_n3017__));
  and1  g2076(.dina(new_new_n7490__), .dinb(new_new_n1381__), .dout(new_new_n3018__));
  or1   g2077(.dina(new_new_n7492__), .dinb(new_new_n1382__), .dout(new_new_n3019__));
  and1  g2078(.dina(new_new_n7489__), .dinb(new_new_n1334__), .dout(new_new_n3020__));
  or1   g2079(.dina(new_new_n7491__), .dinb(new_new_n1333__), .dout(new_new_n3021__));
  and1  g2080(.dina(new_new_n3021__), .dinb(new_new_n3019__), .dout(new_new_n3022__));
  or1   g2081(.dina(new_new_n3020__), .dinb(new_new_n3018__), .dout(new_new_n3023__));
  and1  g2082(.dina(new_new_n1310__), .dinb(new_new_n1247__), .dout(new_new_n3024__));
  or1   g2083(.dina(new_new_n1309__), .dinb(new_new_n1248__), .dout(new_new_n3025__));
  and1  g2084(.dina(new_new_n7813__), .dinb(new_new_n7814__), .dout(new_new_n3026__));
  or1   g2085(.dina(new_new_n7815__), .dinb(new_new_n7816__), .dout(new_new_n3027__));
  and1  g2086(.dina(new_new_n7818__), .dinb(new_new_n7814__), .dout(new_new_n3028__));
  or1   g2087(.dina(new_new_n7820__), .dinb(new_new_n7816__), .dout(new_new_n3029__));
  and1  g2088(.dina(new_new_n7818__), .dinb(new_new_n7813__), .dout(new_new_n3030__));
  or1   g2089(.dina(new_new_n7820__), .dinb(new_new_n7815__), .dout(new_new_n3031__));
  and1  g2090(.dina(new_new_n3031__), .dinb(new_new_n3029__), .dout(new_new_n3032__));
  or1   g2091(.dina(new_new_n3030__), .dinb(new_new_n3028__), .dout(new_new_n3033__));
  and1  g2092(.dina(new_new_n7822__), .dinb(new_new_n6768__), .dout(new_new_n3034__));
  or1   g2093(.dina(new_new_n7824__), .dinb(new_new_n6782__), .dout(new_new_n3035__));
  and1  g2094(.dina(new_new_n7825__), .dinb(new_new_n7826__), .dout(new_new_n3036__));
  or1   g2095(.dina(new_new_n7827__), .dinb(new_new_n7828__), .dout(new_new_n3037__));
  and1  g2096(.dina(new_new_n7830__), .dinb(new_new_n7817__), .dout(new_new_n3038__));
  or1   g2097(.dina(new_new_n7832__), .dinb(new_new_n7819__), .dout(new_new_n3039__));
  and1  g2098(.dina(new_new_n7833__), .dinb(new_new_n7834__), .dout(new_new_n3040__));
  or1   g2099(.dina(new_new_n7835__), .dinb(new_new_n7836__), .dout(new_new_n3041__));
  and1  g2100(.dina(new_new_n7838__), .dinb(new_new_n7834__), .dout(new_new_n3042__));
  or1   g2101(.dina(new_new_n7840__), .dinb(new_new_n7836__), .dout(new_new_n3043__));
  and1  g2102(.dina(new_new_n7838__), .dinb(new_new_n7833__), .dout(new_new_n3044__));
  or1   g2103(.dina(new_new_n7840__), .dinb(new_new_n7835__), .dout(new_new_n3045__));
  and1  g2104(.dina(new_new_n3045__), .dinb(new_new_n3043__), .dout(new_new_n3046__));
  or1   g2105(.dina(new_new_n3044__), .dinb(new_new_n3042__), .dout(new_new_n3047__));
  and1  g2106(.dina(new_new_n7822__), .dinb(new_new_n6809__), .dout(new_new_n3048__));
  or1   g2107(.dina(new_new_n7824__), .dinb(new_new_n6819__), .dout(new_new_n3049__));
  and1  g2108(.dina(new_new_n7841__), .dinb(new_new_n7842__), .dout(new_new_n3050__));
  or1   g2109(.dina(new_new_n7843__), .dinb(new_new_n7844__), .dout(new_new_n3051__));
  and1  g2110(.dina(new_new_n7846__), .dinb(new_new_n7842__), .dout(new_new_n3052__));
  or1   g2111(.dina(new_new_n7848__), .dinb(new_new_n7844__), .dout(new_new_n3053__));
  and1  g2112(.dina(new_new_n7846__), .dinb(new_new_n7841__), .dout(new_new_n3054__));
  or1   g2113(.dina(new_new_n7848__), .dinb(new_new_n7843__), .dout(new_new_n3055__));
  and1  g2114(.dina(new_new_n3055__), .dinb(new_new_n3053__), .dout(new_new_n3056__));
  or1   g2115(.dina(new_new_n3054__), .dinb(new_new_n3052__), .dout(new_new_n3057__));
  and1  g2116(.dina(new_new_n7830__), .dinb(new_new_n7826__), .dout(new_new_n3058__));
  or1   g2117(.dina(new_new_n7832__), .dinb(new_new_n7828__), .dout(new_new_n3059__));
  and1  g2118(.dina(new_new_n7829__), .dinb(new_new_n7825__), .dout(new_new_n3060__));
  or1   g2119(.dina(new_new_n7831__), .dinb(new_new_n7827__), .dout(new_new_n3061__));
  and1  g2120(.dina(new_new_n3061__), .dinb(new_new_n3059__), .dout(new_new_n3062__));
  or1   g2121(.dina(new_new_n3060__), .dinb(new_new_n3058__), .dout(new_new_n3063__));
  and1  g2122(.dina(new_new_n7549__), .dinb(new_new_n7537__), .dout(new_new_n3064__));
  or1   g2123(.dina(new_new_n7551__), .dinb(new_new_n7539__), .dout(new_new_n3065__));
  and1  g2124(.dina(new_new_n7849__), .dinb(new_new_n7850__), .dout(new_new_n3066__));
  or1   g2125(.dina(new_new_n7851__), .dinb(new_new_n7852__), .dout(new_new_n3067__));
  and1  g2126(.dina(new_new_n7854__), .dinb(new_new_n7850__), .dout(new_new_n3068__));
  or1   g2127(.dina(new_new_n7856__), .dinb(new_new_n7852__), .dout(new_new_n3069__));
  and1  g2128(.dina(new_new_n7854__), .dinb(new_new_n7849__), .dout(new_new_n3070__));
  or1   g2129(.dina(new_new_n7856__), .dinb(new_new_n7851__), .dout(new_new_n3071__));
  and1  g2130(.dina(new_new_n3071__), .dinb(new_new_n3069__), .dout(new_new_n3072__));
  or1   g2131(.dina(new_new_n3070__), .dinb(new_new_n3068__), .dout(new_new_n3073__));
  and1  g2132(.dina(new_new_n7542__), .dinb(new_new_n6812__), .dout(new_new_n3074__));
  or1   g2133(.dina(new_new_n7544__), .dinb(new_new_n6822__), .dout(new_new_n3075__));
  and1  g2134(.dina(new_new_n7857__), .dinb(new_new_n7858__), .dout(new_new_n3076__));
  or1   g2135(.dina(new_new_n7859__), .dinb(new_new_n7860__), .dout(new_new_n3077__));
  and1  g2136(.dina(new_new_n7862__), .dinb(new_new_n7853__), .dout(new_new_n3078__));
  or1   g2137(.dina(new_new_n7864__), .dinb(new_new_n7855__), .dout(new_new_n3079__));
  and1  g2138(.dina(new_new_n7865__), .dinb(new_new_n7866__), .dout(new_new_n3080__));
  or1   g2139(.dina(new_new_n7867__), .dinb(new_new_n7868__), .dout(new_new_n3081__));
  and1  g2140(.dina(new_new_n7870__), .dinb(new_new_n7866__), .dout(new_new_n3082__));
  or1   g2141(.dina(new_new_n7872__), .dinb(new_new_n7868__), .dout(new_new_n3083__));
  and1  g2142(.dina(new_new_n7870__), .dinb(new_new_n7865__), .dout(new_new_n3084__));
  or1   g2143(.dina(new_new_n7872__), .dinb(new_new_n7867__), .dout(new_new_n3085__));
  and1  g2144(.dina(new_new_n3085__), .dinb(new_new_n3083__), .dout(new_new_n3086__));
  or1   g2145(.dina(new_new_n3084__), .dinb(new_new_n3082__), .dout(new_new_n3087__));
  and1  g2146(.dina(new_new_n7541__), .dinb(new_new_n6885__), .dout(new_new_n3088__));
  or1   g2147(.dina(new_new_n7543__), .dinb(new_new_n6891__), .dout(new_new_n3089__));
  and1  g2148(.dina(new_new_n7873__), .dinb(new_new_n7874__), .dout(new_new_n3090__));
  or1   g2149(.dina(new_new_n7875__), .dinb(new_new_n7876__), .dout(new_new_n3091__));
  and1  g2150(.dina(new_new_n7878__), .dinb(new_new_n7874__), .dout(new_new_n3092__));
  or1   g2151(.dina(new_new_n7880__), .dinb(new_new_n7876__), .dout(new_new_n3093__));
  and1  g2152(.dina(new_new_n7878__), .dinb(new_new_n7873__), .dout(new_new_n3094__));
  or1   g2153(.dina(new_new_n7880__), .dinb(new_new_n7875__), .dout(new_new_n3095__));
  and1  g2154(.dina(new_new_n3095__), .dinb(new_new_n3093__), .dout(new_new_n3096__));
  or1   g2155(.dina(new_new_n3094__), .dinb(new_new_n3092__), .dout(new_new_n3097__));
  and1  g2156(.dina(new_new_n7862__), .dinb(new_new_n7858__), .dout(new_new_n3098__));
  or1   g2157(.dina(new_new_n7864__), .dinb(new_new_n7860__), .dout(new_new_n3099__));
  and1  g2158(.dina(new_new_n7861__), .dinb(new_new_n7857__), .dout(new_new_n3100__));
  or1   g2159(.dina(new_new_n7863__), .dinb(new_new_n7859__), .dout(new_new_n3101__));
  and1  g2160(.dina(new_new_n3101__), .dinb(new_new_n3099__), .dout(new_new_n3102__));
  or1   g2161(.dina(new_new_n3100__), .dinb(new_new_n3098__), .dout(new_new_n3103__));
  and1  g2162(.dina(new_new_n7565__), .dinb(new_new_n7557__), .dout(new_new_n3104__));
  or1   g2163(.dina(new_new_n7567__), .dinb(new_new_n7559__), .dout(new_new_n3105__));
  and1  g2164(.dina(new_new_n7881__), .dinb(new_new_n7882__), .dout(new_new_n3106__));
  or1   g2165(.dina(new_new_n7883__), .dinb(new_new_n7884__), .dout(new_new_n3107__));
  and1  g2166(.dina(new_new_n7886__), .dinb(new_new_n7882__), .dout(new_new_n3108__));
  or1   g2167(.dina(new_new_n7888__), .dinb(new_new_n7884__), .dout(new_new_n3109__));
  and1  g2168(.dina(new_new_n7886__), .dinb(new_new_n7881__), .dout(new_new_n3110__));
  or1   g2169(.dina(new_new_n7888__), .dinb(new_new_n7883__), .dout(new_new_n3111__));
  and1  g2170(.dina(new_new_n3111__), .dinb(new_new_n3109__), .dout(new_new_n3112__));
  or1   g2171(.dina(new_new_n3110__), .dinb(new_new_n3108__), .dout(new_new_n3113__));
  and1  g2172(.dina(new_new_n6902__), .dinb(new_new_n6885__), .dout(new_new_n3114__));
  or1   g2173(.dina(new_new_n6904__), .dinb(new_new_n6891__), .dout(new_new_n3115__));
  and1  g2174(.dina(new_new_n7889__), .dinb(new_new_n7890__), .dout(new_new_n3116__));
  or1   g2175(.dina(new_new_n7891__), .dinb(new_new_n7892__), .dout(new_new_n3117__));
  and1  g2176(.dina(new_new_n7894__), .dinb(new_new_n7885__), .dout(new_new_n3118__));
  or1   g2177(.dina(new_new_n7896__), .dinb(new_new_n7887__), .dout(new_new_n3119__));
  or1   g2178(.dina(new_new_n3118__), .dinb(new_new_n3096__), .dout(new_new_n3120__));
  and1  g2179(.dina(new_new_n7894__), .dinb(new_new_n7890__), .dout(new_new_n3121__));
  or1   g2180(.dina(new_new_n7896__), .dinb(new_new_n7892__), .dout(new_new_n3122__));
  and1  g2181(.dina(new_new_n7893__), .dinb(new_new_n7889__), .dout(new_new_n3123__));
  or1   g2182(.dina(new_new_n7895__), .dinb(new_new_n7891__), .dout(new_new_n3124__));
  and1  g2183(.dina(new_new_n3124__), .dinb(new_new_n3122__), .dout(new_new_n3125__));
  or1   g2184(.dina(new_new_n3123__), .dinb(new_new_n3121__), .dout(new_new_n3126__));
  and1  g2185(.dina(new_new_n7581__), .dinb(new_new_n7573__), .dout(new_new_n3127__));
  or1   g2186(.dina(new_new_n7583__), .dinb(new_new_n7575__), .dout(new_new_n3128__));
  and1  g2187(.dina(new_new_n7897__), .dinb(new_new_n7898__), .dout(new_new_n3129__));
  or1   g2188(.dina(new_new_n3127__), .dinb(new_new_n3125__), .dout(new_new_n3130__));
  and1  g2189(.dina(new_new_n7899__), .dinb(new_new_n7898__), .dout(new_new_n3131__));
  and1  g2190(.dina(new_new_n7899__), .dinb(new_new_n7897__), .dout(new_new_n3132__));
  or1   g2191(.dina(new_new_n3132__), .dinb(new_new_n3131__), .dout(new_new_n3133__));
  and1  g2192(.dina(new_new_n6999__), .dinb(new_new_n7903__), .dout(new_new_n3134__));
  or1   g2193(.dina(new_new_n7005__), .dinb(new_new_n7918__), .dout(new_new_n3135__));
  and1  g2194(.dina(new_new_n7931__), .dinb(new_new_n7530__), .dout(new_new_n3136__));
  or1   g2195(.dina(new_new_n7932__), .dinb(new_new_n7532__), .dout(new_new_n3137__));
  and1  g2196(.dina(new_new_n7931__), .dinb(new_new_n7529__), .dout(new_new_n3138__));
  or1   g2197(.dina(new_new_n7932__), .dinb(new_new_n7531__), .dout(new_new_n3139__));
  and1  g2198(.dina(new_new_n3139__), .dinb(new_new_n3137__), .dout(new_new_n3140__));
  or1   g2199(.dina(new_new_n3138__), .dinb(new_new_n3136__), .dout(new_new_n3141__));
  and1  g2200(.dina(new_new_n7501__), .dinb(new_new_n6887__), .dout(new_new_n3142__));
  or1   g2201(.dina(new_new_n7503__), .dinb(new_new_n6893__), .dout(new_new_n3143__));
  or1   g2202(.dina(new_new_n3142__), .dinb(new_new_n3140__), .dout(new_new_n3144__));
  and1  g2203(.dina(new_new_n7934__), .dinb(new_new_n7383__), .dout(new_new_n3145__));
  or1   g2204(.dina(new_new_n7935__), .dinb(new_new_n7385__), .dout(new_new_n3146__));
  and1  g2205(.dina(new_new_n7934__), .dinb(new_new_n7382__), .dout(new_new_n3147__));
  or1   g2206(.dina(new_new_n7935__), .dinb(new_new_n7384__), .dout(new_new_n3148__));
  and1  g2207(.dina(new_new_n3148__), .dinb(new_new_n3146__), .dout(new_new_n3149__));
  or1   g2208(.dina(new_new_n3147__), .dinb(new_new_n3145__), .dout(new_new_n3150__));
  and1  g2209(.dina(new_new_n7355__), .dinb(new_new_n6812__), .dout(new_new_n3151__));
  or1   g2210(.dina(new_new_n7356__), .dinb(new_new_n6822__), .dout(new_new_n3152__));
  or1   g2211(.dina(new_new_n3151__), .dinb(new_new_n3149__), .dout(new_new_n3153__));
  and1  g2212(.dina(new_new_n7937__), .dinb(new_new_n7234__), .dout(new_new_n3154__));
  or1   g2213(.dina(new_new_n7938__), .dinb(new_new_n7236__), .dout(new_new_n3155__));
  and1  g2214(.dina(new_new_n7937__), .dinb(new_new_n7233__), .dout(new_new_n3156__));
  or1   g2215(.dina(new_new_n7938__), .dinb(new_new_n7235__), .dout(new_new_n3157__));
  and1  g2216(.dina(new_new_n3157__), .dinb(new_new_n3155__), .dout(new_new_n3158__));
  or1   g2217(.dina(new_new_n3156__), .dinb(new_new_n3154__), .dout(new_new_n3159__));
  and1  g2218(.dina(new_new_n7206__), .dinb(new_new_n6770__), .dout(new_new_n3160__));
  or1   g2219(.dina(new_new_n7207__), .dinb(new_new_n6784__), .dout(new_new_n3161__));
  or1   g2220(.dina(new_new_n3160__), .dinb(new_new_n3158__), .dout(new_new_n3162__));
  and1  g2221(.dina(new_new_n7939__), .dinb(new_new_n7940__), .dout(new_new_n3163__));
  and1  g2222(.dina(new_new_n6860__), .dinb(new_new_n7942__), .dout(new_new_n3164__));
  or1   g2223(.dina(new_new_n6869__), .dinb(new_new_n7945__), .dout(new_new_n3165__));
  and1  g2224(.dina(new_new_n7946__), .dinb(new_new_n7947__), .dout(new_new_n3166__));
  or1   g2225(.dina(new_new_n7948__), .dinb(new_new_n7949__), .dout(new_new_n3167__));
  and1  g2226(.dina(new_new_n7951__), .dinb(new_new_n7947__), .dout(new_new_n3168__));
  or1   g2227(.dina(new_new_n7953__), .dinb(new_new_n7949__), .dout(new_new_n3169__));
  and1  g2228(.dina(new_new_n7951__), .dinb(new_new_n7946__), .dout(new_new_n3170__));
  or1   g2229(.dina(new_new_n7953__), .dinb(new_new_n7948__), .dout(new_new_n3171__));
  and1  g2230(.dina(new_new_n3171__), .dinb(new_new_n3169__), .dout(new_new_n3172__));
  or1   g2231(.dina(new_new_n3170__), .dinb(new_new_n3168__), .dout(new_new_n3173__));
  and1  g2232(.dina(new_new_n6862__), .dinb(new_new_n7955__), .dout(new_new_n3174__));
  or1   g2233(.dina(new_new_n6871__), .dinb(new_new_n7958__), .dout(new_new_n3175__));
  and1  g2234(.dina(new_new_n7959__), .dinb(new_new_n7960__), .dout(new_new_n3176__));
  or1   g2235(.dina(new_new_n7961__), .dinb(new_new_n7962__), .dout(new_new_n3177__));
  and1  g2236(.dina(new_new_n7964__), .dinb(new_new_n7950__), .dout(new_new_n3178__));
  or1   g2237(.dina(new_new_n7966__), .dinb(new_new_n7952__), .dout(new_new_n3179__));
  and1  g2238(.dina(new_new_n7967__), .dinb(new_new_n7968__), .dout(new_new_n3180__));
  or1   g2239(.dina(new_new_n7969__), .dinb(new_new_n7970__), .dout(new_new_n3181__));
  and1  g2240(.dina(new_new_n7972__), .dinb(new_new_n7968__), .dout(new_new_n3182__));
  or1   g2241(.dina(new_new_n7974__), .dinb(new_new_n7970__), .dout(new_new_n3183__));
  and1  g2242(.dina(new_new_n7972__), .dinb(new_new_n7967__), .dout(new_new_n3184__));
  or1   g2243(.dina(new_new_n7974__), .dinb(new_new_n7969__), .dout(new_new_n3185__));
  and1  g2244(.dina(new_new_n3185__), .dinb(new_new_n3183__), .dout(new_new_n3186__));
  or1   g2245(.dina(new_new_n3184__), .dinb(new_new_n3182__), .dout(new_new_n3187__));
  and1  g2246(.dina(new_new_n6943__), .dinb(new_new_n7955__), .dout(new_new_n3188__));
  or1   g2247(.dina(new_new_n6956__), .dinb(new_new_n7958__), .dout(new_new_n3189__));
  and1  g2248(.dina(new_new_n7975__), .dinb(new_new_n7976__), .dout(new_new_n3190__));
  or1   g2249(.dina(new_new_n7977__), .dinb(new_new_n7978__), .dout(new_new_n3191__));
  and1  g2250(.dina(new_new_n7980__), .dinb(new_new_n7976__), .dout(new_new_n3192__));
  or1   g2251(.dina(new_new_n7982__), .dinb(new_new_n7978__), .dout(new_new_n3193__));
  and1  g2252(.dina(new_new_n7980__), .dinb(new_new_n7975__), .dout(new_new_n3194__));
  or1   g2253(.dina(new_new_n7982__), .dinb(new_new_n7977__), .dout(new_new_n3195__));
  and1  g2254(.dina(new_new_n3195__), .dinb(new_new_n3193__), .dout(new_new_n3196__));
  or1   g2255(.dina(new_new_n3194__), .dinb(new_new_n3192__), .dout(new_new_n3197__));
  and1  g2256(.dina(new_new_n7964__), .dinb(new_new_n7960__), .dout(new_new_n3198__));
  or1   g2257(.dina(new_new_n7966__), .dinb(new_new_n7962__), .dout(new_new_n3199__));
  and1  g2258(.dina(new_new_n7963__), .dinb(new_new_n7959__), .dout(new_new_n3200__));
  or1   g2259(.dina(new_new_n7965__), .dinb(new_new_n7961__), .dout(new_new_n3201__));
  and1  g2260(.dina(new_new_n3201__), .dinb(new_new_n3199__), .dout(new_new_n3202__));
  or1   g2261(.dina(new_new_n3200__), .dinb(new_new_n3198__), .dout(new_new_n3203__));
  and1  g2262(.dina(new_new_n1516__), .dinb(new_new_n1508__), .dout(new_new_n3204__));
  or1   g2263(.dina(new_new_n1515__), .dinb(new_new_n1507__), .dout(new_new_n3205__));
  and1  g2264(.dina(new_new_n6862__), .dinb(new_new_n7984__), .dout(new_new_n3206__));
  or1   g2265(.dina(new_new_n6871__), .dinb(new_new_n7987__), .dout(new_new_n3207__));
  and1  g2266(.dina(new_new_n7989__), .dinb(new_new_n7990__), .dout(new_new_n3208__));
  or1   g2267(.dina(new_new_n7991__), .dinb(new_new_n7992__), .dout(new_new_n3209__));
  and1  g2268(.dina(new_new_n7994__), .dinb(new_new_n1451__), .dout(new_new_n3210__));
  or1   g2269(.dina(new_new_n7996__), .dinb(new_new_n1452__), .dout(new_new_n3211__));
  and1  g2270(.dina(new_new_n7997__), .dinb(new_new_n7998__), .dout(new_new_n3212__));
  or1   g2271(.dina(new_new_n7999__), .dinb(new_new_n8000__), .dout(new_new_n3213__));
  and1  g2272(.dina(new_new_n8002__), .dinb(new_new_n7998__), .dout(new_new_n3214__));
  or1   g2273(.dina(new_new_n8004__), .dinb(new_new_n8000__), .dout(new_new_n3215__));
  and1  g2274(.dina(new_new_n8002__), .dinb(new_new_n7997__), .dout(new_new_n3216__));
  or1   g2275(.dina(new_new_n8004__), .dinb(new_new_n7999__), .dout(new_new_n3217__));
  and1  g2276(.dina(new_new_n3217__), .dinb(new_new_n3215__), .dout(new_new_n3218__));
  or1   g2277(.dina(new_new_n3216__), .dinb(new_new_n3214__), .dout(new_new_n3219__));
  and1  g2278(.dina(new_new_n6945__), .dinb(new_new_n7984__), .dout(new_new_n3220__));
  or1   g2279(.dina(new_new_n6958__), .dinb(new_new_n7987__), .dout(new_new_n3221__));
  and1  g2280(.dina(new_new_n8005__), .dinb(new_new_n8006__), .dout(new_new_n3222__));
  or1   g2281(.dina(new_new_n8007__), .dinb(new_new_n8008__), .dout(new_new_n3223__));
  and1  g2282(.dina(new_new_n8010__), .dinb(new_new_n8001__), .dout(new_new_n3224__));
  or1   g2283(.dina(new_new_n8012__), .dinb(new_new_n8003__), .dout(new_new_n3225__));
  and1  g2284(.dina(new_new_n8013__), .dinb(new_new_n8014__), .dout(new_new_n3226__));
  or1   g2285(.dina(new_new_n8015__), .dinb(new_new_n8016__), .dout(new_new_n3227__));
  and1  g2286(.dina(new_new_n8018__), .dinb(new_new_n8014__), .dout(new_new_n3228__));
  or1   g2287(.dina(new_new_n8020__), .dinb(new_new_n8016__), .dout(new_new_n3229__));
  and1  g2288(.dina(new_new_n8018__), .dinb(new_new_n8013__), .dout(new_new_n3230__));
  or1   g2289(.dina(new_new_n8020__), .dinb(new_new_n8015__), .dout(new_new_n3231__));
  and1  g2290(.dina(new_new_n3231__), .dinb(new_new_n3229__), .dout(new_new_n3232__));
  or1   g2291(.dina(new_new_n3230__), .dinb(new_new_n3228__), .dout(new_new_n3233__));
  and1  g2292(.dina(new_new_n7985__), .dinb(new_new_n7020__), .dout(new_new_n3234__));
  or1   g2293(.dina(new_new_n7988__), .dinb(new_new_n7035__), .dout(new_new_n3235__));
  and1  g2294(.dina(new_new_n8021__), .dinb(new_new_n8022__), .dout(new_new_n3236__));
  or1   g2295(.dina(new_new_n8023__), .dinb(new_new_n8024__), .dout(new_new_n3237__));
  and1  g2296(.dina(new_new_n8026__), .dinb(new_new_n8022__), .dout(new_new_n3238__));
  or1   g2297(.dina(new_new_n8028__), .dinb(new_new_n8024__), .dout(new_new_n3239__));
  and1  g2298(.dina(new_new_n8026__), .dinb(new_new_n8021__), .dout(new_new_n3240__));
  or1   g2299(.dina(new_new_n8028__), .dinb(new_new_n8023__), .dout(new_new_n3241__));
  and1  g2300(.dina(new_new_n3241__), .dinb(new_new_n3239__), .dout(new_new_n3242__));
  or1   g2301(.dina(new_new_n3240__), .dinb(new_new_n3238__), .dout(new_new_n3243__));
  and1  g2302(.dina(new_new_n8010__), .dinb(new_new_n8006__), .dout(new_new_n3244__));
  or1   g2303(.dina(new_new_n8012__), .dinb(new_new_n8008__), .dout(new_new_n3245__));
  and1  g2304(.dina(new_new_n8009__), .dinb(new_new_n8005__), .dout(new_new_n3246__));
  or1   g2305(.dina(new_new_n8011__), .dinb(new_new_n8007__), .dout(new_new_n3247__));
  and1  g2306(.dina(new_new_n3247__), .dinb(new_new_n3245__), .dout(new_new_n3248__));
  or1   g2307(.dina(new_new_n3246__), .dinb(new_new_n3244__), .dout(new_new_n3249__));
  and1  g2308(.dina(new_new_n7994__), .dinb(new_new_n7990__), .dout(new_new_n3250__));
  or1   g2309(.dina(new_new_n7996__), .dinb(new_new_n7992__), .dout(new_new_n3251__));
  and1  g2310(.dina(new_new_n7993__), .dinb(new_new_n7989__), .dout(new_new_n3252__));
  or1   g2311(.dina(new_new_n7995__), .dinb(new_new_n7991__), .dout(new_new_n3253__));
  and1  g2312(.dina(new_new_n3253__), .dinb(new_new_n3251__), .dout(new_new_n3254__));
  or1   g2313(.dina(new_new_n3252__), .dinb(new_new_n3250__), .dout(new_new_n3255__));
  and1  g2314(.dina(new_new_n8030__), .dinb(new_new_n1321__), .dout(new_new_n3256__));
  or1   g2315(.dina(new_new_n8032__), .dinb(new_new_n1322__), .dout(new_new_n3257__));
  and1  g2316(.dina(new_new_n8033__), .dinb(new_new_n8034__), .dout(new_new_n3258__));
  or1   g2317(.dina(new_new_n8035__), .dinb(new_new_n8036__), .dout(new_new_n3259__));
  and1  g2318(.dina(new_new_n8038__), .dinb(new_new_n8034__), .dout(new_new_n3260__));
  or1   g2319(.dina(new_new_n8040__), .dinb(new_new_n8036__), .dout(new_new_n3261__));
  and1  g2320(.dina(new_new_n8038__), .dinb(new_new_n8033__), .dout(new_new_n3262__));
  or1   g2321(.dina(new_new_n8040__), .dinb(new_new_n8035__), .dout(new_new_n3263__));
  and1  g2322(.dina(new_new_n3263__), .dinb(new_new_n3261__), .dout(new_new_n3264__));
  or1   g2323(.dina(new_new_n3262__), .dinb(new_new_n3260__), .dout(new_new_n3265__));
  and1  g2324(.dina(new_new_n6945__), .dinb(new_new_n8042__), .dout(new_new_n3266__));
  or1   g2325(.dina(new_new_n6958__), .dinb(new_new_n8045__), .dout(new_new_n3267__));
  and1  g2326(.dina(new_new_n8046__), .dinb(new_new_n8047__), .dout(new_new_n3268__));
  or1   g2327(.dina(new_new_n8048__), .dinb(new_new_n8049__), .dout(new_new_n3269__));
  and1  g2328(.dina(new_new_n8051__), .dinb(new_new_n8037__), .dout(new_new_n3270__));
  or1   g2329(.dina(new_new_n8053__), .dinb(new_new_n8039__), .dout(new_new_n3271__));
  and1  g2330(.dina(new_new_n8054__), .dinb(new_new_n8055__), .dout(new_new_n3272__));
  or1   g2331(.dina(new_new_n8056__), .dinb(new_new_n8057__), .dout(new_new_n3273__));
  and1  g2332(.dina(new_new_n8059__), .dinb(new_new_n8055__), .dout(new_new_n3274__));
  or1   g2333(.dina(new_new_n8061__), .dinb(new_new_n8057__), .dout(new_new_n3275__));
  and1  g2334(.dina(new_new_n8059__), .dinb(new_new_n8054__), .dout(new_new_n3276__));
  or1   g2335(.dina(new_new_n8061__), .dinb(new_new_n8056__), .dout(new_new_n3277__));
  and1  g2336(.dina(new_new_n3277__), .dinb(new_new_n3275__), .dout(new_new_n3278__));
  or1   g2337(.dina(new_new_n3276__), .dinb(new_new_n3274__), .dout(new_new_n3279__));
  and1  g2338(.dina(new_new_n8042__), .dinb(new_new_n7020__), .dout(new_new_n3280__));
  or1   g2339(.dina(new_new_n8045__), .dinb(new_new_n7035__), .dout(new_new_n3281__));
  and1  g2340(.dina(new_new_n8062__), .dinb(new_new_n8063__), .dout(new_new_n3282__));
  or1   g2341(.dina(new_new_n8064__), .dinb(new_new_n8065__), .dout(new_new_n3283__));
  and1  g2342(.dina(new_new_n8067__), .dinb(new_new_n8058__), .dout(new_new_n3284__));
  or1   g2343(.dina(new_new_n8069__), .dinb(new_new_n8060__), .dout(new_new_n3285__));
  and1  g2344(.dina(new_new_n8070__), .dinb(new_new_n8071__), .dout(new_new_n3286__));
  or1   g2345(.dina(new_new_n8072__), .dinb(new_new_n8073__), .dout(new_new_n3287__));
  and1  g2346(.dina(new_new_n8030__), .dinb(new_new_n1475__), .dout(new_new_n3288__));
  or1   g2347(.dina(new_new_n8032__), .dinb(new_new_n1476__), .dout(new_new_n3289__));
  and1  g2348(.dina(new_new_n8029__), .dinb(new_new_n1404__), .dout(new_new_n3290__));
  or1   g2349(.dina(new_new_n8031__), .dinb(new_new_n1403__), .dout(new_new_n3291__));
  and1  g2350(.dina(new_new_n3291__), .dinb(new_new_n3289__), .dout(new_new_n3292__));
  or1   g2351(.dina(new_new_n3290__), .dinb(new_new_n3288__), .dout(new_new_n3293__));
  and1  g2352(.dina(new_new_n1388__), .dinb(new_new_n1301__), .dout(new_new_n3294__));
  or1   g2353(.dina(new_new_n1387__), .dinb(new_new_n1302__), .dout(new_new_n3295__));
  and1  g2354(.dina(new_new_n8074__), .dinb(new_new_n8075__), .dout(new_new_n3296__));
  or1   g2355(.dina(new_new_n8076__), .dinb(new_new_n8077__), .dout(new_new_n3297__));
  and1  g2356(.dina(new_new_n8079__), .dinb(new_new_n8075__), .dout(new_new_n3298__));
  or1   g2357(.dina(new_new_n8081__), .dinb(new_new_n8077__), .dout(new_new_n3299__));
  and1  g2358(.dina(new_new_n8079__), .dinb(new_new_n8074__), .dout(new_new_n3300__));
  or1   g2359(.dina(new_new_n8081__), .dinb(new_new_n8076__), .dout(new_new_n3301__));
  and1  g2360(.dina(new_new_n3301__), .dinb(new_new_n3299__), .dout(new_new_n3302__));
  or1   g2361(.dina(new_new_n3300__), .dinb(new_new_n3298__), .dout(new_new_n3303__));
  and1  g2362(.dina(new_new_n6946__), .dinb(new_new_n8083__), .dout(new_new_n3304__));
  or1   g2363(.dina(new_new_n6959__), .dinb(new_new_n8086__), .dout(new_new_n3305__));
  and1  g2364(.dina(new_new_n8087__), .dinb(new_new_n8088__), .dout(new_new_n3306__));
  or1   g2365(.dina(new_new_n8089__), .dinb(new_new_n8090__), .dout(new_new_n3307__));
  and1  g2366(.dina(new_new_n8092__), .dinb(new_new_n8088__), .dout(new_new_n3308__));
  or1   g2367(.dina(new_new_n8094__), .dinb(new_new_n8090__), .dout(new_new_n3309__));
  and1  g2368(.dina(new_new_n8092__), .dinb(new_new_n8087__), .dout(new_new_n3310__));
  or1   g2369(.dina(new_new_n8094__), .dinb(new_new_n8089__), .dout(new_new_n3311__));
  and1  g2370(.dina(new_new_n3311__), .dinb(new_new_n3309__), .dout(new_new_n3312__));
  or1   g2371(.dina(new_new_n3310__), .dinb(new_new_n3308__), .dout(new_new_n3313__));
  and1  g2372(.dina(new_new_n8095__), .dinb(new_new_n8096__), .dout(new_new_n3314__));
  or1   g2373(.dina(new_new_n8097__), .dinb(new_new_n8098__), .dout(new_new_n3315__));
  and1  g2374(.dina(new_new_n8100__), .dinb(new_new_n8095__), .dout(new_new_n3316__));
  or1   g2375(.dina(new_new_n8102__), .dinb(new_new_n8097__), .dout(new_new_n3317__));
  and1  g2376(.dina(new_new_n8100__), .dinb(new_new_n8096__), .dout(new_new_n3318__));
  or1   g2377(.dina(new_new_n8102__), .dinb(new_new_n8098__), .dout(new_new_n3319__));
  and1  g2378(.dina(new_new_n3319__), .dinb(new_new_n3317__), .dout(new_new_n3320__));
  or1   g2379(.dina(new_new_n3318__), .dinb(new_new_n3316__), .dout(new_new_n3321__));
  and1  g2380(.dina(new_new_n6946__), .dinb(new_new_n8104__), .dout(new_new_n3322__));
  or1   g2381(.dina(new_new_n6959__), .dinb(new_new_n8107__), .dout(new_new_n3323__));
  and1  g2382(.dina(new_new_n8108__), .dinb(new_new_n8109__), .dout(new_new_n3324__));
  or1   g2383(.dina(new_new_n8110__), .dinb(new_new_n8111__), .dout(new_new_n3325__));
  and1  g2384(.dina(new_new_n8113__), .dinb(new_new_n8099__), .dout(new_new_n3326__));
  or1   g2385(.dina(new_new_n8115__), .dinb(new_new_n8101__), .dout(new_new_n3327__));
  and1  g2386(.dina(new_new_n8116__), .dinb(new_new_n8117__), .dout(new_new_n3328__));
  or1   g2387(.dina(new_new_n8118__), .dinb(new_new_n8119__), .dout(new_new_n3329__));
  and1  g2388(.dina(new_new_n8121__), .dinb(new_new_n8117__), .dout(new_new_n3330__));
  or1   g2389(.dina(new_new_n8123__), .dinb(new_new_n8119__), .dout(new_new_n3331__));
  and1  g2390(.dina(new_new_n8121__), .dinb(new_new_n8116__), .dout(new_new_n3332__));
  or1   g2391(.dina(new_new_n8123__), .dinb(new_new_n8118__), .dout(new_new_n3333__));
  and1  g2392(.dina(new_new_n3333__), .dinb(new_new_n3331__), .dout(new_new_n3334__));
  or1   g2393(.dina(new_new_n3332__), .dinb(new_new_n3330__), .dout(new_new_n3335__));
  and1  g2394(.dina(new_new_n8104__), .dinb(new_new_n7022__), .dout(new_new_n3336__));
  or1   g2395(.dina(new_new_n8107__), .dinb(new_new_n7037__), .dout(new_new_n3337__));
  and1  g2396(.dina(new_new_n8124__), .dinb(new_new_n8125__), .dout(new_new_n3338__));
  or1   g2397(.dina(new_new_n8126__), .dinb(new_new_n8127__), .dout(new_new_n3339__));
  and1  g2398(.dina(new_new_n8129__), .dinb(new_new_n8125__), .dout(new_new_n3340__));
  or1   g2399(.dina(new_new_n8131__), .dinb(new_new_n8127__), .dout(new_new_n3341__));
  and1  g2400(.dina(new_new_n8129__), .dinb(new_new_n8124__), .dout(new_new_n3342__));
  or1   g2401(.dina(new_new_n8131__), .dinb(new_new_n8126__), .dout(new_new_n3343__));
  and1  g2402(.dina(new_new_n3343__), .dinb(new_new_n3341__), .dout(new_new_n3344__));
  or1   g2403(.dina(new_new_n3342__), .dinb(new_new_n3340__), .dout(new_new_n3345__));
  and1  g2404(.dina(new_new_n8113__), .dinb(new_new_n8109__), .dout(new_new_n3346__));
  or1   g2405(.dina(new_new_n8115__), .dinb(new_new_n8111__), .dout(new_new_n3347__));
  and1  g2406(.dina(new_new_n8112__), .dinb(new_new_n8108__), .dout(new_new_n3348__));
  or1   g2407(.dina(new_new_n8114__), .dinb(new_new_n8110__), .dout(new_new_n3349__));
  and1  g2408(.dina(new_new_n3349__), .dinb(new_new_n3347__), .dout(new_new_n3350__));
  or1   g2409(.dina(new_new_n3348__), .dinb(new_new_n3346__), .dout(new_new_n3351__));
  and1  g2410(.dina(new_new_n1518__), .dinb(new_new_n1510__), .dout(new_new_n3352__));
  or1   g2411(.dina(new_new_n1517__), .dinb(new_new_n1509__), .dout(new_new_n3353__));
  and1  g2412(.dina(new_new_n6949__), .dinb(new_new_n8133__), .dout(new_new_n3354__));
  or1   g2413(.dina(new_new_n6962__), .dinb(new_new_n8136__), .dout(new_new_n3355__));
  and1  g2414(.dina(new_new_n8138__), .dinb(new_new_n8139__), .dout(new_new_n3356__));
  or1   g2415(.dina(new_new_n8140__), .dinb(new_new_n8141__), .dout(new_new_n3357__));
  and1  g2416(.dina(new_new_n8143__), .dinb(new_new_n1453__), .dout(new_new_n3358__));
  or1   g2417(.dina(new_new_n8145__), .dinb(new_new_n1454__), .dout(new_new_n3359__));
  and1  g2418(.dina(new_new_n8146__), .dinb(new_new_n8147__), .dout(new_new_n3360__));
  or1   g2419(.dina(new_new_n8148__), .dinb(new_new_n8149__), .dout(new_new_n3361__));
  and1  g2420(.dina(new_new_n8151__), .dinb(new_new_n8147__), .dout(new_new_n3362__));
  or1   g2421(.dina(new_new_n8153__), .dinb(new_new_n8149__), .dout(new_new_n3363__));
  and1  g2422(.dina(new_new_n8151__), .dinb(new_new_n8146__), .dout(new_new_n3364__));
  or1   g2423(.dina(new_new_n8153__), .dinb(new_new_n8148__), .dout(new_new_n3365__));
  and1  g2424(.dina(new_new_n3365__), .dinb(new_new_n3363__), .dout(new_new_n3366__));
  or1   g2425(.dina(new_new_n3364__), .dinb(new_new_n3362__), .dout(new_new_n3367__));
  and1  g2426(.dina(new_new_n8133__), .dinb(new_new_n7022__), .dout(new_new_n3368__));
  or1   g2427(.dina(new_new_n8136__), .dinb(new_new_n7037__), .dout(new_new_n3369__));
  and1  g2428(.dina(new_new_n8154__), .dinb(new_new_n8155__), .dout(new_new_n3370__));
  or1   g2429(.dina(new_new_n8156__), .dinb(new_new_n8157__), .dout(new_new_n3371__));
  and1  g2430(.dina(new_new_n8159__), .dinb(new_new_n8150__), .dout(new_new_n3372__));
  or1   g2431(.dina(new_new_n8161__), .dinb(new_new_n8152__), .dout(new_new_n3373__));
  and1  g2432(.dina(new_new_n8162__), .dinb(new_new_n8163__), .dout(new_new_n3374__));
  or1   g2433(.dina(new_new_n8164__), .dinb(new_new_n8165__), .dout(new_new_n3375__));
  and1  g2434(.dina(new_new_n8167__), .dinb(new_new_n8163__), .dout(new_new_n3376__));
  or1   g2435(.dina(new_new_n8169__), .dinb(new_new_n8165__), .dout(new_new_n3377__));
  and1  g2436(.dina(new_new_n8167__), .dinb(new_new_n8162__), .dout(new_new_n3378__));
  or1   g2437(.dina(new_new_n8169__), .dinb(new_new_n8164__), .dout(new_new_n3379__));
  and1  g2438(.dina(new_new_n3379__), .dinb(new_new_n3377__), .dout(new_new_n3380__));
  or1   g2439(.dina(new_new_n3378__), .dinb(new_new_n3376__), .dout(new_new_n3381__));
  and1  g2440(.dina(new_new_n8134__), .dinb(new_new_n7594__), .dout(new_new_n3382__));
  or1   g2441(.dina(new_new_n8137__), .dinb(new_new_n7607__), .dout(new_new_n3383__));
  and1  g2442(.dina(new_new_n8170__), .dinb(new_new_n8171__), .dout(new_new_n3384__));
  or1   g2443(.dina(new_new_n8172__), .dinb(new_new_n8173__), .dout(new_new_n3385__));
  and1  g2444(.dina(new_new_n8175__), .dinb(new_new_n8171__), .dout(new_new_n3386__));
  or1   g2445(.dina(new_new_n8177__), .dinb(new_new_n8173__), .dout(new_new_n3387__));
  and1  g2446(.dina(new_new_n8175__), .dinb(new_new_n8170__), .dout(new_new_n3388__));
  or1   g2447(.dina(new_new_n8177__), .dinb(new_new_n8172__), .dout(new_new_n3389__));
  and1  g2448(.dina(new_new_n3389__), .dinb(new_new_n3387__), .dout(new_new_n3390__));
  or1   g2449(.dina(new_new_n3388__), .dinb(new_new_n3386__), .dout(new_new_n3391__));
  and1  g2450(.dina(new_new_n8159__), .dinb(new_new_n8155__), .dout(new_new_n3392__));
  or1   g2451(.dina(new_new_n8161__), .dinb(new_new_n8157__), .dout(new_new_n3393__));
  and1  g2452(.dina(new_new_n8158__), .dinb(new_new_n8154__), .dout(new_new_n3394__));
  or1   g2453(.dina(new_new_n8160__), .dinb(new_new_n8156__), .dout(new_new_n3395__));
  and1  g2454(.dina(new_new_n3395__), .dinb(new_new_n3393__), .dout(new_new_n3396__));
  or1   g2455(.dina(new_new_n3394__), .dinb(new_new_n3392__), .dout(new_new_n3397__));
  and1  g2456(.dina(new_new_n8143__), .dinb(new_new_n8139__), .dout(new_new_n3398__));
  or1   g2457(.dina(new_new_n8145__), .dinb(new_new_n8141__), .dout(new_new_n3399__));
  and1  g2458(.dina(new_new_n8142__), .dinb(new_new_n8138__), .dout(new_new_n3400__));
  or1   g2459(.dina(new_new_n8144__), .dinb(new_new_n8140__), .dout(new_new_n3401__));
  and1  g2460(.dina(new_new_n3401__), .dinb(new_new_n3399__), .dout(new_new_n3402__));
  or1   g2461(.dina(new_new_n3400__), .dinb(new_new_n3398__), .dout(new_new_n3403__));
  and1  g2462(.dina(new_new_n8179__), .dinb(new_new_n1325__), .dout(new_new_n3404__));
  or1   g2463(.dina(new_new_n8181__), .dinb(new_new_n1326__), .dout(new_new_n3405__));
  and1  g2464(.dina(new_new_n8182__), .dinb(new_new_n8183__), .dout(new_new_n3406__));
  or1   g2465(.dina(new_new_n8184__), .dinb(new_new_n8185__), .dout(new_new_n3407__));
  and1  g2466(.dina(new_new_n8187__), .dinb(new_new_n8183__), .dout(new_new_n3408__));
  or1   g2467(.dina(new_new_n8189__), .dinb(new_new_n8185__), .dout(new_new_n3409__));
  and1  g2468(.dina(new_new_n8187__), .dinb(new_new_n8182__), .dout(new_new_n3410__));
  or1   g2469(.dina(new_new_n8189__), .dinb(new_new_n8184__), .dout(new_new_n3411__));
  and1  g2470(.dina(new_new_n3411__), .dinb(new_new_n3409__), .dout(new_new_n3412__));
  or1   g2471(.dina(new_new_n3410__), .dinb(new_new_n3408__), .dout(new_new_n3413__));
  and1  g2472(.dina(new_new_n8191__), .dinb(new_new_n7023__), .dout(new_new_n3414__));
  or1   g2473(.dina(new_new_n8194__), .dinb(new_new_n7038__), .dout(new_new_n3415__));
  and1  g2474(.dina(new_new_n8195__), .dinb(new_new_n8196__), .dout(new_new_n3416__));
  or1   g2475(.dina(new_new_n8197__), .dinb(new_new_n8198__), .dout(new_new_n3417__));
  and1  g2476(.dina(new_new_n8200__), .dinb(new_new_n8186__), .dout(new_new_n3418__));
  or1   g2477(.dina(new_new_n8202__), .dinb(new_new_n8188__), .dout(new_new_n3419__));
  and1  g2478(.dina(new_new_n8203__), .dinb(new_new_n8204__), .dout(new_new_n3420__));
  or1   g2479(.dina(new_new_n8205__), .dinb(new_new_n8206__), .dout(new_new_n3421__));
  and1  g2480(.dina(new_new_n8208__), .dinb(new_new_n8204__), .dout(new_new_n3422__));
  or1   g2481(.dina(new_new_n8210__), .dinb(new_new_n8206__), .dout(new_new_n3423__));
  and1  g2482(.dina(new_new_n8208__), .dinb(new_new_n8203__), .dout(new_new_n3424__));
  or1   g2483(.dina(new_new_n8210__), .dinb(new_new_n8205__), .dout(new_new_n3425__));
  and1  g2484(.dina(new_new_n3425__), .dinb(new_new_n3423__), .dout(new_new_n3426__));
  or1   g2485(.dina(new_new_n3424__), .dinb(new_new_n3422__), .dout(new_new_n3427__));
  and1  g2486(.dina(new_new_n8191__), .dinb(new_new_n7595__), .dout(new_new_n3428__));
  or1   g2487(.dina(new_new_n8194__), .dinb(new_new_n7608__), .dout(new_new_n3429__));
  and1  g2488(.dina(new_new_n8211__), .dinb(new_new_n8212__), .dout(new_new_n3430__));
  or1   g2489(.dina(new_new_n8213__), .dinb(new_new_n8214__), .dout(new_new_n3431__));
  and1  g2490(.dina(new_new_n8216__), .dinb(new_new_n8207__), .dout(new_new_n3432__));
  or1   g2491(.dina(new_new_n8218__), .dinb(new_new_n8209__), .dout(new_new_n3433__));
  and1  g2492(.dina(new_new_n8219__), .dinb(new_new_n8220__), .dout(new_new_n3434__));
  or1   g2493(.dina(new_new_n8221__), .dinb(new_new_n8222__), .dout(new_new_n3435__));
  and1  g2494(.dina(new_new_n8179__), .dinb(new_new_n1479__), .dout(new_new_n3436__));
  or1   g2495(.dina(new_new_n8181__), .dinb(new_new_n1480__), .dout(new_new_n3437__));
  and1  g2496(.dina(new_new_n8178__), .dinb(new_new_n1406__), .dout(new_new_n3438__));
  or1   g2497(.dina(new_new_n8180__), .dinb(new_new_n1405__), .dout(new_new_n3439__));
  and1  g2498(.dina(new_new_n3439__), .dinb(new_new_n3437__), .dout(new_new_n3440__));
  or1   g2499(.dina(new_new_n3438__), .dinb(new_new_n3436__), .dout(new_new_n3441__));
  and1  g2500(.dina(new_new_n8223__), .dinb(new_new_n8224__), .dout(new_new_n3442__));
  or1   g2501(.dina(new_new_n8225__), .dinb(new_new_n8226__), .dout(new_new_n3443__));
  and1  g2502(.dina(new_new_n8228__), .dinb(new_new_n1393__), .dout(new_new_n3444__));
  or1   g2503(.dina(new_new_n8230__), .dinb(new_new_n1394__), .dout(new_new_n3445__));
  and1  g2504(.dina(new_new_n8231__), .dinb(new_new_n8232__), .dout(new_new_n3446__));
  or1   g2505(.dina(new_new_n8233__), .dinb(new_new_n8234__), .dout(new_new_n3447__));
  and1  g2506(.dina(new_new_n8236__), .dinb(new_new_n8232__), .dout(new_new_n3448__));
  or1   g2507(.dina(new_new_n8238__), .dinb(new_new_n8234__), .dout(new_new_n3449__));
  and1  g2508(.dina(new_new_n8236__), .dinb(new_new_n8231__), .dout(new_new_n3450__));
  or1   g2509(.dina(new_new_n8238__), .dinb(new_new_n8233__), .dout(new_new_n3451__));
  and1  g2510(.dina(new_new_n3451__), .dinb(new_new_n3449__), .dout(new_new_n3452__));
  or1   g2511(.dina(new_new_n3450__), .dinb(new_new_n3448__), .dout(new_new_n3453__));
  and1  g2512(.dina(new_new_n8240__), .dinb(new_new_n7023__), .dout(new_new_n3454__));
  or1   g2513(.dina(new_new_n8243__), .dinb(new_new_n7038__), .dout(new_new_n3455__));
  and1  g2514(.dina(new_new_n8244__), .dinb(new_new_n8245__), .dout(new_new_n3456__));
  or1   g2515(.dina(new_new_n8246__), .dinb(new_new_n8247__), .dout(new_new_n3457__));
  and1  g2516(.dina(new_new_n8249__), .dinb(new_new_n8245__), .dout(new_new_n3458__));
  or1   g2517(.dina(new_new_n8251__), .dinb(new_new_n8247__), .dout(new_new_n3459__));
  and1  g2518(.dina(new_new_n8249__), .dinb(new_new_n8244__), .dout(new_new_n3460__));
  or1   g2519(.dina(new_new_n8251__), .dinb(new_new_n8246__), .dout(new_new_n3461__));
  and1  g2520(.dina(new_new_n3461__), .dinb(new_new_n3459__), .dout(new_new_n3462__));
  or1   g2521(.dina(new_new_n3460__), .dinb(new_new_n3458__), .dout(new_new_n3463__));
  and1  g2522(.dina(new_new_n8228__), .dinb(new_new_n8223__), .dout(new_new_n3464__));
  or1   g2523(.dina(new_new_n8230__), .dinb(new_new_n8225__), .dout(new_new_n3465__));
  and1  g2524(.dina(new_new_n8227__), .dinb(new_new_n8224__), .dout(new_new_n3466__));
  or1   g2525(.dina(new_new_n8229__), .dinb(new_new_n8226__), .dout(new_new_n3467__));
  and1  g2526(.dina(new_new_n3467__), .dinb(new_new_n3465__), .dout(new_new_n3468__));
  or1   g2527(.dina(new_new_n3466__), .dinb(new_new_n3464__), .dout(new_new_n3469__));
  and1  g2528(.dina(new_new_n1520__), .dinb(new_new_n1514__), .dout(new_new_n3470__));
  or1   g2529(.dina(new_new_n1519__), .dinb(new_new_n1513__), .dout(new_new_n3471__));
  and1  g2530(.dina(new_new_n6949__), .dinb(new_new_n8254__), .dout(new_new_n3472__));
  or1   g2531(.dina(new_new_n6962__), .dinb(new_new_n8257__), .dout(new_new_n3473__));
  and1  g2532(.dina(new_new_n8259__), .dinb(new_new_n8260__), .dout(new_new_n3474__));
  or1   g2533(.dina(new_new_n8261__), .dinb(new_new_n8262__), .dout(new_new_n3475__));
  and1  g2534(.dina(new_new_n8264__), .dinb(new_new_n1457__), .dout(new_new_n3476__));
  or1   g2535(.dina(new_new_n8266__), .dinb(new_new_n1458__), .dout(new_new_n3477__));
  and1  g2536(.dina(new_new_n8267__), .dinb(new_new_n8268__), .dout(new_new_n3478__));
  or1   g2537(.dina(new_new_n8269__), .dinb(new_new_n8270__), .dout(new_new_n3479__));
  and1  g2538(.dina(new_new_n8272__), .dinb(new_new_n8268__), .dout(new_new_n3480__));
  or1   g2539(.dina(new_new_n8274__), .dinb(new_new_n8270__), .dout(new_new_n3481__));
  and1  g2540(.dina(new_new_n8272__), .dinb(new_new_n8267__), .dout(new_new_n3482__));
  or1   g2541(.dina(new_new_n8274__), .dinb(new_new_n8269__), .dout(new_new_n3483__));
  and1  g2542(.dina(new_new_n3483__), .dinb(new_new_n3481__), .dout(new_new_n3484__));
  or1   g2543(.dina(new_new_n3482__), .dinb(new_new_n3480__), .dout(new_new_n3485__));
  and1  g2544(.dina(new_new_n8254__), .dinb(new_new_n7026__), .dout(new_new_n3486__));
  or1   g2545(.dina(new_new_n8257__), .dinb(new_new_n7041__), .dout(new_new_n3487__));
  and1  g2546(.dina(new_new_n8275__), .dinb(new_new_n8276__), .dout(new_new_n3488__));
  or1   g2547(.dina(new_new_n8277__), .dinb(new_new_n8278__), .dout(new_new_n3489__));
  and1  g2548(.dina(new_new_n8280__), .dinb(new_new_n8271__), .dout(new_new_n3490__));
  or1   g2549(.dina(new_new_n8282__), .dinb(new_new_n8273__), .dout(new_new_n3491__));
  and1  g2550(.dina(new_new_n8283__), .dinb(new_new_n8284__), .dout(new_new_n3492__));
  or1   g2551(.dina(new_new_n8285__), .dinb(new_new_n8286__), .dout(new_new_n3493__));
  and1  g2552(.dina(new_new_n8288__), .dinb(new_new_n8284__), .dout(new_new_n3494__));
  or1   g2553(.dina(new_new_n8290__), .dinb(new_new_n8286__), .dout(new_new_n3495__));
  and1  g2554(.dina(new_new_n8288__), .dinb(new_new_n8283__), .dout(new_new_n3496__));
  or1   g2555(.dina(new_new_n8290__), .dinb(new_new_n8285__), .dout(new_new_n3497__));
  and1  g2556(.dina(new_new_n3497__), .dinb(new_new_n3495__), .dout(new_new_n3498__));
  or1   g2557(.dina(new_new_n3496__), .dinb(new_new_n3494__), .dout(new_new_n3499__));
  and1  g2558(.dina(new_new_n8253__), .dinb(new_new_n7595__), .dout(new_new_n3500__));
  or1   g2559(.dina(new_new_n8258__), .dinb(new_new_n7608__), .dout(new_new_n3501__));
  and1  g2560(.dina(new_new_n8291__), .dinb(new_new_n8292__), .dout(new_new_n3502__));
  or1   g2561(.dina(new_new_n8293__), .dinb(new_new_n8294__), .dout(new_new_n3503__));
  and1  g2562(.dina(new_new_n8296__), .dinb(new_new_n8292__), .dout(new_new_n3504__));
  or1   g2563(.dina(new_new_n8298__), .dinb(new_new_n8294__), .dout(new_new_n3505__));
  and1  g2564(.dina(new_new_n8296__), .dinb(new_new_n8291__), .dout(new_new_n3506__));
  or1   g2565(.dina(new_new_n8298__), .dinb(new_new_n8293__), .dout(new_new_n3507__));
  and1  g2566(.dina(new_new_n3507__), .dinb(new_new_n3505__), .dout(new_new_n3508__));
  or1   g2567(.dina(new_new_n3506__), .dinb(new_new_n3504__), .dout(new_new_n3509__));
  and1  g2568(.dina(new_new_n8280__), .dinb(new_new_n8276__), .dout(new_new_n3510__));
  or1   g2569(.dina(new_new_n8282__), .dinb(new_new_n8278__), .dout(new_new_n3511__));
  and1  g2570(.dina(new_new_n8279__), .dinb(new_new_n8275__), .dout(new_new_n3512__));
  or1   g2571(.dina(new_new_n8281__), .dinb(new_new_n8277__), .dout(new_new_n3513__));
  and1  g2572(.dina(new_new_n3513__), .dinb(new_new_n3511__), .dout(new_new_n3514__));
  or1   g2573(.dina(new_new_n3512__), .dinb(new_new_n3510__), .dout(new_new_n3515__));
  and1  g2574(.dina(new_new_n8264__), .dinb(new_new_n8260__), .dout(new_new_n3516__));
  or1   g2575(.dina(new_new_n8266__), .dinb(new_new_n8262__), .dout(new_new_n3517__));
  and1  g2576(.dina(new_new_n8263__), .dinb(new_new_n8259__), .dout(new_new_n3518__));
  or1   g2577(.dina(new_new_n8265__), .dinb(new_new_n8261__), .dout(new_new_n3519__));
  and1  g2578(.dina(new_new_n3519__), .dinb(new_new_n3517__), .dout(new_new_n3520__));
  or1   g2579(.dina(new_new_n3518__), .dinb(new_new_n3516__), .dout(new_new_n3521__));
  and1  g2580(.dina(new_new_n8300__), .dinb(new_new_n1472__), .dout(new_new_n3522__));
  or1   g2581(.dina(new_new_n8302__), .dinb(new_new_n1471__), .dout(new_new_n3523__));
  and1  g2582(.dina(new_new_n8300__), .dinb(new_new_n1420__), .dout(new_new_n3524__));
  or1   g2583(.dina(new_new_n8302__), .dinb(new_new_n1419__), .dout(new_new_n3525__));
  and1  g2584(.dina(new_new_n3525__), .dinb(new_new_n3523__), .dout(new_new_n3526__));
  or1   g2585(.dina(new_new_n3524__), .dinb(new_new_n3522__), .dout(new_new_n3527__));
  and1  g2586(.dina(new_new_n6950__), .dinb(new_new_n8305__), .dout(new_new_n3528__));
  or1   g2587(.dina(new_new_n6963__), .dinb(new_new_n8309__), .dout(new_new_n3529__));
  and1  g2588(.dina(new_new_n8311__), .dinb(new_new_n8312__), .dout(new_new_n3530__));
  or1   g2589(.dina(new_new_n8313__), .dinb(new_new_n8314__), .dout(new_new_n3531__));
  and1  g2590(.dina(new_new_n8316__), .dinb(new_new_n8299__), .dout(new_new_n3532__));
  or1   g2591(.dina(new_new_n8318__), .dinb(new_new_n8301__), .dout(new_new_n3533__));
  and1  g2592(.dina(new_new_n8319__), .dinb(new_new_n8320__), .dout(new_new_n3534__));
  or1   g2593(.dina(new_new_n8321__), .dinb(new_new_n8322__), .dout(new_new_n3535__));
  and1  g2594(.dina(new_new_n8324__), .dinb(new_new_n8320__), .dout(new_new_n3536__));
  or1   g2595(.dina(new_new_n8326__), .dinb(new_new_n8322__), .dout(new_new_n3537__));
  and1  g2596(.dina(new_new_n8324__), .dinb(new_new_n8319__), .dout(new_new_n3538__));
  or1   g2597(.dina(new_new_n8326__), .dinb(new_new_n8321__), .dout(new_new_n3539__));
  and1  g2598(.dina(new_new_n3539__), .dinb(new_new_n3537__), .dout(new_new_n3540__));
  or1   g2599(.dina(new_new_n3538__), .dinb(new_new_n3536__), .dout(new_new_n3541__));
  and1  g2600(.dina(new_new_n8305__), .dinb(new_new_n7026__), .dout(new_new_n3542__));
  or1   g2601(.dina(new_new_n8309__), .dinb(new_new_n7041__), .dout(new_new_n3543__));
  and1  g2602(.dina(new_new_n8327__), .dinb(new_new_n8328__), .dout(new_new_n3544__));
  or1   g2603(.dina(new_new_n8329__), .dinb(new_new_n8330__), .dout(new_new_n3545__));
  and1  g2604(.dina(new_new_n8332__), .dinb(new_new_n8323__), .dout(new_new_n3546__));
  or1   g2605(.dina(new_new_n8334__), .dinb(new_new_n8325__), .dout(new_new_n3547__));
  and1  g2606(.dina(new_new_n8335__), .dinb(new_new_n8336__), .dout(new_new_n3548__));
  or1   g2607(.dina(new_new_n8337__), .dinb(new_new_n8338__), .dout(new_new_n3549__));
  and1  g2608(.dina(new_new_n8340__), .dinb(new_new_n8336__), .dout(new_new_n3550__));
  or1   g2609(.dina(new_new_n8342__), .dinb(new_new_n8338__), .dout(new_new_n3551__));
  and1  g2610(.dina(new_new_n8340__), .dinb(new_new_n8335__), .dout(new_new_n3552__));
  or1   g2611(.dina(new_new_n8342__), .dinb(new_new_n8337__), .dout(new_new_n3553__));
  and1  g2612(.dina(new_new_n3553__), .dinb(new_new_n3551__), .dout(new_new_n3554__));
  or1   g2613(.dina(new_new_n3552__), .dinb(new_new_n3550__), .dout(new_new_n3555__));
  and1  g2614(.dina(new_new_n8304__), .dinb(new_new_n7597__), .dout(new_new_n3556__));
  or1   g2615(.dina(new_new_n8308__), .dinb(new_new_n7610__), .dout(new_new_n3557__));
  and1  g2616(.dina(new_new_n8343__), .dinb(new_new_n8344__), .dout(new_new_n3558__));
  or1   g2617(.dina(new_new_n8345__), .dinb(new_new_n8346__), .dout(new_new_n3559__));
  and1  g2618(.dina(new_new_n8348__), .dinb(new_new_n8339__), .dout(new_new_n3560__));
  or1   g2619(.dina(new_new_n8350__), .dinb(new_new_n8341__), .dout(new_new_n3561__));
  and1  g2620(.dina(new_new_n8351__), .dinb(new_new_n8352__), .dout(new_new_n3562__));
  or1   g2621(.dina(new_new_n8353__), .dinb(new_new_n8354__), .dout(new_new_n3563__));
  and1  g2622(.dina(new_new_n8356__), .dinb(new_new_n8352__), .dout(new_new_n3564__));
  or1   g2623(.dina(new_new_n8358__), .dinb(new_new_n8354__), .dout(new_new_n3565__));
  and1  g2624(.dina(new_new_n8356__), .dinb(new_new_n8351__), .dout(new_new_n3566__));
  or1   g2625(.dina(new_new_n8358__), .dinb(new_new_n8353__), .dout(new_new_n3567__));
  and1  g2626(.dina(new_new_n3567__), .dinb(new_new_n3565__), .dout(new_new_n3568__));
  or1   g2627(.dina(new_new_n3566__), .dinb(new_new_n3564__), .dout(new_new_n3569__));
  and1  g2628(.dina(new_new_n8306__), .dinb(new_new_n8362__), .dout(new_new_n3570__));
  or1   g2629(.dina(new_new_n8310__), .dinb(new_new_n8371__), .dout(new_new_n3571__));
  and1  g2630(.dina(new_new_n8377__), .dinb(new_new_n8378__), .dout(new_new_n3572__));
  or1   g2631(.dina(new_new_n8379__), .dinb(new_new_n8380__), .dout(new_new_n3573__));
  and1  g2632(.dina(new_new_n8382__), .dinb(new_new_n8378__), .dout(new_new_n3574__));
  or1   g2633(.dina(new_new_n8384__), .dinb(new_new_n8380__), .dout(new_new_n3575__));
  and1  g2634(.dina(new_new_n8382__), .dinb(new_new_n8377__), .dout(new_new_n3576__));
  or1   g2635(.dina(new_new_n8384__), .dinb(new_new_n8379__), .dout(new_new_n3577__));
  and1  g2636(.dina(new_new_n3577__), .dinb(new_new_n3575__), .dout(new_new_n3578__));
  or1   g2637(.dina(new_new_n3576__), .dinb(new_new_n3574__), .dout(new_new_n3579__));
  and1  g2638(.dina(new_new_n8348__), .dinb(new_new_n8344__), .dout(new_new_n3580__));
  or1   g2639(.dina(new_new_n8350__), .dinb(new_new_n8346__), .dout(new_new_n3581__));
  and1  g2640(.dina(new_new_n8347__), .dinb(new_new_n8343__), .dout(new_new_n3582__));
  or1   g2641(.dina(new_new_n8349__), .dinb(new_new_n8345__), .dout(new_new_n3583__));
  and1  g2642(.dina(new_new_n3583__), .dinb(new_new_n3581__), .dout(new_new_n3584__));
  or1   g2643(.dina(new_new_n3582__), .dinb(new_new_n3580__), .dout(new_new_n3585__));
  and1  g2644(.dina(new_new_n8332__), .dinb(new_new_n8328__), .dout(new_new_n3586__));
  or1   g2645(.dina(new_new_n8334__), .dinb(new_new_n8330__), .dout(new_new_n3587__));
  and1  g2646(.dina(new_new_n8331__), .dinb(new_new_n8327__), .dout(new_new_n3588__));
  or1   g2647(.dina(new_new_n8333__), .dinb(new_new_n8329__), .dout(new_new_n3589__));
  and1  g2648(.dina(new_new_n3589__), .dinb(new_new_n3587__), .dout(new_new_n3590__));
  or1   g2649(.dina(new_new_n3588__), .dinb(new_new_n3586__), .dout(new_new_n3591__));
  and1  g2650(.dina(new_new_n8316__), .dinb(new_new_n8312__), .dout(new_new_n3592__));
  or1   g2651(.dina(new_new_n8318__), .dinb(new_new_n8314__), .dout(new_new_n3593__));
  and1  g2652(.dina(new_new_n8315__), .dinb(new_new_n8311__), .dout(new_new_n3594__));
  or1   g2653(.dina(new_new_n8317__), .dinb(new_new_n8313__), .dout(new_new_n3595__));
  and1  g2654(.dina(new_new_n3595__), .dinb(new_new_n3593__), .dout(new_new_n3596__));
  or1   g2655(.dina(new_new_n3594__), .dinb(new_new_n3592__), .dout(new_new_n3597__));
  and1  g2656(.dina(new_new_n8385__), .dinb(new_new_n8386__), .dout(new_new_n3598__));
  or1   g2657(.dina(new_new_n8387__), .dinb(new_new_n8388__), .dout(new_new_n3599__));
  and1  g2658(.dina(new_new_n8390__), .dinb(new_new_n8385__), .dout(new_new_n3600__));
  or1   g2659(.dina(new_new_n8392__), .dinb(new_new_n8387__), .dout(new_new_n3601__));
  and1  g2660(.dina(new_new_n8390__), .dinb(new_new_n8386__), .dout(new_new_n3602__));
  or1   g2661(.dina(new_new_n8392__), .dinb(new_new_n8388__), .dout(new_new_n3603__));
  and1  g2662(.dina(new_new_n3603__), .dinb(new_new_n3601__), .dout(new_new_n3604__));
  or1   g2663(.dina(new_new_n3602__), .dinb(new_new_n3600__), .dout(new_new_n3605__));
  and1  g2664(.dina(new_new_n6950__), .dinb(new_new_n8395__), .dout(new_new_n3606__));
  or1   g2665(.dina(new_new_n6963__), .dinb(new_new_n8400__), .dout(new_new_n3607__));
  and1  g2666(.dina(new_new_n8402__), .dinb(new_new_n8403__), .dout(new_new_n3608__));
  or1   g2667(.dina(new_new_n8404__), .dinb(new_new_n8405__), .dout(new_new_n3609__));
  and1  g2668(.dina(new_new_n8407__), .dinb(new_new_n8389__), .dout(new_new_n3610__));
  or1   g2669(.dina(new_new_n8409__), .dinb(new_new_n8391__), .dout(new_new_n3611__));
  and1  g2670(.dina(new_new_n8410__), .dinb(new_new_n8411__), .dout(new_new_n3612__));
  or1   g2671(.dina(new_new_n8412__), .dinb(new_new_n8413__), .dout(new_new_n3613__));
  and1  g2672(.dina(new_new_n8415__), .dinb(new_new_n8411__), .dout(new_new_n3614__));
  or1   g2673(.dina(new_new_n8417__), .dinb(new_new_n8413__), .dout(new_new_n3615__));
  and1  g2674(.dina(new_new_n8415__), .dinb(new_new_n8410__), .dout(new_new_n3616__));
  or1   g2675(.dina(new_new_n8417__), .dinb(new_new_n8412__), .dout(new_new_n3617__));
  and1  g2676(.dina(new_new_n3617__), .dinb(new_new_n3615__), .dout(new_new_n3618__));
  or1   g2677(.dina(new_new_n3616__), .dinb(new_new_n3614__), .dout(new_new_n3619__));
  and1  g2678(.dina(new_new_n8395__), .dinb(new_new_n7027__), .dout(new_new_n3620__));
  or1   g2679(.dina(new_new_n8400__), .dinb(new_new_n7042__), .dout(new_new_n3621__));
  and1  g2680(.dina(new_new_n8418__), .dinb(new_new_n8419__), .dout(new_new_n3622__));
  or1   g2681(.dina(new_new_n8420__), .dinb(new_new_n8421__), .dout(new_new_n3623__));
  and1  g2682(.dina(new_new_n8423__), .dinb(new_new_n8414__), .dout(new_new_n3624__));
  or1   g2683(.dina(new_new_n8425__), .dinb(new_new_n8416__), .dout(new_new_n3625__));
  and1  g2684(.dina(new_new_n8426__), .dinb(new_new_n8427__), .dout(new_new_n3626__));
  or1   g2685(.dina(new_new_n8428__), .dinb(new_new_n8429__), .dout(new_new_n3627__));
  and1  g2686(.dina(new_new_n8431__), .dinb(new_new_n8427__), .dout(new_new_n3628__));
  or1   g2687(.dina(new_new_n8433__), .dinb(new_new_n8429__), .dout(new_new_n3629__));
  and1  g2688(.dina(new_new_n8431__), .dinb(new_new_n8426__), .dout(new_new_n3630__));
  or1   g2689(.dina(new_new_n8433__), .dinb(new_new_n8428__), .dout(new_new_n3631__));
  and1  g2690(.dina(new_new_n3631__), .dinb(new_new_n3629__), .dout(new_new_n3632__));
  or1   g2691(.dina(new_new_n3630__), .dinb(new_new_n3628__), .dout(new_new_n3633__));
  and1  g2692(.dina(new_new_n8396__), .dinb(new_new_n7597__), .dout(new_new_n3634__));
  or1   g2693(.dina(new_new_n8399__), .dinb(new_new_n7610__), .dout(new_new_n3635__));
  and1  g2694(.dina(new_new_n8434__), .dinb(new_new_n8435__), .dout(new_new_n3636__));
  or1   g2695(.dina(new_new_n8436__), .dinb(new_new_n8437__), .dout(new_new_n3637__));
  and1  g2696(.dina(new_new_n8439__), .dinb(new_new_n8430__), .dout(new_new_n3638__));
  or1   g2697(.dina(new_new_n8441__), .dinb(new_new_n8432__), .dout(new_new_n3639__));
  and1  g2698(.dina(new_new_n8442__), .dinb(new_new_n8443__), .dout(new_new_n3640__));
  or1   g2699(.dina(new_new_n8444__), .dinb(new_new_n8445__), .dout(new_new_n3641__));
  and1  g2700(.dina(new_new_n8447__), .dinb(new_new_n8443__), .dout(new_new_n3642__));
  or1   g2701(.dina(new_new_n8449__), .dinb(new_new_n8445__), .dout(new_new_n3643__));
  and1  g2702(.dina(new_new_n8447__), .dinb(new_new_n8442__), .dout(new_new_n3644__));
  or1   g2703(.dina(new_new_n8449__), .dinb(new_new_n8444__), .dout(new_new_n3645__));
  and1  g2704(.dina(new_new_n3645__), .dinb(new_new_n3643__), .dout(new_new_n3646__));
  or1   g2705(.dina(new_new_n3644__), .dinb(new_new_n3642__), .dout(new_new_n3647__));
  and1  g2706(.dina(new_new_n8396__), .dinb(new_new_n8362__), .dout(new_new_n3648__));
  or1   g2707(.dina(new_new_n8401__), .dinb(new_new_n8371__), .dout(new_new_n3649__));
  and1  g2708(.dina(new_new_n8450__), .dinb(new_new_n8451__), .dout(new_new_n3650__));
  or1   g2709(.dina(new_new_n8452__), .dinb(new_new_n8453__), .dout(new_new_n3651__));
  and1  g2710(.dina(new_new_n8455__), .dinb(new_new_n8446__), .dout(new_new_n3652__));
  or1   g2711(.dina(new_new_n8457__), .dinb(new_new_n8448__), .dout(new_new_n3653__));
  and1  g2712(.dina(new_new_n8458__), .dinb(new_new_n8459__), .dout(new_new_n3654__));
  or1   g2713(.dina(new_new_n8460__), .dinb(new_new_n8461__), .dout(new_new_n3655__));
  and1  g2714(.dina(new_new_n8462__), .dinb(new_new_n8463__), .dout(new_new_n3656__));
  or1   g2715(.dina(new_new_n8464__), .dinb(new_new_n8465__), .dout(new_new_n3657__));
  and1  g2716(.dina(new_new_n8467__), .dinb(new_new_n8462__), .dout(new_new_n3658__));
  or1   g2717(.dina(new_new_n8469__), .dinb(new_new_n8464__), .dout(new_new_n3659__));
  and1  g2718(.dina(new_new_n8467__), .dinb(new_new_n8463__), .dout(new_new_n3660__));
  or1   g2719(.dina(new_new_n8469__), .dinb(new_new_n8465__), .dout(new_new_n3661__));
  and1  g2720(.dina(new_new_n3661__), .dinb(new_new_n3659__), .dout(new_new_n3662__));
  or1   g2721(.dina(new_new_n3660__), .dinb(new_new_n3658__), .dout(new_new_n3663__));
  and1  g2722(.dina(new_new_n7716__), .dinb(new_new_n1537__), .dout(new_new_n3664__));
  or1   g2723(.dina(new_new_n7718__), .dinb(new_new_n1538__), .dout(new_new_n3665__));
  and1  g2724(.dina(new_new_n8470__), .dinb(new_new_n8471__), .dout(new_new_n3666__));
  or1   g2725(.dina(new_new_n8472__), .dinb(new_new_n8473__), .dout(new_new_n3667__));
  and1  g2726(.dina(new_new_n8475__), .dinb(new_new_n8471__), .dout(new_new_n3668__));
  or1   g2727(.dina(new_new_n8477__), .dinb(new_new_n8473__), .dout(new_new_n3669__));
  and1  g2728(.dina(new_new_n8475__), .dinb(new_new_n8470__), .dout(new_new_n3670__));
  or1   g2729(.dina(new_new_n8477__), .dinb(new_new_n8472__), .dout(new_new_n3671__));
  and1  g2730(.dina(new_new_n3671__), .dinb(new_new_n3669__), .dout(new_new_n3672__));
  or1   g2731(.dina(new_new_n3670__), .dinb(new_new_n3668__), .dout(new_new_n3673__));
  and1  g2732(.dina(new_new_n7085__), .dinb(new_new_n7704__), .dout(new_new_n3674__));
  or1   g2733(.dina(new_new_n7093__), .dinb(new_new_n7710__), .dout(new_new_n3675__));
  and1  g2734(.dina(new_new_n8478__), .dinb(new_new_n8479__), .dout(new_new_n3676__));
  or1   g2735(.dina(new_new_n8480__), .dinb(new_new_n8481__), .dout(new_new_n3677__));
  and1  g2736(.dina(new_new_n8483__), .dinb(new_new_n8479__), .dout(new_new_n3678__));
  or1   g2737(.dina(new_new_n8485__), .dinb(new_new_n8481__), .dout(new_new_n3679__));
  and1  g2738(.dina(new_new_n8483__), .dinb(new_new_n8478__), .dout(new_new_n3680__));
  or1   g2739(.dina(new_new_n8485__), .dinb(new_new_n8480__), .dout(new_new_n3681__));
  and1  g2740(.dina(new_new_n3681__), .dinb(new_new_n3679__), .dout(new_new_n3682__));
  or1   g2741(.dina(new_new_n3680__), .dinb(new_new_n3678__), .dout(new_new_n3683__));
  and1  g2742(.dina(new_new_n7732__), .dinb(new_new_n7724__), .dout(new_new_n3684__));
  or1   g2743(.dina(new_new_n7734__), .dinb(new_new_n7726__), .dout(new_new_n3685__));
  and1  g2744(.dina(new_new_n8486__), .dinb(new_new_n8487__), .dout(new_new_n3686__));
  or1   g2745(.dina(new_new_n8488__), .dinb(new_new_n8489__), .dout(new_new_n3687__));
  and1  g2746(.dina(new_new_n8491__), .dinb(new_new_n8487__), .dout(new_new_n3688__));
  or1   g2747(.dina(new_new_n8493__), .dinb(new_new_n8489__), .dout(new_new_n3689__));
  and1  g2748(.dina(new_new_n8491__), .dinb(new_new_n8486__), .dout(new_new_n3690__));
  or1   g2749(.dina(new_new_n8493__), .dinb(new_new_n8488__), .dout(new_new_n3691__));
  and1  g2750(.dina(new_new_n3691__), .dinb(new_new_n3689__), .dout(new_new_n3692__));
  or1   g2751(.dina(new_new_n3690__), .dinb(new_new_n3688__), .dout(new_new_n3693__));
  and1  g2752(.dina(new_new_n7673__), .dinb(new_new_n7106__), .dout(new_new_n3694__));
  or1   g2753(.dina(new_new_n7688__), .dinb(new_new_n7109__), .dout(new_new_n3695__));
  and1  g2754(.dina(new_new_n8494__), .dinb(new_new_n8495__), .dout(new_new_n3696__));
  or1   g2755(.dina(new_new_n8496__), .dinb(new_new_n8497__), .dout(new_new_n3697__));
  and1  g2756(.dina(new_new_n8499__), .dinb(new_new_n8495__), .dout(new_new_n3698__));
  or1   g2757(.dina(new_new_n8501__), .dinb(new_new_n8497__), .dout(new_new_n3699__));
  and1  g2758(.dina(new_new_n8499__), .dinb(new_new_n8494__), .dout(new_new_n3700__));
  or1   g2759(.dina(new_new_n8501__), .dinb(new_new_n8496__), .dout(new_new_n3701__));
  and1  g2760(.dina(new_new_n3701__), .dinb(new_new_n3699__), .dout(new_new_n3702__));
  or1   g2761(.dina(new_new_n3700__), .dinb(new_new_n3698__), .dout(new_new_n3703__));
  and1  g2762(.dina(new_new_n2907__), .dinb(new_new_n7741__), .dout(new_new_n3704__));
  or1   g2763(.dina(new_new_n8502__), .dinb(new_new_n7743__), .dout(new_new_n3705__));
  and1  g2764(.dina(new_new_n8503__), .dinb(new_new_n8504__), .dout(new_new_n3706__));
  or1   g2765(.dina(new_new_n8505__), .dinb(new_new_n8506__), .dout(new_new_n3707__));
  and1  g2766(.dina(new_new_n8508__), .dinb(new_new_n8504__), .dout(new_new_n3708__));
  or1   g2767(.dina(new_new_n8510__), .dinb(new_new_n8506__), .dout(new_new_n3709__));
  and1  g2768(.dina(new_new_n8508__), .dinb(new_new_n8503__), .dout(new_new_n3710__));
  or1   g2769(.dina(new_new_n8510__), .dinb(new_new_n8505__), .dout(new_new_n3711__));
  and1  g2770(.dina(new_new_n3711__), .dinb(new_new_n3709__), .dout(new_new_n3712__));
  or1   g2771(.dina(new_new_n3710__), .dinb(new_new_n3708__), .dout(new_new_n3713__));
  and1  g2772(.dina(new_new_n6867__), .dinb(new_new_n8363__), .dout(new_new_n3714__));
  or1   g2773(.dina(new_new_n6875__), .dinb(new_new_n8372__), .dout(new_new_n3715__));
  and1  g2774(.dina(new_new_n8511__), .dinb(new_new_n3135__), .dout(new_new_n3716__));
  or1   g2775(.dina(new_new_n3712__), .dinb(new_new_n8512__), .dout(new_new_n3717__));
  and1  g2776(.dina(new_new_n1524__), .dinb(new_new_n1505__), .dout(new_new_n3718__));
  or1   g2777(.dina(new_new_n1523__), .dinb(new_new_n1506__), .dout(new_new_n3719__));
  and1  g2778(.dina(new_new_n7617__), .dinb(new_new_n1323__), .dout(new_new_n3720__));
  or1   g2779(.dina(new_new_n7619__), .dinb(new_new_n1324__), .dout(new_new_n3721__));
  and1  g2780(.dina(new_new_n8513__), .dinb(new_new_n8514__), .dout(new_new_n3722__));
  or1   g2781(.dina(new_new_n8515__), .dinb(new_new_n8516__), .dout(new_new_n3723__));
  and1  g2782(.dina(new_new_n8518__), .dinb(new_new_n8514__), .dout(new_new_n3724__));
  or1   g2783(.dina(new_new_n8520__), .dinb(new_new_n8516__), .dout(new_new_n3725__));
  and1  g2784(.dina(new_new_n8518__), .dinb(new_new_n8513__), .dout(new_new_n3726__));
  or1   g2785(.dina(new_new_n8520__), .dinb(new_new_n8515__), .dout(new_new_n3727__));
  and1  g2786(.dina(new_new_n3727__), .dinb(new_new_n3725__), .dout(new_new_n3728__));
  or1   g2787(.dina(new_new_n3726__), .dinb(new_new_n3724__), .dout(new_new_n3729__));
  and1  g2788(.dina(new_new_n6951__), .dinb(new_new_n8523__), .dout(new_new_n3730__));
  or1   g2789(.dina(new_new_n6964__), .dinb(new_new_n8528__), .dout(new_new_n3731__));
  and1  g2790(.dina(new_new_n8530__), .dinb(new_new_n8531__), .dout(new_new_n3732__));
  or1   g2791(.dina(new_new_n8532__), .dinb(new_new_n8533__), .dout(new_new_n3733__));
  and1  g2792(.dina(new_new_n8535__), .dinb(new_new_n8531__), .dout(new_new_n3734__));
  or1   g2793(.dina(new_new_n8537__), .dinb(new_new_n8533__), .dout(new_new_n3735__));
  and1  g2794(.dina(new_new_n8535__), .dinb(new_new_n8530__), .dout(new_new_n3736__));
  or1   g2795(.dina(new_new_n8537__), .dinb(new_new_n8532__), .dout(new_new_n3737__));
  and1  g2796(.dina(new_new_n3737__), .dinb(new_new_n3735__), .dout(new_new_n3738__));
  or1   g2797(.dina(new_new_n3736__), .dinb(new_new_n3734__), .dout(new_new_n3739__));
  and1  g2798(.dina(new_new_n7641__), .dinb(new_new_n7625__), .dout(new_new_n3740__));
  or1   g2799(.dina(new_new_n7643__), .dinb(new_new_n7627__), .dout(new_new_n3741__));
  and1  g2800(.dina(new_new_n8538__), .dinb(new_new_n8539__), .dout(new_new_n3742__));
  or1   g2801(.dina(new_new_n8540__), .dinb(new_new_n8541__), .dout(new_new_n3743__));
  and1  g2802(.dina(new_new_n8543__), .dinb(new_new_n8539__), .dout(new_new_n3744__));
  or1   g2803(.dina(new_new_n8545__), .dinb(new_new_n8541__), .dout(new_new_n3745__));
  and1  g2804(.dina(new_new_n8543__), .dinb(new_new_n8538__), .dout(new_new_n3746__));
  or1   g2805(.dina(new_new_n8545__), .dinb(new_new_n8540__), .dout(new_new_n3747__));
  and1  g2806(.dina(new_new_n3747__), .dinb(new_new_n3745__), .dout(new_new_n3748__));
  or1   g2807(.dina(new_new_n3746__), .dinb(new_new_n3744__), .dout(new_new_n3749__));
  and1  g2808(.dina(new_new_n7631__), .dinb(new_new_n7027__), .dout(new_new_n3750__));
  or1   g2809(.dina(new_new_n7635__), .dinb(new_new_n7042__), .dout(new_new_n3751__));
  and1  g2810(.dina(new_new_n8546__), .dinb(new_new_n8547__), .dout(new_new_n3752__));
  or1   g2811(.dina(new_new_n8548__), .dinb(new_new_n8549__), .dout(new_new_n3753__));
  and1  g2812(.dina(new_new_n8551__), .dinb(new_new_n8547__), .dout(new_new_n3754__));
  or1   g2813(.dina(new_new_n8553__), .dinb(new_new_n8549__), .dout(new_new_n3755__));
  and1  g2814(.dina(new_new_n8551__), .dinb(new_new_n8546__), .dout(new_new_n3756__));
  or1   g2815(.dina(new_new_n8553__), .dinb(new_new_n8548__), .dout(new_new_n3757__));
  and1  g2816(.dina(new_new_n3757__), .dinb(new_new_n3755__), .dout(new_new_n3758__));
  or1   g2817(.dina(new_new_n3756__), .dinb(new_new_n3754__), .dout(new_new_n3759__));
  and1  g2818(.dina(new_new_n7657__), .dinb(new_new_n7649__), .dout(new_new_n3760__));
  or1   g2819(.dina(new_new_n7659__), .dinb(new_new_n7651__), .dout(new_new_n3761__));
  and1  g2820(.dina(new_new_n8554__), .dinb(new_new_n8555__), .dout(new_new_n3762__));
  or1   g2821(.dina(new_new_n8556__), .dinb(new_new_n8557__), .dout(new_new_n3763__));
  and1  g2822(.dina(new_new_n8559__), .dinb(new_new_n8555__), .dout(new_new_n3764__));
  or1   g2823(.dina(new_new_n8561__), .dinb(new_new_n8557__), .dout(new_new_n3765__));
  and1  g2824(.dina(new_new_n8559__), .dinb(new_new_n8554__), .dout(new_new_n3766__));
  or1   g2825(.dina(new_new_n8561__), .dinb(new_new_n8556__), .dout(new_new_n3767__));
  and1  g2826(.dina(new_new_n3767__), .dinb(new_new_n3765__), .dout(new_new_n3768__));
  or1   g2827(.dina(new_new_n3766__), .dinb(new_new_n3764__), .dout(new_new_n3769__));
  and1  g2828(.dina(new_new_n6970__), .dinb(new_new_n7598__), .dout(new_new_n3770__));
  or1   g2829(.dina(new_new_n6976__), .dinb(new_new_n7611__), .dout(new_new_n3771__));
  and1  g2830(.dina(new_new_n8562__), .dinb(new_new_n8563__), .dout(new_new_n3772__));
  or1   g2831(.dina(new_new_n8564__), .dinb(new_new_n8565__), .dout(new_new_n3773__));
  and1  g2832(.dina(new_new_n8567__), .dinb(new_new_n8563__), .dout(new_new_n3774__));
  or1   g2833(.dina(new_new_n8569__), .dinb(new_new_n8565__), .dout(new_new_n3775__));
  and1  g2834(.dina(new_new_n8567__), .dinb(new_new_n8562__), .dout(new_new_n3776__));
  or1   g2835(.dina(new_new_n8569__), .dinb(new_new_n8564__), .dout(new_new_n3777__));
  and1  g2836(.dina(new_new_n3777__), .dinb(new_new_n3775__), .dout(new_new_n3778__));
  or1   g2837(.dina(new_new_n3776__), .dinb(new_new_n3774__), .dout(new_new_n3779__));
  and1  g2838(.dina(new_new_n2863__), .dinb(new_new_n7666__), .dout(new_new_n3780__));
  or1   g2839(.dina(new_new_n8570__), .dinb(new_new_n7668__), .dout(new_new_n3781__));
  and1  g2840(.dina(new_new_n8571__), .dinb(new_new_n8572__), .dout(new_new_n3782__));
  or1   g2841(.dina(new_new_n8573__), .dinb(new_new_n8574__), .dout(new_new_n3783__));
  and1  g2842(.dina(new_new_n8576__), .dinb(new_new_n8572__), .dout(new_new_n3784__));
  or1   g2843(.dina(new_new_n8578__), .dinb(new_new_n8574__), .dout(new_new_n3785__));
  and1  g2844(.dina(new_new_n8576__), .dinb(new_new_n8571__), .dout(new_new_n3786__));
  or1   g2845(.dina(new_new_n8578__), .dinb(new_new_n8573__), .dout(new_new_n3787__));
  and1  g2846(.dina(new_new_n3787__), .dinb(new_new_n3785__), .dout(new_new_n3788__));
  or1   g2847(.dina(new_new_n3786__), .dinb(new_new_n3784__), .dout(new_new_n3789__));
  or1   g2848(.dina(new_new_n7448__), .dinb(new_new_n6893__), .dout(new_new_n3790__));
  or1   g2849(.dina(new_new_n7300__), .dinb(new_new_n6823__), .dout(new_new_n3791__));
  or1   g2850(.dina(new_new_n7151__), .dinb(new_new_n6784__), .dout(new_new_n3792__));
  or1   g2851(.dina(new_new_n8579__), .dinb(new_new_n3129__), .dout(new_new_n3793__));
  and1  g2852(.dina(new_new_n7230__), .dinb(new_new_n7226__), .dout(new_new_n3794__));
  or1   g2853(.dina(new_new_n7232__), .dinb(new_new_n7228__), .dout(new_new_n3795__));
  and1  g2854(.dina(new_new_n7229__), .dinb(new_new_n7225__), .dout(new_new_n3796__));
  or1   g2855(.dina(new_new_n7231__), .dinb(new_new_n7227__), .dout(new_new_n3797__));
  and1  g2856(.dina(new_new_n3797__), .dinb(new_new_n3795__), .dout(new_new_n3798__));
  or1   g2857(.dina(new_new_n3796__), .dinb(new_new_n3794__), .dout(new_new_n3799__));
  and1  g2858(.dina(new_new_n7761__), .dinb(new_new_n7753__), .dout(new_new_n3800__));
  or1   g2859(.dina(new_new_n7763__), .dinb(new_new_n7755__), .dout(new_new_n3801__));
  and1  g2860(.dina(new_new_n8580__), .dinb(new_new_n8581__), .dout(new_new_n3802__));
  or1   g2861(.dina(new_new_n8582__), .dinb(new_new_n8583__), .dout(new_new_n3803__));
  and1  g2862(.dina(new_new_n8585__), .dinb(new_new_n8581__), .dout(new_new_n3804__));
  or1   g2863(.dina(new_new_n8586__), .dinb(new_new_n8583__), .dout(new_new_n3805__));
  and1  g2864(.dina(new_new_n8585__), .dinb(new_new_n8580__), .dout(new_new_n3806__));
  or1   g2865(.dina(new_new_n8586__), .dinb(new_new_n8582__), .dout(new_new_n3807__));
  and1  g2866(.dina(new_new_n3807__), .dinb(new_new_n3805__), .dout(new_new_n3808__));
  or1   g2867(.dina(new_new_n3806__), .dinb(new_new_n3804__), .dout(new_new_n3809__));
  and1  g2868(.dina(new_new_n7247__), .dinb(new_new_n6770__), .dout(new_new_n3810__));
  or1   g2869(.dina(new_new_n7248__), .dinb(new_new_n6783__), .dout(new_new_n3811__));
  and1  g2870(.dina(new_new_n8587__), .dinb(new_new_n8588__), .dout(new_new_n3812__));
  or1   g2871(.dina(new_new_n8589__), .dinb(new_new_n8590__), .dout(new_new_n3813__));
  and1  g2872(.dina(new_new_n8592__), .dinb(new_new_n8588__), .dout(new_new_n3814__));
  or1   g2873(.dina(new_new_n8593__), .dinb(new_new_n8590__), .dout(new_new_n3815__));
  and1  g2874(.dina(new_new_n8592__), .dinb(new_new_n8587__), .dout(new_new_n3816__));
  or1   g2875(.dina(new_new_n8593__), .dinb(new_new_n8589__), .dout(new_new_n3817__));
  and1  g2876(.dina(new_new_n3817__), .dinb(new_new_n3815__), .dout(new_new_n3818__));
  or1   g2877(.dina(new_new_n3816__), .dinb(new_new_n3814__), .dout(new_new_n3819__));
  and1  g2878(.dina(new_new_n7777__), .dinb(new_new_n7769__), .dout(new_new_n3820__));
  or1   g2879(.dina(new_new_n7779__), .dinb(new_new_n7771__), .dout(new_new_n3821__));
  or1   g2880(.dina(new_new_n3820__), .dinb(new_new_n3818__), .dout(new_new_n3822__));
  and1  g2881(.dina(new_new_n7379__), .dinb(new_new_n7375__), .dout(new_new_n3823__));
  or1   g2882(.dina(new_new_n7381__), .dinb(new_new_n7377__), .dout(new_new_n3824__));
  and1  g2883(.dina(new_new_n7378__), .dinb(new_new_n7374__), .dout(new_new_n3825__));
  or1   g2884(.dina(new_new_n7380__), .dinb(new_new_n7376__), .dout(new_new_n3826__));
  and1  g2885(.dina(new_new_n3826__), .dinb(new_new_n3824__), .dout(new_new_n3827__));
  or1   g2886(.dina(new_new_n3825__), .dinb(new_new_n3823__), .dout(new_new_n3828__));
  and1  g2887(.dina(new_new_n7793__), .dinb(new_new_n7785__), .dout(new_new_n3829__));
  or1   g2888(.dina(new_new_n7795__), .dinb(new_new_n7787__), .dout(new_new_n3830__));
  and1  g2889(.dina(new_new_n8594__), .dinb(new_new_n8595__), .dout(new_new_n3831__));
  or1   g2890(.dina(new_new_n8596__), .dinb(new_new_n8597__), .dout(new_new_n3832__));
  and1  g2891(.dina(new_new_n8599__), .dinb(new_new_n8595__), .dout(new_new_n3833__));
  or1   g2892(.dina(new_new_n8600__), .dinb(new_new_n8597__), .dout(new_new_n3834__));
  and1  g2893(.dina(new_new_n8599__), .dinb(new_new_n8594__), .dout(new_new_n3835__));
  or1   g2894(.dina(new_new_n8600__), .dinb(new_new_n8596__), .dout(new_new_n3836__));
  and1  g2895(.dina(new_new_n3836__), .dinb(new_new_n3834__), .dout(new_new_n3837__));
  or1   g2896(.dina(new_new_n3835__), .dinb(new_new_n3833__), .dout(new_new_n3838__));
  and1  g2897(.dina(new_new_n7396__), .dinb(new_new_n6813__), .dout(new_new_n3839__));
  or1   g2898(.dina(new_new_n7397__), .dinb(new_new_n6823__), .dout(new_new_n3840__));
  and1  g2899(.dina(new_new_n8601__), .dinb(new_new_n8602__), .dout(new_new_n3841__));
  or1   g2900(.dina(new_new_n8603__), .dinb(new_new_n8604__), .dout(new_new_n3842__));
  and1  g2901(.dina(new_new_n8606__), .dinb(new_new_n8602__), .dout(new_new_n3843__));
  or1   g2902(.dina(new_new_n8607__), .dinb(new_new_n8604__), .dout(new_new_n3844__));
  and1  g2903(.dina(new_new_n8606__), .dinb(new_new_n8601__), .dout(new_new_n3845__));
  or1   g2904(.dina(new_new_n8607__), .dinb(new_new_n8603__), .dout(new_new_n3846__));
  and1  g2905(.dina(new_new_n3846__), .dinb(new_new_n3844__), .dout(new_new_n3847__));
  or1   g2906(.dina(new_new_n3845__), .dinb(new_new_n3843__), .dout(new_new_n3848__));
  and1  g2907(.dina(new_new_n7809__), .dinb(new_new_n7801__), .dout(new_new_n3849__));
  or1   g2908(.dina(new_new_n7811__), .dinb(new_new_n7803__), .dout(new_new_n3850__));
  or1   g2909(.dina(new_new_n3849__), .dinb(new_new_n3847__), .dout(new_new_n3851__));
  and1  g2910(.dina(new_new_n7526__), .dinb(new_new_n7522__), .dout(new_new_n3852__));
  or1   g2911(.dina(new_new_n7528__), .dinb(new_new_n7524__), .dout(new_new_n3853__));
  and1  g2912(.dina(new_new_n7525__), .dinb(new_new_n7521__), .dout(new_new_n3854__));
  or1   g2913(.dina(new_new_n7527__), .dinb(new_new_n7523__), .dout(new_new_n3855__));
  and1  g2914(.dina(new_new_n3855__), .dinb(new_new_n3853__), .dout(new_new_n3856__));
  or1   g2915(.dina(new_new_n3854__), .dinb(new_new_n3852__), .dout(new_new_n3857__));
  and1  g2916(.dina(new_new_n7845__), .dinb(new_new_n7837__), .dout(new_new_n3858__));
  or1   g2917(.dina(new_new_n7847__), .dinb(new_new_n7839__), .dout(new_new_n3859__));
  and1  g2918(.dina(new_new_n8608__), .dinb(new_new_n8609__), .dout(new_new_n3860__));
  or1   g2919(.dina(new_new_n8610__), .dinb(new_new_n8611__), .dout(new_new_n3861__));
  and1  g2920(.dina(new_new_n8613__), .dinb(new_new_n8609__), .dout(new_new_n3862__));
  or1   g2921(.dina(new_new_n8614__), .dinb(new_new_n8611__), .dout(new_new_n3863__));
  and1  g2922(.dina(new_new_n8613__), .dinb(new_new_n8608__), .dout(new_new_n3864__));
  or1   g2923(.dina(new_new_n8614__), .dinb(new_new_n8610__), .dout(new_new_n3865__));
  and1  g2924(.dina(new_new_n3865__), .dinb(new_new_n3863__), .dout(new_new_n3866__));
  or1   g2925(.dina(new_new_n3864__), .dinb(new_new_n3862__), .dout(new_new_n3867__));
  and1  g2926(.dina(new_new_n7821__), .dinb(new_new_n6887__), .dout(new_new_n3868__));
  or1   g2927(.dina(new_new_n7823__), .dinb(new_new_n6892__), .dout(new_new_n3869__));
  and1  g2928(.dina(new_new_n8615__), .dinb(new_new_n8616__), .dout(new_new_n3870__));
  or1   g2929(.dina(new_new_n8617__), .dinb(new_new_n8618__), .dout(new_new_n3871__));
  and1  g2930(.dina(new_new_n8620__), .dinb(new_new_n8616__), .dout(new_new_n3872__));
  or1   g2931(.dina(new_new_n8621__), .dinb(new_new_n8618__), .dout(new_new_n3873__));
  and1  g2932(.dina(new_new_n8620__), .dinb(new_new_n8615__), .dout(new_new_n3874__));
  or1   g2933(.dina(new_new_n8621__), .dinb(new_new_n8617__), .dout(new_new_n3875__));
  and1  g2934(.dina(new_new_n3875__), .dinb(new_new_n3873__), .dout(new_new_n3876__));
  or1   g2935(.dina(new_new_n3874__), .dinb(new_new_n3872__), .dout(new_new_n3877__));
  and1  g2936(.dina(new_new_n7877__), .dinb(new_new_n7869__), .dout(new_new_n3878__));
  or1   g2937(.dina(new_new_n7879__), .dinb(new_new_n7871__), .dout(new_new_n3879__));
  or1   g2938(.dina(new_new_n3878__), .dinb(new_new_n3876__), .dout(new_new_n3880__));
  and1  g2939(.dina(new_new_n8623__), .dinb(new_new_n2910__), .dout(new_new_n3881__));
  and1  g2940(.dina(new_new_n8623__), .dinb(new_new_n2912__), .dout(new_new_n3882__));
  or1   g2941(.dina(new_new_n3882__), .dinb(new_new_n3881__), .dout(new_new_n3883__));
  and1  g2942(.dina(new_new_n8625__), .dinb(new_new_n2959__), .dout(new_new_n3884__));
  and1  g2943(.dina(new_new_n8625__), .dinb(new_new_n2961__), .dout(new_new_n3885__));
  or1   g2944(.dina(new_new_n3885__), .dinb(new_new_n3884__), .dout(new_new_n3886__));
  and1  g2945(.dina(new_new_n8627__), .dinb(new_new_n3008__), .dout(new_new_n3887__));
  and1  g2946(.dina(new_new_n8627__), .dinb(new_new_n3010__), .dout(new_new_n3888__));
  or1   g2947(.dina(new_new_n3888__), .dinb(new_new_n3887__), .dout(new_new_n3889__));
  and1  g2948(.dina(new_new_n8629__), .dinb(new_new_n3097__), .dout(new_new_n3890__));
  and1  g2949(.dina(new_new_n8629__), .dinb(new_new_n3119__), .dout(new_new_n3891__));
  or1   g2950(.dina(new_new_n3891__), .dinb(new_new_n3890__), .dout(new_new_n3892__));
  and1  g2951(.dina(new_new_n8630__), .dinb(new_new_n3715__), .dout(new_new_n3893__));
  or1   g2952(.dina(new_new_n3788__), .dinb(new_new_n8631__), .dout(new_new_n3894__));
  and1  g2953(.dina(new_new_n6951__), .dinb(new_new_n7942__), .dout(new_new_n3895__));
  or1   g2954(.dina(new_new_n6964__), .dinb(new_new_n7945__), .dout(new_new_n3896__));
  and1  g2955(.dina(new_new_n7979__), .dinb(new_new_n7971__), .dout(new_new_n3897__));
  or1   g2956(.dina(new_new_n7981__), .dinb(new_new_n7973__), .dout(new_new_n3898__));
  and1  g2957(.dina(new_new_n8632__), .dinb(new_new_n8633__), .dout(new_new_n3899__));
  or1   g2958(.dina(new_new_n8634__), .dinb(new_new_n8635__), .dout(new_new_n3900__));
  and1  g2959(.dina(new_new_n8637__), .dinb(new_new_n8633__), .dout(new_new_n3901__));
  or1   g2960(.dina(new_new_n8639__), .dinb(new_new_n8635__), .dout(new_new_n3902__));
  and1  g2961(.dina(new_new_n8637__), .dinb(new_new_n8632__), .dout(new_new_n3903__));
  or1   g2962(.dina(new_new_n8639__), .dinb(new_new_n8634__), .dout(new_new_n3904__));
  and1  g2963(.dina(new_new_n3904__), .dinb(new_new_n3902__), .dout(new_new_n3905__));
  or1   g2964(.dina(new_new_n3903__), .dinb(new_new_n3901__), .dout(new_new_n3906__));
  and1  g2965(.dina(new_new_n7956__), .dinb(new_new_n7029__), .dout(new_new_n3907__));
  or1   g2966(.dina(new_new_n7957__), .dinb(new_new_n7044__), .dout(new_new_n3908__));
  and1  g2967(.dina(new_new_n8640__), .dinb(new_new_n8641__), .dout(new_new_n3909__));
  or1   g2968(.dina(new_new_n8642__), .dinb(new_new_n8643__), .dout(new_new_n3910__));
  and1  g2969(.dina(new_new_n8645__), .dinb(new_new_n8641__), .dout(new_new_n3911__));
  or1   g2970(.dina(new_new_n8647__), .dinb(new_new_n8643__), .dout(new_new_n3912__));
  and1  g2971(.dina(new_new_n8645__), .dinb(new_new_n8640__), .dout(new_new_n3913__));
  or1   g2972(.dina(new_new_n8647__), .dinb(new_new_n8642__), .dout(new_new_n3914__));
  and1  g2973(.dina(new_new_n3914__), .dinb(new_new_n3912__), .dout(new_new_n3915__));
  or1   g2974(.dina(new_new_n3913__), .dinb(new_new_n3911__), .dout(new_new_n3916__));
  and1  g2975(.dina(new_new_n8025__), .dinb(new_new_n8017__), .dout(new_new_n3917__));
  or1   g2976(.dina(new_new_n8027__), .dinb(new_new_n8019__), .dout(new_new_n3918__));
  or1   g2977(.dina(new_new_n3917__), .dinb(new_new_n3915__), .dout(new_new_n3919__));
  and1  g2978(.dina(new_new_n8051__), .dinb(new_new_n8047__), .dout(new_new_n3920__));
  or1   g2979(.dina(new_new_n8053__), .dinb(new_new_n8049__), .dout(new_new_n3921__));
  and1  g2980(.dina(new_new_n8050__), .dinb(new_new_n8046__), .dout(new_new_n3922__));
  or1   g2981(.dina(new_new_n8052__), .dinb(new_new_n8048__), .dout(new_new_n3923__));
  and1  g2982(.dina(new_new_n3923__), .dinb(new_new_n3921__), .dout(new_new_n3924__));
  or1   g2983(.dina(new_new_n3922__), .dinb(new_new_n3920__), .dout(new_new_n3925__));
  and1  g2984(.dina(new_new_n8091__), .dinb(new_new_n8078__), .dout(new_new_n3926__));
  or1   g2985(.dina(new_new_n8093__), .dinb(new_new_n8080__), .dout(new_new_n3927__));
  and1  g2986(.dina(new_new_n8648__), .dinb(new_new_n8649__), .dout(new_new_n3928__));
  or1   g2987(.dina(new_new_n8650__), .dinb(new_new_n8651__), .dout(new_new_n3929__));
  and1  g2988(.dina(new_new_n8653__), .dinb(new_new_n8649__), .dout(new_new_n3930__));
  or1   g2989(.dina(new_new_n8655__), .dinb(new_new_n8651__), .dout(new_new_n3931__));
  and1  g2990(.dina(new_new_n8653__), .dinb(new_new_n8648__), .dout(new_new_n3932__));
  or1   g2991(.dina(new_new_n8655__), .dinb(new_new_n8650__), .dout(new_new_n3933__));
  and1  g2992(.dina(new_new_n3933__), .dinb(new_new_n3931__), .dout(new_new_n3934__));
  or1   g2993(.dina(new_new_n3932__), .dinb(new_new_n3930__), .dout(new_new_n3935__));
  and1  g2994(.dina(new_new_n8083__), .dinb(new_new_n7029__), .dout(new_new_n3936__));
  or1   g2995(.dina(new_new_n8086__), .dinb(new_new_n7044__), .dout(new_new_n3937__));
  and1  g2996(.dina(new_new_n8656__), .dinb(new_new_n8657__), .dout(new_new_n3938__));
  or1   g2997(.dina(new_new_n8658__), .dinb(new_new_n8659__), .dout(new_new_n3939__));
  and1  g2998(.dina(new_new_n8661__), .dinb(new_new_n8657__), .dout(new_new_n3940__));
  or1   g2999(.dina(new_new_n8663__), .dinb(new_new_n8659__), .dout(new_new_n3941__));
  and1  g3000(.dina(new_new_n8661__), .dinb(new_new_n8656__), .dout(new_new_n3942__));
  or1   g3001(.dina(new_new_n8663__), .dinb(new_new_n8658__), .dout(new_new_n3943__));
  and1  g3002(.dina(new_new_n3943__), .dinb(new_new_n3941__), .dout(new_new_n3944__));
  or1   g3003(.dina(new_new_n3942__), .dinb(new_new_n3940__), .dout(new_new_n3945__));
  and1  g3004(.dina(new_new_n8128__), .dinb(new_new_n8120__), .dout(new_new_n3946__));
  or1   g3005(.dina(new_new_n8130__), .dinb(new_new_n8122__), .dout(new_new_n3947__));
  and1  g3006(.dina(new_new_n8664__), .dinb(new_new_n8665__), .dout(new_new_n3948__));
  or1   g3007(.dina(new_new_n8666__), .dinb(new_new_n8667__), .dout(new_new_n3949__));
  and1  g3008(.dina(new_new_n8669__), .dinb(new_new_n8665__), .dout(new_new_n3950__));
  or1   g3009(.dina(new_new_n8671__), .dinb(new_new_n8667__), .dout(new_new_n3951__));
  and1  g3010(.dina(new_new_n8669__), .dinb(new_new_n8664__), .dout(new_new_n3952__));
  or1   g3011(.dina(new_new_n8671__), .dinb(new_new_n8666__), .dout(new_new_n3953__));
  and1  g3012(.dina(new_new_n3953__), .dinb(new_new_n3951__), .dout(new_new_n3954__));
  or1   g3013(.dina(new_new_n3952__), .dinb(new_new_n3950__), .dout(new_new_n3955__));
  and1  g3014(.dina(new_new_n8105__), .dinb(new_new_n7598__), .dout(new_new_n3956__));
  or1   g3015(.dina(new_new_n8106__), .dinb(new_new_n7611__), .dout(new_new_n3957__));
  and1  g3016(.dina(new_new_n8672__), .dinb(new_new_n8673__), .dout(new_new_n3958__));
  or1   g3017(.dina(new_new_n8674__), .dinb(new_new_n8675__), .dout(new_new_n3959__));
  and1  g3018(.dina(new_new_n8677__), .dinb(new_new_n8673__), .dout(new_new_n3960__));
  or1   g3019(.dina(new_new_n8679__), .dinb(new_new_n8675__), .dout(new_new_n3961__));
  and1  g3020(.dina(new_new_n8677__), .dinb(new_new_n8672__), .dout(new_new_n3962__));
  or1   g3021(.dina(new_new_n8679__), .dinb(new_new_n8674__), .dout(new_new_n3963__));
  and1  g3022(.dina(new_new_n3963__), .dinb(new_new_n3961__), .dout(new_new_n3964__));
  or1   g3023(.dina(new_new_n3962__), .dinb(new_new_n3960__), .dout(new_new_n3965__));
  and1  g3024(.dina(new_new_n8174__), .dinb(new_new_n8166__), .dout(new_new_n3966__));
  or1   g3025(.dina(new_new_n8176__), .dinb(new_new_n8168__), .dout(new_new_n3967__));
  or1   g3026(.dina(new_new_n3966__), .dinb(new_new_n3964__), .dout(new_new_n3968__));
  and1  g3027(.dina(new_new_n8200__), .dinb(new_new_n8196__), .dout(new_new_n3969__));
  or1   g3028(.dina(new_new_n8202__), .dinb(new_new_n8198__), .dout(new_new_n3970__));
  and1  g3029(.dina(new_new_n8199__), .dinb(new_new_n8195__), .dout(new_new_n3971__));
  or1   g3030(.dina(new_new_n8201__), .dinb(new_new_n8197__), .dout(new_new_n3972__));
  and1  g3031(.dina(new_new_n3972__), .dinb(new_new_n3970__), .dout(new_new_n3973__));
  or1   g3032(.dina(new_new_n3971__), .dinb(new_new_n3969__), .dout(new_new_n3974__));
  and1  g3033(.dina(new_new_n8248__), .dinb(new_new_n8235__), .dout(new_new_n3975__));
  or1   g3034(.dina(new_new_n8250__), .dinb(new_new_n8237__), .dout(new_new_n3976__));
  and1  g3035(.dina(new_new_n8680__), .dinb(new_new_n8681__), .dout(new_new_n3977__));
  or1   g3036(.dina(new_new_n8682__), .dinb(new_new_n8683__), .dout(new_new_n3978__));
  and1  g3037(.dina(new_new_n8685__), .dinb(new_new_n8681__), .dout(new_new_n3979__));
  or1   g3038(.dina(new_new_n8687__), .dinb(new_new_n8683__), .dout(new_new_n3980__));
  and1  g3039(.dina(new_new_n8685__), .dinb(new_new_n8680__), .dout(new_new_n3981__));
  or1   g3040(.dina(new_new_n8687__), .dinb(new_new_n8682__), .dout(new_new_n3982__));
  and1  g3041(.dina(new_new_n3982__), .dinb(new_new_n3980__), .dout(new_new_n3983__));
  or1   g3042(.dina(new_new_n3981__), .dinb(new_new_n3979__), .dout(new_new_n3984__));
  and1  g3043(.dina(new_new_n8240__), .dinb(new_new_n7601__), .dout(new_new_n3985__));
  or1   g3044(.dina(new_new_n8243__), .dinb(new_new_n7614__), .dout(new_new_n3986__));
  and1  g3045(.dina(new_new_n8688__), .dinb(new_new_n8689__), .dout(new_new_n3987__));
  or1   g3046(.dina(new_new_n8690__), .dinb(new_new_n8691__), .dout(new_new_n3988__));
  and1  g3047(.dina(new_new_n8693__), .dinb(new_new_n8689__), .dout(new_new_n3989__));
  or1   g3048(.dina(new_new_n8695__), .dinb(new_new_n8691__), .dout(new_new_n3990__));
  and1  g3049(.dina(new_new_n8693__), .dinb(new_new_n8688__), .dout(new_new_n3991__));
  or1   g3050(.dina(new_new_n8695__), .dinb(new_new_n8690__), .dout(new_new_n3992__));
  and1  g3051(.dina(new_new_n3992__), .dinb(new_new_n3990__), .dout(new_new_n3993__));
  or1   g3052(.dina(new_new_n3991__), .dinb(new_new_n3989__), .dout(new_new_n3994__));
  and1  g3053(.dina(new_new_n8295__), .dinb(new_new_n8287__), .dout(new_new_n3995__));
  or1   g3054(.dina(new_new_n8297__), .dinb(new_new_n8289__), .dout(new_new_n3996__));
  and1  g3055(.dina(new_new_n8696__), .dinb(new_new_n8697__), .dout(new_new_n3997__));
  or1   g3056(.dina(new_new_n8698__), .dinb(new_new_n8699__), .dout(new_new_n3998__));
  and1  g3057(.dina(new_new_n8701__), .dinb(new_new_n8697__), .dout(new_new_n3999__));
  or1   g3058(.dina(new_new_n8703__), .dinb(new_new_n8699__), .dout(new_new_n4000__));
  and1  g3059(.dina(new_new_n8701__), .dinb(new_new_n8696__), .dout(new_new_n4001__));
  or1   g3060(.dina(new_new_n8703__), .dinb(new_new_n8698__), .dout(new_new_n4002__));
  and1  g3061(.dina(new_new_n4002__), .dinb(new_new_n4000__), .dout(new_new_n4003__));
  or1   g3062(.dina(new_new_n4001__), .dinb(new_new_n3999__), .dout(new_new_n4004__));
  and1  g3063(.dina(new_new_n8255__), .dinb(new_new_n8363__), .dout(new_new_n4005__));
  or1   g3064(.dina(new_new_n8258__), .dinb(new_new_n8372__), .dout(new_new_n4006__));
  and1  g3065(.dina(new_new_n8704__), .dinb(new_new_n8705__), .dout(new_new_n4007__));
  or1   g3066(.dina(new_new_n8706__), .dinb(new_new_n8707__), .dout(new_new_n4008__));
  and1  g3067(.dina(new_new_n8709__), .dinb(new_new_n8705__), .dout(new_new_n4009__));
  or1   g3068(.dina(new_new_n8711__), .dinb(new_new_n8707__), .dout(new_new_n4010__));
  and1  g3069(.dina(new_new_n8709__), .dinb(new_new_n8704__), .dout(new_new_n4011__));
  or1   g3070(.dina(new_new_n8711__), .dinb(new_new_n8706__), .dout(new_new_n4012__));
  and1  g3071(.dina(new_new_n4012__), .dinb(new_new_n4010__), .dout(new_new_n4013__));
  or1   g3072(.dina(new_new_n4011__), .dinb(new_new_n4009__), .dout(new_new_n4014__));
  and1  g3073(.dina(new_new_n8381__), .dinb(new_new_n8355__), .dout(new_new_n4015__));
  or1   g3074(.dina(new_new_n8383__), .dinb(new_new_n8357__), .dout(new_new_n4016__));
  or1   g3075(.dina(new_new_n4015__), .dinb(new_new_n4013__), .dout(new_new_n4017__));
  and1  g3076(.dina(new_new_n8439__), .dinb(new_new_n8435__), .dout(new_new_n4018__));
  or1   g3077(.dina(new_new_n8441__), .dinb(new_new_n8437__), .dout(new_new_n4019__));
  and1  g3078(.dina(new_new_n8438__), .dinb(new_new_n8434__), .dout(new_new_n4020__));
  or1   g3079(.dina(new_new_n8440__), .dinb(new_new_n8436__), .dout(new_new_n4021__));
  and1  g3080(.dina(new_new_n4021__), .dinb(new_new_n4019__), .dout(new_new_n4022__));
  or1   g3081(.dina(new_new_n4020__), .dinb(new_new_n4018__), .dout(new_new_n4023__));
  and1  g3082(.dina(new_new_n8423__), .dinb(new_new_n8419__), .dout(new_new_n4024__));
  or1   g3083(.dina(new_new_n8425__), .dinb(new_new_n8421__), .dout(new_new_n4025__));
  and1  g3084(.dina(new_new_n8422__), .dinb(new_new_n8418__), .dout(new_new_n4026__));
  or1   g3085(.dina(new_new_n8424__), .dinb(new_new_n8420__), .dout(new_new_n4027__));
  and1  g3086(.dina(new_new_n4027__), .dinb(new_new_n4025__), .dout(new_new_n4028__));
  or1   g3087(.dina(new_new_n4026__), .dinb(new_new_n4024__), .dout(new_new_n4029__));
  and1  g3088(.dina(new_new_n8407__), .dinb(new_new_n8403__), .dout(new_new_n4030__));
  or1   g3089(.dina(new_new_n8409__), .dinb(new_new_n8405__), .dout(new_new_n4031__));
  and1  g3090(.dina(new_new_n8406__), .dinb(new_new_n8402__), .dout(new_new_n4032__));
  or1   g3091(.dina(new_new_n8408__), .dinb(new_new_n8404__), .dout(new_new_n4033__));
  and1  g3092(.dina(new_new_n4033__), .dinb(new_new_n4031__), .dout(new_new_n4034__));
  or1   g3093(.dina(new_new_n4032__), .dinb(new_new_n4030__), .dout(new_new_n4035__));
  and1  g3094(.dina(new_new_n8534__), .dinb(new_new_n8517__), .dout(new_new_n4036__));
  or1   g3095(.dina(new_new_n8536__), .dinb(new_new_n8519__), .dout(new_new_n4037__));
  and1  g3096(.dina(new_new_n8712__), .dinb(new_new_n8713__), .dout(new_new_n4038__));
  or1   g3097(.dina(new_new_n8714__), .dinb(new_new_n8715__), .dout(new_new_n4039__));
  and1  g3098(.dina(new_new_n8717__), .dinb(new_new_n8713__), .dout(new_new_n4040__));
  or1   g3099(.dina(new_new_n8719__), .dinb(new_new_n8715__), .dout(new_new_n4041__));
  and1  g3100(.dina(new_new_n8717__), .dinb(new_new_n8712__), .dout(new_new_n4042__));
  or1   g3101(.dina(new_new_n8719__), .dinb(new_new_n8714__), .dout(new_new_n4043__));
  and1  g3102(.dina(new_new_n4043__), .dinb(new_new_n4041__), .dout(new_new_n4044__));
  or1   g3103(.dina(new_new_n4042__), .dinb(new_new_n4040__), .dout(new_new_n4045__));
  and1  g3104(.dina(new_new_n8523__), .dinb(new_new_n7030__), .dout(new_new_n4046__));
  or1   g3105(.dina(new_new_n8528__), .dinb(new_new_n7045__), .dout(new_new_n4047__));
  and1  g3106(.dina(new_new_n8720__), .dinb(new_new_n8721__), .dout(new_new_n4048__));
  or1   g3107(.dina(new_new_n8722__), .dinb(new_new_n8723__), .dout(new_new_n4049__));
  and1  g3108(.dina(new_new_n8725__), .dinb(new_new_n8716__), .dout(new_new_n4050__));
  or1   g3109(.dina(new_new_n8727__), .dinb(new_new_n8718__), .dout(new_new_n4051__));
  and1  g3110(.dina(new_new_n8728__), .dinb(new_new_n8729__), .dout(new_new_n4052__));
  or1   g3111(.dina(new_new_n8730__), .dinb(new_new_n8731__), .dout(new_new_n4053__));
  and1  g3112(.dina(new_new_n8733__), .dinb(new_new_n8729__), .dout(new_new_n4054__));
  or1   g3113(.dina(new_new_n8735__), .dinb(new_new_n8731__), .dout(new_new_n4055__));
  and1  g3114(.dina(new_new_n8733__), .dinb(new_new_n8728__), .dout(new_new_n4056__));
  or1   g3115(.dina(new_new_n8735__), .dinb(new_new_n8730__), .dout(new_new_n4057__));
  and1  g3116(.dina(new_new_n4057__), .dinb(new_new_n4055__), .dout(new_new_n4058__));
  or1   g3117(.dina(new_new_n4056__), .dinb(new_new_n4054__), .dout(new_new_n4059__));
  and1  g3118(.dina(new_new_n8524__), .dinb(new_new_n7601__), .dout(new_new_n4060__));
  or1   g3119(.dina(new_new_n8527__), .dinb(new_new_n7614__), .dout(new_new_n4061__));
  and1  g3120(.dina(new_new_n8736__), .dinb(new_new_n8737__), .dout(new_new_n4062__));
  or1   g3121(.dina(new_new_n8738__), .dinb(new_new_n8739__), .dout(new_new_n4063__));
  and1  g3122(.dina(new_new_n8741__), .dinb(new_new_n8732__), .dout(new_new_n4064__));
  or1   g3123(.dina(new_new_n8743__), .dinb(new_new_n8734__), .dout(new_new_n4065__));
  and1  g3124(.dina(new_new_n8744__), .dinb(new_new_n8745__), .dout(new_new_n4066__));
  or1   g3125(.dina(new_new_n8746__), .dinb(new_new_n8747__), .dout(new_new_n4067__));
  and1  g3126(.dina(new_new_n8749__), .dinb(new_new_n8745__), .dout(new_new_n4068__));
  or1   g3127(.dina(new_new_n8751__), .dinb(new_new_n8747__), .dout(new_new_n4069__));
  and1  g3128(.dina(new_new_n8749__), .dinb(new_new_n8744__), .dout(new_new_n4070__));
  or1   g3129(.dina(new_new_n8751__), .dinb(new_new_n8746__), .dout(new_new_n4071__));
  and1  g3130(.dina(new_new_n4071__), .dinb(new_new_n4069__), .dout(new_new_n4072__));
  or1   g3131(.dina(new_new_n4070__), .dinb(new_new_n4068__), .dout(new_new_n4073__));
  and1  g3132(.dina(new_new_n8524__), .dinb(new_new_n8364__), .dout(new_new_n4074__));
  or1   g3133(.dina(new_new_n8529__), .dinb(new_new_n8373__), .dout(new_new_n4075__));
  and1  g3134(.dina(new_new_n8752__), .dinb(new_new_n8753__), .dout(new_new_n4076__));
  or1   g3135(.dina(new_new_n8754__), .dinb(new_new_n8755__), .dout(new_new_n4077__));
  and1  g3136(.dina(new_new_n8757__), .dinb(new_new_n8753__), .dout(new_new_n4078__));
  or1   g3137(.dina(new_new_n8759__), .dinb(new_new_n8755__), .dout(new_new_n4079__));
  and1  g3138(.dina(new_new_n8757__), .dinb(new_new_n8752__), .dout(new_new_n4080__));
  or1   g3139(.dina(new_new_n8759__), .dinb(new_new_n8754__), .dout(new_new_n4081__));
  and1  g3140(.dina(new_new_n4081__), .dinb(new_new_n4079__), .dout(new_new_n4082__));
  or1   g3141(.dina(new_new_n4080__), .dinb(new_new_n4078__), .dout(new_new_n4083__));
  and1  g3142(.dina(new_new_n8741__), .dinb(new_new_n8737__), .dout(new_new_n4084__));
  or1   g3143(.dina(new_new_n8743__), .dinb(new_new_n8739__), .dout(new_new_n4085__));
  and1  g3144(.dina(new_new_n8740__), .dinb(new_new_n8736__), .dout(new_new_n4086__));
  or1   g3145(.dina(new_new_n8742__), .dinb(new_new_n8738__), .dout(new_new_n4087__));
  and1  g3146(.dina(new_new_n4087__), .dinb(new_new_n4085__), .dout(new_new_n4088__));
  or1   g3147(.dina(new_new_n4086__), .dinb(new_new_n4084__), .dout(new_new_n4089__));
  and1  g3148(.dina(new_new_n8725__), .dinb(new_new_n8721__), .dout(new_new_n4090__));
  or1   g3149(.dina(new_new_n8727__), .dinb(new_new_n8723__), .dout(new_new_n4091__));
  and1  g3150(.dina(new_new_n8724__), .dinb(new_new_n8720__), .dout(new_new_n4092__));
  or1   g3151(.dina(new_new_n8726__), .dinb(new_new_n8722__), .dout(new_new_n4093__));
  and1  g3152(.dina(new_new_n4093__), .dinb(new_new_n4091__), .dout(new_new_n4094__));
  or1   g3153(.dina(new_new_n4092__), .dinb(new_new_n4090__), .dout(new_new_n4095__));
  and1  g3154(.dina(new_new_n8550__), .dinb(new_new_n8542__), .dout(new_new_n4096__));
  or1   g3155(.dina(new_new_n8552__), .dinb(new_new_n8544__), .dout(new_new_n4097__));
  and1  g3156(.dina(new_new_n8760__), .dinb(new_new_n8761__), .dout(new_new_n4098__));
  or1   g3157(.dina(new_new_n8762__), .dinb(new_new_n8763__), .dout(new_new_n4099__));
  and1  g3158(.dina(new_new_n8765__), .dinb(new_new_n8761__), .dout(new_new_n4100__));
  or1   g3159(.dina(new_new_n8767__), .dinb(new_new_n8763__), .dout(new_new_n4101__));
  and1  g3160(.dina(new_new_n8765__), .dinb(new_new_n8760__), .dout(new_new_n4102__));
  or1   g3161(.dina(new_new_n8767__), .dinb(new_new_n8762__), .dout(new_new_n4103__));
  and1  g3162(.dina(new_new_n4103__), .dinb(new_new_n4101__), .dout(new_new_n4104__));
  or1   g3163(.dina(new_new_n4102__), .dinb(new_new_n4100__), .dout(new_new_n4105__));
  and1  g3164(.dina(new_new_n7630__), .dinb(new_new_n7602__), .dout(new_new_n4106__));
  or1   g3165(.dina(new_new_n7634__), .dinb(new_new_n7615__), .dout(new_new_n4107__));
  and1  g3166(.dina(new_new_n8768__), .dinb(new_new_n8769__), .dout(new_new_n4108__));
  or1   g3167(.dina(new_new_n8770__), .dinb(new_new_n8771__), .dout(new_new_n4109__));
  and1  g3168(.dina(new_new_n8773__), .dinb(new_new_n8764__), .dout(new_new_n4110__));
  or1   g3169(.dina(new_new_n8775__), .dinb(new_new_n8766__), .dout(new_new_n4111__));
  and1  g3170(.dina(new_new_n8776__), .dinb(new_new_n8777__), .dout(new_new_n4112__));
  or1   g3171(.dina(new_new_n8778__), .dinb(new_new_n8779__), .dout(new_new_n4113__));
  and1  g3172(.dina(new_new_n8781__), .dinb(new_new_n8777__), .dout(new_new_n4114__));
  or1   g3173(.dina(new_new_n8783__), .dinb(new_new_n8779__), .dout(new_new_n4115__));
  and1  g3174(.dina(new_new_n8781__), .dinb(new_new_n8776__), .dout(new_new_n4116__));
  or1   g3175(.dina(new_new_n8783__), .dinb(new_new_n8778__), .dout(new_new_n4117__));
  and1  g3176(.dina(new_new_n4117__), .dinb(new_new_n4115__), .dout(new_new_n4118__));
  or1   g3177(.dina(new_new_n4116__), .dinb(new_new_n4114__), .dout(new_new_n4119__));
  and1  g3178(.dina(new_new_n7632__), .dinb(new_new_n8364__), .dout(new_new_n4120__));
  or1   g3179(.dina(new_new_n7636__), .dinb(new_new_n8373__), .dout(new_new_n4121__));
  and1  g3180(.dina(new_new_n8784__), .dinb(new_new_n8785__), .dout(new_new_n4122__));
  or1   g3181(.dina(new_new_n8786__), .dinb(new_new_n8787__), .dout(new_new_n4123__));
  and1  g3182(.dina(new_new_n8789__), .dinb(new_new_n8780__), .dout(new_new_n4124__));
  or1   g3183(.dina(new_new_n8791__), .dinb(new_new_n8782__), .dout(new_new_n4125__));
  or1   g3184(.dina(new_new_n4124__), .dinb(new_new_n4082__), .dout(new_new_n4126__));
  and1  g3185(.dina(new_new_n7087__), .dinb(new_new_n8794__), .dout(new_new_n4127__));
  or1   g3186(.dina(new_new_n7095__), .dinb(new_new_n8797__), .dout(new_new_n4128__));
  and1  g3187(.dina(new_new_n1450__), .dinb(new_new_n1319__), .dout(new_new_n4129__));
  or1   g3188(.dina(new_new_n1449__), .dinb(new_new_n1320__), .dout(new_new_n4130__));
  and1  g3189(.dina(new_new_n8798__), .dinb(new_new_n8799__), .dout(new_new_n4131__));
  or1   g3190(.dina(new_new_n8800__), .dinb(new_new_n8801__), .dout(new_new_n4132__));
  and1  g3191(.dina(new_new_n8803__), .dinb(new_new_n8799__), .dout(new_new_n4133__));
  or1   g3192(.dina(new_new_n8805__), .dinb(new_new_n8801__), .dout(new_new_n4134__));
  and1  g3193(.dina(new_new_n8803__), .dinb(new_new_n8798__), .dout(new_new_n4135__));
  or1   g3194(.dina(new_new_n8805__), .dinb(new_new_n8800__), .dout(new_new_n4136__));
  and1  g3195(.dina(new_new_n4136__), .dinb(new_new_n4134__), .dout(new_new_n4137__));
  or1   g3196(.dina(new_new_n4135__), .dinb(new_new_n4133__), .dout(new_new_n4138__));
  and1  g3197(.dina(new_new_n7674__), .dinb(new_new_n8807__), .dout(new_new_n4139__));
  or1   g3198(.dina(new_new_n7689__), .dinb(new_new_n8810__), .dout(new_new_n4140__));
  and1  g3199(.dina(new_new_n8811__), .dinb(new_new_n8812__), .dout(new_new_n4141__));
  or1   g3200(.dina(new_new_n8813__), .dinb(new_new_n8814__), .dout(new_new_n4142__));
  and1  g3201(.dina(new_new_n8816__), .dinb(new_new_n8812__), .dout(new_new_n4143__));
  or1   g3202(.dina(new_new_n8818__), .dinb(new_new_n8814__), .dout(new_new_n4144__));
  and1  g3203(.dina(new_new_n8816__), .dinb(new_new_n8811__), .dout(new_new_n4145__));
  or1   g3204(.dina(new_new_n8818__), .dinb(new_new_n8813__), .dout(new_new_n4146__));
  and1  g3205(.dina(new_new_n4146__), .dinb(new_new_n4144__), .dout(new_new_n4147__));
  or1   g3206(.dina(new_new_n4145__), .dinb(new_new_n4143__), .dout(new_new_n4148__));
  and1  g3207(.dina(new_new_n8819__), .dinb(new_new_n8820__), .dout(new_new_n4149__));
  or1   g3208(.dina(new_new_n8821__), .dinb(new_new_n8822__), .dout(new_new_n4150__));
  and1  g3209(.dina(new_new_n8824__), .dinb(new_new_n8819__), .dout(new_new_n4151__));
  or1   g3210(.dina(new_new_n8826__), .dinb(new_new_n8821__), .dout(new_new_n4152__));
  and1  g3211(.dina(new_new_n8824__), .dinb(new_new_n8820__), .dout(new_new_n4153__));
  or1   g3212(.dina(new_new_n8826__), .dinb(new_new_n8822__), .dout(new_new_n4154__));
  and1  g3213(.dina(new_new_n4154__), .dinb(new_new_n4152__), .dout(new_new_n4155__));
  or1   g3214(.dina(new_new_n4153__), .dinb(new_new_n4151__), .dout(new_new_n4156__));
  and1  g3215(.dina(new_new_n7674__), .dinb(new_new_n8828__), .dout(new_new_n4157__));
  or1   g3216(.dina(new_new_n7689__), .dinb(new_new_n8831__), .dout(new_new_n4158__));
  and1  g3217(.dina(new_new_n8832__), .dinb(new_new_n8833__), .dout(new_new_n4159__));
  or1   g3218(.dina(new_new_n8834__), .dinb(new_new_n8835__), .dout(new_new_n4160__));
  and1  g3219(.dina(new_new_n8837__), .dinb(new_new_n8823__), .dout(new_new_n4161__));
  or1   g3220(.dina(new_new_n8839__), .dinb(new_new_n8825__), .dout(new_new_n4162__));
  and1  g3221(.dina(new_new_n8840__), .dinb(new_new_n8841__), .dout(new_new_n4163__));
  or1   g3222(.dina(new_new_n8842__), .dinb(new_new_n8843__), .dout(new_new_n4164__));
  and1  g3223(.dina(new_new_n8845__), .dinb(new_new_n8841__), .dout(new_new_n4165__));
  or1   g3224(.dina(new_new_n8847__), .dinb(new_new_n8843__), .dout(new_new_n4166__));
  and1  g3225(.dina(new_new_n8845__), .dinb(new_new_n8840__), .dout(new_new_n4167__));
  or1   g3226(.dina(new_new_n8847__), .dinb(new_new_n8842__), .dout(new_new_n4168__));
  and1  g3227(.dina(new_new_n4168__), .dinb(new_new_n4166__), .dout(new_new_n4169__));
  or1   g3228(.dina(new_new_n4167__), .dinb(new_new_n4165__), .dout(new_new_n4170__));
  and1  g3229(.dina(new_new_n8828__), .dinb(new_new_n7903__), .dout(new_new_n4171__));
  or1   g3230(.dina(new_new_n8831__), .dinb(new_new_n7918__), .dout(new_new_n4172__));
  and1  g3231(.dina(new_new_n8848__), .dinb(new_new_n8849__), .dout(new_new_n4173__));
  or1   g3232(.dina(new_new_n8850__), .dinb(new_new_n8851__), .dout(new_new_n4174__));
  and1  g3233(.dina(new_new_n8853__), .dinb(new_new_n8849__), .dout(new_new_n4175__));
  or1   g3234(.dina(new_new_n8855__), .dinb(new_new_n8851__), .dout(new_new_n4176__));
  and1  g3235(.dina(new_new_n8853__), .dinb(new_new_n8848__), .dout(new_new_n4177__));
  or1   g3236(.dina(new_new_n8855__), .dinb(new_new_n8850__), .dout(new_new_n4178__));
  and1  g3237(.dina(new_new_n4178__), .dinb(new_new_n4176__), .dout(new_new_n4179__));
  or1   g3238(.dina(new_new_n4177__), .dinb(new_new_n4175__), .dout(new_new_n4180__));
  and1  g3239(.dina(new_new_n8837__), .dinb(new_new_n8833__), .dout(new_new_n4181__));
  or1   g3240(.dina(new_new_n8839__), .dinb(new_new_n8835__), .dout(new_new_n4182__));
  and1  g3241(.dina(new_new_n8836__), .dinb(new_new_n8832__), .dout(new_new_n4183__));
  or1   g3242(.dina(new_new_n8838__), .dinb(new_new_n8834__), .dout(new_new_n4184__));
  and1  g3243(.dina(new_new_n4184__), .dinb(new_new_n4182__), .dout(new_new_n4185__));
  or1   g3244(.dina(new_new_n4183__), .dinb(new_new_n4181__), .dout(new_new_n4186__));
  and1  g3245(.dina(new_new_n1584__), .dinb(new_new_n1582__), .dout(new_new_n4187__));
  or1   g3246(.dina(new_new_n1583__), .dinb(new_new_n1581__), .dout(new_new_n4188__));
  and1  g3247(.dina(new_new_n7676__), .dinb(new_new_n8857__), .dout(new_new_n4189__));
  or1   g3248(.dina(new_new_n7691__), .dinb(new_new_n8860__), .dout(new_new_n4190__));
  and1  g3249(.dina(new_new_n8862__), .dinb(new_new_n8863__), .dout(new_new_n4191__));
  or1   g3250(.dina(new_new_n8864__), .dinb(new_new_n8865__), .dout(new_new_n4192__));
  and1  g3251(.dina(new_new_n8867__), .dinb(new_new_n1541__), .dout(new_new_n4193__));
  or1   g3252(.dina(new_new_n8869__), .dinb(new_new_n1542__), .dout(new_new_n4194__));
  and1  g3253(.dina(new_new_n8870__), .dinb(new_new_n8871__), .dout(new_new_n4195__));
  or1   g3254(.dina(new_new_n8872__), .dinb(new_new_n8873__), .dout(new_new_n4196__));
  and1  g3255(.dina(new_new_n8875__), .dinb(new_new_n8871__), .dout(new_new_n4197__));
  or1   g3256(.dina(new_new_n8877__), .dinb(new_new_n8873__), .dout(new_new_n4198__));
  and1  g3257(.dina(new_new_n8875__), .dinb(new_new_n8870__), .dout(new_new_n4199__));
  or1   g3258(.dina(new_new_n8877__), .dinb(new_new_n8872__), .dout(new_new_n4200__));
  and1  g3259(.dina(new_new_n4200__), .dinb(new_new_n4198__), .dout(new_new_n4201__));
  or1   g3260(.dina(new_new_n4199__), .dinb(new_new_n4197__), .dout(new_new_n4202__));
  and1  g3261(.dina(new_new_n8857__), .dinb(new_new_n7904__), .dout(new_new_n4203__));
  or1   g3262(.dina(new_new_n8860__), .dinb(new_new_n7919__), .dout(new_new_n4204__));
  and1  g3263(.dina(new_new_n8878__), .dinb(new_new_n8879__), .dout(new_new_n4205__));
  or1   g3264(.dina(new_new_n8880__), .dinb(new_new_n8881__), .dout(new_new_n4206__));
  and1  g3265(.dina(new_new_n8883__), .dinb(new_new_n8874__), .dout(new_new_n4207__));
  or1   g3266(.dina(new_new_n8885__), .dinb(new_new_n8876__), .dout(new_new_n4208__));
  and1  g3267(.dina(new_new_n8886__), .dinb(new_new_n8887__), .dout(new_new_n4209__));
  or1   g3268(.dina(new_new_n8888__), .dinb(new_new_n8889__), .dout(new_new_n4210__));
  and1  g3269(.dina(new_new_n8891__), .dinb(new_new_n8887__), .dout(new_new_n4211__));
  or1   g3270(.dina(new_new_n8893__), .dinb(new_new_n8889__), .dout(new_new_n4212__));
  and1  g3271(.dina(new_new_n8891__), .dinb(new_new_n8886__), .dout(new_new_n4213__));
  or1   g3272(.dina(new_new_n8893__), .dinb(new_new_n8888__), .dout(new_new_n4214__));
  and1  g3273(.dina(new_new_n4214__), .dinb(new_new_n4212__), .dout(new_new_n4215__));
  or1   g3274(.dina(new_new_n4213__), .dinb(new_new_n4211__), .dout(new_new_n4216__));
  and1  g3275(.dina(new_new_n8858__), .dinb(new_new_n8897__), .dout(new_new_n4217__));
  or1   g3276(.dina(new_new_n8861__), .dinb(new_new_n8911__), .dout(new_new_n4218__));
  and1  g3277(.dina(new_new_n8922__), .dinb(new_new_n8923__), .dout(new_new_n4219__));
  or1   g3278(.dina(new_new_n8924__), .dinb(new_new_n8925__), .dout(new_new_n4220__));
  and1  g3279(.dina(new_new_n8927__), .dinb(new_new_n8923__), .dout(new_new_n4221__));
  or1   g3280(.dina(new_new_n8929__), .dinb(new_new_n8925__), .dout(new_new_n4222__));
  and1  g3281(.dina(new_new_n8927__), .dinb(new_new_n8922__), .dout(new_new_n4223__));
  or1   g3282(.dina(new_new_n8929__), .dinb(new_new_n8924__), .dout(new_new_n4224__));
  and1  g3283(.dina(new_new_n4224__), .dinb(new_new_n4222__), .dout(new_new_n4225__));
  or1   g3284(.dina(new_new_n4223__), .dinb(new_new_n4221__), .dout(new_new_n4226__));
  and1  g3285(.dina(new_new_n8883__), .dinb(new_new_n8879__), .dout(new_new_n4227__));
  or1   g3286(.dina(new_new_n8885__), .dinb(new_new_n8881__), .dout(new_new_n4228__));
  and1  g3287(.dina(new_new_n8882__), .dinb(new_new_n8878__), .dout(new_new_n4229__));
  or1   g3288(.dina(new_new_n8884__), .dinb(new_new_n8880__), .dout(new_new_n4230__));
  and1  g3289(.dina(new_new_n4230__), .dinb(new_new_n4228__), .dout(new_new_n4231__));
  or1   g3290(.dina(new_new_n4229__), .dinb(new_new_n4227__), .dout(new_new_n4232__));
  and1  g3291(.dina(new_new_n8867__), .dinb(new_new_n8863__), .dout(new_new_n4233__));
  or1   g3292(.dina(new_new_n8869__), .dinb(new_new_n8865__), .dout(new_new_n4234__));
  and1  g3293(.dina(new_new_n8866__), .dinb(new_new_n8862__), .dout(new_new_n4235__));
  or1   g3294(.dina(new_new_n8868__), .dinb(new_new_n8864__), .dout(new_new_n4236__));
  and1  g3295(.dina(new_new_n4236__), .dinb(new_new_n4234__), .dout(new_new_n4237__));
  or1   g3296(.dina(new_new_n4235__), .dinb(new_new_n4233__), .dout(new_new_n4238__));
  and1  g3297(.dina(new_new_n8931__), .dinb(new_new_n1552__), .dout(new_new_n4239__));
  or1   g3298(.dina(new_new_n8933__), .dinb(new_new_n1551__), .dout(new_new_n4240__));
  and1  g3299(.dina(new_new_n8931__), .dinb(new_new_n1504__), .dout(new_new_n4241__));
  or1   g3300(.dina(new_new_n8933__), .dinb(new_new_n1503__), .dout(new_new_n4242__));
  and1  g3301(.dina(new_new_n4242__), .dinb(new_new_n4240__), .dout(new_new_n4243__));
  or1   g3302(.dina(new_new_n4241__), .dinb(new_new_n4239__), .dout(new_new_n4244__));
  and1  g3303(.dina(new_new_n7676__), .dinb(new_new_n8936__), .dout(new_new_n4245__));
  or1   g3304(.dina(new_new_n7691__), .dinb(new_new_n8939__), .dout(new_new_n4246__));
  and1  g3305(.dina(new_new_n8941__), .dinb(new_new_n8942__), .dout(new_new_n4247__));
  or1   g3306(.dina(new_new_n8943__), .dinb(new_new_n8944__), .dout(new_new_n4248__));
  and1  g3307(.dina(new_new_n8946__), .dinb(new_new_n8930__), .dout(new_new_n4249__));
  or1   g3308(.dina(new_new_n8948__), .dinb(new_new_n8932__), .dout(new_new_n4250__));
  and1  g3309(.dina(new_new_n8949__), .dinb(new_new_n8950__), .dout(new_new_n4251__));
  or1   g3310(.dina(new_new_n8951__), .dinb(new_new_n8952__), .dout(new_new_n4252__));
  and1  g3311(.dina(new_new_n8954__), .dinb(new_new_n8950__), .dout(new_new_n4253__));
  or1   g3312(.dina(new_new_n8956__), .dinb(new_new_n8952__), .dout(new_new_n4254__));
  and1  g3313(.dina(new_new_n8954__), .dinb(new_new_n8949__), .dout(new_new_n4255__));
  or1   g3314(.dina(new_new_n8956__), .dinb(new_new_n8951__), .dout(new_new_n4256__));
  and1  g3315(.dina(new_new_n4256__), .dinb(new_new_n4254__), .dout(new_new_n4257__));
  or1   g3316(.dina(new_new_n4255__), .dinb(new_new_n4253__), .dout(new_new_n4258__));
  and1  g3317(.dina(new_new_n8936__), .dinb(new_new_n7904__), .dout(new_new_n4259__));
  or1   g3318(.dina(new_new_n8939__), .dinb(new_new_n7919__), .dout(new_new_n4260__));
  and1  g3319(.dina(new_new_n8957__), .dinb(new_new_n8958__), .dout(new_new_n4261__));
  or1   g3320(.dina(new_new_n8959__), .dinb(new_new_n8960__), .dout(new_new_n4262__));
  and1  g3321(.dina(new_new_n8962__), .dinb(new_new_n8953__), .dout(new_new_n4263__));
  or1   g3322(.dina(new_new_n8964__), .dinb(new_new_n8955__), .dout(new_new_n4264__));
  and1  g3323(.dina(new_new_n8965__), .dinb(new_new_n8966__), .dout(new_new_n4265__));
  or1   g3324(.dina(new_new_n8967__), .dinb(new_new_n8968__), .dout(new_new_n4266__));
  and1  g3325(.dina(new_new_n8970__), .dinb(new_new_n8966__), .dout(new_new_n4267__));
  or1   g3326(.dina(new_new_n8972__), .dinb(new_new_n8968__), .dout(new_new_n4268__));
  and1  g3327(.dina(new_new_n8970__), .dinb(new_new_n8965__), .dout(new_new_n4269__));
  or1   g3328(.dina(new_new_n8972__), .dinb(new_new_n8967__), .dout(new_new_n4270__));
  and1  g3329(.dina(new_new_n4270__), .dinb(new_new_n4268__), .dout(new_new_n4271__));
  or1   g3330(.dina(new_new_n4269__), .dinb(new_new_n4267__), .dout(new_new_n4272__));
  and1  g3331(.dina(new_new_n8935__), .dinb(new_new_n8897__), .dout(new_new_n4273__));
  or1   g3332(.dina(new_new_n8940__), .dinb(new_new_n8911__), .dout(new_new_n4274__));
  and1  g3333(.dina(new_new_n8973__), .dinb(new_new_n8974__), .dout(new_new_n4275__));
  or1   g3334(.dina(new_new_n8975__), .dinb(new_new_n8976__), .dout(new_new_n4276__));
  and1  g3335(.dina(new_new_n8978__), .dinb(new_new_n8969__), .dout(new_new_n4277__));
  or1   g3336(.dina(new_new_n8980__), .dinb(new_new_n8971__), .dout(new_new_n4278__));
  and1  g3337(.dina(new_new_n8981__), .dinb(new_new_n8982__), .dout(new_new_n4279__));
  or1   g3338(.dina(new_new_n8983__), .dinb(new_new_n8984__), .dout(new_new_n4280__));
  and1  g3339(.dina(new_new_n8986__), .dinb(new_new_n8071__), .dout(new_new_n4281__));
  or1   g3340(.dina(new_new_n8987__), .dinb(new_new_n8073__), .dout(new_new_n4282__));
  and1  g3341(.dina(new_new_n8986__), .dinb(new_new_n8070__), .dout(new_new_n4283__));
  or1   g3342(.dina(new_new_n8987__), .dinb(new_new_n8072__), .dout(new_new_n4284__));
  and1  g3343(.dina(new_new_n4284__), .dinb(new_new_n4282__), .dout(new_new_n4285__));
  or1   g3344(.dina(new_new_n4283__), .dinb(new_new_n4281__), .dout(new_new_n4286__));
  and1  g3345(.dina(new_new_n8043__), .dinb(new_new_n7602__), .dout(new_new_n4287__));
  or1   g3346(.dina(new_new_n8044__), .dinb(new_new_n7615__), .dout(new_new_n4288__));
  or1   g3347(.dina(new_new_n4287__), .dinb(new_new_n4285__), .dout(new_new_n4289__));
  and1  g3348(.dina(new_new_n8989__), .dinb(new_new_n8220__), .dout(new_new_n4290__));
  or1   g3349(.dina(new_new_n8990__), .dinb(new_new_n8222__), .dout(new_new_n4291__));
  and1  g3350(.dina(new_new_n8989__), .dinb(new_new_n8219__), .dout(new_new_n4292__));
  or1   g3351(.dina(new_new_n8990__), .dinb(new_new_n8221__), .dout(new_new_n4293__));
  and1  g3352(.dina(new_new_n4293__), .dinb(new_new_n4291__), .dout(new_new_n4294__));
  or1   g3353(.dina(new_new_n4292__), .dinb(new_new_n4290__), .dout(new_new_n4295__));
  and1  g3354(.dina(new_new_n8192__), .dinb(new_new_n8366__), .dout(new_new_n4296__));
  or1   g3355(.dina(new_new_n8193__), .dinb(new_new_n8375__), .dout(new_new_n4297__));
  or1   g3356(.dina(new_new_n4296__), .dinb(new_new_n4294__), .dout(new_new_n4298__));
  and1  g3357(.dina(new_new_n8992__), .dinb(new_new_n8459__), .dout(new_new_n4299__));
  or1   g3358(.dina(new_new_n8993__), .dinb(new_new_n8461__), .dout(new_new_n4300__));
  and1  g3359(.dina(new_new_n8992__), .dinb(new_new_n8458__), .dout(new_new_n4301__));
  or1   g3360(.dina(new_new_n8993__), .dinb(new_new_n8460__), .dout(new_new_n4302__));
  and1  g3361(.dina(new_new_n4302__), .dinb(new_new_n4300__), .dout(new_new_n4303__));
  or1   g3362(.dina(new_new_n4301__), .dinb(new_new_n4299__), .dout(new_new_n4304__));
  and1  g3363(.dina(new_new_n8397__), .dinb(new_new_n8995__), .dout(new_new_n4305__));
  or1   g3364(.dina(new_new_n8401__), .dinb(new_new_n8998__), .dout(new_new_n4306__));
  or1   g3365(.dina(new_new_n4305__), .dinb(new_new_n4303__), .dout(new_new_n4307__));
  and1  g3366(.dina(new_new_n8789__), .dinb(new_new_n8785__), .dout(new_new_n4308__));
  or1   g3367(.dina(new_new_n8791__), .dinb(new_new_n8787__), .dout(new_new_n4309__));
  and1  g3368(.dina(new_new_n8788__), .dinb(new_new_n8784__), .dout(new_new_n4310__));
  or1   g3369(.dina(new_new_n8790__), .dinb(new_new_n8786__), .dout(new_new_n4311__));
  and1  g3370(.dina(new_new_n4311__), .dinb(new_new_n4309__), .dout(new_new_n4312__));
  or1   g3371(.dina(new_new_n4310__), .dinb(new_new_n4308__), .dout(new_new_n4313__));
  and1  g3372(.dina(new_new_n8773__), .dinb(new_new_n8769__), .dout(new_new_n4314__));
  or1   g3373(.dina(new_new_n8775__), .dinb(new_new_n8771__), .dout(new_new_n4315__));
  and1  g3374(.dina(new_new_n8772__), .dinb(new_new_n8768__), .dout(new_new_n4316__));
  or1   g3375(.dina(new_new_n8774__), .dinb(new_new_n8770__), .dout(new_new_n4317__));
  and1  g3376(.dina(new_new_n4317__), .dinb(new_new_n4315__), .dout(new_new_n4318__));
  or1   g3377(.dina(new_new_n4316__), .dinb(new_new_n4314__), .dout(new_new_n4319__));
  and1  g3378(.dina(new_new_n8566__), .dinb(new_new_n8558__), .dout(new_new_n4320__));
  or1   g3379(.dina(new_new_n8568__), .dinb(new_new_n8560__), .dout(new_new_n4321__));
  and1  g3380(.dina(new_new_n9000__), .dinb(new_new_n9001__), .dout(new_new_n4322__));
  or1   g3381(.dina(new_new_n9002__), .dinb(new_new_n9003__), .dout(new_new_n4323__));
  and1  g3382(.dina(new_new_n9005__), .dinb(new_new_n9001__), .dout(new_new_n4324__));
  or1   g3383(.dina(new_new_n9007__), .dinb(new_new_n9003__), .dout(new_new_n4325__));
  and1  g3384(.dina(new_new_n9005__), .dinb(new_new_n9000__), .dout(new_new_n4326__));
  or1   g3385(.dina(new_new_n9007__), .dinb(new_new_n9002__), .dout(new_new_n4327__));
  and1  g3386(.dina(new_new_n4327__), .dinb(new_new_n4325__), .dout(new_new_n4328__));
  or1   g3387(.dina(new_new_n4326__), .dinb(new_new_n4324__), .dout(new_new_n4329__));
  and1  g3388(.dina(new_new_n6972__), .dinb(new_new_n8366__), .dout(new_new_n4330__));
  or1   g3389(.dina(new_new_n6976__), .dinb(new_new_n8375__), .dout(new_new_n4331__));
  and1  g3390(.dina(new_new_n9008__), .dinb(new_new_n9009__), .dout(new_new_n4332__));
  or1   g3391(.dina(new_new_n9010__), .dinb(new_new_n9011__), .dout(new_new_n4333__));
  and1  g3392(.dina(new_new_n9013__), .dinb(new_new_n9004__), .dout(new_new_n4334__));
  or1   g3393(.dina(new_new_n9015__), .dinb(new_new_n9006__), .dout(new_new_n4335__));
  or1   g3394(.dina(new_new_n4334__), .dinb(new_new_n4312__), .dout(new_new_n4336__));
  or1   g3395(.dina(new_new_n7005__), .dinb(new_new_n8912__), .dout(new_new_n4337__));
  and1  g3396(.dina(new_new_n9019__), .dinb(new_new_n9029__), .dout(new_new_n4338__));
  or1   g3397(.dina(new_new_n9034__), .dinb(new_new_n9043__), .dout(new_new_n4339__));
  and1  g3398(.dina(new_new_n9047__), .dinb(new_new_n9029__), .dout(new_new_n4340__));
  or1   g3399(.dina(new_new_n9061__), .dinb(new_new_n9043__), .dout(new_new_n4341__));
  and1  g3400(.dina(new_new_n9076__), .dinb(new_new_n9030__), .dout(new_new_n4342__));
  or1   g3401(.dina(new_new_n9091__), .dinb(new_new_n9042__), .dout(new_new_n4343__));
  and1  g3402(.dina(new_new_n9047__), .dinb(new_new_n9104__), .dout(new_new_n4344__));
  or1   g3403(.dina(new_new_n9061__), .dinb(new_new_n9107__), .dout(new_new_n4345__));
  and1  g3404(.dina(new_new_n9109__), .dinb(new_new_n9110__), .dout(new_new_n4346__));
  or1   g3405(.dina(new_new_n9111__), .dinb(new_new_n9112__), .dout(new_new_n4347__));
  and1  g3406(.dina(new_new_n9113__), .dinb(new_new_n9110__), .dout(new_new_n4348__));
  or1   g3407(.dina(new_new_n9114__), .dinb(new_new_n9112__), .dout(new_new_n4349__));
  and1  g3408(.dina(new_new_n9116__), .dinb(new_new_n9117__), .dout(new_new_n4350__));
  or1   g3409(.dina(new_new_n9119__), .dinb(new_new_n9120__), .dout(new_new_n4351__));
  and1  g3410(.dina(new_new_n9122__), .dinb(new_new_n9117__), .dout(new_new_n4352__));
  or1   g3411(.dina(new_new_n9124__), .dinb(new_new_n9120__), .dout(new_new_n4353__));
  and1  g3412(.dina(new_new_n9122__), .dinb(new_new_n9116__), .dout(new_new_n4354__));
  or1   g3413(.dina(new_new_n9124__), .dinb(new_new_n9119__), .dout(new_new_n4355__));
  and1  g3414(.dina(new_new_n4355__), .dinb(new_new_n4353__), .dout(new_new_n4356__));
  or1   g3415(.dina(new_new_n4354__), .dinb(new_new_n4352__), .dout(new_new_n4357__));
  and1  g3416(.dina(new_new_n9019__), .dinb(new_new_n9104__), .dout(new_new_n4358__));
  or1   g3417(.dina(new_new_n9034__), .dinb(new_new_n9107__), .dout(new_new_n4359__));
  and1  g3418(.dina(new_new_n9125__), .dinb(new_new_n9126__), .dout(new_new_n4360__));
  or1   g3419(.dina(new_new_n9127__), .dinb(new_new_n9128__), .dout(new_new_n4361__));
  and1  g3420(.dina(new_new_n9130__), .dinb(new_new_n9121__), .dout(new_new_n4362__));
  or1   g3421(.dina(new_new_n9132__), .dinb(new_new_n9123__), .dout(new_new_n4363__));
  and1  g3422(.dina(new_new_n9133__), .dinb(new_new_n9134__), .dout(new_new_n4364__));
  or1   g3423(.dina(new_new_n9135__), .dinb(new_new_n9136__), .dout(new_new_n4365__));
  and1  g3424(.dina(new_new_n7677__), .dinb(new_new_n8794__), .dout(new_new_n4366__));
  or1   g3425(.dina(new_new_n7692__), .dinb(new_new_n8797__), .dout(new_new_n4367__));
  and1  g3426(.dina(new_new_n8815__), .dinb(new_new_n8802__), .dout(new_new_n4368__));
  or1   g3427(.dina(new_new_n8817__), .dinb(new_new_n8804__), .dout(new_new_n4369__));
  and1  g3428(.dina(new_new_n9137__), .dinb(new_new_n9138__), .dout(new_new_n4370__));
  or1   g3429(.dina(new_new_n9139__), .dinb(new_new_n9140__), .dout(new_new_n4371__));
  and1  g3430(.dina(new_new_n9142__), .dinb(new_new_n9138__), .dout(new_new_n4372__));
  or1   g3431(.dina(new_new_n9144__), .dinb(new_new_n9140__), .dout(new_new_n4373__));
  and1  g3432(.dina(new_new_n9142__), .dinb(new_new_n9137__), .dout(new_new_n4374__));
  or1   g3433(.dina(new_new_n9144__), .dinb(new_new_n9139__), .dout(new_new_n4375__));
  and1  g3434(.dina(new_new_n4375__), .dinb(new_new_n4373__), .dout(new_new_n4376__));
  or1   g3435(.dina(new_new_n4374__), .dinb(new_new_n4372__), .dout(new_new_n4377__));
  and1  g3436(.dina(new_new_n8807__), .dinb(new_new_n7906__), .dout(new_new_n4378__));
  or1   g3437(.dina(new_new_n8810__), .dinb(new_new_n7921__), .dout(new_new_n4379__));
  and1  g3438(.dina(new_new_n9145__), .dinb(new_new_n9146__), .dout(new_new_n4380__));
  or1   g3439(.dina(new_new_n9147__), .dinb(new_new_n9148__), .dout(new_new_n4381__));
  and1  g3440(.dina(new_new_n9150__), .dinb(new_new_n9146__), .dout(new_new_n4382__));
  or1   g3441(.dina(new_new_n9152__), .dinb(new_new_n9148__), .dout(new_new_n4383__));
  and1  g3442(.dina(new_new_n9150__), .dinb(new_new_n9145__), .dout(new_new_n4384__));
  or1   g3443(.dina(new_new_n9152__), .dinb(new_new_n9147__), .dout(new_new_n4385__));
  and1  g3444(.dina(new_new_n4385__), .dinb(new_new_n4383__), .dout(new_new_n4386__));
  or1   g3445(.dina(new_new_n4384__), .dinb(new_new_n4382__), .dout(new_new_n4387__));
  and1  g3446(.dina(new_new_n8852__), .dinb(new_new_n8844__), .dout(new_new_n4388__));
  or1   g3447(.dina(new_new_n8854__), .dinb(new_new_n8846__), .dout(new_new_n4389__));
  and1  g3448(.dina(new_new_n9153__), .dinb(new_new_n9154__), .dout(new_new_n4390__));
  or1   g3449(.dina(new_new_n9155__), .dinb(new_new_n9156__), .dout(new_new_n4391__));
  and1  g3450(.dina(new_new_n9158__), .dinb(new_new_n9154__), .dout(new_new_n4392__));
  or1   g3451(.dina(new_new_n9160__), .dinb(new_new_n9156__), .dout(new_new_n4393__));
  and1  g3452(.dina(new_new_n9158__), .dinb(new_new_n9153__), .dout(new_new_n4394__));
  or1   g3453(.dina(new_new_n9160__), .dinb(new_new_n9155__), .dout(new_new_n4395__));
  and1  g3454(.dina(new_new_n4395__), .dinb(new_new_n4393__), .dout(new_new_n4396__));
  or1   g3455(.dina(new_new_n4394__), .dinb(new_new_n4392__), .dout(new_new_n4397__));
  and1  g3456(.dina(new_new_n8829__), .dinb(new_new_n8898__), .dout(new_new_n4398__));
  or1   g3457(.dina(new_new_n8830__), .dinb(new_new_n8912__), .dout(new_new_n4399__));
  and1  g3458(.dina(new_new_n9161__), .dinb(new_new_n9162__), .dout(new_new_n4400__));
  or1   g3459(.dina(new_new_n9163__), .dinb(new_new_n9164__), .dout(new_new_n4401__));
  and1  g3460(.dina(new_new_n9166__), .dinb(new_new_n9162__), .dout(new_new_n4402__));
  or1   g3461(.dina(new_new_n9168__), .dinb(new_new_n9164__), .dout(new_new_n4403__));
  and1  g3462(.dina(new_new_n9166__), .dinb(new_new_n9161__), .dout(new_new_n4404__));
  or1   g3463(.dina(new_new_n9168__), .dinb(new_new_n9163__), .dout(new_new_n4405__));
  and1  g3464(.dina(new_new_n4405__), .dinb(new_new_n4403__), .dout(new_new_n4406__));
  or1   g3465(.dina(new_new_n4404__), .dinb(new_new_n4402__), .dout(new_new_n4407__));
  and1  g3466(.dina(new_new_n8926__), .dinb(new_new_n8890__), .dout(new_new_n4408__));
  or1   g3467(.dina(new_new_n8928__), .dinb(new_new_n8892__), .dout(new_new_n4409__));
  or1   g3468(.dina(new_new_n4408__), .dinb(new_new_n4406__), .dout(new_new_n4410__));
  and1  g3469(.dina(new_new_n1588__), .dinb(new_new_n1580__), .dout(new_new_n4411__));
  or1   g3470(.dina(new_new_n1587__), .dinb(new_new_n1579__), .dout(new_new_n4412__));
  and1  g3471(.dina(new_new_n7087__), .dinb(new_new_n9171__), .dout(new_new_n4413__));
  or1   g3472(.dina(new_new_n7095__), .dinb(new_new_n9177__), .dout(new_new_n4414__));
  and1  g3473(.dina(new_new_n9179__), .dinb(new_new_n9180__), .dout(new_new_n4415__));
  or1   g3474(.dina(new_new_n9181__), .dinb(new_new_n9182__), .dout(new_new_n4416__));
  and1  g3475(.dina(new_new_n9184__), .dinb(new_new_n9180__), .dout(new_new_n4417__));
  or1   g3476(.dina(new_new_n9186__), .dinb(new_new_n9182__), .dout(new_new_n4418__));
  and1  g3477(.dina(new_new_n9184__), .dinb(new_new_n9179__), .dout(new_new_n4419__));
  or1   g3478(.dina(new_new_n9186__), .dinb(new_new_n9181__), .dout(new_new_n4420__));
  and1  g3479(.dina(new_new_n4420__), .dinb(new_new_n4418__), .dout(new_new_n4421__));
  or1   g3480(.dina(new_new_n4419__), .dinb(new_new_n4417__), .dout(new_new_n4422__));
  and1  g3481(.dina(new_new_n9188__), .dinb(new_new_n1556__), .dout(new_new_n4423__));
  or1   g3482(.dina(new_new_n9190__), .dinb(new_new_n1555__), .dout(new_new_n4424__));
  and1  g3483(.dina(new_new_n9188__), .dinb(new_new_n1502__), .dout(new_new_n4425__));
  or1   g3484(.dina(new_new_n9190__), .dinb(new_new_n1501__), .dout(new_new_n4426__));
  and1  g3485(.dina(new_new_n4426__), .dinb(new_new_n4424__), .dout(new_new_n4427__));
  or1   g3486(.dina(new_new_n4425__), .dinb(new_new_n4423__), .dout(new_new_n4428__));
  and1  g3487(.dina(new_new_n7089__), .dinb(new_new_n9193__), .dout(new_new_n4429__));
  or1   g3488(.dina(new_new_n7097__), .dinb(new_new_n9198__), .dout(new_new_n4430__));
  and1  g3489(.dina(new_new_n9200__), .dinb(new_new_n9201__), .dout(new_new_n4431__));
  or1   g3490(.dina(new_new_n9202__), .dinb(new_new_n9203__), .dout(new_new_n4432__));
  and1  g3491(.dina(new_new_n9205__), .dinb(new_new_n9187__), .dout(new_new_n4433__));
  or1   g3492(.dina(new_new_n9207__), .dinb(new_new_n9189__), .dout(new_new_n4434__));
  and1  g3493(.dina(new_new_n9208__), .dinb(new_new_n9209__), .dout(new_new_n4435__));
  or1   g3494(.dina(new_new_n9210__), .dinb(new_new_n9211__), .dout(new_new_n4436__));
  and1  g3495(.dina(new_new_n9213__), .dinb(new_new_n9209__), .dout(new_new_n4437__));
  or1   g3496(.dina(new_new_n9215__), .dinb(new_new_n9211__), .dout(new_new_n4438__));
  and1  g3497(.dina(new_new_n9213__), .dinb(new_new_n9208__), .dout(new_new_n4439__));
  or1   g3498(.dina(new_new_n9215__), .dinb(new_new_n9210__), .dout(new_new_n4440__));
  and1  g3499(.dina(new_new_n4440__), .dinb(new_new_n4438__), .dout(new_new_n4441__));
  or1   g3500(.dina(new_new_n4439__), .dinb(new_new_n4437__), .dout(new_new_n4442__));
  and1  g3501(.dina(new_new_n7677__), .dinb(new_new_n9193__), .dout(new_new_n4443__));
  or1   g3502(.dina(new_new_n7692__), .dinb(new_new_n9198__), .dout(new_new_n4444__));
  and1  g3503(.dina(new_new_n9216__), .dinb(new_new_n9217__), .dout(new_new_n4445__));
  or1   g3504(.dina(new_new_n9218__), .dinb(new_new_n9219__), .dout(new_new_n4446__));
  and1  g3505(.dina(new_new_n9221__), .dinb(new_new_n9217__), .dout(new_new_n4447__));
  or1   g3506(.dina(new_new_n9223__), .dinb(new_new_n9219__), .dout(new_new_n4448__));
  and1  g3507(.dina(new_new_n9221__), .dinb(new_new_n9216__), .dout(new_new_n4449__));
  or1   g3508(.dina(new_new_n9223__), .dinb(new_new_n9218__), .dout(new_new_n4450__));
  and1  g3509(.dina(new_new_n4450__), .dinb(new_new_n4448__), .dout(new_new_n4451__));
  or1   g3510(.dina(new_new_n4449__), .dinb(new_new_n4447__), .dout(new_new_n4452__));
  and1  g3511(.dina(new_new_n9205__), .dinb(new_new_n9201__), .dout(new_new_n4453__));
  or1   g3512(.dina(new_new_n9207__), .dinb(new_new_n9203__), .dout(new_new_n4454__));
  and1  g3513(.dina(new_new_n9204__), .dinb(new_new_n9200__), .dout(new_new_n4455__));
  or1   g3514(.dina(new_new_n9206__), .dinb(new_new_n9202__), .dout(new_new_n4456__));
  and1  g3515(.dina(new_new_n4456__), .dinb(new_new_n4454__), .dout(new_new_n4457__));
  or1   g3516(.dina(new_new_n4455__), .dinb(new_new_n4453__), .dout(new_new_n4458__));
  and1  g3517(.dina(new_new_n9224__), .dinb(new_new_n9225__), .dout(new_new_n4459__));
  or1   g3518(.dina(new_new_n9226__), .dinb(new_new_n9227__), .dout(new_new_n4460__));
  and1  g3519(.dina(new_new_n9229__), .dinb(new_new_n9224__), .dout(new_new_n4461__));
  or1   g3520(.dina(new_new_n9231__), .dinb(new_new_n9226__), .dout(new_new_n4462__));
  and1  g3521(.dina(new_new_n9229__), .dinb(new_new_n9225__), .dout(new_new_n4463__));
  or1   g3522(.dina(new_new_n9231__), .dinb(new_new_n9227__), .dout(new_new_n4464__));
  and1  g3523(.dina(new_new_n4464__), .dinb(new_new_n4462__), .dout(new_new_n4465__));
  or1   g3524(.dina(new_new_n4463__), .dinb(new_new_n4461__), .dout(new_new_n4466__));
  and1  g3525(.dina(new_new_n7089__), .dinb(new_new_n9234__), .dout(new_new_n4467__));
  or1   g3526(.dina(new_new_n7097__), .dinb(new_new_n9239__), .dout(new_new_n4468__));
  and1  g3527(.dina(new_new_n9241__), .dinb(new_new_n9242__), .dout(new_new_n4469__));
  or1   g3528(.dina(new_new_n9243__), .dinb(new_new_n9244__), .dout(new_new_n4470__));
  and1  g3529(.dina(new_new_n9246__), .dinb(new_new_n9228__), .dout(new_new_n4471__));
  or1   g3530(.dina(new_new_n9248__), .dinb(new_new_n9230__), .dout(new_new_n4472__));
  and1  g3531(.dina(new_new_n9249__), .dinb(new_new_n9250__), .dout(new_new_n4473__));
  or1   g3532(.dina(new_new_n9251__), .dinb(new_new_n9252__), .dout(new_new_n4474__));
  and1  g3533(.dina(new_new_n9254__), .dinb(new_new_n9250__), .dout(new_new_n4475__));
  or1   g3534(.dina(new_new_n9256__), .dinb(new_new_n9252__), .dout(new_new_n4476__));
  and1  g3535(.dina(new_new_n9254__), .dinb(new_new_n9249__), .dout(new_new_n4477__));
  or1   g3536(.dina(new_new_n9256__), .dinb(new_new_n9251__), .dout(new_new_n4478__));
  and1  g3537(.dina(new_new_n4478__), .dinb(new_new_n4476__), .dout(new_new_n4479__));
  or1   g3538(.dina(new_new_n4477__), .dinb(new_new_n4475__), .dout(new_new_n4480__));
  and1  g3539(.dina(new_new_n7680__), .dinb(new_new_n9234__), .dout(new_new_n4481__));
  or1   g3540(.dina(new_new_n7695__), .dinb(new_new_n9239__), .dout(new_new_n4482__));
  and1  g3541(.dina(new_new_n9257__), .dinb(new_new_n9258__), .dout(new_new_n4483__));
  or1   g3542(.dina(new_new_n9259__), .dinb(new_new_n9260__), .dout(new_new_n4484__));
  and1  g3543(.dina(new_new_n9262__), .dinb(new_new_n9253__), .dout(new_new_n4485__));
  or1   g3544(.dina(new_new_n9264__), .dinb(new_new_n9255__), .dout(new_new_n4486__));
  and1  g3545(.dina(new_new_n9265__), .dinb(new_new_n9266__), .dout(new_new_n4487__));
  or1   g3546(.dina(new_new_n9267__), .dinb(new_new_n9268__), .dout(new_new_n4488__));
  and1  g3547(.dina(new_new_n9270__), .dinb(new_new_n9266__), .dout(new_new_n4489__));
  or1   g3548(.dina(new_new_n9272__), .dinb(new_new_n9268__), .dout(new_new_n4490__));
  and1  g3549(.dina(new_new_n9270__), .dinb(new_new_n9265__), .dout(new_new_n4491__));
  or1   g3550(.dina(new_new_n9272__), .dinb(new_new_n9267__), .dout(new_new_n4492__));
  and1  g3551(.dina(new_new_n4492__), .dinb(new_new_n4490__), .dout(new_new_n4493__));
  or1   g3552(.dina(new_new_n4491__), .dinb(new_new_n4489__), .dout(new_new_n4494__));
  and1  g3553(.dina(new_new_n9235__), .dinb(new_new_n7906__), .dout(new_new_n4495__));
  or1   g3554(.dina(new_new_n9238__), .dinb(new_new_n7921__), .dout(new_new_n4496__));
  and1  g3555(.dina(new_new_n9273__), .dinb(new_new_n9274__), .dout(new_new_n4497__));
  or1   g3556(.dina(new_new_n9275__), .dinb(new_new_n9276__), .dout(new_new_n4498__));
  and1  g3557(.dina(new_new_n9278__), .dinb(new_new_n9274__), .dout(new_new_n4499__));
  or1   g3558(.dina(new_new_n9280__), .dinb(new_new_n9276__), .dout(new_new_n4500__));
  and1  g3559(.dina(new_new_n9278__), .dinb(new_new_n9273__), .dout(new_new_n4501__));
  or1   g3560(.dina(new_new_n9280__), .dinb(new_new_n9275__), .dout(new_new_n4502__));
  and1  g3561(.dina(new_new_n4502__), .dinb(new_new_n4500__), .dout(new_new_n4503__));
  or1   g3562(.dina(new_new_n4501__), .dinb(new_new_n4499__), .dout(new_new_n4504__));
  and1  g3563(.dina(new_new_n9262__), .dinb(new_new_n9258__), .dout(new_new_n4505__));
  or1   g3564(.dina(new_new_n9264__), .dinb(new_new_n9260__), .dout(new_new_n4506__));
  and1  g3565(.dina(new_new_n9261__), .dinb(new_new_n9257__), .dout(new_new_n4507__));
  or1   g3566(.dina(new_new_n9263__), .dinb(new_new_n9259__), .dout(new_new_n4508__));
  and1  g3567(.dina(new_new_n4508__), .dinb(new_new_n4506__), .dout(new_new_n4509__));
  or1   g3568(.dina(new_new_n4507__), .dinb(new_new_n4505__), .dout(new_new_n4510__));
  and1  g3569(.dina(new_new_n9246__), .dinb(new_new_n9242__), .dout(new_new_n4511__));
  or1   g3570(.dina(new_new_n9248__), .dinb(new_new_n9244__), .dout(new_new_n4512__));
  and1  g3571(.dina(new_new_n9245__), .dinb(new_new_n9241__), .dout(new_new_n4513__));
  or1   g3572(.dina(new_new_n9247__), .dinb(new_new_n9243__), .dout(new_new_n4514__));
  and1  g3573(.dina(new_new_n4514__), .dinb(new_new_n4512__), .dout(new_new_n4515__));
  or1   g3574(.dina(new_new_n4513__), .dinb(new_new_n4511__), .dout(new_new_n4516__));
  and1  g3575(.dina(new_new_n1590__), .dinb(new_new_n1575__), .dout(new_new_n4517__));
  or1   g3576(.dina(new_new_n1589__), .dinb(new_new_n1576__), .dout(new_new_n4518__));
  and1  g3577(.dina(new_new_n9282__), .dinb(new_new_n1395__), .dout(new_new_n4519__));
  or1   g3578(.dina(new_new_n9284__), .dinb(new_new_n1396__), .dout(new_new_n4520__));
  and1  g3579(.dina(new_new_n9285__), .dinb(new_new_n9286__), .dout(new_new_n4521__));
  or1   g3580(.dina(new_new_n9287__), .dinb(new_new_n9288__), .dout(new_new_n4522__));
  and1  g3581(.dina(new_new_n9290__), .dinb(new_new_n9286__), .dout(new_new_n4523__));
  or1   g3582(.dina(new_new_n9292__), .dinb(new_new_n9288__), .dout(new_new_n4524__));
  and1  g3583(.dina(new_new_n9290__), .dinb(new_new_n9285__), .dout(new_new_n4525__));
  or1   g3584(.dina(new_new_n9292__), .dinb(new_new_n9287__), .dout(new_new_n4526__));
  and1  g3585(.dina(new_new_n4526__), .dinb(new_new_n4524__), .dout(new_new_n4527__));
  or1   g3586(.dina(new_new_n4525__), .dinb(new_new_n4523__), .dout(new_new_n4528__));
  and1  g3587(.dina(new_new_n7090__), .dinb(new_new_n9295__), .dout(new_new_n4529__));
  or1   g3588(.dina(new_new_n7098__), .dinb(new_new_n9300__), .dout(new_new_n4530__));
  and1  g3589(.dina(new_new_n9302__), .dinb(new_new_n9303__), .dout(new_new_n4531__));
  or1   g3590(.dina(new_new_n9304__), .dinb(new_new_n9305__), .dout(new_new_n4532__));
  and1  g3591(.dina(new_new_n9307__), .dinb(new_new_n9289__), .dout(new_new_n4533__));
  or1   g3592(.dina(new_new_n9309__), .dinb(new_new_n9291__), .dout(new_new_n4534__));
  and1  g3593(.dina(new_new_n9310__), .dinb(new_new_n9311__), .dout(new_new_n4535__));
  or1   g3594(.dina(new_new_n9312__), .dinb(new_new_n9313__), .dout(new_new_n4536__));
  and1  g3595(.dina(new_new_n9315__), .dinb(new_new_n9311__), .dout(new_new_n4537__));
  or1   g3596(.dina(new_new_n9317__), .dinb(new_new_n9313__), .dout(new_new_n4538__));
  and1  g3597(.dina(new_new_n9315__), .dinb(new_new_n9310__), .dout(new_new_n4539__));
  or1   g3598(.dina(new_new_n9317__), .dinb(new_new_n9312__), .dout(new_new_n4540__));
  and1  g3599(.dina(new_new_n4540__), .dinb(new_new_n4538__), .dout(new_new_n4541__));
  or1   g3600(.dina(new_new_n4539__), .dinb(new_new_n4537__), .dout(new_new_n4542__));
  and1  g3601(.dina(new_new_n7680__), .dinb(new_new_n9295__), .dout(new_new_n4543__));
  or1   g3602(.dina(new_new_n7695__), .dinb(new_new_n9300__), .dout(new_new_n4544__));
  and1  g3603(.dina(new_new_n9318__), .dinb(new_new_n9319__), .dout(new_new_n4545__));
  or1   g3604(.dina(new_new_n9320__), .dinb(new_new_n9321__), .dout(new_new_n4546__));
  and1  g3605(.dina(new_new_n9323__), .dinb(new_new_n9314__), .dout(new_new_n4547__));
  or1   g3606(.dina(new_new_n9325__), .dinb(new_new_n9316__), .dout(new_new_n4548__));
  and1  g3607(.dina(new_new_n9326__), .dinb(new_new_n9327__), .dout(new_new_n4549__));
  or1   g3608(.dina(new_new_n9328__), .dinb(new_new_n9329__), .dout(new_new_n4550__));
  and1  g3609(.dina(new_new_n9331__), .dinb(new_new_n9327__), .dout(new_new_n4551__));
  or1   g3610(.dina(new_new_n9333__), .dinb(new_new_n9329__), .dout(new_new_n4552__));
  and1  g3611(.dina(new_new_n9331__), .dinb(new_new_n9326__), .dout(new_new_n4553__));
  or1   g3612(.dina(new_new_n9333__), .dinb(new_new_n9328__), .dout(new_new_n4554__));
  and1  g3613(.dina(new_new_n4554__), .dinb(new_new_n4552__), .dout(new_new_n4555__));
  or1   g3614(.dina(new_new_n4553__), .dinb(new_new_n4551__), .dout(new_new_n4556__));
  and1  g3615(.dina(new_new_n9296__), .dinb(new_new_n7907__), .dout(new_new_n4557__));
  or1   g3616(.dina(new_new_n9299__), .dinb(new_new_n7922__), .dout(new_new_n4558__));
  and1  g3617(.dina(new_new_n9334__), .dinb(new_new_n9335__), .dout(new_new_n4559__));
  or1   g3618(.dina(new_new_n9336__), .dinb(new_new_n9337__), .dout(new_new_n4560__));
  and1  g3619(.dina(new_new_n9339__), .dinb(new_new_n9330__), .dout(new_new_n4561__));
  or1   g3620(.dina(new_new_n9341__), .dinb(new_new_n9332__), .dout(new_new_n4562__));
  and1  g3621(.dina(new_new_n9342__), .dinb(new_new_n9343__), .dout(new_new_n4563__));
  or1   g3622(.dina(new_new_n9344__), .dinb(new_new_n9345__), .dout(new_new_n4564__));
  and1  g3623(.dina(new_new_n9347__), .dinb(new_new_n9343__), .dout(new_new_n4565__));
  or1   g3624(.dina(new_new_n9349__), .dinb(new_new_n9345__), .dout(new_new_n4566__));
  and1  g3625(.dina(new_new_n9347__), .dinb(new_new_n9342__), .dout(new_new_n4567__));
  or1   g3626(.dina(new_new_n9349__), .dinb(new_new_n9344__), .dout(new_new_n4568__));
  and1  g3627(.dina(new_new_n4568__), .dinb(new_new_n4566__), .dout(new_new_n4569__));
  or1   g3628(.dina(new_new_n4567__), .dinb(new_new_n4565__), .dout(new_new_n4570__));
  and1  g3629(.dina(new_new_n9296__), .dinb(new_new_n8898__), .dout(new_new_n4571__));
  or1   g3630(.dina(new_new_n9301__), .dinb(new_new_n8914__), .dout(new_new_n4572__));
  and1  g3631(.dina(new_new_n9350__), .dinb(new_new_n9351__), .dout(new_new_n4573__));
  or1   g3632(.dina(new_new_n9352__), .dinb(new_new_n9353__), .dout(new_new_n4574__));
  and1  g3633(.dina(new_new_n9355__), .dinb(new_new_n9351__), .dout(new_new_n4575__));
  or1   g3634(.dina(new_new_n9357__), .dinb(new_new_n9353__), .dout(new_new_n4576__));
  and1  g3635(.dina(new_new_n9355__), .dinb(new_new_n9350__), .dout(new_new_n4577__));
  or1   g3636(.dina(new_new_n9357__), .dinb(new_new_n9352__), .dout(new_new_n4578__));
  and1  g3637(.dina(new_new_n4578__), .dinb(new_new_n4576__), .dout(new_new_n4579__));
  or1   g3638(.dina(new_new_n4577__), .dinb(new_new_n4575__), .dout(new_new_n4580__));
  and1  g3639(.dina(new_new_n9339__), .dinb(new_new_n9335__), .dout(new_new_n4581__));
  or1   g3640(.dina(new_new_n9341__), .dinb(new_new_n9337__), .dout(new_new_n4582__));
  and1  g3641(.dina(new_new_n9338__), .dinb(new_new_n9334__), .dout(new_new_n4583__));
  or1   g3642(.dina(new_new_n9340__), .dinb(new_new_n9336__), .dout(new_new_n4584__));
  and1  g3643(.dina(new_new_n4584__), .dinb(new_new_n4582__), .dout(new_new_n4585__));
  or1   g3644(.dina(new_new_n4583__), .dinb(new_new_n4581__), .dout(new_new_n4586__));
  and1  g3645(.dina(new_new_n9323__), .dinb(new_new_n9319__), .dout(new_new_n4587__));
  or1   g3646(.dina(new_new_n9325__), .dinb(new_new_n9321__), .dout(new_new_n4588__));
  and1  g3647(.dina(new_new_n9322__), .dinb(new_new_n9318__), .dout(new_new_n4589__));
  or1   g3648(.dina(new_new_n9324__), .dinb(new_new_n9320__), .dout(new_new_n4590__));
  and1  g3649(.dina(new_new_n4590__), .dinb(new_new_n4588__), .dout(new_new_n4591__));
  or1   g3650(.dina(new_new_n4589__), .dinb(new_new_n4587__), .dout(new_new_n4592__));
  and1  g3651(.dina(new_new_n9307__), .dinb(new_new_n9303__), .dout(new_new_n4593__));
  or1   g3652(.dina(new_new_n9309__), .dinb(new_new_n9305__), .dout(new_new_n4594__));
  and1  g3653(.dina(new_new_n9306__), .dinb(new_new_n9302__), .dout(new_new_n4595__));
  or1   g3654(.dina(new_new_n9308__), .dinb(new_new_n9304__), .dout(new_new_n4596__));
  and1  g3655(.dina(new_new_n4596__), .dinb(new_new_n4594__), .dout(new_new_n4597__));
  or1   g3656(.dina(new_new_n4595__), .dinb(new_new_n4593__), .dout(new_new_n4598__));
  and1  g3657(.dina(new_new_n9282__), .dinb(new_new_n1557__), .dout(new_new_n4599__));
  or1   g3658(.dina(new_new_n9284__), .dinb(new_new_n1558__), .dout(new_new_n4600__));
  and1  g3659(.dina(new_new_n9281__), .dinb(new_new_n1492__), .dout(new_new_n4601__));
  or1   g3660(.dina(new_new_n9283__), .dinb(new_new_n1491__), .dout(new_new_n4602__));
  and1  g3661(.dina(new_new_n4602__), .dinb(new_new_n4600__), .dout(new_new_n4603__));
  or1   g3662(.dina(new_new_n4601__), .dinb(new_new_n4599__), .dout(new_new_n4604__));
  and1  g3663(.dina(new_new_n8466__), .dinb(new_new_n1467__), .dout(new_new_n4605__));
  or1   g3664(.dina(new_new_n8468__), .dinb(new_new_n1468__), .dout(new_new_n4606__));
  and1  g3665(.dina(new_new_n9358__), .dinb(new_new_n9359__), .dout(new_new_n4607__));
  or1   g3666(.dina(new_new_n9360__), .dinb(new_new_n9361__), .dout(new_new_n4608__));
  and1  g3667(.dina(new_new_n9363__), .dinb(new_new_n9359__), .dout(new_new_n4609__));
  or1   g3668(.dina(new_new_n9365__), .dinb(new_new_n9361__), .dout(new_new_n4610__));
  and1  g3669(.dina(new_new_n9363__), .dinb(new_new_n9358__), .dout(new_new_n4611__));
  or1   g3670(.dina(new_new_n9365__), .dinb(new_new_n9360__), .dout(new_new_n4612__));
  and1  g3671(.dina(new_new_n4612__), .dinb(new_new_n4610__), .dout(new_new_n4613__));
  or1   g3672(.dina(new_new_n4611__), .dinb(new_new_n4609__), .dout(new_new_n4614__));
  and1  g3673(.dina(new_new_n7090__), .dinb(new_new_n9368__), .dout(new_new_n4615__));
  or1   g3674(.dina(new_new_n7098__), .dinb(new_new_n9372__), .dout(new_new_n4616__));
  and1  g3675(.dina(new_new_n9374__), .dinb(new_new_n9375__), .dout(new_new_n4617__));
  or1   g3676(.dina(new_new_n9376__), .dinb(new_new_n9377__), .dout(new_new_n4618__));
  and1  g3677(.dina(new_new_n9379__), .dinb(new_new_n9362__), .dout(new_new_n4619__));
  or1   g3678(.dina(new_new_n9381__), .dinb(new_new_n9364__), .dout(new_new_n4620__));
  and1  g3679(.dina(new_new_n9382__), .dinb(new_new_n9383__), .dout(new_new_n4621__));
  or1   g3680(.dina(new_new_n9384__), .dinb(new_new_n9385__), .dout(new_new_n4622__));
  and1  g3681(.dina(new_new_n9387__), .dinb(new_new_n9383__), .dout(new_new_n4623__));
  or1   g3682(.dina(new_new_n9389__), .dinb(new_new_n9385__), .dout(new_new_n4624__));
  and1  g3683(.dina(new_new_n9387__), .dinb(new_new_n9382__), .dout(new_new_n4625__));
  or1   g3684(.dina(new_new_n9389__), .dinb(new_new_n9384__), .dout(new_new_n4626__));
  and1  g3685(.dina(new_new_n4626__), .dinb(new_new_n4624__), .dout(new_new_n4627__));
  or1   g3686(.dina(new_new_n4625__), .dinb(new_new_n4623__), .dout(new_new_n4628__));
  and1  g3687(.dina(new_new_n7681__), .dinb(new_new_n9368__), .dout(new_new_n4629__));
  or1   g3688(.dina(new_new_n7696__), .dinb(new_new_n9372__), .dout(new_new_n4630__));
  and1  g3689(.dina(new_new_n9390__), .dinb(new_new_n9391__), .dout(new_new_n4631__));
  or1   g3690(.dina(new_new_n9392__), .dinb(new_new_n9393__), .dout(new_new_n4632__));
  and1  g3691(.dina(new_new_n9395__), .dinb(new_new_n9386__), .dout(new_new_n4633__));
  or1   g3692(.dina(new_new_n9397__), .dinb(new_new_n9388__), .dout(new_new_n4634__));
  and1  g3693(.dina(new_new_n9398__), .dinb(new_new_n9399__), .dout(new_new_n4635__));
  or1   g3694(.dina(new_new_n9400__), .dinb(new_new_n9401__), .dout(new_new_n4636__));
  and1  g3695(.dina(new_new_n9403__), .dinb(new_new_n9399__), .dout(new_new_n4637__));
  or1   g3696(.dina(new_new_n9405__), .dinb(new_new_n9401__), .dout(new_new_n4638__));
  and1  g3697(.dina(new_new_n9403__), .dinb(new_new_n9398__), .dout(new_new_n4639__));
  or1   g3698(.dina(new_new_n9405__), .dinb(new_new_n9400__), .dout(new_new_n4640__));
  and1  g3699(.dina(new_new_n4640__), .dinb(new_new_n4638__), .dout(new_new_n4641__));
  or1   g3700(.dina(new_new_n4639__), .dinb(new_new_n4637__), .dout(new_new_n4642__));
  and1  g3701(.dina(new_new_n9367__), .dinb(new_new_n7907__), .dout(new_new_n4643__));
  or1   g3702(.dina(new_new_n9371__), .dinb(new_new_n7922__), .dout(new_new_n4644__));
  and1  g3703(.dina(new_new_n9406__), .dinb(new_new_n9407__), .dout(new_new_n4645__));
  or1   g3704(.dina(new_new_n9408__), .dinb(new_new_n9409__), .dout(new_new_n4646__));
  and1  g3705(.dina(new_new_n9411__), .dinb(new_new_n9402__), .dout(new_new_n4647__));
  or1   g3706(.dina(new_new_n9413__), .dinb(new_new_n9404__), .dout(new_new_n4648__));
  and1  g3707(.dina(new_new_n9414__), .dinb(new_new_n9415__), .dout(new_new_n4649__));
  or1   g3708(.dina(new_new_n9416__), .dinb(new_new_n9417__), .dout(new_new_n4650__));
  and1  g3709(.dina(new_new_n9419__), .dinb(new_new_n9415__), .dout(new_new_n4651__));
  or1   g3710(.dina(new_new_n9421__), .dinb(new_new_n9417__), .dout(new_new_n4652__));
  and1  g3711(.dina(new_new_n9419__), .dinb(new_new_n9414__), .dout(new_new_n4653__));
  or1   g3712(.dina(new_new_n9421__), .dinb(new_new_n9416__), .dout(new_new_n4654__));
  and1  g3713(.dina(new_new_n4654__), .dinb(new_new_n4652__), .dout(new_new_n4655__));
  or1   g3714(.dina(new_new_n4653__), .dinb(new_new_n4651__), .dout(new_new_n4656__));
  and1  g3715(.dina(new_new_n9369__), .dinb(new_new_n8900__), .dout(new_new_n4657__));
  or1   g3716(.dina(new_new_n9373__), .dinb(new_new_n8914__), .dout(new_new_n4658__));
  and1  g3717(.dina(new_new_n9422__), .dinb(new_new_n9423__), .dout(new_new_n4659__));
  or1   g3718(.dina(new_new_n9424__), .dinb(new_new_n9425__), .dout(new_new_n4660__));
  and1  g3719(.dina(new_new_n9427__), .dinb(new_new_n9418__), .dout(new_new_n4661__));
  or1   g3720(.dina(new_new_n9429__), .dinb(new_new_n9420__), .dout(new_new_n4662__));
  or1   g3721(.dina(new_new_n4661__), .dinb(new_new_n4579__), .dout(new_new_n4663__));
  and1  g3722(.dina(new_new_n8962__), .dinb(new_new_n8958__), .dout(new_new_n4664__));
  or1   g3723(.dina(new_new_n8964__), .dinb(new_new_n8960__), .dout(new_new_n4665__));
  and1  g3724(.dina(new_new_n8961__), .dinb(new_new_n8957__), .dout(new_new_n4666__));
  or1   g3725(.dina(new_new_n8963__), .dinb(new_new_n8959__), .dout(new_new_n4667__));
  and1  g3726(.dina(new_new_n4667__), .dinb(new_new_n4665__), .dout(new_new_n4668__));
  or1   g3727(.dina(new_new_n4666__), .dinb(new_new_n4664__), .dout(new_new_n4669__));
  and1  g3728(.dina(new_new_n8946__), .dinb(new_new_n8942__), .dout(new_new_n4670__));
  or1   g3729(.dina(new_new_n8948__), .dinb(new_new_n8944__), .dout(new_new_n4671__));
  and1  g3730(.dina(new_new_n8945__), .dinb(new_new_n8941__), .dout(new_new_n4672__));
  or1   g3731(.dina(new_new_n8947__), .dinb(new_new_n8943__), .dout(new_new_n4673__));
  and1  g3732(.dina(new_new_n4673__), .dinb(new_new_n4671__), .dout(new_new_n4674__));
  or1   g3733(.dina(new_new_n4672__), .dinb(new_new_n4670__), .dout(new_new_n4675__));
  and1  g3734(.dina(new_new_n9430__), .dinb(new_new_n9431__), .dout(new_new_n4676__));
  or1   g3735(.dina(new_new_n9432__), .dinb(new_new_n9433__), .dout(new_new_n4677__));
  and1  g3736(.dina(new_new_n9435__), .dinb(new_new_n9430__), .dout(new_new_n4678__));
  or1   g3737(.dina(new_new_n9437__), .dinb(new_new_n9432__), .dout(new_new_n4679__));
  and1  g3738(.dina(new_new_n9435__), .dinb(new_new_n9431__), .dout(new_new_n4680__));
  or1   g3739(.dina(new_new_n9437__), .dinb(new_new_n9433__), .dout(new_new_n4681__));
  and1  g3740(.dina(new_new_n4681__), .dinb(new_new_n4679__), .dout(new_new_n4682__));
  or1   g3741(.dina(new_new_n4680__), .dinb(new_new_n4678__), .dout(new_new_n4683__));
  and1  g3742(.dina(new_new_n7681__), .dinb(new_new_n9440__), .dout(new_new_n4684__));
  or1   g3743(.dina(new_new_n7696__), .dinb(new_new_n9443__), .dout(new_new_n4685__));
  and1  g3744(.dina(new_new_n9445__), .dinb(new_new_n9446__), .dout(new_new_n4686__));
  or1   g3745(.dina(new_new_n9447__), .dinb(new_new_n9448__), .dout(new_new_n4687__));
  and1  g3746(.dina(new_new_n9450__), .dinb(new_new_n9434__), .dout(new_new_n4688__));
  or1   g3747(.dina(new_new_n9452__), .dinb(new_new_n9436__), .dout(new_new_n4689__));
  and1  g3748(.dina(new_new_n9453__), .dinb(new_new_n9454__), .dout(new_new_n4690__));
  or1   g3749(.dina(new_new_n9455__), .dinb(new_new_n9456__), .dout(new_new_n4691__));
  and1  g3750(.dina(new_new_n9458__), .dinb(new_new_n9454__), .dout(new_new_n4692__));
  or1   g3751(.dina(new_new_n9460__), .dinb(new_new_n9456__), .dout(new_new_n4693__));
  and1  g3752(.dina(new_new_n9458__), .dinb(new_new_n9453__), .dout(new_new_n4694__));
  or1   g3753(.dina(new_new_n9460__), .dinb(new_new_n9455__), .dout(new_new_n4695__));
  and1  g3754(.dina(new_new_n4695__), .dinb(new_new_n4693__), .dout(new_new_n4696__));
  or1   g3755(.dina(new_new_n4694__), .dinb(new_new_n4692__), .dout(new_new_n4697__));
  and1  g3756(.dina(new_new_n9440__), .dinb(new_new_n7910__), .dout(new_new_n4698__));
  or1   g3757(.dina(new_new_n9443__), .dinb(new_new_n7925__), .dout(new_new_n4699__));
  and1  g3758(.dina(new_new_n9461__), .dinb(new_new_n9462__), .dout(new_new_n4700__));
  or1   g3759(.dina(new_new_n9463__), .dinb(new_new_n9464__), .dout(new_new_n4701__));
  and1  g3760(.dina(new_new_n9466__), .dinb(new_new_n9457__), .dout(new_new_n4702__));
  or1   g3761(.dina(new_new_n9468__), .dinb(new_new_n9459__), .dout(new_new_n4703__));
  and1  g3762(.dina(new_new_n9469__), .dinb(new_new_n9470__), .dout(new_new_n4704__));
  or1   g3763(.dina(new_new_n9471__), .dinb(new_new_n9472__), .dout(new_new_n4705__));
  and1  g3764(.dina(new_new_n9474__), .dinb(new_new_n9470__), .dout(new_new_n4706__));
  or1   g3765(.dina(new_new_n9476__), .dinb(new_new_n9472__), .dout(new_new_n4707__));
  and1  g3766(.dina(new_new_n9474__), .dinb(new_new_n9469__), .dout(new_new_n4708__));
  or1   g3767(.dina(new_new_n9476__), .dinb(new_new_n9471__), .dout(new_new_n4709__));
  and1  g3768(.dina(new_new_n4709__), .dinb(new_new_n4707__), .dout(new_new_n4710__));
  or1   g3769(.dina(new_new_n4708__), .dinb(new_new_n4706__), .dout(new_new_n4711__));
  and1  g3770(.dina(new_new_n9439__), .dinb(new_new_n8900__), .dout(new_new_n4712__));
  or1   g3771(.dina(new_new_n9444__), .dinb(new_new_n8915__), .dout(new_new_n4713__));
  and1  g3772(.dina(new_new_n9477__), .dinb(new_new_n9478__), .dout(new_new_n4714__));
  or1   g3773(.dina(new_new_n9479__), .dinb(new_new_n9480__), .dout(new_new_n4715__));
  and1  g3774(.dina(new_new_n9482__), .dinb(new_new_n9478__), .dout(new_new_n4716__));
  or1   g3775(.dina(new_new_n9484__), .dinb(new_new_n9480__), .dout(new_new_n4717__));
  and1  g3776(.dina(new_new_n9482__), .dinb(new_new_n9477__), .dout(new_new_n4718__));
  or1   g3777(.dina(new_new_n9484__), .dinb(new_new_n9479__), .dout(new_new_n4719__));
  and1  g3778(.dina(new_new_n4719__), .dinb(new_new_n4717__), .dout(new_new_n4720__));
  or1   g3779(.dina(new_new_n4718__), .dinb(new_new_n4716__), .dout(new_new_n4721__));
  and1  g3780(.dina(new_new_n9466__), .dinb(new_new_n9462__), .dout(new_new_n4722__));
  or1   g3781(.dina(new_new_n9468__), .dinb(new_new_n9464__), .dout(new_new_n4723__));
  and1  g3782(.dina(new_new_n9465__), .dinb(new_new_n9461__), .dout(new_new_n4724__));
  or1   g3783(.dina(new_new_n9467__), .dinb(new_new_n9463__), .dout(new_new_n4725__));
  and1  g3784(.dina(new_new_n4725__), .dinb(new_new_n4723__), .dout(new_new_n4726__));
  or1   g3785(.dina(new_new_n4724__), .dinb(new_new_n4722__), .dout(new_new_n4727__));
  and1  g3786(.dina(new_new_n9450__), .dinb(new_new_n9446__), .dout(new_new_n4728__));
  or1   g3787(.dina(new_new_n9452__), .dinb(new_new_n9448__), .dout(new_new_n4729__));
  and1  g3788(.dina(new_new_n9449__), .dinb(new_new_n9445__), .dout(new_new_n4730__));
  or1   g3789(.dina(new_new_n9451__), .dinb(new_new_n9447__), .dout(new_new_n4731__));
  and1  g3790(.dina(new_new_n4731__), .dinb(new_new_n4729__), .dout(new_new_n4732__));
  or1   g3791(.dina(new_new_n4730__), .dinb(new_new_n4728__), .dout(new_new_n4733__));
  and1  g3792(.dina(new_new_n1592__), .dinb(new_new_n1573__), .dout(new_new_n4734__));
  or1   g3793(.dina(new_new_n1591__), .dinb(new_new_n1574__), .dout(new_new_n4735__));
  and1  g3794(.dina(new_new_n9486__), .dinb(new_new_n1397__), .dout(new_new_n4736__));
  or1   g3795(.dina(new_new_n9488__), .dinb(new_new_n1398__), .dout(new_new_n4737__));
  and1  g3796(.dina(new_new_n9489__), .dinb(new_new_n9490__), .dout(new_new_n4738__));
  or1   g3797(.dina(new_new_n9491__), .dinb(new_new_n9492__), .dout(new_new_n4739__));
  and1  g3798(.dina(new_new_n9494__), .dinb(new_new_n9490__), .dout(new_new_n4740__));
  or1   g3799(.dina(new_new_n9496__), .dinb(new_new_n9492__), .dout(new_new_n4741__));
  and1  g3800(.dina(new_new_n9494__), .dinb(new_new_n9489__), .dout(new_new_n4742__));
  or1   g3801(.dina(new_new_n9496__), .dinb(new_new_n9491__), .dout(new_new_n4743__));
  and1  g3802(.dina(new_new_n4743__), .dinb(new_new_n4741__), .dout(new_new_n4744__));
  or1   g3803(.dina(new_new_n4742__), .dinb(new_new_n4740__), .dout(new_new_n4745__));
  and1  g3804(.dina(new_new_n7683__), .dinb(new_new_n9499__), .dout(new_new_n4746__));
  or1   g3805(.dina(new_new_n7698__), .dinb(new_new_n9502__), .dout(new_new_n4747__));
  and1  g3806(.dina(new_new_n9504__), .dinb(new_new_n9505__), .dout(new_new_n4748__));
  or1   g3807(.dina(new_new_n9506__), .dinb(new_new_n9507__), .dout(new_new_n4749__));
  and1  g3808(.dina(new_new_n9509__), .dinb(new_new_n9493__), .dout(new_new_n4750__));
  or1   g3809(.dina(new_new_n9511__), .dinb(new_new_n9495__), .dout(new_new_n4751__));
  and1  g3810(.dina(new_new_n9512__), .dinb(new_new_n9513__), .dout(new_new_n4752__));
  or1   g3811(.dina(new_new_n9514__), .dinb(new_new_n9515__), .dout(new_new_n4753__));
  and1  g3812(.dina(new_new_n9517__), .dinb(new_new_n9513__), .dout(new_new_n4754__));
  or1   g3813(.dina(new_new_n9519__), .dinb(new_new_n9515__), .dout(new_new_n4755__));
  and1  g3814(.dina(new_new_n9517__), .dinb(new_new_n9512__), .dout(new_new_n4756__));
  or1   g3815(.dina(new_new_n9519__), .dinb(new_new_n9514__), .dout(new_new_n4757__));
  and1  g3816(.dina(new_new_n4757__), .dinb(new_new_n4755__), .dout(new_new_n4758__));
  or1   g3817(.dina(new_new_n4756__), .dinb(new_new_n4754__), .dout(new_new_n4759__));
  and1  g3818(.dina(new_new_n9499__), .dinb(new_new_n7910__), .dout(new_new_n4760__));
  or1   g3819(.dina(new_new_n9502__), .dinb(new_new_n7925__), .dout(new_new_n4761__));
  and1  g3820(.dina(new_new_n9520__), .dinb(new_new_n9521__), .dout(new_new_n4762__));
  or1   g3821(.dina(new_new_n9522__), .dinb(new_new_n9523__), .dout(new_new_n4763__));
  and1  g3822(.dina(new_new_n9525__), .dinb(new_new_n9516__), .dout(new_new_n4764__));
  or1   g3823(.dina(new_new_n9527__), .dinb(new_new_n9518__), .dout(new_new_n4765__));
  and1  g3824(.dina(new_new_n9528__), .dinb(new_new_n9529__), .dout(new_new_n4766__));
  or1   g3825(.dina(new_new_n9530__), .dinb(new_new_n9531__), .dout(new_new_n4767__));
  and1  g3826(.dina(new_new_n9533__), .dinb(new_new_n9529__), .dout(new_new_n4768__));
  or1   g3827(.dina(new_new_n9535__), .dinb(new_new_n9531__), .dout(new_new_n4769__));
  and1  g3828(.dina(new_new_n9533__), .dinb(new_new_n9528__), .dout(new_new_n4770__));
  or1   g3829(.dina(new_new_n9535__), .dinb(new_new_n9530__), .dout(new_new_n4771__));
  and1  g3830(.dina(new_new_n4771__), .dinb(new_new_n4769__), .dout(new_new_n4772__));
  or1   g3831(.dina(new_new_n4770__), .dinb(new_new_n4768__), .dout(new_new_n4773__));
  and1  g3832(.dina(new_new_n9498__), .dinb(new_new_n8901__), .dout(new_new_n4774__));
  or1   g3833(.dina(new_new_n9503__), .dinb(new_new_n8915__), .dout(new_new_n4775__));
  and1  g3834(.dina(new_new_n9536__), .dinb(new_new_n9537__), .dout(new_new_n4776__));
  or1   g3835(.dina(new_new_n9538__), .dinb(new_new_n9539__), .dout(new_new_n4777__));
  and1  g3836(.dina(new_new_n9541__), .dinb(new_new_n9532__), .dout(new_new_n4778__));
  or1   g3837(.dina(new_new_n9543__), .dinb(new_new_n9534__), .dout(new_new_n4779__));
  and1  g3838(.dina(new_new_n9544__), .dinb(new_new_n9545__), .dout(new_new_n4780__));
  or1   g3839(.dina(new_new_n9546__), .dinb(new_new_n9547__), .dout(new_new_n4781__));
  and1  g3840(.dina(new_new_n9549__), .dinb(new_new_n9545__), .dout(new_new_n4782__));
  or1   g3841(.dina(new_new_n9551__), .dinb(new_new_n9547__), .dout(new_new_n4783__));
  and1  g3842(.dina(new_new_n9549__), .dinb(new_new_n9544__), .dout(new_new_n4784__));
  or1   g3843(.dina(new_new_n9551__), .dinb(new_new_n9546__), .dout(new_new_n4785__));
  and1  g3844(.dina(new_new_n4785__), .dinb(new_new_n4783__), .dout(new_new_n4786__));
  or1   g3845(.dina(new_new_n4784__), .dinb(new_new_n4782__), .dout(new_new_n4787__));
  and1  g3846(.dina(new_new_n9500__), .dinb(new_new_n9555__), .dout(new_new_n4788__));
  or1   g3847(.dina(new_new_n9503__), .dinb(new_new_n9564__), .dout(new_new_n4789__));
  and1  g3848(.dina(new_new_n9570__), .dinb(new_new_n9571__), .dout(new_new_n4790__));
  or1   g3849(.dina(new_new_n9572__), .dinb(new_new_n9573__), .dout(new_new_n4791__));
  and1  g3850(.dina(new_new_n9575__), .dinb(new_new_n9571__), .dout(new_new_n4792__));
  or1   g3851(.dina(new_new_n9577__), .dinb(new_new_n9573__), .dout(new_new_n4793__));
  and1  g3852(.dina(new_new_n9575__), .dinb(new_new_n9570__), .dout(new_new_n4794__));
  or1   g3853(.dina(new_new_n9577__), .dinb(new_new_n9572__), .dout(new_new_n4795__));
  and1  g3854(.dina(new_new_n4795__), .dinb(new_new_n4793__), .dout(new_new_n4796__));
  or1   g3855(.dina(new_new_n4794__), .dinb(new_new_n4792__), .dout(new_new_n4797__));
  and1  g3856(.dina(new_new_n9541__), .dinb(new_new_n9537__), .dout(new_new_n4798__));
  or1   g3857(.dina(new_new_n9543__), .dinb(new_new_n9539__), .dout(new_new_n4799__));
  and1  g3858(.dina(new_new_n9540__), .dinb(new_new_n9536__), .dout(new_new_n4800__));
  or1   g3859(.dina(new_new_n9542__), .dinb(new_new_n9538__), .dout(new_new_n4801__));
  and1  g3860(.dina(new_new_n4801__), .dinb(new_new_n4799__), .dout(new_new_n4802__));
  or1   g3861(.dina(new_new_n4800__), .dinb(new_new_n4798__), .dout(new_new_n4803__));
  and1  g3862(.dina(new_new_n9525__), .dinb(new_new_n9521__), .dout(new_new_n4804__));
  or1   g3863(.dina(new_new_n9527__), .dinb(new_new_n9523__), .dout(new_new_n4805__));
  and1  g3864(.dina(new_new_n9524__), .dinb(new_new_n9520__), .dout(new_new_n4806__));
  or1   g3865(.dina(new_new_n9526__), .dinb(new_new_n9522__), .dout(new_new_n4807__));
  and1  g3866(.dina(new_new_n4807__), .dinb(new_new_n4805__), .dout(new_new_n4808__));
  or1   g3867(.dina(new_new_n4806__), .dinb(new_new_n4804__), .dout(new_new_n4809__));
  and1  g3868(.dina(new_new_n9509__), .dinb(new_new_n9505__), .dout(new_new_n4810__));
  or1   g3869(.dina(new_new_n9511__), .dinb(new_new_n9507__), .dout(new_new_n4811__));
  and1  g3870(.dina(new_new_n9508__), .dinb(new_new_n9504__), .dout(new_new_n4812__));
  or1   g3871(.dina(new_new_n9510__), .dinb(new_new_n9506__), .dout(new_new_n4813__));
  and1  g3872(.dina(new_new_n4813__), .dinb(new_new_n4811__), .dout(new_new_n4814__));
  or1   g3873(.dina(new_new_n4812__), .dinb(new_new_n4810__), .dout(new_new_n4815__));
  and1  g3874(.dina(new_new_n9486__), .dinb(new_new_n1559__), .dout(new_new_n4816__));
  or1   g3875(.dina(new_new_n9488__), .dinb(new_new_n1560__), .dout(new_new_n4817__));
  and1  g3876(.dina(new_new_n9485__), .dinb(new_new_n1490__), .dout(new_new_n4818__));
  or1   g3877(.dina(new_new_n9487__), .dinb(new_new_n1489__), .dout(new_new_n4819__));
  and1  g3878(.dina(new_new_n4819__), .dinb(new_new_n4817__), .dout(new_new_n4820__));
  or1   g3879(.dina(new_new_n4818__), .dinb(new_new_n4816__), .dout(new_new_n4821__));
  and1  g3880(.dina(new_new_n9578__), .dinb(new_new_n9579__), .dout(new_new_n4822__));
  or1   g3881(.dina(new_new_n9580__), .dinb(new_new_n9581__), .dout(new_new_n4823__));
  and1  g3882(.dina(new_new_n9583__), .dinb(new_new_n1469__), .dout(new_new_n4824__));
  or1   g3883(.dina(new_new_n9585__), .dinb(new_new_n1470__), .dout(new_new_n4825__));
  and1  g3884(.dina(new_new_n9586__), .dinb(new_new_n9587__), .dout(new_new_n4826__));
  or1   g3885(.dina(new_new_n9588__), .dinb(new_new_n9589__), .dout(new_new_n4827__));
  and1  g3886(.dina(new_new_n9591__), .dinb(new_new_n9587__), .dout(new_new_n4828__));
  or1   g3887(.dina(new_new_n9593__), .dinb(new_new_n9589__), .dout(new_new_n4829__));
  and1  g3888(.dina(new_new_n9591__), .dinb(new_new_n9586__), .dout(new_new_n4830__));
  or1   g3889(.dina(new_new_n9593__), .dinb(new_new_n9588__), .dout(new_new_n4831__));
  and1  g3890(.dina(new_new_n4831__), .dinb(new_new_n4829__), .dout(new_new_n4832__));
  or1   g3891(.dina(new_new_n4830__), .dinb(new_new_n4828__), .dout(new_new_n4833__));
  and1  g3892(.dina(new_new_n7683__), .dinb(new_new_n9596__), .dout(new_new_n4834__));
  or1   g3893(.dina(new_new_n7698__), .dinb(new_new_n9600__), .dout(new_new_n4835__));
  and1  g3894(.dina(new_new_n9602__), .dinb(new_new_n9603__), .dout(new_new_n4836__));
  or1   g3895(.dina(new_new_n9604__), .dinb(new_new_n9605__), .dout(new_new_n4837__));
  and1  g3896(.dina(new_new_n9607__), .dinb(new_new_n9590__), .dout(new_new_n4838__));
  or1   g3897(.dina(new_new_n9609__), .dinb(new_new_n9592__), .dout(new_new_n4839__));
  and1  g3898(.dina(new_new_n9610__), .dinb(new_new_n9611__), .dout(new_new_n4840__));
  or1   g3899(.dina(new_new_n9612__), .dinb(new_new_n9613__), .dout(new_new_n4841__));
  and1  g3900(.dina(new_new_n9615__), .dinb(new_new_n9611__), .dout(new_new_n4842__));
  or1   g3901(.dina(new_new_n9617__), .dinb(new_new_n9613__), .dout(new_new_n4843__));
  and1  g3902(.dina(new_new_n9615__), .dinb(new_new_n9610__), .dout(new_new_n4844__));
  or1   g3903(.dina(new_new_n9617__), .dinb(new_new_n9612__), .dout(new_new_n4845__));
  and1  g3904(.dina(new_new_n4845__), .dinb(new_new_n4843__), .dout(new_new_n4846__));
  or1   g3905(.dina(new_new_n4844__), .dinb(new_new_n4842__), .dout(new_new_n4847__));
  and1  g3906(.dina(new_new_n9596__), .dinb(new_new_n7911__), .dout(new_new_n4848__));
  or1   g3907(.dina(new_new_n9600__), .dinb(new_new_n7926__), .dout(new_new_n4849__));
  and1  g3908(.dina(new_new_n9618__), .dinb(new_new_n9619__), .dout(new_new_n4850__));
  or1   g3909(.dina(new_new_n9620__), .dinb(new_new_n9621__), .dout(new_new_n4851__));
  and1  g3910(.dina(new_new_n9623__), .dinb(new_new_n9614__), .dout(new_new_n4852__));
  or1   g3911(.dina(new_new_n9625__), .dinb(new_new_n9616__), .dout(new_new_n4853__));
  and1  g3912(.dina(new_new_n9626__), .dinb(new_new_n9627__), .dout(new_new_n4854__));
  or1   g3913(.dina(new_new_n9628__), .dinb(new_new_n9629__), .dout(new_new_n4855__));
  and1  g3914(.dina(new_new_n9631__), .dinb(new_new_n9627__), .dout(new_new_n4856__));
  or1   g3915(.dina(new_new_n9633__), .dinb(new_new_n9629__), .dout(new_new_n4857__));
  and1  g3916(.dina(new_new_n9631__), .dinb(new_new_n9626__), .dout(new_new_n4858__));
  or1   g3917(.dina(new_new_n9633__), .dinb(new_new_n9628__), .dout(new_new_n4859__));
  and1  g3918(.dina(new_new_n4859__), .dinb(new_new_n4857__), .dout(new_new_n4860__));
  or1   g3919(.dina(new_new_n4858__), .dinb(new_new_n4856__), .dout(new_new_n4861__));
  and1  g3920(.dina(new_new_n9595__), .dinb(new_new_n8901__), .dout(new_new_n4862__));
  or1   g3921(.dina(new_new_n9599__), .dinb(new_new_n8918__), .dout(new_new_n4863__));
  and1  g3922(.dina(new_new_n9634__), .dinb(new_new_n9635__), .dout(new_new_n4864__));
  or1   g3923(.dina(new_new_n9636__), .dinb(new_new_n9637__), .dout(new_new_n4865__));
  and1  g3924(.dina(new_new_n9639__), .dinb(new_new_n9630__), .dout(new_new_n4866__));
  or1   g3925(.dina(new_new_n9641__), .dinb(new_new_n9632__), .dout(new_new_n4867__));
  and1  g3926(.dina(new_new_n9642__), .dinb(new_new_n9643__), .dout(new_new_n4868__));
  or1   g3927(.dina(new_new_n9644__), .dinb(new_new_n9645__), .dout(new_new_n4869__));
  and1  g3928(.dina(new_new_n9647__), .dinb(new_new_n9643__), .dout(new_new_n4870__));
  or1   g3929(.dina(new_new_n9649__), .dinb(new_new_n9645__), .dout(new_new_n4871__));
  and1  g3930(.dina(new_new_n9647__), .dinb(new_new_n9642__), .dout(new_new_n4872__));
  or1   g3931(.dina(new_new_n9649__), .dinb(new_new_n9644__), .dout(new_new_n4873__));
  and1  g3932(.dina(new_new_n4873__), .dinb(new_new_n4871__), .dout(new_new_n4874__));
  or1   g3933(.dina(new_new_n4872__), .dinb(new_new_n4870__), .dout(new_new_n4875__));
  and1  g3934(.dina(new_new_n9597__), .dinb(new_new_n9555__), .dout(new_new_n4876__));
  or1   g3935(.dina(new_new_n9601__), .dinb(new_new_n9564__), .dout(new_new_n4877__));
  and1  g3936(.dina(new_new_n9650__), .dinb(new_new_n9651__), .dout(new_new_n4878__));
  or1   g3937(.dina(new_new_n9652__), .dinb(new_new_n9653__), .dout(new_new_n4879__));
  and1  g3938(.dina(new_new_n9655__), .dinb(new_new_n9646__), .dout(new_new_n4880__));
  or1   g3939(.dina(new_new_n9657__), .dinb(new_new_n9648__), .dout(new_new_n4881__));
  or1   g3940(.dina(new_new_n4880__), .dinb(new_new_n4796__), .dout(new_new_n4882__));
  and1  g3941(.dina(new_new_n9379__), .dinb(new_new_n9375__), .dout(new_new_n4883__));
  or1   g3942(.dina(new_new_n9381__), .dinb(new_new_n9377__), .dout(new_new_n4884__));
  and1  g3943(.dina(new_new_n9378__), .dinb(new_new_n9374__), .dout(new_new_n4885__));
  or1   g3944(.dina(new_new_n9380__), .dinb(new_new_n9376__), .dout(new_new_n4886__));
  and1  g3945(.dina(new_new_n4886__), .dinb(new_new_n4884__), .dout(new_new_n4887__));
  or1   g3946(.dina(new_new_n4885__), .dinb(new_new_n4883__), .dout(new_new_n4888__));
  and1  g3947(.dina(new_new_n8482__), .dinb(new_new_n8474__), .dout(new_new_n4889__));
  or1   g3948(.dina(new_new_n8484__), .dinb(new_new_n8476__), .dout(new_new_n4890__));
  and1  g3949(.dina(new_new_n9658__), .dinb(new_new_n9659__), .dout(new_new_n4891__));
  or1   g3950(.dina(new_new_n9660__), .dinb(new_new_n9661__), .dout(new_new_n4892__));
  and1  g3951(.dina(new_new_n9663__), .dinb(new_new_n9659__), .dout(new_new_n4893__));
  or1   g3952(.dina(new_new_n9665__), .dinb(new_new_n9661__), .dout(new_new_n4894__));
  and1  g3953(.dina(new_new_n9663__), .dinb(new_new_n9658__), .dout(new_new_n4895__));
  or1   g3954(.dina(new_new_n9665__), .dinb(new_new_n9660__), .dout(new_new_n4896__));
  and1  g3955(.dina(new_new_n4896__), .dinb(new_new_n4894__), .dout(new_new_n4897__));
  or1   g3956(.dina(new_new_n4895__), .dinb(new_new_n4893__), .dout(new_new_n4898__));
  and1  g3957(.dina(new_new_n7684__), .dinb(new_new_n7705__), .dout(new_new_n4899__));
  or1   g3958(.dina(new_new_n7699__), .dinb(new_new_n7709__), .dout(new_new_n4900__));
  and1  g3959(.dina(new_new_n9666__), .dinb(new_new_n9667__), .dout(new_new_n4901__));
  or1   g3960(.dina(new_new_n9668__), .dinb(new_new_n9669__), .dout(new_new_n4902__));
  and1  g3961(.dina(new_new_n9671__), .dinb(new_new_n9667__), .dout(new_new_n4903__));
  or1   g3962(.dina(new_new_n9673__), .dinb(new_new_n9669__), .dout(new_new_n4904__));
  and1  g3963(.dina(new_new_n9671__), .dinb(new_new_n9666__), .dout(new_new_n4905__));
  or1   g3964(.dina(new_new_n9673__), .dinb(new_new_n9668__), .dout(new_new_n4906__));
  and1  g3965(.dina(new_new_n4906__), .dinb(new_new_n4904__), .dout(new_new_n4907__));
  or1   g3966(.dina(new_new_n4905__), .dinb(new_new_n4903__), .dout(new_new_n4908__));
  and1  g3967(.dina(new_new_n8498__), .dinb(new_new_n8490__), .dout(new_new_n4909__));
  or1   g3968(.dina(new_new_n8500__), .dinb(new_new_n8492__), .dout(new_new_n4910__));
  and1  g3969(.dina(new_new_n9674__), .dinb(new_new_n9675__), .dout(new_new_n4911__));
  or1   g3970(.dina(new_new_n9676__), .dinb(new_new_n9677__), .dout(new_new_n4912__));
  and1  g3971(.dina(new_new_n9679__), .dinb(new_new_n9675__), .dout(new_new_n4913__));
  or1   g3972(.dina(new_new_n9681__), .dinb(new_new_n9677__), .dout(new_new_n4914__));
  and1  g3973(.dina(new_new_n9679__), .dinb(new_new_n9674__), .dout(new_new_n4915__));
  or1   g3974(.dina(new_new_n9681__), .dinb(new_new_n9676__), .dout(new_new_n4916__));
  and1  g3975(.dina(new_new_n4916__), .dinb(new_new_n4914__), .dout(new_new_n4917__));
  or1   g3976(.dina(new_new_n4915__), .dinb(new_new_n4913__), .dout(new_new_n4918__));
  and1  g3977(.dina(new_new_n7106__), .dinb(new_new_n7911__), .dout(new_new_n4919__));
  or1   g3978(.dina(new_new_n7111__), .dinb(new_new_n7926__), .dout(new_new_n4920__));
  and1  g3979(.dina(new_new_n9682__), .dinb(new_new_n9683__), .dout(new_new_n4921__));
  or1   g3980(.dina(new_new_n9684__), .dinb(new_new_n9685__), .dout(new_new_n4922__));
  and1  g3981(.dina(new_new_n9687__), .dinb(new_new_n9683__), .dout(new_new_n4923__));
  or1   g3982(.dina(new_new_n9689__), .dinb(new_new_n9685__), .dout(new_new_n4924__));
  and1  g3983(.dina(new_new_n9687__), .dinb(new_new_n9682__), .dout(new_new_n4925__));
  or1   g3984(.dina(new_new_n9689__), .dinb(new_new_n9684__), .dout(new_new_n4926__));
  and1  g3985(.dina(new_new_n4926__), .dinb(new_new_n4924__), .dout(new_new_n4927__));
  or1   g3986(.dina(new_new_n4925__), .dinb(new_new_n4923__), .dout(new_new_n4928__));
  and1  g3987(.dina(new_new_n3717__), .dinb(new_new_n8507__), .dout(new_new_n4929__));
  or1   g3988(.dina(new_new_n9690__), .dinb(new_new_n8509__), .dout(new_new_n4930__));
  and1  g3989(.dina(new_new_n9691__), .dinb(new_new_n9692__), .dout(new_new_n4931__));
  or1   g3990(.dina(new_new_n4929__), .dinb(new_new_n4927__), .dout(new_new_n4932__));
  and1  g3991(.dina(new_new_n9693__), .dinb(new_new_n9692__), .dout(new_new_n4933__));
  and1  g3992(.dina(new_new_n9693__), .dinb(new_new_n9691__), .dout(new_new_n4934__));
  or1   g3993(.dina(new_new_n4934__), .dinb(new_new_n4933__), .dout(new_new_n4935__));
  or1   g3994(.dina(new_new_n7988__), .dinb(new_new_n7616__), .dout(new_new_n4936__));
  or1   g3995(.dina(new_new_n8137__), .dinb(new_new_n8376__), .dout(new_new_n4937__));
  or1   g3996(.dina(new_new_n8310__), .dinb(new_new_n8998__), .dout(new_new_n4938__));
  or1   g3997(.dina(new_new_n7636__), .dinb(new_new_n8999__), .dout(new_new_n4939__));
  and1  g3998(.dina(new_new_n8591__), .dinb(new_new_n8584__), .dout(new_new_n4940__));
  and1  g3999(.dina(new_new_n8605__), .dinb(new_new_n8598__), .dout(new_new_n4941__));
  and1  g4000(.dina(new_new_n8619__), .dinb(new_new_n8612__), .dout(new_new_n4942__));
  and1  g4001(.dina(new_new_n9695__), .dinb(new_new_n3821__), .dout(new_new_n4943__));
  and1  g4002(.dina(new_new_n9697__), .dinb(new_new_n3850__), .dout(new_new_n4944__));
  and1  g4003(.dina(new_new_n9699__), .dinb(new_new_n3879__), .dout(new_new_n4945__));
  and1  g4004(.dina(new_new_n9699__), .dinb(new_new_n3877__), .dout(new_new_n4946__));
  and1  g4005(.dina(new_new_n9697__), .dinb(new_new_n3848__), .dout(new_new_n4947__));
  and1  g4006(.dina(new_new_n9695__), .dinb(new_new_n3819__), .dout(new_new_n4948__));
  and1  g4007(.dina(new_new_n9700__), .dinb(new_new_n9701__), .dout(new_new_n4949__));
  and1  g4008(.dina(new_new_n9702__), .dinb(new_new_n9703__), .dout(new_new_n4950__));
  and1  g4009(.dina(new_new_n9704__), .dinb(new_new_n9705__), .dout(new_new_n4951__));
  and1  g4010(.dina(new_new_n9706__), .dinb(new_new_n9707__), .dout(new_new_n4952__));
  and1  g4011(.dina(new_new_n9709__), .dinb(new_new_n3141__), .dout(new_new_n4953__));
  and1  g4012(.dina(new_new_n9709__), .dinb(new_new_n3143__), .dout(new_new_n4954__));
  or1   g4013(.dina(new_new_n4954__), .dinb(new_new_n4953__), .dout(new_new_n4955__));
  and1  g4014(.dina(new_new_n9711__), .dinb(new_new_n3150__), .dout(new_new_n4956__));
  and1  g4015(.dina(new_new_n9711__), .dinb(new_new_n3152__), .dout(new_new_n4957__));
  or1   g4016(.dina(new_new_n4957__), .dinb(new_new_n4956__), .dout(new_new_n4958__));
  and1  g4017(.dina(new_new_n9713__), .dinb(new_new_n3159__), .dout(new_new_n4959__));
  and1  g4018(.dina(new_new_n9713__), .dinb(new_new_n3161__), .dout(new_new_n4960__));
  or1   g4019(.dina(new_new_n4960__), .dinb(new_new_n4959__), .dout(new_new_n4961__));
  and1  g4020(.dina(new_new_n7943__), .dinb(new_new_n7030__), .dout(new_new_n4962__));
  or1   g4021(.dina(new_new_n7944__), .dinb(new_new_n7045__), .dout(new_new_n4963__));
  and1  g4022(.dina(new_new_n8644__), .dinb(new_new_n8636__), .dout(new_new_n4964__));
  or1   g4023(.dina(new_new_n8646__), .dinb(new_new_n8638__), .dout(new_new_n4965__));
  or1   g4024(.dina(new_new_n4964__), .dinb(new_new_n4962__), .dout(new_new_n4966__));
  and1  g4025(.dina(new_new_n8067__), .dinb(new_new_n8063__), .dout(new_new_n4967__));
  or1   g4026(.dina(new_new_n8069__), .dinb(new_new_n8065__), .dout(new_new_n4968__));
  and1  g4027(.dina(new_new_n8066__), .dinb(new_new_n8062__), .dout(new_new_n4969__));
  or1   g4028(.dina(new_new_n8068__), .dinb(new_new_n8064__), .dout(new_new_n4970__));
  and1  g4029(.dina(new_new_n4970__), .dinb(new_new_n4968__), .dout(new_new_n4971__));
  or1   g4030(.dina(new_new_n4969__), .dinb(new_new_n4967__), .dout(new_new_n4972__));
  and1  g4031(.dina(new_new_n8660__), .dinb(new_new_n8652__), .dout(new_new_n4973__));
  or1   g4032(.dina(new_new_n8662__), .dinb(new_new_n8654__), .dout(new_new_n4974__));
  and1  g4033(.dina(new_new_n9714__), .dinb(new_new_n9715__), .dout(new_new_n4975__));
  or1   g4034(.dina(new_new_n9716__), .dinb(new_new_n9717__), .dout(new_new_n4976__));
  and1  g4035(.dina(new_new_n9719__), .dinb(new_new_n9715__), .dout(new_new_n4977__));
  or1   g4036(.dina(new_new_n9720__), .dinb(new_new_n9717__), .dout(new_new_n4978__));
  and1  g4037(.dina(new_new_n9719__), .dinb(new_new_n9714__), .dout(new_new_n4979__));
  or1   g4038(.dina(new_new_n9720__), .dinb(new_new_n9716__), .dout(new_new_n4980__));
  and1  g4039(.dina(new_new_n4980__), .dinb(new_new_n4978__), .dout(new_new_n4981__));
  or1   g4040(.dina(new_new_n4979__), .dinb(new_new_n4977__), .dout(new_new_n4982__));
  and1  g4041(.dina(new_new_n8084__), .dinb(new_new_n7603__), .dout(new_new_n4983__));
  or1   g4042(.dina(new_new_n8085__), .dinb(new_new_n7616__), .dout(new_new_n4984__));
  and1  g4043(.dina(new_new_n9721__), .dinb(new_new_n9722__), .dout(new_new_n4985__));
  or1   g4044(.dina(new_new_n9723__), .dinb(new_new_n9724__), .dout(new_new_n4986__));
  and1  g4045(.dina(new_new_n9726__), .dinb(new_new_n9722__), .dout(new_new_n4987__));
  or1   g4046(.dina(new_new_n9727__), .dinb(new_new_n9724__), .dout(new_new_n4988__));
  and1  g4047(.dina(new_new_n9726__), .dinb(new_new_n9721__), .dout(new_new_n4989__));
  or1   g4048(.dina(new_new_n9727__), .dinb(new_new_n9723__), .dout(new_new_n4990__));
  and1  g4049(.dina(new_new_n4990__), .dinb(new_new_n4988__), .dout(new_new_n4991__));
  or1   g4050(.dina(new_new_n4989__), .dinb(new_new_n4987__), .dout(new_new_n4992__));
  and1  g4051(.dina(new_new_n8676__), .dinb(new_new_n8668__), .dout(new_new_n4993__));
  or1   g4052(.dina(new_new_n8678__), .dinb(new_new_n8670__), .dout(new_new_n4994__));
  or1   g4053(.dina(new_new_n4993__), .dinb(new_new_n4991__), .dout(new_new_n4995__));
  and1  g4054(.dina(new_new_n8216__), .dinb(new_new_n8212__), .dout(new_new_n4996__));
  or1   g4055(.dina(new_new_n8218__), .dinb(new_new_n8214__), .dout(new_new_n4997__));
  and1  g4056(.dina(new_new_n8215__), .dinb(new_new_n8211__), .dout(new_new_n4998__));
  or1   g4057(.dina(new_new_n8217__), .dinb(new_new_n8213__), .dout(new_new_n4999__));
  and1  g4058(.dina(new_new_n4999__), .dinb(new_new_n4997__), .dout(new_new_n5000__));
  or1   g4059(.dina(new_new_n4998__), .dinb(new_new_n4996__), .dout(new_new_n5001__));
  and1  g4060(.dina(new_new_n8692__), .dinb(new_new_n8684__), .dout(new_new_n5002__));
  or1   g4061(.dina(new_new_n8694__), .dinb(new_new_n8686__), .dout(new_new_n5003__));
  and1  g4062(.dina(new_new_n9728__), .dinb(new_new_n9729__), .dout(new_new_n5004__));
  or1   g4063(.dina(new_new_n9730__), .dinb(new_new_n9731__), .dout(new_new_n5005__));
  and1  g4064(.dina(new_new_n9733__), .dinb(new_new_n9729__), .dout(new_new_n5006__));
  or1   g4065(.dina(new_new_n9734__), .dinb(new_new_n9731__), .dout(new_new_n5007__));
  and1  g4066(.dina(new_new_n9733__), .dinb(new_new_n9728__), .dout(new_new_n5008__));
  or1   g4067(.dina(new_new_n9734__), .dinb(new_new_n9730__), .dout(new_new_n5009__));
  and1  g4068(.dina(new_new_n5009__), .dinb(new_new_n5007__), .dout(new_new_n5010__));
  or1   g4069(.dina(new_new_n5008__), .dinb(new_new_n5006__), .dout(new_new_n5011__));
  and1  g4070(.dina(new_new_n8241__), .dinb(new_new_n8367__), .dout(new_new_n5012__));
  or1   g4071(.dina(new_new_n8242__), .dinb(new_new_n8376__), .dout(new_new_n5013__));
  and1  g4072(.dina(new_new_n9735__), .dinb(new_new_n9736__), .dout(new_new_n5014__));
  or1   g4073(.dina(new_new_n9737__), .dinb(new_new_n9738__), .dout(new_new_n5015__));
  and1  g4074(.dina(new_new_n9740__), .dinb(new_new_n9736__), .dout(new_new_n5016__));
  or1   g4075(.dina(new_new_n9741__), .dinb(new_new_n9738__), .dout(new_new_n5017__));
  and1  g4076(.dina(new_new_n9740__), .dinb(new_new_n9735__), .dout(new_new_n5018__));
  or1   g4077(.dina(new_new_n9741__), .dinb(new_new_n9737__), .dout(new_new_n5019__));
  and1  g4078(.dina(new_new_n5019__), .dinb(new_new_n5017__), .dout(new_new_n5020__));
  or1   g4079(.dina(new_new_n5018__), .dinb(new_new_n5016__), .dout(new_new_n5021__));
  and1  g4080(.dina(new_new_n8708__), .dinb(new_new_n8700__), .dout(new_new_n5022__));
  or1   g4081(.dina(new_new_n8710__), .dinb(new_new_n8702__), .dout(new_new_n5023__));
  or1   g4082(.dina(new_new_n5022__), .dinb(new_new_n5020__), .dout(new_new_n5024__));
  and1  g4083(.dina(new_new_n9013__), .dinb(new_new_n9009__), .dout(new_new_n5025__));
  or1   g4084(.dina(new_new_n9015__), .dinb(new_new_n9011__), .dout(new_new_n5026__));
  and1  g4085(.dina(new_new_n9012__), .dinb(new_new_n9008__), .dout(new_new_n5027__));
  or1   g4086(.dina(new_new_n9014__), .dinb(new_new_n9010__), .dout(new_new_n5028__));
  and1  g4087(.dina(new_new_n5028__), .dinb(new_new_n5026__), .dout(new_new_n5029__));
  or1   g4088(.dina(new_new_n5027__), .dinb(new_new_n5025__), .dout(new_new_n5030__));
  and1  g4089(.dina(new_new_n3894__), .dinb(new_new_n8575__), .dout(new_new_n5031__));
  or1   g4090(.dina(new_new_n9742__), .dinb(new_new_n8577__), .dout(new_new_n5032__));
  or1   g4091(.dina(new_new_n5031__), .dinb(new_new_n5029__), .dout(new_new_n5033__));
  and1  g4092(.dina(new_new_n9744__), .dinb(new_new_n3916__), .dout(new_new_n5034__));
  and1  g4093(.dina(new_new_n9744__), .dinb(new_new_n3918__), .dout(new_new_n5035__));
  or1   g4094(.dina(new_new_n5035__), .dinb(new_new_n5034__), .dout(new_new_n5036__));
  and1  g4095(.dina(new_new_n9746__), .dinb(new_new_n3965__), .dout(new_new_n5037__));
  and1  g4096(.dina(new_new_n9746__), .dinb(new_new_n3967__), .dout(new_new_n5038__));
  or1   g4097(.dina(new_new_n5038__), .dinb(new_new_n5037__), .dout(new_new_n5039__));
  and1  g4098(.dina(new_new_n9748__), .dinb(new_new_n4014__), .dout(new_new_n5040__));
  and1  g4099(.dina(new_new_n9748__), .dinb(new_new_n4016__), .dout(new_new_n5041__));
  or1   g4100(.dina(new_new_n5041__), .dinb(new_new_n5040__), .dout(new_new_n5042__));
  and1  g4101(.dina(new_new_n9750__), .dinb(new_new_n4083__), .dout(new_new_n5043__));
  and1  g4102(.dina(new_new_n9750__), .dinb(new_new_n4125__), .dout(new_new_n5044__));
  or1   g4103(.dina(new_new_n5044__), .dinb(new_new_n5043__), .dout(new_new_n5045__));
  and1  g4104(.dina(new_new_n9752__), .dinb(new_new_n8982__), .dout(new_new_n5046__));
  or1   g4105(.dina(new_new_n9753__), .dinb(new_new_n8984__), .dout(new_new_n5047__));
  and1  g4106(.dina(new_new_n9752__), .dinb(new_new_n8981__), .dout(new_new_n5048__));
  or1   g4107(.dina(new_new_n9753__), .dinb(new_new_n8983__), .dout(new_new_n5049__));
  and1  g4108(.dina(new_new_n5049__), .dinb(new_new_n5047__), .dout(new_new_n5050__));
  or1   g4109(.dina(new_new_n5048__), .dinb(new_new_n5046__), .dout(new_new_n5051__));
  and1  g4110(.dina(new_new_n8937__), .dinb(new_new_n9556__), .dout(new_new_n5052__));
  or1   g4111(.dina(new_new_n8940__), .dinb(new_new_n9565__), .dout(new_new_n5053__));
  or1   g4112(.dina(new_new_n5052__), .dinb(new_new_n5050__), .dout(new_new_n5054__));
  and1  g4113(.dina(new_new_n9754__), .dinb(new_new_n9755__), .dout(new_new_n5055__));
  and1  g4114(.dina(new_new_n9427__), .dinb(new_new_n9423__), .dout(new_new_n5056__));
  or1   g4115(.dina(new_new_n9429__), .dinb(new_new_n9425__), .dout(new_new_n5057__));
  and1  g4116(.dina(new_new_n9426__), .dinb(new_new_n9422__), .dout(new_new_n5058__));
  or1   g4117(.dina(new_new_n9428__), .dinb(new_new_n9424__), .dout(new_new_n5059__));
  and1  g4118(.dina(new_new_n5059__), .dinb(new_new_n5057__), .dout(new_new_n5060__));
  or1   g4119(.dina(new_new_n5058__), .dinb(new_new_n5056__), .dout(new_new_n5061__));
  and1  g4120(.dina(new_new_n9411__), .dinb(new_new_n9407__), .dout(new_new_n5062__));
  or1   g4121(.dina(new_new_n9413__), .dinb(new_new_n9409__), .dout(new_new_n5063__));
  and1  g4122(.dina(new_new_n9410__), .dinb(new_new_n9406__), .dout(new_new_n5064__));
  or1   g4123(.dina(new_new_n9412__), .dinb(new_new_n9408__), .dout(new_new_n5065__));
  and1  g4124(.dina(new_new_n5065__), .dinb(new_new_n5063__), .dout(new_new_n5066__));
  or1   g4125(.dina(new_new_n5064__), .dinb(new_new_n5062__), .dout(new_new_n5067__));
  and1  g4126(.dina(new_new_n9395__), .dinb(new_new_n9391__), .dout(new_new_n5068__));
  or1   g4127(.dina(new_new_n9397__), .dinb(new_new_n9393__), .dout(new_new_n5069__));
  and1  g4128(.dina(new_new_n9394__), .dinb(new_new_n9390__), .dout(new_new_n5070__));
  or1   g4129(.dina(new_new_n9396__), .dinb(new_new_n9392__), .dout(new_new_n5071__));
  and1  g4130(.dina(new_new_n5071__), .dinb(new_new_n5069__), .dout(new_new_n5072__));
  or1   g4131(.dina(new_new_n5070__), .dinb(new_new_n5068__), .dout(new_new_n5073__));
  and1  g4132(.dina(new_new_n9670__), .dinb(new_new_n9662__), .dout(new_new_n5074__));
  or1   g4133(.dina(new_new_n9672__), .dinb(new_new_n9664__), .dout(new_new_n5075__));
  and1  g4134(.dina(new_new_n9756__), .dinb(new_new_n9757__), .dout(new_new_n5076__));
  or1   g4135(.dina(new_new_n9758__), .dinb(new_new_n9759__), .dout(new_new_n5077__));
  and1  g4136(.dina(new_new_n9761__), .dinb(new_new_n9757__), .dout(new_new_n5078__));
  or1   g4137(.dina(new_new_n9763__), .dinb(new_new_n9759__), .dout(new_new_n5079__));
  and1  g4138(.dina(new_new_n9761__), .dinb(new_new_n9756__), .dout(new_new_n5080__));
  or1   g4139(.dina(new_new_n9763__), .dinb(new_new_n9758__), .dout(new_new_n5081__));
  and1  g4140(.dina(new_new_n5081__), .dinb(new_new_n5079__), .dout(new_new_n5082__));
  or1   g4141(.dina(new_new_n5080__), .dinb(new_new_n5078__), .dout(new_new_n5083__));
  and1  g4142(.dina(new_new_n7705__), .dinb(new_new_n7913__), .dout(new_new_n5084__));
  or1   g4143(.dina(new_new_n7711__), .dinb(new_new_n7928__), .dout(new_new_n5085__));
  and1  g4144(.dina(new_new_n9764__), .dinb(new_new_n9765__), .dout(new_new_n5086__));
  or1   g4145(.dina(new_new_n9766__), .dinb(new_new_n9767__), .dout(new_new_n5087__));
  and1  g4146(.dina(new_new_n9769__), .dinb(new_new_n9760__), .dout(new_new_n5088__));
  or1   g4147(.dina(new_new_n9771__), .dinb(new_new_n9762__), .dout(new_new_n5089__));
  and1  g4148(.dina(new_new_n9772__), .dinb(new_new_n9773__), .dout(new_new_n5090__));
  or1   g4149(.dina(new_new_n9774__), .dinb(new_new_n9775__), .dout(new_new_n5091__));
  and1  g4150(.dina(new_new_n9777__), .dinb(new_new_n9773__), .dout(new_new_n5092__));
  or1   g4151(.dina(new_new_n9779__), .dinb(new_new_n9775__), .dout(new_new_n5093__));
  and1  g4152(.dina(new_new_n9777__), .dinb(new_new_n9772__), .dout(new_new_n5094__));
  or1   g4153(.dina(new_new_n9779__), .dinb(new_new_n9774__), .dout(new_new_n5095__));
  and1  g4154(.dina(new_new_n5095__), .dinb(new_new_n5093__), .dout(new_new_n5096__));
  or1   g4155(.dina(new_new_n5094__), .dinb(new_new_n5092__), .dout(new_new_n5097__));
  and1  g4156(.dina(new_new_n7707__), .dinb(new_new_n8904__), .dout(new_new_n5098__));
  or1   g4157(.dina(new_new_n7711__), .dinb(new_new_n8918__), .dout(new_new_n5099__));
  and1  g4158(.dina(new_new_n9780__), .dinb(new_new_n9781__), .dout(new_new_n5100__));
  or1   g4159(.dina(new_new_n9782__), .dinb(new_new_n9783__), .dout(new_new_n5101__));
  and1  g4160(.dina(new_new_n9785__), .dinb(new_new_n9776__), .dout(new_new_n5102__));
  or1   g4161(.dina(new_new_n9787__), .dinb(new_new_n9778__), .dout(new_new_n5103__));
  or1   g4162(.dina(new_new_n5102__), .dinb(new_new_n5060__), .dout(new_new_n5104__));
  and1  g4163(.dina(new_new_n9655__), .dinb(new_new_n9651__), .dout(new_new_n5105__));
  or1   g4164(.dina(new_new_n9657__), .dinb(new_new_n9653__), .dout(new_new_n5106__));
  and1  g4165(.dina(new_new_n9654__), .dinb(new_new_n9650__), .dout(new_new_n5107__));
  or1   g4166(.dina(new_new_n9656__), .dinb(new_new_n9652__), .dout(new_new_n5108__));
  and1  g4167(.dina(new_new_n5108__), .dinb(new_new_n5106__), .dout(new_new_n5109__));
  or1   g4168(.dina(new_new_n5107__), .dinb(new_new_n5105__), .dout(new_new_n5110__));
  and1  g4169(.dina(new_new_n9639__), .dinb(new_new_n9635__), .dout(new_new_n5111__));
  or1   g4170(.dina(new_new_n9641__), .dinb(new_new_n9637__), .dout(new_new_n5112__));
  and1  g4171(.dina(new_new_n9638__), .dinb(new_new_n9634__), .dout(new_new_n5113__));
  or1   g4172(.dina(new_new_n9640__), .dinb(new_new_n9636__), .dout(new_new_n5114__));
  and1  g4173(.dina(new_new_n5114__), .dinb(new_new_n5112__), .dout(new_new_n5115__));
  or1   g4174(.dina(new_new_n5113__), .dinb(new_new_n5111__), .dout(new_new_n5116__));
  and1  g4175(.dina(new_new_n9623__), .dinb(new_new_n9619__), .dout(new_new_n5117__));
  or1   g4176(.dina(new_new_n9625__), .dinb(new_new_n9621__), .dout(new_new_n5118__));
  and1  g4177(.dina(new_new_n9622__), .dinb(new_new_n9618__), .dout(new_new_n5119__));
  or1   g4178(.dina(new_new_n9624__), .dinb(new_new_n9620__), .dout(new_new_n5120__));
  and1  g4179(.dina(new_new_n5120__), .dinb(new_new_n5118__), .dout(new_new_n5121__));
  or1   g4180(.dina(new_new_n5119__), .dinb(new_new_n5117__), .dout(new_new_n5122__));
  and1  g4181(.dina(new_new_n9607__), .dinb(new_new_n9603__), .dout(new_new_n5123__));
  or1   g4182(.dina(new_new_n9609__), .dinb(new_new_n9605__), .dout(new_new_n5124__));
  and1  g4183(.dina(new_new_n9606__), .dinb(new_new_n9602__), .dout(new_new_n5125__));
  or1   g4184(.dina(new_new_n9608__), .dinb(new_new_n9604__), .dout(new_new_n5126__));
  and1  g4185(.dina(new_new_n5126__), .dinb(new_new_n5124__), .dout(new_new_n5127__));
  or1   g4186(.dina(new_new_n5125__), .dinb(new_new_n5123__), .dout(new_new_n5128__));
  and1  g4187(.dina(new_new_n9583__), .dinb(new_new_n9578__), .dout(new_new_n5129__));
  or1   g4188(.dina(new_new_n9585__), .dinb(new_new_n9580__), .dout(new_new_n5130__));
  and1  g4189(.dina(new_new_n9582__), .dinb(new_new_n9579__), .dout(new_new_n5131__));
  or1   g4190(.dina(new_new_n9584__), .dinb(new_new_n9581__), .dout(new_new_n5132__));
  and1  g4191(.dina(new_new_n5132__), .dinb(new_new_n5130__), .dout(new_new_n5133__));
  or1   g4192(.dina(new_new_n5131__), .dinb(new_new_n5129__), .dout(new_new_n5134__));
  and1  g4193(.dina(new_new_n9183__), .dinb(new_new_n1539__), .dout(new_new_n5135__));
  or1   g4194(.dina(new_new_n9185__), .dinb(new_new_n1540__), .dout(new_new_n5136__));
  and1  g4195(.dina(new_new_n9788__), .dinb(new_new_n9789__), .dout(new_new_n5137__));
  or1   g4196(.dina(new_new_n9790__), .dinb(new_new_n9791__), .dout(new_new_n5138__));
  and1  g4197(.dina(new_new_n9793__), .dinb(new_new_n9789__), .dout(new_new_n5139__));
  or1   g4198(.dina(new_new_n9795__), .dinb(new_new_n9791__), .dout(new_new_n5140__));
  and1  g4199(.dina(new_new_n9793__), .dinb(new_new_n9788__), .dout(new_new_n5141__));
  or1   g4200(.dina(new_new_n9795__), .dinb(new_new_n9790__), .dout(new_new_n5142__));
  and1  g4201(.dina(new_new_n5142__), .dinb(new_new_n5140__), .dout(new_new_n5143__));
  or1   g4202(.dina(new_new_n5141__), .dinb(new_new_n5139__), .dout(new_new_n5144__));
  and1  g4203(.dina(new_new_n7684__), .dinb(new_new_n9171__), .dout(new_new_n5145__));
  or1   g4204(.dina(new_new_n7699__), .dinb(new_new_n9177__), .dout(new_new_n5146__));
  and1  g4205(.dina(new_new_n9796__), .dinb(new_new_n9797__), .dout(new_new_n5147__));
  or1   g4206(.dina(new_new_n9798__), .dinb(new_new_n9799__), .dout(new_new_n5148__));
  and1  g4207(.dina(new_new_n9801__), .dinb(new_new_n9792__), .dout(new_new_n5149__));
  or1   g4208(.dina(new_new_n9803__), .dinb(new_new_n9794__), .dout(new_new_n5150__));
  and1  g4209(.dina(new_new_n9804__), .dinb(new_new_n9805__), .dout(new_new_n5151__));
  or1   g4210(.dina(new_new_n9806__), .dinb(new_new_n9807__), .dout(new_new_n5152__));
  and1  g4211(.dina(new_new_n9809__), .dinb(new_new_n9805__), .dout(new_new_n5153__));
  or1   g4212(.dina(new_new_n9811__), .dinb(new_new_n9807__), .dout(new_new_n5154__));
  and1  g4213(.dina(new_new_n9809__), .dinb(new_new_n9804__), .dout(new_new_n5155__));
  or1   g4214(.dina(new_new_n9811__), .dinb(new_new_n9806__), .dout(new_new_n5156__));
  and1  g4215(.dina(new_new_n5156__), .dinb(new_new_n5154__), .dout(new_new_n5157__));
  or1   g4216(.dina(new_new_n5155__), .dinb(new_new_n5153__), .dout(new_new_n5158__));
  and1  g4217(.dina(new_new_n9172__), .dinb(new_new_n7913__), .dout(new_new_n5159__));
  or1   g4218(.dina(new_new_n9176__), .dinb(new_new_n7928__), .dout(new_new_n5160__));
  and1  g4219(.dina(new_new_n9812__), .dinb(new_new_n9813__), .dout(new_new_n5161__));
  or1   g4220(.dina(new_new_n9814__), .dinb(new_new_n9815__), .dout(new_new_n5162__));
  and1  g4221(.dina(new_new_n9817__), .dinb(new_new_n9808__), .dout(new_new_n5163__));
  or1   g4222(.dina(new_new_n9819__), .dinb(new_new_n9810__), .dout(new_new_n5164__));
  and1  g4223(.dina(new_new_n9820__), .dinb(new_new_n9821__), .dout(new_new_n5165__));
  or1   g4224(.dina(new_new_n9822__), .dinb(new_new_n9823__), .dout(new_new_n5166__));
  and1  g4225(.dina(new_new_n9825__), .dinb(new_new_n9821__), .dout(new_new_n5167__));
  or1   g4226(.dina(new_new_n9827__), .dinb(new_new_n9823__), .dout(new_new_n5168__));
  and1  g4227(.dina(new_new_n9825__), .dinb(new_new_n9820__), .dout(new_new_n5169__));
  or1   g4228(.dina(new_new_n9827__), .dinb(new_new_n9822__), .dout(new_new_n5170__));
  and1  g4229(.dina(new_new_n5170__), .dinb(new_new_n5168__), .dout(new_new_n5171__));
  or1   g4230(.dina(new_new_n5169__), .dinb(new_new_n5167__), .dout(new_new_n5172__));
  and1  g4231(.dina(new_new_n9172__), .dinb(new_new_n8904__), .dout(new_new_n5173__));
  or1   g4232(.dina(new_new_n9178__), .dinb(new_new_n8919__), .dout(new_new_n5174__));
  and1  g4233(.dina(new_new_n9828__), .dinb(new_new_n9829__), .dout(new_new_n5175__));
  or1   g4234(.dina(new_new_n9830__), .dinb(new_new_n9831__), .dout(new_new_n5176__));
  and1  g4235(.dina(new_new_n9833__), .dinb(new_new_n9824__), .dout(new_new_n5177__));
  or1   g4236(.dina(new_new_n9835__), .dinb(new_new_n9826__), .dout(new_new_n5178__));
  and1  g4237(.dina(new_new_n9836__), .dinb(new_new_n9837__), .dout(new_new_n5179__));
  or1   g4238(.dina(new_new_n9838__), .dinb(new_new_n9839__), .dout(new_new_n5180__));
  and1  g4239(.dina(new_new_n9841__), .dinb(new_new_n9837__), .dout(new_new_n5181__));
  or1   g4240(.dina(new_new_n9843__), .dinb(new_new_n9839__), .dout(new_new_n5182__));
  and1  g4241(.dina(new_new_n9841__), .dinb(new_new_n9836__), .dout(new_new_n5183__));
  or1   g4242(.dina(new_new_n9843__), .dinb(new_new_n9838__), .dout(new_new_n5184__));
  and1  g4243(.dina(new_new_n5184__), .dinb(new_new_n5182__), .dout(new_new_n5185__));
  or1   g4244(.dina(new_new_n5183__), .dinb(new_new_n5181__), .dout(new_new_n5186__));
  and1  g4245(.dina(new_new_n9174__), .dinb(new_new_n9556__), .dout(new_new_n5187__));
  or1   g4246(.dina(new_new_n9178__), .dinb(new_new_n9565__), .dout(new_new_n5188__));
  and1  g4247(.dina(new_new_n9844__), .dinb(new_new_n9845__), .dout(new_new_n5189__));
  or1   g4248(.dina(new_new_n9846__), .dinb(new_new_n9847__), .dout(new_new_n5190__));
  and1  g4249(.dina(new_new_n9849__), .dinb(new_new_n9840__), .dout(new_new_n5191__));
  or1   g4250(.dina(new_new_n9851__), .dinb(new_new_n9842__), .dout(new_new_n5192__));
  or1   g4251(.dina(new_new_n5191__), .dinb(new_new_n5109__), .dout(new_new_n5193__));
  and1  g4252(.dina(new_new_n9076__), .dinb(new_new_n9853__), .dout(new_new_n5194__));
  or1   g4253(.dina(new_new_n9091__), .dinb(new_new_n9856__), .dout(new_new_n5195__));
  and1  g4254(.dina(new_new_n9048__), .dinb(new_new_n9858__), .dout(new_new_n5196__));
  or1   g4255(.dina(new_new_n9062__), .dinb(new_new_n9861__), .dout(new_new_n5197__));
  and1  g4256(.dina(new_new_n9862__), .dinb(new_new_n9863__), .dout(new_new_n5198__));
  or1   g4257(.dina(new_new_n9864__), .dinb(new_new_n9865__), .dout(new_new_n5199__));
  and1  g4258(.dina(new_new_n9866__), .dinb(new_new_n9863__), .dout(new_new_n5200__));
  or1   g4259(.dina(new_new_n9867__), .dinb(new_new_n9865__), .dout(new_new_n5201__));
  and1  g4260(.dina(new_new_n9866__), .dinb(new_new_n9862__), .dout(new_new_n5202__));
  or1   g4261(.dina(new_new_n9867__), .dinb(new_new_n9864__), .dout(new_new_n5203__));
  and1  g4262(.dina(new_new_n5203__), .dinb(new_new_n9869__), .dout(new_new_n5204__));
  or1   g4263(.dina(new_new_n5202__), .dinb(new_new_n9871__), .dout(new_new_n5205__));
  and1  g4264(.dina(new_new_n9077__), .dinb(new_new_n9858__), .dout(new_new_n5206__));
  or1   g4265(.dina(new_new_n9092__), .dinb(new_new_n9861__), .dout(new_new_n5207__));
  and1  g4266(.dina(new_new_n9048__), .dinb(new_new_n9873__), .dout(new_new_n5208__));
  or1   g4267(.dina(new_new_n9062__), .dinb(new_new_n9875__), .dout(new_new_n5209__));
  and1  g4268(.dina(new_new_n9876__), .dinb(new_new_n9877__), .dout(new_new_n5210__));
  or1   g4269(.dina(new_new_n9878__), .dinb(new_new_n9879__), .dout(new_new_n5211__));
  and1  g4270(.dina(new_new_n9880__), .dinb(new_new_n9877__), .dout(new_new_n5212__));
  or1   g4271(.dina(new_new_n9881__), .dinb(new_new_n9879__), .dout(new_new_n5213__));
  or1   g4272(.dina(new_new_n9882__), .dinb(new_new_n5204__), .dout(new_new_n5214__));
  and1  g4273(.dina(new_new_n9077__), .dinb(new_new_n9885__), .dout(new_new_n5215__));
  or1   g4274(.dina(new_new_n9092__), .dinb(new_new_n9888__), .dout(new_new_n5216__));
  and1  g4275(.dina(new_new_n9050__), .dinb(new_new_n9892__), .dout(new_new_n5217__));
  or1   g4276(.dina(new_new_n9064__), .dinb(new_new_n9895__), .dout(new_new_n5218__));
  and1  g4277(.dina(new_new_n9897__), .dinb(new_new_n9898__), .dout(new_new_n5219__));
  or1   g4278(.dina(new_new_n9899__), .dinb(new_new_n9900__), .dout(new_new_n5220__));
  and1  g4279(.dina(new_new_n9901__), .dinb(new_new_n9898__), .dout(new_new_n5221__));
  or1   g4280(.dina(new_new_n9902__), .dinb(new_new_n9900__), .dout(new_new_n5222__));
  and1  g4281(.dina(new_new_n9901__), .dinb(new_new_n9897__), .dout(new_new_n5223__));
  or1   g4282(.dina(new_new_n9902__), .dinb(new_new_n9899__), .dout(new_new_n5224__));
  and1  g4283(.dina(new_new_n5224__), .dinb(new_new_n9904__), .dout(new_new_n5225__));
  or1   g4284(.dina(new_new_n5223__), .dinb(new_new_n9906__), .dout(new_new_n5226__));
  and1  g4285(.dina(new_new_n9079__), .dinb(new_new_n9892__), .dout(new_new_n5227__));
  or1   g4286(.dina(new_new_n9094__), .dinb(new_new_n9895__), .dout(new_new_n5228__));
  and1  g4287(.dina(new_new_n9050__), .dinb(new_new_n9909__), .dout(new_new_n5229__));
  or1   g4288(.dina(new_new_n9064__), .dinb(new_new_n9912__), .dout(new_new_n5230__));
  and1  g4289(.dina(new_new_n9914__), .dinb(new_new_n9915__), .dout(new_new_n5231__));
  or1   g4290(.dina(new_new_n9916__), .dinb(new_new_n9917__), .dout(new_new_n5232__));
  and1  g4291(.dina(new_new_n9918__), .dinb(new_new_n9915__), .dout(new_new_n5233__));
  or1   g4292(.dina(new_new_n9919__), .dinb(new_new_n9917__), .dout(new_new_n5234__));
  and1  g4293(.dina(new_new_n9921__), .dinb(new_new_n9922__), .dout(new_new_n5235__));
  or1   g4294(.dina(new_new_n9924__), .dinb(new_new_n9925__), .dout(new_new_n5236__));
  and1  g4295(.dina(new_new_n9927__), .dinb(new_new_n9922__), .dout(new_new_n5237__));
  or1   g4296(.dina(new_new_n9929__), .dinb(new_new_n9925__), .dout(new_new_n5238__));
  and1  g4297(.dina(new_new_n9927__), .dinb(new_new_n9921__), .dout(new_new_n5239__));
  or1   g4298(.dina(new_new_n9929__), .dinb(new_new_n9924__), .dout(new_new_n5240__));
  and1  g4299(.dina(new_new_n5240__), .dinb(new_new_n5238__), .dout(new_new_n5241__));
  or1   g4300(.dina(new_new_n5239__), .dinb(new_new_n5237__), .dout(new_new_n5242__));
  and1  g4301(.dina(new_new_n9020__), .dinb(new_new_n9909__), .dout(new_new_n5243__));
  or1   g4302(.dina(new_new_n9035__), .dinb(new_new_n9912__), .dout(new_new_n5244__));
  and1  g4303(.dina(new_new_n9930__), .dinb(new_new_n9931__), .dout(new_new_n5245__));
  or1   g4304(.dina(new_new_n9932__), .dinb(new_new_n9933__), .dout(new_new_n5246__));
  and1  g4305(.dina(new_new_n9935__), .dinb(new_new_n9931__), .dout(new_new_n5247__));
  or1   g4306(.dina(new_new_n9937__), .dinb(new_new_n9933__), .dout(new_new_n5248__));
  and1  g4307(.dina(new_new_n9935__), .dinb(new_new_n9930__), .dout(new_new_n5249__));
  or1   g4308(.dina(new_new_n9937__), .dinb(new_new_n9932__), .dout(new_new_n5250__));
  and1  g4309(.dina(new_new_n5250__), .dinb(new_new_n5248__), .dout(new_new_n5251__));
  or1   g4310(.dina(new_new_n5249__), .dinb(new_new_n5247__), .dout(new_new_n5252__));
  and1  g4311(.dina(new_new_n9918__), .dinb(new_new_n9914__), .dout(new_new_n5253__));
  or1   g4312(.dina(new_new_n9919__), .dinb(new_new_n9916__), .dout(new_new_n5254__));
  and1  g4313(.dina(new_new_n5254__), .dinb(new_new_n9920__), .dout(new_new_n5255__));
  or1   g4314(.dina(new_new_n5253__), .dinb(new_new_n9923__), .dout(new_new_n5256__));
  and1  g4315(.dina(new_new_n9079__), .dinb(new_new_n9908__), .dout(new_new_n5257__));
  or1   g4316(.dina(new_new_n9094__), .dinb(new_new_n9913__), .dout(new_new_n5258__));
  and1  g4317(.dina(new_new_n9051__), .dinb(new_new_n9939__), .dout(new_new_n5259__));
  or1   g4318(.dina(new_new_n9065__), .dinb(new_new_n9942__), .dout(new_new_n5260__));
  and1  g4319(.dina(new_new_n9944__), .dinb(new_new_n9945__), .dout(new_new_n5261__));
  or1   g4320(.dina(new_new_n9946__), .dinb(new_new_n9947__), .dout(new_new_n5262__));
  and1  g4321(.dina(new_new_n9948__), .dinb(new_new_n9945__), .dout(new_new_n5263__));
  or1   g4322(.dina(new_new_n9949__), .dinb(new_new_n9947__), .dout(new_new_n5264__));
  and1  g4323(.dina(new_new_n9951__), .dinb(new_new_n9952__), .dout(new_new_n5265__));
  or1   g4324(.dina(new_new_n9954__), .dinb(new_new_n9955__), .dout(new_new_n5266__));
  and1  g4325(.dina(new_new_n9957__), .dinb(new_new_n9952__), .dout(new_new_n5267__));
  or1   g4326(.dina(new_new_n9959__), .dinb(new_new_n9955__), .dout(new_new_n5268__));
  and1  g4327(.dina(new_new_n9957__), .dinb(new_new_n9951__), .dout(new_new_n5269__));
  or1   g4328(.dina(new_new_n9959__), .dinb(new_new_n9954__), .dout(new_new_n5270__));
  and1  g4329(.dina(new_new_n5270__), .dinb(new_new_n5268__), .dout(new_new_n5271__));
  or1   g4330(.dina(new_new_n5269__), .dinb(new_new_n5267__), .dout(new_new_n5272__));
  and1  g4331(.dina(new_new_n9020__), .dinb(new_new_n9939__), .dout(new_new_n5273__));
  or1   g4332(.dina(new_new_n9035__), .dinb(new_new_n9942__), .dout(new_new_n5274__));
  and1  g4333(.dina(new_new_n9960__), .dinb(new_new_n9961__), .dout(new_new_n5275__));
  or1   g4334(.dina(new_new_n9962__), .dinb(new_new_n9963__), .dout(new_new_n5276__));
  and1  g4335(.dina(new_new_n9965__), .dinb(new_new_n9956__), .dout(new_new_n5277__));
  or1   g4336(.dina(new_new_n9967__), .dinb(new_new_n9958__), .dout(new_new_n5278__));
  or1   g4337(.dina(new_new_n5277__), .dinb(new_new_n5251__), .dout(new_new_n5279__));
  and1  g4338(.dina(new_new_n6972__), .dinb(new_new_n8995__), .dout(new_new_n5280__));
  or1   g4339(.dina(new_new_n8861__), .dinb(new_new_n9566__), .dout(new_new_n5281__));
  or1   g4340(.dina(new_new_n9601__), .dinb(new_new_n902__), .dout(new_new_n5282__));
  or1   g4341(.dina(new_new_n9373__), .dinb(new_new_n9566__), .dout(new_new_n5283__));
  or1   g4342(.dina(new_new_n9065__), .dinb(new_new_n810__), .dout(new_new_n5284__));
  and1  g4343(.dina(new_new_n9725__), .dinb(new_new_n9718__), .dout(new_new_n5285__));
  and1  g4344(.dina(new_new_n9739__), .dinb(new_new_n9732__), .dout(new_new_n5286__));
  and1  g4345(.dina(new_new_n8455__), .dinb(new_new_n8451__), .dout(new_new_n5287__));
  or1   g4346(.dina(new_new_n8457__), .dinb(new_new_n8453__), .dout(new_new_n5288__));
  and1  g4347(.dina(new_new_n8454__), .dinb(new_new_n8450__), .dout(new_new_n5289__));
  or1   g4348(.dina(new_new_n8456__), .dinb(new_new_n8452__), .dout(new_new_n5290__));
  and1  g4349(.dina(new_new_n5290__), .dinb(new_new_n5288__), .dout(new_new_n5291__));
  or1   g4350(.dina(new_new_n5289__), .dinb(new_new_n5287__), .dout(new_new_n5292__));
  and1  g4351(.dina(new_new_n8756__), .dinb(new_new_n8748__), .dout(new_new_n5293__));
  or1   g4352(.dina(new_new_n8758__), .dinb(new_new_n8750__), .dout(new_new_n5294__));
  and1  g4353(.dina(new_new_n9968__), .dinb(new_new_n9969__), .dout(new_new_n5295__));
  or1   g4354(.dina(new_new_n9970__), .dinb(new_new_n9971__), .dout(new_new_n5296__));
  and1  g4355(.dina(new_new_n9973__), .dinb(new_new_n9969__), .dout(new_new_n5297__));
  or1   g4356(.dina(new_new_n9974__), .dinb(new_new_n9971__), .dout(new_new_n5298__));
  and1  g4357(.dina(new_new_n9973__), .dinb(new_new_n9968__), .dout(new_new_n5299__));
  or1   g4358(.dina(new_new_n9974__), .dinb(new_new_n9970__), .dout(new_new_n5300__));
  and1  g4359(.dina(new_new_n5300__), .dinb(new_new_n5298__), .dout(new_new_n5301__));
  or1   g4360(.dina(new_new_n5299__), .dinb(new_new_n5297__), .dout(new_new_n5302__));
  and1  g4361(.dina(new_new_n8525__), .dinb(new_new_n8996__), .dout(new_new_n5303__));
  or1   g4362(.dina(new_new_n8529__), .dinb(new_new_n8999__), .dout(new_new_n5304__));
  or1   g4363(.dina(new_new_n5303__), .dinb(new_new_n5301__), .dout(new_new_n5305__));
  and1  g4364(.dina(new_new_n9976__), .dinb(new_new_n9972__), .dout(new_new_n5306__));
  or1   g4365(.dina(new_new_n9977__), .dinb(new_new_n4931__), .dout(new_new_n5307__));
  and1  g4366(.dina(new_new_n9817__), .dinb(new_new_n9813__), .dout(new_new_n5308__));
  or1   g4367(.dina(new_new_n9819__), .dinb(new_new_n9815__), .dout(new_new_n5309__));
  and1  g4368(.dina(new_new_n9816__), .dinb(new_new_n9812__), .dout(new_new_n5310__));
  or1   g4369(.dina(new_new_n9818__), .dinb(new_new_n9814__), .dout(new_new_n5311__));
  and1  g4370(.dina(new_new_n5311__), .dinb(new_new_n5309__), .dout(new_new_n5312__));
  or1   g4371(.dina(new_new_n5310__), .dinb(new_new_n5308__), .dout(new_new_n5313__));
  and1  g4372(.dina(new_new_n9801__), .dinb(new_new_n9797__), .dout(new_new_n5314__));
  or1   g4373(.dina(new_new_n9803__), .dinb(new_new_n9799__), .dout(new_new_n5315__));
  and1  g4374(.dina(new_new_n9800__), .dinb(new_new_n9796__), .dout(new_new_n5316__));
  or1   g4375(.dina(new_new_n9802__), .dinb(new_new_n9798__), .dout(new_new_n5317__));
  and1  g4376(.dina(new_new_n5317__), .dinb(new_new_n5315__), .dout(new_new_n5318__));
  or1   g4377(.dina(new_new_n5316__), .dinb(new_new_n5314__), .dout(new_new_n5319__));
  and1  g4378(.dina(new_new_n9220__), .dinb(new_new_n9212__), .dout(new_new_n5320__));
  or1   g4379(.dina(new_new_n9222__), .dinb(new_new_n9214__), .dout(new_new_n5321__));
  and1  g4380(.dina(new_new_n9978__), .dinb(new_new_n9979__), .dout(new_new_n5322__));
  or1   g4381(.dina(new_new_n9980__), .dinb(new_new_n9981__), .dout(new_new_n5323__));
  and1  g4382(.dina(new_new_n9983__), .dinb(new_new_n9979__), .dout(new_new_n5324__));
  or1   g4383(.dina(new_new_n9985__), .dinb(new_new_n9981__), .dout(new_new_n5325__));
  and1  g4384(.dina(new_new_n9983__), .dinb(new_new_n9978__), .dout(new_new_n5326__));
  or1   g4385(.dina(new_new_n9985__), .dinb(new_new_n9980__), .dout(new_new_n5327__));
  and1  g4386(.dina(new_new_n5327__), .dinb(new_new_n5325__), .dout(new_new_n5328__));
  or1   g4387(.dina(new_new_n5326__), .dinb(new_new_n5324__), .dout(new_new_n5329__));
  and1  g4388(.dina(new_new_n9194__), .dinb(new_new_n7914__), .dout(new_new_n5330__));
  or1   g4389(.dina(new_new_n9197__), .dinb(new_new_n7929__), .dout(new_new_n5331__));
  and1  g4390(.dina(new_new_n9986__), .dinb(new_new_n9987__), .dout(new_new_n5332__));
  or1   g4391(.dina(new_new_n9988__), .dinb(new_new_n9989__), .dout(new_new_n5333__));
  and1  g4392(.dina(new_new_n9991__), .dinb(new_new_n9982__), .dout(new_new_n5334__));
  or1   g4393(.dina(new_new_n9993__), .dinb(new_new_n9984__), .dout(new_new_n5335__));
  and1  g4394(.dina(new_new_n9994__), .dinb(new_new_n9995__), .dout(new_new_n5336__));
  or1   g4395(.dina(new_new_n9996__), .dinb(new_new_n9997__), .dout(new_new_n5337__));
  and1  g4396(.dina(new_new_n9999__), .dinb(new_new_n9995__), .dout(new_new_n5338__));
  or1   g4397(.dina(new_new_n10001__), .dinb(new_new_n9997__), .dout(new_new_n5339__));
  and1  g4398(.dina(new_new_n9999__), .dinb(new_new_n9994__), .dout(new_new_n5340__));
  or1   g4399(.dina(new_new_n10001__), .dinb(new_new_n9996__), .dout(new_new_n5341__));
  and1  g4400(.dina(new_new_n5341__), .dinb(new_new_n5339__), .dout(new_new_n5342__));
  or1   g4401(.dina(new_new_n5340__), .dinb(new_new_n5338__), .dout(new_new_n5343__));
  and1  g4402(.dina(new_new_n9194__), .dinb(new_new_n8905__), .dout(new_new_n5344__));
  or1   g4403(.dina(new_new_n9199__), .dinb(new_new_n8919__), .dout(new_new_n5345__));
  and1  g4404(.dina(new_new_n10002__), .dinb(new_new_n10003__), .dout(new_new_n5346__));
  or1   g4405(.dina(new_new_n10004__), .dinb(new_new_n10005__), .dout(new_new_n5347__));
  and1  g4406(.dina(new_new_n10007__), .dinb(new_new_n10003__), .dout(new_new_n5348__));
  or1   g4407(.dina(new_new_n10009__), .dinb(new_new_n10005__), .dout(new_new_n5349__));
  and1  g4408(.dina(new_new_n10007__), .dinb(new_new_n10002__), .dout(new_new_n5350__));
  or1   g4409(.dina(new_new_n10009__), .dinb(new_new_n10004__), .dout(new_new_n5351__));
  and1  g4410(.dina(new_new_n5351__), .dinb(new_new_n5349__), .dout(new_new_n5352__));
  or1   g4411(.dina(new_new_n5350__), .dinb(new_new_n5348__), .dout(new_new_n5353__));
  and1  g4412(.dina(new_new_n9991__), .dinb(new_new_n9987__), .dout(new_new_n5354__));
  or1   g4413(.dina(new_new_n9993__), .dinb(new_new_n9989__), .dout(new_new_n5355__));
  and1  g4414(.dina(new_new_n9990__), .dinb(new_new_n9986__), .dout(new_new_n5356__));
  or1   g4415(.dina(new_new_n9992__), .dinb(new_new_n9988__), .dout(new_new_n5357__));
  and1  g4416(.dina(new_new_n5357__), .dinb(new_new_n5355__), .dout(new_new_n5358__));
  or1   g4417(.dina(new_new_n5356__), .dinb(new_new_n5354__), .dout(new_new_n5359__));
  and1  g4418(.dina(new_new_n9277__), .dinb(new_new_n9269__), .dout(new_new_n5360__));
  or1   g4419(.dina(new_new_n9279__), .dinb(new_new_n9271__), .dout(new_new_n5361__));
  and1  g4420(.dina(new_new_n10010__), .dinb(new_new_n10011__), .dout(new_new_n5362__));
  or1   g4421(.dina(new_new_n10012__), .dinb(new_new_n10013__), .dout(new_new_n5363__));
  and1  g4422(.dina(new_new_n10015__), .dinb(new_new_n10011__), .dout(new_new_n5364__));
  or1   g4423(.dina(new_new_n10017__), .dinb(new_new_n10013__), .dout(new_new_n5365__));
  and1  g4424(.dina(new_new_n10015__), .dinb(new_new_n10010__), .dout(new_new_n5366__));
  or1   g4425(.dina(new_new_n10017__), .dinb(new_new_n10012__), .dout(new_new_n5367__));
  and1  g4426(.dina(new_new_n5367__), .dinb(new_new_n5365__), .dout(new_new_n5368__));
  or1   g4427(.dina(new_new_n5366__), .dinb(new_new_n5364__), .dout(new_new_n5369__));
  and1  g4428(.dina(new_new_n9235__), .dinb(new_new_n8905__), .dout(new_new_n5370__));
  or1   g4429(.dina(new_new_n9240__), .dinb(new_new_n8921__), .dout(new_new_n5371__));
  and1  g4430(.dina(new_new_n10018__), .dinb(new_new_n10019__), .dout(new_new_n5372__));
  or1   g4431(.dina(new_new_n10020__), .dinb(new_new_n10021__), .dout(new_new_n5373__));
  and1  g4432(.dina(new_new_n10023__), .dinb(new_new_n10014__), .dout(new_new_n5374__));
  or1   g4433(.dina(new_new_n10025__), .dinb(new_new_n10016__), .dout(new_new_n5375__));
  and1  g4434(.dina(new_new_n10026__), .dinb(new_new_n10027__), .dout(new_new_n5376__));
  or1   g4435(.dina(new_new_n10028__), .dinb(new_new_n10029__), .dout(new_new_n5377__));
  and1  g4436(.dina(new_new_n10031__), .dinb(new_new_n10027__), .dout(new_new_n5378__));
  or1   g4437(.dina(new_new_n10032__), .dinb(new_new_n10029__), .dout(new_new_n5379__));
  and1  g4438(.dina(new_new_n10031__), .dinb(new_new_n10026__), .dout(new_new_n5380__));
  or1   g4439(.dina(new_new_n10032__), .dinb(new_new_n10028__), .dout(new_new_n5381__));
  and1  g4440(.dina(new_new_n5381__), .dinb(new_new_n5379__), .dout(new_new_n5382__));
  or1   g4441(.dina(new_new_n5380__), .dinb(new_new_n5378__), .dout(new_new_n5383__));
  and1  g4442(.dina(new_new_n9236__), .dinb(new_new_n9557__), .dout(new_new_n5384__));
  or1   g4443(.dina(new_new_n9240__), .dinb(new_new_n9568__), .dout(new_new_n5385__));
  or1   g4444(.dina(new_new_n5384__), .dinb(new_new_n5382__), .dout(new_new_n5386__));
  and1  g4445(.dina(new_new_n10034__), .dinb(new_new_n10030__), .dout(new_new_n5387__));
  and1  g4446(.dina(new_new_n10036__), .dinb(new_new_n4963__), .dout(new_new_n5388__));
  and1  g4447(.dina(new_new_n9976__), .dinb(new_new_n5304__), .dout(new_new_n5389__));
  and1  g4448(.dina(new_new_n10036__), .dinb(new_new_n4965__), .dout(new_new_n5390__));
  and1  g4449(.dina(new_new_n10038__), .dinb(new_new_n4994__), .dout(new_new_n5391__));
  and1  g4450(.dina(new_new_n10040__), .dinb(new_new_n5023__), .dout(new_new_n5392__));
  and1  g4451(.dina(new_new_n10042__), .dinb(new_new_n5032__), .dout(new_new_n5393__));
  and1  g4452(.dina(new_new_n10038__), .dinb(new_new_n4992__), .dout(new_new_n5394__));
  and1  g4453(.dina(new_new_n10040__), .dinb(new_new_n5021__), .dout(new_new_n5395__));
  and1  g4454(.dina(new_new_n10042__), .dinb(new_new_n5030__), .dout(new_new_n5396__));
  and1  g4455(.dina(new_new_n9975__), .dinb(new_new_n5302__), .dout(new_new_n5397__));
  and1  g4456(.dina(new_new_n10043__), .dinb(new_new_n10044__), .dout(new_new_n5398__));
  and1  g4457(.dina(new_new_n10045__), .dinb(new_new_n10046__), .dout(new_new_n5399__));
  and1  g4458(.dina(new_new_n10047__), .dinb(new_new_n10048__), .dout(new_new_n5400__));
  and1  g4459(.dina(new_new_n10049__), .dinb(new_new_n10050__), .dout(new_new_n5401__));
  and1  g4460(.dina(new_new_n10052__), .dinb(new_new_n9134__), .dout(new_new_n5402__));
  or1   g4461(.dina(new_new_n10053__), .dinb(new_new_n9136__), .dout(new_new_n5403__));
  and1  g4462(.dina(new_new_n10052__), .dinb(new_new_n9133__), .dout(new_new_n5404__));
  or1   g4463(.dina(new_new_n10053__), .dinb(new_new_n9135__), .dout(new_new_n5405__));
  and1  g4464(.dina(new_new_n5405__), .dinb(new_new_n5403__), .dout(new_new_n5406__));
  or1   g4465(.dina(new_new_n5404__), .dinb(new_new_n5402__), .dout(new_new_n5407__));
  and1  g4466(.dina(new_new_n10056__), .dinb(new_new_n9103__), .dout(new_new_n5408__));
  or1   g4467(.dina(new_new_n10062__), .dinb(new_new_n9108__), .dout(new_new_n5409__));
  or1   g4468(.dina(new_new_n5408__), .dinb(new_new_n5406__), .dout(new_new_n5410__));
  and1  g4469(.dina(new_new_n8793__), .dinb(new_new_n7914__), .dout(new_new_n5411__));
  or1   g4470(.dina(new_new_n8796__), .dinb(new_new_n7929__), .dout(new_new_n5412__));
  and1  g4471(.dina(new_new_n9149__), .dinb(new_new_n9141__), .dout(new_new_n5413__));
  or1   g4472(.dina(new_new_n9151__), .dinb(new_new_n9143__), .dout(new_new_n5414__));
  and1  g4473(.dina(new_new_n10065__), .dinb(new_new_n10066__), .dout(new_new_n5415__));
  or1   g4474(.dina(new_new_n10067__), .dinb(new_new_n10068__), .dout(new_new_n5416__));
  and1  g4475(.dina(new_new_n10070__), .dinb(new_new_n10066__), .dout(new_new_n5417__));
  or1   g4476(.dina(new_new_n10071__), .dinb(new_new_n10068__), .dout(new_new_n5418__));
  and1  g4477(.dina(new_new_n10070__), .dinb(new_new_n10065__), .dout(new_new_n5419__));
  or1   g4478(.dina(new_new_n10071__), .dinb(new_new_n10067__), .dout(new_new_n5420__));
  and1  g4479(.dina(new_new_n5420__), .dinb(new_new_n5418__), .dout(new_new_n5421__));
  or1   g4480(.dina(new_new_n5419__), .dinb(new_new_n5417__), .dout(new_new_n5422__));
  and1  g4481(.dina(new_new_n8808__), .dinb(new_new_n8907__), .dout(new_new_n5423__));
  or1   g4482(.dina(new_new_n8809__), .dinb(new_new_n8921__), .dout(new_new_n5424__));
  and1  g4483(.dina(new_new_n10072__), .dinb(new_new_n10073__), .dout(new_new_n5425__));
  or1   g4484(.dina(new_new_n10074__), .dinb(new_new_n10075__), .dout(new_new_n5426__));
  and1  g4485(.dina(new_new_n10077__), .dinb(new_new_n10073__), .dout(new_new_n5427__));
  or1   g4486(.dina(new_new_n10078__), .dinb(new_new_n10075__), .dout(new_new_n5428__));
  and1  g4487(.dina(new_new_n10077__), .dinb(new_new_n10072__), .dout(new_new_n5429__));
  or1   g4488(.dina(new_new_n10078__), .dinb(new_new_n10074__), .dout(new_new_n5430__));
  and1  g4489(.dina(new_new_n5430__), .dinb(new_new_n5428__), .dout(new_new_n5431__));
  or1   g4490(.dina(new_new_n5429__), .dinb(new_new_n5427__), .dout(new_new_n5432__));
  and1  g4491(.dina(new_new_n9165__), .dinb(new_new_n9157__), .dout(new_new_n5433__));
  or1   g4492(.dina(new_new_n9167__), .dinb(new_new_n9159__), .dout(new_new_n5434__));
  or1   g4493(.dina(new_new_n5433__), .dinb(new_new_n5431__), .dout(new_new_n5435__));
  and1  g4494(.dina(new_new_n8978__), .dinb(new_new_n8974__), .dout(new_new_n5436__));
  or1   g4495(.dina(new_new_n8980__), .dinb(new_new_n8976__), .dout(new_new_n5437__));
  and1  g4496(.dina(new_new_n8977__), .dinb(new_new_n8973__), .dout(new_new_n5438__));
  or1   g4497(.dina(new_new_n8979__), .dinb(new_new_n8975__), .dout(new_new_n5439__));
  and1  g4498(.dina(new_new_n5439__), .dinb(new_new_n5437__), .dout(new_new_n5440__));
  or1   g4499(.dina(new_new_n5438__), .dinb(new_new_n5436__), .dout(new_new_n5441__));
  and1  g4500(.dina(new_new_n9481__), .dinb(new_new_n9473__), .dout(new_new_n5442__));
  or1   g4501(.dina(new_new_n9483__), .dinb(new_new_n9475__), .dout(new_new_n5443__));
  and1  g4502(.dina(new_new_n10079__), .dinb(new_new_n10080__), .dout(new_new_n5444__));
  or1   g4503(.dina(new_new_n10081__), .dinb(new_new_n10082__), .dout(new_new_n5445__));
  and1  g4504(.dina(new_new_n10084__), .dinb(new_new_n10080__), .dout(new_new_n5446__));
  or1   g4505(.dina(new_new_n10085__), .dinb(new_new_n10082__), .dout(new_new_n5447__));
  and1  g4506(.dina(new_new_n10084__), .dinb(new_new_n10079__), .dout(new_new_n5448__));
  or1   g4507(.dina(new_new_n10085__), .dinb(new_new_n10081__), .dout(new_new_n5449__));
  and1  g4508(.dina(new_new_n5449__), .dinb(new_new_n5447__), .dout(new_new_n5450__));
  or1   g4509(.dina(new_new_n5448__), .dinb(new_new_n5446__), .dout(new_new_n5451__));
  and1  g4510(.dina(new_new_n9441__), .dinb(new_new_n9557__), .dout(new_new_n5452__));
  or1   g4511(.dina(new_new_n9444__), .dinb(new_new_n9568__), .dout(new_new_n5453__));
  and1  g4512(.dina(new_new_n10086__), .dinb(new_new_n10087__), .dout(new_new_n5454__));
  or1   g4513(.dina(new_new_n10088__), .dinb(new_new_n10089__), .dout(new_new_n5455__));
  and1  g4514(.dina(new_new_n10091__), .dinb(new_new_n10087__), .dout(new_new_n5456__));
  or1   g4515(.dina(new_new_n10092__), .dinb(new_new_n10089__), .dout(new_new_n5457__));
  and1  g4516(.dina(new_new_n10091__), .dinb(new_new_n10086__), .dout(new_new_n5458__));
  or1   g4517(.dina(new_new_n10092__), .dinb(new_new_n10088__), .dout(new_new_n5459__));
  and1  g4518(.dina(new_new_n5459__), .dinb(new_new_n5457__), .dout(new_new_n5460__));
  or1   g4519(.dina(new_new_n5458__), .dinb(new_new_n5456__), .dout(new_new_n5461__));
  and1  g4520(.dina(new_new_n9574__), .dinb(new_new_n9548__), .dout(new_new_n5462__));
  or1   g4521(.dina(new_new_n9576__), .dinb(new_new_n9550__), .dout(new_new_n5463__));
  or1   g4522(.dina(new_new_n5462__), .dinb(new_new_n5460__), .dout(new_new_n5464__));
  and1  g4523(.dina(new_new_n9785__), .dinb(new_new_n9781__), .dout(new_new_n5465__));
  or1   g4524(.dina(new_new_n9787__), .dinb(new_new_n9783__), .dout(new_new_n5466__));
  and1  g4525(.dina(new_new_n9784__), .dinb(new_new_n9780__), .dout(new_new_n5467__));
  or1   g4526(.dina(new_new_n9786__), .dinb(new_new_n9782__), .dout(new_new_n5468__));
  and1  g4527(.dina(new_new_n5468__), .dinb(new_new_n5466__), .dout(new_new_n5469__));
  or1   g4528(.dina(new_new_n5467__), .dinb(new_new_n5465__), .dout(new_new_n5470__));
  and1  g4529(.dina(new_new_n9769__), .dinb(new_new_n9765__), .dout(new_new_n5471__));
  or1   g4530(.dina(new_new_n9771__), .dinb(new_new_n9767__), .dout(new_new_n5472__));
  and1  g4531(.dina(new_new_n9768__), .dinb(new_new_n9764__), .dout(new_new_n5473__));
  or1   g4532(.dina(new_new_n9770__), .dinb(new_new_n9766__), .dout(new_new_n5474__));
  and1  g4533(.dina(new_new_n5474__), .dinb(new_new_n5472__), .dout(new_new_n5475__));
  or1   g4534(.dina(new_new_n5473__), .dinb(new_new_n5471__), .dout(new_new_n5476__));
  and1  g4535(.dina(new_new_n9686__), .dinb(new_new_n9678__), .dout(new_new_n5477__));
  or1   g4536(.dina(new_new_n9688__), .dinb(new_new_n9680__), .dout(new_new_n5478__));
  and1  g4537(.dina(new_new_n10093__), .dinb(new_new_n10094__), .dout(new_new_n5479__));
  or1   g4538(.dina(new_new_n10095__), .dinb(new_new_n10096__), .dout(new_new_n5480__));
  and1  g4539(.dina(new_new_n10098__), .dinb(new_new_n10094__), .dout(new_new_n5481__));
  or1   g4540(.dina(new_new_n10100__), .dinb(new_new_n10096__), .dout(new_new_n5482__));
  and1  g4541(.dina(new_new_n10098__), .dinb(new_new_n10093__), .dout(new_new_n5483__));
  or1   g4542(.dina(new_new_n10100__), .dinb(new_new_n10095__), .dout(new_new_n5484__));
  and1  g4543(.dina(new_new_n5484__), .dinb(new_new_n5482__), .dout(new_new_n5485__));
  or1   g4544(.dina(new_new_n5483__), .dinb(new_new_n5481__), .dout(new_new_n5486__));
  and1  g4545(.dina(new_new_n7107__), .dinb(new_new_n8907__), .dout(new_new_n5487__));
  or1   g4546(.dina(new_new_n7111__), .dinb(new_new_n8920__), .dout(new_new_n5488__));
  and1  g4547(.dina(new_new_n10101__), .dinb(new_new_n10102__), .dout(new_new_n5489__));
  or1   g4548(.dina(new_new_n5487__), .dinb(new_new_n5485__), .dout(new_new_n5490__));
  and1  g4549(.dina(new_new_n10104__), .dinb(new_new_n10097__), .dout(new_new_n5491__));
  or1   g4550(.dina(new_new_n5489__), .dinb(new_new_n10099__), .dout(new_new_n5492__));
  or1   g4551(.dina(new_new_n5491__), .dinb(new_new_n5469__), .dout(new_new_n5493__));
  and1  g4552(.dina(new_new_n9849__), .dinb(new_new_n9845__), .dout(new_new_n5494__));
  or1   g4553(.dina(new_new_n9851__), .dinb(new_new_n9847__), .dout(new_new_n5495__));
  and1  g4554(.dina(new_new_n9848__), .dinb(new_new_n9844__), .dout(new_new_n5496__));
  or1   g4555(.dina(new_new_n9850__), .dinb(new_new_n9846__), .dout(new_new_n5497__));
  and1  g4556(.dina(new_new_n5497__), .dinb(new_new_n5495__), .dout(new_new_n5498__));
  or1   g4557(.dina(new_new_n5496__), .dinb(new_new_n5494__), .dout(new_new_n5499__));
  and1  g4558(.dina(new_new_n9833__), .dinb(new_new_n9829__), .dout(new_new_n5500__));
  or1   g4559(.dina(new_new_n9835__), .dinb(new_new_n9831__), .dout(new_new_n5501__));
  and1  g4560(.dina(new_new_n9832__), .dinb(new_new_n9828__), .dout(new_new_n5502__));
  or1   g4561(.dina(new_new_n9834__), .dinb(new_new_n9830__), .dout(new_new_n5503__));
  and1  g4562(.dina(new_new_n5503__), .dinb(new_new_n5501__), .dout(new_new_n5504__));
  or1   g4563(.dina(new_new_n5502__), .dinb(new_new_n5500__), .dout(new_new_n5505__));
  and1  g4564(.dina(new_new_n10006__), .dinb(new_new_n9998__), .dout(new_new_n5506__));
  or1   g4565(.dina(new_new_n10008__), .dinb(new_new_n10000__), .dout(new_new_n5507__));
  and1  g4566(.dina(new_new_n10105__), .dinb(new_new_n10106__), .dout(new_new_n5508__));
  or1   g4567(.dina(new_new_n10107__), .dinb(new_new_n10108__), .dout(new_new_n5509__));
  and1  g4568(.dina(new_new_n10110__), .dinb(new_new_n10106__), .dout(new_new_n5510__));
  or1   g4569(.dina(new_new_n10112__), .dinb(new_new_n10108__), .dout(new_new_n5511__));
  and1  g4570(.dina(new_new_n10110__), .dinb(new_new_n10105__), .dout(new_new_n5512__));
  or1   g4571(.dina(new_new_n10112__), .dinb(new_new_n10107__), .dout(new_new_n5513__));
  and1  g4572(.dina(new_new_n5513__), .dinb(new_new_n5511__), .dout(new_new_n5514__));
  or1   g4573(.dina(new_new_n5512__), .dinb(new_new_n5510__), .dout(new_new_n5515__));
  and1  g4574(.dina(new_new_n9195__), .dinb(new_new_n9559__), .dout(new_new_n5516__));
  or1   g4575(.dina(new_new_n9199__), .dinb(new_new_n9569__), .dout(new_new_n5517__));
  and1  g4576(.dina(new_new_n5517__), .dinb(new_new_n5515__), .dout(new_new_n5518__));
  or1   g4577(.dina(new_new_n10113__), .dinb(new_new_n10114__), .dout(new_new_n5519__));
  and1  g4578(.dina(new_new_n5519__), .dinb(new_new_n10109__), .dout(new_new_n5520__));
  or1   g4579(.dina(new_new_n10116__), .dinb(new_new_n10111__), .dout(new_new_n5521__));
  or1   g4580(.dina(new_new_n5520__), .dinb(new_new_n5498__), .dout(new_new_n5522__));
  and1  g4581(.dina(new_new_n10118__), .dinb(new_new_n4286__), .dout(new_new_n5523__));
  and1  g4582(.dina(new_new_n10118__), .dinb(new_new_n4288__), .dout(new_new_n5524__));
  or1   g4583(.dina(new_new_n5524__), .dinb(new_new_n5523__), .dout(new_new_n5525__));
  and1  g4584(.dina(new_new_n10120__), .dinb(new_new_n4295__), .dout(new_new_n5526__));
  and1  g4585(.dina(new_new_n10120__), .dinb(new_new_n4297__), .dout(new_new_n5527__));
  or1   g4586(.dina(new_new_n5527__), .dinb(new_new_n5526__), .dout(new_new_n5528__));
  and1  g4587(.dina(new_new_n10122__), .dinb(new_new_n4304__), .dout(new_new_n5529__));
  and1  g4588(.dina(new_new_n10122__), .dinb(new_new_n4306__), .dout(new_new_n5530__));
  or1   g4589(.dina(new_new_n5530__), .dinb(new_new_n5529__), .dout(new_new_n5531__));
  and1  g4590(.dina(new_new_n10124__), .dinb(new_new_n4313__), .dout(new_new_n5532__));
  and1  g4591(.dina(new_new_n10124__), .dinb(new_new_n4335__), .dout(new_new_n5533__));
  or1   g4592(.dina(new_new_n5533__), .dinb(new_new_n5532__), .dout(new_new_n5534__));
  and1  g4593(.dina(new_new_n9880__), .dinb(new_new_n9876__), .dout(new_new_n5535__));
  or1   g4594(.dina(new_new_n9881__), .dinb(new_new_n9878__), .dout(new_new_n5536__));
  and1  g4595(.dina(new_new_n5536__), .dinb(new_new_n10125__), .dout(new_new_n5537__));
  or1   g4596(.dina(new_new_n5535__), .dinb(new_new_n9882__), .dout(new_new_n5538__));
  and1  g4597(.dina(new_new_n9080__), .dinb(new_new_n9873__), .dout(new_new_n5539__));
  or1   g4598(.dina(new_new_n9095__), .dinb(new_new_n9875__), .dout(new_new_n5540__));
  and1  g4599(.dina(new_new_n9051__), .dinb(new_new_n10127__), .dout(new_new_n5541__));
  or1   g4600(.dina(new_new_n9068__), .dinb(new_new_n10129__), .dout(new_new_n5542__));
  and1  g4601(.dina(new_new_n10130__), .dinb(new_new_n10131__), .dout(new_new_n5543__));
  or1   g4602(.dina(new_new_n10132__), .dinb(new_new_n10133__), .dout(new_new_n5544__));
  and1  g4603(.dina(new_new_n10134__), .dinb(new_new_n10131__), .dout(new_new_n5545__));
  or1   g4604(.dina(new_new_n10135__), .dinb(new_new_n10133__), .dout(new_new_n5546__));
  or1   g4605(.dina(new_new_n10136__), .dinb(new_new_n5537__), .dout(new_new_n5547__));
  and1  g4606(.dina(new_new_n9965__), .dinb(new_new_n9961__), .dout(new_new_n5548__));
  or1   g4607(.dina(new_new_n9967__), .dinb(new_new_n9963__), .dout(new_new_n5549__));
  and1  g4608(.dina(new_new_n9964__), .dinb(new_new_n9960__), .dout(new_new_n5550__));
  or1   g4609(.dina(new_new_n9966__), .dinb(new_new_n9962__), .dout(new_new_n5551__));
  and1  g4610(.dina(new_new_n5551__), .dinb(new_new_n5549__), .dout(new_new_n5552__));
  or1   g4611(.dina(new_new_n5550__), .dinb(new_new_n5548__), .dout(new_new_n5553__));
  and1  g4612(.dina(new_new_n9948__), .dinb(new_new_n9944__), .dout(new_new_n5554__));
  or1   g4613(.dina(new_new_n9949__), .dinb(new_new_n9946__), .dout(new_new_n5555__));
  and1  g4614(.dina(new_new_n5555__), .dinb(new_new_n9950__), .dout(new_new_n5556__));
  or1   g4615(.dina(new_new_n5554__), .dinb(new_new_n9953__), .dout(new_new_n5557__));
  and1  g4616(.dina(new_new_n9080__), .dinb(new_new_n9940__), .dout(new_new_n5558__));
  or1   g4617(.dina(new_new_n9095__), .dinb(new_new_n9943__), .dout(new_new_n5559__));
  and1  g4618(.dina(new_new_n9054__), .dinb(new_new_n10139__), .dout(new_new_n5560__));
  or1   g4619(.dina(new_new_n9068__), .dinb(new_new_n10142__), .dout(new_new_n5561__));
  and1  g4620(.dina(new_new_n10143__), .dinb(new_new_n10144__), .dout(new_new_n5562__));
  or1   g4621(.dina(new_new_n10145__), .dinb(new_new_n10146__), .dout(new_new_n5563__));
  and1  g4622(.dina(new_new_n10147__), .dinb(new_new_n10144__), .dout(new_new_n5564__));
  or1   g4623(.dina(new_new_n10148__), .dinb(new_new_n10146__), .dout(new_new_n5565__));
  and1  g4624(.dina(new_new_n10150__), .dinb(new_new_n10151__), .dout(new_new_n5566__));
  or1   g4625(.dina(new_new_n10153__), .dinb(new_new_n10154__), .dout(new_new_n5567__));
  and1  g4626(.dina(new_new_n10156__), .dinb(new_new_n10151__), .dout(new_new_n5568__));
  or1   g4627(.dina(new_new_n10158__), .dinb(new_new_n10154__), .dout(new_new_n5569__));
  and1  g4628(.dina(new_new_n10156__), .dinb(new_new_n10150__), .dout(new_new_n5570__));
  or1   g4629(.dina(new_new_n10158__), .dinb(new_new_n10153__), .dout(new_new_n5571__));
  and1  g4630(.dina(new_new_n5571__), .dinb(new_new_n5569__), .dout(new_new_n5572__));
  or1   g4631(.dina(new_new_n5570__), .dinb(new_new_n5568__), .dout(new_new_n5573__));
  and1  g4632(.dina(new_new_n9022__), .dinb(new_new_n10139__), .dout(new_new_n5574__));
  or1   g4633(.dina(new_new_n9037__), .dinb(new_new_n10142__), .dout(new_new_n5575__));
  and1  g4634(.dina(new_new_n10159__), .dinb(new_new_n10160__), .dout(new_new_n5576__));
  or1   g4635(.dina(new_new_n10161__), .dinb(new_new_n10162__), .dout(new_new_n5577__));
  and1  g4636(.dina(new_new_n10164__), .dinb(new_new_n10155__), .dout(new_new_n5578__));
  or1   g4637(.dina(new_new_n10166__), .dinb(new_new_n10157__), .dout(new_new_n5579__));
  or1   g4638(.dina(new_new_n5578__), .dinb(new_new_n5552__), .dout(new_new_n5580__));
  or1   g4639(.dina(new_new_n10116__), .dinb(new_new_n10114__), .dout(new_new_n5581__));
  or1   g4640(.dina(new_new_n10115__), .dinb(new_new_n10113__), .dout(new_new_n5582__));
  and1  g4641(.dina(new_new_n5582__), .dinb(new_new_n5581__), .dout(new_new_n5583__));
  and1  g4642(.dina(new_new_n10104__), .dinb(new_new_n10102__), .dout(new_new_n5584__));
  and1  g4643(.dina(new_new_n10103__), .dinb(new_new_n10101__), .dout(new_new_n5585__));
  or1   g4644(.dina(new_new_n5585__), .dinb(new_new_n5584__), .dout(new_new_n5586__));
  and1  g4645(.dina(new_new_n10168__), .dinb(new_new_n4407__), .dout(new_new_n5587__));
  and1  g4646(.dina(new_new_n10168__), .dinb(new_new_n4409__), .dout(new_new_n5588__));
  or1   g4647(.dina(new_new_n5588__), .dinb(new_new_n5587__), .dout(new_new_n5589__));
  and1  g4648(.dina(new_new_n10170__), .dinb(new_new_n4580__), .dout(new_new_n5590__));
  and1  g4649(.dina(new_new_n10170__), .dinb(new_new_n4662__), .dout(new_new_n5591__));
  or1   g4650(.dina(new_new_n5591__), .dinb(new_new_n5590__), .dout(new_new_n5592__));
  and1  g4651(.dina(new_new_n10172__), .dinb(new_new_n4797__), .dout(new_new_n5593__));
  and1  g4652(.dina(new_new_n10172__), .dinb(new_new_n4881__), .dout(new_new_n5594__));
  or1   g4653(.dina(new_new_n5594__), .dinb(new_new_n5593__), .dout(new_new_n5595__));
  and1  g4654(.dina(new_new_n9083__), .dinb(new_new_n10174__), .dout(new_new_n5596__));
  or1   g4655(.dina(new_new_n9098__), .dinb(new_new_n10175__), .dout(new_new_n5597__));
  and1  g4656(.dina(new_new_n8795__), .dinb(new_new_n8906__), .dout(new_new_n5598__));
  and1  g4657(.dina(new_new_n9174__), .dinb(new_new_n10176__), .dout(new_new_n5599__));
  and1  g4658(.dina(new_new_n7707__), .dinb(new_new_n9559__), .dout(new_new_n5600__));
  or1   g4659(.dina(new_new_n10062__), .dinb(new_new_n9943__), .dout(new_new_n5601__));
  or1   g4660(.dina(new_new_n9037__), .dinb(new_new_n9874__), .dout(new_new_n5602__));
  and1  g4661(.dina(new_new_n10076__), .dinb(new_new_n10069__), .dout(new_new_n5603__));
  and1  g4662(.dina(new_new_n10090__), .dinb(new_new_n10083__), .dout(new_new_n5604__));
  and1  g4663(.dina(new_new_n10023__), .dinb(new_new_n10019__), .dout(new_new_n5605__));
  or1   g4664(.dina(new_new_n10025__), .dinb(new_new_n10021__), .dout(new_new_n5606__));
  and1  g4665(.dina(new_new_n10022__), .dinb(new_new_n10018__), .dout(new_new_n5607__));
  or1   g4666(.dina(new_new_n10024__), .dinb(new_new_n10020__), .dout(new_new_n5608__));
  and1  g4667(.dina(new_new_n5608__), .dinb(new_new_n5606__), .dout(new_new_n5609__));
  or1   g4668(.dina(new_new_n5607__), .dinb(new_new_n5605__), .dout(new_new_n5610__));
  and1  g4669(.dina(new_new_n9354__), .dinb(new_new_n9346__), .dout(new_new_n5611__));
  or1   g4670(.dina(new_new_n9356__), .dinb(new_new_n9348__), .dout(new_new_n5612__));
  and1  g4671(.dina(new_new_n10177__), .dinb(new_new_n10178__), .dout(new_new_n5613__));
  or1   g4672(.dina(new_new_n10179__), .dinb(new_new_n10180__), .dout(new_new_n5614__));
  and1  g4673(.dina(new_new_n10182__), .dinb(new_new_n10178__), .dout(new_new_n5615__));
  or1   g4674(.dina(new_new_n10183__), .dinb(new_new_n10180__), .dout(new_new_n5616__));
  and1  g4675(.dina(new_new_n10182__), .dinb(new_new_n10177__), .dout(new_new_n5617__));
  or1   g4676(.dina(new_new_n10183__), .dinb(new_new_n10179__), .dout(new_new_n5618__));
  and1  g4677(.dina(new_new_n5618__), .dinb(new_new_n5616__), .dout(new_new_n5619__));
  or1   g4678(.dina(new_new_n5617__), .dinb(new_new_n5615__), .dout(new_new_n5620__));
  and1  g4679(.dina(new_new_n9297__), .dinb(new_new_n9560__), .dout(new_new_n5621__));
  or1   g4680(.dina(new_new_n9301__), .dinb(new_new_n9569__), .dout(new_new_n5622__));
  or1   g4681(.dina(new_new_n5621__), .dinb(new_new_n5619__), .dout(new_new_n5623__));
  and1  g4682(.dina(new_new_n10185__), .dinb(new_new_n10181__), .dout(new_new_n5624__));
  and1  g4683(.dina(new_new_n9083__), .dinb(new_new_n10187__), .dout(new_new_n5625__));
  or1   g4684(.dina(new_new_n9098__), .dinb(new_new_n10188__), .dout(new_new_n5626__));
  and1  g4685(.dina(new_new_n9054__), .dinb(new_new_n10174__), .dout(new_new_n5627__));
  or1   g4686(.dina(new_new_n9069__), .dinb(new_new_n10175__), .dout(new_new_n5628__));
  and1  g4687(.dina(new_new_n5628__), .dinb(new_new_n5625__), .dout(new_new_n5629__));
  or1   g4688(.dina(new_new_n10189__), .dinb(new_new_n5626__), .dout(new_new_n5630__));
  and1  g4689(.dina(new_new_n9084__), .dinb(new_new_n10138__), .dout(new_new_n5631__));
  or1   g4690(.dina(new_new_n9099__), .dinb(new_new_n10141__), .dout(new_new_n5632__));
  and1  g4691(.dina(new_new_n9055__), .dinb(new_new_n10191__), .dout(new_new_n5633__));
  or1   g4692(.dina(new_new_n9069__), .dinb(new_new_n10194__), .dout(new_new_n5634__));
  and1  g4693(.dina(new_new_n10195__), .dinb(new_new_n10196__), .dout(new_new_n5635__));
  or1   g4694(.dina(new_new_n10197__), .dinb(new_new_n10198__), .dout(new_new_n5636__));
  and1  g4695(.dina(new_new_n10199__), .dinb(new_new_n10196__), .dout(new_new_n5637__));
  or1   g4696(.dina(new_new_n10200__), .dinb(new_new_n10198__), .dout(new_new_n5638__));
  and1  g4697(.dina(new_new_n10199__), .dinb(new_new_n10195__), .dout(new_new_n5639__));
  or1   g4698(.dina(new_new_n10200__), .dinb(new_new_n10197__), .dout(new_new_n5640__));
  and1  g4699(.dina(new_new_n5640__), .dinb(new_new_n10202__), .dout(new_new_n5641__));
  or1   g4700(.dina(new_new_n5639__), .dinb(new_new_n10204__), .dout(new_new_n5642__));
  and1  g4701(.dina(new_new_n9084__), .dinb(new_new_n10191__), .dout(new_new_n5643__));
  or1   g4702(.dina(new_new_n9099__), .dinb(new_new_n10194__), .dout(new_new_n5644__));
  and1  g4703(.dina(new_new_n9055__), .dinb(new_new_n9853__), .dout(new_new_n5645__));
  or1   g4704(.dina(new_new_n9071__), .dinb(new_new_n9856__), .dout(new_new_n5646__));
  and1  g4705(.dina(new_new_n10205__), .dinb(new_new_n10206__), .dout(new_new_n5647__));
  or1   g4706(.dina(new_new_n10207__), .dinb(new_new_n10208__), .dout(new_new_n5648__));
  and1  g4707(.dina(new_new_n10209__), .dinb(new_new_n10206__), .dout(new_new_n5649__));
  or1   g4708(.dina(new_new_n10210__), .dinb(new_new_n10208__), .dout(new_new_n5650__));
  and1  g4709(.dina(new_new_n10212__), .dinb(new_new_n10213__), .dout(new_new_n5651__));
  or1   g4710(.dina(new_new_n10215__), .dinb(new_new_n10216__), .dout(new_new_n5652__));
  and1  g4711(.dina(new_new_n10218__), .dinb(new_new_n10213__), .dout(new_new_n5653__));
  or1   g4712(.dina(new_new_n10219__), .dinb(new_new_n10216__), .dout(new_new_n5654__));
  and1  g4713(.dina(new_new_n10218__), .dinb(new_new_n10212__), .dout(new_new_n5655__));
  or1   g4714(.dina(new_new_n10219__), .dinb(new_new_n10215__), .dout(new_new_n5656__));
  and1  g4715(.dina(new_new_n5656__), .dinb(new_new_n5654__), .dout(new_new_n5657__));
  or1   g4716(.dina(new_new_n5655__), .dinb(new_new_n5653__), .dout(new_new_n5658__));
  and1  g4717(.dina(new_new_n9022__), .dinb(new_new_n9854__), .dout(new_new_n5659__));
  or1   g4718(.dina(new_new_n9038__), .dinb(new_new_n9855__), .dout(new_new_n5660__));
  or1   g4719(.dina(new_new_n5659__), .dinb(new_new_n5657__), .dout(new_new_n5661__));
  and1  g4720(.dina(new_new_n10221__), .dinb(new_new_n10217__), .dout(new_new_n5662__));
  and1  g4721(.dina(new_new_n9086__), .dinb(new_new_n9105__), .dout(new_new_n5663__));
  or1   g4722(.dina(new_new_n9101__), .dinb(new_new_n9108__), .dout(new_new_n5664__));
  and1  g4723(.dina(new_new_n9057__), .dinb(new_new_n10224__), .dout(new_new_n5665__));
  or1   g4724(.dina(new_new_n9071__), .dinb(new_new_n10227__), .dout(new_new_n5666__));
  and1  g4725(.dina(new_new_n10229__), .dinb(new_new_n10230__), .dout(new_new_n5667__));
  or1   g4726(.dina(new_new_n10231__), .dinb(new_new_n10232__), .dout(new_new_n5668__));
  and1  g4727(.dina(new_new_n10233__), .dinb(new_new_n10230__), .dout(new_new_n5669__));
  or1   g4728(.dina(new_new_n10234__), .dinb(new_new_n10232__), .dout(new_new_n5670__));
  and1  g4729(.dina(new_new_n10233__), .dinb(new_new_n10229__), .dout(new_new_n5671__));
  or1   g4730(.dina(new_new_n10234__), .dinb(new_new_n10231__), .dout(new_new_n5672__));
  and1  g4731(.dina(new_new_n5672__), .dinb(new_new_n10236__), .dout(new_new_n5673__));
  or1   g4732(.dina(new_new_n5671__), .dinb(new_new_n10238__), .dout(new_new_n5674__));
  and1  g4733(.dina(new_new_n9086__), .dinb(new_new_n10224__), .dout(new_new_n5675__));
  or1   g4734(.dina(new_new_n9101__), .dinb(new_new_n10227__), .dout(new_new_n5676__));
  and1  g4735(.dina(new_new_n9057__), .dinb(new_new_n9885__), .dout(new_new_n5677__));
  or1   g4736(.dina(new_new_n9072__), .dinb(new_new_n9888__), .dout(new_new_n5678__));
  and1  g4737(.dina(new_new_n10239__), .dinb(new_new_n10240__), .dout(new_new_n5679__));
  or1   g4738(.dina(new_new_n10241__), .dinb(new_new_n10242__), .dout(new_new_n5680__));
  and1  g4739(.dina(new_new_n10243__), .dinb(new_new_n10240__), .dout(new_new_n5681__));
  or1   g4740(.dina(new_new_n10244__), .dinb(new_new_n10242__), .dout(new_new_n5682__));
  and1  g4741(.dina(new_new_n10246__), .dinb(new_new_n10247__), .dout(new_new_n5683__));
  or1   g4742(.dina(new_new_n10249__), .dinb(new_new_n10250__), .dout(new_new_n5684__));
  and1  g4743(.dina(new_new_n10252__), .dinb(new_new_n10247__), .dout(new_new_n5685__));
  or1   g4744(.dina(new_new_n10254__), .dinb(new_new_n10250__), .dout(new_new_n5686__));
  and1  g4745(.dina(new_new_n10252__), .dinb(new_new_n10246__), .dout(new_new_n5687__));
  or1   g4746(.dina(new_new_n10254__), .dinb(new_new_n10249__), .dout(new_new_n5688__));
  and1  g4747(.dina(new_new_n5688__), .dinb(new_new_n5686__), .dout(new_new_n5689__));
  or1   g4748(.dina(new_new_n5687__), .dinb(new_new_n5685__), .dout(new_new_n5690__));
  and1  g4749(.dina(new_new_n9023__), .dinb(new_new_n9884__), .dout(new_new_n5691__));
  or1   g4750(.dina(new_new_n9038__), .dinb(new_new_n9889__), .dout(new_new_n5692__));
  and1  g4751(.dina(new_new_n10255__), .dinb(new_new_n10256__), .dout(new_new_n5693__));
  or1   g4752(.dina(new_new_n10257__), .dinb(new_new_n10258__), .dout(new_new_n5694__));
  and1  g4753(.dina(new_new_n10260__), .dinb(new_new_n10256__), .dout(new_new_n5695__));
  or1   g4754(.dina(new_new_n10262__), .dinb(new_new_n10258__), .dout(new_new_n5696__));
  and1  g4755(.dina(new_new_n10260__), .dinb(new_new_n10255__), .dout(new_new_n5697__));
  or1   g4756(.dina(new_new_n10262__), .dinb(new_new_n10257__), .dout(new_new_n5698__));
  and1  g4757(.dina(new_new_n5698__), .dinb(new_new_n5696__), .dout(new_new_n5699__));
  or1   g4758(.dina(new_new_n5697__), .dinb(new_new_n5695__), .dout(new_new_n5700__));
  and1  g4759(.dina(new_new_n10243__), .dinb(new_new_n10239__), .dout(new_new_n5701__));
  or1   g4760(.dina(new_new_n10244__), .dinb(new_new_n10241__), .dout(new_new_n5702__));
  and1  g4761(.dina(new_new_n5702__), .dinb(new_new_n10245__), .dout(new_new_n5703__));
  or1   g4762(.dina(new_new_n5701__), .dinb(new_new_n10248__), .dout(new_new_n5704__));
  and1  g4763(.dina(new_new_n10263__), .dinb(new_new_n9904__), .dout(new_new_n5705__));
  or1   g4764(.dina(new_new_n10264__), .dinb(new_new_n9906__), .dout(new_new_n5706__));
  and1  g4765(.dina(new_new_n10266__), .dinb(new_new_n10263__), .dout(new_new_n5707__));
  or1   g4766(.dina(new_new_n10268__), .dinb(new_new_n10264__), .dout(new_new_n5708__));
  and1  g4767(.dina(new_new_n10266__), .dinb(new_new_n9903__), .dout(new_new_n5709__));
  or1   g4768(.dina(new_new_n10268__), .dinb(new_new_n9905__), .dout(new_new_n5710__));
  and1  g4769(.dina(new_new_n5710__), .dinb(new_new_n5708__), .dout(new_new_n5711__));
  or1   g4770(.dina(new_new_n5709__), .dinb(new_new_n5707__), .dout(new_new_n5712__));
  and1  g4771(.dina(new_new_n9023__), .dinb(new_new_n9891__), .dout(new_new_n5713__));
  or1   g4772(.dina(new_new_n9040__), .dinb(new_new_n9896__), .dout(new_new_n5714__));
  and1  g4773(.dina(new_new_n10269__), .dinb(new_new_n10270__), .dout(new_new_n5715__));
  or1   g4774(.dina(new_new_n10271__), .dinb(new_new_n10272__), .dout(new_new_n5716__));
  and1  g4775(.dina(new_new_n10274__), .dinb(new_new_n10265__), .dout(new_new_n5717__));
  or1   g4776(.dina(new_new_n10276__), .dinb(new_new_n10267__), .dout(new_new_n5718__));
  and1  g4777(.dina(new_new_n10277__), .dinb(new_new_n10278__), .dout(new_new_n5719__));
  or1   g4778(.dina(new_new_n10279__), .dinb(new_new_n10280__), .dout(new_new_n5720__));
  and1  g4779(.dina(new_new_n10282__), .dinb(new_new_n10278__), .dout(new_new_n5721__));
  or1   g4780(.dina(new_new_n10283__), .dinb(new_new_n10280__), .dout(new_new_n5722__));
  and1  g4781(.dina(new_new_n10282__), .dinb(new_new_n10277__), .dout(new_new_n5723__));
  or1   g4782(.dina(new_new_n10283__), .dinb(new_new_n10279__), .dout(new_new_n5724__));
  and1  g4783(.dina(new_new_n5724__), .dinb(new_new_n5722__), .dout(new_new_n5725__));
  or1   g4784(.dina(new_new_n5723__), .dinb(new_new_n5721__), .dout(new_new_n5726__));
  and1  g4785(.dina(new_new_n10056__), .dinb(new_new_n9893__), .dout(new_new_n5727__));
  or1   g4786(.dina(new_new_n10063__), .dinb(new_new_n9896__), .dout(new_new_n5728__));
  or1   g4787(.dina(new_new_n5727__), .dinb(new_new_n5725__), .dout(new_new_n5729__));
  and1  g4788(.dina(new_new_n10285__), .dinb(new_new_n10281__), .dout(new_new_n5730__));
  and1  g4789(.dina(new_new_n10185__), .dinb(new_new_n5622__), .dout(new_new_n5731__));
  and1  g4790(.dina(new_new_n10287__), .dinb(new_new_n5434__), .dout(new_new_n5732__));
  and1  g4791(.dina(new_new_n10289__), .dinb(new_new_n5463__), .dout(new_new_n5733__));
  and1  g4792(.dina(new_new_n10291__), .dinb(new_new_n5492__), .dout(new_new_n5734__));
  and1  g4793(.dina(new_new_n10293__), .dinb(new_new_n5521__), .dout(new_new_n5735__));
  and1  g4794(.dina(new_new_n10287__), .dinb(new_new_n5432__), .dout(new_new_n5736__));
  and1  g4795(.dina(new_new_n10289__), .dinb(new_new_n5461__), .dout(new_new_n5737__));
  and1  g4796(.dina(new_new_n10293__), .dinb(new_new_n5499__), .dout(new_new_n5738__));
  and1  g4797(.dina(new_new_n10291__), .dinb(new_new_n5470__), .dout(new_new_n5739__));
  and1  g4798(.dina(new_new_n10184__), .dinb(new_new_n5620__), .dout(new_new_n5740__));
  and1  g4799(.dina(new_new_n10294__), .dinb(new_new_n10295__), .dout(new_new_n5741__));
  and1  g4800(.dina(new_new_n10296__), .dinb(new_new_n10297__), .dout(new_new_n5742__));
  and1  g4801(.dina(new_new_n10298__), .dinb(new_new_n10299__), .dout(new_new_n5743__));
  and1  g4802(.dina(new_new_n10300__), .dinb(new_new_n10301__), .dout(new_new_n5744__));
  and1  g4803(.dina(new_new_n10302__), .dinb(new_new_n10303__), .dout(new_new_n5745__));
  or1   g4804(.dina(new_new_n10304__), .dinb(new_new_n10305__), .dout(new_new_n5746__));
  and1  g4805(.dina(new_new_n10134__), .dinb(new_new_n10130__), .dout(new_new_n5747__));
  or1   g4806(.dina(new_new_n10135__), .dinb(new_new_n10132__), .dout(new_new_n5748__));
  and1  g4807(.dina(new_new_n5748__), .dinb(new_new_n10306__), .dout(new_new_n5749__));
  or1   g4808(.dina(new_new_n5747__), .dinb(new_new_n10136__), .dout(new_new_n5750__));
  and1  g4809(.dina(new_new_n9087__), .dinb(new_new_n10127__), .dout(new_new_n5751__));
  or1   g4810(.dina(new_new_n9100__), .dinb(new_new_n10129__), .dout(new_new_n5752__));
  and1  g4811(.dina(new_new_n9056__), .dinb(new_new_n10187__), .dout(new_new_n5753__));
  or1   g4812(.dina(new_new_n9072__), .dinb(new_new_n10188__), .dout(new_new_n5754__));
  and1  g4813(.dina(new_new_n10307__), .dinb(new_new_n10308__), .dout(new_new_n5755__));
  or1   g4814(.dina(new_new_n5753__), .dinb(new_new_n10309__), .dout(new_new_n5756__));
  and1  g4815(.dina(new_new_n10310__), .dinb(new_new_n10308__), .dout(new_new_n5757__));
  or1   g4816(.dina(new_new_n5755__), .dinb(new_new_n10309__), .dout(new_new_n5758__));
  or1   g4817(.dina(new_new_n10311__), .dinb(new_new_n5749__), .dout(new_new_n5759__));
  and1  g4818(.dina(new_new_n10164__), .dinb(new_new_n10160__), .dout(new_new_n5760__));
  or1   g4819(.dina(new_new_n10166__), .dinb(new_new_n10162__), .dout(new_new_n5761__));
  and1  g4820(.dina(new_new_n10163__), .dinb(new_new_n10159__), .dout(new_new_n5762__));
  or1   g4821(.dina(new_new_n10165__), .dinb(new_new_n10161__), .dout(new_new_n5763__));
  and1  g4822(.dina(new_new_n5763__), .dinb(new_new_n5761__), .dout(new_new_n5764__));
  or1   g4823(.dina(new_new_n5762__), .dinb(new_new_n5760__), .dout(new_new_n5765__));
  and1  g4824(.dina(new_new_n10147__), .dinb(new_new_n10143__), .dout(new_new_n5766__));
  or1   g4825(.dina(new_new_n10148__), .dinb(new_new_n10145__), .dout(new_new_n5767__));
  and1  g4826(.dina(new_new_n5767__), .dinb(new_new_n10149__), .dout(new_new_n5768__));
  or1   g4827(.dina(new_new_n5766__), .dinb(new_new_n10152__), .dout(new_new_n5769__));
  and1  g4828(.dina(new_new_n10312__), .dinb(new_new_n10202__), .dout(new_new_n5770__));
  or1   g4829(.dina(new_new_n10313__), .dinb(new_new_n10204__), .dout(new_new_n5771__));
  and1  g4830(.dina(new_new_n10315__), .dinb(new_new_n10312__), .dout(new_new_n5772__));
  or1   g4831(.dina(new_new_n10317__), .dinb(new_new_n10313__), .dout(new_new_n5773__));
  and1  g4832(.dina(new_new_n10315__), .dinb(new_new_n10201__), .dout(new_new_n5774__));
  or1   g4833(.dina(new_new_n10317__), .dinb(new_new_n10203__), .dout(new_new_n5775__));
  and1  g4834(.dina(new_new_n5775__), .dinb(new_new_n5773__), .dout(new_new_n5776__));
  or1   g4835(.dina(new_new_n5774__), .dinb(new_new_n5772__), .dout(new_new_n5777__));
  and1  g4836(.dina(new_new_n9026__), .dinb(new_new_n10192__), .dout(new_new_n5778__));
  or1   g4837(.dina(new_new_n9040__), .dinb(new_new_n10193__), .dout(new_new_n5779__));
  and1  g4838(.dina(new_new_n5779__), .dinb(new_new_n5777__), .dout(new_new_n5780__));
  or1   g4839(.dina(new_new_n10318__), .dinb(new_new_n10319__), .dout(new_new_n5781__));
  and1  g4840(.dina(new_new_n5781__), .dinb(new_new_n10314__), .dout(new_new_n5782__));
  or1   g4841(.dina(new_new_n10321__), .dinb(new_new_n10316__), .dout(new_new_n5783__));
  or1   g4842(.dina(new_new_n5782__), .dinb(new_new_n5764__), .dout(new_new_n5784__));
  and1  g4843(.dina(new_new_n9130__), .dinb(new_new_n9126__), .dout(new_new_n5785__));
  or1   g4844(.dina(new_new_n9132__), .dinb(new_new_n9128__), .dout(new_new_n5786__));
  and1  g4845(.dina(new_new_n9129__), .dinb(new_new_n9125__), .dout(new_new_n5787__));
  or1   g4846(.dina(new_new_n9131__), .dinb(new_new_n9127__), .dout(new_new_n5788__));
  and1  g4847(.dina(new_new_n5788__), .dinb(new_new_n5786__), .dout(new_new_n5789__));
  or1   g4848(.dina(new_new_n5787__), .dinb(new_new_n5785__), .dout(new_new_n5790__));
  and1  g4849(.dina(new_new_n9113__), .dinb(new_new_n9109__), .dout(new_new_n5791__));
  or1   g4850(.dina(new_new_n9114__), .dinb(new_new_n9111__), .dout(new_new_n5792__));
  and1  g4851(.dina(new_new_n5792__), .dinb(new_new_n9115__), .dout(new_new_n5793__));
  or1   g4852(.dina(new_new_n5791__), .dinb(new_new_n9118__), .dout(new_new_n5794__));
  and1  g4853(.dina(new_new_n10322__), .dinb(new_new_n10236__), .dout(new_new_n5795__));
  or1   g4854(.dina(new_new_n10323__), .dinb(new_new_n10238__), .dout(new_new_n5796__));
  and1  g4855(.dina(new_new_n10325__), .dinb(new_new_n10322__), .dout(new_new_n5797__));
  or1   g4856(.dina(new_new_n10327__), .dinb(new_new_n10323__), .dout(new_new_n5798__));
  and1  g4857(.dina(new_new_n10325__), .dinb(new_new_n10235__), .dout(new_new_n5799__));
  or1   g4858(.dina(new_new_n10327__), .dinb(new_new_n10237__), .dout(new_new_n5800__));
  and1  g4859(.dina(new_new_n5800__), .dinb(new_new_n5798__), .dout(new_new_n5801__));
  or1   g4860(.dina(new_new_n5799__), .dinb(new_new_n5797__), .dout(new_new_n5802__));
  and1  g4861(.dina(new_new_n9026__), .dinb(new_new_n10223__), .dout(new_new_n5803__));
  or1   g4862(.dina(new_new_n9041__), .dinb(new_new_n10228__), .dout(new_new_n5804__));
  and1  g4863(.dina(new_new_n10328__), .dinb(new_new_n10329__), .dout(new_new_n5805__));
  or1   g4864(.dina(new_new_n10330__), .dinb(new_new_n10331__), .dout(new_new_n5806__));
  and1  g4865(.dina(new_new_n10333__), .dinb(new_new_n10324__), .dout(new_new_n5807__));
  or1   g4866(.dina(new_new_n10335__), .dinb(new_new_n10326__), .dout(new_new_n5808__));
  and1  g4867(.dina(new_new_n10336__), .dinb(new_new_n10337__), .dout(new_new_n5809__));
  or1   g4868(.dina(new_new_n10338__), .dinb(new_new_n10339__), .dout(new_new_n5810__));
  and1  g4869(.dina(new_new_n10341__), .dinb(new_new_n10337__), .dout(new_new_n5811__));
  or1   g4870(.dina(new_new_n10342__), .dinb(new_new_n10339__), .dout(new_new_n5812__));
  and1  g4871(.dina(new_new_n10341__), .dinb(new_new_n10336__), .dout(new_new_n5813__));
  or1   g4872(.dina(new_new_n10342__), .dinb(new_new_n10338__), .dout(new_new_n5814__));
  and1  g4873(.dina(new_new_n5814__), .dinb(new_new_n5812__), .dout(new_new_n5815__));
  or1   g4874(.dina(new_new_n5813__), .dinb(new_new_n5811__), .dout(new_new_n5816__));
  and1  g4875(.dina(new_new_n10057__), .dinb(new_new_n10225__), .dout(new_new_n5817__));
  or1   g4876(.dina(new_new_n10063__), .dinb(new_new_n10228__), .dout(new_new_n5818__));
  and1  g4877(.dina(new_new_n10343__), .dinb(new_new_n10344__), .dout(new_new_n5819__));
  or1   g4878(.dina(new_new_n10345__), .dinb(new_new_n10346__), .dout(new_new_n5820__));
  and1  g4879(.dina(new_new_n10348__), .dinb(new_new_n10344__), .dout(new_new_n5821__));
  or1   g4880(.dina(new_new_n10349__), .dinb(new_new_n10346__), .dout(new_new_n5822__));
  and1  g4881(.dina(new_new_n10348__), .dinb(new_new_n10343__), .dout(new_new_n5823__));
  or1   g4882(.dina(new_new_n10349__), .dinb(new_new_n10345__), .dout(new_new_n5824__));
  and1  g4883(.dina(new_new_n5824__), .dinb(new_new_n5822__), .dout(new_new_n5825__));
  or1   g4884(.dina(new_new_n5823__), .dinb(new_new_n5821__), .dout(new_new_n5826__));
  and1  g4885(.dina(new_new_n10333__), .dinb(new_new_n10329__), .dout(new_new_n5827__));
  or1   g4886(.dina(new_new_n10335__), .dinb(new_new_n10331__), .dout(new_new_n5828__));
  and1  g4887(.dina(new_new_n10332__), .dinb(new_new_n10328__), .dout(new_new_n5829__));
  or1   g4888(.dina(new_new_n10334__), .dinb(new_new_n10330__), .dout(new_new_n5830__));
  and1  g4889(.dina(new_new_n5830__), .dinb(new_new_n5828__), .dout(new_new_n5831__));
  or1   g4890(.dina(new_new_n5829__), .dinb(new_new_n5827__), .dout(new_new_n5832__));
  and1  g4891(.dina(new_new_n10259__), .dinb(new_new_n10251__), .dout(new_new_n5833__));
  or1   g4892(.dina(new_new_n10261__), .dinb(new_new_n10253__), .dout(new_new_n5834__));
  and1  g4893(.dina(new_new_n10350__), .dinb(new_new_n10351__), .dout(new_new_n5835__));
  or1   g4894(.dina(new_new_n10352__), .dinb(new_new_n10353__), .dout(new_new_n5836__));
  and1  g4895(.dina(new_new_n10355__), .dinb(new_new_n10351__), .dout(new_new_n5837__));
  or1   g4896(.dina(new_new_n10357__), .dinb(new_new_n10353__), .dout(new_new_n5838__));
  and1  g4897(.dina(new_new_n10355__), .dinb(new_new_n10350__), .dout(new_new_n5839__));
  or1   g4898(.dina(new_new_n10357__), .dinb(new_new_n10352__), .dout(new_new_n5840__));
  and1  g4899(.dina(new_new_n5840__), .dinb(new_new_n5838__), .dout(new_new_n5841__));
  or1   g4900(.dina(new_new_n5839__), .dinb(new_new_n5837__), .dout(new_new_n5842__));
  and1  g4901(.dina(new_new_n10057__), .dinb(new_new_n9886__), .dout(new_new_n5843__));
  or1   g4902(.dina(new_new_n10064__), .dinb(new_new_n9889__), .dout(new_new_n5844__));
  and1  g4903(.dina(new_new_n5844__), .dinb(new_new_n5842__), .dout(new_new_n5845__));
  or1   g4904(.dina(new_new_n10358__), .dinb(new_new_n10359__), .dout(new_new_n5846__));
  and1  g4905(.dina(new_new_n5846__), .dinb(new_new_n10354__), .dout(new_new_n5847__));
  or1   g4906(.dina(new_new_n10361__), .dinb(new_new_n10356__), .dout(new_new_n5848__));
  or1   g4907(.dina(new_new_n5847__), .dinb(new_new_n5825__), .dout(new_new_n5849__));
  and1  g4908(.dina(new_new_n10363__), .dinb(new_new_n5051__), .dout(new_new_n5850__));
  and1  g4909(.dina(new_new_n10363__), .dinb(new_new_n5053__), .dout(new_new_n5851__));
  or1   g4910(.dina(new_new_n5851__), .dinb(new_new_n5850__), .dout(new_new_n5852__));
  and1  g4911(.dina(new_new_n10034__), .dinb(new_new_n5383__), .dout(new_new_n5853__));
  and1  g4912(.dina(new_new_n10033__), .dinb(new_new_n5385__), .dout(new_new_n5854__));
  or1   g4913(.dina(new_new_n5854__), .dinb(new_new_n5853__), .dout(new_new_n5855__));
  and1  g4914(.dina(new_new_n10365__), .dinb(new_new_n5061__), .dout(new_new_n5856__));
  and1  g4915(.dina(new_new_n10365__), .dinb(new_new_n5103__), .dout(new_new_n5857__));
  or1   g4916(.dina(new_new_n5857__), .dinb(new_new_n5856__), .dout(new_new_n5858__));
  and1  g4917(.dina(new_new_n10367__), .dinb(new_new_n5110__), .dout(new_new_n5859__));
  and1  g4918(.dina(new_new_n10367__), .dinb(new_new_n5192__), .dout(new_new_n5860__));
  or1   g4919(.dina(new_new_n5860__), .dinb(new_new_n5859__), .dout(new_new_n5861__));
  or1   g4920(.dina(new_new_n10361__), .dinb(new_new_n10359__), .dout(new_new_n5862__));
  or1   g4921(.dina(new_new_n10360__), .dinb(new_new_n10358__), .dout(new_new_n5863__));
  and1  g4922(.dina(new_new_n5863__), .dinb(new_new_n5862__), .dout(new_new_n5864__));
  and1  g4923(.dina(new_new_n10310__), .dinb(new_new_n10307__), .dout(new_new_n5865__));
  or1   g4924(.dina(new_new_n5865__), .dinb(new_new_n10311__), .dout(new_new_n5866__));
  or1   g4925(.dina(new_new_n10321__), .dinb(new_new_n10319__), .dout(new_new_n5867__));
  or1   g4926(.dina(new_new_n10320__), .dinb(new_new_n10318__), .dout(new_new_n5868__));
  and1  g4927(.dina(new_new_n5868__), .dinb(new_new_n5867__), .dout(new_new_n5869__));
  and1  g4928(.dina(new_new_n10369__), .dinb(new_new_n5205__), .dout(new_new_n5870__));
  and1  g4929(.dina(new_new_n10369__), .dinb(new_new_n10125__), .dout(new_new_n5871__));
  or1   g4930(.dina(new_new_n5871__), .dinb(new_new_n5870__), .dout(new_new_n5872__));
  and1  g4931(.dina(new_new_n10371__), .dinb(new_new_n5252__), .dout(new_new_n5873__));
  and1  g4932(.dina(new_new_n10371__), .dinb(new_new_n5278__), .dout(new_new_n5874__));
  or1   g4933(.dina(new_new_n5874__), .dinb(new_new_n5873__), .dout(new_new_n5875__));
  and1  g4934(.dina(new_new_n10059__), .dinb(new_new_n10140__), .dout(new_new_n5876__));
  and1  g4935(.dina(new_new_n9025__), .dinb(new_new_n10128__), .dout(new_new_n5877__));
  and1  g4936(.dina(new_new_n10347__), .dinb(new_new_n10340__), .dout(new_new_n5878__));
  or1   g4937(.dina(new_new_n10372__), .dinb(new_new_n5597__), .dout(new_new_n5879__));
  and1  g4938(.dina(new_new_n10209__), .dinb(new_new_n10205__), .dout(new_new_n5880__));
  or1   g4939(.dina(new_new_n10210__), .dinb(new_new_n10207__), .dout(new_new_n5881__));
  and1  g4940(.dina(new_new_n5881__), .dinb(new_new_n10211__), .dout(new_new_n5882__));
  or1   g4941(.dina(new_new_n5880__), .dinb(new_new_n10214__), .dout(new_new_n5883__));
  and1  g4942(.dina(new_new_n10373__), .dinb(new_new_n9869__), .dout(new_new_n5884__));
  or1   g4943(.dina(new_new_n10374__), .dinb(new_new_n9871__), .dout(new_new_n5885__));
  and1  g4944(.dina(new_new_n10376__), .dinb(new_new_n10373__), .dout(new_new_n5886__));
  or1   g4945(.dina(new_new_n10377__), .dinb(new_new_n10374__), .dout(new_new_n5887__));
  and1  g4946(.dina(new_new_n10376__), .dinb(new_new_n9868__), .dout(new_new_n5888__));
  or1   g4947(.dina(new_new_n10377__), .dinb(new_new_n9870__), .dout(new_new_n5889__));
  and1  g4948(.dina(new_new_n5889__), .dinb(new_new_n5887__), .dout(new_new_n5890__));
  or1   g4949(.dina(new_new_n5888__), .dinb(new_new_n5886__), .dout(new_new_n5891__));
  and1  g4950(.dina(new_new_n9027__), .dinb(new_new_n9859__), .dout(new_new_n5892__));
  or1   g4951(.dina(new_new_n9041__), .dinb(new_new_n9860__), .dout(new_new_n5893__));
  or1   g4952(.dina(new_new_n5892__), .dinb(new_new_n5890__), .dout(new_new_n5894__));
  and1  g4953(.dina(new_new_n10379__), .dinb(new_new_n10375__), .dout(new_new_n5895__));
  and1  g4954(.dina(new_new_n10274__), .dinb(new_new_n10270__), .dout(new_new_n5896__));
  or1   g4955(.dina(new_new_n10276__), .dinb(new_new_n10272__), .dout(new_new_n5897__));
  and1  g4956(.dina(new_new_n10273__), .dinb(new_new_n10269__), .dout(new_new_n5898__));
  or1   g4957(.dina(new_new_n10275__), .dinb(new_new_n10271__), .dout(new_new_n5899__));
  and1  g4958(.dina(new_new_n5899__), .dinb(new_new_n5897__), .dout(new_new_n5900__));
  or1   g4959(.dina(new_new_n5898__), .dinb(new_new_n5896__), .dout(new_new_n5901__));
  and1  g4960(.dina(new_new_n9934__), .dinb(new_new_n9926__), .dout(new_new_n5902__));
  or1   g4961(.dina(new_new_n9936__), .dinb(new_new_n9928__), .dout(new_new_n5903__));
  and1  g4962(.dina(new_new_n10380__), .dinb(new_new_n10381__), .dout(new_new_n5904__));
  or1   g4963(.dina(new_new_n10382__), .dinb(new_new_n10383__), .dout(new_new_n5905__));
  and1  g4964(.dina(new_new_n10385__), .dinb(new_new_n10381__), .dout(new_new_n5906__));
  or1   g4965(.dina(new_new_n10386__), .dinb(new_new_n10383__), .dout(new_new_n5907__));
  and1  g4966(.dina(new_new_n10385__), .dinb(new_new_n10380__), .dout(new_new_n5908__));
  or1   g4967(.dina(new_new_n10386__), .dinb(new_new_n10382__), .dout(new_new_n5909__));
  and1  g4968(.dina(new_new_n5909__), .dinb(new_new_n5907__), .dout(new_new_n5910__));
  or1   g4969(.dina(new_new_n5908__), .dinb(new_new_n5906__), .dout(new_new_n5911__));
  and1  g4970(.dina(new_new_n10059__), .dinb(new_new_n9910__), .dout(new_new_n5912__));
  or1   g4971(.dina(new_new_n10064__), .dinb(new_new_n9913__), .dout(new_new_n5913__));
  or1   g4972(.dina(new_new_n5912__), .dinb(new_new_n5910__), .dout(new_new_n5914__));
  and1  g4973(.dina(new_new_n10388__), .dinb(new_new_n10384__), .dout(new_new_n5915__));
  and1  g4974(.dina(new_new_n10388__), .dinb(new_new_n5913__), .dout(new_new_n5916__));
  and1  g4975(.dina(new_new_n10379__), .dinb(new_new_n5893__), .dout(new_new_n5917__));
  and1  g4976(.dina(new_new_n10390__), .dinb(new_new_n5758__), .dout(new_new_n5918__));
  and1  g4977(.dina(new_new_n10392__), .dinb(new_new_n5783__), .dout(new_new_n5919__));
  and1  g4978(.dina(new_new_n10394__), .dinb(new_new_n5848__), .dout(new_new_n5920__));
  and1  g4979(.dina(new_new_n10394__), .dinb(new_new_n5826__), .dout(new_new_n5921__));
  and1  g4980(.dina(new_new_n10390__), .dinb(new_new_n5750__), .dout(new_new_n5922__));
  and1  g4981(.dina(new_new_n10392__), .dinb(new_new_n5765__), .dout(new_new_n5923__));
  and1  g4982(.dina(new_new_n10378__), .dinb(new_new_n5891__), .dout(new_new_n5924__));
  and1  g4983(.dina(new_new_n10387__), .dinb(new_new_n5911__), .dout(new_new_n5925__));
  and1  g4984(.dina(new_new_n10395__), .dinb(new_new_n10396__), .dout(new_new_n5926__));
  and1  g4985(.dina(new_new_n10397__), .dinb(new_new_n10398__), .dout(new_new_n5927__));
  and1  g4986(.dina(new_new_n10399__), .dinb(new_new_n10401__), .dout(new_new_n5928__));
  or1   g4987(.dina(new_new_n10402__), .dinb(new_new_n10403__), .dout(new_new_n5929__));
  or1   g4988(.dina(new_new_n10404__), .dinb(new_new_n10405__), .dout(new_new_n5930__));
  and1  g4989(.dina(new_new_n10407__), .dinb(new_new_n5407__), .dout(new_new_n5931__));
  and1  g4990(.dina(new_new_n10407__), .dinb(new_new_n5409__), .dout(new_new_n5932__));
  or1   g4991(.dina(new_new_n5932__), .dinb(new_new_n5931__), .dout(new_new_n5933__));
  or1   g4992(.dina(new_new_n10189__), .dinb(new_new_n5627__), .dout(new_new_n5934__));
  and1  g4993(.dina(new_new_n5934__), .dinb(new_new_n10401__), .dout(new_new_n5935__));
  and1  g4994(.dina(new_new_n10285__), .dinb(new_new_n5726__), .dout(new_new_n5936__));
  and1  g4995(.dina(new_new_n10284__), .dinb(new_new_n5728__), .dout(new_new_n5937__));
  or1   g4996(.dina(new_new_n5937__), .dinb(new_new_n5936__), .dout(new_new_n5938__));
  and1  g4997(.dina(new_new_n10221__), .dinb(new_new_n5658__), .dout(new_new_n5939__));
  and1  g4998(.dina(new_new_n10220__), .dinb(new_new_n5660__), .dout(new_new_n5940__));
  or1   g4999(.dina(new_new_n5940__), .dinb(new_new_n5939__), .dout(new_new_n5941__));
  and1  g5000(.dina(new_new_n10409__), .dinb(new_new_n5538__), .dout(new_new_n5942__));
  and1  g5001(.dina(new_new_n10409__), .dinb(new_new_n10306__), .dout(new_new_n5943__));
  or1   g5002(.dina(new_new_n5943__), .dinb(new_new_n5942__), .dout(new_new_n5944__));
  and1  g5003(.dina(new_new_n10411__), .dinb(new_new_n5553__), .dout(new_new_n5945__));
  and1  g5004(.dina(new_new_n10411__), .dinb(new_new_n5579__), .dout(new_new_n5946__));
  or1   g5005(.dina(new_new_n5946__), .dinb(new_new_n5945__), .dout(new_new_n5947__));
  buf1  g5006(.din(new_new_n1617__), .dout(G6257));
  buf1  g5007(.din(new_new_n1620__), .dout(G6258));
  buf1  g5008(.din(new_new_n1623__), .dout(G6259));
  buf1  g5009(.din(new_new_n1626__), .dout(G6260));
  buf1  g5010(.din(new_new_n1629__), .dout(G6261));
  buf1  g5011(.din(new_new_n1632__), .dout(G6262));
  buf1  g5012(.din(new_new_n1635__), .dout(G6263));
  buf1  g5013(.din(new_new_n1638__), .dout(G6264));
  buf1  g5014(.din(new_new_n1641__), .dout(G6265));
  buf1  g5015(.din(new_new_n1644__), .dout(G6266));
  buf1  g5016(.din(new_new_n1647__), .dout(G6267));
  buf1  g5017(.din(new_new_n1650__), .dout(G6268));
  buf1  g5018(.din(new_new_n1653__), .dout(G6269));
  buf1  g5019(.din(new_new_n1656__), .dout(G6270));
  buf1  g5020(.din(new_new_n1659__), .dout(G6271));
  buf1  g5021(.din(new_new_n1662__), .dout(G6272));
  buf1  g5022(.din(new_new_n1664__), .dout(G6273));
  buf1  g5023(.din(new_new_n1667__), .dout(G6274));
  buf1  g5024(.din(new_new_n1670__), .dout(G6275));
  buf1  g5025(.din(new_new_n1679__), .dout(G6276));
  buf1  g5026(.din(new_new_n1694__), .dout(G6277));
  buf1  g5027(.din(new_new_n1717__), .dout(G6278));
  buf1  g5028(.din(new_new_n1746__), .dout(G6279));
  buf1  g5029(.din(new_new_n1781__), .dout(G6280));
  buf1  g5030(.din(new_new_n1824__), .dout(G6281));
  buf1  g5031(.din(new_new_n1873__), .dout(G6282));
  buf1  g5032(.din(new_new_n1928__), .dout(G6283));
  buf1  g5033(.din(new_new_n1991__), .dout(G6284));
  buf1  g5034(.din(new_new_n2050__), .dout(G6285));
  buf1  g5035(.din(new_new_n2089__), .dout(G6286));
  buf1  g5036(.din(new_new_n2105__), .dout(G6287));
  not1  g5037(.din(new_new_n2108__), .dout(G6288));
  buf1  g5038(.din(new_new_n6741__), .dout(n19409));
  buf1  g5039(.din(new_new_n7417__), .dout(n19412));
  buf1  g5040(.din(new_new_n7396__), .dout(n19415));
  buf1  g5041(.din(new_new_n7355__), .dout(n19418));
  buf1  g5042(.din(new_new_n7297__), .dout(n19421));
  buf1  g5043(.din(new_new_n7268__), .dout(n19424));
  buf1  g5044(.din(new_new_n7247__), .dout(n19427));
  buf1  g5045(.din(new_new_n7206__), .dout(n19430));
  buf1  g5046(.din(new_new_n7148__), .dout(n19433));
  buf1  g5047(.din(new_new_n7136__), .dout(n19436));
  buf1  g5048(.din(new_new_n999__), .dout(n19439));
  buf1  g5049(.din(new_new_n851__), .dout(n19442));
  buf1  g5050(.din(new_new_n853__), .dout(n19445));
  buf1  g5051(.din(new_new_n855__), .dout(n19448));
  buf1  g5052(.din(new_new_n857__), .dout(n19451));
  buf1  g5053(.din(new_new_n859__), .dout(n19454));
  buf1  g5054(.din(new_new_n903__), .dout(n19457));
  buf1  g5055(.din(new_new_n861__), .dout(n19460));
  buf1  g5056(.din(new_new_n907__), .dout(n19463));
  buf1  g5057(.din(new_new_n863__), .dout(n19466));
  buf1  g5058(.din(new_new_n911__), .dout(n19469));
  buf1  g5059(.din(new_new_n865__), .dout(n19472));
  buf1  g5060(.din(new_new_n915__), .dout(n19475));
  buf1  g5061(.din(new_new_n867__), .dout(n19478));
  buf1  g5062(.din(new_new_n919__), .dout(n19481));
  buf1  g5063(.din(new_new_n921__), .dout(n19484));
  buf1  g5064(.din(new_new_n6769__), .dout(n19487));
  buf1  g5065(.din(new_new_n869__), .dout(n19490));
  buf1  g5066(.din(new_new_n927__), .dout(n19493));
  buf1  g5067(.din(new_new_n929__), .dout(n19496));
  buf1  g5068(.din(new_new_n6813__), .dout(n19499));
  buf1  g5069(.din(new_new_n871__), .dout(n19502));
  buf1  g5070(.din(new_new_n935__), .dout(n19505));
  buf1  g5071(.din(new_new_n937__), .dout(n19508));
  buf1  g5072(.din(new_new_n6886__), .dout(n19511));
  buf1  g5073(.din(new_new_n1043__), .dout(n19514));
  buf1  g5074(.din(new_new_n1045__), .dout(n19517));
  buf1  g5075(.din(new_new_n1047__), .dout(n19520));
  buf1  g5076(.din(new_new_n1053__), .dout(n19523));
  buf1  g5077(.din(new_new_n1057__), .dout(n19526));
  buf1  g5078(.din(new_new_n1059__), .dout(n19529));
  buf1  g5079(.din(new_new_n1061__), .dout(n19532));
  buf1  g5080(.din(new_new_n1063__), .dout(n19535));
  buf1  g5081(.din(new_new_n1065__), .dout(n19538));
  buf1  g5082(.din(new_new_n1071__), .dout(n19541));
  buf1  g5083(.din(new_new_n1075__), .dout(n19544));
  buf1  g5084(.din(new_new_n1077__), .dout(n19547));
  buf1  g5085(.din(new_new_n1079__), .dout(n19550));
  buf1  g5086(.din(new_new_n1081__), .dout(n19553));
  buf1  g5087(.din(new_new_n1083__), .dout(n19556));
  buf1  g5088(.din(new_new_n1095__), .dout(n19559));
  buf1  g5089(.din(new_new_n1099__), .dout(n19562));
  buf1  g5090(.din(new_new_n1105__), .dout(n19565));
  buf1  g5091(.din(new_new_n1117__), .dout(n19568));
  buf1  g5092(.din(new_new_n1121__), .dout(n19571));
  buf1  g5093(.din(new_new_n1125__), .dout(n19574));
  buf1  g5094(.din(new_new_n1139__), .dout(n19577));
  buf1  g5095(.din(new_new_n1143__), .dout(n19580));
  buf1  g5096(.din(new_new_n1149__), .dout(n19583));
  buf1  g5097(.din(new_new_n1161__), .dout(n19586));
  buf1  g5098(.din(new_new_n1165__), .dout(n19589));
  buf1  g5099(.din(new_new_n1167__), .dout(n19592));
  buf1  g5100(.din(new_new_n7943__), .dout(n19595));
  buf1  g5101(.din(new_new_n1091__), .dout(n19598));
  buf1  g5102(.din(new_new_n1189__), .dout(n19601));
  buf1  g5103(.din(new_new_n7956__), .dout(n19604));
  buf1  g5104(.din(new_new_n1193__), .dout(n19607));
  buf1  g5105(.din(new_new_n7985__), .dout(n19610));
  buf1  g5106(.din(new_new_n8043__), .dout(n19613));
  buf1  g5107(.din(new_new_n1199__), .dout(n19616));
  buf1  g5108(.din(new_new_n8084__), .dout(n19619));
  buf1  g5109(.din(new_new_n8105__), .dout(n19622));
  buf1  g5110(.din(new_new_n8134__), .dout(n19625));
  buf1  g5111(.din(new_new_n8192__), .dout(n19628));
  buf1  g5112(.din(new_new_n8241__), .dout(n19631));
  buf1  g5113(.din(new_new_n8255__), .dout(n19634));
  buf1  g5114(.din(new_new_n8306__), .dout(n19637));
  buf1  g5115(.din(new_new_n1257__), .dout(n19640));
  buf1  g5116(.din(new_new_n8397__), .dout(n19643));
  buf1  g5117(.din(new_new_n1261__), .dout(n19646));
  buf1  g5118(.din(new_new_n8525__), .dout(n19649));
  buf1  g5119(.din(new_new_n7632__), .dout(n19652));
  buf1  g5120(.din(new_new_n1291__), .dout(n19655));
  buf1  g5121(.din(new_new_n6971__), .dout(n19658));
  buf1  g5122(.din(new_new_n6867__), .dout(n19661));
  buf1  g5123(.din(new_new_n1147__), .dout(n19664));
  buf1  g5124(.din(new_new_n1151__), .dout(n19667));
  buf1  g5125(.din(new_new_n1153__), .dout(n19670));
  buf1  g5126(.din(new_new_n6756__), .dout(n19673));
  buf1  g5127(.din(new_new_n6755__), .dout(n19676));
  buf1  g5128(.din(new_new_n1157__), .dout(n19679));
  buf1  g5129(.din(new_new_n6793__), .dout(n19682));
  buf1  g5130(.din(new_new_n1159__), .dout(n19685));
  buf1  g5131(.din(new_new_n1163__), .dout(n19688));
  buf1  g5132(.din(new_new_n1169__), .dout(n19691));
  buf1  g5133(.din(new_new_n1171__), .dout(n19694));
  buf1  g5134(.din(new_new_n1181__), .dout(n19697));
  buf1  g5135(.din(new_new_n6803__), .dout(n19700));
  buf1  g5136(.din(new_new_n6802__), .dout(n19703));
  buf1  g5137(.din(new_new_n1197__), .dout(n19706));
  buf1  g5138(.din(new_new_n6848__), .dout(n19709));
  buf1  g5139(.din(new_new_n1201__), .dout(n19712));
  buf1  g5140(.din(new_new_n1205__), .dout(n19715));
  buf1  g5141(.din(new_new_n1233__), .dout(n19718));
  buf1  g5142(.din(new_new_n1251__), .dout(n19721));
  buf1  g5143(.din(new_new_n1259__), .dout(n19724));
  buf1  g5144(.din(new_new_n6858__), .dout(n19727));
  buf1  g5145(.din(new_new_n6857__), .dout(n19730));
  buf1  g5146(.din(new_new_n8795__), .dout(n19733));
  buf1  g5147(.din(new_new_n1187__), .dout(n19736));
  buf1  g5148(.din(new_new_n8808__), .dout(n19739));
  buf1  g5149(.din(new_new_n1317__), .dout(n19742));
  buf1  g5150(.din(new_new_n6930__), .dout(n19745));
  buf1  g5151(.din(new_new_n1327__), .dout(n19748));
  buf1  g5152(.din(new_new_n8829__), .dout(n19751));
  buf1  g5153(.din(new_new_n8858__), .dout(n19754));
  buf1  g5154(.din(new_new_n1389__), .dout(n19757));
  buf1  g5155(.din(new_new_n8937__), .dout(n19760));
  buf1  g5156(.din(new_new_n9441__), .dout(n19763));
  buf1  g5157(.din(new_new_n9500__), .dout(n19766));
  buf1  g5158(.din(new_new_n9597__), .dout(n19769));
  buf1  g5159(.din(new_new_n9173__), .dout(n19772));
  buf1  g5160(.din(new_new_n6881__), .dout(n19775));
  buf1  g5161(.din(new_new_n9195__), .dout(n19778));
  buf1  g5162(.din(new_new_n6880__), .dout(n19781));
  buf1  g5163(.din(new_new_n9236__), .dout(n19784));
  buf1  g5164(.din(new_new_n6985__), .dout(n19787));
  buf1  g5165(.din(new_new_n9297__), .dout(n19790));
  buf1  g5166(.din(new_new_n9369__), .dout(n19793));
  buf1  g5167(.din(new_new_n7706__), .dout(n19796));
  buf1  g5168(.din(new_new_n6966__), .dout(n19799));
  buf1  g5169(.din(new_new_n6965__), .dout(n19802));
  buf1  g5170(.din(new_new_n7107__), .dout(n19805));
  buf1  g5171(.din(new_new_n6995__), .dout(n19808));
  buf1  g5172(.din(new_new_n7585__), .dout(n19811));
  buf1  g5173(.din(new_new_n6994__), .dout(n19814));
  buf1  g5174(.din(new_new_n6999__), .dout(n19817));
  buf1  g5175(.din(new_new_n1409__), .dout(n19820));
  buf1  g5176(.din(new_new_n7072__), .dout(n19823));
  buf1  g5177(.din(new_new_n1481__), .dout(n19826));
  buf1  g5178(.din(new_new_n1531__), .dout(n19829));
  buf1  g5179(.din(new_new_n7603__), .dout(n19832));
  buf1  g5180(.din(new_new_n7047__), .dout(n19835));
  buf1  g5181(.din(new_new_n7046__), .dout(n19838));
  buf1  g5182(.din(new_new_n7082__), .dout(n19841));
  buf1  g5183(.din(new_new_n7120__), .dout(n19844));
  buf1  g5184(.din(new_new_n7081__), .dout(n19847));
  buf1  g5185(.din(new_new_n7661__), .dout(n19850));
  buf1  g5186(.din(new_new_n7590__), .dout(n19853));
  buf1  g5187(.din(new_new_n7589__), .dout(n19856));
  buf1  g5188(.din(new_new_n7936__), .dout(n19859));
  buf1  g5189(.din(new_new_n7933__), .dout(n19862));
  buf1  g5190(.din(new_new_n7930__), .dout(n19865));
  buf1  g5191(.din(new_new_n7748__), .dout(n19868));
  buf1  g5192(.din(new_new_n7736__), .dout(n19871));
  buf1  g5193(.din(new_new_n8367__), .dout(n19874));
  buf1  g5194(.din(new_new_n9030__), .dout(n19877));
  buf1  g5195(.din(new_new_n9087__), .dout(n19880));
  buf1  g5196(.din(new_new_n7701__), .dout(n19883));
  buf1  g5197(.din(new_new_n7747__), .dout(n19886));
  buf1  g5198(.din(new_new_n7700__), .dout(n19889));
  buf1  g5199(.din(new_new_n9105__), .dout(n19892));
  buf1  g5200(.din(new_new_n7746__), .dout(n19895));
  buf1  g5201(.din(new_new_n8570__), .dout(n19898));
  buf1  g5202(.din(new_new_n7745__), .dout(n19901));
  buf1  g5203(.din(new_new_n10225__), .dout(n19904));
  buf1  g5204(.din(new_new_n8502__), .dout(n19907));
  buf1  g5205(.din(new_new_n9886__), .dout(n19910));
  buf1  g5206(.din(new_new_n9893__), .dout(n19913));
  not1  g5207(.din(new_new_n7940__), .dout(n19916));
  buf1  g5208(.din(new_new_n8622__), .dout(n19919));
  buf1  g5209(.din(new_new_n8624__), .dout(n19922));
  buf1  g5210(.din(new_new_n8626__), .dout(n19925));
  buf1  g5211(.din(new_new_n8628__), .dout(n19928));
  buf1  g5212(.din(new_new_n7939__), .dout(n19931));
  buf1  g5213(.din(new_new_n9910__), .dout(n19934));
  buf1  g5214(.din(new_new_n9940__), .dout(n19937));
  buf1  g5215(.din(new_new_n10140__), .dout(n19940));
  buf1  g5216(.din(new_new_n10192__), .dout(n19943));
  buf1  g5217(.din(new_new_n9027__), .dout(n19946));
  buf1  g5218(.din(new_new_n8512__), .dout(n19949));
  not1  g5219(.din(new_new_n9708__), .dout(n19952));
  not1  g5220(.din(new_new_n9710__), .dout(n19955));
  not1  g5221(.din(new_new_n9712__), .dout(n19958));
  buf1  g5222(.din(new_new_n8579__), .dout(n19961));
  buf1  g5223(.din(new_new_n8985__), .dout(n19964));
  buf1  g5224(.din(new_new_n8988__), .dout(n19967));
  buf1  g5225(.din(new_new_n8991__), .dout(n19970));
  buf1  g5226(.din(new_new_n9560__), .dout(n19973));
  buf1  g5227(.din(new_new_n8511__), .dout(n19976));
  buf1  g5228(.din(new_new_n9854__), .dout(n19979));
  buf1  g5229(.din(new_new_n8996__), .dout(n19982));
  buf1  g5230(.din(new_new_n8631__), .dout(n19985));
  buf1  g5231(.din(new_new_n9690__), .dout(n19988));
  buf1  g5232(.din(new_new_n8630__), .dout(n19991));
  buf1  g5233(.din(new_new_n9859__), .dout(n19994));
  buf1  g5234(.din(new_new_n9872__), .dout(n19997));
  buf1  g5235(.din(new_new_n10128__), .dout(n20000));
  not1  g5236(.din(new_new_n9701__), .dout(n20003));
  not1  g5237(.din(new_new_n9703__), .dout(n20006));
  not1  g5238(.din(new_new_n9705__), .dout(n20009));
  not1  g5239(.din(new_new_n9707__), .dout(n20012));
  buf1  g5240(.din(new_new_n9694__), .dout(n20015));
  buf1  g5241(.din(new_new_n9696__), .dout(n20018));
  buf1  g5242(.din(new_new_n9698__), .dout(n20021));
  buf1  g5243(.din(new_new_n9704__), .dout(n20024));
  buf1  g5244(.din(new_new_n9702__), .dout(n20027));
  buf1  g5245(.din(new_new_n9700__), .dout(n20030));
  buf1  g5246(.din(new_new_n9706__), .dout(n20033));
  buf1  g5247(.din(new_new_n9742__), .dout(n20036));
  buf1  g5248(.din(new_new_n9743__), .dout(n20039));
  buf1  g5249(.din(new_new_n9745__), .dout(n20042));
  buf1  g5250(.din(new_new_n9747__), .dout(n20045));
  buf1  g5251(.din(new_new_n9749__), .dout(n20048));
  buf1  g5252(.din(new_new_n9751__), .dout(n20051));
  buf1  g5253(.din(new_new_n10186__), .dout(n20054));
  not1  g5254(.din(new_new_n10117__), .dout(n20057));
  not1  g5255(.din(new_new_n10119__), .dout(n20060));
  not1  g5256(.din(new_new_n10121__), .dout(n20063));
  buf1  g5257(.din(new_new_n10123__), .dout(n20066));
  buf1  g5258(.din(new_new_n10173__), .dout(n20069));
  buf1  g5259(.din(new_new_n10058__), .dout(n20072));
  not1  g5260(.din(new_new_n9755__), .dout(n20075));
  buf1  g5261(.din(new_new_n10051__), .dout(n20078));
  buf1  g5262(.din(new_new_n10167__), .dout(n20081));
  buf1  g5263(.din(new_new_n10169__), .dout(n20084));
  buf1  g5264(.din(new_new_n10171__), .dout(n20087));
  buf1  g5265(.din(new_new_n9754__), .dout(n20090));
  not1  g5266(.din(new_new_n10044__), .dout(n20093));
  not1  g5267(.din(new_new_n10046__), .dout(n20096));
  not1  g5268(.din(new_new_n10048__), .dout(n20099));
  not1  g5269(.din(new_new_n10050__), .dout(n20102));
  buf1  g5270(.din(new_new_n4940__), .dout(n20105));
  buf1  g5271(.din(new_new_n4941__), .dout(n20108));
  buf1  g5272(.din(new_new_n4942__), .dout(n20111));
  buf1  g5273(.din(new_new_n4943__), .dout(n20114));
  buf1  g5274(.din(new_new_n4944__), .dout(n20117));
  buf1  g5275(.din(new_new_n4945__), .dout(n20120));
  buf1  g5276(.din(new_new_n4946__), .dout(n20123));
  buf1  g5277(.din(new_new_n4947__), .dout(n20126));
  buf1  g5278(.din(new_new_n4948__), .dout(n20129));
  buf1  g5279(.din(new_new_n4949__), .dout(n20132));
  buf1  g5280(.din(new_new_n4950__), .dout(n20135));
  buf1  g5281(.din(new_new_n4951__), .dout(n20138));
  buf1  g5282(.din(new_new_n4952__), .dout(n20141));
  not1  g5283(.din(new_new_n4955__), .dout(n20144));
  not1  g5284(.din(new_new_n4958__), .dout(n20147));
  not1  g5285(.din(new_new_n4961__), .dout(n20150));
  buf1  g5286(.din(new_new_n10035__), .dout(n20153));
  buf1  g5287(.din(new_new_n10037__), .dout(n20156));
  buf1  g5288(.din(new_new_n10039__), .dout(n20159));
  buf1  g5289(.din(new_new_n10041__), .dout(n20162));
  buf1  g5290(.din(new_new_n10043__), .dout(n20165));
  buf1  g5291(.din(new_new_n10045__), .dout(n20168));
  buf1  g5292(.din(new_new_n10047__), .dout(n20171));
  buf1  g5293(.din(new_new_n10049__), .dout(n20174));
  buf1  g5294(.din(new_new_n10176__), .dout(n20177));
  not1  g5295(.din(new_new_n10362__), .dout(n20180));
  buf1  g5296(.din(new_new_n9977__), .dout(n20183));
  buf1  g5297(.din(new_new_n10364__), .dout(n20186));
  buf1  g5298(.din(new_new_n10366__), .dout(n20189));
  buf1  g5299(.din(new_new_n10368__), .dout(n20192));
  buf1  g5300(.din(new_new_n10370__), .dout(n20195));
  buf1  g5301(.din(new_new_n809__), .dout(n20198));
  buf1  g5302(.din(new_new_n5280__), .dout(n20201));
  not1  g5303(.din(new_new_n10295__), .dout(n20204));
  not1  g5304(.din(new_new_n10297__), .dout(n20207));
  not1  g5305(.din(new_new_n10299__), .dout(n20210));
  not1  g5306(.din(new_new_n10301__), .dout(n20213));
  buf1  g5307(.din(new_new_n5285__), .dout(n20216));
  buf1  g5308(.din(new_new_n5286__), .dout(n20219));
  buf1  g5309(.din(new_new_n5306__), .dout(n20222));
  not1  g5310(.din(new_new_n10303__), .dout(n20225));
  buf1  g5311(.din(new_new_n10305__), .dout(n20228));
  buf1  g5312(.din(new_new_n5388__), .dout(n20231));
  not1  g5313(.din(new_new_n5389__), .dout(n20234));
  buf1  g5314(.din(new_new_n5390__), .dout(n20237));
  buf1  g5315(.din(new_new_n5391__), .dout(n20240));
  buf1  g5316(.din(new_new_n5392__), .dout(n20243));
  buf1  g5317(.din(new_new_n5393__), .dout(n20246));
  buf1  g5318(.din(new_new_n5394__), .dout(n20249));
  buf1  g5319(.din(new_new_n5395__), .dout(n20252));
  buf1  g5320(.din(new_new_n5396__), .dout(n20255));
  buf1  g5321(.din(new_new_n5397__), .dout(n20258));
  buf1  g5322(.din(new_new_n5398__), .dout(n20261));
  buf1  g5323(.din(new_new_n5399__), .dout(n20264));
  buf1  g5324(.din(new_new_n5400__), .dout(n20267));
  buf1  g5325(.din(new_new_n5401__), .dout(n20270));
  not1  g5326(.din(new_new_n10406__), .dout(n20273));
  buf1  g5327(.din(new_new_n10286__), .dout(n20276));
  buf1  g5328(.din(new_new_n10288__), .dout(n20279));
  buf1  g5329(.din(new_new_n10290__), .dout(n20282));
  buf1  g5330(.din(new_new_n10292__), .dout(n20285));
  not1  g5331(.din(new_new_n5525__), .dout(n20288));
  not1  g5332(.din(new_new_n5528__), .dout(n20291));
  not1  g5333(.din(new_new_n5531__), .dout(n20294));
  buf1  g5334(.din(new_new_n5534__), .dout(n20297));
  buf1  g5335(.din(new_new_n10408__), .dout(n20300));
  buf1  g5336(.din(new_new_n10410__), .dout(n20303));
  buf1  g5337(.din(new_new_n10304__), .dout(n20306));
  not1  g5338(.din(new_new_n10302__), .dout(n20309));
  buf1  g5339(.din(new_new_n10294__), .dout(n20312));
  buf1  g5340(.din(new_new_n10298__), .dout(n20315));
  buf1  g5341(.din(new_new_n10296__), .dout(n20318));
  buf1  g5342(.din(new_new_n10300__), .dout(n20321));
  buf1  g5343(.din(new_new_n5598__), .dout(n20324));
  buf1  g5344(.din(new_new_n5599__), .dout(n20327));
  buf1  g5345(.din(new_new_n5600__), .dout(n20330));
  not1  g5346(.din(new_new_n10396__), .dout(n20333));
  not1  g5347(.din(new_new_n10398__), .dout(n20336));
  buf1  g5348(.din(new_new_n5603__), .dout(n20339));
  buf1  g5349(.din(new_new_n5604__), .dout(n20342));
  buf1  g5350(.din(new_new_n5624__), .dout(n20345));
  not1  g5351(.din(new_new_n10400__), .dout(n20348));
  buf1  g5352(.din(new_new_n10403__), .dout(n20351));
  buf1  g5353(.din(new_new_n10405__), .dout(n20354));
  not1  g5354(.din(new_new_n5731__), .dout(n20357));
  buf1  g5355(.din(new_new_n5732__), .dout(n20360));
  buf1  g5356(.din(new_new_n5733__), .dout(n20363));
  buf1  g5357(.din(new_new_n5734__), .dout(n20366));
  buf1  g5358(.din(new_new_n5735__), .dout(n20369));
  buf1  g5359(.din(new_new_n5736__), .dout(n20372));
  buf1  g5360(.din(new_new_n5737__), .dout(n20375));
  buf1  g5361(.din(new_new_n5738__), .dout(n20378));
  buf1  g5362(.din(new_new_n5739__), .dout(n20381));
  buf1  g5363(.din(new_new_n5740__), .dout(n20384));
  buf1  g5364(.din(new_new_n5741__), .dout(n20387));
  buf1  g5365(.din(new_new_n5742__), .dout(n20390));
  buf1  g5366(.din(new_new_n5743__), .dout(n20393));
  buf1  g5367(.din(new_new_n10372__), .dout(n20396));
  not1  g5368(.din(new_new_n5745__), .dout(n20399));
  buf1  g5369(.din(new_new_n5746__), .dout(n20402));
  buf1  g5370(.din(new_new_n10389__), .dout(n20405));
  buf1  g5371(.din(new_new_n10391__), .dout(n20408));
  buf1  g5372(.din(new_new_n10393__), .dout(n20411));
  not1  g5373(.din(new_new_n5852__), .dout(n20414));
  not1  g5374(.din(new_new_n5855__), .dout(n20417));
  buf1  g5375(.din(new_new_n5858__), .dout(n20420));
  buf1  g5376(.din(new_new_n5861__), .dout(n20423));
  buf1  g5377(.din(new_new_n10404__), .dout(n20426));
  not1  g5378(.din(new_new_n10399__), .dout(n20429));
  buf1  g5379(.din(new_new_n10402__), .dout(n20432));
  buf1  g5380(.din(new_new_n10397__), .dout(n20435));
  buf1  g5381(.din(new_new_n10395__), .dout(n20438));
  buf1  g5382(.din(new_new_n5876__), .dout(n20441));
  buf1  g5383(.din(new_new_n5877__), .dout(n20444));
  buf1  g5384(.din(new_new_n5878__), .dout(n20447));
  not1  g5385(.din(new_new_n5879__), .dout(n20450));
  buf1  g5386(.din(new_new_n5895__), .dout(n20453));
  buf1  g5387(.din(new_new_n5915__), .dout(n20456));
  not1  g5388(.din(new_new_n5916__), .dout(n20459));
  not1  g5389(.din(new_new_n5917__), .dout(n20462));
  buf1  g5390(.din(new_new_n5918__), .dout(n20465));
  buf1  g5391(.din(new_new_n5919__), .dout(n20468));
  buf1  g5392(.din(new_new_n5920__), .dout(n20471));
  buf1  g5393(.din(new_new_n5921__), .dout(n20474));
  buf1  g5394(.din(new_new_n5922__), .dout(n20477));
  buf1  g5395(.din(new_new_n5923__), .dout(n20480));
  buf1  g5396(.din(new_new_n5924__), .dout(n20483));
  buf1  g5397(.din(new_new_n5925__), .dout(n20486));
  buf1  g5398(.din(new_new_n5926__), .dout(n20489));
  buf1  g5399(.din(new_new_n5927__), .dout(n20492));
  not1  g5400(.din(new_new_n5928__), .dout(n20495));
  buf1  g5401(.din(new_new_n5929__), .dout(n20498));
  buf1  g5402(.din(new_new_n5930__), .dout(n20501));
  not1  g5403(.din(new_new_n5933__), .dout(n20504));
  buf1  g5404(.din(new_new_n5935__), .dout(n20507));
  not1  g5405(.din(new_new_n5938__), .dout(n20510));
  not1  g5406(.din(new_new_n5941__), .dout(n20513));
  buf1  g5407(.din(new_new_n5944__), .dout(n20516));
  buf1  g5408(.din(new_new_n5947__), .dout(n20519));
  buf1  g5409(.din(new_new_n849__), .dout(n20522));
  buf1  g5410(.din(new_new_n947__), .dout(new_new_n6352__));
  buf1  g5411(.din(new_new_n953__), .dout(new_new_n6353__));
  buf1  g5412(.din(new_new_n959__), .dout(new_new_n6354__));
  buf1  g5413(.din(new_new_n965__), .dout(new_new_n6355__));
  buf1  g5414(.din(new_new_n971__), .dout(new_new_n6356__));
  buf1  g5415(.din(new_new_n977__), .dout(new_new_n6357__));
  buf1  g5416(.din(new_new_n983__), .dout(new_new_n6358__));
  buf1  g5417(.din(new_new_n989__), .dout(new_new_n6359__));
  buf1  g5418(.din(new_new_n995__), .dout(new_new_n6360__));
  buf1  g5419(.din(new_new_n1011__), .dout(new_new_n6361__));
  buf1  g5420(.din(new_new_n1037__), .dout(new_new_n6362__));
  buf1  g5421(.din(new_new_n1055__), .dout(new_new_n6363__));
  buf1  g5422(.din(new_new_n1073__), .dout(new_new_n6364__));
  buf1  g5423(.din(new_new_n1097__), .dout(new_new_n6365__));
  buf1  g5424(.din(new_new_n1141__), .dout(new_new_n6366__));
  buf1  g5425(.din(new_new_n1191__), .dout(new_new_n6367__));
  buf1  g5426(.din(new_new_n1241__), .dout(new_new_n6368__));
  buf1  g5427(.din(new_new_n1361__), .dout(new_new_n6369__));
  buf1  g5428(.din(new_new_n6369__), .dout(new_new_n6370__));
  buf1  g5429(.din(new_new_n1673__), .dout(new_new_n6371__));
  buf1  g5430(.din(new_new_n1671__), .dout(new_new_n6372__));
  buf1  g5431(.din(new_new_n1675__), .dout(new_new_n6373__));
  buf1  g5432(.din(new_new_n6373__), .dout(new_new_n6374__));
  buf1  g5433(.din(new_new_n1364__), .dout(new_new_n6375__));
  buf1  g5434(.din(new_new_n1342__), .dout(new_new_n6376__));
  buf1  g5435(.din(new_new_n1363__), .dout(new_new_n6377__));
  buf1  g5436(.din(new_new_n1341__), .dout(new_new_n6378__));
  buf1  g5437(.din(new_new_n1681__), .dout(new_new_n6379__));
  buf1  g5438(.din(new_new_n6379__), .dout(new_new_n6380__));
  buf1  g5439(.din(new_new_n1680__), .dout(new_new_n6381__));
  buf1  g5440(.din(new_new_n6381__), .dout(new_new_n6382__));
  buf1  g5441(.din(new_new_n1688__), .dout(new_new_n6383__));
  buf1  g5442(.din(new_new_n1686__), .dout(new_new_n6384__));
  buf1  g5443(.din(new_new_n1690__), .dout(new_new_n6385__));
  buf1  g5444(.din(new_new_n6385__), .dout(new_new_n6386__));
  buf1  g5445(.din(new_new_n1356__), .dout(new_new_n6387__));
  buf1  g5446(.din(new_new_n6387__), .dout(new_new_n6388__));
  buf1  g5447(.din(new_new_n1355__), .dout(new_new_n6389__));
  buf1  g5448(.din(new_new_n6389__), .dout(new_new_n6390__));
  buf1  g5449(.din(new_new_n1702__), .dout(new_new_n6391__));
  buf1  g5450(.din(new_new_n1700__), .dout(new_new_n6392__));
  buf1  g5451(.din(new_new_n1701__), .dout(new_new_n6393__));
  buf1  g5452(.din(new_new_n1699__), .dout(new_new_n6394__));
  buf1  g5453(.din(new_new_n1704__), .dout(new_new_n6395__));
  buf1  g5454(.din(new_new_n6395__), .dout(new_new_n6396__));
  buf1  g5455(.din(new_new_n1703__), .dout(new_new_n6397__));
  buf1  g5456(.din(new_new_n6397__), .dout(new_new_n6398__));
  buf1  g5457(.din(new_new_n1711__), .dout(new_new_n6399__));
  buf1  g5458(.din(new_new_n1709__), .dout(new_new_n6400__));
  buf1  g5459(.din(new_new_n1713__), .dout(new_new_n6401__));
  buf1  g5460(.din(new_new_n6401__), .dout(new_new_n6402__));
  buf1  g5461(.din(new_new_n941__), .dout(new_new_n6403__));
  buf1  g5462(.din(new_new_n6403__), .dout(new_new_n6404__));
  buf1  g5463(.din(new_new_n6404__), .dout(new_new_n6405__));
  buf1  g5464(.din(new_new_n6405__), .dout(new_new_n6406__));
  buf1  g5465(.din(new_new_n6404__), .dout(new_new_n6407__));
  buf1  g5466(.din(new_new_n6403__), .dout(new_new_n6408__));
  buf1  g5467(.din(new_new_n6408__), .dout(new_new_n6409__));
  buf1  g5468(.din(new_new_n6408__), .dout(new_new_n6410__));
  buf1  g5469(.din(new_new_n942__), .dout(new_new_n6411__));
  buf1  g5470(.din(new_new_n6411__), .dout(new_new_n6412__));
  buf1  g5471(.din(new_new_n6412__), .dout(new_new_n6413__));
  buf1  g5472(.din(new_new_n6413__), .dout(new_new_n6414__));
  buf1  g5473(.din(new_new_n6412__), .dout(new_new_n6415__));
  buf1  g5474(.din(new_new_n6411__), .dout(new_new_n6416__));
  buf1  g5475(.din(new_new_n6416__), .dout(new_new_n6417__));
  buf1  g5476(.din(new_new_n6416__), .dout(new_new_n6418__));
  buf1  g5477(.din(new_new_n1721__), .dout(new_new_n6419__));
  buf1  g5478(.din(new_new_n1719__), .dout(new_new_n6420__));
  buf1  g5479(.din(new_new_n1720__), .dout(new_new_n6421__));
  buf1  g5480(.din(new_new_n1718__), .dout(new_new_n6422__));
  buf1  g5481(.din(new_new_n1723__), .dout(new_new_n6423__));
  buf1  g5482(.din(new_new_n6423__), .dout(new_new_n6424__));
  buf1  g5483(.din(new_new_n1722__), .dout(new_new_n6425__));
  buf1  g5484(.din(new_new_n6425__), .dout(new_new_n6426__));
  buf1  g5485(.din(new_new_n1731__), .dout(new_new_n6427__));
  buf1  g5486(.din(new_new_n1729__), .dout(new_new_n6428__));
  buf1  g5487(.din(new_new_n1730__), .dout(new_new_n6429__));
  buf1  g5488(.din(new_new_n1728__), .dout(new_new_n6430__));
  buf1  g5489(.din(new_new_n1733__), .dout(new_new_n6431__));
  buf1  g5490(.din(new_new_n6431__), .dout(new_new_n6432__));
  buf1  g5491(.din(new_new_n1732__), .dout(new_new_n6433__));
  buf1  g5492(.din(new_new_n6433__), .dout(new_new_n6434__));
  buf1  g5493(.din(new_new_n1740__), .dout(new_new_n6435__));
  buf1  g5494(.din(new_new_n1738__), .dout(new_new_n6436__));
  buf1  g5495(.din(new_new_n1742__), .dout(new_new_n6437__));
  buf1  g5496(.din(new_new_n6437__), .dout(new_new_n6438__));
  buf1  g5497(.din(new_new_n1366__), .dout(new_new_n6439__));
  buf1  g5498(.din(new_new_n1340__), .dout(new_new_n6440__));
  buf1  g5499(.din(new_new_n1365__), .dout(new_new_n6441__));
  buf1  g5500(.din(new_new_n1339__), .dout(new_new_n6442__));
  buf1  g5501(.din(new_new_n1748__), .dout(new_new_n6443__));
  buf1  g5502(.din(new_new_n6443__), .dout(new_new_n6444__));
  buf1  g5503(.din(new_new_n1747__), .dout(new_new_n6445__));
  buf1  g5504(.din(new_new_n6445__), .dout(new_new_n6446__));
  buf1  g5505(.din(new_new_n1756__), .dout(new_new_n6447__));
  buf1  g5506(.din(new_new_n1754__), .dout(new_new_n6448__));
  buf1  g5507(.din(new_new_n1755__), .dout(new_new_n6449__));
  buf1  g5508(.din(new_new_n1753__), .dout(new_new_n6450__));
  buf1  g5509(.din(new_new_n1758__), .dout(new_new_n6451__));
  buf1  g5510(.din(new_new_n6451__), .dout(new_new_n6452__));
  buf1  g5511(.din(new_new_n1757__), .dout(new_new_n6453__));
  buf1  g5512(.din(new_new_n6453__), .dout(new_new_n6454__));
  buf1  g5513(.din(new_new_n1766__), .dout(new_new_n6455__));
  buf1  g5514(.din(new_new_n1764__), .dout(new_new_n6456__));
  buf1  g5515(.din(new_new_n1765__), .dout(new_new_n6457__));
  buf1  g5516(.din(new_new_n1763__), .dout(new_new_n6458__));
  buf1  g5517(.din(new_new_n1768__), .dout(new_new_n6459__));
  buf1  g5518(.din(new_new_n6459__), .dout(new_new_n6460__));
  buf1  g5519(.din(new_new_n1767__), .dout(new_new_n6461__));
  buf1  g5520(.din(new_new_n6461__), .dout(new_new_n6462__));
  buf1  g5521(.din(new_new_n1775__), .dout(new_new_n6463__));
  buf1  g5522(.din(new_new_n1773__), .dout(new_new_n6464__));
  buf1  g5523(.din(new_new_n1777__), .dout(new_new_n6465__));
  buf1  g5524(.din(new_new_n6465__), .dout(new_new_n6466__));
  buf1  g5525(.din(new_new_n1358__), .dout(new_new_n6467__));
  buf1  g5526(.din(new_new_n6467__), .dout(new_new_n6468__));
  buf1  g5527(.din(new_new_n1357__), .dout(new_new_n6469__));
  buf1  g5528(.din(new_new_n6469__), .dout(new_new_n6470__));
  buf1  g5529(.din(new_new_n1789__), .dout(new_new_n6471__));
  buf1  g5530(.din(new_new_n1787__), .dout(new_new_n6472__));
  buf1  g5531(.din(new_new_n1788__), .dout(new_new_n6473__));
  buf1  g5532(.din(new_new_n1786__), .dout(new_new_n6474__));
  buf1  g5533(.din(new_new_n1791__), .dout(new_new_n6475__));
  buf1  g5534(.din(new_new_n6475__), .dout(new_new_n6476__));
  buf1  g5535(.din(new_new_n1790__), .dout(new_new_n6477__));
  buf1  g5536(.din(new_new_n6477__), .dout(new_new_n6478__));
  buf1  g5537(.din(new_new_n1799__), .dout(new_new_n6479__));
  buf1  g5538(.din(new_new_n1797__), .dout(new_new_n6480__));
  buf1  g5539(.din(new_new_n1798__), .dout(new_new_n6481__));
  buf1  g5540(.din(new_new_n1796__), .dout(new_new_n6482__));
  buf1  g5541(.din(new_new_n1801__), .dout(new_new_n6483__));
  buf1  g5542(.din(new_new_n6483__), .dout(new_new_n6484__));
  buf1  g5543(.din(new_new_n1800__), .dout(new_new_n6485__));
  buf1  g5544(.din(new_new_n6485__), .dout(new_new_n6486__));
  buf1  g5545(.din(new_new_n1809__), .dout(new_new_n6487__));
  buf1  g5546(.din(new_new_n1807__), .dout(new_new_n6488__));
  buf1  g5547(.din(new_new_n1808__), .dout(new_new_n6489__));
  buf1  g5548(.din(new_new_n1806__), .dout(new_new_n6490__));
  buf1  g5549(.din(new_new_n1811__), .dout(new_new_n6491__));
  buf1  g5550(.din(new_new_n6491__), .dout(new_new_n6492__));
  buf1  g5551(.din(new_new_n1810__), .dout(new_new_n6493__));
  buf1  g5552(.din(new_new_n6493__), .dout(new_new_n6494__));
  buf1  g5553(.din(new_new_n1818__), .dout(new_new_n6495__));
  buf1  g5554(.din(new_new_n1816__), .dout(new_new_n6496__));
  buf1  g5555(.din(new_new_n1820__), .dout(new_new_n6497__));
  buf1  g5556(.din(new_new_n6497__), .dout(new_new_n6498__));
  buf1  g5557(.din(new_new_n933__), .dout(new_new_n6499__));
  buf1  g5558(.din(new_new_n6499__), .dout(new_new_n6500__));
  buf1  g5559(.din(new_new_n6500__), .dout(new_new_n6501__));
  buf1  g5560(.din(new_new_n6499__), .dout(new_new_n6502__));
  buf1  g5561(.din(new_new_n883__), .dout(new_new_n6503__));
  buf1  g5562(.din(new_new_n934__), .dout(new_new_n6504__));
  buf1  g5563(.din(new_new_n6504__), .dout(new_new_n6505__));
  buf1  g5564(.din(new_new_n6505__), .dout(new_new_n6506__));
  buf1  g5565(.din(new_new_n6504__), .dout(new_new_n6507__));
  buf1  g5566(.din(new_new_n884__), .dout(new_new_n6508__));
  buf1  g5567(.din(new_new_n1828__), .dout(new_new_n6509__));
  buf1  g5568(.din(new_new_n1826__), .dout(new_new_n6510__));
  buf1  g5569(.din(new_new_n1827__), .dout(new_new_n6511__));
  buf1  g5570(.din(new_new_n1825__), .dout(new_new_n6512__));
  buf1  g5571(.din(new_new_n1830__), .dout(new_new_n6513__));
  buf1  g5572(.din(new_new_n6513__), .dout(new_new_n6514__));
  buf1  g5573(.din(new_new_n1829__), .dout(new_new_n6515__));
  buf1  g5574(.din(new_new_n6515__), .dout(new_new_n6516__));
  buf1  g5575(.din(new_new_n1838__), .dout(new_new_n6517__));
  buf1  g5576(.din(new_new_n1836__), .dout(new_new_n6518__));
  buf1  g5577(.din(new_new_n1837__), .dout(new_new_n6519__));
  buf1  g5578(.din(new_new_n1835__), .dout(new_new_n6520__));
  buf1  g5579(.din(new_new_n1840__), .dout(new_new_n6521__));
  buf1  g5580(.din(new_new_n6521__), .dout(new_new_n6522__));
  buf1  g5581(.din(new_new_n1839__), .dout(new_new_n6523__));
  buf1  g5582(.din(new_new_n6523__), .dout(new_new_n6524__));
  buf1  g5583(.din(new_new_n1848__), .dout(new_new_n6525__));
  buf1  g5584(.din(new_new_n1846__), .dout(new_new_n6526__));
  buf1  g5585(.din(new_new_n1847__), .dout(new_new_n6527__));
  buf1  g5586(.din(new_new_n1845__), .dout(new_new_n6528__));
  buf1  g5587(.din(new_new_n1850__), .dout(new_new_n6529__));
  buf1  g5588(.din(new_new_n6529__), .dout(new_new_n6530__));
  buf1  g5589(.din(new_new_n1849__), .dout(new_new_n6531__));
  buf1  g5590(.din(new_new_n6531__), .dout(new_new_n6532__));
  buf1  g5591(.din(new_new_n1858__), .dout(new_new_n6533__));
  buf1  g5592(.din(new_new_n1856__), .dout(new_new_n6534__));
  buf1  g5593(.din(new_new_n1857__), .dout(new_new_n6535__));
  buf1  g5594(.din(new_new_n1855__), .dout(new_new_n6536__));
  buf1  g5595(.din(new_new_n1860__), .dout(new_new_n6537__));
  buf1  g5596(.din(new_new_n6537__), .dout(new_new_n6538__));
  buf1  g5597(.din(new_new_n1859__), .dout(new_new_n6539__));
  buf1  g5598(.din(new_new_n6539__), .dout(new_new_n6540__));
  buf1  g5599(.din(new_new_n1867__), .dout(new_new_n6541__));
  buf1  g5600(.din(new_new_n1865__), .dout(new_new_n6542__));
  buf1  g5601(.din(new_new_n1869__), .dout(new_new_n6543__));
  buf1  g5602(.din(new_new_n6543__), .dout(new_new_n6544__));
  buf1  g5603(.din(new_new_n1368__), .dout(new_new_n6545__));
  buf1  g5604(.din(new_new_n1338__), .dout(new_new_n6546__));
  buf1  g5605(.din(new_new_n1367__), .dout(new_new_n6547__));
  buf1  g5606(.din(new_new_n1337__), .dout(new_new_n6548__));
  buf1  g5607(.din(new_new_n1875__), .dout(new_new_n6549__));
  buf1  g5608(.din(new_new_n6549__), .dout(new_new_n6550__));
  buf1  g5609(.din(new_new_n1874__), .dout(new_new_n6551__));
  buf1  g5610(.din(new_new_n6551__), .dout(new_new_n6552__));
  buf1  g5611(.din(new_new_n885__), .dout(new_new_n6553__));
  buf1  g5612(.din(new_new_n886__), .dout(new_new_n6554__));
  buf1  g5613(.din(new_new_n1883__), .dout(new_new_n6555__));
  buf1  g5614(.din(new_new_n1881__), .dout(new_new_n6556__));
  buf1  g5615(.din(new_new_n1882__), .dout(new_new_n6557__));
  buf1  g5616(.din(new_new_n1880__), .dout(new_new_n6558__));
  buf1  g5617(.din(new_new_n1885__), .dout(new_new_n6559__));
  buf1  g5618(.din(new_new_n6559__), .dout(new_new_n6560__));
  buf1  g5619(.din(new_new_n1884__), .dout(new_new_n6561__));
  buf1  g5620(.din(new_new_n6561__), .dout(new_new_n6562__));
  buf1  g5621(.din(new_new_n1893__), .dout(new_new_n6563__));
  buf1  g5622(.din(new_new_n1891__), .dout(new_new_n6564__));
  buf1  g5623(.din(new_new_n1892__), .dout(new_new_n6565__));
  buf1  g5624(.din(new_new_n1890__), .dout(new_new_n6566__));
  buf1  g5625(.din(new_new_n1895__), .dout(new_new_n6567__));
  buf1  g5626(.din(new_new_n6567__), .dout(new_new_n6568__));
  buf1  g5627(.din(new_new_n1894__), .dout(new_new_n6569__));
  buf1  g5628(.din(new_new_n6569__), .dout(new_new_n6570__));
  buf1  g5629(.din(new_new_n1903__), .dout(new_new_n6571__));
  buf1  g5630(.din(new_new_n1901__), .dout(new_new_n6572__));
  buf1  g5631(.din(new_new_n1902__), .dout(new_new_n6573__));
  buf1  g5632(.din(new_new_n1900__), .dout(new_new_n6574__));
  buf1  g5633(.din(new_new_n1905__), .dout(new_new_n6575__));
  buf1  g5634(.din(new_new_n6575__), .dout(new_new_n6576__));
  buf1  g5635(.din(new_new_n1904__), .dout(new_new_n6577__));
  buf1  g5636(.din(new_new_n6577__), .dout(new_new_n6578__));
  buf1  g5637(.din(new_new_n1913__), .dout(new_new_n6579__));
  buf1  g5638(.din(new_new_n1911__), .dout(new_new_n6580__));
  buf1  g5639(.din(new_new_n1912__), .dout(new_new_n6581__));
  buf1  g5640(.din(new_new_n1910__), .dout(new_new_n6582__));
  buf1  g5641(.din(new_new_n1915__), .dout(new_new_n6583__));
  buf1  g5642(.din(new_new_n6583__), .dout(new_new_n6584__));
  buf1  g5643(.din(new_new_n1914__), .dout(new_new_n6585__));
  buf1  g5644(.din(new_new_n6585__), .dout(new_new_n6586__));
  buf1  g5645(.din(new_new_n1922__), .dout(new_new_n6587__));
  buf1  g5646(.din(new_new_n1920__), .dout(new_new_n6588__));
  buf1  g5647(.din(new_new_n1924__), .dout(new_new_n6589__));
  buf1  g5648(.din(new_new_n6589__), .dout(new_new_n6590__));
  buf1  g5649(.din(new_new_n1360__), .dout(new_new_n6591__));
  buf1  g5650(.din(new_new_n6591__), .dout(new_new_n6592__));
  buf1  g5651(.din(new_new_n1359__), .dout(new_new_n6593__));
  buf1  g5652(.din(new_new_n6593__), .dout(new_new_n6594__));
  buf1  g5653(.din(new_new_n1936__), .dout(new_new_n6595__));
  buf1  g5654(.din(new_new_n1934__), .dout(new_new_n6596__));
  buf1  g5655(.din(new_new_n1935__), .dout(new_new_n6597__));
  buf1  g5656(.din(new_new_n1933__), .dout(new_new_n6598__));
  buf1  g5657(.din(new_new_n1938__), .dout(new_new_n6599__));
  buf1  g5658(.din(new_new_n6599__), .dout(new_new_n6600__));
  buf1  g5659(.din(new_new_n1937__), .dout(new_new_n6601__));
  buf1  g5660(.din(new_new_n6601__), .dout(new_new_n6602__));
  buf1  g5661(.din(new_new_n887__), .dout(new_new_n6603__));
  buf1  g5662(.din(new_new_n888__), .dout(new_new_n6604__));
  buf1  g5663(.din(new_new_n1946__), .dout(new_new_n6605__));
  buf1  g5664(.din(new_new_n1944__), .dout(new_new_n6606__));
  buf1  g5665(.din(new_new_n1945__), .dout(new_new_n6607__));
  buf1  g5666(.din(new_new_n1943__), .dout(new_new_n6608__));
  buf1  g5667(.din(new_new_n1948__), .dout(new_new_n6609__));
  buf1  g5668(.din(new_new_n6609__), .dout(new_new_n6610__));
  buf1  g5669(.din(new_new_n1947__), .dout(new_new_n6611__));
  buf1  g5670(.din(new_new_n6611__), .dout(new_new_n6612__));
  buf1  g5671(.din(new_new_n1956__), .dout(new_new_n6613__));
  buf1  g5672(.din(new_new_n1954__), .dout(new_new_n6614__));
  buf1  g5673(.din(new_new_n1955__), .dout(new_new_n6615__));
  buf1  g5674(.din(new_new_n1953__), .dout(new_new_n6616__));
  buf1  g5675(.din(new_new_n1958__), .dout(new_new_n6617__));
  buf1  g5676(.din(new_new_n6617__), .dout(new_new_n6618__));
  buf1  g5677(.din(new_new_n1957__), .dout(new_new_n6619__));
  buf1  g5678(.din(new_new_n6619__), .dout(new_new_n6620__));
  buf1  g5679(.din(new_new_n1966__), .dout(new_new_n6621__));
  buf1  g5680(.din(new_new_n1964__), .dout(new_new_n6622__));
  buf1  g5681(.din(new_new_n1965__), .dout(new_new_n6623__));
  buf1  g5682(.din(new_new_n1963__), .dout(new_new_n6624__));
  buf1  g5683(.din(new_new_n1968__), .dout(new_new_n6625__));
  buf1  g5684(.din(new_new_n6625__), .dout(new_new_n6626__));
  buf1  g5685(.din(new_new_n1967__), .dout(new_new_n6627__));
  buf1  g5686(.din(new_new_n6627__), .dout(new_new_n6628__));
  buf1  g5687(.din(new_new_n1976__), .dout(new_new_n6629__));
  buf1  g5688(.din(new_new_n1974__), .dout(new_new_n6630__));
  buf1  g5689(.din(new_new_n1975__), .dout(new_new_n6631__));
  buf1  g5690(.din(new_new_n1973__), .dout(new_new_n6632__));
  buf1  g5691(.din(new_new_n1978__), .dout(new_new_n6633__));
  buf1  g5692(.din(new_new_n6633__), .dout(new_new_n6634__));
  buf1  g5693(.din(new_new_n1977__), .dout(new_new_n6635__));
  buf1  g5694(.din(new_new_n6635__), .dout(new_new_n6636__));
  buf1  g5695(.din(new_new_n1985__), .dout(new_new_n6637__));
  buf1  g5696(.din(new_new_n1983__), .dout(new_new_n6638__));
  buf1  g5697(.din(new_new_n1987__), .dout(new_new_n6639__));
  buf1  g5698(.din(new_new_n6639__), .dout(new_new_n6640__));
  buf1  g5699(.din(new_new_n891__), .dout(new_new_n6641__));
  buf1  g5700(.din(new_new_n6641__), .dout(new_new_n6642__));
  buf1  g5701(.din(new_new_n892__), .dout(new_new_n6643__));
  buf1  g5702(.din(new_new_n6643__), .dout(new_new_n6644__));
  buf1  g5703(.din(new_new_n1995__), .dout(new_new_n6645__));
  buf1  g5704(.din(new_new_n1993__), .dout(new_new_n6646__));
  buf1  g5705(.din(new_new_n1994__), .dout(new_new_n6647__));
  buf1  g5706(.din(new_new_n1992__), .dout(new_new_n6648__));
  buf1  g5707(.din(new_new_n1997__), .dout(new_new_n6649__));
  buf1  g5708(.din(new_new_n6649__), .dout(new_new_n6650__));
  buf1  g5709(.din(new_new_n1996__), .dout(new_new_n6651__));
  buf1  g5710(.din(new_new_n6651__), .dout(new_new_n6652__));
  buf1  g5711(.din(new_new_n889__), .dout(new_new_n6653__));
  buf1  g5712(.din(new_new_n890__), .dout(new_new_n6654__));
  buf1  g5713(.din(new_new_n2005__), .dout(new_new_n6655__));
  buf1  g5714(.din(new_new_n2003__), .dout(new_new_n6656__));
  buf1  g5715(.din(new_new_n2004__), .dout(new_new_n6657__));
  buf1  g5716(.din(new_new_n2002__), .dout(new_new_n6658__));
  buf1  g5717(.din(new_new_n2007__), .dout(new_new_n6659__));
  buf1  g5718(.din(new_new_n6659__), .dout(new_new_n6660__));
  buf1  g5719(.din(new_new_n2006__), .dout(new_new_n6661__));
  buf1  g5720(.din(new_new_n6661__), .dout(new_new_n6662__));
  buf1  g5721(.din(new_new_n2015__), .dout(new_new_n6663__));
  buf1  g5722(.din(new_new_n2013__), .dout(new_new_n6664__));
  buf1  g5723(.din(new_new_n2014__), .dout(new_new_n6665__));
  buf1  g5724(.din(new_new_n2012__), .dout(new_new_n6666__));
  buf1  g5725(.din(new_new_n2017__), .dout(new_new_n6667__));
  buf1  g5726(.din(new_new_n6667__), .dout(new_new_n6668__));
  buf1  g5727(.din(new_new_n2016__), .dout(new_new_n6669__));
  buf1  g5728(.din(new_new_n6669__), .dout(new_new_n6670__));
  buf1  g5729(.din(new_new_n2025__), .dout(new_new_n6671__));
  buf1  g5730(.din(new_new_n2023__), .dout(new_new_n6672__));
  buf1  g5731(.din(new_new_n2024__), .dout(new_new_n6673__));
  buf1  g5732(.din(new_new_n2022__), .dout(new_new_n6674__));
  buf1  g5733(.din(new_new_n2027__), .dout(new_new_n6675__));
  buf1  g5734(.din(new_new_n6675__), .dout(new_new_n6676__));
  buf1  g5735(.din(new_new_n2026__), .dout(new_new_n6677__));
  buf1  g5736(.din(new_new_n6677__), .dout(new_new_n6678__));
  buf1  g5737(.din(new_new_n2035__), .dout(new_new_n6679__));
  buf1  g5738(.din(new_new_n2033__), .dout(new_new_n6680__));
  buf1  g5739(.din(new_new_n2034__), .dout(new_new_n6681__));
  buf1  g5740(.din(new_new_n2032__), .dout(new_new_n6682__));
  buf1  g5741(.din(new_new_n2037__), .dout(new_new_n6683__));
  buf1  g5742(.din(new_new_n6683__), .dout(new_new_n6684__));
  buf1  g5743(.din(new_new_n2036__), .dout(new_new_n6685__));
  buf1  g5744(.din(new_new_n6685__), .dout(new_new_n6686__));
  buf1  g5745(.din(new_new_n2044__), .dout(new_new_n6687__));
  buf1  g5746(.din(new_new_n2042__), .dout(new_new_n6688__));
  buf1  g5747(.din(new_new_n2046__), .dout(new_new_n6689__));
  buf1  g5748(.din(new_new_n6689__), .dout(new_new_n6690__));
  buf1  g5749(.din(new_new_n2054__), .dout(new_new_n6691__));
  buf1  g5750(.din(new_new_n2052__), .dout(new_new_n6692__));
  buf1  g5751(.din(new_new_n2053__), .dout(new_new_n6693__));
  buf1  g5752(.din(new_new_n2051__), .dout(new_new_n6694__));
  buf1  g5753(.din(new_new_n2056__), .dout(new_new_n6695__));
  buf1  g5754(.din(new_new_n6695__), .dout(new_new_n6696__));
  buf1  g5755(.din(new_new_n2055__), .dout(new_new_n6697__));
  buf1  g5756(.din(new_new_n6697__), .dout(new_new_n6698__));
  buf1  g5757(.din(new_new_n2064__), .dout(new_new_n6699__));
  buf1  g5758(.din(new_new_n2062__), .dout(new_new_n6700__));
  buf1  g5759(.din(new_new_n2063__), .dout(new_new_n6701__));
  buf1  g5760(.din(new_new_n2061__), .dout(new_new_n6702__));
  buf1  g5761(.din(new_new_n2066__), .dout(new_new_n6703__));
  buf1  g5762(.din(new_new_n6703__), .dout(new_new_n6704__));
  buf1  g5763(.din(new_new_n2065__), .dout(new_new_n6705__));
  buf1  g5764(.din(new_new_n6705__), .dout(new_new_n6706__));
  buf1  g5765(.din(new_new_n2074__), .dout(new_new_n6707__));
  buf1  g5766(.din(new_new_n2072__), .dout(new_new_n6708__));
  buf1  g5767(.din(new_new_n2073__), .dout(new_new_n6709__));
  buf1  g5768(.din(new_new_n2071__), .dout(new_new_n6710__));
  buf1  g5769(.din(new_new_n2076__), .dout(new_new_n6711__));
  buf1  g5770(.din(new_new_n6711__), .dout(new_new_n6712__));
  buf1  g5771(.din(new_new_n2075__), .dout(new_new_n6713__));
  buf1  g5772(.din(new_new_n6713__), .dout(new_new_n6714__));
  buf1  g5773(.din(new_new_n2083__), .dout(new_new_n6715__));
  buf1  g5774(.din(new_new_n2081__), .dout(new_new_n6716__));
  buf1  g5775(.din(new_new_n2085__), .dout(new_new_n6717__));
  buf1  g5776(.din(new_new_n6717__), .dout(new_new_n6718__));
  buf1  g5777(.din(new_new_n2093__), .dout(new_new_n6719__));
  buf1  g5778(.din(new_new_n2091__), .dout(new_new_n6720__));
  buf1  g5779(.din(new_new_n2092__), .dout(new_new_n6721__));
  buf1  g5780(.din(new_new_n2090__), .dout(new_new_n6722__));
  buf1  g5781(.din(new_new_n2095__), .dout(new_new_n6723__));
  buf1  g5782(.din(new_new_n6723__), .dout(new_new_n6724__));
  buf1  g5783(.din(new_new_n2094__), .dout(new_new_n6725__));
  buf1  g5784(.din(new_new_n2104__), .dout(new_new_n6726__));
  buf1  g5785(.din(new_new_n6726__), .dout(new_new_n6727__));
  buf1  g5786(.din(new_new_n1255__), .dout(new_new_n6728__));
  buf1  g5787(.din(new_new_n6728__), .dout(new_new_n6729__));
  buf1  g5788(.din(new_new_n6729__), .dout(new_new_n6730__));
  buf1  g5789(.din(new_new_n6730__), .dout(new_new_n6731__));
  buf1  g5790(.din(new_new_n6730__), .dout(new_new_n6732__));
  buf1  g5791(.din(new_new_n6729__), .dout(new_new_n6733__));
  buf1  g5792(.din(new_new_n6733__), .dout(new_new_n6734__));
  buf1  g5793(.din(new_new_n6728__), .dout(new_new_n6735__));
  buf1  g5794(.din(new_new_n6735__), .dout(new_new_n6736__));
  buf1  g5795(.din(new_new_n6735__), .dout(new_new_n6737__));
  buf1  g5796(.din(new_new_n1041__), .dout(new_new_n6738__));
  buf1  g5797(.din(new_new_n6738__), .dout(new_new_n6739__));
  buf1  g5798(.din(new_new_n6739__), .dout(new_new_n6740__));
  buf1  g5799(.din(new_new_n6738__), .dout(new_new_n6741__));
  buf1  g5800(.din(new_new_n1256__), .dout(new_new_n6742__));
  buf1  g5801(.din(new_new_n6742__), .dout(new_new_n6743__));
  buf1  g5802(.din(new_new_n6743__), .dout(new_new_n6744__));
  buf1  g5803(.din(new_new_n6744__), .dout(new_new_n6745__));
  buf1  g5804(.din(new_new_n6744__), .dout(new_new_n6746__));
  buf1  g5805(.din(new_new_n6743__), .dout(new_new_n6747__));
  buf1  g5806(.din(new_new_n6747__), .dout(new_new_n6748__));
  buf1  g5807(.din(new_new_n6742__), .dout(new_new_n6749__));
  buf1  g5808(.din(new_new_n6749__), .dout(new_new_n6750__));
  buf1  g5809(.din(new_new_n6749__), .dout(new_new_n6751__));
  buf1  g5810(.din(new_new_n1042__), .dout(new_new_n6752__));
  buf1  g5811(.din(new_new_n6752__), .dout(new_new_n6753__));
  buf1  g5812(.din(new_new_n6752__), .dout(new_new_n6754__));
  buf1  g5813(.din(new_new_n2112__), .dout(new_new_n6755__));
  buf1  g5814(.din(new_new_n2109__), .dout(new_new_n6756__));
  buf1  g5815(.din(new_new_n923__), .dout(new_new_n6757__));
  buf1  g5816(.din(new_new_n6757__), .dout(new_new_n6758__));
  buf1  g5817(.din(new_new_n6758__), .dout(new_new_n6759__));
  buf1  g5818(.din(new_new_n6759__), .dout(new_new_n6760__));
  buf1  g5819(.din(new_new_n6759__), .dout(new_new_n6761__));
  buf1  g5820(.din(new_new_n6758__), .dout(new_new_n6762__));
  buf1  g5821(.din(new_new_n6762__), .dout(new_new_n6763__));
  buf1  g5822(.din(new_new_n6762__), .dout(new_new_n6764__));
  buf1  g5823(.din(new_new_n6757__), .dout(new_new_n6765__));
  buf1  g5824(.din(new_new_n6765__), .dout(new_new_n6766__));
  buf1  g5825(.din(new_new_n6766__), .dout(new_new_n6767__));
  buf1  g5826(.din(new_new_n6766__), .dout(new_new_n6768__));
  buf1  g5827(.din(new_new_n6765__), .dout(new_new_n6769__));
  buf1  g5828(.din(new_new_n6769__), .dout(new_new_n6770__));
  buf1  g5829(.din(new_new_n924__), .dout(new_new_n6771__));
  buf1  g5830(.din(new_new_n6771__), .dout(new_new_n6772__));
  buf1  g5831(.din(new_new_n6772__), .dout(new_new_n6773__));
  buf1  g5832(.din(new_new_n6773__), .dout(new_new_n6774__));
  buf1  g5833(.din(new_new_n6773__), .dout(new_new_n6775__));
  buf1  g5834(.din(new_new_n6772__), .dout(new_new_n6776__));
  buf1  g5835(.din(new_new_n6776__), .dout(new_new_n6777__));
  buf1  g5836(.din(new_new_n6776__), .dout(new_new_n6778__));
  buf1  g5837(.din(new_new_n6771__), .dout(new_new_n6779__));
  buf1  g5838(.din(new_new_n6779__), .dout(new_new_n6780__));
  buf1  g5839(.din(new_new_n6780__), .dout(new_new_n6781__));
  buf1  g5840(.din(new_new_n6780__), .dout(new_new_n6782__));
  buf1  g5841(.din(new_new_n6779__), .dout(new_new_n6783__));
  buf1  g5842(.din(new_new_n6783__), .dout(new_new_n6784__));
  buf1  g5843(.din(new_new_n1465__), .dout(new_new_n6785__));
  buf1  g5844(.din(new_new_n1402__), .dout(new_new_n6786__));
  buf1  g5845(.din(new_new_n1466__), .dout(new_new_n6787__));
  buf1  g5846(.din(new_new_n1401__), .dout(new_new_n6788__));
  buf1  g5847(.din(new_new_n2118__), .dout(new_new_n6789__));
  buf1  g5848(.din(new_new_n6789__), .dout(new_new_n6790__));
  buf1  g5849(.din(new_new_n2117__), .dout(new_new_n6791__));
  buf1  g5850(.din(new_new_n6791__), .dout(new_new_n6792__));
  buf1  g5851(.din(new_new_n2113__), .dout(new_new_n6793__));
  buf1  g5852(.din(new_new_n2126__), .dout(new_new_n6794__));
  buf1  g5853(.din(new_new_n2124__), .dout(new_new_n6795__));
  buf1  g5854(.din(new_new_n2125__), .dout(new_new_n6796__));
  buf1  g5855(.din(new_new_n2123__), .dout(new_new_n6797__));
  buf1  g5856(.din(new_new_n2128__), .dout(new_new_n6798__));
  buf1  g5857(.din(new_new_n6798__), .dout(new_new_n6799__));
  buf1  g5858(.din(new_new_n2127__), .dout(new_new_n6800__));
  buf1  g5859(.din(new_new_n6800__), .dout(new_new_n6801__));
  buf1  g5860(.din(new_new_n2134__), .dout(new_new_n6802__));
  buf1  g5861(.din(new_new_n2115__), .dout(new_new_n6803__));
  buf1  g5862(.din(new_new_n931__), .dout(new_new_n6804__));
  buf1  g5863(.din(new_new_n6804__), .dout(new_new_n6805__));
  buf1  g5864(.din(new_new_n6805__), .dout(new_new_n6806__));
  buf1  g5865(.din(new_new_n6806__), .dout(new_new_n6807__));
  buf1  g5866(.din(new_new_n6806__), .dout(new_new_n6808__));
  buf1  g5867(.din(new_new_n6805__), .dout(new_new_n6809__));
  buf1  g5868(.din(new_new_n6809__), .dout(new_new_n6810__));
  buf1  g5869(.din(new_new_n6804__), .dout(new_new_n6811__));
  buf1  g5870(.din(new_new_n6811__), .dout(new_new_n6812__));
  buf1  g5871(.din(new_new_n6811__), .dout(new_new_n6813__));
  buf1  g5872(.din(new_new_n932__), .dout(new_new_n6814__));
  buf1  g5873(.din(new_new_n6814__), .dout(new_new_n6815__));
  buf1  g5874(.din(new_new_n6815__), .dout(new_new_n6816__));
  buf1  g5875(.din(new_new_n6816__), .dout(new_new_n6817__));
  buf1  g5876(.din(new_new_n6816__), .dout(new_new_n6818__));
  buf1  g5877(.din(new_new_n6815__), .dout(new_new_n6819__));
  buf1  g5878(.din(new_new_n6819__), .dout(new_new_n6820__));
  buf1  g5879(.din(new_new_n6814__), .dout(new_new_n6821__));
  buf1  g5880(.din(new_new_n6821__), .dout(new_new_n6822__));
  buf1  g5881(.din(new_new_n6821__), .dout(new_new_n6823__));
  buf1  g5882(.din(new_new_n1448__), .dout(new_new_n6824__));
  buf1  g5883(.din(new_new_n6824__), .dout(new_new_n6825__));
  buf1  g5884(.din(new_new_n1447__), .dout(new_new_n6826__));
  buf1  g5885(.din(new_new_n6826__), .dout(new_new_n6827__));
  buf1  g5886(.din(new_new_n2146__), .dout(new_new_n6828__));
  buf1  g5887(.din(new_new_n2144__), .dout(new_new_n6829__));
  buf1  g5888(.din(new_new_n2145__), .dout(new_new_n6830__));
  buf1  g5889(.din(new_new_n2143__), .dout(new_new_n6831__));
  buf1  g5890(.din(new_new_n2148__), .dout(new_new_n6832__));
  buf1  g5891(.din(new_new_n6832__), .dout(new_new_n6833__));
  buf1  g5892(.din(new_new_n2147__), .dout(new_new_n6834__));
  buf1  g5893(.din(new_new_n6834__), .dout(new_new_n6835__));
  buf1  g5894(.din(new_new_n1039__), .dout(new_new_n6836__));
  buf1  g5895(.din(new_new_n6836__), .dout(new_new_n6837__));
  buf1  g5896(.din(new_new_n1040__), .dout(new_new_n6838__));
  buf1  g5897(.din(new_new_n6838__), .dout(new_new_n6839__));
  buf1  g5898(.din(new_new_n2156__), .dout(new_new_n6840__));
  buf1  g5899(.din(new_new_n2154__), .dout(new_new_n6841__));
  buf1  g5900(.din(new_new_n2155__), .dout(new_new_n6842__));
  buf1  g5901(.din(new_new_n2153__), .dout(new_new_n6843__));
  buf1  g5902(.din(new_new_n2158__), .dout(new_new_n6844__));
  buf1  g5903(.din(new_new_n6844__), .dout(new_new_n6845__));
  buf1  g5904(.din(new_new_n2157__), .dout(new_new_n6846__));
  buf1  g5905(.din(new_new_n6846__), .dout(new_new_n6847__));
  buf1  g5906(.din(new_new_n2135__), .dout(new_new_n6848__));
  buf1  g5907(.din(new_new_n2166__), .dout(new_new_n6849__));
  buf1  g5908(.din(new_new_n2164__), .dout(new_new_n6850__));
  buf1  g5909(.din(new_new_n2165__), .dout(new_new_n6851__));
  buf1  g5910(.din(new_new_n2163__), .dout(new_new_n6852__));
  buf1  g5911(.din(new_new_n2168__), .dout(new_new_n6853__));
  buf1  g5912(.din(new_new_n6853__), .dout(new_new_n6854__));
  buf1  g5913(.din(new_new_n2167__), .dout(new_new_n6855__));
  buf1  g5914(.din(new_new_n6855__), .dout(new_new_n6856__));
  buf1  g5915(.din(new_new_n2174__), .dout(new_new_n6857__));
  buf1  g5916(.din(new_new_n2137__), .dout(new_new_n6858__));
  buf1  g5917(.din(new_new_n1249__), .dout(new_new_n6859__));
  buf1  g5918(.din(new_new_n6859__), .dout(new_new_n6860__));
  buf1  g5919(.din(new_new_n6860__), .dout(new_new_n6861__));
  buf1  g5920(.din(new_new_n6859__), .dout(new_new_n6862__));
  buf1  g5921(.din(new_new_n1145__), .dout(new_new_n6863__));
  buf1  g5922(.din(new_new_n6863__), .dout(new_new_n6864__));
  buf1  g5923(.din(new_new_n6864__), .dout(new_new_n6865__));
  buf1  g5924(.din(new_new_n6864__), .dout(new_new_n6866__));
  buf1  g5925(.din(new_new_n6863__), .dout(new_new_n6867__));
  buf1  g5926(.din(new_new_n1250__), .dout(new_new_n6868__));
  buf1  g5927(.din(new_new_n6868__), .dout(new_new_n6869__));
  buf1  g5928(.din(new_new_n6869__), .dout(new_new_n6870__));
  buf1  g5929(.din(new_new_n6868__), .dout(new_new_n6871__));
  buf1  g5930(.din(new_new_n1146__), .dout(new_new_n6872__));
  buf1  g5931(.din(new_new_n6872__), .dout(new_new_n6873__));
  buf1  g5932(.din(new_new_n6873__), .dout(new_new_n6874__));
  buf1  g5933(.din(new_new_n6872__), .dout(new_new_n6875__));
  buf1  g5934(.din(new_new_n1533__), .dout(new_new_n6876__));
  buf1  g5935(.din(new_new_n6876__), .dout(new_new_n6877__));
  buf1  g5936(.din(new_new_n1534__), .dout(new_new_n6878__));
  buf1  g5937(.din(new_new_n6878__), .dout(new_new_n6879__));
  buf1  g5938(.din(new_new_n2184__), .dout(new_new_n6880__));
  buf1  g5939(.din(new_new_n2177__), .dout(new_new_n6881__));
  buf1  g5940(.din(new_new_n939__), .dout(new_new_n6882__));
  buf1  g5941(.din(new_new_n6882__), .dout(new_new_n6883__));
  buf1  g5942(.din(new_new_n6883__), .dout(new_new_n6884__));
  buf1  g5943(.din(new_new_n6883__), .dout(new_new_n6885__));
  buf1  g5944(.din(new_new_n6882__), .dout(new_new_n6886__));
  buf1  g5945(.din(new_new_n6886__), .dout(new_new_n6887__));
  buf1  g5946(.din(new_new_n940__), .dout(new_new_n6888__));
  buf1  g5947(.din(new_new_n6888__), .dout(new_new_n6889__));
  buf1  g5948(.din(new_new_n6889__), .dout(new_new_n6890__));
  buf1  g5949(.din(new_new_n6889__), .dout(new_new_n6891__));
  buf1  g5950(.din(new_new_n6888__), .dout(new_new_n6892__));
  buf1  g5951(.din(new_new_n6892__), .dout(new_new_n6893__));
  buf1  g5952(.din(new_new_n2192__), .dout(new_new_n6894__));
  buf1  g5953(.din(new_new_n2190__), .dout(new_new_n6895__));
  buf1  g5954(.din(new_new_n2191__), .dout(new_new_n6896__));
  buf1  g5955(.din(new_new_n2189__), .dout(new_new_n6897__));
  buf1  g5956(.din(new_new_n2194__), .dout(new_new_n6898__));
  buf1  g5957(.din(new_new_n6898__), .dout(new_new_n6899__));
  buf1  g5958(.din(new_new_n2193__), .dout(new_new_n6900__));
  buf1  g5959(.din(new_new_n6900__), .dout(new_new_n6901__));
  buf1  g5960(.din(new_new_n1035__), .dout(new_new_n6902__));
  buf1  g5961(.din(new_new_n6902__), .dout(new_new_n6903__));
  buf1  g5962(.din(new_new_n1036__), .dout(new_new_n6904__));
  buf1  g5963(.din(new_new_n6904__), .dout(new_new_n6905__));
  buf1  g5964(.din(new_new_n2202__), .dout(new_new_n6906__));
  buf1  g5965(.din(new_new_n2200__), .dout(new_new_n6907__));
  buf1  g5966(.din(new_new_n2201__), .dout(new_new_n6908__));
  buf1  g5967(.din(new_new_n2199__), .dout(new_new_n6909__));
  buf1  g5968(.din(new_new_n2204__), .dout(new_new_n6910__));
  buf1  g5969(.din(new_new_n6910__), .dout(new_new_n6911__));
  buf1  g5970(.din(new_new_n2203__), .dout(new_new_n6912__));
  buf1  g5971(.din(new_new_n6912__), .dout(new_new_n6913__));
  buf1  g5972(.din(new_new_n2212__), .dout(new_new_n6914__));
  buf1  g5973(.din(new_new_n2210__), .dout(new_new_n6915__));
  buf1  g5974(.din(new_new_n2211__), .dout(new_new_n6916__));
  buf1  g5975(.din(new_new_n2209__), .dout(new_new_n6917__));
  buf1  g5976(.din(new_new_n2214__), .dout(new_new_n6918__));
  buf1  g5977(.din(new_new_n6918__), .dout(new_new_n6919__));
  buf1  g5978(.din(new_new_n2213__), .dout(new_new_n6920__));
  buf1  g5979(.din(new_new_n6920__), .dout(new_new_n6921__));
  buf1  g5980(.din(new_new_n2222__), .dout(new_new_n6922__));
  buf1  g5981(.din(new_new_n2220__), .dout(new_new_n6923__));
  buf1  g5982(.din(new_new_n2221__), .dout(new_new_n6924__));
  buf1  g5983(.din(new_new_n2219__), .dout(new_new_n6925__));
  buf1  g5984(.din(new_new_n2224__), .dout(new_new_n6926__));
  buf1  g5985(.din(new_new_n6926__), .dout(new_new_n6927__));
  buf1  g5986(.din(new_new_n2223__), .dout(new_new_n6928__));
  buf1  g5987(.din(new_new_n6928__), .dout(new_new_n6929__));
  buf1  g5988(.din(new_new_n2175__), .dout(new_new_n6930__));
  buf1  g5989(.din(new_new_n2232__), .dout(new_new_n6931__));
  buf1  g5990(.din(new_new_n2230__), .dout(new_new_n6932__));
  buf1  g5991(.din(new_new_n2231__), .dout(new_new_n6933__));
  buf1  g5992(.din(new_new_n2229__), .dout(new_new_n6934__));
  buf1  g5993(.din(new_new_n2234__), .dout(new_new_n6935__));
  buf1  g5994(.din(new_new_n6935__), .dout(new_new_n6936__));
  buf1  g5995(.din(new_new_n2233__), .dout(new_new_n6937__));
  buf1  g5996(.din(new_new_n6937__), .dout(new_new_n6938__));
  buf1  g5997(.din(new_new_n1385__), .dout(new_new_n6939__));
  buf1  g5998(.din(new_new_n6939__), .dout(new_new_n6940__));
  buf1  g5999(.din(new_new_n6940__), .dout(new_new_n6941__));
  buf1  g6000(.din(new_new_n6941__), .dout(new_new_n6942__));
  buf1  g6001(.din(new_new_n6941__), .dout(new_new_n6943__));
  buf1  g6002(.din(new_new_n6940__), .dout(new_new_n6944__));
  buf1  g6003(.din(new_new_n6944__), .dout(new_new_n6945__));
  buf1  g6004(.din(new_new_n6944__), .dout(new_new_n6946__));
  buf1  g6005(.din(new_new_n6939__), .dout(new_new_n6947__));
  buf1  g6006(.din(new_new_n6947__), .dout(new_new_n6948__));
  buf1  g6007(.din(new_new_n6948__), .dout(new_new_n6949__));
  buf1  g6008(.din(new_new_n6948__), .dout(new_new_n6950__));
  buf1  g6009(.din(new_new_n6947__), .dout(new_new_n6951__));
  buf1  g6010(.din(new_new_n1386__), .dout(new_new_n6952__));
  buf1  g6011(.din(new_new_n6952__), .dout(new_new_n6953__));
  buf1  g6012(.din(new_new_n6953__), .dout(new_new_n6954__));
  buf1  g6013(.din(new_new_n6954__), .dout(new_new_n6955__));
  buf1  g6014(.din(new_new_n6954__), .dout(new_new_n6956__));
  buf1  g6015(.din(new_new_n6953__), .dout(new_new_n6957__));
  buf1  g6016(.din(new_new_n6957__), .dout(new_new_n6958__));
  buf1  g6017(.din(new_new_n6957__), .dout(new_new_n6959__));
  buf1  g6018(.din(new_new_n6952__), .dout(new_new_n6960__));
  buf1  g6019(.din(new_new_n6960__), .dout(new_new_n6961__));
  buf1  g6020(.din(new_new_n6961__), .dout(new_new_n6962__));
  buf1  g6021(.din(new_new_n6961__), .dout(new_new_n6963__));
  buf1  g6022(.din(new_new_n6960__), .dout(new_new_n6964__));
  buf1  g6023(.din(new_new_n2240__), .dout(new_new_n6965__));
  buf1  g6024(.din(new_new_n2187__), .dout(new_new_n6966__));
  buf1  g6025(.din(new_new_n1137__), .dout(new_new_n6967__));
  buf1  g6026(.din(new_new_n6967__), .dout(new_new_n6968__));
  buf1  g6027(.din(new_new_n6968__), .dout(new_new_n6969__));
  buf1  g6028(.din(new_new_n6968__), .dout(new_new_n6970__));
  buf1  g6029(.din(new_new_n6967__), .dout(new_new_n6971__));
  buf1  g6030(.din(new_new_n6971__), .dout(new_new_n6972__));
  buf1  g6031(.din(new_new_n1138__), .dout(new_new_n6973__));
  buf1  g6032(.din(new_new_n6973__), .dout(new_new_n6974__));
  buf1  g6033(.din(new_new_n6974__), .dout(new_new_n6975__));
  buf1  g6034(.din(new_new_n6973__), .dout(new_new_n6976__));
  buf1  g6035(.din(new_new_n2248__), .dout(new_new_n6977__));
  buf1  g6036(.din(new_new_n2246__), .dout(new_new_n6978__));
  buf1  g6037(.din(new_new_n2247__), .dout(new_new_n6979__));
  buf1  g6038(.din(new_new_n2245__), .dout(new_new_n6980__));
  buf1  g6039(.din(new_new_n2250__), .dout(new_new_n6981__));
  buf1  g6040(.din(new_new_n6981__), .dout(new_new_n6982__));
  buf1  g6041(.din(new_new_n2249__), .dout(new_new_n6983__));
  buf1  g6042(.din(new_new_n6983__), .dout(new_new_n6984__));
  buf1  g6043(.din(new_new_n2185__), .dout(new_new_n6985__));
  buf1  g6044(.din(new_new_n2258__), .dout(new_new_n6986__));
  buf1  g6045(.din(new_new_n2256__), .dout(new_new_n6987__));
  buf1  g6046(.din(new_new_n2257__), .dout(new_new_n6988__));
  buf1  g6047(.din(new_new_n2255__), .dout(new_new_n6989__));
  buf1  g6048(.din(new_new_n2260__), .dout(new_new_n6990__));
  buf1  g6049(.din(new_new_n6990__), .dout(new_new_n6991__));
  buf1  g6050(.din(new_new_n2259__), .dout(new_new_n6992__));
  buf1  g6051(.din(new_new_n6992__), .dout(new_new_n6993__));
  buf1  g6052(.din(new_new_n2266__), .dout(new_new_n6994__));
  buf1  g6053(.din(new_new_n2241__), .dout(new_new_n6995__));
  buf1  g6054(.din(new_new_n1399__), .dout(new_new_n6996__));
  buf1  g6055(.din(new_new_n6996__), .dout(new_new_n6997__));
  buf1  g6056(.din(new_new_n6997__), .dout(new_new_n6998__));
  buf1  g6057(.din(new_new_n6996__), .dout(new_new_n6999__));
  buf1  g6058(.din(new_new_n1231__), .dout(new_new_n7000__));
  buf1  g6059(.din(new_new_n7000__), .dout(new_new_n7001__));
  buf1  g6060(.din(new_new_n1400__), .dout(new_new_n7002__));
  buf1  g6061(.din(new_new_n7002__), .dout(new_new_n7003__));
  buf1  g6062(.din(new_new_n7003__), .dout(new_new_n7004__));
  buf1  g6063(.din(new_new_n7002__), .dout(new_new_n7005__));
  buf1  g6064(.din(new_new_n1232__), .dout(new_new_n7006__));
  buf1  g6065(.din(new_new_n7006__), .dout(new_new_n7007__));
  buf1  g6066(.din(new_new_n1606__), .dout(new_new_n7008__));
  buf1  g6067(.din(new_new_n1568__), .dout(new_new_n7009__));
  buf1  g6068(.din(new_new_n1605__), .dout(new_new_n7010__));
  buf1  g6069(.din(new_new_n1567__), .dout(new_new_n7011__));
  buf1  g6070(.din(new_new_n2272__), .dout(new_new_n7012__));
  buf1  g6071(.din(new_new_n7012__), .dout(new_new_n7013__));
  buf1  g6072(.din(new_new_n2271__), .dout(new_new_n7014__));
  buf1  g6073(.din(new_new_n7014__), .dout(new_new_n7015__));
  buf1  g6074(.din(new_new_n905__), .dout(new_new_n7016__));
  buf1  g6075(.din(new_new_n7016__), .dout(new_new_n7017__));
  buf1  g6076(.din(new_new_n7017__), .dout(new_new_n7018__));
  buf1  g6077(.din(new_new_n7018__), .dout(new_new_n7019__));
  buf1  g6078(.din(new_new_n7018__), .dout(new_new_n7020__));
  buf1  g6079(.din(new_new_n7017__), .dout(new_new_n7021__));
  buf1  g6080(.din(new_new_n7021__), .dout(new_new_n7022__));
  buf1  g6081(.din(new_new_n7021__), .dout(new_new_n7023__));
  buf1  g6082(.din(new_new_n7016__), .dout(new_new_n7024__));
  buf1  g6083(.din(new_new_n7024__), .dout(new_new_n7025__));
  buf1  g6084(.din(new_new_n7025__), .dout(new_new_n7026__));
  buf1  g6085(.din(new_new_n7025__), .dout(new_new_n7027__));
  buf1  g6086(.din(new_new_n7024__), .dout(new_new_n7028__));
  buf1  g6087(.din(new_new_n7028__), .dout(new_new_n7029__));
  buf1  g6088(.din(new_new_n7028__), .dout(new_new_n7030__));
  buf1  g6089(.din(new_new_n906__), .dout(new_new_n7031__));
  buf1  g6090(.din(new_new_n7031__), .dout(new_new_n7032__));
  buf1  g6091(.din(new_new_n7032__), .dout(new_new_n7033__));
  buf1  g6092(.din(new_new_n7033__), .dout(new_new_n7034__));
  buf1  g6093(.din(new_new_n7033__), .dout(new_new_n7035__));
  buf1  g6094(.din(new_new_n7032__), .dout(new_new_n7036__));
  buf1  g6095(.din(new_new_n7036__), .dout(new_new_n7037__));
  buf1  g6096(.din(new_new_n7036__), .dout(new_new_n7038__));
  buf1  g6097(.din(new_new_n7031__), .dout(new_new_n7039__));
  buf1  g6098(.din(new_new_n7039__), .dout(new_new_n7040__));
  buf1  g6099(.din(new_new_n7040__), .dout(new_new_n7041__));
  buf1  g6100(.din(new_new_n7040__), .dout(new_new_n7042__));
  buf1  g6101(.din(new_new_n7039__), .dout(new_new_n7043__));
  buf1  g6102(.din(new_new_n7043__), .dout(new_new_n7044__));
  buf1  g6103(.din(new_new_n7043__), .dout(new_new_n7045__));
  buf1  g6104(.din(new_new_n2278__), .dout(new_new_n7046__));
  buf1  g6105(.din(new_new_n2269__), .dout(new_new_n7047__));
  buf1  g6106(.din(new_new_n1547__), .dout(new_new_n7048__));
  buf1  g6107(.din(new_new_n1488__), .dout(new_new_n7049__));
  buf1  g6108(.din(new_new_n1548__), .dout(new_new_n7050__));
  buf1  g6109(.din(new_new_n1487__), .dout(new_new_n7051__));
  buf1  g6110(.din(new_new_n2284__), .dout(new_new_n7052__));
  buf1  g6111(.din(new_new_n7052__), .dout(new_new_n7053__));
  buf1  g6112(.din(new_new_n2283__), .dout(new_new_n7054__));
  buf1  g6113(.din(new_new_n7054__), .dout(new_new_n7055__));
  buf1  g6114(.din(new_new_n2292__), .dout(new_new_n7056__));
  buf1  g6115(.din(new_new_n2290__), .dout(new_new_n7057__));
  buf1  g6116(.din(new_new_n2291__), .dout(new_new_n7058__));
  buf1  g6117(.din(new_new_n2289__), .dout(new_new_n7059__));
  buf1  g6118(.din(new_new_n2294__), .dout(new_new_n7060__));
  buf1  g6119(.din(new_new_n7060__), .dout(new_new_n7061__));
  buf1  g6120(.din(new_new_n2293__), .dout(new_new_n7062__));
  buf1  g6121(.din(new_new_n7062__), .dout(new_new_n7063__));
  buf1  g6122(.din(new_new_n2302__), .dout(new_new_n7064__));
  buf1  g6123(.din(new_new_n2300__), .dout(new_new_n7065__));
  buf1  g6124(.din(new_new_n2301__), .dout(new_new_n7066__));
  buf1  g6125(.din(new_new_n2299__), .dout(new_new_n7067__));
  buf1  g6126(.din(new_new_n2304__), .dout(new_new_n7068__));
  buf1  g6127(.din(new_new_n7068__), .dout(new_new_n7069__));
  buf1  g6128(.din(new_new_n2303__), .dout(new_new_n7070__));
  buf1  g6129(.din(new_new_n7070__), .dout(new_new_n7071__));
  buf1  g6130(.din(new_new_n2267__), .dout(new_new_n7072__));
  buf1  g6131(.din(new_new_n2312__), .dout(new_new_n7073__));
  buf1  g6132(.din(new_new_n2310__), .dout(new_new_n7074__));
  buf1  g6133(.din(new_new_n2311__), .dout(new_new_n7075__));
  buf1  g6134(.din(new_new_n2309__), .dout(new_new_n7076__));
  buf1  g6135(.din(new_new_n2314__), .dout(new_new_n7077__));
  buf1  g6136(.din(new_new_n7077__), .dout(new_new_n7078__));
  buf1  g6137(.din(new_new_n2313__), .dout(new_new_n7079__));
  buf1  g6138(.din(new_new_n7079__), .dout(new_new_n7080__));
  buf1  g6139(.din(new_new_n2320__), .dout(new_new_n7081__));
  buf1  g6140(.din(new_new_n2279__), .dout(new_new_n7082__));
  buf1  g6141(.din(new_new_n1315__), .dout(new_new_n7083__));
  buf1  g6142(.din(new_new_n7083__), .dout(new_new_n7084__));
  buf1  g6143(.din(new_new_n7084__), .dout(new_new_n7085__));
  buf1  g6144(.din(new_new_n7085__), .dout(new_new_n7086__));
  buf1  g6145(.din(new_new_n7084__), .dout(new_new_n7087__));
  buf1  g6146(.din(new_new_n7083__), .dout(new_new_n7088__));
  buf1  g6147(.din(new_new_n7088__), .dout(new_new_n7089__));
  buf1  g6148(.din(new_new_n7088__), .dout(new_new_n7090__));
  buf1  g6149(.din(new_new_n1316__), .dout(new_new_n7091__));
  buf1  g6150(.din(new_new_n7091__), .dout(new_new_n7092__));
  buf1  g6151(.din(new_new_n7092__), .dout(new_new_n7093__));
  buf1  g6152(.din(new_new_n7093__), .dout(new_new_n7094__));
  buf1  g6153(.din(new_new_n7092__), .dout(new_new_n7095__));
  buf1  g6154(.din(new_new_n7091__), .dout(new_new_n7096__));
  buf1  g6155(.din(new_new_n7096__), .dout(new_new_n7097__));
  buf1  g6156(.din(new_new_n7096__), .dout(new_new_n7098__));
  buf1  g6157(.din(new_new_n1597__), .dout(new_new_n7099__));
  buf1  g6158(.din(new_new_n7099__), .dout(new_new_n7100__));
  buf1  g6159(.din(new_new_n1598__), .dout(new_new_n7101__));
  buf1  g6160(.din(new_new_n7101__), .dout(new_new_n7102__));
  buf1  g6161(.din(new_new_n1313__), .dout(new_new_n7103__));
  buf1  g6162(.din(new_new_n7103__), .dout(new_new_n7104__));
  buf1  g6163(.din(new_new_n7104__), .dout(new_new_n7105__));
  buf1  g6164(.din(new_new_n7104__), .dout(new_new_n7106__));
  buf1  g6165(.din(new_new_n7103__), .dout(new_new_n7107__));
  buf1  g6166(.din(new_new_n1314__), .dout(new_new_n7108__));
  buf1  g6167(.din(new_new_n7108__), .dout(new_new_n7109__));
  buf1  g6168(.din(new_new_n7109__), .dout(new_new_n7110__));
  buf1  g6169(.din(new_new_n7108__), .dout(new_new_n7111__));
  buf1  g6170(.din(new_new_n2332__), .dout(new_new_n7112__));
  buf1  g6171(.din(new_new_n2330__), .dout(new_new_n7113__));
  buf1  g6172(.din(new_new_n2331__), .dout(new_new_n7114__));
  buf1  g6173(.din(new_new_n2329__), .dout(new_new_n7115__));
  buf1  g6174(.din(new_new_n2334__), .dout(new_new_n7116__));
  buf1  g6175(.din(new_new_n7116__), .dout(new_new_n7117__));
  buf1  g6176(.din(new_new_n2333__), .dout(new_new_n7118__));
  buf1  g6177(.din(new_new_n7118__), .dout(new_new_n7119__));
  buf1  g6178(.din(new_new_n2281__), .dout(new_new_n7120__));
  buf1  g6179(.din(new_new_n2342__), .dout(new_new_n7121__));
  buf1  g6180(.din(new_new_n2340__), .dout(new_new_n7122__));
  buf1  g6181(.din(new_new_n2341__), .dout(new_new_n7123__));
  buf1  g6182(.din(new_new_n2339__), .dout(new_new_n7124__));
  buf1  g6183(.din(new_new_n2344__), .dout(new_new_n7125__));
  buf1  g6184(.din(new_new_n7125__), .dout(new_new_n7126__));
  buf1  g6185(.din(new_new_n2343__), .dout(new_new_n7127__));
  buf1  g6186(.din(new_new_n7127__), .dout(new_new_n7128__));
  buf1  g6187(.din(new_new_n1183__), .dout(new_new_n7129__));
  buf1  g6188(.din(new_new_n7129__), .dout(new_new_n7130__));
  buf1  g6189(.din(new_new_n7130__), .dout(new_new_n7131__));
  buf1  g6190(.din(new_new_n7130__), .dout(new_new_n7132__));
  buf1  g6191(.din(new_new_n7129__), .dout(new_new_n7133__));
  buf1  g6192(.din(new_new_n997__), .dout(new_new_n7134__));
  buf1  g6193(.din(new_new_n7134__), .dout(new_new_n7135__));
  buf1  g6194(.din(new_new_n7134__), .dout(new_new_n7136__));
  buf1  g6195(.din(new_new_n1184__), .dout(new_new_n7137__));
  buf1  g6196(.din(new_new_n7137__), .dout(new_new_n7138__));
  buf1  g6197(.din(new_new_n7138__), .dout(new_new_n7139__));
  buf1  g6198(.din(new_new_n7138__), .dout(new_new_n7140__));
  buf1  g6199(.din(new_new_n7137__), .dout(new_new_n7141__));
  buf1  g6200(.din(new_new_n998__), .dout(new_new_n7142__));
  buf1  g6201(.din(new_new_n7142__), .dout(new_new_n7143__));
  buf1  g6202(.din(new_new_n1155__), .dout(new_new_n7144__));
  buf1  g6203(.din(new_new_n1156__), .dout(new_new_n7145__));
  buf1  g6204(.din(new_new_n1003__), .dout(new_new_n7146__));
  buf1  g6205(.din(new_new_n7146__), .dout(new_new_n7147__));
  buf1  g6206(.din(new_new_n7146__), .dout(new_new_n7148__));
  buf1  g6207(.din(new_new_n1004__), .dout(new_new_n7149__));
  buf1  g6208(.din(new_new_n7149__), .dout(new_new_n7150__));
  buf1  g6209(.din(new_new_n7149__), .dout(new_new_n7151__));
  buf1  g6210(.din(new_new_n2358__), .dout(new_new_n7152__));
  buf1  g6211(.din(new_new_n2356__), .dout(new_new_n7153__));
  buf1  g6212(.din(new_new_n2357__), .dout(new_new_n7154__));
  buf1  g6213(.din(new_new_n2355__), .dout(new_new_n7155__));
  buf1  g6214(.din(new_new_n2360__), .dout(new_new_n7156__));
  buf1  g6215(.din(new_new_n7156__), .dout(new_new_n7157__));
  buf1  g6216(.din(new_new_n2359__), .dout(new_new_n7158__));
  buf1  g6217(.din(new_new_n7158__), .dout(new_new_n7159__));
  buf1  g6218(.din(new_new_n2362__), .dout(new_new_n7160__));
  buf1  g6219(.din(new_new_n2354__), .dout(new_new_n7161__));
  buf1  g6220(.din(new_new_n2361__), .dout(new_new_n7162__));
  buf1  g6221(.din(new_new_n2353__), .dout(new_new_n7163__));
  buf1  g6222(.din(new_new_n2364__), .dout(new_new_n7164__));
  buf1  g6223(.din(new_new_n7164__), .dout(new_new_n7165__));
  buf1  g6224(.din(new_new_n2363__), .dout(new_new_n7166__));
  buf1  g6225(.din(new_new_n7166__), .dout(new_new_n7167__));
  buf1  g6226(.din(new_new_n2372__), .dout(new_new_n7168__));
  buf1  g6227(.din(new_new_n2370__), .dout(new_new_n7169__));
  buf1  g6228(.din(new_new_n2371__), .dout(new_new_n7170__));
  buf1  g6229(.din(new_new_n2369__), .dout(new_new_n7171__));
  buf1  g6230(.din(new_new_n2374__), .dout(new_new_n7172__));
  buf1  g6231(.din(new_new_n7172__), .dout(new_new_n7173__));
  buf1  g6232(.din(new_new_n2373__), .dout(new_new_n7174__));
  buf1  g6233(.din(new_new_n7174__), .dout(new_new_n7175__));
  buf1  g6234(.din(new_new_n2376__), .dout(new_new_n7176__));
  buf1  g6235(.din(new_new_n2352__), .dout(new_new_n7177__));
  buf1  g6236(.din(new_new_n2375__), .dout(new_new_n7178__));
  buf1  g6237(.din(new_new_n2351__), .dout(new_new_n7179__));
  buf1  g6238(.din(new_new_n2378__), .dout(new_new_n7180__));
  buf1  g6239(.din(new_new_n7180__), .dout(new_new_n7181__));
  buf1  g6240(.din(new_new_n2377__), .dout(new_new_n7182__));
  buf1  g6241(.din(new_new_n7182__), .dout(new_new_n7183__));
  buf1  g6242(.din(new_new_n2386__), .dout(new_new_n7184__));
  buf1  g6243(.din(new_new_n2384__), .dout(new_new_n7185__));
  buf1  g6244(.din(new_new_n2385__), .dout(new_new_n7186__));
  buf1  g6245(.din(new_new_n2383__), .dout(new_new_n7187__));
  buf1  g6246(.din(new_new_n2388__), .dout(new_new_n7188__));
  buf1  g6247(.din(new_new_n7188__), .dout(new_new_n7189__));
  buf1  g6248(.din(new_new_n2387__), .dout(new_new_n7190__));
  buf1  g6249(.din(new_new_n7190__), .dout(new_new_n7191__));
  buf1  g6250(.din(new_new_n1442__), .dout(new_new_n7192__));
  buf1  g6251(.din(new_new_n7192__), .dout(new_new_n7193__));
  buf1  g6252(.din(new_new_n1441__), .dout(new_new_n7194__));
  buf1  g6253(.din(new_new_n7194__), .dout(new_new_n7195__));
  buf1  g6254(.din(new_new_n2408__), .dout(new_new_n7196__));
  buf1  g6255(.din(new_new_n2406__), .dout(new_new_n7197__));
  buf1  g6256(.din(new_new_n2407__), .dout(new_new_n7198__));
  buf1  g6257(.din(new_new_n2405__), .dout(new_new_n7199__));
  buf1  g6258(.din(new_new_n2410__), .dout(new_new_n7200__));
  buf1  g6259(.din(new_new_n7200__), .dout(new_new_n7201__));
  buf1  g6260(.din(new_new_n2409__), .dout(new_new_n7202__));
  buf1  g6261(.din(new_new_n7202__), .dout(new_new_n7203__));
  buf1  g6262(.din(new_new_n1007__), .dout(new_new_n7204__));
  buf1  g6263(.din(new_new_n7204__), .dout(new_new_n7205__));
  buf1  g6264(.din(new_new_n7204__), .dout(new_new_n7206__));
  buf1  g6265(.din(new_new_n1008__), .dout(new_new_n7207__));
  buf1  g6266(.din(new_new_n7207__), .dout(new_new_n7208__));
  buf1  g6267(.din(new_new_n2418__), .dout(new_new_n7209__));
  buf1  g6268(.din(new_new_n2416__), .dout(new_new_n7210__));
  buf1  g6269(.din(new_new_n2417__), .dout(new_new_n7211__));
  buf1  g6270(.din(new_new_n2415__), .dout(new_new_n7212__));
  buf1  g6271(.din(new_new_n2420__), .dout(new_new_n7213__));
  buf1  g6272(.din(new_new_n7213__), .dout(new_new_n7214__));
  buf1  g6273(.din(new_new_n2419__), .dout(new_new_n7215__));
  buf1  g6274(.din(new_new_n7215__), .dout(new_new_n7216__));
  buf1  g6275(.din(new_new_n2422__), .dout(new_new_n7217__));
  buf1  g6276(.din(new_new_n2400__), .dout(new_new_n7218__));
  buf1  g6277(.din(new_new_n2421__), .dout(new_new_n7219__));
  buf1  g6278(.din(new_new_n2399__), .dout(new_new_n7220__));
  buf1  g6279(.din(new_new_n2424__), .dout(new_new_n7221__));
  buf1  g6280(.din(new_new_n7221__), .dout(new_new_n7222__));
  buf1  g6281(.din(new_new_n2423__), .dout(new_new_n7223__));
  buf1  g6282(.din(new_new_n7223__), .dout(new_new_n7224__));
  buf1  g6283(.din(new_new_n2432__), .dout(new_new_n7225__));
  buf1  g6284(.din(new_new_n2430__), .dout(new_new_n7226__));
  buf1  g6285(.din(new_new_n2431__), .dout(new_new_n7227__));
  buf1  g6286(.din(new_new_n2429__), .dout(new_new_n7228__));
  buf1  g6287(.din(new_new_n2434__), .dout(new_new_n7229__));
  buf1  g6288(.din(new_new_n7229__), .dout(new_new_n7230__));
  buf1  g6289(.din(new_new_n2433__), .dout(new_new_n7231__));
  buf1  g6290(.din(new_new_n7231__), .dout(new_new_n7232__));
  buf1  g6291(.din(new_new_n2436__), .dout(new_new_n7233__));
  buf1  g6292(.din(new_new_n2394__), .dout(new_new_n7234__));
  buf1  g6293(.din(new_new_n2435__), .dout(new_new_n7235__));
  buf1  g6294(.din(new_new_n2393__), .dout(new_new_n7236__));
  buf1  g6295(.din(new_new_n2446__), .dout(new_new_n7237__));
  buf1  g6296(.din(new_new_n2444__), .dout(new_new_n7238__));
  buf1  g6297(.din(new_new_n2445__), .dout(new_new_n7239__));
  buf1  g6298(.din(new_new_n2443__), .dout(new_new_n7240__));
  buf1  g6299(.din(new_new_n2448__), .dout(new_new_n7241__));
  buf1  g6300(.din(new_new_n7241__), .dout(new_new_n7242__));
  buf1  g6301(.din(new_new_n2447__), .dout(new_new_n7243__));
  buf1  g6302(.din(new_new_n7243__), .dout(new_new_n7244__));
  buf1  g6303(.din(new_new_n1009__), .dout(new_new_n7245__));
  buf1  g6304(.din(new_new_n7245__), .dout(new_new_n7246__));
  buf1  g6305(.din(new_new_n7245__), .dout(new_new_n7247__));
  buf1  g6306(.din(new_new_n1010__), .dout(new_new_n7248__));
  buf1  g6307(.din(new_new_n7248__), .dout(new_new_n7249__));
  buf1  g6308(.din(new_new_n2456__), .dout(new_new_n7250__));
  buf1  g6309(.din(new_new_n2454__), .dout(new_new_n7251__));
  buf1  g6310(.din(new_new_n2455__), .dout(new_new_n7252__));
  buf1  g6311(.din(new_new_n2453__), .dout(new_new_n7253__));
  buf1  g6312(.din(new_new_n2458__), .dout(new_new_n7254__));
  buf1  g6313(.din(new_new_n7254__), .dout(new_new_n7255__));
  buf1  g6314(.din(new_new_n2457__), .dout(new_new_n7256__));
  buf1  g6315(.din(new_new_n7256__), .dout(new_new_n7257__));
  buf1  g6316(.din(new_new_n1460__), .dout(new_new_n7258__));
  buf1  g6317(.din(new_new_n1412__), .dout(new_new_n7259__));
  buf1  g6318(.din(new_new_n1459__), .dout(new_new_n7260__));
  buf1  g6319(.din(new_new_n1411__), .dout(new_new_n7261__));
  buf1  g6320(.din(new_new_n2466__), .dout(new_new_n7262__));
  buf1  g6321(.din(new_new_n7262__), .dout(new_new_n7263__));
  buf1  g6322(.din(new_new_n2465__), .dout(new_new_n7264__));
  buf1  g6323(.din(new_new_n7264__), .dout(new_new_n7265__));
  buf1  g6324(.din(new_new_n1013__), .dout(new_new_n7266__));
  buf1  g6325(.din(new_new_n7266__), .dout(new_new_n7267__));
  buf1  g6326(.din(new_new_n7266__), .dout(new_new_n7268__));
  buf1  g6327(.din(new_new_n1014__), .dout(new_new_n7269__));
  buf1  g6328(.din(new_new_n7269__), .dout(new_new_n7270__));
  buf1  g6329(.din(new_new_n2474__), .dout(new_new_n7271__));
  buf1  g6330(.din(new_new_n2472__), .dout(new_new_n7272__));
  buf1  g6331(.din(new_new_n2473__), .dout(new_new_n7273__));
  buf1  g6332(.din(new_new_n2471__), .dout(new_new_n7274__));
  buf1  g6333(.din(new_new_n2476__), .dout(new_new_n7275__));
  buf1  g6334(.din(new_new_n7275__), .dout(new_new_n7276__));
  buf1  g6335(.din(new_new_n2475__), .dout(new_new_n7277__));
  buf1  g6336(.din(new_new_n7277__), .dout(new_new_n7278__));
  buf1  g6337(.din(new_new_n2478__), .dout(new_new_n7279__));
  buf1  g6338(.din(new_new_n2464__), .dout(new_new_n7280__));
  buf1  g6339(.din(new_new_n2477__), .dout(new_new_n7281__));
  buf1  g6340(.din(new_new_n2463__), .dout(new_new_n7282__));
  buf1  g6341(.din(new_new_n2480__), .dout(new_new_n7283__));
  buf1  g6342(.din(new_new_n7283__), .dout(new_new_n7284__));
  buf1  g6343(.din(new_new_n2479__), .dout(new_new_n7285__));
  buf1  g6344(.din(new_new_n7285__), .dout(new_new_n7286__));
  buf1  g6345(.din(new_new_n2488__), .dout(new_new_n7287__));
  buf1  g6346(.din(new_new_n2486__), .dout(new_new_n7288__));
  buf1  g6347(.din(new_new_n2487__), .dout(new_new_n7289__));
  buf1  g6348(.din(new_new_n2485__), .dout(new_new_n7290__));
  buf1  g6349(.din(new_new_n2490__), .dout(new_new_n7291__));
  buf1  g6350(.din(new_new_n7291__), .dout(new_new_n7292__));
  buf1  g6351(.din(new_new_n2489__), .dout(new_new_n7293__));
  buf1  g6352(.din(new_new_n7293__), .dout(new_new_n7294__));
  buf1  g6353(.din(new_new_n1015__), .dout(new_new_n7295__));
  buf1  g6354(.din(new_new_n7295__), .dout(new_new_n7296__));
  buf1  g6355(.din(new_new_n7295__), .dout(new_new_n7297__));
  buf1  g6356(.din(new_new_n1016__), .dout(new_new_n7298__));
  buf1  g6357(.din(new_new_n7298__), .dout(new_new_n7299__));
  buf1  g6358(.din(new_new_n7298__), .dout(new_new_n7300__));
  buf1  g6359(.din(new_new_n2506__), .dout(new_new_n7301__));
  buf1  g6360(.din(new_new_n2504__), .dout(new_new_n7302__));
  buf1  g6361(.din(new_new_n2505__), .dout(new_new_n7303__));
  buf1  g6362(.din(new_new_n2503__), .dout(new_new_n7304__));
  buf1  g6363(.din(new_new_n2508__), .dout(new_new_n7305__));
  buf1  g6364(.din(new_new_n7305__), .dout(new_new_n7306__));
  buf1  g6365(.din(new_new_n2507__), .dout(new_new_n7307__));
  buf1  g6366(.din(new_new_n7307__), .dout(new_new_n7308__));
  buf1  g6367(.din(new_new_n2510__), .dout(new_new_n7309__));
  buf1  g6368(.din(new_new_n2502__), .dout(new_new_n7310__));
  buf1  g6369(.din(new_new_n2509__), .dout(new_new_n7311__));
  buf1  g6370(.din(new_new_n2501__), .dout(new_new_n7312__));
  buf1  g6371(.din(new_new_n2512__), .dout(new_new_n7313__));
  buf1  g6372(.din(new_new_n7313__), .dout(new_new_n7314__));
  buf1  g6373(.din(new_new_n2511__), .dout(new_new_n7315__));
  buf1  g6374(.din(new_new_n7315__), .dout(new_new_n7316__));
  buf1  g6375(.din(new_new_n2520__), .dout(new_new_n7317__));
  buf1  g6376(.din(new_new_n2518__), .dout(new_new_n7318__));
  buf1  g6377(.din(new_new_n2519__), .dout(new_new_n7319__));
  buf1  g6378(.din(new_new_n2517__), .dout(new_new_n7320__));
  buf1  g6379(.din(new_new_n2522__), .dout(new_new_n7321__));
  buf1  g6380(.din(new_new_n7321__), .dout(new_new_n7322__));
  buf1  g6381(.din(new_new_n2521__), .dout(new_new_n7323__));
  buf1  g6382(.din(new_new_n7323__), .dout(new_new_n7324__));
  buf1  g6383(.din(new_new_n2524__), .dout(new_new_n7325__));
  buf1  g6384(.din(new_new_n2496__), .dout(new_new_n7326__));
  buf1  g6385(.din(new_new_n2523__), .dout(new_new_n7327__));
  buf1  g6386(.din(new_new_n2495__), .dout(new_new_n7328__));
  buf1  g6387(.din(new_new_n2526__), .dout(new_new_n7329__));
  buf1  g6388(.din(new_new_n7329__), .dout(new_new_n7330__));
  buf1  g6389(.din(new_new_n2525__), .dout(new_new_n7331__));
  buf1  g6390(.din(new_new_n7331__), .dout(new_new_n7332__));
  buf1  g6391(.din(new_new_n2534__), .dout(new_new_n7333__));
  buf1  g6392(.din(new_new_n2532__), .dout(new_new_n7334__));
  buf1  g6393(.din(new_new_n2533__), .dout(new_new_n7335__));
  buf1  g6394(.din(new_new_n2531__), .dout(new_new_n7336__));
  buf1  g6395(.din(new_new_n2536__), .dout(new_new_n7337__));
  buf1  g6396(.din(new_new_n7337__), .dout(new_new_n7338__));
  buf1  g6397(.din(new_new_n2535__), .dout(new_new_n7339__));
  buf1  g6398(.din(new_new_n7339__), .dout(new_new_n7340__));
  buf1  g6399(.din(new_new_n1444__), .dout(new_new_n7341__));
  buf1  g6400(.din(new_new_n7341__), .dout(new_new_n7342__));
  buf1  g6401(.din(new_new_n1443__), .dout(new_new_n7343__));
  buf1  g6402(.din(new_new_n7343__), .dout(new_new_n7344__));
  buf1  g6403(.din(new_new_n2556__), .dout(new_new_n7345__));
  buf1  g6404(.din(new_new_n2554__), .dout(new_new_n7346__));
  buf1  g6405(.din(new_new_n2555__), .dout(new_new_n7347__));
  buf1  g6406(.din(new_new_n2553__), .dout(new_new_n7348__));
  buf1  g6407(.din(new_new_n2558__), .dout(new_new_n7349__));
  buf1  g6408(.din(new_new_n7349__), .dout(new_new_n7350__));
  buf1  g6409(.din(new_new_n2557__), .dout(new_new_n7351__));
  buf1  g6410(.din(new_new_n7351__), .dout(new_new_n7352__));
  buf1  g6411(.din(new_new_n1017__), .dout(new_new_n7353__));
  buf1  g6412(.din(new_new_n7353__), .dout(new_new_n7354__));
  buf1  g6413(.din(new_new_n7353__), .dout(new_new_n7355__));
  buf1  g6414(.din(new_new_n1018__), .dout(new_new_n7356__));
  buf1  g6415(.din(new_new_n7356__), .dout(new_new_n7357__));
  buf1  g6416(.din(new_new_n2566__), .dout(new_new_n7358__));
  buf1  g6417(.din(new_new_n2564__), .dout(new_new_n7359__));
  buf1  g6418(.din(new_new_n2565__), .dout(new_new_n7360__));
  buf1  g6419(.din(new_new_n2563__), .dout(new_new_n7361__));
  buf1  g6420(.din(new_new_n2568__), .dout(new_new_n7362__));
  buf1  g6421(.din(new_new_n7362__), .dout(new_new_n7363__));
  buf1  g6422(.din(new_new_n2567__), .dout(new_new_n7364__));
  buf1  g6423(.din(new_new_n7364__), .dout(new_new_n7365__));
  buf1  g6424(.din(new_new_n2570__), .dout(new_new_n7366__));
  buf1  g6425(.din(new_new_n2548__), .dout(new_new_n7367__));
  buf1  g6426(.din(new_new_n2569__), .dout(new_new_n7368__));
  buf1  g6427(.din(new_new_n2547__), .dout(new_new_n7369__));
  buf1  g6428(.din(new_new_n2572__), .dout(new_new_n7370__));
  buf1  g6429(.din(new_new_n7370__), .dout(new_new_n7371__));
  buf1  g6430(.din(new_new_n2571__), .dout(new_new_n7372__));
  buf1  g6431(.din(new_new_n7372__), .dout(new_new_n7373__));
  buf1  g6432(.din(new_new_n2580__), .dout(new_new_n7374__));
  buf1  g6433(.din(new_new_n2578__), .dout(new_new_n7375__));
  buf1  g6434(.din(new_new_n2579__), .dout(new_new_n7376__));
  buf1  g6435(.din(new_new_n2577__), .dout(new_new_n7377__));
  buf1  g6436(.din(new_new_n2582__), .dout(new_new_n7378__));
  buf1  g6437(.din(new_new_n7378__), .dout(new_new_n7379__));
  buf1  g6438(.din(new_new_n2581__), .dout(new_new_n7380__));
  buf1  g6439(.din(new_new_n7380__), .dout(new_new_n7381__));
  buf1  g6440(.din(new_new_n2584__), .dout(new_new_n7382__));
  buf1  g6441(.din(new_new_n2542__), .dout(new_new_n7383__));
  buf1  g6442(.din(new_new_n2583__), .dout(new_new_n7384__));
  buf1  g6443(.din(new_new_n2541__), .dout(new_new_n7385__));
  buf1  g6444(.din(new_new_n2594__), .dout(new_new_n7386__));
  buf1  g6445(.din(new_new_n2592__), .dout(new_new_n7387__));
  buf1  g6446(.din(new_new_n2593__), .dout(new_new_n7388__));
  buf1  g6447(.din(new_new_n2591__), .dout(new_new_n7389__));
  buf1  g6448(.din(new_new_n2596__), .dout(new_new_n7390__));
  buf1  g6449(.din(new_new_n7390__), .dout(new_new_n7391__));
  buf1  g6450(.din(new_new_n2595__), .dout(new_new_n7392__));
  buf1  g6451(.din(new_new_n7392__), .dout(new_new_n7393__));
  buf1  g6452(.din(new_new_n1019__), .dout(new_new_n7394__));
  buf1  g6453(.din(new_new_n7394__), .dout(new_new_n7395__));
  buf1  g6454(.din(new_new_n7394__), .dout(new_new_n7396__));
  buf1  g6455(.din(new_new_n1020__), .dout(new_new_n7397__));
  buf1  g6456(.din(new_new_n7397__), .dout(new_new_n7398__));
  buf1  g6457(.din(new_new_n2604__), .dout(new_new_n7399__));
  buf1  g6458(.din(new_new_n2602__), .dout(new_new_n7400__));
  buf1  g6459(.din(new_new_n2603__), .dout(new_new_n7401__));
  buf1  g6460(.din(new_new_n2601__), .dout(new_new_n7402__));
  buf1  g6461(.din(new_new_n2606__), .dout(new_new_n7403__));
  buf1  g6462(.din(new_new_n7403__), .dout(new_new_n7404__));
  buf1  g6463(.din(new_new_n2605__), .dout(new_new_n7405__));
  buf1  g6464(.din(new_new_n7405__), .dout(new_new_n7406__));
  buf1  g6465(.din(new_new_n1462__), .dout(new_new_n7407__));
  buf1  g6466(.din(new_new_n1414__), .dout(new_new_n7408__));
  buf1  g6467(.din(new_new_n1461__), .dout(new_new_n7409__));
  buf1  g6468(.din(new_new_n1413__), .dout(new_new_n7410__));
  buf1  g6469(.din(new_new_n2614__), .dout(new_new_n7411__));
  buf1  g6470(.din(new_new_n7411__), .dout(new_new_n7412__));
  buf1  g6471(.din(new_new_n2613__), .dout(new_new_n7413__));
  buf1  g6472(.din(new_new_n7413__), .dout(new_new_n7414__));
  buf1  g6473(.din(new_new_n1021__), .dout(new_new_n7415__));
  buf1  g6474(.din(new_new_n7415__), .dout(new_new_n7416__));
  buf1  g6475(.din(new_new_n7415__), .dout(new_new_n7417__));
  buf1  g6476(.din(new_new_n1022__), .dout(new_new_n7418__));
  buf1  g6477(.din(new_new_n7418__), .dout(new_new_n7419__));
  buf1  g6478(.din(new_new_n2622__), .dout(new_new_n7420__));
  buf1  g6479(.din(new_new_n2620__), .dout(new_new_n7421__));
  buf1  g6480(.din(new_new_n2621__), .dout(new_new_n7422__));
  buf1  g6481(.din(new_new_n2619__), .dout(new_new_n7423__));
  buf1  g6482(.din(new_new_n2624__), .dout(new_new_n7424__));
  buf1  g6483(.din(new_new_n7424__), .dout(new_new_n7425__));
  buf1  g6484(.din(new_new_n2623__), .dout(new_new_n7426__));
  buf1  g6485(.din(new_new_n7426__), .dout(new_new_n7427__));
  buf1  g6486(.din(new_new_n2626__), .dout(new_new_n7428__));
  buf1  g6487(.din(new_new_n2612__), .dout(new_new_n7429__));
  buf1  g6488(.din(new_new_n2625__), .dout(new_new_n7430__));
  buf1  g6489(.din(new_new_n2611__), .dout(new_new_n7431__));
  buf1  g6490(.din(new_new_n2628__), .dout(new_new_n7432__));
  buf1  g6491(.din(new_new_n7432__), .dout(new_new_n7433__));
  buf1  g6492(.din(new_new_n2627__), .dout(new_new_n7434__));
  buf1  g6493(.din(new_new_n7434__), .dout(new_new_n7435__));
  buf1  g6494(.din(new_new_n2636__), .dout(new_new_n7436__));
  buf1  g6495(.din(new_new_n2634__), .dout(new_new_n7437__));
  buf1  g6496(.din(new_new_n2635__), .dout(new_new_n7438__));
  buf1  g6497(.din(new_new_n2633__), .dout(new_new_n7439__));
  buf1  g6498(.din(new_new_n2638__), .dout(new_new_n7440__));
  buf1  g6499(.din(new_new_n7440__), .dout(new_new_n7441__));
  buf1  g6500(.din(new_new_n2637__), .dout(new_new_n7442__));
  buf1  g6501(.din(new_new_n7442__), .dout(new_new_n7443__));
  buf1  g6502(.din(new_new_n1023__), .dout(new_new_n7444__));
  buf1  g6503(.din(new_new_n7444__), .dout(new_new_n7445__));
  buf1  g6504(.din(new_new_n1024__), .dout(new_new_n7446__));
  buf1  g6505(.din(new_new_n7446__), .dout(new_new_n7447__));
  buf1  g6506(.din(new_new_n7446__), .dout(new_new_n7448__));
  buf1  g6507(.din(new_new_n2654__), .dout(new_new_n7449__));
  buf1  g6508(.din(new_new_n2652__), .dout(new_new_n7450__));
  buf1  g6509(.din(new_new_n2653__), .dout(new_new_n7451__));
  buf1  g6510(.din(new_new_n2651__), .dout(new_new_n7452__));
  buf1  g6511(.din(new_new_n2656__), .dout(new_new_n7453__));
  buf1  g6512(.din(new_new_n7453__), .dout(new_new_n7454__));
  buf1  g6513(.din(new_new_n2655__), .dout(new_new_n7455__));
  buf1  g6514(.din(new_new_n7455__), .dout(new_new_n7456__));
  buf1  g6515(.din(new_new_n2658__), .dout(new_new_n7457__));
  buf1  g6516(.din(new_new_n2650__), .dout(new_new_n7458__));
  buf1  g6517(.din(new_new_n2657__), .dout(new_new_n7459__));
  buf1  g6518(.din(new_new_n2649__), .dout(new_new_n7460__));
  buf1  g6519(.din(new_new_n2660__), .dout(new_new_n7461__));
  buf1  g6520(.din(new_new_n7461__), .dout(new_new_n7462__));
  buf1  g6521(.din(new_new_n2659__), .dout(new_new_n7463__));
  buf1  g6522(.din(new_new_n7463__), .dout(new_new_n7464__));
  buf1  g6523(.din(new_new_n2668__), .dout(new_new_n7465__));
  buf1  g6524(.din(new_new_n2666__), .dout(new_new_n7466__));
  buf1  g6525(.din(new_new_n2667__), .dout(new_new_n7467__));
  buf1  g6526(.din(new_new_n2665__), .dout(new_new_n7468__));
  buf1  g6527(.din(new_new_n2670__), .dout(new_new_n7469__));
  buf1  g6528(.din(new_new_n7469__), .dout(new_new_n7470__));
  buf1  g6529(.din(new_new_n2669__), .dout(new_new_n7471__));
  buf1  g6530(.din(new_new_n7471__), .dout(new_new_n7472__));
  buf1  g6531(.din(new_new_n2672__), .dout(new_new_n7473__));
  buf1  g6532(.din(new_new_n2644__), .dout(new_new_n7474__));
  buf1  g6533(.din(new_new_n2671__), .dout(new_new_n7475__));
  buf1  g6534(.din(new_new_n2643__), .dout(new_new_n7476__));
  buf1  g6535(.din(new_new_n2674__), .dout(new_new_n7477__));
  buf1  g6536(.din(new_new_n7477__), .dout(new_new_n7478__));
  buf1  g6537(.din(new_new_n2673__), .dout(new_new_n7479__));
  buf1  g6538(.din(new_new_n7479__), .dout(new_new_n7480__));
  buf1  g6539(.din(new_new_n2682__), .dout(new_new_n7481__));
  buf1  g6540(.din(new_new_n2680__), .dout(new_new_n7482__));
  buf1  g6541(.din(new_new_n2681__), .dout(new_new_n7483__));
  buf1  g6542(.din(new_new_n2679__), .dout(new_new_n7484__));
  buf1  g6543(.din(new_new_n2684__), .dout(new_new_n7485__));
  buf1  g6544(.din(new_new_n7485__), .dout(new_new_n7486__));
  buf1  g6545(.din(new_new_n2683__), .dout(new_new_n7487__));
  buf1  g6546(.din(new_new_n7487__), .dout(new_new_n7488__));
  buf1  g6547(.din(new_new_n1446__), .dout(new_new_n7489__));
  buf1  g6548(.din(new_new_n7489__), .dout(new_new_n7490__));
  buf1  g6549(.din(new_new_n1445__), .dout(new_new_n7491__));
  buf1  g6550(.din(new_new_n7491__), .dout(new_new_n7492__));
  buf1  g6551(.din(new_new_n2704__), .dout(new_new_n7493__));
  buf1  g6552(.din(new_new_n2702__), .dout(new_new_n7494__));
  buf1  g6553(.din(new_new_n2703__), .dout(new_new_n7495__));
  buf1  g6554(.din(new_new_n2701__), .dout(new_new_n7496__));
  buf1  g6555(.din(new_new_n2706__), .dout(new_new_n7497__));
  buf1  g6556(.din(new_new_n7497__), .dout(new_new_n7498__));
  buf1  g6557(.din(new_new_n2705__), .dout(new_new_n7499__));
  buf1  g6558(.din(new_new_n7499__), .dout(new_new_n7500__));
  buf1  g6559(.din(new_new_n1025__), .dout(new_new_n7501__));
  buf1  g6560(.din(new_new_n7501__), .dout(new_new_n7502__));
  buf1  g6561(.din(new_new_n1026__), .dout(new_new_n7503__));
  buf1  g6562(.din(new_new_n7503__), .dout(new_new_n7504__));
  buf1  g6563(.din(new_new_n2714__), .dout(new_new_n7505__));
  buf1  g6564(.din(new_new_n2712__), .dout(new_new_n7506__));
  buf1  g6565(.din(new_new_n2713__), .dout(new_new_n7507__));
  buf1  g6566(.din(new_new_n2711__), .dout(new_new_n7508__));
  buf1  g6567(.din(new_new_n2716__), .dout(new_new_n7509__));
  buf1  g6568(.din(new_new_n7509__), .dout(new_new_n7510__));
  buf1  g6569(.din(new_new_n2715__), .dout(new_new_n7511__));
  buf1  g6570(.din(new_new_n7511__), .dout(new_new_n7512__));
  buf1  g6571(.din(new_new_n2718__), .dout(new_new_n7513__));
  buf1  g6572(.din(new_new_n2696__), .dout(new_new_n7514__));
  buf1  g6573(.din(new_new_n2717__), .dout(new_new_n7515__));
  buf1  g6574(.din(new_new_n2695__), .dout(new_new_n7516__));
  buf1  g6575(.din(new_new_n2720__), .dout(new_new_n7517__));
  buf1  g6576(.din(new_new_n7517__), .dout(new_new_n7518__));
  buf1  g6577(.din(new_new_n2719__), .dout(new_new_n7519__));
  buf1  g6578(.din(new_new_n7519__), .dout(new_new_n7520__));
  buf1  g6579(.din(new_new_n2728__), .dout(new_new_n7521__));
  buf1  g6580(.din(new_new_n2726__), .dout(new_new_n7522__));
  buf1  g6581(.din(new_new_n2727__), .dout(new_new_n7523__));
  buf1  g6582(.din(new_new_n2725__), .dout(new_new_n7524__));
  buf1  g6583(.din(new_new_n2730__), .dout(new_new_n7525__));
  buf1  g6584(.din(new_new_n7525__), .dout(new_new_n7526__));
  buf1  g6585(.din(new_new_n2729__), .dout(new_new_n7527__));
  buf1  g6586(.din(new_new_n7527__), .dout(new_new_n7528__));
  buf1  g6587(.din(new_new_n2732__), .dout(new_new_n7529__));
  buf1  g6588(.din(new_new_n2690__), .dout(new_new_n7530__));
  buf1  g6589(.din(new_new_n2731__), .dout(new_new_n7531__));
  buf1  g6590(.din(new_new_n2689__), .dout(new_new_n7532__));
  buf1  g6591(.din(new_new_n1464__), .dout(new_new_n7533__));
  buf1  g6592(.din(new_new_n1416__), .dout(new_new_n7534__));
  buf1  g6593(.din(new_new_n1463__), .dout(new_new_n7535__));
  buf1  g6594(.din(new_new_n1415__), .dout(new_new_n7536__));
  buf1  g6595(.din(new_new_n2736__), .dout(new_new_n7537__));
  buf1  g6596(.din(new_new_n7537__), .dout(new_new_n7538__));
  buf1  g6597(.din(new_new_n2735__), .dout(new_new_n7539__));
  buf1  g6598(.din(new_new_n7539__), .dout(new_new_n7540__));
  buf1  g6599(.din(new_new_n1033__), .dout(new_new_n7541__));
  buf1  g6600(.din(new_new_n7541__), .dout(new_new_n7542__));
  buf1  g6601(.din(new_new_n1034__), .dout(new_new_n7543__));
  buf1  g6602(.din(new_new_n7543__), .dout(new_new_n7544__));
  buf1  g6603(.din(new_new_n2744__), .dout(new_new_n7545__));
  buf1  g6604(.din(new_new_n2742__), .dout(new_new_n7546__));
  buf1  g6605(.din(new_new_n2743__), .dout(new_new_n7547__));
  buf1  g6606(.din(new_new_n2741__), .dout(new_new_n7548__));
  buf1  g6607(.din(new_new_n2746__), .dout(new_new_n7549__));
  buf1  g6608(.din(new_new_n7549__), .dout(new_new_n7550__));
  buf1  g6609(.din(new_new_n2745__), .dout(new_new_n7551__));
  buf1  g6610(.din(new_new_n7551__), .dout(new_new_n7552__));
  buf1  g6611(.din(new_new_n2754__), .dout(new_new_n7553__));
  buf1  g6612(.din(new_new_n2752__), .dout(new_new_n7554__));
  buf1  g6613(.din(new_new_n2753__), .dout(new_new_n7555__));
  buf1  g6614(.din(new_new_n2751__), .dout(new_new_n7556__));
  buf1  g6615(.din(new_new_n2756__), .dout(new_new_n7557__));
  buf1  g6616(.din(new_new_n7557__), .dout(new_new_n7558__));
  buf1  g6617(.din(new_new_n2755__), .dout(new_new_n7559__));
  buf1  g6618(.din(new_new_n7559__), .dout(new_new_n7560__));
  buf1  g6619(.din(new_new_n2764__), .dout(new_new_n7561__));
  buf1  g6620(.din(new_new_n2762__), .dout(new_new_n7562__));
  buf1  g6621(.din(new_new_n2763__), .dout(new_new_n7563__));
  buf1  g6622(.din(new_new_n2761__), .dout(new_new_n7564__));
  buf1  g6623(.din(new_new_n2766__), .dout(new_new_n7565__));
  buf1  g6624(.din(new_new_n7565__), .dout(new_new_n7566__));
  buf1  g6625(.din(new_new_n2765__), .dout(new_new_n7567__));
  buf1  g6626(.din(new_new_n7567__), .dout(new_new_n7568__));
  buf1  g6627(.din(new_new_n2774__), .dout(new_new_n7569__));
  buf1  g6628(.din(new_new_n2772__), .dout(new_new_n7570__));
  buf1  g6629(.din(new_new_n2773__), .dout(new_new_n7571__));
  buf1  g6630(.din(new_new_n2771__), .dout(new_new_n7572__));
  buf1  g6631(.din(new_new_n2776__), .dout(new_new_n7573__));
  buf1  g6632(.din(new_new_n7573__), .dout(new_new_n7574__));
  buf1  g6633(.din(new_new_n2775__), .dout(new_new_n7575__));
  buf1  g6634(.din(new_new_n7575__), .dout(new_new_n7576__));
  buf1  g6635(.din(new_new_n2784__), .dout(new_new_n7577__));
  buf1  g6636(.din(new_new_n2782__), .dout(new_new_n7578__));
  buf1  g6637(.din(new_new_n2783__), .dout(new_new_n7579__));
  buf1  g6638(.din(new_new_n2781__), .dout(new_new_n7580__));
  buf1  g6639(.din(new_new_n2786__), .dout(new_new_n7581__));
  buf1  g6640(.din(new_new_n7581__), .dout(new_new_n7582__));
  buf1  g6641(.din(new_new_n2785__), .dout(new_new_n7583__));
  buf1  g6642(.din(new_new_n7583__), .dout(new_new_n7584__));
  buf1  g6643(.din(new_new_n2243__), .dout(new_new_n7585__));
  buf1  g6644(.din(new_new_n2794__), .dout(new_new_n7586__));
  buf1  g6645(.din(new_new_n2792__), .dout(new_new_n7587__));
  buf1  g6646(.din(new_new_n2796__), .dout(new_new_n7588__));
  buf1  g6647(.din(new_new_n2350__), .dout(new_new_n7589__));
  buf1  g6648(.din(new_new_n2323__), .dout(new_new_n7590__));
  buf1  g6649(.din(new_new_n909__), .dout(new_new_n7591__));
  buf1  g6650(.din(new_new_n7591__), .dout(new_new_n7592__));
  buf1  g6651(.din(new_new_n7592__), .dout(new_new_n7593__));
  buf1  g6652(.din(new_new_n7593__), .dout(new_new_n7594__));
  buf1  g6653(.din(new_new_n7593__), .dout(new_new_n7595__));
  buf1  g6654(.din(new_new_n7592__), .dout(new_new_n7596__));
  buf1  g6655(.din(new_new_n7596__), .dout(new_new_n7597__));
  buf1  g6656(.din(new_new_n7596__), .dout(new_new_n7598__));
  buf1  g6657(.din(new_new_n7591__), .dout(new_new_n7599__));
  buf1  g6658(.din(new_new_n7599__), .dout(new_new_n7600__));
  buf1  g6659(.din(new_new_n7600__), .dout(new_new_n7601__));
  buf1  g6660(.din(new_new_n7600__), .dout(new_new_n7602__));
  buf1  g6661(.din(new_new_n7599__), .dout(new_new_n7603__));
  buf1  g6662(.din(new_new_n910__), .dout(new_new_n7604__));
  buf1  g6663(.din(new_new_n7604__), .dout(new_new_n7605__));
  buf1  g6664(.din(new_new_n7605__), .dout(new_new_n7606__));
  buf1  g6665(.din(new_new_n7606__), .dout(new_new_n7607__));
  buf1  g6666(.din(new_new_n7606__), .dout(new_new_n7608__));
  buf1  g6667(.din(new_new_n7605__), .dout(new_new_n7609__));
  buf1  g6668(.din(new_new_n7609__), .dout(new_new_n7610__));
  buf1  g6669(.din(new_new_n7609__), .dout(new_new_n7611__));
  buf1  g6670(.din(new_new_n7604__), .dout(new_new_n7612__));
  buf1  g6671(.din(new_new_n7612__), .dout(new_new_n7613__));
  buf1  g6672(.din(new_new_n7613__), .dout(new_new_n7614__));
  buf1  g6673(.din(new_new_n7613__), .dout(new_new_n7615__));
  buf1  g6674(.din(new_new_n7612__), .dout(new_new_n7616__));
  buf1  g6675(.din(new_new_n1530__), .dout(new_new_n7617__));
  buf1  g6676(.din(new_new_n7617__), .dout(new_new_n7618__));
  buf1  g6677(.din(new_new_n1529__), .dout(new_new_n7619__));
  buf1  g6678(.din(new_new_n7619__), .dout(new_new_n7620__));
  buf1  g6679(.din(new_new_n2811__), .dout(new_new_n7621__));
  buf1  g6680(.din(new_new_n2809__), .dout(new_new_n7622__));
  buf1  g6681(.din(new_new_n2810__), .dout(new_new_n7623__));
  buf1  g6682(.din(new_new_n2808__), .dout(new_new_n7624__));
  buf1  g6683(.din(new_new_n2813__), .dout(new_new_n7625__));
  buf1  g6684(.din(new_new_n7625__), .dout(new_new_n7626__));
  buf1  g6685(.din(new_new_n2812__), .dout(new_new_n7627__));
  buf1  g6686(.din(new_new_n7627__), .dout(new_new_n7628__));
  buf1  g6687(.din(new_new_n1131__), .dout(new_new_n7629__));
  buf1  g6688(.din(new_new_n7629__), .dout(new_new_n7630__));
  buf1  g6689(.din(new_new_n7630__), .dout(new_new_n7631__));
  buf1  g6690(.din(new_new_n7629__), .dout(new_new_n7632__));
  buf1  g6691(.din(new_new_n1132__), .dout(new_new_n7633__));
  buf1  g6692(.din(new_new_n7633__), .dout(new_new_n7634__));
  buf1  g6693(.din(new_new_n7634__), .dout(new_new_n7635__));
  buf1  g6694(.din(new_new_n7633__), .dout(new_new_n7636__));
  buf1  g6695(.din(new_new_n2821__), .dout(new_new_n7637__));
  buf1  g6696(.din(new_new_n2819__), .dout(new_new_n7638__));
  buf1  g6697(.din(new_new_n2820__), .dout(new_new_n7639__));
  buf1  g6698(.din(new_new_n2818__), .dout(new_new_n7640__));
  buf1  g6699(.din(new_new_n2823__), .dout(new_new_n7641__));
  buf1  g6700(.din(new_new_n7641__), .dout(new_new_n7642__));
  buf1  g6701(.din(new_new_n2822__), .dout(new_new_n7643__));
  buf1  g6702(.din(new_new_n7643__), .dout(new_new_n7644__));
  buf1  g6703(.din(new_new_n2831__), .dout(new_new_n7645__));
  buf1  g6704(.din(new_new_n2829__), .dout(new_new_n7646__));
  buf1  g6705(.din(new_new_n2830__), .dout(new_new_n7647__));
  buf1  g6706(.din(new_new_n2828__), .dout(new_new_n7648__));
  buf1  g6707(.din(new_new_n2833__), .dout(new_new_n7649__));
  buf1  g6708(.din(new_new_n7649__), .dout(new_new_n7650__));
  buf1  g6709(.din(new_new_n2832__), .dout(new_new_n7651__));
  buf1  g6710(.din(new_new_n7651__), .dout(new_new_n7652__));
  buf1  g6711(.din(new_new_n2841__), .dout(new_new_n7653__));
  buf1  g6712(.din(new_new_n2839__), .dout(new_new_n7654__));
  buf1  g6713(.din(new_new_n2840__), .dout(new_new_n7655__));
  buf1  g6714(.din(new_new_n2838__), .dout(new_new_n7656__));
  buf1  g6715(.din(new_new_n2843__), .dout(new_new_n7657__));
  buf1  g6716(.din(new_new_n7657__), .dout(new_new_n7658__));
  buf1  g6717(.din(new_new_n2842__), .dout(new_new_n7659__));
  buf1  g6718(.din(new_new_n7659__), .dout(new_new_n7660__));
  buf1  g6719(.din(new_new_n2321__), .dout(new_new_n7661__));
  buf1  g6720(.din(new_new_n2851__), .dout(new_new_n7662__));
  buf1  g6721(.din(new_new_n2849__), .dout(new_new_n7663__));
  buf1  g6722(.din(new_new_n2850__), .dout(new_new_n7664__));
  buf1  g6723(.din(new_new_n2848__), .dout(new_new_n7665__));
  buf1  g6724(.din(new_new_n2853__), .dout(new_new_n7666__));
  buf1  g6725(.din(new_new_n7666__), .dout(new_new_n7667__));
  buf1  g6726(.din(new_new_n2852__), .dout(new_new_n7668__));
  buf1  g6727(.din(new_new_n7668__), .dout(new_new_n7669__));
  buf1  g6728(.din(new_new_n1615__), .dout(new_new_n7670__));
  buf1  g6729(.din(new_new_n7670__), .dout(new_new_n7671__));
  buf1  g6730(.din(new_new_n7671__), .dout(new_new_n7672__));
  buf1  g6731(.din(new_new_n7672__), .dout(new_new_n7673__));
  buf1  g6732(.din(new_new_n7672__), .dout(new_new_n7674__));
  buf1  g6733(.din(new_new_n7671__), .dout(new_new_n7675__));
  buf1  g6734(.din(new_new_n7675__), .dout(new_new_n7676__));
  buf1  g6735(.din(new_new_n7675__), .dout(new_new_n7677__));
  buf1  g6736(.din(new_new_n7670__), .dout(new_new_n7678__));
  buf1  g6737(.din(new_new_n7678__), .dout(new_new_n7679__));
  buf1  g6738(.din(new_new_n7679__), .dout(new_new_n7680__));
  buf1  g6739(.din(new_new_n7679__), .dout(new_new_n7681__));
  buf1  g6740(.din(new_new_n7678__), .dout(new_new_n7682__));
  buf1  g6741(.din(new_new_n7682__), .dout(new_new_n7683__));
  buf1  g6742(.din(new_new_n7682__), .dout(new_new_n7684__));
  buf1  g6743(.din(new_new_n1616__), .dout(new_new_n7685__));
  buf1  g6744(.din(new_new_n7685__), .dout(new_new_n7686__));
  buf1  g6745(.din(new_new_n7686__), .dout(new_new_n7687__));
  buf1  g6746(.din(new_new_n7687__), .dout(new_new_n7688__));
  buf1  g6747(.din(new_new_n7687__), .dout(new_new_n7689__));
  buf1  g6748(.din(new_new_n7686__), .dout(new_new_n7690__));
  buf1  g6749(.din(new_new_n7690__), .dout(new_new_n7691__));
  buf1  g6750(.din(new_new_n7690__), .dout(new_new_n7692__));
  buf1  g6751(.din(new_new_n7685__), .dout(new_new_n7693__));
  buf1  g6752(.din(new_new_n7693__), .dout(new_new_n7694__));
  buf1  g6753(.din(new_new_n7694__), .dout(new_new_n7695__));
  buf1  g6754(.din(new_new_n7694__), .dout(new_new_n7696__));
  buf1  g6755(.din(new_new_n7693__), .dout(new_new_n7697__));
  buf1  g6756(.din(new_new_n7697__), .dout(new_new_n7698__));
  buf1  g6757(.din(new_new_n7697__), .dout(new_new_n7699__));
  buf1  g6758(.din(new_new_n2859__), .dout(new_new_n7700__));
  buf1  g6759(.din(new_new_n2802__), .dout(new_new_n7701__));
  buf1  g6760(.din(new_new_n1303__), .dout(new_new_n7702__));
  buf1  g6761(.din(new_new_n7702__), .dout(new_new_n7703__));
  buf1  g6762(.din(new_new_n7703__), .dout(new_new_n7704__));
  buf1  g6763(.din(new_new_n7703__), .dout(new_new_n7705__));
  buf1  g6764(.din(new_new_n7702__), .dout(new_new_n7706__));
  buf1  g6765(.din(new_new_n7706__), .dout(new_new_n7707__));
  buf1  g6766(.din(new_new_n1304__), .dout(new_new_n7708__));
  buf1  g6767(.din(new_new_n7708__), .dout(new_new_n7709__));
  buf1  g6768(.din(new_new_n7709__), .dout(new_new_n7710__));
  buf1  g6769(.din(new_new_n7708__), .dout(new_new_n7711__));
  buf1  g6770(.din(new_new_n2867__), .dout(new_new_n7712__));
  buf1  g6771(.din(new_new_n2865__), .dout(new_new_n7713__));
  buf1  g6772(.din(new_new_n2866__), .dout(new_new_n7714__));
  buf1  g6773(.din(new_new_n2864__), .dout(new_new_n7715__));
  buf1  g6774(.din(new_new_n2869__), .dout(new_new_n7716__));
  buf1  g6775(.din(new_new_n7716__), .dout(new_new_n7717__));
  buf1  g6776(.din(new_new_n2868__), .dout(new_new_n7718__));
  buf1  g6777(.din(new_new_n7718__), .dout(new_new_n7719__));
  buf1  g6778(.din(new_new_n2877__), .dout(new_new_n7720__));
  buf1  g6779(.din(new_new_n2875__), .dout(new_new_n7721__));
  buf1  g6780(.din(new_new_n2876__), .dout(new_new_n7722__));
  buf1  g6781(.din(new_new_n2874__), .dout(new_new_n7723__));
  buf1  g6782(.din(new_new_n2879__), .dout(new_new_n7724__));
  buf1  g6783(.din(new_new_n7724__), .dout(new_new_n7725__));
  buf1  g6784(.din(new_new_n2878__), .dout(new_new_n7726__));
  buf1  g6785(.din(new_new_n7726__), .dout(new_new_n7727__));
  buf1  g6786(.din(new_new_n2887__), .dout(new_new_n7728__));
  buf1  g6787(.din(new_new_n2885__), .dout(new_new_n7729__));
  buf1  g6788(.din(new_new_n2886__), .dout(new_new_n7730__));
  buf1  g6789(.din(new_new_n2884__), .dout(new_new_n7731__));
  buf1  g6790(.din(new_new_n2889__), .dout(new_new_n7732__));
  buf1  g6791(.din(new_new_n7732__), .dout(new_new_n7733__));
  buf1  g6792(.din(new_new_n2888__), .dout(new_new_n7734__));
  buf1  g6793(.din(new_new_n7734__), .dout(new_new_n7735__));
  buf1  g6794(.din(new_new_n2800__), .dout(new_new_n7736__));
  buf1  g6795(.din(new_new_n2897__), .dout(new_new_n7737__));
  buf1  g6796(.din(new_new_n2895__), .dout(new_new_n7738__));
  buf1  g6797(.din(new_new_n2896__), .dout(new_new_n7739__));
  buf1  g6798(.din(new_new_n2894__), .dout(new_new_n7740__));
  buf1  g6799(.din(new_new_n2899__), .dout(new_new_n7741__));
  buf1  g6800(.din(new_new_n7741__), .dout(new_new_n7742__));
  buf1  g6801(.din(new_new_n2898__), .dout(new_new_n7743__));
  buf1  g6802(.din(new_new_n7743__), .dout(new_new_n7744__));
  buf1  g6803(.din(new_new_n2905__), .dout(new_new_n7745__));
  buf1  g6804(.din(new_new_n2860__), .dout(new_new_n7746__));
  buf1  g6805(.din(new_new_n2799__), .dout(new_new_n7747__));
  buf1  g6806(.din(new_new_n7747__), .dout(new_new_n7748__));
  buf1  g6807(.din(new_new_n2921__), .dout(new_new_n7749__));
  buf1  g6808(.din(new_new_n2919__), .dout(new_new_n7750__));
  buf1  g6809(.din(new_new_n2920__), .dout(new_new_n7751__));
  buf1  g6810(.din(new_new_n2918__), .dout(new_new_n7752__));
  buf1  g6811(.din(new_new_n2923__), .dout(new_new_n7753__));
  buf1  g6812(.din(new_new_n7753__), .dout(new_new_n7754__));
  buf1  g6813(.din(new_new_n2922__), .dout(new_new_n7755__));
  buf1  g6814(.din(new_new_n7755__), .dout(new_new_n7756__));
  buf1  g6815(.din(new_new_n2931__), .dout(new_new_n7757__));
  buf1  g6816(.din(new_new_n2929__), .dout(new_new_n7758__));
  buf1  g6817(.din(new_new_n2930__), .dout(new_new_n7759__));
  buf1  g6818(.din(new_new_n2928__), .dout(new_new_n7760__));
  buf1  g6819(.din(new_new_n2933__), .dout(new_new_n7761__));
  buf1  g6820(.din(new_new_n7761__), .dout(new_new_n7762__));
  buf1  g6821(.din(new_new_n2932__), .dout(new_new_n7763__));
  buf1  g6822(.din(new_new_n7763__), .dout(new_new_n7764__));
  buf1  g6823(.din(new_new_n2941__), .dout(new_new_n7765__));
  buf1  g6824(.din(new_new_n2939__), .dout(new_new_n7766__));
  buf1  g6825(.din(new_new_n2940__), .dout(new_new_n7767__));
  buf1  g6826(.din(new_new_n2938__), .dout(new_new_n7768__));
  buf1  g6827(.din(new_new_n2943__), .dout(new_new_n7769__));
  buf1  g6828(.din(new_new_n7769__), .dout(new_new_n7770__));
  buf1  g6829(.din(new_new_n2942__), .dout(new_new_n7771__));
  buf1  g6830(.din(new_new_n7771__), .dout(new_new_n7772__));
  buf1  g6831(.din(new_new_n2951__), .dout(new_new_n7773__));
  buf1  g6832(.din(new_new_n2949__), .dout(new_new_n7774__));
  buf1  g6833(.din(new_new_n2950__), .dout(new_new_n7775__));
  buf1  g6834(.din(new_new_n2948__), .dout(new_new_n7776__));
  buf1  g6835(.din(new_new_n2953__), .dout(new_new_n7777__));
  buf1  g6836(.din(new_new_n7777__), .dout(new_new_n7778__));
  buf1  g6837(.din(new_new_n2952__), .dout(new_new_n7779__));
  buf1  g6838(.din(new_new_n7779__), .dout(new_new_n7780__));
  buf1  g6839(.din(new_new_n2970__), .dout(new_new_n7781__));
  buf1  g6840(.din(new_new_n2968__), .dout(new_new_n7782__));
  buf1  g6841(.din(new_new_n2969__), .dout(new_new_n7783__));
  buf1  g6842(.din(new_new_n2967__), .dout(new_new_n7784__));
  buf1  g6843(.din(new_new_n2972__), .dout(new_new_n7785__));
  buf1  g6844(.din(new_new_n7785__), .dout(new_new_n7786__));
  buf1  g6845(.din(new_new_n2971__), .dout(new_new_n7787__));
  buf1  g6846(.din(new_new_n7787__), .dout(new_new_n7788__));
  buf1  g6847(.din(new_new_n2980__), .dout(new_new_n7789__));
  buf1  g6848(.din(new_new_n2978__), .dout(new_new_n7790__));
  buf1  g6849(.din(new_new_n2979__), .dout(new_new_n7791__));
  buf1  g6850(.din(new_new_n2977__), .dout(new_new_n7792__));
  buf1  g6851(.din(new_new_n2982__), .dout(new_new_n7793__));
  buf1  g6852(.din(new_new_n7793__), .dout(new_new_n7794__));
  buf1  g6853(.din(new_new_n2981__), .dout(new_new_n7795__));
  buf1  g6854(.din(new_new_n7795__), .dout(new_new_n7796__));
  buf1  g6855(.din(new_new_n2990__), .dout(new_new_n7797__));
  buf1  g6856(.din(new_new_n2988__), .dout(new_new_n7798__));
  buf1  g6857(.din(new_new_n2989__), .dout(new_new_n7799__));
  buf1  g6858(.din(new_new_n2987__), .dout(new_new_n7800__));
  buf1  g6859(.din(new_new_n2992__), .dout(new_new_n7801__));
  buf1  g6860(.din(new_new_n7801__), .dout(new_new_n7802__));
  buf1  g6861(.din(new_new_n2991__), .dout(new_new_n7803__));
  buf1  g6862(.din(new_new_n7803__), .dout(new_new_n7804__));
  buf1  g6863(.din(new_new_n3000__), .dout(new_new_n7805__));
  buf1  g6864(.din(new_new_n2998__), .dout(new_new_n7806__));
  buf1  g6865(.din(new_new_n2999__), .dout(new_new_n7807__));
  buf1  g6866(.din(new_new_n2997__), .dout(new_new_n7808__));
  buf1  g6867(.din(new_new_n3002__), .dout(new_new_n7809__));
  buf1  g6868(.din(new_new_n7809__), .dout(new_new_n7810__));
  buf1  g6869(.din(new_new_n3001__), .dout(new_new_n7811__));
  buf1  g6870(.din(new_new_n7811__), .dout(new_new_n7812__));
  buf1  g6871(.din(new_new_n3025__), .dout(new_new_n7813__));
  buf1  g6872(.din(new_new_n3023__), .dout(new_new_n7814__));
  buf1  g6873(.din(new_new_n3024__), .dout(new_new_n7815__));
  buf1  g6874(.din(new_new_n3022__), .dout(new_new_n7816__));
  buf1  g6875(.din(new_new_n3027__), .dout(new_new_n7817__));
  buf1  g6876(.din(new_new_n7817__), .dout(new_new_n7818__));
  buf1  g6877(.din(new_new_n3026__), .dout(new_new_n7819__));
  buf1  g6878(.din(new_new_n7819__), .dout(new_new_n7820__));
  buf1  g6879(.din(new_new_n1029__), .dout(new_new_n7821__));
  buf1  g6880(.din(new_new_n7821__), .dout(new_new_n7822__));
  buf1  g6881(.din(new_new_n1030__), .dout(new_new_n7823__));
  buf1  g6882(.din(new_new_n7823__), .dout(new_new_n7824__));
  buf1  g6883(.din(new_new_n3035__), .dout(new_new_n7825__));
  buf1  g6884(.din(new_new_n3033__), .dout(new_new_n7826__));
  buf1  g6885(.din(new_new_n3034__), .dout(new_new_n7827__));
  buf1  g6886(.din(new_new_n3032__), .dout(new_new_n7828__));
  buf1  g6887(.din(new_new_n3037__), .dout(new_new_n7829__));
  buf1  g6888(.din(new_new_n7829__), .dout(new_new_n7830__));
  buf1  g6889(.din(new_new_n3036__), .dout(new_new_n7831__));
  buf1  g6890(.din(new_new_n7831__), .dout(new_new_n7832__));
  buf1  g6891(.din(new_new_n3039__), .dout(new_new_n7833__));
  buf1  g6892(.din(new_new_n3017__), .dout(new_new_n7834__));
  buf1  g6893(.din(new_new_n3038__), .dout(new_new_n7835__));
  buf1  g6894(.din(new_new_n3016__), .dout(new_new_n7836__));
  buf1  g6895(.din(new_new_n3041__), .dout(new_new_n7837__));
  buf1  g6896(.din(new_new_n7837__), .dout(new_new_n7838__));
  buf1  g6897(.din(new_new_n3040__), .dout(new_new_n7839__));
  buf1  g6898(.din(new_new_n7839__), .dout(new_new_n7840__));
  buf1  g6899(.din(new_new_n3049__), .dout(new_new_n7841__));
  buf1  g6900(.din(new_new_n3047__), .dout(new_new_n7842__));
  buf1  g6901(.din(new_new_n3048__), .dout(new_new_n7843__));
  buf1  g6902(.din(new_new_n3046__), .dout(new_new_n7844__));
  buf1  g6903(.din(new_new_n3051__), .dout(new_new_n7845__));
  buf1  g6904(.din(new_new_n7845__), .dout(new_new_n7846__));
  buf1  g6905(.din(new_new_n3050__), .dout(new_new_n7847__));
  buf1  g6906(.din(new_new_n7847__), .dout(new_new_n7848__));
  buf1  g6907(.din(new_new_n3065__), .dout(new_new_n7849__));
  buf1  g6908(.din(new_new_n3063__), .dout(new_new_n7850__));
  buf1  g6909(.din(new_new_n3064__), .dout(new_new_n7851__));
  buf1  g6910(.din(new_new_n3062__), .dout(new_new_n7852__));
  buf1  g6911(.din(new_new_n3067__), .dout(new_new_n7853__));
  buf1  g6912(.din(new_new_n7853__), .dout(new_new_n7854__));
  buf1  g6913(.din(new_new_n3066__), .dout(new_new_n7855__));
  buf1  g6914(.din(new_new_n7855__), .dout(new_new_n7856__));
  buf1  g6915(.din(new_new_n3075__), .dout(new_new_n7857__));
  buf1  g6916(.din(new_new_n3073__), .dout(new_new_n7858__));
  buf1  g6917(.din(new_new_n3074__), .dout(new_new_n7859__));
  buf1  g6918(.din(new_new_n3072__), .dout(new_new_n7860__));
  buf1  g6919(.din(new_new_n3077__), .dout(new_new_n7861__));
  buf1  g6920(.din(new_new_n7861__), .dout(new_new_n7862__));
  buf1  g6921(.din(new_new_n3076__), .dout(new_new_n7863__));
  buf1  g6922(.din(new_new_n7863__), .dout(new_new_n7864__));
  buf1  g6923(.din(new_new_n3079__), .dout(new_new_n7865__));
  buf1  g6924(.din(new_new_n3057__), .dout(new_new_n7866__));
  buf1  g6925(.din(new_new_n3078__), .dout(new_new_n7867__));
  buf1  g6926(.din(new_new_n3056__), .dout(new_new_n7868__));
  buf1  g6927(.din(new_new_n3081__), .dout(new_new_n7869__));
  buf1  g6928(.din(new_new_n7869__), .dout(new_new_n7870__));
  buf1  g6929(.din(new_new_n3080__), .dout(new_new_n7871__));
  buf1  g6930(.din(new_new_n7871__), .dout(new_new_n7872__));
  buf1  g6931(.din(new_new_n3089__), .dout(new_new_n7873__));
  buf1  g6932(.din(new_new_n3087__), .dout(new_new_n7874__));
  buf1  g6933(.din(new_new_n3088__), .dout(new_new_n7875__));
  buf1  g6934(.din(new_new_n3086__), .dout(new_new_n7876__));
  buf1  g6935(.din(new_new_n3091__), .dout(new_new_n7877__));
  buf1  g6936(.din(new_new_n7877__), .dout(new_new_n7878__));
  buf1  g6937(.din(new_new_n3090__), .dout(new_new_n7879__));
  buf1  g6938(.din(new_new_n7879__), .dout(new_new_n7880__));
  buf1  g6939(.din(new_new_n3105__), .dout(new_new_n7881__));
  buf1  g6940(.din(new_new_n3103__), .dout(new_new_n7882__));
  buf1  g6941(.din(new_new_n3104__), .dout(new_new_n7883__));
  buf1  g6942(.din(new_new_n3102__), .dout(new_new_n7884__));
  buf1  g6943(.din(new_new_n3107__), .dout(new_new_n7885__));
  buf1  g6944(.din(new_new_n7885__), .dout(new_new_n7886__));
  buf1  g6945(.din(new_new_n3106__), .dout(new_new_n7887__));
  buf1  g6946(.din(new_new_n7887__), .dout(new_new_n7888__));
  buf1  g6947(.din(new_new_n3115__), .dout(new_new_n7889__));
  buf1  g6948(.din(new_new_n3113__), .dout(new_new_n7890__));
  buf1  g6949(.din(new_new_n3114__), .dout(new_new_n7891__));
  buf1  g6950(.din(new_new_n3112__), .dout(new_new_n7892__));
  buf1  g6951(.din(new_new_n3117__), .dout(new_new_n7893__));
  buf1  g6952(.din(new_new_n7893__), .dout(new_new_n7894__));
  buf1  g6953(.din(new_new_n3116__), .dout(new_new_n7895__));
  buf1  g6954(.din(new_new_n7895__), .dout(new_new_n7896__));
  buf1  g6955(.din(new_new_n3128__), .dout(new_new_n7897__));
  buf1  g6956(.din(new_new_n3126__), .dout(new_new_n7898__));
  buf1  g6957(.din(new_new_n3130__), .dout(new_new_n7899__));
  buf1  g6958(.din(new_new_n895__), .dout(new_new_n7900__));
  buf1  g6959(.din(new_new_n7900__), .dout(new_new_n7901__));
  buf1  g6960(.din(new_new_n7901__), .dout(new_new_n7902__));
  buf1  g6961(.din(new_new_n7902__), .dout(new_new_n7903__));
  buf1  g6962(.din(new_new_n7902__), .dout(new_new_n7904__));
  buf1  g6963(.din(new_new_n7901__), .dout(new_new_n7905__));
  buf1  g6964(.din(new_new_n7905__), .dout(new_new_n7906__));
  buf1  g6965(.din(new_new_n7905__), .dout(new_new_n7907__));
  buf1  g6966(.din(new_new_n7900__), .dout(new_new_n7908__));
  buf1  g6967(.din(new_new_n7908__), .dout(new_new_n7909__));
  buf1  g6968(.din(new_new_n7909__), .dout(new_new_n7910__));
  buf1  g6969(.din(new_new_n7909__), .dout(new_new_n7911__));
  buf1  g6970(.din(new_new_n7908__), .dout(new_new_n7912__));
  buf1  g6971(.din(new_new_n7912__), .dout(new_new_n7913__));
  buf1  g6972(.din(new_new_n7912__), .dout(new_new_n7914__));
  buf1  g6973(.din(new_new_n896__), .dout(new_new_n7915__));
  buf1  g6974(.din(new_new_n7915__), .dout(new_new_n7916__));
  buf1  g6975(.din(new_new_n7916__), .dout(new_new_n7917__));
  buf1  g6976(.din(new_new_n7917__), .dout(new_new_n7918__));
  buf1  g6977(.din(new_new_n7917__), .dout(new_new_n7919__));
  buf1  g6978(.din(new_new_n7916__), .dout(new_new_n7920__));
  buf1  g6979(.din(new_new_n7920__), .dout(new_new_n7921__));
  buf1  g6980(.din(new_new_n7920__), .dout(new_new_n7922__));
  buf1  g6981(.din(new_new_n7915__), .dout(new_new_n7923__));
  buf1  g6982(.din(new_new_n7923__), .dout(new_new_n7924__));
  buf1  g6983(.din(new_new_n7924__), .dout(new_new_n7925__));
  buf1  g6984(.din(new_new_n7924__), .dout(new_new_n7926__));
  buf1  g6985(.din(new_new_n7923__), .dout(new_new_n7927__));
  buf1  g6986(.din(new_new_n7927__), .dout(new_new_n7928__));
  buf1  g6987(.din(new_new_n7927__), .dout(new_new_n7929__));
  buf1  g6988(.din(new_new_n2734__), .dout(new_new_n7930__));
  buf1  g6989(.din(new_new_n7930__), .dout(new_new_n7931__));
  buf1  g6990(.din(new_new_n2733__), .dout(new_new_n7932__));
  buf1  g6991(.din(new_new_n2586__), .dout(new_new_n7933__));
  buf1  g6992(.din(new_new_n7933__), .dout(new_new_n7934__));
  buf1  g6993(.din(new_new_n2585__), .dout(new_new_n7935__));
  buf1  g6994(.din(new_new_n2438__), .dout(new_new_n7936__));
  buf1  g6995(.din(new_new_n7936__), .dout(new_new_n7937__));
  buf1  g6996(.din(new_new_n2437__), .dout(new_new_n7938__));
  buf1  g6997(.din(new_new_n3133__), .dout(new_new_n7939__));
  buf1  g6998(.din(new_new_n2908__), .dout(new_new_n7940__));
  buf1  g6999(.din(new_new_n1089__), .dout(new_new_n7941__));
  buf1  g7000(.din(new_new_n7941__), .dout(new_new_n7942__));
  buf1  g7001(.din(new_new_n7941__), .dout(new_new_n7943__));
  buf1  g7002(.din(new_new_n1090__), .dout(new_new_n7944__));
  buf1  g7003(.din(new_new_n7944__), .dout(new_new_n7945__));
  buf1  g7004(.din(new_new_n1494__), .dout(new_new_n7946__));
  buf1  g7005(.din(new_new_n1484__), .dout(new_new_n7947__));
  buf1  g7006(.din(new_new_n1493__), .dout(new_new_n7948__));
  buf1  g7007(.din(new_new_n1483__), .dout(new_new_n7949__));
  buf1  g7008(.din(new_new_n3167__), .dout(new_new_n7950__));
  buf1  g7009(.din(new_new_n7950__), .dout(new_new_n7951__));
  buf1  g7010(.din(new_new_n3166__), .dout(new_new_n7952__));
  buf1  g7011(.din(new_new_n7952__), .dout(new_new_n7953__));
  buf1  g7012(.din(new_new_n1093__), .dout(new_new_n7954__));
  buf1  g7013(.din(new_new_n7954__), .dout(new_new_n7955__));
  buf1  g7014(.din(new_new_n7954__), .dout(new_new_n7956__));
  buf1  g7015(.din(new_new_n1094__), .dout(new_new_n7957__));
  buf1  g7016(.din(new_new_n7957__), .dout(new_new_n7958__));
  buf1  g7017(.din(new_new_n3175__), .dout(new_new_n7959__));
  buf1  g7018(.din(new_new_n3173__), .dout(new_new_n7960__));
  buf1  g7019(.din(new_new_n3174__), .dout(new_new_n7961__));
  buf1  g7020(.din(new_new_n3172__), .dout(new_new_n7962__));
  buf1  g7021(.din(new_new_n3177__), .dout(new_new_n7963__));
  buf1  g7022(.din(new_new_n7963__), .dout(new_new_n7964__));
  buf1  g7023(.din(new_new_n3176__), .dout(new_new_n7965__));
  buf1  g7024(.din(new_new_n7965__), .dout(new_new_n7966__));
  buf1  g7025(.din(new_new_n3179__), .dout(new_new_n7967__));
  buf1  g7026(.din(new_new_n3165__), .dout(new_new_n7968__));
  buf1  g7027(.din(new_new_n3178__), .dout(new_new_n7969__));
  buf1  g7028(.din(new_new_n3164__), .dout(new_new_n7970__));
  buf1  g7029(.din(new_new_n3181__), .dout(new_new_n7971__));
  buf1  g7030(.din(new_new_n7971__), .dout(new_new_n7972__));
  buf1  g7031(.din(new_new_n3180__), .dout(new_new_n7973__));
  buf1  g7032(.din(new_new_n7973__), .dout(new_new_n7974__));
  buf1  g7033(.din(new_new_n3189__), .dout(new_new_n7975__));
  buf1  g7034(.din(new_new_n3187__), .dout(new_new_n7976__));
  buf1  g7035(.din(new_new_n3188__), .dout(new_new_n7977__));
  buf1  g7036(.din(new_new_n3186__), .dout(new_new_n7978__));
  buf1  g7037(.din(new_new_n3191__), .dout(new_new_n7979__));
  buf1  g7038(.din(new_new_n7979__), .dout(new_new_n7980__));
  buf1  g7039(.din(new_new_n3190__), .dout(new_new_n7981__));
  buf1  g7040(.din(new_new_n7981__), .dout(new_new_n7982__));
  buf1  g7041(.din(new_new_n1101__), .dout(new_new_n7983__));
  buf1  g7042(.din(new_new_n7983__), .dout(new_new_n7984__));
  buf1  g7043(.din(new_new_n7983__), .dout(new_new_n7985__));
  buf1  g7044(.din(new_new_n1102__), .dout(new_new_n7986__));
  buf1  g7045(.din(new_new_n7986__), .dout(new_new_n7987__));
  buf1  g7046(.din(new_new_n7986__), .dout(new_new_n7988__));
  buf1  g7047(.din(new_new_n3207__), .dout(new_new_n7989__));
  buf1  g7048(.din(new_new_n3205__), .dout(new_new_n7990__));
  buf1  g7049(.din(new_new_n3206__), .dout(new_new_n7991__));
  buf1  g7050(.din(new_new_n3204__), .dout(new_new_n7992__));
  buf1  g7051(.din(new_new_n3209__), .dout(new_new_n7993__));
  buf1  g7052(.din(new_new_n7993__), .dout(new_new_n7994__));
  buf1  g7053(.din(new_new_n3208__), .dout(new_new_n7995__));
  buf1  g7054(.din(new_new_n7995__), .dout(new_new_n7996__));
  buf1  g7055(.din(new_new_n3211__), .dout(new_new_n7997__));
  buf1  g7056(.din(new_new_n3203__), .dout(new_new_n7998__));
  buf1  g7057(.din(new_new_n3210__), .dout(new_new_n7999__));
  buf1  g7058(.din(new_new_n3202__), .dout(new_new_n8000__));
  buf1  g7059(.din(new_new_n3213__), .dout(new_new_n8001__));
  buf1  g7060(.din(new_new_n8001__), .dout(new_new_n8002__));
  buf1  g7061(.din(new_new_n3212__), .dout(new_new_n8003__));
  buf1  g7062(.din(new_new_n8003__), .dout(new_new_n8004__));
  buf1  g7063(.din(new_new_n3221__), .dout(new_new_n8005__));
  buf1  g7064(.din(new_new_n3219__), .dout(new_new_n8006__));
  buf1  g7065(.din(new_new_n3220__), .dout(new_new_n8007__));
  buf1  g7066(.din(new_new_n3218__), .dout(new_new_n8008__));
  buf1  g7067(.din(new_new_n3223__), .dout(new_new_n8009__));
  buf1  g7068(.din(new_new_n8009__), .dout(new_new_n8010__));
  buf1  g7069(.din(new_new_n3222__), .dout(new_new_n8011__));
  buf1  g7070(.din(new_new_n8011__), .dout(new_new_n8012__));
  buf1  g7071(.din(new_new_n3225__), .dout(new_new_n8013__));
  buf1  g7072(.din(new_new_n3197__), .dout(new_new_n8014__));
  buf1  g7073(.din(new_new_n3224__), .dout(new_new_n8015__));
  buf1  g7074(.din(new_new_n3196__), .dout(new_new_n8016__));
  buf1  g7075(.din(new_new_n3227__), .dout(new_new_n8017__));
  buf1  g7076(.din(new_new_n8017__), .dout(new_new_n8018__));
  buf1  g7077(.din(new_new_n3226__), .dout(new_new_n8019__));
  buf1  g7078(.din(new_new_n8019__), .dout(new_new_n8020__));
  buf1  g7079(.din(new_new_n3235__), .dout(new_new_n8021__));
  buf1  g7080(.din(new_new_n3233__), .dout(new_new_n8022__));
  buf1  g7081(.din(new_new_n3234__), .dout(new_new_n8023__));
  buf1  g7082(.din(new_new_n3232__), .dout(new_new_n8024__));
  buf1  g7083(.din(new_new_n3237__), .dout(new_new_n8025__));
  buf1  g7084(.din(new_new_n8025__), .dout(new_new_n8026__));
  buf1  g7085(.din(new_new_n3236__), .dout(new_new_n8027__));
  buf1  g7086(.din(new_new_n8027__), .dout(new_new_n8028__));
  buf1  g7087(.din(new_new_n1526__), .dout(new_new_n8029__));
  buf1  g7088(.din(new_new_n8029__), .dout(new_new_n8030__));
  buf1  g7089(.din(new_new_n1525__), .dout(new_new_n8031__));
  buf1  g7090(.din(new_new_n8031__), .dout(new_new_n8032__));
  buf1  g7091(.din(new_new_n3257__), .dout(new_new_n8033__));
  buf1  g7092(.din(new_new_n3255__), .dout(new_new_n8034__));
  buf1  g7093(.din(new_new_n3256__), .dout(new_new_n8035__));
  buf1  g7094(.din(new_new_n3254__), .dout(new_new_n8036__));
  buf1  g7095(.din(new_new_n3259__), .dout(new_new_n8037__));
  buf1  g7096(.din(new_new_n8037__), .dout(new_new_n8038__));
  buf1  g7097(.din(new_new_n3258__), .dout(new_new_n8039__));
  buf1  g7098(.din(new_new_n8039__), .dout(new_new_n8040__));
  buf1  g7099(.din(new_new_n1103__), .dout(new_new_n8041__));
  buf1  g7100(.din(new_new_n8041__), .dout(new_new_n8042__));
  buf1  g7101(.din(new_new_n8041__), .dout(new_new_n8043__));
  buf1  g7102(.din(new_new_n1104__), .dout(new_new_n8044__));
  buf1  g7103(.din(new_new_n8044__), .dout(new_new_n8045__));
  buf1  g7104(.din(new_new_n3267__), .dout(new_new_n8046__));
  buf1  g7105(.din(new_new_n3265__), .dout(new_new_n8047__));
  buf1  g7106(.din(new_new_n3266__), .dout(new_new_n8048__));
  buf1  g7107(.din(new_new_n3264__), .dout(new_new_n8049__));
  buf1  g7108(.din(new_new_n3269__), .dout(new_new_n8050__));
  buf1  g7109(.din(new_new_n8050__), .dout(new_new_n8051__));
  buf1  g7110(.din(new_new_n3268__), .dout(new_new_n8052__));
  buf1  g7111(.din(new_new_n8052__), .dout(new_new_n8053__));
  buf1  g7112(.din(new_new_n3271__), .dout(new_new_n8054__));
  buf1  g7113(.din(new_new_n3249__), .dout(new_new_n8055__));
  buf1  g7114(.din(new_new_n3270__), .dout(new_new_n8056__));
  buf1  g7115(.din(new_new_n3248__), .dout(new_new_n8057__));
  buf1  g7116(.din(new_new_n3273__), .dout(new_new_n8058__));
  buf1  g7117(.din(new_new_n8058__), .dout(new_new_n8059__));
  buf1  g7118(.din(new_new_n3272__), .dout(new_new_n8060__));
  buf1  g7119(.din(new_new_n8060__), .dout(new_new_n8061__));
  buf1  g7120(.din(new_new_n3281__), .dout(new_new_n8062__));
  buf1  g7121(.din(new_new_n3279__), .dout(new_new_n8063__));
  buf1  g7122(.din(new_new_n3280__), .dout(new_new_n8064__));
  buf1  g7123(.din(new_new_n3278__), .dout(new_new_n8065__));
  buf1  g7124(.din(new_new_n3283__), .dout(new_new_n8066__));
  buf1  g7125(.din(new_new_n8066__), .dout(new_new_n8067__));
  buf1  g7126(.din(new_new_n3282__), .dout(new_new_n8068__));
  buf1  g7127(.din(new_new_n8068__), .dout(new_new_n8069__));
  buf1  g7128(.din(new_new_n3285__), .dout(new_new_n8070__));
  buf1  g7129(.din(new_new_n3243__), .dout(new_new_n8071__));
  buf1  g7130(.din(new_new_n3284__), .dout(new_new_n8072__));
  buf1  g7131(.din(new_new_n3242__), .dout(new_new_n8073__));
  buf1  g7132(.din(new_new_n3295__), .dout(new_new_n8074__));
  buf1  g7133(.din(new_new_n3293__), .dout(new_new_n8075__));
  buf1  g7134(.din(new_new_n3294__), .dout(new_new_n8076__));
  buf1  g7135(.din(new_new_n3292__), .dout(new_new_n8077__));
  buf1  g7136(.din(new_new_n3297__), .dout(new_new_n8078__));
  buf1  g7137(.din(new_new_n8078__), .dout(new_new_n8079__));
  buf1  g7138(.din(new_new_n3296__), .dout(new_new_n8080__));
  buf1  g7139(.din(new_new_n8080__), .dout(new_new_n8081__));
  buf1  g7140(.din(new_new_n1107__), .dout(new_new_n8082__));
  buf1  g7141(.din(new_new_n8082__), .dout(new_new_n8083__));
  buf1  g7142(.din(new_new_n8082__), .dout(new_new_n8084__));
  buf1  g7143(.din(new_new_n1108__), .dout(new_new_n8085__));
  buf1  g7144(.din(new_new_n8085__), .dout(new_new_n8086__));
  buf1  g7145(.din(new_new_n3305__), .dout(new_new_n8087__));
  buf1  g7146(.din(new_new_n3303__), .dout(new_new_n8088__));
  buf1  g7147(.din(new_new_n3304__), .dout(new_new_n8089__));
  buf1  g7148(.din(new_new_n3302__), .dout(new_new_n8090__));
  buf1  g7149(.din(new_new_n3307__), .dout(new_new_n8091__));
  buf1  g7150(.din(new_new_n8091__), .dout(new_new_n8092__));
  buf1  g7151(.din(new_new_n3306__), .dout(new_new_n8093__));
  buf1  g7152(.din(new_new_n8093__), .dout(new_new_n8094__));
  buf1  g7153(.din(new_new_n1544__), .dout(new_new_n8095__));
  buf1  g7154(.din(new_new_n1496__), .dout(new_new_n8096__));
  buf1  g7155(.din(new_new_n1543__), .dout(new_new_n8097__));
  buf1  g7156(.din(new_new_n1495__), .dout(new_new_n8098__));
  buf1  g7157(.din(new_new_n3315__), .dout(new_new_n8099__));
  buf1  g7158(.din(new_new_n8099__), .dout(new_new_n8100__));
  buf1  g7159(.din(new_new_n3314__), .dout(new_new_n8101__));
  buf1  g7160(.din(new_new_n8101__), .dout(new_new_n8102__));
  buf1  g7161(.din(new_new_n1109__), .dout(new_new_n8103__));
  buf1  g7162(.din(new_new_n8103__), .dout(new_new_n8104__));
  buf1  g7163(.din(new_new_n8103__), .dout(new_new_n8105__));
  buf1  g7164(.din(new_new_n1110__), .dout(new_new_n8106__));
  buf1  g7165(.din(new_new_n8106__), .dout(new_new_n8107__));
  buf1  g7166(.din(new_new_n3323__), .dout(new_new_n8108__));
  buf1  g7167(.din(new_new_n3321__), .dout(new_new_n8109__));
  buf1  g7168(.din(new_new_n3322__), .dout(new_new_n8110__));
  buf1  g7169(.din(new_new_n3320__), .dout(new_new_n8111__));
  buf1  g7170(.din(new_new_n3325__), .dout(new_new_n8112__));
  buf1  g7171(.din(new_new_n8112__), .dout(new_new_n8113__));
  buf1  g7172(.din(new_new_n3324__), .dout(new_new_n8114__));
  buf1  g7173(.din(new_new_n8114__), .dout(new_new_n8115__));
  buf1  g7174(.din(new_new_n3327__), .dout(new_new_n8116__));
  buf1  g7175(.din(new_new_n3313__), .dout(new_new_n8117__));
  buf1  g7176(.din(new_new_n3326__), .dout(new_new_n8118__));
  buf1  g7177(.din(new_new_n3312__), .dout(new_new_n8119__));
  buf1  g7178(.din(new_new_n3329__), .dout(new_new_n8120__));
  buf1  g7179(.din(new_new_n8120__), .dout(new_new_n8121__));
  buf1  g7180(.din(new_new_n3328__), .dout(new_new_n8122__));
  buf1  g7181(.din(new_new_n8122__), .dout(new_new_n8123__));
  buf1  g7182(.din(new_new_n3337__), .dout(new_new_n8124__));
  buf1  g7183(.din(new_new_n3335__), .dout(new_new_n8125__));
  buf1  g7184(.din(new_new_n3336__), .dout(new_new_n8126__));
  buf1  g7185(.din(new_new_n3334__), .dout(new_new_n8127__));
  buf1  g7186(.din(new_new_n3339__), .dout(new_new_n8128__));
  buf1  g7187(.din(new_new_n8128__), .dout(new_new_n8129__));
  buf1  g7188(.din(new_new_n3338__), .dout(new_new_n8130__));
  buf1  g7189(.din(new_new_n8130__), .dout(new_new_n8131__));
  buf1  g7190(.din(new_new_n1111__), .dout(new_new_n8132__));
  buf1  g7191(.din(new_new_n8132__), .dout(new_new_n8133__));
  buf1  g7192(.din(new_new_n8132__), .dout(new_new_n8134__));
  buf1  g7193(.din(new_new_n1112__), .dout(new_new_n8135__));
  buf1  g7194(.din(new_new_n8135__), .dout(new_new_n8136__));
  buf1  g7195(.din(new_new_n8135__), .dout(new_new_n8137__));
  buf1  g7196(.din(new_new_n3355__), .dout(new_new_n8138__));
  buf1  g7197(.din(new_new_n3353__), .dout(new_new_n8139__));
  buf1  g7198(.din(new_new_n3354__), .dout(new_new_n8140__));
  buf1  g7199(.din(new_new_n3352__), .dout(new_new_n8141__));
  buf1  g7200(.din(new_new_n3357__), .dout(new_new_n8142__));
  buf1  g7201(.din(new_new_n8142__), .dout(new_new_n8143__));
  buf1  g7202(.din(new_new_n3356__), .dout(new_new_n8144__));
  buf1  g7203(.din(new_new_n8144__), .dout(new_new_n8145__));
  buf1  g7204(.din(new_new_n3359__), .dout(new_new_n8146__));
  buf1  g7205(.din(new_new_n3351__), .dout(new_new_n8147__));
  buf1  g7206(.din(new_new_n3358__), .dout(new_new_n8148__));
  buf1  g7207(.din(new_new_n3350__), .dout(new_new_n8149__));
  buf1  g7208(.din(new_new_n3361__), .dout(new_new_n8150__));
  buf1  g7209(.din(new_new_n8150__), .dout(new_new_n8151__));
  buf1  g7210(.din(new_new_n3360__), .dout(new_new_n8152__));
  buf1  g7211(.din(new_new_n8152__), .dout(new_new_n8153__));
  buf1  g7212(.din(new_new_n3369__), .dout(new_new_n8154__));
  buf1  g7213(.din(new_new_n3367__), .dout(new_new_n8155__));
  buf1  g7214(.din(new_new_n3368__), .dout(new_new_n8156__));
  buf1  g7215(.din(new_new_n3366__), .dout(new_new_n8157__));
  buf1  g7216(.din(new_new_n3371__), .dout(new_new_n8158__));
  buf1  g7217(.din(new_new_n8158__), .dout(new_new_n8159__));
  buf1  g7218(.din(new_new_n3370__), .dout(new_new_n8160__));
  buf1  g7219(.din(new_new_n8160__), .dout(new_new_n8161__));
  buf1  g7220(.din(new_new_n3373__), .dout(new_new_n8162__));
  buf1  g7221(.din(new_new_n3345__), .dout(new_new_n8163__));
  buf1  g7222(.din(new_new_n3372__), .dout(new_new_n8164__));
  buf1  g7223(.din(new_new_n3344__), .dout(new_new_n8165__));
  buf1  g7224(.din(new_new_n3375__), .dout(new_new_n8166__));
  buf1  g7225(.din(new_new_n8166__), .dout(new_new_n8167__));
  buf1  g7226(.din(new_new_n3374__), .dout(new_new_n8168__));
  buf1  g7227(.din(new_new_n8168__), .dout(new_new_n8169__));
  buf1  g7228(.din(new_new_n3383__), .dout(new_new_n8170__));
  buf1  g7229(.din(new_new_n3381__), .dout(new_new_n8171__));
  buf1  g7230(.din(new_new_n3382__), .dout(new_new_n8172__));
  buf1  g7231(.din(new_new_n3380__), .dout(new_new_n8173__));
  buf1  g7232(.din(new_new_n3385__), .dout(new_new_n8174__));
  buf1  g7233(.din(new_new_n8174__), .dout(new_new_n8175__));
  buf1  g7234(.din(new_new_n3384__), .dout(new_new_n8176__));
  buf1  g7235(.din(new_new_n8176__), .dout(new_new_n8177__));
  buf1  g7236(.din(new_new_n1528__), .dout(new_new_n8178__));
  buf1  g7237(.din(new_new_n8178__), .dout(new_new_n8179__));
  buf1  g7238(.din(new_new_n1527__), .dout(new_new_n8180__));
  buf1  g7239(.din(new_new_n8180__), .dout(new_new_n8181__));
  buf1  g7240(.din(new_new_n3405__), .dout(new_new_n8182__));
  buf1  g7241(.din(new_new_n3403__), .dout(new_new_n8183__));
  buf1  g7242(.din(new_new_n3404__), .dout(new_new_n8184__));
  buf1  g7243(.din(new_new_n3402__), .dout(new_new_n8185__));
  buf1  g7244(.din(new_new_n3407__), .dout(new_new_n8186__));
  buf1  g7245(.din(new_new_n8186__), .dout(new_new_n8187__));
  buf1  g7246(.din(new_new_n3406__), .dout(new_new_n8188__));
  buf1  g7247(.din(new_new_n8188__), .dout(new_new_n8189__));
  buf1  g7248(.din(new_new_n1113__), .dout(new_new_n8190__));
  buf1  g7249(.din(new_new_n8190__), .dout(new_new_n8191__));
  buf1  g7250(.din(new_new_n8190__), .dout(new_new_n8192__));
  buf1  g7251(.din(new_new_n1114__), .dout(new_new_n8193__));
  buf1  g7252(.din(new_new_n8193__), .dout(new_new_n8194__));
  buf1  g7253(.din(new_new_n3415__), .dout(new_new_n8195__));
  buf1  g7254(.din(new_new_n3413__), .dout(new_new_n8196__));
  buf1  g7255(.din(new_new_n3414__), .dout(new_new_n8197__));
  buf1  g7256(.din(new_new_n3412__), .dout(new_new_n8198__));
  buf1  g7257(.din(new_new_n3417__), .dout(new_new_n8199__));
  buf1  g7258(.din(new_new_n8199__), .dout(new_new_n8200__));
  buf1  g7259(.din(new_new_n3416__), .dout(new_new_n8201__));
  buf1  g7260(.din(new_new_n8201__), .dout(new_new_n8202__));
  buf1  g7261(.din(new_new_n3419__), .dout(new_new_n8203__));
  buf1  g7262(.din(new_new_n3397__), .dout(new_new_n8204__));
  buf1  g7263(.din(new_new_n3418__), .dout(new_new_n8205__));
  buf1  g7264(.din(new_new_n3396__), .dout(new_new_n8206__));
  buf1  g7265(.din(new_new_n3421__), .dout(new_new_n8207__));
  buf1  g7266(.din(new_new_n8207__), .dout(new_new_n8208__));
  buf1  g7267(.din(new_new_n3420__), .dout(new_new_n8209__));
  buf1  g7268(.din(new_new_n8209__), .dout(new_new_n8210__));
  buf1  g7269(.din(new_new_n3429__), .dout(new_new_n8211__));
  buf1  g7270(.din(new_new_n3427__), .dout(new_new_n8212__));
  buf1  g7271(.din(new_new_n3428__), .dout(new_new_n8213__));
  buf1  g7272(.din(new_new_n3426__), .dout(new_new_n8214__));
  buf1  g7273(.din(new_new_n3431__), .dout(new_new_n8215__));
  buf1  g7274(.din(new_new_n8215__), .dout(new_new_n8216__));
  buf1  g7275(.din(new_new_n3430__), .dout(new_new_n8217__));
  buf1  g7276(.din(new_new_n8217__), .dout(new_new_n8218__));
  buf1  g7277(.din(new_new_n3433__), .dout(new_new_n8219__));
  buf1  g7278(.din(new_new_n3391__), .dout(new_new_n8220__));
  buf1  g7279(.din(new_new_n3432__), .dout(new_new_n8221__));
  buf1  g7280(.din(new_new_n3390__), .dout(new_new_n8222__));
  buf1  g7281(.din(new_new_n1549__), .dout(new_new_n8223__));
  buf1  g7282(.din(new_new_n1486__), .dout(new_new_n8224__));
  buf1  g7283(.din(new_new_n1550__), .dout(new_new_n8225__));
  buf1  g7284(.din(new_new_n1485__), .dout(new_new_n8226__));
  buf1  g7285(.din(new_new_n3443__), .dout(new_new_n8227__));
  buf1  g7286(.din(new_new_n8227__), .dout(new_new_n8228__));
  buf1  g7287(.din(new_new_n3442__), .dout(new_new_n8229__));
  buf1  g7288(.din(new_new_n8229__), .dout(new_new_n8230__));
  buf1  g7289(.din(new_new_n3445__), .dout(new_new_n8231__));
  buf1  g7290(.din(new_new_n3441__), .dout(new_new_n8232__));
  buf1  g7291(.din(new_new_n3444__), .dout(new_new_n8233__));
  buf1  g7292(.din(new_new_n3440__), .dout(new_new_n8234__));
  buf1  g7293(.din(new_new_n3447__), .dout(new_new_n8235__));
  buf1  g7294(.din(new_new_n8235__), .dout(new_new_n8236__));
  buf1  g7295(.din(new_new_n3446__), .dout(new_new_n8237__));
  buf1  g7296(.din(new_new_n8237__), .dout(new_new_n8238__));
  buf1  g7297(.din(new_new_n1115__), .dout(new_new_n8239__));
  buf1  g7298(.din(new_new_n8239__), .dout(new_new_n8240__));
  buf1  g7299(.din(new_new_n8239__), .dout(new_new_n8241__));
  buf1  g7300(.din(new_new_n1116__), .dout(new_new_n8242__));
  buf1  g7301(.din(new_new_n8242__), .dout(new_new_n8243__));
  buf1  g7302(.din(new_new_n3455__), .dout(new_new_n8244__));
  buf1  g7303(.din(new_new_n3453__), .dout(new_new_n8245__));
  buf1  g7304(.din(new_new_n3454__), .dout(new_new_n8246__));
  buf1  g7305(.din(new_new_n3452__), .dout(new_new_n8247__));
  buf1  g7306(.din(new_new_n3457__), .dout(new_new_n8248__));
  buf1  g7307(.din(new_new_n8248__), .dout(new_new_n8249__));
  buf1  g7308(.din(new_new_n3456__), .dout(new_new_n8250__));
  buf1  g7309(.din(new_new_n8250__), .dout(new_new_n8251__));
  buf1  g7310(.din(new_new_n1119__), .dout(new_new_n8252__));
  buf1  g7311(.din(new_new_n8252__), .dout(new_new_n8253__));
  buf1  g7312(.din(new_new_n8253__), .dout(new_new_n8254__));
  buf1  g7313(.din(new_new_n8252__), .dout(new_new_n8255__));
  buf1  g7314(.din(new_new_n1120__), .dout(new_new_n8256__));
  buf1  g7315(.din(new_new_n8256__), .dout(new_new_n8257__));
  buf1  g7316(.din(new_new_n8256__), .dout(new_new_n8258__));
  buf1  g7317(.din(new_new_n3473__), .dout(new_new_n8259__));
  buf1  g7318(.din(new_new_n3471__), .dout(new_new_n8260__));
  buf1  g7319(.din(new_new_n3472__), .dout(new_new_n8261__));
  buf1  g7320(.din(new_new_n3470__), .dout(new_new_n8262__));
  buf1  g7321(.din(new_new_n3475__), .dout(new_new_n8263__));
  buf1  g7322(.din(new_new_n8263__), .dout(new_new_n8264__));
  buf1  g7323(.din(new_new_n3474__), .dout(new_new_n8265__));
  buf1  g7324(.din(new_new_n8265__), .dout(new_new_n8266__));
  buf1  g7325(.din(new_new_n3477__), .dout(new_new_n8267__));
  buf1  g7326(.din(new_new_n3469__), .dout(new_new_n8268__));
  buf1  g7327(.din(new_new_n3476__), .dout(new_new_n8269__));
  buf1  g7328(.din(new_new_n3468__), .dout(new_new_n8270__));
  buf1  g7329(.din(new_new_n3479__), .dout(new_new_n8271__));
  buf1  g7330(.din(new_new_n8271__), .dout(new_new_n8272__));
  buf1  g7331(.din(new_new_n3478__), .dout(new_new_n8273__));
  buf1  g7332(.din(new_new_n8273__), .dout(new_new_n8274__));
  buf1  g7333(.din(new_new_n3487__), .dout(new_new_n8275__));
  buf1  g7334(.din(new_new_n3485__), .dout(new_new_n8276__));
  buf1  g7335(.din(new_new_n3486__), .dout(new_new_n8277__));
  buf1  g7336(.din(new_new_n3484__), .dout(new_new_n8278__));
  buf1  g7337(.din(new_new_n3489__), .dout(new_new_n8279__));
  buf1  g7338(.din(new_new_n8279__), .dout(new_new_n8280__));
  buf1  g7339(.din(new_new_n3488__), .dout(new_new_n8281__));
  buf1  g7340(.din(new_new_n8281__), .dout(new_new_n8282__));
  buf1  g7341(.din(new_new_n3491__), .dout(new_new_n8283__));
  buf1  g7342(.din(new_new_n3463__), .dout(new_new_n8284__));
  buf1  g7343(.din(new_new_n3490__), .dout(new_new_n8285__));
  buf1  g7344(.din(new_new_n3462__), .dout(new_new_n8286__));
  buf1  g7345(.din(new_new_n3493__), .dout(new_new_n8287__));
  buf1  g7346(.din(new_new_n8287__), .dout(new_new_n8288__));
  buf1  g7347(.din(new_new_n3492__), .dout(new_new_n8289__));
  buf1  g7348(.din(new_new_n8289__), .dout(new_new_n8290__));
  buf1  g7349(.din(new_new_n3501__), .dout(new_new_n8291__));
  buf1  g7350(.din(new_new_n3499__), .dout(new_new_n8292__));
  buf1  g7351(.din(new_new_n3500__), .dout(new_new_n8293__));
  buf1  g7352(.din(new_new_n3498__), .dout(new_new_n8294__));
  buf1  g7353(.din(new_new_n3503__), .dout(new_new_n8295__));
  buf1  g7354(.din(new_new_n8295__), .dout(new_new_n8296__));
  buf1  g7355(.din(new_new_n3502__), .dout(new_new_n8297__));
  buf1  g7356(.din(new_new_n8297__), .dout(new_new_n8298__));
  buf1  g7357(.din(new_new_n1535__), .dout(new_new_n8299__));
  buf1  g7358(.din(new_new_n8299__), .dout(new_new_n8300__));
  buf1  g7359(.din(new_new_n1536__), .dout(new_new_n8301__));
  buf1  g7360(.din(new_new_n8301__), .dout(new_new_n8302__));
  buf1  g7361(.din(new_new_n1123__), .dout(new_new_n8303__));
  buf1  g7362(.din(new_new_n8303__), .dout(new_new_n8304__));
  buf1  g7363(.din(new_new_n8304__), .dout(new_new_n8305__));
  buf1  g7364(.din(new_new_n8303__), .dout(new_new_n8306__));
  buf1  g7365(.din(new_new_n1124__), .dout(new_new_n8307__));
  buf1  g7366(.din(new_new_n8307__), .dout(new_new_n8308__));
  buf1  g7367(.din(new_new_n8308__), .dout(new_new_n8309__));
  buf1  g7368(.din(new_new_n8307__), .dout(new_new_n8310__));
  buf1  g7369(.din(new_new_n3529__), .dout(new_new_n8311__));
  buf1  g7370(.din(new_new_n3527__), .dout(new_new_n8312__));
  buf1  g7371(.din(new_new_n3528__), .dout(new_new_n8313__));
  buf1  g7372(.din(new_new_n3526__), .dout(new_new_n8314__));
  buf1  g7373(.din(new_new_n3531__), .dout(new_new_n8315__));
  buf1  g7374(.din(new_new_n8315__), .dout(new_new_n8316__));
  buf1  g7375(.din(new_new_n3530__), .dout(new_new_n8317__));
  buf1  g7376(.din(new_new_n8317__), .dout(new_new_n8318__));
  buf1  g7377(.din(new_new_n3533__), .dout(new_new_n8319__));
  buf1  g7378(.din(new_new_n3521__), .dout(new_new_n8320__));
  buf1  g7379(.din(new_new_n3532__), .dout(new_new_n8321__));
  buf1  g7380(.din(new_new_n3520__), .dout(new_new_n8322__));
  buf1  g7381(.din(new_new_n3535__), .dout(new_new_n8323__));
  buf1  g7382(.din(new_new_n8323__), .dout(new_new_n8324__));
  buf1  g7383(.din(new_new_n3534__), .dout(new_new_n8325__));
  buf1  g7384(.din(new_new_n8325__), .dout(new_new_n8326__));
  buf1  g7385(.din(new_new_n3543__), .dout(new_new_n8327__));
  buf1  g7386(.din(new_new_n3541__), .dout(new_new_n8328__));
  buf1  g7387(.din(new_new_n3542__), .dout(new_new_n8329__));
  buf1  g7388(.din(new_new_n3540__), .dout(new_new_n8330__));
  buf1  g7389(.din(new_new_n3545__), .dout(new_new_n8331__));
  buf1  g7390(.din(new_new_n8331__), .dout(new_new_n8332__));
  buf1  g7391(.din(new_new_n3544__), .dout(new_new_n8333__));
  buf1  g7392(.din(new_new_n8333__), .dout(new_new_n8334__));
  buf1  g7393(.din(new_new_n3547__), .dout(new_new_n8335__));
  buf1  g7394(.din(new_new_n3515__), .dout(new_new_n8336__));
  buf1  g7395(.din(new_new_n3546__), .dout(new_new_n8337__));
  buf1  g7396(.din(new_new_n3514__), .dout(new_new_n8338__));
  buf1  g7397(.din(new_new_n3549__), .dout(new_new_n8339__));
  buf1  g7398(.din(new_new_n8339__), .dout(new_new_n8340__));
  buf1  g7399(.din(new_new_n3548__), .dout(new_new_n8341__));
  buf1  g7400(.din(new_new_n8341__), .dout(new_new_n8342__));
  buf1  g7401(.din(new_new_n3557__), .dout(new_new_n8343__));
  buf1  g7402(.din(new_new_n3555__), .dout(new_new_n8344__));
  buf1  g7403(.din(new_new_n3556__), .dout(new_new_n8345__));
  buf1  g7404(.din(new_new_n3554__), .dout(new_new_n8346__));
  buf1  g7405(.din(new_new_n3559__), .dout(new_new_n8347__));
  buf1  g7406(.din(new_new_n8347__), .dout(new_new_n8348__));
  buf1  g7407(.din(new_new_n3558__), .dout(new_new_n8349__));
  buf1  g7408(.din(new_new_n8349__), .dout(new_new_n8350__));
  buf1  g7409(.din(new_new_n3561__), .dout(new_new_n8351__));
  buf1  g7410(.din(new_new_n3509__), .dout(new_new_n8352__));
  buf1  g7411(.din(new_new_n3560__), .dout(new_new_n8353__));
  buf1  g7412(.din(new_new_n3508__), .dout(new_new_n8354__));
  buf1  g7413(.din(new_new_n3563__), .dout(new_new_n8355__));
  buf1  g7414(.din(new_new_n8355__), .dout(new_new_n8356__));
  buf1  g7415(.din(new_new_n3562__), .dout(new_new_n8357__));
  buf1  g7416(.din(new_new_n8357__), .dout(new_new_n8358__));
  buf1  g7417(.din(new_new_n913__), .dout(new_new_n8359__));
  buf1  g7418(.din(new_new_n8359__), .dout(new_new_n8360__));
  buf1  g7419(.din(new_new_n8360__), .dout(new_new_n8361__));
  buf1  g7420(.din(new_new_n8361__), .dout(new_new_n8362__));
  buf1  g7421(.din(new_new_n8361__), .dout(new_new_n8363__));
  buf1  g7422(.din(new_new_n8360__), .dout(new_new_n8364__));
  buf1  g7423(.din(new_new_n8359__), .dout(new_new_n8365__));
  buf1  g7424(.din(new_new_n8365__), .dout(new_new_n8366__));
  buf1  g7425(.din(new_new_n8365__), .dout(new_new_n8367__));
  buf1  g7426(.din(new_new_n914__), .dout(new_new_n8368__));
  buf1  g7427(.din(new_new_n8368__), .dout(new_new_n8369__));
  buf1  g7428(.din(new_new_n8369__), .dout(new_new_n8370__));
  buf1  g7429(.din(new_new_n8370__), .dout(new_new_n8371__));
  buf1  g7430(.din(new_new_n8370__), .dout(new_new_n8372__));
  buf1  g7431(.din(new_new_n8369__), .dout(new_new_n8373__));
  buf1  g7432(.din(new_new_n8368__), .dout(new_new_n8374__));
  buf1  g7433(.din(new_new_n8374__), .dout(new_new_n8375__));
  buf1  g7434(.din(new_new_n8374__), .dout(new_new_n8376__));
  buf1  g7435(.din(new_new_n3571__), .dout(new_new_n8377__));
  buf1  g7436(.din(new_new_n3569__), .dout(new_new_n8378__));
  buf1  g7437(.din(new_new_n3570__), .dout(new_new_n8379__));
  buf1  g7438(.din(new_new_n3568__), .dout(new_new_n8380__));
  buf1  g7439(.din(new_new_n3573__), .dout(new_new_n8381__));
  buf1  g7440(.din(new_new_n8381__), .dout(new_new_n8382__));
  buf1  g7441(.din(new_new_n3572__), .dout(new_new_n8383__));
  buf1  g7442(.din(new_new_n8383__), .dout(new_new_n8384__));
  buf1  g7443(.din(new_new_n1546__), .dout(new_new_n8385__));
  buf1  g7444(.din(new_new_n1498__), .dout(new_new_n8386__));
  buf1  g7445(.din(new_new_n1545__), .dout(new_new_n8387__));
  buf1  g7446(.din(new_new_n1497__), .dout(new_new_n8388__));
  buf1  g7447(.din(new_new_n3599__), .dout(new_new_n8389__));
  buf1  g7448(.din(new_new_n8389__), .dout(new_new_n8390__));
  buf1  g7449(.din(new_new_n3598__), .dout(new_new_n8391__));
  buf1  g7450(.din(new_new_n8391__), .dout(new_new_n8392__));
  buf1  g7451(.din(new_new_n1127__), .dout(new_new_n8393__));
  buf1  g7452(.din(new_new_n8393__), .dout(new_new_n8394__));
  buf1  g7453(.din(new_new_n8394__), .dout(new_new_n8395__));
  buf1  g7454(.din(new_new_n8394__), .dout(new_new_n8396__));
  buf1  g7455(.din(new_new_n8393__), .dout(new_new_n8397__));
  buf1  g7456(.din(new_new_n1128__), .dout(new_new_n8398__));
  buf1  g7457(.din(new_new_n8398__), .dout(new_new_n8399__));
  buf1  g7458(.din(new_new_n8399__), .dout(new_new_n8400__));
  buf1  g7459(.din(new_new_n8398__), .dout(new_new_n8401__));
  buf1  g7460(.din(new_new_n3607__), .dout(new_new_n8402__));
  buf1  g7461(.din(new_new_n3605__), .dout(new_new_n8403__));
  buf1  g7462(.din(new_new_n3606__), .dout(new_new_n8404__));
  buf1  g7463(.din(new_new_n3604__), .dout(new_new_n8405__));
  buf1  g7464(.din(new_new_n3609__), .dout(new_new_n8406__));
  buf1  g7465(.din(new_new_n8406__), .dout(new_new_n8407__));
  buf1  g7466(.din(new_new_n3608__), .dout(new_new_n8408__));
  buf1  g7467(.din(new_new_n8408__), .dout(new_new_n8409__));
  buf1  g7468(.din(new_new_n3611__), .dout(new_new_n8410__));
  buf1  g7469(.din(new_new_n3597__), .dout(new_new_n8411__));
  buf1  g7470(.din(new_new_n3610__), .dout(new_new_n8412__));
  buf1  g7471(.din(new_new_n3596__), .dout(new_new_n8413__));
  buf1  g7472(.din(new_new_n3613__), .dout(new_new_n8414__));
  buf1  g7473(.din(new_new_n8414__), .dout(new_new_n8415__));
  buf1  g7474(.din(new_new_n3612__), .dout(new_new_n8416__));
  buf1  g7475(.din(new_new_n8416__), .dout(new_new_n8417__));
  buf1  g7476(.din(new_new_n3621__), .dout(new_new_n8418__));
  buf1  g7477(.din(new_new_n3619__), .dout(new_new_n8419__));
  buf1  g7478(.din(new_new_n3620__), .dout(new_new_n8420__));
  buf1  g7479(.din(new_new_n3618__), .dout(new_new_n8421__));
  buf1  g7480(.din(new_new_n3623__), .dout(new_new_n8422__));
  buf1  g7481(.din(new_new_n8422__), .dout(new_new_n8423__));
  buf1  g7482(.din(new_new_n3622__), .dout(new_new_n8424__));
  buf1  g7483(.din(new_new_n8424__), .dout(new_new_n8425__));
  buf1  g7484(.din(new_new_n3625__), .dout(new_new_n8426__));
  buf1  g7485(.din(new_new_n3591__), .dout(new_new_n8427__));
  buf1  g7486(.din(new_new_n3624__), .dout(new_new_n8428__));
  buf1  g7487(.din(new_new_n3590__), .dout(new_new_n8429__));
  buf1  g7488(.din(new_new_n3627__), .dout(new_new_n8430__));
  buf1  g7489(.din(new_new_n8430__), .dout(new_new_n8431__));
  buf1  g7490(.din(new_new_n3626__), .dout(new_new_n8432__));
  buf1  g7491(.din(new_new_n8432__), .dout(new_new_n8433__));
  buf1  g7492(.din(new_new_n3635__), .dout(new_new_n8434__));
  buf1  g7493(.din(new_new_n3633__), .dout(new_new_n8435__));
  buf1  g7494(.din(new_new_n3634__), .dout(new_new_n8436__));
  buf1  g7495(.din(new_new_n3632__), .dout(new_new_n8437__));
  buf1  g7496(.din(new_new_n3637__), .dout(new_new_n8438__));
  buf1  g7497(.din(new_new_n8438__), .dout(new_new_n8439__));
  buf1  g7498(.din(new_new_n3636__), .dout(new_new_n8440__));
  buf1  g7499(.din(new_new_n8440__), .dout(new_new_n8441__));
  buf1  g7500(.din(new_new_n3639__), .dout(new_new_n8442__));
  buf1  g7501(.din(new_new_n3585__), .dout(new_new_n8443__));
  buf1  g7502(.din(new_new_n3638__), .dout(new_new_n8444__));
  buf1  g7503(.din(new_new_n3584__), .dout(new_new_n8445__));
  buf1  g7504(.din(new_new_n3641__), .dout(new_new_n8446__));
  buf1  g7505(.din(new_new_n8446__), .dout(new_new_n8447__));
  buf1  g7506(.din(new_new_n3640__), .dout(new_new_n8448__));
  buf1  g7507(.din(new_new_n8448__), .dout(new_new_n8449__));
  buf1  g7508(.din(new_new_n3649__), .dout(new_new_n8450__));
  buf1  g7509(.din(new_new_n3647__), .dout(new_new_n8451__));
  buf1  g7510(.din(new_new_n3648__), .dout(new_new_n8452__));
  buf1  g7511(.din(new_new_n3646__), .dout(new_new_n8453__));
  buf1  g7512(.din(new_new_n3651__), .dout(new_new_n8454__));
  buf1  g7513(.din(new_new_n8454__), .dout(new_new_n8455__));
  buf1  g7514(.din(new_new_n3650__), .dout(new_new_n8456__));
  buf1  g7515(.din(new_new_n8456__), .dout(new_new_n8457__));
  buf1  g7516(.din(new_new_n3653__), .dout(new_new_n8458__));
  buf1  g7517(.din(new_new_n3579__), .dout(new_new_n8459__));
  buf1  g7518(.din(new_new_n3652__), .dout(new_new_n8460__));
  buf1  g7519(.din(new_new_n3578__), .dout(new_new_n8461__));
  buf1  g7520(.din(new_new_n1611__), .dout(new_new_n8462__));
  buf1  g7521(.din(new_new_n1564__), .dout(new_new_n8463__));
  buf1  g7522(.din(new_new_n1612__), .dout(new_new_n8464__));
  buf1  g7523(.din(new_new_n1563__), .dout(new_new_n8465__));
  buf1  g7524(.din(new_new_n3657__), .dout(new_new_n8466__));
  buf1  g7525(.din(new_new_n8466__), .dout(new_new_n8467__));
  buf1  g7526(.din(new_new_n3656__), .dout(new_new_n8468__));
  buf1  g7527(.din(new_new_n8468__), .dout(new_new_n8469__));
  buf1  g7528(.din(new_new_n3665__), .dout(new_new_n8470__));
  buf1  g7529(.din(new_new_n3663__), .dout(new_new_n8471__));
  buf1  g7530(.din(new_new_n3664__), .dout(new_new_n8472__));
  buf1  g7531(.din(new_new_n3662__), .dout(new_new_n8473__));
  buf1  g7532(.din(new_new_n3667__), .dout(new_new_n8474__));
  buf1  g7533(.din(new_new_n8474__), .dout(new_new_n8475__));
  buf1  g7534(.din(new_new_n3666__), .dout(new_new_n8476__));
  buf1  g7535(.din(new_new_n8476__), .dout(new_new_n8477__));
  buf1  g7536(.din(new_new_n3675__), .dout(new_new_n8478__));
  buf1  g7537(.din(new_new_n3673__), .dout(new_new_n8479__));
  buf1  g7538(.din(new_new_n3674__), .dout(new_new_n8480__));
  buf1  g7539(.din(new_new_n3672__), .dout(new_new_n8481__));
  buf1  g7540(.din(new_new_n3677__), .dout(new_new_n8482__));
  buf1  g7541(.din(new_new_n8482__), .dout(new_new_n8483__));
  buf1  g7542(.din(new_new_n3676__), .dout(new_new_n8484__));
  buf1  g7543(.din(new_new_n8484__), .dout(new_new_n8485__));
  buf1  g7544(.din(new_new_n3685__), .dout(new_new_n8486__));
  buf1  g7545(.din(new_new_n3683__), .dout(new_new_n8487__));
  buf1  g7546(.din(new_new_n3684__), .dout(new_new_n8488__));
  buf1  g7547(.din(new_new_n3682__), .dout(new_new_n8489__));
  buf1  g7548(.din(new_new_n3687__), .dout(new_new_n8490__));
  buf1  g7549(.din(new_new_n8490__), .dout(new_new_n8491__));
  buf1  g7550(.din(new_new_n3686__), .dout(new_new_n8492__));
  buf1  g7551(.din(new_new_n8492__), .dout(new_new_n8493__));
  buf1  g7552(.din(new_new_n3695__), .dout(new_new_n8494__));
  buf1  g7553(.din(new_new_n3693__), .dout(new_new_n8495__));
  buf1  g7554(.din(new_new_n3694__), .dout(new_new_n8496__));
  buf1  g7555(.din(new_new_n3692__), .dout(new_new_n8497__));
  buf1  g7556(.din(new_new_n3697__), .dout(new_new_n8498__));
  buf1  g7557(.din(new_new_n8498__), .dout(new_new_n8499__));
  buf1  g7558(.din(new_new_n3696__), .dout(new_new_n8500__));
  buf1  g7559(.din(new_new_n8500__), .dout(new_new_n8501__));
  buf1  g7560(.din(new_new_n2906__), .dout(new_new_n8502__));
  buf1  g7561(.din(new_new_n3705__), .dout(new_new_n8503__));
  buf1  g7562(.din(new_new_n3703__), .dout(new_new_n8504__));
  buf1  g7563(.din(new_new_n3704__), .dout(new_new_n8505__));
  buf1  g7564(.din(new_new_n3702__), .dout(new_new_n8506__));
  buf1  g7565(.din(new_new_n3707__), .dout(new_new_n8507__));
  buf1  g7566(.din(new_new_n8507__), .dout(new_new_n8508__));
  buf1  g7567(.din(new_new_n3706__), .dout(new_new_n8509__));
  buf1  g7568(.din(new_new_n8509__), .dout(new_new_n8510__));
  buf1  g7569(.din(new_new_n3713__), .dout(new_new_n8511__));
  buf1  g7570(.din(new_new_n3134__), .dout(new_new_n8512__));
  buf1  g7571(.din(new_new_n3721__), .dout(new_new_n8513__));
  buf1  g7572(.din(new_new_n3719__), .dout(new_new_n8514__));
  buf1  g7573(.din(new_new_n3720__), .dout(new_new_n8515__));
  buf1  g7574(.din(new_new_n3718__), .dout(new_new_n8516__));
  buf1  g7575(.din(new_new_n3723__), .dout(new_new_n8517__));
  buf1  g7576(.din(new_new_n8517__), .dout(new_new_n8518__));
  buf1  g7577(.din(new_new_n3722__), .dout(new_new_n8519__));
  buf1  g7578(.din(new_new_n8519__), .dout(new_new_n8520__));
  buf1  g7579(.din(new_new_n1129__), .dout(new_new_n8521__));
  buf1  g7580(.din(new_new_n8521__), .dout(new_new_n8522__));
  buf1  g7581(.din(new_new_n8522__), .dout(new_new_n8523__));
  buf1  g7582(.din(new_new_n8522__), .dout(new_new_n8524__));
  buf1  g7583(.din(new_new_n8521__), .dout(new_new_n8525__));
  buf1  g7584(.din(new_new_n1130__), .dout(new_new_n8526__));
  buf1  g7585(.din(new_new_n8526__), .dout(new_new_n8527__));
  buf1  g7586(.din(new_new_n8527__), .dout(new_new_n8528__));
  buf1  g7587(.din(new_new_n8526__), .dout(new_new_n8529__));
  buf1  g7588(.din(new_new_n3731__), .dout(new_new_n8530__));
  buf1  g7589(.din(new_new_n3729__), .dout(new_new_n8531__));
  buf1  g7590(.din(new_new_n3730__), .dout(new_new_n8532__));
  buf1  g7591(.din(new_new_n3728__), .dout(new_new_n8533__));
  buf1  g7592(.din(new_new_n3733__), .dout(new_new_n8534__));
  buf1  g7593(.din(new_new_n8534__), .dout(new_new_n8535__));
  buf1  g7594(.din(new_new_n3732__), .dout(new_new_n8536__));
  buf1  g7595(.din(new_new_n8536__), .dout(new_new_n8537__));
  buf1  g7596(.din(new_new_n3741__), .dout(new_new_n8538__));
  buf1  g7597(.din(new_new_n3739__), .dout(new_new_n8539__));
  buf1  g7598(.din(new_new_n3740__), .dout(new_new_n8540__));
  buf1  g7599(.din(new_new_n3738__), .dout(new_new_n8541__));
  buf1  g7600(.din(new_new_n3743__), .dout(new_new_n8542__));
  buf1  g7601(.din(new_new_n8542__), .dout(new_new_n8543__));
  buf1  g7602(.din(new_new_n3742__), .dout(new_new_n8544__));
  buf1  g7603(.din(new_new_n8544__), .dout(new_new_n8545__));
  buf1  g7604(.din(new_new_n3751__), .dout(new_new_n8546__));
  buf1  g7605(.din(new_new_n3749__), .dout(new_new_n8547__));
  buf1  g7606(.din(new_new_n3750__), .dout(new_new_n8548__));
  buf1  g7607(.din(new_new_n3748__), .dout(new_new_n8549__));
  buf1  g7608(.din(new_new_n3753__), .dout(new_new_n8550__));
  buf1  g7609(.din(new_new_n8550__), .dout(new_new_n8551__));
  buf1  g7610(.din(new_new_n3752__), .dout(new_new_n8552__));
  buf1  g7611(.din(new_new_n8552__), .dout(new_new_n8553__));
  buf1  g7612(.din(new_new_n3761__), .dout(new_new_n8554__));
  buf1  g7613(.din(new_new_n3759__), .dout(new_new_n8555__));
  buf1  g7614(.din(new_new_n3760__), .dout(new_new_n8556__));
  buf1  g7615(.din(new_new_n3758__), .dout(new_new_n8557__));
  buf1  g7616(.din(new_new_n3763__), .dout(new_new_n8558__));
  buf1  g7617(.din(new_new_n8558__), .dout(new_new_n8559__));
  buf1  g7618(.din(new_new_n3762__), .dout(new_new_n8560__));
  buf1  g7619(.din(new_new_n8560__), .dout(new_new_n8561__));
  buf1  g7620(.din(new_new_n3771__), .dout(new_new_n8562__));
  buf1  g7621(.din(new_new_n3769__), .dout(new_new_n8563__));
  buf1  g7622(.din(new_new_n3770__), .dout(new_new_n8564__));
  buf1  g7623(.din(new_new_n3768__), .dout(new_new_n8565__));
  buf1  g7624(.din(new_new_n3773__), .dout(new_new_n8566__));
  buf1  g7625(.din(new_new_n8566__), .dout(new_new_n8567__));
  buf1  g7626(.din(new_new_n3772__), .dout(new_new_n8568__));
  buf1  g7627(.din(new_new_n8568__), .dout(new_new_n8569__));
  buf1  g7628(.din(new_new_n2862__), .dout(new_new_n8570__));
  buf1  g7629(.din(new_new_n3781__), .dout(new_new_n8571__));
  buf1  g7630(.din(new_new_n3779__), .dout(new_new_n8572__));
  buf1  g7631(.din(new_new_n3780__), .dout(new_new_n8573__));
  buf1  g7632(.din(new_new_n3778__), .dout(new_new_n8574__));
  buf1  g7633(.din(new_new_n3783__), .dout(new_new_n8575__));
  buf1  g7634(.din(new_new_n8575__), .dout(new_new_n8576__));
  buf1  g7635(.din(new_new_n3782__), .dout(new_new_n8577__));
  buf1  g7636(.din(new_new_n8577__), .dout(new_new_n8578__));
  buf1  g7637(.din(new_new_n3163__), .dout(new_new_n8579__));
  buf1  g7638(.din(new_new_n3801__), .dout(new_new_n8580__));
  buf1  g7639(.din(new_new_n3799__), .dout(new_new_n8581__));
  buf1  g7640(.din(new_new_n3800__), .dout(new_new_n8582__));
  buf1  g7641(.din(new_new_n3798__), .dout(new_new_n8583__));
  buf1  g7642(.din(new_new_n3803__), .dout(new_new_n8584__));
  buf1  g7643(.din(new_new_n8584__), .dout(new_new_n8585__));
  buf1  g7644(.din(new_new_n3802__), .dout(new_new_n8586__));
  buf1  g7645(.din(new_new_n3811__), .dout(new_new_n8587__));
  buf1  g7646(.din(new_new_n3809__), .dout(new_new_n8588__));
  buf1  g7647(.din(new_new_n3810__), .dout(new_new_n8589__));
  buf1  g7648(.din(new_new_n3808__), .dout(new_new_n8590__));
  buf1  g7649(.din(new_new_n3813__), .dout(new_new_n8591__));
  buf1  g7650(.din(new_new_n8591__), .dout(new_new_n8592__));
  buf1  g7651(.din(new_new_n3812__), .dout(new_new_n8593__));
  buf1  g7652(.din(new_new_n3830__), .dout(new_new_n8594__));
  buf1  g7653(.din(new_new_n3828__), .dout(new_new_n8595__));
  buf1  g7654(.din(new_new_n3829__), .dout(new_new_n8596__));
  buf1  g7655(.din(new_new_n3827__), .dout(new_new_n8597__));
  buf1  g7656(.din(new_new_n3832__), .dout(new_new_n8598__));
  buf1  g7657(.din(new_new_n8598__), .dout(new_new_n8599__));
  buf1  g7658(.din(new_new_n3831__), .dout(new_new_n8600__));
  buf1  g7659(.din(new_new_n3840__), .dout(new_new_n8601__));
  buf1  g7660(.din(new_new_n3838__), .dout(new_new_n8602__));
  buf1  g7661(.din(new_new_n3839__), .dout(new_new_n8603__));
  buf1  g7662(.din(new_new_n3837__), .dout(new_new_n8604__));
  buf1  g7663(.din(new_new_n3842__), .dout(new_new_n8605__));
  buf1  g7664(.din(new_new_n8605__), .dout(new_new_n8606__));
  buf1  g7665(.din(new_new_n3841__), .dout(new_new_n8607__));
  buf1  g7666(.din(new_new_n3859__), .dout(new_new_n8608__));
  buf1  g7667(.din(new_new_n3857__), .dout(new_new_n8609__));
  buf1  g7668(.din(new_new_n3858__), .dout(new_new_n8610__));
  buf1  g7669(.din(new_new_n3856__), .dout(new_new_n8611__));
  buf1  g7670(.din(new_new_n3861__), .dout(new_new_n8612__));
  buf1  g7671(.din(new_new_n8612__), .dout(new_new_n8613__));
  buf1  g7672(.din(new_new_n3860__), .dout(new_new_n8614__));
  buf1  g7673(.din(new_new_n3869__), .dout(new_new_n8615__));
  buf1  g7674(.din(new_new_n3867__), .dout(new_new_n8616__));
  buf1  g7675(.din(new_new_n3868__), .dout(new_new_n8617__));
  buf1  g7676(.din(new_new_n3866__), .dout(new_new_n8618__));
  buf1  g7677(.din(new_new_n3871__), .dout(new_new_n8619__));
  buf1  g7678(.din(new_new_n8619__), .dout(new_new_n8620__));
  buf1  g7679(.din(new_new_n3870__), .dout(new_new_n8621__));
  buf1  g7680(.din(new_new_n2913__), .dout(new_new_n8622__));
  buf1  g7681(.din(new_new_n8622__), .dout(new_new_n8623__));
  buf1  g7682(.din(new_new_n2962__), .dout(new_new_n8624__));
  buf1  g7683(.din(new_new_n8624__), .dout(new_new_n8625__));
  buf1  g7684(.din(new_new_n3011__), .dout(new_new_n8626__));
  buf1  g7685(.din(new_new_n8626__), .dout(new_new_n8627__));
  buf1  g7686(.din(new_new_n3120__), .dout(new_new_n8628__));
  buf1  g7687(.din(new_new_n8628__), .dout(new_new_n8629__));
  buf1  g7688(.din(new_new_n3789__), .dout(new_new_n8630__));
  buf1  g7689(.din(new_new_n3714__), .dout(new_new_n8631__));
  buf1  g7690(.din(new_new_n3898__), .dout(new_new_n8632__));
  buf1  g7691(.din(new_new_n3896__), .dout(new_new_n8633__));
  buf1  g7692(.din(new_new_n3897__), .dout(new_new_n8634__));
  buf1  g7693(.din(new_new_n3895__), .dout(new_new_n8635__));
  buf1  g7694(.din(new_new_n3900__), .dout(new_new_n8636__));
  buf1  g7695(.din(new_new_n8636__), .dout(new_new_n8637__));
  buf1  g7696(.din(new_new_n3899__), .dout(new_new_n8638__));
  buf1  g7697(.din(new_new_n8638__), .dout(new_new_n8639__));
  buf1  g7698(.din(new_new_n3908__), .dout(new_new_n8640__));
  buf1  g7699(.din(new_new_n3906__), .dout(new_new_n8641__));
  buf1  g7700(.din(new_new_n3907__), .dout(new_new_n8642__));
  buf1  g7701(.din(new_new_n3905__), .dout(new_new_n8643__));
  buf1  g7702(.din(new_new_n3910__), .dout(new_new_n8644__));
  buf1  g7703(.din(new_new_n8644__), .dout(new_new_n8645__));
  buf1  g7704(.din(new_new_n3909__), .dout(new_new_n8646__));
  buf1  g7705(.din(new_new_n8646__), .dout(new_new_n8647__));
  buf1  g7706(.din(new_new_n3927__), .dout(new_new_n8648__));
  buf1  g7707(.din(new_new_n3925__), .dout(new_new_n8649__));
  buf1  g7708(.din(new_new_n3926__), .dout(new_new_n8650__));
  buf1  g7709(.din(new_new_n3924__), .dout(new_new_n8651__));
  buf1  g7710(.din(new_new_n3929__), .dout(new_new_n8652__));
  buf1  g7711(.din(new_new_n8652__), .dout(new_new_n8653__));
  buf1  g7712(.din(new_new_n3928__), .dout(new_new_n8654__));
  buf1  g7713(.din(new_new_n8654__), .dout(new_new_n8655__));
  buf1  g7714(.din(new_new_n3937__), .dout(new_new_n8656__));
  buf1  g7715(.din(new_new_n3935__), .dout(new_new_n8657__));
  buf1  g7716(.din(new_new_n3936__), .dout(new_new_n8658__));
  buf1  g7717(.din(new_new_n3934__), .dout(new_new_n8659__));
  buf1  g7718(.din(new_new_n3939__), .dout(new_new_n8660__));
  buf1  g7719(.din(new_new_n8660__), .dout(new_new_n8661__));
  buf1  g7720(.din(new_new_n3938__), .dout(new_new_n8662__));
  buf1  g7721(.din(new_new_n8662__), .dout(new_new_n8663__));
  buf1  g7722(.din(new_new_n3947__), .dout(new_new_n8664__));
  buf1  g7723(.din(new_new_n3945__), .dout(new_new_n8665__));
  buf1  g7724(.din(new_new_n3946__), .dout(new_new_n8666__));
  buf1  g7725(.din(new_new_n3944__), .dout(new_new_n8667__));
  buf1  g7726(.din(new_new_n3949__), .dout(new_new_n8668__));
  buf1  g7727(.din(new_new_n8668__), .dout(new_new_n8669__));
  buf1  g7728(.din(new_new_n3948__), .dout(new_new_n8670__));
  buf1  g7729(.din(new_new_n8670__), .dout(new_new_n8671__));
  buf1  g7730(.din(new_new_n3957__), .dout(new_new_n8672__));
  buf1  g7731(.din(new_new_n3955__), .dout(new_new_n8673__));
  buf1  g7732(.din(new_new_n3956__), .dout(new_new_n8674__));
  buf1  g7733(.din(new_new_n3954__), .dout(new_new_n8675__));
  buf1  g7734(.din(new_new_n3959__), .dout(new_new_n8676__));
  buf1  g7735(.din(new_new_n8676__), .dout(new_new_n8677__));
  buf1  g7736(.din(new_new_n3958__), .dout(new_new_n8678__));
  buf1  g7737(.din(new_new_n8678__), .dout(new_new_n8679__));
  buf1  g7738(.din(new_new_n3976__), .dout(new_new_n8680__));
  buf1  g7739(.din(new_new_n3974__), .dout(new_new_n8681__));
  buf1  g7740(.din(new_new_n3975__), .dout(new_new_n8682__));
  buf1  g7741(.din(new_new_n3973__), .dout(new_new_n8683__));
  buf1  g7742(.din(new_new_n3978__), .dout(new_new_n8684__));
  buf1  g7743(.din(new_new_n8684__), .dout(new_new_n8685__));
  buf1  g7744(.din(new_new_n3977__), .dout(new_new_n8686__));
  buf1  g7745(.din(new_new_n8686__), .dout(new_new_n8687__));
  buf1  g7746(.din(new_new_n3986__), .dout(new_new_n8688__));
  buf1  g7747(.din(new_new_n3984__), .dout(new_new_n8689__));
  buf1  g7748(.din(new_new_n3985__), .dout(new_new_n8690__));
  buf1  g7749(.din(new_new_n3983__), .dout(new_new_n8691__));
  buf1  g7750(.din(new_new_n3988__), .dout(new_new_n8692__));
  buf1  g7751(.din(new_new_n8692__), .dout(new_new_n8693__));
  buf1  g7752(.din(new_new_n3987__), .dout(new_new_n8694__));
  buf1  g7753(.din(new_new_n8694__), .dout(new_new_n8695__));
  buf1  g7754(.din(new_new_n3996__), .dout(new_new_n8696__));
  buf1  g7755(.din(new_new_n3994__), .dout(new_new_n8697__));
  buf1  g7756(.din(new_new_n3995__), .dout(new_new_n8698__));
  buf1  g7757(.din(new_new_n3993__), .dout(new_new_n8699__));
  buf1  g7758(.din(new_new_n3998__), .dout(new_new_n8700__));
  buf1  g7759(.din(new_new_n8700__), .dout(new_new_n8701__));
  buf1  g7760(.din(new_new_n3997__), .dout(new_new_n8702__));
  buf1  g7761(.din(new_new_n8702__), .dout(new_new_n8703__));
  buf1  g7762(.din(new_new_n4006__), .dout(new_new_n8704__));
  buf1  g7763(.din(new_new_n4004__), .dout(new_new_n8705__));
  buf1  g7764(.din(new_new_n4005__), .dout(new_new_n8706__));
  buf1  g7765(.din(new_new_n4003__), .dout(new_new_n8707__));
  buf1  g7766(.din(new_new_n4008__), .dout(new_new_n8708__));
  buf1  g7767(.din(new_new_n8708__), .dout(new_new_n8709__));
  buf1  g7768(.din(new_new_n4007__), .dout(new_new_n8710__));
  buf1  g7769(.din(new_new_n8710__), .dout(new_new_n8711__));
  buf1  g7770(.din(new_new_n4037__), .dout(new_new_n8712__));
  buf1  g7771(.din(new_new_n4035__), .dout(new_new_n8713__));
  buf1  g7772(.din(new_new_n4036__), .dout(new_new_n8714__));
  buf1  g7773(.din(new_new_n4034__), .dout(new_new_n8715__));
  buf1  g7774(.din(new_new_n4039__), .dout(new_new_n8716__));
  buf1  g7775(.din(new_new_n8716__), .dout(new_new_n8717__));
  buf1  g7776(.din(new_new_n4038__), .dout(new_new_n8718__));
  buf1  g7777(.din(new_new_n8718__), .dout(new_new_n8719__));
  buf1  g7778(.din(new_new_n4047__), .dout(new_new_n8720__));
  buf1  g7779(.din(new_new_n4045__), .dout(new_new_n8721__));
  buf1  g7780(.din(new_new_n4046__), .dout(new_new_n8722__));
  buf1  g7781(.din(new_new_n4044__), .dout(new_new_n8723__));
  buf1  g7782(.din(new_new_n4049__), .dout(new_new_n8724__));
  buf1  g7783(.din(new_new_n8724__), .dout(new_new_n8725__));
  buf1  g7784(.din(new_new_n4048__), .dout(new_new_n8726__));
  buf1  g7785(.din(new_new_n8726__), .dout(new_new_n8727__));
  buf1  g7786(.din(new_new_n4051__), .dout(new_new_n8728__));
  buf1  g7787(.din(new_new_n4029__), .dout(new_new_n8729__));
  buf1  g7788(.din(new_new_n4050__), .dout(new_new_n8730__));
  buf1  g7789(.din(new_new_n4028__), .dout(new_new_n8731__));
  buf1  g7790(.din(new_new_n4053__), .dout(new_new_n8732__));
  buf1  g7791(.din(new_new_n8732__), .dout(new_new_n8733__));
  buf1  g7792(.din(new_new_n4052__), .dout(new_new_n8734__));
  buf1  g7793(.din(new_new_n8734__), .dout(new_new_n8735__));
  buf1  g7794(.din(new_new_n4061__), .dout(new_new_n8736__));
  buf1  g7795(.din(new_new_n4059__), .dout(new_new_n8737__));
  buf1  g7796(.din(new_new_n4060__), .dout(new_new_n8738__));
  buf1  g7797(.din(new_new_n4058__), .dout(new_new_n8739__));
  buf1  g7798(.din(new_new_n4063__), .dout(new_new_n8740__));
  buf1  g7799(.din(new_new_n8740__), .dout(new_new_n8741__));
  buf1  g7800(.din(new_new_n4062__), .dout(new_new_n8742__));
  buf1  g7801(.din(new_new_n8742__), .dout(new_new_n8743__));
  buf1  g7802(.din(new_new_n4065__), .dout(new_new_n8744__));
  buf1  g7803(.din(new_new_n4023__), .dout(new_new_n8745__));
  buf1  g7804(.din(new_new_n4064__), .dout(new_new_n8746__));
  buf1  g7805(.din(new_new_n4022__), .dout(new_new_n8747__));
  buf1  g7806(.din(new_new_n4067__), .dout(new_new_n8748__));
  buf1  g7807(.din(new_new_n8748__), .dout(new_new_n8749__));
  buf1  g7808(.din(new_new_n4066__), .dout(new_new_n8750__));
  buf1  g7809(.din(new_new_n8750__), .dout(new_new_n8751__));
  buf1  g7810(.din(new_new_n4075__), .dout(new_new_n8752__));
  buf1  g7811(.din(new_new_n4073__), .dout(new_new_n8753__));
  buf1  g7812(.din(new_new_n4074__), .dout(new_new_n8754__));
  buf1  g7813(.din(new_new_n4072__), .dout(new_new_n8755__));
  buf1  g7814(.din(new_new_n4077__), .dout(new_new_n8756__));
  buf1  g7815(.din(new_new_n8756__), .dout(new_new_n8757__));
  buf1  g7816(.din(new_new_n4076__), .dout(new_new_n8758__));
  buf1  g7817(.din(new_new_n8758__), .dout(new_new_n8759__));
  buf1  g7818(.din(new_new_n4097__), .dout(new_new_n8760__));
  buf1  g7819(.din(new_new_n4095__), .dout(new_new_n8761__));
  buf1  g7820(.din(new_new_n4096__), .dout(new_new_n8762__));
  buf1  g7821(.din(new_new_n4094__), .dout(new_new_n8763__));
  buf1  g7822(.din(new_new_n4099__), .dout(new_new_n8764__));
  buf1  g7823(.din(new_new_n8764__), .dout(new_new_n8765__));
  buf1  g7824(.din(new_new_n4098__), .dout(new_new_n8766__));
  buf1  g7825(.din(new_new_n8766__), .dout(new_new_n8767__));
  buf1  g7826(.din(new_new_n4107__), .dout(new_new_n8768__));
  buf1  g7827(.din(new_new_n4105__), .dout(new_new_n8769__));
  buf1  g7828(.din(new_new_n4106__), .dout(new_new_n8770__));
  buf1  g7829(.din(new_new_n4104__), .dout(new_new_n8771__));
  buf1  g7830(.din(new_new_n4109__), .dout(new_new_n8772__));
  buf1  g7831(.din(new_new_n8772__), .dout(new_new_n8773__));
  buf1  g7832(.din(new_new_n4108__), .dout(new_new_n8774__));
  buf1  g7833(.din(new_new_n8774__), .dout(new_new_n8775__));
  buf1  g7834(.din(new_new_n4111__), .dout(new_new_n8776__));
  buf1  g7835(.din(new_new_n4089__), .dout(new_new_n8777__));
  buf1  g7836(.din(new_new_n4110__), .dout(new_new_n8778__));
  buf1  g7837(.din(new_new_n4088__), .dout(new_new_n8779__));
  buf1  g7838(.din(new_new_n4113__), .dout(new_new_n8780__));
  buf1  g7839(.din(new_new_n8780__), .dout(new_new_n8781__));
  buf1  g7840(.din(new_new_n4112__), .dout(new_new_n8782__));
  buf1  g7841(.din(new_new_n8782__), .dout(new_new_n8783__));
  buf1  g7842(.din(new_new_n4121__), .dout(new_new_n8784__));
  buf1  g7843(.din(new_new_n4119__), .dout(new_new_n8785__));
  buf1  g7844(.din(new_new_n4120__), .dout(new_new_n8786__));
  buf1  g7845(.din(new_new_n4118__), .dout(new_new_n8787__));
  buf1  g7846(.din(new_new_n4123__), .dout(new_new_n8788__));
  buf1  g7847(.din(new_new_n8788__), .dout(new_new_n8789__));
  buf1  g7848(.din(new_new_n4122__), .dout(new_new_n8790__));
  buf1  g7849(.din(new_new_n8790__), .dout(new_new_n8791__));
  buf1  g7850(.din(new_new_n1185__), .dout(new_new_n8792__));
  buf1  g7851(.din(new_new_n8792__), .dout(new_new_n8793__));
  buf1  g7852(.din(new_new_n8793__), .dout(new_new_n8794__));
  buf1  g7853(.din(new_new_n8792__), .dout(new_new_n8795__));
  buf1  g7854(.din(new_new_n1186__), .dout(new_new_n8796__));
  buf1  g7855(.din(new_new_n8796__), .dout(new_new_n8797__));
  buf1  g7856(.din(new_new_n4130__), .dout(new_new_n8798__));
  buf1  g7857(.din(new_new_n4128__), .dout(new_new_n8799__));
  buf1  g7858(.din(new_new_n4129__), .dout(new_new_n8800__));
  buf1  g7859(.din(new_new_n4127__), .dout(new_new_n8801__));
  buf1  g7860(.din(new_new_n4132__), .dout(new_new_n8802__));
  buf1  g7861(.din(new_new_n8802__), .dout(new_new_n8803__));
  buf1  g7862(.din(new_new_n4131__), .dout(new_new_n8804__));
  buf1  g7863(.din(new_new_n8804__), .dout(new_new_n8805__));
  buf1  g7864(.din(new_new_n1195__), .dout(new_new_n8806__));
  buf1  g7865(.din(new_new_n8806__), .dout(new_new_n8807__));
  buf1  g7866(.din(new_new_n8806__), .dout(new_new_n8808__));
  buf1  g7867(.din(new_new_n1196__), .dout(new_new_n8809__));
  buf1  g7868(.din(new_new_n8809__), .dout(new_new_n8810__));
  buf1  g7869(.din(new_new_n4140__), .dout(new_new_n8811__));
  buf1  g7870(.din(new_new_n4138__), .dout(new_new_n8812__));
  buf1  g7871(.din(new_new_n4139__), .dout(new_new_n8813__));
  buf1  g7872(.din(new_new_n4137__), .dout(new_new_n8814__));
  buf1  g7873(.din(new_new_n4142__), .dout(new_new_n8815__));
  buf1  g7874(.din(new_new_n8815__), .dout(new_new_n8816__));
  buf1  g7875(.din(new_new_n4141__), .dout(new_new_n8817__));
  buf1  g7876(.din(new_new_n8817__), .dout(new_new_n8818__));
  buf1  g7877(.din(new_new_n1604__), .dout(new_new_n8819__));
  buf1  g7878(.din(new_new_n1566__), .dout(new_new_n8820__));
  buf1  g7879(.din(new_new_n1603__), .dout(new_new_n8821__));
  buf1  g7880(.din(new_new_n1565__), .dout(new_new_n8822__));
  buf1  g7881(.din(new_new_n4150__), .dout(new_new_n8823__));
  buf1  g7882(.din(new_new_n8823__), .dout(new_new_n8824__));
  buf1  g7883(.din(new_new_n4149__), .dout(new_new_n8825__));
  buf1  g7884(.din(new_new_n8825__), .dout(new_new_n8826__));
  buf1  g7885(.din(new_new_n1203__), .dout(new_new_n8827__));
  buf1  g7886(.din(new_new_n8827__), .dout(new_new_n8828__));
  buf1  g7887(.din(new_new_n8827__), .dout(new_new_n8829__));
  buf1  g7888(.din(new_new_n1204__), .dout(new_new_n8830__));
  buf1  g7889(.din(new_new_n8830__), .dout(new_new_n8831__));
  buf1  g7890(.din(new_new_n4158__), .dout(new_new_n8832__));
  buf1  g7891(.din(new_new_n4156__), .dout(new_new_n8833__));
  buf1  g7892(.din(new_new_n4157__), .dout(new_new_n8834__));
  buf1  g7893(.din(new_new_n4155__), .dout(new_new_n8835__));
  buf1  g7894(.din(new_new_n4160__), .dout(new_new_n8836__));
  buf1  g7895(.din(new_new_n8836__), .dout(new_new_n8837__));
  buf1  g7896(.din(new_new_n4159__), .dout(new_new_n8838__));
  buf1  g7897(.din(new_new_n8838__), .dout(new_new_n8839__));
  buf1  g7898(.din(new_new_n4162__), .dout(new_new_n8840__));
  buf1  g7899(.din(new_new_n4148__), .dout(new_new_n8841__));
  buf1  g7900(.din(new_new_n4161__), .dout(new_new_n8842__));
  buf1  g7901(.din(new_new_n4147__), .dout(new_new_n8843__));
  buf1  g7902(.din(new_new_n4164__), .dout(new_new_n8844__));
  buf1  g7903(.din(new_new_n8844__), .dout(new_new_n8845__));
  buf1  g7904(.din(new_new_n4163__), .dout(new_new_n8846__));
  buf1  g7905(.din(new_new_n8846__), .dout(new_new_n8847__));
  buf1  g7906(.din(new_new_n4172__), .dout(new_new_n8848__));
  buf1  g7907(.din(new_new_n4170__), .dout(new_new_n8849__));
  buf1  g7908(.din(new_new_n4171__), .dout(new_new_n8850__));
  buf1  g7909(.din(new_new_n4169__), .dout(new_new_n8851__));
  buf1  g7910(.din(new_new_n4174__), .dout(new_new_n8852__));
  buf1  g7911(.din(new_new_n8852__), .dout(new_new_n8853__));
  buf1  g7912(.din(new_new_n4173__), .dout(new_new_n8854__));
  buf1  g7913(.din(new_new_n8854__), .dout(new_new_n8855__));
  buf1  g7914(.din(new_new_n1207__), .dout(new_new_n8856__));
  buf1  g7915(.din(new_new_n8856__), .dout(new_new_n8857__));
  buf1  g7916(.din(new_new_n8856__), .dout(new_new_n8858__));
  buf1  g7917(.din(new_new_n1208__), .dout(new_new_n8859__));
  buf1  g7918(.din(new_new_n8859__), .dout(new_new_n8860__));
  buf1  g7919(.din(new_new_n8859__), .dout(new_new_n8861__));
  buf1  g7920(.din(new_new_n4190__), .dout(new_new_n8862__));
  buf1  g7921(.din(new_new_n4188__), .dout(new_new_n8863__));
  buf1  g7922(.din(new_new_n4189__), .dout(new_new_n8864__));
  buf1  g7923(.din(new_new_n4187__), .dout(new_new_n8865__));
  buf1  g7924(.din(new_new_n4192__), .dout(new_new_n8866__));
  buf1  g7925(.din(new_new_n8866__), .dout(new_new_n8867__));
  buf1  g7926(.din(new_new_n4191__), .dout(new_new_n8868__));
  buf1  g7927(.din(new_new_n8868__), .dout(new_new_n8869__));
  buf1  g7928(.din(new_new_n4194__), .dout(new_new_n8870__));
  buf1  g7929(.din(new_new_n4186__), .dout(new_new_n8871__));
  buf1  g7930(.din(new_new_n4193__), .dout(new_new_n8872__));
  buf1  g7931(.din(new_new_n4185__), .dout(new_new_n8873__));
  buf1  g7932(.din(new_new_n4196__), .dout(new_new_n8874__));
  buf1  g7933(.din(new_new_n8874__), .dout(new_new_n8875__));
  buf1  g7934(.din(new_new_n4195__), .dout(new_new_n8876__));
  buf1  g7935(.din(new_new_n8876__), .dout(new_new_n8877__));
  buf1  g7936(.din(new_new_n4204__), .dout(new_new_n8878__));
  buf1  g7937(.din(new_new_n4202__), .dout(new_new_n8879__));
  buf1  g7938(.din(new_new_n4203__), .dout(new_new_n8880__));
  buf1  g7939(.din(new_new_n4201__), .dout(new_new_n8881__));
  buf1  g7940(.din(new_new_n4206__), .dout(new_new_n8882__));
  buf1  g7941(.din(new_new_n8882__), .dout(new_new_n8883__));
  buf1  g7942(.din(new_new_n4205__), .dout(new_new_n8884__));
  buf1  g7943(.din(new_new_n8884__), .dout(new_new_n8885__));
  buf1  g7944(.din(new_new_n4208__), .dout(new_new_n8886__));
  buf1  g7945(.din(new_new_n4180__), .dout(new_new_n8887__));
  buf1  g7946(.din(new_new_n4207__), .dout(new_new_n8888__));
  buf1  g7947(.din(new_new_n4179__), .dout(new_new_n8889__));
  buf1  g7948(.din(new_new_n4210__), .dout(new_new_n8890__));
  buf1  g7949(.din(new_new_n8890__), .dout(new_new_n8891__));
  buf1  g7950(.din(new_new_n4209__), .dout(new_new_n8892__));
  buf1  g7951(.din(new_new_n8892__), .dout(new_new_n8893__));
  buf1  g7952(.din(new_new_n897__), .dout(new_new_n8894__));
  buf1  g7953(.din(new_new_n8894__), .dout(new_new_n8895__));
  buf1  g7954(.din(new_new_n8895__), .dout(new_new_n8896__));
  buf1  g7955(.din(new_new_n8896__), .dout(new_new_n8897__));
  buf1  g7956(.din(new_new_n8896__), .dout(new_new_n8898__));
  buf1  g7957(.din(new_new_n8895__), .dout(new_new_n8899__));
  buf1  g7958(.din(new_new_n8899__), .dout(new_new_n8900__));
  buf1  g7959(.din(new_new_n8899__), .dout(new_new_n8901__));
  buf1  g7960(.din(new_new_n8894__), .dout(new_new_n8902__));
  buf1  g7961(.din(new_new_n8902__), .dout(new_new_n8903__));
  buf1  g7962(.din(new_new_n8903__), .dout(new_new_n8904__));
  buf1  g7963(.din(new_new_n8903__), .dout(new_new_n8905__));
  buf1  g7964(.din(new_new_n8902__), .dout(new_new_n8906__));
  buf1  g7965(.din(new_new_n8906__), .dout(new_new_n8907__));
  buf1  g7966(.din(new_new_n898__), .dout(new_new_n8908__));
  buf1  g7967(.din(new_new_n8908__), .dout(new_new_n8909__));
  buf1  g7968(.din(new_new_n8909__), .dout(new_new_n8910__));
  buf1  g7969(.din(new_new_n8910__), .dout(new_new_n8911__));
  buf1  g7970(.din(new_new_n8910__), .dout(new_new_n8912__));
  buf1  g7971(.din(new_new_n8909__), .dout(new_new_n8913__));
  buf1  g7972(.din(new_new_n8913__), .dout(new_new_n8914__));
  buf1  g7973(.din(new_new_n8913__), .dout(new_new_n8915__));
  buf1  g7974(.din(new_new_n8908__), .dout(new_new_n8916__));
  buf1  g7975(.din(new_new_n8916__), .dout(new_new_n8917__));
  buf1  g7976(.din(new_new_n8917__), .dout(new_new_n8918__));
  buf1  g7977(.din(new_new_n8917__), .dout(new_new_n8919__));
  buf1  g7978(.din(new_new_n8916__), .dout(new_new_n8920__));
  buf1  g7979(.din(new_new_n8920__), .dout(new_new_n8921__));
  buf1  g7980(.din(new_new_n4218__), .dout(new_new_n8922__));
  buf1  g7981(.din(new_new_n4216__), .dout(new_new_n8923__));
  buf1  g7982(.din(new_new_n4217__), .dout(new_new_n8924__));
  buf1  g7983(.din(new_new_n4215__), .dout(new_new_n8925__));
  buf1  g7984(.din(new_new_n4220__), .dout(new_new_n8926__));
  buf1  g7985(.din(new_new_n8926__), .dout(new_new_n8927__));
  buf1  g7986(.din(new_new_n4219__), .dout(new_new_n8928__));
  buf1  g7987(.din(new_new_n8928__), .dout(new_new_n8929__));
  buf1  g7988(.din(new_new_n1601__), .dout(new_new_n8930__));
  buf1  g7989(.din(new_new_n8930__), .dout(new_new_n8931__));
  buf1  g7990(.din(new_new_n1602__), .dout(new_new_n8932__));
  buf1  g7991(.din(new_new_n8932__), .dout(new_new_n8933__));
  buf1  g7992(.din(new_new_n1209__), .dout(new_new_n8934__));
  buf1  g7993(.din(new_new_n8934__), .dout(new_new_n8935__));
  buf1  g7994(.din(new_new_n8935__), .dout(new_new_n8936__));
  buf1  g7995(.din(new_new_n8934__), .dout(new_new_n8937__));
  buf1  g7996(.din(new_new_n1210__), .dout(new_new_n8938__));
  buf1  g7997(.din(new_new_n8938__), .dout(new_new_n8939__));
  buf1  g7998(.din(new_new_n8938__), .dout(new_new_n8940__));
  buf1  g7999(.din(new_new_n4246__), .dout(new_new_n8941__));
  buf1  g8000(.din(new_new_n4244__), .dout(new_new_n8942__));
  buf1  g8001(.din(new_new_n4245__), .dout(new_new_n8943__));
  buf1  g8002(.din(new_new_n4243__), .dout(new_new_n8944__));
  buf1  g8003(.din(new_new_n4248__), .dout(new_new_n8945__));
  buf1  g8004(.din(new_new_n8945__), .dout(new_new_n8946__));
  buf1  g8005(.din(new_new_n4247__), .dout(new_new_n8947__));
  buf1  g8006(.din(new_new_n8947__), .dout(new_new_n8948__));
  buf1  g8007(.din(new_new_n4250__), .dout(new_new_n8949__));
  buf1  g8008(.din(new_new_n4238__), .dout(new_new_n8950__));
  buf1  g8009(.din(new_new_n4249__), .dout(new_new_n8951__));
  buf1  g8010(.din(new_new_n4237__), .dout(new_new_n8952__));
  buf1  g8011(.din(new_new_n4252__), .dout(new_new_n8953__));
  buf1  g8012(.din(new_new_n8953__), .dout(new_new_n8954__));
  buf1  g8013(.din(new_new_n4251__), .dout(new_new_n8955__));
  buf1  g8014(.din(new_new_n8955__), .dout(new_new_n8956__));
  buf1  g8015(.din(new_new_n4260__), .dout(new_new_n8957__));
  buf1  g8016(.din(new_new_n4258__), .dout(new_new_n8958__));
  buf1  g8017(.din(new_new_n4259__), .dout(new_new_n8959__));
  buf1  g8018(.din(new_new_n4257__), .dout(new_new_n8960__));
  buf1  g8019(.din(new_new_n4262__), .dout(new_new_n8961__));
  buf1  g8020(.din(new_new_n8961__), .dout(new_new_n8962__));
  buf1  g8021(.din(new_new_n4261__), .dout(new_new_n8963__));
  buf1  g8022(.din(new_new_n8963__), .dout(new_new_n8964__));
  buf1  g8023(.din(new_new_n4264__), .dout(new_new_n8965__));
  buf1  g8024(.din(new_new_n4232__), .dout(new_new_n8966__));
  buf1  g8025(.din(new_new_n4263__), .dout(new_new_n8967__));
  buf1  g8026(.din(new_new_n4231__), .dout(new_new_n8968__));
  buf1  g8027(.din(new_new_n4266__), .dout(new_new_n8969__));
  buf1  g8028(.din(new_new_n8969__), .dout(new_new_n8970__));
  buf1  g8029(.din(new_new_n4265__), .dout(new_new_n8971__));
  buf1  g8030(.din(new_new_n8971__), .dout(new_new_n8972__));
  buf1  g8031(.din(new_new_n4274__), .dout(new_new_n8973__));
  buf1  g8032(.din(new_new_n4272__), .dout(new_new_n8974__));
  buf1  g8033(.din(new_new_n4273__), .dout(new_new_n8975__));
  buf1  g8034(.din(new_new_n4271__), .dout(new_new_n8976__));
  buf1  g8035(.din(new_new_n4276__), .dout(new_new_n8977__));
  buf1  g8036(.din(new_new_n8977__), .dout(new_new_n8978__));
  buf1  g8037(.din(new_new_n4275__), .dout(new_new_n8979__));
  buf1  g8038(.din(new_new_n8979__), .dout(new_new_n8980__));
  buf1  g8039(.din(new_new_n4278__), .dout(new_new_n8981__));
  buf1  g8040(.din(new_new_n4226__), .dout(new_new_n8982__));
  buf1  g8041(.din(new_new_n4277__), .dout(new_new_n8983__));
  buf1  g8042(.din(new_new_n4225__), .dout(new_new_n8984__));
  buf1  g8043(.din(new_new_n3287__), .dout(new_new_n8985__));
  buf1  g8044(.din(new_new_n8985__), .dout(new_new_n8986__));
  buf1  g8045(.din(new_new_n3286__), .dout(new_new_n8987__));
  buf1  g8046(.din(new_new_n3435__), .dout(new_new_n8988__));
  buf1  g8047(.din(new_new_n8988__), .dout(new_new_n8989__));
  buf1  g8048(.din(new_new_n3434__), .dout(new_new_n8990__));
  buf1  g8049(.din(new_new_n3655__), .dout(new_new_n8991__));
  buf1  g8050(.din(new_new_n8991__), .dout(new_new_n8992__));
  buf1  g8051(.din(new_new_n3654__), .dout(new_new_n8993__));
  buf1  g8052(.din(new_new_n917__), .dout(new_new_n8994__));
  buf1  g8053(.din(new_new_n8994__), .dout(new_new_n8995__));
  buf1  g8054(.din(new_new_n8994__), .dout(new_new_n8996__));
  buf1  g8055(.din(new_new_n918__), .dout(new_new_n8997__));
  buf1  g8056(.din(new_new_n8997__), .dout(new_new_n8998__));
  buf1  g8057(.din(new_new_n8997__), .dout(new_new_n8999__));
  buf1  g8058(.din(new_new_n4321__), .dout(new_new_n9000__));
  buf1  g8059(.din(new_new_n4319__), .dout(new_new_n9001__));
  buf1  g8060(.din(new_new_n4320__), .dout(new_new_n9002__));
  buf1  g8061(.din(new_new_n4318__), .dout(new_new_n9003__));
  buf1  g8062(.din(new_new_n4323__), .dout(new_new_n9004__));
  buf1  g8063(.din(new_new_n9004__), .dout(new_new_n9005__));
  buf1  g8064(.din(new_new_n4322__), .dout(new_new_n9006__));
  buf1  g8065(.din(new_new_n9006__), .dout(new_new_n9007__));
  buf1  g8066(.din(new_new_n4331__), .dout(new_new_n9008__));
  buf1  g8067(.din(new_new_n4329__), .dout(new_new_n9009__));
  buf1  g8068(.din(new_new_n4330__), .dout(new_new_n9010__));
  buf1  g8069(.din(new_new_n4328__), .dout(new_new_n9011__));
  buf1  g8070(.din(new_new_n4333__), .dout(new_new_n9012__));
  buf1  g8071(.din(new_new_n9012__), .dout(new_new_n9013__));
  buf1  g8072(.din(new_new_n4332__), .dout(new_new_n9014__));
  buf1  g8073(.din(new_new_n9014__), .dout(new_new_n9015__));
  buf1  g8074(.din(new_new_n845__), .dout(new_new_n9016__));
  buf1  g8075(.din(new_new_n9016__), .dout(new_new_n9017__));
  buf1  g8076(.din(new_new_n9017__), .dout(new_new_n9018__));
  buf1  g8077(.din(new_new_n9018__), .dout(new_new_n9019__));
  buf1  g8078(.din(new_new_n9018__), .dout(new_new_n9020__));
  buf1  g8079(.din(new_new_n9017__), .dout(new_new_n9021__));
  buf1  g8080(.din(new_new_n9021__), .dout(new_new_n9022__));
  buf1  g8081(.din(new_new_n9021__), .dout(new_new_n9023__));
  buf1  g8082(.din(new_new_n9016__), .dout(new_new_n9024__));
  buf1  g8083(.din(new_new_n9024__), .dout(new_new_n9025__));
  buf1  g8084(.din(new_new_n9025__), .dout(new_new_n9026__));
  buf1  g8085(.din(new_new_n9024__), .dout(new_new_n9027__));
  buf1  g8086(.din(new_new_n839__), .dout(new_new_n9028__));
  buf1  g8087(.din(new_new_n9028__), .dout(new_new_n9029__));
  buf1  g8088(.din(new_new_n9028__), .dout(new_new_n9030__));
  buf1  g8089(.din(new_new_n846__), .dout(new_new_n9031__));
  buf1  g8090(.din(new_new_n9031__), .dout(new_new_n9032__));
  buf1  g8091(.din(new_new_n9032__), .dout(new_new_n9033__));
  buf1  g8092(.din(new_new_n9033__), .dout(new_new_n9034__));
  buf1  g8093(.din(new_new_n9033__), .dout(new_new_n9035__));
  buf1  g8094(.din(new_new_n9032__), .dout(new_new_n9036__));
  buf1  g8095(.din(new_new_n9036__), .dout(new_new_n9037__));
  buf1  g8096(.din(new_new_n9036__), .dout(new_new_n9038__));
  buf1  g8097(.din(new_new_n9031__), .dout(new_new_n9039__));
  buf1  g8098(.din(new_new_n9039__), .dout(new_new_n9040__));
  buf1  g8099(.din(new_new_n9039__), .dout(new_new_n9041__));
  buf1  g8100(.din(new_new_n840__), .dout(new_new_n9042__));
  buf1  g8101(.din(new_new_n9042__), .dout(new_new_n9043__));
  buf1  g8102(.din(new_new_n843__), .dout(new_new_n9044__));
  buf1  g8103(.din(new_new_n9044__), .dout(new_new_n9045__));
  buf1  g8104(.din(new_new_n9045__), .dout(new_new_n9046__));
  buf1  g8105(.din(new_new_n9046__), .dout(new_new_n9047__));
  buf1  g8106(.din(new_new_n9046__), .dout(new_new_n9048__));
  buf1  g8107(.din(new_new_n9045__), .dout(new_new_n9049__));
  buf1  g8108(.din(new_new_n9049__), .dout(new_new_n9050__));
  buf1  g8109(.din(new_new_n9049__), .dout(new_new_n9051__));
  buf1  g8110(.din(new_new_n9044__), .dout(new_new_n9052__));
  buf1  g8111(.din(new_new_n9052__), .dout(new_new_n9053__));
  buf1  g8112(.din(new_new_n9053__), .dout(new_new_n9054__));
  buf1  g8113(.din(new_new_n9053__), .dout(new_new_n9055__));
  buf1  g8114(.din(new_new_n9052__), .dout(new_new_n9056__));
  buf1  g8115(.din(new_new_n9056__), .dout(new_new_n9057__));
  buf1  g8116(.din(new_new_n844__), .dout(new_new_n9058__));
  buf1  g8117(.din(new_new_n9058__), .dout(new_new_n9059__));
  buf1  g8118(.din(new_new_n9059__), .dout(new_new_n9060__));
  buf1  g8119(.din(new_new_n9060__), .dout(new_new_n9061__));
  buf1  g8120(.din(new_new_n9060__), .dout(new_new_n9062__));
  buf1  g8121(.din(new_new_n9059__), .dout(new_new_n9063__));
  buf1  g8122(.din(new_new_n9063__), .dout(new_new_n9064__));
  buf1  g8123(.din(new_new_n9063__), .dout(new_new_n9065__));
  buf1  g8124(.din(new_new_n9058__), .dout(new_new_n9066__));
  buf1  g8125(.din(new_new_n9066__), .dout(new_new_n9067__));
  buf1  g8126(.din(new_new_n9067__), .dout(new_new_n9068__));
  buf1  g8127(.din(new_new_n9067__), .dout(new_new_n9069__));
  buf1  g8128(.din(new_new_n9066__), .dout(new_new_n9070__));
  buf1  g8129(.din(new_new_n9070__), .dout(new_new_n9071__));
  buf1  g8130(.din(new_new_n9070__), .dout(new_new_n9072__));
  buf1  g8131(.din(new_new_n841__), .dout(new_new_n9073__));
  buf1  g8132(.din(new_new_n9073__), .dout(new_new_n9074__));
  buf1  g8133(.din(new_new_n9074__), .dout(new_new_n9075__));
  buf1  g8134(.din(new_new_n9075__), .dout(new_new_n9076__));
  buf1  g8135(.din(new_new_n9075__), .dout(new_new_n9077__));
  buf1  g8136(.din(new_new_n9074__), .dout(new_new_n9078__));
  buf1  g8137(.din(new_new_n9078__), .dout(new_new_n9079__));
  buf1  g8138(.din(new_new_n9078__), .dout(new_new_n9080__));
  buf1  g8139(.din(new_new_n9073__), .dout(new_new_n9081__));
  buf1  g8140(.din(new_new_n9081__), .dout(new_new_n9082__));
  buf1  g8141(.din(new_new_n9082__), .dout(new_new_n9083__));
  buf1  g8142(.din(new_new_n9082__), .dout(new_new_n9084__));
  buf1  g8143(.din(new_new_n9081__), .dout(new_new_n9085__));
  buf1  g8144(.din(new_new_n9085__), .dout(new_new_n9086__));
  buf1  g8145(.din(new_new_n9085__), .dout(new_new_n9087__));
  buf1  g8146(.din(new_new_n842__), .dout(new_new_n9088__));
  buf1  g8147(.din(new_new_n9088__), .dout(new_new_n9089__));
  buf1  g8148(.din(new_new_n9089__), .dout(new_new_n9090__));
  buf1  g8149(.din(new_new_n9090__), .dout(new_new_n9091__));
  buf1  g8150(.din(new_new_n9090__), .dout(new_new_n9092__));
  buf1  g8151(.din(new_new_n9089__), .dout(new_new_n9093__));
  buf1  g8152(.din(new_new_n9093__), .dout(new_new_n9094__));
  buf1  g8153(.din(new_new_n9093__), .dout(new_new_n9095__));
  buf1  g8154(.din(new_new_n9088__), .dout(new_new_n9096__));
  buf1  g8155(.din(new_new_n9096__), .dout(new_new_n9097__));
  buf1  g8156(.din(new_new_n9097__), .dout(new_new_n9098__));
  buf1  g8157(.din(new_new_n9097__), .dout(new_new_n9099__));
  buf1  g8158(.din(new_new_n9096__), .dout(new_new_n9100__));
  buf1  g8159(.din(new_new_n9100__), .dout(new_new_n9101__));
  buf1  g8160(.din(new_new_n837__), .dout(new_new_n9102__));
  buf1  g8161(.din(new_new_n9102__), .dout(new_new_n9103__));
  buf1  g8162(.din(new_new_n9103__), .dout(new_new_n9104__));
  buf1  g8163(.din(new_new_n9102__), .dout(new_new_n9105__));
  buf1  g8164(.din(new_new_n838__), .dout(new_new_n9106__));
  buf1  g8165(.din(new_new_n9106__), .dout(new_new_n9107__));
  buf1  g8166(.din(new_new_n9106__), .dout(new_new_n9108__));
  buf1  g8167(.din(new_new_n4345__), .dout(new_new_n9109__));
  buf1  g8168(.din(new_new_n4342__), .dout(new_new_n9110__));
  buf1  g8169(.din(new_new_n4344__), .dout(new_new_n9111__));
  buf1  g8170(.din(new_new_n4343__), .dout(new_new_n9112__));
  buf1  g8171(.din(new_new_n4347__), .dout(new_new_n9113__));
  buf1  g8172(.din(new_new_n4346__), .dout(new_new_n9114__));
  buf1  g8173(.din(new_new_n4349__), .dout(new_new_n9115__));
  buf1  g8174(.din(new_new_n9115__), .dout(new_new_n9116__));
  buf1  g8175(.din(new_new_n4341__), .dout(new_new_n9117__));
  buf1  g8176(.din(new_new_n4348__), .dout(new_new_n9118__));
  buf1  g8177(.din(new_new_n9118__), .dout(new_new_n9119__));
  buf1  g8178(.din(new_new_n4340__), .dout(new_new_n9120__));
  buf1  g8179(.din(new_new_n4351__), .dout(new_new_n9121__));
  buf1  g8180(.din(new_new_n9121__), .dout(new_new_n9122__));
  buf1  g8181(.din(new_new_n4350__), .dout(new_new_n9123__));
  buf1  g8182(.din(new_new_n9123__), .dout(new_new_n9124__));
  buf1  g8183(.din(new_new_n4359__), .dout(new_new_n9125__));
  buf1  g8184(.din(new_new_n4357__), .dout(new_new_n9126__));
  buf1  g8185(.din(new_new_n4358__), .dout(new_new_n9127__));
  buf1  g8186(.din(new_new_n4356__), .dout(new_new_n9128__));
  buf1  g8187(.din(new_new_n4361__), .dout(new_new_n9129__));
  buf1  g8188(.din(new_new_n9129__), .dout(new_new_n9130__));
  buf1  g8189(.din(new_new_n4360__), .dout(new_new_n9131__));
  buf1  g8190(.din(new_new_n9131__), .dout(new_new_n9132__));
  buf1  g8191(.din(new_new_n4363__), .dout(new_new_n9133__));
  buf1  g8192(.din(new_new_n4339__), .dout(new_new_n9134__));
  buf1  g8193(.din(new_new_n4362__), .dout(new_new_n9135__));
  buf1  g8194(.din(new_new_n4338__), .dout(new_new_n9136__));
  buf1  g8195(.din(new_new_n4369__), .dout(new_new_n9137__));
  buf1  g8196(.din(new_new_n4367__), .dout(new_new_n9138__));
  buf1  g8197(.din(new_new_n4368__), .dout(new_new_n9139__));
  buf1  g8198(.din(new_new_n4366__), .dout(new_new_n9140__));
  buf1  g8199(.din(new_new_n4371__), .dout(new_new_n9141__));
  buf1  g8200(.din(new_new_n9141__), .dout(new_new_n9142__));
  buf1  g8201(.din(new_new_n4370__), .dout(new_new_n9143__));
  buf1  g8202(.din(new_new_n9143__), .dout(new_new_n9144__));
  buf1  g8203(.din(new_new_n4379__), .dout(new_new_n9145__));
  buf1  g8204(.din(new_new_n4377__), .dout(new_new_n9146__));
  buf1  g8205(.din(new_new_n4378__), .dout(new_new_n9147__));
  buf1  g8206(.din(new_new_n4376__), .dout(new_new_n9148__));
  buf1  g8207(.din(new_new_n4381__), .dout(new_new_n9149__));
  buf1  g8208(.din(new_new_n9149__), .dout(new_new_n9150__));
  buf1  g8209(.din(new_new_n4380__), .dout(new_new_n9151__));
  buf1  g8210(.din(new_new_n9151__), .dout(new_new_n9152__));
  buf1  g8211(.din(new_new_n4389__), .dout(new_new_n9153__));
  buf1  g8212(.din(new_new_n4387__), .dout(new_new_n9154__));
  buf1  g8213(.din(new_new_n4388__), .dout(new_new_n9155__));
  buf1  g8214(.din(new_new_n4386__), .dout(new_new_n9156__));
  buf1  g8215(.din(new_new_n4391__), .dout(new_new_n9157__));
  buf1  g8216(.din(new_new_n9157__), .dout(new_new_n9158__));
  buf1  g8217(.din(new_new_n4390__), .dout(new_new_n9159__));
  buf1  g8218(.din(new_new_n9159__), .dout(new_new_n9160__));
  buf1  g8219(.din(new_new_n4399__), .dout(new_new_n9161__));
  buf1  g8220(.din(new_new_n4397__), .dout(new_new_n9162__));
  buf1  g8221(.din(new_new_n4398__), .dout(new_new_n9163__));
  buf1  g8222(.din(new_new_n4396__), .dout(new_new_n9164__));
  buf1  g8223(.din(new_new_n4401__), .dout(new_new_n9165__));
  buf1  g8224(.din(new_new_n9165__), .dout(new_new_n9166__));
  buf1  g8225(.din(new_new_n4400__), .dout(new_new_n9167__));
  buf1  g8226(.din(new_new_n9167__), .dout(new_new_n9168__));
  buf1  g8227(.din(new_new_n1229__), .dout(new_new_n9169__));
  buf1  g8228(.din(new_new_n9169__), .dout(new_new_n9170__));
  buf1  g8229(.din(new_new_n9170__), .dout(new_new_n9171__));
  buf1  g8230(.din(new_new_n9170__), .dout(new_new_n9172__));
  buf1  g8231(.din(new_new_n9169__), .dout(new_new_n9173__));
  buf1  g8232(.din(new_new_n9173__), .dout(new_new_n9174__));
  buf1  g8233(.din(new_new_n1230__), .dout(new_new_n9175__));
  buf1  g8234(.din(new_new_n9175__), .dout(new_new_n9176__));
  buf1  g8235(.din(new_new_n9176__), .dout(new_new_n9177__));
  buf1  g8236(.din(new_new_n9175__), .dout(new_new_n9178__));
  buf1  g8237(.din(new_new_n4414__), .dout(new_new_n9179__));
  buf1  g8238(.din(new_new_n4412__), .dout(new_new_n9180__));
  buf1  g8239(.din(new_new_n4413__), .dout(new_new_n9181__));
  buf1  g8240(.din(new_new_n4411__), .dout(new_new_n9182__));
  buf1  g8241(.din(new_new_n4416__), .dout(new_new_n9183__));
  buf1  g8242(.din(new_new_n9183__), .dout(new_new_n9184__));
  buf1  g8243(.din(new_new_n4415__), .dout(new_new_n9185__));
  buf1  g8244(.din(new_new_n9185__), .dout(new_new_n9186__));
  buf1  g8245(.din(new_new_n1599__), .dout(new_new_n9187__));
  buf1  g8246(.din(new_new_n9187__), .dout(new_new_n9188__));
  buf1  g8247(.din(new_new_n1600__), .dout(new_new_n9189__));
  buf1  g8248(.din(new_new_n9189__), .dout(new_new_n9190__));
  buf1  g8249(.din(new_new_n1253__), .dout(new_new_n9191__));
  buf1  g8250(.din(new_new_n9191__), .dout(new_new_n9192__));
  buf1  g8251(.din(new_new_n9192__), .dout(new_new_n9193__));
  buf1  g8252(.din(new_new_n9192__), .dout(new_new_n9194__));
  buf1  g8253(.din(new_new_n9191__), .dout(new_new_n9195__));
  buf1  g8254(.din(new_new_n1254__), .dout(new_new_n9196__));
  buf1  g8255(.din(new_new_n9196__), .dout(new_new_n9197__));
  buf1  g8256(.din(new_new_n9197__), .dout(new_new_n9198__));
  buf1  g8257(.din(new_new_n9196__), .dout(new_new_n9199__));
  buf1  g8258(.din(new_new_n4430__), .dout(new_new_n9200__));
  buf1  g8259(.din(new_new_n4428__), .dout(new_new_n9201__));
  buf1  g8260(.din(new_new_n4429__), .dout(new_new_n9202__));
  buf1  g8261(.din(new_new_n4427__), .dout(new_new_n9203__));
  buf1  g8262(.din(new_new_n4432__), .dout(new_new_n9204__));
  buf1  g8263(.din(new_new_n9204__), .dout(new_new_n9205__));
  buf1  g8264(.din(new_new_n4431__), .dout(new_new_n9206__));
  buf1  g8265(.din(new_new_n9206__), .dout(new_new_n9207__));
  buf1  g8266(.din(new_new_n4434__), .dout(new_new_n9208__));
  buf1  g8267(.din(new_new_n4422__), .dout(new_new_n9209__));
  buf1  g8268(.din(new_new_n4433__), .dout(new_new_n9210__));
  buf1  g8269(.din(new_new_n4421__), .dout(new_new_n9211__));
  buf1  g8270(.din(new_new_n4436__), .dout(new_new_n9212__));
  buf1  g8271(.din(new_new_n9212__), .dout(new_new_n9213__));
  buf1  g8272(.din(new_new_n4435__), .dout(new_new_n9214__));
  buf1  g8273(.din(new_new_n9214__), .dout(new_new_n9215__));
  buf1  g8274(.din(new_new_n4444__), .dout(new_new_n9216__));
  buf1  g8275(.din(new_new_n4442__), .dout(new_new_n9217__));
  buf1  g8276(.din(new_new_n4443__), .dout(new_new_n9218__));
  buf1  g8277(.din(new_new_n4441__), .dout(new_new_n9219__));
  buf1  g8278(.din(new_new_n4446__), .dout(new_new_n9220__));
  buf1  g8279(.din(new_new_n9220__), .dout(new_new_n9221__));
  buf1  g8280(.din(new_new_n4445__), .dout(new_new_n9222__));
  buf1  g8281(.din(new_new_n9222__), .dout(new_new_n9223__));
  buf1  g8282(.din(new_new_n1610__), .dout(new_new_n9224__));
  buf1  g8283(.din(new_new_n1570__), .dout(new_new_n9225__));
  buf1  g8284(.din(new_new_n1609__), .dout(new_new_n9226__));
  buf1  g8285(.din(new_new_n1569__), .dout(new_new_n9227__));
  buf1  g8286(.din(new_new_n4460__), .dout(new_new_n9228__));
  buf1  g8287(.din(new_new_n9228__), .dout(new_new_n9229__));
  buf1  g8288(.din(new_new_n4459__), .dout(new_new_n9230__));
  buf1  g8289(.din(new_new_n9230__), .dout(new_new_n9231__));
  buf1  g8290(.din(new_new_n1263__), .dout(new_new_n9232__));
  buf1  g8291(.din(new_new_n9232__), .dout(new_new_n9233__));
  buf1  g8292(.din(new_new_n9233__), .dout(new_new_n9234__));
  buf1  g8293(.din(new_new_n9233__), .dout(new_new_n9235__));
  buf1  g8294(.din(new_new_n9232__), .dout(new_new_n9236__));
  buf1  g8295(.din(new_new_n1264__), .dout(new_new_n9237__));
  buf1  g8296(.din(new_new_n9237__), .dout(new_new_n9238__));
  buf1  g8297(.din(new_new_n9238__), .dout(new_new_n9239__));
  buf1  g8298(.din(new_new_n9237__), .dout(new_new_n9240__));
  buf1  g8299(.din(new_new_n4468__), .dout(new_new_n9241__));
  buf1  g8300(.din(new_new_n4466__), .dout(new_new_n9242__));
  buf1  g8301(.din(new_new_n4467__), .dout(new_new_n9243__));
  buf1  g8302(.din(new_new_n4465__), .dout(new_new_n9244__));
  buf1  g8303(.din(new_new_n4470__), .dout(new_new_n9245__));
  buf1  g8304(.din(new_new_n9245__), .dout(new_new_n9246__));
  buf1  g8305(.din(new_new_n4469__), .dout(new_new_n9247__));
  buf1  g8306(.din(new_new_n9247__), .dout(new_new_n9248__));
  buf1  g8307(.din(new_new_n4472__), .dout(new_new_n9249__));
  buf1  g8308(.din(new_new_n4458__), .dout(new_new_n9250__));
  buf1  g8309(.din(new_new_n4471__), .dout(new_new_n9251__));
  buf1  g8310(.din(new_new_n4457__), .dout(new_new_n9252__));
  buf1  g8311(.din(new_new_n4474__), .dout(new_new_n9253__));
  buf1  g8312(.din(new_new_n9253__), .dout(new_new_n9254__));
  buf1  g8313(.din(new_new_n4473__), .dout(new_new_n9255__));
  buf1  g8314(.din(new_new_n9255__), .dout(new_new_n9256__));
  buf1  g8315(.din(new_new_n4482__), .dout(new_new_n9257__));
  buf1  g8316(.din(new_new_n4480__), .dout(new_new_n9258__));
  buf1  g8317(.din(new_new_n4481__), .dout(new_new_n9259__));
  buf1  g8318(.din(new_new_n4479__), .dout(new_new_n9260__));
  buf1  g8319(.din(new_new_n4484__), .dout(new_new_n9261__));
  buf1  g8320(.din(new_new_n9261__), .dout(new_new_n9262__));
  buf1  g8321(.din(new_new_n4483__), .dout(new_new_n9263__));
  buf1  g8322(.din(new_new_n9263__), .dout(new_new_n9264__));
  buf1  g8323(.din(new_new_n4486__), .dout(new_new_n9265__));
  buf1  g8324(.din(new_new_n4452__), .dout(new_new_n9266__));
  buf1  g8325(.din(new_new_n4485__), .dout(new_new_n9267__));
  buf1  g8326(.din(new_new_n4451__), .dout(new_new_n9268__));
  buf1  g8327(.din(new_new_n4488__), .dout(new_new_n9269__));
  buf1  g8328(.din(new_new_n9269__), .dout(new_new_n9270__));
  buf1  g8329(.din(new_new_n4487__), .dout(new_new_n9271__));
  buf1  g8330(.din(new_new_n9271__), .dout(new_new_n9272__));
  buf1  g8331(.din(new_new_n4496__), .dout(new_new_n9273__));
  buf1  g8332(.din(new_new_n4494__), .dout(new_new_n9274__));
  buf1  g8333(.din(new_new_n4495__), .dout(new_new_n9275__));
  buf1  g8334(.din(new_new_n4493__), .dout(new_new_n9276__));
  buf1  g8335(.din(new_new_n4498__), .dout(new_new_n9277__));
  buf1  g8336(.din(new_new_n9277__), .dout(new_new_n9278__));
  buf1  g8337(.din(new_new_n4497__), .dout(new_new_n9279__));
  buf1  g8338(.din(new_new_n9279__), .dout(new_new_n9280__));
  buf1  g8339(.din(new_new_n1596__), .dout(new_new_n9281__));
  buf1  g8340(.din(new_new_n9281__), .dout(new_new_n9282__));
  buf1  g8341(.din(new_new_n1595__), .dout(new_new_n9283__));
  buf1  g8342(.din(new_new_n9283__), .dout(new_new_n9284__));
  buf1  g8343(.din(new_new_n4520__), .dout(new_new_n9285__));
  buf1  g8344(.din(new_new_n4518__), .dout(new_new_n9286__));
  buf1  g8345(.din(new_new_n4519__), .dout(new_new_n9287__));
  buf1  g8346(.din(new_new_n4517__), .dout(new_new_n9288__));
  buf1  g8347(.din(new_new_n4522__), .dout(new_new_n9289__));
  buf1  g8348(.din(new_new_n9289__), .dout(new_new_n9290__));
  buf1  g8349(.din(new_new_n4521__), .dout(new_new_n9291__));
  buf1  g8350(.din(new_new_n9291__), .dout(new_new_n9292__));
  buf1  g8351(.din(new_new_n1265__), .dout(new_new_n9293__));
  buf1  g8352(.din(new_new_n9293__), .dout(new_new_n9294__));
  buf1  g8353(.din(new_new_n9294__), .dout(new_new_n9295__));
  buf1  g8354(.din(new_new_n9294__), .dout(new_new_n9296__));
  buf1  g8355(.din(new_new_n9293__), .dout(new_new_n9297__));
  buf1  g8356(.din(new_new_n1266__), .dout(new_new_n9298__));
  buf1  g8357(.din(new_new_n9298__), .dout(new_new_n9299__));
  buf1  g8358(.din(new_new_n9299__), .dout(new_new_n9300__));
  buf1  g8359(.din(new_new_n9298__), .dout(new_new_n9301__));
  buf1  g8360(.din(new_new_n4530__), .dout(new_new_n9302__));
  buf1  g8361(.din(new_new_n4528__), .dout(new_new_n9303__));
  buf1  g8362(.din(new_new_n4529__), .dout(new_new_n9304__));
  buf1  g8363(.din(new_new_n4527__), .dout(new_new_n9305__));
  buf1  g8364(.din(new_new_n4532__), .dout(new_new_n9306__));
  buf1  g8365(.din(new_new_n9306__), .dout(new_new_n9307__));
  buf1  g8366(.din(new_new_n4531__), .dout(new_new_n9308__));
  buf1  g8367(.din(new_new_n9308__), .dout(new_new_n9309__));
  buf1  g8368(.din(new_new_n4534__), .dout(new_new_n9310__));
  buf1  g8369(.din(new_new_n4516__), .dout(new_new_n9311__));
  buf1  g8370(.din(new_new_n4533__), .dout(new_new_n9312__));
  buf1  g8371(.din(new_new_n4515__), .dout(new_new_n9313__));
  buf1  g8372(.din(new_new_n4536__), .dout(new_new_n9314__));
  buf1  g8373(.din(new_new_n9314__), .dout(new_new_n9315__));
  buf1  g8374(.din(new_new_n4535__), .dout(new_new_n9316__));
  buf1  g8375(.din(new_new_n9316__), .dout(new_new_n9317__));
  buf1  g8376(.din(new_new_n4544__), .dout(new_new_n9318__));
  buf1  g8377(.din(new_new_n4542__), .dout(new_new_n9319__));
  buf1  g8378(.din(new_new_n4543__), .dout(new_new_n9320__));
  buf1  g8379(.din(new_new_n4541__), .dout(new_new_n9321__));
  buf1  g8380(.din(new_new_n4546__), .dout(new_new_n9322__));
  buf1  g8381(.din(new_new_n9322__), .dout(new_new_n9323__));
  buf1  g8382(.din(new_new_n4545__), .dout(new_new_n9324__));
  buf1  g8383(.din(new_new_n9324__), .dout(new_new_n9325__));
  buf1  g8384(.din(new_new_n4548__), .dout(new_new_n9326__));
  buf1  g8385(.din(new_new_n4510__), .dout(new_new_n9327__));
  buf1  g8386(.din(new_new_n4547__), .dout(new_new_n9328__));
  buf1  g8387(.din(new_new_n4509__), .dout(new_new_n9329__));
  buf1  g8388(.din(new_new_n4550__), .dout(new_new_n9330__));
  buf1  g8389(.din(new_new_n9330__), .dout(new_new_n9331__));
  buf1  g8390(.din(new_new_n4549__), .dout(new_new_n9332__));
  buf1  g8391(.din(new_new_n9332__), .dout(new_new_n9333__));
  buf1  g8392(.din(new_new_n4558__), .dout(new_new_n9334__));
  buf1  g8393(.din(new_new_n4556__), .dout(new_new_n9335__));
  buf1  g8394(.din(new_new_n4557__), .dout(new_new_n9336__));
  buf1  g8395(.din(new_new_n4555__), .dout(new_new_n9337__));
  buf1  g8396(.din(new_new_n4560__), .dout(new_new_n9338__));
  buf1  g8397(.din(new_new_n9338__), .dout(new_new_n9339__));
  buf1  g8398(.din(new_new_n4559__), .dout(new_new_n9340__));
  buf1  g8399(.din(new_new_n9340__), .dout(new_new_n9341__));
  buf1  g8400(.din(new_new_n4562__), .dout(new_new_n9342__));
  buf1  g8401(.din(new_new_n4504__), .dout(new_new_n9343__));
  buf1  g8402(.din(new_new_n4561__), .dout(new_new_n9344__));
  buf1  g8403(.din(new_new_n4503__), .dout(new_new_n9345__));
  buf1  g8404(.din(new_new_n4564__), .dout(new_new_n9346__));
  buf1  g8405(.din(new_new_n9346__), .dout(new_new_n9347__));
  buf1  g8406(.din(new_new_n4563__), .dout(new_new_n9348__));
  buf1  g8407(.din(new_new_n9348__), .dout(new_new_n9349__));
  buf1  g8408(.din(new_new_n4572__), .dout(new_new_n9350__));
  buf1  g8409(.din(new_new_n4570__), .dout(new_new_n9351__));
  buf1  g8410(.din(new_new_n4571__), .dout(new_new_n9352__));
  buf1  g8411(.din(new_new_n4569__), .dout(new_new_n9353__));
  buf1  g8412(.din(new_new_n4574__), .dout(new_new_n9354__));
  buf1  g8413(.din(new_new_n9354__), .dout(new_new_n9355__));
  buf1  g8414(.din(new_new_n4573__), .dout(new_new_n9356__));
  buf1  g8415(.din(new_new_n9356__), .dout(new_new_n9357__));
  buf1  g8416(.din(new_new_n4606__), .dout(new_new_n9358__));
  buf1  g8417(.din(new_new_n4604__), .dout(new_new_n9359__));
  buf1  g8418(.din(new_new_n4605__), .dout(new_new_n9360__));
  buf1  g8419(.din(new_new_n4603__), .dout(new_new_n9361__));
  buf1  g8420(.din(new_new_n4608__), .dout(new_new_n9362__));
  buf1  g8421(.din(new_new_n9362__), .dout(new_new_n9363__));
  buf1  g8422(.din(new_new_n4607__), .dout(new_new_n9364__));
  buf1  g8423(.din(new_new_n9364__), .dout(new_new_n9365__));
  buf1  g8424(.din(new_new_n1267__), .dout(new_new_n9366__));
  buf1  g8425(.din(new_new_n9366__), .dout(new_new_n9367__));
  buf1  g8426(.din(new_new_n9367__), .dout(new_new_n9368__));
  buf1  g8427(.din(new_new_n9366__), .dout(new_new_n9369__));
  buf1  g8428(.din(new_new_n1268__), .dout(new_new_n9370__));
  buf1  g8429(.din(new_new_n9370__), .dout(new_new_n9371__));
  buf1  g8430(.din(new_new_n9371__), .dout(new_new_n9372__));
  buf1  g8431(.din(new_new_n9370__), .dout(new_new_n9373__));
  buf1  g8432(.din(new_new_n4616__), .dout(new_new_n9374__));
  buf1  g8433(.din(new_new_n4614__), .dout(new_new_n9375__));
  buf1  g8434(.din(new_new_n4615__), .dout(new_new_n9376__));
  buf1  g8435(.din(new_new_n4613__), .dout(new_new_n9377__));
  buf1  g8436(.din(new_new_n4618__), .dout(new_new_n9378__));
  buf1  g8437(.din(new_new_n9378__), .dout(new_new_n9379__));
  buf1  g8438(.din(new_new_n4617__), .dout(new_new_n9380__));
  buf1  g8439(.din(new_new_n9380__), .dout(new_new_n9381__));
  buf1  g8440(.din(new_new_n4620__), .dout(new_new_n9382__));
  buf1  g8441(.din(new_new_n4598__), .dout(new_new_n9383__));
  buf1  g8442(.din(new_new_n4619__), .dout(new_new_n9384__));
  buf1  g8443(.din(new_new_n4597__), .dout(new_new_n9385__));
  buf1  g8444(.din(new_new_n4622__), .dout(new_new_n9386__));
  buf1  g8445(.din(new_new_n9386__), .dout(new_new_n9387__));
  buf1  g8446(.din(new_new_n4621__), .dout(new_new_n9388__));
  buf1  g8447(.din(new_new_n9388__), .dout(new_new_n9389__));
  buf1  g8448(.din(new_new_n4630__), .dout(new_new_n9390__));
  buf1  g8449(.din(new_new_n4628__), .dout(new_new_n9391__));
  buf1  g8450(.din(new_new_n4629__), .dout(new_new_n9392__));
  buf1  g8451(.din(new_new_n4627__), .dout(new_new_n9393__));
  buf1  g8452(.din(new_new_n4632__), .dout(new_new_n9394__));
  buf1  g8453(.din(new_new_n9394__), .dout(new_new_n9395__));
  buf1  g8454(.din(new_new_n4631__), .dout(new_new_n9396__));
  buf1  g8455(.din(new_new_n9396__), .dout(new_new_n9397__));
  buf1  g8456(.din(new_new_n4634__), .dout(new_new_n9398__));
  buf1  g8457(.din(new_new_n4592__), .dout(new_new_n9399__));
  buf1  g8458(.din(new_new_n4633__), .dout(new_new_n9400__));
  buf1  g8459(.din(new_new_n4591__), .dout(new_new_n9401__));
  buf1  g8460(.din(new_new_n4636__), .dout(new_new_n9402__));
  buf1  g8461(.din(new_new_n9402__), .dout(new_new_n9403__));
  buf1  g8462(.din(new_new_n4635__), .dout(new_new_n9404__));
  buf1  g8463(.din(new_new_n9404__), .dout(new_new_n9405__));
  buf1  g8464(.din(new_new_n4644__), .dout(new_new_n9406__));
  buf1  g8465(.din(new_new_n4642__), .dout(new_new_n9407__));
  buf1  g8466(.din(new_new_n4643__), .dout(new_new_n9408__));
  buf1  g8467(.din(new_new_n4641__), .dout(new_new_n9409__));
  buf1  g8468(.din(new_new_n4646__), .dout(new_new_n9410__));
  buf1  g8469(.din(new_new_n9410__), .dout(new_new_n9411__));
  buf1  g8470(.din(new_new_n4645__), .dout(new_new_n9412__));
  buf1  g8471(.din(new_new_n9412__), .dout(new_new_n9413__));
  buf1  g8472(.din(new_new_n4648__), .dout(new_new_n9414__));
  buf1  g8473(.din(new_new_n4586__), .dout(new_new_n9415__));
  buf1  g8474(.din(new_new_n4647__), .dout(new_new_n9416__));
  buf1  g8475(.din(new_new_n4585__), .dout(new_new_n9417__));
  buf1  g8476(.din(new_new_n4650__), .dout(new_new_n9418__));
  buf1  g8477(.din(new_new_n9418__), .dout(new_new_n9419__));
  buf1  g8478(.din(new_new_n4649__), .dout(new_new_n9420__));
  buf1  g8479(.din(new_new_n9420__), .dout(new_new_n9421__));
  buf1  g8480(.din(new_new_n4658__), .dout(new_new_n9422__));
  buf1  g8481(.din(new_new_n4656__), .dout(new_new_n9423__));
  buf1  g8482(.din(new_new_n4657__), .dout(new_new_n9424__));
  buf1  g8483(.din(new_new_n4655__), .dout(new_new_n9425__));
  buf1  g8484(.din(new_new_n4660__), .dout(new_new_n9426__));
  buf1  g8485(.din(new_new_n9426__), .dout(new_new_n9427__));
  buf1  g8486(.din(new_new_n4659__), .dout(new_new_n9428__));
  buf1  g8487(.din(new_new_n9428__), .dout(new_new_n9429__));
  buf1  g8488(.din(new_new_n1608__), .dout(new_new_n9430__));
  buf1  g8489(.din(new_new_n1572__), .dout(new_new_n9431__));
  buf1  g8490(.din(new_new_n1607__), .dout(new_new_n9432__));
  buf1  g8491(.din(new_new_n1571__), .dout(new_new_n9433__));
  buf1  g8492(.din(new_new_n4677__), .dout(new_new_n9434__));
  buf1  g8493(.din(new_new_n9434__), .dout(new_new_n9435__));
  buf1  g8494(.din(new_new_n4676__), .dout(new_new_n9436__));
  buf1  g8495(.din(new_new_n9436__), .dout(new_new_n9437__));
  buf1  g8496(.din(new_new_n1223__), .dout(new_new_n9438__));
  buf1  g8497(.din(new_new_n9438__), .dout(new_new_n9439__));
  buf1  g8498(.din(new_new_n9439__), .dout(new_new_n9440__));
  buf1  g8499(.din(new_new_n9438__), .dout(new_new_n9441__));
  buf1  g8500(.din(new_new_n1224__), .dout(new_new_n9442__));
  buf1  g8501(.din(new_new_n9442__), .dout(new_new_n9443__));
  buf1  g8502(.din(new_new_n9442__), .dout(new_new_n9444__));
  buf1  g8503(.din(new_new_n4685__), .dout(new_new_n9445__));
  buf1  g8504(.din(new_new_n4683__), .dout(new_new_n9446__));
  buf1  g8505(.din(new_new_n4684__), .dout(new_new_n9447__));
  buf1  g8506(.din(new_new_n4682__), .dout(new_new_n9448__));
  buf1  g8507(.din(new_new_n4687__), .dout(new_new_n9449__));
  buf1  g8508(.din(new_new_n9449__), .dout(new_new_n9450__));
  buf1  g8509(.din(new_new_n4686__), .dout(new_new_n9451__));
  buf1  g8510(.din(new_new_n9451__), .dout(new_new_n9452__));
  buf1  g8511(.din(new_new_n4689__), .dout(new_new_n9453__));
  buf1  g8512(.din(new_new_n4675__), .dout(new_new_n9454__));
  buf1  g8513(.din(new_new_n4688__), .dout(new_new_n9455__));
  buf1  g8514(.din(new_new_n4674__), .dout(new_new_n9456__));
  buf1  g8515(.din(new_new_n4691__), .dout(new_new_n9457__));
  buf1  g8516(.din(new_new_n9457__), .dout(new_new_n9458__));
  buf1  g8517(.din(new_new_n4690__), .dout(new_new_n9459__));
  buf1  g8518(.din(new_new_n9459__), .dout(new_new_n9460__));
  buf1  g8519(.din(new_new_n4699__), .dout(new_new_n9461__));
  buf1  g8520(.din(new_new_n4697__), .dout(new_new_n9462__));
  buf1  g8521(.din(new_new_n4698__), .dout(new_new_n9463__));
  buf1  g8522(.din(new_new_n4696__), .dout(new_new_n9464__));
  buf1  g8523(.din(new_new_n4701__), .dout(new_new_n9465__));
  buf1  g8524(.din(new_new_n9465__), .dout(new_new_n9466__));
  buf1  g8525(.din(new_new_n4700__), .dout(new_new_n9467__));
  buf1  g8526(.din(new_new_n9467__), .dout(new_new_n9468__));
  buf1  g8527(.din(new_new_n4703__), .dout(new_new_n9469__));
  buf1  g8528(.din(new_new_n4669__), .dout(new_new_n9470__));
  buf1  g8529(.din(new_new_n4702__), .dout(new_new_n9471__));
  buf1  g8530(.din(new_new_n4668__), .dout(new_new_n9472__));
  buf1  g8531(.din(new_new_n4705__), .dout(new_new_n9473__));
  buf1  g8532(.din(new_new_n9473__), .dout(new_new_n9474__));
  buf1  g8533(.din(new_new_n4704__), .dout(new_new_n9475__));
  buf1  g8534(.din(new_new_n9475__), .dout(new_new_n9476__));
  buf1  g8535(.din(new_new_n4713__), .dout(new_new_n9477__));
  buf1  g8536(.din(new_new_n4711__), .dout(new_new_n9478__));
  buf1  g8537(.din(new_new_n4712__), .dout(new_new_n9479__));
  buf1  g8538(.din(new_new_n4710__), .dout(new_new_n9480__));
  buf1  g8539(.din(new_new_n4715__), .dout(new_new_n9481__));
  buf1  g8540(.din(new_new_n9481__), .dout(new_new_n9482__));
  buf1  g8541(.din(new_new_n4714__), .dout(new_new_n9483__));
  buf1  g8542(.din(new_new_n9483__), .dout(new_new_n9484__));
  buf1  g8543(.din(new_new_n1594__), .dout(new_new_n9485__));
  buf1  g8544(.din(new_new_n9485__), .dout(new_new_n9486__));
  buf1  g8545(.din(new_new_n1593__), .dout(new_new_n9487__));
  buf1  g8546(.din(new_new_n9487__), .dout(new_new_n9488__));
  buf1  g8547(.din(new_new_n4737__), .dout(new_new_n9489__));
  buf1  g8548(.din(new_new_n4735__), .dout(new_new_n9490__));
  buf1  g8549(.din(new_new_n4736__), .dout(new_new_n9491__));
  buf1  g8550(.din(new_new_n4734__), .dout(new_new_n9492__));
  buf1  g8551(.din(new_new_n4739__), .dout(new_new_n9493__));
  buf1  g8552(.din(new_new_n9493__), .dout(new_new_n9494__));
  buf1  g8553(.din(new_new_n4738__), .dout(new_new_n9495__));
  buf1  g8554(.din(new_new_n9495__), .dout(new_new_n9496__));
  buf1  g8555(.din(new_new_n1225__), .dout(new_new_n9497__));
  buf1  g8556(.din(new_new_n9497__), .dout(new_new_n9498__));
  buf1  g8557(.din(new_new_n9498__), .dout(new_new_n9499__));
  buf1  g8558(.din(new_new_n9497__), .dout(new_new_n9500__));
  buf1  g8559(.din(new_new_n1226__), .dout(new_new_n9501__));
  buf1  g8560(.din(new_new_n9501__), .dout(new_new_n9502__));
  buf1  g8561(.din(new_new_n9501__), .dout(new_new_n9503__));
  buf1  g8562(.din(new_new_n4747__), .dout(new_new_n9504__));
  buf1  g8563(.din(new_new_n4745__), .dout(new_new_n9505__));
  buf1  g8564(.din(new_new_n4746__), .dout(new_new_n9506__));
  buf1  g8565(.din(new_new_n4744__), .dout(new_new_n9507__));
  buf1  g8566(.din(new_new_n4749__), .dout(new_new_n9508__));
  buf1  g8567(.din(new_new_n9508__), .dout(new_new_n9509__));
  buf1  g8568(.din(new_new_n4748__), .dout(new_new_n9510__));
  buf1  g8569(.din(new_new_n9510__), .dout(new_new_n9511__));
  buf1  g8570(.din(new_new_n4751__), .dout(new_new_n9512__));
  buf1  g8571(.din(new_new_n4733__), .dout(new_new_n9513__));
  buf1  g8572(.din(new_new_n4750__), .dout(new_new_n9514__));
  buf1  g8573(.din(new_new_n4732__), .dout(new_new_n9515__));
  buf1  g8574(.din(new_new_n4753__), .dout(new_new_n9516__));
  buf1  g8575(.din(new_new_n9516__), .dout(new_new_n9517__));
  buf1  g8576(.din(new_new_n4752__), .dout(new_new_n9518__));
  buf1  g8577(.din(new_new_n9518__), .dout(new_new_n9519__));
  buf1  g8578(.din(new_new_n4761__), .dout(new_new_n9520__));
  buf1  g8579(.din(new_new_n4759__), .dout(new_new_n9521__));
  buf1  g8580(.din(new_new_n4760__), .dout(new_new_n9522__));
  buf1  g8581(.din(new_new_n4758__), .dout(new_new_n9523__));
  buf1  g8582(.din(new_new_n4763__), .dout(new_new_n9524__));
  buf1  g8583(.din(new_new_n9524__), .dout(new_new_n9525__));
  buf1  g8584(.din(new_new_n4762__), .dout(new_new_n9526__));
  buf1  g8585(.din(new_new_n9526__), .dout(new_new_n9527__));
  buf1  g8586(.din(new_new_n4765__), .dout(new_new_n9528__));
  buf1  g8587(.din(new_new_n4727__), .dout(new_new_n9529__));
  buf1  g8588(.din(new_new_n4764__), .dout(new_new_n9530__));
  buf1  g8589(.din(new_new_n4726__), .dout(new_new_n9531__));
  buf1  g8590(.din(new_new_n4767__), .dout(new_new_n9532__));
  buf1  g8591(.din(new_new_n9532__), .dout(new_new_n9533__));
  buf1  g8592(.din(new_new_n4766__), .dout(new_new_n9534__));
  buf1  g8593(.din(new_new_n9534__), .dout(new_new_n9535__));
  buf1  g8594(.din(new_new_n4775__), .dout(new_new_n9536__));
  buf1  g8595(.din(new_new_n4773__), .dout(new_new_n9537__));
  buf1  g8596(.din(new_new_n4774__), .dout(new_new_n9538__));
  buf1  g8597(.din(new_new_n4772__), .dout(new_new_n9539__));
  buf1  g8598(.din(new_new_n4777__), .dout(new_new_n9540__));
  buf1  g8599(.din(new_new_n9540__), .dout(new_new_n9541__));
  buf1  g8600(.din(new_new_n4776__), .dout(new_new_n9542__));
  buf1  g8601(.din(new_new_n9542__), .dout(new_new_n9543__));
  buf1  g8602(.din(new_new_n4779__), .dout(new_new_n9544__));
  buf1  g8603(.din(new_new_n4721__), .dout(new_new_n9545__));
  buf1  g8604(.din(new_new_n4778__), .dout(new_new_n9546__));
  buf1  g8605(.din(new_new_n4720__), .dout(new_new_n9547__));
  buf1  g8606(.din(new_new_n4781__), .dout(new_new_n9548__));
  buf1  g8607(.din(new_new_n9548__), .dout(new_new_n9549__));
  buf1  g8608(.din(new_new_n4780__), .dout(new_new_n9550__));
  buf1  g8609(.din(new_new_n9550__), .dout(new_new_n9551__));
  buf1  g8610(.din(new_new_n899__), .dout(new_new_n9552__));
  buf1  g8611(.din(new_new_n9552__), .dout(new_new_n9553__));
  buf1  g8612(.din(new_new_n9553__), .dout(new_new_n9554__));
  buf1  g8613(.din(new_new_n9554__), .dout(new_new_n9555__));
  buf1  g8614(.din(new_new_n9554__), .dout(new_new_n9556__));
  buf1  g8615(.din(new_new_n9553__), .dout(new_new_n9557__));
  buf1  g8616(.din(new_new_n9552__), .dout(new_new_n9558__));
  buf1  g8617(.din(new_new_n9558__), .dout(new_new_n9559__));
  buf1  g8618(.din(new_new_n9558__), .dout(new_new_n9560__));
  buf1  g8619(.din(new_new_n900__), .dout(new_new_n9561__));
  buf1  g8620(.din(new_new_n9561__), .dout(new_new_n9562__));
  buf1  g8621(.din(new_new_n9562__), .dout(new_new_n9563__));
  buf1  g8622(.din(new_new_n9563__), .dout(new_new_n9564__));
  buf1  g8623(.din(new_new_n9563__), .dout(new_new_n9565__));
  buf1  g8624(.din(new_new_n9562__), .dout(new_new_n9566__));
  buf1  g8625(.din(new_new_n9561__), .dout(new_new_n9567__));
  buf1  g8626(.din(new_new_n9567__), .dout(new_new_n9568__));
  buf1  g8627(.din(new_new_n9567__), .dout(new_new_n9569__));
  buf1  g8628(.din(new_new_n4789__), .dout(new_new_n9570__));
  buf1  g8629(.din(new_new_n4787__), .dout(new_new_n9571__));
  buf1  g8630(.din(new_new_n4788__), .dout(new_new_n9572__));
  buf1  g8631(.din(new_new_n4786__), .dout(new_new_n9573__));
  buf1  g8632(.din(new_new_n4791__), .dout(new_new_n9574__));
  buf1  g8633(.din(new_new_n9574__), .dout(new_new_n9575__));
  buf1  g8634(.din(new_new_n4790__), .dout(new_new_n9576__));
  buf1  g8635(.din(new_new_n9576__), .dout(new_new_n9577__));
  buf1  g8636(.din(new_new_n1613__), .dout(new_new_n9578__));
  buf1  g8637(.din(new_new_n1562__), .dout(new_new_n9579__));
  buf1  g8638(.din(new_new_n1614__), .dout(new_new_n9580__));
  buf1  g8639(.din(new_new_n1561__), .dout(new_new_n9581__));
  buf1  g8640(.din(new_new_n4823__), .dout(new_new_n9582__));
  buf1  g8641(.din(new_new_n9582__), .dout(new_new_n9583__));
  buf1  g8642(.din(new_new_n4822__), .dout(new_new_n9584__));
  buf1  g8643(.din(new_new_n9584__), .dout(new_new_n9585__));
  buf1  g8644(.din(new_new_n4825__), .dout(new_new_n9586__));
  buf1  g8645(.din(new_new_n4821__), .dout(new_new_n9587__));
  buf1  g8646(.din(new_new_n4824__), .dout(new_new_n9588__));
  buf1  g8647(.din(new_new_n4820__), .dout(new_new_n9589__));
  buf1  g8648(.din(new_new_n4827__), .dout(new_new_n9590__));
  buf1  g8649(.din(new_new_n9590__), .dout(new_new_n9591__));
  buf1  g8650(.din(new_new_n4826__), .dout(new_new_n9592__));
  buf1  g8651(.din(new_new_n9592__), .dout(new_new_n9593__));
  buf1  g8652(.din(new_new_n1227__), .dout(new_new_n9594__));
  buf1  g8653(.din(new_new_n9594__), .dout(new_new_n9595__));
  buf1  g8654(.din(new_new_n9595__), .dout(new_new_n9596__));
  buf1  g8655(.din(new_new_n9594__), .dout(new_new_n9597__));
  buf1  g8656(.din(new_new_n1228__), .dout(new_new_n9598__));
  buf1  g8657(.din(new_new_n9598__), .dout(new_new_n9599__));
  buf1  g8658(.din(new_new_n9599__), .dout(new_new_n9600__));
  buf1  g8659(.din(new_new_n9598__), .dout(new_new_n9601__));
  buf1  g8660(.din(new_new_n4835__), .dout(new_new_n9602__));
  buf1  g8661(.din(new_new_n4833__), .dout(new_new_n9603__));
  buf1  g8662(.din(new_new_n4834__), .dout(new_new_n9604__));
  buf1  g8663(.din(new_new_n4832__), .dout(new_new_n9605__));
  buf1  g8664(.din(new_new_n4837__), .dout(new_new_n9606__));
  buf1  g8665(.din(new_new_n9606__), .dout(new_new_n9607__));
  buf1  g8666(.din(new_new_n4836__), .dout(new_new_n9608__));
  buf1  g8667(.din(new_new_n9608__), .dout(new_new_n9609__));
  buf1  g8668(.din(new_new_n4839__), .dout(new_new_n9610__));
  buf1  g8669(.din(new_new_n4815__), .dout(new_new_n9611__));
  buf1  g8670(.din(new_new_n4838__), .dout(new_new_n9612__));
  buf1  g8671(.din(new_new_n4814__), .dout(new_new_n9613__));
  buf1  g8672(.din(new_new_n4841__), .dout(new_new_n9614__));
  buf1  g8673(.din(new_new_n9614__), .dout(new_new_n9615__));
  buf1  g8674(.din(new_new_n4840__), .dout(new_new_n9616__));
  buf1  g8675(.din(new_new_n9616__), .dout(new_new_n9617__));
  buf1  g8676(.din(new_new_n4849__), .dout(new_new_n9618__));
  buf1  g8677(.din(new_new_n4847__), .dout(new_new_n9619__));
  buf1  g8678(.din(new_new_n4848__), .dout(new_new_n9620__));
  buf1  g8679(.din(new_new_n4846__), .dout(new_new_n9621__));
  buf1  g8680(.din(new_new_n4851__), .dout(new_new_n9622__));
  buf1  g8681(.din(new_new_n9622__), .dout(new_new_n9623__));
  buf1  g8682(.din(new_new_n4850__), .dout(new_new_n9624__));
  buf1  g8683(.din(new_new_n9624__), .dout(new_new_n9625__));
  buf1  g8684(.din(new_new_n4853__), .dout(new_new_n9626__));
  buf1  g8685(.din(new_new_n4809__), .dout(new_new_n9627__));
  buf1  g8686(.din(new_new_n4852__), .dout(new_new_n9628__));
  buf1  g8687(.din(new_new_n4808__), .dout(new_new_n9629__));
  buf1  g8688(.din(new_new_n4855__), .dout(new_new_n9630__));
  buf1  g8689(.din(new_new_n9630__), .dout(new_new_n9631__));
  buf1  g8690(.din(new_new_n4854__), .dout(new_new_n9632__));
  buf1  g8691(.din(new_new_n9632__), .dout(new_new_n9633__));
  buf1  g8692(.din(new_new_n4863__), .dout(new_new_n9634__));
  buf1  g8693(.din(new_new_n4861__), .dout(new_new_n9635__));
  buf1  g8694(.din(new_new_n4862__), .dout(new_new_n9636__));
  buf1  g8695(.din(new_new_n4860__), .dout(new_new_n9637__));
  buf1  g8696(.din(new_new_n4865__), .dout(new_new_n9638__));
  buf1  g8697(.din(new_new_n9638__), .dout(new_new_n9639__));
  buf1  g8698(.din(new_new_n4864__), .dout(new_new_n9640__));
  buf1  g8699(.din(new_new_n9640__), .dout(new_new_n9641__));
  buf1  g8700(.din(new_new_n4867__), .dout(new_new_n9642__));
  buf1  g8701(.din(new_new_n4803__), .dout(new_new_n9643__));
  buf1  g8702(.din(new_new_n4866__), .dout(new_new_n9644__));
  buf1  g8703(.din(new_new_n4802__), .dout(new_new_n9645__));
  buf1  g8704(.din(new_new_n4869__), .dout(new_new_n9646__));
  buf1  g8705(.din(new_new_n9646__), .dout(new_new_n9647__));
  buf1  g8706(.din(new_new_n4868__), .dout(new_new_n9648__));
  buf1  g8707(.din(new_new_n9648__), .dout(new_new_n9649__));
  buf1  g8708(.din(new_new_n4877__), .dout(new_new_n9650__));
  buf1  g8709(.din(new_new_n4875__), .dout(new_new_n9651__));
  buf1  g8710(.din(new_new_n4876__), .dout(new_new_n9652__));
  buf1  g8711(.din(new_new_n4874__), .dout(new_new_n9653__));
  buf1  g8712(.din(new_new_n4879__), .dout(new_new_n9654__));
  buf1  g8713(.din(new_new_n9654__), .dout(new_new_n9655__));
  buf1  g8714(.din(new_new_n4878__), .dout(new_new_n9656__));
  buf1  g8715(.din(new_new_n9656__), .dout(new_new_n9657__));
  buf1  g8716(.din(new_new_n4890__), .dout(new_new_n9658__));
  buf1  g8717(.din(new_new_n4888__), .dout(new_new_n9659__));
  buf1  g8718(.din(new_new_n4889__), .dout(new_new_n9660__));
  buf1  g8719(.din(new_new_n4887__), .dout(new_new_n9661__));
  buf1  g8720(.din(new_new_n4892__), .dout(new_new_n9662__));
  buf1  g8721(.din(new_new_n9662__), .dout(new_new_n9663__));
  buf1  g8722(.din(new_new_n4891__), .dout(new_new_n9664__));
  buf1  g8723(.din(new_new_n9664__), .dout(new_new_n9665__));
  buf1  g8724(.din(new_new_n4900__), .dout(new_new_n9666__));
  buf1  g8725(.din(new_new_n4898__), .dout(new_new_n9667__));
  buf1  g8726(.din(new_new_n4899__), .dout(new_new_n9668__));
  buf1  g8727(.din(new_new_n4897__), .dout(new_new_n9669__));
  buf1  g8728(.din(new_new_n4902__), .dout(new_new_n9670__));
  buf1  g8729(.din(new_new_n9670__), .dout(new_new_n9671__));
  buf1  g8730(.din(new_new_n4901__), .dout(new_new_n9672__));
  buf1  g8731(.din(new_new_n9672__), .dout(new_new_n9673__));
  buf1  g8732(.din(new_new_n4910__), .dout(new_new_n9674__));
  buf1  g8733(.din(new_new_n4908__), .dout(new_new_n9675__));
  buf1  g8734(.din(new_new_n4909__), .dout(new_new_n9676__));
  buf1  g8735(.din(new_new_n4907__), .dout(new_new_n9677__));
  buf1  g8736(.din(new_new_n4912__), .dout(new_new_n9678__));
  buf1  g8737(.din(new_new_n9678__), .dout(new_new_n9679__));
  buf1  g8738(.din(new_new_n4911__), .dout(new_new_n9680__));
  buf1  g8739(.din(new_new_n9680__), .dout(new_new_n9681__));
  buf1  g8740(.din(new_new_n4920__), .dout(new_new_n9682__));
  buf1  g8741(.din(new_new_n4918__), .dout(new_new_n9683__));
  buf1  g8742(.din(new_new_n4919__), .dout(new_new_n9684__));
  buf1  g8743(.din(new_new_n4917__), .dout(new_new_n9685__));
  buf1  g8744(.din(new_new_n4922__), .dout(new_new_n9686__));
  buf1  g8745(.din(new_new_n9686__), .dout(new_new_n9687__));
  buf1  g8746(.din(new_new_n4921__), .dout(new_new_n9688__));
  buf1  g8747(.din(new_new_n9688__), .dout(new_new_n9689__));
  buf1  g8748(.din(new_new_n3716__), .dout(new_new_n9690__));
  buf1  g8749(.din(new_new_n4930__), .dout(new_new_n9691__));
  buf1  g8750(.din(new_new_n4928__), .dout(new_new_n9692__));
  buf1  g8751(.din(new_new_n4932__), .dout(new_new_n9693__));
  buf1  g8752(.din(new_new_n3822__), .dout(new_new_n9694__));
  buf1  g8753(.din(new_new_n9694__), .dout(new_new_n9695__));
  buf1  g8754(.din(new_new_n3851__), .dout(new_new_n9696__));
  buf1  g8755(.din(new_new_n9696__), .dout(new_new_n9697__));
  buf1  g8756(.din(new_new_n3880__), .dout(new_new_n9698__));
  buf1  g8757(.din(new_new_n9698__), .dout(new_new_n9699__));
  buf1  g8758(.din(new_new_n3889__), .dout(new_new_n9700__));
  buf1  g8759(.din(new_new_n3790__), .dout(new_new_n9701__));
  buf1  g8760(.din(new_new_n3886__), .dout(new_new_n9702__));
  buf1  g8761(.din(new_new_n3791__), .dout(new_new_n9703__));
  buf1  g8762(.din(new_new_n3883__), .dout(new_new_n9704__));
  buf1  g8763(.din(new_new_n3792__), .dout(new_new_n9705__));
  buf1  g8764(.din(new_new_n3892__), .dout(new_new_n9706__));
  buf1  g8765(.din(new_new_n3793__), .dout(new_new_n9707__));
  buf1  g8766(.din(new_new_n3144__), .dout(new_new_n9708__));
  buf1  g8767(.din(new_new_n9708__), .dout(new_new_n9709__));
  buf1  g8768(.din(new_new_n3153__), .dout(new_new_n9710__));
  buf1  g8769(.din(new_new_n9710__), .dout(new_new_n9711__));
  buf1  g8770(.din(new_new_n3162__), .dout(new_new_n9712__));
  buf1  g8771(.din(new_new_n9712__), .dout(new_new_n9713__));
  buf1  g8772(.din(new_new_n4974__), .dout(new_new_n9714__));
  buf1  g8773(.din(new_new_n4972__), .dout(new_new_n9715__));
  buf1  g8774(.din(new_new_n4973__), .dout(new_new_n9716__));
  buf1  g8775(.din(new_new_n4971__), .dout(new_new_n9717__));
  buf1  g8776(.din(new_new_n4976__), .dout(new_new_n9718__));
  buf1  g8777(.din(new_new_n9718__), .dout(new_new_n9719__));
  buf1  g8778(.din(new_new_n4975__), .dout(new_new_n9720__));
  buf1  g8779(.din(new_new_n4984__), .dout(new_new_n9721__));
  buf1  g8780(.din(new_new_n4982__), .dout(new_new_n9722__));
  buf1  g8781(.din(new_new_n4983__), .dout(new_new_n9723__));
  buf1  g8782(.din(new_new_n4981__), .dout(new_new_n9724__));
  buf1  g8783(.din(new_new_n4986__), .dout(new_new_n9725__));
  buf1  g8784(.din(new_new_n9725__), .dout(new_new_n9726__));
  buf1  g8785(.din(new_new_n4985__), .dout(new_new_n9727__));
  buf1  g8786(.din(new_new_n5003__), .dout(new_new_n9728__));
  buf1  g8787(.din(new_new_n5001__), .dout(new_new_n9729__));
  buf1  g8788(.din(new_new_n5002__), .dout(new_new_n9730__));
  buf1  g8789(.din(new_new_n5000__), .dout(new_new_n9731__));
  buf1  g8790(.din(new_new_n5005__), .dout(new_new_n9732__));
  buf1  g8791(.din(new_new_n9732__), .dout(new_new_n9733__));
  buf1  g8792(.din(new_new_n5004__), .dout(new_new_n9734__));
  buf1  g8793(.din(new_new_n5013__), .dout(new_new_n9735__));
  buf1  g8794(.din(new_new_n5011__), .dout(new_new_n9736__));
  buf1  g8795(.din(new_new_n5012__), .dout(new_new_n9737__));
  buf1  g8796(.din(new_new_n5010__), .dout(new_new_n9738__));
  buf1  g8797(.din(new_new_n5015__), .dout(new_new_n9739__));
  buf1  g8798(.din(new_new_n9739__), .dout(new_new_n9740__));
  buf1  g8799(.din(new_new_n5014__), .dout(new_new_n9741__));
  buf1  g8800(.din(new_new_n3893__), .dout(new_new_n9742__));
  buf1  g8801(.din(new_new_n3919__), .dout(new_new_n9743__));
  buf1  g8802(.din(new_new_n9743__), .dout(new_new_n9744__));
  buf1  g8803(.din(new_new_n3968__), .dout(new_new_n9745__));
  buf1  g8804(.din(new_new_n9745__), .dout(new_new_n9746__));
  buf1  g8805(.din(new_new_n4017__), .dout(new_new_n9747__));
  buf1  g8806(.din(new_new_n9747__), .dout(new_new_n9748__));
  buf1  g8807(.din(new_new_n4126__), .dout(new_new_n9749__));
  buf1  g8808(.din(new_new_n9749__), .dout(new_new_n9750__));
  buf1  g8809(.din(new_new_n4280__), .dout(new_new_n9751__));
  buf1  g8810(.din(new_new_n9751__), .dout(new_new_n9752__));
  buf1  g8811(.din(new_new_n4279__), .dout(new_new_n9753__));
  buf1  g8812(.din(new_new_n4935__), .dout(new_new_n9754__));
  buf1  g8813(.din(new_new_n4337__), .dout(new_new_n9755__));
  buf1  g8814(.din(new_new_n5075__), .dout(new_new_n9756__));
  buf1  g8815(.din(new_new_n5073__), .dout(new_new_n9757__));
  buf1  g8816(.din(new_new_n5074__), .dout(new_new_n9758__));
  buf1  g8817(.din(new_new_n5072__), .dout(new_new_n9759__));
  buf1  g8818(.din(new_new_n5077__), .dout(new_new_n9760__));
  buf1  g8819(.din(new_new_n9760__), .dout(new_new_n9761__));
  buf1  g8820(.din(new_new_n5076__), .dout(new_new_n9762__));
  buf1  g8821(.din(new_new_n9762__), .dout(new_new_n9763__));
  buf1  g8822(.din(new_new_n5085__), .dout(new_new_n9764__));
  buf1  g8823(.din(new_new_n5083__), .dout(new_new_n9765__));
  buf1  g8824(.din(new_new_n5084__), .dout(new_new_n9766__));
  buf1  g8825(.din(new_new_n5082__), .dout(new_new_n9767__));
  buf1  g8826(.din(new_new_n5087__), .dout(new_new_n9768__));
  buf1  g8827(.din(new_new_n9768__), .dout(new_new_n9769__));
  buf1  g8828(.din(new_new_n5086__), .dout(new_new_n9770__));
  buf1  g8829(.din(new_new_n9770__), .dout(new_new_n9771__));
  buf1  g8830(.din(new_new_n5089__), .dout(new_new_n9772__));
  buf1  g8831(.din(new_new_n5067__), .dout(new_new_n9773__));
  buf1  g8832(.din(new_new_n5088__), .dout(new_new_n9774__));
  buf1  g8833(.din(new_new_n5066__), .dout(new_new_n9775__));
  buf1  g8834(.din(new_new_n5091__), .dout(new_new_n9776__));
  buf1  g8835(.din(new_new_n9776__), .dout(new_new_n9777__));
  buf1  g8836(.din(new_new_n5090__), .dout(new_new_n9778__));
  buf1  g8837(.din(new_new_n9778__), .dout(new_new_n9779__));
  buf1  g8838(.din(new_new_n5099__), .dout(new_new_n9780__));
  buf1  g8839(.din(new_new_n5097__), .dout(new_new_n9781__));
  buf1  g8840(.din(new_new_n5098__), .dout(new_new_n9782__));
  buf1  g8841(.din(new_new_n5096__), .dout(new_new_n9783__));
  buf1  g8842(.din(new_new_n5101__), .dout(new_new_n9784__));
  buf1  g8843(.din(new_new_n9784__), .dout(new_new_n9785__));
  buf1  g8844(.din(new_new_n5100__), .dout(new_new_n9786__));
  buf1  g8845(.din(new_new_n9786__), .dout(new_new_n9787__));
  buf1  g8846(.din(new_new_n5136__), .dout(new_new_n9788__));
  buf1  g8847(.din(new_new_n5134__), .dout(new_new_n9789__));
  buf1  g8848(.din(new_new_n5135__), .dout(new_new_n9790__));
  buf1  g8849(.din(new_new_n5133__), .dout(new_new_n9791__));
  buf1  g8850(.din(new_new_n5138__), .dout(new_new_n9792__));
  buf1  g8851(.din(new_new_n9792__), .dout(new_new_n9793__));
  buf1  g8852(.din(new_new_n5137__), .dout(new_new_n9794__));
  buf1  g8853(.din(new_new_n9794__), .dout(new_new_n9795__));
  buf1  g8854(.din(new_new_n5146__), .dout(new_new_n9796__));
  buf1  g8855(.din(new_new_n5144__), .dout(new_new_n9797__));
  buf1  g8856(.din(new_new_n5145__), .dout(new_new_n9798__));
  buf1  g8857(.din(new_new_n5143__), .dout(new_new_n9799__));
  buf1  g8858(.din(new_new_n5148__), .dout(new_new_n9800__));
  buf1  g8859(.din(new_new_n9800__), .dout(new_new_n9801__));
  buf1  g8860(.din(new_new_n5147__), .dout(new_new_n9802__));
  buf1  g8861(.din(new_new_n9802__), .dout(new_new_n9803__));
  buf1  g8862(.din(new_new_n5150__), .dout(new_new_n9804__));
  buf1  g8863(.din(new_new_n5128__), .dout(new_new_n9805__));
  buf1  g8864(.din(new_new_n5149__), .dout(new_new_n9806__));
  buf1  g8865(.din(new_new_n5127__), .dout(new_new_n9807__));
  buf1  g8866(.din(new_new_n5152__), .dout(new_new_n9808__));
  buf1  g8867(.din(new_new_n9808__), .dout(new_new_n9809__));
  buf1  g8868(.din(new_new_n5151__), .dout(new_new_n9810__));
  buf1  g8869(.din(new_new_n9810__), .dout(new_new_n9811__));
  buf1  g8870(.din(new_new_n5160__), .dout(new_new_n9812__));
  buf1  g8871(.din(new_new_n5158__), .dout(new_new_n9813__));
  buf1  g8872(.din(new_new_n5159__), .dout(new_new_n9814__));
  buf1  g8873(.din(new_new_n5157__), .dout(new_new_n9815__));
  buf1  g8874(.din(new_new_n5162__), .dout(new_new_n9816__));
  buf1  g8875(.din(new_new_n9816__), .dout(new_new_n9817__));
  buf1  g8876(.din(new_new_n5161__), .dout(new_new_n9818__));
  buf1  g8877(.din(new_new_n9818__), .dout(new_new_n9819__));
  buf1  g8878(.din(new_new_n5164__), .dout(new_new_n9820__));
  buf1  g8879(.din(new_new_n5122__), .dout(new_new_n9821__));
  buf1  g8880(.din(new_new_n5163__), .dout(new_new_n9822__));
  buf1  g8881(.din(new_new_n5121__), .dout(new_new_n9823__));
  buf1  g8882(.din(new_new_n5166__), .dout(new_new_n9824__));
  buf1  g8883(.din(new_new_n9824__), .dout(new_new_n9825__));
  buf1  g8884(.din(new_new_n5165__), .dout(new_new_n9826__));
  buf1  g8885(.din(new_new_n9826__), .dout(new_new_n9827__));
  buf1  g8886(.din(new_new_n5174__), .dout(new_new_n9828__));
  buf1  g8887(.din(new_new_n5172__), .dout(new_new_n9829__));
  buf1  g8888(.din(new_new_n5173__), .dout(new_new_n9830__));
  buf1  g8889(.din(new_new_n5171__), .dout(new_new_n9831__));
  buf1  g8890(.din(new_new_n5176__), .dout(new_new_n9832__));
  buf1  g8891(.din(new_new_n9832__), .dout(new_new_n9833__));
  buf1  g8892(.din(new_new_n5175__), .dout(new_new_n9834__));
  buf1  g8893(.din(new_new_n9834__), .dout(new_new_n9835__));
  buf1  g8894(.din(new_new_n5178__), .dout(new_new_n9836__));
  buf1  g8895(.din(new_new_n5116__), .dout(new_new_n9837__));
  buf1  g8896(.din(new_new_n5177__), .dout(new_new_n9838__));
  buf1  g8897(.din(new_new_n5115__), .dout(new_new_n9839__));
  buf1  g8898(.din(new_new_n5180__), .dout(new_new_n9840__));
  buf1  g8899(.din(new_new_n9840__), .dout(new_new_n9841__));
  buf1  g8900(.din(new_new_n5179__), .dout(new_new_n9842__));
  buf1  g8901(.din(new_new_n9842__), .dout(new_new_n9843__));
  buf1  g8902(.din(new_new_n5188__), .dout(new_new_n9844__));
  buf1  g8903(.din(new_new_n5186__), .dout(new_new_n9845__));
  buf1  g8904(.din(new_new_n5187__), .dout(new_new_n9846__));
  buf1  g8905(.din(new_new_n5185__), .dout(new_new_n9847__));
  buf1  g8906(.din(new_new_n5190__), .dout(new_new_n9848__));
  buf1  g8907(.din(new_new_n9848__), .dout(new_new_n9849__));
  buf1  g8908(.din(new_new_n5189__), .dout(new_new_n9850__));
  buf1  g8909(.din(new_new_n9850__), .dout(new_new_n9851__));
  buf1  g8910(.din(new_new_n821__), .dout(new_new_n9852__));
  buf1  g8911(.din(new_new_n9852__), .dout(new_new_n9853__));
  buf1  g8912(.din(new_new_n9852__), .dout(new_new_n9854__));
  buf1  g8913(.din(new_new_n822__), .dout(new_new_n9855__));
  buf1  g8914(.din(new_new_n9855__), .dout(new_new_n9856__));
  buf1  g8915(.din(new_new_n819__), .dout(new_new_n9857__));
  buf1  g8916(.din(new_new_n9857__), .dout(new_new_n9858__));
  buf1  g8917(.din(new_new_n9857__), .dout(new_new_n9859__));
  buf1  g8918(.din(new_new_n820__), .dout(new_new_n9860__));
  buf1  g8919(.din(new_new_n9860__), .dout(new_new_n9861__));
  buf1  g8920(.din(new_new_n5197__), .dout(new_new_n9862__));
  buf1  g8921(.din(new_new_n5194__), .dout(new_new_n9863__));
  buf1  g8922(.din(new_new_n5196__), .dout(new_new_n9864__));
  buf1  g8923(.din(new_new_n5195__), .dout(new_new_n9865__));
  buf1  g8924(.din(new_new_n5199__), .dout(new_new_n9866__));
  buf1  g8925(.din(new_new_n5198__), .dout(new_new_n9867__));
  buf1  g8926(.din(new_new_n5201__), .dout(new_new_n9868__));
  buf1  g8927(.din(new_new_n9868__), .dout(new_new_n9869__));
  buf1  g8928(.din(new_new_n5200__), .dout(new_new_n9870__));
  buf1  g8929(.din(new_new_n9870__), .dout(new_new_n9871__));
  buf1  g8930(.din(new_new_n817__), .dout(new_new_n9872__));
  buf1  g8931(.din(new_new_n9872__), .dout(new_new_n9873__));
  buf1  g8932(.din(new_new_n818__), .dout(new_new_n9874__));
  buf1  g8933(.din(new_new_n9874__), .dout(new_new_n9875__));
  buf1  g8934(.din(new_new_n5209__), .dout(new_new_n9876__));
  buf1  g8935(.din(new_new_n5206__), .dout(new_new_n9877__));
  buf1  g8936(.din(new_new_n5208__), .dout(new_new_n9878__));
  buf1  g8937(.din(new_new_n5207__), .dout(new_new_n9879__));
  buf1  g8938(.din(new_new_n5211__), .dout(new_new_n9880__));
  buf1  g8939(.din(new_new_n5210__), .dout(new_new_n9881__));
  buf1  g8940(.din(new_new_n5212__), .dout(new_new_n9882__));
  buf1  g8941(.din(new_new_n833__), .dout(new_new_n9883__));
  buf1  g8942(.din(new_new_n9883__), .dout(new_new_n9884__));
  buf1  g8943(.din(new_new_n9884__), .dout(new_new_n9885__));
  buf1  g8944(.din(new_new_n9883__), .dout(new_new_n9886__));
  buf1  g8945(.din(new_new_n834__), .dout(new_new_n9887__));
  buf1  g8946(.din(new_new_n9887__), .dout(new_new_n9888__));
  buf1  g8947(.din(new_new_n9887__), .dout(new_new_n9889__));
  buf1  g8948(.din(new_new_n831__), .dout(new_new_n9890__));
  buf1  g8949(.din(new_new_n9890__), .dout(new_new_n9891__));
  buf1  g8950(.din(new_new_n9891__), .dout(new_new_n9892__));
  buf1  g8951(.din(new_new_n9890__), .dout(new_new_n9893__));
  buf1  g8952(.din(new_new_n832__), .dout(new_new_n9894__));
  buf1  g8953(.din(new_new_n9894__), .dout(new_new_n9895__));
  buf1  g8954(.din(new_new_n9894__), .dout(new_new_n9896__));
  buf1  g8955(.din(new_new_n5218__), .dout(new_new_n9897__));
  buf1  g8956(.din(new_new_n5215__), .dout(new_new_n9898__));
  buf1  g8957(.din(new_new_n5217__), .dout(new_new_n9899__));
  buf1  g8958(.din(new_new_n5216__), .dout(new_new_n9900__));
  buf1  g8959(.din(new_new_n5220__), .dout(new_new_n9901__));
  buf1  g8960(.din(new_new_n5219__), .dout(new_new_n9902__));
  buf1  g8961(.din(new_new_n5222__), .dout(new_new_n9903__));
  buf1  g8962(.din(new_new_n9903__), .dout(new_new_n9904__));
  buf1  g8963(.din(new_new_n5221__), .dout(new_new_n9905__));
  buf1  g8964(.din(new_new_n9905__), .dout(new_new_n9906__));
  buf1  g8965(.din(new_new_n829__), .dout(new_new_n9907__));
  buf1  g8966(.din(new_new_n9907__), .dout(new_new_n9908__));
  buf1  g8967(.din(new_new_n9908__), .dout(new_new_n9909__));
  buf1  g8968(.din(new_new_n9907__), .dout(new_new_n9910__));
  buf1  g8969(.din(new_new_n830__), .dout(new_new_n9911__));
  buf1  g8970(.din(new_new_n9911__), .dout(new_new_n9912__));
  buf1  g8971(.din(new_new_n9911__), .dout(new_new_n9913__));
  buf1  g8972(.din(new_new_n5230__), .dout(new_new_n9914__));
  buf1  g8973(.din(new_new_n5227__), .dout(new_new_n9915__));
  buf1  g8974(.din(new_new_n5229__), .dout(new_new_n9916__));
  buf1  g8975(.din(new_new_n5228__), .dout(new_new_n9917__));
  buf1  g8976(.din(new_new_n5232__), .dout(new_new_n9918__));
  buf1  g8977(.din(new_new_n5231__), .dout(new_new_n9919__));
  buf1  g8978(.din(new_new_n5234__), .dout(new_new_n9920__));
  buf1  g8979(.din(new_new_n9920__), .dout(new_new_n9921__));
  buf1  g8980(.din(new_new_n5226__), .dout(new_new_n9922__));
  buf1  g8981(.din(new_new_n5233__), .dout(new_new_n9923__));
  buf1  g8982(.din(new_new_n9923__), .dout(new_new_n9924__));
  buf1  g8983(.din(new_new_n5225__), .dout(new_new_n9925__));
  buf1  g8984(.din(new_new_n5236__), .dout(new_new_n9926__));
  buf1  g8985(.din(new_new_n9926__), .dout(new_new_n9927__));
  buf1  g8986(.din(new_new_n5235__), .dout(new_new_n9928__));
  buf1  g8987(.din(new_new_n9928__), .dout(new_new_n9929__));
  buf1  g8988(.din(new_new_n5244__), .dout(new_new_n9930__));
  buf1  g8989(.din(new_new_n5242__), .dout(new_new_n9931__));
  buf1  g8990(.din(new_new_n5243__), .dout(new_new_n9932__));
  buf1  g8991(.din(new_new_n5241__), .dout(new_new_n9933__));
  buf1  g8992(.din(new_new_n5246__), .dout(new_new_n9934__));
  buf1  g8993(.din(new_new_n9934__), .dout(new_new_n9935__));
  buf1  g8994(.din(new_new_n5245__), .dout(new_new_n9936__));
  buf1  g8995(.din(new_new_n9936__), .dout(new_new_n9937__));
  buf1  g8996(.din(new_new_n827__), .dout(new_new_n9938__));
  buf1  g8997(.din(new_new_n9938__), .dout(new_new_n9939__));
  buf1  g8998(.din(new_new_n9938__), .dout(new_new_n9940__));
  buf1  g8999(.din(new_new_n828__), .dout(new_new_n9941__));
  buf1  g9000(.din(new_new_n9941__), .dout(new_new_n9942__));
  buf1  g9001(.din(new_new_n9941__), .dout(new_new_n9943__));
  buf1  g9002(.din(new_new_n5260__), .dout(new_new_n9944__));
  buf1  g9003(.din(new_new_n5257__), .dout(new_new_n9945__));
  buf1  g9004(.din(new_new_n5259__), .dout(new_new_n9946__));
  buf1  g9005(.din(new_new_n5258__), .dout(new_new_n9947__));
  buf1  g9006(.din(new_new_n5262__), .dout(new_new_n9948__));
  buf1  g9007(.din(new_new_n5261__), .dout(new_new_n9949__));
  buf1  g9008(.din(new_new_n5264__), .dout(new_new_n9950__));
  buf1  g9009(.din(new_new_n9950__), .dout(new_new_n9951__));
  buf1  g9010(.din(new_new_n5256__), .dout(new_new_n9952__));
  buf1  g9011(.din(new_new_n5263__), .dout(new_new_n9953__));
  buf1  g9012(.din(new_new_n9953__), .dout(new_new_n9954__));
  buf1  g9013(.din(new_new_n5255__), .dout(new_new_n9955__));
  buf1  g9014(.din(new_new_n5266__), .dout(new_new_n9956__));
  buf1  g9015(.din(new_new_n9956__), .dout(new_new_n9957__));
  buf1  g9016(.din(new_new_n5265__), .dout(new_new_n9958__));
  buf1  g9017(.din(new_new_n9958__), .dout(new_new_n9959__));
  buf1  g9018(.din(new_new_n5274__), .dout(new_new_n9960__));
  buf1  g9019(.din(new_new_n5272__), .dout(new_new_n9961__));
  buf1  g9020(.din(new_new_n5273__), .dout(new_new_n9962__));
  buf1  g9021(.din(new_new_n5271__), .dout(new_new_n9963__));
  buf1  g9022(.din(new_new_n5276__), .dout(new_new_n9964__));
  buf1  g9023(.din(new_new_n9964__), .dout(new_new_n9965__));
  buf1  g9024(.din(new_new_n5275__), .dout(new_new_n9966__));
  buf1  g9025(.din(new_new_n9966__), .dout(new_new_n9967__));
  buf1  g9026(.din(new_new_n5294__), .dout(new_new_n9968__));
  buf1  g9027(.din(new_new_n5292__), .dout(new_new_n9969__));
  buf1  g9028(.din(new_new_n5293__), .dout(new_new_n9970__));
  buf1  g9029(.din(new_new_n5291__), .dout(new_new_n9971__));
  buf1  g9030(.din(new_new_n5296__), .dout(new_new_n9972__));
  buf1  g9031(.din(new_new_n9972__), .dout(new_new_n9973__));
  buf1  g9032(.din(new_new_n5295__), .dout(new_new_n9974__));
  buf1  g9033(.din(new_new_n5305__), .dout(new_new_n9975__));
  buf1  g9034(.din(new_new_n9975__), .dout(new_new_n9976__));
  buf1  g9035(.din(new_new_n5055__), .dout(new_new_n9977__));
  buf1  g9036(.din(new_new_n5321__), .dout(new_new_n9978__));
  buf1  g9037(.din(new_new_n5319__), .dout(new_new_n9979__));
  buf1  g9038(.din(new_new_n5320__), .dout(new_new_n9980__));
  buf1  g9039(.din(new_new_n5318__), .dout(new_new_n9981__));
  buf1  g9040(.din(new_new_n5323__), .dout(new_new_n9982__));
  buf1  g9041(.din(new_new_n9982__), .dout(new_new_n9983__));
  buf1  g9042(.din(new_new_n5322__), .dout(new_new_n9984__));
  buf1  g9043(.din(new_new_n9984__), .dout(new_new_n9985__));
  buf1  g9044(.din(new_new_n5331__), .dout(new_new_n9986__));
  buf1  g9045(.din(new_new_n5329__), .dout(new_new_n9987__));
  buf1  g9046(.din(new_new_n5330__), .dout(new_new_n9988__));
  buf1  g9047(.din(new_new_n5328__), .dout(new_new_n9989__));
  buf1  g9048(.din(new_new_n5333__), .dout(new_new_n9990__));
  buf1  g9049(.din(new_new_n9990__), .dout(new_new_n9991__));
  buf1  g9050(.din(new_new_n5332__), .dout(new_new_n9992__));
  buf1  g9051(.din(new_new_n9992__), .dout(new_new_n9993__));
  buf1  g9052(.din(new_new_n5335__), .dout(new_new_n9994__));
  buf1  g9053(.din(new_new_n5313__), .dout(new_new_n9995__));
  buf1  g9054(.din(new_new_n5334__), .dout(new_new_n9996__));
  buf1  g9055(.din(new_new_n5312__), .dout(new_new_n9997__));
  buf1  g9056(.din(new_new_n5337__), .dout(new_new_n9998__));
  buf1  g9057(.din(new_new_n9998__), .dout(new_new_n9999__));
  buf1  g9058(.din(new_new_n5336__), .dout(new_new_n10000__));
  buf1  g9059(.din(new_new_n10000__), .dout(new_new_n10001__));
  buf1  g9060(.din(new_new_n5345__), .dout(new_new_n10002__));
  buf1  g9061(.din(new_new_n5343__), .dout(new_new_n10003__));
  buf1  g9062(.din(new_new_n5344__), .dout(new_new_n10004__));
  buf1  g9063(.din(new_new_n5342__), .dout(new_new_n10005__));
  buf1  g9064(.din(new_new_n5347__), .dout(new_new_n10006__));
  buf1  g9065(.din(new_new_n10006__), .dout(new_new_n10007__));
  buf1  g9066(.din(new_new_n5346__), .dout(new_new_n10008__));
  buf1  g9067(.din(new_new_n10008__), .dout(new_new_n10009__));
  buf1  g9068(.din(new_new_n5361__), .dout(new_new_n10010__));
  buf1  g9069(.din(new_new_n5359__), .dout(new_new_n10011__));
  buf1  g9070(.din(new_new_n5360__), .dout(new_new_n10012__));
  buf1  g9071(.din(new_new_n5358__), .dout(new_new_n10013__));
  buf1  g9072(.din(new_new_n5363__), .dout(new_new_n10014__));
  buf1  g9073(.din(new_new_n10014__), .dout(new_new_n10015__));
  buf1  g9074(.din(new_new_n5362__), .dout(new_new_n10016__));
  buf1  g9075(.din(new_new_n10016__), .dout(new_new_n10017__));
  buf1  g9076(.din(new_new_n5371__), .dout(new_new_n10018__));
  buf1  g9077(.din(new_new_n5369__), .dout(new_new_n10019__));
  buf1  g9078(.din(new_new_n5370__), .dout(new_new_n10020__));
  buf1  g9079(.din(new_new_n5368__), .dout(new_new_n10021__));
  buf1  g9080(.din(new_new_n5373__), .dout(new_new_n10022__));
  buf1  g9081(.din(new_new_n10022__), .dout(new_new_n10023__));
  buf1  g9082(.din(new_new_n5372__), .dout(new_new_n10024__));
  buf1  g9083(.din(new_new_n10024__), .dout(new_new_n10025__));
  buf1  g9084(.din(new_new_n5375__), .dout(new_new_n10026__));
  buf1  g9085(.din(new_new_n5353__), .dout(new_new_n10027__));
  buf1  g9086(.din(new_new_n5374__), .dout(new_new_n10028__));
  buf1  g9087(.din(new_new_n5352__), .dout(new_new_n10029__));
  buf1  g9088(.din(new_new_n5377__), .dout(new_new_n10030__));
  buf1  g9089(.din(new_new_n10030__), .dout(new_new_n10031__));
  buf1  g9090(.din(new_new_n5376__), .dout(new_new_n10032__));
  buf1  g9091(.din(new_new_n5386__), .dout(new_new_n10033__));
  buf1  g9092(.din(new_new_n10033__), .dout(new_new_n10034__));
  buf1  g9093(.din(new_new_n4966__), .dout(new_new_n10035__));
  buf1  g9094(.din(new_new_n10035__), .dout(new_new_n10036__));
  buf1  g9095(.din(new_new_n4995__), .dout(new_new_n10037__));
  buf1  g9096(.din(new_new_n10037__), .dout(new_new_n10038__));
  buf1  g9097(.din(new_new_n5024__), .dout(new_new_n10039__));
  buf1  g9098(.din(new_new_n10039__), .dout(new_new_n10040__));
  buf1  g9099(.din(new_new_n5033__), .dout(new_new_n10041__));
  buf1  g9100(.din(new_new_n10041__), .dout(new_new_n10042__));
  buf1  g9101(.din(new_new_n5036__), .dout(new_new_n10043__));
  buf1  g9102(.din(new_new_n4936__), .dout(new_new_n10044__));
  buf1  g9103(.din(new_new_n5039__), .dout(new_new_n10045__));
  buf1  g9104(.din(new_new_n4937__), .dout(new_new_n10046__));
  buf1  g9105(.din(new_new_n5042__), .dout(new_new_n10047__));
  buf1  g9106(.din(new_new_n4938__), .dout(new_new_n10048__));
  buf1  g9107(.din(new_new_n5045__), .dout(new_new_n10049__));
  buf1  g9108(.din(new_new_n4939__), .dout(new_new_n10050__));
  buf1  g9109(.din(new_new_n4365__), .dout(new_new_n10051__));
  buf1  g9110(.din(new_new_n10051__), .dout(new_new_n10052__));
  buf1  g9111(.din(new_new_n4364__), .dout(new_new_n10053__));
  buf1  g9112(.din(new_new_n847__), .dout(new_new_n10054__));
  buf1  g9113(.din(new_new_n10054__), .dout(new_new_n10055__));
  buf1  g9114(.din(new_new_n10055__), .dout(new_new_n10056__));
  buf1  g9115(.din(new_new_n10055__), .dout(new_new_n10057__));
  buf1  g9116(.din(new_new_n10054__), .dout(new_new_n10058__));
  buf1  g9117(.din(new_new_n10058__), .dout(new_new_n10059__));
  buf1  g9118(.din(new_new_n848__), .dout(new_new_n10060__));
  buf1  g9119(.din(new_new_n10060__), .dout(new_new_n10061__));
  buf1  g9120(.din(new_new_n10061__), .dout(new_new_n10062__));
  buf1  g9121(.din(new_new_n10061__), .dout(new_new_n10063__));
  buf1  g9122(.din(new_new_n10060__), .dout(new_new_n10064__));
  buf1  g9123(.din(new_new_n5414__), .dout(new_new_n10065__));
  buf1  g9124(.din(new_new_n5412__), .dout(new_new_n10066__));
  buf1  g9125(.din(new_new_n5413__), .dout(new_new_n10067__));
  buf1  g9126(.din(new_new_n5411__), .dout(new_new_n10068__));
  buf1  g9127(.din(new_new_n5416__), .dout(new_new_n10069__));
  buf1  g9128(.din(new_new_n10069__), .dout(new_new_n10070__));
  buf1  g9129(.din(new_new_n5415__), .dout(new_new_n10071__));
  buf1  g9130(.din(new_new_n5424__), .dout(new_new_n10072__));
  buf1  g9131(.din(new_new_n5422__), .dout(new_new_n10073__));
  buf1  g9132(.din(new_new_n5423__), .dout(new_new_n10074__));
  buf1  g9133(.din(new_new_n5421__), .dout(new_new_n10075__));
  buf1  g9134(.din(new_new_n5426__), .dout(new_new_n10076__));
  buf1  g9135(.din(new_new_n10076__), .dout(new_new_n10077__));
  buf1  g9136(.din(new_new_n5425__), .dout(new_new_n10078__));
  buf1  g9137(.din(new_new_n5443__), .dout(new_new_n10079__));
  buf1  g9138(.din(new_new_n5441__), .dout(new_new_n10080__));
  buf1  g9139(.din(new_new_n5442__), .dout(new_new_n10081__));
  buf1  g9140(.din(new_new_n5440__), .dout(new_new_n10082__));
  buf1  g9141(.din(new_new_n5445__), .dout(new_new_n10083__));
  buf1  g9142(.din(new_new_n10083__), .dout(new_new_n10084__));
  buf1  g9143(.din(new_new_n5444__), .dout(new_new_n10085__));
  buf1  g9144(.din(new_new_n5453__), .dout(new_new_n10086__));
  buf1  g9145(.din(new_new_n5451__), .dout(new_new_n10087__));
  buf1  g9146(.din(new_new_n5452__), .dout(new_new_n10088__));
  buf1  g9147(.din(new_new_n5450__), .dout(new_new_n10089__));
  buf1  g9148(.din(new_new_n5455__), .dout(new_new_n10090__));
  buf1  g9149(.din(new_new_n10090__), .dout(new_new_n10091__));
  buf1  g9150(.din(new_new_n5454__), .dout(new_new_n10092__));
  buf1  g9151(.din(new_new_n5478__), .dout(new_new_n10093__));
  buf1  g9152(.din(new_new_n5476__), .dout(new_new_n10094__));
  buf1  g9153(.din(new_new_n5477__), .dout(new_new_n10095__));
  buf1  g9154(.din(new_new_n5475__), .dout(new_new_n10096__));
  buf1  g9155(.din(new_new_n5480__), .dout(new_new_n10097__));
  buf1  g9156(.din(new_new_n10097__), .dout(new_new_n10098__));
  buf1  g9157(.din(new_new_n5479__), .dout(new_new_n10099__));
  buf1  g9158(.din(new_new_n10099__), .dout(new_new_n10100__));
  buf1  g9159(.din(new_new_n5488__), .dout(new_new_n10101__));
  buf1  g9160(.din(new_new_n5486__), .dout(new_new_n10102__));
  buf1  g9161(.din(new_new_n5490__), .dout(new_new_n10103__));
  buf1  g9162(.din(new_new_n10103__), .dout(new_new_n10104__));
  buf1  g9163(.din(new_new_n5507__), .dout(new_new_n10105__));
  buf1  g9164(.din(new_new_n5505__), .dout(new_new_n10106__));
  buf1  g9165(.din(new_new_n5506__), .dout(new_new_n10107__));
  buf1  g9166(.din(new_new_n5504__), .dout(new_new_n10108__));
  buf1  g9167(.din(new_new_n5509__), .dout(new_new_n10109__));
  buf1  g9168(.din(new_new_n10109__), .dout(new_new_n10110__));
  buf1  g9169(.din(new_new_n5508__), .dout(new_new_n10111__));
  buf1  g9170(.din(new_new_n10111__), .dout(new_new_n10112__));
  buf1  g9171(.din(new_new_n5516__), .dout(new_new_n10113__));
  buf1  g9172(.din(new_new_n5514__), .dout(new_new_n10114__));
  buf1  g9173(.din(new_new_n5518__), .dout(new_new_n10115__));
  buf1  g9174(.din(new_new_n10115__), .dout(new_new_n10116__));
  buf1  g9175(.din(new_new_n4289__), .dout(new_new_n10117__));
  buf1  g9176(.din(new_new_n10117__), .dout(new_new_n10118__));
  buf1  g9177(.din(new_new_n4298__), .dout(new_new_n10119__));
  buf1  g9178(.din(new_new_n10119__), .dout(new_new_n10120__));
  buf1  g9179(.din(new_new_n4307__), .dout(new_new_n10121__));
  buf1  g9180(.din(new_new_n10121__), .dout(new_new_n10122__));
  buf1  g9181(.din(new_new_n4336__), .dout(new_new_n10123__));
  buf1  g9182(.din(new_new_n10123__), .dout(new_new_n10124__));
  buf1  g9183(.din(new_new_n5213__), .dout(new_new_n10125__));
  buf1  g9184(.din(new_new_n815__), .dout(new_new_n10126__));
  buf1  g9185(.din(new_new_n10126__), .dout(new_new_n10127__));
  buf1  g9186(.din(new_new_n10126__), .dout(new_new_n10128__));
  buf1  g9187(.din(new_new_n816__), .dout(new_new_n10129__));
  buf1  g9188(.din(new_new_n5542__), .dout(new_new_n10130__));
  buf1  g9189(.din(new_new_n5539__), .dout(new_new_n10131__));
  buf1  g9190(.din(new_new_n5541__), .dout(new_new_n10132__));
  buf1  g9191(.din(new_new_n5540__), .dout(new_new_n10133__));
  buf1  g9192(.din(new_new_n5544__), .dout(new_new_n10134__));
  buf1  g9193(.din(new_new_n5543__), .dout(new_new_n10135__));
  buf1  g9194(.din(new_new_n5545__), .dout(new_new_n10136__));
  buf1  g9195(.din(new_new_n825__), .dout(new_new_n10137__));
  buf1  g9196(.din(new_new_n10137__), .dout(new_new_n10138__));
  buf1  g9197(.din(new_new_n10138__), .dout(new_new_n10139__));
  buf1  g9198(.din(new_new_n10137__), .dout(new_new_n10140__));
  buf1  g9199(.din(new_new_n826__), .dout(new_new_n10141__));
  buf1  g9200(.din(new_new_n10141__), .dout(new_new_n10142__));
  buf1  g9201(.din(new_new_n5561__), .dout(new_new_n10143__));
  buf1  g9202(.din(new_new_n5558__), .dout(new_new_n10144__));
  buf1  g9203(.din(new_new_n5560__), .dout(new_new_n10145__));
  buf1  g9204(.din(new_new_n5559__), .dout(new_new_n10146__));
  buf1  g9205(.din(new_new_n5563__), .dout(new_new_n10147__));
  buf1  g9206(.din(new_new_n5562__), .dout(new_new_n10148__));
  buf1  g9207(.din(new_new_n5565__), .dout(new_new_n10149__));
  buf1  g9208(.din(new_new_n10149__), .dout(new_new_n10150__));
  buf1  g9209(.din(new_new_n5557__), .dout(new_new_n10151__));
  buf1  g9210(.din(new_new_n5564__), .dout(new_new_n10152__));
  buf1  g9211(.din(new_new_n10152__), .dout(new_new_n10153__));
  buf1  g9212(.din(new_new_n5556__), .dout(new_new_n10154__));
  buf1  g9213(.din(new_new_n5567__), .dout(new_new_n10155__));
  buf1  g9214(.din(new_new_n10155__), .dout(new_new_n10156__));
  buf1  g9215(.din(new_new_n5566__), .dout(new_new_n10157__));
  buf1  g9216(.din(new_new_n10157__), .dout(new_new_n10158__));
  buf1  g9217(.din(new_new_n5575__), .dout(new_new_n10159__));
  buf1  g9218(.din(new_new_n5573__), .dout(new_new_n10160__));
  buf1  g9219(.din(new_new_n5574__), .dout(new_new_n10161__));
  buf1  g9220(.din(new_new_n5572__), .dout(new_new_n10162__));
  buf1  g9221(.din(new_new_n5577__), .dout(new_new_n10163__));
  buf1  g9222(.din(new_new_n10163__), .dout(new_new_n10164__));
  buf1  g9223(.din(new_new_n5576__), .dout(new_new_n10165__));
  buf1  g9224(.din(new_new_n10165__), .dout(new_new_n10166__));
  buf1  g9225(.din(new_new_n4410__), .dout(new_new_n10167__));
  buf1  g9226(.din(new_new_n10167__), .dout(new_new_n10168__));
  buf1  g9227(.din(new_new_n4663__), .dout(new_new_n10169__));
  buf1  g9228(.din(new_new_n10169__), .dout(new_new_n10170__));
  buf1  g9229(.din(new_new_n4882__), .dout(new_new_n10171__));
  buf1  g9230(.din(new_new_n10171__), .dout(new_new_n10172__));
  buf1  g9231(.din(new_new_n811__), .dout(new_new_n10173__));
  buf1  g9232(.din(new_new_n10173__), .dout(new_new_n10174__));
  buf1  g9233(.din(new_new_n812__), .dout(new_new_n10175__));
  buf1  g9234(.din(new_new_n901__), .dout(new_new_n10176__));
  buf1  g9235(.din(new_new_n5612__), .dout(new_new_n10177__));
  buf1  g9236(.din(new_new_n5610__), .dout(new_new_n10178__));
  buf1  g9237(.din(new_new_n5611__), .dout(new_new_n10179__));
  buf1  g9238(.din(new_new_n5609__), .dout(new_new_n10180__));
  buf1  g9239(.din(new_new_n5614__), .dout(new_new_n10181__));
  buf1  g9240(.din(new_new_n10181__), .dout(new_new_n10182__));
  buf1  g9241(.din(new_new_n5613__), .dout(new_new_n10183__));
  buf1  g9242(.din(new_new_n5623__), .dout(new_new_n10184__));
  buf1  g9243(.din(new_new_n10184__), .dout(new_new_n10185__));
  buf1  g9244(.din(new_new_n813__), .dout(new_new_n10186__));
  buf1  g9245(.din(new_new_n10186__), .dout(new_new_n10187__));
  buf1  g9246(.din(new_new_n814__), .dout(new_new_n10188__));
  buf1  g9247(.din(new_new_n5629__), .dout(new_new_n10189__));
  buf1  g9248(.din(new_new_n823__), .dout(new_new_n10190__));
  buf1  g9249(.din(new_new_n10190__), .dout(new_new_n10191__));
  buf1  g9250(.din(new_new_n10190__), .dout(new_new_n10192__));
  buf1  g9251(.din(new_new_n824__), .dout(new_new_n10193__));
  buf1  g9252(.din(new_new_n10193__), .dout(new_new_n10194__));
  buf1  g9253(.din(new_new_n5634__), .dout(new_new_n10195__));
  buf1  g9254(.din(new_new_n5631__), .dout(new_new_n10196__));
  buf1  g9255(.din(new_new_n5633__), .dout(new_new_n10197__));
  buf1  g9256(.din(new_new_n5632__), .dout(new_new_n10198__));
  buf1  g9257(.din(new_new_n5636__), .dout(new_new_n10199__));
  buf1  g9258(.din(new_new_n5635__), .dout(new_new_n10200__));
  buf1  g9259(.din(new_new_n5638__), .dout(new_new_n10201__));
  buf1  g9260(.din(new_new_n10201__), .dout(new_new_n10202__));
  buf1  g9261(.din(new_new_n5637__), .dout(new_new_n10203__));
  buf1  g9262(.din(new_new_n10203__), .dout(new_new_n10204__));
  buf1  g9263(.din(new_new_n5646__), .dout(new_new_n10205__));
  buf1  g9264(.din(new_new_n5643__), .dout(new_new_n10206__));
  buf1  g9265(.din(new_new_n5645__), .dout(new_new_n10207__));
  buf1  g9266(.din(new_new_n5644__), .dout(new_new_n10208__));
  buf1  g9267(.din(new_new_n5648__), .dout(new_new_n10209__));
  buf1  g9268(.din(new_new_n5647__), .dout(new_new_n10210__));
  buf1  g9269(.din(new_new_n5650__), .dout(new_new_n10211__));
  buf1  g9270(.din(new_new_n10211__), .dout(new_new_n10212__));
  buf1  g9271(.din(new_new_n5642__), .dout(new_new_n10213__));
  buf1  g9272(.din(new_new_n5649__), .dout(new_new_n10214__));
  buf1  g9273(.din(new_new_n10214__), .dout(new_new_n10215__));
  buf1  g9274(.din(new_new_n5641__), .dout(new_new_n10216__));
  buf1  g9275(.din(new_new_n5652__), .dout(new_new_n10217__));
  buf1  g9276(.din(new_new_n10217__), .dout(new_new_n10218__));
  buf1  g9277(.din(new_new_n5651__), .dout(new_new_n10219__));
  buf1  g9278(.din(new_new_n5661__), .dout(new_new_n10220__));
  buf1  g9279(.din(new_new_n10220__), .dout(new_new_n10221__));
  buf1  g9280(.din(new_new_n835__), .dout(new_new_n10222__));
  buf1  g9281(.din(new_new_n10222__), .dout(new_new_n10223__));
  buf1  g9282(.din(new_new_n10223__), .dout(new_new_n10224__));
  buf1  g9283(.din(new_new_n10222__), .dout(new_new_n10225__));
  buf1  g9284(.din(new_new_n836__), .dout(new_new_n10226__));
  buf1  g9285(.din(new_new_n10226__), .dout(new_new_n10227__));
  buf1  g9286(.din(new_new_n10226__), .dout(new_new_n10228__));
  buf1  g9287(.din(new_new_n5666__), .dout(new_new_n10229__));
  buf1  g9288(.din(new_new_n5663__), .dout(new_new_n10230__));
  buf1  g9289(.din(new_new_n5665__), .dout(new_new_n10231__));
  buf1  g9290(.din(new_new_n5664__), .dout(new_new_n10232__));
  buf1  g9291(.din(new_new_n5668__), .dout(new_new_n10233__));
  buf1  g9292(.din(new_new_n5667__), .dout(new_new_n10234__));
  buf1  g9293(.din(new_new_n5670__), .dout(new_new_n10235__));
  buf1  g9294(.din(new_new_n10235__), .dout(new_new_n10236__));
  buf1  g9295(.din(new_new_n5669__), .dout(new_new_n10237__));
  buf1  g9296(.din(new_new_n10237__), .dout(new_new_n10238__));
  buf1  g9297(.din(new_new_n5678__), .dout(new_new_n10239__));
  buf1  g9298(.din(new_new_n5675__), .dout(new_new_n10240__));
  buf1  g9299(.din(new_new_n5677__), .dout(new_new_n10241__));
  buf1  g9300(.din(new_new_n5676__), .dout(new_new_n10242__));
  buf1  g9301(.din(new_new_n5680__), .dout(new_new_n10243__));
  buf1  g9302(.din(new_new_n5679__), .dout(new_new_n10244__));
  buf1  g9303(.din(new_new_n5682__), .dout(new_new_n10245__));
  buf1  g9304(.din(new_new_n10245__), .dout(new_new_n10246__));
  buf1  g9305(.din(new_new_n5674__), .dout(new_new_n10247__));
  buf1  g9306(.din(new_new_n5681__), .dout(new_new_n10248__));
  buf1  g9307(.din(new_new_n10248__), .dout(new_new_n10249__));
  buf1  g9308(.din(new_new_n5673__), .dout(new_new_n10250__));
  buf1  g9309(.din(new_new_n5684__), .dout(new_new_n10251__));
  buf1  g9310(.din(new_new_n10251__), .dout(new_new_n10252__));
  buf1  g9311(.din(new_new_n5683__), .dout(new_new_n10253__));
  buf1  g9312(.din(new_new_n10253__), .dout(new_new_n10254__));
  buf1  g9313(.din(new_new_n5692__), .dout(new_new_n10255__));
  buf1  g9314(.din(new_new_n5690__), .dout(new_new_n10256__));
  buf1  g9315(.din(new_new_n5691__), .dout(new_new_n10257__));
  buf1  g9316(.din(new_new_n5689__), .dout(new_new_n10258__));
  buf1  g9317(.din(new_new_n5694__), .dout(new_new_n10259__));
  buf1  g9318(.din(new_new_n10259__), .dout(new_new_n10260__));
  buf1  g9319(.din(new_new_n5693__), .dout(new_new_n10261__));
  buf1  g9320(.din(new_new_n10261__), .dout(new_new_n10262__));
  buf1  g9321(.din(new_new_n5704__), .dout(new_new_n10263__));
  buf1  g9322(.din(new_new_n5703__), .dout(new_new_n10264__));
  buf1  g9323(.din(new_new_n5706__), .dout(new_new_n10265__));
  buf1  g9324(.din(new_new_n10265__), .dout(new_new_n10266__));
  buf1  g9325(.din(new_new_n5705__), .dout(new_new_n10267__));
  buf1  g9326(.din(new_new_n10267__), .dout(new_new_n10268__));
  buf1  g9327(.din(new_new_n5714__), .dout(new_new_n10269__));
  buf1  g9328(.din(new_new_n5712__), .dout(new_new_n10270__));
  buf1  g9329(.din(new_new_n5713__), .dout(new_new_n10271__));
  buf1  g9330(.din(new_new_n5711__), .dout(new_new_n10272__));
  buf1  g9331(.din(new_new_n5716__), .dout(new_new_n10273__));
  buf1  g9332(.din(new_new_n10273__), .dout(new_new_n10274__));
  buf1  g9333(.din(new_new_n5715__), .dout(new_new_n10275__));
  buf1  g9334(.din(new_new_n10275__), .dout(new_new_n10276__));
  buf1  g9335(.din(new_new_n5718__), .dout(new_new_n10277__));
  buf1  g9336(.din(new_new_n5700__), .dout(new_new_n10278__));
  buf1  g9337(.din(new_new_n5717__), .dout(new_new_n10279__));
  buf1  g9338(.din(new_new_n5699__), .dout(new_new_n10280__));
  buf1  g9339(.din(new_new_n5720__), .dout(new_new_n10281__));
  buf1  g9340(.din(new_new_n10281__), .dout(new_new_n10282__));
  buf1  g9341(.din(new_new_n5719__), .dout(new_new_n10283__));
  buf1  g9342(.din(new_new_n5729__), .dout(new_new_n10284__));
  buf1  g9343(.din(new_new_n10284__), .dout(new_new_n10285__));
  buf1  g9344(.din(new_new_n5435__), .dout(new_new_n10286__));
  buf1  g9345(.din(new_new_n10286__), .dout(new_new_n10287__));
  buf1  g9346(.din(new_new_n5464__), .dout(new_new_n10288__));
  buf1  g9347(.din(new_new_n10288__), .dout(new_new_n10289__));
  buf1  g9348(.din(new_new_n5493__), .dout(new_new_n10290__));
  buf1  g9349(.din(new_new_n10290__), .dout(new_new_n10291__));
  buf1  g9350(.din(new_new_n5522__), .dout(new_new_n10292__));
  buf1  g9351(.din(new_new_n10292__), .dout(new_new_n10293__));
  buf1  g9352(.din(new_new_n5589__), .dout(new_new_n10294__));
  buf1  g9353(.din(new_new_n5281__), .dout(new_new_n10295__));
  buf1  g9354(.din(new_new_n5595__), .dout(new_new_n10296__));
  buf1  g9355(.din(new_new_n5282__), .dout(new_new_n10297__));
  buf1  g9356(.din(new_new_n5592__), .dout(new_new_n10298__));
  buf1  g9357(.din(new_new_n5283__), .dout(new_new_n10299__));
  buf1  g9358(.din(new_new_n5596__), .dout(new_new_n10300__));
  buf1  g9359(.din(new_new_n5284__), .dout(new_new_n10301__));
  buf1  g9360(.din(new_new_n5586__), .dout(new_new_n10302__));
  buf1  g9361(.din(new_new_n5307__), .dout(new_new_n10303__));
  buf1  g9362(.din(new_new_n5583__), .dout(new_new_n10304__));
  buf1  g9363(.din(new_new_n5387__), .dout(new_new_n10305__));
  buf1  g9364(.din(new_new_n5546__), .dout(new_new_n10306__));
  buf1  g9365(.din(new_new_n5754__), .dout(new_new_n10307__));
  buf1  g9366(.din(new_new_n5751__), .dout(new_new_n10308__));
  buf1  g9367(.din(new_new_n5752__), .dout(new_new_n10309__));
  buf1  g9368(.din(new_new_n5756__), .dout(new_new_n10310__));
  buf1  g9369(.din(new_new_n5757__), .dout(new_new_n10311__));
  buf1  g9370(.din(new_new_n5769__), .dout(new_new_n10312__));
  buf1  g9371(.din(new_new_n5768__), .dout(new_new_n10313__));
  buf1  g9372(.din(new_new_n5771__), .dout(new_new_n10314__));
  buf1  g9373(.din(new_new_n10314__), .dout(new_new_n10315__));
  buf1  g9374(.din(new_new_n5770__), .dout(new_new_n10316__));
  buf1  g9375(.din(new_new_n10316__), .dout(new_new_n10317__));
  buf1  g9376(.din(new_new_n5778__), .dout(new_new_n10318__));
  buf1  g9377(.din(new_new_n5776__), .dout(new_new_n10319__));
  buf1  g9378(.din(new_new_n5780__), .dout(new_new_n10320__));
  buf1  g9379(.din(new_new_n10320__), .dout(new_new_n10321__));
  buf1  g9380(.din(new_new_n5794__), .dout(new_new_n10322__));
  buf1  g9381(.din(new_new_n5793__), .dout(new_new_n10323__));
  buf1  g9382(.din(new_new_n5796__), .dout(new_new_n10324__));
  buf1  g9383(.din(new_new_n10324__), .dout(new_new_n10325__));
  buf1  g9384(.din(new_new_n5795__), .dout(new_new_n10326__));
  buf1  g9385(.din(new_new_n10326__), .dout(new_new_n10327__));
  buf1  g9386(.din(new_new_n5804__), .dout(new_new_n10328__));
  buf1  g9387(.din(new_new_n5802__), .dout(new_new_n10329__));
  buf1  g9388(.din(new_new_n5803__), .dout(new_new_n10330__));
  buf1  g9389(.din(new_new_n5801__), .dout(new_new_n10331__));
  buf1  g9390(.din(new_new_n5806__), .dout(new_new_n10332__));
  buf1  g9391(.din(new_new_n10332__), .dout(new_new_n10333__));
  buf1  g9392(.din(new_new_n5805__), .dout(new_new_n10334__));
  buf1  g9393(.din(new_new_n10334__), .dout(new_new_n10335__));
  buf1  g9394(.din(new_new_n5808__), .dout(new_new_n10336__));
  buf1  g9395(.din(new_new_n5790__), .dout(new_new_n10337__));
  buf1  g9396(.din(new_new_n5807__), .dout(new_new_n10338__));
  buf1  g9397(.din(new_new_n5789__), .dout(new_new_n10339__));
  buf1  g9398(.din(new_new_n5810__), .dout(new_new_n10340__));
  buf1  g9399(.din(new_new_n10340__), .dout(new_new_n10341__));
  buf1  g9400(.din(new_new_n5809__), .dout(new_new_n10342__));
  buf1  g9401(.din(new_new_n5818__), .dout(new_new_n10343__));
  buf1  g9402(.din(new_new_n5816__), .dout(new_new_n10344__));
  buf1  g9403(.din(new_new_n5817__), .dout(new_new_n10345__));
  buf1  g9404(.din(new_new_n5815__), .dout(new_new_n10346__));
  buf1  g9405(.din(new_new_n5820__), .dout(new_new_n10347__));
  buf1  g9406(.din(new_new_n10347__), .dout(new_new_n10348__));
  buf1  g9407(.din(new_new_n5819__), .dout(new_new_n10349__));
  buf1  g9408(.din(new_new_n5834__), .dout(new_new_n10350__));
  buf1  g9409(.din(new_new_n5832__), .dout(new_new_n10351__));
  buf1  g9410(.din(new_new_n5833__), .dout(new_new_n10352__));
  buf1  g9411(.din(new_new_n5831__), .dout(new_new_n10353__));
  buf1  g9412(.din(new_new_n5836__), .dout(new_new_n10354__));
  buf1  g9413(.din(new_new_n10354__), .dout(new_new_n10355__));
  buf1  g9414(.din(new_new_n5835__), .dout(new_new_n10356__));
  buf1  g9415(.din(new_new_n10356__), .dout(new_new_n10357__));
  buf1  g9416(.din(new_new_n5843__), .dout(new_new_n10358__));
  buf1  g9417(.din(new_new_n5841__), .dout(new_new_n10359__));
  buf1  g9418(.din(new_new_n5845__), .dout(new_new_n10360__));
  buf1  g9419(.din(new_new_n10360__), .dout(new_new_n10361__));
  buf1  g9420(.din(new_new_n5054__), .dout(new_new_n10362__));
  buf1  g9421(.din(new_new_n10362__), .dout(new_new_n10363__));
  buf1  g9422(.din(new_new_n5104__), .dout(new_new_n10364__));
  buf1  g9423(.din(new_new_n10364__), .dout(new_new_n10365__));
  buf1  g9424(.din(new_new_n5193__), .dout(new_new_n10366__));
  buf1  g9425(.din(new_new_n10366__), .dout(new_new_n10367__));
  buf1  g9426(.din(new_new_n5214__), .dout(new_new_n10368__));
  buf1  g9427(.din(new_new_n10368__), .dout(new_new_n10369__));
  buf1  g9428(.din(new_new_n5279__), .dout(new_new_n10370__));
  buf1  g9429(.din(new_new_n10370__), .dout(new_new_n10371__));
  buf1  g9430(.din(new_new_n5744__), .dout(new_new_n10372__));
  buf1  g9431(.din(new_new_n5883__), .dout(new_new_n10373__));
  buf1  g9432(.din(new_new_n5882__), .dout(new_new_n10374__));
  buf1  g9433(.din(new_new_n5885__), .dout(new_new_n10375__));
  buf1  g9434(.din(new_new_n10375__), .dout(new_new_n10376__));
  buf1  g9435(.din(new_new_n5884__), .dout(new_new_n10377__));
  buf1  g9436(.din(new_new_n5894__), .dout(new_new_n10378__));
  buf1  g9437(.din(new_new_n10378__), .dout(new_new_n10379__));
  buf1  g9438(.din(new_new_n5903__), .dout(new_new_n10380__));
  buf1  g9439(.din(new_new_n5901__), .dout(new_new_n10381__));
  buf1  g9440(.din(new_new_n5902__), .dout(new_new_n10382__));
  buf1  g9441(.din(new_new_n5900__), .dout(new_new_n10383__));
  buf1  g9442(.din(new_new_n5905__), .dout(new_new_n10384__));
  buf1  g9443(.din(new_new_n10384__), .dout(new_new_n10385__));
  buf1  g9444(.din(new_new_n5904__), .dout(new_new_n10386__));
  buf1  g9445(.din(new_new_n5914__), .dout(new_new_n10387__));
  buf1  g9446(.din(new_new_n10387__), .dout(new_new_n10388__));
  buf1  g9447(.din(new_new_n5759__), .dout(new_new_n10389__));
  buf1  g9448(.din(new_new_n10389__), .dout(new_new_n10390__));
  buf1  g9449(.din(new_new_n5784__), .dout(new_new_n10391__));
  buf1  g9450(.din(new_new_n10391__), .dout(new_new_n10392__));
  buf1  g9451(.din(new_new_n5849__), .dout(new_new_n10393__));
  buf1  g9452(.din(new_new_n10393__), .dout(new_new_n10394__));
  buf1  g9453(.din(new_new_n5875__), .dout(new_new_n10395__));
  buf1  g9454(.din(new_new_n5601__), .dout(new_new_n10396__));
  buf1  g9455(.din(new_new_n5872__), .dout(new_new_n10397__));
  buf1  g9456(.din(new_new_n5602__), .dout(new_new_n10398__));
  buf1  g9457(.din(new_new_n5866__), .dout(new_new_n10399__));
  buf1  g9458(.din(new_new_n5630__), .dout(new_new_n10400__));
  buf1  g9459(.din(new_new_n10400__), .dout(new_new_n10401__));
  buf1  g9460(.din(new_new_n5869__), .dout(new_new_n10402__));
  buf1  g9461(.din(new_new_n5662__), .dout(new_new_n10403__));
  buf1  g9462(.din(new_new_n5864__), .dout(new_new_n10404__));
  buf1  g9463(.din(new_new_n5730__), .dout(new_new_n10405__));
  buf1  g9464(.din(new_new_n5410__), .dout(new_new_n10406__));
  buf1  g9465(.din(new_new_n10406__), .dout(new_new_n10407__));
  buf1  g9466(.din(new_new_n5547__), .dout(new_new_n10408__));
  buf1  g9467(.din(new_new_n10408__), .dout(new_new_n10409__));
  buf1  g9468(.din(new_new_n5580__), .dout(new_new_n10410__));
  buf1  g9469(.din(new_new_n10410__), .dout(new_new_n10411__));
  always @ (posedge clock) begin
    n2491_lo <= n19409;
    n2575_lo <= n19412;
    n2587_lo <= n19415;
    n2599_lo <= n19418;
    n2611_lo <= n19421;
    n2623_lo <= n19424;
    n2635_lo <= n19427;
    n2647_lo <= n19430;
    n2659_lo <= n19433;
    n2671_lo <= n19436;
    n2683_lo <= n19439;
    n2734_lo <= n19442;
    n2746_lo <= n19445;
    n2758_lo <= n19448;
    n2770_lo <= n19451;
    n2782_lo <= n19454;
    n2785_lo <= n19457;
    n2794_lo <= n19460;
    n2797_lo <= n19463;
    n2806_lo <= n19466;
    n2809_lo <= n19469;
    n2818_lo <= n19472;
    n2821_lo <= n19475;
    n2830_lo <= n19478;
    n2833_lo <= n19481;
    n2836_lo <= n19484;
    n2839_lo <= n19487;
    n2842_lo <= n19490;
    n2845_lo <= n19493;
    n2848_lo <= n19496;
    n2851_lo <= n19499;
    n2854_lo <= n19502;
    n2857_lo <= n19505;
    n2860_lo <= n19508;
    n2863_lo <= n19511;
    n4871_o2 <= n19514;
    n4893_o2 <= n19517;
    n4938_o2 <= n19520;
    n5056_o2 <= n19523;
    n5100_o2 <= n19526;
    n5122_o2 <= n19529;
    n5254_o2 <= n19532;
    n5276_o2 <= n19535;
    n5316_o2 <= n19538;
    n5434_o2 <= n19541;
    n5473_o2 <= n19544;
    n5494_o2 <= n19547;
    n5620_o2 <= n19550;
    n5643_o2 <= n19553;
    n5682_o2 <= n19556;
    n5798_o2 <= n19559;
    n5839_o2 <= n19562;
    n5867_o2 <= n19565;
    n6052_o2 <= n19568;
    n6087_o2 <= n19571;
    n6153_o2 <= n19574;
    n6408_o2 <= n19577;
    n6454_o2 <= n19580;
    n6509_o2 <= n19583;
    n6775_o2 <= n19586;
    n6818_o2 <= n19589;
    n6892_o2 <= n19592;
    n5779_o2 <= n19595;
    n5780_o2 <= n19598;
    n7156_o2 <= n19601;
    n5792_o2 <= n19604;
    n7205_o2 <= n19607;
    n5842_o2 <= n19610;
    n5863_o2 <= n19613;
    n7263_o2 <= n19616;
    n5881_o2 <= n19619;
    n5930_o2 <= n19622;
    n5959_o2 <= n19625;
    n5981_o2 <= n19628;
    n6042_o2 <= n19631;
    n6075_o2 <= n19634;
    n6103_o2 <= n19637;
    n7610_o2 <= n19640;
    n6169_o2 <= n19643;
    n7665_o2 <= n19646;
    n6205_o2 <= n19649;
    n6239_o2 <= n19652;
    n7788_o2 <= n19655;
    n6309_o2 <= n19658;
    n6461_o2 <= n19661;
    n6476_o2 <= n19664;
    n325_inv <= n19667;
    n6545_o2 <= n19670;
    G578_o2 <= n19673;
    G5106_o2 <= n19676;
    n6713_o2 <= n19679;
    G5164_o2 <= n19682;
    n343_inv <= n19685;
    n6810_o2 <= n19688;
    n6973_o2 <= n19691;
    n352_inv <= n19694;
    n7053_o2 <= n19697;
    G581_o2 <= n19700;
    G5467_o2 <= n19703;
    n7231_o2 <= n19706;
    G5527_o2 <= n19709;
    n370_inv <= n19712;
    n7304_o2 <= n19715;
    n7530_o2 <= n19718;
    n379_inv <= n19721;
    n7653_o2 <= n19724;
    G584_o2 <= n19727;
    G5820_o2 <= n19730;
    n7148_o2 <= n19733;
    n7149_o2 <= n19736;
    n7224_o2 <= n19739;
    n7916_o2 <= n19742;
    G5868_o2 <= n19745;
    n406_inv <= n19748;
    n7280_o2 <= n19751;
    n7313_o2 <= n19754;
    n8056_o2 <= n19757;
    n7323_o2 <= n19760;
    n7398_o2 <= n19763;
    n7459_o2 <= n19766;
    n7501_o2 <= n19769;
    n7518_o2 <= n19772;
    G563_o2 <= n19775;
    n7606_o2 <= n19778;
    n439_inv <= n19781;
    n7675_o2 <= n19784;
    G3410_o2 <= n19787;
    n7722_o2 <= n19790;
    n7747_o2 <= n19793;
    n7835_o2 <= n19796;
    G587_o2 <= n19799;
    G6046_o2 <= n19802;
    n7909_o2 <= n19805;
    G566_o2 <= n19808;
    G6070_o2 <= n19811;
    n472_inv <= n19814;
    n8086_o2 <= n19817;
    n8093_o2 <= n19820;
    G3752_o2 <= n19823;
    n484_inv <= n19826;
    n8199_o2 <= n19829;
    n2800_lo_buf_o2 <= n19832;
    G548_o2 <= n19835;
    n496_inv <= n19838;
    G569_o2 <= n19841;
    G1761_o2 <= n19844;
    n505_inv <= n19847;
    G4101_o2 <= n19850;
    G551_o2 <= n19853;
    n514_inv <= n19856;
    G4743_o2 <= n19859;
    G5271_o2 <= n19862;
    G5790_o2 <= n19865;
    G6122_o2 <= n19868;
    G2082_o2 <= n19871;
    n2812_lo_buf_o2 <= n19874;
    n2668_lo_buf_o2 <= n19877;
    n2680_lo_buf_o2 <= n19880;
    G572_o2 <= n19883;
    G6125_o2 <= n19886;
    n547_inv <= n19889;
    n2656_lo_buf_o2 <= n19892;
    G554_o2 <= n19895;
    G4452_o2 <= n19898;
    n559_inv <= n19901;
    n2644_lo_buf_o2 <= n19904;
    G2410_o2 <= n19907;
    n2632_lo_buf_o2 <= n19910;
    n2620_lo_buf_o2 <= n19913;
    G6131_o2 <= n19916;
    G4693_o2 <= n19919;
    G5209_o2 <= n19922;
    G5741_o2 <= n19925;
    G6082_o2 <= n19928;
    G6119_o2 <= n19931;
    n2608_lo_buf_o2 <= n19934;
    n2596_lo_buf_o2 <= n19937;
    n2584_lo_buf_o2 <= n19940;
    n2572_lo_buf_o2 <= n19943;
    n2704_lo_buf_o2 <= n19946;
    G557_o2 <= n19949;
    G5936_o2 <= n19952;
    G5442_o2 <= n19955;
    G4926_o2 <= n19958;
    G6134_o2 <= n19961;
    G3929_o2 <= n19964;
    G4425_o2 <= n19967;
    G4947_o2 <= n19970;
    n2764_lo_buf_o2 <= n19973;
    n634_inv <= n19976;
    n2560_lo_buf_o2 <= n19979;
    n2824_lo_buf_o2 <= n19982;
    G575_o2 <= n19985;
    G2740_o2 <= n19988;
    n649_inv <= n19991;
    n2548_lo_buf_o2 <= n19994;
    n2536_lo_buf_o2 <= n19997;
    n2524_lo_buf_o2 <= n20000;
    G875_o2 <= n20003;
    G1064_o2 <= n20006;
    G1253_o2 <= n20009;
    G6140_o2 <= n20012;
    G5151_o2 <= n20015;
    G5686_o2 <= n20018;
    G6061_o2 <= n20021;
    G4803_o2 <= n20024;
    G5332_o2 <= n20027;
    G5844_o2 <= n20030;
    G6114_o2 <= n20033;
    G4806_o2 <= n20036;
    G3881_o2 <= n20039;
    G4370_o2 <= n20042;
    G4896_o2 <= n20045;
    G5001_o2 <= n20048;
    G3121_o2 <= n20051;
    n2512_lo_buf_o2 <= n20054;
    G4085_o2 <= n20057;
    G4605_o2 <= n20060;
    G5118_o2 <= n20063;
    G4997_o2 <= n20066;
    n2500_lo_buf_o2 <= n20069;
    n2716_lo_buf_o2 <= n20072;
    G560_o2 <= n20075;
    G1895_o2 <= n20078;
    G3064_o2 <= n20081;
    G3269_o2 <= n20084;
    G3569_o2 <= n20087;
    n748_inv <= n20090;
    G1196_o2 <= n20093;
    G1007_o2 <= n20096;
    G818_o2 <= n20099;
    G674_o2 <= n20102;
    G5041_o2 <= n20105;
    G5562_o2 <= n20108;
    G6005_o2 <= n20111;
    G5214_o2 <= n20114;
    G5746_o2 <= n20117;
    G6087_o2 <= n20120;
    G6086_o2 <= n20123;
    G5745_o2 <= n20126;
    G5213_o2 <= n20129;
    G5893_o2 <= n20132;
    G5391_o2 <= n20135;
    G4864_o2 <= n20138;
    G6143_o2 <= n20141;
    G6008_o2 <= n20144;
    G5565_o2 <= n20147;
    G5044_o2 <= n20150;
    G3813_o2 <= n20153;
    G4325_o2 <= n20156;
    G4834_o2 <= n20159;
    G4993_o2 <= n20162;
    G3989_o2 <= n20165;
    G4490_o2 <= n20168;
    G5011_o2 <= n20171;
    G5112_o2 <= n20174;
    n2776_lo_buf_o2 <= n20177;
    G3298_o2 <= n20180;
    G3073_o2 <= n20183;
    G3265_o2 <= n20186;
    G3624_o2 <= n20189;
    G1642_o2 <= n20192;
    G1980_o2 <= n20195;
    n2488_lo_buf_o2 <= n20198;
    G626_o2 <= n20201;
    G1139_o2 <= n20204;
    G950_o2 <= n20207;
    G707_o2 <= n20210;
    G545_o2 <= n20213;
    G4217_o2 <= n20216;
    G4716_o2 <= n20219;
    G5244_o2 <= n20222;
    G3136_o2 <= n20225;
    G3499_o2 <= n20228;
    G3885_o2 <= n20231;
    G5243_o2 <= n20234;
    G3886_o2 <= n20237;
    G4375_o2 <= n20240;
    G4901_o2 <= n20243;
    G5054_o2 <= n20246;
    G4374_o2 <= n20249;
    G4900_o2 <= n20252;
    G5053_o2 <= n20255;
    G5242_o2 <= n20258;
    G4034_o2 <= n20261;
    G4556_o2 <= n20264;
    G5064_o2 <= n20267;
    G5172_o2 <= n20270;
    G2030_o2 <= n20273;
    G3016_o2 <= n20276;
    G3520_o2 <= n20279;
    G3261_o2 <= n20282;
    G3620_o2 <= n20285;
    G4220_o2 <= n20288;
    G4719_o2 <= n20291;
    G5247_o2 <= n20294;
    G5109_o2 <= n20297;
    G1638_o2 <= n20300;
    G1976_o2 <= n20303;
    G3560_o2 <= n20306;
    G3205_o2 <= n20309;
    G3193_o2 <= n20312;
    G3367_o2 <= n20315;
    G3670_o2 <= n20318;
    n979_inv <= n20321;
    G1280_o2 <= n20324;
    G902_o2 <= n20327;
    G659_o2 <= n20330;
    G983_o2 <= n20333;
    G740_o2 <= n20336;
    G2917_o2 <= n20339;
    G3391_o2 <= n20342;
    G3494_o2 <= n20345;
    G1512_o2 <= n20348;
    G1854_o2 <= n20351;
    G2203_o2 <= n20354;
    G3493_o2 <= n20357;
    G3069_o2 <= n20360;
    G3574_o2 <= n20363;
    G3319_o2 <= n20366;
    G3667_o2 <= n20369;
    G3068_o2 <= n20372;
    G3573_o2 <= n20375;
    G3666_o2 <= n20378;
    G3318_o2 <= n20381;
    G3492_o2 <= n20384;
    G3241_o2 <= n20387;
    G3722_o2 <= n20390;
    G3422_o2 <= n20393;
    G1445_o2 <= n20396;
    G3257_o2 <= n20399;
    G3616_o2 <= n20402;
    G1634_o2 <= n20405;
    G1972_o2 <= n20408;
    G2256_o2 <= n20411;
    G3394_o2 <= n20414;
    G3557_o2 <= n20417;
    G3364_o2 <= n20420;
    G3719_o2 <= n20423;
    G2253_o2 <= n20426;
    G1583_o2 <= n20429;
    G1917_o2 <= n20432;
    G1727_o2 <= n20435;
    G2061_o2 <= n20438;
    G935_o2 <= n20441;
    G692_o2 <= n20444;
    G2136_o2 <= n20447;
    G1507_o2 <= n20450;
    G1849_o2 <= n20453;
    G2198_o2 <= n20456;
    G2197_o2 <= n20459;
    G1848_o2 <= n20462;
    G1689_o2 <= n20465;
    G2016_o2 <= n20468;
    G2314_o2 <= n20471;
    G2313_o2 <= n20474;
    G1688_o2 <= n20477;
    G2015_o2 <= n20480;
    G1847_o2 <= n20483;
    G2196_o2 <= n20486;
    G2118_o2 <= n20489;
    G1777_o2 <= n20492;
    G1630_o2 <= n20495;
    G1968_o2 <= n20498;
    G2309_o2 <= n20501;
    G2139_o2 <= n20504;
    G1580_o2 <= n20507;
    G2250_o2 <= n20510;
    G1914_o2 <= n20513;
    G1724_o2 <= n20516;
    G2058_o2 <= n20519;
    n2728_lo_buf_o2 <= n20522;
  end
  initial begin
    n2491_lo <= 1'b0;
    n2575_lo <= 1'b0;
    n2587_lo <= 1'b0;
    n2599_lo <= 1'b0;
    n2611_lo <= 1'b0;
    n2623_lo <= 1'b0;
    n2635_lo <= 1'b0;
    n2647_lo <= 1'b0;
    n2659_lo <= 1'b0;
    n2671_lo <= 1'b0;
    n2683_lo <= 1'b0;
    n2734_lo <= 1'b0;
    n2746_lo <= 1'b0;
    n2758_lo <= 1'b0;
    n2770_lo <= 1'b0;
    n2782_lo <= 1'b0;
    n2785_lo <= 1'b0;
    n2794_lo <= 1'b0;
    n2797_lo <= 1'b0;
    n2806_lo <= 1'b0;
    n2809_lo <= 1'b0;
    n2818_lo <= 1'b0;
    n2821_lo <= 1'b0;
    n2830_lo <= 1'b0;
    n2833_lo <= 1'b0;
    n2836_lo <= 1'b0;
    n2839_lo <= 1'b0;
    n2842_lo <= 1'b0;
    n2845_lo <= 1'b0;
    n2848_lo <= 1'b0;
    n2851_lo <= 1'b0;
    n2854_lo <= 1'b0;
    n2857_lo <= 1'b0;
    n2860_lo <= 1'b0;
    n2863_lo <= 1'b0;
    n4871_o2 <= 1'b0;
    n4893_o2 <= 1'b0;
    n4938_o2 <= 1'b0;
    n5056_o2 <= 1'b0;
    n5100_o2 <= 1'b0;
    n5122_o2 <= 1'b0;
    n5254_o2 <= 1'b0;
    n5276_o2 <= 1'b0;
    n5316_o2 <= 1'b0;
    n5434_o2 <= 1'b0;
    n5473_o2 <= 1'b0;
    n5494_o2 <= 1'b0;
    n5620_o2 <= 1'b0;
    n5643_o2 <= 1'b0;
    n5682_o2 <= 1'b0;
    n5798_o2 <= 1'b0;
    n5839_o2 <= 1'b0;
    n5867_o2 <= 1'b0;
    n6052_o2 <= 1'b0;
    n6087_o2 <= 1'b0;
    n6153_o2 <= 1'b0;
    n6408_o2 <= 1'b0;
    n6454_o2 <= 1'b0;
    n6509_o2 <= 1'b0;
    n6775_o2 <= 1'b0;
    n6818_o2 <= 1'b0;
    n6892_o2 <= 1'b0;
    n5779_o2 <= 1'b0;
    n5780_o2 <= 1'b0;
    n7156_o2 <= 1'b0;
    n5792_o2 <= 1'b0;
    n7205_o2 <= 1'b0;
    n5842_o2 <= 1'b0;
    n5863_o2 <= 1'b0;
    n7263_o2 <= 1'b0;
    n5881_o2 <= 1'b0;
    n5930_o2 <= 1'b0;
    n5959_o2 <= 1'b0;
    n5981_o2 <= 1'b0;
    n6042_o2 <= 1'b0;
    n6075_o2 <= 1'b0;
    n6103_o2 <= 1'b0;
    n7610_o2 <= 1'b0;
    n6169_o2 <= 1'b0;
    n7665_o2 <= 1'b0;
    n6205_o2 <= 1'b0;
    n6239_o2 <= 1'b0;
    n7788_o2 <= 1'b0;
    n6309_o2 <= 1'b0;
    n6461_o2 <= 1'b0;
    n6476_o2 <= 1'b0;
    n325_inv <= 1'b0;
    n6545_o2 <= 1'b0;
    G578_o2 <= 1'b0;
    G5106_o2 <= 1'b0;
    n6713_o2 <= 1'b0;
    G5164_o2 <= 1'b0;
    n343_inv <= 1'b0;
    n6810_o2 <= 1'b0;
    n6973_o2 <= 1'b0;
    n352_inv <= 1'b0;
    n7053_o2 <= 1'b0;
    G581_o2 <= 1'b0;
    G5467_o2 <= 1'b0;
    n7231_o2 <= 1'b0;
    G5527_o2 <= 1'b0;
    n370_inv <= 1'b0;
    n7304_o2 <= 1'b0;
    n7530_o2 <= 1'b0;
    n379_inv <= 1'b0;
    n7653_o2 <= 1'b0;
    G584_o2 <= 1'b0;
    G5820_o2 <= 1'b0;
    n7148_o2 <= 1'b0;
    n7149_o2 <= 1'b0;
    n7224_o2 <= 1'b0;
    n7916_o2 <= 1'b0;
    G5868_o2 <= 1'b0;
    n406_inv <= 1'b0;
    n7280_o2 <= 1'b0;
    n7313_o2 <= 1'b0;
    n8056_o2 <= 1'b0;
    n7323_o2 <= 1'b0;
    n7398_o2 <= 1'b0;
    n7459_o2 <= 1'b0;
    n7501_o2 <= 1'b0;
    n7518_o2 <= 1'b0;
    G563_o2 <= 1'b0;
    n7606_o2 <= 1'b0;
    n439_inv <= 1'b0;
    n7675_o2 <= 1'b0;
    G3410_o2 <= 1'b0;
    n7722_o2 <= 1'b0;
    n7747_o2 <= 1'b0;
    n7835_o2 <= 1'b0;
    G587_o2 <= 1'b0;
    G6046_o2 <= 1'b0;
    n7909_o2 <= 1'b0;
    G566_o2 <= 1'b0;
    G6070_o2 <= 1'b0;
    n472_inv <= 1'b0;
    n8086_o2 <= 1'b0;
    n8093_o2 <= 1'b0;
    G3752_o2 <= 1'b0;
    n484_inv <= 1'b0;
    n8199_o2 <= 1'b0;
    n2800_lo_buf_o2 <= 1'b0;
    G548_o2 <= 1'b0;
    n496_inv <= 1'b0;
    G569_o2 <= 1'b0;
    G1761_o2 <= 1'b0;
    n505_inv <= 1'b0;
    G4101_o2 <= 1'b0;
    G551_o2 <= 1'b0;
    n514_inv <= 1'b0;
    G4743_o2 <= 1'b0;
    G5271_o2 <= 1'b0;
    G5790_o2 <= 1'b0;
    G6122_o2 <= 1'b0;
    G2082_o2 <= 1'b0;
    n2812_lo_buf_o2 <= 1'b0;
    n2668_lo_buf_o2 <= 1'b0;
    n2680_lo_buf_o2 <= 1'b0;
    G572_o2 <= 1'b0;
    G6125_o2 <= 1'b0;
    n547_inv <= 1'b0;
    n2656_lo_buf_o2 <= 1'b0;
    G554_o2 <= 1'b0;
    G4452_o2 <= 1'b0;
    n559_inv <= 1'b0;
    n2644_lo_buf_o2 <= 1'b0;
    G2410_o2 <= 1'b0;
    n2632_lo_buf_o2 <= 1'b0;
    n2620_lo_buf_o2 <= 1'b0;
    G6131_o2 <= 1'b0;
    G4693_o2 <= 1'b0;
    G5209_o2 <= 1'b0;
    G5741_o2 <= 1'b0;
    G6082_o2 <= 1'b0;
    G6119_o2 <= 1'b0;
    n2608_lo_buf_o2 <= 1'b0;
    n2596_lo_buf_o2 <= 1'b0;
    n2584_lo_buf_o2 <= 1'b0;
    n2572_lo_buf_o2 <= 1'b0;
    n2704_lo_buf_o2 <= 1'b0;
    G557_o2 <= 1'b0;
    G5936_o2 <= 1'b0;
    G5442_o2 <= 1'b0;
    G4926_o2 <= 1'b0;
    G6134_o2 <= 1'b0;
    G3929_o2 <= 1'b0;
    G4425_o2 <= 1'b0;
    G4947_o2 <= 1'b0;
    n2764_lo_buf_o2 <= 1'b0;
    n634_inv <= 1'b0;
    n2560_lo_buf_o2 <= 1'b0;
    n2824_lo_buf_o2 <= 1'b0;
    G575_o2 <= 1'b0;
    G2740_o2 <= 1'b0;
    n649_inv <= 1'b0;
    n2548_lo_buf_o2 <= 1'b0;
    n2536_lo_buf_o2 <= 1'b0;
    n2524_lo_buf_o2 <= 1'b0;
    G875_o2 <= 1'b0;
    G1064_o2 <= 1'b0;
    G1253_o2 <= 1'b0;
    G6140_o2 <= 1'b0;
    G5151_o2 <= 1'b0;
    G5686_o2 <= 1'b0;
    G6061_o2 <= 1'b0;
    G4803_o2 <= 1'b0;
    G5332_o2 <= 1'b0;
    G5844_o2 <= 1'b0;
    G6114_o2 <= 1'b0;
    G4806_o2 <= 1'b0;
    G3881_o2 <= 1'b0;
    G4370_o2 <= 1'b0;
    G4896_o2 <= 1'b0;
    G5001_o2 <= 1'b0;
    G3121_o2 <= 1'b0;
    n2512_lo_buf_o2 <= 1'b0;
    G4085_o2 <= 1'b0;
    G4605_o2 <= 1'b0;
    G5118_o2 <= 1'b0;
    G4997_o2 <= 1'b0;
    n2500_lo_buf_o2 <= 1'b0;
    n2716_lo_buf_o2 <= 1'b0;
    G560_o2 <= 1'b0;
    G1895_o2 <= 1'b0;
    G3064_o2 <= 1'b0;
    G3269_o2 <= 1'b0;
    G3569_o2 <= 1'b0;
    n748_inv <= 1'b0;
    G1196_o2 <= 1'b0;
    G1007_o2 <= 1'b0;
    G818_o2 <= 1'b0;
    G674_o2 <= 1'b0;
    G5041_o2 <= 1'b0;
    G5562_o2 <= 1'b0;
    G6005_o2 <= 1'b0;
    G5214_o2 <= 1'b0;
    G5746_o2 <= 1'b0;
    G6087_o2 <= 1'b0;
    G6086_o2 <= 1'b0;
    G5745_o2 <= 1'b0;
    G5213_o2 <= 1'b0;
    G5893_o2 <= 1'b0;
    G5391_o2 <= 1'b0;
    G4864_o2 <= 1'b0;
    G6143_o2 <= 1'b0;
    G6008_o2 <= 1'b0;
    G5565_o2 <= 1'b0;
    G5044_o2 <= 1'b0;
    G3813_o2 <= 1'b0;
    G4325_o2 <= 1'b0;
    G4834_o2 <= 1'b0;
    G4993_o2 <= 1'b0;
    G3989_o2 <= 1'b0;
    G4490_o2 <= 1'b0;
    G5011_o2 <= 1'b0;
    G5112_o2 <= 1'b0;
    n2776_lo_buf_o2 <= 1'b0;
    G3298_o2 <= 1'b0;
    G3073_o2 <= 1'b0;
    G3265_o2 <= 1'b0;
    G3624_o2 <= 1'b0;
    G1642_o2 <= 1'b0;
    G1980_o2 <= 1'b0;
    n2488_lo_buf_o2 <= 1'b0;
    G626_o2 <= 1'b0;
    G1139_o2 <= 1'b0;
    G950_o2 <= 1'b0;
    G707_o2 <= 1'b0;
    G545_o2 <= 1'b0;
    G4217_o2 <= 1'b0;
    G4716_o2 <= 1'b0;
    G5244_o2 <= 1'b0;
    G3136_o2 <= 1'b0;
    G3499_o2 <= 1'b0;
    G3885_o2 <= 1'b0;
    G5243_o2 <= 1'b0;
    G3886_o2 <= 1'b0;
    G4375_o2 <= 1'b0;
    G4901_o2 <= 1'b0;
    G5054_o2 <= 1'b0;
    G4374_o2 <= 1'b0;
    G4900_o2 <= 1'b0;
    G5053_o2 <= 1'b0;
    G5242_o2 <= 1'b0;
    G4034_o2 <= 1'b0;
    G4556_o2 <= 1'b0;
    G5064_o2 <= 1'b0;
    G5172_o2 <= 1'b0;
    G2030_o2 <= 1'b0;
    G3016_o2 <= 1'b0;
    G3520_o2 <= 1'b0;
    G3261_o2 <= 1'b0;
    G3620_o2 <= 1'b0;
    G4220_o2 <= 1'b0;
    G4719_o2 <= 1'b0;
    G5247_o2 <= 1'b0;
    G5109_o2 <= 1'b0;
    G1638_o2 <= 1'b0;
    G1976_o2 <= 1'b0;
    G3560_o2 <= 1'b0;
    G3205_o2 <= 1'b0;
    G3193_o2 <= 1'b0;
    G3367_o2 <= 1'b0;
    G3670_o2 <= 1'b0;
    n979_inv <= 1'b0;
    G1280_o2 <= 1'b0;
    G902_o2 <= 1'b0;
    G659_o2 <= 1'b0;
    G983_o2 <= 1'b0;
    G740_o2 <= 1'b0;
    G2917_o2 <= 1'b0;
    G3391_o2 <= 1'b0;
    G3494_o2 <= 1'b0;
    G1512_o2 <= 1'b0;
    G1854_o2 <= 1'b0;
    G2203_o2 <= 1'b0;
    G3493_o2 <= 1'b0;
    G3069_o2 <= 1'b0;
    G3574_o2 <= 1'b0;
    G3319_o2 <= 1'b0;
    G3667_o2 <= 1'b0;
    G3068_o2 <= 1'b0;
    G3573_o2 <= 1'b0;
    G3666_o2 <= 1'b0;
    G3318_o2 <= 1'b0;
    G3492_o2 <= 1'b0;
    G3241_o2 <= 1'b0;
    G3722_o2 <= 1'b0;
    G3422_o2 <= 1'b0;
    G1445_o2 <= 1'b0;
    G3257_o2 <= 1'b0;
    G3616_o2 <= 1'b0;
    G1634_o2 <= 1'b0;
    G1972_o2 <= 1'b0;
    G2256_o2 <= 1'b0;
    G3394_o2 <= 1'b0;
    G3557_o2 <= 1'b0;
    G3364_o2 <= 1'b0;
    G3719_o2 <= 1'b0;
    G2253_o2 <= 1'b0;
    G1583_o2 <= 1'b0;
    G1917_o2 <= 1'b0;
    G1727_o2 <= 1'b0;
    G2061_o2 <= 1'b0;
    G935_o2 <= 1'b0;
    G692_o2 <= 1'b0;
    G2136_o2 <= 1'b0;
    G1507_o2 <= 1'b0;
    G1849_o2 <= 1'b0;
    G2198_o2 <= 1'b0;
    G2197_o2 <= 1'b0;
    G1848_o2 <= 1'b0;
    G1689_o2 <= 1'b0;
    G2016_o2 <= 1'b0;
    G2314_o2 <= 1'b0;
    G2313_o2 <= 1'b0;
    G1688_o2 <= 1'b0;
    G2015_o2 <= 1'b0;
    G1847_o2 <= 1'b0;
    G2196_o2 <= 1'b0;
    G2118_o2 <= 1'b0;
    G1777_o2 <= 1'b0;
    G1630_o2 <= 1'b0;
    G1968_o2 <= 1'b0;
    G2309_o2 <= 1'b0;
    G2139_o2 <= 1'b0;
    G1580_o2 <= 1'b0;
    G2250_o2 <= 1'b0;
    G1914_o2 <= 1'b0;
    G1724_o2 <= 1'b0;
    G2058_o2 <= 1'b0;
    n2728_lo_buf_o2 <= 1'b0;
  end
endmodule


