
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  n621_lo,
  n630_lo,
  n633_lo,
  n642_lo,
  n645_lo,
  n654_lo,
  n657_lo,
  n666_lo,
  n669_lo,
  n678_lo,
  n681_lo,
  n690_lo,
  n693_lo,
  n702_lo,
  n705_lo,
  n714_lo,
  n717_lo,
  n726_lo,
  n729_lo,
  n738_lo,
  n741_lo,
  n750_lo,
  n753_lo,
  n762_lo,
  n765_lo,
  n774_lo,
  n777_lo,
  n786_lo,
  n789_lo,
  n798_lo,
  n801_lo,
  n810_lo,
  n813_lo,
  n822_lo,
  n825_lo,
  n834_lo,
  n837_lo,
  n846_lo,
  n849_lo,
  n858_lo,
  n861_lo,
  n870_lo,
  n873_lo,
  n882_lo,
  n885_lo,
  n894_lo,
  n897_lo,
  n906_lo,
  n909_lo,
  n918_lo,
  n921_lo,
  n930_lo,
  n933_lo,
  n942_lo,
  n945_lo,
  n954_lo,
  n957_lo,
  n966_lo,
  n969_lo,
  n978_lo,
  n981_lo,
  n990_lo,
  n993_lo,
  n1002_lo,
  n1005_lo,
  n1017_lo,
  n1029_lo,
  n1041_lo,
  n1053_lo,
  n1065_lo,
  n1077_lo,
  n1089_lo,
  n1101_lo,
  n602_o2,
  n639_o2,
  n678_o2,
  n658_o2,
  n783_o2,
  n802_o2,
  n726_o2,
  n763_o2,
  n1644_o2,
  n1645_o2,
  n1646_o2,
  n1647_o2,
  n1648_o2,
  n1649_o2,
  n1650_o2,
  n1651_o2,
  n1652_o2,
  n1653_o2,
  n1654_o2,
  n1655_o2,
  n1656_o2,
  n1657_o2,
  n1658_o2,
  n1659_o2,
  n1660_o2,
  n1661_o2,
  n1662_o2,
  n1663_o2,
  n1664_o2,
  n1665_o2,
  n1666_o2,
  n1667_o2,
  n1668_o2,
  n1669_o2,
  n1670_o2,
  n1671_o2,
  n1672_o2,
  n1673_o2,
  n1674_o2,
  n1675_o2,
  n685_o2,
  n680_o2,
  n822_o2,
  n843_o2,
  n842_o2,
  n681_o2,
  n684_o2,
  n686_o2,
  n823_o2,
  n683_o2,
  n688_o2,
  n803_o2,
  n862_o2,
  n764_o2,
  n863_o2,
  n886_o2,
  lo002_buf_o2,
  lo006_buf_o2,
  lo010_buf_o2,
  lo014_buf_o2,
  lo018_buf_o2,
  lo022_buf_o2,
  lo026_buf_o2,
  lo030_buf_o2,
  lo034_buf_o2,
  lo038_buf_o2,
  lo042_buf_o2,
  lo046_buf_o2,
  lo050_buf_o2,
  lo054_buf_o2,
  lo058_buf_o2,
  lo062_buf_o2,
  lo066_buf_o2,
  lo070_buf_o2,
  lo074_buf_o2,
  lo078_buf_o2,
  lo082_buf_o2,
  lo086_buf_o2,
  lo090_buf_o2,
  lo094_buf_o2,
  lo098_buf_o2,
  lo102_buf_o2,
  lo106_buf_o2,
  lo110_buf_o2,
  lo114_buf_o2,
  lo118_buf_o2,
  lo122_buf_o2,
  lo126_buf_o2,
  n600_o2,
  n601_o2,
  n637_o2,
  n638_o2,
  n676_o2,
  n677_o2,
  n656_o2,
  n657_o2,
  n781_o2,
  n782_o2,
  n800_o2,
  n801_o2,
  n724_o2,
  n725_o2,
  n761_o2,
  n762_o2,
  lo129_buf_o2,
  lo133_buf_o2,
  lo137_buf_o2,
  lo141_buf_o2,
  lo145_buf_o2,
  lo149_buf_o2,
  lo153_buf_o2,
  lo157_buf_o2,
  lo161_buf_o2,
  n571_o2,
  n708_o2,
  n608_o2,
  n665_o2,
  n705_o2,
  n645_o2,
  n745_o2,
  n742_o2,
  n568_o2,
  n717_o2,
  n605_o2,
  n662_o2,
  n714_o2,
  n642_o2,
  n754_o2,
  n751_o2,
  n584_o2,
  n770_o2,
  n789_o2,
  n581_o2,
  n695_o2,
  n732_o2,
  n593_o2,
  n590_o2,
  n630_o2,
  n767_o2,
  n786_o2,
  n627_o2,
  n692_o2,
  n729_o2,
  n621_o2,
  n618_o2,
  G1324,
  G1325,
  G1326,
  G1327,
  G1328,
  G1329,
  G1330,
  G1331,
  G1332,
  G1333,
  G1334,
  G1335,
  G1336,
  G1337,
  G1338,
  G1339,
  G1340,
  G1341,
  G1342,
  G1343,
  G1344,
  G1345,
  G1346,
  G1347,
  G1348,
  G1349,
  G1350,
  G1351,
  G1352,
  G1353,
  G1354,
  G1355,
  n1699_li000_li000,
  n1708_li003_li003,
  n1711_li004_li004,
  n1720_li007_li007,
  n1723_li008_li008,
  n1732_li011_li011,
  n1735_li012_li012,
  n1744_li015_li015,
  n1747_li016_li016,
  n1756_li019_li019,
  n1759_li020_li020,
  n1768_li023_li023,
  n1771_li024_li024,
  n1780_li027_li027,
  n1783_li028_li028,
  n1792_li031_li031,
  n1795_li032_li032,
  n1804_li035_li035,
  n1807_li036_li036,
  n1816_li039_li039,
  n1819_li040_li040,
  n1828_li043_li043,
  n1831_li044_li044,
  n1840_li047_li047,
  n1843_li048_li048,
  n1852_li051_li051,
  n1855_li052_li052,
  n1864_li055_li055,
  n1867_li056_li056,
  n1876_li059_li059,
  n1879_li060_li060,
  n1888_li063_li063,
  n1891_li064_li064,
  n1900_li067_li067,
  n1903_li068_li068,
  n1912_li071_li071,
  n1915_li072_li072,
  n1924_li075_li075,
  n1927_li076_li076,
  n1936_li079_li079,
  n1939_li080_li080,
  n1948_li083_li083,
  n1951_li084_li084,
  n1960_li087_li087,
  n1963_li088_li088,
  n1972_li091_li091,
  n1975_li092_li092,
  n1984_li095_li095,
  n1987_li096_li096,
  n1996_li099_li099,
  n1999_li100_li100,
  n2008_li103_li103,
  n2011_li104_li104,
  n2020_li107_li107,
  n2023_li108_li108,
  n2032_li111_li111,
  n2035_li112_li112,
  n2044_li115_li115,
  n2047_li116_li116,
  n2056_li119_li119,
  n2059_li120_li120,
  n2068_li123_li123,
  n2071_li124_li124,
  n2080_li127_li127,
  n2083_li128_li128,
  n2095_li132_li132,
  n2107_li136_li136,
  n2119_li140_li140,
  n2131_li144_li144,
  n2143_li148_li148,
  n2155_li152_li152,
  n2167_li156_li156,
  n2179_li160_li160,
  n602_i2,
  n639_i2,
  n678_i2,
  n658_i2,
  n783_i2,
  n802_i2,
  n726_i2,
  n763_i2,
  n1644_i2,
  n1645_i2,
  n1646_i2,
  n1647_i2,
  n1648_i2,
  n1649_i2,
  n1650_i2,
  n1651_i2,
  n1652_i2,
  n1653_i2,
  n1654_i2,
  n1655_i2,
  n1656_i2,
  n1657_i2,
  n1658_i2,
  n1659_i2,
  n1660_i2,
  n1661_i2,
  n1662_i2,
  n1663_i2,
  n1664_i2,
  n1665_i2,
  n1666_i2,
  n1667_i2,
  n1668_i2,
  n1669_i2,
  n1670_i2,
  n1671_i2,
  n1672_i2,
  n1673_i2,
  n1674_i2,
  n1675_i2,
  n685_i2,
  n680_i2,
  n822_i2,
  n843_i2,
  n842_i2,
  n681_i2,
  n684_i2,
  n686_i2,
  n823_i2,
  n683_i2,
  n688_i2,
  n803_i2,
  n862_i2,
  n764_i2,
  n863_i2,
  n886_i2,
  lo002_buf_i2,
  lo006_buf_i2,
  lo010_buf_i2,
  lo014_buf_i2,
  lo018_buf_i2,
  lo022_buf_i2,
  lo026_buf_i2,
  lo030_buf_i2,
  lo034_buf_i2,
  lo038_buf_i2,
  lo042_buf_i2,
  lo046_buf_i2,
  lo050_buf_i2,
  lo054_buf_i2,
  lo058_buf_i2,
  lo062_buf_i2,
  lo066_buf_i2,
  lo070_buf_i2,
  lo074_buf_i2,
  lo078_buf_i2,
  lo082_buf_i2,
  lo086_buf_i2,
  lo090_buf_i2,
  lo094_buf_i2,
  lo098_buf_i2,
  lo102_buf_i2,
  lo106_buf_i2,
  lo110_buf_i2,
  lo114_buf_i2,
  lo118_buf_i2,
  lo122_buf_i2,
  lo126_buf_i2,
  n600_i2,
  n601_i2,
  n637_i2,
  n638_i2,
  n676_i2,
  n677_i2,
  n656_i2,
  n657_i2,
  n781_i2,
  n782_i2,
  n800_i2,
  n801_i2,
  n724_i2,
  n725_i2,
  n761_i2,
  n762_i2,
  lo129_buf_i2,
  lo133_buf_i2,
  lo137_buf_i2,
  lo141_buf_i2,
  lo145_buf_i2,
  lo149_buf_i2,
  lo153_buf_i2,
  lo157_buf_i2,
  lo161_buf_i2,
  n571_i2,
  n708_i2,
  n608_i2,
  n665_i2,
  n705_i2,
  n645_i2,
  n745_i2,
  n742_i2,
  n568_i2,
  n717_i2,
  n605_i2,
  n662_i2,
  n714_i2,
  n642_i2,
  n754_i2,
  n751_i2,
  n584_i2,
  n770_i2,
  n789_i2,
  n581_i2,
  n695_i2,
  n732_i2,
  n593_i2,
  n590_i2,
  n630_i2,
  n767_i2,
  n786_i2,
  n627_i2,
  n692_i2,
  n729_i2,
  n621_i2,
  n618_i2
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input n621_lo;input n630_lo;input n633_lo;input n642_lo;input n645_lo;input n654_lo;input n657_lo;input n666_lo;input n669_lo;input n678_lo;input n681_lo;input n690_lo;input n693_lo;input n702_lo;input n705_lo;input n714_lo;input n717_lo;input n726_lo;input n729_lo;input n738_lo;input n741_lo;input n750_lo;input n753_lo;input n762_lo;input n765_lo;input n774_lo;input n777_lo;input n786_lo;input n789_lo;input n798_lo;input n801_lo;input n810_lo;input n813_lo;input n822_lo;input n825_lo;input n834_lo;input n837_lo;input n846_lo;input n849_lo;input n858_lo;input n861_lo;input n870_lo;input n873_lo;input n882_lo;input n885_lo;input n894_lo;input n897_lo;input n906_lo;input n909_lo;input n918_lo;input n921_lo;input n930_lo;input n933_lo;input n942_lo;input n945_lo;input n954_lo;input n957_lo;input n966_lo;input n969_lo;input n978_lo;input n981_lo;input n990_lo;input n993_lo;input n1002_lo;input n1005_lo;input n1017_lo;input n1029_lo;input n1041_lo;input n1053_lo;input n1065_lo;input n1077_lo;input n1089_lo;input n1101_lo;input n602_o2;input n639_o2;input n678_o2;input n658_o2;input n783_o2;input n802_o2;input n726_o2;input n763_o2;input n1644_o2;input n1645_o2;input n1646_o2;input n1647_o2;input n1648_o2;input n1649_o2;input n1650_o2;input n1651_o2;input n1652_o2;input n1653_o2;input n1654_o2;input n1655_o2;input n1656_o2;input n1657_o2;input n1658_o2;input n1659_o2;input n1660_o2;input n1661_o2;input n1662_o2;input n1663_o2;input n1664_o2;input n1665_o2;input n1666_o2;input n1667_o2;input n1668_o2;input n1669_o2;input n1670_o2;input n1671_o2;input n1672_o2;input n1673_o2;input n1674_o2;input n1675_o2;input n685_o2;input n680_o2;input n822_o2;input n843_o2;input n842_o2;input n681_o2;input n684_o2;input n686_o2;input n823_o2;input n683_o2;input n688_o2;input n803_o2;input n862_o2;input n764_o2;input n863_o2;input n886_o2;input lo002_buf_o2;input lo006_buf_o2;input lo010_buf_o2;input lo014_buf_o2;input lo018_buf_o2;input lo022_buf_o2;input lo026_buf_o2;input lo030_buf_o2;input lo034_buf_o2;input lo038_buf_o2;input lo042_buf_o2;input lo046_buf_o2;input lo050_buf_o2;input lo054_buf_o2;input lo058_buf_o2;input lo062_buf_o2;input lo066_buf_o2;input lo070_buf_o2;input lo074_buf_o2;input lo078_buf_o2;input lo082_buf_o2;input lo086_buf_o2;input lo090_buf_o2;input lo094_buf_o2;input lo098_buf_o2;input lo102_buf_o2;input lo106_buf_o2;input lo110_buf_o2;input lo114_buf_o2;input lo118_buf_o2;input lo122_buf_o2;input lo126_buf_o2;input n600_o2;input n601_o2;input n637_o2;input n638_o2;input n676_o2;input n677_o2;input n656_o2;input n657_o2;input n781_o2;input n782_o2;input n800_o2;input n801_o2;input n724_o2;input n725_o2;input n761_o2;input n762_o2;input lo129_buf_o2;input lo133_buf_o2;input lo137_buf_o2;input lo141_buf_o2;input lo145_buf_o2;input lo149_buf_o2;input lo153_buf_o2;input lo157_buf_o2;input lo161_buf_o2;input n571_o2;input n708_o2;input n608_o2;input n665_o2;input n705_o2;input n645_o2;input n745_o2;input n742_o2;input n568_o2;input n717_o2;input n605_o2;input n662_o2;input n714_o2;input n642_o2;input n754_o2;input n751_o2;input n584_o2;input n770_o2;input n789_o2;input n581_o2;input n695_o2;input n732_o2;input n593_o2;input n590_o2;input n630_o2;input n767_o2;input n786_o2;input n627_o2;input n692_o2;input n729_o2;input n621_o2;input n618_o2;
  output G1324;output G1325;output G1326;output G1327;output G1328;output G1329;output G1330;output G1331;output G1332;output G1333;output G1334;output G1335;output G1336;output G1337;output G1338;output G1339;output G1340;output G1341;output G1342;output G1343;output G1344;output G1345;output G1346;output G1347;output G1348;output G1349;output G1350;output G1351;output G1352;output G1353;output G1354;output G1355;output n1699_li000_li000;output n1708_li003_li003;output n1711_li004_li004;output n1720_li007_li007;output n1723_li008_li008;output n1732_li011_li011;output n1735_li012_li012;output n1744_li015_li015;output n1747_li016_li016;output n1756_li019_li019;output n1759_li020_li020;output n1768_li023_li023;output n1771_li024_li024;output n1780_li027_li027;output n1783_li028_li028;output n1792_li031_li031;output n1795_li032_li032;output n1804_li035_li035;output n1807_li036_li036;output n1816_li039_li039;output n1819_li040_li040;output n1828_li043_li043;output n1831_li044_li044;output n1840_li047_li047;output n1843_li048_li048;output n1852_li051_li051;output n1855_li052_li052;output n1864_li055_li055;output n1867_li056_li056;output n1876_li059_li059;output n1879_li060_li060;output n1888_li063_li063;output n1891_li064_li064;output n1900_li067_li067;output n1903_li068_li068;output n1912_li071_li071;output n1915_li072_li072;output n1924_li075_li075;output n1927_li076_li076;output n1936_li079_li079;output n1939_li080_li080;output n1948_li083_li083;output n1951_li084_li084;output n1960_li087_li087;output n1963_li088_li088;output n1972_li091_li091;output n1975_li092_li092;output n1984_li095_li095;output n1987_li096_li096;output n1996_li099_li099;output n1999_li100_li100;output n2008_li103_li103;output n2011_li104_li104;output n2020_li107_li107;output n2023_li108_li108;output n2032_li111_li111;output n2035_li112_li112;output n2044_li115_li115;output n2047_li116_li116;output n2056_li119_li119;output n2059_li120_li120;output n2068_li123_li123;output n2071_li124_li124;output n2080_li127_li127;output n2083_li128_li128;output n2095_li132_li132;output n2107_li136_li136;output n2119_li140_li140;output n2131_li144_li144;output n2143_li148_li148;output n2155_li152_li152;output n2167_li156_li156;output n2179_li160_li160;output n602_i2;output n639_i2;output n678_i2;output n658_i2;output n783_i2;output n802_i2;output n726_i2;output n763_i2;output n1644_i2;output n1645_i2;output n1646_i2;output n1647_i2;output n1648_i2;output n1649_i2;output n1650_i2;output n1651_i2;output n1652_i2;output n1653_i2;output n1654_i2;output n1655_i2;output n1656_i2;output n1657_i2;output n1658_i2;output n1659_i2;output n1660_i2;output n1661_i2;output n1662_i2;output n1663_i2;output n1664_i2;output n1665_i2;output n1666_i2;output n1667_i2;output n1668_i2;output n1669_i2;output n1670_i2;output n1671_i2;output n1672_i2;output n1673_i2;output n1674_i2;output n1675_i2;output n685_i2;output n680_i2;output n822_i2;output n843_i2;output n842_i2;output n681_i2;output n684_i2;output n686_i2;output n823_i2;output n683_i2;output n688_i2;output n803_i2;output n862_i2;output n764_i2;output n863_i2;output n886_i2;output lo002_buf_i2;output lo006_buf_i2;output lo010_buf_i2;output lo014_buf_i2;output lo018_buf_i2;output lo022_buf_i2;output lo026_buf_i2;output lo030_buf_i2;output lo034_buf_i2;output lo038_buf_i2;output lo042_buf_i2;output lo046_buf_i2;output lo050_buf_i2;output lo054_buf_i2;output lo058_buf_i2;output lo062_buf_i2;output lo066_buf_i2;output lo070_buf_i2;output lo074_buf_i2;output lo078_buf_i2;output lo082_buf_i2;output lo086_buf_i2;output lo090_buf_i2;output lo094_buf_i2;output lo098_buf_i2;output lo102_buf_i2;output lo106_buf_i2;output lo110_buf_i2;output lo114_buf_i2;output lo118_buf_i2;output lo122_buf_i2;output lo126_buf_i2;output n600_i2;output n601_i2;output n637_i2;output n638_i2;output n676_i2;output n677_i2;output n656_i2;output n657_i2;output n781_i2;output n782_i2;output n800_i2;output n801_i2;output n724_i2;output n725_i2;output n761_i2;output n762_i2;output lo129_buf_i2;output lo133_buf_i2;output lo137_buf_i2;output lo141_buf_i2;output lo145_buf_i2;output lo149_buf_i2;output lo153_buf_i2;output lo157_buf_i2;output lo161_buf_i2;output n571_i2;output n708_i2;output n608_i2;output n665_i2;output n705_i2;output n645_i2;output n745_i2;output n742_i2;output n568_i2;output n717_i2;output n605_i2;output n662_i2;output n714_i2;output n642_i2;output n754_i2;output n751_i2;output n584_i2;output n770_i2;output n789_i2;output n581_i2;output n695_i2;output n732_i2;output n593_i2;output n590_i2;output n630_i2;output n767_i2;output n786_i2;output n627_i2;output n692_i2;output n729_i2;output n621_i2;output n618_i2;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire n621_lo_p;
  wire n621_lo_n;
  wire n630_lo_p;
  wire n630_lo_n;
  wire n633_lo_p;
  wire n633_lo_n;
  wire n642_lo_p;
  wire n642_lo_n;
  wire n645_lo_p;
  wire n645_lo_n;
  wire n654_lo_p;
  wire n654_lo_n;
  wire n657_lo_p;
  wire n657_lo_n;
  wire n666_lo_p;
  wire n666_lo_n;
  wire n669_lo_p;
  wire n669_lo_n;
  wire n678_lo_p;
  wire n678_lo_n;
  wire n681_lo_p;
  wire n681_lo_n;
  wire n690_lo_p;
  wire n690_lo_n;
  wire n693_lo_p;
  wire n693_lo_n;
  wire n702_lo_p;
  wire n702_lo_n;
  wire n705_lo_p;
  wire n705_lo_n;
  wire n714_lo_p;
  wire n714_lo_n;
  wire n717_lo_p;
  wire n717_lo_n;
  wire n726_lo_p;
  wire n726_lo_n;
  wire n729_lo_p;
  wire n729_lo_n;
  wire n738_lo_p;
  wire n738_lo_n;
  wire n741_lo_p;
  wire n741_lo_n;
  wire n750_lo_p;
  wire n750_lo_n;
  wire n753_lo_p;
  wire n753_lo_n;
  wire n762_lo_p;
  wire n762_lo_n;
  wire n765_lo_p;
  wire n765_lo_n;
  wire n774_lo_p;
  wire n774_lo_n;
  wire n777_lo_p;
  wire n777_lo_n;
  wire n786_lo_p;
  wire n786_lo_n;
  wire n789_lo_p;
  wire n789_lo_n;
  wire n798_lo_p;
  wire n798_lo_n;
  wire n801_lo_p;
  wire n801_lo_n;
  wire n810_lo_p;
  wire n810_lo_n;
  wire n813_lo_p;
  wire n813_lo_n;
  wire n822_lo_p;
  wire n822_lo_n;
  wire n825_lo_p;
  wire n825_lo_n;
  wire n834_lo_p;
  wire n834_lo_n;
  wire n837_lo_p;
  wire n837_lo_n;
  wire n846_lo_p;
  wire n846_lo_n;
  wire n849_lo_p;
  wire n849_lo_n;
  wire n858_lo_p;
  wire n858_lo_n;
  wire n861_lo_p;
  wire n861_lo_n;
  wire n870_lo_p;
  wire n870_lo_n;
  wire n873_lo_p;
  wire n873_lo_n;
  wire n882_lo_p;
  wire n882_lo_n;
  wire n885_lo_p;
  wire n885_lo_n;
  wire n894_lo_p;
  wire n894_lo_n;
  wire n897_lo_p;
  wire n897_lo_n;
  wire n906_lo_p;
  wire n906_lo_n;
  wire n909_lo_p;
  wire n909_lo_n;
  wire n918_lo_p;
  wire n918_lo_n;
  wire n921_lo_p;
  wire n921_lo_n;
  wire n930_lo_p;
  wire n930_lo_n;
  wire n933_lo_p;
  wire n933_lo_n;
  wire n942_lo_p;
  wire n942_lo_n;
  wire n945_lo_p;
  wire n945_lo_n;
  wire n954_lo_p;
  wire n954_lo_n;
  wire n957_lo_p;
  wire n957_lo_n;
  wire n966_lo_p;
  wire n966_lo_n;
  wire n969_lo_p;
  wire n969_lo_n;
  wire n978_lo_p;
  wire n978_lo_n;
  wire n981_lo_p;
  wire n981_lo_n;
  wire n990_lo_p;
  wire n990_lo_n;
  wire n993_lo_p;
  wire n993_lo_n;
  wire n1002_lo_p;
  wire n1002_lo_n;
  wire n1005_lo_p;
  wire n1005_lo_n;
  wire n1017_lo_p;
  wire n1017_lo_n;
  wire n1029_lo_p;
  wire n1029_lo_n;
  wire n1041_lo_p;
  wire n1041_lo_n;
  wire n1053_lo_p;
  wire n1053_lo_n;
  wire n1065_lo_p;
  wire n1065_lo_n;
  wire n1077_lo_p;
  wire n1077_lo_n;
  wire n1089_lo_p;
  wire n1089_lo_n;
  wire n1101_lo_p;
  wire n1101_lo_n;
  wire n602_o2_p;
  wire n602_o2_n;
  wire n639_o2_p;
  wire n639_o2_n;
  wire n678_o2_p;
  wire n678_o2_n;
  wire n658_o2_p;
  wire n658_o2_n;
  wire n783_o2_p;
  wire n783_o2_n;
  wire n802_o2_p;
  wire n802_o2_n;
  wire n726_o2_p;
  wire n726_o2_n;
  wire n763_o2_p;
  wire n763_o2_n;
  wire n1644_o2_p;
  wire n1644_o2_n;
  wire n1645_o2_p;
  wire n1645_o2_n;
  wire n1646_o2_p;
  wire n1646_o2_n;
  wire n1647_o2_p;
  wire n1647_o2_n;
  wire n1648_o2_p;
  wire n1648_o2_n;
  wire n1649_o2_p;
  wire n1649_o2_n;
  wire n1650_o2_p;
  wire n1650_o2_n;
  wire n1651_o2_p;
  wire n1651_o2_n;
  wire n1652_o2_p;
  wire n1652_o2_n;
  wire n1653_o2_p;
  wire n1653_o2_n;
  wire n1654_o2_p;
  wire n1654_o2_n;
  wire n1655_o2_p;
  wire n1655_o2_n;
  wire n1656_o2_p;
  wire n1656_o2_n;
  wire n1657_o2_p;
  wire n1657_o2_n;
  wire n1658_o2_p;
  wire n1658_o2_n;
  wire n1659_o2_p;
  wire n1659_o2_n;
  wire n1660_o2_p;
  wire n1660_o2_n;
  wire n1661_o2_p;
  wire n1661_o2_n;
  wire n1662_o2_p;
  wire n1662_o2_n;
  wire n1663_o2_p;
  wire n1663_o2_n;
  wire n1664_o2_p;
  wire n1664_o2_n;
  wire n1665_o2_p;
  wire n1665_o2_n;
  wire n1666_o2_p;
  wire n1666_o2_n;
  wire n1667_o2_p;
  wire n1667_o2_n;
  wire n1668_o2_p;
  wire n1668_o2_n;
  wire n1669_o2_p;
  wire n1669_o2_n;
  wire n1670_o2_p;
  wire n1670_o2_n;
  wire n1671_o2_p;
  wire n1671_o2_n;
  wire n1672_o2_p;
  wire n1672_o2_n;
  wire n1673_o2_p;
  wire n1673_o2_n;
  wire n1674_o2_p;
  wire n1674_o2_n;
  wire n1675_o2_p;
  wire n1675_o2_n;
  wire n685_o2_p;
  wire n685_o2_n;
  wire n680_o2_p;
  wire n680_o2_n;
  wire n822_o2_p;
  wire n822_o2_n;
  wire n843_o2_p;
  wire n843_o2_n;
  wire n842_o2_p;
  wire n842_o2_n;
  wire n681_o2_p;
  wire n681_o2_n;
  wire n684_o2_p;
  wire n684_o2_n;
  wire n686_o2_p;
  wire n686_o2_n;
  wire n823_o2_p;
  wire n823_o2_n;
  wire n683_o2_p;
  wire n683_o2_n;
  wire n688_o2_p;
  wire n688_o2_n;
  wire n803_o2_p;
  wire n803_o2_n;
  wire n862_o2_p;
  wire n862_o2_n;
  wire n764_o2_p;
  wire n764_o2_n;
  wire n863_o2_p;
  wire n863_o2_n;
  wire n886_o2_p;
  wire n886_o2_n;
  wire lo002_buf_o2_p;
  wire lo002_buf_o2_n;
  wire lo006_buf_o2_p;
  wire lo006_buf_o2_n;
  wire lo010_buf_o2_p;
  wire lo010_buf_o2_n;
  wire lo014_buf_o2_p;
  wire lo014_buf_o2_n;
  wire lo018_buf_o2_p;
  wire lo018_buf_o2_n;
  wire lo022_buf_o2_p;
  wire lo022_buf_o2_n;
  wire lo026_buf_o2_p;
  wire lo026_buf_o2_n;
  wire lo030_buf_o2_p;
  wire lo030_buf_o2_n;
  wire lo034_buf_o2_p;
  wire lo034_buf_o2_n;
  wire lo038_buf_o2_p;
  wire lo038_buf_o2_n;
  wire lo042_buf_o2_p;
  wire lo042_buf_o2_n;
  wire lo046_buf_o2_p;
  wire lo046_buf_o2_n;
  wire lo050_buf_o2_p;
  wire lo050_buf_o2_n;
  wire lo054_buf_o2_p;
  wire lo054_buf_o2_n;
  wire lo058_buf_o2_p;
  wire lo058_buf_o2_n;
  wire lo062_buf_o2_p;
  wire lo062_buf_o2_n;
  wire lo066_buf_o2_p;
  wire lo066_buf_o2_n;
  wire lo070_buf_o2_p;
  wire lo070_buf_o2_n;
  wire lo074_buf_o2_p;
  wire lo074_buf_o2_n;
  wire lo078_buf_o2_p;
  wire lo078_buf_o2_n;
  wire lo082_buf_o2_p;
  wire lo082_buf_o2_n;
  wire lo086_buf_o2_p;
  wire lo086_buf_o2_n;
  wire lo090_buf_o2_p;
  wire lo090_buf_o2_n;
  wire lo094_buf_o2_p;
  wire lo094_buf_o2_n;
  wire lo098_buf_o2_p;
  wire lo098_buf_o2_n;
  wire lo102_buf_o2_p;
  wire lo102_buf_o2_n;
  wire lo106_buf_o2_p;
  wire lo106_buf_o2_n;
  wire lo110_buf_o2_p;
  wire lo110_buf_o2_n;
  wire lo114_buf_o2_p;
  wire lo114_buf_o2_n;
  wire lo118_buf_o2_p;
  wire lo118_buf_o2_n;
  wire lo122_buf_o2_p;
  wire lo122_buf_o2_n;
  wire lo126_buf_o2_p;
  wire lo126_buf_o2_n;
  wire n600_o2_p;
  wire n600_o2_n;
  wire n601_o2_p;
  wire n601_o2_n;
  wire n637_o2_p;
  wire n637_o2_n;
  wire n638_o2_p;
  wire n638_o2_n;
  wire n676_o2_p;
  wire n676_o2_n;
  wire n677_o2_p;
  wire n677_o2_n;
  wire n656_o2_p;
  wire n656_o2_n;
  wire n657_o2_p;
  wire n657_o2_n;
  wire n781_o2_p;
  wire n781_o2_n;
  wire n782_o2_p;
  wire n782_o2_n;
  wire n800_o2_p;
  wire n800_o2_n;
  wire n801_o2_p;
  wire n801_o2_n;
  wire n724_o2_p;
  wire n724_o2_n;
  wire n725_o2_p;
  wire n725_o2_n;
  wire n761_o2_p;
  wire n761_o2_n;
  wire n762_o2_p;
  wire n762_o2_n;
  wire lo129_buf_o2_p;
  wire lo129_buf_o2_n;
  wire lo133_buf_o2_p;
  wire lo133_buf_o2_n;
  wire lo137_buf_o2_p;
  wire lo137_buf_o2_n;
  wire lo141_buf_o2_p;
  wire lo141_buf_o2_n;
  wire lo145_buf_o2_p;
  wire lo145_buf_o2_n;
  wire lo149_buf_o2_p;
  wire lo149_buf_o2_n;
  wire lo153_buf_o2_p;
  wire lo153_buf_o2_n;
  wire lo157_buf_o2_p;
  wire lo157_buf_o2_n;
  wire lo161_buf_o2_p;
  wire lo161_buf_o2_n;
  wire n571_o2_p;
  wire n571_o2_n;
  wire n708_o2_p;
  wire n708_o2_n;
  wire n608_o2_p;
  wire n608_o2_n;
  wire n665_o2_p;
  wire n665_o2_n;
  wire n705_o2_p;
  wire n705_o2_n;
  wire n645_o2_p;
  wire n645_o2_n;
  wire n745_o2_p;
  wire n745_o2_n;
  wire n742_o2_p;
  wire n742_o2_n;
  wire n568_o2_p;
  wire n568_o2_n;
  wire n717_o2_p;
  wire n717_o2_n;
  wire n605_o2_p;
  wire n605_o2_n;
  wire n662_o2_p;
  wire n662_o2_n;
  wire n714_o2_p;
  wire n714_o2_n;
  wire n642_o2_p;
  wire n642_o2_n;
  wire n754_o2_p;
  wire n754_o2_n;
  wire n751_o2_p;
  wire n751_o2_n;
  wire n584_o2_p;
  wire n584_o2_n;
  wire n770_o2_p;
  wire n770_o2_n;
  wire n789_o2_p;
  wire n789_o2_n;
  wire n581_o2_p;
  wire n581_o2_n;
  wire n695_o2_p;
  wire n695_o2_n;
  wire n732_o2_p;
  wire n732_o2_n;
  wire n593_o2_p;
  wire n593_o2_n;
  wire n590_o2_p;
  wire n590_o2_n;
  wire n630_o2_p;
  wire n630_o2_n;
  wire n767_o2_p;
  wire n767_o2_n;
  wire n786_o2_p;
  wire n786_o2_n;
  wire n627_o2_p;
  wire n627_o2_n;
  wire n692_o2_p;
  wire n692_o2_n;
  wire n729_o2_p;
  wire n729_o2_n;
  wire n621_o2_p;
  wire n621_o2_n;
  wire n618_o2_p;
  wire n618_o2_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g260_n_spl_;
  wire g260_n_spl_0;
  wire g260_n_spl_1;
  wire g260_p_spl_;
  wire g260_p_spl_0;
  wire g260_p_spl_1;
  wire n602_o2_p_spl_;
  wire n602_o2_p_spl_0;
  wire n602_o2_p_spl_1;
  wire g262_p_spl_;
  wire g262_p_spl_0;
  wire g262_p_spl_1;
  wire n602_o2_n_spl_;
  wire n602_o2_n_spl_0;
  wire n602_o2_n_spl_1;
  wire g262_n_spl_;
  wire g262_n_spl_0;
  wire g262_n_spl_1;
  wire n639_o2_p_spl_;
  wire n639_o2_p_spl_0;
  wire n639_o2_p_spl_00;
  wire n639_o2_p_spl_1;
  wire n639_o2_n_spl_;
  wire n639_o2_n_spl_0;
  wire n639_o2_n_spl_00;
  wire n639_o2_n_spl_1;
  wire n678_o2_p_spl_;
  wire n678_o2_p_spl_0;
  wire n678_o2_p_spl_00;
  wire n678_o2_p_spl_01;
  wire n678_o2_p_spl_1;
  wire n678_o2_n_spl_;
  wire n678_o2_n_spl_0;
  wire n678_o2_n_spl_00;
  wire n678_o2_n_spl_01;
  wire n678_o2_n_spl_1;
  wire n658_o2_p_spl_;
  wire n658_o2_p_spl_0;
  wire n658_o2_p_spl_1;
  wire n658_o2_n_spl_;
  wire n658_o2_n_spl_0;
  wire n658_o2_n_spl_1;
  wire g280_p_spl_;
  wire g280_p_spl_0;
  wire g280_p_spl_1;
  wire g280_n_spl_;
  wire g280_n_spl_0;
  wire g280_n_spl_1;
  wire g298_p_spl_;
  wire g298_p_spl_0;
  wire g298_p_spl_1;
  wire g298_n_spl_;
  wire g298_n_spl_0;
  wire g298_n_spl_1;
  wire g316_p_spl_;
  wire g316_p_spl_0;
  wire g316_p_spl_1;
  wire g316_n_spl_;
  wire g316_n_spl_0;
  wire g316_n_spl_1;
  wire n886_o2_p_spl_;
  wire n886_o2_p_spl_0;
  wire n886_o2_p_spl_1;
  wire n886_o2_n_spl_;
  wire n886_o2_n_spl_0;
  wire n886_o2_n_spl_1;
  wire n783_o2_p_spl_;
  wire n783_o2_p_spl_0;
  wire n783_o2_p_spl_1;
  wire g334_p_spl_;
  wire g334_p_spl_0;
  wire g334_p_spl_1;
  wire n783_o2_n_spl_;
  wire n783_o2_n_spl_0;
  wire n783_o2_n_spl_1;
  wire g334_n_spl_;
  wire g334_n_spl_0;
  wire g334_n_spl_1;
  wire n802_o2_p_spl_;
  wire n802_o2_p_spl_0;
  wire n802_o2_p_spl_1;
  wire n802_o2_n_spl_;
  wire n802_o2_n_spl_0;
  wire n802_o2_n_spl_1;
  wire n726_o2_p_spl_;
  wire n726_o2_p_spl_0;
  wire n726_o2_p_spl_1;
  wire n726_o2_n_spl_;
  wire n726_o2_n_spl_0;
  wire n726_o2_n_spl_1;
  wire n763_o2_p_spl_;
  wire n763_o2_p_spl_0;
  wire n763_o2_p_spl_1;
  wire n763_o2_n_spl_;
  wire n763_o2_n_spl_0;
  wire n763_o2_n_spl_1;
  wire g352_p_spl_;
  wire g352_p_spl_0;
  wire g352_p_spl_1;
  wire g352_n_spl_;
  wire g352_n_spl_0;
  wire g352_n_spl_1;
  wire g370_p_spl_;
  wire g370_p_spl_0;
  wire g370_p_spl_1;
  wire g370_n_spl_;
  wire g370_n_spl_0;
  wire g370_n_spl_1;
  wire g388_p_spl_;
  wire g388_p_spl_0;
  wire g388_p_spl_1;
  wire g388_n_spl_;
  wire g388_n_spl_0;
  wire g388_n_spl_1;
  wire g406_n_spl_;
  wire g406_n_spl_0;
  wire g407_n_spl_;
  wire g407_n_spl_0;
  wire g409_p_spl_;
  wire g409_p_spl_0;
  wire g412_p_spl_;
  wire g412_p_spl_0;
  wire g409_n_spl_;
  wire g409_n_spl_0;
  wire g412_n_spl_;
  wire g412_n_spl_0;
  wire g410_p_spl_;
  wire g410_p_spl_0;
  wire g411_p_spl_;
  wire g411_p_spl_0;
  wire g405_n_spl_;
  wire g405_n_spl_0;
  wire g414_n_spl_;
  wire g408_n_spl_;
  wire g408_n_spl_0;
  wire g419_n_spl_;
  wire g413_n_spl_;
  wire g410_n_spl_;
  wire g410_n_spl_0;
  wire g411_n_spl_;
  wire g411_n_spl_0;
  wire g418_n_spl_;
  wire g420_n_spl_;
  wire g421_n_spl_;
  wire g415_n_spl_;
  wire g416_n_spl_;
  wire g422_n_spl_;
  wire g417_n_spl_;
  wire n571_o2_p_spl_;
  wire n568_o2_n_spl_;
  wire n571_o2_n_spl_;
  wire n568_o2_p_spl_;
  wire lo161_buf_o2_p_spl_;
  wire lo161_buf_o2_p_spl_0;
  wire lo161_buf_o2_p_spl_00;
  wire lo161_buf_o2_p_spl_01;
  wire lo161_buf_o2_p_spl_1;
  wire lo161_buf_o2_p_spl_10;
  wire lo161_buf_o2_p_spl_11;
  wire lo161_buf_o2_n_spl_;
  wire lo161_buf_o2_n_spl_0;
  wire lo161_buf_o2_n_spl_00;
  wire lo161_buf_o2_n_spl_01;
  wire lo161_buf_o2_n_spl_1;
  wire lo161_buf_o2_n_spl_10;
  wire lo161_buf_o2_n_spl_11;
  wire n584_o2_p_spl_;
  wire n581_o2_n_spl_;
  wire n584_o2_n_spl_;
  wire n581_o2_p_spl_;
  wire n593_o2_p_spl_;
  wire n590_o2_n_spl_;
  wire n593_o2_n_spl_;
  wire n590_o2_p_spl_;
  wire g446_p_spl_;
  wire g449_n_spl_;
  wire g446_n_spl_;
  wire g449_p_spl_;
  wire g443_n_spl_;
  wire g452_n_spl_;
  wire n608_o2_p_spl_;
  wire n605_o2_n_spl_;
  wire n608_o2_n_spl_;
  wire n605_o2_p_spl_;
  wire n621_o2_p_spl_;
  wire n618_o2_n_spl_;
  wire n621_o2_n_spl_;
  wire n618_o2_p_spl_;
  wire n630_o2_p_spl_;
  wire n627_o2_n_spl_;
  wire n630_o2_n_spl_;
  wire n627_o2_p_spl_;
  wire g464_p_spl_;
  wire g467_n_spl_;
  wire g464_n_spl_;
  wire g467_p_spl_;
  wire g461_n_spl_;
  wire g470_n_spl_;
  wire n665_o2_p_spl_;
  wire n662_o2_n_spl_;
  wire n665_o2_n_spl_;
  wire n662_o2_p_spl_;
  wire g479_n_spl_;
  wire g482_n_spl_;
  wire n645_o2_p_spl_;
  wire n642_o2_n_spl_;
  wire n645_o2_n_spl_;
  wire n642_o2_p_spl_;
  wire g491_n_spl_;
  wire g494_n_spl_;
  wire n770_o2_p_spl_;
  wire n767_o2_n_spl_;
  wire n770_o2_n_spl_;
  wire n767_o2_p_spl_;
  wire n708_o2_p_spl_;
  wire n705_o2_n_spl_;
  wire n708_o2_n_spl_;
  wire n705_o2_p_spl_;
  wire n745_o2_p_spl_;
  wire n742_o2_n_spl_;
  wire n745_o2_n_spl_;
  wire n742_o2_p_spl_;
  wire g506_p_spl_;
  wire g509_n_spl_;
  wire g506_n_spl_;
  wire g509_p_spl_;
  wire g503_n_spl_;
  wire g512_n_spl_;
  wire n789_o2_p_spl_;
  wire n786_o2_n_spl_;
  wire n789_o2_n_spl_;
  wire n786_o2_p_spl_;
  wire n717_o2_p_spl_;
  wire n714_o2_n_spl_;
  wire n717_o2_n_spl_;
  wire n714_o2_p_spl_;
  wire n754_o2_p_spl_;
  wire n751_o2_n_spl_;
  wire n754_o2_n_spl_;
  wire n751_o2_p_spl_;
  wire g524_p_spl_;
  wire g527_n_spl_;
  wire g524_n_spl_;
  wire g527_p_spl_;
  wire g521_n_spl_;
  wire g530_n_spl_;
  wire n695_o2_p_spl_;
  wire n692_o2_n_spl_;
  wire n695_o2_n_spl_;
  wire n692_o2_p_spl_;
  wire g539_n_spl_;
  wire g542_n_spl_;
  wire n732_o2_p_spl_;
  wire n729_o2_n_spl_;
  wire n732_o2_n_spl_;
  wire n729_o2_p_spl_;
  wire g551_n_spl_;
  wire g554_n_spl_;
  wire n621_lo_p_spl_;
  wire n621_lo_p_spl_0;
  wire n669_lo_p_spl_;
  wire n669_lo_p_spl_0;
  wire n621_lo_n_spl_;
  wire n669_lo_n_spl_;
  wire n633_lo_p_spl_;
  wire n633_lo_p_spl_0;
  wire n633_lo_n_spl_;
  wire n681_lo_p_spl_;
  wire n681_lo_p_spl_0;
  wire n681_lo_n_spl_;
  wire n645_lo_p_spl_;
  wire n645_lo_p_spl_0;
  wire n693_lo_p_spl_;
  wire n693_lo_p_spl_0;
  wire n645_lo_n_spl_;
  wire n693_lo_n_spl_;
  wire n657_lo_n_spl_;
  wire n657_lo_p_spl_;
  wire n657_lo_p_spl_0;
  wire n705_lo_p_spl_;
  wire n705_lo_p_spl_0;
  wire n705_lo_n_spl_;
  wire n717_lo_p_spl_;
  wire n717_lo_p_spl_0;
  wire n765_lo_n_spl_;
  wire n717_lo_n_spl_;
  wire n765_lo_p_spl_;
  wire n765_lo_p_spl_0;
  wire n729_lo_p_spl_;
  wire n729_lo_p_spl_0;
  wire n729_lo_n_spl_;
  wire n777_lo_n_spl_;
  wire n777_lo_p_spl_;
  wire n777_lo_p_spl_0;
  wire n741_lo_p_spl_;
  wire n741_lo_p_spl_0;
  wire n789_lo_n_spl_;
  wire n741_lo_n_spl_;
  wire n789_lo_p_spl_;
  wire n789_lo_p_spl_0;
  wire n753_lo_n_spl_;
  wire n753_lo_p_spl_;
  wire n753_lo_p_spl_0;
  wire n801_lo_n_spl_;
  wire n801_lo_p_spl_;
  wire n801_lo_p_spl_0;
  wire n813_lo_p_spl_;
  wire n813_lo_p_spl_0;
  wire n825_lo_p_spl_;
  wire n825_lo_p_spl_0;
  wire n813_lo_n_spl_;
  wire n825_lo_n_spl_;
  wire n861_lo_p_spl_;
  wire n861_lo_p_spl_0;
  wire n861_lo_n_spl_;
  wire n873_lo_p_spl_;
  wire n873_lo_p_spl_0;
  wire n873_lo_n_spl_;
  wire n837_lo_p_spl_;
  wire n837_lo_p_spl_0;
  wire n849_lo_n_spl_;
  wire n837_lo_n_spl_;
  wire n849_lo_p_spl_;
  wire n849_lo_p_spl_0;
  wire n885_lo_p_spl_;
  wire n885_lo_p_spl_0;
  wire n885_lo_n_spl_;
  wire n897_lo_p_spl_;
  wire n897_lo_p_spl_0;
  wire n897_lo_n_spl_;
  wire n909_lo_p_spl_;
  wire n909_lo_p_spl_0;
  wire n921_lo_p_spl_;
  wire n921_lo_p_spl_0;
  wire n909_lo_n_spl_;
  wire n921_lo_n_spl_;
  wire n957_lo_n_spl_;
  wire n957_lo_p_spl_;
  wire n957_lo_p_spl_0;
  wire n969_lo_n_spl_;
  wire n969_lo_p_spl_;
  wire n969_lo_p_spl_0;
  wire n933_lo_p_spl_;
  wire n933_lo_p_spl_0;
  wire n945_lo_n_spl_;
  wire n933_lo_n_spl_;
  wire n945_lo_p_spl_;
  wire n945_lo_p_spl_0;
  wire n981_lo_n_spl_;
  wire n981_lo_p_spl_;
  wire n981_lo_p_spl_0;
  wire n993_lo_n_spl_;
  wire n993_lo_p_spl_;
  wire n993_lo_p_spl_0;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    G37_p,
    G37
  );


  not

  (
    G37_n,
    G37
  );


  buf

  (
    G38_p,
    G38
  );


  not

  (
    G38_n,
    G38
  );


  buf

  (
    G39_p,
    G39
  );


  not

  (
    G39_n,
    G39
  );


  buf

  (
    G40_p,
    G40
  );


  not

  (
    G40_n,
    G40
  );


  buf

  (
    G41_p,
    G41
  );


  not

  (
    G41_n,
    G41
  );


  buf

  (
    n621_lo_p,
    n621_lo
  );


  not

  (
    n621_lo_n,
    n621_lo
  );


  buf

  (
    n630_lo_p,
    n630_lo
  );


  not

  (
    n630_lo_n,
    n630_lo
  );


  buf

  (
    n633_lo_p,
    n633_lo
  );


  not

  (
    n633_lo_n,
    n633_lo
  );


  buf

  (
    n642_lo_p,
    n642_lo
  );


  not

  (
    n642_lo_n,
    n642_lo
  );


  buf

  (
    n645_lo_p,
    n645_lo
  );


  not

  (
    n645_lo_n,
    n645_lo
  );


  buf

  (
    n654_lo_p,
    n654_lo
  );


  not

  (
    n654_lo_n,
    n654_lo
  );


  buf

  (
    n657_lo_p,
    n657_lo
  );


  not

  (
    n657_lo_n,
    n657_lo
  );


  buf

  (
    n666_lo_p,
    n666_lo
  );


  not

  (
    n666_lo_n,
    n666_lo
  );


  buf

  (
    n669_lo_p,
    n669_lo
  );


  not

  (
    n669_lo_n,
    n669_lo
  );


  buf

  (
    n678_lo_p,
    n678_lo
  );


  not

  (
    n678_lo_n,
    n678_lo
  );


  buf

  (
    n681_lo_p,
    n681_lo
  );


  not

  (
    n681_lo_n,
    n681_lo
  );


  buf

  (
    n690_lo_p,
    n690_lo
  );


  not

  (
    n690_lo_n,
    n690_lo
  );


  buf

  (
    n693_lo_p,
    n693_lo
  );


  not

  (
    n693_lo_n,
    n693_lo
  );


  buf

  (
    n702_lo_p,
    n702_lo
  );


  not

  (
    n702_lo_n,
    n702_lo
  );


  buf

  (
    n705_lo_p,
    n705_lo
  );


  not

  (
    n705_lo_n,
    n705_lo
  );


  buf

  (
    n714_lo_p,
    n714_lo
  );


  not

  (
    n714_lo_n,
    n714_lo
  );


  buf

  (
    n717_lo_p,
    n717_lo
  );


  not

  (
    n717_lo_n,
    n717_lo
  );


  buf

  (
    n726_lo_p,
    n726_lo
  );


  not

  (
    n726_lo_n,
    n726_lo
  );


  buf

  (
    n729_lo_p,
    n729_lo
  );


  not

  (
    n729_lo_n,
    n729_lo
  );


  buf

  (
    n738_lo_p,
    n738_lo
  );


  not

  (
    n738_lo_n,
    n738_lo
  );


  buf

  (
    n741_lo_p,
    n741_lo
  );


  not

  (
    n741_lo_n,
    n741_lo
  );


  buf

  (
    n750_lo_p,
    n750_lo
  );


  not

  (
    n750_lo_n,
    n750_lo
  );


  buf

  (
    n753_lo_p,
    n753_lo
  );


  not

  (
    n753_lo_n,
    n753_lo
  );


  buf

  (
    n762_lo_p,
    n762_lo
  );


  not

  (
    n762_lo_n,
    n762_lo
  );


  buf

  (
    n765_lo_p,
    n765_lo
  );


  not

  (
    n765_lo_n,
    n765_lo
  );


  buf

  (
    n774_lo_p,
    n774_lo
  );


  not

  (
    n774_lo_n,
    n774_lo
  );


  buf

  (
    n777_lo_p,
    n777_lo
  );


  not

  (
    n777_lo_n,
    n777_lo
  );


  buf

  (
    n786_lo_p,
    n786_lo
  );


  not

  (
    n786_lo_n,
    n786_lo
  );


  buf

  (
    n789_lo_p,
    n789_lo
  );


  not

  (
    n789_lo_n,
    n789_lo
  );


  buf

  (
    n798_lo_p,
    n798_lo
  );


  not

  (
    n798_lo_n,
    n798_lo
  );


  buf

  (
    n801_lo_p,
    n801_lo
  );


  not

  (
    n801_lo_n,
    n801_lo
  );


  buf

  (
    n810_lo_p,
    n810_lo
  );


  not

  (
    n810_lo_n,
    n810_lo
  );


  buf

  (
    n813_lo_p,
    n813_lo
  );


  not

  (
    n813_lo_n,
    n813_lo
  );


  buf

  (
    n822_lo_p,
    n822_lo
  );


  not

  (
    n822_lo_n,
    n822_lo
  );


  buf

  (
    n825_lo_p,
    n825_lo
  );


  not

  (
    n825_lo_n,
    n825_lo
  );


  buf

  (
    n834_lo_p,
    n834_lo
  );


  not

  (
    n834_lo_n,
    n834_lo
  );


  buf

  (
    n837_lo_p,
    n837_lo
  );


  not

  (
    n837_lo_n,
    n837_lo
  );


  buf

  (
    n846_lo_p,
    n846_lo
  );


  not

  (
    n846_lo_n,
    n846_lo
  );


  buf

  (
    n849_lo_p,
    n849_lo
  );


  not

  (
    n849_lo_n,
    n849_lo
  );


  buf

  (
    n858_lo_p,
    n858_lo
  );


  not

  (
    n858_lo_n,
    n858_lo
  );


  buf

  (
    n861_lo_p,
    n861_lo
  );


  not

  (
    n861_lo_n,
    n861_lo
  );


  buf

  (
    n870_lo_p,
    n870_lo
  );


  not

  (
    n870_lo_n,
    n870_lo
  );


  buf

  (
    n873_lo_p,
    n873_lo
  );


  not

  (
    n873_lo_n,
    n873_lo
  );


  buf

  (
    n882_lo_p,
    n882_lo
  );


  not

  (
    n882_lo_n,
    n882_lo
  );


  buf

  (
    n885_lo_p,
    n885_lo
  );


  not

  (
    n885_lo_n,
    n885_lo
  );


  buf

  (
    n894_lo_p,
    n894_lo
  );


  not

  (
    n894_lo_n,
    n894_lo
  );


  buf

  (
    n897_lo_p,
    n897_lo
  );


  not

  (
    n897_lo_n,
    n897_lo
  );


  buf

  (
    n906_lo_p,
    n906_lo
  );


  not

  (
    n906_lo_n,
    n906_lo
  );


  buf

  (
    n909_lo_p,
    n909_lo
  );


  not

  (
    n909_lo_n,
    n909_lo
  );


  buf

  (
    n918_lo_p,
    n918_lo
  );


  not

  (
    n918_lo_n,
    n918_lo
  );


  buf

  (
    n921_lo_p,
    n921_lo
  );


  not

  (
    n921_lo_n,
    n921_lo
  );


  buf

  (
    n930_lo_p,
    n930_lo
  );


  not

  (
    n930_lo_n,
    n930_lo
  );


  buf

  (
    n933_lo_p,
    n933_lo
  );


  not

  (
    n933_lo_n,
    n933_lo
  );


  buf

  (
    n942_lo_p,
    n942_lo
  );


  not

  (
    n942_lo_n,
    n942_lo
  );


  buf

  (
    n945_lo_p,
    n945_lo
  );


  not

  (
    n945_lo_n,
    n945_lo
  );


  buf

  (
    n954_lo_p,
    n954_lo
  );


  not

  (
    n954_lo_n,
    n954_lo
  );


  buf

  (
    n957_lo_p,
    n957_lo
  );


  not

  (
    n957_lo_n,
    n957_lo
  );


  buf

  (
    n966_lo_p,
    n966_lo
  );


  not

  (
    n966_lo_n,
    n966_lo
  );


  buf

  (
    n969_lo_p,
    n969_lo
  );


  not

  (
    n969_lo_n,
    n969_lo
  );


  buf

  (
    n978_lo_p,
    n978_lo
  );


  not

  (
    n978_lo_n,
    n978_lo
  );


  buf

  (
    n981_lo_p,
    n981_lo
  );


  not

  (
    n981_lo_n,
    n981_lo
  );


  buf

  (
    n990_lo_p,
    n990_lo
  );


  not

  (
    n990_lo_n,
    n990_lo
  );


  buf

  (
    n993_lo_p,
    n993_lo
  );


  not

  (
    n993_lo_n,
    n993_lo
  );


  buf

  (
    n1002_lo_p,
    n1002_lo
  );


  not

  (
    n1002_lo_n,
    n1002_lo
  );


  buf

  (
    n1005_lo_p,
    n1005_lo
  );


  not

  (
    n1005_lo_n,
    n1005_lo
  );


  buf

  (
    n1017_lo_p,
    n1017_lo
  );


  not

  (
    n1017_lo_n,
    n1017_lo
  );


  buf

  (
    n1029_lo_p,
    n1029_lo
  );


  not

  (
    n1029_lo_n,
    n1029_lo
  );


  buf

  (
    n1041_lo_p,
    n1041_lo
  );


  not

  (
    n1041_lo_n,
    n1041_lo
  );


  buf

  (
    n1053_lo_p,
    n1053_lo
  );


  not

  (
    n1053_lo_n,
    n1053_lo
  );


  buf

  (
    n1065_lo_p,
    n1065_lo
  );


  not

  (
    n1065_lo_n,
    n1065_lo
  );


  buf

  (
    n1077_lo_p,
    n1077_lo
  );


  not

  (
    n1077_lo_n,
    n1077_lo
  );


  buf

  (
    n1089_lo_p,
    n1089_lo
  );


  not

  (
    n1089_lo_n,
    n1089_lo
  );


  buf

  (
    n1101_lo_p,
    n1101_lo
  );


  not

  (
    n1101_lo_n,
    n1101_lo
  );


  buf

  (
    n602_o2_p,
    n602_o2
  );


  not

  (
    n602_o2_n,
    n602_o2
  );


  buf

  (
    n639_o2_p,
    n639_o2
  );


  not

  (
    n639_o2_n,
    n639_o2
  );


  buf

  (
    n678_o2_p,
    n678_o2
  );


  not

  (
    n678_o2_n,
    n678_o2
  );


  buf

  (
    n658_o2_p,
    n658_o2
  );


  not

  (
    n658_o2_n,
    n658_o2
  );


  buf

  (
    n783_o2_p,
    n783_o2
  );


  not

  (
    n783_o2_n,
    n783_o2
  );


  buf

  (
    n802_o2_p,
    n802_o2
  );


  not

  (
    n802_o2_n,
    n802_o2
  );


  buf

  (
    n726_o2_p,
    n726_o2
  );


  not

  (
    n726_o2_n,
    n726_o2
  );


  buf

  (
    n763_o2_p,
    n763_o2
  );


  not

  (
    n763_o2_n,
    n763_o2
  );


  buf

  (
    n1644_o2_p,
    n1644_o2
  );


  not

  (
    n1644_o2_n,
    n1644_o2
  );


  buf

  (
    n1645_o2_p,
    n1645_o2
  );


  not

  (
    n1645_o2_n,
    n1645_o2
  );


  buf

  (
    n1646_o2_p,
    n1646_o2
  );


  not

  (
    n1646_o2_n,
    n1646_o2
  );


  buf

  (
    n1647_o2_p,
    n1647_o2
  );


  not

  (
    n1647_o2_n,
    n1647_o2
  );


  buf

  (
    n1648_o2_p,
    n1648_o2
  );


  not

  (
    n1648_o2_n,
    n1648_o2
  );


  buf

  (
    n1649_o2_p,
    n1649_o2
  );


  not

  (
    n1649_o2_n,
    n1649_o2
  );


  buf

  (
    n1650_o2_p,
    n1650_o2
  );


  not

  (
    n1650_o2_n,
    n1650_o2
  );


  buf

  (
    n1651_o2_p,
    n1651_o2
  );


  not

  (
    n1651_o2_n,
    n1651_o2
  );


  buf

  (
    n1652_o2_p,
    n1652_o2
  );


  not

  (
    n1652_o2_n,
    n1652_o2
  );


  buf

  (
    n1653_o2_p,
    n1653_o2
  );


  not

  (
    n1653_o2_n,
    n1653_o2
  );


  buf

  (
    n1654_o2_p,
    n1654_o2
  );


  not

  (
    n1654_o2_n,
    n1654_o2
  );


  buf

  (
    n1655_o2_p,
    n1655_o2
  );


  not

  (
    n1655_o2_n,
    n1655_o2
  );


  buf

  (
    n1656_o2_p,
    n1656_o2
  );


  not

  (
    n1656_o2_n,
    n1656_o2
  );


  buf

  (
    n1657_o2_p,
    n1657_o2
  );


  not

  (
    n1657_o2_n,
    n1657_o2
  );


  buf

  (
    n1658_o2_p,
    n1658_o2
  );


  not

  (
    n1658_o2_n,
    n1658_o2
  );


  buf

  (
    n1659_o2_p,
    n1659_o2
  );


  not

  (
    n1659_o2_n,
    n1659_o2
  );


  buf

  (
    n1660_o2_p,
    n1660_o2
  );


  not

  (
    n1660_o2_n,
    n1660_o2
  );


  buf

  (
    n1661_o2_p,
    n1661_o2
  );


  not

  (
    n1661_o2_n,
    n1661_o2
  );


  buf

  (
    n1662_o2_p,
    n1662_o2
  );


  not

  (
    n1662_o2_n,
    n1662_o2
  );


  buf

  (
    n1663_o2_p,
    n1663_o2
  );


  not

  (
    n1663_o2_n,
    n1663_o2
  );


  buf

  (
    n1664_o2_p,
    n1664_o2
  );


  not

  (
    n1664_o2_n,
    n1664_o2
  );


  buf

  (
    n1665_o2_p,
    n1665_o2
  );


  not

  (
    n1665_o2_n,
    n1665_o2
  );


  buf

  (
    n1666_o2_p,
    n1666_o2
  );


  not

  (
    n1666_o2_n,
    n1666_o2
  );


  buf

  (
    n1667_o2_p,
    n1667_o2
  );


  not

  (
    n1667_o2_n,
    n1667_o2
  );


  buf

  (
    n1668_o2_p,
    n1668_o2
  );


  not

  (
    n1668_o2_n,
    n1668_o2
  );


  buf

  (
    n1669_o2_p,
    n1669_o2
  );


  not

  (
    n1669_o2_n,
    n1669_o2
  );


  buf

  (
    n1670_o2_p,
    n1670_o2
  );


  not

  (
    n1670_o2_n,
    n1670_o2
  );


  buf

  (
    n1671_o2_p,
    n1671_o2
  );


  not

  (
    n1671_o2_n,
    n1671_o2
  );


  buf

  (
    n1672_o2_p,
    n1672_o2
  );


  not

  (
    n1672_o2_n,
    n1672_o2
  );


  buf

  (
    n1673_o2_p,
    n1673_o2
  );


  not

  (
    n1673_o2_n,
    n1673_o2
  );


  buf

  (
    n1674_o2_p,
    n1674_o2
  );


  not

  (
    n1674_o2_n,
    n1674_o2
  );


  buf

  (
    n1675_o2_p,
    n1675_o2
  );


  not

  (
    n1675_o2_n,
    n1675_o2
  );


  buf

  (
    n685_o2_p,
    n685_o2
  );


  not

  (
    n685_o2_n,
    n685_o2
  );


  buf

  (
    n680_o2_p,
    n680_o2
  );


  not

  (
    n680_o2_n,
    n680_o2
  );


  buf

  (
    n822_o2_p,
    n822_o2
  );


  not

  (
    n822_o2_n,
    n822_o2
  );


  buf

  (
    n843_o2_p,
    n843_o2
  );


  not

  (
    n843_o2_n,
    n843_o2
  );


  buf

  (
    n842_o2_p,
    n842_o2
  );


  not

  (
    n842_o2_n,
    n842_o2
  );


  buf

  (
    n681_o2_p,
    n681_o2
  );


  not

  (
    n681_o2_n,
    n681_o2
  );


  buf

  (
    n684_o2_p,
    n684_o2
  );


  not

  (
    n684_o2_n,
    n684_o2
  );


  buf

  (
    n686_o2_p,
    n686_o2
  );


  not

  (
    n686_o2_n,
    n686_o2
  );


  buf

  (
    n823_o2_p,
    n823_o2
  );


  not

  (
    n823_o2_n,
    n823_o2
  );


  buf

  (
    n683_o2_p,
    n683_o2
  );


  not

  (
    n683_o2_n,
    n683_o2
  );


  buf

  (
    n688_o2_p,
    n688_o2
  );


  not

  (
    n688_o2_n,
    n688_o2
  );


  buf

  (
    n803_o2_p,
    n803_o2
  );


  not

  (
    n803_o2_n,
    n803_o2
  );


  buf

  (
    n862_o2_p,
    n862_o2
  );


  not

  (
    n862_o2_n,
    n862_o2
  );


  buf

  (
    n764_o2_p,
    n764_o2
  );


  not

  (
    n764_o2_n,
    n764_o2
  );


  buf

  (
    n863_o2_p,
    n863_o2
  );


  not

  (
    n863_o2_n,
    n863_o2
  );


  buf

  (
    n886_o2_p,
    n886_o2
  );


  not

  (
    n886_o2_n,
    n886_o2
  );


  buf

  (
    lo002_buf_o2_p,
    lo002_buf_o2
  );


  not

  (
    lo002_buf_o2_n,
    lo002_buf_o2
  );


  buf

  (
    lo006_buf_o2_p,
    lo006_buf_o2
  );


  not

  (
    lo006_buf_o2_n,
    lo006_buf_o2
  );


  buf

  (
    lo010_buf_o2_p,
    lo010_buf_o2
  );


  not

  (
    lo010_buf_o2_n,
    lo010_buf_o2
  );


  buf

  (
    lo014_buf_o2_p,
    lo014_buf_o2
  );


  not

  (
    lo014_buf_o2_n,
    lo014_buf_o2
  );


  buf

  (
    lo018_buf_o2_p,
    lo018_buf_o2
  );


  not

  (
    lo018_buf_o2_n,
    lo018_buf_o2
  );


  buf

  (
    lo022_buf_o2_p,
    lo022_buf_o2
  );


  not

  (
    lo022_buf_o2_n,
    lo022_buf_o2
  );


  buf

  (
    lo026_buf_o2_p,
    lo026_buf_o2
  );


  not

  (
    lo026_buf_o2_n,
    lo026_buf_o2
  );


  buf

  (
    lo030_buf_o2_p,
    lo030_buf_o2
  );


  not

  (
    lo030_buf_o2_n,
    lo030_buf_o2
  );


  buf

  (
    lo034_buf_o2_p,
    lo034_buf_o2
  );


  not

  (
    lo034_buf_o2_n,
    lo034_buf_o2
  );


  buf

  (
    lo038_buf_o2_p,
    lo038_buf_o2
  );


  not

  (
    lo038_buf_o2_n,
    lo038_buf_o2
  );


  buf

  (
    lo042_buf_o2_p,
    lo042_buf_o2
  );


  not

  (
    lo042_buf_o2_n,
    lo042_buf_o2
  );


  buf

  (
    lo046_buf_o2_p,
    lo046_buf_o2
  );


  not

  (
    lo046_buf_o2_n,
    lo046_buf_o2
  );


  buf

  (
    lo050_buf_o2_p,
    lo050_buf_o2
  );


  not

  (
    lo050_buf_o2_n,
    lo050_buf_o2
  );


  buf

  (
    lo054_buf_o2_p,
    lo054_buf_o2
  );


  not

  (
    lo054_buf_o2_n,
    lo054_buf_o2
  );


  buf

  (
    lo058_buf_o2_p,
    lo058_buf_o2
  );


  not

  (
    lo058_buf_o2_n,
    lo058_buf_o2
  );


  buf

  (
    lo062_buf_o2_p,
    lo062_buf_o2
  );


  not

  (
    lo062_buf_o2_n,
    lo062_buf_o2
  );


  buf

  (
    lo066_buf_o2_p,
    lo066_buf_o2
  );


  not

  (
    lo066_buf_o2_n,
    lo066_buf_o2
  );


  buf

  (
    lo070_buf_o2_p,
    lo070_buf_o2
  );


  not

  (
    lo070_buf_o2_n,
    lo070_buf_o2
  );


  buf

  (
    lo074_buf_o2_p,
    lo074_buf_o2
  );


  not

  (
    lo074_buf_o2_n,
    lo074_buf_o2
  );


  buf

  (
    lo078_buf_o2_p,
    lo078_buf_o2
  );


  not

  (
    lo078_buf_o2_n,
    lo078_buf_o2
  );


  buf

  (
    lo082_buf_o2_p,
    lo082_buf_o2
  );


  not

  (
    lo082_buf_o2_n,
    lo082_buf_o2
  );


  buf

  (
    lo086_buf_o2_p,
    lo086_buf_o2
  );


  not

  (
    lo086_buf_o2_n,
    lo086_buf_o2
  );


  buf

  (
    lo090_buf_o2_p,
    lo090_buf_o2
  );


  not

  (
    lo090_buf_o2_n,
    lo090_buf_o2
  );


  buf

  (
    lo094_buf_o2_p,
    lo094_buf_o2
  );


  not

  (
    lo094_buf_o2_n,
    lo094_buf_o2
  );


  buf

  (
    lo098_buf_o2_p,
    lo098_buf_o2
  );


  not

  (
    lo098_buf_o2_n,
    lo098_buf_o2
  );


  buf

  (
    lo102_buf_o2_p,
    lo102_buf_o2
  );


  not

  (
    lo102_buf_o2_n,
    lo102_buf_o2
  );


  buf

  (
    lo106_buf_o2_p,
    lo106_buf_o2
  );


  not

  (
    lo106_buf_o2_n,
    lo106_buf_o2
  );


  buf

  (
    lo110_buf_o2_p,
    lo110_buf_o2
  );


  not

  (
    lo110_buf_o2_n,
    lo110_buf_o2
  );


  buf

  (
    lo114_buf_o2_p,
    lo114_buf_o2
  );


  not

  (
    lo114_buf_o2_n,
    lo114_buf_o2
  );


  buf

  (
    lo118_buf_o2_p,
    lo118_buf_o2
  );


  not

  (
    lo118_buf_o2_n,
    lo118_buf_o2
  );


  buf

  (
    lo122_buf_o2_p,
    lo122_buf_o2
  );


  not

  (
    lo122_buf_o2_n,
    lo122_buf_o2
  );


  buf

  (
    lo126_buf_o2_p,
    lo126_buf_o2
  );


  not

  (
    lo126_buf_o2_n,
    lo126_buf_o2
  );


  buf

  (
    n600_o2_p,
    n600_o2
  );


  not

  (
    n600_o2_n,
    n600_o2
  );


  buf

  (
    n601_o2_p,
    n601_o2
  );


  not

  (
    n601_o2_n,
    n601_o2
  );


  buf

  (
    n637_o2_p,
    n637_o2
  );


  not

  (
    n637_o2_n,
    n637_o2
  );


  buf

  (
    n638_o2_p,
    n638_o2
  );


  not

  (
    n638_o2_n,
    n638_o2
  );


  buf

  (
    n676_o2_p,
    n676_o2
  );


  not

  (
    n676_o2_n,
    n676_o2
  );


  buf

  (
    n677_o2_p,
    n677_o2
  );


  not

  (
    n677_o2_n,
    n677_o2
  );


  buf

  (
    n656_o2_p,
    n656_o2
  );


  not

  (
    n656_o2_n,
    n656_o2
  );


  buf

  (
    n657_o2_p,
    n657_o2
  );


  not

  (
    n657_o2_n,
    n657_o2
  );


  buf

  (
    n781_o2_p,
    n781_o2
  );


  not

  (
    n781_o2_n,
    n781_o2
  );


  buf

  (
    n782_o2_p,
    n782_o2
  );


  not

  (
    n782_o2_n,
    n782_o2
  );


  buf

  (
    n800_o2_p,
    n800_o2
  );


  not

  (
    n800_o2_n,
    n800_o2
  );


  buf

  (
    n801_o2_p,
    n801_o2
  );


  not

  (
    n801_o2_n,
    n801_o2
  );


  buf

  (
    n724_o2_p,
    n724_o2
  );


  not

  (
    n724_o2_n,
    n724_o2
  );


  buf

  (
    n725_o2_p,
    n725_o2
  );


  not

  (
    n725_o2_n,
    n725_o2
  );


  buf

  (
    n761_o2_p,
    n761_o2
  );


  not

  (
    n761_o2_n,
    n761_o2
  );


  buf

  (
    n762_o2_p,
    n762_o2
  );


  not

  (
    n762_o2_n,
    n762_o2
  );


  buf

  (
    lo129_buf_o2_p,
    lo129_buf_o2
  );


  not

  (
    lo129_buf_o2_n,
    lo129_buf_o2
  );


  buf

  (
    lo133_buf_o2_p,
    lo133_buf_o2
  );


  not

  (
    lo133_buf_o2_n,
    lo133_buf_o2
  );


  buf

  (
    lo137_buf_o2_p,
    lo137_buf_o2
  );


  not

  (
    lo137_buf_o2_n,
    lo137_buf_o2
  );


  buf

  (
    lo141_buf_o2_p,
    lo141_buf_o2
  );


  not

  (
    lo141_buf_o2_n,
    lo141_buf_o2
  );


  buf

  (
    lo145_buf_o2_p,
    lo145_buf_o2
  );


  not

  (
    lo145_buf_o2_n,
    lo145_buf_o2
  );


  buf

  (
    lo149_buf_o2_p,
    lo149_buf_o2
  );


  not

  (
    lo149_buf_o2_n,
    lo149_buf_o2
  );


  buf

  (
    lo153_buf_o2_p,
    lo153_buf_o2
  );


  not

  (
    lo153_buf_o2_n,
    lo153_buf_o2
  );


  buf

  (
    lo157_buf_o2_p,
    lo157_buf_o2
  );


  not

  (
    lo157_buf_o2_n,
    lo157_buf_o2
  );


  buf

  (
    lo161_buf_o2_p,
    lo161_buf_o2
  );


  not

  (
    lo161_buf_o2_n,
    lo161_buf_o2
  );


  buf

  (
    n571_o2_p,
    n571_o2
  );


  not

  (
    n571_o2_n,
    n571_o2
  );


  buf

  (
    n708_o2_p,
    n708_o2
  );


  not

  (
    n708_o2_n,
    n708_o2
  );


  buf

  (
    n608_o2_p,
    n608_o2
  );


  not

  (
    n608_o2_n,
    n608_o2
  );


  buf

  (
    n665_o2_p,
    n665_o2
  );


  not

  (
    n665_o2_n,
    n665_o2
  );


  buf

  (
    n705_o2_p,
    n705_o2
  );


  not

  (
    n705_o2_n,
    n705_o2
  );


  buf

  (
    n645_o2_p,
    n645_o2
  );


  not

  (
    n645_o2_n,
    n645_o2
  );


  buf

  (
    n745_o2_p,
    n745_o2
  );


  not

  (
    n745_o2_n,
    n745_o2
  );


  buf

  (
    n742_o2_p,
    n742_o2
  );


  not

  (
    n742_o2_n,
    n742_o2
  );


  buf

  (
    n568_o2_p,
    n568_o2
  );


  not

  (
    n568_o2_n,
    n568_o2
  );


  buf

  (
    n717_o2_p,
    n717_o2
  );


  not

  (
    n717_o2_n,
    n717_o2
  );


  buf

  (
    n605_o2_p,
    n605_o2
  );


  not

  (
    n605_o2_n,
    n605_o2
  );


  buf

  (
    n662_o2_p,
    n662_o2
  );


  not

  (
    n662_o2_n,
    n662_o2
  );


  buf

  (
    n714_o2_p,
    n714_o2
  );


  not

  (
    n714_o2_n,
    n714_o2
  );


  buf

  (
    n642_o2_p,
    n642_o2
  );


  not

  (
    n642_o2_n,
    n642_o2
  );


  buf

  (
    n754_o2_p,
    n754_o2
  );


  not

  (
    n754_o2_n,
    n754_o2
  );


  buf

  (
    n751_o2_p,
    n751_o2
  );


  not

  (
    n751_o2_n,
    n751_o2
  );


  buf

  (
    n584_o2_p,
    n584_o2
  );


  not

  (
    n584_o2_n,
    n584_o2
  );


  buf

  (
    n770_o2_p,
    n770_o2
  );


  not

  (
    n770_o2_n,
    n770_o2
  );


  buf

  (
    n789_o2_p,
    n789_o2
  );


  not

  (
    n789_o2_n,
    n789_o2
  );


  buf

  (
    n581_o2_p,
    n581_o2
  );


  not

  (
    n581_o2_n,
    n581_o2
  );


  buf

  (
    n695_o2_p,
    n695_o2
  );


  not

  (
    n695_o2_n,
    n695_o2
  );


  buf

  (
    n732_o2_p,
    n732_o2
  );


  not

  (
    n732_o2_n,
    n732_o2
  );


  buf

  (
    n593_o2_p,
    n593_o2
  );


  not

  (
    n593_o2_n,
    n593_o2
  );


  buf

  (
    n590_o2_p,
    n590_o2
  );


  not

  (
    n590_o2_n,
    n590_o2
  );


  buf

  (
    n630_o2_p,
    n630_o2
  );


  not

  (
    n630_o2_n,
    n630_o2
  );


  buf

  (
    n767_o2_p,
    n767_o2
  );


  not

  (
    n767_o2_n,
    n767_o2
  );


  buf

  (
    n786_o2_p,
    n786_o2
  );


  not

  (
    n786_o2_n,
    n786_o2
  );


  buf

  (
    n627_o2_p,
    n627_o2
  );


  not

  (
    n627_o2_n,
    n627_o2
  );


  buf

  (
    n692_o2_p,
    n692_o2
  );


  not

  (
    n692_o2_n,
    n692_o2
  );


  buf

  (
    n729_o2_p,
    n729_o2
  );


  not

  (
    n729_o2_n,
    n729_o2
  );


  buf

  (
    n621_o2_p,
    n621_o2
  );


  not

  (
    n621_o2_n,
    n621_o2
  );


  buf

  (
    n618_o2_p,
    n618_o2
  );


  not

  (
    n618_o2_n,
    n618_o2
  );


  and

  (
    g260_p,
    n683_o2_n,
    n688_o2_n
  );


  or

  (
    g260_n,
    n683_o2_p,
    n688_o2_p
  );


  and

  (
    g261_p,
    n803_o2_p,
    n764_o2_p
  );


  or

  (
    g261_n,
    n803_o2_n,
    n764_o2_n
  );


  and

  (
    g262_p,
    g260_n_spl_0,
    g261_p
  );


  or

  (
    g262_n,
    g260_p_spl_0,
    g261_n
  );


  and

  (
    g263_p,
    n602_o2_p_spl_0,
    g262_p_spl_0
  );


  or

  (
    g263_n,
    n602_o2_n_spl_0,
    g262_n_spl_0
  );


  or

  (
    g264_n,
    n630_lo_n,
    g263_p
  );


  or

  (
    g265_n,
    n630_lo_p,
    g263_n
  );


  and

  (
    g266_p,
    g264_n,
    g265_n
  );


  and

  (
    g267_p,
    n639_o2_p_spl_00,
    g262_p_spl_0
  );


  or

  (
    g267_n,
    n639_o2_n_spl_00,
    g262_n_spl_0
  );


  or

  (
    g268_n,
    n642_lo_n,
    g267_p
  );


  or

  (
    g269_n,
    n642_lo_p,
    g267_n
  );


  and

  (
    g270_p,
    g268_n,
    g269_n
  );


  and

  (
    g271_p,
    n678_o2_p_spl_00,
    g262_p_spl_1
  );


  or

  (
    g271_n,
    n678_o2_n_spl_00,
    g262_n_spl_1
  );


  or

  (
    g272_n,
    n654_lo_n,
    g271_p
  );


  or

  (
    g273_n,
    n654_lo_p,
    g271_n
  );


  and

  (
    g274_p,
    g272_n,
    g273_n
  );


  and

  (
    g275_p,
    n658_o2_p_spl_0,
    g262_p_spl_1
  );


  or

  (
    g275_n,
    n658_o2_n_spl_0,
    g262_n_spl_1
  );


  or

  (
    g276_n,
    n666_lo_n,
    g275_p
  );


  or

  (
    g277_n,
    n666_lo_p,
    g275_n
  );


  and

  (
    g278_p,
    g276_n,
    g277_n
  );


  and

  (
    g279_p,
    n822_o2_p,
    n823_o2_n
  );


  or

  (
    g279_n,
    n822_o2_n,
    n823_o2_p
  );


  and

  (
    g280_p,
    g260_n_spl_0,
    g279_p
  );


  or

  (
    g280_n,
    g260_p_spl_0,
    g279_n
  );


  and

  (
    g281_p,
    n602_o2_p_spl_0,
    g280_p_spl_0
  );


  or

  (
    g281_n,
    n602_o2_n_spl_0,
    g280_n_spl_0
  );


  or

  (
    g282_n,
    n678_lo_n,
    g281_p
  );


  or

  (
    g283_n,
    n678_lo_p,
    g281_n
  );


  and

  (
    g284_p,
    g282_n,
    g283_n
  );


  and

  (
    g285_p,
    n639_o2_p_spl_00,
    g280_p_spl_0
  );


  or

  (
    g285_n,
    n639_o2_n_spl_00,
    g280_n_spl_0
  );


  or

  (
    g286_n,
    n690_lo_n,
    g285_p
  );


  or

  (
    g287_n,
    n690_lo_p,
    g285_n
  );


  and

  (
    g288_p,
    g286_n,
    g287_n
  );


  and

  (
    g289_p,
    n678_o2_p_spl_00,
    g280_p_spl_1
  );


  or

  (
    g289_n,
    n678_o2_n_spl_00,
    g280_n_spl_1
  );


  or

  (
    g290_n,
    n702_lo_n,
    g289_p
  );


  or

  (
    g291_n,
    n702_lo_p,
    g289_n
  );


  and

  (
    g292_p,
    g290_n,
    g291_n
  );


  and

  (
    g293_p,
    n658_o2_p_spl_0,
    g280_p_spl_1
  );


  or

  (
    g293_n,
    n658_o2_n_spl_0,
    g280_n_spl_1
  );


  or

  (
    g294_n,
    n714_lo_n,
    g293_p
  );


  or

  (
    g295_n,
    n714_lo_p,
    g293_n
  );


  and

  (
    g296_p,
    g294_n,
    g295_n
  );


  and

  (
    g297_p,
    n843_o2_n,
    n842_o2_p
  );


  or

  (
    g297_n,
    n843_o2_p,
    n842_o2_n
  );


  and

  (
    g298_p,
    g260_n_spl_1,
    g297_p
  );


  or

  (
    g298_n,
    g260_p_spl_1,
    g297_n
  );


  and

  (
    g299_p,
    n602_o2_p_spl_1,
    g298_p_spl_0
  );


  or

  (
    g299_n,
    n602_o2_n_spl_1,
    g298_n_spl_0
  );


  or

  (
    g300_n,
    n726_lo_n,
    g299_p
  );


  or

  (
    g301_n,
    n726_lo_p,
    g299_n
  );


  and

  (
    g302_p,
    g300_n,
    g301_n
  );


  and

  (
    g303_p,
    n639_o2_p_spl_0,
    g298_p_spl_0
  );


  or

  (
    g303_n,
    n639_o2_n_spl_0,
    g298_n_spl_0
  );


  or

  (
    g304_n,
    n738_lo_n,
    g303_p
  );


  or

  (
    g305_n,
    n738_lo_p,
    g303_n
  );


  and

  (
    g306_p,
    g304_n,
    g305_n
  );


  and

  (
    g307_p,
    n678_o2_p_spl_01,
    g298_p_spl_1
  );


  or

  (
    g307_n,
    n678_o2_n_spl_01,
    g298_n_spl_1
  );


  or

  (
    g308_n,
    n750_lo_n,
    g307_p
  );


  or

  (
    g309_n,
    n750_lo_p,
    g307_n
  );


  and

  (
    g310_p,
    g308_n,
    g309_n
  );


  and

  (
    g311_p,
    n658_o2_p_spl_1,
    g298_p_spl_1
  );


  or

  (
    g311_n,
    n658_o2_n_spl_1,
    g298_n_spl_1
  );


  or

  (
    g312_n,
    n762_lo_n,
    g311_p
  );


  or

  (
    g313_n,
    n762_lo_p,
    g311_n
  );


  and

  (
    g314_p,
    g312_n,
    g313_n
  );


  and

  (
    g315_p,
    n862_o2_p,
    n863_o2_p
  );


  or

  (
    g315_n,
    n862_o2_n,
    n863_o2_n
  );


  and

  (
    g316_p,
    g260_n_spl_1,
    g315_p
  );


  or

  (
    g316_n,
    g260_p_spl_1,
    g315_n
  );


  and

  (
    g317_p,
    n602_o2_p_spl_1,
    g316_p_spl_0
  );


  or

  (
    g317_n,
    n602_o2_n_spl_1,
    g316_n_spl_0
  );


  or

  (
    g318_n,
    n774_lo_n,
    g317_p
  );


  or

  (
    g319_n,
    n774_lo_p,
    g317_n
  );


  and

  (
    g320_p,
    g318_n,
    g319_n
  );


  and

  (
    g321_p,
    n639_o2_p_spl_1,
    g316_p_spl_0
  );


  or

  (
    g321_n,
    n639_o2_n_spl_1,
    g316_n_spl_0
  );


  or

  (
    g322_n,
    n786_lo_n,
    g321_p
  );


  or

  (
    g323_n,
    n786_lo_p,
    g321_n
  );


  and

  (
    g324_p,
    g322_n,
    g323_n
  );


  and

  (
    g325_p,
    n678_o2_p_spl_01,
    g316_p_spl_1
  );


  or

  (
    g325_n,
    n678_o2_n_spl_01,
    g316_n_spl_1
  );


  or

  (
    g326_n,
    n798_lo_n,
    g325_p
  );


  or

  (
    g327_n,
    n798_lo_p,
    g325_n
  );


  and

  (
    g328_p,
    g326_n,
    g327_n
  );


  and

  (
    g329_p,
    n658_o2_p_spl_1,
    g316_p_spl_1
  );


  or

  (
    g329_n,
    n658_o2_n_spl_1,
    g316_n_spl_1
  );


  or

  (
    g330_n,
    n810_lo_n,
    g329_p
  );


  or

  (
    g331_n,
    n810_lo_p,
    g329_n
  );


  and

  (
    g332_p,
    g330_n,
    g331_n
  );


  and

  (
    g333_p,
    n686_o2_p,
    n886_o2_p_spl_0
  );


  or

  (
    g333_n,
    n686_o2_n,
    n886_o2_n_spl_0
  );


  and

  (
    g334_p,
    n678_o2_p_spl_1,
    g333_p
  );


  or

  (
    g334_n,
    n678_o2_n_spl_1,
    g333_n
  );


  and

  (
    g335_p,
    n783_o2_p_spl_0,
    g334_p_spl_0
  );


  or

  (
    g335_n,
    n783_o2_n_spl_0,
    g334_n_spl_0
  );


  or

  (
    g336_n,
    n822_lo_n,
    g335_p
  );


  or

  (
    g337_n,
    n822_lo_p,
    g335_n
  );


  and

  (
    g338_p,
    g336_n,
    g337_n
  );


  and

  (
    g339_p,
    n802_o2_p_spl_0,
    g334_p_spl_0
  );


  or

  (
    g339_n,
    n802_o2_n_spl_0,
    g334_n_spl_0
  );


  or

  (
    g340_n,
    n834_lo_n,
    g339_p
  );


  or

  (
    g341_n,
    n834_lo_p,
    g339_n
  );


  and

  (
    g342_p,
    g340_n,
    g341_n
  );


  and

  (
    g343_p,
    n726_o2_p_spl_0,
    g334_p_spl_1
  );


  or

  (
    g343_n,
    n726_o2_n_spl_0,
    g334_n_spl_1
  );


  or

  (
    g344_n,
    n846_lo_n,
    g343_p
  );


  or

  (
    g345_n,
    n846_lo_p,
    g343_n
  );


  and

  (
    g346_p,
    g344_n,
    g345_n
  );


  and

  (
    g347_p,
    n763_o2_p_spl_0,
    g334_p_spl_1
  );


  or

  (
    g347_n,
    n763_o2_n_spl_0,
    g334_n_spl_1
  );


  or

  (
    g348_n,
    n858_lo_n,
    g347_p
  );


  or

  (
    g349_n,
    n858_lo_p,
    g347_n
  );


  and

  (
    g350_p,
    g348_n,
    g349_n
  );


  and

  (
    g351_p,
    n685_o2_p,
    n680_o2_p
  );


  or

  (
    g351_n,
    n685_o2_n,
    n680_o2_n
  );


  and

  (
    g352_p,
    n886_o2_p_spl_0,
    g351_p
  );


  or

  (
    g352_n,
    n886_o2_n_spl_0,
    g351_n
  );


  and

  (
    g353_p,
    n783_o2_p_spl_0,
    g352_p_spl_0
  );


  or

  (
    g353_n,
    n783_o2_n_spl_0,
    g352_n_spl_0
  );


  or

  (
    g354_n,
    n870_lo_n,
    g353_p
  );


  or

  (
    g355_n,
    n870_lo_p,
    g353_n
  );


  and

  (
    g356_p,
    g354_n,
    g355_n
  );


  and

  (
    g357_p,
    n802_o2_p_spl_0,
    g352_p_spl_0
  );


  or

  (
    g357_n,
    n802_o2_n_spl_0,
    g352_n_spl_0
  );


  or

  (
    g358_n,
    n882_lo_n,
    g357_p
  );


  or

  (
    g359_n,
    n882_lo_p,
    g357_n
  );


  and

  (
    g360_p,
    g358_n,
    g359_n
  );


  and

  (
    g361_p,
    n726_o2_p_spl_0,
    g352_p_spl_1
  );


  or

  (
    g361_n,
    n726_o2_n_spl_0,
    g352_n_spl_1
  );


  or

  (
    g362_n,
    n894_lo_n,
    g361_p
  );


  or

  (
    g363_n,
    n894_lo_p,
    g361_n
  );


  and

  (
    g364_p,
    g362_n,
    g363_n
  );


  and

  (
    g365_p,
    n763_o2_p_spl_0,
    g352_p_spl_1
  );


  or

  (
    g365_n,
    n763_o2_n_spl_0,
    g352_n_spl_1
  );


  or

  (
    g366_n,
    n906_lo_n,
    g365_p
  );


  or

  (
    g367_n,
    n906_lo_p,
    g365_n
  );


  and

  (
    g368_p,
    g366_n,
    g367_n
  );


  and

  (
    g369_p,
    n678_o2_p_spl_1,
    n684_o2_p
  );


  or

  (
    g369_n,
    n678_o2_n_spl_1,
    n684_o2_n
  );


  and

  (
    g370_p,
    n886_o2_p_spl_1,
    g369_p
  );


  or

  (
    g370_n,
    n886_o2_n_spl_1,
    g369_n
  );


  and

  (
    g371_p,
    n783_o2_p_spl_1,
    g370_p_spl_0
  );


  or

  (
    g371_n,
    n783_o2_n_spl_1,
    g370_n_spl_0
  );


  or

  (
    g372_n,
    n918_lo_n,
    g371_p
  );


  or

  (
    g373_n,
    n918_lo_p,
    g371_n
  );


  and

  (
    g374_p,
    g372_n,
    g373_n
  );


  and

  (
    g375_p,
    n802_o2_p_spl_1,
    g370_p_spl_0
  );


  or

  (
    g375_n,
    n802_o2_n_spl_1,
    g370_n_spl_0
  );


  or

  (
    g376_n,
    n930_lo_n,
    g375_p
  );


  or

  (
    g377_n,
    n930_lo_p,
    g375_n
  );


  and

  (
    g378_p,
    g376_n,
    g377_n
  );


  and

  (
    g379_p,
    n726_o2_p_spl_1,
    g370_p_spl_1
  );


  or

  (
    g379_n,
    n726_o2_n_spl_1,
    g370_n_spl_1
  );


  or

  (
    g380_n,
    n942_lo_n,
    g379_p
  );


  or

  (
    g381_n,
    n942_lo_p,
    g379_n
  );


  and

  (
    g382_p,
    g380_n,
    g381_n
  );


  and

  (
    g383_p,
    n763_o2_p_spl_1,
    g370_p_spl_1
  );


  or

  (
    g383_n,
    n763_o2_n_spl_1,
    g370_n_spl_1
  );


  or

  (
    g384_n,
    n954_lo_n,
    g383_p
  );


  or

  (
    g385_n,
    n954_lo_p,
    g383_n
  );


  and

  (
    g386_p,
    g384_n,
    g385_n
  );


  and

  (
    g387_p,
    n639_o2_p_spl_1,
    n681_o2_p
  );


  or

  (
    g387_n,
    n639_o2_n_spl_1,
    n681_o2_n
  );


  and

  (
    g388_p,
    n886_o2_p_spl_1,
    g387_p
  );


  or

  (
    g388_n,
    n886_o2_n_spl_1,
    g387_n
  );


  and

  (
    g389_p,
    n783_o2_p_spl_1,
    g388_p_spl_0
  );


  or

  (
    g389_n,
    n783_o2_n_spl_1,
    g388_n_spl_0
  );


  or

  (
    g390_n,
    n966_lo_n,
    g389_p
  );


  or

  (
    g391_n,
    n966_lo_p,
    g389_n
  );


  and

  (
    g392_p,
    g390_n,
    g391_n
  );


  and

  (
    g393_p,
    n802_o2_p_spl_1,
    g388_p_spl_0
  );


  or

  (
    g393_n,
    n802_o2_n_spl_1,
    g388_n_spl_0
  );


  or

  (
    g394_n,
    n978_lo_n,
    g393_p
  );


  or

  (
    g395_n,
    n978_lo_p,
    g393_n
  );


  and

  (
    g396_p,
    g394_n,
    g395_n
  );


  and

  (
    g397_p,
    n726_o2_p_spl_1,
    g388_p_spl_1
  );


  or

  (
    g397_n,
    n726_o2_n_spl_1,
    g388_n_spl_1
  );


  or

  (
    g398_n,
    n990_lo_n,
    g397_p
  );


  or

  (
    g399_n,
    n990_lo_p,
    g397_n
  );


  and

  (
    g400_p,
    g398_n,
    g399_n
  );


  and

  (
    g401_p,
    n763_o2_p_spl_1,
    g388_p_spl_1
  );


  or

  (
    g401_n,
    n763_o2_n_spl_1,
    g388_n_spl_1
  );


  or

  (
    g402_n,
    n1002_lo_n,
    g401_p
  );


  or

  (
    g403_n,
    n1002_lo_p,
    g401_n
  );


  and

  (
    g404_p,
    g402_n,
    g403_n
  );


  and

  (
    g405_p,
    n600_o2_n,
    n601_o2_n
  );


  or

  (
    g405_n,
    n600_o2_p,
    n601_o2_p
  );


  and

  (
    g406_p,
    n637_o2_n,
    n638_o2_n
  );


  or

  (
    g406_n,
    n637_o2_p,
    n638_o2_p
  );


  and

  (
    g407_p,
    n676_o2_n,
    n677_o2_n
  );


  or

  (
    g407_n,
    n676_o2_p,
    n677_o2_p
  );


  and

  (
    g408_p,
    n656_o2_n,
    n657_o2_n
  );


  or

  (
    g408_n,
    n656_o2_p,
    n657_o2_p
  );


  and

  (
    g409_p,
    n781_o2_n,
    n782_o2_n
  );


  or

  (
    g409_n,
    n781_o2_p,
    n782_o2_p
  );


  and

  (
    g410_p,
    n800_o2_n,
    n801_o2_n
  );


  or

  (
    g410_n,
    n800_o2_p,
    n801_o2_p
  );


  and

  (
    g411_p,
    n724_o2_n,
    n725_o2_n
  );


  or

  (
    g411_n,
    n724_o2_p,
    n725_o2_p
  );


  and

  (
    g412_p,
    n761_o2_n,
    n762_o2_n
  );


  or

  (
    g412_n,
    n761_o2_p,
    n762_o2_p
  );


  or

  (
    g413_n,
    g405_p,
    g406_n_spl_0
  );


  or

  (
    g414_n,
    g407_n_spl_0,
    g408_p
  );


  or

  (
    g415_n,
    g409_p_spl_0,
    g412_p_spl_0
  );


  and

  (
    g416_p,
    g409_p_spl_0,
    g412_p_spl_0
  );


  or

  (
    g416_n,
    g409_n_spl_0,
    g412_n_spl_0
  );


  or

  (
    g417_n,
    g410_p_spl_0,
    g411_p_spl_0
  );


  or

  (
    g418_n,
    g405_n_spl_0,
    g414_n_spl_
  );


  or

  (
    g419_n,
    g405_n_spl_0,
    g408_n_spl_0
  );


  or

  (
    g420_n,
    g406_p,
    g419_n_spl_
  );


  or

  (
    g421_n,
    g408_n_spl_0,
    g413_n_spl_
  );


  and

  (
    g422_p,
    g410_p_spl_0,
    g411_p_spl_0
  );


  or

  (
    g422_n,
    g410_n_spl_0,
    g411_n_spl_0
  );


  or

  (
    g423_n,
    g407_p,
    g419_n_spl_
  );


  and

  (
    g424_p,
    g418_n_spl_,
    g423_n
  );


  or

  (
    g425_n,
    g406_n_spl_0,
    g424_p
  );


  and

  (
    g426_p,
    g420_n_spl_,
    g421_n_spl_
  );


  or

  (
    g427_n,
    g407_n_spl_0,
    g426_p
  );


  and

  (
    g428_p,
    g409_n_spl_0,
    g410_p_spl_
  );


  and

  (
    g429_p,
    g409_p_spl_,
    g410_n_spl_0
  );


  and

  (
    g430_p,
    g411_n_spl_0,
    g412_p_spl_
  );


  and

  (
    g431_p,
    g411_p_spl_,
    g412_n_spl_0
  );


  and

  (
    g432_p,
    g415_n_spl_,
    g416_n_spl_
  );


  or

  (
    g433_n,
    g422_n_spl_,
    g432_p
  );


  and

  (
    g434_p,
    g416_p,
    g417_n_spl_
  );


  or

  (
    g435_n,
    g422_p,
    g434_p
  );


  and

  (
    g436_p,
    g433_n,
    g435_n
  );


  and

  (
    g437_p,
    n571_o2_p_spl_,
    n568_o2_n_spl_
  );


  or

  (
    g437_n,
    n571_o2_n_spl_,
    n568_o2_p_spl_
  );


  and

  (
    g438_p,
    n571_o2_n_spl_,
    n568_o2_p_spl_
  );


  or

  (
    g438_n,
    n571_o2_p_spl_,
    n568_o2_n_spl_
  );


  and

  (
    g439_p,
    g437_n,
    g438_n
  );


  or

  (
    g439_n,
    g437_p,
    g438_p
  );


  and

  (
    g440_p,
    lo129_buf_o2_p,
    lo161_buf_o2_p_spl_00
  );


  or

  (
    g440_n,
    lo129_buf_o2_n,
    lo161_buf_o2_n_spl_00
  );


  and

  (
    g441_p,
    g439_n,
    g440_p
  );


  and

  (
    g442_p,
    g439_p,
    g440_n
  );


  or

  (
    g443_n,
    g441_p,
    g442_p
  );


  and

  (
    g444_p,
    n584_o2_p_spl_,
    n581_o2_n_spl_
  );


  or

  (
    g444_n,
    n584_o2_n_spl_,
    n581_o2_p_spl_
  );


  and

  (
    g445_p,
    n584_o2_n_spl_,
    n581_o2_p_spl_
  );


  or

  (
    g445_n,
    n584_o2_p_spl_,
    n581_o2_n_spl_
  );


  and

  (
    g446_p,
    g444_n,
    g445_n
  );


  or

  (
    g446_n,
    g444_p,
    g445_p
  );


  and

  (
    g447_p,
    n593_o2_p_spl_,
    n590_o2_n_spl_
  );


  or

  (
    g447_n,
    n593_o2_n_spl_,
    n590_o2_p_spl_
  );


  and

  (
    g448_p,
    n593_o2_n_spl_,
    n590_o2_p_spl_
  );


  or

  (
    g448_n,
    n593_o2_p_spl_,
    n590_o2_n_spl_
  );


  and

  (
    g449_p,
    g447_n,
    g448_n
  );


  or

  (
    g449_n,
    g447_p,
    g448_p
  );


  and

  (
    g450_p,
    g446_p_spl_,
    g449_n_spl_
  );


  and

  (
    g451_p,
    g446_n_spl_,
    g449_p_spl_
  );


  or

  (
    g452_n,
    g450_p,
    g451_p
  );


  and

  (
    g453_p,
    g443_n_spl_,
    g452_n_spl_
  );


  or

  (
    g454_n,
    g443_n_spl_,
    g452_n_spl_
  );


  and

  (
    g455_p,
    n608_o2_p_spl_,
    n605_o2_n_spl_
  );


  or

  (
    g455_n,
    n608_o2_n_spl_,
    n605_o2_p_spl_
  );


  and

  (
    g456_p,
    n608_o2_n_spl_,
    n605_o2_p_spl_
  );


  or

  (
    g456_n,
    n608_o2_p_spl_,
    n605_o2_n_spl_
  );


  and

  (
    g457_p,
    g455_n,
    g456_n
  );


  or

  (
    g457_n,
    g455_p,
    g456_p
  );


  and

  (
    g458_p,
    lo133_buf_o2_p,
    lo161_buf_o2_p_spl_00
  );


  or

  (
    g458_n,
    lo133_buf_o2_n,
    lo161_buf_o2_n_spl_00
  );


  and

  (
    g459_p,
    g457_n,
    g458_p
  );


  and

  (
    g460_p,
    g457_p,
    g458_n
  );


  or

  (
    g461_n,
    g459_p,
    g460_p
  );


  and

  (
    g462_p,
    n621_o2_p_spl_,
    n618_o2_n_spl_
  );


  or

  (
    g462_n,
    n621_o2_n_spl_,
    n618_o2_p_spl_
  );


  and

  (
    g463_p,
    n621_o2_n_spl_,
    n618_o2_p_spl_
  );


  or

  (
    g463_n,
    n621_o2_p_spl_,
    n618_o2_n_spl_
  );


  and

  (
    g464_p,
    g462_n,
    g463_n
  );


  or

  (
    g464_n,
    g462_p,
    g463_p
  );


  and

  (
    g465_p,
    n630_o2_p_spl_,
    n627_o2_n_spl_
  );


  or

  (
    g465_n,
    n630_o2_n_spl_,
    n627_o2_p_spl_
  );


  and

  (
    g466_p,
    n630_o2_n_spl_,
    n627_o2_p_spl_
  );


  or

  (
    g466_n,
    n630_o2_p_spl_,
    n627_o2_n_spl_
  );


  and

  (
    g467_p,
    g465_n,
    g466_n
  );


  or

  (
    g467_n,
    g465_p,
    g466_p
  );


  and

  (
    g468_p,
    g464_p_spl_,
    g467_n_spl_
  );


  and

  (
    g469_p,
    g464_n_spl_,
    g467_p_spl_
  );


  or

  (
    g470_n,
    g468_p,
    g469_p
  );


  and

  (
    g471_p,
    g461_n_spl_,
    g470_n_spl_
  );


  or

  (
    g472_n,
    g461_n_spl_,
    g470_n_spl_
  );


  and

  (
    g473_p,
    n665_o2_p_spl_,
    n662_o2_n_spl_
  );


  or

  (
    g473_n,
    n665_o2_n_spl_,
    n662_o2_p_spl_
  );


  and

  (
    g474_p,
    n665_o2_n_spl_,
    n662_o2_p_spl_
  );


  or

  (
    g474_n,
    n665_o2_p_spl_,
    n662_o2_n_spl_
  );


  and

  (
    g475_p,
    g473_n,
    g474_n
  );


  or

  (
    g475_n,
    g473_p,
    g474_p
  );


  and

  (
    g476_p,
    lo137_buf_o2_p,
    lo161_buf_o2_p_spl_01
  );


  or

  (
    g476_n,
    lo137_buf_o2_n,
    lo161_buf_o2_n_spl_01
  );


  and

  (
    g477_p,
    g475_n,
    g476_p
  );


  and

  (
    g478_p,
    g475_p,
    g476_n
  );


  or

  (
    g479_n,
    g477_p,
    g478_p
  );


  and

  (
    g480_p,
    g446_p_spl_,
    g467_n_spl_
  );


  and

  (
    g481_p,
    g446_n_spl_,
    g467_p_spl_
  );


  or

  (
    g482_n,
    g480_p,
    g481_p
  );


  and

  (
    g483_p,
    g479_n_spl_,
    g482_n_spl_
  );


  or

  (
    g484_n,
    g479_n_spl_,
    g482_n_spl_
  );


  and

  (
    g485_p,
    n645_o2_p_spl_,
    n642_o2_n_spl_
  );


  or

  (
    g485_n,
    n645_o2_n_spl_,
    n642_o2_p_spl_
  );


  and

  (
    g486_p,
    n645_o2_n_spl_,
    n642_o2_p_spl_
  );


  or

  (
    g486_n,
    n645_o2_p_spl_,
    n642_o2_n_spl_
  );


  and

  (
    g487_p,
    g485_n,
    g486_n
  );


  or

  (
    g487_n,
    g485_p,
    g486_p
  );


  and

  (
    g488_p,
    lo141_buf_o2_p,
    lo161_buf_o2_p_spl_01
  );


  or

  (
    g488_n,
    lo141_buf_o2_n,
    lo161_buf_o2_n_spl_01
  );


  and

  (
    g489_p,
    g487_n,
    g488_p
  );


  and

  (
    g490_p,
    g487_p,
    g488_n
  );


  or

  (
    g491_n,
    g489_p,
    g490_p
  );


  and

  (
    g492_p,
    g449_p_spl_,
    g464_n_spl_
  );


  and

  (
    g493_p,
    g449_n_spl_,
    g464_p_spl_
  );


  or

  (
    g494_n,
    g492_p,
    g493_p
  );


  and

  (
    g495_p,
    g491_n_spl_,
    g494_n_spl_
  );


  or

  (
    g496_n,
    g491_n_spl_,
    g494_n_spl_
  );


  and

  (
    g497_p,
    n770_o2_p_spl_,
    n767_o2_n_spl_
  );


  or

  (
    g497_n,
    n770_o2_n_spl_,
    n767_o2_p_spl_
  );


  and

  (
    g498_p,
    n770_o2_n_spl_,
    n767_o2_p_spl_
  );


  or

  (
    g498_n,
    n770_o2_p_spl_,
    n767_o2_n_spl_
  );


  and

  (
    g499_p,
    g497_n,
    g498_n
  );


  or

  (
    g499_n,
    g497_p,
    g498_p
  );


  and

  (
    g500_p,
    lo145_buf_o2_p,
    lo161_buf_o2_p_spl_10
  );


  or

  (
    g500_n,
    lo145_buf_o2_n,
    lo161_buf_o2_n_spl_10
  );


  and

  (
    g501_p,
    g499_n,
    g500_p
  );


  and

  (
    g502_p,
    g499_p,
    g500_n
  );


  or

  (
    g503_n,
    g501_p,
    g502_p
  );


  and

  (
    g504_p,
    n708_o2_p_spl_,
    n705_o2_n_spl_
  );


  or

  (
    g504_n,
    n708_o2_n_spl_,
    n705_o2_p_spl_
  );


  and

  (
    g505_p,
    n708_o2_n_spl_,
    n705_o2_p_spl_
  );


  or

  (
    g505_n,
    n708_o2_p_spl_,
    n705_o2_n_spl_
  );


  and

  (
    g506_p,
    g504_n,
    g505_n
  );


  or

  (
    g506_n,
    g504_p,
    g505_p
  );


  and

  (
    g507_p,
    n745_o2_p_spl_,
    n742_o2_n_spl_
  );


  or

  (
    g507_n,
    n745_o2_n_spl_,
    n742_o2_p_spl_
  );


  and

  (
    g508_p,
    n745_o2_n_spl_,
    n742_o2_p_spl_
  );


  or

  (
    g508_n,
    n745_o2_p_spl_,
    n742_o2_n_spl_
  );


  and

  (
    g509_p,
    g507_n,
    g508_n
  );


  or

  (
    g509_n,
    g507_p,
    g508_p
  );


  and

  (
    g510_p,
    g506_p_spl_,
    g509_n_spl_
  );


  and

  (
    g511_p,
    g506_n_spl_,
    g509_p_spl_
  );


  or

  (
    g512_n,
    g510_p,
    g511_p
  );


  and

  (
    g513_p,
    g503_n_spl_,
    g512_n_spl_
  );


  or

  (
    g514_n,
    g503_n_spl_,
    g512_n_spl_
  );


  and

  (
    g515_p,
    n789_o2_p_spl_,
    n786_o2_n_spl_
  );


  or

  (
    g515_n,
    n789_o2_n_spl_,
    n786_o2_p_spl_
  );


  and

  (
    g516_p,
    n789_o2_n_spl_,
    n786_o2_p_spl_
  );


  or

  (
    g516_n,
    n789_o2_p_spl_,
    n786_o2_n_spl_
  );


  and

  (
    g517_p,
    g515_n,
    g516_n
  );


  or

  (
    g517_n,
    g515_p,
    g516_p
  );


  and

  (
    g518_p,
    lo149_buf_o2_p,
    lo161_buf_o2_p_spl_10
  );


  or

  (
    g518_n,
    lo149_buf_o2_n,
    lo161_buf_o2_n_spl_10
  );


  and

  (
    g519_p,
    g517_n,
    g518_p
  );


  and

  (
    g520_p,
    g517_p,
    g518_n
  );


  or

  (
    g521_n,
    g519_p,
    g520_p
  );


  and

  (
    g522_p,
    n717_o2_p_spl_,
    n714_o2_n_spl_
  );


  or

  (
    g522_n,
    n717_o2_n_spl_,
    n714_o2_p_spl_
  );


  and

  (
    g523_p,
    n717_o2_n_spl_,
    n714_o2_p_spl_
  );


  or

  (
    g523_n,
    n717_o2_p_spl_,
    n714_o2_n_spl_
  );


  and

  (
    g524_p,
    g522_n,
    g523_n
  );


  or

  (
    g524_n,
    g522_p,
    g523_p
  );


  and

  (
    g525_p,
    n754_o2_p_spl_,
    n751_o2_n_spl_
  );


  or

  (
    g525_n,
    n754_o2_n_spl_,
    n751_o2_p_spl_
  );


  and

  (
    g526_p,
    n754_o2_n_spl_,
    n751_o2_p_spl_
  );


  or

  (
    g526_n,
    n754_o2_p_spl_,
    n751_o2_n_spl_
  );


  and

  (
    g527_p,
    g525_n,
    g526_n
  );


  or

  (
    g527_n,
    g525_p,
    g526_p
  );


  and

  (
    g528_p,
    g524_p_spl_,
    g527_n_spl_
  );


  and

  (
    g529_p,
    g524_n_spl_,
    g527_p_spl_
  );


  or

  (
    g530_n,
    g528_p,
    g529_p
  );


  and

  (
    g531_p,
    g521_n_spl_,
    g530_n_spl_
  );


  or

  (
    g532_n,
    g521_n_spl_,
    g530_n_spl_
  );


  and

  (
    g533_p,
    n695_o2_p_spl_,
    n692_o2_n_spl_
  );


  or

  (
    g533_n,
    n695_o2_n_spl_,
    n692_o2_p_spl_
  );


  and

  (
    g534_p,
    n695_o2_n_spl_,
    n692_o2_p_spl_
  );


  or

  (
    g534_n,
    n695_o2_p_spl_,
    n692_o2_n_spl_
  );


  and

  (
    g535_p,
    g533_n,
    g534_n
  );


  or

  (
    g535_n,
    g533_p,
    g534_p
  );


  and

  (
    g536_p,
    lo153_buf_o2_p,
    lo161_buf_o2_p_spl_11
  );


  or

  (
    g536_n,
    lo153_buf_o2_n,
    lo161_buf_o2_n_spl_11
  );


  and

  (
    g537_p,
    g535_n,
    g536_p
  );


  and

  (
    g538_p,
    g535_p,
    g536_n
  );


  or

  (
    g539_n,
    g537_p,
    g538_p
  );


  and

  (
    g540_p,
    g506_p_spl_,
    g524_n_spl_
  );


  and

  (
    g541_p,
    g506_n_spl_,
    g524_p_spl_
  );


  or

  (
    g542_n,
    g540_p,
    g541_p
  );


  and

  (
    g543_p,
    g539_n_spl_,
    g542_n_spl_
  );


  or

  (
    g544_n,
    g539_n_spl_,
    g542_n_spl_
  );


  and

  (
    g545_p,
    n732_o2_p_spl_,
    n729_o2_n_spl_
  );


  or

  (
    g545_n,
    n732_o2_n_spl_,
    n729_o2_p_spl_
  );


  and

  (
    g546_p,
    n732_o2_n_spl_,
    n729_o2_p_spl_
  );


  or

  (
    g546_n,
    n732_o2_p_spl_,
    n729_o2_n_spl_
  );


  and

  (
    g547_p,
    g545_n,
    g546_n
  );


  or

  (
    g547_n,
    g545_p,
    g546_p
  );


  and

  (
    g548_p,
    lo157_buf_o2_p,
    lo161_buf_o2_p_spl_11
  );


  or

  (
    g548_n,
    lo157_buf_o2_n,
    lo161_buf_o2_n_spl_11
  );


  and

  (
    g549_p,
    g547_n,
    g548_p
  );


  and

  (
    g550_p,
    g547_p,
    g548_n
  );


  or

  (
    g551_n,
    g549_p,
    g550_p
  );


  and

  (
    g552_p,
    g509_p_spl_,
    g527_n_spl_
  );


  and

  (
    g553_p,
    g509_n_spl_,
    g527_p_spl_
  );


  or

  (
    g554_n,
    g552_p,
    g553_p
  );


  and

  (
    g555_p,
    g551_n_spl_,
    g554_n_spl_
  );


  or

  (
    g556_n,
    g551_n_spl_,
    g554_n_spl_
  );


  or

  (
    g557_n,
    n621_lo_p_spl_0,
    n669_lo_p_spl_0
  );


  or

  (
    g558_n,
    n621_lo_n_spl_,
    n669_lo_n_spl_
  );


  and

  (
    g559_p,
    g557_n,
    g558_n
  );


  or

  (
    g560_n,
    n621_lo_p_spl_0,
    n633_lo_p_spl_0
  );


  or

  (
    g561_n,
    n621_lo_n_spl_,
    n633_lo_n_spl_
  );


  and

  (
    g562_p,
    g560_n,
    g561_n
  );


  or

  (
    g563_n,
    n633_lo_p_spl_0,
    n681_lo_p_spl_0
  );


  or

  (
    g564_n,
    n633_lo_n_spl_,
    n681_lo_n_spl_
  );


  and

  (
    g565_p,
    g563_n,
    g564_n
  );


  or

  (
    g566_n,
    n645_lo_p_spl_0,
    n693_lo_p_spl_0
  );


  or

  (
    g567_n,
    n645_lo_n_spl_,
    n693_lo_n_spl_
  );


  and

  (
    g568_p,
    g566_n,
    g567_n
  );


  and

  (
    g569_p,
    n645_lo_p_spl_0,
    n657_lo_n_spl_
  );


  and

  (
    g570_p,
    n645_lo_n_spl_,
    n657_lo_p_spl_0
  );


  or

  (
    g571_n,
    g569_p,
    g570_p
  );


  or

  (
    g572_n,
    n657_lo_p_spl_0,
    n705_lo_p_spl_0
  );


  or

  (
    g573_n,
    n657_lo_n_spl_,
    n705_lo_n_spl_
  );


  and

  (
    g574_p,
    g572_n,
    g573_n
  );


  or

  (
    g575_n,
    n669_lo_p_spl_0,
    n681_lo_p_spl_0
  );


  or

  (
    g576_n,
    n669_lo_n_spl_,
    n681_lo_n_spl_
  );


  and

  (
    g577_p,
    g575_n,
    g576_n
  );


  and

  (
    g578_p,
    n693_lo_p_spl_0,
    n705_lo_n_spl_
  );


  and

  (
    g579_p,
    n693_lo_n_spl_,
    n705_lo_p_spl_0
  );


  or

  (
    g580_n,
    g578_p,
    g579_p
  );


  and

  (
    g581_p,
    n717_lo_p_spl_0,
    n765_lo_n_spl_
  );


  and

  (
    g582_p,
    n717_lo_n_spl_,
    n765_lo_p_spl_0
  );


  or

  (
    g583_n,
    g581_p,
    g582_p
  );


  or

  (
    g584_n,
    n717_lo_p_spl_0,
    n729_lo_p_spl_0
  );


  or

  (
    g585_n,
    n717_lo_n_spl_,
    n729_lo_n_spl_
  );


  and

  (
    g586_p,
    g584_n,
    g585_n
  );


  and

  (
    g587_p,
    n729_lo_p_spl_0,
    n777_lo_n_spl_
  );


  and

  (
    g588_p,
    n729_lo_n_spl_,
    n777_lo_p_spl_0
  );


  or

  (
    g589_n,
    g587_p,
    g588_p
  );


  and

  (
    g590_p,
    n741_lo_p_spl_0,
    n789_lo_n_spl_
  );


  and

  (
    g591_p,
    n741_lo_n_spl_,
    n789_lo_p_spl_0
  );


  or

  (
    g592_n,
    g590_p,
    g591_p
  );


  and

  (
    g593_p,
    n741_lo_p_spl_0,
    n753_lo_n_spl_
  );


  and

  (
    g594_p,
    n741_lo_n_spl_,
    n753_lo_p_spl_0
  );


  or

  (
    g595_n,
    g593_p,
    g594_p
  );


  and

  (
    g596_p,
    n753_lo_p_spl_0,
    n801_lo_n_spl_
  );


  and

  (
    g597_p,
    n753_lo_n_spl_,
    n801_lo_p_spl_0
  );


  or

  (
    g598_n,
    g596_p,
    g597_p
  );


  or

  (
    g599_n,
    n765_lo_p_spl_0,
    n777_lo_p_spl_0
  );


  or

  (
    g600_n,
    n765_lo_n_spl_,
    n777_lo_n_spl_
  );


  and

  (
    g601_p,
    g599_n,
    g600_n
  );


  and

  (
    g602_p,
    n789_lo_p_spl_0,
    n801_lo_n_spl_
  );


  and

  (
    g603_p,
    n789_lo_n_spl_,
    n801_lo_p_spl_0
  );


  or

  (
    g604_n,
    g602_p,
    g603_p
  );


  or

  (
    g605_n,
    n813_lo_p_spl_0,
    n825_lo_p_spl_0
  );


  or

  (
    g606_n,
    n813_lo_n_spl_,
    n825_lo_n_spl_
  );


  and

  (
    g607_p,
    g605_n,
    g606_n
  );


  or

  (
    g608_n,
    n813_lo_p_spl_0,
    n861_lo_p_spl_0
  );


  or

  (
    g609_n,
    n813_lo_n_spl_,
    n861_lo_n_spl_
  );


  and

  (
    g610_p,
    g608_n,
    g609_n
  );


  or

  (
    g611_n,
    n825_lo_p_spl_0,
    n873_lo_p_spl_0
  );


  or

  (
    g612_n,
    n825_lo_n_spl_,
    n873_lo_n_spl_
  );


  and

  (
    g613_p,
    g611_n,
    g612_n
  );


  and

  (
    g614_p,
    n837_lo_p_spl_0,
    n849_lo_n_spl_
  );


  and

  (
    g615_p,
    n837_lo_n_spl_,
    n849_lo_p_spl_0
  );


  or

  (
    g616_n,
    g614_p,
    g615_p
  );


  or

  (
    g617_n,
    n837_lo_p_spl_0,
    n885_lo_p_spl_0
  );


  or

  (
    g618_n,
    n837_lo_n_spl_,
    n885_lo_n_spl_
  );


  and

  (
    g619_p,
    g617_n,
    g618_n
  );


  or

  (
    g620_n,
    n849_lo_p_spl_0,
    n897_lo_p_spl_0
  );


  or

  (
    g621_n,
    n849_lo_n_spl_,
    n897_lo_n_spl_
  );


  and

  (
    g622_p,
    g620_n,
    g621_n
  );


  or

  (
    g623_n,
    n861_lo_p_spl_0,
    n873_lo_p_spl_0
  );


  or

  (
    g624_n,
    n861_lo_n_spl_,
    n873_lo_n_spl_
  );


  and

  (
    g625_p,
    g623_n,
    g624_n
  );


  and

  (
    g626_p,
    n885_lo_p_spl_0,
    n897_lo_n_spl_
  );


  and

  (
    g627_p,
    n885_lo_n_spl_,
    n897_lo_p_spl_0
  );


  or

  (
    g628_n,
    g626_p,
    g627_p
  );


  or

  (
    g629_n,
    n909_lo_p_spl_0,
    n921_lo_p_spl_0
  );


  or

  (
    g630_n,
    n909_lo_n_spl_,
    n921_lo_n_spl_
  );


  and

  (
    g631_p,
    g629_n,
    g630_n
  );


  and

  (
    g632_p,
    n909_lo_p_spl_0,
    n957_lo_n_spl_
  );


  and

  (
    g633_p,
    n909_lo_n_spl_,
    n957_lo_p_spl_0
  );


  or

  (
    g634_n,
    g632_p,
    g633_p
  );


  and

  (
    g635_p,
    n921_lo_p_spl_0,
    n969_lo_n_spl_
  );


  and

  (
    g636_p,
    n921_lo_n_spl_,
    n969_lo_p_spl_0
  );


  or

  (
    g637_n,
    g635_p,
    g636_p
  );


  and

  (
    g638_p,
    n933_lo_p_spl_0,
    n945_lo_n_spl_
  );


  and

  (
    g639_p,
    n933_lo_n_spl_,
    n945_lo_p_spl_0
  );


  or

  (
    g640_n,
    g638_p,
    g639_p
  );


  and

  (
    g641_p,
    n933_lo_p_spl_0,
    n981_lo_n_spl_
  );


  and

  (
    g642_p,
    n933_lo_n_spl_,
    n981_lo_p_spl_0
  );


  or

  (
    g643_n,
    g641_p,
    g642_p
  );


  and

  (
    g644_p,
    n945_lo_p_spl_0,
    n993_lo_n_spl_
  );


  and

  (
    g645_p,
    n945_lo_n_spl_,
    n993_lo_p_spl_0
  );


  or

  (
    g646_n,
    g644_p,
    g645_p
  );


  or

  (
    g647_n,
    n957_lo_p_spl_0,
    n969_lo_p_spl_0
  );


  or

  (
    g648_n,
    n957_lo_n_spl_,
    n969_lo_n_spl_
  );


  and

  (
    g649_p,
    g647_n,
    g648_n
  );


  and

  (
    g650_p,
    n981_lo_p_spl_0,
    n993_lo_n_spl_
  );


  and

  (
    g651_p,
    n981_lo_n_spl_,
    n993_lo_p_spl_0
  );


  or

  (
    g652_n,
    g650_p,
    g651_p
  );


  buf

  (
    G1324,
    g266_p
  );


  buf

  (
    G1325,
    g270_p
  );


  buf

  (
    G1326,
    g274_p
  );


  buf

  (
    G1327,
    g278_p
  );


  buf

  (
    G1328,
    g284_p
  );


  buf

  (
    G1329,
    g288_p
  );


  buf

  (
    G1330,
    g292_p
  );


  buf

  (
    G1331,
    g296_p
  );


  buf

  (
    G1332,
    g302_p
  );


  buf

  (
    G1333,
    g306_p
  );


  buf

  (
    G1334,
    g310_p
  );


  buf

  (
    G1335,
    g314_p
  );


  buf

  (
    G1336,
    g320_p
  );


  buf

  (
    G1337,
    g324_p
  );


  buf

  (
    G1338,
    g328_p
  );


  buf

  (
    G1339,
    g332_p
  );


  buf

  (
    G1340,
    g338_p
  );


  buf

  (
    G1341,
    g342_p
  );


  buf

  (
    G1342,
    g346_p
  );


  buf

  (
    G1343,
    g350_p
  );


  buf

  (
    G1344,
    g356_p
  );


  buf

  (
    G1345,
    g360_p
  );


  buf

  (
    G1346,
    g364_p
  );


  buf

  (
    G1347,
    g368_p
  );


  buf

  (
    G1348,
    g374_p
  );


  buf

  (
    G1349,
    g378_p
  );


  buf

  (
    G1350,
    g382_p
  );


  buf

  (
    G1351,
    g386_p
  );


  buf

  (
    G1352,
    g392_p
  );


  buf

  (
    G1353,
    g396_p
  );


  buf

  (
    G1354,
    g400_p
  );


  buf

  (
    G1355,
    g404_p
  );


  buf

  (
    n1699_li000_li000,
    G1_p
  );


  buf

  (
    n1708_li003_li003,
    n1644_o2_p
  );


  buf

  (
    n1711_li004_li004,
    G2_p
  );


  buf

  (
    n1720_li007_li007,
    n1645_o2_p
  );


  buf

  (
    n1723_li008_li008,
    G3_p
  );


  buf

  (
    n1732_li011_li011,
    n1646_o2_p
  );


  buf

  (
    n1735_li012_li012,
    G4_p
  );


  buf

  (
    n1744_li015_li015,
    n1647_o2_p
  );


  buf

  (
    n1747_li016_li016,
    G5_p
  );


  buf

  (
    n1756_li019_li019,
    n1648_o2_p
  );


  buf

  (
    n1759_li020_li020,
    G6_p
  );


  buf

  (
    n1768_li023_li023,
    n1649_o2_p
  );


  buf

  (
    n1771_li024_li024,
    G7_p
  );


  buf

  (
    n1780_li027_li027,
    n1650_o2_p
  );


  buf

  (
    n1783_li028_li028,
    G8_p
  );


  buf

  (
    n1792_li031_li031,
    n1651_o2_p
  );


  buf

  (
    n1795_li032_li032,
    G9_p
  );


  buf

  (
    n1804_li035_li035,
    n1652_o2_p
  );


  buf

  (
    n1807_li036_li036,
    G10_p
  );


  buf

  (
    n1816_li039_li039,
    n1653_o2_p
  );


  buf

  (
    n1819_li040_li040,
    G11_p
  );


  buf

  (
    n1828_li043_li043,
    n1654_o2_p
  );


  buf

  (
    n1831_li044_li044,
    G12_p
  );


  buf

  (
    n1840_li047_li047,
    n1655_o2_p
  );


  buf

  (
    n1843_li048_li048,
    G13_p
  );


  buf

  (
    n1852_li051_li051,
    n1656_o2_p
  );


  buf

  (
    n1855_li052_li052,
    G14_p
  );


  buf

  (
    n1864_li055_li055,
    n1657_o2_p
  );


  buf

  (
    n1867_li056_li056,
    G15_p
  );


  buf

  (
    n1876_li059_li059,
    n1658_o2_p
  );


  buf

  (
    n1879_li060_li060,
    G16_p
  );


  buf

  (
    n1888_li063_li063,
    n1659_o2_p
  );


  buf

  (
    n1891_li064_li064,
    G17_p
  );


  buf

  (
    n1900_li067_li067,
    n1660_o2_p
  );


  buf

  (
    n1903_li068_li068,
    G18_p
  );


  buf

  (
    n1912_li071_li071,
    n1661_o2_p
  );


  buf

  (
    n1915_li072_li072,
    G19_p
  );


  buf

  (
    n1924_li075_li075,
    n1662_o2_p
  );


  buf

  (
    n1927_li076_li076,
    G20_p
  );


  buf

  (
    n1936_li079_li079,
    n1663_o2_p
  );


  buf

  (
    n1939_li080_li080,
    G21_p
  );


  buf

  (
    n1948_li083_li083,
    n1664_o2_p
  );


  buf

  (
    n1951_li084_li084,
    G22_p
  );


  buf

  (
    n1960_li087_li087,
    n1665_o2_p
  );


  buf

  (
    n1963_li088_li088,
    G23_p
  );


  buf

  (
    n1972_li091_li091,
    n1666_o2_p
  );


  buf

  (
    n1975_li092_li092,
    G24_p
  );


  buf

  (
    n1984_li095_li095,
    n1667_o2_p
  );


  buf

  (
    n1987_li096_li096,
    G25_p
  );


  buf

  (
    n1996_li099_li099,
    n1668_o2_p
  );


  buf

  (
    n1999_li100_li100,
    G26_p
  );


  buf

  (
    n2008_li103_li103,
    n1669_o2_p
  );


  buf

  (
    n2011_li104_li104,
    G27_p
  );


  buf

  (
    n2020_li107_li107,
    n1670_o2_p
  );


  buf

  (
    n2023_li108_li108,
    G28_p
  );


  buf

  (
    n2032_li111_li111,
    n1671_o2_p
  );


  buf

  (
    n2035_li112_li112,
    G29_p
  );


  buf

  (
    n2044_li115_li115,
    n1672_o2_p
  );


  buf

  (
    n2047_li116_li116,
    G30_p
  );


  buf

  (
    n2056_li119_li119,
    n1673_o2_p
  );


  buf

  (
    n2059_li120_li120,
    G31_p
  );


  buf

  (
    n2068_li123_li123,
    n1674_o2_p
  );


  buf

  (
    n2071_li124_li124,
    G32_p
  );


  buf

  (
    n2080_li127_li127,
    n1675_o2_p
  );


  buf

  (
    n2083_li128_li128,
    G33_p
  );


  buf

  (
    n2095_li132_li132,
    G34_p
  );


  buf

  (
    n2107_li136_li136,
    G35_p
  );


  buf

  (
    n2119_li140_li140,
    G36_p
  );


  buf

  (
    n2131_li144_li144,
    G37_p
  );


  buf

  (
    n2143_li148_li148,
    G38_p
  );


  buf

  (
    n2155_li152_li152,
    G39_p
  );


  buf

  (
    n2167_li156_li156,
    G40_p
  );


  buf

  (
    n2179_li160_li160,
    G41_p
  );


  buf

  (
    n602_i2,
    g405_n_spl_
  );


  buf

  (
    n639_i2,
    g406_n_spl_
  );


  buf

  (
    n678_i2,
    g407_n_spl_
  );


  buf

  (
    n658_i2,
    g408_n_spl_
  );


  buf

  (
    n783_i2,
    g409_n_spl_
  );


  buf

  (
    n802_i2,
    g410_n_spl_
  );


  buf

  (
    n726_i2,
    g411_n_spl_
  );


  buf

  (
    n763_i2,
    g412_n_spl_
  );


  buf

  (
    n1644_i2,
    lo002_buf_o2_p
  );


  buf

  (
    n1645_i2,
    lo006_buf_o2_p
  );


  buf

  (
    n1646_i2,
    lo010_buf_o2_p
  );


  buf

  (
    n1647_i2,
    lo014_buf_o2_p
  );


  buf

  (
    n1648_i2,
    lo018_buf_o2_p
  );


  buf

  (
    n1649_i2,
    lo022_buf_o2_p
  );


  buf

  (
    n1650_i2,
    lo026_buf_o2_p
  );


  buf

  (
    n1651_i2,
    lo030_buf_o2_p
  );


  buf

  (
    n1652_i2,
    lo034_buf_o2_p
  );


  buf

  (
    n1653_i2,
    lo038_buf_o2_p
  );


  buf

  (
    n1654_i2,
    lo042_buf_o2_p
  );


  buf

  (
    n1655_i2,
    lo046_buf_o2_p
  );


  buf

  (
    n1656_i2,
    lo050_buf_o2_p
  );


  buf

  (
    n1657_i2,
    lo054_buf_o2_p
  );


  buf

  (
    n1658_i2,
    lo058_buf_o2_p
  );


  buf

  (
    n1659_i2,
    lo062_buf_o2_p
  );


  buf

  (
    n1660_i2,
    lo066_buf_o2_p
  );


  buf

  (
    n1661_i2,
    lo070_buf_o2_p
  );


  buf

  (
    n1662_i2,
    lo074_buf_o2_p
  );


  buf

  (
    n1663_i2,
    lo078_buf_o2_p
  );


  buf

  (
    n1664_i2,
    lo082_buf_o2_p
  );


  buf

  (
    n1665_i2,
    lo086_buf_o2_p
  );


  buf

  (
    n1666_i2,
    lo090_buf_o2_p
  );


  buf

  (
    n1667_i2,
    lo094_buf_o2_p
  );


  buf

  (
    n1668_i2,
    lo098_buf_o2_p
  );


  buf

  (
    n1669_i2,
    lo102_buf_o2_p
  );


  buf

  (
    n1670_i2,
    lo106_buf_o2_p
  );


  buf

  (
    n1671_i2,
    lo110_buf_o2_p
  );


  buf

  (
    n1672_i2,
    lo114_buf_o2_p
  );


  buf

  (
    n1673_i2,
    lo118_buf_o2_p
  );


  buf

  (
    n1674_i2,
    lo122_buf_o2_p
  );


  buf

  (
    n1675_i2,
    lo126_buf_o2_p
  );


  not

  (
    n685_i2,
    g413_n_spl_
  );


  not

  (
    n680_i2,
    g414_n_spl_
  );


  not

  (
    n822_i2,
    g415_n_spl_
  );


  buf

  (
    n843_i2,
    g416_n_spl_
  );


  not

  (
    n842_i2,
    g417_n_spl_
  );


  not

  (
    n681_i2,
    g418_n_spl_
  );


  not

  (
    n684_i2,
    g420_n_spl_
  );


  not

  (
    n686_i2,
    g421_n_spl_
  );


  buf

  (
    n823_i2,
    g422_n_spl_
  );


  not

  (
    n683_i2,
    g425_n
  );


  not

  (
    n688_i2,
    g427_n
  );


  buf

  (
    n803_i2,
    g428_p
  );


  buf

  (
    n862_i2,
    g429_p
  );


  buf

  (
    n764_i2,
    g430_p
  );


  buf

  (
    n863_i2,
    g431_p
  );


  buf

  (
    n886_i2,
    g436_p
  );


  buf

  (
    lo002_buf_i2,
    n621_lo_p_spl_
  );


  buf

  (
    lo006_buf_i2,
    n633_lo_p_spl_
  );


  buf

  (
    lo010_buf_i2,
    n645_lo_p_spl_
  );


  buf

  (
    lo014_buf_i2,
    n657_lo_p_spl_
  );


  buf

  (
    lo018_buf_i2,
    n669_lo_p_spl_
  );


  buf

  (
    lo022_buf_i2,
    n681_lo_p_spl_
  );


  buf

  (
    lo026_buf_i2,
    n693_lo_p_spl_
  );


  buf

  (
    lo030_buf_i2,
    n705_lo_p_spl_
  );


  buf

  (
    lo034_buf_i2,
    n717_lo_p_spl_
  );


  buf

  (
    lo038_buf_i2,
    n729_lo_p_spl_
  );


  buf

  (
    lo042_buf_i2,
    n741_lo_p_spl_
  );


  buf

  (
    lo046_buf_i2,
    n753_lo_p_spl_
  );


  buf

  (
    lo050_buf_i2,
    n765_lo_p_spl_
  );


  buf

  (
    lo054_buf_i2,
    n777_lo_p_spl_
  );


  buf

  (
    lo058_buf_i2,
    n789_lo_p_spl_
  );


  buf

  (
    lo062_buf_i2,
    n801_lo_p_spl_
  );


  buf

  (
    lo066_buf_i2,
    n813_lo_p_spl_
  );


  buf

  (
    lo070_buf_i2,
    n825_lo_p_spl_
  );


  buf

  (
    lo074_buf_i2,
    n837_lo_p_spl_
  );


  buf

  (
    lo078_buf_i2,
    n849_lo_p_spl_
  );


  buf

  (
    lo082_buf_i2,
    n861_lo_p_spl_
  );


  buf

  (
    lo086_buf_i2,
    n873_lo_p_spl_
  );


  buf

  (
    lo090_buf_i2,
    n885_lo_p_spl_
  );


  buf

  (
    lo094_buf_i2,
    n897_lo_p_spl_
  );


  buf

  (
    lo098_buf_i2,
    n909_lo_p_spl_
  );


  buf

  (
    lo102_buf_i2,
    n921_lo_p_spl_
  );


  buf

  (
    lo106_buf_i2,
    n933_lo_p_spl_
  );


  buf

  (
    lo110_buf_i2,
    n945_lo_p_spl_
  );


  buf

  (
    lo114_buf_i2,
    n957_lo_p_spl_
  );


  buf

  (
    lo118_buf_i2,
    n969_lo_p_spl_
  );


  buf

  (
    lo122_buf_i2,
    n981_lo_p_spl_
  );


  buf

  (
    lo126_buf_i2,
    n993_lo_p_spl_
  );


  buf

  (
    n600_i2,
    g453_p
  );


  not

  (
    n601_i2,
    g454_n
  );


  buf

  (
    n637_i2,
    g471_p
  );


  not

  (
    n638_i2,
    g472_n
  );


  buf

  (
    n676_i2,
    g483_p
  );


  not

  (
    n677_i2,
    g484_n
  );


  buf

  (
    n656_i2,
    g495_p
  );


  not

  (
    n657_i2,
    g496_n
  );


  buf

  (
    n781_i2,
    g513_p
  );


  not

  (
    n782_i2,
    g514_n
  );


  buf

  (
    n800_i2,
    g531_p
  );


  not

  (
    n801_i2,
    g532_n
  );


  buf

  (
    n724_i2,
    g543_p
  );


  not

  (
    n725_i2,
    g544_n
  );


  buf

  (
    n761_i2,
    g555_p
  );


  not

  (
    n762_i2,
    g556_n
  );


  buf

  (
    lo129_buf_i2,
    n1005_lo_p
  );


  buf

  (
    lo133_buf_i2,
    n1017_lo_p
  );


  buf

  (
    lo137_buf_i2,
    n1029_lo_p
  );


  buf

  (
    lo141_buf_i2,
    n1041_lo_p
  );


  buf

  (
    lo145_buf_i2,
    n1053_lo_p
  );


  buf

  (
    lo149_buf_i2,
    n1065_lo_p
  );


  buf

  (
    lo153_buf_i2,
    n1077_lo_p
  );


  buf

  (
    lo157_buf_i2,
    n1089_lo_p
  );


  buf

  (
    lo161_buf_i2,
    n1101_lo_p
  );


  buf

  (
    n571_i2,
    g559_p
  );


  buf

  (
    n708_i2,
    g562_p
  );


  buf

  (
    n608_i2,
    g565_p
  );


  buf

  (
    n665_i2,
    g568_p
  );


  buf

  (
    n705_i2,
    g571_n
  );


  buf

  (
    n645_i2,
    g574_p
  );


  buf

  (
    n745_i2,
    g577_p
  );


  buf

  (
    n742_i2,
    g580_n
  );


  buf

  (
    n568_i2,
    g583_n
  );


  buf

  (
    n717_i2,
    g586_p
  );


  buf

  (
    n605_i2,
    g589_n
  );


  buf

  (
    n662_i2,
    g592_n
  );


  buf

  (
    n714_i2,
    g595_n
  );


  buf

  (
    n642_i2,
    g598_n
  );


  buf

  (
    n754_i2,
    g601_p
  );


  buf

  (
    n751_i2,
    g604_n
  );


  buf

  (
    n584_i2,
    g607_p
  );


  buf

  (
    n770_i2,
    g610_p
  );


  buf

  (
    n789_i2,
    g613_p
  );


  buf

  (
    n581_i2,
    g616_n
  );


  buf

  (
    n695_i2,
    g619_p
  );


  buf

  (
    n732_i2,
    g622_p
  );


  buf

  (
    n593_i2,
    g625_p
  );


  buf

  (
    n590_i2,
    g628_n
  );


  buf

  (
    n630_i2,
    g631_p
  );


  buf

  (
    n767_i2,
    g634_n
  );


  buf

  (
    n786_i2,
    g637_n
  );


  buf

  (
    n627_i2,
    g640_n
  );


  buf

  (
    n692_i2,
    g643_n
  );


  buf

  (
    n729_i2,
    g646_n
  );


  buf

  (
    n621_i2,
    g649_p
  );


  buf

  (
    n618_i2,
    g652_n
  );


  buf

  (
    g260_n_spl_,
    g260_n
  );


  buf

  (
    g260_n_spl_0,
    g260_n_spl_
  );


  buf

  (
    g260_n_spl_1,
    g260_n_spl_
  );


  buf

  (
    g260_p_spl_,
    g260_p
  );


  buf

  (
    g260_p_spl_0,
    g260_p_spl_
  );


  buf

  (
    g260_p_spl_1,
    g260_p_spl_
  );


  buf

  (
    n602_o2_p_spl_,
    n602_o2_p
  );


  buf

  (
    n602_o2_p_spl_0,
    n602_o2_p_spl_
  );


  buf

  (
    n602_o2_p_spl_1,
    n602_o2_p_spl_
  );


  buf

  (
    g262_p_spl_,
    g262_p
  );


  buf

  (
    g262_p_spl_0,
    g262_p_spl_
  );


  buf

  (
    g262_p_spl_1,
    g262_p_spl_
  );


  buf

  (
    n602_o2_n_spl_,
    n602_o2_n
  );


  buf

  (
    n602_o2_n_spl_0,
    n602_o2_n_spl_
  );


  buf

  (
    n602_o2_n_spl_1,
    n602_o2_n_spl_
  );


  buf

  (
    g262_n_spl_,
    g262_n
  );


  buf

  (
    g262_n_spl_0,
    g262_n_spl_
  );


  buf

  (
    g262_n_spl_1,
    g262_n_spl_
  );


  buf

  (
    n639_o2_p_spl_,
    n639_o2_p
  );


  buf

  (
    n639_o2_p_spl_0,
    n639_o2_p_spl_
  );


  buf

  (
    n639_o2_p_spl_00,
    n639_o2_p_spl_0
  );


  buf

  (
    n639_o2_p_spl_1,
    n639_o2_p_spl_
  );


  buf

  (
    n639_o2_n_spl_,
    n639_o2_n
  );


  buf

  (
    n639_o2_n_spl_0,
    n639_o2_n_spl_
  );


  buf

  (
    n639_o2_n_spl_00,
    n639_o2_n_spl_0
  );


  buf

  (
    n639_o2_n_spl_1,
    n639_o2_n_spl_
  );


  buf

  (
    n678_o2_p_spl_,
    n678_o2_p
  );


  buf

  (
    n678_o2_p_spl_0,
    n678_o2_p_spl_
  );


  buf

  (
    n678_o2_p_spl_00,
    n678_o2_p_spl_0
  );


  buf

  (
    n678_o2_p_spl_01,
    n678_o2_p_spl_0
  );


  buf

  (
    n678_o2_p_spl_1,
    n678_o2_p_spl_
  );


  buf

  (
    n678_o2_n_spl_,
    n678_o2_n
  );


  buf

  (
    n678_o2_n_spl_0,
    n678_o2_n_spl_
  );


  buf

  (
    n678_o2_n_spl_00,
    n678_o2_n_spl_0
  );


  buf

  (
    n678_o2_n_spl_01,
    n678_o2_n_spl_0
  );


  buf

  (
    n678_o2_n_spl_1,
    n678_o2_n_spl_
  );


  buf

  (
    n658_o2_p_spl_,
    n658_o2_p
  );


  buf

  (
    n658_o2_p_spl_0,
    n658_o2_p_spl_
  );


  buf

  (
    n658_o2_p_spl_1,
    n658_o2_p_spl_
  );


  buf

  (
    n658_o2_n_spl_,
    n658_o2_n
  );


  buf

  (
    n658_o2_n_spl_0,
    n658_o2_n_spl_
  );


  buf

  (
    n658_o2_n_spl_1,
    n658_o2_n_spl_
  );


  buf

  (
    g280_p_spl_,
    g280_p
  );


  buf

  (
    g280_p_spl_0,
    g280_p_spl_
  );


  buf

  (
    g280_p_spl_1,
    g280_p_spl_
  );


  buf

  (
    g280_n_spl_,
    g280_n
  );


  buf

  (
    g280_n_spl_0,
    g280_n_spl_
  );


  buf

  (
    g280_n_spl_1,
    g280_n_spl_
  );


  buf

  (
    g298_p_spl_,
    g298_p
  );


  buf

  (
    g298_p_spl_0,
    g298_p_spl_
  );


  buf

  (
    g298_p_spl_1,
    g298_p_spl_
  );


  buf

  (
    g298_n_spl_,
    g298_n
  );


  buf

  (
    g298_n_spl_0,
    g298_n_spl_
  );


  buf

  (
    g298_n_spl_1,
    g298_n_spl_
  );


  buf

  (
    g316_p_spl_,
    g316_p
  );


  buf

  (
    g316_p_spl_0,
    g316_p_spl_
  );


  buf

  (
    g316_p_spl_1,
    g316_p_spl_
  );


  buf

  (
    g316_n_spl_,
    g316_n
  );


  buf

  (
    g316_n_spl_0,
    g316_n_spl_
  );


  buf

  (
    g316_n_spl_1,
    g316_n_spl_
  );


  buf

  (
    n886_o2_p_spl_,
    n886_o2_p
  );


  buf

  (
    n886_o2_p_spl_0,
    n886_o2_p_spl_
  );


  buf

  (
    n886_o2_p_spl_1,
    n886_o2_p_spl_
  );


  buf

  (
    n886_o2_n_spl_,
    n886_o2_n
  );


  buf

  (
    n886_o2_n_spl_0,
    n886_o2_n_spl_
  );


  buf

  (
    n886_o2_n_spl_1,
    n886_o2_n_spl_
  );


  buf

  (
    n783_o2_p_spl_,
    n783_o2_p
  );


  buf

  (
    n783_o2_p_spl_0,
    n783_o2_p_spl_
  );


  buf

  (
    n783_o2_p_spl_1,
    n783_o2_p_spl_
  );


  buf

  (
    g334_p_spl_,
    g334_p
  );


  buf

  (
    g334_p_spl_0,
    g334_p_spl_
  );


  buf

  (
    g334_p_spl_1,
    g334_p_spl_
  );


  buf

  (
    n783_o2_n_spl_,
    n783_o2_n
  );


  buf

  (
    n783_o2_n_spl_0,
    n783_o2_n_spl_
  );


  buf

  (
    n783_o2_n_spl_1,
    n783_o2_n_spl_
  );


  buf

  (
    g334_n_spl_,
    g334_n
  );


  buf

  (
    g334_n_spl_0,
    g334_n_spl_
  );


  buf

  (
    g334_n_spl_1,
    g334_n_spl_
  );


  buf

  (
    n802_o2_p_spl_,
    n802_o2_p
  );


  buf

  (
    n802_o2_p_spl_0,
    n802_o2_p_spl_
  );


  buf

  (
    n802_o2_p_spl_1,
    n802_o2_p_spl_
  );


  buf

  (
    n802_o2_n_spl_,
    n802_o2_n
  );


  buf

  (
    n802_o2_n_spl_0,
    n802_o2_n_spl_
  );


  buf

  (
    n802_o2_n_spl_1,
    n802_o2_n_spl_
  );


  buf

  (
    n726_o2_p_spl_,
    n726_o2_p
  );


  buf

  (
    n726_o2_p_spl_0,
    n726_o2_p_spl_
  );


  buf

  (
    n726_o2_p_spl_1,
    n726_o2_p_spl_
  );


  buf

  (
    n726_o2_n_spl_,
    n726_o2_n
  );


  buf

  (
    n726_o2_n_spl_0,
    n726_o2_n_spl_
  );


  buf

  (
    n726_o2_n_spl_1,
    n726_o2_n_spl_
  );


  buf

  (
    n763_o2_p_spl_,
    n763_o2_p
  );


  buf

  (
    n763_o2_p_spl_0,
    n763_o2_p_spl_
  );


  buf

  (
    n763_o2_p_spl_1,
    n763_o2_p_spl_
  );


  buf

  (
    n763_o2_n_spl_,
    n763_o2_n
  );


  buf

  (
    n763_o2_n_spl_0,
    n763_o2_n_spl_
  );


  buf

  (
    n763_o2_n_spl_1,
    n763_o2_n_spl_
  );


  buf

  (
    g352_p_spl_,
    g352_p
  );


  buf

  (
    g352_p_spl_0,
    g352_p_spl_
  );


  buf

  (
    g352_p_spl_1,
    g352_p_spl_
  );


  buf

  (
    g352_n_spl_,
    g352_n
  );


  buf

  (
    g352_n_spl_0,
    g352_n_spl_
  );


  buf

  (
    g352_n_spl_1,
    g352_n_spl_
  );


  buf

  (
    g370_p_spl_,
    g370_p
  );


  buf

  (
    g370_p_spl_0,
    g370_p_spl_
  );


  buf

  (
    g370_p_spl_1,
    g370_p_spl_
  );


  buf

  (
    g370_n_spl_,
    g370_n
  );


  buf

  (
    g370_n_spl_0,
    g370_n_spl_
  );


  buf

  (
    g370_n_spl_1,
    g370_n_spl_
  );


  buf

  (
    g388_p_spl_,
    g388_p
  );


  buf

  (
    g388_p_spl_0,
    g388_p_spl_
  );


  buf

  (
    g388_p_spl_1,
    g388_p_spl_
  );


  buf

  (
    g388_n_spl_,
    g388_n
  );


  buf

  (
    g388_n_spl_0,
    g388_n_spl_
  );


  buf

  (
    g388_n_spl_1,
    g388_n_spl_
  );


  buf

  (
    g406_n_spl_,
    g406_n
  );


  buf

  (
    g406_n_spl_0,
    g406_n_spl_
  );


  buf

  (
    g407_n_spl_,
    g407_n
  );


  buf

  (
    g407_n_spl_0,
    g407_n_spl_
  );


  buf

  (
    g409_p_spl_,
    g409_p
  );


  buf

  (
    g409_p_spl_0,
    g409_p_spl_
  );


  buf

  (
    g412_p_spl_,
    g412_p
  );


  buf

  (
    g412_p_spl_0,
    g412_p_spl_
  );


  buf

  (
    g409_n_spl_,
    g409_n
  );


  buf

  (
    g409_n_spl_0,
    g409_n_spl_
  );


  buf

  (
    g412_n_spl_,
    g412_n
  );


  buf

  (
    g412_n_spl_0,
    g412_n_spl_
  );


  buf

  (
    g410_p_spl_,
    g410_p
  );


  buf

  (
    g410_p_spl_0,
    g410_p_spl_
  );


  buf

  (
    g411_p_spl_,
    g411_p
  );


  buf

  (
    g411_p_spl_0,
    g411_p_spl_
  );


  buf

  (
    g405_n_spl_,
    g405_n
  );


  buf

  (
    g405_n_spl_0,
    g405_n_spl_
  );


  buf

  (
    g414_n_spl_,
    g414_n
  );


  buf

  (
    g408_n_spl_,
    g408_n
  );


  buf

  (
    g408_n_spl_0,
    g408_n_spl_
  );


  buf

  (
    g419_n_spl_,
    g419_n
  );


  buf

  (
    g413_n_spl_,
    g413_n
  );


  buf

  (
    g410_n_spl_,
    g410_n
  );


  buf

  (
    g410_n_spl_0,
    g410_n_spl_
  );


  buf

  (
    g411_n_spl_,
    g411_n
  );


  buf

  (
    g411_n_spl_0,
    g411_n_spl_
  );


  buf

  (
    g418_n_spl_,
    g418_n
  );


  buf

  (
    g420_n_spl_,
    g420_n
  );


  buf

  (
    g421_n_spl_,
    g421_n
  );


  buf

  (
    g415_n_spl_,
    g415_n
  );


  buf

  (
    g416_n_spl_,
    g416_n
  );


  buf

  (
    g422_n_spl_,
    g422_n
  );


  buf

  (
    g417_n_spl_,
    g417_n
  );


  buf

  (
    n571_o2_p_spl_,
    n571_o2_p
  );


  buf

  (
    n568_o2_n_spl_,
    n568_o2_n
  );


  buf

  (
    n571_o2_n_spl_,
    n571_o2_n
  );


  buf

  (
    n568_o2_p_spl_,
    n568_o2_p
  );


  buf

  (
    lo161_buf_o2_p_spl_,
    lo161_buf_o2_p
  );


  buf

  (
    lo161_buf_o2_p_spl_0,
    lo161_buf_o2_p_spl_
  );


  buf

  (
    lo161_buf_o2_p_spl_00,
    lo161_buf_o2_p_spl_0
  );


  buf

  (
    lo161_buf_o2_p_spl_01,
    lo161_buf_o2_p_spl_0
  );


  buf

  (
    lo161_buf_o2_p_spl_1,
    lo161_buf_o2_p_spl_
  );


  buf

  (
    lo161_buf_o2_p_spl_10,
    lo161_buf_o2_p_spl_1
  );


  buf

  (
    lo161_buf_o2_p_spl_11,
    lo161_buf_o2_p_spl_1
  );


  buf

  (
    lo161_buf_o2_n_spl_,
    lo161_buf_o2_n
  );


  buf

  (
    lo161_buf_o2_n_spl_0,
    lo161_buf_o2_n_spl_
  );


  buf

  (
    lo161_buf_o2_n_spl_00,
    lo161_buf_o2_n_spl_0
  );


  buf

  (
    lo161_buf_o2_n_spl_01,
    lo161_buf_o2_n_spl_0
  );


  buf

  (
    lo161_buf_o2_n_spl_1,
    lo161_buf_o2_n_spl_
  );


  buf

  (
    lo161_buf_o2_n_spl_10,
    lo161_buf_o2_n_spl_1
  );


  buf

  (
    lo161_buf_o2_n_spl_11,
    lo161_buf_o2_n_spl_1
  );


  buf

  (
    n584_o2_p_spl_,
    n584_o2_p
  );


  buf

  (
    n581_o2_n_spl_,
    n581_o2_n
  );


  buf

  (
    n584_o2_n_spl_,
    n584_o2_n
  );


  buf

  (
    n581_o2_p_spl_,
    n581_o2_p
  );


  buf

  (
    n593_o2_p_spl_,
    n593_o2_p
  );


  buf

  (
    n590_o2_n_spl_,
    n590_o2_n
  );


  buf

  (
    n593_o2_n_spl_,
    n593_o2_n
  );


  buf

  (
    n590_o2_p_spl_,
    n590_o2_p
  );


  buf

  (
    g446_p_spl_,
    g446_p
  );


  buf

  (
    g449_n_spl_,
    g449_n
  );


  buf

  (
    g446_n_spl_,
    g446_n
  );


  buf

  (
    g449_p_spl_,
    g449_p
  );


  buf

  (
    g443_n_spl_,
    g443_n
  );


  buf

  (
    g452_n_spl_,
    g452_n
  );


  buf

  (
    n608_o2_p_spl_,
    n608_o2_p
  );


  buf

  (
    n605_o2_n_spl_,
    n605_o2_n
  );


  buf

  (
    n608_o2_n_spl_,
    n608_o2_n
  );


  buf

  (
    n605_o2_p_spl_,
    n605_o2_p
  );


  buf

  (
    n621_o2_p_spl_,
    n621_o2_p
  );


  buf

  (
    n618_o2_n_spl_,
    n618_o2_n
  );


  buf

  (
    n621_o2_n_spl_,
    n621_o2_n
  );


  buf

  (
    n618_o2_p_spl_,
    n618_o2_p
  );


  buf

  (
    n630_o2_p_spl_,
    n630_o2_p
  );


  buf

  (
    n627_o2_n_spl_,
    n627_o2_n
  );


  buf

  (
    n630_o2_n_spl_,
    n630_o2_n
  );


  buf

  (
    n627_o2_p_spl_,
    n627_o2_p
  );


  buf

  (
    g464_p_spl_,
    g464_p
  );


  buf

  (
    g467_n_spl_,
    g467_n
  );


  buf

  (
    g464_n_spl_,
    g464_n
  );


  buf

  (
    g467_p_spl_,
    g467_p
  );


  buf

  (
    g461_n_spl_,
    g461_n
  );


  buf

  (
    g470_n_spl_,
    g470_n
  );


  buf

  (
    n665_o2_p_spl_,
    n665_o2_p
  );


  buf

  (
    n662_o2_n_spl_,
    n662_o2_n
  );


  buf

  (
    n665_o2_n_spl_,
    n665_o2_n
  );


  buf

  (
    n662_o2_p_spl_,
    n662_o2_p
  );


  buf

  (
    g479_n_spl_,
    g479_n
  );


  buf

  (
    g482_n_spl_,
    g482_n
  );


  buf

  (
    n645_o2_p_spl_,
    n645_o2_p
  );


  buf

  (
    n642_o2_n_spl_,
    n642_o2_n
  );


  buf

  (
    n645_o2_n_spl_,
    n645_o2_n
  );


  buf

  (
    n642_o2_p_spl_,
    n642_o2_p
  );


  buf

  (
    g491_n_spl_,
    g491_n
  );


  buf

  (
    g494_n_spl_,
    g494_n
  );


  buf

  (
    n770_o2_p_spl_,
    n770_o2_p
  );


  buf

  (
    n767_o2_n_spl_,
    n767_o2_n
  );


  buf

  (
    n770_o2_n_spl_,
    n770_o2_n
  );


  buf

  (
    n767_o2_p_spl_,
    n767_o2_p
  );


  buf

  (
    n708_o2_p_spl_,
    n708_o2_p
  );


  buf

  (
    n705_o2_n_spl_,
    n705_o2_n
  );


  buf

  (
    n708_o2_n_spl_,
    n708_o2_n
  );


  buf

  (
    n705_o2_p_spl_,
    n705_o2_p
  );


  buf

  (
    n745_o2_p_spl_,
    n745_o2_p
  );


  buf

  (
    n742_o2_n_spl_,
    n742_o2_n
  );


  buf

  (
    n745_o2_n_spl_,
    n745_o2_n
  );


  buf

  (
    n742_o2_p_spl_,
    n742_o2_p
  );


  buf

  (
    g506_p_spl_,
    g506_p
  );


  buf

  (
    g509_n_spl_,
    g509_n
  );


  buf

  (
    g506_n_spl_,
    g506_n
  );


  buf

  (
    g509_p_spl_,
    g509_p
  );


  buf

  (
    g503_n_spl_,
    g503_n
  );


  buf

  (
    g512_n_spl_,
    g512_n
  );


  buf

  (
    n789_o2_p_spl_,
    n789_o2_p
  );


  buf

  (
    n786_o2_n_spl_,
    n786_o2_n
  );


  buf

  (
    n789_o2_n_spl_,
    n789_o2_n
  );


  buf

  (
    n786_o2_p_spl_,
    n786_o2_p
  );


  buf

  (
    n717_o2_p_spl_,
    n717_o2_p
  );


  buf

  (
    n714_o2_n_spl_,
    n714_o2_n
  );


  buf

  (
    n717_o2_n_spl_,
    n717_o2_n
  );


  buf

  (
    n714_o2_p_spl_,
    n714_o2_p
  );


  buf

  (
    n754_o2_p_spl_,
    n754_o2_p
  );


  buf

  (
    n751_o2_n_spl_,
    n751_o2_n
  );


  buf

  (
    n754_o2_n_spl_,
    n754_o2_n
  );


  buf

  (
    n751_o2_p_spl_,
    n751_o2_p
  );


  buf

  (
    g524_p_spl_,
    g524_p
  );


  buf

  (
    g527_n_spl_,
    g527_n
  );


  buf

  (
    g524_n_spl_,
    g524_n
  );


  buf

  (
    g527_p_spl_,
    g527_p
  );


  buf

  (
    g521_n_spl_,
    g521_n
  );


  buf

  (
    g530_n_spl_,
    g530_n
  );


  buf

  (
    n695_o2_p_spl_,
    n695_o2_p
  );


  buf

  (
    n692_o2_n_spl_,
    n692_o2_n
  );


  buf

  (
    n695_o2_n_spl_,
    n695_o2_n
  );


  buf

  (
    n692_o2_p_spl_,
    n692_o2_p
  );


  buf

  (
    g539_n_spl_,
    g539_n
  );


  buf

  (
    g542_n_spl_,
    g542_n
  );


  buf

  (
    n732_o2_p_spl_,
    n732_o2_p
  );


  buf

  (
    n729_o2_n_spl_,
    n729_o2_n
  );


  buf

  (
    n732_o2_n_spl_,
    n732_o2_n
  );


  buf

  (
    n729_o2_p_spl_,
    n729_o2_p
  );


  buf

  (
    g551_n_spl_,
    g551_n
  );


  buf

  (
    g554_n_spl_,
    g554_n
  );


  buf

  (
    n621_lo_p_spl_,
    n621_lo_p
  );


  buf

  (
    n621_lo_p_spl_0,
    n621_lo_p_spl_
  );


  buf

  (
    n669_lo_p_spl_,
    n669_lo_p
  );


  buf

  (
    n669_lo_p_spl_0,
    n669_lo_p_spl_
  );


  buf

  (
    n621_lo_n_spl_,
    n621_lo_n
  );


  buf

  (
    n669_lo_n_spl_,
    n669_lo_n
  );


  buf

  (
    n633_lo_p_spl_,
    n633_lo_p
  );


  buf

  (
    n633_lo_p_spl_0,
    n633_lo_p_spl_
  );


  buf

  (
    n633_lo_n_spl_,
    n633_lo_n
  );


  buf

  (
    n681_lo_p_spl_,
    n681_lo_p
  );


  buf

  (
    n681_lo_p_spl_0,
    n681_lo_p_spl_
  );


  buf

  (
    n681_lo_n_spl_,
    n681_lo_n
  );


  buf

  (
    n645_lo_p_spl_,
    n645_lo_p
  );


  buf

  (
    n645_lo_p_spl_0,
    n645_lo_p_spl_
  );


  buf

  (
    n693_lo_p_spl_,
    n693_lo_p
  );


  buf

  (
    n693_lo_p_spl_0,
    n693_lo_p_spl_
  );


  buf

  (
    n645_lo_n_spl_,
    n645_lo_n
  );


  buf

  (
    n693_lo_n_spl_,
    n693_lo_n
  );


  buf

  (
    n657_lo_n_spl_,
    n657_lo_n
  );


  buf

  (
    n657_lo_p_spl_,
    n657_lo_p
  );


  buf

  (
    n657_lo_p_spl_0,
    n657_lo_p_spl_
  );


  buf

  (
    n705_lo_p_spl_,
    n705_lo_p
  );


  buf

  (
    n705_lo_p_spl_0,
    n705_lo_p_spl_
  );


  buf

  (
    n705_lo_n_spl_,
    n705_lo_n
  );


  buf

  (
    n717_lo_p_spl_,
    n717_lo_p
  );


  buf

  (
    n717_lo_p_spl_0,
    n717_lo_p_spl_
  );


  buf

  (
    n765_lo_n_spl_,
    n765_lo_n
  );


  buf

  (
    n717_lo_n_spl_,
    n717_lo_n
  );


  buf

  (
    n765_lo_p_spl_,
    n765_lo_p
  );


  buf

  (
    n765_lo_p_spl_0,
    n765_lo_p_spl_
  );


  buf

  (
    n729_lo_p_spl_,
    n729_lo_p
  );


  buf

  (
    n729_lo_p_spl_0,
    n729_lo_p_spl_
  );


  buf

  (
    n729_lo_n_spl_,
    n729_lo_n
  );


  buf

  (
    n777_lo_n_spl_,
    n777_lo_n
  );


  buf

  (
    n777_lo_p_spl_,
    n777_lo_p
  );


  buf

  (
    n777_lo_p_spl_0,
    n777_lo_p_spl_
  );


  buf

  (
    n741_lo_p_spl_,
    n741_lo_p
  );


  buf

  (
    n741_lo_p_spl_0,
    n741_lo_p_spl_
  );


  buf

  (
    n789_lo_n_spl_,
    n789_lo_n
  );


  buf

  (
    n741_lo_n_spl_,
    n741_lo_n
  );


  buf

  (
    n789_lo_p_spl_,
    n789_lo_p
  );


  buf

  (
    n789_lo_p_spl_0,
    n789_lo_p_spl_
  );


  buf

  (
    n753_lo_n_spl_,
    n753_lo_n
  );


  buf

  (
    n753_lo_p_spl_,
    n753_lo_p
  );


  buf

  (
    n753_lo_p_spl_0,
    n753_lo_p_spl_
  );


  buf

  (
    n801_lo_n_spl_,
    n801_lo_n
  );


  buf

  (
    n801_lo_p_spl_,
    n801_lo_p
  );


  buf

  (
    n801_lo_p_spl_0,
    n801_lo_p_spl_
  );


  buf

  (
    n813_lo_p_spl_,
    n813_lo_p
  );


  buf

  (
    n813_lo_p_spl_0,
    n813_lo_p_spl_
  );


  buf

  (
    n825_lo_p_spl_,
    n825_lo_p
  );


  buf

  (
    n825_lo_p_spl_0,
    n825_lo_p_spl_
  );


  buf

  (
    n813_lo_n_spl_,
    n813_lo_n
  );


  buf

  (
    n825_lo_n_spl_,
    n825_lo_n
  );


  buf

  (
    n861_lo_p_spl_,
    n861_lo_p
  );


  buf

  (
    n861_lo_p_spl_0,
    n861_lo_p_spl_
  );


  buf

  (
    n861_lo_n_spl_,
    n861_lo_n
  );


  buf

  (
    n873_lo_p_spl_,
    n873_lo_p
  );


  buf

  (
    n873_lo_p_spl_0,
    n873_lo_p_spl_
  );


  buf

  (
    n873_lo_n_spl_,
    n873_lo_n
  );


  buf

  (
    n837_lo_p_spl_,
    n837_lo_p
  );


  buf

  (
    n837_lo_p_spl_0,
    n837_lo_p_spl_
  );


  buf

  (
    n849_lo_n_spl_,
    n849_lo_n
  );


  buf

  (
    n837_lo_n_spl_,
    n837_lo_n
  );


  buf

  (
    n849_lo_p_spl_,
    n849_lo_p
  );


  buf

  (
    n849_lo_p_spl_0,
    n849_lo_p_spl_
  );


  buf

  (
    n885_lo_p_spl_,
    n885_lo_p
  );


  buf

  (
    n885_lo_p_spl_0,
    n885_lo_p_spl_
  );


  buf

  (
    n885_lo_n_spl_,
    n885_lo_n
  );


  buf

  (
    n897_lo_p_spl_,
    n897_lo_p
  );


  buf

  (
    n897_lo_p_spl_0,
    n897_lo_p_spl_
  );


  buf

  (
    n897_lo_n_spl_,
    n897_lo_n
  );


  buf

  (
    n909_lo_p_spl_,
    n909_lo_p
  );


  buf

  (
    n909_lo_p_spl_0,
    n909_lo_p_spl_
  );


  buf

  (
    n921_lo_p_spl_,
    n921_lo_p
  );


  buf

  (
    n921_lo_p_spl_0,
    n921_lo_p_spl_
  );


  buf

  (
    n909_lo_n_spl_,
    n909_lo_n
  );


  buf

  (
    n921_lo_n_spl_,
    n921_lo_n
  );


  buf

  (
    n957_lo_n_spl_,
    n957_lo_n
  );


  buf

  (
    n957_lo_p_spl_,
    n957_lo_p
  );


  buf

  (
    n957_lo_p_spl_0,
    n957_lo_p_spl_
  );


  buf

  (
    n969_lo_n_spl_,
    n969_lo_n
  );


  buf

  (
    n969_lo_p_spl_,
    n969_lo_p
  );


  buf

  (
    n969_lo_p_spl_0,
    n969_lo_p_spl_
  );


  buf

  (
    n933_lo_p_spl_,
    n933_lo_p
  );


  buf

  (
    n933_lo_p_spl_0,
    n933_lo_p_spl_
  );


  buf

  (
    n945_lo_n_spl_,
    n945_lo_n
  );


  buf

  (
    n933_lo_n_spl_,
    n933_lo_n
  );


  buf

  (
    n945_lo_p_spl_,
    n945_lo_p
  );


  buf

  (
    n945_lo_p_spl_0,
    n945_lo_p_spl_
  );


  buf

  (
    n981_lo_n_spl_,
    n981_lo_n
  );


  buf

  (
    n981_lo_p_spl_,
    n981_lo_p
  );


  buf

  (
    n981_lo_p_spl_0,
    n981_lo_p_spl_
  );


  buf

  (
    n993_lo_n_spl_,
    n993_lo_n
  );


  buf

  (
    n993_lo_p_spl_,
    n993_lo_p
  );


  buf

  (
    n993_lo_p_spl_0,
    n993_lo_p_spl_
  );


endmodule
