
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G426,
  G427,
  G428,
  G429,
  G430,
  G431,
  G432
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;
  output G426;output G427;output G428;output G429;output G430;output G431;output G432;
  wire new_n44_;wire new_n45_;wire new_n46_;wire new_n47_;wire new_n48_;wire new_n49_;wire new_n50_;wire new_n51_;wire new_n52_;wire new_n53_;wire new_n54_;wire new_n55_;wire new_n56_;wire new_n57_;wire new_n58_;wire new_n59_;wire new_n60_;wire new_n62_;wire new_n63_;wire new_n64_;wire new_n65_;wire new_n66_;wire new_n67_;wire new_n68_;wire new_n69_;wire new_n70_;wire new_n71_;wire new_n72_;wire new_n73_;wire new_n74_;wire new_n75_;wire new_n76_;wire new_n77_;wire new_n78_;wire new_n79_;wire new_n80_;wire new_n81_;wire new_n82_;wire new_n83_;wire new_n84_;wire new_n85_;wire new_n86_;wire new_n87_;wire new_n88_;wire new_n89_;wire new_n90_;wire new_n91_;wire new_n92_;wire new_n93_;wire new_n94_;wire new_n95_;wire new_n96_;wire new_n98_;wire new_n99_;wire new_n100_;wire new_n101_;wire new_n102_;wire new_n103_;wire new_n104_;wire new_n105_;wire new_n106_;wire new_n107_;wire new_n108_;wire new_n109_;wire new_n110_;wire new_n111_;wire new_n112_;wire new_n113_;wire new_n114_;wire new_n115_;wire new_n116_;wire new_n117_;wire new_n118_;wire new_n119_;wire new_n120_;wire new_n121_;wire new_n122_;wire new_n123_;wire new_n124_;wire new_n125_;wire new_n126_;wire new_n127_;wire new_n128_;wire new_n129_;wire new_n130_;wire new_n131_;wire new_n132_;wire new_n134_;wire new_n135_;wire new_n136_;wire new_n137_;wire new_n138_;wire new_n139_;wire new_n140_;wire new_n141_;wire new_n142_;wire new_n143_;wire new_n144_;wire new_n145_;wire new_n147_;wire new_n148_;wire new_n149_;wire new_n150_;wire new_n151_;wire new_n152_;wire new_n153_;wire new_n154_;wire new_n155_;wire new_n156_;wire new_n157_;wire new_n158_;wire new_n160_;wire new_n161_;wire new_n162_;wire new_n163_;wire new_n165_;wire new_n166_;wire new_n167_;wire new_n168_;
  wire G30_spl_;
  wire G28_spl_;
  wire G16_spl_;
  wire G18_spl_;
  wire G20_spl_;
  wire G22_spl_;
  wire G1_spl_;
  wire G2_spl_;
  wire G4_spl_;
  wire G6_spl_;
  wire G26_spl_;
  wire G24_spl_;
  wire G34_spl_;
  wire G32_spl_;
  wire G14_spl_;
  wire G12_spl_;
  wire G10_spl_;
  wire G8_spl_;
  wire new_n54__spl_;
  wire new_n59__spl_;
  wire new_n60__spl_;
  wire new_n60__spl_0;
  wire new_n60__spl_00;
  wire new_n60__spl_000;
  wire new_n60__spl_01;
  wire new_n60__spl_1;
  wire new_n60__spl_10;
  wire new_n60__spl_11;
  wire new_n63__spl_;
  wire G23_spl_;
  wire G11_spl_;
  wire new_n66__spl_;
  wire G3_spl_;
  wire new_n69__spl_;
  wire G7_spl_;
  wire new_n72__spl_;
  wire G31_spl_;
  wire new_n75__spl_;
  wire new_n78__spl_;
  wire G19_spl_;
  wire new_n81__spl_;
  wire G15_spl_;
  wire new_n84__spl_;
  wire G35_spl_;
  wire new_n87__spl_;
  wire G27_spl_;
  wire new_n90__spl_;
  wire new_n95__spl_;
  wire new_n96__spl_;
  wire new_n96__spl_0;
  wire new_n96__spl_00;
  wire new_n96__spl_000;
  wire new_n96__spl_01;
  wire new_n96__spl_1;
  wire new_n96__spl_10;
  wire new_n96__spl_11;
  wire new_n99__spl_;
  wire G25_spl_;
  wire G13_spl_;
  wire new_n102__spl_;
  wire G5_spl_;
  wire new_n105__spl_;
  wire G9_spl_;
  wire new_n108__spl_;
  wire G33_spl_;
  wire new_n111__spl_;
  wire new_n114__spl_;
  wire G21_spl_;
  wire new_n117__spl_;
  wire G17_spl_;
  wire new_n120__spl_;
  wire G36_spl_;
  wire new_n123__spl_;
  wire G29_spl_;
  wire new_n126__spl_;
  wire new_n131__spl_;
  wire new_n132__spl_;
  wire new_n132__spl_0;
  wire new_n132__spl_00;
  wire new_n132__spl_000;
  wire new_n132__spl_01;
  wire new_n132__spl_1;
  wire new_n132__spl_10;
  wire new_n132__spl_11;
  wire new_n137__spl_;
  wire new_n139__spl_;
  wire new_n139__spl_0;
  wire new_n144__spl_;
  wire new_n140__spl_;
  wire new_n145__spl_;
  wire new_n145__spl_0;
  wire new_n150__spl_;
  wire new_n153__spl_;
  wire new_n153__spl_0;
  wire new_n155__spl_;
  wire new_n161__spl_;

  anb1
  g000
  (
    .dina(G30_spl_),
    .dinb(G28_spl_),
    .dout(new_n44_)
  );


  anb2
  g001
  (
    .dina(G16_spl_),
    .dinb(G18_spl_),
    .dout(new_n45_)
  );


  anb2
  g002
  (
    .dina(G20_spl_),
    .dinb(G22_spl_),
    .dout(new_n46_)
  );


  anb2
  g003
  (
    .dina(G1_spl_),
    .dinb(G2_spl_),
    .dout(new_n47_)
  );


  anb2
  g004
  (
    .dina(G4_spl_),
    .dinb(G6_spl_),
    .dout(new_n48_)
  );


  anb1
  g005
  (
    .dina(G26_spl_),
    .dinb(G24_spl_),
    .dout(new_n49_)
  );


  anb1
  g006
  (
    .dina(G34_spl_),
    .dinb(G32_spl_),
    .dout(new_n50_)
  );


  anb1
  g007
  (
    .dina(G14_spl_),
    .dinb(G12_spl_),
    .dout(new_n51_)
  );


  anb1
  g008
  (
    .dina(G10_spl_),
    .dinb(G8_spl_),
    .dout(new_n52_)
  );


  anb1
  g009
  (
    .dina(new_n48_),
    .dinb(new_n49_),
    .dout(new_n53_)
  );


  anb2
  g010
  (
    .dina(new_n52_),
    .dinb(new_n53_),
    .dout(new_n54_)
  );


  anb1
  g011
  (
    .dina(new_n45_),
    .dinb(new_n51_),
    .dout(new_n55_)
  );


  anb2
  g012
  (
    .dina(new_n44_),
    .dinb(new_n47_),
    .dout(new_n56_)
  );


  anb1
  g013
  (
    .dina(new_n46_),
    .dinb(new_n50_),
    .dout(new_n57_)
  );


  anb2
  g014
  (
    .dina(new_n56_),
    .dinb(new_n57_),
    .dout(new_n58_)
  );


  anb1
  g015
  (
    .dina(new_n55_),
    .dinb(new_n58_),
    .dout(new_n59_)
  );


  nab1
  g016
  (
    .dina(new_n54__spl_),
    .dinb(new_n59__spl_),
    .dout(new_n60_)
  );


  anb2
  g017
  (
    .dina(new_n54__spl_),
    .dinb(new_n59__spl_),
    .dout(G426)
  );


  anb1
  g018
  (
    .dina(G20_spl_),
    .dinb(new_n60__spl_000),
    .dout(new_n62_)
  );


  anb1
  g019
  (
    .dina(G22_spl_),
    .dinb(new_n62_),
    .dout(new_n63_)
  );


  anb1
  g020
  (
    .dina(new_n63__spl_),
    .dinb(G23_spl_),
    .dout(new_n64_)
  );


  anb1
  g021
  (
    .dina(G8_spl_),
    .dinb(new_n60__spl_000),
    .dout(new_n65_)
  );


  anb1
  g022
  (
    .dina(G10_spl_),
    .dinb(new_n65_),
    .dout(new_n66_)
  );


  anb2
  g023
  (
    .dina(G11_spl_),
    .dinb(new_n66__spl_),
    .dout(new_n67_)
  );


  anb1
  g024
  (
    .dina(G1_spl_),
    .dinb(new_n60__spl_00),
    .dout(new_n68_)
  );


  anb1
  g025
  (
    .dina(G2_spl_),
    .dinb(new_n68_),
    .dout(new_n69_)
  );


  anb2
  g026
  (
    .dina(G3_spl_),
    .dinb(new_n69__spl_),
    .dout(new_n70_)
  );


  anb1
  g027
  (
    .dina(G4_spl_),
    .dinb(new_n60__spl_01),
    .dout(new_n71_)
  );


  anb1
  g028
  (
    .dina(G6_spl_),
    .dinb(new_n71_),
    .dout(new_n72_)
  );


  anb2
  g029
  (
    .dina(G7_spl_),
    .dinb(new_n72__spl_),
    .dout(new_n73_)
  );


  anb1
  g030
  (
    .dina(G28_spl_),
    .dinb(new_n60__spl_01),
    .dout(new_n74_)
  );


  anb1
  g031
  (
    .dina(G30_spl_),
    .dinb(new_n74_),
    .dout(new_n75_)
  );


  anb2
  g032
  (
    .dina(G31_spl_),
    .dinb(new_n75__spl_),
    .dout(new_n76_)
  );


  anb1
  g033
  (
    .dina(G16_spl_),
    .dinb(new_n60__spl_10),
    .dout(new_n77_)
  );


  anb1
  g034
  (
    .dina(G18_spl_),
    .dinb(new_n77_),
    .dout(new_n78_)
  );


  anb1
  g035
  (
    .dina(new_n78__spl_),
    .dinb(G19_spl_),
    .dout(new_n79_)
  );


  anb1
  g036
  (
    .dina(G12_spl_),
    .dinb(new_n60__spl_10),
    .dout(new_n80_)
  );


  anb1
  g037
  (
    .dina(G14_spl_),
    .dinb(new_n80_),
    .dout(new_n81_)
  );


  anb1
  g038
  (
    .dina(new_n81__spl_),
    .dinb(G15_spl_),
    .dout(new_n82_)
  );


  anb1
  g039
  (
    .dina(G32_spl_),
    .dinb(new_n60__spl_11),
    .dout(new_n83_)
  );


  anb1
  g040
  (
    .dina(G34_spl_),
    .dinb(new_n83_),
    .dout(new_n84_)
  );


  anb1
  g041
  (
    .dina(new_n84__spl_),
    .dinb(G35_spl_),
    .dout(new_n85_)
  );


  anb1
  g042
  (
    .dina(G24_spl_),
    .dinb(new_n60__spl_11),
    .dout(new_n86_)
  );


  anb1
  g043
  (
    .dina(G26_spl_),
    .dinb(new_n86_),
    .dout(new_n87_)
  );


  anb1
  g044
  (
    .dina(new_n87__spl_),
    .dinb(G27_spl_),
    .dout(new_n88_)
  );


  anb1
  g045
  (
    .dina(new_n76_),
    .dinb(new_n79_),
    .dout(new_n89_)
  );


  anb2
  g046
  (
    .dina(new_n88_),
    .dinb(new_n89_),
    .dout(new_n90_)
  );


  anb1
  g047
  (
    .dina(new_n67_),
    .dinb(new_n85_),
    .dout(new_n91_)
  );


  anb2
  g048
  (
    .dina(new_n64_),
    .dinb(new_n73_),
    .dout(new_n92_)
  );


  anb1
  g049
  (
    .dina(new_n70_),
    .dinb(new_n82_),
    .dout(new_n93_)
  );


  anb2
  g050
  (
    .dina(new_n92_),
    .dinb(new_n93_),
    .dout(new_n94_)
  );


  anb1
  g051
  (
    .dina(new_n91_),
    .dinb(new_n94_),
    .dout(new_n95_)
  );


  nab1
  g052
  (
    .dina(new_n90__spl_),
    .dinb(new_n95__spl_),
    .dout(new_n96_)
  );


  anb2
  g053
  (
    .dina(new_n90__spl_),
    .dinb(new_n95__spl_),
    .dout(G427)
  );


  anb1
  g054
  (
    .dina(G23_spl_),
    .dinb(new_n96__spl_000),
    .dout(new_n98_)
  );


  anb1
  g055
  (
    .dina(new_n63__spl_),
    .dinb(new_n98_),
    .dout(new_n99_)
  );


  anb1
  g056
  (
    .dina(new_n99__spl_),
    .dinb(G25_spl_),
    .dout(new_n100_)
  );


  anb1
  g057
  (
    .dina(G11_spl_),
    .dinb(new_n96__spl_000),
    .dout(new_n101_)
  );


  anb1
  g058
  (
    .dina(new_n66__spl_),
    .dinb(new_n101_),
    .dout(new_n102_)
  );


  anb2
  g059
  (
    .dina(G13_spl_),
    .dinb(new_n102__spl_),
    .dout(new_n103_)
  );


  anb1
  g060
  (
    .dina(G3_spl_),
    .dinb(new_n96__spl_00),
    .dout(new_n104_)
  );


  anb1
  g061
  (
    .dina(new_n69__spl_),
    .dinb(new_n104_),
    .dout(new_n105_)
  );


  anb2
  g062
  (
    .dina(G5_spl_),
    .dinb(new_n105__spl_),
    .dout(new_n106_)
  );


  anb1
  g063
  (
    .dina(G7_spl_),
    .dinb(new_n96__spl_01),
    .dout(new_n107_)
  );


  anb1
  g064
  (
    .dina(new_n72__spl_),
    .dinb(new_n107_),
    .dout(new_n108_)
  );


  anb2
  g065
  (
    .dina(G9_spl_),
    .dinb(new_n108__spl_),
    .dout(new_n109_)
  );


  anb1
  g066
  (
    .dina(G31_spl_),
    .dinb(new_n96__spl_01),
    .dout(new_n110_)
  );


  anb1
  g067
  (
    .dina(new_n75__spl_),
    .dinb(new_n110_),
    .dout(new_n111_)
  );


  anb2
  g068
  (
    .dina(G33_spl_),
    .dinb(new_n111__spl_),
    .dout(new_n112_)
  );


  anb1
  g069
  (
    .dina(G19_spl_),
    .dinb(new_n96__spl_10),
    .dout(new_n113_)
  );


  anb1
  g070
  (
    .dina(new_n78__spl_),
    .dinb(new_n113_),
    .dout(new_n114_)
  );


  anb1
  g071
  (
    .dina(new_n114__spl_),
    .dinb(G21_spl_),
    .dout(new_n115_)
  );


  anb1
  g072
  (
    .dina(G15_spl_),
    .dinb(new_n96__spl_10),
    .dout(new_n116_)
  );


  anb1
  g073
  (
    .dina(new_n81__spl_),
    .dinb(new_n116_),
    .dout(new_n117_)
  );


  anb1
  g074
  (
    .dina(new_n117__spl_),
    .dinb(G17_spl_),
    .dout(new_n118_)
  );


  anb1
  g075
  (
    .dina(G35_spl_),
    .dinb(new_n96__spl_11),
    .dout(new_n119_)
  );


  anb1
  g076
  (
    .dina(new_n84__spl_),
    .dinb(new_n119_),
    .dout(new_n120_)
  );


  anb1
  g077
  (
    .dina(new_n120__spl_),
    .dinb(G36_spl_),
    .dout(new_n121_)
  );


  anb1
  g078
  (
    .dina(G27_spl_),
    .dinb(new_n96__spl_11),
    .dout(new_n122_)
  );


  anb1
  g079
  (
    .dina(new_n87__spl_),
    .dinb(new_n122_),
    .dout(new_n123_)
  );


  anb1
  g080
  (
    .dina(new_n123__spl_),
    .dinb(G29_spl_),
    .dout(new_n124_)
  );


  anb1
  g081
  (
    .dina(new_n112_),
    .dinb(new_n115_),
    .dout(new_n125_)
  );


  anb2
  g082
  (
    .dina(new_n124_),
    .dinb(new_n125_),
    .dout(new_n126_)
  );


  anb1
  g083
  (
    .dina(new_n103_),
    .dinb(new_n121_),
    .dout(new_n127_)
  );


  anb2
  g084
  (
    .dina(new_n100_),
    .dinb(new_n109_),
    .dout(new_n128_)
  );


  anb1
  g085
  (
    .dina(new_n106_),
    .dinb(new_n118_),
    .dout(new_n129_)
  );


  anb2
  g086
  (
    .dina(new_n128_),
    .dinb(new_n129_),
    .dout(new_n130_)
  );


  anb1
  g087
  (
    .dina(new_n127_),
    .dinb(new_n130_),
    .dout(new_n131_)
  );


  nab1
  g088
  (
    .dina(new_n126__spl_),
    .dinb(new_n131__spl_),
    .dout(new_n132_)
  );


  anb2
  g089
  (
    .dina(new_n126__spl_),
    .dinb(new_n131__spl_),
    .dout(G428)
  );


  anb1
  g090
  (
    .dina(G5_spl_),
    .dinb(new_n132__spl_000),
    .dout(new_n134_)
  );


  anb2
  g091
  (
    .dina(new_n134_),
    .dinb(new_n105__spl_),
    .dout(new_n135_)
  );


  anb1
  g092
  (
    .dina(G9_spl_),
    .dinb(new_n132__spl_000),
    .dout(new_n136_)
  );


  anb2
  g093
  (
    .dina(new_n136_),
    .dinb(new_n108__spl_),
    .dout(new_n137_)
  );


  anb1
  g094
  (
    .dina(G13_spl_),
    .dinb(new_n132__spl_00),
    .dout(new_n138_)
  );


  anb1
  g095
  (
    .dina(new_n102__spl_),
    .dinb(new_n138_),
    .dout(new_n139_)
  );


  anb1
  g096
  (
    .dina(new_n137__spl_),
    .dinb(new_n139__spl_0),
    .dout(new_n140_)
  );


  anb1
  g097
  (
    .dina(G21_spl_),
    .dinb(new_n132__spl_01),
    .dout(new_n141_)
  );


  anb2
  g098
  (
    .dina(new_n141_),
    .dinb(new_n114__spl_),
    .dout(new_n142_)
  );


  anb1
  g099
  (
    .dina(G17_spl_),
    .dinb(new_n132__spl_01),
    .dout(new_n143_)
  );


  anb2
  g100
  (
    .dina(new_n143_),
    .dinb(new_n117__spl_),
    .dout(new_n144_)
  );


  and1
  g101
  (
    .dina(new_n142_),
    .dinb(new_n144__spl_),
    .dout(new_n145_)
  );


  nor2
  g102
  (
    .dina(new_n140__spl_),
    .dinb(new_n145__spl_0),
    .dout(G430)
  );


  anb1
  g103
  (
    .dina(G36_spl_),
    .dinb(new_n132__spl_10),
    .dout(new_n147_)
  );


  anb2
  g104
  (
    .dina(new_n147_),
    .dinb(new_n120__spl_),
    .dout(new_n148_)
  );


  anb1
  g105
  (
    .dina(G33_spl_),
    .dinb(new_n132__spl_10),
    .dout(new_n149_)
  );


  anb2
  g106
  (
    .dina(new_n149_),
    .dinb(new_n111__spl_),
    .dout(new_n150_)
  );


  and1
  g107
  (
    .dina(new_n148_),
    .dinb(new_n150__spl_),
    .dout(new_n151_)
  );


  anb1
  g108
  (
    .dina(G29_spl_),
    .dinb(new_n132__spl_11),
    .dout(new_n152_)
  );


  anb2
  g109
  (
    .dina(new_n152_),
    .dinb(new_n123__spl_),
    .dout(new_n153_)
  );


  anb1
  g110
  (
    .dina(G25_spl_),
    .dinb(new_n132__spl_11),
    .dout(new_n154_)
  );


  anb1
  g111
  (
    .dina(new_n99__spl_),
    .dinb(new_n154_),
    .dout(new_n155_)
  );


  nab2
  g112
  (
    .dina(new_n153__spl_0),
    .dinb(new_n155__spl_),
    .dout(new_n156_)
  );


  anb1
  g113
  (
    .dina(new_n151_),
    .dinb(new_n156_),
    .dout(new_n157_)
  );


  nab1
  g114
  (
    .dina(G430),
    .dinb(new_n157_),
    .dout(new_n158_)
  );


  anb1
  g115
  (
    .dina(new_n135_),
    .dinb(new_n158_),
    .dout(G429)
  );


  anb2
  g116
  (
    .dina(new_n139__spl_0),
    .dinb(new_n155__spl_),
    .dout(new_n160_)
  );


  anb1
  g117
  (
    .dina(new_n145__spl_0),
    .dinb(new_n160_),
    .dout(new_n161_)
  );


  anb1
  g118
  (
    .dina(new_n145__spl_),
    .dinb(new_n153__spl_0),
    .dout(new_n162_)
  );


  anb1
  g119
  (
    .dina(new_n140__spl_),
    .dinb(new_n162_),
    .dout(new_n163_)
  );


  anb2
  g120
  (
    .dina(new_n161__spl_),
    .dinb(new_n163_),
    .dout(G431)
  );


  anb1
  g121
  (
    .dina(new_n153__spl_),
    .dinb(new_n150__spl_),
    .dout(new_n165_)
  );


  nab2
  g122
  (
    .dina(new_n144__spl_),
    .dinb(new_n165_),
    .dout(new_n166_)
  );


  nab1
  g123
  (
    .dina(new_n139__spl_),
    .dinb(new_n166_),
    .dout(new_n167_)
  );


  anb1
  g124
  (
    .dina(new_n137__spl_),
    .dinb(new_n161__spl_),
    .dout(new_n168_)
  );


  anb2
  g125
  (
    .dina(new_n167_),
    .dinb(new_n168_),
    .dout(G432)
  );


  splt
  gG30
  (
    .dout(G30_spl_),
    .din(G30)
  );


  splt
  gG28
  (
    .dout(G28_spl_),
    .din(G28)
  );


  splt
  gG16
  (
    .dout(G16_spl_),
    .din(G16)
  );


  splt
  gG18
  (
    .dout(G18_spl_),
    .din(G18)
  );


  splt
  gG20
  (
    .dout(G20_spl_),
    .din(G20)
  );


  splt
  gG22
  (
    .dout(G22_spl_),
    .din(G22)
  );


  splt
  gG1
  (
    .dout(G1_spl_),
    .din(G1)
  );


  splt
  gG2
  (
    .dout(G2_spl_),
    .din(G2)
  );


  splt
  gG4
  (
    .dout(G4_spl_),
    .din(G4)
  );


  splt
  gG6
  (
    .dout(G6_spl_),
    .din(G6)
  );


  splt
  gG26
  (
    .dout(G26_spl_),
    .din(G26)
  );


  splt
  gG24
  (
    .dout(G24_spl_),
    .din(G24)
  );


  splt
  gG34
  (
    .dout(G34_spl_),
    .din(G34)
  );


  splt
  gG32
  (
    .dout(G32_spl_),
    .din(G32)
  );


  splt
  gG14
  (
    .dout(G14_spl_),
    .din(G14)
  );


  splt
  gG12
  (
    .dout(G12_spl_),
    .din(G12)
  );


  splt
  gG10
  (
    .dout(G10_spl_),
    .din(G10)
  );


  splt
  gG8
  (
    .dout(G8_spl_),
    .din(G8)
  );


  splt
  gnew_n54_
  (
    .dout(new_n54__spl_),
    .din(new_n54_)
  );


  splt
  gnew_n59_
  (
    .dout(new_n59__spl_),
    .din(new_n59_)
  );


  splt
  gnew_n60_
  (
    .dout(new_n60__spl_),
    .din(new_n60_)
  );


  splt
  gnew_n60__spl_
  (
    .dout(new_n60__spl_0),
    .din(new_n60__spl_)
  );


  splt
  gnew_n60__spl_0
  (
    .dout(new_n60__spl_00),
    .din(new_n60__spl_0)
  );


  splt
  gnew_n60__spl_00
  (
    .dout(new_n60__spl_000),
    .din(new_n60__spl_00)
  );


  splt
  gnew_n60__spl_0
  (
    .dout(new_n60__spl_01),
    .din(new_n60__spl_0)
  );


  splt
  gnew_n60__spl_
  (
    .dout(new_n60__spl_1),
    .din(new_n60__spl_)
  );


  splt
  gnew_n60__spl_1
  (
    .dout(new_n60__spl_10),
    .din(new_n60__spl_1)
  );


  splt
  gnew_n60__spl_1
  (
    .dout(new_n60__spl_11),
    .din(new_n60__spl_1)
  );


  splt
  gnew_n63_
  (
    .dout(new_n63__spl_),
    .din(new_n63_)
  );


  splt
  gG23
  (
    .dout(G23_spl_),
    .din(G23)
  );


  splt
  gG11
  (
    .dout(G11_spl_),
    .din(G11)
  );


  splt
  gnew_n66_
  (
    .dout(new_n66__spl_),
    .din(new_n66_)
  );


  splt
  gG3
  (
    .dout(G3_spl_),
    .din(G3)
  );


  splt
  gnew_n69_
  (
    .dout(new_n69__spl_),
    .din(new_n69_)
  );


  splt
  gG7
  (
    .dout(G7_spl_),
    .din(G7)
  );


  splt
  gnew_n72_
  (
    .dout(new_n72__spl_),
    .din(new_n72_)
  );


  splt
  gG31
  (
    .dout(G31_spl_),
    .din(G31)
  );


  splt
  gnew_n75_
  (
    .dout(new_n75__spl_),
    .din(new_n75_)
  );


  splt
  gnew_n78_
  (
    .dout(new_n78__spl_),
    .din(new_n78_)
  );


  splt
  gG19
  (
    .dout(G19_spl_),
    .din(G19)
  );


  splt
  gnew_n81_
  (
    .dout(new_n81__spl_),
    .din(new_n81_)
  );


  splt
  gG15
  (
    .dout(G15_spl_),
    .din(G15)
  );


  splt
  gnew_n84_
  (
    .dout(new_n84__spl_),
    .din(new_n84_)
  );


  splt
  gG35
  (
    .dout(G35_spl_),
    .din(G35)
  );


  splt
  gnew_n87_
  (
    .dout(new_n87__spl_),
    .din(new_n87_)
  );


  splt
  gG27
  (
    .dout(G27_spl_),
    .din(G27)
  );


  splt
  gnew_n90_
  (
    .dout(new_n90__spl_),
    .din(new_n90_)
  );


  splt
  gnew_n95_
  (
    .dout(new_n95__spl_),
    .din(new_n95_)
  );


  splt
  gnew_n96_
  (
    .dout(new_n96__spl_),
    .din(new_n96_)
  );


  splt
  gnew_n96__spl_
  (
    .dout(new_n96__spl_0),
    .din(new_n96__spl_)
  );


  splt
  gnew_n96__spl_0
  (
    .dout(new_n96__spl_00),
    .din(new_n96__spl_0)
  );


  splt
  gnew_n96__spl_00
  (
    .dout(new_n96__spl_000),
    .din(new_n96__spl_00)
  );


  splt
  gnew_n96__spl_0
  (
    .dout(new_n96__spl_01),
    .din(new_n96__spl_0)
  );


  splt
  gnew_n96__spl_
  (
    .dout(new_n96__spl_1),
    .din(new_n96__spl_)
  );


  splt
  gnew_n96__spl_1
  (
    .dout(new_n96__spl_10),
    .din(new_n96__spl_1)
  );


  splt
  gnew_n96__spl_1
  (
    .dout(new_n96__spl_11),
    .din(new_n96__spl_1)
  );


  splt
  gnew_n99_
  (
    .dout(new_n99__spl_),
    .din(new_n99_)
  );


  splt
  gG25
  (
    .dout(G25_spl_),
    .din(G25)
  );


  splt
  gG13
  (
    .dout(G13_spl_),
    .din(G13)
  );


  splt
  gnew_n102_
  (
    .dout(new_n102__spl_),
    .din(new_n102_)
  );


  splt
  gG5
  (
    .dout(G5_spl_),
    .din(G5)
  );


  splt
  gnew_n105_
  (
    .dout(new_n105__spl_),
    .din(new_n105_)
  );


  splt
  gG9
  (
    .dout(G9_spl_),
    .din(G9)
  );


  splt
  gnew_n108_
  (
    .dout(new_n108__spl_),
    .din(new_n108_)
  );


  splt
  gG33
  (
    .dout(G33_spl_),
    .din(G33)
  );


  splt
  gnew_n111_
  (
    .dout(new_n111__spl_),
    .din(new_n111_)
  );


  splt
  gnew_n114_
  (
    .dout(new_n114__spl_),
    .din(new_n114_)
  );


  splt
  gG21
  (
    .dout(G21_spl_),
    .din(G21)
  );


  splt
  gnew_n117_
  (
    .dout(new_n117__spl_),
    .din(new_n117_)
  );


  splt
  gG17
  (
    .dout(G17_spl_),
    .din(G17)
  );


  splt
  gnew_n120_
  (
    .dout(new_n120__spl_),
    .din(new_n120_)
  );


  splt
  gG36
  (
    .dout(G36_spl_),
    .din(G36)
  );


  splt
  gnew_n123_
  (
    .dout(new_n123__spl_),
    .din(new_n123_)
  );


  splt
  gG29
  (
    .dout(G29_spl_),
    .din(G29)
  );


  splt
  gnew_n126_
  (
    .dout(new_n126__spl_),
    .din(new_n126_)
  );


  splt
  gnew_n131_
  (
    .dout(new_n131__spl_),
    .din(new_n131_)
  );


  splt
  gnew_n132_
  (
    .dout(new_n132__spl_),
    .din(new_n132_)
  );


  splt
  gnew_n132__spl_
  (
    .dout(new_n132__spl_0),
    .din(new_n132__spl_)
  );


  splt
  gnew_n132__spl_0
  (
    .dout(new_n132__spl_00),
    .din(new_n132__spl_0)
  );


  splt
  gnew_n132__spl_00
  (
    .dout(new_n132__spl_000),
    .din(new_n132__spl_00)
  );


  splt
  gnew_n132__spl_0
  (
    .dout(new_n132__spl_01),
    .din(new_n132__spl_0)
  );


  splt
  gnew_n132__spl_
  (
    .dout(new_n132__spl_1),
    .din(new_n132__spl_)
  );


  splt
  gnew_n132__spl_1
  (
    .dout(new_n132__spl_10),
    .din(new_n132__spl_1)
  );


  splt
  gnew_n132__spl_1
  (
    .dout(new_n132__spl_11),
    .din(new_n132__spl_1)
  );


  splt
  gnew_n137_
  (
    .dout(new_n137__spl_),
    .din(new_n137_)
  );


  splt
  gnew_n139_
  (
    .dout(new_n139__spl_),
    .din(new_n139_)
  );


  splt
  gnew_n139__spl_
  (
    .dout(new_n139__spl_0),
    .din(new_n139__spl_)
  );


  splt
  gnew_n144_
  (
    .dout(new_n144__spl_),
    .din(new_n144_)
  );


  splt
  gnew_n140_
  (
    .dout(new_n140__spl_),
    .din(new_n140_)
  );


  splt
  gnew_n145_
  (
    .dout(new_n145__spl_),
    .din(new_n145_)
  );


  splt
  gnew_n145__spl_
  (
    .dout(new_n145__spl_0),
    .din(new_n145__spl_)
  );


  splt
  gnew_n150_
  (
    .dout(new_n150__spl_),
    .din(new_n150_)
  );


  splt
  gnew_n153_
  (
    .dout(new_n153__spl_),
    .din(new_n153_)
  );


  splt
  gnew_n153__spl_
  (
    .dout(new_n153__spl_0),
    .din(new_n153__spl_)
  );


  splt
  gnew_n155_
  (
    .dout(new_n155__spl_),
    .din(new_n155_)
  );


  splt
  gnew_n161_
  (
    .dout(new_n161__spl_),
    .din(new_n161_)
  );


endmodule
