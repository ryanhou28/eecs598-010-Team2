module c5315(G1,G10,G100,G101,G102,G103,G104,G105,G106,G107,G108,G109,G11,
  G110,G111,G112,G113,G114,G115,G116,G117,G118,G119,G12,G120,G121,G122,G123,
  G124,G125,G126,G127,G128,G129,G13,G130,G131,G132,G133,G134,G135,G136,G137,
  G138,G139,G14,G140,G141,G142,G143,G144,G145,G146,G147,G148,G149,G15,G150,
  G151,G152,G153,G154,G155,G156,G157,G158,G159,G16,G160,G161,G162,G163,G164,
  G165,G166,G167,G168,G169,G17,G170,G171,G172,G173,G174,G175,G176,G177,G178,
  G18,G19,G2,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G3,G30,G31,G32,G33,G34,
  G35,G36,G37,G38,G39,G4,G40,G41,G42,G43,G44,G45,G46,G47,G48,G49,G5,G50,G51,
  G5193,G5194,G5195,G5196,G5197,G5198,G5199,G52,G5200,G5201,G5202,G5203,G5204,
  G5205,G5206,G5207,G5208,G5209,G5210,G5211,G5212,G5213,G5214,G5215,G5216,
  G5217,G5218,G5219,G5220,G5221,G5222,G5223,G5224,G5225,G5226,G5227,G5228,
  G5229,G5230,G5231,G5232,G5233,G5234,G5235,G5236,G5237,G5238,G5239,G5240,
  G5241,G5242,G5243,G5244,G5245,G5246,G5247,G5248,G5249,G5250,G5251,G5252,
  G5253,G5254,G5255,G5256,G5257,G5258,G5259,G5260,G5261,G5262,G5263,G5264,
  G5265,G5266,G5267,G5268,G5269,G5270,G5271,G5272,G5273,G5274,G5275,G5276,
  G5277,G5278,G5279,G5280,G5281,G5282,G5283,G5284,G5285,G5286,G5287,G5288,
  G5289,G5290,G5291,G5292,G5293,G5294,G5295,G5296,G5297,G5298,G5299,G53,G5300,
  G5301,G5302,G5303,G5304,G5305,G5306,G5307,G5308,G5309,G5310,G5311,G5312,
  G5313,G5314,G5315,G54,G55,G56,G57,G58,G59,G6,G60,G61,G62,G63,G64,G65,G66,G67,
  G68,G69,G7,G70,G71,G72,G73,G74,G75,G76,G77,G78,G79,G8,G80,G81,G82,G83,G84,
  G85,G86,G87,G88,G89,G9,G90,G91,G92,G93,G94,G95,G96,G97,G98,G99);
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
  G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,
  G40,G41,G42,G43,G44,G45,G46,G47,G48,G49,G50,G51,G52,G53,G54,G55,G56,G57,G58,
  G59,G60,G61,G62,G63,G64,G65,G66,G67,G68,G69,G70,G71,G72,G73,G74,G75,G76,G77,
  G78,G79,G80,G81,G82,G83,G84,G85,G86,G87,G88,G89,G90,G91,G92,G93,G94,G95,G96,
  G97,G98,G99,G100,G101,G102,G103,G104,G105,G106,G107,G108,G109,G110,G111,G112,
  G113,G114,G115,G116,G117,G118,G119,G120,G121,G122,G123,G124,G125,G126,G127,
  G128,G129,G130,G131,G132,G133,G134,G135,G136,G137,G138,G139,G140,G141,G142,
  G143,G144,G145,G146,G147,G148,G149,G150,G151,G152,G153,G154,G155,G156,G157,
  G158,G159,G160,G161,G162,G163,G164,G165,G166,G167,G168,G169,G170,G171,G172,
  G173,G174,G175,G176,G177,G178;
output G5193,G5194,G5195,G5196,G5197,G5198,G5199,G5200,G5201,G5202,G5203,G5204,
  G5205,G5206,G5207,G5208,G5209,G5210,G5211,G5212,G5213,G5214,G5215,G5216,
  G5217,G5218,G5219,G5220,G5221,G5222,G5223,G5224,G5225,G5226,G5227,G5228,
  G5229,G5230,G5231,G5232,G5233,G5234,G5235,G5236,G5237,G5238,G5239,G5240,
  G5241,G5242,G5243,G5244,G5245,G5246,G5247,G5248,G5249,G5250,G5251,G5252,
  G5253,G5254,G5255,G5256,G5257,G5258,G5259,G5260,G5261,G5262,G5263,G5264,
  G5265,G5266,G5267,G5268,G5269,G5270,G5271,G5272,G5273,G5274,G5275,G5276,
  G5277,G5278,G5279,G5280,G5281,G5282,G5283,G5284,G5285,G5286,G5287,G5288,
  G5289,G5290,G5291,G5292,G5293,G5294,G5295,G5296,G5297,G5298,G5299,G5300,
  G5301,G5302,G5303,G5304,G5305,G5306,G5307,G5308,G5309,G5310,G5311,G5312,
  G5313,G5314,G5315;

  wire G632,G633,G634,G647,G659,G671,G684,G685,G686,G687,G688,G689,G690,G694,
    G706,G718,G730,G742,G746,G749,G752,G756,G768,G780,G792,G804,G813,G825,G836,
    G848,G860,G872,G884,G896,G908,G911,G914,G917,G920,G923,G926,G929,G932,G935,
    G938,G941,G944,G947,G950,G953,G956,G963,G970,G976,G980,G983,G993,G996,G999,
    G1002,G1005,G1008,G1011,G1014,G1017,G1020,G1023,G1026,G1029,G1032,G1035,
    G1038,G1041,G1044,G1047,G1050,G1053,G1060,G1067,G1070,G1075,G1081,G1084,
    G1087,G1090,G1093,G1096,G1099,G1102,G1105,G1108,G1111,G1114,G1117,G1120,
    G1123,G1126,G1129,G1132,G1135,G1138,G1141,G1144,G1147,G1150,G1162,G1172,
    G1184,G1196,G1208,G1214,G1218,G1230,G1242,G1245,G1248,G1256,G1264,G1272,
    G1280,G1287,G1294,G1301,G1308,G1311,G1314,G1317,G1320,G1323,G1326,G1329,
    G1332,G1335,G1338,G1341,G1344,G1347,G1350,G1353,G1356,G1359,G1362,G1365,
    G1368,G1371,G1374,G1377,G1380,G1383,G1386,G1389,G1392,G1395,G1398,G1401,
    G1404,G1407,G1410,G1413,G1416,G1419,G1422,G1425,G1428,G1431,G1434,G1437,
    G1440,G1443,G1446,G1449,G1452,G1455,G1458,G1459,G1460,G1461,G1462,G1463,
    G1464,G1465,G1466,G1467,G1468,G1469,G1470,G1471,G1472,G1473,G1474,G1475,
    G1476,G1477,G1478,G1479,G1480,G1481,G1482,G1483,G1484,G1485,G1486,G1487,
    G1488,G1489,G1490,G1491,G1492,G1493,G1494,G1495,G1496,G1497,G1498,G1499,
    G1500,G1501,G1502,G1503,G1504,G1505,G1506,G1507,G1508,G1509,G1510,G1511,
    G1512,G1513,G1514,G1515,G1516,G1517,G1518,G1519,G1520,G1526,G1537,G1548,
    G1554,G1565,G1576,G1577,G1582,G1583,G1584,G1585,G1586,G1587,G1588,G1589,
    G1590,G1591,G1592,G1593,G1594,G1595,G1601,G1612,G1623,G1629,G1640,G1651,
    G1652,G1663,G1674,G1685,G1696,G1697,G1698,G1699,G1700,G1701,G1702,G1703,
    G1704,G1705,G1706,G1707,G1708,G1709,G1710,G1711,G1712,G1713,G1714,G1715,
    G1716,G1717,G1718,G1719,G1720,G1721,G1722,G1723,G1724,G1725,G1726,G1727,
    G1728,G1734,G1740,G1741,G1742,G1743,G1744,G1745,G1746,G1747,G1748,G1749,
    G1750,G1755,G1764,G1774,G1775,G1776,G1777,G1778,G1779,G1780,G1781,G1782,
    G1783,G1784,G1785,G1786,G1787,G1788,G1789,G1790,G1791,G1792,G1793,G1794,
    G1795,G1796,G1797,G1798,G1799,G1800,G1801,G1802,G1803,G1804,G1805,G1806,
    G1807,G1808,G1809,G1810,G1811,G1812,G1813,G1814,G1815,G1821,G1827,G1828,
    G1829,G1830,G1831,G1832,G1833,G1834,G1835,G1836,G1837,G1842,G1843,G1844,
    G1845,G1846,G1847,G1848,G1849,G1850,G1851,G1852,G1853,G1854,G1855,G1856,
    G1857,G1858,G1859,G1860,G1861,G1862,G1863,G1864,G1865,G1866,G1867,G1868,
    G1869,G1870,G1871,G1872,G1873,G1876,G1879,G1880,G1883,G1886,G1887,G1888,
    G1889,G1890,G1891,G1892,G1893,G1894,G1895,G1896,G1897,G1898,G1899,G1900,
    G1901,G1902,G1903,G1904,G1905,G1906,G1907,G1908,G1911,G1914,G1925,G1936,
    G1941,G1944,G1945,G1946,G1947,G1948,G1959,G1970,G1981,G1992,G2003,G2014,
    G2015,G2016,G2017,G2018,G2019,G2020,G2031,G2042,G2053,G2064,G2067,G2068,
    G2069,G2070,G2071,G2072,G2073,G2076,G2077,G2078,G2079,G2080,G2081,G2082,
    G2083,G2084,G2085,G2086,G2087,G2088,G2089,G2090,G2091,G2092,G2093,G2094,
    G2095,G2096,G2097,G2098,G2099,G2100,G2101,G2102,G2103,G2104,G2105,G2108,
    G2109,G2110,G2111,G2112,G2113,G2114,G2115,G2116,G2117,G2118,G2119,G2120,
    G2121,G2122,G2123,G2124,G2125,G2126,G2127,G2128,G2129,G2130,G2131,G2132,
    G2133,G2134,G2135,G2136,G2137,G2138,G2139,G2140,G2141,G2142,G2143,G2144,
    G2145,G2146,G2147,G2148,G2149,G2150,G2151,G2152,G2153,G2154,G2155,G2156,
    G2157,G2158,G2159,G2160,G2161,G2162,G2163,G2164,G2165,G2166,G2167,G2168,
    G2169,G2170,G2171,G2172,G2173,G2174,G2175,G2176,G2177,G2178,G2179,G2180,
    G2181,G2182,G2183,G2184,G2185,G2186,G2187,G2188,G2189,G2190,G2191,G2192,
    G2193,G2194,G2195,G2196,G2197,G2198,G2199,G2200,G2201,G2202,G2203,G2204,
    G2205,G2206,G2207,G2208,G2209,G2210,G2211,G2212,G2213,G2214,G2215,G2216,
    G2217,G2218,G2219,G2220,G2221,G2222,G2223,G2224,G2225,G2226,G2227,G2228,
    G2229,G2230,G2231,G2240,G2241,G2242,G2243,G2244,G2245,G2248,G2249,G2250,
    G2251,G2252,G2253,G2254,G2255,G2256,G2257,G2258,G2259,G2260,G2261,G2262,
    G2263,G2264,G2265,G2266,G2267,G2268,G2269,G2270,G2271,G2277,G2278,G2279,
    G2280,G2281,G2282,G2283,G2284,G2285,G2286,G2287,G2288,G2289,G2290,G2291,
    G2292,G2293,G2294,G2295,G2296,G2297,G2298,G2299,G2300,G2301,G2302,G2303,
    G2304,G2305,G2306,G2307,G2308,G2309,G2310,G2314,G2318,G2319,G2320,G2321,
    G2322,G2323,G2324,G2325,G2326,G2327,G2328,G2332,G2336,G2339,G2340,G2341,
    G2342,G2343,G2344,G2345,G2346,G2347,G2348,G2349,G2352,G2355,G2358,G2361,
    G2362,G2363,G2366,G2367,G2368,G2369,G2370,G2371,G2372,G2373,G2374,G2375,
    G2376,G2377,G2378,G2379,G2386,G2392,G2398,G2404,G2410,G2418,G2424,G2430,
    G2436,G2437,G2438,G2441,G2442,G2443,G2444,G2445,G2446,G2447,G2448,G2454,
    G2460,G2466,G2472,G2480,G2486,G2492,G2499,G2500,G2501,G2502,G2503,G2504,
    G2505,G2506,G2507,G2508,G2511,G2512,G2513,G2514,G2515,G2516,G2517,G2520,
    G2523,G2526,G2527,G2528,G2529,G2530,G2531,G2532,G2533,G2534,G2535,G2536,
    G2537,G2538,G2539,G2540,G2543,G2547,G2550,G2553,G2556,G2559,G2562,G2565,
    G2568,G2571,G2574,G2577,G2580,G2583,G2586,G2589,G2590,G2591,G2592,G2593,
    G2596,G2599,G2600,G2601,G2602,G2603,G2606,G2609,G2612,G2615,G2618,G2621,
    G2624,G2625,G2626,G2629,G2632,G2635,G2638,G2641,G2644,G2647,G2650,G2653,
    G2656,G2659,G2662,G2663,G2666,G2667,G2668,G2669,G2670,G2671,G2672,G2673,
    G2674,G2675,G2679,G2685,G2692,G2693,G2696,G2700,G2705,G2711,G2715,G2720,
    G2726,G2727,G2731,G2737,G2744,G2752,G2759,G2770,G2774,G2780,G2787,G2788,
    G2792,G2797,G2804,G2810,G2817,G2828,G2832,G2837,G2843,G2844,G2850,G2857,
    G2865,G2872,G2875,G2876,G2877,G2878,G2879,G2883,G2887,G2888,G2891,G2894,
    G2897,G2900,G2903,G2906,G2909,G2912,G2915,G2918,G2921,G2924,G2927,G2930,
    G2933,G2936,G2939,G2942,G2945,G2948,G2951,G2954,G2957,G2960,G2963,G2966,
    G2969,G2972,G2975,G2978,G2981,G2984,G2987,G2990,G2993,G2996,G2999,G3002,
    G3005,G3008,G3011,G3014,G3017,G3020,G3023,G3026,G3029,G3032,G3035,G3038,
    G3039,G3040,G3041,G3042,G3043,G3044,G3045,G3046,G3047,G3048,G3049,G3050,
    G3051,G3052,G3053,G3054,G3055,G3056,G3057,G3058,G3059,G3060,G3063,G3064,
    G3065,G3066,G3067,G3068,G3069,G3070,G3071,G3072,G3073,G3074,G3075,G3076,
    G3077,G3078,G3079,G3080,G3081,G3082,G3083,G3084,G3085,G3086,G3087,G3088,
    G3089,G3090,G3091,G3092,G3093,G3094,G3097,G3098,G3099,G3100,G3101,G3102,
    G3103,G3104,G3105,G3106,G3107,G3108,G3109,G3110,G3111,G3112,G3113,G3114,
    G3115,G3116,G3117,G3118,G3119,G3120,G3121,G3122,G3123,G3124,G3125,G3126,
    G3127,G3128,G3129,G3130,G3131,G3132,G3133,G3134,G3135,G3136,G3137,G3138,
    G3139,G3140,G3141,G3142,G3143,G3144,G3145,G3146,G3147,G3148,G3149,G3150,
    G3151,G3152,G3153,G3154,G3155,G3156,G3157,G3158,G3159,G3160,G3161,G3162,
    G3163,G3164,G3165,G3166,G3167,G3168,G3169,G3170,G3171,G3172,G3173,G3174,
    G3175,G3176,G3177,G3178,G3179,G3180,G3181,G3182,G3183,G3184,G3185,G3186,
    G3187,G3188,G3189,G3190,G3191,G3192,G3195,G3196,G3197,G3198,G3199,G3202,
    G3203,G3204,G3205,G3206,G3207,G3208,G3211,G3214,G3215,G3218,G3219,G3222,
    G3225,G3228,G3231,G3234,G3237,G3240,G3241,G3244,G3247,G3250,G3253,G3256,
    G3259,G3262,G3265,G3266,G3267,G3268,G3269,G3270,G3271,G3272,G3273,G3274,
    G3275,G3276,G3277,G3280,G3281,G3282,G3283,G3284,G3285,G3286,G3287,G3288,
    G3289,G3290,G3291,G3292,G3293,G3294,G3295,G3296,G3297,G3298,G3299,G3300,
    G3301,G3302,G3303,G3313,G3314,G3315,G3316,G3317,G3331,G3332,G3333,G3334,
    G3335,G3336,G3337,G3338,G3339,G3340,G3341,G3342,G3343,G3344,G3348,G3351,
    G3355,G3358,G3359,G3360,G3363,G3364,G3365,G3366,G3367,G3368,G3369,G3370,
    G3371,G3374,G3377,G3380,G3383,G3386,G3393,G3404,G3415,G3421,G3428,G3438,
    G3449,G3459,G3466,G3467,G3474,G3485,G3495,G3503,G3517,G3533,G3546,G3552,
    G3559,G3570,G3576,G3583,G3594,G3604,G3605,G3606,G3607,G3608,G3609,G3610,
    G3611,G3621,G3629,G3645,G3658,G3664,G3665,G3666,G3670,G3674,G3677,G3681,
    G3685,G3688,G3689,G3690,G3691,G3692,G3693,G3694,G3695,G3696,G3697,G3700,
    G3703,G3706,G3709,G3710,G3713,G3714,G3715,G3716,G3717,G3718,G3719,G3720,
    G3723,G3726,G3729,G3732,G3735,G3738,G3739,G3742,G3745,G3748,G3751,G3752,
    G3753,G3754,G3755,G3756,G3757,G3758,G3759,G3760,G3761,G3762,G3763,G3764,
    G3765,G3768,G3769,G3770,G3771,G3772,G3773,G3774,G3775,G3776,G3779,G3780,
    G3781,G3782,G3783,G3784,G3785,G3786,G3787,G3788,G3789,G3790,G3791,G3792,
    G3793,G3796,G3797,G3798,G3799,G3800,G3801,G3802,G3805,G3806,G3807,G3808,
    G3809,G3810,G3811,G3812,G3813,G3814,G3815,G3816,G3817,G3818,G3819,G3820,
    G3821,G3822,G3823,G3824,G3825,G3828,G3829,G3830,G3831,G3832,G3833,G3834,
    G3837,G3838,G3839,G3840,G3841,G3842,G3843,G3844,G3845,G3846,G3847,G3848,
    G3849,G3852,G3855,G3856,G3857,G3858,G3859,G3862,G3863,G3864,G3865,G3866,
    G3867,G3868,G3869,G3870,G3871,G3872,G3873,G3874,G3875,G3876,G3877,G3878,
    G3879,G3882,G3885,G3888,G3891,G3894,G3897,G3900,G3903,G3904,G3905,G3906,
    G3909,G3912,G3915,G3918,G3921,G3924,G3927,G3930,G3933,G3936,G3939,G3942,
    G3945,G3948,G3951,G3954,G3957,G3960,G3963,G3966,G3969,G3972,G3975,G3978,
    G3981,G3984,G3987,G3990,G3993,G3996,G3999,G4002,G4005,G4008,G4011,G4014,
    G4017,G4020,G4023,G4026,G4029,G4032,G4035,G4038,G4039,G4040,G4041,G4042,
    G4043,G4044,G4045,G4046,G4047,G4048,G4051,G4054,G4058,G4061,G4064,G4065,
    G4068,G4072,G4075,G4076,G4077,G4080,G4081,G4082,G4083,G4084,G4085,G4086,
    G4087,G4088,G4089,G4092,G4095,G4098,G4101,G4104,G4107,G4110,G4113,G4116,
    G4119,G4122,G4125,G4128,G4131,G4134,G4137,G4140,G4143,G4146,G4149,G4152,
    G4155,G4158,G4161,G4164,G4167,G4170,G4173,G4174,G4175,G4176,G4177,G4180,
    G4183,G4184,G4185,G4186,G4187,G4188,G4189,G4190,G4191,G4192,G4193,G4194,
    G4195,G4196,G4197,G4198,G4199,G4200,G4201,G4202,G4203,G4204,G4205,G4206,
    G4207,G4208,G4209,G4210,G4211,G4212,G4213,G4214,G4215,G4216,G4217,G4218,
    G4219,G4220,G4221,G4222,G4223,G4224,G4225,G4226,G4227,G4230,G4231,G4232,
    G4233,G4234,G4235,G4236,G4237,G4238,G4239,G4240,G4241,G4242,G4243,G4244,
    G4245,G4246,G4247,G4248,G4249,G4250,G4251,G4252,G4253,G4254,G4257,G4260,
    G4261,G4262,G4263,G4264,G4265,G4266,G4267,G4268,G4269,G4270,G4271,G4272,
    G4273,G4274,G4275,G4276,G4282,G4283,G4284,G4285,G4286,G4287,G4288,G4289,
    G4290,G4293,G4294,G4295,G4296,G4297,G4298,G4299,G4300,G4301,G4302,G4303,
    G4309,G4310,G4311,G4312,G4313,G4314,G4315,G4316,G4319,G4320,G4321,G4322,
    G4323,G4329,G4330,G4331,G4332,G4333,G4334,G4335,G4336,G4339,G4340,G4343,
    G4344,G4345,G4346,G4349,G4350,G4351,G4352,G4355,G4356,G4359,G4360,G4363,
    G4364,G4367,G4368,G4369,G4370,G4371,G4374,G4375,G4376,G4377,G4378,G4381,
    G4382,G4383,G4384,G4385,G4386,G4387,G4388,G4389,G4390,G4391,G4392,G4393,
    G4394,G4395,G4396,G4397,G4398,G4399,G4400,G4403,G4404,G4405,G4406,G4407,
    G4408,G4409,G4413,G4414,G4415,G4416,G4417,G4420,G4423,G4424,G4425,G4426,
    G4427,G4428,G4429,G4430,G4431,G4432,G4437,G4440,G4443,G4446,G4449,G4450,
    G4453,G4454,G4455,G4456,G4457,G4458,G4463,G4466,G4469,G4472,G4473,G4476,
    G4477,G4478,G4479,G4480,G4483,G4484,G4487,G4488,G4489,G4490,G4491,G4492,
    G4493,G4494,G4497,G4498,G4501,G4504,G4507,G4508,G4509,G4510,G4511,G4512,
    G4513,G4514,G4515,G4516,G4517,G4518,G4519,G4520,G4521,G4522,G4523,G4524,
    G4525,G4526,G4527,G4528,G4529,G4530,G4531,G4532,G4533,G4534,G4535,G4536,
    G4537,G4538,G4539,G4540,G4541,G4542,G4543,G4544,G4545,G4546,G4547,G4548,
    G4549,G4550,G4551,G4552,G4553,G4554,G4560,G4561,G4562,G4568,G4569,G4570,
    G4571,G4572,G4573,G4576,G4579,G4580,G4581,G4582,G4583,G4586,G4589,G4592,
    G4593,G4594,G4597,G4600,G4603,G4606,G4613,G4616,G4619,G4622,G4623,G4624,
    G4630,G4636,G4642,G4648,G4654,G4655,G4658,G4664,G4670,G4671,G4672,G4673,
    G4674,G4675,G4676,G4677,G4678,G4679,G4680,G4681,G4684,G4687,G4690,G4691,
    G4692,G4693,G4694,G4697,G4700,G4701,G4702,G4703,G4704,G4705,G4706,G4709,
    G4710,G4711,G4712,G4713,G4714,G4715,G4716,G4717,G4718,G4719,G4720,G4721,
    G4722,G4723,G4724,G4725,G4726,G4727,G4728,G4729,G4730,G4731,G4732,G4733,
    G4734,G4735,G4736,G4737,G4738,G4739,G4740,G4741,G4742,G4743,G4744,G4745,
    G4746,G4747,G4748,G4749,G4750,G4751,G4752,G4753,G4754,G4755,G4756,G4757,
    G4758,G4761,G4762,G4763,G4764,G4765,G4766,G4767,G4768,G4769,G4770,G4771,
    G4772,G4773,G4774,G4775,G4776,G4777,G4778,G4779,G4780,G4786,G4792,G4798,
    G4804,G4810,G4816,G4822,G4828,G4831,G4834,G4835,G4836,G4837,G4838,G4841,
    G4844,G4847,G4848,G4849,G4850,G4851,G4852,G4853,G4854,G4855,G4856,G4857,
    G4858,G4859,G4860,G4861,G4862,G4863,G4864,G4865,G4866,G4867,G4868,G4869,
    G4870,G4871,G4872,G4873,G4874,G4875,G4876,G4877,G4878,G4879,G4880,G4881,
    G4882,G4883,G4884,G4885,G4886,G4887,G4888,G4889,G4890,G4891,G4892,G4895,
    G4898,G4899,G4900,G4901,G4902,G4903,G4904,G4907,G4908,G4909,G4910,G4911,
    G4912,G4913,G4914,G4915,G4916,G4917,G4918,G4919,G4920,G4923,G4926,G4927,
    G4928,G4929,G4930,G4933,G4936,G4939,G4940,G4941,G4942,G4943,G4944,G4945,
    G4946,G4947,G4948,G4951,G4954,G4955,G4956,G4957,G4958,G4959,G4960,G4963,
    G4964,G4965,G4966,G4967,G4968,G4971,G4974,G4975,G4976,G4977,G4978,G4981,
    G4984,G4987,G4988,G4989,G4990,G4991,G4992,G4993,G4994,G4995,G4996,G4999,
    G5002,G5003,G5004,G5005,G5006,G5007,G5008,G5011,G5012,G5013,G5014,G5015,
    G5016,G5019,G5022,G5023,G5024,G5025,G5026,G5029,G5032,G5035,G5036,G5037,
    G5038,G5039,G5040,G5041,G5042,G5043,G5044,G5045,G5046,G5047,G5048,G5051,
    G5054,G5055,G5056,G5059,G5060,G5061,G5062,G5063,G5064,G5067,G5070,G5073,
    G5076,G5077,G5078,G5079,G5080,G5083,G5084,G5085,G5086,G5087,G5088,G5089,
    G5090,G5091,G5092,G5093,G5094,G5095,G5096,G5097,G5098,G5101,G5104,G5107,
    G5108,G5111,G5114,G5115,G5116,G5117,G5118,G5119,G5120,G5121,G5122,G5123,
    G5124,G5125,G5126,G5127,G5128,G5129,G5130,G5131,G5132,G5133,G5134,G5135,
    G5138,G5141,G5142,G5143,G5144,G5145,G5146,G5147,G5150,G5153,G5154,G5155,
    G5156,G5157,G5158,G5159,G5162,G5165,G5166,G5167,G5168,G5169,G5172,G5175,
    G5178,G5181,G5182,G5183,G5184,G5185,G5186,G5187,G5188,G5189,G5190,G5191,
    G5192;

  and (G632,G62,G178);
  not (G633,G164);
  not (G634,G166);
  not (G647,G167);
  not (G659,G168);
  not (G671,G169);
  nand (G684,G134,G1);
  not (G685,G165);
  not (G686,G632);
  and (G687,G633,G11);
  and (G688,G136,G154);
  and (G689,G136,G155,G154,G153);
  not (G690,G157);
  not (G694,G158);
  not (G706,G159);
  not (G718,G158);
  not (G730,G159);
  not (G742,G64);
  not (G746,G64);
  not (G749,G66);
  not (G752,G162);
  not (G756,G160);
  not (G768,G161);
  not (G780,G160);
  not (G792,G161);
  not (G804,G102);
  not (G813,G101);
  not (G825,G101);
  not (G836,G100);
  not (G848,G100);
  not (G860,G173);
  not (G872,G172);
  not (G884,G174);
  not (G896,G175);
  not (G908,G90);
  not (G911,G90);
  not (G914,G92);
  not (G917,G92);
  not (G920,G94);
  not (G923,G94);
  not (G926,G96);
  not (G929,G96);
  not (G932,G103);
  not (G935,G103);
  not (G938,G105);
  not (G941,G105);
  not (G944,G107);
  not (G947,G107);
  not (G950,G109);
  not (G953,G109);
  not (G956,G124);
  not (G963,G124);
  not (G970,G88);
  and (G976,G11,G12);
  not (G980,G1);
  not (G983,G163);
  not (G993,G113);
  not (G996,G115);
  not (G999,G117);
  not (G1002,G117);
  not (G1005,G119);
  not (G1008,G119);
  not (G1011,G121);
  not (G1014,G121);
  not (G1017,G126);
  not (G1020,G126);
  not (G1023,G128);
  not (G1026,G128);
  not (G1029,G103);
  not (G1032,G103);
  not (G1035,G105);
  not (G1038,G105);
  not (G1041,G107);
  not (G1044,G107);
  not (G1047,G109);
  not (G1050,G109);
  not (G1053,G123);
  not (G1060,G123);
  not (G1067,G152);
  and (G1070,G12,G11);
  not (G1075,G163);
  not (G1081,G121);
  not (G1084,G121);
  not (G1087,G126);
  not (G1090,G126);
  not (G1093,G128);
  not (G1096,G128);
  not (G1099,G113);
  not (G1102,G115);
  not (G1105,G117);
  not (G1108,G117);
  not (G1111,G119);
  not (G1114,G119);
  not (G1117,G130);
  not (G1120,G130);
  not (G1123,G90);
  not (G1126,G90);
  not (G1129,G92);
  not (G1132,G92);
  not (G1135,G94);
  not (G1138,G94);
  not (G1141,G96);
  not (G1144,G96);
  not (G1147,G121);
  not (G1150,G98);
  not (G1162,G98);
  not (G1172,G102);
  not (G1184,G173);
  not (G1196,G172);
  not (G1208,G177);
  not (G1214,G176);
  not (G1218,G174);
  not (G1230,G175);
  not (G1242,G170);
  not (G1245,G171);
  not (G1248,G176);
  not (G1256,G177);
  not (G1264,G176);
  not (G1272,G177);
  not (G1280,G176);
  not (G1287,G177);
  not (G1294,G176);
  not (G1301,G177);
  not (G1308,G114);
  not (G1311,G142);
  not (G1314,G143);
  not (G1317,G144);
  not (G1320,G140);
  not (G1323,G141);
  not (G1326,G137);
  not (G1329,G138);
  not (G1332,G139);
  not (G1335,G135);
  not (G1338,G2);
  not (G1341,G142);
  not (G1344,G143);
  not (G1347,G144);
  not (G1350,G141);
  not (G1353,G137);
  not (G1356,G138);
  not (G1359,G139);
  not (G1362,G140);
  not (G1365,G135);
  not (G1368,G145);
  not (G1371,G146);
  not (G1374,G147);
  not (G1377,G148);
  not (G1380,G149);
  not (G1383,G150);
  not (G1386,G21);
  not (G1389,G145);
  not (G1392,G147);
  not (G1395,G148);
  not (G1398,G149);
  not (G1401,G150);
  not (G1404,G146);
  not (G1407,G130);
  not (G1410,G132);
  not (G1413,G126);
  not (G1416,G128);
  not (G1419,G117);
  not (G1422,G119);
  not (G1425,G113);
  not (G1428,G115);
  not (G1431,G109);
  not (G1434,G111);
  not (G1437,G105);
  not (G1440,G107);
  not (G1443,G96);
  not (G1446,G103);
  not (G1449,G92);
  not (G1452,G94);
  not (G1455,G90);
  and (G1458,G671,G148);
  or (G1459,G634,G148);
  and (G1460,G76,G694,G706);
  and (G1461,G77,G694,G706);
  and (G1462,G75,G694,G706);
  and (G1463,G74,G694,G706);
  and (G1464,G73,G694,G706);
  and (G1465,G81,G718,G730);
  and (G1466,G72,G718,G730);
  and (G1467,G70,G718,G730);
  and (G1468,G68,G718,G730);
  and (G1469,G76,G756,G768);
  and (G1470,G77,G756,G768);
  and (G1471,G75,G756,G768);
  and (G1472,G74,G756,G768);
  and (G1473,G73,G756,G768);
  and (G1474,G81,G780,G792);
  and (G1475,G72,G780,G792);
  and (G1476,G70,G780,G792);
  and (G1477,G68,G780,G792);
  and (G1478,G41,G1218,G1230);
  and (G1479,G22,G860,G872);
  and (G1480,G41,G1184,G1196);
  and (G1481,G18,G1184,G1196);
  and (G1482,G40,G1184,G1196);
  and (G1483,G15,G1184,G1196);
  and (G1484,G14,G1184,G1196);
  and (G1485,G6,G860,G872);
  and (G1486,G5,G860,G872);
  and (G1487,G25,G860,G872);
  and (G1488,G23,G860,G872);
  and (G1489,G18,G1218,G1230);
  and (G1490,G40,G1218,G1230);
  and (G1491,G15,G1218,G1230);
  and (G1492,G14,G1218,G1230);
  and (G1493,G6,G884,G896);
  and (G1494,G5,G884,G896);
  and (G1495,G25,G884,G896);
  and (G1496,G23,G884,G896);
  and (G1497,G54,G1245,G170);
  and (G1498,G1264,G1272);
  and (G1499,G22,G884,G896);
  and (G1500,G1248,G1256);
  not (G1501,G1311);
  not (G1502,G1314);
  not (G1503,G1317);
  not (G1504,G1320);
  not (G1505,G1323);
  not (G1506,G1326);
  not (G1507,G1329);
  not (G1508,G1332);
  not (G1509,G1335);
  not (G1510,G1338);
  not (G1511,G1341);
  not (G1512,G1344);
  not (G1513,G1347);
  not (G1514,G1350);
  not (G1515,G1353);
  not (G1516,G1356);
  not (G1517,G1359);
  not (G1518,G1362);
  not (G1519,G1365);
  not (G1520,G742);
  not (G1526,G694);
  not (G1537,G706);
  not (G1548,G742);
  not (G1554,G718);
  not (G1565,G730);
  and (G1576,G79,G718,G730);
  not (G1577,G980);
  not (G1582,G1368);
  not (G1583,G1371);
  not (G1584,G1374);
  not (G1585,G1377);
  not (G1586,G1380);
  not (G1587,G1383);
  not (G1588,G1386);
  not (G1589,G1389);
  not (G1590,G1392);
  not (G1591,G1395);
  not (G1592,G1398);
  not (G1593,G1401);
  not (G1594,G1404);
  not (G1595,G746);
  not (G1601,G756);
  not (G1612,G768);
  not (G1623,G746);
  not (G1629,G780);
  not (G1640,G792);
  and (G1651,G79,G780,G792);
  not (G1652,G860);
  not (G1663,G872);
  not (G1674,G884);
  not (G1685,G896);
  not (G1696,G908);
  not (G1697,G911);
  not (G1698,G914);
  not (G1699,G917);
  not (G1700,G920);
  not (G1701,G923);
  not (G1702,G926);
  not (G1703,G929);
  and (G1704,G671,G143,G911);
  and (G1705,G671,G144,G917);
  and (G1706,G671,G140,G923);
  and (G1707,G671,G141,G929);
  and (G1708,G634,G908);
  and (G1709,G634,G914);
  and (G1710,G634,G920);
  and (G1711,G634,G926);
  not (G1712,G932);
  not (G1713,G935);
  not (G1714,G938);
  not (G1715,G941);
  not (G1716,G944);
  not (G1717,G947);
  not (G1718,G950);
  not (G1719,G953);
  and (G1720,G671,G137,G935);
  and (G1721,G671,G138,G941);
  and (G1722,G671,G139,G947);
  and (G1723,G671,G135,G953);
  and (G1724,G634,G932);
  and (G1725,G634,G938);
  and (G1726,G634,G944);
  and (G1727,G634,G950);
  not (G1728,G956);
  not (G1734,G963);
  and (G1740,G112,G956);
  and (G1741,G110,G956);
  and (G1742,G108,G956);
  and (G1743,G106,G956);
  and (G1744,G104,G956);
  and (G1745,G97,G963);
  and (G1746,G95,G963);
  and (G1747,G93,G963);
  and (G1748,G91,G963);
  and (G1749,G89,G963);
  not (G1750,G749);
  not (G1755,G983);
  not (G1764,G976);
  not (G1774,G993);
  not (G1775,G996);
  not (G1776,G999);
  not (G1777,G1002);
  not (G1778,G1005);
  not (G1779,G1008);
  and (G1780,G836,G996);
  and (G1781,G836,G145,G1002);
  and (G1782,G836,G146,G1008);
  and (G1783,G1150,G993);
  and (G1784,G1150,G999);
  and (G1785,G1150,G1005);
  not (G1786,G1011);
  not (G1787,G1014);
  not (G1788,G1017);
  not (G1789,G1020);
  not (G1790,G1023);
  not (G1791,G1026);
  and (G1792,G671,G147,G1014);
  not (G1793,G1458);
  and (G1794,G671,G149,G1020);
  and (G1795,G671,G150,G1026);
  and (G1796,G634,G1011);
  and (G1797,G634,G1017);
  and (G1798,G634,G1023);
  not (G1799,G1029);
  not (G1800,G1032);
  not (G1801,G1035);
  not (G1802,G1038);
  not (G1803,G1041);
  not (G1804,G1044);
  not (G1805,G1047);
  not (G1806,G1050);
  and (G1807,G836,G137,G1032);
  and (G1808,G836,G138,G1038);
  and (G1809,G836,G139,G1044);
  and (G1810,G836,G135,G1050);
  and (G1811,G1150,G1029);
  and (G1812,G1150,G1035);
  and (G1813,G1150,G1041);
  and (G1814,G1150,G1047);
  not (G1815,G1053);
  not (G1821,G1060);
  and (G1827,G133,G1053);
  and (G1828,G131,G1053);
  and (G1829,G129,G1053);
  and (G1830,G127,G1053);
  and (G1831,G125,G1053);
  and (G1832,G122,G1060);
  and (G1833,G120,G1060);
  and (G1834,G118,G1060);
  and (G1835,G116,G1060);
  and (G1836,G114,G1060);
  not (G1837,G1075);
  and (G1842,G32,G1075);
  and (G1843,G33,G1075);
  and (G1844,G35,G1075);
  and (G1845,G35,G1075);
  not (G1846,G1081);
  not (G1847,G1084);
  not (G1848,G1087);
  not (G1849,G1090);
  not (G1850,G1093);
  not (G1851,G1096);
  and (G1852,G848,G147,G1084);
  and (G1853,G848,G148);
  and (G1854,G848,G149,G1090);
  and (G1855,G848,G150,G1096);
  and (G1856,G1162,G1081);
  or (G1857,G1162,G148);
  and (G1858,G1162,G1087);
  and (G1859,G1162,G1093);
  not (G1860,G1099);
  not (G1861,G1102);
  not (G1862,G1105);
  not (G1863,G1108);
  not (G1864,G1111);
  not (G1865,G1114);
  and (G1866,G848,G1102);
  and (G1867,G848,G145,G1108);
  and (G1868,G848,G146,G1114);
  and (G1869,G1162,G1099);
  and (G1870,G1162,G1105);
  and (G1871,G1162,G1111);
  not (G1872,G1117);
  not (G1873,G970);
  not (G1876,G970);
  not (G1879,G1120);
  not (G1880,G970);
  not (G1883,G970);
  and (G1886,G848,G1117);
  and (G1887,G848,G1120);
  not (G1888,G1123);
  not (G1889,G1126);
  not (G1890,G1129);
  not (G1891,G1132);
  not (G1892,G1135);
  not (G1893,G1138);
  not (G1894,G1141);
  not (G1895,G1144);
  and (G1896,G836,G143,G1126);
  and (G1897,G836,G144,G1132);
  and (G1898,G836,G140,G1138);
  and (G1899,G836,G141,G1144);
  and (G1900,G1150,G1123);
  and (G1901,G1150,G1129);
  and (G1902,G1150,G1135);
  and (G1903,G1150,G1141);
  not (G1904,G1407);
  not (G1905,G1410);
  not (G1906,G1413);
  not (G1907,G1416);
  not (G1908,G1147);
  not (G1911,G1147);
  not (G1914,G1184);
  not (G1925,G1196);
  not (G1936,G1208);
  not (G1941,G1214);
  and (G1944,G38,G1208);
  and (G1945,G37,G1208);
  and (G1946,G38,G1208);
  and (G1947,G37,G1208);
  not (G1948,G1218);
  not (G1959,G1230);
  not (G1970,G1248);
  not (G1981,G1256);
  not (G1992,G1264);
  not (G2003,G1272);
  not (G2014,G1431);
  not (G2015,G1434);
  not (G2016,G1437);
  not (G2017,G1440);
  not (G2018,G1443);
  not (G2019,G1446);
  not (G2020,G1280);
  not (G2031,G1287);
  not (G2042,G1294);
  not (G2053,G1301);
  not (G2064,G1308);
  not (G2067,G1419);
  not (G2068,G1422);
  not (G2069,G1425);
  not (G2070,G1428);
  not (G2071,G1449);
  not (G2072,G1452);
  not (G2073,G970);
  not (G2076,G1455);
  and (G2077,G143,G659,G1697);
  and (G2078,G144,G659,G1699);
  and (G2079,G140,G659,G1701);
  and (G2080,G141,G659,G1703);
  and (G2081,G647,G1696);
  and (G2082,G647,G1698);
  and (G2083,G647,G1700);
  and (G2084,G647,G1702);
  and (G2085,G137,G659,G1713);
  and (G2086,G138,G659,G1715);
  and (G2087,G139,G659,G1717);
  and (G2088,G135,G659,G1719);
  and (G2089,G647,G1712);
  and (G2090,G647,G1714);
  and (G2091,G647,G1716);
  and (G2092,G647,G1718);
  and (G2093,G813,G1775);
  and (G2094,G145,G813,G1777);
  and (G2095,G146,G813,G1779);
  and (G2096,G1172,G1774);
  and (G2097,G1172,G1776);
  and (G2098,G1172,G1778);
  and (G2099,G147,G659,G1787);
  and (G2100,G149,G659,G1789);
  and (G2101,G150,G659,G1791);
  and (G2102,G647,G1786);
  and (G2103,G647,G1788);
  and (G2104,G647,G1790);
  and (G2105,G1793,G1459);
  and (G2108,G137,G813,G1800);
  and (G2109,G138,G813,G1802);
  and (G2110,G139,G813,G1804);
  and (G2111,G135,G813,G1806);
  and (G2112,G1172,G1799);
  and (G2113,G1172,G1801);
  and (G2114,G1172,G1803);
  and (G2115,G1172,G1805);
  and (G2116,G147,G825,G1847);
  not (G2117,G1853);
  and (G2118,G149,G825,G1849);
  and (G2119,G150,G825,G1851);
  and (G2120,G804,G1846);
  and (G2121,G804,G1848);
  and (G2122,G804,G1850);
  and (G2123,G825,G1861);
  and (G2124,G145,G825,G1863);
  and (G2125,G146,G825,G1865);
  and (G2126,G804,G1860);
  and (G2127,G804,G1862);
  and (G2128,G804,G1864);
  and (G2129,G825,G1872);
  and (G2130,G825,G1879);
  and (G2131,G143,G813,G1889);
  and (G2132,G144,G813,G1891);
  and (G2133,G140,G813,G1893);
  and (G2134,G141,G813,G1895);
  and (G2135,G1172,G1888);
  and (G2136,G1172,G1890);
  and (G2137,G1172,G1892);
  and (G2138,G1172,G1894);
  nand (G2139,G1410,G1904);
  nand (G2140,G1407,G1905);
  nand (G2141,G1416,G1906);
  nand (G2142,G1413,G1907);
  nand (G2143,G1434,G2014);
  nand (G2144,G1431,G2015);
  nand (G2145,G1440,G2016);
  nand (G2146,G1437,G2017);
  nand (G2147,G1446,G2018);
  nand (G2148,G1443,G2019);
  nand (G2149,G1422,G2067);
  nand (G2150,G1419,G2068);
  nand (G2151,G1428,G2069);
  nand (G2152,G1425,G2070);
  nand (G2153,G1452,G2071);
  nand (G2154,G1449,G2072);
  and (G2155,G1755,G1764);
  and (G2156,G983,G1764);
  and (G2157,G86,G1526,G706);
  and (G2158,G87,G1526,G706);
  and (G2159,G85,G1526,G706);
  and (G2160,G84,G1526,G706);
  and (G2161,G83,G1526,G706);
  and (G2162,G80,G1554,G730);
  and (G2163,G82,G1554,G730);
  and (G2164,G71,G1554,G730);
  and (G2165,G69,G1554,G730);
  and (G2166,G1755,G1764);
  and (G2167,G983,G1764);
  and (G2168,G86,G1601,G768);
  and (G2169,G87,G1601,G768);
  and (G2170,G85,G1601,G768);
  and (G2171,G84,G1601,G768);
  and (G2172,G83,G1601,G768);
  and (G2173,G80,G1629,G792);
  and (G2174,G82,G1629,G792);
  and (G2175,G71,G1629,G792);
  and (G2176,G69,G1629,G792);
  and (G2177,G1755,G1764);
  and (G2178,G983,G1764);
  and (G2179,G42,G1948,G1230);
  and (G2180,G1755,G1764);
  and (G2181,G983,G1764);
  and (G2182,G3,G1652,G872);
  and (G2183,G42,G1914,G1196);
  and (G2184,G17,G1914,G1196);
  and (G2185,G39,G1914,G1196);
  and (G2186,G36,G1914,G1196);
  and (G2187,G16,G1914,G1196);
  and (G2188,G27,G1652,G872);
  and (G2189,G26,G1652,G872);
  and (G2190,G24,G1652,G872);
  and (G2191,G4,G1652,G872);
  and (G2192,G17,G1948,G1230);
  and (G2193,G39,G1948,G1230);
  and (G2194,G36,G1948,G1230);
  and (G2195,G16,G1948,G1230);
  and (G2196,G27,G1674,G896);
  and (G2197,G26,G1674,G896);
  and (G2198,G24,G1674,G896);
  and (G2199,G4,G1674,G896);
  and (G2200,G51,G1992,G1272);
  and (G2201,G3,G1674,G896);
  and (G2202,G49,G1970,G1256);
  and (G2203,G78,G1554,G730);
  and (G2204,G78,G1629,G792);
  or (G2205,G1704,G2077);
  or (G2206,G1705,G2078);
  or (G2207,G1706,G2079);
  or (G2208,G1707,G2080);
  or (G2209,G1708,G2081,G143);
  or (G2210,G1709,G2082,G144);
  or (G2211,G1710,G2083,G140);
  or (G2212,G1711,G2084,G141);
  or (G2213,G1720,G2085);
  or (G2214,G1721,G2086);
  or (G2215,G1722,G2087);
  or (G2216,G1723,G2088);
  or (G2217,G1724,G2089,G137);
  or (G2218,G1725,G2090,G138);
  or (G2219,G1726,G2091,G139);
  or (G2220,G1727,G2092,G135);
  and (G2221,G111,G1728);
  and (G2222,G109,G1728);
  and (G2223,G107,G1728);
  and (G2224,G105,G1728);
  and (G2225,G103,G1728);
  and (G2226,G96,G1734);
  and (G2227,G94,G1734);
  and (G2228,G92,G1734);
  and (G2229,G90,G1734);
  and (G2230,G88,G1734);
  not (G2231,G1764);
  or (G2240,G1780,G2093);
  or (G2241,G1781,G2094);
  or (G2242,G1782,G2095);
  or (G2243,G1784,G2097,G145);
  or (G2244,G1785,G2098,G146);
  or (G2245,G1783,G2096);
  or (G2248,G1792,G2099);
  or (G2249,G1794,G2100);
  or (G2250,G1795,G2101);
  or (G2251,G1796,G2102,G147);
  or (G2252,G1797,G2103,G149);
  or (G2253,G1798,G2104,G150);
  or (G2254,G1807,G2108);
  or (G2255,G1808,G2109);
  or (G2256,G1809,G2110);
  or (G2257,G1810,G2111);
  or (G2258,G1811,G2112,G137);
  or (G2259,G1812,G2113,G138);
  or (G2260,G1813,G2114,G139);
  or (G2261,G1814,G2115,G135);
  and (G2262,G132,G1815);
  and (G2263,G130,G1815);
  and (G2264,G128,G1815);
  and (G2265,G126,G1815);
  and (G2266,G121,G1821);
  and (G2267,G119,G1821);
  and (G2268,G117,G1821);
  and (G2269,G115,G1821);
  and (G2270,G113,G1821);
  or (G2271,G1815,G1831);
  and (G2277,G32,G1837);
  and (G2278,G34,G1837);
  and (G2279,G13,G1837);
  and (G2280,G13,G1837);
  or (G2281,G1852,G2116);
  or (G2282,G1854,G2118);
  or (G2283,G1855,G2119);
  or (G2284,G1856,G2120,G147);
  or (G2285,G1858,G2121,G149);
  or (G2286,G1859,G2122,G150);
  or (G2287,G1866,G2123);
  or (G2288,G1867,G2124);
  or (G2289,G1868,G2125);
  or (G2290,G1870,G2127,G145);
  or (G2291,G1871,G2128,G146);
  not (G2292,G1873);
  not (G2293,G1876);
  not (G2294,G1880);
  not (G2295,G1883);
  or (G2296,G1886,G2129);
  and (G2297,G848,G142,G1876);
  or (G2298,G1887,G2130);
  and (G2299,G848,G142,G1883);
  and (G2300,G1162,G1873);
  and (G2301,G1162,G1880);
  or (G2302,G1896,G2131);
  or (G2303,G1897,G2132);
  or (G2304,G1898,G2133);
  or (G2305,G1899,G2134);
  or (G2306,G1900,G2135,G143);
  or (G2307,G1901,G2136,G144);
  or (G2308,G1902,G2137,G140);
  or (G2309,G1903,G2138,G141);
  nand (G2310,G2139,G2140);
  nand (G2314,G2141,G2142);
  not (G2318,G1908);
  not (G2319,G1911);
  and (G2320,G48,G1970,G1256);
  and (G2321,G55,G1970,G1256);
  and (G2322,G56,G1970,G1256);
  and (G2323,G57,G1970,G1256);
  and (G2324,G60,G1992,G1272);
  and (G2325,G58,G1992,G1272);
  and (G2326,G50,G1992,G1272);
  and (G2327,G59,G1992,G1272);
  nand (G2328,G2143,G2144);
  nand (G2332,G2145,G2146);
  nand (G2336,G2147,G2148);
  and (G2339,G53,G2020,G1287);
  and (G2340,G44,G2020,G1287);
  and (G2341,G20,G2020,G1287);
  and (G2342,G45,G2020,G1287);
  and (G2343,G46,G2020,G1287);
  and (G2344,G19,G2042,G1301);
  and (G2345,G43,G2042,G1301);
  and (G2346,G47,G2042,G1301);
  and (G2347,G52,G2042,G1301);
  and (G2348,G54,G2042,G1301);
  nand (G2349,G2151,G2152);
  nand (G2352,G2149,G2150);
  and (G2355,G2117,G1857);
  or (G2358,G1869,G2126);
  not (G2361,G2073);
  nand (G2362,G2073,G2076);
  nand (G2363,G2153,G2154);
  not (G2366,G2105);
  or (G2367,G2278,G1843);
  or (G2368,G2279,G1844);
  or (G2369,G2280,G1845);
  or (G2370,G2277,G1842);
  not (G2371,G2205);
  not (G2372,G2206);
  not (G2373,G2207);
  not (G2374,G2208);
  not (G2375,G2213);
  not (G2376,G2214);
  not (G2377,G2215);
  not (G2378,G2216);
  or (G2379,G2222,G1741);
  or (G2386,G2223,G1742);
  or (G2392,G2224,G1743);
  or (G2398,G2225,G1744);
  or (G2404,G2226,G1745);
  or (G2410,G2227,G1746);
  or (G2418,G2228,G1747);
  or (G2424,G2229,G1748);
  or (G2430,G2230,G1749);
  not (G2436,G2241);
  not (G2437,G2242);
  not (G2438,G2240);
  not (G2441,G2248);
  not (G2442,G2249);
  not (G2443,G2250);
  not (G2444,G2254);
  not (G2445,G2255);
  not (G2446,G2256);
  not (G2447,G2257);
  or (G2448,G2263,G1828);
  or (G2454,G2264,G1829);
  or (G2460,G2265,G1830);
  or (G2466,G2266,G1832);
  or (G2472,G2267,G1833);
  or (G2480,G2268,G1834);
  or (G2486,G2269,G1835);
  or (G2492,G2270,G1836);
  not (G2499,G2281);
  not (G2500,G2282);
  not (G2501,G2283);
  not (G2502,G2288);
  not (G2503,G2289);
  and (G2504,G142,G825,G2293);
  and (G2505,G142,G825,G2295);
  and (G2506,G804,G2292);
  and (G2507,G804,G2294);
  not (G2508,G2296);
  not (G2511,G2298);
  not (G2512,G2302);
  not (G2513,G2303);
  not (G2514,G2304);
  not (G2515,G2305);
  and (G2516,G2105,G1992,G2003);
  or (G2517,G2262,G1827);
  or (G2520,G2221,G1740);
  not (G2523,G2287);
  nand (G2526,G1455,G2361);
  not (G2527,G2245);
  and (G2528,G2367,G1070);
  and (G2529,G8,G1755,G2231);
  and (G2530,G9,G983,G2231);
  and (G2531,G10,G1755,G2231);
  and (G2532,G30,G983,G2231);
  and (G2533,G2368,G1070);
  and (G2534,G28,G1755,G2231);
  and (G2535,G7,G983,G2231);
  and (G2536,G31,G1755,G2231);
  and (G2537,G29,G983,G2231);
  and (G2538,G2369,G1070);
  and (G2539,G2370,G1070);
  and (G2540,G2271,G148);
  and (G2543,G148,G2271);
  and (G2547,G2371,G2209);
  and (G2550,G2372,G2210);
  and (G2553,G2373,G2211);
  and (G2556,G2374,G2212);
  and (G2559,G2375,G2217);
  and (G2562,G2376,G2218);
  and (G2565,G2377,G2219);
  and (G2568,G2378,G2220);
  and (G2571,G2436,G2243);
  and (G2574,G2437,G2244);
  not (G2577,G2245);
  and (G2580,G2441,G2251);
  and (G2583,G2442,G2252);
  and (G2586,G2443,G2253);
  or (G2589,G2297,G2504);
  or (G2590,G2299,G2505);
  or (G2591,G2300,G2506,G142);
  or (G2592,G2301,G2507,G142);
  not (G2593,G2310);
  not (G2596,G2314);
  and (G2599,G2314,G2310,G1908);
  and (G2600,G2511,G1992,G2003);
  and (G2601,G2447,G2261);
  not (G2602,G2355);
  not (G2603,G2328);
  not (G2606,G2332);
  not (G2609,G2336);
  not (G2612,G2336);
  not (G2615,G2271);
  not (G2618,G2271);
  not (G2621,G2271);
  not (G2624,G2349);
  not (G2625,G2352);
  and (G2626,G2445,G2259);
  and (G2629,G2446,G2260);
  and (G2632,G2515,G2309);
  and (G2635,G2444,G2258);
  and (G2638,G2513,G2307);
  and (G2641,G2514,G2308);
  and (G2644,G2512,G2306);
  and (G2647,G2500,G2285);
  and (G2650,G2501,G2286);
  and (G2653,G2499,G2284);
  and (G2656,G2502,G2290);
  and (G2659,G2503,G2291);
  not (G2662,G2358);
  nand (G2663,G2526,G2362);
  not (G2666,G2363);
  and (G2667,G142,G2430);
  not (G2668,G2438);
  not (G2669,G2508);
  and (G2670,G2430,G142);
  or (G2671,G2529,G2530,G2155,G2156);
  or (G2672,G2531,G2532,G2166,G2167);
  or (G2673,G2534,G2535,G2177,G2178);
  or (G2674,G2536,G2537,G2180,G2181);
  and (G2675,G2424,G143);
  and (G2679,G2418,G144);
  and (G2685,G140,G2410);
  and (G2692,G2404,G141);
  and (G2693,G2398,G137);
  and (G2696,G2392,G138);
  and (G2700,G2386,G139);
  and (G2705,G2379,G135);
  and (G2711,G143,G2424);
  and (G2715,G144,G2418);
  and (G2720,G140,G2410);
  and (G2726,G141,G2404);
  and (G2727,G137,G2398);
  and (G2731,G138,G2392);
  and (G2737,G139,G2386);
  and (G2744,G135,G2379);
  not (G2752,G2492);
  not (G2759,G2486);
  not (G2770,G2486);
  and (G2774,G2480,G145);
  and (G2780,G146,G2472);
  and (G2787,G2466,G147);
  and (G2788,G2460,G149);
  and (G2792,G2454,G150);
  not (G2797,G2448);
  not (G2804,G2448);
  not (G2810,G2492);
  not (G2817,G2486);
  not (G2828,G2486);
  and (G2832,G145,G2480);
  and (G2837,G146,G2472);
  and (G2843,G147,G2466);
  and (G2844,G149,G2460);
  and (G2850,G150,G2454);
  not (G2857,G2448);
  not (G2865,G2448);
  not (G2872,G2492);
  not (G2875,G2589);
  not (G2876,G2590);
  not (G2877,G2517);
  not (G2878,G2520);
  not (G2879,G2601);
  not (G2883,G2508);
  and (G2887,G2438,G2042,G2053);
  not (G2888,G2430);
  not (G2891,G2424);
  not (G2894,G2418);
  not (G2897,G2410);
  not (G2900,G2404);
  not (G2903,G2398);
  not (G2906,G2392);
  not (G2909,G2386);
  not (G2912,G2379);
  nor (G2915,G140,G2410);
  not (G2918,G2430);
  not (G2921,G2424);
  not (G2924,G2418);
  not (G2927,G2404);
  not (G2930,G2398);
  not (G2933,G2392);
  not (G2936,G2386);
  not (G2939,G2410);
  not (G2942,G2379);
  nor (G2945,G140,G2410);
  nor (G2948,G135,G2379);
  not (G2951,G2480);
  not (G2954,G2472);
  not (G2957,G2466);
  not (G2960,G2460);
  not (G2963,G2454);
  nor (G2966,G146,G2472);
  not (G2969,G2480);
  not (G2972,G2466);
  not (G2975,G2460);
  not (G2978,G2454);
  not (G2981,G2472);
  nor (G2984,G146,G2472);
  not (G2987,G2454);
  not (G2990,G2460);
  not (G2993,G2448);
  not (G2996,G2466);
  not (G2999,G2480);
  not (G3002,G2472);
  not (G3005,G2492);
  not (G3008,G2486);
  not (G3011,G2410);
  not (G3014,G2404);
  not (G3017,G2424);
  not (G3020,G2418);
  not (G3023,G2430);
  not (G3026,G2386);
  not (G3029,G2379);
  not (G3032,G2398);
  not (G3035,G2392);
  nand (G3038,G2352,G2624);
  nand (G3039,G2349,G2625);
  not (G3040,G2523);
  nand (G3041,G2523,G2662);
  not (G3042,G2574);
  not (G3043,G2571);
  not (G3044,G2586);
  not (G3045,G2583);
  not (G3046,G2580);
  not (G3047,G2556);
  not (G3048,G2553);
  not (G3049,G2550);
  not (G3050,G2547);
  not (G3051,G2568);
  not (G3052,G2565);
  not (G3053,G2562);
  not (G3054,G2559);
  and (G3055,G2577,G1245,G1242);
  not (G3056,G2615);
  nand (G3057,G2615,G1585);
  nand (G3058,G2618,G1591);
  not (G3059,G2618);
  and (G3060,G2875,G2591);
  and (G3063,G2876,G2592);
  not (G3064,G2621);
  and (G3065,G2593,G2314,G2318);
  and (G3066,G2310,G2596,G2319);
  and (G3067,G2596,G2593,G1911);
  and (G3068,G2568,G1970,G1981);
  and (G3069,G2565,G1970,G1981);
  and (G3070,G2562,G1970,G1981);
  and (G3071,G2559,G1970,G1981);
  and (G3072,G2586,G1992,G2003);
  and (G3073,G2583,G1992,G2003);
  not (G3074,G2626);
  not (G3075,G2629);
  not (G3076,G2632);
  not (G3077,G2635);
  not (G3078,G2647);
  not (G3079,G2650);
  not (G3080,G2653);
  nand (G3081,G2653,G2602);
  not (G3082,G2609);
  not (G3083,G2612);
  and (G3084,G2332,G2328,G2609);
  and (G3085,G2606,G2603,G2612);
  and (G3086,G2556,G2020,G2031);
  and (G3087,G2553,G2020,G2031);
  and (G3088,G2550,G2020,G2031);
  and (G3089,G2547,G2020,G2031);
  and (G3090,G2580,G2042,G2053);
  and (G3091,G2574,G2042,G2053);
  and (G3092,G2571,G2042,G2053);
  and (G3093,G2577,G2042,G2053);
  nand (G3094,G3038,G3039);
  not (G3097,G2638);
  not (G3098,G2641);
  not (G3099,G2644);
  not (G3100,G2656);
  not (G3101,G2659);
  nand (G3102,G2358,G3040);
  not (G3103,G2663);
  nand (G3104,G2663,G2666);
  and (G3105,G3042,G3043,G2668,G2527);
  and (G3106,G3044,G3045,G2366,G3046);
  and (G3107,G3047,G3048,G3049,G3050);
  and (G3108,G3051,G3052,G3053,G3054);
  and (G3109,G2752,G2770);
  and (G3110,G2759,G2752,G2774);
  and (G3111,G2810,G2828);
  and (G3112,G2817,G2810,G2832);
  not (G3113,G2888);
  nand (G3114,G2888,G1501);
  not (G3115,G2891);
  nand (G3116,G2891,G1502);
  not (G3117,G2894);
  nand (G3118,G2894,G1503);
  not (G3119,G2897);
  nand (G3120,G2897,G1504);
  not (G3121,G2900);
  nand (G3122,G2900,G1505);
  not (G3123,G2903);
  nand (G3124,G2903,G1506);
  not (G3125,G2906);
  nand (G3126,G2906,G1507);
  not (G3127,G2909);
  nand (G3128,G2909,G1508);
  not (G3129,G2912);
  nand (G3130,G2912,G1509);
  not (G3131,G2915);
  nand (G3132,G2918,G1511);
  not (G3133,G2918);
  nand (G3134,G2921,G1512);
  not (G3135,G2921);
  nand (G3136,G2924,G1513);
  not (G3137,G2924);
  nand (G3138,G2927,G1514);
  not (G3139,G2927);
  nand (G3140,G2930,G1515);
  not (G3141,G2930);
  nand (G3142,G2933,G1516);
  not (G3143,G2933);
  nand (G3144,G2936,G1517);
  not (G3145,G2936);
  nand (G3146,G2939,G1518);
  not (G3147,G2939);
  nand (G3148,G2942,G1519);
  not (G3149,G2942);
  not (G3150,G2951);
  nand (G3151,G2951,G1582);
  not (G3152,G2954);
  nand (G3153,G2954,G1583);
  not (G3154,G2957);
  nand (G3155,G2957,G1584);
  nand (G3156,G1377,G3056);
  not (G3157,G2960);
  nand (G3158,G2960,G1586);
  not (G3159,G2963);
  nand (G3160,G2963,G1587);
  and (G3161,G2759,G2774);
  and (G3162,G2759,G2774);
  and (G3163,G21,G2797);
  not (G3164,G2966);
  nand (G3165,G2969,G1589);
  not (G3166,G2969);
  nand (G3167,G2972,G1590);
  not (G3168,G2972);
  nand (G3169,G1395,G3059);
  nand (G3170,G2975,G1592);
  not (G3171,G2975);
  nand (G3172,G2978,G1593);
  not (G3173,G2978);
  nand (G3174,G2981,G1594);
  not (G3175,G2981);
  and (G3176,G2817,G2832);
  and (G3177,G2817,G2832);
  not (G3178,G2987);
  not (G3179,G2990);
  nand (G3180,G2993,G2877);
  not (G3181,G2993);
  not (G3182,G2996);
  nand (G3183,G2996,G3064);
  not (G3184,G3011);
  not (G3185,G3014);
  not (G3186,G3017);
  not (G3187,G3020);
  nand (G3188,G3023,G2878);
  not (G3189,G3023);
  nor (G3190,G3065,G2599);
  nor (G3191,G3066,G3067);
  not (G3192,G2879);
  nand (G3195,G2629,G3074);
  nand (G3196,G2626,G3075);
  nand (G3197,G2635,G3076);
  nand (G3198,G2632,G3077);
  not (G3199,G2883);
  nand (G3202,G2650,G3078);
  nand (G3203,G2647,G3079);
  nand (G3204,G2355,G3080);
  and (G3205,G2603,G2332,G3082);
  and (G3206,G2328,G2606,G3083);
  and (G3207,G3063,G2020,G2031);
  not (G3208,G2872);
  not (G3211,G2685);
  not (G3214,G2945);
  not (G3215,G2720);
  not (G3218,G2948);
  not (G3219,G2744);
  not (G3222,G2797);
  not (G3225,G2752);
  not (G3228,G2752);
  not (G3231,G2759);
  not (G3234,G2759);
  not (G3237,G2780);
  not (G3240,G2984);
  not (G3241,G2810);
  not (G3244,G2817);
  not (G3247,G2837);
  not (G3250,G2810);
  not (G3253,G2817);
  not (G3256,G2865);
  not (G3259,G2857);
  not (G3262,G2865);
  not (G3265,G2999);
  not (G3266,G3002);
  not (G3267,G3005);
  not (G3268,G3008);
  not (G3269,G3026);
  not (G3270,G3029);
  not (G3271,G3032);
  not (G3272,G3035);
  nand (G3273,G2641,G3097);
  nand (G3274,G2638,G3098);
  nand (G3275,G2659,G3100);
  nand (G3276,G2656,G3101);
  nand (G3277,G3041,G3102);
  nand (G3280,G2363,G3103);
  not (G3281,G3060);
  nand (G3282,G1311,G3113);
  nand (G3283,G1314,G3115);
  nand (G3284,G1317,G3117);
  nand (G3285,G1320,G3119);
  nand (G3286,G1323,G3121);
  nand (G3287,G1326,G3123);
  nand (G3288,G1329,G3125);
  nand (G3289,G1332,G3127);
  nand (G3290,G1335,G3129);
  nand (G3291,G1341,G3133);
  nand (G3292,G1344,G3135);
  nand (G3293,G1347,G3137);
  nand (G3294,G1350,G3139);
  nand (G3295,G1353,G3141);
  nand (G3296,G1356,G3143);
  nand (G3297,G1359,G3145);
  nand (G3298,G1362,G3147);
  nand (G3299,G1365,G3149);
  nand (G3300,G1368,G3150);
  nand (G3301,G1371,G3152);
  nand (G3302,G1374,G3154);
  nand (G3303,G3156,G3057);
  nand (G3313,G1380,G3157);
  nand (G3314,G1383,G3159);
  nand (G3315,G1389,G3166);
  nand (G3316,G1392,G3168);
  nand (G3317,G3058,G3169);
  nand (G3331,G1398,G3171);
  nand (G3332,G1401,G3173);
  nand (G3333,G1404,G3175);
  nand (G3334,G2990,G3178);
  nand (G3335,G2987,G3179);
  nand (G3336,G2517,G3181);
  nand (G3337,G2621,G3182);
  nand (G3338,G3014,G3184);
  nand (G3339,G3011,G3185);
  nand (G3340,G3020,G3186);
  nand (G3341,G3017,G3187);
  nand (G3342,G2520,G3189);
  not (G3343,G3094);
  nand (G3344,G3195,G3196);
  nand (G3348,G3197,G3198);
  nand (G3351,G3202,G3203);
  nand (G3355,G3204,G3081);
  nor (G3358,G3205,G3084);
  nor (G3359,G3206,G3085);
  or (G3360,G2804,G3163);
  nand (G3363,G3002,G3265);
  nand (G3364,G2999,G3266);
  nand (G3365,G3008,G3267);
  nand (G3366,G3005,G3268);
  nand (G3367,G3029,G3269);
  nand (G3368,G3026,G3270);
  nand (G3369,G3035,G3271);
  nand (G3370,G3032,G3272);
  nand (G3371,G3191,G3190);
  not (G3374,G3060);
  nand (G3377,G3273,G3274);
  nand (G3380,G3275,G3276);
  nand (G3383,G3280,G3104);
  nand (G3386,G3282,G3114);
  nand (G3393,G3283,G3116);
  nand (G3404,G3284,G3118);
  nand (G3415,G3285,G3120);
  nand (G3421,G3286,G3122);
  nand (G3428,G3287,G3124);
  nand (G3438,G3288,G3126);
  nand (G3449,G3289,G3128);
  nand (G3459,G3290,G3130);
  not (G3466,G3211);
  nand (G3467,G3132,G3291);
  nand (G3474,G3134,G3292);
  nand (G3485,G3136,G3293);
  nand (G3495,G3138,G3294);
  nand (G3503,G3140,G3295);
  nand (G3517,G3142,G3296);
  nand (G3533,G3144,G3297);
  nand (G3546,G3146,G3298);
  nand (G3552,G3148,G3299);
  nand (G3559,G3300,G3151);
  nand (G3570,G3301,G3153);
  nand (G3576,G3302,G3155);
  nand (G3583,G3313,G3158);
  nand (G3594,G3314,G3160);
  nand (G3604,G3222,G1588);
  not (G3605,G3222);
  not (G3606,G3225);
  not (G3607,G3228);
  not (G3608,G3231);
  not (G3609,G3234);
  not (G3610,G3237);
  nand (G3611,G3165,G3315);
  nand (G3621,G3167,G3316);
  nand (G3629,G3170,G3331);
  nand (G3645,G3172,G3332);
  nand (G3658,G3174,G3333);
  not (G3664,G3244);
  not (G3665,G3253);
  nand (G3666,G3334,G3335);
  nand (G3670,G3180,G3336);
  nand (G3674,G3337,G3183);
  nand (G3677,G3338,G3339);
  nand (G3681,G3340,G3341);
  nand (G3685,G3188,G3342);
  and (G3688,G3208,G2872);
  not (G3689,G3215);
  not (G3690,G3219);
  not (G3691,G3241);
  not (G3692,G3247);
  not (G3693,G3250);
  not (G3694,G3256);
  not (G3695,G3259);
  not (G3696,G3262);
  nand (G3697,G3365,G3366);
  nand (G3700,G3363,G3364);
  nand (G3703,G3369,G3370);
  nand (G3706,G3367,G3368);
  not (G3709,G3277);
  nand (G3710,G3359,G3358);
  and (G3713,G3303,G2788);
  nand (G3714,G1386,G3605);
  not (G3715,G3360);
  and (G3716,G3317,G2844);
  and (G3717,G3317,G2844);
  not (G3718,G3371);
  nand (G3719,G3371,G3343);
  not (G3720,G3344);
  not (G3723,G3351);
  not (G3726,G3348);
  not (G3729,G3348);
  not (G3732,G3355);
  not (G3735,G3355);
  not (G3738,G3383);
  or (G3739,G3208,G3688);
  not (G3742,G3303);
  not (G3745,G3317);
  not (G3748,G3317);
  not (G3751,G3374);
  nand (G3752,G3374,G3099);
  not (G3753,G3377);
  not (G3754,G3380);
  nand (G3755,G3380,G3709);
  and (G3756,G3467,G2711);
  and (G3757,G3474,G3467,G2715);
  and (G3758,G3485,G3467,G2720,G3474);
  and (G3759,G3559,G2752,G2780,G2759);
  and (G3760,G3386,G2675);
  and (G3761,G3393,G3386,G2679);
  and (G3762,G3404,G3386,G2685,G3393);
  and (G3763,G3611,G2810,G2837,G2817);
  not (G3764,G3415);
  and (G3765,G3393,G3415,G3404,G3386);
  and (G3768,G3393,G2679);
  and (G3769,G3404,G2685,G3393);
  and (G3770,G3415,G3404,G3393);
  and (G3771,G3393,G2679);
  and (G3772,G2685,G3404,G3393);
  and (G3773,G3404,G2685);
  and (G3774,G3415,G3404);
  and (G3775,G3404,G2685);
  and (G3776,G3428,G3459,G3438,G3421,G3449);
  and (G3779,G3421,G2693);
  and (G3780,G3428,G3421,G2696);
  and (G3781,G3438,G3421,G2700,G3428);
  and (G3782,G3449,G3438,G3421,G2705,G3428);
  and (G3783,G3428,G2696);
  and (G3784,G3438,G2700,G3428);
  and (G3785,G3449,G3438,G2705,G3428);
  and (G3786,G2,G3459,G3438,G3449,G3428);
  and (G3787,G2700,G3438);
  and (G3788,G3449,G3438,G2705);
  and (G3789,G2,G3459,G3438,G3449);
  and (G3790,G3449,G2705);
  and (G3791,G2,G3459,G3449);
  and (G3792,G2,G3459);
  and (G3793,G3546,G3485,G3474,G3467);
  and (G3796,G3474,G2715);
  and (G3797,G3485,G2720,G3474);
  and (G3798,G3546,G3485,G3474);
  and (G3799,G3474,G2715);
  and (G3800,G3485,G2720,G3474);
  and (G3801,G3485,G2720);
  and (G3802,G3552,G3533,G3517,G3503,G3495);
  and (G3805,G3495,G2727);
  and (G3806,G3503,G3495,G2731);
  and (G3807,G3517,G3495,G2737,G3503);
  and (G3808,G3533,G3517,G3495,G2744,G3503);
  and (G3809,G3503,G2731);
  and (G3810,G3517,G2737,G3503);
  and (G3811,G3533,G3517,G2744,G3503);
  and (G3812,G3552,G3517,G3503,G3533);
  and (G3813,G3503,G2731);
  and (G3814,G3517,G2737,G3503);
  and (G3815,G3533,G3517,G2744,G3503);
  and (G3816,G3517,G2737);
  and (G3817,G3533,G3517,G2744);
  and (G3818,G3552,G3517,G3533);
  and (G3819,G3517,G2737);
  and (G3820,G3533,G3517,G2744);
  and (G3821,G3533,G2744);
  and (G3822,G3546,G3485);
  and (G3823,G3552,G3533);
  not (G3824,G3570);
  and (G3825,G2759,G3570,G3559,G2752);
  and (G3828,G3559,G2780,G2759);
  and (G3829,G3570,G3559,G2759);
  and (G3830,G2780,G3559,G2759);
  and (G3831,G3559,G2780);
  and (G3832,G3570,G3559);
  and (G3833,G3559,G2780);
  and (G3834,G3303,G2797,G3583,G3576,G3594);
  and (G3837,G3576,G2540);
  and (G3838,G3303,G3576,G2788);
  and (G3839,G3583,G3576,G2792,G3303);
  and (G3840,G3594,G3583,G3576,G2804,G3303);
  and (G3841,G3583,G2792,G3303);
  and (G3842,G3594,G3583,G2804,G3303);
  and (G3843,G21,G2797,G3583,G3594,G3303);
  and (G3844,G2792,G3583);
  and (G3845,G3594,G3583,G2804);
  and (G3846,G21,G2797,G3583,G3594);
  and (G3847,G3594,G2804);
  and (G3848,G21,G2797,G3594);
  nand (G3849,G3604,G3714);
  and (G3852,G3658,G3611,G2817,G2810);
  and (G3855,G3611,G2837,G2817);
  and (G3856,G3658,G3611,G2817);
  and (G3857,G3611,G2837,G2817);
  and (G3858,G3611,G2837);
  and (G3859,G2865,G3645,G3629,G3317,G3621);
  and (G3862,G3621,G2543);
  and (G3863,G3317,G3621,G2844);
  and (G3864,G3629,G3621,G2850,G3317);
  and (G3865,G3645,G3629,G3621,G2857,G3317);
  and (G3866,G3629,G2850,G3317);
  and (G3867,G3645,G3629,G2857,G3317);
  and (G3868,G2865,G3629,G3317,G3645);
  and (G3869,G3629,G2850,G3317);
  and (G3870,G3645,G3629,G2857,G3317);
  and (G3871,G3629,G2850);
  and (G3872,G3645,G3629,G2857);
  and (G3873,G2865,G3629,G3645);
  and (G3874,G3629,G2850);
  and (G3875,G3645,G3629,G2857);
  and (G3876,G3645,G2857);
  and (G3877,G3658,G3611);
  and (G3878,G2865,G3645);
  not (G3879,G3666);
  not (G3882,G3670);
  not (G3885,G3677);
  not (G3888,G3681);
  not (G3891,G3674);
  not (G3894,G3674);
  not (G3897,G3685);
  not (G3900,G3685);
  nand (G3903,G3094,G3718);
  not (G3904,G3710);
  nand (G3905,G3710,G3738);
  not (G3906,G3459);
  not (G3909,G3386);
  not (G3912,G3386);
  not (G3915,G3393);
  not (G3918,G3393);
  not (G3921,G3404);
  not (G3924,G3404);
  not (G3927,G3421);
  not (G3930,G3428);
  not (G3933,G3438);
  not (G3936,G3449);
  not (G3939,G3546);
  not (G3942,G3485);
  not (G3945,G3467);
  not (G3948,G3474);
  not (G3951,G3546);
  not (G3954,G3485);
  not (G3957,G3467);
  not (G3960,G3474);
  not (G3963,G3552);
  not (G3966,G3533);
  not (G3969,G3495);
  not (G3972,G3517);
  not (G3975,G3503);
  not (G3978,G3503);
  not (G3981,G3552);
  not (G3984,G3533);
  not (G3987,G3495);
  not (G3990,G3517);
  not (G3993,G3559);
  not (G3996,G3559);
  not (G3999,G3576);
  not (G4002,G3583);
  not (G4005,G3594);
  not (G4008,G3658);
  not (G4011,G3611);
  not (G4014,G3658);
  not (G4017,G3611);
  not (G4020,G3645);
  not (G4023,G3621);
  not (G4026,G3629);
  not (G4029,G3645);
  not (G4032,G3621);
  not (G4035,G3629);
  not (G4038,G3697);
  not (G4039,G3700);
  not (G4040,G3703);
  not (G4041,G3706);
  nand (G4042,G2644,G3751);
  nand (G4043,G3277,G3754);
  or (G4044,G2667,G3756,G3757,G3758);
  or (G4045,G2492,G3109,G3110,G3759);
  or (G4046,G2670,G3760,G3761,G3762);
  or (G4047,G2492,G3111,G3112,G3763);
  or (G4048,G2692,G3779,G3780,G3781,G3782);
  or (G4051,G2715,G3801);
  or (G4054,G2726,G3805,G3806,G3807,G3808);
  or (G4058,G2737,G3821);
  or (G4061,G2787,G3837,G3838,G3839,G3840);
  not (G4064,G3742);
  or (G4065,G2832,G3858);
  or (G4068,G2843,G3862,G3863,G3864,G3865);
  or (G4072,G2850,G3876);
  not (G4075,G3745);
  not (G4076,G3748);
  nand (G4077,G3903,G3719);
  not (G4080,G3726);
  not (G4081,G3729);
  not (G4082,G3732);
  not (G4083,G3735);
  and (G4084,G3344,G2879,G3726);
  and (G4085,G3720,G3192,G3729);
  and (G4086,G3351,G2883,G3732);
  and (G4087,G3723,G3199,G3735);
  nand (G4088,G3383,G3904);
  nand (G4089,G3739,G61);
  or (G4092,G2675,G3768,G3769,G3770);
  nor (G4095,G2675,G3771,G3772);
  or (G4098,G2679,G3773,G3774);
  nor (G4101,G2679,G3775);
  or (G4104,G2693,G3783,G3784,G3785,G3786);
  or (G4107,G2696,G3787,G3788,G3789);
  or (G4110,G2700,G3790,G3791);
  or (G4113,G2705,G3792);
  or (G4116,G2711,G3796,G3797,G3798);
  nor (G4119,G2711,G3799,G3800);
  or (G4122,G2731,G3816,G3817,G3818);
  or (G4125,G2727,G3809,G3810,G3811,G3812);
  nor (G4128,G2731,G3819,G3820);
  nor (G4131,G2727,G3813,G3814,G3815);
  or (G4134,G2770,G3161,G3828,G3829);
  nor (G4137,G2770,G3162,G3830);
  or (G4140,G2774,G3831,G3832);
  nor (G4143,G2774,G3833);
  or (G4146,G2540,G3713,G3841,G3842,G3843);
  or (G4149,G2788,G3844,G3845,G3846);
  or (G4152,G2792,G3847,G3848);
  or (G4155,G2828,G3176,G3855,G3856);
  nor (G4158,G2828,G3177,G3857);
  or (G4161,G2844,G3871,G3872,G3873);
  or (G4164,G2543,G3716,G3866,G3867,G3868);
  nor (G4167,G2844,G3874,G3875);
  nor (G4170,G2543,G3717,G3869,G3870);
  nand (G4173,G3700,G4038);
  nand (G4174,G3697,G4039);
  nand (G4175,G3706,G4040);
  nand (G4176,G3703,G4041);
  nand (G4177,G4042,G3752);
  nand (G4180,G3755,G4043);
  not (G4183,G3849);
  nand (G4184,G3906,G1510);
  not (G4185,G3906);
  not (G4186,G3909);
  not (G4187,G3912);
  not (G4188,G3915);
  not (G4189,G3918);
  nand (G4190,G3921,G3131);
  not (G4191,G3921);
  nand (G4192,G3924,G3466);
  not (G4193,G3924);
  and (G4194,G3776,G2);
  not (G4195,G3927);
  not (G4196,G3930);
  not (G4197,G3933);
  not (G4198,G3936);
  not (G4199,G3802);
  not (G4200,G3948);
  not (G4201,G3960);
  not (G4202,G3975);
  not (G4203,G3978);
  nand (G4204,G3993,G3164);
  not (G4205,G3993);
  nand (G4206,G3996,G3610);
  not (G4207,G3996);
  and (G4208,G3834,G21);
  not (G4209,G3999);
  not (G4210,G4002);
  nand (G4211,G4005,G3715);
  not (G4212,G4005);
  not (G4213,G3859);
  not (G4214,G3891);
  not (G4215,G3894);
  not (G4216,G3897);
  not (G4217,G3900);
  and (G4218,G3670,G3666,G3891);
  and (G4219,G3882,G3879,G3894);
  and (G4220,G3681,G3677,G3897);
  and (G4221,G3888,G3885,G3900);
  and (G4222,G3849,G1264,G2003);
  and (G4223,G3192,G3344,G4080);
  and (G4224,G2879,G3720,G4081);
  and (G4225,G3199,G3351,G4082);
  and (G4226,G2883,G3723,G4083);
  nand (G4227,G4088,G3905);
  not (G4230,G3939);
  not (G4231,G3942);
  not (G4232,G3945);
  not (G4233,G3951);
  not (G4234,G3954);
  not (G4235,G3957);
  not (G4236,G3963);
  not (G4237,G3966);
  not (G4238,G3969);
  not (G4239,G3972);
  not (G4240,G3990);
  not (G4241,G3981);
  not (G4242,G3984);
  not (G4243,G3987);
  not (G4244,G4008);
  not (G4245,G4011);
  not (G4246,G4014);
  not (G4247,G4017);
  not (G4248,G4020);
  not (G4249,G4023);
  not (G4250,G4026);
  not (G4251,G4035);
  not (G4252,G4029);
  not (G4253,G4032);
  nand (G4254,G4173,G4174);
  nand (G4257,G4175,G4176);
  and (G4260,G3793,G4054);
  and (G4261,G4061,G3825);
  and (G4262,G4048,G3765);
  and (G4263,G3852,G4068);
  not (G4264,G4077);
  nand (G4265,G1338,G4185);
  not (G4266,G4092);
  nand (G4267,G4092,G4186);
  not (G4268,G4095);
  nand (G4269,G4095,G4187);
  not (G4270,G4098);
  nand (G4271,G4098,G4188);
  not (G4272,G4101);
  nand (G4273,G4101,G4189);
  nand (G4274,G2915,G4191);
  nand (G4275,G3211,G4193);
  or (G4276,G4048,G4194);
  not (G4282,G4104);
  nand (G4283,G4104,G4195);
  not (G4284,G4107);
  nand (G4285,G4107,G4196);
  not (G4286,G4110);
  nand (G4287,G4110,G4197);
  not (G4288,G4113);
  nand (G4289,G4113,G4198);
  not (G4290,G4054);
  not (G4293,G4134);
  nand (G4294,G4134,G3606);
  not (G4295,G4137);
  nand (G4296,G4137,G3607);
  not (G4297,G4140);
  nand (G4298,G4140,G3608);
  not (G4299,G4143);
  nand (G4300,G4143,G3609);
  nand (G4301,G2966,G4205);
  nand (G4302,G3237,G4207);
  or (G4303,G4061,G4208);
  not (G4309,G4146);
  nand (G4310,G4146,G4209);
  not (G4311,G4149);
  nand (G4312,G4149,G4064);
  not (G4313,G4152);
  nand (G4314,G4152,G4210);
  nand (G4315,G3360,G4212);
  not (G4316,G4068);
  and (G4319,G3879,G3670,G4214);
  and (G4320,G3666,G3882,G4215);
  and (G4321,G3885,G3681,G4216);
  and (G4322,G3677,G3888,G4217);
  or (G4323,G2600,G4222,G2324);
  nor (G4329,G4223,G4084);
  nor (G4330,G4224,G4085);
  nor (G4331,G4225,G4086);
  nor (G4332,G4226,G4087);
  not (G4333,G4180);
  and (G4334,G3739,G4089);
  and (G4335,G4089,G61);
  or (G4336,G4051,G3822);
  not (G4339,G4116);
  not (G4340,G4051);
  not (G4343,G4119);
  not (G4344,G4122);
  nand (G4345,G4122,G3218);
  or (G4346,G4058,G3823);
  not (G4349,G4125);
  not (G4350,G4128);
  nand (G4351,G4128,G3690);
  not (G4352,G4058);
  not (G4355,G4131);
  or (G4356,G4065,G3877);
  not (G4359,G4155);
  not (G4360,G4065);
  not (G4363,G4158);
  or (G4364,G4072,G3878);
  not (G4367,G4161);
  not (G4368,G4164);
  not (G4369,G4167);
  nand (G4370,G4167,G3695);
  not (G4371,G4072);
  not (G4374,G4170);
  not (G4375,G4177);
  nand (G4376,G4177,G3753);
  not (G4377,G4227);
  nand (G4378,G4184,G4265);
  nand (G4381,G3909,G4266);
  nand (G4382,G3912,G4268);
  nand (G4383,G3915,G4270);
  nand (G4384,G3918,G4272);
  nand (G4385,G4190,G4274);
  nand (G4386,G4192,G4275);
  nand (G4387,G3927,G4282);
  nand (G4388,G3930,G4284);
  nand (G4389,G3933,G4286);
  nand (G4390,G3936,G4288);
  nand (G4391,G3225,G4293);
  nand (G4392,G3228,G4295);
  nand (G4393,G3231,G4297);
  nand (G4394,G3234,G4299);
  nand (G4395,G4204,G4301);
  nand (G4396,G4206,G4302);
  nand (G4397,G3999,G4309);
  nand (G4398,G3742,G4311);
  nand (G4399,G4002,G4313);
  nand (G4400,G4211,G4315);
  nor (G4403,G4319,G4218);
  nor (G4404,G4320,G4219);
  nor (G4405,G4321,G4220);
  nor (G4406,G4322,G4221);
  not (G4407,G4254);
  not (G4408,G4257);
  or (G4409,G4334,G4335);
  nand (G4413,G2948,G4344);
  nand (G4414,G3219,G4350);
  nand (G4415,G3259,G4369);
  nand (G4416,G3377,G4375);
  nand (G4417,G4330,G4329);
  nand (G4420,G4332,G4331);
  and (G4423,G4323,G1554,G1565);
  and (G4424,G4323,G1629,G1640);
  and (G4425,G4323,G1652,G1663);
  and (G4426,G4323,G1674,G1685);
  nand (G4427,G4381,G4267);
  nand (G4428,G4382,G4269);
  nand (G4429,G4383,G4271);
  nand (G4430,G4384,G4273);
  not (G4431,G4385);
  not (G4432,G4276);
  nand (G4437,G4387,G4283);
  nand (G4440,G4388,G4285);
  nand (G4443,G4389,G4287);
  nand (G4446,G4390,G4289);
  and (G4449,G4276,G3764);
  and (G4450,G4290,G4199);
  nand (G4453,G4391,G4294);
  nand (G4454,G4392,G4296);
  nand (G4455,G4393,G4298);
  nand (G4456,G4394,G4300);
  not (G4457,G4395);
  not (G4458,G4303);
  nand (G4463,G4397,G4310);
  nand (G4466,G4398,G4312);
  nand (G4469,G4399,G4314);
  and (G4472,G4303,G3824);
  and (G4473,G4316,G4213);
  not (G4476,G4336);
  nand (G4477,G4336,G3214);
  not (G4478,G4340);
  nand (G4479,G4340,G3689);
  nand (G4480,G4345,G4413);
  not (G4483,G4346);
  nand (G4484,G4351,G4414);
  not (G4487,G4352);
  not (G4488,G4356);
  nand (G4489,G4356,G3240);
  not (G4490,G4360);
  nand (G4491,G4360,G3692);
  not (G4492,G4364);
  nand (G4493,G4364,G4367);
  nand (G4494,G4370,G4415);
  not (G4497,G4371);
  nand (G4498,G4404,G4403);
  nand (G4501,G4406,G4405);
  nand (G4504,G4416,G4376);
  not (G4507,G4378);
  not (G4508,G4400);
  and (G4509,G4409,G171,G1242);
  not (G4510,G4428);
  not (G4511,G4430);
  and (G4512,G4276,G4427);
  and (G4513,G4276,G4429);
  and (G4514,G4276,G4431);
  not (G4515,G4454);
  not (G4516,G4456);
  and (G4517,G4303,G4453);
  and (G4518,G4303,G4455);
  and (G4519,G4303,G4457);
  and (G4520,G4378,G1248,G1981);
  and (G4521,G4400,G1264,G2003);
  not (G4522,G4417);
  not (G4523,G4420);
  nand (G4524,G4420,G4333);
  nand (G4525,G2945,G4476);
  nand (G4526,G3215,G4478);
  nand (G4527,G2984,G4488);
  nand (G4528,G3247,G4490);
  nand (G4529,G4161,G4492);
  not (G4530,G4446);
  not (G4531,G4443);
  not (G4532,G4440);
  not (G4533,G4437);
  not (G4534,G4469);
  not (G4535,G4466);
  not (G4536,G4463);
  and (G4537,G4510,G4432);
  and (G4538,G4511,G4432);
  and (G4539,G4386,G4432);
  and (G4540,G3415,G4432);
  not (G4541,G4450);
  and (G4542,G4515,G4458);
  and (G4543,G4516,G4458);
  and (G4544,G4396,G4458);
  and (G4545,G3570,G4458);
  not (G4546,G4473);
  not (G4547,G4498);
  nand (G4548,G4498,G4407);
  not (G4549,G4501);
  nand (G4550,G4501,G4408);
  and (G4551,G4446,G1248,G1981);
  and (G4552,G4443,G1248,G1981);
  and (G4553,G4440,G1248,G1981);
  or (G4554,G3068,G4520,G2320);
  and (G4560,G4469,G1264,G2003);
  and (G4561,G4466,G1264,G2003);
  or (G4562,G3072,G4521,G2325);
  nand (G4568,G4504,G4522);
  not (G4569,G4504);
  nand (G4570,G4180,G4523);
  and (G4571,G4437,G1280,G2031);
  and (G4572,G4463,G1294,G2053);
  nand (G4573,G4477,G4525);
  nand (G4576,G4479,G4526);
  not (G4579,G4480);
  nand (G4580,G4480,G4483);
  not (G4581,G4484);
  nand (G4582,G4484,G4487);
  nand (G4583,G4489,G4527);
  nand (G4586,G4491,G4528);
  nand (G4589,G4493,G4529);
  not (G4592,G4494);
  nand (G4593,G4494,G4497);
  or (G4594,G4537,G4512);
  or (G4597,G4538,G4513);
  or (G4600,G4539,G4514);
  or (G4603,G4540,G4449);
  or (G4606,G4542,G4517);
  or (G4613,G4543,G4518);
  or (G4616,G4544,G4519);
  or (G4619,G4545,G4472);
  nand (G4622,G4254,G4547);
  nand (G4623,G4257,G4549);
  or (G4624,G3069,G4551,G2321);
  or (G4630,G3070,G4552,G2322);
  or (G4636,G3071,G4553,G2323);
  or (G4642,G3073,G4560,G2326);
  or (G4648,G2516,G4561,G2327);
  nand (G4654,G4417,G4569);
  nand (G4655,G4570,G4524);
  or (G4658,G3086,G4571,G2339);
  or (G4664,G3090,G4572,G2344);
  nand (G4670,G4346,G4579);
  nand (G4671,G4352,G4581);
  nand (G4672,G4371,G4592);
  and (G4673,G4554,G718,G1565);
  and (G4674,G4562,G1554,G1565);
  and (G4675,G4554,G780,G1640);
  and (G4676,G4562,G1629,G1640);
  and (G4677,G4554,G860,G1663);
  and (G4678,G4562,G1652,G1663);
  and (G4679,G4562,G1674,G1685);
  and (G4680,G4554,G884,G1685);
  nand (G4681,G4622,G4548);
  nand (G4684,G4623,G4550);
  nand (G4687,G4568,G4654);
  not (G4690,G4573);
  nand (G4691,G4573,G4339);
  not (G4692,G4576);
  nand (G4693,G4576,G4343);
  nand (G4694,G4670,G4580);
  nand (G4697,G4671,G4582);
  not (G4700,G4583);
  nand (G4701,G4583,G4359);
  not (G4702,G4586);
  nand (G4703,G4586,G4363);
  not (G4704,G4589);
  nand (G4705,G4589,G4368);
  nand (G4706,G4672,G4593);
  not (G4709,G4603);
  not (G4710,G4600);
  not (G4711,G4597);
  not (G4712,G4594);
  not (G4713,G4619);
  not (G4714,G4616);
  not (G4715,G4613);
  not (G4716,G4606);
  and (G4717,G4664,G1526,G1537);
  and (G4718,G4658,G694,G1537);
  or (G4719,G4423,G4673,G2162,G1465);
  and (G4720,G4624,G718,G1565);
  and (G4721,G4642,G1554,G1565);
  and (G4722,G4630,G718,G1565);
  and (G4723,G4648,G1554,G1565);
  and (G4724,G4636,G718,G1565);
  and (G4725,G4664,G1601,G1612);
  and (G4726,G4658,G756,G1612);
  or (G4727,G4424,G4675,G2173,G1474);
  and (G4728,G4624,G780,G1640);
  and (G4729,G4642,G1629,G1640);
  and (G4730,G4630,G780,G1640);
  and (G4731,G4648,G1629,G1640);
  and (G4732,G4636,G780,G1640);
  and (G4733,G4664,G1914,G1925);
  and (G4734,G4658,G1184,G1925);
  and (G4735,G4648,G1652,G1663);
  and (G4736,G4636,G860,G1663);
  and (G4737,G4642,G1652,G1663);
  and (G4738,G4630,G860,G1663);
  and (G4739,G4624,G860,G1663);
  and (G4740,G4664,G1948,G1959);
  and (G4741,G4658,G1218,G1959);
  and (G4742,G4648,G1674,G1685);
  and (G4743,G4636,G884,G1685);
  and (G4744,G4642,G1674,G1685);
  and (G4745,G4630,G884,G1685);
  and (G4746,G4624,G884,G1685);
  and (G4747,G4606,G171,G170);
  not (G4748,G4655);
  and (G4749,G4655,G1941);
  and (G4750,G4603,G1280,G2031);
  and (G4751,G4600,G1280,G2031);
  and (G4752,G4597,G1280,G2031);
  and (G4753,G4594,G1280,G2031);
  and (G4754,G4619,G1294,G2053);
  and (G4755,G4616,G1294,G2053);
  and (G4756,G4613,G1294,G2053);
  and (G4757,G4606,G1294,G2053);
  nand (G4758,G4409,G4606);
  nand (G4761,G4116,G4690);
  nand (G4762,G4119,G4692);
  nand (G4763,G4155,G4700);
  nand (G4764,G4158,G4702);
  nand (G4765,G4164,G4704);
  or (G4766,G4717,G4718,G2157,G1460);
  or (G4767,G4674,G4720,G2163,G1466);
  or (G4768,G4721,G4722,G2164,G1467);
  or (G4769,G4723,G4724,G2165,G1468);
  or (G4770,G4725,G4726,G2168,G1469);
  or (G4771,G4676,G4728,G2174,G1475);
  or (G4772,G4729,G4730,G2175,G1476);
  or (G4773,G4731,G4732,G2176,G1477);
  or (G4774,G3055,G4509,G1497,G4747);
  and (G4775,G4748,G1992,G2003);
  not (G4776,G4681);
  not (G4777,G4684);
  not (G4778,G4687);
  and (G4779,G4687,G1941);
  or (G4780,G3087,G4750,G2340);
  or (G4786,G3088,G4751,G2341);
  or (G4792,G3089,G4752,G2342);
  or (G4798,G3207,G4753,G2343);
  or (G4804,G3091,G4754,G2345);
  or (G4810,G3092,G4755,G2346);
  or (G4816,G2887,G4756,G2347);
  or (G4822,G3093,G4757,G2348);
  nand (G4828,G4761,G4691);
  nand (G4831,G4762,G4693);
  not (G4834,G4694);
  nand (G4835,G4694,G4349);
  not (G4836,G4697);
  nand (G4837,G4697,G4355);
  nand (G4838,G4763,G4701);
  nand (G4841,G4764,G4703);
  nand (G4844,G4765,G4705);
  not (G4847,G4706);
  nand (G4848,G4706,G4374);
  and (G4849,G4409,G4758);
  and (G4850,G4758,G4606);
  and (G4851,G156,G4776,G4777,G4264,G4377);
  and (G4852,G4778,G1970,G1981);
  nand (G4853,G4125,G4834);
  nand (G4854,G4131,G4836);
  nand (G4855,G4170,G4847);
  and (G4856,G4804,G1526,G1537);
  and (G4857,G4780,G694,G1537);
  and (G4858,G4810,G1526,G1537);
  and (G4859,G4786,G694,G1537);
  and (G4860,G4816,G1526,G1537);
  and (G4861,G4792,G694,G1537);
  and (G4862,G4822,G1526,G1537);
  and (G4863,G4798,G694,G1537);
  and (G4864,G4804,G1601,G1612);
  and (G4865,G4780,G756,G1612);
  and (G4866,G4810,G1601,G1612);
  and (G4867,G4786,G756,G1612);
  and (G4868,G4816,G1601,G1612);
  and (G4869,G4792,G756,G1612);
  and (G4870,G4822,G1601,G1612);
  and (G4871,G4798,G756,G1612);
  and (G4872,G4822,G1948,G1959);
  and (G4873,G4798,G1218,G1959);
  and (G4874,G4822,G1914,G1925);
  and (G4875,G4798,G1184,G1925);
  and (G4876,G4816,G1914,G1925);
  and (G4877,G4792,G1184,G1925);
  and (G4878,G4810,G1914,G1925);
  and (G4879,G4786,G1184,G1925);
  and (G4880,G4804,G1914,G1925);
  and (G4881,G4780,G1184,G1925);
  and (G4882,G4816,G1948,G1959);
  and (G4883,G4792,G1218,G1959);
  and (G4884,G4810,G1948,G1959);
  and (G4885,G4786,G1218,G1959);
  and (G4886,G4804,G1948,G1959);
  and (G4887,G4780,G1218,G1959);
  not (G4888,G4828);
  nand (G4889,G4828,G4230);
  not (G4890,G4831);
  nand (G4891,G4831,G4233);
  nand (G4892,G4853,G4835);
  nand (G4895,G4854,G4837);
  not (G4898,G4838);
  nand (G4899,G4838,G4244);
  not (G4900,G4841);
  nand (G4901,G4841,G4246);
  not (G4902,G4844);
  nand (G4903,G4844,G3694);
  nand (G4904,G4855,G4848);
  or (G4907,G4856,G4857,G2158,G1461);
  or (G4908,G4858,G4859,G2159,G1462);
  or (G4909,G4860,G4861,G2160,G1463);
  or (G4910,G4862,G4863,G2161,G1464);
  or (G4911,G4864,G4865,G2169,G1470);
  or (G4912,G4866,G4867,G2170,G1471);
  or (G4913,G4868,G4869,G2171,G1472);
  or (G4914,G4870,G4871,G2172,G1473);
  nand (G4915,G3939,G4888);
  nand (G4916,G3951,G4890);
  nand (G4917,G4008,G4898);
  nand (G4918,G4014,G4900);
  nand (G4919,G3256,G4902);
  nand (G4920,G4915,G4889);
  nand (G4923,G4916,G4891);
  not (G4926,G4892);
  nand (G4927,G4892,G4236);
  not (G4928,G4895);
  nand (G4929,G4895,G4241);
  nand (G4930,G4917,G4899);
  nand (G4933,G4918,G4901);
  nand (G4936,G4919,G4903);
  not (G4939,G4904);
  nand (G4940,G4904,G3696);
  nand (G4941,G3963,G4926);
  nand (G4942,G3981,G4928);
  nand (G4943,G3262,G4939);
  not (G4944,G4920);
  nand (G4945,G4920,G4231);
  not (G4946,G4923);
  nand (G4947,G4923,G4234);
  nand (G4948,G4941,G4927);
  nand (G4951,G4942,G4929);
  not (G4954,G4930);
  nand (G4955,G4930,G4245);
  not (G4956,G4933);
  nand (G4957,G4933,G4247);
  not (G4958,G4936);
  nand (G4959,G4936,G4248);
  nand (G4960,G4943,G4940);
  nand (G4963,G3942,G4944);
  nand (G4964,G3954,G4946);
  nand (G4965,G4011,G4954);
  nand (G4966,G4017,G4956);
  nand (G4967,G4020,G4958);
  nand (G4968,G4963,G4945);
  nand (G4971,G4964,G4947);
  not (G4974,G4948);
  nand (G4975,G4948,G4237);
  not (G4976,G4951);
  nand (G4977,G4951,G4242);
  nand (G4978,G4965,G4955);
  nand (G4981,G4966,G4957);
  nand (G4984,G4967,G4959);
  not (G4987,G4960);
  nand (G4988,G4960,G4252);
  nand (G4989,G3966,G4974);
  nand (G4990,G3984,G4976);
  nand (G4991,G4029,G4987);
  not (G4992,G4968);
  nand (G4993,G4968,G4232);
  not (G4994,G4971);
  nand (G4995,G4971,G4235);
  nand (G4996,G4989,G4975);
  nand (G4999,G4990,G4977);
  not (G5002,G4978);
  nand (G5003,G4978,G3691);
  not (G5004,G4981);
  nand (G5005,G4981,G3693);
  not (G5006,G4984);
  nand (G5007,G4984,G4249);
  nand (G5008,G4991,G4988);
  nand (G5011,G3945,G4992);
  nand (G5012,G3957,G4994);
  nand (G5013,G3241,G5002);
  nand (G5014,G3250,G5004);
  nand (G5015,G4023,G5006);
  nand (G5016,G5011,G4993);
  nand (G5019,G5012,G4995);
  not (G5022,G4996);
  nand (G5023,G4996,G4238);
  not (G5024,G4999);
  nand (G5025,G4999,G4243);
  nand (G5026,G5013,G5003);
  nand (G5029,G5014,G5005);
  nand (G5032,G5015,G5007);
  not (G5035,G5008);
  nand (G5036,G5008,G4253);
  nand (G5037,G3969,G5022);
  nand (G5038,G3987,G5024);
  nand (G5039,G4032,G5035);
  not (G5040,G5016);
  nand (G5041,G5016,G4200);
  not (G5042,G5019);
  nand (G5043,G5019,G4201);
  not (G5044,G5026);
  nand (G5045,G5026,G3664);
  not (G5046,G5029);
  nand (G5047,G5029,G3665);
  nand (G5048,G5037,G5023);
  nand (G5051,G5038,G5025);
  not (G5054,G5032);
  nand (G5055,G5032,G4250);
  nand (G5056,G5039,G5036);
  nand (G5059,G3948,G5040);
  nand (G5060,G3960,G5042);
  nand (G5061,G3244,G5044);
  nand (G5062,G3253,G5046);
  nand (G5063,G4026,G5054);
  nand (G5064,G5059,G5041);
  nand (G5067,G5060,G5043);
  nand (G5070,G5061,G5045);
  nand (G5073,G5062,G5047);
  not (G5076,G5048);
  nand (G5077,G5048,G4239);
  not (G5078,G5051);
  nand (G5079,G5051,G4240);
  nand (G5080,G5063,G5055);
  not (G5083,G5056);
  nand (G5084,G5056,G4251);
  nand (G5085,G3972,G5076);
  nand (G5086,G3990,G5078);
  nand (G5087,G4035,G5083);
  and (G5088,G5067,G4290,G690);
  and (G5089,G5064,G4054,G690);
  and (G5090,G5067,G4450,G157);
  and (G5091,G5064,G4541,G157);
  not (G5092,G5080);
  nand (G5093,G5080,G4075);
  and (G5094,G5073,G4316,G752);
  and (G5095,G5070,G4068,G752);
  and (G5096,G5073,G4473,G162);
  and (G5097,G5070,G4546,G162);
  nand (G5098,G5085,G5077);
  nand (G5101,G5086,G5079);
  nand (G5104,G5087,G5084);
  nand (G5107,G3745,G5092);
  or (G5108,G5088,G5089,G5090,G5091);
  or (G5111,G5094,G5095,G5096,G5097);
  not (G5114,G5098);
  nand (G5115,G5098,G4202);
  not (G5116,G5101);
  nand (G5117,G5101,G4203);
  nand (G5118,G5107,G5093);
  not (G5119,G5104);
  nand (G5120,G5104,G4076);
  nand (G5121,G3975,G5114);
  nand (G5122,G3978,G5116);
  not (G5123,G5108);
  nand (G5124,G3748,G5119);
  and (G5125,G162,G5118);
  not (G5126,G5111);
  nand (G5127,G5121,G5115);
  nand (G5128,G5122,G5117);
  nand (G5129,G5124,G5120);
  not (G5130,G5128);
  and (G5131,G157,G5127);
  not (G5132,G5129);
  and (G5133,G5130,G690);
  and (G5134,G5132,G752);
  or (G5135,G5133,G5131);
  or (G5138,G5134,G5125);
  nand (G5141,G5135,G5123);
  not (G5142,G5135);
  nand (G5143,G5138,G5126);
  not (G5144,G5138);
  nand (G5145,G5108,G5142);
  nand (G5146,G5111,G5144);
  nand (G5147,G5141,G5145);
  nand (G5150,G5143,G5146);
  and (G5153,G5150,G1264,G2003);
  and (G5154,G5147,G1248,G1981);
  not (G5155,G5147);
  not (G5156,G5150);
  and (G5157,G5155,G1214);
  and (G5158,G5156,G1214);
  or (G5159,G4779,G5157);
  or (G5162,G4749,G5158);
  and (G5165,G5159,G1936);
  and (G5166,G5162,G1936);
  and (G5167,G5159,G1936);
  and (G5168,G5162,G1936);
  or (G5169,G5165,G1944);
  or (G5172,G5166,G1945);
  or (G5175,G5167,G1946);
  or (G5178,G5168,G1947);
  and (G5181,G5178,G1652,G1663);
  and (G5182,G5175,G860,G1663);
  and (G5183,G5178,G1674,G1685);
  and (G5184,G5175,G884,G1685);
  and (G5185,G5172,G1554,G1565);
  and (G5186,G5169,G718,G1565);
  and (G5187,G5172,G1629,G1640);
  and (G5188,G5169,G780,G1640);
  or (G5189,G5185,G5186,G2203,G1576);
  or (G5190,G5187,G5188,G2204,G1651);
  and (G5191,G5189,G1548);
  and (G5192,G5190,G1623);
  not (G5193,G66);
  not (G5194,G113);
  not (G5195,G165);
  not (G5196,G151);
  not (G5197,G127);
  not (G5198,G131);
  and (G5199,G153,G156);
  not (G5200,G152);
  not (G5201,G151);
  not (G5202,G151);
  not (G5203,G125);
  not (G5204,G129);
  and (G5205,G66,G67);
  not (G5206,G99);
  not (G5207,G153);
  not (G5208,G156);
  not (G5209,G155);
  not (G5210,G684);
  and (G5211,G63,G685);
  not (G5212,G687);
  not (G5213,G688);
  not (G5214,G742);
  not (G5215,G749);
  not (G5216,G980);
  not (G5217,G1067);
  not (G5218,G1308);
  not (G5219,G1067);
  nand (G5220,G976,G65);
  not (G5221,G976);
  not (G5222,G1577);
  not (G5223,G1577);
  not (G5224,G1577);
  not (G5225,G1577);
  not (G5226,G2064);
  not (G5227,G2064);
  not (G5228,G2528);
  not (G5229,G2533);
  not (G5230,G2538);
  not (G5231,G2539);
  and (G5232,G2671,G1750);
  and (G5233,G2672,G1750);
  and (G5234,G2673,G1750);
  and (G5235,G2674,G1750);
  and (G5236,G3105,G3106,G2669);
  and (G5237,G3107,G3108,G3281);
  and (G5238,G3793,G3802);
  and (G5239,G3825,G3834);
  and (G5240,G3852,G3859);
  and (G5241,G3765,G3776);
  not (G5242,G4077);
  not (G5243,G4227);
  or (G5244,G4044,G4260);
  or (G5245,G4045,G4261);
  or (G5246,G4046,G4262);
  or (G5247,G4047,G4263);
  not (G5248,G4323);
  not (G5249,G4562);
  not (G5250,G4554);
  not (G5251,G4606);
  or (G5252,G4425,G4677,G2182,G1479);
  not (G5253,G4664);
  not (G5254,G4648);
  not (G5255,G4642);
  or (G5256,G4426,G4680,G2201,G1499);
  not (G5257,G4658);
  not (G5258,G4636);
  not (G5259,G4630);
  not (G5260,G4624);
  not (G5261,G4681);
  not (G5262,G4684);
  and (G5263,G4507,G4530,G4531,G4532,G4533,G4709,G4710,G4711,G4712);
  and (G5264,G4183,G4508,G4534,G4535,G4536,G4713,G4714,G4715,G4716);
  and (G5265,G4719,G1548);
  and (G5266,G4727,G1623);
  or (G5267,G4733,G4734,G2187,G1484);
  or (G5268,G4735,G4736,G2188,G1485);
  or (G5269,G4737,G4738,G2189,G1486);
  or (G5270,G4678,G4739,G2190,G1487);
  or (G5271,G4740,G4741,G2195,G1492);
  or (G5272,G4742,G4743,G2196,G1493);
  or (G5273,G4744,G4745,G2197,G1494);
  or (G5274,G4679,G4746,G2198,G1495);
  and (G5275,G4766,G1520);
  and (G5276,G4767,G1548);
  and (G5277,G4768,G1548);
  and (G5278,G4769,G1548);
  and (G5279,G4770,G1595);
  and (G5280,G4771,G1623);
  and (G5281,G4772,G1623);
  and (G5282,G4773,G1623);
  and (G5283,G686,G4774);
  or (G5284,G4849,G4850);
  not (G5285,G4822);
  not (G5286,G4816);
  not (G5287,G4810);
  not (G5288,G4804);
  and (G5289,G689,G4851,G99);
  not (G5290,G4798);
  not (G5291,G4792);
  not (G5292,G4786);
  not (G5293,G4780);
  or (G5294,G4872,G4873,G2179,G1478);
  or (G5295,G4874,G4875,G2183,G1480);
  or (G5296,G4876,G4877,G2184,G1481);
  or (G5297,G4878,G4879,G2185,G1482);
  or (G5298,G4880,G4881,G2186,G1483);
  or (G5299,G4882,G4883,G2192,G1489);
  or (G5300,G4884,G4885,G2193,G1490);
  or (G5301,G4886,G4887,G2194,G1491);
  and (G5302,G4907,G1520);
  and (G5303,G4908,G1520);
  and (G5304,G4909,G1520);
  and (G5305,G4910,G1520);
  and (G5306,G4911,G1595);
  and (G5307,G4912,G1595);
  and (G5308,G4913,G1595);
  and (G5309,G4914,G1595);
  or (G5310,G4775,G5153,G2200,G1498);
  or (G5311,G4852,G5154,G2202,G1500);
  or (G5312,G5181,G5182,G2191,G1488);
  or (G5313,G5183,G5184,G2199,G1496);
  not (G5314,G5191);
  not (G5315,G5192);

endmodule
