// Benchmark "mymod" written by ABC on Sun Oct 29 19:31:54 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58,
    G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70, G71, G72,
    G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86,
    G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G109, G110, G111, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G124,
    G125, G126, G127, G128, G129, G130, G131, G132, G133, G134, G135, G136,
    G137, G138, G139, G140, G141, G142, G143, G144, G145, G146, G147, G148,
    G149, G150, G151, G152, G153, G154, G155, G156, G157,
    G2531, G2532, G2533, G2534, G2535, G2536, G2537, G2538, G2539, G2540,
    G2541, G2542, G2543, G2544, G2545, G2546, G2547, G2548, G2549, G2550,
    G2551, G2552, G2553, G2554, G2555, G2556, G2557, G2558, G2559, G2560,
    G2561, G2562, G2563, G2564, G2565, G2566, G2567, G2568, G2569, G2570,
    G2571, G2572, G2573, G2574, G2575, G2576, G2577, G2578, G2579, G2580,
    G2581, G2582, G2583, G2584, G2585, G2586, G2587, G2588, G2589, G2590,
    G2591, G2592, G2593, G2594  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70,
    G71, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98,
    G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G110,
    G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G133, G134,
    G135, G136, G137, G138, G139, G140, G141, G142, G143, G144, G145, G146,
    G147, G148, G149, G150, G151, G152, G153, G154, G155, G156, G157;
  output G2531, G2532, G2533, G2534, G2535, G2536, G2537, G2538, G2539, G2540,
    G2541, G2542, G2543, G2544, G2545, G2546, G2547, G2548, G2549, G2550,
    G2551, G2552, G2553, G2554, G2555, G2556, G2557, G2558, G2559, G2560,
    G2561, G2562, G2563, G2564, G2565, G2566, G2567, G2568, G2569, G2570,
    G2571, G2572, G2573, G2574, G2575, G2576, G2577, G2578, G2579, G2580,
    G2581, G2582, G2583, G2584, G2585, G2586, G2587, G2588, G2589, G2590,
    G2591, G2592, G2593, G2594;
  reg n1416_lo, n1419_lo, n1422_lo, n1425_lo, n1428_lo, n1431_lo, n1434_lo,
    n1437_lo, n1440_lo, n1443_lo, n1446_lo, n1449_lo, n1452_lo, n1455_lo,
    n1458_lo, n1464_lo, n1467_lo, n1470_lo, n1476_lo, n1479_lo, n1482_lo,
    n1488_lo, n1491_lo, n1494_lo, n1497_lo, n1500_lo, n1512_lo, n1515_lo,
    n1518_lo, n1521_lo, n1524_lo, n1527_lo, n1530_lo, n1533_lo, n1536_lo,
    n1539_lo, n1542_lo, n1545_lo, n1548_lo, n1551_lo, n1554_lo, n1560_lo,
    n1563_lo, n1566_lo, n1572_lo, n1575_lo, n1578_lo, n1584_lo, n1587_lo,
    n1590_lo, n1596_lo, n1599_lo, n1602_lo, n1608_lo, n1611_lo, n1614_lo,
    n1620_lo, n1623_lo, n1626_lo, n1632_lo, n1635_lo, n1638_lo, n1644_lo,
    n1647_lo, n1650_lo, n1656_lo, n1659_lo, n1662_lo, n1668_lo, n1671_lo,
    n1674_lo, n1677_lo, n1680_lo, n1683_lo, n1686_lo, n1692_lo, n1695_lo,
    n1698_lo, n1704_lo, n1707_lo, n1710_lo, n1716_lo, n1719_lo, n1722_lo,
    n1728_lo, n1731_lo, n1734_lo, n1740_lo, n1743_lo, n1746_lo, n1749_lo,
    n1752_lo, n1755_lo, n1758_lo, n1761_lo, n1764_lo, n1776_lo, n1779_lo,
    n1788_lo, n1791_lo, n1794_lo, n1797_lo, n1800_lo, n1812_lo, n1824_lo,
    n1836_lo, n1848_lo, n1860_lo, n1872_lo, n1884_lo, n1896_lo, n1899_lo,
    n1908_lo, n1911_lo, n1920_lo, n1923_lo, n1926_lo, n1929_lo, n1932_lo,
    n1944_lo, n1956_lo, n1968_lo, n1980_lo, n1992_lo, n2004_lo, n2016_lo,
    n2019_lo, n2028_lo, n2031_lo, n2040_lo, n2043_lo, n2046_lo, n2049_lo,
    n2052_lo, n2064_lo, n2076_lo, n2088_lo, n2100_lo, n2112_lo, n2124_lo,
    n2136_lo, n2148_lo, n2151_lo, n2160_lo, n2163_lo, n2172_lo, n2175_lo,
    n2178_lo, n2181_lo, n2184_lo, n2196_lo, n2208_lo, n2220_lo, n2232_lo,
    n2244_lo, n2256_lo, n2268_lo, n2280_lo, n2283_lo, n2292_lo, n2295_lo,
    n2298_lo, n2301_lo, n2304_lo, n2316_lo, n2319_lo, n2322_lo, n2325_lo,
    n2328_lo, n2331_lo, n2340_lo, n2343_lo, n2376_lo, n2379_lo, n2388_lo,
    n2400_lo, n2412_lo, n2415_lo, n2424_lo, n2436_lo, n2439_lo, n2442_lo,
    n2445_lo, n2448_lo, n2451_lo, n2460_lo, n2463_lo, n2496_lo, n2499_lo,
    n2508_lo, n2520_lo, n2532_lo, n2535_lo, n2544_lo, n2556_lo, n2559_lo,
    n2562_lo, n2565_lo, n2568_lo, n2571_lo, n2580_lo, n2583_lo, n2616_lo,
    n2619_lo, n2628_lo, n2640_lo, n2652_lo, n2655_lo, n2664_lo, n2676_lo,
    n2679_lo, n2682_lo, n2685_lo, n2688_lo, n2691_lo, n2700_lo, n2703_lo,
    n2736_lo, n2739_lo, n2748_lo, n2760_lo, n2772_lo, n2775_lo, n2784_lo,
    n2787_lo, n2790_lo, n2793_lo, n2796_lo, n2799_lo, n2802_lo, n2805_lo,
    n2808_lo, n2820_lo, n2823_lo, n2826_lo, n2832_lo, n2835_lo, n2838_lo,
    n2841_lo, n2844_lo, n2856_lo, n2859_lo, n2862_lo, n2865_lo, n2868_lo,
    n2871_lo, n2874_lo, n2877_lo, n2880_lo, n2883_lo, n2886_lo, n2889_lo,
    n2892_lo, n2895_lo, n2898_lo, n2901_lo, n2904_lo, n2907_lo, n2916_lo,
    n2928_lo, n2940_lo, n2952_lo, n2955_lo, n2964_lo, n2976_lo, n2988_lo,
    n2991_lo, n3000_lo, n3003_lo, n3012_lo, n3015_lo, n3024_lo, n3027_lo,
    n3036_lo, n3039_lo, n3048_lo, n3051_lo, n3054_lo, n3057_lo, n3060_lo,
    n3072_lo, n3081_lo, n3084_lo, n3087_lo, n3093_lo, n3096_lo, n3105_lo,
    n3108_lo, n3117_lo, n3120_lo, n3123_lo, n3126_lo, n3129_lo, n3132_lo,
    n3135_lo, n3138_lo, n3141_lo, n3168_lo, n3171_lo, n3174_lo, n3177_lo,
    n3180_lo, n3183_lo, n3192_lo, n3195_lo, n3204_lo, n3207_lo, n3216_lo,
    n3219_lo, n3228_lo, n3231_lo, n3240_lo, n3243_lo, n3252_lo, n3255_lo,
    n3258_lo, n3264_lo, n3267_lo, n3270_lo, n3276_lo, n3279_lo, n3282_lo,
    n3288_lo, n3291_lo, n3294_lo, n4537_o2, n4538_o2, n4710_o2, n4711_o2,
    n1211_inv, n1214_inv, n1217_inv, n1220_inv, n4927_o2, n4928_o2,
    n1229_inv, n1232_inv, n1235_inv, n5178_o2, n5179_o2, n5477_o2,
    n5478_o2, n5479_o2, n5222_o2, n5223_o2, n5553_o2, n5554_o2, G491_o2,
    n2922_lo_buf_o2, n2946_lo_buf_o2, n2970_lo_buf_o2, n2982_lo_buf_o2,
    n3066_lo_buf_o2, n3078_lo_buf_o2, n3102_lo_buf_o2, n3114_lo_buf_o2,
    G1321_o2, G1033_o2, G1030_o2, G1072_o2, n1304_inv, n1307_inv,
    n2958_lo_buf_o2, n2994_lo_buf_o2, n3006_lo_buf_o2, n3030_lo_buf_o2,
    n3042_lo_buf_o2, n3090_lo_buf_o2, n1328_inv, n1331_inv, n1334_inv,
    n1337_inv, n1340_inv, n1343_inv, n1346_inv, n1349_inv, G1036_o2,
    G1062_o2, G1067_o2, G1014_o2, n1364_inv, n1367_inv, n3018_lo_buf_o2,
    G766_o2, n1376_inv, n1379_inv, n1382_inv, n1385_inv, n1388_inv,
    n1391_inv, G1017_o2, G1008_o2, n1400_inv, n1403_inv, n2910_lo_buf_o2,
    n1409_inv, G2138_o2, G2147_o2, n1418_inv, G1137_o2, G1329_o2, G374_o2,
    G386_o2, G663_o2, G674_o2, G578_o2, G575_o2, G2505_o2, n1448_inv,
    G987_o2, G984_o2, G1862_o2, G1859_o2, G1260_o2, G1865_o2, G2073_o2,
    G1402_o2, G2048_o2, G2276_o2, n1481_inv, G2141_o2, G2008_o2, G2011_o2,
    G2150_o2, G2026_o2, G2029_o2, G2023_o2, G2041_o2, G2017_o2, G2020_o2,
    G2035_o2, G2038_o2, G2228_o2, G2231_o2, G2234_o2, G2237_o2, G1904_o2,
    G1907_o2, G1928_o2, G1931_o2, G1893_o2, G1896_o2, G1899_o2, G1937_o2,
    G1940_o2, G1943_o2, G1336_o2, G1996_o2, G1999_o2, G2002_o2, G2005_o2,
    G2014_o2, G2032_o2, G1076_o2, G1002_o2, G998_o2, G1890_o2, G1934_o2,
    G1044_o2, G1039_o2, n1770_lo_buf_o2, G342_o2, G354_o2, G1193_o2,
    n3234_lo_buf_o2, n3246_lo_buf_o2, G783_o2, G786_o2, G792_o2, G795_o2,
    G815_o2, G818_o2, G824_o2, G827_o2, G789_o2, G798_o2, G801_o2, G807_o2,
    G812_o2, G821_o2, G804_o2, G780_o2, G1231_o2, G1572_o2, G1377_o2,
    G1253_o2, G1359_o2, G1258_o2, G1367_o2, G1358_o2, G1366_o2, G2057_o2,
    G2117_o2, G2118_o2, G1254_o2, G1259_o2, G2058_o2, G405_o2, G417_o2,
    G1269_o2, G1275_o2, G1287_o2, G1266_o2, G1272_o2, G1278_o2, G1281_o2,
    G1284_o2, G1290_o2, G1293_o2, G1299_o2, G1305_o2, G1296_o2, G1302_o2,
    G1308_o2, G1311_o2, G811_o2, G810_o2, G1728_o2, G2512_o2, G1114_o2,
    G1113_o2, G1992_o2, G1991_o2, G1426_o2, G1966_o2, G2211_o2, G1509_o2,
    G2153_o2, G2329_o2, G1540_o2, G2167_o2, G2191_o2, G1234_o2, G1132_o2,
    G1129_o2, G2088_o2, G2106_o2, G1314_o2, G636_o2, G647_o2,
    n3186_lo_buf_o2, n3198_lo_buf_o2, n3210_lo_buf_o2, n3222_lo_buf_o2,
    G1225_o2, G1342_o2, G1222_o2, G1228_o2, G1348_o2, G1345_o2, G1351_o2,
    G2242_o2, G2260_o2, G1374_o2, G1537_o2, G301_o2, G313_o2, G2365_o2,
    G2255_o2, G2253_o2, G2395_o2, G2272_o2, G2270_o2, G2245_o2, G2262_o2,
    G2249_o2, G2247_o2, G2266_o2, G2264_o2, G2403_o2, G2401_o2, G2410_o2,
    G2408_o2, G2306_o2, G2305_o2, G2314_o2, G2313_o2, G2303_o2, G2302_o2,
    G2301_o2, G2311_o2, G2310_o2, G2309_o2, G2404_o2, G2411_o2, G2420_o2,
    G2419_o2, G2433_o2, G2432_o2, G402_o2, G403_o2, G1053_o2, G1049_o2,
    n2003_inv, G1364_o2, G1079_o2, G1478_o2, G707_o2, G718_o2, G2417_o2,
    G2414_o2, G2431_o2, G2428_o2, G1653_o2, G2213_o2, G2221_o2, G2250_o2,
    G2267_o2, G1365_o2, G1368_o2, G1371_o2, G2218_o2, G2225_o2,
    n1503_lo_buf_o2, n1863_lo_buf_o2, n1887_lo_buf_o2, n1983_lo_buf_o2,
    n2007_lo_buf_o2, n2115_lo_buf_o2, n2139_lo_buf_o2, n2247_lo_buf_o2,
    n2271_lo_buf_o2, n2919_lo_buf_o2, n2943_lo_buf_o2, n2967_lo_buf_o2,
    n2979_lo_buf_o2, n3063_lo_buf_o2, n3075_lo_buf_o2, n3099_lo_buf_o2,
    n3111_lo_buf_o2, G878_o2, G875_o2, G661_o2, G660_o2, G879_o2, G876_o2,
    G1320_o2, G941_o2, G732_o2, G942_o2, G1493_o2, G1498_o2, G877_o2,
    G874_o2, n1806_lo_buf_o2, n1878_lo_buf_o2, n1938_lo_buf_o2,
    n1998_lo_buf_o2, n2058_lo_buf_o2, n2130_lo_buf_o2, n2190_lo_buf_o2,
    n2262_lo_buf_o2, n2310_lo_buf_o2, n2406_lo_buf_o2, n2430_lo_buf_o2,
    n2526_lo_buf_o2, n2550_lo_buf_o2, n2646_lo_buf_o2, n2670_lo_buf_o2,
    n2766_lo_buf_o2, G603_o2, G614_o2, G1026_o2, G1021_o2, G940_o2,
    G1636_o2, G1684_o2, n2352_lo_buf_o2, n2364_lo_buf_o2, n2472_lo_buf_o2,
    n2484_lo_buf_o2, n2592_lo_buf_o2, n2604_lo_buf_o2, n2712_lo_buf_o2,
    n2724_lo_buf_o2, n3150_lo_buf_o2, n3162_lo_buf_o2;
  wire new_new_n1576__, new_new_n1578__, new_new_n1580__, new_new_n1582__,
    new_new_n1584__, new_new_n1586__, new_new_n1588__, new_new_n1590__,
    new_new_n1592__, new_new_n1594__, new_new_n1596__, new_new_n1598__,
    new_new_n1600__, new_new_n1602__, new_new_n1604__, new_new_n1606__,
    new_new_n1608__, new_new_n1610__, new_new_n1612__, new_new_n1614__,
    new_new_n1616__, new_new_n1618__, new_new_n1620__, new_new_n1622__,
    new_new_n1624__, new_new_n1626__, new_new_n1628__, new_new_n1630__,
    new_new_n1632__, new_new_n1634__, new_new_n1636__, new_new_n1638__,
    new_new_n1640__, new_new_n1642__, new_new_n1644__, new_new_n1646__,
    new_new_n1648__, new_new_n1650__, new_new_n1652__, new_new_n1654__,
    new_new_n1656__, new_new_n1658__, new_new_n1660__, new_new_n1662__,
    new_new_n1664__, new_new_n1666__, new_new_n1668__, new_new_n1670__,
    new_new_n1672__, new_new_n1674__, new_new_n1676__, new_new_n1678__,
    new_new_n1680__, new_new_n1682__, new_new_n1684__, new_new_n1686__,
    new_new_n1688__, new_new_n1690__, new_new_n1692__, new_new_n1694__,
    new_new_n1696__, new_new_n1698__, new_new_n1700__, new_new_n1702__,
    new_new_n1704__, new_new_n1706__, new_new_n1708__, new_new_n1710__,
    new_new_n1712__, new_new_n1714__, new_new_n1716__, new_new_n1718__,
    new_new_n1720__, new_new_n1722__, new_new_n1724__, new_new_n1726__,
    new_new_n1728__, new_new_n1730__, new_new_n1732__, new_new_n1734__,
    new_new_n1736__, new_new_n1738__, new_new_n1740__, new_new_n1742__,
    new_new_n1744__, new_new_n1746__, new_new_n1748__, new_new_n1750__,
    new_new_n1752__, new_new_n1754__, new_new_n1756__, new_new_n1758__,
    new_new_n1760__, new_new_n1762__, new_new_n1764__, new_new_n1766__,
    new_new_n1768__, new_new_n1770__, new_new_n1772__, new_new_n1774__,
    new_new_n1776__, new_new_n1778__, new_new_n1780__, new_new_n1782__,
    new_new_n1784__, new_new_n1786__, new_new_n1788__, new_new_n1790__,
    new_new_n1792__, new_new_n1794__, new_new_n1796__, new_new_n1798__,
    new_new_n1800__, new_new_n1802__, new_new_n1804__, new_new_n1806__,
    new_new_n1808__, new_new_n1810__, new_new_n1812__, new_new_n1814__,
    new_new_n1816__, new_new_n1818__, new_new_n1820__, new_new_n1822__,
    new_new_n1824__, new_new_n1826__, new_new_n1828__, new_new_n1830__,
    new_new_n1832__, new_new_n1834__, new_new_n1836__, new_new_n1838__,
    new_new_n1840__, new_new_n1842__, new_new_n1844__, new_new_n1846__,
    new_new_n1848__, new_new_n1850__, new_new_n1852__, new_new_n1854__,
    new_new_n1856__, new_new_n1858__, new_new_n1860__, new_new_n1862__,
    new_new_n1864__, new_new_n1866__, new_new_n1868__, new_new_n1870__,
    new_new_n1872__, new_new_n1874__, new_new_n1876__, new_new_n1878__,
    new_new_n1880__, new_new_n1882__, new_new_n1884__, new_new_n1886__,
    new_new_n1888__, new_new_n1890__, new_new_n1892__, new_new_n1894__,
    new_new_n1896__, new_new_n1898__, new_new_n1900__, new_new_n1902__,
    new_new_n1905__, new_new_n1906__, new_new_n1908__, new_new_n1910__,
    new_new_n1912__, new_new_n1914__, new_new_n1916__, new_new_n1918__,
    new_new_n1920__, new_new_n1922__, new_new_n1924__, new_new_n1926__,
    new_new_n1928__, new_new_n1930__, new_new_n1932__, new_new_n1934__,
    new_new_n1936__, new_new_n1939__, new_new_n1940__, new_new_n1942__,
    new_new_n1944__, new_new_n1946__, new_new_n1949__, new_new_n1950__,
    new_new_n1952__, new_new_n1954__, new_new_n1956__, new_new_n1958__,
    new_new_n1960__, new_new_n1962__, new_new_n1965__, new_new_n1966__,
    new_new_n1968__, new_new_n1970__, new_new_n1971__, new_new_n1972__,
    new_new_n1974__, new_new_n1976__, new_new_n1978__, new_new_n1980__,
    new_new_n1982__, new_new_n1984__, new_new_n1986__, new_new_n1988__,
    new_new_n1990__, new_new_n1992__, new_new_n1994__, new_new_n1996__,
    new_new_n1998__, new_new_n2000__, new_new_n2002__, new_new_n2004__,
    new_new_n2006__, new_new_n2008__, new_new_n2010__, new_new_n2012__,
    new_new_n2014__, new_new_n2016__, new_new_n2018__, new_new_n2020__,
    new_new_n2022__, new_new_n2024__, new_new_n2026__, new_new_n2028__,
    new_new_n2030__, new_new_n2033__, new_new_n2034__, new_new_n2036__,
    new_new_n2038__, new_new_n2039__, new_new_n2040__, new_new_n2042__,
    new_new_n2044__, new_new_n2046__, new_new_n2048__, new_new_n2050__,
    new_new_n2052__, new_new_n2054__, new_new_n2056__, new_new_n2058__,
    new_new_n2060__, new_new_n2062__, new_new_n2064__, new_new_n2066__,
    new_new_n2068__, new_new_n2071__, new_new_n2072__, new_new_n2074__,
    new_new_n2076__, new_new_n2079__, new_new_n2080__, new_new_n2081__,
    new_new_n2082__, new_new_n2084__, new_new_n2086__, new_new_n2088__,
    new_new_n2090__, new_new_n2093__, new_new_n2094__, new_new_n2096__,
    new_new_n2098__, new_new_n2100__, new_new_n2102__, new_new_n2104__,
    new_new_n2106__, new_new_n2108__, new_new_n2110__, new_new_n2112__,
    new_new_n2114__, new_new_n2116__, new_new_n2118__, new_new_n2120__,
    new_new_n2122__, new_new_n2125__, new_new_n2126__, new_new_n2128__,
    new_new_n2130__, new_new_n2132__, new_new_n2134__, new_new_n2136__,
    new_new_n2138__, new_new_n2140__, new_new_n2142__, new_new_n2144__,
    new_new_n2146__, new_new_n2148__, new_new_n2150__, new_new_n2152__,
    new_new_n2155__, new_new_n2156__, new_new_n2158__, new_new_n2160__,
    new_new_n2162__, new_new_n2164__, new_new_n2166__, new_new_n2168__,
    new_new_n2170__, new_new_n2172__, new_new_n2174__, new_new_n2176__,
    new_new_n2178__, new_new_n2180__, new_new_n2182__, new_new_n2184__,
    new_new_n2187__, new_new_n2188__, new_new_n2190__, new_new_n2192__,
    new_new_n2194__, new_new_n2196__, new_new_n2198__, new_new_n2200__,
    new_new_n2202__, new_new_n2204__, new_new_n2206__, new_new_n2208__,
    new_new_n2210__, new_new_n2212__, new_new_n2214__, new_new_n2216__,
    new_new_n2218__, new_new_n2220__, new_new_n2222__, new_new_n2225__,
    new_new_n2226__, new_new_n2228__, new_new_n2230__, new_new_n2232__,
    new_new_n2234__, new_new_n2236__, new_new_n2238__, new_new_n2240__,
    new_new_n2242__, new_new_n2244__, new_new_n2246__, new_new_n2248__,
    new_new_n2250__, new_new_n2252__, new_new_n2255__, new_new_n2256__,
    new_new_n2258__, new_new_n2260__, new_new_n2262__, new_new_n2264__,
    new_new_n2266__, new_new_n2268__, new_new_n2270__, new_new_n2272__,
    new_new_n2274__, new_new_n2276__, new_new_n2278__, new_new_n2280__,
    new_new_n2282__, new_new_n2285__, new_new_n2286__, new_new_n2288__,
    new_new_n2290__, new_new_n2292__, new_new_n2294__, new_new_n2296__,
    new_new_n2298__, new_new_n2300__, new_new_n2302__, new_new_n2304__,
    new_new_n2306__, new_new_n2308__, new_new_n2310__, new_new_n2312__,
    new_new_n2315__, new_new_n2316__, new_new_n2318__, new_new_n2320__,
    new_new_n2322__, new_new_n2324__, new_new_n2326__, new_new_n2328__,
    new_new_n2330__, new_new_n2332__, new_new_n2334__, new_new_n2336__,
    new_new_n2338__, new_new_n2340__, new_new_n2342__, new_new_n2343__,
    new_new_n2344__, new_new_n2346__, new_new_n2348__, new_new_n2351__,
    new_new_n2352__, new_new_n2353__, new_new_n2354__, new_new_n2356__,
    new_new_n2358__, new_new_n2359__, new_new_n2360__, new_new_n2362__,
    new_new_n2364__, new_new_n2366__, new_new_n2367__, new_new_n2368__,
    new_new_n2369__, new_new_n2370__, new_new_n2372__, new_new_n2374__,
    new_new_n2376__, new_new_n2377__, new_new_n2378__, new_new_n2380__,
    new_new_n2382__, new_new_n2384__, new_new_n2385__, new_new_n2386__,
    new_new_n2388__, new_new_n2390__, new_new_n2392__, new_new_n2393__,
    new_new_n2394__, new_new_n2396__, new_new_n2398__, new_new_n2401__,
    new_new_n2402__, new_new_n2404__, new_new_n2406__, new_new_n2408__,
    new_new_n2410__, new_new_n2412__, new_new_n2414__, new_new_n2415__,
    new_new_n2416__, new_new_n2418__, new_new_n2420__, new_new_n2422__,
    new_new_n2424__, new_new_n2426__, new_new_n2428__, new_new_n2430__,
    new_new_n2431__, new_new_n2432__, new_new_n2434__, new_new_n2435__,
    new_new_n2436__, new_new_n2438__, new_new_n2439__, new_new_n2440__,
    new_new_n2442__, new_new_n2444__, new_new_n2447__, new_new_n2448__,
    new_new_n2450__, new_new_n2453__, new_new_n2454__, new_new_n2456__,
    new_new_n2457__, new_new_n2459__, new_new_n2460__, new_new_n2463__,
    new_new_n2464__, new_new_n2467__, new_new_n2468__, new_new_n2470__,
    new_new_n2472__, new_new_n2474__, new_new_n2475__, new_new_n2476__,
    new_new_n2478__, new_new_n2480__, new_new_n2482__, new_new_n2483__,
    new_new_n2484__, new_new_n2486__, new_new_n2488__, new_new_n2490__,
    new_new_n2491__, new_new_n2492__, new_new_n2494__, new_new_n2496__,
    new_new_n2498__, new_new_n2500__, new_new_n2502__, new_new_n2504__,
    new_new_n2506__, new_new_n2508__, new_new_n2510__, new_new_n2512__,
    new_new_n2514__, new_new_n2516__, new_new_n2518__, new_new_n2520__,
    new_new_n2521__, new_new_n2522__, new_new_n2524__, new_new_n2526__,
    new_new_n2527__, new_new_n2528__, new_new_n2530__, new_new_n2532__,
    new_new_n2533__, new_new_n2534__, new_new_n2536__, new_new_n2538__,
    new_new_n2539__, new_new_n2541__, new_new_n2543__, new_new_n2545__,
    new_new_n2547__, new_new_n2548__, new_new_n2550__, new_new_n2552__,
    new_new_n2554__, new_new_n2557__, new_new_n2558__, new_new_n2559__,
    new_new_n2560__, new_new_n2562__, new_new_n2564__, new_new_n2566__,
    new_new_n2567__, new_new_n2568__, new_new_n2569__, new_new_n2570__,
    new_new_n2571__, new_new_n2573__, new_new_n2574__, new_new_n2575__,
    new_new_n2576__, new_new_n2577__, new_new_n2578__, new_new_n2580__,
    new_new_n2582__, new_new_n2584__, new_new_n2586__, new_new_n2587__,
    new_new_n2588__, new_new_n2589__, new_new_n2590__, new_new_n2591__,
    new_new_n2592__, new_new_n2593__, new_new_n2594__, new_new_n2595__,
    new_new_n2596__, new_new_n2597__, new_new_n2598__, new_new_n2599__,
    new_new_n2600__, new_new_n2601__, new_new_n2602__, new_new_n2603__,
    new_new_n2604__, new_new_n2606__, new_new_n2608__, new_new_n2610__,
    new_new_n2612__, new_new_n2614__, new_new_n2615__, new_new_n2616__,
    new_new_n2617__, new_new_n2618__, new_new_n2619__, new_new_n2620__,
    new_new_n2621__, new_new_n2622__, new_new_n2623__, new_new_n2624__,
    new_new_n2625__, new_new_n2626__, new_new_n2628__, new_new_n2630__,
    new_new_n2632__, new_new_n2634__, new_new_n2636__, new_new_n2638__,
    new_new_n2640__, new_new_n2642__, new_new_n2644__, new_new_n2646__,
    new_new_n2648__, new_new_n2650__, new_new_n2652__, new_new_n2654__,
    new_new_n2655__, new_new_n2657__, new_new_n2658__, new_new_n2660__,
    new_new_n2662__, new_new_n2664__, new_new_n2666__, new_new_n2668__,
    new_new_n2670__, new_new_n2672__, new_new_n2673__, new_new_n2674__,
    new_new_n2676__, new_new_n2678__, new_new_n2679__, new_new_n2680__,
    new_new_n2682__, new_new_n2683__, new_new_n2684__, new_new_n2685__,
    new_new_n2686__, new_new_n2688__, new_new_n2689__, new_new_n2690__,
    new_new_n2691__, new_new_n2692__, new_new_n2693__, new_new_n2694__,
    new_new_n2695__, new_new_n2696__, new_new_n2697__, new_new_n2698__,
    new_new_n2699__, new_new_n2700__, new_new_n2701__, new_new_n2702__,
    new_new_n2703__, new_new_n2705__, new_new_n2706__, new_new_n2707__,
    new_new_n2708__, new_new_n2709__, new_new_n2710__, new_new_n2711__,
    new_new_n2712__, new_new_n2713__, new_new_n2714__, new_new_n2715__,
    new_new_n2717__, new_new_n2718__, new_new_n2721__, new_new_n2722__,
    new_new_n2725__, new_new_n2726__, new_new_n2728__, new_new_n2730__,
    new_new_n2731__, new_new_n2732__, new_new_n2733__, new_new_n2734__,
    new_new_n2735__, new_new_n2736__, new_new_n2737__, new_new_n2738__,
    new_new_n2739__, new_new_n2740__, new_new_n2741__, new_new_n2742__,
    new_new_n2744__, new_new_n2746__, new_new_n2748__, new_new_n2750__,
    new_new_n2752__, new_new_n2754__, new_new_n2755__, new_new_n2756__,
    new_new_n2757__, new_new_n2758__, new_new_n2759__, new_new_n2760__,
    new_new_n2761__, new_new_n2762__, new_new_n2763__, new_new_n2764__,
    new_new_n2765__, new_new_n2766__, new_new_n2767__, new_new_n2768__,
    new_new_n2769__, new_new_n2771__, new_new_n2773__, new_new_n2775__,
    new_new_n2777__, new_new_n2779__, new_new_n2781__, new_new_n2782__,
    new_new_n2783__, new_new_n2784__, new_new_n2785__, new_new_n2786__,
    new_new_n2787__, new_new_n2788__, new_new_n2789__, new_new_n2790__,
    new_new_n2791__, new_new_n2792__, new_new_n2794__, new_new_n2796__,
    new_new_n2798__, new_new_n2799__, new_new_n2800__, new_new_n2803__,
    new_new_n2805__, new_new_n2806__, new_new_n2808__, new_new_n2810__,
    new_new_n2811__, new_new_n2813__, new_new_n2815__, new_new_n2816__,
    new_new_n2817__, new_new_n2818__, new_new_n2819__, new_new_n2820__,
    new_new_n2821__, new_new_n2822__, new_new_n2823__, new_new_n2824__,
    new_new_n2825__, new_new_n2826__, new_new_n2827__, new_new_n2828__,
    new_new_n2829__, new_new_n2830__, new_new_n2831__, new_new_n2832__,
    new_new_n2833__, new_new_n2834__, new_new_n2835__, new_new_n2836__,
    new_new_n2837__, new_new_n2838__, new_new_n2839__, new_new_n2840__,
    new_new_n2841__, new_new_n2842__, new_new_n2843__, new_new_n2844__,
    new_new_n2845__, new_new_n2846__, new_new_n2847__, new_new_n2848__,
    new_new_n2849__, new_new_n2850__, new_new_n2851__, new_new_n2852__,
    new_new_n2853__, new_new_n2854__, new_new_n2855__, new_new_n2856__,
    new_new_n2857__, new_new_n2858__, new_new_n2859__, new_new_n2860__,
    new_new_n2861__, new_new_n2862__, new_new_n2863__, new_new_n2864__,
    new_new_n2865__, new_new_n2866__, new_new_n2867__, new_new_n2868__,
    new_new_n2869__, new_new_n2870__, new_new_n2871__, new_new_n2872__,
    new_new_n2873__, new_new_n2874__, new_new_n2875__, new_new_n2876__,
    new_new_n2877__, new_new_n2878__, new_new_n2879__, new_new_n2880__,
    new_new_n2881__, new_new_n2882__, new_new_n2883__, new_new_n2885__,
    new_new_n2887__, new_new_n2888__, new_new_n2889__, new_new_n2890__,
    new_new_n2891__, new_new_n2892__, new_new_n2893__, new_new_n2894__,
    new_new_n2895__, new_new_n2896__, new_new_n2897__, new_new_n2898__,
    new_new_n2899__, new_new_n2900__, new_new_n2901__, new_new_n2902__,
    new_new_n2903__, new_new_n2904__, new_new_n2905__, new_new_n2906__,
    new_new_n2907__, new_new_n2908__, new_new_n2909__, new_new_n2910__,
    new_new_n2911__, new_new_n2912__, new_new_n2913__, new_new_n2914__,
    new_new_n2915__, new_new_n2916__, new_new_n2917__, new_new_n2918__,
    new_new_n2919__, new_new_n2920__, new_new_n2921__, new_new_n2922__,
    new_new_n2923__, new_new_n2924__, new_new_n2925__, new_new_n2926__,
    new_new_n2928__, new_new_n2929__, new_new_n2930__, new_new_n2931__,
    new_new_n2932__, new_new_n2933__, new_new_n2934__, new_new_n2935__,
    new_new_n2936__, new_new_n2939__, new_new_n2940__, new_new_n2943__,
    new_new_n2944__, new_new_n2947__, new_new_n2948__, new_new_n2949__,
    new_new_n2951__, new_new_n2953__, new_new_n2954__, new_new_n2955__,
    new_new_n2956__, new_new_n2957__, new_new_n2958__, new_new_n2959__,
    new_new_n2960__, new_new_n2962__, new_new_n2964__, new_new_n2965__,
    new_new_n2966__, new_new_n2968__, new_new_n2970__, new_new_n2971__,
    new_new_n2972__, new_new_n2973__, new_new_n2974__, new_new_n2975__,
    new_new_n2976__, new_new_n2977__, new_new_n2978__, new_new_n2979__,
    new_new_n2980__, new_new_n2981__, new_new_n2982__, new_new_n2983__,
    new_new_n2984__, new_new_n2985__, new_new_n2986__, new_new_n2987__,
    new_new_n2988__, new_new_n2989__, new_new_n2990__, new_new_n2991__,
    new_new_n2992__, new_new_n2993__, new_new_n2994__, new_new_n2995__,
    new_new_n2996__, new_new_n2997__, new_new_n2998__, new_new_n2999__,
    new_new_n3000__, new_new_n3001__, new_new_n3002__, new_new_n3003__,
    new_new_n3004__, new_new_n3005__, new_new_n3006__, new_new_n3007__,
    new_new_n3008__, new_new_n3009__, new_new_n3010__, new_new_n3011__,
    new_new_n3012__, new_new_n3013__, new_new_n3014__, new_new_n3015__,
    new_new_n3017__, new_new_n3019__, new_new_n3021__, new_new_n3023__,
    new_new_n3025__, new_new_n3027__, new_new_n3028__, new_new_n3029__,
    new_new_n3030__, new_new_n3031__, new_new_n3032__, new_new_n3033__,
    new_new_n3034__, new_new_n3035__, new_new_n3036__, new_new_n3037__,
    new_new_n3038__, new_new_n3039__, new_new_n3040__, new_new_n3041__,
    new_new_n3042__, new_new_n3043__, new_new_n3044__, new_new_n3046__,
    new_new_n3048__, new_new_n3050__, new_new_n3052__, new_new_n3054__,
    new_new_n3056__, new_new_n3057__, new_new_n3058__, new_new_n3059__,
    new_new_n3060__, new_new_n3061__, new_new_n3062__, new_new_n3063__,
    new_new_n3064__, new_new_n3065__, new_new_n3066__, new_new_n3067__,
    new_new_n3068__, new_new_n3069__, new_new_n3070__, new_new_n3071__,
    new_new_n3072__, new_new_n3073__, new_new_n3074__, new_new_n3075__,
    new_new_n3076__, new_new_n3077__, new_new_n3078__, new_new_n3079__,
    new_new_n3080__, new_new_n3081__, new_new_n3082__, new_new_n3083__,
    new_new_n3084__, new_new_n3086__, new_new_n3088__, new_new_n3089__,
    new_new_n3090__, new_new_n3091__, new_new_n3092__, new_new_n3093__,
    new_new_n3094__, new_new_n3095__, new_new_n3096__, new_new_n3097__,
    new_new_n3098__, new_new_n3099__, new_new_n3100__, new_new_n3101__,
    new_new_n3102__, new_new_n3104__, new_new_n3106__, new_new_n3107__,
    new_new_n3108__, new_new_n3109__, new_new_n3110__, new_new_n3111__,
    new_new_n3113__, new_new_n3115__, new_new_n3117__, new_new_n3118__,
    new_new_n3119__, new_new_n3120__, new_new_n3121__, new_new_n3122__,
    new_new_n3123__, new_new_n3124__, new_new_n3125__, new_new_n3126__,
    new_new_n3127__, new_new_n3128__, new_new_n3129__, new_new_n3130__,
    new_new_n3131__, new_new_n3132__, new_new_n3133__, new_new_n3134__,
    new_new_n3135__, new_new_n3136__, new_new_n3137__, new_new_n3138__,
    new_new_n3140__, new_new_n3142__, new_new_n3143__, new_new_n3144__,
    new_new_n3145__, new_new_n3146__, new_new_n3148__, new_new_n3150__,
    new_new_n3152__, new_new_n3154__, new_new_n3156__, new_new_n3158__,
    new_new_n3160__, new_new_n3162__, new_new_n3163__, new_new_n3164__,
    new_new_n3166__, new_new_n3168__, new_new_n3170__, new_new_n3171__,
    new_new_n3172__, new_new_n3173__, new_new_n3174__, new_new_n3176__,
    new_new_n3178__, new_new_n3180__, new_new_n3181__, new_new_n3182__,
    new_new_n3184__, new_new_n3185__, new_new_n3186__, new_new_n3188__,
    new_new_n3189__, new_new_n3190__, new_new_n3192__, new_new_n3193__,
    new_new_n3194__, new_new_n3196__, new_new_n3198__, new_new_n3200__,
    new_new_n3202__, new_new_n3204__, new_new_n3206__, new_new_n3208__,
    new_new_n3210__, new_new_n3211__, new_new_n3212__, new_new_n3213__,
    new_new_n3214__, new_new_n3216__, new_new_n3218__, new_new_n3220__,
    new_new_n3221__, new_new_n3222__, new_new_n3223__, new_new_n3224__,
    new_new_n3227__, new_new_n3228__, new_new_n3231__, new_new_n3232__,
    new_new_n3235__, new_new_n3236__, new_new_n3239__, new_new_n3240__,
    new_new_n3241__, new_new_n3242__, new_new_n3243__, new_new_n3244__,
    new_new_n3245__, new_new_n3246__, new_new_n3247__, new_new_n3248__,
    new_new_n3249__, new_new_n3250__, new_new_n3251__, new_new_n3252__,
    new_new_n3253__, new_new_n3254__, new_new_n3255__, new_new_n3256__,
    new_new_n3257__, new_new_n3258__, new_new_n3259__, new_new_n3260__,
    new_new_n3261__, new_new_n3262__, new_new_n3263__, new_new_n3264__,
    new_new_n3265__, new_new_n3266__, new_new_n3267__, new_new_n3268__,
    new_new_n3269__, new_new_n3270__, new_new_n3271__, new_new_n3272__,
    new_new_n3273__, new_new_n3274__, new_new_n3275__, new_new_n3276__,
    new_new_n3277__, new_new_n3278__, new_new_n3279__, new_new_n3280__,
    new_new_n3281__, new_new_n3282__, new_new_n3283__, new_new_n3284__,
    new_new_n3285__, new_new_n3286__, new_new_n3287__, new_new_n3288__,
    new_new_n3289__, new_new_n3290__, new_new_n3291__, new_new_n3292__,
    new_new_n3293__, new_new_n3294__, new_new_n3295__, new_new_n3296__,
    new_new_n3297__, new_new_n3298__, new_new_n3299__, new_new_n3300__,
    new_new_n3301__, new_new_n3302__, new_new_n3303__, new_new_n3304__,
    new_new_n3305__, new_new_n3306__, new_new_n3307__, new_new_n3308__,
    new_new_n3309__, new_new_n3310__, new_new_n3311__, new_new_n3312__,
    new_new_n3313__, new_new_n3314__, new_new_n3315__, new_new_n3316__,
    new_new_n3317__, new_new_n3318__, new_new_n3319__, new_new_n3320__,
    new_new_n3321__, new_new_n3322__, new_new_n3323__, new_new_n3324__,
    new_new_n3325__, new_new_n3326__, new_new_n3327__, new_new_n3328__,
    new_new_n3329__, new_new_n3330__, new_new_n3331__, new_new_n3332__,
    new_new_n3333__, new_new_n3334__, new_new_n3335__, new_new_n3336__,
    new_new_n3337__, new_new_n3338__, new_new_n3339__, new_new_n3340__,
    new_new_n3341__, new_new_n3342__, new_new_n3343__, new_new_n3344__,
    new_new_n3345__, new_new_n3346__, new_new_n3347__, new_new_n3348__,
    new_new_n3349__, new_new_n3350__, new_new_n3351__, new_new_n3352__,
    new_new_n3353__, new_new_n3354__, new_new_n3355__, new_new_n3356__,
    new_new_n3357__, new_new_n3358__, new_new_n3359__, new_new_n3360__,
    new_new_n3361__, new_new_n3362__, new_new_n3363__, new_new_n3364__,
    new_new_n3365__, new_new_n3366__, new_new_n3367__, new_new_n3368__,
    new_new_n3369__, new_new_n3370__, new_new_n3371__, new_new_n3372__,
    new_new_n3373__, new_new_n3374__, new_new_n3375__, new_new_n3376__,
    new_new_n3377__, new_new_n3378__, new_new_n3379__, new_new_n3380__,
    new_new_n3381__, new_new_n3382__, new_new_n3383__, new_new_n3384__,
    new_new_n3385__, new_new_n3386__, new_new_n3387__, new_new_n3388__,
    new_new_n3389__, new_new_n3390__, new_new_n3391__, new_new_n3392__,
    new_new_n3393__, new_new_n3394__, new_new_n3395__, new_new_n3396__,
    new_new_n3397__, new_new_n3398__, new_new_n3399__, new_new_n3400__,
    new_new_n3401__, new_new_n3402__, new_new_n3403__, new_new_n3404__,
    new_new_n3405__, new_new_n3406__, new_new_n3407__, new_new_n3408__,
    new_new_n3409__, new_new_n3410__, new_new_n3411__, new_new_n3412__,
    new_new_n3413__, new_new_n3414__, new_new_n3415__, new_new_n3416__,
    new_new_n3417__, new_new_n3418__, new_new_n3419__, new_new_n3420__,
    new_new_n3421__, new_new_n3422__, new_new_n3423__, new_new_n3424__,
    new_new_n3425__, new_new_n3426__, new_new_n3427__, new_new_n3428__,
    new_new_n3429__, new_new_n3430__, new_new_n3431__, new_new_n3432__,
    new_new_n3433__, new_new_n3434__, new_new_n3435__, new_new_n3436__,
    new_new_n3437__, new_new_n3438__, new_new_n3439__, new_new_n3440__,
    new_new_n3441__, new_new_n3442__, new_new_n3443__, new_new_n3444__,
    new_new_n3445__, new_new_n3446__, new_new_n3447__, new_new_n3448__,
    new_new_n3449__, new_new_n3450__, new_new_n3451__, new_new_n3452__,
    new_new_n3453__, new_new_n3454__, new_new_n3455__, new_new_n3456__,
    new_new_n3457__, new_new_n3458__, new_new_n3459__, new_new_n3460__,
    new_new_n3461__, new_new_n3462__, new_new_n3463__, new_new_n3464__,
    new_new_n3465__, new_new_n3466__, new_new_n3467__, new_new_n3468__,
    new_new_n3469__, new_new_n3470__, new_new_n3471__, new_new_n3472__,
    new_new_n3473__, new_new_n3474__, new_new_n3475__, new_new_n3476__,
    new_new_n3477__, new_new_n3478__, new_new_n3479__, new_new_n3480__,
    new_new_n3481__, new_new_n3482__, new_new_n3483__, new_new_n3484__,
    new_new_n3485__, new_new_n3486__, new_new_n3487__, new_new_n3488__,
    new_new_n3489__, new_new_n3490__, new_new_n3491__, new_new_n3492__,
    new_new_n3493__, new_new_n3494__, new_new_n3495__, new_new_n3496__,
    new_new_n3497__, new_new_n3498__, new_new_n3499__, new_new_n3500__,
    new_new_n3501__, new_new_n3502__, new_new_n3503__, new_new_n3504__,
    new_new_n3505__, new_new_n3506__, new_new_n3507__, new_new_n3508__,
    new_new_n3509__, new_new_n3510__, new_new_n3511__, new_new_n3512__,
    new_new_n3513__, new_new_n3514__, new_new_n3515__, new_new_n3516__,
    new_new_n3517__, new_new_n3518__, new_new_n3519__, new_new_n3520__,
    new_new_n3521__, new_new_n3522__, new_new_n3523__, new_new_n3524__,
    new_new_n3525__, new_new_n3526__, new_new_n3527__, new_new_n3528__,
    new_new_n3529__, new_new_n3530__, new_new_n3531__, new_new_n3532__,
    new_new_n3533__, new_new_n3534__, new_new_n3535__, new_new_n3536__,
    new_new_n3537__, new_new_n3538__, new_new_n3539__, new_new_n3540__,
    new_new_n3541__, new_new_n3542__, new_new_n3543__, new_new_n3544__,
    new_new_n3545__, new_new_n3546__, new_new_n3547__, new_new_n3548__,
    new_new_n3549__, new_new_n3550__, new_new_n3551__, new_new_n3552__,
    new_new_n3553__, new_new_n3554__, new_new_n3555__, new_new_n3556__,
    new_new_n3557__, new_new_n3558__, new_new_n3559__, new_new_n3560__,
    new_new_n3561__, new_new_n3562__, new_new_n3563__, new_new_n3564__,
    new_new_n3565__, new_new_n3566__, new_new_n3567__, new_new_n3568__,
    new_new_n3569__, new_new_n3570__, new_new_n3571__, new_new_n3572__,
    new_new_n3573__, new_new_n3574__, new_new_n3575__, new_new_n3576__,
    new_new_n3577__, new_new_n3578__, new_new_n3579__, new_new_n3580__,
    new_new_n3581__, new_new_n3582__, new_new_n3583__, new_new_n3584__,
    new_new_n3585__, new_new_n3586__, new_new_n3587__, new_new_n3588__,
    new_new_n3589__, new_new_n3590__, new_new_n3591__, new_new_n3592__,
    new_new_n3593__, new_new_n3594__, new_new_n3595__, new_new_n3596__,
    new_new_n3597__, new_new_n3598__, new_new_n3599__, new_new_n3600__,
    new_new_n3601__, new_new_n3602__, new_new_n3603__, new_new_n3604__,
    new_new_n3605__, new_new_n3606__, new_new_n3607__, new_new_n3608__,
    new_new_n3609__, new_new_n3610__, new_new_n3611__, new_new_n3612__,
    new_new_n3613__, new_new_n3614__, new_new_n3615__, new_new_n3616__,
    new_new_n3617__, new_new_n3618__, new_new_n3619__, new_new_n3620__,
    new_new_n3621__, new_new_n3622__, new_new_n3623__, new_new_n3624__,
    new_new_n3625__, new_new_n3626__, new_new_n3627__, new_new_n3628__,
    new_new_n3629__, new_new_n3630__, new_new_n3631__, new_new_n3632__,
    new_new_n3633__, new_new_n3634__, new_new_n3635__, new_new_n3636__,
    new_new_n3637__, new_new_n3638__, new_new_n3639__, new_new_n3640__,
    new_new_n3641__, new_new_n3642__, new_new_n3643__, new_new_n3644__,
    new_new_n3645__, new_new_n3646__, new_new_n3647__, new_new_n3648__,
    new_new_n3649__, new_new_n3650__, new_new_n3651__, new_new_n3652__,
    new_new_n3653__, new_new_n3654__, new_new_n3655__, new_new_n3656__,
    new_new_n3657__, new_new_n3658__, new_new_n3659__, new_new_n3660__,
    new_new_n3661__, new_new_n3662__, new_new_n3663__, new_new_n3664__,
    new_new_n3665__, new_new_n3666__, new_new_n3667__, new_new_n3668__,
    new_new_n3669__, new_new_n3670__, new_new_n3671__, new_new_n3672__,
    new_new_n3673__, new_new_n3674__, new_new_n3675__, new_new_n3676__,
    new_new_n3677__, new_new_n3678__, new_new_n3679__, new_new_n3680__,
    new_new_n3681__, new_new_n3682__, new_new_n3683__, new_new_n3684__,
    new_new_n3685__, new_new_n3686__, new_new_n3687__, new_new_n3688__,
    new_new_n3689__, new_new_n3690__, new_new_n3691__, new_new_n3692__,
    new_new_n3693__, new_new_n3694__, new_new_n3695__, new_new_n3696__,
    new_new_n3697__, new_new_n3698__, new_new_n3699__, new_new_n3700__,
    new_new_n3701__, new_new_n3702__, new_new_n3703__, new_new_n3704__,
    new_new_n3705__, new_new_n3706__, new_new_n3707__, new_new_n3708__,
    new_new_n3709__, new_new_n3710__, new_new_n3711__, new_new_n3712__,
    new_new_n3713__, new_new_n3714__, new_new_n3715__, new_new_n3716__,
    new_new_n3717__, new_new_n3718__, new_new_n3719__, new_new_n3720__,
    new_new_n3721__, new_new_n3722__, new_new_n3723__, new_new_n3724__,
    new_new_n3725__, new_new_n3726__, new_new_n3727__, new_new_n3728__,
    new_new_n3729__, new_new_n3730__, new_new_n3731__, new_new_n3732__,
    new_new_n3733__, new_new_n3734__, new_new_n3735__, new_new_n3736__,
    new_new_n3737__, new_new_n3738__, new_new_n3739__, new_new_n3740__,
    new_new_n3741__, new_new_n3742__, new_new_n3743__, new_new_n3744__,
    new_new_n3745__, new_new_n3746__, new_new_n3747__, new_new_n3748__,
    new_new_n3749__, new_new_n3750__, new_new_n3751__, new_new_n3752__,
    new_new_n3753__, new_new_n3754__, new_new_n3755__, new_new_n3756__,
    new_new_n3757__, new_new_n3758__, new_new_n3759__, new_new_n3760__,
    new_new_n3761__, new_new_n3762__, new_new_n3763__, new_new_n3764__,
    new_new_n3765__, new_new_n3766__, new_new_n3767__, new_new_n3768__,
    new_new_n3769__, new_new_n3770__, new_new_n3771__, new_new_n3772__,
    new_new_n3773__, new_new_n3774__, new_new_n3775__, new_new_n3776__,
    new_new_n3777__, new_new_n3778__, new_new_n3779__, new_new_n3780__,
    new_new_n3781__, new_new_n3782__, new_new_n3783__, new_new_n3784__,
    new_new_n3785__, new_new_n3786__, new_new_n3787__, new_new_n3788__,
    new_new_n3789__, new_new_n3790__, new_new_n3791__, new_new_n3792__,
    new_new_n3793__, new_new_n3794__, new_new_n3795__, new_new_n3796__,
    new_new_n3797__, new_new_n3798__, new_new_n3799__, new_new_n3800__,
    new_new_n3801__, new_new_n3802__, new_new_n3803__, new_new_n3804__,
    new_new_n3805__, new_new_n3806__, new_new_n3807__, new_new_n3808__,
    new_new_n3809__, new_new_n3810__, new_new_n3811__, new_new_n3812__,
    new_new_n3813__, new_new_n3814__, new_new_n3815__, new_new_n3816__,
    new_new_n3817__, new_new_n3818__, new_new_n3819__, new_new_n3820__,
    new_new_n3821__, new_new_n3822__, new_new_n3823__, new_new_n3824__,
    new_new_n3825__, new_new_n3826__, new_new_n3827__, new_new_n3828__,
    new_new_n3829__, new_new_n3830__, new_new_n3831__, new_new_n3832__,
    new_new_n3833__, new_new_n3834__, new_new_n3835__, new_new_n3836__,
    new_new_n3837__, new_new_n3838__, new_new_n3839__, new_new_n3840__,
    new_new_n3841__, new_new_n3842__, new_new_n3843__, new_new_n3844__,
    new_new_n3845__, new_new_n3846__, new_new_n3847__, new_new_n3848__,
    new_new_n3849__, new_new_n3850__, new_new_n3851__, new_new_n3852__,
    new_new_n3853__, new_new_n3854__, new_new_n3855__, new_new_n3856__,
    new_new_n3857__, new_new_n3858__, new_new_n3859__, new_new_n3860__,
    new_new_n3861__, new_new_n3862__, new_new_n3863__, new_new_n3864__,
    new_new_n3865__, new_new_n3866__, new_new_n3867__, new_new_n3868__,
    new_new_n3869__, new_new_n3870__, new_new_n3871__, new_new_n3872__,
    new_new_n3873__, new_new_n3874__, new_new_n3875__, new_new_n3876__,
    new_new_n3877__, new_new_n3878__, new_new_n3879__, new_new_n3880__,
    new_new_n3881__, new_new_n3882__, new_new_n3883__, new_new_n3884__,
    new_new_n3885__, new_new_n3886__, new_new_n3887__, new_new_n3888__,
    new_new_n3889__, new_new_n3890__, new_new_n3891__, new_new_n3892__,
    new_new_n3893__, new_new_n3894__, new_new_n3895__, new_new_n3896__,
    new_new_n3897__, new_new_n3898__, new_new_n3899__, new_new_n3900__,
    new_new_n3901__, new_new_n3902__, new_new_n3903__, new_new_n3904__,
    new_new_n3905__, new_new_n3906__, new_new_n3907__, new_new_n3908__,
    new_new_n3909__, new_new_n3910__, new_new_n3911__, new_new_n3912__,
    new_new_n3913__, new_new_n3914__, new_new_n3915__, new_new_n3916__,
    new_new_n3917__, new_new_n3918__, new_new_n3919__, new_new_n3920__,
    new_new_n3921__, new_new_n3922__, new_new_n3923__, new_new_n3924__,
    new_new_n3925__, new_new_n3926__, new_new_n3927__, new_new_n3928__,
    new_new_n3929__, new_new_n3930__, new_new_n3931__, new_new_n3932__,
    new_new_n3933__, new_new_n3934__, new_new_n3935__, new_new_n3936__,
    new_new_n3937__, new_new_n3938__, new_new_n3939__, new_new_n3940__,
    new_new_n3941__, new_new_n3942__, new_new_n3943__, new_new_n3944__,
    new_new_n3945__, new_new_n3946__, new_new_n3947__, new_new_n3948__,
    new_new_n3949__, new_new_n3950__, new_new_n3951__, new_new_n3952__,
    new_new_n3953__, new_new_n3954__, new_new_n3955__, new_new_n3956__,
    new_new_n3957__, new_new_n3958__, new_new_n3959__, new_new_n3960__,
    new_new_n3961__, new_new_n3962__, new_new_n3963__, new_new_n3964__,
    new_new_n3965__, new_new_n3966__, new_new_n3967__, new_new_n3968__,
    new_new_n3969__, new_new_n3970__, new_new_n3971__, new_new_n3972__,
    new_new_n3973__, new_new_n3974__, new_new_n3975__, new_new_n3976__,
    new_new_n3977__, new_new_n3978__, new_new_n3979__, new_new_n3980__,
    new_new_n3981__, new_new_n3982__, new_new_n3983__, new_new_n3984__,
    new_new_n3985__, new_new_n3986__, new_new_n3987__, new_new_n3988__,
    new_new_n3989__, new_new_n3990__, new_new_n3991__, new_new_n3992__,
    new_new_n3993__, new_new_n3994__, new_new_n3995__, new_new_n3996__,
    new_new_n3997__, new_new_n3998__, new_new_n3999__, new_new_n4000__,
    new_new_n4001__, new_new_n4002__, new_new_n4003__, new_new_n4004__,
    new_new_n4005__, new_new_n4006__, new_new_n4007__, new_new_n4008__,
    new_new_n4009__, new_new_n4010__, new_new_n4011__, new_new_n4012__,
    new_new_n4013__, new_new_n4014__, new_new_n4015__, new_new_n4016__,
    new_new_n4017__, new_new_n4018__, new_new_n4019__, new_new_n4020__,
    new_new_n4021__, new_new_n4022__, new_new_n4023__, new_new_n4024__,
    new_new_n4025__, new_new_n4026__, new_new_n4027__, new_new_n4028__,
    new_new_n4029__, new_new_n4030__, new_new_n4031__, new_new_n4032__,
    new_new_n4033__, new_new_n4034__, new_new_n4035__, new_new_n4036__,
    new_new_n4037__, new_new_n4038__, new_new_n4039__, new_new_n4040__,
    new_new_n4041__, new_new_n4042__, new_new_n4043__, new_new_n4044__,
    new_new_n4045__, new_new_n4046__, new_new_n4047__, new_new_n4048__,
    new_new_n4049__, new_new_n4050__, new_new_n4051__, new_new_n4052__,
    new_new_n4053__, new_new_n4054__, new_new_n4055__, new_new_n4056__,
    new_new_n4057__, new_new_n4058__, new_new_n4059__, new_new_n4060__,
    new_new_n4061__, new_new_n4062__, new_new_n4063__, new_new_n4064__,
    new_new_n4065__, new_new_n4066__, new_new_n4067__, new_new_n4068__,
    new_new_n4069__, new_new_n4070__, new_new_n4071__, new_new_n4072__,
    new_new_n4073__, new_new_n4074__, new_new_n4075__, new_new_n4076__,
    new_new_n4077__, new_new_n4078__, new_new_n4079__, new_new_n4080__,
    new_new_n4081__, new_new_n4082__, new_new_n4083__, new_new_n4084__,
    new_new_n4085__, new_new_n4086__, new_new_n4087__, new_new_n4088__,
    new_new_n4089__, new_new_n4090__, new_new_n4091__, new_new_n4092__,
    new_new_n4093__, new_new_n4094__, new_new_n4095__, new_new_n4096__,
    new_new_n4097__, new_new_n4098__, new_new_n4099__, new_new_n4100__,
    new_new_n4101__, new_new_n4102__, new_new_n4103__, new_new_n4104__,
    new_new_n4105__, new_new_n4106__, new_new_n4107__, new_new_n4108__,
    new_new_n4109__, new_new_n4110__, new_new_n4111__, new_new_n4112__,
    new_new_n4113__, new_new_n4114__, new_new_n4115__, new_new_n4116__,
    new_new_n4117__, new_new_n4118__, new_new_n4119__, new_new_n4120__,
    new_new_n4121__, new_new_n4122__, new_new_n4123__, new_new_n4124__,
    new_new_n4125__, new_new_n4126__, new_new_n4127__, new_new_n4128__,
    new_new_n4129__, new_new_n4130__, new_new_n4131__, new_new_n4132__,
    new_new_n4133__, new_new_n4134__, new_new_n4135__, new_new_n4136__,
    new_new_n4137__, new_new_n4138__, new_new_n4139__, new_new_n4140__,
    new_new_n4141__, new_new_n4142__, new_new_n4143__, new_new_n4144__,
    new_new_n4145__, new_new_n4146__, new_new_n4147__, new_new_n4148__,
    new_new_n4149__, new_new_n4150__, new_new_n4151__, new_new_n4152__,
    new_new_n4153__, new_new_n4154__, new_new_n4155__, new_new_n4156__,
    new_new_n4157__, new_new_n4158__, new_new_n4159__, new_new_n4160__,
    new_new_n4161__, new_new_n4162__, new_new_n4163__, new_new_n4164__,
    new_new_n4165__, new_new_n4166__, new_new_n4167__, new_new_n4168__,
    new_new_n4169__, new_new_n4170__, new_new_n4171__, new_new_n4172__,
    new_new_n4173__, new_new_n4174__, new_new_n4175__, new_new_n4176__,
    new_new_n4177__, new_new_n4178__, new_new_n4179__, new_new_n4180__,
    new_new_n4181__, new_new_n4182__, new_new_n4183__, new_new_n4184__,
    new_new_n4185__, new_new_n4186__, new_new_n4187__, new_new_n4188__,
    new_new_n4189__, new_new_n4190__, new_new_n4191__, new_new_n4192__,
    new_new_n4193__, new_new_n4194__, new_new_n4195__, new_new_n4196__,
    new_new_n4197__, new_new_n4198__, new_new_n4199__, new_new_n4200__,
    new_new_n4201__, new_new_n4202__, new_new_n4203__, new_new_n4204__,
    new_new_n4205__, new_new_n4206__, new_new_n4207__, new_new_n4208__,
    new_new_n4209__, new_new_n4210__, new_new_n4211__, new_new_n4212__,
    new_new_n4213__, new_new_n4214__, new_new_n4215__, new_new_n4216__,
    new_new_n4217__, new_new_n4218__, new_new_n4219__, new_new_n4220__,
    new_new_n4221__, new_new_n4222__, new_new_n4223__, new_new_n4224__,
    new_new_n4225__, new_new_n4226__, new_new_n4227__, new_new_n4228__,
    new_new_n4229__, new_new_n4230__, new_new_n4231__, new_new_n4232__,
    new_new_n4233__, new_new_n4234__, new_new_n4235__, new_new_n4236__,
    new_new_n4237__, new_new_n4238__, new_new_n4239__, new_new_n4240__,
    new_new_n4241__, new_new_n4242__, new_new_n4243__, new_new_n4244__,
    new_new_n4245__, new_new_n4246__, new_new_n4247__, new_new_n4248__,
    new_new_n4249__, new_new_n4250__, new_new_n4251__, new_new_n4252__,
    new_new_n4253__, new_new_n4254__, new_new_n4255__, new_new_n4256__,
    new_new_n4257__, new_new_n4258__, new_new_n4259__, new_new_n4260__,
    new_new_n4261__, new_new_n4262__, new_new_n4263__, new_new_n4264__,
    new_new_n4265__, new_new_n4266__, new_new_n4267__, new_new_n4268__,
    new_new_n4269__, new_new_n4270__, new_new_n4271__, new_new_n4272__,
    new_new_n4273__, new_new_n4274__, new_new_n4275__, new_new_n4276__,
    new_new_n4277__, new_new_n4278__, new_new_n4279__, new_new_n4280__,
    new_new_n4281__, new_new_n4282__, new_new_n4283__, new_new_n4284__,
    new_new_n4285__, new_new_n4286__, new_new_n4287__, new_new_n4288__,
    new_new_n4289__, new_new_n4290__, new_new_n4291__, new_new_n4292__,
    new_new_n4293__, new_new_n4294__, new_new_n4295__, new_new_n4296__,
    new_new_n4297__, new_new_n4298__, new_new_n4299__, new_new_n4300__,
    new_new_n4301__, new_new_n4302__, new_new_n4303__, new_new_n4304__,
    new_new_n4305__, new_new_n5047__, new_new_n5048__, new_new_n5049__,
    new_new_n5050__, new_new_n5051__, new_new_n5052__, new_new_n5053__,
    new_new_n5054__, new_new_n5055__, new_new_n5056__, new_new_n5057__,
    new_new_n5058__, new_new_n5059__, new_new_n5060__, new_new_n5061__,
    new_new_n5062__, new_new_n5063__, new_new_n5064__, new_new_n5065__,
    new_new_n5066__, new_new_n5067__, new_new_n5068__, new_new_n5069__,
    new_new_n5070__, new_new_n5071__, new_new_n5072__, new_new_n5073__,
    new_new_n5074__, new_new_n5075__, new_new_n5076__, new_new_n5077__,
    new_new_n5078__, new_new_n5079__, new_new_n5080__, new_new_n5081__,
    new_new_n5082__, new_new_n5083__, new_new_n5084__, new_new_n5085__,
    new_new_n5086__, new_new_n5087__, new_new_n5088__, new_new_n5089__,
    new_new_n5090__, new_new_n5091__, new_new_n5092__, new_new_n5093__,
    new_new_n5094__, new_new_n5095__, new_new_n5096__, new_new_n5097__,
    new_new_n5098__, new_new_n5099__, new_new_n5100__, new_new_n5101__,
    new_new_n5102__, new_new_n5103__, new_new_n5104__, new_new_n5105__,
    new_new_n5106__, new_new_n5107__, new_new_n5108__, new_new_n5109__,
    new_new_n5110__, new_new_n5111__, new_new_n5112__, new_new_n5113__,
    new_new_n5114__, new_new_n5115__, new_new_n5116__, new_new_n5117__,
    new_new_n5118__, new_new_n5119__, new_new_n5120__, new_new_n5121__,
    new_new_n5122__, new_new_n5123__, new_new_n5124__, new_new_n5125__,
    new_new_n5126__, new_new_n5127__, new_new_n5128__, new_new_n5129__,
    new_new_n5130__, new_new_n5131__, new_new_n5132__, new_new_n5133__,
    new_new_n5134__, new_new_n5135__, new_new_n5136__, new_new_n5137__,
    new_new_n5138__, new_new_n5139__, new_new_n5140__, new_new_n5141__,
    new_new_n5142__, new_new_n5143__, new_new_n5144__, new_new_n5145__,
    new_new_n5146__, new_new_n5147__, new_new_n5148__, new_new_n5149__,
    new_new_n5150__, new_new_n5151__, new_new_n5152__, new_new_n5153__,
    new_new_n5154__, new_new_n5155__, new_new_n5156__, new_new_n5157__,
    new_new_n5158__, new_new_n5159__, new_new_n5160__, new_new_n5161__,
    new_new_n5162__, new_new_n5163__, new_new_n5164__, new_new_n5165__,
    new_new_n5166__, new_new_n5167__, new_new_n5168__, new_new_n5169__,
    new_new_n5170__, new_new_n5171__, new_new_n5172__, new_new_n5173__,
    new_new_n5174__, new_new_n5175__, new_new_n5176__, new_new_n5177__,
    new_new_n5178__, new_new_n5179__, new_new_n5180__, new_new_n5181__,
    new_new_n5182__, new_new_n5183__, new_new_n5184__, new_new_n5185__,
    new_new_n5186__, new_new_n5187__, new_new_n5188__, new_new_n5189__,
    new_new_n5190__, new_new_n5191__, new_new_n5192__, new_new_n5193__,
    new_new_n5194__, new_new_n5195__, new_new_n5196__, new_new_n5197__,
    new_new_n5198__, new_new_n5199__, new_new_n5200__, new_new_n5201__,
    new_new_n5202__, new_new_n5203__, new_new_n5204__, new_new_n5205__,
    new_new_n5206__, new_new_n5207__, new_new_n5208__, new_new_n5209__,
    new_new_n5210__, new_new_n5211__, new_new_n5212__, new_new_n5213__,
    new_new_n5214__, new_new_n5215__, new_new_n5216__, new_new_n5217__,
    new_new_n5218__, new_new_n5219__, new_new_n5220__, new_new_n5221__,
    new_new_n5222__, new_new_n5223__, new_new_n5224__, new_new_n5225__,
    new_new_n5226__, new_new_n5227__, new_new_n5228__, new_new_n5229__,
    new_new_n5230__, new_new_n5231__, new_new_n5232__, new_new_n5233__,
    new_new_n5234__, new_new_n5235__, new_new_n5236__, new_new_n5237__,
    new_new_n5238__, new_new_n5239__, new_new_n5240__, new_new_n5241__,
    new_new_n5242__, new_new_n5243__, new_new_n5244__, new_new_n5245__,
    new_new_n5246__, new_new_n5247__, new_new_n5248__, new_new_n5249__,
    new_new_n5250__, new_new_n5251__, new_new_n5252__, new_new_n5253__,
    new_new_n5254__, new_new_n5255__, new_new_n5256__, new_new_n5257__,
    new_new_n5258__, new_new_n5259__, new_new_n5260__, new_new_n5261__,
    new_new_n5262__, new_new_n5263__, new_new_n5264__, new_new_n5265__,
    new_new_n5266__, new_new_n5267__, new_new_n5268__, new_new_n5269__,
    new_new_n5270__, new_new_n5271__, new_new_n5272__, new_new_n5273__,
    new_new_n5274__, new_new_n5275__, new_new_n5276__, new_new_n5277__,
    new_new_n5278__, new_new_n5279__, new_new_n5280__, new_new_n5281__,
    new_new_n5282__, new_new_n5283__, new_new_n5284__, new_new_n5285__,
    new_new_n5286__, new_new_n5287__, new_new_n5288__, new_new_n5289__,
    new_new_n5290__, new_new_n5291__, new_new_n5292__, new_new_n5293__,
    new_new_n5294__, new_new_n5295__, new_new_n5296__, new_new_n5297__,
    new_new_n5298__, new_new_n5299__, new_new_n5300__, new_new_n5301__,
    new_new_n5302__, new_new_n5303__, new_new_n5304__, new_new_n5305__,
    new_new_n5306__, new_new_n5307__, new_new_n5308__, new_new_n5309__,
    new_new_n5310__, new_new_n5311__, new_new_n5312__, new_new_n5313__,
    new_new_n5314__, new_new_n5315__, new_new_n5316__, new_new_n5317__,
    new_new_n5318__, new_new_n5319__, new_new_n5320__, new_new_n5321__,
    new_new_n5322__, new_new_n5323__, new_new_n5324__, new_new_n5325__,
    new_new_n5326__, new_new_n5327__, new_new_n5328__, new_new_n5329__,
    new_new_n5330__, new_new_n5331__, new_new_n5332__, new_new_n5333__,
    new_new_n5334__, new_new_n5335__, new_new_n5336__, new_new_n5337__,
    new_new_n5338__, new_new_n5339__, new_new_n5340__, new_new_n5341__,
    new_new_n5342__, new_new_n5343__, new_new_n5344__, new_new_n5345__,
    new_new_n5346__, new_new_n5347__, new_new_n5348__, new_new_n5349__,
    new_new_n5350__, new_new_n5351__, new_new_n5352__, new_new_n5353__,
    new_new_n5354__, new_new_n5355__, new_new_n5356__, new_new_n5357__,
    new_new_n5358__, new_new_n5359__, new_new_n5360__, new_new_n5361__,
    new_new_n5362__, new_new_n5363__, new_new_n5364__, new_new_n5365__,
    new_new_n5366__, new_new_n5367__, new_new_n5368__, new_new_n5369__,
    new_new_n5370__, new_new_n5371__, new_new_n5372__, new_new_n5373__,
    new_new_n5374__, new_new_n5375__, new_new_n5376__, new_new_n5377__,
    new_new_n5378__, new_new_n5379__, new_new_n5380__, new_new_n5381__,
    new_new_n5382__, new_new_n5383__, new_new_n5384__, new_new_n5385__,
    new_new_n5386__, new_new_n5387__, new_new_n5388__, new_new_n5389__,
    new_new_n5390__, new_new_n5391__, new_new_n5392__, new_new_n5393__,
    new_new_n5394__, new_new_n5395__, new_new_n5396__, new_new_n5397__,
    new_new_n5398__, new_new_n5399__, new_new_n5400__, new_new_n5401__,
    new_new_n5402__, new_new_n5403__, new_new_n5404__, new_new_n5405__,
    new_new_n5406__, new_new_n5407__, new_new_n5408__, new_new_n5409__,
    new_new_n5410__, new_new_n5411__, new_new_n5412__, new_new_n5413__,
    new_new_n5414__, new_new_n5415__, new_new_n5416__, new_new_n5417__,
    new_new_n5418__, new_new_n5419__, new_new_n5420__, new_new_n5421__,
    new_new_n5422__, new_new_n5423__, new_new_n5424__, new_new_n5425__,
    new_new_n5426__, new_new_n5427__, new_new_n5428__, new_new_n5429__,
    new_new_n5430__, new_new_n5431__, new_new_n5432__, new_new_n5433__,
    new_new_n5434__, new_new_n5435__, new_new_n5436__, new_new_n5437__,
    new_new_n5438__, new_new_n5439__, new_new_n5440__, new_new_n5441__,
    new_new_n5442__, new_new_n5443__, new_new_n5444__, new_new_n5445__,
    new_new_n5446__, new_new_n5447__, new_new_n5448__, new_new_n5449__,
    new_new_n5450__, new_new_n5451__, new_new_n5452__, new_new_n5453__,
    new_new_n5454__, new_new_n5455__, new_new_n5456__, new_new_n5457__,
    new_new_n5458__, new_new_n5459__, new_new_n5460__, new_new_n5461__,
    new_new_n5462__, new_new_n5463__, new_new_n5464__, new_new_n5465__,
    new_new_n5466__, new_new_n5467__, new_new_n5468__, new_new_n5469__,
    new_new_n5470__, new_new_n5471__, new_new_n5472__, new_new_n5473__,
    new_new_n5474__, new_new_n5475__, new_new_n5476__, new_new_n5477__,
    new_new_n5478__, new_new_n5479__, new_new_n5480__, new_new_n5481__,
    new_new_n5482__, new_new_n5483__, new_new_n5484__, new_new_n5485__,
    new_new_n5486__, new_new_n5487__, new_new_n5488__, new_new_n5489__,
    new_new_n5490__, new_new_n5491__, new_new_n5492__, new_new_n5493__,
    new_new_n5494__, new_new_n5495__, new_new_n5496__, new_new_n5497__,
    new_new_n5498__, new_new_n5499__, new_new_n5500__, new_new_n5501__,
    new_new_n5502__, new_new_n5503__, new_new_n5504__, new_new_n5505__,
    new_new_n5506__, new_new_n5507__, new_new_n5508__, new_new_n5509__,
    new_new_n5510__, new_new_n5511__, new_new_n5512__, new_new_n5513__,
    new_new_n5514__, new_new_n5515__, new_new_n5516__, new_new_n5517__,
    new_new_n5518__, new_new_n5519__, new_new_n5520__, new_new_n5521__,
    new_new_n5522__, new_new_n5523__, new_new_n5524__, new_new_n5525__,
    new_new_n5526__, new_new_n5527__, new_new_n5528__, new_new_n5529__,
    new_new_n5530__, new_new_n5531__, new_new_n5532__, new_new_n5533__,
    new_new_n5534__, new_new_n5535__, new_new_n5536__, new_new_n5537__,
    new_new_n5538__, new_new_n5539__, new_new_n5540__, new_new_n5541__,
    new_new_n5542__, new_new_n5543__, new_new_n5544__, new_new_n5545__,
    new_new_n5546__, new_new_n5547__, new_new_n5548__, new_new_n5549__,
    new_new_n5550__, new_new_n5551__, new_new_n5552__, new_new_n5553__,
    new_new_n5554__, new_new_n5555__, new_new_n5556__, new_new_n5557__,
    new_new_n5558__, new_new_n5559__, new_new_n5560__, new_new_n5561__,
    new_new_n5562__, new_new_n5563__, new_new_n5564__, new_new_n5565__,
    new_new_n5566__, new_new_n5567__, new_new_n5568__, new_new_n5569__,
    new_new_n5570__, new_new_n5571__, new_new_n5572__, new_new_n5573__,
    new_new_n5574__, new_new_n5575__, new_new_n5576__, new_new_n5577__,
    new_new_n5578__, new_new_n5579__, new_new_n5580__, new_new_n5581__,
    new_new_n5582__, new_new_n5583__, new_new_n5584__, new_new_n5585__,
    new_new_n5586__, new_new_n5587__, new_new_n5588__, new_new_n5589__,
    new_new_n5590__, new_new_n5591__, new_new_n5592__, new_new_n5593__,
    new_new_n5594__, new_new_n5595__, new_new_n5596__, new_new_n5597__,
    new_new_n5598__, new_new_n5599__, new_new_n5600__, new_new_n5601__,
    new_new_n5602__, new_new_n5603__, new_new_n5604__, new_new_n5605__,
    new_new_n5606__, new_new_n5607__, new_new_n5608__, new_new_n5609__,
    new_new_n5610__, new_new_n5611__, new_new_n5612__, new_new_n5613__,
    new_new_n5614__, new_new_n5615__, new_new_n5616__, new_new_n5617__,
    new_new_n5618__, new_new_n5619__, new_new_n5620__, new_new_n5621__,
    new_new_n5622__, new_new_n5623__, new_new_n5624__, new_new_n5625__,
    new_new_n5626__, new_new_n5627__, new_new_n5628__, new_new_n5629__,
    new_new_n5630__, new_new_n5631__, new_new_n5632__, new_new_n5633__,
    new_new_n5634__, new_new_n5635__, new_new_n5636__, new_new_n5637__,
    new_new_n5638__, new_new_n5639__, new_new_n5640__, new_new_n5641__,
    new_new_n5642__, new_new_n5643__, new_new_n5644__, new_new_n5645__,
    new_new_n5646__, new_new_n5647__, new_new_n5648__, new_new_n5649__,
    new_new_n5650__, new_new_n5651__, new_new_n5652__, new_new_n5653__,
    new_new_n5654__, new_new_n5655__, new_new_n5656__, new_new_n5657__,
    new_new_n5658__, new_new_n5659__, new_new_n5660__, new_new_n5661__,
    new_new_n5662__, new_new_n5663__, new_new_n5664__, new_new_n5665__,
    new_new_n5666__, new_new_n5667__, new_new_n5668__, new_new_n5669__,
    new_new_n5670__, new_new_n5671__, new_new_n5672__, new_new_n5673__,
    new_new_n5674__, new_new_n5675__, new_new_n5676__, new_new_n5677__,
    new_new_n5678__, new_new_n5679__, new_new_n5680__, new_new_n5681__,
    new_new_n5682__, new_new_n5683__, new_new_n5684__, new_new_n5685__,
    new_new_n5686__, new_new_n5687__, new_new_n5688__, new_new_n5689__,
    new_new_n5690__, new_new_n5691__, new_new_n5692__, new_new_n5693__,
    new_new_n5694__, new_new_n5695__, new_new_n5696__, new_new_n5697__,
    new_new_n5698__, new_new_n5699__, new_new_n5700__, new_new_n5701__,
    new_new_n5702__, new_new_n5703__, new_new_n5704__, new_new_n5705__,
    new_new_n5706__, new_new_n5707__, new_new_n5708__, new_new_n5709__,
    new_new_n5710__, new_new_n5711__, new_new_n5712__, new_new_n5713__,
    new_new_n5714__, new_new_n5715__, new_new_n5716__, new_new_n5717__,
    new_new_n5718__, new_new_n5719__, new_new_n5720__, new_new_n5721__,
    new_new_n5722__, new_new_n5723__, new_new_n5724__, new_new_n5725__,
    new_new_n5726__, new_new_n5727__, new_new_n5728__, new_new_n5729__,
    new_new_n5730__, new_new_n5731__, new_new_n5732__, new_new_n5733__,
    new_new_n5734__, new_new_n5735__, new_new_n5736__, new_new_n5737__,
    new_new_n5738__, new_new_n5739__, new_new_n5740__, new_new_n5741__,
    new_new_n5742__, new_new_n5743__, new_new_n5744__, new_new_n5745__,
    new_new_n5746__, new_new_n5747__, new_new_n5748__, new_new_n5749__,
    new_new_n5750__, new_new_n5751__, new_new_n5752__, new_new_n5753__,
    new_new_n5754__, new_new_n5755__, new_new_n5756__, new_new_n5757__,
    new_new_n5758__, new_new_n5759__, new_new_n5760__, new_new_n5761__,
    new_new_n5762__, new_new_n5763__, new_new_n5764__, new_new_n5765__,
    new_new_n5766__, new_new_n5767__, new_new_n5768__, new_new_n5769__,
    new_new_n5770__, new_new_n5771__, new_new_n5772__, new_new_n5773__,
    new_new_n5774__, new_new_n5775__, new_new_n5776__, new_new_n5777__,
    new_new_n5778__, new_new_n5779__, new_new_n5780__, new_new_n5781__,
    new_new_n5782__, new_new_n5783__, new_new_n5784__, new_new_n5785__,
    new_new_n5786__, new_new_n5787__, new_new_n5788__, new_new_n5789__,
    new_new_n5790__, n8268, n8271, n8274, n8277, n8280, n8283, n8286,
    n8289, n8292, n8295, n8298, n8301, n8304, n8307, n8310, n8313, n8316,
    n8319, n8322, n8325, n8328, n8331, n8334, n8337, n8340, n8343, n8346,
    n8349, n8352, n8355, n8358, n8361, n8364, n8367, n8370, n8373, n8376,
    n8379, n8382, n8385, n8388, n8391, n8394, n8397, n8400, n8403, n8406,
    n8409, n8412, n8415, n8418, n8421, n8424, n8427, n8430, n8433, n8436,
    n8439, n8442, n8445, n8448, n8451, n8454, n8457, n8460, n8463, n8466,
    n8469, n8472, n8475, n8478, n8481, n8484, n8487, n8490, n8493, n8496,
    n8499, n8502, n8505, n8508, n8511, n8514, n8517, n8520, n8523, n8526,
    n8529, n8532, n8535, n8538, n8541, n8544, n8547, n8550, n8553, n8556,
    n8559, n8562, n8565, n8568, n8571, n8574, n8577, n8580, n8583, n8586,
    n8589, n8592, n8595, n8598, n8601, n8604, n8607, n8610, n8613, n8616,
    n8619, n8622, n8625, n8628, n8631, n8634, n8637, n8640, n8643, n8646,
    n8649, n8652, n8655, n8658, n8661, n8664, n8667, n8670, n8673, n8676,
    n8679, n8682, n8685, n8688, n8691, n8694, n8697, n8700, n8703, n8706,
    n8709, n8712, n8715, n8718, n8721, n8724, n8727, n8730, n8733, n8736,
    n8739, n8742, n8745, n8748, n8751, n8754, n8757, n8760, n8763, n8766,
    n8769, n8772, n8775, n8778, n8781, n8784, n8787, n8790, n8793, n8796,
    n8799, n8802, n8805, n8808, n8811, n8814, n8817, n8820, n8823, n8826,
    n8829, n8832, n8835, n8838, n8841, n8844, n8847, n8850, n8853, n8856,
    n8859, n8862, n8865, n8868, n8871, n8874, n8877, n8880, n8883, n8886,
    n8889, n8892, n8895, n8898, n8901, n8904, n8907, n8910, n8913, n8916,
    n8919, n8922, n8925, n8928, n8931, n8934, n8937, n8940, n8943, n8946,
    n8949, n8952, n8955, n8958, n8961, n8964, n8967, n8970, n8973, n8976,
    n8979, n8982, n8985, n8988, n8991, n8994, n8997, n9000, n9003, n9006,
    n9009, n9012, n9015, n9018, n9021, n9024, n9027, n9030, n9033, n9036,
    n9039, n9042, n9045, n9048, n9051, n9054, n9057, n9060, n9063, n9066,
    n9069, n9072, n9075, n9078, n9081, n9084, n9087, n9090, n9093, n9096,
    n9099, n9102, n9105, n9108, n9111, n9114, n9117, n9120, n9123, n9126,
    n9129, n9132, n9135, n9138, n9141, n9144, n9147, n9150, n9153, n9156,
    n9159, n9162, n9165, n9168, n9171, n9174, n9177, n9180, n9183, n9186,
    n9189, n9192, n9195, n9198, n9201, n9204, n9207, n9210, n9213, n9216,
    n9219, n9222, n9225, n9228, n9231, n9234, n9237, n9240, n9243, n9246,
    n9249, n9252, n9255, n9258, n9261, n9264, n9267, n9270, n9273, n9276,
    n9279, n9282, n9285, n9288, n9291, n9294, n9297, n9300, n9303, n9306,
    n9309, n9312, n9315, n9318, n9321, n9324, n9327, n9330, n9333, n9336,
    n9339, n9342, n9345, n9348, n9351, n9354, n9357, n9360, n9363, n9366,
    n9369, n9372, n9375, n9378, n9381, n9384, n9387, n9390, n9393, n9396,
    n9399, n9402, n9405, n9408, n9411, n9414, n9417, n9420, n9423, n9426,
    n9429, n9432, n9435, n9438, n9441, n9444, n9447, n9450, n9453, n9456,
    n9459, n9462, n9465, n9468, n9471, n9474, n9477, n9480, n9483, n9486,
    n9489, n9492, n9495, n9498, n9501, n9504, n9507, n9510, n9513, n9516,
    n9519, n9522, n9525, n9528, n9531, n9534, n9537, n9540, n9543, n9546,
    n9549, n9552, n9555, n9558, n9561, n9564, n9567, n9570, n9573, n9576,
    n9579, n9582, n9585, n9588, n9591, n9594, n9597, n9600, n9603, n9606,
    n9609, n9612, n9615, n9618, n9621, n9624, n9627, n9630, n9633, n9636,
    n9639, n9642, n9645, n9648, n9651, n9654, n9657, n9660, n9663, n9666,
    n9669, n9672, n9675, n9678, n9681, n9684, n9687, n9690, n9693, n9696,
    n9699, n9702, n9705, n9708, n9711, n9714, n9717, n9720, n9723, n9726,
    n9729, n9732, n9735, n9738, n9741, n9744, n9747, n9750, n9753, n9756,
    n9759, n9762, n9765, n9768, n9771, n9774, n9777, n9780, n9783, n9786,
    n9789, n9792, n9795, n9798, n9801, n9804, n9807, n9810, n9813, n9816,
    n9819, n9822, n9825, n9828, n9831, n9834, n9837, n9840, n9843, n9846,
    n9849, n9852, n9855, n9858, n9861, n9864, n9867, n9870, n9873, n9876,
    n9879, n9882, n9885, n9888, n9891, n9894, n9897, n9900, n9903, n9906,
    n9909, n9912, n9915, n9918, n9921, n9924, n9927, n9930, n9933, n9936,
    n9939, n9942, n9945, n9948, n9951, n9954, n9957, n9960, n9963, n9966,
    n9969, n9972, n9975, n9978, n9981, n9984, n9987, n9990, n9993, n9996,
    n9999, n10002, n10005, n10008, n10011, n10014, n10017, n10020, n10023,
    n10026, n10029, n10032, n10035, n10038, n10041, n10044, n10047, n10050,
    n10053, n10056, n10059, n10062, n10065, n10068, n10071, n10074, n10077,
    n10080, n10083, n10086, n10089, n10092, n10095, n10098, n10101, n10104,
    n10107, n10110, n10113, n10116, n10119, n10122, n10125, n10128, n10131,
    n10134, n10137, n10140, n10143, n10146, n10149, n10152, n10155, n10158,
    n10161, n10164, n10167, n10170, n10173, n10176, n10179, n10182, n10185,
    n10188, n10191, n10194, n10197, n10200, n10203, n10206, n10209, n10212,
    n10215, n10218, n10221, n10224, n10227, n10230, n10233, n10236, n10239,
    n10242, n10245, n10248, n10251, n10254, n10257, n10260, n10263, n10266,
    n10269, n10272, n10275, n10278, n10281, n10284, n10287, n10290, n10293,
    n10296;
  buf1  g0000(.din(G1), .dout(new_new_n1576__));
  buf1  g0001(.din(G2), .dout(new_new_n1578__));
  buf1  g0002(.din(G3), .dout(new_new_n1580__));
  buf1  g0003(.din(G4), .dout(new_new_n1582__));
  buf1  g0004(.din(G5), .dout(new_new_n1584__));
  buf1  g0005(.din(G6), .dout(new_new_n1586__));
  buf1  g0006(.din(G7), .dout(new_new_n1588__));
  buf1  g0007(.din(G8), .dout(new_new_n1590__));
  buf1  g0008(.din(G9), .dout(new_new_n1592__));
  buf1  g0009(.din(G10), .dout(new_new_n1594__));
  buf1  g0010(.din(G11), .dout(new_new_n1596__));
  buf1  g0011(.din(G12), .dout(new_new_n1598__));
  buf1  g0012(.din(G13), .dout(new_new_n1600__));
  buf1  g0013(.din(G14), .dout(new_new_n1602__));
  buf1  g0014(.din(G15), .dout(new_new_n1604__));
  buf1  g0015(.din(G16), .dout(new_new_n1606__));
  buf1  g0016(.din(G17), .dout(new_new_n1608__));
  buf1  g0017(.din(G18), .dout(new_new_n1610__));
  buf1  g0018(.din(G19), .dout(new_new_n1612__));
  buf1  g0019(.din(G20), .dout(new_new_n1614__));
  buf1  g0020(.din(G21), .dout(new_new_n1616__));
  buf1  g0021(.din(G22), .dout(new_new_n1618__));
  buf1  g0022(.din(G23), .dout(new_new_n1620__));
  buf1  g0023(.din(G24), .dout(new_new_n1622__));
  buf1  g0024(.din(G25), .dout(new_new_n1624__));
  buf1  g0025(.din(G26), .dout(new_new_n1626__));
  buf1  g0026(.din(G27), .dout(new_new_n1628__));
  buf1  g0027(.din(G28), .dout(new_new_n1630__));
  buf1  g0028(.din(G29), .dout(new_new_n1632__));
  buf1  g0029(.din(G30), .dout(new_new_n1634__));
  buf1  g0030(.din(G31), .dout(new_new_n1636__));
  buf1  g0031(.din(G32), .dout(new_new_n1638__));
  buf1  g0032(.din(G33), .dout(new_new_n1640__));
  buf1  g0033(.din(G34), .dout(new_new_n1642__));
  buf1  g0034(.din(G35), .dout(new_new_n1644__));
  buf1  g0035(.din(G36), .dout(new_new_n1646__));
  buf1  g0036(.din(G37), .dout(new_new_n1648__));
  buf1  g0037(.din(G38), .dout(new_new_n1650__));
  buf1  g0038(.din(G39), .dout(new_new_n1652__));
  buf1  g0039(.din(G40), .dout(new_new_n1654__));
  buf1  g0040(.din(G41), .dout(new_new_n1656__));
  buf1  g0041(.din(G42), .dout(new_new_n1658__));
  buf1  g0042(.din(G43), .dout(new_new_n1660__));
  buf1  g0043(.din(G44), .dout(new_new_n1662__));
  buf1  g0044(.din(G45), .dout(new_new_n1664__));
  buf1  g0045(.din(G46), .dout(new_new_n1666__));
  buf1  g0046(.din(G47), .dout(new_new_n1668__));
  buf1  g0047(.din(G48), .dout(new_new_n1670__));
  buf1  g0048(.din(G49), .dout(new_new_n1672__));
  buf1  g0049(.din(G50), .dout(new_new_n1674__));
  buf1  g0050(.din(G51), .dout(new_new_n1676__));
  buf1  g0051(.din(G52), .dout(new_new_n1678__));
  buf1  g0052(.din(G53), .dout(new_new_n1680__));
  buf1  g0053(.din(G54), .dout(new_new_n1682__));
  buf1  g0054(.din(G55), .dout(new_new_n1684__));
  buf1  g0055(.din(G56), .dout(new_new_n1686__));
  buf1  g0056(.din(G57), .dout(new_new_n1688__));
  buf1  g0057(.din(G58), .dout(new_new_n1690__));
  buf1  g0058(.din(G59), .dout(new_new_n1692__));
  buf1  g0059(.din(G60), .dout(new_new_n1694__));
  buf1  g0060(.din(G61), .dout(new_new_n1696__));
  buf1  g0061(.din(G62), .dout(new_new_n1698__));
  buf1  g0062(.din(G63), .dout(new_new_n1700__));
  buf1  g0063(.din(G64), .dout(new_new_n1702__));
  buf1  g0064(.din(G65), .dout(new_new_n1704__));
  buf1  g0065(.din(G66), .dout(new_new_n1706__));
  buf1  g0066(.din(G67), .dout(new_new_n1708__));
  buf1  g0067(.din(G68), .dout(new_new_n1710__));
  buf1  g0068(.din(G69), .dout(new_new_n1712__));
  buf1  g0069(.din(G70), .dout(new_new_n1714__));
  buf1  g0070(.din(G71), .dout(new_new_n1716__));
  buf1  g0071(.din(G72), .dout(new_new_n1718__));
  buf1  g0072(.din(G73), .dout(new_new_n1720__));
  buf1  g0073(.din(G74), .dout(new_new_n1722__));
  buf1  g0074(.din(G75), .dout(new_new_n1724__));
  buf1  g0075(.din(G76), .dout(new_new_n1726__));
  buf1  g0076(.din(G77), .dout(new_new_n1728__));
  buf1  g0077(.din(G78), .dout(new_new_n1730__));
  buf1  g0078(.din(G79), .dout(new_new_n1732__));
  buf1  g0079(.din(G80), .dout(new_new_n1734__));
  buf1  g0080(.din(G81), .dout(new_new_n1736__));
  buf1  g0081(.din(G82), .dout(new_new_n1738__));
  buf1  g0082(.din(G83), .dout(new_new_n1740__));
  buf1  g0083(.din(G84), .dout(new_new_n1742__));
  buf1  g0084(.din(G85), .dout(new_new_n1744__));
  buf1  g0085(.din(G86), .dout(new_new_n1746__));
  buf1  g0086(.din(G87), .dout(new_new_n1748__));
  buf1  g0087(.din(G88), .dout(new_new_n1750__));
  buf1  g0088(.din(G89), .dout(new_new_n1752__));
  buf1  g0089(.din(G90), .dout(new_new_n1754__));
  buf1  g0090(.din(G91), .dout(new_new_n1756__));
  buf1  g0091(.din(G92), .dout(new_new_n1758__));
  buf1  g0092(.din(G93), .dout(new_new_n1760__));
  buf1  g0093(.din(G94), .dout(new_new_n1762__));
  buf1  g0094(.din(G95), .dout(new_new_n1764__));
  buf1  g0095(.din(G96), .dout(new_new_n1766__));
  buf1  g0096(.din(G97), .dout(new_new_n1768__));
  buf1  g0097(.din(G98), .dout(new_new_n1770__));
  buf1  g0098(.din(G99), .dout(new_new_n1772__));
  buf1  g0099(.din(G100), .dout(new_new_n1774__));
  buf1  g0100(.din(G101), .dout(new_new_n1776__));
  buf1  g0101(.din(G102), .dout(new_new_n1778__));
  buf1  g0102(.din(G103), .dout(new_new_n1780__));
  buf1  g0103(.din(G104), .dout(new_new_n1782__));
  buf1  g0104(.din(G105), .dout(new_new_n1784__));
  buf1  g0105(.din(G106), .dout(new_new_n1786__));
  buf1  g0106(.din(G107), .dout(new_new_n1788__));
  buf1  g0107(.din(G108), .dout(new_new_n1790__));
  buf1  g0108(.din(G109), .dout(new_new_n1792__));
  buf1  g0109(.din(G110), .dout(new_new_n1794__));
  buf1  g0110(.din(G111), .dout(new_new_n1796__));
  buf1  g0111(.din(G112), .dout(new_new_n1798__));
  buf1  g0112(.din(G113), .dout(new_new_n1800__));
  buf1  g0113(.din(G114), .dout(new_new_n1802__));
  buf1  g0114(.din(G115), .dout(new_new_n1804__));
  buf1  g0115(.din(G116), .dout(new_new_n1806__));
  buf1  g0116(.din(G117), .dout(new_new_n1808__));
  buf1  g0117(.din(G118), .dout(new_new_n1810__));
  buf1  g0118(.din(G119), .dout(new_new_n1812__));
  buf1  g0119(.din(G120), .dout(new_new_n1814__));
  buf1  g0120(.din(G121), .dout(new_new_n1816__));
  buf1  g0121(.din(G122), .dout(new_new_n1818__));
  buf1  g0122(.din(G123), .dout(new_new_n1820__));
  buf1  g0123(.din(G124), .dout(new_new_n1822__));
  buf1  g0124(.din(G125), .dout(new_new_n1824__));
  buf1  g0125(.din(G126), .dout(new_new_n1826__));
  buf1  g0126(.din(G127), .dout(new_new_n1828__));
  buf1  g0127(.din(G128), .dout(new_new_n1830__));
  buf1  g0128(.din(G129), .dout(new_new_n1832__));
  buf1  g0129(.din(G130), .dout(new_new_n1834__));
  buf1  g0130(.din(G131), .dout(new_new_n1836__));
  buf1  g0131(.din(G132), .dout(new_new_n1838__));
  buf1  g0132(.din(G133), .dout(new_new_n1840__));
  buf1  g0133(.din(G134), .dout(new_new_n1842__));
  buf1  g0134(.din(G135), .dout(new_new_n1844__));
  buf1  g0135(.din(G136), .dout(new_new_n1846__));
  buf1  g0136(.din(G137), .dout(new_new_n1848__));
  buf1  g0137(.din(G138), .dout(new_new_n1850__));
  buf1  g0138(.din(G139), .dout(new_new_n1852__));
  buf1  g0139(.din(G140), .dout(new_new_n1854__));
  buf1  g0140(.din(G141), .dout(new_new_n1856__));
  buf1  g0141(.din(G142), .dout(new_new_n1858__));
  buf1  g0142(.din(G143), .dout(new_new_n1860__));
  buf1  g0143(.din(G144), .dout(new_new_n1862__));
  buf1  g0144(.din(G145), .dout(new_new_n1864__));
  buf1  g0145(.din(G146), .dout(new_new_n1866__));
  buf1  g0146(.din(G147), .dout(new_new_n1868__));
  buf1  g0147(.din(G148), .dout(new_new_n1870__));
  buf1  g0148(.din(G149), .dout(new_new_n1872__));
  buf1  g0149(.din(G150), .dout(new_new_n1874__));
  buf1  g0150(.din(G151), .dout(new_new_n1876__));
  buf1  g0151(.din(G152), .dout(new_new_n1878__));
  buf1  g0152(.din(G153), .dout(new_new_n1880__));
  buf1  g0153(.din(G154), .dout(new_new_n1882__));
  buf1  g0154(.din(G155), .dout(new_new_n1884__));
  buf1  g0155(.din(G156), .dout(new_new_n1886__));
  buf1  g0156(.din(G157), .dout(new_new_n1888__));
  buf1  g0157(.din(n1416_lo), .dout(new_new_n1890__));
  buf1  g0158(.din(n1419_lo), .dout(new_new_n1892__));
  buf1  g0159(.din(n1422_lo), .dout(new_new_n1894__));
  buf1  g0160(.din(n1425_lo), .dout(new_new_n1896__));
  buf1  g0161(.din(n1428_lo), .dout(new_new_n1898__));
  buf1  g0162(.din(n1431_lo), .dout(new_new_n1900__));
  buf1  g0163(.din(n1434_lo), .dout(new_new_n1902__));
  not1  g0164(.din(n1437_lo), .dout(new_new_n1905__));
  buf1  g0165(.din(n1440_lo), .dout(new_new_n1906__));
  buf1  g0166(.din(n1443_lo), .dout(new_new_n1908__));
  buf1  g0167(.din(n1446_lo), .dout(new_new_n1910__));
  buf1  g0168(.din(n1449_lo), .dout(new_new_n1912__));
  buf1  g0169(.din(n1452_lo), .dout(new_new_n1914__));
  buf1  g0170(.din(n1455_lo), .dout(new_new_n1916__));
  buf1  g0171(.din(n1458_lo), .dout(new_new_n1918__));
  buf1  g0172(.din(n1464_lo), .dout(new_new_n1920__));
  buf1  g0173(.din(n1467_lo), .dout(new_new_n1922__));
  buf1  g0174(.din(n1470_lo), .dout(new_new_n1924__));
  buf1  g0175(.din(n1476_lo), .dout(new_new_n1926__));
  buf1  g0176(.din(n1479_lo), .dout(new_new_n1928__));
  buf1  g0177(.din(n1482_lo), .dout(new_new_n1930__));
  buf1  g0178(.din(n1488_lo), .dout(new_new_n1932__));
  buf1  g0179(.din(n1491_lo), .dout(new_new_n1934__));
  buf1  g0180(.din(n1494_lo), .dout(new_new_n1936__));
  not1  g0181(.din(n1497_lo), .dout(new_new_n1939__));
  buf1  g0182(.din(n1500_lo), .dout(new_new_n1940__));
  buf1  g0183(.din(n1512_lo), .dout(new_new_n1942__));
  buf1  g0184(.din(n1515_lo), .dout(new_new_n1944__));
  buf1  g0185(.din(n1518_lo), .dout(new_new_n1946__));
  not1  g0186(.din(n1521_lo), .dout(new_new_n1949__));
  buf1  g0187(.din(n1524_lo), .dout(new_new_n1950__));
  buf1  g0188(.din(n1527_lo), .dout(new_new_n1952__));
  buf1  g0189(.din(n1530_lo), .dout(new_new_n1954__));
  buf1  g0190(.din(n1533_lo), .dout(new_new_n1956__));
  buf1  g0191(.din(n1536_lo), .dout(new_new_n1958__));
  buf1  g0192(.din(n1539_lo), .dout(new_new_n1960__));
  buf1  g0193(.din(n1542_lo), .dout(new_new_n1962__));
  not1  g0194(.din(n1545_lo), .dout(new_new_n1965__));
  buf1  g0195(.din(n1548_lo), .dout(new_new_n1966__));
  buf1  g0196(.din(n1551_lo), .dout(new_new_n1968__));
  buf1  g0197(.din(n1554_lo), .dout(new_new_n1970__));
  not1  g0198(.din(n1554_lo), .dout(new_new_n1971__));
  buf1  g0199(.din(n1560_lo), .dout(new_new_n1972__));
  buf1  g0200(.din(n1563_lo), .dout(new_new_n1974__));
  buf1  g0201(.din(n1566_lo), .dout(new_new_n1976__));
  buf1  g0202(.din(n1572_lo), .dout(new_new_n1978__));
  buf1  g0203(.din(n1575_lo), .dout(new_new_n1980__));
  buf1  g0204(.din(n1578_lo), .dout(new_new_n1982__));
  buf1  g0205(.din(n1584_lo), .dout(new_new_n1984__));
  buf1  g0206(.din(n1587_lo), .dout(new_new_n1986__));
  buf1  g0207(.din(n1590_lo), .dout(new_new_n1988__));
  buf1  g0208(.din(n1596_lo), .dout(new_new_n1990__));
  buf1  g0209(.din(n1599_lo), .dout(new_new_n1992__));
  buf1  g0210(.din(n1602_lo), .dout(new_new_n1994__));
  buf1  g0211(.din(n1608_lo), .dout(new_new_n1996__));
  buf1  g0212(.din(n1611_lo), .dout(new_new_n1998__));
  buf1  g0213(.din(n1614_lo), .dout(new_new_n2000__));
  buf1  g0214(.din(n1620_lo), .dout(new_new_n2002__));
  buf1  g0215(.din(n1623_lo), .dout(new_new_n2004__));
  buf1  g0216(.din(n1626_lo), .dout(new_new_n2006__));
  buf1  g0217(.din(n1632_lo), .dout(new_new_n2008__));
  buf1  g0218(.din(n1635_lo), .dout(new_new_n2010__));
  buf1  g0219(.din(n1638_lo), .dout(new_new_n2012__));
  buf1  g0220(.din(n1644_lo), .dout(new_new_n2014__));
  buf1  g0221(.din(n1647_lo), .dout(new_new_n2016__));
  buf1  g0222(.din(n1650_lo), .dout(new_new_n2018__));
  buf1  g0223(.din(n1656_lo), .dout(new_new_n2020__));
  buf1  g0224(.din(n1659_lo), .dout(new_new_n2022__));
  buf1  g0225(.din(n1662_lo), .dout(new_new_n2024__));
  buf1  g0226(.din(n1668_lo), .dout(new_new_n2026__));
  buf1  g0227(.din(n1671_lo), .dout(new_new_n2028__));
  buf1  g0228(.din(n1674_lo), .dout(new_new_n2030__));
  not1  g0229(.din(n1677_lo), .dout(new_new_n2033__));
  buf1  g0230(.din(n1680_lo), .dout(new_new_n2034__));
  buf1  g0231(.din(n1683_lo), .dout(new_new_n2036__));
  buf1  g0232(.din(n1686_lo), .dout(new_new_n2038__));
  not1  g0233(.din(n1686_lo), .dout(new_new_n2039__));
  buf1  g0234(.din(n1692_lo), .dout(new_new_n2040__));
  buf1  g0235(.din(n1695_lo), .dout(new_new_n2042__));
  buf1  g0236(.din(n1698_lo), .dout(new_new_n2044__));
  buf1  g0237(.din(n1704_lo), .dout(new_new_n2046__));
  buf1  g0238(.din(n1707_lo), .dout(new_new_n2048__));
  buf1  g0239(.din(n1710_lo), .dout(new_new_n2050__));
  buf1  g0240(.din(n1716_lo), .dout(new_new_n2052__));
  buf1  g0241(.din(n1719_lo), .dout(new_new_n2054__));
  buf1  g0242(.din(n1722_lo), .dout(new_new_n2056__));
  buf1  g0243(.din(n1728_lo), .dout(new_new_n2058__));
  buf1  g0244(.din(n1731_lo), .dout(new_new_n2060__));
  buf1  g0245(.din(n1734_lo), .dout(new_new_n2062__));
  buf1  g0246(.din(n1740_lo), .dout(new_new_n2064__));
  buf1  g0247(.din(n1743_lo), .dout(new_new_n2066__));
  buf1  g0248(.din(n1746_lo), .dout(new_new_n2068__));
  not1  g0249(.din(n1749_lo), .dout(new_new_n2071__));
  buf1  g0250(.din(n1752_lo), .dout(new_new_n2072__));
  buf1  g0251(.din(n1755_lo), .dout(new_new_n2074__));
  buf1  g0252(.din(n1758_lo), .dout(new_new_n2076__));
  not1  g0253(.din(n1761_lo), .dout(new_new_n2079__));
  buf1  g0254(.din(n1764_lo), .dout(new_new_n2080__));
  not1  g0255(.din(n1764_lo), .dout(new_new_n2081__));
  buf1  g0256(.din(n1776_lo), .dout(new_new_n2082__));
  buf1  g0257(.din(n1779_lo), .dout(new_new_n2084__));
  buf1  g0258(.din(n1788_lo), .dout(new_new_n2086__));
  buf1  g0259(.din(n1791_lo), .dout(new_new_n2088__));
  buf1  g0260(.din(n1794_lo), .dout(new_new_n2090__));
  not1  g0261(.din(n1797_lo), .dout(new_new_n2093__));
  buf1  g0262(.din(n1800_lo), .dout(new_new_n2094__));
  buf1  g0263(.din(n1812_lo), .dout(new_new_n2096__));
  buf1  g0264(.din(n1824_lo), .dout(new_new_n2098__));
  buf1  g0265(.din(n1836_lo), .dout(new_new_n2100__));
  buf1  g0266(.din(n1848_lo), .dout(new_new_n2102__));
  buf1  g0267(.din(n1860_lo), .dout(new_new_n2104__));
  buf1  g0268(.din(n1872_lo), .dout(new_new_n2106__));
  buf1  g0269(.din(n1884_lo), .dout(new_new_n2108__));
  buf1  g0270(.din(n1896_lo), .dout(new_new_n2110__));
  buf1  g0271(.din(n1899_lo), .dout(new_new_n2112__));
  buf1  g0272(.din(n1908_lo), .dout(new_new_n2114__));
  buf1  g0273(.din(n1911_lo), .dout(new_new_n2116__));
  buf1  g0274(.din(n1920_lo), .dout(new_new_n2118__));
  buf1  g0275(.din(n1923_lo), .dout(new_new_n2120__));
  buf1  g0276(.din(n1926_lo), .dout(new_new_n2122__));
  not1  g0277(.din(n1929_lo), .dout(new_new_n2125__));
  buf1  g0278(.din(n1932_lo), .dout(new_new_n2126__));
  buf1  g0279(.din(n1944_lo), .dout(new_new_n2128__));
  buf1  g0280(.din(n1956_lo), .dout(new_new_n2130__));
  buf1  g0281(.din(n1968_lo), .dout(new_new_n2132__));
  buf1  g0282(.din(n1980_lo), .dout(new_new_n2134__));
  buf1  g0283(.din(n1992_lo), .dout(new_new_n2136__));
  buf1  g0284(.din(n2004_lo), .dout(new_new_n2138__));
  buf1  g0285(.din(n2016_lo), .dout(new_new_n2140__));
  buf1  g0286(.din(n2019_lo), .dout(new_new_n2142__));
  buf1  g0287(.din(n2028_lo), .dout(new_new_n2144__));
  buf1  g0288(.din(n2031_lo), .dout(new_new_n2146__));
  buf1  g0289(.din(n2040_lo), .dout(new_new_n2148__));
  buf1  g0290(.din(n2043_lo), .dout(new_new_n2150__));
  buf1  g0291(.din(n2046_lo), .dout(new_new_n2152__));
  not1  g0292(.din(n2049_lo), .dout(new_new_n2155__));
  buf1  g0293(.din(n2052_lo), .dout(new_new_n2156__));
  buf1  g0294(.din(n2064_lo), .dout(new_new_n2158__));
  buf1  g0295(.din(n2076_lo), .dout(new_new_n2160__));
  buf1  g0296(.din(n2088_lo), .dout(new_new_n2162__));
  buf1  g0297(.din(n2100_lo), .dout(new_new_n2164__));
  buf1  g0298(.din(n2112_lo), .dout(new_new_n2166__));
  buf1  g0299(.din(n2124_lo), .dout(new_new_n2168__));
  buf1  g0300(.din(n2136_lo), .dout(new_new_n2170__));
  buf1  g0301(.din(n2148_lo), .dout(new_new_n2172__));
  buf1  g0302(.din(n2151_lo), .dout(new_new_n2174__));
  buf1  g0303(.din(n2160_lo), .dout(new_new_n2176__));
  buf1  g0304(.din(n2163_lo), .dout(new_new_n2178__));
  buf1  g0305(.din(n2172_lo), .dout(new_new_n2180__));
  buf1  g0306(.din(n2175_lo), .dout(new_new_n2182__));
  buf1  g0307(.din(n2178_lo), .dout(new_new_n2184__));
  not1  g0308(.din(n2181_lo), .dout(new_new_n2187__));
  buf1  g0309(.din(n2184_lo), .dout(new_new_n2188__));
  buf1  g0310(.din(n2196_lo), .dout(new_new_n2190__));
  buf1  g0311(.din(n2208_lo), .dout(new_new_n2192__));
  buf1  g0312(.din(n2220_lo), .dout(new_new_n2194__));
  buf1  g0313(.din(n2232_lo), .dout(new_new_n2196__));
  buf1  g0314(.din(n2244_lo), .dout(new_new_n2198__));
  buf1  g0315(.din(n2256_lo), .dout(new_new_n2200__));
  buf1  g0316(.din(n2268_lo), .dout(new_new_n2202__));
  buf1  g0317(.din(n2280_lo), .dout(new_new_n2204__));
  buf1  g0318(.din(n2283_lo), .dout(new_new_n2206__));
  buf1  g0319(.din(n2292_lo), .dout(new_new_n2208__));
  buf1  g0320(.din(n2295_lo), .dout(new_new_n2210__));
  buf1  g0321(.din(n2298_lo), .dout(new_new_n2212__));
  buf1  g0322(.din(n2301_lo), .dout(new_new_n2214__));
  buf1  g0323(.din(n2304_lo), .dout(new_new_n2216__));
  buf1  g0324(.din(n2316_lo), .dout(new_new_n2218__));
  buf1  g0325(.din(n2319_lo), .dout(new_new_n2220__));
  buf1  g0326(.din(n2322_lo), .dout(new_new_n2222__));
  not1  g0327(.din(n2325_lo), .dout(new_new_n2225__));
  buf1  g0328(.din(n2328_lo), .dout(new_new_n2226__));
  buf1  g0329(.din(n2331_lo), .dout(new_new_n2228__));
  buf1  g0330(.din(n2340_lo), .dout(new_new_n2230__));
  buf1  g0331(.din(n2343_lo), .dout(new_new_n2232__));
  buf1  g0332(.din(n2376_lo), .dout(new_new_n2234__));
  buf1  g0333(.din(n2379_lo), .dout(new_new_n2236__));
  buf1  g0334(.din(n2388_lo), .dout(new_new_n2238__));
  buf1  g0335(.din(n2400_lo), .dout(new_new_n2240__));
  buf1  g0336(.din(n2412_lo), .dout(new_new_n2242__));
  buf1  g0337(.din(n2415_lo), .dout(new_new_n2244__));
  buf1  g0338(.din(n2424_lo), .dout(new_new_n2246__));
  buf1  g0339(.din(n2436_lo), .dout(new_new_n2248__));
  buf1  g0340(.din(n2439_lo), .dout(new_new_n2250__));
  buf1  g0341(.din(n2442_lo), .dout(new_new_n2252__));
  not1  g0342(.din(n2445_lo), .dout(new_new_n2255__));
  buf1  g0343(.din(n2448_lo), .dout(new_new_n2256__));
  buf1  g0344(.din(n2451_lo), .dout(new_new_n2258__));
  buf1  g0345(.din(n2460_lo), .dout(new_new_n2260__));
  buf1  g0346(.din(n2463_lo), .dout(new_new_n2262__));
  buf1  g0347(.din(n2496_lo), .dout(new_new_n2264__));
  buf1  g0348(.din(n2499_lo), .dout(new_new_n2266__));
  buf1  g0349(.din(n2508_lo), .dout(new_new_n2268__));
  buf1  g0350(.din(n2520_lo), .dout(new_new_n2270__));
  buf1  g0351(.din(n2532_lo), .dout(new_new_n2272__));
  buf1  g0352(.din(n2535_lo), .dout(new_new_n2274__));
  buf1  g0353(.din(n2544_lo), .dout(new_new_n2276__));
  buf1  g0354(.din(n2556_lo), .dout(new_new_n2278__));
  buf1  g0355(.din(n2559_lo), .dout(new_new_n2280__));
  buf1  g0356(.din(n2562_lo), .dout(new_new_n2282__));
  not1  g0357(.din(n2565_lo), .dout(new_new_n2285__));
  buf1  g0358(.din(n2568_lo), .dout(new_new_n2286__));
  buf1  g0359(.din(n2571_lo), .dout(new_new_n2288__));
  buf1  g0360(.din(n2580_lo), .dout(new_new_n2290__));
  buf1  g0361(.din(n2583_lo), .dout(new_new_n2292__));
  buf1  g0362(.din(n2616_lo), .dout(new_new_n2294__));
  buf1  g0363(.din(n2619_lo), .dout(new_new_n2296__));
  buf1  g0364(.din(n2628_lo), .dout(new_new_n2298__));
  buf1  g0365(.din(n2640_lo), .dout(new_new_n2300__));
  buf1  g0366(.din(n2652_lo), .dout(new_new_n2302__));
  buf1  g0367(.din(n2655_lo), .dout(new_new_n2304__));
  buf1  g0368(.din(n2664_lo), .dout(new_new_n2306__));
  buf1  g0369(.din(n2676_lo), .dout(new_new_n2308__));
  buf1  g0370(.din(n2679_lo), .dout(new_new_n2310__));
  buf1  g0371(.din(n2682_lo), .dout(new_new_n2312__));
  not1  g0372(.din(n2685_lo), .dout(new_new_n2315__));
  buf1  g0373(.din(n2688_lo), .dout(new_new_n2316__));
  buf1  g0374(.din(n2691_lo), .dout(new_new_n2318__));
  buf1  g0375(.din(n2700_lo), .dout(new_new_n2320__));
  buf1  g0376(.din(n2703_lo), .dout(new_new_n2322__));
  buf1  g0377(.din(n2736_lo), .dout(new_new_n2324__));
  buf1  g0378(.din(n2739_lo), .dout(new_new_n2326__));
  buf1  g0379(.din(n2748_lo), .dout(new_new_n2328__));
  buf1  g0380(.din(n2760_lo), .dout(new_new_n2330__));
  buf1  g0381(.din(n2772_lo), .dout(new_new_n2332__));
  buf1  g0382(.din(n2775_lo), .dout(new_new_n2334__));
  buf1  g0383(.din(n2784_lo), .dout(new_new_n2336__));
  buf1  g0384(.din(n2787_lo), .dout(new_new_n2338__));
  buf1  g0385(.din(n2790_lo), .dout(new_new_n2340__));
  buf1  g0386(.din(n2793_lo), .dout(new_new_n2342__));
  not1  g0387(.din(n2793_lo), .dout(new_new_n2343__));
  buf1  g0388(.din(n2796_lo), .dout(new_new_n2344__));
  buf1  g0389(.din(n2799_lo), .dout(new_new_n2346__));
  buf1  g0390(.din(n2802_lo), .dout(new_new_n2348__));
  not1  g0391(.din(n2805_lo), .dout(new_new_n2351__));
  buf1  g0392(.din(n2808_lo), .dout(new_new_n2352__));
  not1  g0393(.din(n2808_lo), .dout(new_new_n2353__));
  buf1  g0394(.din(n2820_lo), .dout(new_new_n2354__));
  buf1  g0395(.din(n2823_lo), .dout(new_new_n2356__));
  buf1  g0396(.din(n2826_lo), .dout(new_new_n2358__));
  not1  g0397(.din(n2826_lo), .dout(new_new_n2359__));
  buf1  g0398(.din(n2832_lo), .dout(new_new_n2360__));
  buf1  g0399(.din(n2835_lo), .dout(new_new_n2362__));
  buf1  g0400(.din(n2838_lo), .dout(new_new_n2364__));
  buf1  g0401(.din(n2841_lo), .dout(new_new_n2366__));
  not1  g0402(.din(n2841_lo), .dout(new_new_n2367__));
  buf1  g0403(.din(n2844_lo), .dout(new_new_n2368__));
  not1  g0404(.din(n2844_lo), .dout(new_new_n2369__));
  buf1  g0405(.din(n2856_lo), .dout(new_new_n2370__));
  buf1  g0406(.din(n2859_lo), .dout(new_new_n2372__));
  buf1  g0407(.din(n2862_lo), .dout(new_new_n2374__));
  buf1  g0408(.din(n2865_lo), .dout(new_new_n2376__));
  not1  g0409(.din(n2865_lo), .dout(new_new_n2377__));
  buf1  g0410(.din(n2868_lo), .dout(new_new_n2378__));
  buf1  g0411(.din(n2871_lo), .dout(new_new_n2380__));
  buf1  g0412(.din(n2874_lo), .dout(new_new_n2382__));
  buf1  g0413(.din(n2877_lo), .dout(new_new_n2384__));
  not1  g0414(.din(n2877_lo), .dout(new_new_n2385__));
  buf1  g0415(.din(n2880_lo), .dout(new_new_n2386__));
  buf1  g0416(.din(n2883_lo), .dout(new_new_n2388__));
  buf1  g0417(.din(n2886_lo), .dout(new_new_n2390__));
  buf1  g0418(.din(n2889_lo), .dout(new_new_n2392__));
  not1  g0419(.din(n2889_lo), .dout(new_new_n2393__));
  buf1  g0420(.din(n2892_lo), .dout(new_new_n2394__));
  buf1  g0421(.din(n2895_lo), .dout(new_new_n2396__));
  buf1  g0422(.din(n2898_lo), .dout(new_new_n2398__));
  not1  g0423(.din(n2901_lo), .dout(new_new_n2401__));
  buf1  g0424(.din(n2904_lo), .dout(new_new_n2402__));
  buf1  g0425(.din(n2907_lo), .dout(new_new_n2404__));
  buf1  g0426(.din(n2916_lo), .dout(new_new_n2406__));
  buf1  g0427(.din(n2928_lo), .dout(new_new_n2408__));
  buf1  g0428(.din(n2940_lo), .dout(new_new_n2410__));
  buf1  g0429(.din(n2952_lo), .dout(new_new_n2412__));
  buf1  g0430(.din(n2955_lo), .dout(new_new_n2414__));
  not1  g0431(.din(n2955_lo), .dout(new_new_n2415__));
  buf1  g0432(.din(n2964_lo), .dout(new_new_n2416__));
  buf1  g0433(.din(n2976_lo), .dout(new_new_n2418__));
  buf1  g0434(.din(n2988_lo), .dout(new_new_n2420__));
  buf1  g0435(.din(n2991_lo), .dout(new_new_n2422__));
  buf1  g0436(.din(n3000_lo), .dout(new_new_n2424__));
  buf1  g0437(.din(n3003_lo), .dout(new_new_n2426__));
  buf1  g0438(.din(n3012_lo), .dout(new_new_n2428__));
  buf1  g0439(.din(n3015_lo), .dout(new_new_n2430__));
  not1  g0440(.din(n3015_lo), .dout(new_new_n2431__));
  buf1  g0441(.din(n3024_lo), .dout(new_new_n2432__));
  buf1  g0442(.din(n3027_lo), .dout(new_new_n2434__));
  not1  g0443(.din(n3027_lo), .dout(new_new_n2435__));
  buf1  g0444(.din(n3036_lo), .dout(new_new_n2436__));
  buf1  g0445(.din(n3039_lo), .dout(new_new_n2438__));
  not1  g0446(.din(n3039_lo), .dout(new_new_n2439__));
  buf1  g0447(.din(n3048_lo), .dout(new_new_n2440__));
  buf1  g0448(.din(n3051_lo), .dout(new_new_n2442__));
  buf1  g0449(.din(n3054_lo), .dout(new_new_n2444__));
  not1  g0450(.din(n3057_lo), .dout(new_new_n2447__));
  buf1  g0451(.din(n3060_lo), .dout(new_new_n2448__));
  buf1  g0452(.din(n3072_lo), .dout(new_new_n2450__));
  not1  g0453(.din(n3081_lo), .dout(new_new_n2453__));
  buf1  g0454(.din(n3084_lo), .dout(new_new_n2454__));
  buf1  g0455(.din(n3087_lo), .dout(new_new_n2456__));
  not1  g0456(.din(n3087_lo), .dout(new_new_n2457__));
  not1  g0457(.din(n3093_lo), .dout(new_new_n2459__));
  buf1  g0458(.din(n3096_lo), .dout(new_new_n2460__));
  not1  g0459(.din(n3105_lo), .dout(new_new_n2463__));
  buf1  g0460(.din(n3108_lo), .dout(new_new_n2464__));
  not1  g0461(.din(n3117_lo), .dout(new_new_n2467__));
  buf1  g0462(.din(n3120_lo), .dout(new_new_n2468__));
  buf1  g0463(.din(n3123_lo), .dout(new_new_n2470__));
  buf1  g0464(.din(n3126_lo), .dout(new_new_n2472__));
  buf1  g0465(.din(n3129_lo), .dout(new_new_n2474__));
  not1  g0466(.din(n3129_lo), .dout(new_new_n2475__));
  buf1  g0467(.din(n3132_lo), .dout(new_new_n2476__));
  buf1  g0468(.din(n3135_lo), .dout(new_new_n2478__));
  buf1  g0469(.din(n3138_lo), .dout(new_new_n2480__));
  buf1  g0470(.din(n3141_lo), .dout(new_new_n2482__));
  not1  g0471(.din(n3141_lo), .dout(new_new_n2483__));
  buf1  g0472(.din(n3168_lo), .dout(new_new_n2484__));
  buf1  g0473(.din(n3171_lo), .dout(new_new_n2486__));
  buf1  g0474(.din(n3174_lo), .dout(new_new_n2488__));
  buf1  g0475(.din(n3177_lo), .dout(new_new_n2490__));
  not1  g0476(.din(n3177_lo), .dout(new_new_n2491__));
  buf1  g0477(.din(n3180_lo), .dout(new_new_n2492__));
  buf1  g0478(.din(n3183_lo), .dout(new_new_n2494__));
  buf1  g0479(.din(n3192_lo), .dout(new_new_n2496__));
  buf1  g0480(.din(n3195_lo), .dout(new_new_n2498__));
  buf1  g0481(.din(n3204_lo), .dout(new_new_n2500__));
  buf1  g0482(.din(n3207_lo), .dout(new_new_n2502__));
  buf1  g0483(.din(n3216_lo), .dout(new_new_n2504__));
  buf1  g0484(.din(n3219_lo), .dout(new_new_n2506__));
  buf1  g0485(.din(n3228_lo), .dout(new_new_n2508__));
  buf1  g0486(.din(n3231_lo), .dout(new_new_n2510__));
  buf1  g0487(.din(n3240_lo), .dout(new_new_n2512__));
  buf1  g0488(.din(n3243_lo), .dout(new_new_n2514__));
  buf1  g0489(.din(n3252_lo), .dout(new_new_n2516__));
  buf1  g0490(.din(n3255_lo), .dout(new_new_n2518__));
  buf1  g0491(.din(n3258_lo), .dout(new_new_n2520__));
  not1  g0492(.din(n3258_lo), .dout(new_new_n2521__));
  buf1  g0493(.din(n3264_lo), .dout(new_new_n2522__));
  buf1  g0494(.din(n3267_lo), .dout(new_new_n2524__));
  buf1  g0495(.din(n3270_lo), .dout(new_new_n2526__));
  not1  g0496(.din(n3270_lo), .dout(new_new_n2527__));
  buf1  g0497(.din(n3276_lo), .dout(new_new_n2528__));
  buf1  g0498(.din(n3279_lo), .dout(new_new_n2530__));
  buf1  g0499(.din(n3282_lo), .dout(new_new_n2532__));
  not1  g0500(.din(n3282_lo), .dout(new_new_n2533__));
  buf1  g0501(.din(n3288_lo), .dout(new_new_n2534__));
  buf1  g0502(.din(n3291_lo), .dout(new_new_n2536__));
  buf1  g0503(.din(n3294_lo), .dout(new_new_n2538__));
  not1  g0504(.din(n3294_lo), .dout(new_new_n2539__));
  not1  g0505(.din(n4537_o2), .dout(new_new_n2541__));
  not1  g0506(.din(n4538_o2), .dout(new_new_n2543__));
  not1  g0507(.din(n4710_o2), .dout(new_new_n2545__));
  not1  g0508(.din(n4711_o2), .dout(new_new_n2547__));
  buf1  g0509(.din(n1211_inv), .dout(new_new_n2548__));
  buf1  g0510(.din(n1214_inv), .dout(new_new_n2550__));
  buf1  g0511(.din(n1217_inv), .dout(new_new_n2552__));
  buf1  g0512(.din(n1220_inv), .dout(new_new_n2554__));
  not1  g0513(.din(n4927_o2), .dout(new_new_n2557__));
  buf1  g0514(.din(n4928_o2), .dout(new_new_n2558__));
  not1  g0515(.din(n4928_o2), .dout(new_new_n2559__));
  buf1  g0516(.din(n1229_inv), .dout(new_new_n2560__));
  buf1  g0517(.din(n1232_inv), .dout(new_new_n2562__));
  buf1  g0518(.din(n1235_inv), .dout(new_new_n2564__));
  buf1  g0519(.din(n5178_o2), .dout(new_new_n2566__));
  not1  g0520(.din(n5178_o2), .dout(new_new_n2567__));
  buf1  g0521(.din(n5179_o2), .dout(new_new_n2568__));
  not1  g0522(.din(n5179_o2), .dout(new_new_n2569__));
  buf1  g0523(.din(n5477_o2), .dout(new_new_n2570__));
  not1  g0524(.din(n5477_o2), .dout(new_new_n2571__));
  not1  g0525(.din(n5478_o2), .dout(new_new_n2573__));
  buf1  g0526(.din(n5479_o2), .dout(new_new_n2574__));
  not1  g0527(.din(n5479_o2), .dout(new_new_n2575__));
  buf1  g0528(.din(n5222_o2), .dout(new_new_n2576__));
  not1  g0529(.din(n5222_o2), .dout(new_new_n2577__));
  buf1  g0530(.din(n5223_o2), .dout(new_new_n2578__));
  buf1  g0531(.din(n5553_o2), .dout(new_new_n2580__));
  buf1  g0532(.din(n5554_o2), .dout(new_new_n2582__));
  buf1  g0533(.din(G491_o2), .dout(new_new_n2584__));
  buf1  g0534(.din(n2922_lo_buf_o2), .dout(new_new_n2586__));
  not1  g0535(.din(n2922_lo_buf_o2), .dout(new_new_n2587__));
  buf1  g0536(.din(n2946_lo_buf_o2), .dout(new_new_n2588__));
  not1  g0537(.din(n2946_lo_buf_o2), .dout(new_new_n2589__));
  buf1  g0538(.din(n2970_lo_buf_o2), .dout(new_new_n2590__));
  not1  g0539(.din(n2970_lo_buf_o2), .dout(new_new_n2591__));
  buf1  g0540(.din(n2982_lo_buf_o2), .dout(new_new_n2592__));
  not1  g0541(.din(n2982_lo_buf_o2), .dout(new_new_n2593__));
  buf1  g0542(.din(n3066_lo_buf_o2), .dout(new_new_n2594__));
  not1  g0543(.din(n3066_lo_buf_o2), .dout(new_new_n2595__));
  buf1  g0544(.din(n3078_lo_buf_o2), .dout(new_new_n2596__));
  not1  g0545(.din(n3078_lo_buf_o2), .dout(new_new_n2597__));
  buf1  g0546(.din(n3102_lo_buf_o2), .dout(new_new_n2598__));
  not1  g0547(.din(n3102_lo_buf_o2), .dout(new_new_n2599__));
  buf1  g0548(.din(n3114_lo_buf_o2), .dout(new_new_n2600__));
  not1  g0549(.din(n3114_lo_buf_o2), .dout(new_new_n2601__));
  buf1  g0550(.din(G1321_o2), .dout(new_new_n2602__));
  not1  g0551(.din(G1321_o2), .dout(new_new_n2603__));
  buf1  g0552(.din(G1033_o2), .dout(new_new_n2604__));
  buf1  g0553(.din(G1030_o2), .dout(new_new_n2606__));
  buf1  g0554(.din(G1072_o2), .dout(new_new_n2608__));
  buf1  g0555(.din(n1304_inv), .dout(new_new_n2610__));
  buf1  g0556(.din(n1307_inv), .dout(new_new_n2612__));
  buf1  g0557(.din(n2958_lo_buf_o2), .dout(new_new_n2614__));
  not1  g0558(.din(n2958_lo_buf_o2), .dout(new_new_n2615__));
  buf1  g0559(.din(n2994_lo_buf_o2), .dout(new_new_n2616__));
  not1  g0560(.din(n2994_lo_buf_o2), .dout(new_new_n2617__));
  buf1  g0561(.din(n3006_lo_buf_o2), .dout(new_new_n2618__));
  not1  g0562(.din(n3006_lo_buf_o2), .dout(new_new_n2619__));
  buf1  g0563(.din(n3030_lo_buf_o2), .dout(new_new_n2620__));
  not1  g0564(.din(n3030_lo_buf_o2), .dout(new_new_n2621__));
  buf1  g0565(.din(n3042_lo_buf_o2), .dout(new_new_n2622__));
  not1  g0566(.din(n3042_lo_buf_o2), .dout(new_new_n2623__));
  buf1  g0567(.din(n3090_lo_buf_o2), .dout(new_new_n2624__));
  not1  g0568(.din(n3090_lo_buf_o2), .dout(new_new_n2625__));
  buf1  g0569(.din(n1328_inv), .dout(new_new_n2626__));
  buf1  g0570(.din(n1331_inv), .dout(new_new_n2628__));
  buf1  g0571(.din(n1334_inv), .dout(new_new_n2630__));
  buf1  g0572(.din(n1337_inv), .dout(new_new_n2632__));
  buf1  g0573(.din(n1340_inv), .dout(new_new_n2634__));
  buf1  g0574(.din(n1343_inv), .dout(new_new_n2636__));
  buf1  g0575(.din(n1346_inv), .dout(new_new_n2638__));
  buf1  g0576(.din(n1349_inv), .dout(new_new_n2640__));
  buf1  g0577(.din(G1036_o2), .dout(new_new_n2642__));
  buf1  g0578(.din(G1062_o2), .dout(new_new_n2644__));
  buf1  g0579(.din(G1067_o2), .dout(new_new_n2646__));
  buf1  g0580(.din(G1014_o2), .dout(new_new_n2648__));
  buf1  g0581(.din(n1364_inv), .dout(new_new_n2650__));
  buf1  g0582(.din(n1367_inv), .dout(new_new_n2652__));
  buf1  g0583(.din(n3018_lo_buf_o2), .dout(new_new_n2654__));
  not1  g0584(.din(n3018_lo_buf_o2), .dout(new_new_n2655__));
  not1  g0585(.din(G766_o2), .dout(new_new_n2657__));
  buf1  g0586(.din(n1376_inv), .dout(new_new_n2658__));
  buf1  g0587(.din(n1379_inv), .dout(new_new_n2660__));
  buf1  g0588(.din(n1382_inv), .dout(new_new_n2662__));
  buf1  g0589(.din(n1385_inv), .dout(new_new_n2664__));
  buf1  g0590(.din(n1388_inv), .dout(new_new_n2666__));
  buf1  g0591(.din(n1391_inv), .dout(new_new_n2668__));
  buf1  g0592(.din(G1017_o2), .dout(new_new_n2670__));
  buf1  g0593(.din(G1008_o2), .dout(new_new_n2672__));
  not1  g0594(.din(G1008_o2), .dout(new_new_n2673__));
  buf1  g0595(.din(n1400_inv), .dout(new_new_n2674__));
  buf1  g0596(.din(n1403_inv), .dout(new_new_n2676__));
  buf1  g0597(.din(n2910_lo_buf_o2), .dout(new_new_n2678__));
  not1  g0598(.din(n2910_lo_buf_o2), .dout(new_new_n2679__));
  buf1  g0599(.din(n1409_inv), .dout(new_new_n2680__));
  buf1  g0600(.din(G2138_o2), .dout(new_new_n2682__));
  not1  g0601(.din(G2138_o2), .dout(new_new_n2683__));
  buf1  g0602(.din(G2147_o2), .dout(new_new_n2684__));
  not1  g0603(.din(G2147_o2), .dout(new_new_n2685__));
  buf1  g0604(.din(n1418_inv), .dout(new_new_n2686__));
  buf1  g0605(.din(G1137_o2), .dout(new_new_n2688__));
  not1  g0606(.din(G1137_o2), .dout(new_new_n2689__));
  buf1  g0607(.din(G1329_o2), .dout(new_new_n2690__));
  not1  g0608(.din(G1329_o2), .dout(new_new_n2691__));
  buf1  g0609(.din(G374_o2), .dout(new_new_n2692__));
  not1  g0610(.din(G374_o2), .dout(new_new_n2693__));
  buf1  g0611(.din(G386_o2), .dout(new_new_n2694__));
  not1  g0612(.din(G386_o2), .dout(new_new_n2695__));
  buf1  g0613(.din(G663_o2), .dout(new_new_n2696__));
  not1  g0614(.din(G663_o2), .dout(new_new_n2697__));
  buf1  g0615(.din(G674_o2), .dout(new_new_n2698__));
  not1  g0616(.din(G674_o2), .dout(new_new_n2699__));
  buf1  g0617(.din(G578_o2), .dout(new_new_n2700__));
  not1  g0618(.din(G578_o2), .dout(new_new_n2701__));
  buf1  g0619(.din(G575_o2), .dout(new_new_n2702__));
  not1  g0620(.din(G575_o2), .dout(new_new_n2703__));
  not1  g0621(.din(G2505_o2), .dout(new_new_n2705__));
  buf1  g0622(.din(n1448_inv), .dout(new_new_n2706__));
  not1  g0623(.din(n1448_inv), .dout(new_new_n2707__));
  buf1  g0624(.din(G987_o2), .dout(new_new_n2708__));
  not1  g0625(.din(G987_o2), .dout(new_new_n2709__));
  buf1  g0626(.din(G984_o2), .dout(new_new_n2710__));
  not1  g0627(.din(G984_o2), .dout(new_new_n2711__));
  buf1  g0628(.din(G1862_o2), .dout(new_new_n2712__));
  not1  g0629(.din(G1862_o2), .dout(new_new_n2713__));
  buf1  g0630(.din(G1859_o2), .dout(new_new_n2714__));
  not1  g0631(.din(G1859_o2), .dout(new_new_n2715__));
  not1  g0632(.din(G1260_o2), .dout(new_new_n2717__));
  buf1  g0633(.din(G1865_o2), .dout(new_new_n2718__));
  not1  g0634(.din(G2073_o2), .dout(new_new_n2721__));
  buf1  g0635(.din(G1402_o2), .dout(new_new_n2722__));
  not1  g0636(.din(G2048_o2), .dout(new_new_n2725__));
  buf1  g0637(.din(G2276_o2), .dout(new_new_n2726__));
  buf1  g0638(.din(n1481_inv), .dout(new_new_n2728__));
  buf1  g0639(.din(G2141_o2), .dout(new_new_n2730__));
  not1  g0640(.din(G2141_o2), .dout(new_new_n2731__));
  buf1  g0641(.din(G2008_o2), .dout(new_new_n2732__));
  not1  g0642(.din(G2008_o2), .dout(new_new_n2733__));
  buf1  g0643(.din(G2011_o2), .dout(new_new_n2734__));
  not1  g0644(.din(G2011_o2), .dout(new_new_n2735__));
  buf1  g0645(.din(G2150_o2), .dout(new_new_n2736__));
  not1  g0646(.din(G2150_o2), .dout(new_new_n2737__));
  buf1  g0647(.din(G2026_o2), .dout(new_new_n2738__));
  not1  g0648(.din(G2026_o2), .dout(new_new_n2739__));
  buf1  g0649(.din(G2029_o2), .dout(new_new_n2740__));
  not1  g0650(.din(G2029_o2), .dout(new_new_n2741__));
  buf1  g0651(.din(G2023_o2), .dout(new_new_n2742__));
  buf1  g0652(.din(G2041_o2), .dout(new_new_n2744__));
  buf1  g0653(.din(G2017_o2), .dout(new_new_n2746__));
  buf1  g0654(.din(G2020_o2), .dout(new_new_n2748__));
  buf1  g0655(.din(G2035_o2), .dout(new_new_n2750__));
  buf1  g0656(.din(G2038_o2), .dout(new_new_n2752__));
  buf1  g0657(.din(G2228_o2), .dout(new_new_n2754__));
  not1  g0658(.din(G2228_o2), .dout(new_new_n2755__));
  buf1  g0659(.din(G2231_o2), .dout(new_new_n2756__));
  not1  g0660(.din(G2231_o2), .dout(new_new_n2757__));
  buf1  g0661(.din(G2234_o2), .dout(new_new_n2758__));
  not1  g0662(.din(G2234_o2), .dout(new_new_n2759__));
  buf1  g0663(.din(G2237_o2), .dout(new_new_n2760__));
  not1  g0664(.din(G2237_o2), .dout(new_new_n2761__));
  buf1  g0665(.din(G1904_o2), .dout(new_new_n2762__));
  not1  g0666(.din(G1904_o2), .dout(new_new_n2763__));
  buf1  g0667(.din(G1907_o2), .dout(new_new_n2764__));
  not1  g0668(.din(G1907_o2), .dout(new_new_n2765__));
  buf1  g0669(.din(G1928_o2), .dout(new_new_n2766__));
  not1  g0670(.din(G1928_o2), .dout(new_new_n2767__));
  buf1  g0671(.din(G1931_o2), .dout(new_new_n2768__));
  not1  g0672(.din(G1931_o2), .dout(new_new_n2769__));
  not1  g0673(.din(G1893_o2), .dout(new_new_n2771__));
  not1  g0674(.din(G1896_o2), .dout(new_new_n2773__));
  not1  g0675(.din(G1899_o2), .dout(new_new_n2775__));
  not1  g0676(.din(G1937_o2), .dout(new_new_n2777__));
  not1  g0677(.din(G1940_o2), .dout(new_new_n2779__));
  not1  g0678(.din(G1943_o2), .dout(new_new_n2781__));
  buf1  g0679(.din(G1336_o2), .dout(new_new_n2782__));
  not1  g0680(.din(G1336_o2), .dout(new_new_n2783__));
  buf1  g0681(.din(G1996_o2), .dout(new_new_n2784__));
  not1  g0682(.din(G1996_o2), .dout(new_new_n2785__));
  buf1  g0683(.din(G1999_o2), .dout(new_new_n2786__));
  not1  g0684(.din(G1999_o2), .dout(new_new_n2787__));
  buf1  g0685(.din(G2002_o2), .dout(new_new_n2788__));
  not1  g0686(.din(G2002_o2), .dout(new_new_n2789__));
  buf1  g0687(.din(G2005_o2), .dout(new_new_n2790__));
  not1  g0688(.din(G2005_o2), .dout(new_new_n2791__));
  buf1  g0689(.din(G2014_o2), .dout(new_new_n2792__));
  buf1  g0690(.din(G2032_o2), .dout(new_new_n2794__));
  buf1  g0691(.din(G1076_o2), .dout(new_new_n2796__));
  buf1  g0692(.din(G1002_o2), .dout(new_new_n2798__));
  not1  g0693(.din(G1002_o2), .dout(new_new_n2799__));
  buf1  g0694(.din(G998_o2), .dout(new_new_n2800__));
  not1  g0695(.din(G1890_o2), .dout(new_new_n2803__));
  not1  g0696(.din(G1934_o2), .dout(new_new_n2805__));
  buf1  g0697(.din(G1044_o2), .dout(new_new_n2806__));
  buf1  g0698(.din(G1039_o2), .dout(new_new_n2808__));
  buf1  g0699(.din(n1770_lo_buf_o2), .dout(new_new_n2810__));
  not1  g0700(.din(n1770_lo_buf_o2), .dout(new_new_n2811__));
  not1  g0701(.din(G342_o2), .dout(new_new_n2813__));
  not1  g0702(.din(G354_o2), .dout(new_new_n2815__));
  buf1  g0703(.din(G1193_o2), .dout(new_new_n2816__));
  not1  g0704(.din(G1193_o2), .dout(new_new_n2817__));
  buf1  g0705(.din(n3234_lo_buf_o2), .dout(new_new_n2818__));
  not1  g0706(.din(n3234_lo_buf_o2), .dout(new_new_n2819__));
  buf1  g0707(.din(n3246_lo_buf_o2), .dout(new_new_n2820__));
  not1  g0708(.din(n3246_lo_buf_o2), .dout(new_new_n2821__));
  buf1  g0709(.din(G783_o2), .dout(new_new_n2822__));
  not1  g0710(.din(G783_o2), .dout(new_new_n2823__));
  buf1  g0711(.din(G786_o2), .dout(new_new_n2824__));
  not1  g0712(.din(G786_o2), .dout(new_new_n2825__));
  buf1  g0713(.din(G792_o2), .dout(new_new_n2826__));
  not1  g0714(.din(G792_o2), .dout(new_new_n2827__));
  buf1  g0715(.din(G795_o2), .dout(new_new_n2828__));
  not1  g0716(.din(G795_o2), .dout(new_new_n2829__));
  buf1  g0717(.din(G815_o2), .dout(new_new_n2830__));
  not1  g0718(.din(G815_o2), .dout(new_new_n2831__));
  buf1  g0719(.din(G818_o2), .dout(new_new_n2832__));
  not1  g0720(.din(G818_o2), .dout(new_new_n2833__));
  buf1  g0721(.din(G824_o2), .dout(new_new_n2834__));
  not1  g0722(.din(G824_o2), .dout(new_new_n2835__));
  buf1  g0723(.din(G827_o2), .dout(new_new_n2836__));
  not1  g0724(.din(G827_o2), .dout(new_new_n2837__));
  buf1  g0725(.din(G789_o2), .dout(new_new_n2838__));
  not1  g0726(.din(G789_o2), .dout(new_new_n2839__));
  buf1  g0727(.din(G798_o2), .dout(new_new_n2840__));
  not1  g0728(.din(G798_o2), .dout(new_new_n2841__));
  buf1  g0729(.din(G801_o2), .dout(new_new_n2842__));
  not1  g0730(.din(G801_o2), .dout(new_new_n2843__));
  buf1  g0731(.din(G807_o2), .dout(new_new_n2844__));
  not1  g0732(.din(G807_o2), .dout(new_new_n2845__));
  buf1  g0733(.din(G812_o2), .dout(new_new_n2846__));
  not1  g0734(.din(G812_o2), .dout(new_new_n2847__));
  buf1  g0735(.din(G821_o2), .dout(new_new_n2848__));
  not1  g0736(.din(G821_o2), .dout(new_new_n2849__));
  buf1  g0737(.din(G804_o2), .dout(new_new_n2850__));
  not1  g0738(.din(G804_o2), .dout(new_new_n2851__));
  buf1  g0739(.din(G780_o2), .dout(new_new_n2852__));
  not1  g0740(.din(G780_o2), .dout(new_new_n2853__));
  buf1  g0741(.din(G1231_o2), .dout(new_new_n2854__));
  not1  g0742(.din(G1231_o2), .dout(new_new_n2855__));
  buf1  g0743(.din(G1572_o2), .dout(new_new_n2856__));
  not1  g0744(.din(G1572_o2), .dout(new_new_n2857__));
  buf1  g0745(.din(G1377_o2), .dout(new_new_n2858__));
  not1  g0746(.din(G1377_o2), .dout(new_new_n2859__));
  buf1  g0747(.din(G1253_o2), .dout(new_new_n2860__));
  not1  g0748(.din(G1253_o2), .dout(new_new_n2861__));
  buf1  g0749(.din(G1359_o2), .dout(new_new_n2862__));
  not1  g0750(.din(G1359_o2), .dout(new_new_n2863__));
  buf1  g0751(.din(G1258_o2), .dout(new_new_n2864__));
  not1  g0752(.din(G1258_o2), .dout(new_new_n2865__));
  buf1  g0753(.din(G1367_o2), .dout(new_new_n2866__));
  not1  g0754(.din(G1367_o2), .dout(new_new_n2867__));
  buf1  g0755(.din(G1358_o2), .dout(new_new_n2868__));
  not1  g0756(.din(G1358_o2), .dout(new_new_n2869__));
  buf1  g0757(.din(G1366_o2), .dout(new_new_n2870__));
  not1  g0758(.din(G1366_o2), .dout(new_new_n2871__));
  buf1  g0759(.din(G2057_o2), .dout(new_new_n2872__));
  not1  g0760(.din(G2057_o2), .dout(new_new_n2873__));
  buf1  g0761(.din(G2117_o2), .dout(new_new_n2874__));
  not1  g0762(.din(G2117_o2), .dout(new_new_n2875__));
  buf1  g0763(.din(G2118_o2), .dout(new_new_n2876__));
  not1  g0764(.din(G2118_o2), .dout(new_new_n2877__));
  buf1  g0765(.din(G1254_o2), .dout(new_new_n2878__));
  not1  g0766(.din(G1254_o2), .dout(new_new_n2879__));
  buf1  g0767(.din(G1259_o2), .dout(new_new_n2880__));
  not1  g0768(.din(G1259_o2), .dout(new_new_n2881__));
  buf1  g0769(.din(G2058_o2), .dout(new_new_n2882__));
  not1  g0770(.din(G2058_o2), .dout(new_new_n2883__));
  not1  g0771(.din(G405_o2), .dout(new_new_n2885__));
  not1  g0772(.din(G417_o2), .dout(new_new_n2887__));
  buf1  g0773(.din(G1269_o2), .dout(new_new_n2888__));
  not1  g0774(.din(G1269_o2), .dout(new_new_n2889__));
  buf1  g0775(.din(G1275_o2), .dout(new_new_n2890__));
  not1  g0776(.din(G1275_o2), .dout(new_new_n2891__));
  buf1  g0777(.din(G1287_o2), .dout(new_new_n2892__));
  not1  g0778(.din(G1287_o2), .dout(new_new_n2893__));
  buf1  g0779(.din(G1266_o2), .dout(new_new_n2894__));
  not1  g0780(.din(G1266_o2), .dout(new_new_n2895__));
  buf1  g0781(.din(G1272_o2), .dout(new_new_n2896__));
  not1  g0782(.din(G1272_o2), .dout(new_new_n2897__));
  buf1  g0783(.din(G1278_o2), .dout(new_new_n2898__));
  not1  g0784(.din(G1278_o2), .dout(new_new_n2899__));
  buf1  g0785(.din(G1281_o2), .dout(new_new_n2900__));
  not1  g0786(.din(G1281_o2), .dout(new_new_n2901__));
  buf1  g0787(.din(G1284_o2), .dout(new_new_n2902__));
  not1  g0788(.din(G1284_o2), .dout(new_new_n2903__));
  buf1  g0789(.din(G1290_o2), .dout(new_new_n2904__));
  not1  g0790(.din(G1290_o2), .dout(new_new_n2905__));
  buf1  g0791(.din(G1293_o2), .dout(new_new_n2906__));
  not1  g0792(.din(G1293_o2), .dout(new_new_n2907__));
  buf1  g0793(.din(G1299_o2), .dout(new_new_n2908__));
  not1  g0794(.din(G1299_o2), .dout(new_new_n2909__));
  buf1  g0795(.din(G1305_o2), .dout(new_new_n2910__));
  not1  g0796(.din(G1305_o2), .dout(new_new_n2911__));
  buf1  g0797(.din(G1296_o2), .dout(new_new_n2912__));
  not1  g0798(.din(G1296_o2), .dout(new_new_n2913__));
  buf1  g0799(.din(G1302_o2), .dout(new_new_n2914__));
  not1  g0800(.din(G1302_o2), .dout(new_new_n2915__));
  buf1  g0801(.din(G1308_o2), .dout(new_new_n2916__));
  not1  g0802(.din(G1308_o2), .dout(new_new_n2917__));
  buf1  g0803(.din(G1311_o2), .dout(new_new_n2918__));
  not1  g0804(.din(G1311_o2), .dout(new_new_n2919__));
  buf1  g0805(.din(G811_o2), .dout(new_new_n2920__));
  not1  g0806(.din(G811_o2), .dout(new_new_n2921__));
  buf1  g0807(.din(G810_o2), .dout(new_new_n2922__));
  not1  g0808(.din(G810_o2), .dout(new_new_n2923__));
  buf1  g0809(.din(G1728_o2), .dout(new_new_n2924__));
  not1  g0810(.din(G1728_o2), .dout(new_new_n2925__));
  buf1  g0811(.din(G2512_o2), .dout(new_new_n2926__));
  buf1  g0812(.din(G1114_o2), .dout(new_new_n2928__));
  not1  g0813(.din(G1114_o2), .dout(new_new_n2929__));
  buf1  g0814(.din(G1113_o2), .dout(new_new_n2930__));
  not1  g0815(.din(G1113_o2), .dout(new_new_n2931__));
  buf1  g0816(.din(G1992_o2), .dout(new_new_n2932__));
  not1  g0817(.din(G1992_o2), .dout(new_new_n2933__));
  buf1  g0818(.din(G1991_o2), .dout(new_new_n2934__));
  not1  g0819(.din(G1991_o2), .dout(new_new_n2935__));
  buf1  g0820(.din(G1426_o2), .dout(new_new_n2936__));
  not1  g0821(.din(G1966_o2), .dout(new_new_n2939__));
  buf1  g0822(.din(G2211_o2), .dout(new_new_n2940__));
  not1  g0823(.din(G1509_o2), .dout(new_new_n2943__));
  buf1  g0824(.din(G2153_o2), .dout(new_new_n2944__));
  not1  g0825(.din(G2329_o2), .dout(new_new_n2947__));
  buf1  g0826(.din(G1540_o2), .dout(new_new_n2948__));
  not1  g0827(.din(G1540_o2), .dout(new_new_n2949__));
  not1  g0828(.din(G2167_o2), .dout(new_new_n2951__));
  not1  g0829(.din(G2191_o2), .dout(new_new_n2953__));
  buf1  g0830(.din(G1234_o2), .dout(new_new_n2954__));
  not1  g0831(.din(G1234_o2), .dout(new_new_n2955__));
  buf1  g0832(.din(G1132_o2), .dout(new_new_n2956__));
  not1  g0833(.din(G1132_o2), .dout(new_new_n2957__));
  buf1  g0834(.din(G1129_o2), .dout(new_new_n2958__));
  not1  g0835(.din(G1129_o2), .dout(new_new_n2959__));
  buf1  g0836(.din(G2088_o2), .dout(new_new_n2960__));
  buf1  g0837(.din(G2106_o2), .dout(new_new_n2962__));
  buf1  g0838(.din(G1314_o2), .dout(new_new_n2964__));
  not1  g0839(.din(G1314_o2), .dout(new_new_n2965__));
  buf1  g0840(.din(G636_o2), .dout(new_new_n2966__));
  buf1  g0841(.din(G647_o2), .dout(new_new_n2968__));
  buf1  g0842(.din(n3186_lo_buf_o2), .dout(new_new_n2970__));
  not1  g0843(.din(n3186_lo_buf_o2), .dout(new_new_n2971__));
  buf1  g0844(.din(n3198_lo_buf_o2), .dout(new_new_n2972__));
  not1  g0845(.din(n3198_lo_buf_o2), .dout(new_new_n2973__));
  buf1  g0846(.din(n3210_lo_buf_o2), .dout(new_new_n2974__));
  not1  g0847(.din(n3210_lo_buf_o2), .dout(new_new_n2975__));
  buf1  g0848(.din(n3222_lo_buf_o2), .dout(new_new_n2976__));
  not1  g0849(.din(n3222_lo_buf_o2), .dout(new_new_n2977__));
  buf1  g0850(.din(G1225_o2), .dout(new_new_n2978__));
  not1  g0851(.din(G1225_o2), .dout(new_new_n2979__));
  buf1  g0852(.din(G1342_o2), .dout(new_new_n2980__));
  not1  g0853(.din(G1342_o2), .dout(new_new_n2981__));
  buf1  g0854(.din(G1222_o2), .dout(new_new_n2982__));
  not1  g0855(.din(G1222_o2), .dout(new_new_n2983__));
  buf1  g0856(.din(G1228_o2), .dout(new_new_n2984__));
  not1  g0857(.din(G1228_o2), .dout(new_new_n2985__));
  buf1  g0858(.din(G1348_o2), .dout(new_new_n2986__));
  not1  g0859(.din(G1348_o2), .dout(new_new_n2987__));
  buf1  g0860(.din(G1345_o2), .dout(new_new_n2988__));
  not1  g0861(.din(G1345_o2), .dout(new_new_n2989__));
  buf1  g0862(.din(G1351_o2), .dout(new_new_n2990__));
  not1  g0863(.din(G1351_o2), .dout(new_new_n2991__));
  buf1  g0864(.din(G2242_o2), .dout(new_new_n2992__));
  not1  g0865(.din(G2242_o2), .dout(new_new_n2993__));
  buf1  g0866(.din(G2260_o2), .dout(new_new_n2994__));
  not1  g0867(.din(G2260_o2), .dout(new_new_n2995__));
  buf1  g0868(.din(G1374_o2), .dout(new_new_n2996__));
  not1  g0869(.din(G1374_o2), .dout(new_new_n2997__));
  buf1  g0870(.din(G1537_o2), .dout(new_new_n2998__));
  not1  g0871(.din(G1537_o2), .dout(new_new_n2999__));
  buf1  g0872(.din(G301_o2), .dout(new_new_n3000__));
  not1  g0873(.din(G301_o2), .dout(new_new_n3001__));
  buf1  g0874(.din(G313_o2), .dout(new_new_n3002__));
  not1  g0875(.din(G313_o2), .dout(new_new_n3003__));
  buf1  g0876(.din(G2365_o2), .dout(new_new_n3004__));
  not1  g0877(.din(G2365_o2), .dout(new_new_n3005__));
  buf1  g0878(.din(G2255_o2), .dout(new_new_n3006__));
  not1  g0879(.din(G2255_o2), .dout(new_new_n3007__));
  buf1  g0880(.din(G2253_o2), .dout(new_new_n3008__));
  not1  g0881(.din(G2253_o2), .dout(new_new_n3009__));
  buf1  g0882(.din(G2395_o2), .dout(new_new_n3010__));
  not1  g0883(.din(G2395_o2), .dout(new_new_n3011__));
  buf1  g0884(.din(G2272_o2), .dout(new_new_n3012__));
  not1  g0885(.din(G2272_o2), .dout(new_new_n3013__));
  buf1  g0886(.din(G2270_o2), .dout(new_new_n3014__));
  not1  g0887(.din(G2270_o2), .dout(new_new_n3015__));
  not1  g0888(.din(G2245_o2), .dout(new_new_n3017__));
  not1  g0889(.din(G2262_o2), .dout(new_new_n3019__));
  not1  g0890(.din(G2249_o2), .dout(new_new_n3021__));
  not1  g0891(.din(G2247_o2), .dout(new_new_n3023__));
  not1  g0892(.din(G2266_o2), .dout(new_new_n3025__));
  not1  g0893(.din(G2264_o2), .dout(new_new_n3027__));
  buf1  g0894(.din(G2403_o2), .dout(new_new_n3028__));
  not1  g0895(.din(G2403_o2), .dout(new_new_n3029__));
  buf1  g0896(.din(G2401_o2), .dout(new_new_n3030__));
  not1  g0897(.din(G2401_o2), .dout(new_new_n3031__));
  buf1  g0898(.din(G2410_o2), .dout(new_new_n3032__));
  not1  g0899(.din(G2410_o2), .dout(new_new_n3033__));
  buf1  g0900(.din(G2408_o2), .dout(new_new_n3034__));
  not1  g0901(.din(G2408_o2), .dout(new_new_n3035__));
  buf1  g0902(.din(G2306_o2), .dout(new_new_n3036__));
  not1  g0903(.din(G2306_o2), .dout(new_new_n3037__));
  buf1  g0904(.din(G2305_o2), .dout(new_new_n3038__));
  not1  g0905(.din(G2305_o2), .dout(new_new_n3039__));
  buf1  g0906(.din(G2314_o2), .dout(new_new_n3040__));
  not1  g0907(.din(G2314_o2), .dout(new_new_n3041__));
  buf1  g0908(.din(G2313_o2), .dout(new_new_n3042__));
  not1  g0909(.din(G2313_o2), .dout(new_new_n3043__));
  buf1  g0910(.din(G2303_o2), .dout(new_new_n3044__));
  buf1  g0911(.din(G2302_o2), .dout(new_new_n3046__));
  buf1  g0912(.din(G2301_o2), .dout(new_new_n3048__));
  buf1  g0913(.din(G2311_o2), .dout(new_new_n3050__));
  buf1  g0914(.din(G2310_o2), .dout(new_new_n3052__));
  buf1  g0915(.din(G2309_o2), .dout(new_new_n3054__));
  buf1  g0916(.din(G2404_o2), .dout(new_new_n3056__));
  not1  g0917(.din(G2404_o2), .dout(new_new_n3057__));
  buf1  g0918(.din(G2411_o2), .dout(new_new_n3058__));
  not1  g0919(.din(G2411_o2), .dout(new_new_n3059__));
  buf1  g0920(.din(G2420_o2), .dout(new_new_n3060__));
  not1  g0921(.din(G2420_o2), .dout(new_new_n3061__));
  buf1  g0922(.din(G2419_o2), .dout(new_new_n3062__));
  not1  g0923(.din(G2419_o2), .dout(new_new_n3063__));
  buf1  g0924(.din(G2433_o2), .dout(new_new_n3064__));
  not1  g0925(.din(G2433_o2), .dout(new_new_n3065__));
  buf1  g0926(.din(G2432_o2), .dout(new_new_n3066__));
  not1  g0927(.din(G2432_o2), .dout(new_new_n3067__));
  buf1  g0928(.din(G402_o2), .dout(new_new_n3068__));
  not1  g0929(.din(G402_o2), .dout(new_new_n3069__));
  buf1  g0930(.din(G403_o2), .dout(new_new_n3070__));
  not1  g0931(.din(G403_o2), .dout(new_new_n3071__));
  buf1  g0932(.din(G1053_o2), .dout(new_new_n3072__));
  not1  g0933(.din(G1053_o2), .dout(new_new_n3073__));
  buf1  g0934(.din(G1049_o2), .dout(new_new_n3074__));
  not1  g0935(.din(G1049_o2), .dout(new_new_n3075__));
  buf1  g0936(.din(n2003_inv), .dout(new_new_n3076__));
  not1  g0937(.din(n2003_inv), .dout(new_new_n3077__));
  buf1  g0938(.din(G1364_o2), .dout(new_new_n3078__));
  not1  g0939(.din(G1364_o2), .dout(new_new_n3079__));
  buf1  g0940(.din(G1079_o2), .dout(new_new_n3080__));
  not1  g0941(.din(G1079_o2), .dout(new_new_n3081__));
  buf1  g0942(.din(G1478_o2), .dout(new_new_n3082__));
  not1  g0943(.din(G1478_o2), .dout(new_new_n3083__));
  buf1  g0944(.din(G707_o2), .dout(new_new_n3084__));
  buf1  g0945(.din(G718_o2), .dout(new_new_n3086__));
  buf1  g0946(.din(G2417_o2), .dout(new_new_n3088__));
  not1  g0947(.din(G2417_o2), .dout(new_new_n3089__));
  buf1  g0948(.din(G2414_o2), .dout(new_new_n3090__));
  not1  g0949(.din(G2414_o2), .dout(new_new_n3091__));
  buf1  g0950(.din(G2431_o2), .dout(new_new_n3092__));
  not1  g0951(.din(G2431_o2), .dout(new_new_n3093__));
  buf1  g0952(.din(G2428_o2), .dout(new_new_n3094__));
  not1  g0953(.din(G2428_o2), .dout(new_new_n3095__));
  buf1  g0954(.din(G1653_o2), .dout(new_new_n3096__));
  not1  g0955(.din(G1653_o2), .dout(new_new_n3097__));
  buf1  g0956(.din(G2213_o2), .dout(new_new_n3098__));
  not1  g0957(.din(G2213_o2), .dout(new_new_n3099__));
  buf1  g0958(.din(G2221_o2), .dout(new_new_n3100__));
  not1  g0959(.din(G2221_o2), .dout(new_new_n3101__));
  buf1  g0960(.din(G2250_o2), .dout(new_new_n3102__));
  buf1  g0961(.din(G2267_o2), .dout(new_new_n3104__));
  buf1  g0962(.din(G1365_o2), .dout(new_new_n3106__));
  not1  g0963(.din(G1365_o2), .dout(new_new_n3107__));
  buf1  g0964(.din(G1368_o2), .dout(new_new_n3108__));
  not1  g0965(.din(G1368_o2), .dout(new_new_n3109__));
  buf1  g0966(.din(G1371_o2), .dout(new_new_n3110__));
  not1  g0967(.din(G1371_o2), .dout(new_new_n3111__));
  not1  g0968(.din(G2218_o2), .dout(new_new_n3113__));
  not1  g0969(.din(G2225_o2), .dout(new_new_n3115__));
  not1  g0970(.din(n1503_lo_buf_o2), .dout(new_new_n3117__));
  buf1  g0971(.din(n1863_lo_buf_o2), .dout(new_new_n3118__));
  not1  g0972(.din(n1863_lo_buf_o2), .dout(new_new_n3119__));
  buf1  g0973(.din(n1887_lo_buf_o2), .dout(new_new_n3120__));
  not1  g0974(.din(n1887_lo_buf_o2), .dout(new_new_n3121__));
  buf1  g0975(.din(n1983_lo_buf_o2), .dout(new_new_n3122__));
  not1  g0976(.din(n1983_lo_buf_o2), .dout(new_new_n3123__));
  buf1  g0977(.din(n2007_lo_buf_o2), .dout(new_new_n3124__));
  not1  g0978(.din(n2007_lo_buf_o2), .dout(new_new_n3125__));
  buf1  g0979(.din(n2115_lo_buf_o2), .dout(new_new_n3126__));
  not1  g0980(.din(n2115_lo_buf_o2), .dout(new_new_n3127__));
  buf1  g0981(.din(n2139_lo_buf_o2), .dout(new_new_n3128__));
  not1  g0982(.din(n2139_lo_buf_o2), .dout(new_new_n3129__));
  buf1  g0983(.din(n2247_lo_buf_o2), .dout(new_new_n3130__));
  not1  g0984(.din(n2247_lo_buf_o2), .dout(new_new_n3131__));
  buf1  g0985(.din(n2271_lo_buf_o2), .dout(new_new_n3132__));
  not1  g0986(.din(n2271_lo_buf_o2), .dout(new_new_n3133__));
  buf1  g0987(.din(n2919_lo_buf_o2), .dout(new_new_n3134__));
  not1  g0988(.din(n2919_lo_buf_o2), .dout(new_new_n3135__));
  buf1  g0989(.din(n2943_lo_buf_o2), .dout(new_new_n3136__));
  not1  g0990(.din(n2943_lo_buf_o2), .dout(new_new_n3137__));
  buf1  g0991(.din(n2967_lo_buf_o2), .dout(new_new_n3138__));
  buf1  g0992(.din(n2979_lo_buf_o2), .dout(new_new_n3140__));
  buf1  g0993(.din(n3063_lo_buf_o2), .dout(new_new_n3142__));
  not1  g0994(.din(n3063_lo_buf_o2), .dout(new_new_n3143__));
  buf1  g0995(.din(n3075_lo_buf_o2), .dout(new_new_n3144__));
  not1  g0996(.din(n3075_lo_buf_o2), .dout(new_new_n3145__));
  buf1  g0997(.din(n3099_lo_buf_o2), .dout(new_new_n3146__));
  buf1  g0998(.din(n3111_lo_buf_o2), .dout(new_new_n3148__));
  buf1  g0999(.din(G878_o2), .dout(new_new_n3150__));
  buf1  g1000(.din(G875_o2), .dout(new_new_n3152__));
  buf1  g1001(.din(G661_o2), .dout(new_new_n3154__));
  buf1  g1002(.din(G660_o2), .dout(new_new_n3156__));
  buf1  g1003(.din(G879_o2), .dout(new_new_n3158__));
  buf1  g1004(.din(G876_o2), .dout(new_new_n3160__));
  buf1  g1005(.din(G1320_o2), .dout(new_new_n3162__));
  not1  g1006(.din(G1320_o2), .dout(new_new_n3163__));
  buf1  g1007(.din(G941_o2), .dout(new_new_n3164__));
  buf1  g1008(.din(G732_o2), .dout(new_new_n3166__));
  buf1  g1009(.din(G942_o2), .dout(new_new_n3168__));
  buf1  g1010(.din(G1493_o2), .dout(new_new_n3170__));
  not1  g1011(.din(G1493_o2), .dout(new_new_n3171__));
  buf1  g1012(.din(G1498_o2), .dout(new_new_n3172__));
  not1  g1013(.din(G1498_o2), .dout(new_new_n3173__));
  buf1  g1014(.din(G877_o2), .dout(new_new_n3174__));
  buf1  g1015(.din(G874_o2), .dout(new_new_n3176__));
  buf1  g1016(.din(n1806_lo_buf_o2), .dout(new_new_n3178__));
  buf1  g1017(.din(n1878_lo_buf_o2), .dout(new_new_n3180__));
  not1  g1018(.din(n1878_lo_buf_o2), .dout(new_new_n3181__));
  buf1  g1019(.din(n1938_lo_buf_o2), .dout(new_new_n3182__));
  buf1  g1020(.din(n1998_lo_buf_o2), .dout(new_new_n3184__));
  not1  g1021(.din(n1998_lo_buf_o2), .dout(new_new_n3185__));
  buf1  g1022(.din(n2058_lo_buf_o2), .dout(new_new_n3186__));
  buf1  g1023(.din(n2130_lo_buf_o2), .dout(new_new_n3188__));
  not1  g1024(.din(n2130_lo_buf_o2), .dout(new_new_n3189__));
  buf1  g1025(.din(n2190_lo_buf_o2), .dout(new_new_n3190__));
  buf1  g1026(.din(n2262_lo_buf_o2), .dout(new_new_n3192__));
  not1  g1027(.din(n2262_lo_buf_o2), .dout(new_new_n3193__));
  buf1  g1028(.din(n2310_lo_buf_o2), .dout(new_new_n3194__));
  buf1  g1029(.din(n2406_lo_buf_o2), .dout(new_new_n3196__));
  buf1  g1030(.din(n2430_lo_buf_o2), .dout(new_new_n3198__));
  buf1  g1031(.din(n2526_lo_buf_o2), .dout(new_new_n3200__));
  buf1  g1032(.din(n2550_lo_buf_o2), .dout(new_new_n3202__));
  buf1  g1033(.din(n2646_lo_buf_o2), .dout(new_new_n3204__));
  buf1  g1034(.din(n2670_lo_buf_o2), .dout(new_new_n3206__));
  buf1  g1035(.din(n2766_lo_buf_o2), .dout(new_new_n3208__));
  buf1  g1036(.din(G603_o2), .dout(new_new_n3210__));
  not1  g1037(.din(G603_o2), .dout(new_new_n3211__));
  buf1  g1038(.din(G614_o2), .dout(new_new_n3212__));
  not1  g1039(.din(G614_o2), .dout(new_new_n3213__));
  buf1  g1040(.din(G1026_o2), .dout(new_new_n3214__));
  buf1  g1041(.din(G1021_o2), .dout(new_new_n3216__));
  buf1  g1042(.din(G940_o2), .dout(new_new_n3218__));
  buf1  g1043(.din(G1636_o2), .dout(new_new_n3220__));
  not1  g1044(.din(G1636_o2), .dout(new_new_n3221__));
  buf1  g1045(.din(G1684_o2), .dout(new_new_n3222__));
  not1  g1046(.din(G1684_o2), .dout(new_new_n3223__));
  buf1  g1047(.din(n2352_lo_buf_o2), .dout(new_new_n3224__));
  not1  g1048(.din(n2364_lo_buf_o2), .dout(new_new_n3227__));
  buf1  g1049(.din(n2472_lo_buf_o2), .dout(new_new_n3228__));
  not1  g1050(.din(n2484_lo_buf_o2), .dout(new_new_n3231__));
  buf1  g1051(.din(n2592_lo_buf_o2), .dout(new_new_n3232__));
  not1  g1052(.din(n2604_lo_buf_o2), .dout(new_new_n3235__));
  buf1  g1053(.din(n2712_lo_buf_o2), .dout(new_new_n3236__));
  not1  g1054(.din(n2724_lo_buf_o2), .dout(new_new_n3239__));
  buf1  g1055(.din(n3150_lo_buf_o2), .dout(new_new_n3240__));
  not1  g1056(.din(n3150_lo_buf_o2), .dout(new_new_n3241__));
  buf1  g1057(.din(n3162_lo_buf_o2), .dout(new_new_n3242__));
  not1  g1058(.din(n3162_lo_buf_o2), .dout(new_new_n3243__));
  or1   g1059(.dina(new_new_n2467__), .dinb(new_new_n2463__), .dout(new_new_n3244__));
  or1   g1060(.dina(new_new_n3244__), .dinb(new_new_n2459__), .dout(new_new_n3245__));
  or1   g1061(.dina(new_new_n3245__), .dinb(new_new_n2453__), .dout(new_new_n3246__));
  or1   g1062(.dina(new_new_n1965__), .dinb(new_new_n1905__), .dout(new_new_n3247__));
  or1   g1063(.dina(new_new_n3247__), .dinb(new_new_n5047__), .dout(new_new_n3248__));
  and1  g1064(.dina(new_new_n5049__), .dinb(new_new_n2214__), .dout(new_new_n3249__));
  or1   g1065(.dina(new_new_n5047__), .dinb(new_new_n1939__), .dout(new_new_n3250__));
  or1   g1066(.dina(new_new_n5052__), .dinb(new_new_n2367__), .dout(new_new_n3251__));
  or1   g1067(.dina(new_new_n5052__), .dinb(new_new_n2491__), .dout(new_new_n3252__));
  or1   g1068(.dina(new_new_n5053__), .dinb(new_new_n5054__), .dout(new_new_n3253__));
  or1   g1069(.dina(new_new_n3253__), .dinb(new_new_n5055__), .dout(new_new_n3254__));
  or1   g1070(.dina(new_new_n3254__), .dinb(new_new_n5056__), .dout(new_new_n3255__));
  or1   g1071(.dina(new_new_n5057__), .dinb(new_new_n5058__), .dout(new_new_n3256__));
  or1   g1072(.dina(new_new_n3256__), .dinb(new_new_n5059__), .dout(new_new_n3257__));
  or1   g1073(.dina(new_new_n3257__), .dinb(new_new_n5060__), .dout(new_new_n3258__));
  or1   g1074(.dina(new_new_n5061__), .dinb(new_new_n5062__), .dout(new_new_n3259__));
  and1  g1075(.dina(new_new_n5061__), .dinb(new_new_n2490__), .dout(new_new_n3260__));
  and1  g1076(.dina(new_new_n5062__), .dinb(new_new_n2366__), .dout(new_new_n3261__));
  or1   g1077(.dina(new_new_n3261__), .dinb(new_new_n3260__), .dout(new_new_n3262__));
  and1  g1078(.dina(new_new_n2566__), .dinb(new_new_n5064__), .dout(new_new_n3263__));
  or1   g1079(.dina(new_new_n3263__), .dinb(new_new_n5066__), .dout(new_new_n3264__));
  or1   g1080(.dina(new_new_n2376__), .dinb(new_new_n2351__), .dout(new_new_n3265__));
  or1   g1081(.dina(new_new_n5067__), .dinb(new_new_n2071__), .dout(new_new_n3266__));
  or1   g1082(.dina(new_new_n3266__), .dinb(new_new_n5069__), .dout(new_new_n3267__));
  and1  g1083(.dina(new_new_n1912__), .dinb(new_new_n1896__), .dout(new_new_n3268__));
  or1   g1084(.dina(new_new_n5067__), .dinb(new_new_n5069__), .dout(new_new_n3269__));
  or1   g1085(.dina(new_new_n3269__), .dinb(new_new_n3268__), .dout(new_new_n3270__));
  or1   g1086(.dina(new_new_n2559__), .dinb(new_new_n5073__), .dout(new_new_n3271__));
  or1   g1087(.dina(new_new_n5075__), .dinb(new_new_n5078__), .dout(new_new_n3272__));
  and1  g1088(.dina(new_new_n3272__), .dinb(new_new_n3271__), .dout(new_new_n3273__));
  or1   g1089(.dina(new_new_n5080__), .dinb(new_new_n5073__), .dout(new_new_n3274__));
  or1   g1090(.dina(new_new_n5081__), .dinb(new_new_n5078__), .dout(new_new_n3275__));
  and1  g1091(.dina(new_new_n3275__), .dinb(new_new_n3274__), .dout(new_new_n3276__));
  and1  g1092(.dina(new_new_n2602__), .dinb(new_new_n5066__), .dout(new_new_n3277__));
  and1  g1093(.dina(new_new_n2558__), .dinb(new_new_n5064__), .dout(new_new_n3278__));
  or1   g1094(.dina(new_new_n3278__), .dinb(new_new_n3277__), .dout(new_new_n3279__));
  or1   g1095(.dina(new_new_n2567__), .dinb(new_new_n5072__), .dout(new_new_n3280__));
  or1   g1096(.dina(new_new_n2603__), .dinb(new_new_n5077__), .dout(new_new_n3281__));
  and1  g1097(.dina(new_new_n3281__), .dinb(new_new_n3280__), .dout(new_new_n3282__));
  or1   g1098(.dina(new_new_n2574__), .dinb(new_new_n2482__), .dout(new_new_n3283__));
  and1  g1099(.dina(new_new_n5082__), .dinb(new_new_n2483__), .dout(new_new_n3284__));
  and1  g1100(.dina(new_new_n5082__), .dinb(new_new_n2575__), .dout(new_new_n3285__));
  or1   g1101(.dina(new_new_n3285__), .dinb(new_new_n3284__), .dout(new_new_n3286__));
  or1   g1102(.dina(new_new_n5083__), .dinb(new_new_n2474__), .dout(new_new_n3287__));
  and1  g1103(.dina(new_new_n5084__), .dinb(new_new_n2475__), .dout(new_new_n3288__));
  and1  g1104(.dina(new_new_n5084__), .dinb(new_new_n2570__), .dout(new_new_n3289__));
  or1   g1105(.dina(new_new_n3289__), .dinb(new_new_n3288__), .dout(new_new_n3290__));
  or1   g1106(.dina(new_new_n3290__), .dinb(new_new_n3286__), .dout(new_new_n3291__));
  or1   g1107(.dina(new_new_n2943__), .dinb(new_new_n2717__), .dout(new_new_n3292__));
  or1   g1108(.dina(new_new_n2936__), .dinb(new_new_n2722__), .dout(new_new_n3293__));
  and1  g1109(.dina(new_new_n3293__), .dinb(new_new_n3292__), .dout(new_new_n3294__));
  and1  g1110(.dina(new_new_n3294__), .dinb(new_new_n1956__), .dout(new_new_n3295__));
  and1  g1111(.dina(new_new_n2922__), .dinb(new_new_n2701__), .dout(new_new_n3296__));
  or1   g1112(.dina(new_new_n2923__), .dinb(new_new_n2700__), .dout(new_new_n3297__));
  and1  g1113(.dina(new_new_n2920__), .dinb(new_new_n2703__), .dout(new_new_n3298__));
  or1   g1114(.dina(new_new_n2921__), .dinb(new_new_n2702__), .dout(new_new_n3299__));
  and1  g1115(.dina(new_new_n3299__), .dinb(new_new_n3297__), .dout(new_new_n3300__));
  or1   g1116(.dina(new_new_n3298__), .dinb(new_new_n3296__), .dout(new_new_n3301__));
  and1  g1117(.dina(new_new_n2881__), .dinb(new_new_n2867__), .dout(new_new_n3302__));
  or1   g1118(.dina(new_new_n2880__), .dinb(new_new_n2866__), .dout(new_new_n3303__));
  and1  g1119(.dina(new_new_n2871__), .dinb(new_new_n2865__), .dout(new_new_n3304__));
  or1   g1120(.dina(new_new_n2870__), .dinb(new_new_n2864__), .dout(new_new_n3305__));
  and1  g1121(.dina(new_new_n3304__), .dinb(new_new_n3302__), .dout(new_new_n3306__));
  or1   g1122(.dina(new_new_n3305__), .dinb(new_new_n3303__), .dout(new_new_n3307__));
  or1   g1123(.dina(new_new_n3307__), .dinb(new_new_n3300__), .dout(new_new_n3308__));
  or1   g1124(.dina(new_new_n3306__), .dinb(new_new_n3301__), .dout(new_new_n3309__));
  and1  g1125(.dina(new_new_n3309__), .dinb(new_new_n3308__), .dout(new_new_n3310__));
  and1  g1126(.dina(new_new_n2931__), .dinb(new_new_n2708__), .dout(new_new_n3311__));
  or1   g1127(.dina(new_new_n2930__), .dinb(new_new_n2709__), .dout(new_new_n3312__));
  and1  g1128(.dina(new_new_n2929__), .dinb(new_new_n2710__), .dout(new_new_n3313__));
  or1   g1129(.dina(new_new_n2928__), .dinb(new_new_n2711__), .dout(new_new_n3314__));
  and1  g1130(.dina(new_new_n3314__), .dinb(new_new_n3312__), .dout(new_new_n3315__));
  or1   g1131(.dina(new_new_n3313__), .dinb(new_new_n3311__), .dout(new_new_n3316__));
  and1  g1132(.dina(new_new_n2879__), .dinb(new_new_n2863__), .dout(new_new_n3317__));
  or1   g1133(.dina(new_new_n2878__), .dinb(new_new_n2862__), .dout(new_new_n3318__));
  and1  g1134(.dina(new_new_n2869__), .dinb(new_new_n2861__), .dout(new_new_n3319__));
  or1   g1135(.dina(new_new_n2868__), .dinb(new_new_n2860__), .dout(new_new_n3320__));
  and1  g1136(.dina(new_new_n3319__), .dinb(new_new_n3317__), .dout(new_new_n3321__));
  or1   g1137(.dina(new_new_n3320__), .dinb(new_new_n3318__), .dout(new_new_n3322__));
  or1   g1138(.dina(new_new_n3322__), .dinb(new_new_n3315__), .dout(new_new_n3323__));
  or1   g1139(.dina(new_new_n3321__), .dinb(new_new_n3316__), .dout(new_new_n3324__));
  and1  g1140(.dina(new_new_n3324__), .dinb(new_new_n3323__), .dout(new_new_n3325__));
  and1  g1141(.dina(new_new_n2906__), .dinb(new_new_n2845__), .dout(new_new_n3326__));
  and1  g1142(.dina(new_new_n2907__), .dinb(new_new_n2844__), .dout(new_new_n3327__));
  or1   g1143(.dina(new_new_n3327__), .dinb(new_new_n3326__), .dout(new_new_n3328__));
  and1  g1144(.dina(new_new_n2904__), .dinb(new_new_n2851__), .dout(new_new_n3329__));
  and1  g1145(.dina(new_new_n2905__), .dinb(new_new_n2850__), .dout(new_new_n3330__));
  or1   g1146(.dina(new_new_n3330__), .dinb(new_new_n3329__), .dout(new_new_n3331__));
  and1  g1147(.dina(new_new_n2892__), .dinb(new_new_n2843__), .dout(new_new_n3332__));
  and1  g1148(.dina(new_new_n2893__), .dinb(new_new_n2842__), .dout(new_new_n3333__));
  or1   g1149(.dina(new_new_n3333__), .dinb(new_new_n3332__), .dout(new_new_n3334__));
  and1  g1150(.dina(new_new_n2902__), .dinb(new_new_n2841__), .dout(new_new_n3335__));
  and1  g1151(.dina(new_new_n2903__), .dinb(new_new_n2840__), .dout(new_new_n3336__));
  or1   g1152(.dina(new_new_n3336__), .dinb(new_new_n3335__), .dout(new_new_n3337__));
  and1  g1153(.dina(new_new_n2900__), .dinb(new_new_n2829__), .dout(new_new_n3338__));
  and1  g1154(.dina(new_new_n2901__), .dinb(new_new_n2828__), .dout(new_new_n3339__));
  or1   g1155(.dina(new_new_n3339__), .dinb(new_new_n3338__), .dout(new_new_n3340__));
  or1   g1156(.dina(new_new_n3331__), .dinb(new_new_n3328__), .dout(new_new_n3341__));
  or1   g1157(.dina(new_new_n3341__), .dinb(new_new_n3334__), .dout(new_new_n3342__));
  or1   g1158(.dina(new_new_n3342__), .dinb(new_new_n3337__), .dout(new_new_n3343__));
  or1   g1159(.dina(new_new_n3343__), .dinb(new_new_n3340__), .dout(new_new_n3344__));
  and1  g1160(.dina(new_new_n2898__), .dinb(new_new_n2827__), .dout(new_new_n3345__));
  and1  g1161(.dina(new_new_n2899__), .dinb(new_new_n2826__), .dout(new_new_n3346__));
  or1   g1162(.dina(new_new_n3346__), .dinb(new_new_n3345__), .dout(new_new_n3347__));
  and1  g1163(.dina(new_new_n2890__), .dinb(new_new_n2839__), .dout(new_new_n3348__));
  and1  g1164(.dina(new_new_n2891__), .dinb(new_new_n2838__), .dout(new_new_n3349__));
  or1   g1165(.dina(new_new_n3349__), .dinb(new_new_n3348__), .dout(new_new_n3350__));
  and1  g1166(.dina(new_new_n2896__), .dinb(new_new_n2825__), .dout(new_new_n3351__));
  and1  g1167(.dina(new_new_n2897__), .dinb(new_new_n2824__), .dout(new_new_n3352__));
  or1   g1168(.dina(new_new_n3352__), .dinb(new_new_n3351__), .dout(new_new_n3353__));
  and1  g1169(.dina(new_new_n2888__), .dinb(new_new_n2823__), .dout(new_new_n3354__));
  and1  g1170(.dina(new_new_n2889__), .dinb(new_new_n2822__), .dout(new_new_n3355__));
  or1   g1171(.dina(new_new_n3355__), .dinb(new_new_n3354__), .dout(new_new_n3356__));
  and1  g1172(.dina(new_new_n2894__), .dinb(new_new_n2853__), .dout(new_new_n3357__));
  and1  g1173(.dina(new_new_n2895__), .dinb(new_new_n2852__), .dout(new_new_n3358__));
  or1   g1174(.dina(new_new_n3358__), .dinb(new_new_n3357__), .dout(new_new_n3359__));
  or1   g1175(.dina(new_new_n3350__), .dinb(new_new_n3347__), .dout(new_new_n3360__));
  or1   g1176(.dina(new_new_n3360__), .dinb(new_new_n3353__), .dout(new_new_n3361__));
  or1   g1177(.dina(new_new_n3361__), .dinb(new_new_n3356__), .dout(new_new_n3362__));
  or1   g1178(.dina(new_new_n3362__), .dinb(new_new_n3359__), .dout(new_new_n3363__));
  or1   g1179(.dina(new_new_n3363__), .dinb(new_new_n3344__), .dout(new_new_n3364__));
  or1   g1180(.dina(new_new_n2657__), .dinb(new_new_n2033__), .dout(new_new_n3365__));
  or1   g1181(.dina(new_new_n2584__), .dinb(new_new_n5083__), .dout(new_new_n3366__));
  and1  g1182(.dina(new_new_n3366__), .dinb(new_new_n3365__), .dout(new_new_n3367__));
  and1  g1183(.dina(new_new_n2918__), .dinb(new_new_n2837__), .dout(new_new_n3368__));
  and1  g1184(.dina(new_new_n2919__), .dinb(new_new_n2836__), .dout(new_new_n3369__));
  or1   g1185(.dina(new_new_n3369__), .dinb(new_new_n3368__), .dout(new_new_n3370__));
  or1   g1186(.dina(new_new_n3370__), .dinb(new_new_n3367__), .dout(new_new_n3371__));
  and1  g1187(.dina(new_new_n2916__), .dinb(new_new_n2835__), .dout(new_new_n3372__));
  and1  g1188(.dina(new_new_n2917__), .dinb(new_new_n2834__), .dout(new_new_n3373__));
  or1   g1189(.dina(new_new_n3373__), .dinb(new_new_n3372__), .dout(new_new_n3374__));
  and1  g1190(.dina(new_new_n2910__), .dinb(new_new_n2849__), .dout(new_new_n3375__));
  and1  g1191(.dina(new_new_n2911__), .dinb(new_new_n2848__), .dout(new_new_n3376__));
  or1   g1192(.dina(new_new_n3376__), .dinb(new_new_n3375__), .dout(new_new_n3377__));
  and1  g1193(.dina(new_new_n2914__), .dinb(new_new_n2833__), .dout(new_new_n3378__));
  and1  g1194(.dina(new_new_n2915__), .dinb(new_new_n2832__), .dout(new_new_n3379__));
  or1   g1195(.dina(new_new_n3379__), .dinb(new_new_n3378__), .dout(new_new_n3380__));
  and1  g1196(.dina(new_new_n2908__), .dinb(new_new_n2831__), .dout(new_new_n3381__));
  and1  g1197(.dina(new_new_n2909__), .dinb(new_new_n2830__), .dout(new_new_n3382__));
  or1   g1198(.dina(new_new_n3382__), .dinb(new_new_n3381__), .dout(new_new_n3383__));
  and1  g1199(.dina(new_new_n2912__), .dinb(new_new_n2847__), .dout(new_new_n3384__));
  and1  g1200(.dina(new_new_n2913__), .dinb(new_new_n2846__), .dout(new_new_n3385__));
  or1   g1201(.dina(new_new_n3385__), .dinb(new_new_n3384__), .dout(new_new_n3386__));
  or1   g1202(.dina(new_new_n3377__), .dinb(new_new_n3374__), .dout(new_new_n3387__));
  or1   g1203(.dina(new_new_n3387__), .dinb(new_new_n3380__), .dout(new_new_n3388__));
  or1   g1204(.dina(new_new_n3388__), .dinb(new_new_n3383__), .dout(new_new_n3389__));
  or1   g1205(.dina(new_new_n3389__), .dinb(new_new_n3386__), .dout(new_new_n3390__));
  or1   g1206(.dina(new_new_n3390__), .dinb(new_new_n3371__), .dout(new_new_n3391__));
  or1   g1207(.dina(new_new_n5074__), .dinb(new_new_n5085__), .dout(new_new_n3392__));
  or1   g1208(.dina(new_new_n5079__), .dinb(new_new_n5085__), .dout(new_new_n3393__));
  and1  g1209(.dina(new_new_n3393__), .dinb(new_new_n3392__), .dout(new_new_n3394__));
  or1   g1210(.dina(new_new_n3391__), .dinb(new_new_n3364__), .dout(new_new_n3395__));
  or1   g1211(.dina(new_new_n3395__), .dinb(new_new_n3394__), .dout(new_new_n3396__));
  and1  g1212(.dina(new_new_n5086__), .dinb(new_new_n5087__), .dout(new_new_n3397__));
  or1   g1213(.dina(new_new_n5088__), .dinb(new_new_n5089__), .dout(new_new_n3398__));
  and1  g1214(.dina(new_new_n5088__), .dinb(new_new_n5089__), .dout(new_new_n3399__));
  or1   g1215(.dina(new_new_n5086__), .dinb(new_new_n5087__), .dout(new_new_n3400__));
  and1  g1216(.dina(new_new_n3400__), .dinb(new_new_n3398__), .dout(new_new_n3401__));
  or1   g1217(.dina(new_new_n3399__), .dinb(new_new_n3397__), .dout(new_new_n3402__));
  and1  g1218(.dina(new_new_n3402__), .dinb(new_new_n2569__), .dout(new_new_n3403__));
  and1  g1219(.dina(new_new_n3401__), .dinb(new_new_n5091__), .dout(new_new_n3404__));
  or1   g1220(.dina(new_new_n3404__), .dinb(new_new_n3403__), .dout(new_new_n3405__));
  and1  g1221(.dina(new_new_n3405__), .dinb(new_new_n5065__), .dout(new_new_n3406__));
  and1  g1222(.dina(new_new_n5091__), .dinb(new_new_n5063__), .dout(new_new_n3407__));
  or1   g1223(.dina(new_new_n3407__), .dinb(new_new_n3406__), .dout(new_new_n3408__));
  or1   g1224(.dina(new_new_n2944__), .dinb(new_new_n2718__), .dout(new_new_n3409__));
  or1   g1225(.dina(new_new_n2939__), .dinb(new_new_n2725__), .dout(new_new_n3410__));
  and1  g1226(.dina(new_new_n3410__), .dinb(new_new_n3409__), .dout(new_new_n3411__));
  and1  g1227(.dina(new_new_n3411__), .dinb(new_new_n5092__), .dout(new_new_n3412__));
  or1   g1228(.dina(new_new_n5090__), .dinb(new_new_n5074__), .dout(new_new_n3413__));
  and1  g1229(.dina(new_new_n2935__), .dinb(new_new_n2712__), .dout(new_new_n3414__));
  or1   g1230(.dina(new_new_n2934__), .dinb(new_new_n2713__), .dout(new_new_n3415__));
  and1  g1231(.dina(new_new_n2933__), .dinb(new_new_n2714__), .dout(new_new_n3416__));
  or1   g1232(.dina(new_new_n2932__), .dinb(new_new_n2715__), .dout(new_new_n3417__));
  and1  g1233(.dina(new_new_n3417__), .dinb(new_new_n3415__), .dout(new_new_n3418__));
  or1   g1234(.dina(new_new_n3416__), .dinb(new_new_n3414__), .dout(new_new_n3419__));
  and1  g1235(.dina(new_new_n2883__), .dinb(new_new_n2876__), .dout(new_new_n3420__));
  or1   g1236(.dina(new_new_n2882__), .dinb(new_new_n2877__), .dout(new_new_n3421__));
  and1  g1237(.dina(new_new_n2875__), .dinb(new_new_n2873__), .dout(new_new_n3422__));
  or1   g1238(.dina(new_new_n2874__), .dinb(new_new_n2872__), .dout(new_new_n3423__));
  and1  g1239(.dina(new_new_n3422__), .dinb(new_new_n3420__), .dout(new_new_n3424__));
  or1   g1240(.dina(new_new_n3423__), .dinb(new_new_n3421__), .dout(new_new_n3425__));
  or1   g1241(.dina(new_new_n3425__), .dinb(new_new_n3418__), .dout(new_new_n3426__));
  or1   g1242(.dina(new_new_n3424__), .dinb(new_new_n3419__), .dout(new_new_n3427__));
  and1  g1243(.dina(new_new_n3427__), .dinb(new_new_n3426__), .dout(new_new_n3428__));
  or1   g1244(.dina(new_new_n3428__), .dinb(new_new_n5079__), .dout(new_new_n3429__));
  and1  g1245(.dina(new_new_n3429__), .dinb(new_new_n3413__), .dout(new_new_n3430__));
  or1   g1246(.dina(new_new_n2947__), .dinb(new_new_n2721__), .dout(new_new_n3431__));
  or1   g1247(.dina(new_new_n2940__), .dinb(new_new_n2726__), .dout(new_new_n3432__));
  and1  g1248(.dina(new_new_n3432__), .dinb(new_new_n3431__), .dout(new_new_n3433__));
  and1  g1249(.dina(new_new_n3433__), .dinb(new_new_n5092__), .dout(new_new_n3434__));
  and1  g1250(.dina(new_new_n5093__), .dinb(new_new_n2707__), .dout(new_new_n3435__));
  and1  g1251(.dina(new_new_n5093__), .dinb(new_new_n2705__), .dout(new_new_n3436__));
  or1   g1252(.dina(new_new_n3436__), .dinb(new_new_n3435__), .dout(new_new_n3437__));
  or1   g1253(.dina(new_new_n5094__), .dinb(new_new_n5095__), .dout(new_new_n3438__));
  or1   g1254(.dina(new_new_n3438__), .dinb(new_new_n5096__), .dout(new_new_n3439__));
  or1   g1255(.dina(new_new_n5097__), .dinb(new_new_n5098__), .dout(new_new_n3440__));
  or1   g1256(.dina(new_new_n3440__), .dinb(new_new_n5099__), .dout(new_new_n3441__));
  or1   g1257(.dina(new_new_n3441__), .dinb(new_new_n3439__), .dout(new_new_n3442__));
  or1   g1258(.dina(new_new_n3442__), .dinb(new_new_n5070__), .dout(new_new_n3443__));
  and1  g1259(.dina(new_new_n5100__), .dinb(new_new_n2359__), .dout(new_new_n3444__));
  or1   g1260(.dina(new_new_n5102__), .dinb(new_new_n2358__), .dout(new_new_n3445__));
  or1   g1261(.dina(new_new_n3174__), .dinb(new_new_n3150__), .dout(new_new_n3446__));
  or1   g1262(.dina(new_new_n3446__), .dinb(new_new_n3158__), .dout(new_new_n3447__));
  or1   g1263(.dina(new_new_n3447__), .dinb(new_new_n3154__), .dout(new_new_n3448__));
  or1   g1264(.dina(new_new_n3176__), .dinb(new_new_n3152__), .dout(new_new_n3449__));
  or1   g1265(.dina(new_new_n3449__), .dinb(new_new_n3160__), .dout(new_new_n3450__));
  or1   g1266(.dina(new_new_n3450__), .dinb(new_new_n3156__), .dout(new_new_n3451__));
  or1   g1267(.dina(new_new_n3218__), .dinb(new_new_n3164__), .dout(new_new_n3452__));
  or1   g1268(.dina(new_new_n3452__), .dinb(new_new_n3168__), .dout(new_new_n3453__));
  or1   g1269(.dina(new_new_n3453__), .dinb(new_new_n3166__), .dout(new_new_n3454__));
  and1  g1270(.dina(new_new_n3190__), .dinb(new_new_n5104__), .dout(new_new_n3455__));
  and1  g1271(.dina(new_new_n3455__), .dinb(new_new_n5105__), .dout(new_new_n3456__));
  and1  g1272(.dina(new_new_n3178__), .dinb(new_new_n5106__), .dout(new_new_n3457__));
  and1  g1273(.dina(new_new_n3457__), .dinb(new_new_n5105__), .dout(new_new_n3458__));
  and1  g1274(.dina(new_new_n3182__), .dinb(new_new_n5104__), .dout(new_new_n3459__));
  and1  g1275(.dina(new_new_n3459__), .dinb(new_new_n5107__), .dout(new_new_n3460__));
  and1  g1276(.dina(new_new_n3186__), .dinb(new_new_n5106__), .dout(new_new_n3461__));
  and1  g1277(.dina(new_new_n3461__), .dinb(new_new_n5107__), .dout(new_new_n3462__));
  or1   g1278(.dina(new_new_n3458__), .dinb(new_new_n3456__), .dout(new_new_n3463__));
  or1   g1279(.dina(new_new_n3463__), .dinb(new_new_n3460__), .dout(new_new_n3464__));
  or1   g1280(.dina(new_new_n3464__), .dinb(new_new_n3462__), .dout(new_new_n3465__));
  and1  g1281(.dina(new_new_n3206__), .dinb(new_new_n5110__), .dout(new_new_n3466__));
  and1  g1282(.dina(new_new_n3466__), .dinb(new_new_n5117__), .dout(new_new_n3467__));
  and1  g1283(.dina(new_new_n3194__), .dinb(new_new_n5124__), .dout(new_new_n3468__));
  and1  g1284(.dina(new_new_n3468__), .dinb(new_new_n5117__), .dout(new_new_n3469__));
  and1  g1285(.dina(new_new_n3202__), .dinb(new_new_n5110__), .dout(new_new_n3470__));
  and1  g1286(.dina(new_new_n3470__), .dinb(new_new_n5131__), .dout(new_new_n3471__));
  and1  g1287(.dina(new_new_n3198__), .dinb(new_new_n5124__), .dout(new_new_n3472__));
  and1  g1288(.dina(new_new_n3472__), .dinb(new_new_n5131__), .dout(new_new_n3473__));
  or1   g1289(.dina(new_new_n3469__), .dinb(new_new_n3467__), .dout(new_new_n3474__));
  or1   g1290(.dina(new_new_n3474__), .dinb(new_new_n3471__), .dout(new_new_n3475__));
  or1   g1291(.dina(new_new_n3475__), .dinb(new_new_n3473__), .dout(new_new_n3476__));
  and1  g1292(.dina(new_new_n3208__), .dinb(new_new_n5111__), .dout(new_new_n3477__));
  and1  g1293(.dina(new_new_n3477__), .dinb(new_new_n5118__), .dout(new_new_n3478__));
  and1  g1294(.dina(new_new_n3196__), .dinb(new_new_n5125__), .dout(new_new_n3479__));
  and1  g1295(.dina(new_new_n3479__), .dinb(new_new_n5118__), .dout(new_new_n3480__));
  and1  g1296(.dina(new_new_n3204__), .dinb(new_new_n5111__), .dout(new_new_n3481__));
  and1  g1297(.dina(new_new_n3481__), .dinb(new_new_n5132__), .dout(new_new_n3482__));
  and1  g1298(.dina(new_new_n3200__), .dinb(new_new_n5125__), .dout(new_new_n3483__));
  and1  g1299(.dina(new_new_n3483__), .dinb(new_new_n5132__), .dout(new_new_n3484__));
  or1   g1300(.dina(new_new_n3480__), .dinb(new_new_n3478__), .dout(new_new_n3485__));
  or1   g1301(.dina(new_new_n3485__), .dinb(new_new_n3482__), .dout(new_new_n3486__));
  or1   g1302(.dina(new_new_n3486__), .dinb(new_new_n3484__), .dout(new_new_n3487__));
  and1  g1303(.dina(new_new_n5139__), .dinb(new_new_n3192__), .dout(new_new_n3488__));
  or1   g1304(.dina(new_new_n5147__), .dinb(new_new_n3193__), .dout(new_new_n3489__));
  and1  g1305(.dina(new_new_n3488__), .dinb(new_new_n5153__), .dout(new_new_n3490__));
  or1   g1306(.dina(new_new_n3489__), .dinb(new_new_n5161__), .dout(new_new_n3491__));
  and1  g1307(.dina(new_new_n3180__), .dinb(new_new_n5167__), .dout(new_new_n3492__));
  or1   g1308(.dina(new_new_n3181__), .dinb(new_new_n5175__), .dout(new_new_n3493__));
  and1  g1309(.dina(new_new_n3492__), .dinb(new_new_n5153__), .dout(new_new_n3494__));
  or1   g1310(.dina(new_new_n3493__), .dinb(new_new_n5161__), .dout(new_new_n3495__));
  and1  g1311(.dina(new_new_n5139__), .dinb(new_new_n3184__), .dout(new_new_n3496__));
  or1   g1312(.dina(new_new_n5147__), .dinb(new_new_n3185__), .dout(new_new_n3497__));
  and1  g1313(.dina(new_new_n3496__), .dinb(new_new_n5181__), .dout(new_new_n3498__));
  or1   g1314(.dina(new_new_n3497__), .dinb(new_new_n5189__), .dout(new_new_n3499__));
  and1  g1315(.dina(new_new_n3188__), .dinb(new_new_n5167__), .dout(new_new_n3500__));
  or1   g1316(.dina(new_new_n3189__), .dinb(new_new_n5175__), .dout(new_new_n3501__));
  and1  g1317(.dina(new_new_n3500__), .dinb(new_new_n5181__), .dout(new_new_n3502__));
  or1   g1318(.dina(new_new_n3501__), .dinb(new_new_n5189__), .dout(new_new_n3503__));
  and1  g1319(.dina(new_new_n3495__), .dinb(new_new_n3491__), .dout(new_new_n3504__));
  or1   g1320(.dina(new_new_n3494__), .dinb(new_new_n3490__), .dout(new_new_n3505__));
  and1  g1321(.dina(new_new_n3504__), .dinb(new_new_n3499__), .dout(new_new_n3506__));
  or1   g1322(.dina(new_new_n3505__), .dinb(new_new_n3498__), .dout(new_new_n3507__));
  and1  g1323(.dina(new_new_n3506__), .dinb(new_new_n3503__), .dout(new_new_n3508__));
  or1   g1324(.dina(new_new_n3507__), .dinb(new_new_n3502__), .dout(new_new_n3509__));
  and1  g1325(.dina(new_new_n5140__), .dinb(new_new_n3130__), .dout(new_new_n3510__));
  or1   g1326(.dina(new_new_n5148__), .dinb(new_new_n3131__), .dout(new_new_n3511__));
  and1  g1327(.dina(new_new_n3510__), .dinb(new_new_n5154__), .dout(new_new_n3512__));
  or1   g1328(.dina(new_new_n3511__), .dinb(new_new_n5162__), .dout(new_new_n3513__));
  and1  g1329(.dina(new_new_n3118__), .dinb(new_new_n5168__), .dout(new_new_n3514__));
  or1   g1330(.dina(new_new_n3119__), .dinb(new_new_n5176__), .dout(new_new_n3515__));
  and1  g1331(.dina(new_new_n3514__), .dinb(new_new_n5154__), .dout(new_new_n3516__));
  or1   g1332(.dina(new_new_n3515__), .dinb(new_new_n5162__), .dout(new_new_n3517__));
  and1  g1333(.dina(new_new_n5140__), .dinb(new_new_n3122__), .dout(new_new_n3518__));
  or1   g1334(.dina(new_new_n5148__), .dinb(new_new_n3123__), .dout(new_new_n3519__));
  and1  g1335(.dina(new_new_n3518__), .dinb(new_new_n5182__), .dout(new_new_n3520__));
  or1   g1336(.dina(new_new_n3519__), .dinb(new_new_n5190__), .dout(new_new_n3521__));
  and1  g1337(.dina(new_new_n3126__), .dinb(new_new_n5168__), .dout(new_new_n3522__));
  or1   g1338(.dina(new_new_n3127__), .dinb(new_new_n5176__), .dout(new_new_n3523__));
  and1  g1339(.dina(new_new_n3522__), .dinb(new_new_n5182__), .dout(new_new_n3524__));
  or1   g1340(.dina(new_new_n3523__), .dinb(new_new_n5190__), .dout(new_new_n3525__));
  and1  g1341(.dina(new_new_n3517__), .dinb(new_new_n3513__), .dout(new_new_n3526__));
  or1   g1342(.dina(new_new_n3516__), .dinb(new_new_n3512__), .dout(new_new_n3527__));
  and1  g1343(.dina(new_new_n3526__), .dinb(new_new_n3521__), .dout(new_new_n3528__));
  or1   g1344(.dina(new_new_n3527__), .dinb(new_new_n3520__), .dout(new_new_n3529__));
  and1  g1345(.dina(new_new_n3528__), .dinb(new_new_n3525__), .dout(new_new_n3530__));
  or1   g1346(.dina(new_new_n3529__), .dinb(new_new_n3524__), .dout(new_new_n3531__));
  and1  g1347(.dina(new_new_n5141__), .dinb(new_new_n3132__), .dout(new_new_n3532__));
  or1   g1348(.dina(new_new_n5149__), .dinb(new_new_n3133__), .dout(new_new_n3533__));
  and1  g1349(.dina(new_new_n3532__), .dinb(new_new_n5155__), .dout(new_new_n3534__));
  or1   g1350(.dina(new_new_n3533__), .dinb(new_new_n5163__), .dout(new_new_n3535__));
  and1  g1351(.dina(new_new_n3120__), .dinb(new_new_n5169__), .dout(new_new_n3536__));
  or1   g1352(.dina(new_new_n3121__), .dinb(new_new_n5177__), .dout(new_new_n3537__));
  and1  g1353(.dina(new_new_n3536__), .dinb(new_new_n5155__), .dout(new_new_n3538__));
  or1   g1354(.dina(new_new_n3537__), .dinb(new_new_n5163__), .dout(new_new_n3539__));
  and1  g1355(.dina(new_new_n5141__), .dinb(new_new_n3124__), .dout(new_new_n3540__));
  or1   g1356(.dina(new_new_n5149__), .dinb(new_new_n3125__), .dout(new_new_n3541__));
  and1  g1357(.dina(new_new_n3540__), .dinb(new_new_n5183__), .dout(new_new_n3542__));
  or1   g1358(.dina(new_new_n3541__), .dinb(new_new_n5191__), .dout(new_new_n3543__));
  and1  g1359(.dina(new_new_n3128__), .dinb(new_new_n5169__), .dout(new_new_n3544__));
  or1   g1360(.dina(new_new_n3129__), .dinb(new_new_n5177__), .dout(new_new_n3545__));
  and1  g1361(.dina(new_new_n3544__), .dinb(new_new_n5183__), .dout(new_new_n3546__));
  or1   g1362(.dina(new_new_n3545__), .dinb(new_new_n5191__), .dout(new_new_n3547__));
  and1  g1363(.dina(new_new_n3539__), .dinb(new_new_n3535__), .dout(new_new_n3548__));
  or1   g1364(.dina(new_new_n3538__), .dinb(new_new_n3534__), .dout(new_new_n3549__));
  and1  g1365(.dina(new_new_n3548__), .dinb(new_new_n3543__), .dout(new_new_n3550__));
  or1   g1366(.dina(new_new_n3549__), .dinb(new_new_n3542__), .dout(new_new_n3551__));
  and1  g1367(.dina(new_new_n3550__), .dinb(new_new_n3547__), .dout(new_new_n3552__));
  or1   g1368(.dina(new_new_n3551__), .dinb(new_new_n3546__), .dout(new_new_n3553__));
  and1  g1369(.dina(new_new_n5195__), .dinb(new_new_n5202__), .dout(new_new_n3554__));
  or1   g1370(.dina(new_new_n5206__), .dinb(new_new_n5214__), .dout(new_new_n3555__));
  and1  g1371(.dina(new_new_n5206__), .dinb(new_new_n5216__), .dout(new_new_n3556__));
  or1   g1372(.dina(new_new_n5195__), .dinb(new_new_n5218__), .dout(new_new_n3557__));
  and1  g1373(.dina(new_new_n3557__), .dinb(new_new_n3555__), .dout(new_new_n3558__));
  or1   g1374(.dina(new_new_n3556__), .dinb(new_new_n3554__), .dout(new_new_n3559__));
  and1  g1375(.dina(new_new_n5223__), .dinb(new_new_n5202__), .dout(new_new_n3560__));
  or1   g1376(.dina(new_new_n5233__), .dinb(new_new_n5214__), .dout(new_new_n3561__));
  and1  g1377(.dina(new_new_n5233__), .dinb(new_new_n5216__), .dout(new_new_n3562__));
  or1   g1378(.dina(new_new_n5223__), .dinb(new_new_n5218__), .dout(new_new_n3563__));
  and1  g1379(.dina(new_new_n3563__), .dinb(new_new_n3561__), .dout(new_new_n3564__));
  or1   g1380(.dina(new_new_n3562__), .dinb(new_new_n3560__), .dout(new_new_n3565__));
  and1  g1381(.dina(new_new_n2775__), .dinb(new_new_n2742__), .dout(new_new_n3566__));
  or1   g1382(.dina(new_new_n3048__), .dinb(new_new_n3017__), .dout(new_new_n3567__));
  and1  g1383(.dina(new_new_n2773__), .dinb(new_new_n2748__), .dout(new_new_n3568__));
  and1  g1384(.dina(new_new_n3568__), .dinb(new_new_n5241__), .dout(new_new_n3569__));
  or1   g1385(.dina(new_new_n3046__), .dinb(new_new_n3023__), .dout(new_new_n3570__));
  and1  g1386(.dina(new_new_n2771__), .dinb(new_new_n2746__), .dout(new_new_n3571__));
  and1  g1387(.dina(new_new_n5244__), .dinb(new_new_n5241__), .dout(new_new_n3572__));
  and1  g1388(.dina(new_new_n3572__), .dinb(new_new_n3571__), .dout(new_new_n3573__));
  or1   g1389(.dina(new_new_n3044__), .dinb(new_new_n3021__), .dout(new_new_n3574__));
  and1  g1390(.dina(new_new_n2803__), .dinb(new_new_n2792__), .dout(new_new_n3575__));
  and1  g1391(.dina(new_new_n5245__), .dinb(new_new_n5242__), .dout(new_new_n3576__));
  and1  g1392(.dina(new_new_n3576__), .dinb(new_new_n3575__), .dout(new_new_n3577__));
  and1  g1393(.dina(new_new_n3577__), .dinb(new_new_n5244__), .dout(new_new_n3578__));
  or1   g1394(.dina(new_new_n3569__), .dinb(new_new_n3566__), .dout(new_new_n3579__));
  or1   g1395(.dina(new_new_n3579__), .dinb(new_new_n3573__), .dout(new_new_n3580__));
  or1   g1396(.dina(new_new_n3580__), .dinb(new_new_n3578__), .dout(new_new_n3581__));
  and1  g1397(.dina(new_new_n2765__), .dinb(new_new_n2734__), .dout(new_new_n3582__));
  or1   g1398(.dina(new_new_n2764__), .dinb(new_new_n2735__), .dout(new_new_n3583__));
  and1  g1399(.dina(new_new_n3039__), .dinb(new_new_n3008__), .dout(new_new_n3584__));
  or1   g1400(.dina(new_new_n3038__), .dinb(new_new_n3009__), .dout(new_new_n3585__));
  and1  g1401(.dina(new_new_n2763__), .dinb(new_new_n2732__), .dout(new_new_n3586__));
  or1   g1402(.dina(new_new_n2762__), .dinb(new_new_n2733__), .dout(new_new_n3587__));
  and1  g1403(.dina(new_new_n3586__), .dinb(new_new_n5248__), .dout(new_new_n3588__));
  or1   g1404(.dina(new_new_n3587__), .dinb(new_new_n5252__), .dout(new_new_n3589__));
  and1  g1405(.dina(new_new_n3037__), .dinb(new_new_n3006__), .dout(new_new_n3590__));
  or1   g1406(.dina(new_new_n3036__), .dinb(new_new_n3007__), .dout(new_new_n3591__));
  and1  g1407(.dina(new_new_n2787__), .dinb(new_new_n2756__), .dout(new_new_n3592__));
  or1   g1408(.dina(new_new_n2786__), .dinb(new_new_n2757__), .dout(new_new_n3593__));
  and1  g1409(.dina(new_new_n5255__), .dinb(new_new_n5248__), .dout(new_new_n3594__));
  or1   g1410(.dina(new_new_n5258__), .dinb(new_new_n5252__), .dout(new_new_n3595__));
  and1  g1411(.dina(new_new_n3594__), .dinb(new_new_n3592__), .dout(new_new_n3596__));
  or1   g1412(.dina(new_new_n3595__), .dinb(new_new_n3593__), .dout(new_new_n3597__));
  and1  g1413(.dina(new_new_n3063__), .dinb(new_new_n3030__), .dout(new_new_n3598__));
  or1   g1414(.dina(new_new_n3062__), .dinb(new_new_n3031__), .dout(new_new_n3599__));
  and1  g1415(.dina(new_new_n2785__), .dinb(new_new_n2754__), .dout(new_new_n3600__));
  or1   g1416(.dina(new_new_n2784__), .dinb(new_new_n2755__), .dout(new_new_n3601__));
  and1  g1417(.dina(new_new_n5261__), .dinb(new_new_n5247__), .dout(new_new_n3602__));
  or1   g1418(.dina(new_new_n5263__), .dinb(new_new_n5251__), .dout(new_new_n3603__));
  and1  g1419(.dina(new_new_n3602__), .dinb(new_new_n3600__), .dout(new_new_n3604__));
  or1   g1420(.dina(new_new_n3603__), .dinb(new_new_n3601__), .dout(new_new_n3605__));
  and1  g1421(.dina(new_new_n3604__), .dinb(new_new_n5255__), .dout(new_new_n3606__));
  or1   g1422(.dina(new_new_n3605__), .dinb(new_new_n5258__), .dout(new_new_n3607__));
  and1  g1423(.dina(new_new_n3061__), .dinb(new_new_n3028__), .dout(new_new_n3608__));
  or1   g1424(.dina(new_new_n3060__), .dinb(new_new_n3029__), .dout(new_new_n3609__));
  and1  g1425(.dina(new_new_n5264__), .dinb(new_new_n2731__), .dout(new_new_n3610__));
  or1   g1426(.dina(new_new_n5265__), .dinb(new_new_n2730__), .dout(new_new_n3611__));
  and1  g1427(.dina(new_new_n5266__), .dinb(new_new_n5261__), .dout(new_new_n3612__));
  or1   g1428(.dina(new_new_n5267__), .dinb(new_new_n5263__), .dout(new_new_n3613__));
  and1  g1429(.dina(new_new_n3612__), .dinb(new_new_n5249__), .dout(new_new_n3614__));
  or1   g1430(.dina(new_new_n3613__), .dinb(new_new_n5253__), .dout(new_new_n3615__));
  and1  g1431(.dina(new_new_n3614__), .dinb(new_new_n3610__), .dout(new_new_n3616__));
  or1   g1432(.dina(new_new_n3615__), .dinb(new_new_n3611__), .dout(new_new_n3617__));
  and1  g1433(.dina(new_new_n3616__), .dinb(new_new_n5256__), .dout(new_new_n3618__));
  or1   g1434(.dina(new_new_n3617__), .dinb(new_new_n5259__), .dout(new_new_n3619__));
  and1  g1435(.dina(new_new_n3589__), .dinb(new_new_n3583__), .dout(new_new_n3620__));
  or1   g1436(.dina(new_new_n3588__), .dinb(new_new_n3582__), .dout(new_new_n3621__));
  and1  g1437(.dina(new_new_n3620__), .dinb(new_new_n3597__), .dout(new_new_n3622__));
  or1   g1438(.dina(new_new_n3621__), .dinb(new_new_n3596__), .dout(new_new_n3623__));
  and1  g1439(.dina(new_new_n3622__), .dinb(new_new_n3607__), .dout(new_new_n3624__));
  or1   g1440(.dina(new_new_n3623__), .dinb(new_new_n3606__), .dout(new_new_n3625__));
  and1  g1441(.dina(new_new_n3624__), .dinb(new_new_n3619__), .dout(new_new_n3626__));
  or1   g1442(.dina(new_new_n3625__), .dinb(new_new_n3618__), .dout(new_new_n3627__));
  and1  g1443(.dina(new_new_n3056__), .dinb(new_new_n3005__), .dout(new_new_n3628__));
  or1   g1444(.dina(new_new_n3057__), .dinb(new_new_n3004__), .dout(new_new_n3629__));
  and1  g1445(.dina(new_new_n3629__), .dinb(new_new_n5256__), .dout(new_new_n3630__));
  or1   g1446(.dina(new_new_n3628__), .dinb(new_new_n5259__), .dout(new_new_n3631__));
  and1  g1447(.dina(new_new_n3630__), .dinb(new_new_n5260__), .dout(new_new_n3632__));
  or1   g1448(.dina(new_new_n3631__), .dinb(new_new_n5262__), .dout(new_new_n3633__));
  and1  g1449(.dina(new_new_n3632__), .dinb(new_new_n5249__), .dout(new_new_n3634__));
  or1   g1450(.dina(new_new_n3633__), .dinb(new_new_n5253__), .dout(new_new_n3635__));
  and1  g1451(.dina(new_new_n3634__), .dinb(new_new_n5266__), .dout(new_new_n3636__));
  or1   g1452(.dina(new_new_n3635__), .dinb(new_new_n5267__), .dout(new_new_n3637__));
  and1  g1453(.dina(new_new_n5269__), .dinb(new_new_n2683__), .dout(new_new_n3638__));
  or1   g1454(.dina(new_new_n5271__), .dinb(new_new_n2682__), .dout(new_new_n3639__));
  and1  g1455(.dina(new_new_n5272__), .dinb(new_new_n2993__), .dout(new_new_n3640__));
  or1   g1456(.dina(new_new_n5273__), .dinb(new_new_n2992__), .dout(new_new_n3641__));
  and1  g1457(.dina(new_new_n5272__), .dinb(new_new_n3088__), .dout(new_new_n3642__));
  or1   g1458(.dina(new_new_n5273__), .dinb(new_new_n3089__), .dout(new_new_n3643__));
  and1  g1459(.dina(new_new_n3642__), .dinb(new_new_n3099__), .dout(new_new_n3644__));
  or1   g1460(.dina(new_new_n3643__), .dinb(new_new_n3098__), .dout(new_new_n3645__));
  and1  g1461(.dina(new_new_n3641__), .dinb(new_new_n3639__), .dout(new_new_n3646__));
  or1   g1462(.dina(new_new_n3640__), .dinb(new_new_n3638__), .dout(new_new_n3647__));
  and1  g1463(.dina(new_new_n3646__), .dinb(new_new_n3645__), .dout(new_new_n3648__));
  or1   g1464(.dina(new_new_n3647__), .dinb(new_new_n3644__), .dout(new_new_n3649__));
  and1  g1465(.dina(new_new_n3649__), .dinb(new_new_n3636__), .dout(new_new_n3650__));
  or1   g1466(.dina(new_new_n3648__), .dinb(new_new_n3637__), .dout(new_new_n3651__));
  and1  g1467(.dina(new_new_n3651__), .dinb(new_new_n3626__), .dout(new_new_n3652__));
  or1   g1468(.dina(new_new_n3650__), .dinb(new_new_n3627__), .dout(new_new_n3653__));
  and1  g1469(.dina(new_new_n3652__), .dinb(new_new_n5274__), .dout(new_new_n3654__));
  and1  g1470(.dina(new_new_n3102__), .dinb(new_new_n2960__), .dout(new_new_n3655__));
  and1  g1471(.dina(new_new_n3113__), .dinb(new_new_n2951__), .dout(new_new_n3656__));
  or1   g1472(.dina(new_new_n3656__), .dinb(new_new_n3655__), .dout(new_new_n3657__));
  and1  g1473(.dina(new_new_n3657__), .dinb(new_new_n5243__), .dout(new_new_n3658__));
  and1  g1474(.dina(new_new_n3658__), .dinb(new_new_n5245__), .dout(new_new_n3659__));
  and1  g1475(.dina(new_new_n3659__), .dinb(new_new_n5242__), .dout(new_new_n3660__));
  or1   g1476(.dina(new_new_n3660__), .dinb(new_new_n5274__), .dout(new_new_n3661__));
  and1  g1477(.dina(new_new_n3661__), .dinb(new_new_n3653__), .dout(new_new_n3662__));
  or1   g1478(.dina(new_new_n3662__), .dinb(new_new_n3654__), .dout(new_new_n3663__));
  and1  g1479(.dina(new_new_n2781__), .dinb(new_new_n2744__), .dout(new_new_n3664__));
  or1   g1480(.dina(new_new_n3054__), .dinb(new_new_n3019__), .dout(new_new_n3665__));
  and1  g1481(.dina(new_new_n2779__), .dinb(new_new_n2752__), .dout(new_new_n3666__));
  and1  g1482(.dina(new_new_n3666__), .dinb(new_new_n5276__), .dout(new_new_n3667__));
  or1   g1483(.dina(new_new_n3052__), .dinb(new_new_n3027__), .dout(new_new_n3668__));
  and1  g1484(.dina(new_new_n2777__), .dinb(new_new_n2750__), .dout(new_new_n3669__));
  and1  g1485(.dina(new_new_n5279__), .dinb(new_new_n5276__), .dout(new_new_n3670__));
  and1  g1486(.dina(new_new_n3670__), .dinb(new_new_n3669__), .dout(new_new_n3671__));
  or1   g1487(.dina(new_new_n3050__), .dinb(new_new_n3025__), .dout(new_new_n3672__));
  and1  g1488(.dina(new_new_n2805__), .dinb(new_new_n2794__), .dout(new_new_n3673__));
  and1  g1489(.dina(new_new_n5280__), .dinb(new_new_n5277__), .dout(new_new_n3674__));
  and1  g1490(.dina(new_new_n3674__), .dinb(new_new_n3673__), .dout(new_new_n3675__));
  and1  g1491(.dina(new_new_n3675__), .dinb(new_new_n5279__), .dout(new_new_n3676__));
  or1   g1492(.dina(new_new_n3667__), .dinb(new_new_n3664__), .dout(new_new_n3677__));
  or1   g1493(.dina(new_new_n3677__), .dinb(new_new_n3671__), .dout(new_new_n3678__));
  or1   g1494(.dina(new_new_n3678__), .dinb(new_new_n3676__), .dout(new_new_n3679__));
  and1  g1495(.dina(new_new_n2769__), .dinb(new_new_n2740__), .dout(new_new_n3680__));
  or1   g1496(.dina(new_new_n2768__), .dinb(new_new_n2741__), .dout(new_new_n3681__));
  and1  g1497(.dina(new_new_n3043__), .dinb(new_new_n3014__), .dout(new_new_n3682__));
  or1   g1498(.dina(new_new_n3042__), .dinb(new_new_n3015__), .dout(new_new_n3683__));
  and1  g1499(.dina(new_new_n2767__), .dinb(new_new_n2738__), .dout(new_new_n3684__));
  or1   g1500(.dina(new_new_n2766__), .dinb(new_new_n2739__), .dout(new_new_n3685__));
  and1  g1501(.dina(new_new_n3684__), .dinb(new_new_n5283__), .dout(new_new_n3686__));
  or1   g1502(.dina(new_new_n3685__), .dinb(new_new_n5287__), .dout(new_new_n3687__));
  and1  g1503(.dina(new_new_n3041__), .dinb(new_new_n3012__), .dout(new_new_n3688__));
  or1   g1504(.dina(new_new_n3040__), .dinb(new_new_n3013__), .dout(new_new_n3689__));
  and1  g1505(.dina(new_new_n2791__), .dinb(new_new_n2760__), .dout(new_new_n3690__));
  or1   g1506(.dina(new_new_n2790__), .dinb(new_new_n2761__), .dout(new_new_n3691__));
  and1  g1507(.dina(new_new_n5290__), .dinb(new_new_n5283__), .dout(new_new_n3692__));
  or1   g1508(.dina(new_new_n5293__), .dinb(new_new_n5287__), .dout(new_new_n3693__));
  and1  g1509(.dina(new_new_n3692__), .dinb(new_new_n3690__), .dout(new_new_n3694__));
  or1   g1510(.dina(new_new_n3693__), .dinb(new_new_n3691__), .dout(new_new_n3695__));
  and1  g1511(.dina(new_new_n3067__), .dinb(new_new_n3034__), .dout(new_new_n3696__));
  or1   g1512(.dina(new_new_n3066__), .dinb(new_new_n3035__), .dout(new_new_n3697__));
  and1  g1513(.dina(new_new_n2789__), .dinb(new_new_n2758__), .dout(new_new_n3698__));
  or1   g1514(.dina(new_new_n2788__), .dinb(new_new_n2759__), .dout(new_new_n3699__));
  and1  g1515(.dina(new_new_n5296__), .dinb(new_new_n5282__), .dout(new_new_n3700__));
  or1   g1516(.dina(new_new_n5298__), .dinb(new_new_n5286__), .dout(new_new_n3701__));
  and1  g1517(.dina(new_new_n3700__), .dinb(new_new_n3698__), .dout(new_new_n3702__));
  or1   g1518(.dina(new_new_n3701__), .dinb(new_new_n3699__), .dout(new_new_n3703__));
  and1  g1519(.dina(new_new_n3702__), .dinb(new_new_n5290__), .dout(new_new_n3704__));
  or1   g1520(.dina(new_new_n3703__), .dinb(new_new_n5293__), .dout(new_new_n3705__));
  and1  g1521(.dina(new_new_n3065__), .dinb(new_new_n3032__), .dout(new_new_n3706__));
  or1   g1522(.dina(new_new_n3064__), .dinb(new_new_n3033__), .dout(new_new_n3707__));
  and1  g1523(.dina(new_new_n5264__), .dinb(new_new_n2737__), .dout(new_new_n3708__));
  or1   g1524(.dina(new_new_n5265__), .dinb(new_new_n2736__), .dout(new_new_n3709__));
  and1  g1525(.dina(new_new_n5299__), .dinb(new_new_n5296__), .dout(new_new_n3710__));
  or1   g1526(.dina(new_new_n5300__), .dinb(new_new_n5298__), .dout(new_new_n3711__));
  and1  g1527(.dina(new_new_n3710__), .dinb(new_new_n5284__), .dout(new_new_n3712__));
  or1   g1528(.dina(new_new_n3711__), .dinb(new_new_n5288__), .dout(new_new_n3713__));
  and1  g1529(.dina(new_new_n3712__), .dinb(new_new_n3708__), .dout(new_new_n3714__));
  or1   g1530(.dina(new_new_n3713__), .dinb(new_new_n3709__), .dout(new_new_n3715__));
  and1  g1531(.dina(new_new_n3714__), .dinb(new_new_n5291__), .dout(new_new_n3716__));
  or1   g1532(.dina(new_new_n3715__), .dinb(new_new_n5294__), .dout(new_new_n3717__));
  and1  g1533(.dina(new_new_n3687__), .dinb(new_new_n3681__), .dout(new_new_n3718__));
  or1   g1534(.dina(new_new_n3686__), .dinb(new_new_n3680__), .dout(new_new_n3719__));
  and1  g1535(.dina(new_new_n3718__), .dinb(new_new_n3695__), .dout(new_new_n3720__));
  or1   g1536(.dina(new_new_n3719__), .dinb(new_new_n3694__), .dout(new_new_n3721__));
  and1  g1537(.dina(new_new_n3720__), .dinb(new_new_n3705__), .dout(new_new_n3722__));
  or1   g1538(.dina(new_new_n3721__), .dinb(new_new_n3704__), .dout(new_new_n3723__));
  and1  g1539(.dina(new_new_n3722__), .dinb(new_new_n3717__), .dout(new_new_n3724__));
  or1   g1540(.dina(new_new_n3723__), .dinb(new_new_n3716__), .dout(new_new_n3725__));
  and1  g1541(.dina(new_new_n3058__), .dinb(new_new_n3011__), .dout(new_new_n3726__));
  or1   g1542(.dina(new_new_n3059__), .dinb(new_new_n3010__), .dout(new_new_n3727__));
  and1  g1543(.dina(new_new_n3727__), .dinb(new_new_n5291__), .dout(new_new_n3728__));
  or1   g1544(.dina(new_new_n3726__), .dinb(new_new_n5294__), .dout(new_new_n3729__));
  and1  g1545(.dina(new_new_n3728__), .dinb(new_new_n5295__), .dout(new_new_n3730__));
  or1   g1546(.dina(new_new_n3729__), .dinb(new_new_n5297__), .dout(new_new_n3731__));
  and1  g1547(.dina(new_new_n3730__), .dinb(new_new_n5284__), .dout(new_new_n3732__));
  or1   g1548(.dina(new_new_n3731__), .dinb(new_new_n5288__), .dout(new_new_n3733__));
  and1  g1549(.dina(new_new_n3732__), .dinb(new_new_n5299__), .dout(new_new_n3734__));
  or1   g1550(.dina(new_new_n3733__), .dinb(new_new_n5300__), .dout(new_new_n3735__));
  and1  g1551(.dina(new_new_n5269__), .dinb(new_new_n2685__), .dout(new_new_n3736__));
  or1   g1552(.dina(new_new_n5271__), .dinb(new_new_n2684__), .dout(new_new_n3737__));
  and1  g1553(.dina(new_new_n5301__), .dinb(new_new_n2995__), .dout(new_new_n3738__));
  or1   g1554(.dina(new_new_n5302__), .dinb(new_new_n2994__), .dout(new_new_n3739__));
  and1  g1555(.dina(new_new_n5301__), .dinb(new_new_n3092__), .dout(new_new_n3740__));
  or1   g1556(.dina(new_new_n5302__), .dinb(new_new_n3093__), .dout(new_new_n3741__));
  and1  g1557(.dina(new_new_n3740__), .dinb(new_new_n3101__), .dout(new_new_n3742__));
  or1   g1558(.dina(new_new_n3741__), .dinb(new_new_n3100__), .dout(new_new_n3743__));
  and1  g1559(.dina(new_new_n3739__), .dinb(new_new_n3737__), .dout(new_new_n3744__));
  or1   g1560(.dina(new_new_n3738__), .dinb(new_new_n3736__), .dout(new_new_n3745__));
  and1  g1561(.dina(new_new_n3744__), .dinb(new_new_n3743__), .dout(new_new_n3746__));
  or1   g1562(.dina(new_new_n3745__), .dinb(new_new_n3742__), .dout(new_new_n3747__));
  and1  g1563(.dina(new_new_n3747__), .dinb(new_new_n3734__), .dout(new_new_n3748__));
  or1   g1564(.dina(new_new_n3746__), .dinb(new_new_n3735__), .dout(new_new_n3749__));
  and1  g1565(.dina(new_new_n3749__), .dinb(new_new_n3724__), .dout(new_new_n3750__));
  or1   g1566(.dina(new_new_n3748__), .dinb(new_new_n3725__), .dout(new_new_n3751__));
  and1  g1567(.dina(new_new_n3750__), .dinb(new_new_n5303__), .dout(new_new_n3752__));
  and1  g1568(.dina(new_new_n3104__), .dinb(new_new_n2962__), .dout(new_new_n3753__));
  and1  g1569(.dina(new_new_n3115__), .dinb(new_new_n2953__), .dout(new_new_n3754__));
  or1   g1570(.dina(new_new_n3754__), .dinb(new_new_n3753__), .dout(new_new_n3755__));
  and1  g1571(.dina(new_new_n3755__), .dinb(new_new_n5278__), .dout(new_new_n3756__));
  and1  g1572(.dina(new_new_n3756__), .dinb(new_new_n5280__), .dout(new_new_n3757__));
  and1  g1573(.dina(new_new_n3757__), .dinb(new_new_n5277__), .dout(new_new_n3758__));
  or1   g1574(.dina(new_new_n3758__), .dinb(new_new_n5303__), .dout(new_new_n3759__));
  and1  g1575(.dina(new_new_n3759__), .dinb(new_new_n3751__), .dout(new_new_n3760__));
  or1   g1576(.dina(new_new_n3760__), .dinb(new_new_n3752__), .dout(new_new_n3761__));
  and1  g1577(.dina(new_new_n2654__), .dinb(new_new_n2619__), .dout(new_new_n3762__));
  and1  g1578(.dina(new_new_n2655__), .dinb(new_new_n2618__), .dout(new_new_n3763__));
  or1   g1579(.dina(new_new_n3763__), .dinb(new_new_n3762__), .dout(new_new_n3764__));
  and1  g1580(.dina(new_new_n2622__), .dinb(new_new_n2621__), .dout(new_new_n3765__));
  and1  g1581(.dina(new_new_n2623__), .dinb(new_new_n2620__), .dout(new_new_n3766__));
  or1   g1582(.dina(new_new_n3766__), .dinb(new_new_n3765__), .dout(new_new_n3767__));
  and1  g1583(.dina(new_new_n5304__), .dinb(new_new_n5305__), .dout(new_new_n3768__));
  or1   g1584(.dina(new_new_n5306__), .dinb(new_new_n5307__), .dout(new_new_n3769__));
  and1  g1585(.dina(new_new_n5306__), .dinb(new_new_n5307__), .dout(new_new_n3770__));
  or1   g1586(.dina(new_new_n5304__), .dinb(new_new_n5305__), .dout(new_new_n3771__));
  and1  g1587(.dina(new_new_n3771__), .dinb(new_new_n3769__), .dout(new_new_n3772__));
  or1   g1588(.dina(new_new_n3770__), .dinb(new_new_n3768__), .dout(new_new_n3773__));
  and1  g1589(.dina(new_new_n5308__), .dinb(new_new_n5309__), .dout(new_new_n3774__));
  or1   g1590(.dina(new_new_n5310__), .dinb(new_new_n5311__), .dout(new_new_n3775__));
  and1  g1591(.dina(new_new_n5310__), .dinb(new_new_n5311__), .dout(new_new_n3776__));
  or1   g1592(.dina(new_new_n5308__), .dinb(new_new_n5309__), .dout(new_new_n3777__));
  and1  g1593(.dina(new_new_n3777__), .dinb(new_new_n3775__), .dout(new_new_n3778__));
  or1   g1594(.dina(new_new_n3776__), .dinb(new_new_n3774__), .dout(new_new_n3779__));
  and1  g1595(.dina(new_new_n5312__), .dinb(new_new_n5313__), .dout(new_new_n3780__));
  or1   g1596(.dina(new_new_n5314__), .dinb(new_new_n5315__), .dout(new_new_n3781__));
  and1  g1597(.dina(new_new_n5314__), .dinb(new_new_n5315__), .dout(new_new_n3782__));
  or1   g1598(.dina(new_new_n5312__), .dinb(new_new_n5313__), .dout(new_new_n3783__));
  and1  g1599(.dina(new_new_n3783__), .dinb(new_new_n3781__), .dout(new_new_n3784__));
  or1   g1600(.dina(new_new_n3782__), .dinb(new_new_n3780__), .dout(new_new_n3785__));
  and1  g1601(.dina(new_new_n5316__), .dinb(new_new_n5317__), .dout(new_new_n3786__));
  or1   g1602(.dina(new_new_n5318__), .dinb(new_new_n5319__), .dout(new_new_n3787__));
  and1  g1603(.dina(new_new_n5318__), .dinb(new_new_n5319__), .dout(new_new_n3788__));
  or1   g1604(.dina(new_new_n5316__), .dinb(new_new_n5317__), .dout(new_new_n3789__));
  and1  g1605(.dina(new_new_n3789__), .dinb(new_new_n3787__), .dout(new_new_n3790__));
  or1   g1606(.dina(new_new_n3788__), .dinb(new_new_n3786__), .dout(new_new_n3791__));
  and1  g1607(.dina(new_new_n3790__), .dinb(new_new_n3785__), .dout(new_new_n3792__));
  and1  g1608(.dina(new_new_n3791__), .dinb(new_new_n3784__), .dout(new_new_n3793__));
  or1   g1609(.dina(new_new_n3793__), .dinb(new_new_n3792__), .dout(new_new_n3794__));
  and1  g1610(.dina(new_new_n5321__), .dinb(new_new_n5323__), .dout(new_new_n3795__));
  or1   g1611(.dina(new_new_n5324__), .dinb(new_new_n5326__), .dout(new_new_n3796__));
  and1  g1612(.dina(new_new_n5324__), .dinb(new_new_n5326__), .dout(new_new_n3797__));
  or1   g1613(.dina(new_new_n5321__), .dinb(new_new_n5323__), .dout(new_new_n3798__));
  and1  g1614(.dina(new_new_n3798__), .dinb(new_new_n3796__), .dout(new_new_n3799__));
  or1   g1615(.dina(new_new_n3797__), .dinb(new_new_n3795__), .dout(new_new_n3800__));
  and1  g1616(.dina(new_new_n5328__), .dinb(new_new_n5329__), .dout(new_new_n3801__));
  or1   g1617(.dina(new_new_n5331__), .dinb(new_new_n5333__), .dout(new_new_n3802__));
  and1  g1618(.dina(new_new_n5331__), .dinb(new_new_n5333__), .dout(new_new_n3803__));
  or1   g1619(.dina(new_new_n5328__), .dinb(new_new_n5329__), .dout(new_new_n3804__));
  and1  g1620(.dina(new_new_n3804__), .dinb(new_new_n3802__), .dout(new_new_n3805__));
  or1   g1621(.dina(new_new_n3803__), .dinb(new_new_n3801__), .dout(new_new_n3806__));
  or1   g1622(.dina(new_new_n3806__), .dinb(new_new_n3799__), .dout(new_new_n3807__));
  or1   g1623(.dina(new_new_n3805__), .dinb(new_new_n3800__), .dout(new_new_n3808__));
  and1  g1624(.dina(new_new_n3808__), .dinb(new_new_n3807__), .dout(new_new_n3809__));
  and1  g1625(.dina(new_new_n3778__), .dinb(new_new_n5335__), .dout(new_new_n3810__));
  and1  g1626(.dina(new_new_n5337__), .dinb(new_new_n3772__), .dout(new_new_n3811__));
  or1   g1627(.dina(new_new_n3811__), .dinb(new_new_n3810__), .dout(new_new_n3812__));
  and1  g1628(.dina(new_new_n5338__), .dinb(new_new_n5339__), .dout(new_new_n3813__));
  or1   g1629(.dina(new_new_n5340__), .dinb(new_new_n5341__), .dout(new_new_n3814__));
  and1  g1630(.dina(new_new_n5340__), .dinb(new_new_n5341__), .dout(new_new_n3815__));
  or1   g1631(.dina(new_new_n5338__), .dinb(new_new_n5339__), .dout(new_new_n3816__));
  and1  g1632(.dina(new_new_n3816__), .dinb(new_new_n3814__), .dout(new_new_n3817__));
  or1   g1633(.dina(new_new_n3815__), .dinb(new_new_n3813__), .dout(new_new_n3818__));
  and1  g1634(.dina(new_new_n5342__), .dinb(new_new_n5343__), .dout(new_new_n3819__));
  or1   g1635(.dina(new_new_n5344__), .dinb(new_new_n5345__), .dout(new_new_n3820__));
  and1  g1636(.dina(new_new_n5344__), .dinb(new_new_n5345__), .dout(new_new_n3821__));
  or1   g1637(.dina(new_new_n5342__), .dinb(new_new_n5343__), .dout(new_new_n3822__));
  and1  g1638(.dina(new_new_n3822__), .dinb(new_new_n3820__), .dout(new_new_n3823__));
  or1   g1639(.dina(new_new_n3821__), .dinb(new_new_n3819__), .dout(new_new_n3824__));
  and1  g1640(.dina(new_new_n3069__), .dinb(new_new_n2820__), .dout(new_new_n3825__));
  or1   g1641(.dina(new_new_n3068__), .dinb(new_new_n2821__), .dout(new_new_n3826__));
  and1  g1642(.dina(new_new_n3071__), .dinb(new_new_n2818__), .dout(new_new_n3827__));
  or1   g1643(.dina(new_new_n3070__), .dinb(new_new_n2819__), .dout(new_new_n3828__));
  and1  g1644(.dina(new_new_n3828__), .dinb(new_new_n3826__), .dout(new_new_n3829__));
  or1   g1645(.dina(new_new_n3827__), .dinb(new_new_n3825__), .dout(new_new_n3830__));
  or1   g1646(.dina(new_new_n5346__), .dinb(new_new_n5347__), .dout(new_new_n3831__));
  or1   g1647(.dina(new_new_n3831__), .dinb(new_new_n5348__), .dout(new_new_n3832__));
  or1   g1648(.dina(new_new_n5346__), .dinb(new_new_n5349__), .dout(new_new_n3833__));
  or1   g1649(.dina(new_new_n3833__), .dinb(new_new_n5350__), .dout(new_new_n3834__));
  and1  g1650(.dina(new_new_n3834__), .dinb(new_new_n3832__), .dout(new_new_n3835__));
  or1   g1651(.dina(new_new_n5351__), .dinb(new_new_n5349__), .dout(new_new_n3836__));
  or1   g1652(.dina(new_new_n3836__), .dinb(new_new_n5348__), .dout(new_new_n3837__));
  or1   g1653(.dina(new_new_n5351__), .dinb(new_new_n5347__), .dout(new_new_n3838__));
  or1   g1654(.dina(new_new_n3838__), .dinb(new_new_n5350__), .dout(new_new_n3839__));
  and1  g1655(.dina(new_new_n3839__), .dinb(new_new_n3837__), .dout(new_new_n3840__));
  and1  g1656(.dina(new_new_n3840__), .dinb(new_new_n3835__), .dout(new_new_n3841__));
  and1  g1657(.dina(new_new_n5352__), .dinb(new_new_n5353__), .dout(new_new_n3842__));
  or1   g1658(.dina(new_new_n5354__), .dinb(new_new_n5355__), .dout(new_new_n3843__));
  and1  g1659(.dina(new_new_n5354__), .dinb(new_new_n5355__), .dout(new_new_n3844__));
  or1   g1660(.dina(new_new_n5352__), .dinb(new_new_n5353__), .dout(new_new_n3845__));
  and1  g1661(.dina(new_new_n3845__), .dinb(new_new_n3843__), .dout(new_new_n3846__));
  or1   g1662(.dina(new_new_n3844__), .dinb(new_new_n3842__), .dout(new_new_n3847__));
  and1  g1663(.dina(new_new_n5356__), .dinb(new_new_n5357__), .dout(new_new_n3848__));
  or1   g1664(.dina(new_new_n5358__), .dinb(new_new_n5359__), .dout(new_new_n3849__));
  and1  g1665(.dina(new_new_n5358__), .dinb(new_new_n5359__), .dout(new_new_n3850__));
  or1   g1666(.dina(new_new_n5356__), .dinb(new_new_n5357__), .dout(new_new_n3851__));
  and1  g1667(.dina(new_new_n3851__), .dinb(new_new_n3849__), .dout(new_new_n3852__));
  or1   g1668(.dina(new_new_n3850__), .dinb(new_new_n3848__), .dout(new_new_n3853__));
  and1  g1669(.dina(new_new_n3078__), .dinb(new_new_n2955__), .dout(new_new_n3854__));
  or1   g1670(.dina(new_new_n3079__), .dinb(new_new_n2954__), .dout(new_new_n3855__));
  and1  g1671(.dina(new_new_n3106__), .dinb(new_new_n2855__), .dout(new_new_n3856__));
  or1   g1672(.dina(new_new_n3107__), .dinb(new_new_n2854__), .dout(new_new_n3857__));
  and1  g1673(.dina(new_new_n3857__), .dinb(new_new_n3855__), .dout(new_new_n3858__));
  or1   g1674(.dina(new_new_n3856__), .dinb(new_new_n3854__), .dout(new_new_n3859__));
  and1  g1675(.dina(new_new_n5360__), .dinb(new_new_n5361__), .dout(new_new_n3860__));
  and1  g1676(.dina(new_new_n3860__), .dinb(new_new_n5362__), .dout(new_new_n3861__));
  and1  g1677(.dina(new_new_n5360__), .dinb(new_new_n5363__), .dout(new_new_n3862__));
  and1  g1678(.dina(new_new_n3862__), .dinb(new_new_n5364__), .dout(new_new_n3863__));
  or1   g1679(.dina(new_new_n3863__), .dinb(new_new_n3861__), .dout(new_new_n3864__));
  and1  g1680(.dina(new_new_n5365__), .dinb(new_new_n5363__), .dout(new_new_n3865__));
  and1  g1681(.dina(new_new_n3865__), .dinb(new_new_n5362__), .dout(new_new_n3866__));
  and1  g1682(.dina(new_new_n5365__), .dinb(new_new_n5361__), .dout(new_new_n3867__));
  and1  g1683(.dina(new_new_n3867__), .dinb(new_new_n5364__), .dout(new_new_n3868__));
  or1   g1684(.dina(new_new_n3868__), .dinb(new_new_n3866__), .dout(new_new_n3869__));
  or1   g1685(.dina(new_new_n3869__), .dinb(new_new_n3864__), .dout(new_new_n3870__));
  and1  g1686(.dina(new_new_n5366__), .dinb(new_new_n5367__), .dout(new_new_n3871__));
  or1   g1687(.dina(new_new_n5368__), .dinb(new_new_n5369__), .dout(new_new_n3872__));
  and1  g1688(.dina(new_new_n5368__), .dinb(new_new_n5369__), .dout(new_new_n3873__));
  or1   g1689(.dina(new_new_n5366__), .dinb(new_new_n5367__), .dout(new_new_n3874__));
  and1  g1690(.dina(new_new_n3874__), .dinb(new_new_n3872__), .dout(new_new_n3875__));
  or1   g1691(.dina(new_new_n3873__), .dinb(new_new_n3871__), .dout(new_new_n3876__));
  and1  g1692(.dina(new_new_n5370__), .dinb(new_new_n5371__), .dout(new_new_n3877__));
  or1   g1693(.dina(new_new_n5372__), .dinb(new_new_n5373__), .dout(new_new_n3878__));
  and1  g1694(.dina(new_new_n5372__), .dinb(new_new_n5373__), .dout(new_new_n3879__));
  or1   g1695(.dina(new_new_n5370__), .dinb(new_new_n5371__), .dout(new_new_n3880__));
  and1  g1696(.dina(new_new_n3880__), .dinb(new_new_n3878__), .dout(new_new_n3881__));
  or1   g1697(.dina(new_new_n3879__), .dinb(new_new_n3877__), .dout(new_new_n3882__));
  and1  g1698(.dina(new_new_n3083__), .dinb(new_new_n2949__), .dout(new_new_n3883__));
  or1   g1699(.dina(new_new_n3082__), .dinb(new_new_n2948__), .dout(new_new_n3884__));
  and1  g1700(.dina(new_new_n3096__), .dinb(new_new_n2858__), .dout(new_new_n3885__));
  or1   g1701(.dina(new_new_n3097__), .dinb(new_new_n2859__), .dout(new_new_n3886__));
  and1  g1702(.dina(new_new_n3886__), .dinb(new_new_n3884__), .dout(new_new_n3887__));
  or1   g1703(.dina(new_new_n3885__), .dinb(new_new_n3883__), .dout(new_new_n3888__));
  or1   g1704(.dina(new_new_n5374__), .dinb(new_new_n5375__), .dout(new_new_n3889__));
  or1   g1705(.dina(new_new_n3889__), .dinb(new_new_n5376__), .dout(new_new_n3890__));
  or1   g1706(.dina(new_new_n5374__), .dinb(new_new_n5377__), .dout(new_new_n3891__));
  or1   g1707(.dina(new_new_n3891__), .dinb(new_new_n5378__), .dout(new_new_n3892__));
  and1  g1708(.dina(new_new_n3892__), .dinb(new_new_n3890__), .dout(new_new_n3893__));
  or1   g1709(.dina(new_new_n5379__), .dinb(new_new_n5377__), .dout(new_new_n3894__));
  or1   g1710(.dina(new_new_n3894__), .dinb(new_new_n5376__), .dout(new_new_n3895__));
  or1   g1711(.dina(new_new_n5379__), .dinb(new_new_n5375__), .dout(new_new_n3896__));
  or1   g1712(.dina(new_new_n3896__), .dinb(new_new_n5378__), .dout(new_new_n3897__));
  and1  g1713(.dina(new_new_n3897__), .dinb(new_new_n3895__), .dout(new_new_n3898__));
  and1  g1714(.dina(new_new_n3898__), .dinb(new_new_n3893__), .dout(new_new_n3899__));
  and1  g1715(.dina(new_new_n5196__), .dinb(new_new_n5380__), .dout(new_new_n3900__));
  and1  g1716(.dina(new_new_n5207__), .dinb(new_new_n5381__), .dout(new_new_n3901__));
  or1   g1717(.dina(new_new_n3901__), .dinb(new_new_n3900__), .dout(new_new_n3902__));
  or1   g1718(.dina(new_new_n5196__), .dinb(new_new_n5383__), .dout(new_new_n3903__));
  or1   g1719(.dina(new_new_n3903__), .dinb(new_new_n5388__), .dout(new_new_n3904__));
  or1   g1720(.dina(new_new_n5198__), .dinb(new_new_n5401__), .dout(new_new_n3905__));
  or1   g1721(.dina(new_new_n3905__), .dinb(new_new_n5388__), .dout(new_new_n3906__));
  and1  g1722(.dina(new_new_n5224__), .dinb(new_new_n5380__), .dout(new_new_n3907__));
  and1  g1723(.dina(new_new_n5234__), .dinb(new_new_n5381__), .dout(new_new_n3908__));
  or1   g1724(.dina(new_new_n3908__), .dinb(new_new_n3907__), .dout(new_new_n3909__));
  or1   g1725(.dina(new_new_n5224__), .dinb(new_new_n5383__), .dout(new_new_n3910__));
  or1   g1726(.dina(new_new_n3910__), .dinb(new_new_n5389__), .dout(new_new_n3911__));
  or1   g1727(.dina(new_new_n5226__), .dinb(new_new_n5401__), .dout(new_new_n3912__));
  or1   g1728(.dina(new_new_n3912__), .dinb(new_new_n5389__), .dout(new_new_n3913__));
  or1   g1729(.dina(new_new_n5198__), .dinb(new_new_n5405__), .dout(new_new_n3914__));
  and1  g1730(.dina(new_new_n2817__), .dinb(new_new_n2810__), .dout(new_new_n3915__));
  or1   g1731(.dina(new_new_n2816__), .dinb(new_new_n2811__), .dout(new_new_n3916__));
  and1  g1732(.dina(new_new_n3915__), .dinb(new_new_n3163__), .dout(new_new_n3917__));
  or1   g1733(.dina(new_new_n3916__), .dinb(new_new_n3162__), .dout(new_new_n3918__));
  or1   g1734(.dina(new_new_n5409__), .dinb(new_new_n3914__), .dout(new_new_n3919__));
  or1   g1735(.dina(new_new_n5226__), .dinb(new_new_n5405__), .dout(new_new_n3920__));
  or1   g1736(.dina(new_new_n3920__), .dinb(new_new_n5409__), .dout(new_new_n3921__));
  and1  g1737(.dina(new_new_n5207__), .dinb(new_new_n5411__), .dout(new_new_n3922__));
  and1  g1738(.dina(new_new_n3922__), .dinb(new_new_n5414__), .dout(new_new_n3923__));
  and1  g1739(.dina(new_new_n5209__), .dinb(new_new_n5419__), .dout(new_new_n3924__));
  and1  g1740(.dina(new_new_n3924__), .dinb(new_new_n5414__), .dout(new_new_n3925__));
  and1  g1741(.dina(new_new_n5234__), .dinb(new_new_n5411__), .dout(new_new_n3926__));
  and1  g1742(.dina(new_new_n3926__), .dinb(new_new_n5415__), .dout(new_new_n3927__));
  and1  g1743(.dina(new_new_n5236__), .dinb(new_new_n5419__), .dout(new_new_n3928__));
  and1  g1744(.dina(new_new_n3928__), .dinb(new_new_n5415__), .dout(new_new_n3929__));
  or1   g1745(.dina(new_new_n5209__), .dinb(new_new_n5421__), .dout(new_new_n3930__));
  or1   g1746(.dina(new_new_n5197__), .dinb(new_new_n5424__), .dout(new_new_n3931__));
  and1  g1747(.dina(new_new_n3931__), .dinb(new_new_n3930__), .dout(new_new_n3932__));
  or1   g1748(.dina(new_new_n3932__), .dinb(new_new_n5391__), .dout(new_new_n3933__));
  or1   g1749(.dina(new_new_n5208__), .dinb(new_new_n5427__), .dout(new_new_n3934__));
  or1   g1750(.dina(new_new_n5200__), .dinb(new_new_n5430__), .dout(new_new_n3935__));
  and1  g1751(.dina(new_new_n3935__), .dinb(new_new_n3934__), .dout(new_new_n3936__));
  or1   g1752(.dina(new_new_n3936__), .dinb(new_new_n5391__), .dout(new_new_n3937__));
  or1   g1753(.dina(new_new_n5236__), .dinb(new_new_n5421__), .dout(new_new_n3938__));
  or1   g1754(.dina(new_new_n5225__), .dinb(new_new_n5424__), .dout(new_new_n3939__));
  and1  g1755(.dina(new_new_n3939__), .dinb(new_new_n3938__), .dout(new_new_n3940__));
  or1   g1756(.dina(new_new_n3940__), .dinb(new_new_n5392__), .dout(new_new_n3941__));
  or1   g1757(.dina(new_new_n5235__), .dinb(new_new_n5427__), .dout(new_new_n3942__));
  or1   g1758(.dina(new_new_n5228__), .dinb(new_new_n5430__), .dout(new_new_n3943__));
  and1  g1759(.dina(new_new_n3943__), .dinb(new_new_n3942__), .dout(new_new_n3944__));
  or1   g1760(.dina(new_new_n3944__), .dinb(new_new_n5392__), .dout(new_new_n3945__));
  or1   g1761(.dina(new_new_n5434__), .dinb(new_new_n5437__), .dout(new_new_n3946__));
  or1   g1762(.dina(new_new_n3946__), .dinb(new_new_n5395__), .dout(new_new_n3947__));
  or1   g1763(.dina(new_new_n5441__), .dinb(new_new_n5437__), .dout(new_new_n3948__));
  or1   g1764(.dina(new_new_n3948__), .dinb(new_new_n5395__), .dout(new_new_n3949__));
  or1   g1765(.dina(new_new_n5434__), .dinb(new_new_n5444__), .dout(new_new_n3950__));
  or1   g1766(.dina(new_new_n3950__), .dinb(new_new_n5396__), .dout(new_new_n3951__));
  or1   g1767(.dina(new_new_n5441__), .dinb(new_new_n5444__), .dout(new_new_n3952__));
  or1   g1768(.dina(new_new_n3952__), .dinb(new_new_n5396__), .dout(new_new_n3953__));
  and1  g1769(.dina(new_new_n5447__), .dinb(new_new_n5448__), .dout(new_new_n3954__));
  and1  g1770(.dina(new_new_n3954__), .dinb(new_new_n5417__), .dout(new_new_n3955__));
  and1  g1771(.dina(new_new_n5450__), .dinb(new_new_n5448__), .dout(new_new_n3956__));
  and1  g1772(.dina(new_new_n3956__), .dinb(new_new_n5417__), .dout(new_new_n3957__));
  or1   g1773(.dina(new_new_n5452__), .dinb(new_new_n5453__), .dout(new_new_n3958__));
  or1   g1774(.dina(new_new_n3958__), .dinb(new_new_n5410__), .dout(new_new_n3959__));
  or1   g1775(.dina(new_new_n5456__), .dinb(new_new_n5438__), .dout(new_new_n3960__));
  or1   g1776(.dina(new_new_n5456__), .dinb(new_new_n5461__), .dout(new_new_n3961__));
  and1  g1777(.dina(new_new_n3961__), .dinb(new_new_n3960__), .dout(new_new_n3962__));
  or1   g1778(.dina(new_new_n3962__), .dinb(new_new_n5398__), .dout(new_new_n3963__));
  or1   g1779(.dina(new_new_n5464__), .dinb(new_new_n5438__), .dout(new_new_n3964__));
  or1   g1780(.dina(new_new_n5464__), .dinb(new_new_n5461__), .dout(new_new_n3965__));
  and1  g1781(.dina(new_new_n3965__), .dinb(new_new_n3964__), .dout(new_new_n3966__));
  or1   g1782(.dina(new_new_n3966__), .dinb(new_new_n5398__), .dout(new_new_n3967__));
  or1   g1783(.dina(new_new_n5457__), .dinb(new_new_n5445__), .dout(new_new_n3968__));
  or1   g1784(.dina(new_new_n5457__), .dinb(new_new_n5468__), .dout(new_new_n3969__));
  and1  g1785(.dina(new_new_n3969__), .dinb(new_new_n3968__), .dout(new_new_n3970__));
  or1   g1786(.dina(new_new_n3970__), .dinb(new_new_n5399__), .dout(new_new_n3971__));
  or1   g1787(.dina(new_new_n5465__), .dinb(new_new_n5445__), .dout(new_new_n3972__));
  or1   g1788(.dina(new_new_n5465__), .dinb(new_new_n5468__), .dout(new_new_n3973__));
  and1  g1789(.dina(new_new_n3973__), .dinb(new_new_n3972__), .dout(new_new_n3974__));
  or1   g1790(.dina(new_new_n3974__), .dinb(new_new_n5399__), .dout(new_new_n3975__));
  and1  g1791(.dina(new_new_n5211__), .dinb(new_new_n5469__), .dout(new_new_n3976__));
  and1  g1792(.dina(new_new_n3976__), .dinb(new_new_n5418__), .dout(new_new_n3977__));
  and1  g1793(.dina(new_new_n5238__), .dinb(new_new_n5469__), .dout(new_new_n3978__));
  and1  g1794(.dina(new_new_n3978__), .dinb(new_new_n5418__), .dout(new_new_n3979__));
  and1  g1795(.dina(new_new_n5113__), .dinb(new_new_n2326__), .dout(new_new_n3980__));
  and1  g1796(.dina(new_new_n3980__), .dinb(new_new_n5120__), .dout(new_new_n3981__));
  and1  g1797(.dina(new_new_n5127__), .dinb(new_new_n2236__), .dout(new_new_n3982__));
  and1  g1798(.dina(new_new_n3982__), .dinb(new_new_n5120__), .dout(new_new_n3983__));
  and1  g1799(.dina(new_new_n5113__), .dinb(new_new_n2296__), .dout(new_new_n3984__));
  and1  g1800(.dina(new_new_n3984__), .dinb(new_new_n5134__), .dout(new_new_n3985__));
  and1  g1801(.dina(new_new_n5127__), .dinb(new_new_n2266__), .dout(new_new_n3986__));
  and1  g1802(.dina(new_new_n3986__), .dinb(new_new_n5134__), .dout(new_new_n3987__));
  or1   g1803(.dina(new_new_n3983__), .dinb(new_new_n3981__), .dout(new_new_n3988__));
  or1   g1804(.dina(new_new_n3988__), .dinb(new_new_n3985__), .dout(new_new_n3989__));
  or1   g1805(.dina(new_new_n3989__), .dinb(new_new_n3987__), .dout(new_new_n3990__));
  and1  g1806(.dina(new_new_n5143__), .dinb(new_new_n2178__), .dout(new_new_n3991__));
  and1  g1807(.dina(new_new_n3991__), .dinb(new_new_n5157__), .dout(new_new_n3992__));
  and1  g1808(.dina(new_new_n5171__), .dinb(new_new_n2084__), .dout(new_new_n3993__));
  and1  g1809(.dina(new_new_n3993__), .dinb(new_new_n5157__), .dout(new_new_n3994__));
  and1  g1810(.dina(new_new_n5143__), .dinb(new_new_n2116__), .dout(new_new_n3995__));
  and1  g1811(.dina(new_new_n3995__), .dinb(new_new_n5185__), .dout(new_new_n3996__));
  and1  g1812(.dina(new_new_n5171__), .dinb(new_new_n2146__), .dout(new_new_n3997__));
  and1  g1813(.dina(new_new_n3997__), .dinb(new_new_n5185__), .dout(new_new_n3998__));
  or1   g1814(.dina(new_new_n3994__), .dinb(new_new_n3992__), .dout(new_new_n3999__));
  or1   g1815(.dina(new_new_n3999__), .dinb(new_new_n3996__), .dout(new_new_n4000__));
  or1   g1816(.dina(new_new_n4000__), .dinb(new_new_n3998__), .dout(new_new_n4001__));
  and1  g1817(.dina(new_new_n5144__), .dinb(new_new_n2206__), .dout(new_new_n4002__));
  and1  g1818(.dina(new_new_n4002__), .dinb(new_new_n5158__), .dout(new_new_n4003__));
  and1  g1819(.dina(new_new_n5172__), .dinb(new_new_n2112__), .dout(new_new_n4004__));
  and1  g1820(.dina(new_new_n4004__), .dinb(new_new_n5158__), .dout(new_new_n4005__));
  and1  g1821(.dina(new_new_n5144__), .dinb(new_new_n2142__), .dout(new_new_n4006__));
  and1  g1822(.dina(new_new_n4006__), .dinb(new_new_n5186__), .dout(new_new_n4007__));
  and1  g1823(.dina(new_new_n5172__), .dinb(new_new_n2174__), .dout(new_new_n4008__));
  and1  g1824(.dina(new_new_n4008__), .dinb(new_new_n5186__), .dout(new_new_n4009__));
  or1   g1825(.dina(new_new_n4005__), .dinb(new_new_n4003__), .dout(new_new_n4010__));
  or1   g1826(.dina(new_new_n4010__), .dinb(new_new_n4007__), .dout(new_new_n4011__));
  or1   g1827(.dina(new_new_n4011__), .dinb(new_new_n4009__), .dout(new_new_n4012__));
  or1   g1828(.dina(new_new_n5471__), .dinb(new_new_n5453__), .dout(new_new_n4013__));
  or1   g1829(.dina(new_new_n4013__), .dinb(new_new_n5410__), .dout(new_new_n4014__));
  and1  g1830(.dina(new_new_n5476__), .dinb(new_new_n3236__), .dout(new_new_n4015__));
  and1  g1831(.dina(new_new_n4015__), .dinb(new_new_n5485__), .dout(new_new_n4016__));
  and1  g1832(.dina(new_new_n5493__), .dinb(new_new_n3224__), .dout(new_new_n4017__));
  and1  g1833(.dina(new_new_n4017__), .dinb(new_new_n5485__), .dout(new_new_n4018__));
  and1  g1834(.dina(new_new_n5476__), .dinb(new_new_n3232__), .dout(new_new_n4019__));
  and1  g1835(.dina(new_new_n4019__), .dinb(new_new_n5498__), .dout(new_new_n4020__));
  and1  g1836(.dina(new_new_n5493__), .dinb(new_new_n3228__), .dout(new_new_n4021__));
  and1  g1837(.dina(new_new_n4021__), .dinb(new_new_n5498__), .dout(new_new_n4022__));
  or1   g1838(.dina(new_new_n4018__), .dinb(new_new_n4016__), .dout(new_new_n4023__));
  or1   g1839(.dina(new_new_n4023__), .dinb(new_new_n4020__), .dout(new_new_n4024__));
  or1   g1840(.dina(new_new_n4024__), .dinb(new_new_n4022__), .dout(new_new_n4025__));
  or1   g1841(.dina(new_new_n5494__), .dinb(new_new_n3239__), .dout(new_new_n4026__));
  or1   g1842(.dina(new_new_n4026__), .dinb(new_new_n5499__), .dout(new_new_n4027__));
  or1   g1843(.dina(new_new_n5477__), .dinb(new_new_n3227__), .dout(new_new_n4028__));
  or1   g1844(.dina(new_new_n4028__), .dinb(new_new_n5499__), .dout(new_new_n4029__));
  or1   g1845(.dina(new_new_n5494__), .dinb(new_new_n3235__), .dout(new_new_n4030__));
  or1   g1846(.dina(new_new_n4030__), .dinb(new_new_n5486__), .dout(new_new_n4031__));
  or1   g1847(.dina(new_new_n5477__), .dinb(new_new_n3231__), .dout(new_new_n4032__));
  or1   g1848(.dina(new_new_n4032__), .dinb(new_new_n5486__), .dout(new_new_n4033__));
  and1  g1849(.dina(new_new_n4029__), .dinb(new_new_n4027__), .dout(new_new_n4034__));
  and1  g1850(.dina(new_new_n4034__), .dinb(new_new_n4031__), .dout(new_new_n4035__));
  and1  g1851(.dina(new_new_n4035__), .dinb(new_new_n4033__), .dout(new_new_n4036__));
  and1  g1852(.dina(new_new_n5501__), .dinb(new_new_n5502__), .dout(new_new_n4037__));
  or1   g1853(.dina(new_new_n5503__), .dinb(new_new_n5504__), .dout(new_new_n4038__));
  and1  g1854(.dina(new_new_n5503__), .dinb(new_new_n5504__), .dout(new_new_n4039__));
  or1   g1855(.dina(new_new_n5501__), .dinb(new_new_n5502__), .dout(new_new_n4040__));
  and1  g1856(.dina(new_new_n4040__), .dinb(new_new_n4038__), .dout(new_new_n4041__));
  or1   g1857(.dina(new_new_n4039__), .dinb(new_new_n4037__), .dout(new_new_n4042__));
  and1  g1858(.dina(new_new_n5505__), .dinb(new_new_n5506__), .dout(new_new_n4043__));
  or1   g1859(.dina(new_new_n5507__), .dinb(new_new_n5508__), .dout(new_new_n4044__));
  and1  g1860(.dina(new_new_n5507__), .dinb(new_new_n5508__), .dout(new_new_n4045__));
  or1   g1861(.dina(new_new_n5505__), .dinb(new_new_n5506__), .dout(new_new_n4046__));
  and1  g1862(.dina(new_new_n4046__), .dinb(new_new_n4044__), .dout(new_new_n4047__));
  or1   g1863(.dina(new_new_n4045__), .dinb(new_new_n4043__), .dout(new_new_n4048__));
  and1  g1864(.dina(new_new_n2616__), .dinb(new_new_n2593__), .dout(new_new_n4049__));
  and1  g1865(.dina(new_new_n2617__), .dinb(new_new_n2592__), .dout(new_new_n4050__));
  or1   g1866(.dina(new_new_n4050__), .dinb(new_new_n4049__), .dout(new_new_n4051__));
  or1   g1867(.dina(new_new_n5509__), .dinb(new_new_n5510__), .dout(new_new_n4052__));
  or1   g1868(.dina(new_new_n4052__), .dinb(new_new_n5512__), .dout(new_new_n4053__));
  and1  g1869(.dina(new_new_n5514__), .dinb(new_new_n5510__), .dout(new_new_n4054__));
  and1  g1870(.dina(new_new_n4054__), .dinb(new_new_n5512__), .dout(new_new_n4055__));
  and1  g1871(.dina(new_new_n5516__), .dinb(new_new_n5517__), .dout(new_new_n4056__));
  or1   g1872(.dina(new_new_n5518__), .dinb(new_new_n5520__), .dout(new_new_n4057__));
  and1  g1873(.dina(new_new_n5518__), .dinb(new_new_n5520__), .dout(new_new_n4058__));
  or1   g1874(.dina(new_new_n5516__), .dinb(new_new_n5517__), .dout(new_new_n4059__));
  and1  g1875(.dina(new_new_n4059__), .dinb(new_new_n4057__), .dout(new_new_n4060__));
  or1   g1876(.dina(new_new_n4058__), .dinb(new_new_n4056__), .dout(new_new_n4061__));
  and1  g1877(.dina(new_new_n5521__), .dinb(new_new_n5522__), .dout(new_new_n4062__));
  or1   g1878(.dina(new_new_n5523__), .dinb(new_new_n5524__), .dout(new_new_n4063__));
  and1  g1879(.dina(new_new_n5523__), .dinb(new_new_n5524__), .dout(new_new_n4064__));
  or1   g1880(.dina(new_new_n5521__), .dinb(new_new_n5522__), .dout(new_new_n4065__));
  and1  g1881(.dina(new_new_n4065__), .dinb(new_new_n4063__), .dout(new_new_n4066__));
  or1   g1882(.dina(new_new_n4064__), .dinb(new_new_n4062__), .dout(new_new_n4067__));
  and1  g1883(.dina(new_new_n5525__), .dinb(new_new_n2599__), .dout(new_new_n4068__));
  and1  g1884(.dina(new_new_n2601__), .dinb(new_new_n5526__), .dout(new_new_n4069__));
  or1   g1885(.dina(new_new_n4069__), .dinb(new_new_n4068__), .dout(new_new_n4070__));
  or1   g1886(.dina(new_new_n5527__), .dinb(new_new_n5528__), .dout(new_new_n4071__));
  or1   g1887(.dina(new_new_n4071__), .dinb(new_new_n5530__), .dout(new_new_n4072__));
  and1  g1888(.dina(new_new_n5532__), .dinb(new_new_n5528__), .dout(new_new_n4073__));
  and1  g1889(.dina(new_new_n4073__), .dinb(new_new_n5530__), .dout(new_new_n4074__));
  and1  g1890(.dina(new_new_n5509__), .dinb(new_new_n5533__), .dout(new_new_n4075__));
  and1  g1891(.dina(new_new_n4075__), .dinb(new_new_n5513__), .dout(new_new_n4076__));
  and1  g1892(.dina(new_new_n5527__), .dinb(new_new_n5534__), .dout(new_new_n4077__));
  and1  g1893(.dina(new_new_n4077__), .dinb(new_new_n5531__), .dout(new_new_n4078__));
  and1  g1894(.dina(new_new_n5535__), .dinb(new_new_n5536__), .dout(new_new_n4079__));
  or1   g1895(.dina(new_new_n5537__), .dinb(new_new_n5538__), .dout(new_new_n4080__));
  and1  g1896(.dina(new_new_n5537__), .dinb(new_new_n5538__), .dout(new_new_n4081__));
  or1   g1897(.dina(new_new_n5535__), .dinb(new_new_n5536__), .dout(new_new_n4082__));
  and1  g1898(.dina(new_new_n4082__), .dinb(new_new_n4080__), .dout(new_new_n4083__));
  or1   g1899(.dina(new_new_n4081__), .dinb(new_new_n4079__), .dout(new_new_n4084__));
  and1  g1900(.dina(new_new_n5268__), .dinb(new_new_n2688__), .dout(new_new_n4085__));
  and1  g1901(.dina(new_new_n5270__), .dinb(new_new_n2689__), .dout(new_new_n4086__));
  or1   g1902(.dina(new_new_n4086__), .dinb(new_new_n4085__), .dout(new_new_n4087__));
  or1   g1903(.dina(new_new_n5539__), .dinb(new_new_n5541__), .dout(new_new_n4088__));
  or1   g1904(.dina(new_new_n4088__), .dinb(new_new_n5544__), .dout(new_new_n4089__));
  and1  g1905(.dina(new_new_n5546__), .dinb(new_new_n5541__), .dout(new_new_n4090__));
  and1  g1906(.dina(new_new_n4090__), .dinb(new_new_n5544__), .dout(new_new_n4091__));
  and1  g1907(.dina(new_new_n5539__), .dinb(new_new_n5547__), .dout(new_new_n4092__));
  and1  g1908(.dina(new_new_n4092__), .dinb(new_new_n5545__), .dout(new_new_n4093__));
  or1   g1909(.dina(new_new_n5514__), .dinb(new_new_n5533__), .dout(new_new_n4094__));
  or1   g1910(.dina(new_new_n4094__), .dinb(new_new_n5513__), .dout(new_new_n4095__));
  or1   g1911(.dina(new_new_n5532__), .dinb(new_new_n5534__), .dout(new_new_n4096__));
  or1   g1912(.dina(new_new_n4096__), .dinb(new_new_n5531__), .dout(new_new_n4097__));
  or1   g1913(.dina(new_new_n5546__), .dinb(new_new_n5547__), .dout(new_new_n4098__));
  or1   g1914(.dina(new_new_n4098__), .dinb(new_new_n5545__), .dout(new_new_n4099__));
  and1  g1915(.dina(new_new_n5551__), .dinb(new_new_n1918__), .dout(new_new_n4100__));
  and1  g1916(.dina(new_new_n5102__), .dinb(new_new_n5559__), .dout(new_new_n4101__));
  or1   g1917(.dina(new_new_n4101__), .dinb(new_new_n4100__), .dout(new_new_n4102__));
  and1  g1918(.dina(new_new_n5551__), .dinb(new_new_n1924__), .dout(new_new_n4103__));
  and1  g1919(.dina(new_new_n5564__), .dinb(new_new_n5559__), .dout(new_new_n4104__));
  or1   g1920(.dina(new_new_n4104__), .dinb(new_new_n4103__), .dout(new_new_n4105__));
  and1  g1921(.dina(new_new_n5550__), .dinb(new_new_n1930__), .dout(new_new_n4106__));
  and1  g1922(.dina(new_new_n2604__), .dinb(new_new_n5558__), .dout(new_new_n4107__));
  or1   g1923(.dina(new_new_n4107__), .dinb(new_new_n4106__), .dout(new_new_n4108__));
  and1  g1924(.dina(new_new_n1976__), .dinb(new_new_n5552__), .dout(new_new_n4109__));
  and1  g1925(.dina(new_new_n5566__), .dinb(new_new_n5560__), .dout(new_new_n4110__));
  or1   g1926(.dina(new_new_n4110__), .dinb(new_new_n4109__), .dout(new_new_n4111__));
  and1  g1927(.dina(new_new_n1982__), .dinb(new_new_n5552__), .dout(new_new_n4112__));
  and1  g1928(.dina(new_new_n2648__), .dinb(new_new_n5560__), .dout(new_new_n4113__));
  or1   g1929(.dina(new_new_n4113__), .dinb(new_new_n4112__), .dout(new_new_n4114__));
  and1  g1930(.dina(new_new_n1988__), .dinb(new_new_n5554__), .dout(new_new_n4115__));
  and1  g1931(.dina(new_new_n5567__), .dinb(new_new_n5562__), .dout(new_new_n4116__));
  or1   g1932(.dina(new_new_n4116__), .dinb(new_new_n4115__), .dout(new_new_n4117__));
  and1  g1933(.dina(new_new_n1994__), .dinb(new_new_n5554__), .dout(new_new_n4118__));
  and1  g1934(.dina(new_new_n5568__), .dinb(new_new_n5562__), .dout(new_new_n4119__));
  or1   g1935(.dina(new_new_n4119__), .dinb(new_new_n4118__), .dout(new_new_n4120__));
  and1  g1936(.dina(new_new_n2000__), .dinb(new_new_n5555__), .dout(new_new_n4121__));
  and1  g1937(.dina(new_new_n2606__), .dinb(new_new_n5563__), .dout(new_new_n4122__));
  or1   g1938(.dina(new_new_n4122__), .dinb(new_new_n4121__), .dout(new_new_n4123__));
  and1  g1939(.dina(new_new_n2006__), .dinb(new_new_n5555__), .dout(new_new_n4124__));
  and1  g1940(.dina(new_new_n2642__), .dinb(new_new_n5563__), .dout(new_new_n4125__));
  or1   g1941(.dina(new_new_n4125__), .dinb(new_new_n4124__), .dout(new_new_n4126__));
  and1  g1942(.dina(new_new_n5572__), .dinb(new_new_n2012__), .dout(new_new_n4127__));
  and1  g1943(.dina(new_new_n2644__), .dinb(new_new_n5579__), .dout(new_new_n4128__));
  or1   g1944(.dina(new_new_n4128__), .dinb(new_new_n4127__), .dout(new_new_n4129__));
  and1  g1945(.dina(new_new_n5572__), .dinb(new_new_n2018__), .dout(new_new_n4130__));
  and1  g1946(.dina(new_new_n2608__), .dinb(new_new_n5579__), .dout(new_new_n4131__));
  or1   g1947(.dina(new_new_n4131__), .dinb(new_new_n4130__), .dout(new_new_n4132__));
  and1  g1948(.dina(new_new_n5571__), .dinb(new_new_n2024__), .dout(new_new_n4133__));
  and1  g1949(.dina(new_new_n5583__), .dinb(new_new_n5580__), .dout(new_new_n4134__));
  or1   g1950(.dina(new_new_n4134__), .dinb(new_new_n4133__), .dout(new_new_n4135__));
  and1  g1951(.dina(new_new_n2044__), .dinb(new_new_n5573__), .dout(new_new_n4136__));
  and1  g1952(.dina(new_new_n2646__), .dinb(new_new_n5580__), .dout(new_new_n4137__));
  or1   g1953(.dina(new_new_n4137__), .dinb(new_new_n4136__), .dout(new_new_n4138__));
  and1  g1954(.dina(new_new_n2050__), .dinb(new_new_n5573__), .dout(new_new_n4139__));
  and1  g1955(.dina(new_new_n2796__), .dinb(new_new_n5582__), .dout(new_new_n4140__));
  or1   g1956(.dina(new_new_n4140__), .dinb(new_new_n4139__), .dout(new_new_n4141__));
  and1  g1957(.dina(new_new_n2056__), .dinb(new_new_n5575__), .dout(new_new_n4142__));
  and1  g1958(.dina(new_new_n5327__), .dinb(new_new_n5582__), .dout(new_new_n4143__));
  or1   g1959(.dina(new_new_n4143__), .dinb(new_new_n4142__), .dout(new_new_n4144__));
  and1  g1960(.dina(new_new_n2062__), .dinb(new_new_n5575__), .dout(new_new_n4145__));
  and1  g1961(.dina(new_new_n5322__), .dinb(new_new_n5581__), .dout(new_new_n4146__));
  or1   g1962(.dina(new_new_n4146__), .dinb(new_new_n4145__), .dout(new_new_n4147__));
  or1   g1963(.dina(new_new_n5566__), .dinb(new_new_n5103__), .dout(new_new_n4148__));
  or1   g1964(.dina(new_new_n2799__), .dinb(new_new_n5100__), .dout(new_new_n4149__));
  and1  g1965(.dina(new_new_n4149__), .dinb(new_new_n4148__), .dout(new_new_n4150__));
  and1  g1966(.dina(new_new_n5584__), .dinb(new_new_n5585__), .dout(new_new_n4151__));
  or1   g1967(.dina(new_new_n5586__), .dinb(new_new_n2408__), .dout(new_new_n4152__));
  or1   g1968(.dina(new_new_n5587__), .dinb(new_new_n5589__), .dout(new_new_n4153__));
  or1   g1969(.dina(new_new_n4153__), .dinb(new_new_n2081__), .dout(new_new_n4154__));
  and1  g1970(.dina(new_new_n5200__), .dinb(new_new_n5590__), .dout(new_new_n4155__));
  or1   g1971(.dina(new_new_n5211__), .dinb(new_new_n5406__), .dout(new_new_n4156__));
  and1  g1972(.dina(new_new_n5212__), .dinb(new_new_n5591__), .dout(new_new_n4157__));
  or1   g1973(.dina(new_new_n5201__), .dinb(new_new_n5593__), .dout(new_new_n4158__));
  and1  g1974(.dina(new_new_n4158__), .dinb(new_new_n4156__), .dout(new_new_n4159__));
  or1   g1975(.dina(new_new_n4157__), .dinb(new_new_n4155__), .dout(new_new_n4160__));
  or1   g1976(.dina(new_new_n5595__), .dinb(new_new_n5598__), .dout(new_new_n4161__));
  and1  g1977(.dina(new_new_n5228__), .dinb(new_new_n5590__), .dout(new_new_n4162__));
  or1   g1978(.dina(new_new_n5238__), .dinb(new_new_n5406__), .dout(new_new_n4163__));
  and1  g1979(.dina(new_new_n5239__), .dinb(new_new_n5591__), .dout(new_new_n4164__));
  or1   g1980(.dina(new_new_n5229__), .dinb(new_new_n5593__), .dout(new_new_n4165__));
  and1  g1981(.dina(new_new_n4165__), .dinb(new_new_n4163__), .dout(new_new_n4166__));
  or1   g1982(.dina(new_new_n4164__), .dinb(new_new_n4162__), .dout(new_new_n4167__));
  or1   g1983(.dina(new_new_n5602__), .dinb(new_new_n5598__), .dout(new_new_n4168__));
  or1   g1984(.dina(new_new_n5604__), .dinb(new_new_n5606__), .dout(new_new_n4169__));
  and1  g1985(.dina(new_new_n5609__), .dinb(new_new_n5611__), .dout(new_new_n4170__));
  and1  g1986(.dina(new_new_n5613__), .dinb(new_new_n5615__), .dout(new_new_n4171__));
  or1   g1987(.dina(new_new_n5617__), .dinb(new_new_n5606__), .dout(new_new_n4172__));
  and1  g1988(.dina(new_new_n5619__), .dinb(new_new_n5621__), .dout(new_new_n4173__));
  and1  g1989(.dina(new_new_n5623__), .dinb(new_new_n5625__), .dout(new_new_n4174__));
  and1  g1990(.dina(new_new_n5628__), .dinb(new_new_n5632__), .dout(new_new_n4175__));
  and1  g1991(.dina(new_new_n5628__), .dinb(new_new_n5634__), .dout(new_new_n4176__));
  or1   g1992(.dina(new_new_n5637__), .dinb(new_new_n5641__), .dout(new_new_n4177__));
  or1   g1993(.dina(new_new_n5644__), .dinb(new_new_n5648__), .dout(new_new_n4178__));
  or1   g1994(.dina(new_new_n5637__), .dinb(new_new_n5650__), .dout(new_new_n4179__));
  or1   g1995(.dina(new_new_n5644__), .dinb(new_new_n5652__), .dout(new_new_n4180__));
  and1  g1996(.dina(new_new_n5654__), .dinb(new_new_n5656__), .dout(new_new_n4181__));
  and1  g1997(.dina(new_new_n5658__), .dinb(new_new_n5660__), .dout(new_new_n4182__));
  and1  g1998(.dina(new_new_n5662__), .dinb(new_new_n5664__), .dout(new_new_n4183__));
  and1  g1999(.dina(new_new_n5666__), .dinb(new_new_n5668__), .dout(new_new_n4184__));
  or1   g2000(.dina(new_new_n5609__), .dinb(new_new_n5611__), .dout(new_new_n4185__));
  or1   g2001(.dina(new_new_n5613__), .dinb(new_new_n5615__), .dout(new_new_n4186__));
  or1   g2002(.dina(new_new_n5619__), .dinb(new_new_n5621__), .dout(new_new_n4187__));
  or1   g2003(.dina(new_new_n5623__), .dinb(new_new_n5625__), .dout(new_new_n4188__));
  and1  g2004(.dina(new_new_n5638__), .dinb(new_new_n5641__), .dout(new_new_n4189__));
  and1  g2005(.dina(new_new_n5645__), .dinb(new_new_n5648__), .dout(new_new_n4190__));
  or1   g2006(.dina(new_new_n5629__), .dinb(new_new_n5632__), .dout(new_new_n4191__));
  and1  g2007(.dina(new_new_n5638__), .dinb(new_new_n5650__), .dout(new_new_n4192__));
  and1  g2008(.dina(new_new_n5645__), .dinb(new_new_n5652__), .dout(new_new_n4193__));
  or1   g2009(.dina(new_new_n5629__), .dinb(new_new_n5634__), .dout(new_new_n4194__));
  and1  g2010(.dina(new_new_n5604__), .dinb(new_new_n5607__), .dout(new_new_n4195__));
  and1  g2011(.dina(new_new_n5617__), .dinb(new_new_n5607__), .dout(new_new_n4196__));
  or1   g2012(.dina(new_new_n5654__), .dinb(new_new_n5656__), .dout(new_new_n4197__));
  or1   g2013(.dina(new_new_n5658__), .dinb(new_new_n5660__), .dout(new_new_n4198__));
  or1   g2014(.dina(new_new_n5662__), .dinb(new_new_n5664__), .dout(new_new_n4199__));
  or1   g2015(.dina(new_new_n5666__), .dinb(new_new_n5668__), .dout(new_new_n4200__));
  and1  g2016(.dina(new_new_n5670__), .dinb(new_new_n2318__), .dout(new_new_n4201__));
  and1  g2017(.dina(new_new_n4201__), .dinb(new_new_n5673__), .dout(new_new_n4202__));
  and1  g2018(.dina(new_new_n5676__), .dinb(new_new_n2228__), .dout(new_new_n4203__));
  and1  g2019(.dina(new_new_n4203__), .dinb(new_new_n5673__), .dout(new_new_n4204__));
  and1  g2020(.dina(new_new_n5670__), .dinb(new_new_n2288__), .dout(new_new_n4205__));
  and1  g2021(.dina(new_new_n4205__), .dinb(new_new_n5679__), .dout(new_new_n4206__));
  and1  g2022(.dina(new_new_n5676__), .dinb(new_new_n2258__), .dout(new_new_n4207__));
  and1  g2023(.dina(new_new_n4207__), .dinb(new_new_n5679__), .dout(new_new_n4208__));
  or1   g2024(.dina(new_new_n4204__), .dinb(new_new_n4202__), .dout(new_new_n4209__));
  or1   g2025(.dina(new_new_n4209__), .dinb(new_new_n4206__), .dout(new_new_n4210__));
  or1   g2026(.dina(new_new_n4210__), .dinb(new_new_n4208__), .dout(new_new_n4211__));
  and1  g2027(.dina(new_new_n5671__), .dinb(new_new_n2322__), .dout(new_new_n4212__));
  and1  g2028(.dina(new_new_n4212__), .dinb(new_new_n5674__), .dout(new_new_n4213__));
  and1  g2029(.dina(new_new_n5677__), .dinb(new_new_n2232__), .dout(new_new_n4214__));
  and1  g2030(.dina(new_new_n4214__), .dinb(new_new_n5674__), .dout(new_new_n4215__));
  and1  g2031(.dina(new_new_n5671__), .dinb(new_new_n2292__), .dout(new_new_n4216__));
  and1  g2032(.dina(new_new_n4216__), .dinb(new_new_n5680__), .dout(new_new_n4217__));
  and1  g2033(.dina(new_new_n5677__), .dinb(new_new_n2262__), .dout(new_new_n4218__));
  and1  g2034(.dina(new_new_n4218__), .dinb(new_new_n5680__), .dout(new_new_n4219__));
  or1   g2035(.dina(new_new_n4215__), .dinb(new_new_n4213__), .dout(new_new_n4220__));
  or1   g2036(.dina(new_new_n4220__), .dinb(new_new_n4217__), .dout(new_new_n4221__));
  or1   g2037(.dina(new_new_n4221__), .dinb(new_new_n4219__), .dout(new_new_n4222__));
  or1   g2038(.dina(new_new_n5681__), .dinb(new_new_n5682__), .dout(new_new_n4223__));
  or1   g2039(.dina(new_new_n5681__), .dinb(new_new_n5683__), .dout(new_new_n4224__));
  or1   g2040(.dina(new_new_n5682__), .dinb(new_new_n5684__), .dout(new_new_n4225__));
  or1   g2041(.dina(new_new_n5684__), .dinb(new_new_n5683__), .dout(new_new_n4226__));
  and1  g2042(.dina(new_new_n4224__), .dinb(new_new_n4223__), .dout(new_new_n4227__));
  and1  g2043(.dina(new_new_n4227__), .dinb(new_new_n4225__), .dout(new_new_n4228__));
  and1  g2044(.dina(new_new_n4228__), .dinb(new_new_n4226__), .dout(new_new_n4229__));
  and1  g2045(.dina(new_new_n5114__), .dinb(new_new_n2334__), .dout(new_new_n4230__));
  and1  g2046(.dina(new_new_n4230__), .dinb(new_new_n5121__), .dout(new_new_n4231__));
  and1  g2047(.dina(new_new_n5128__), .dinb(new_new_n2244__), .dout(new_new_n4232__));
  and1  g2048(.dina(new_new_n4232__), .dinb(new_new_n5121__), .dout(new_new_n4233__));
  and1  g2049(.dina(new_new_n5114__), .dinb(new_new_n2304__), .dout(new_new_n4234__));
  and1  g2050(.dina(new_new_n4234__), .dinb(new_new_n5135__), .dout(new_new_n4235__));
  and1  g2051(.dina(new_new_n5128__), .dinb(new_new_n2274__), .dout(new_new_n4236__));
  and1  g2052(.dina(new_new_n4236__), .dinb(new_new_n5135__), .dout(new_new_n4237__));
  or1   g2053(.dina(new_new_n4233__), .dinb(new_new_n4231__), .dout(new_new_n4238__));
  or1   g2054(.dina(new_new_n4238__), .dinb(new_new_n4235__), .dout(new_new_n4239__));
  or1   g2055(.dina(new_new_n4239__), .dinb(new_new_n4237__), .dout(new_new_n4240__));
  and1  g2056(.dina(new_new_n4160__), .dinb(new_new_n5599__), .dout(new_new_n4241__));
  and1  g2057(.dina(new_new_n5595__), .dinb(new_new_n5685__), .dout(new_new_n4242__));
  or1   g2058(.dina(new_new_n4242__), .dinb(new_new_n4241__), .dout(new_new_n4243__));
  or1   g2059(.dina(new_new_n5686__), .dinb(new_new_n5689__), .dout(new_new_n4244__));
  or1   g2060(.dina(new_new_n3559__), .dinb(new_new_n5692__), .dout(new_new_n4245__));
  and1  g2061(.dina(new_new_n4245__), .dinb(new_new_n4244__), .dout(new_new_n4246__));
  and1  g2062(.dina(new_new_n4167__), .dinb(new_new_n5599__), .dout(new_new_n4247__));
  and1  g2063(.dina(new_new_n5602__), .dinb(new_new_n5685__), .dout(new_new_n4248__));
  or1   g2064(.dina(new_new_n4248__), .dinb(new_new_n4247__), .dout(new_new_n4249__));
  or1   g2065(.dina(new_new_n5693__), .dinb(new_new_n5689__), .dout(new_new_n4250__));
  or1   g2066(.dina(new_new_n3565__), .dinb(new_new_n5692__), .dout(new_new_n4251__));
  and1  g2067(.dina(new_new_n4251__), .dinb(new_new_n4250__), .dout(new_new_n4252__));
  or1   g2068(.dina(new_new_n5212__), .dinb(new_new_n5695__), .dout(new_new_n4253__));
  or1   g2069(.dina(new_new_n5201__), .dinb(new_new_n5698__), .dout(new_new_n4254__));
  and1  g2070(.dina(new_new_n4254__), .dinb(new_new_n4253__), .dout(new_new_n4255__));
  or1   g2071(.dina(new_new_n4255__), .dinb(new_new_n5702__), .dout(new_new_n4256__));
  or1   g2072(.dina(new_new_n5239__), .dinb(new_new_n5695__), .dout(new_new_n4257__));
  or1   g2073(.dina(new_new_n5229__), .dinb(new_new_n5698__), .dout(new_new_n4258__));
  and1  g2074(.dina(new_new_n4258__), .dinb(new_new_n4257__), .dout(new_new_n4259__));
  or1   g2075(.dina(new_new_n4259__), .dinb(new_new_n5702__), .dout(new_new_n4260__));
  and1  g2076(.dina(new_new_n5706__), .dinb(new_new_n2096__), .dout(new_new_n4261__));
  and1  g2077(.dina(new_new_n4261__), .dinb(new_new_n5714__), .dout(new_new_n4262__));
  and1  g2078(.dina(new_new_n5706__), .dinb(new_new_n2098__), .dout(new_new_n4263__));
  and1  g2079(.dina(new_new_n4263__), .dinb(new_new_n5714__), .dout(new_new_n4264__));
  and1  g2080(.dina(new_new_n5707__), .dinb(new_new_n2158__), .dout(new_new_n4265__));
  and1  g2081(.dina(new_new_n4265__), .dinb(new_new_n5724__), .dout(new_new_n4266__));
  and1  g2082(.dina(new_new_n5707__), .dinb(new_new_n2160__), .dout(new_new_n4267__));
  and1  g2083(.dina(new_new_n4267__), .dinb(new_new_n5724__), .dout(new_new_n4268__));
  and1  g2084(.dina(new_new_n5732__), .dinb(new_new_n2128__), .dout(new_new_n4269__));
  and1  g2085(.dina(new_new_n4269__), .dinb(new_new_n5725__), .dout(new_new_n4270__));
  and1  g2086(.dina(new_new_n5725__), .dinb(new_new_n5732__), .dout(new_new_n4271__));
  and1  g2087(.dina(new_new_n5495__), .dinb(new_new_n2238__), .dout(new_new_n4272__));
  and1  g2088(.dina(new_new_n4272__), .dinb(new_new_n5487__), .dout(new_new_n4273__));
  and1  g2089(.dina(new_new_n5495__), .dinb(new_new_n2268__), .dout(new_new_n4274__));
  and1  g2090(.dina(new_new_n4274__), .dinb(new_new_n5500__), .dout(new_new_n4275__));
  and1  g2091(.dina(new_new_n5478__), .dinb(new_new_n2298__), .dout(new_new_n4276__));
  and1  g2092(.dina(new_new_n4276__), .dinb(new_new_n5500__), .dout(new_new_n4277__));
  and1  g2093(.dina(new_new_n5733__), .dinb(new_new_n2190__), .dout(new_new_n4278__));
  and1  g2094(.dina(new_new_n4278__), .dinb(new_new_n5715__), .dout(new_new_n4279__));
  and1  g2095(.dina(new_new_n5733__), .dinb(new_new_n2192__), .dout(new_new_n4280__));
  and1  g2096(.dina(new_new_n4280__), .dinb(new_new_n5715__), .dout(new_new_n4281__));
  and1  g2097(.dina(new_new_n5735__), .dinb(new_new_n2194__), .dout(new_new_n4282__));
  and1  g2098(.dina(new_new_n4282__), .dinb(new_new_n5717__), .dout(new_new_n4283__));
  and1  g2099(.dina(new_new_n5709__), .dinb(new_new_n2100__), .dout(new_new_n4284__));
  and1  g2100(.dina(new_new_n4284__), .dinb(new_new_n5717__), .dout(new_new_n4285__));
  and1  g2101(.dina(new_new_n5735__), .dinb(new_new_n2130__), .dout(new_new_n4286__));
  and1  g2102(.dina(new_new_n4286__), .dinb(new_new_n5727__), .dout(new_new_n4287__));
  and1  g2103(.dina(new_new_n5709__), .dinb(new_new_n2162__), .dout(new_new_n4288__));
  and1  g2104(.dina(new_new_n4288__), .dinb(new_new_n5727__), .dout(new_new_n4289__));
  or1   g2105(.dina(new_new_n4285__), .dinb(new_new_n4283__), .dout(new_new_n4290__));
  or1   g2106(.dina(new_new_n4290__), .dinb(new_new_n4287__), .dout(new_new_n4291__));
  or1   g2107(.dina(new_new_n4291__), .dinb(new_new_n4289__), .dout(new_new_n4292__));
  and1  g2108(.dina(new_new_n5736__), .dinb(new_new_n2196__), .dout(new_new_n4293__));
  and1  g2109(.dina(new_new_n4293__), .dinb(new_new_n5718__), .dout(new_new_n4294__));
  and1  g2110(.dina(new_new_n5710__), .dinb(new_new_n2102__), .dout(new_new_n4295__));
  and1  g2111(.dina(new_new_n4295__), .dinb(new_new_n5718__), .dout(new_new_n4296__));
  and1  g2112(.dina(new_new_n5736__), .dinb(new_new_n2132__), .dout(new_new_n4297__));
  and1  g2113(.dina(new_new_n4297__), .dinb(new_new_n5728__), .dout(new_new_n4298__));
  and1  g2114(.dina(new_new_n5710__), .dinb(new_new_n2164__), .dout(new_new_n4299__));
  and1  g2115(.dina(new_new_n4299__), .dinb(new_new_n5728__), .dout(new_new_n4300__));
  or1   g2116(.dina(new_new_n4296__), .dinb(new_new_n4294__), .dout(new_new_n4301__));
  or1   g2117(.dina(new_new_n4301__), .dinb(new_new_n4298__), .dout(new_new_n4302__));
  or1   g2118(.dina(new_new_n4302__), .dinb(new_new_n4300__), .dout(new_new_n4303__));
  and1  g2119(.dina(new_new_n5478__), .dinb(new_new_n2328__), .dout(new_new_n4304__));
  and1  g2120(.dina(new_new_n4304__), .dinb(new_new_n5487__), .dout(new_new_n4305__));
  buf1  g2121(.din(new_new_n5049__), .dout(G2531));
  buf1  g2122(.din(new_new_n5050__), .dout(G2532));
  buf1  g2123(.din(G2532), .dout(G2533));
  buf1  g2124(.din(new_new_n5740__), .dout(G2534));
  buf1  g2125(.din(G2534), .dout(G2535));
  buf1  g2126(.din(new_new_n5742__), .dout(G2536));
  buf1  g2127(.din(G2536), .dout(G2537));
  buf1  g2128(.din(new_new_n5741__), .dout(G2538));
  buf1  g2129(.din(new_new_n5060__), .dout(G2539));
  buf1  g2130(.din(new_new_n5057__), .dout(G2540));
  buf1  g2131(.din(new_new_n5058__), .dout(G2541));
  buf1  g2132(.din(new_new_n5059__), .dout(G2542));
  buf1  g2133(.din(new_new_n5056__), .dout(G2543));
  buf1  g2134(.din(new_new_n5053__), .dout(G2544));
  buf1  g2135(.din(new_new_n5054__), .dout(G2545));
  buf1  g2136(.din(new_new_n5055__), .dout(G2546));
  buf1  g2137(.din(new_new_n3246__), .dout(G2547));
  buf1  g2138(.din(new_new_n3248__), .dout(G2548));
  buf1  g2139(.din(new_new_n2342__), .dout(G2549));
  buf1  g2140(.din(new_new_n3249__), .dout(G2550));
  buf1  g2141(.din(new_new_n5051__), .dout(G2551));
  buf1  g2142(.din(new_new_n3251__), .dout(G2552));
  buf1  g2143(.din(new_new_n3252__), .dout(G2553));
  buf1  g2144(.din(new_new_n5743__), .dout(G2554));
  buf1  g2145(.din(G2554), .dout(G2555));
  buf1  g2146(.din(new_new_n5070__), .dout(G2556));
  buf1  g2147(.din(new_new_n2541__), .dout(G2557));
  buf1  g2148(.din(new_new_n2573__), .dout(G2558));
  buf1  g2149(.din(new_new_n2543__), .dout(G2559));
  buf1  g2150(.din(new_new_n2545__), .dout(G2560));
  buf1  g2151(.din(new_new_n5081__), .dout(G2561));
  buf1  g2152(.din(new_new_n2557__), .dout(G2562));
  buf1  g2153(.din(new_new_n3264__), .dout(G2563));
  buf1  g2154(.din(new_new_n3267__), .dout(G2564));
  buf1  g2155(.din(new_new_n3270__), .dout(G2565));
  buf1  g2156(.din(new_new_n5080__), .dout(G2566));
  buf1  g2157(.din(new_new_n5075__), .dout(G2567));
  buf1  g2158(.din(new_new_n2550__), .dout(G2568));
  buf1  g2159(.din(new_new_n2548__), .dout(G2569));
  buf1  g2160(.din(new_new_n2554__), .dout(G2570));
  buf1  g2161(.din(new_new_n2552__), .dout(G2571));
  buf1  g2162(.din(new_new_n2560__), .dout(G2572));
  buf1  g2163(.din(new_new_n5744__), .dout(G2573));
  buf1  g2164(.din(G2573), .dout(G2574));
  buf1  g2165(.din(new_new_n5745__), .dout(G2575));
  buf1  g2166(.din(G2575), .dout(G2576));
  buf1  g2167(.din(new_new_n3279__), .dout(G2577));
  buf1  g2168(.din(new_new_n5746__), .dout(G2578));
  buf1  g2169(.din(G2578), .dout(G2579));
  buf1  g2170(.din(new_new_n3291__), .dout(G2580));
  not1  g2171(.din(new_new_n5098__), .dout(G2581));
  buf1  g2172(.din(new_new_n5096__), .dout(G2582));
  buf1  g2173(.din(new_new_n5097__), .dout(G2583));
  buf1  g2174(.din(new_new_n5747__), .dout(G2584));
  buf1  g2175(.din(G2584), .dout(G2585));
  buf1  g2176(.din(new_new_n3408__), .dout(G2586));
  not1  g2177(.din(new_new_n5095__), .dout(G2587));
  buf1  g2178(.din(new_new_n5748__), .dout(G2588));
  buf1  g2179(.din(G2588), .dout(G2589));
  not1  g2180(.din(new_new_n5094__), .dout(G2590));
  buf1  g2181(.din(new_new_n2706__), .dout(G2591));
  buf1  g2182(.din(new_new_n5099__), .dout(G2592));
  buf1  g2183(.din(new_new_n5749__), .dout(G2593));
  buf1  g2184(.din(G2593), .dout(G2594));
  buf1  g2185(.din(new_new_n1576__), .dout(n8268));
  buf1  g2186(.din(new_new_n1890__), .dout(n8271));
  buf1  g2187(.din(new_new_n1892__), .dout(n8274));
  buf1  g2188(.din(new_new_n1894__), .dout(n8277));
  buf1  g2189(.din(new_new_n1578__), .dout(n8280));
  buf1  g2190(.din(new_new_n1898__), .dout(n8283));
  buf1  g2191(.din(new_new_n1900__), .dout(n8286));
  buf1  g2192(.din(new_new_n1902__), .dout(n8289));
  buf1  g2193(.din(new_new_n1580__), .dout(n8292));
  buf1  g2194(.din(new_new_n1906__), .dout(n8295));
  buf1  g2195(.din(new_new_n1908__), .dout(n8298));
  buf1  g2196(.din(new_new_n1910__), .dout(n8301));
  buf1  g2197(.din(new_new_n1582__), .dout(n8304));
  buf1  g2198(.din(new_new_n1914__), .dout(n8307));
  buf1  g2199(.din(new_new_n1916__), .dout(n8310));
  buf1  g2200(.din(new_new_n1584__), .dout(n8313));
  buf1  g2201(.din(new_new_n1920__), .dout(n8316));
  buf1  g2202(.din(new_new_n1922__), .dout(n8319));
  buf1  g2203(.din(new_new_n1586__), .dout(n8322));
  buf1  g2204(.din(new_new_n1926__), .dout(n8325));
  buf1  g2205(.din(new_new_n1928__), .dout(n8328));
  buf1  g2206(.din(new_new_n1588__), .dout(n8331));
  buf1  g2207(.din(new_new_n1932__), .dout(n8334));
  buf1  g2208(.din(new_new_n1934__), .dout(n8337));
  buf1  g2209(.din(new_new_n1936__), .dout(n8340));
  buf1  g2210(.din(new_new_n1590__), .dout(n8343));
  buf1  g2211(.din(new_new_n1592__), .dout(n8346));
  buf1  g2212(.din(new_new_n1942__), .dout(n8349));
  buf1  g2213(.din(new_new_n1944__), .dout(n8352));
  buf1  g2214(.din(new_new_n1946__), .dout(n8355));
  buf1  g2215(.din(new_new_n1594__), .dout(n8358));
  buf1  g2216(.din(new_new_n1950__), .dout(n8361));
  buf1  g2217(.din(new_new_n1952__), .dout(n8364));
  buf1  g2218(.din(new_new_n1954__), .dout(n8367));
  buf1  g2219(.din(new_new_n1596__), .dout(n8370));
  buf1  g2220(.din(new_new_n1958__), .dout(n8373));
  buf1  g2221(.din(new_new_n1960__), .dout(n8376));
  buf1  g2222(.din(new_new_n1962__), .dout(n8379));
  buf1  g2223(.din(new_new_n1598__), .dout(n8382));
  buf1  g2224(.din(new_new_n1966__), .dout(n8385));
  buf1  g2225(.din(new_new_n1968__), .dout(n8388));
  buf1  g2226(.din(new_new_n1600__), .dout(n8391));
  buf1  g2227(.din(new_new_n1972__), .dout(n8394));
  buf1  g2228(.din(new_new_n1974__), .dout(n8397));
  buf1  g2229(.din(new_new_n1602__), .dout(n8400));
  buf1  g2230(.din(new_new_n1978__), .dout(n8403));
  buf1  g2231(.din(new_new_n1980__), .dout(n8406));
  buf1  g2232(.din(new_new_n1604__), .dout(n8409));
  buf1  g2233(.din(new_new_n1984__), .dout(n8412));
  buf1  g2234(.din(new_new_n1986__), .dout(n8415));
  buf1  g2235(.din(new_new_n1606__), .dout(n8418));
  buf1  g2236(.din(new_new_n1990__), .dout(n8421));
  buf1  g2237(.din(new_new_n1992__), .dout(n8424));
  buf1  g2238(.din(new_new_n1608__), .dout(n8427));
  buf1  g2239(.din(new_new_n1996__), .dout(n8430));
  buf1  g2240(.din(new_new_n1998__), .dout(n8433));
  buf1  g2241(.din(new_new_n1610__), .dout(n8436));
  buf1  g2242(.din(new_new_n2002__), .dout(n8439));
  buf1  g2243(.din(new_new_n2004__), .dout(n8442));
  buf1  g2244(.din(new_new_n1612__), .dout(n8445));
  buf1  g2245(.din(new_new_n2008__), .dout(n8448));
  buf1  g2246(.din(new_new_n2010__), .dout(n8451));
  buf1  g2247(.din(new_new_n1614__), .dout(n8454));
  buf1  g2248(.din(new_new_n2014__), .dout(n8457));
  buf1  g2249(.din(new_new_n2016__), .dout(n8460));
  buf1  g2250(.din(new_new_n1616__), .dout(n8463));
  buf1  g2251(.din(new_new_n2020__), .dout(n8466));
  buf1  g2252(.din(new_new_n2022__), .dout(n8469));
  buf1  g2253(.din(new_new_n1618__), .dout(n8472));
  buf1  g2254(.din(new_new_n2026__), .dout(n8475));
  buf1  g2255(.din(new_new_n2028__), .dout(n8478));
  buf1  g2256(.din(new_new_n2030__), .dout(n8481));
  buf1  g2257(.din(new_new_n1620__), .dout(n8484));
  buf1  g2258(.din(new_new_n2034__), .dout(n8487));
  buf1  g2259(.din(new_new_n2036__), .dout(n8490));
  buf1  g2260(.din(new_new_n1622__), .dout(n8493));
  buf1  g2261(.din(new_new_n2040__), .dout(n8496));
  buf1  g2262(.din(new_new_n2042__), .dout(n8499));
  buf1  g2263(.din(new_new_n1624__), .dout(n8502));
  buf1  g2264(.din(new_new_n2046__), .dout(n8505));
  buf1  g2265(.din(new_new_n2048__), .dout(n8508));
  buf1  g2266(.din(new_new_n1626__), .dout(n8511));
  buf1  g2267(.din(new_new_n2052__), .dout(n8514));
  buf1  g2268(.din(new_new_n2054__), .dout(n8517));
  buf1  g2269(.din(new_new_n1628__), .dout(n8520));
  buf1  g2270(.din(new_new_n2058__), .dout(n8523));
  buf1  g2271(.din(new_new_n2060__), .dout(n8526));
  buf1  g2272(.din(new_new_n1630__), .dout(n8529));
  buf1  g2273(.din(new_new_n2064__), .dout(n8532));
  buf1  g2274(.din(new_new_n2066__), .dout(n8535));
  buf1  g2275(.din(new_new_n2068__), .dout(n8538));
  buf1  g2276(.din(new_new_n1632__), .dout(n8541));
  buf1  g2277(.din(new_new_n2072__), .dout(n8544));
  buf1  g2278(.din(new_new_n2074__), .dout(n8547));
  buf1  g2279(.din(new_new_n2076__), .dout(n8550));
  buf1  g2280(.din(new_new_n1634__), .dout(n8553));
  buf1  g2281(.din(new_new_n1636__), .dout(n8556));
  buf1  g2282(.din(new_new_n2082__), .dout(n8559));
  buf1  g2283(.din(new_new_n1638__), .dout(n8562));
  buf1  g2284(.din(new_new_n2086__), .dout(n8565));
  buf1  g2285(.din(new_new_n2088__), .dout(n8568));
  buf1  g2286(.din(new_new_n2090__), .dout(n8571));
  buf1  g2287(.din(new_new_n1640__), .dout(n8574));
  buf1  g2288(.din(new_new_n1642__), .dout(n8577));
  buf1  g2289(.din(new_new_n1644__), .dout(n8580));
  buf1  g2290(.din(new_new_n1646__), .dout(n8583));
  buf1  g2291(.din(new_new_n1648__), .dout(n8586));
  buf1  g2292(.din(new_new_n1650__), .dout(n8589));
  buf1  g2293(.din(new_new_n1652__), .dout(n8592));
  buf1  g2294(.din(new_new_n1654__), .dout(n8595));
  buf1  g2295(.din(new_new_n1656__), .dout(n8598));
  buf1  g2296(.din(new_new_n2110__), .dout(n8601));
  buf1  g2297(.din(new_new_n1658__), .dout(n8604));
  buf1  g2298(.din(new_new_n2114__), .dout(n8607));
  buf1  g2299(.din(new_new_n1660__), .dout(n8610));
  buf1  g2300(.din(new_new_n2118__), .dout(n8613));
  buf1  g2301(.din(new_new_n2120__), .dout(n8616));
  buf1  g2302(.din(new_new_n2122__), .dout(n8619));
  buf1  g2303(.din(new_new_n1662__), .dout(n8622));
  buf1  g2304(.din(new_new_n1664__), .dout(n8625));
  buf1  g2305(.din(new_new_n1666__), .dout(n8628));
  buf1  g2306(.din(new_new_n1668__), .dout(n8631));
  buf1  g2307(.din(new_new_n1670__), .dout(n8634));
  buf1  g2308(.din(new_new_n1672__), .dout(n8637));
  buf1  g2309(.din(new_new_n1674__), .dout(n8640));
  buf1  g2310(.din(new_new_n1676__), .dout(n8643));
  buf1  g2311(.din(new_new_n2140__), .dout(n8646));
  buf1  g2312(.din(new_new_n1678__), .dout(n8649));
  buf1  g2313(.din(new_new_n2144__), .dout(n8652));
  buf1  g2314(.din(new_new_n1680__), .dout(n8655));
  buf1  g2315(.din(new_new_n2148__), .dout(n8658));
  buf1  g2316(.din(new_new_n2150__), .dout(n8661));
  buf1  g2317(.din(new_new_n2152__), .dout(n8664));
  buf1  g2318(.din(new_new_n1682__), .dout(n8667));
  buf1  g2319(.din(new_new_n1684__), .dout(n8670));
  buf1  g2320(.din(new_new_n1686__), .dout(n8673));
  buf1  g2321(.din(new_new_n1688__), .dout(n8676));
  buf1  g2322(.din(new_new_n1690__), .dout(n8679));
  buf1  g2323(.din(new_new_n1692__), .dout(n8682));
  buf1  g2324(.din(new_new_n1694__), .dout(n8685));
  buf1  g2325(.din(new_new_n1696__), .dout(n8688));
  buf1  g2326(.din(new_new_n1698__), .dout(n8691));
  buf1  g2327(.din(new_new_n2172__), .dout(n8694));
  buf1  g2328(.din(new_new_n1700__), .dout(n8697));
  buf1  g2329(.din(new_new_n2176__), .dout(n8700));
  buf1  g2330(.din(new_new_n1702__), .dout(n8703));
  buf1  g2331(.din(new_new_n2180__), .dout(n8706));
  buf1  g2332(.din(new_new_n2182__), .dout(n8709));
  buf1  g2333(.din(new_new_n2184__), .dout(n8712));
  buf1  g2334(.din(new_new_n1704__), .dout(n8715));
  buf1  g2335(.din(new_new_n1706__), .dout(n8718));
  buf1  g2336(.din(new_new_n1708__), .dout(n8721));
  buf1  g2337(.din(new_new_n1710__), .dout(n8724));
  buf1  g2338(.din(new_new_n1712__), .dout(n8727));
  buf1  g2339(.din(new_new_n1714__), .dout(n8730));
  buf1  g2340(.din(new_new_n1716__), .dout(n8733));
  buf1  g2341(.din(new_new_n1718__), .dout(n8736));
  buf1  g2342(.din(new_new_n1720__), .dout(n8739));
  buf1  g2343(.din(new_new_n2204__), .dout(n8742));
  buf1  g2344(.din(new_new_n1722__), .dout(n8745));
  buf1  g2345(.din(new_new_n2208__), .dout(n8748));
  buf1  g2346(.din(new_new_n2210__), .dout(n8751));
  buf1  g2347(.din(new_new_n2212__), .dout(n8754));
  buf1  g2348(.din(new_new_n1724__), .dout(n8757));
  buf1  g2349(.din(new_new_n1726__), .dout(n8760));
  buf1  g2350(.din(new_new_n2218__), .dout(n8763));
  buf1  g2351(.din(new_new_n2220__), .dout(n8766));
  buf1  g2352(.din(new_new_n2222__), .dout(n8769));
  buf1  g2353(.din(new_new_n1728__), .dout(n8772));
  buf1  g2354(.din(new_new_n2226__), .dout(n8775));
  buf1  g2355(.din(new_new_n1730__), .dout(n8778));
  buf1  g2356(.din(new_new_n2230__), .dout(n8781));
  buf1  g2357(.din(new_new_n1736__), .dout(n8784));
  buf1  g2358(.din(new_new_n2234__), .dout(n8787));
  buf1  g2359(.din(new_new_n1738__), .dout(n8790));
  buf1  g2360(.din(new_new_n1740__), .dout(n8793));
  buf1  g2361(.din(new_new_n1742__), .dout(n8796));
  buf1  g2362(.din(new_new_n2242__), .dout(n8799));
  buf1  g2363(.din(new_new_n1744__), .dout(n8802));
  buf1  g2364(.din(new_new_n1746__), .dout(n8805));
  buf1  g2365(.din(new_new_n2248__), .dout(n8808));
  buf1  g2366(.din(new_new_n2250__), .dout(n8811));
  buf1  g2367(.din(new_new_n2252__), .dout(n8814));
  buf1  g2368(.din(new_new_n1748__), .dout(n8817));
  buf1  g2369(.din(new_new_n2256__), .dout(n8820));
  buf1  g2370(.din(new_new_n1750__), .dout(n8823));
  buf1  g2371(.din(new_new_n2260__), .dout(n8826));
  buf1  g2372(.din(new_new_n1756__), .dout(n8829));
  buf1  g2373(.din(new_new_n2264__), .dout(n8832));
  buf1  g2374(.din(new_new_n1758__), .dout(n8835));
  buf1  g2375(.din(new_new_n1760__), .dout(n8838));
  buf1  g2376(.din(new_new_n1762__), .dout(n8841));
  buf1  g2377(.din(new_new_n2272__), .dout(n8844));
  buf1  g2378(.din(new_new_n1764__), .dout(n8847));
  buf1  g2379(.din(new_new_n1766__), .dout(n8850));
  buf1  g2380(.din(new_new_n2278__), .dout(n8853));
  buf1  g2381(.din(new_new_n2280__), .dout(n8856));
  buf1  g2382(.din(new_new_n2282__), .dout(n8859));
  buf1  g2383(.din(new_new_n1768__), .dout(n8862));
  buf1  g2384(.din(new_new_n2286__), .dout(n8865));
  buf1  g2385(.din(new_new_n1770__), .dout(n8868));
  buf1  g2386(.din(new_new_n2290__), .dout(n8871));
  buf1  g2387(.din(new_new_n1776__), .dout(n8874));
  buf1  g2388(.din(new_new_n2294__), .dout(n8877));
  buf1  g2389(.din(new_new_n1778__), .dout(n8880));
  buf1  g2390(.din(new_new_n1780__), .dout(n8883));
  buf1  g2391(.din(new_new_n1782__), .dout(n8886));
  buf1  g2392(.din(new_new_n2302__), .dout(n8889));
  buf1  g2393(.din(new_new_n1784__), .dout(n8892));
  buf1  g2394(.din(new_new_n1786__), .dout(n8895));
  buf1  g2395(.din(new_new_n2308__), .dout(n8898));
  buf1  g2396(.din(new_new_n2310__), .dout(n8901));
  buf1  g2397(.din(new_new_n2312__), .dout(n8904));
  buf1  g2398(.din(new_new_n1788__), .dout(n8907));
  buf1  g2399(.din(new_new_n2316__), .dout(n8910));
  buf1  g2400(.din(new_new_n1790__), .dout(n8913));
  buf1  g2401(.din(new_new_n2320__), .dout(n8916));
  buf1  g2402(.din(new_new_n1796__), .dout(n8919));
  buf1  g2403(.din(new_new_n2324__), .dout(n8922));
  buf1  g2404(.din(new_new_n1798__), .dout(n8925));
  buf1  g2405(.din(new_new_n1800__), .dout(n8928));
  buf1  g2406(.din(new_new_n1802__), .dout(n8931));
  buf1  g2407(.din(new_new_n2332__), .dout(n8934));
  buf1  g2408(.din(new_new_n1804__), .dout(n8937));
  buf1  g2409(.din(new_new_n2336__), .dout(n8940));
  buf1  g2410(.din(new_new_n2338__), .dout(n8943));
  buf1  g2411(.din(new_new_n2340__), .dout(n8946));
  buf1  g2412(.din(new_new_n1806__), .dout(n8949));
  buf1  g2413(.din(new_new_n2344__), .dout(n8952));
  buf1  g2414(.din(new_new_n2346__), .dout(n8955));
  buf1  g2415(.din(new_new_n2348__), .dout(n8958));
  buf1  g2416(.din(new_new_n1808__), .dout(n8961));
  buf1  g2417(.din(new_new_n1810__), .dout(n8964));
  buf1  g2418(.din(new_new_n2354__), .dout(n8967));
  buf1  g2419(.din(new_new_n2356__), .dout(n8970));
  buf1  g2420(.din(new_new_n1812__), .dout(n8973));
  buf1  g2421(.din(new_new_n2360__), .dout(n8976));
  buf1  g2422(.din(new_new_n2362__), .dout(n8979));
  buf1  g2423(.din(new_new_n2364__), .dout(n8982));
  buf1  g2424(.din(new_new_n1814__), .dout(n8985));
  buf1  g2425(.din(new_new_n1816__), .dout(n8988));
  buf1  g2426(.din(new_new_n2370__), .dout(n8991));
  buf1  g2427(.din(new_new_n2372__), .dout(n8994));
  buf1  g2428(.din(new_new_n2374__), .dout(n8997));
  buf1  g2429(.din(new_new_n1818__), .dout(n9000));
  buf1  g2430(.din(new_new_n2378__), .dout(n9003));
  buf1  g2431(.din(new_new_n2380__), .dout(n9006));
  buf1  g2432(.din(new_new_n2382__), .dout(n9009));
  buf1  g2433(.din(new_new_n1820__), .dout(n9012));
  buf1  g2434(.din(new_new_n2386__), .dout(n9015));
  buf1  g2435(.din(new_new_n2388__), .dout(n9018));
  buf1  g2436(.din(new_new_n2390__), .dout(n9021));
  buf1  g2437(.din(new_new_n1822__), .dout(n9024));
  buf1  g2438(.din(new_new_n2394__), .dout(n9027));
  buf1  g2439(.din(new_new_n2396__), .dout(n9030));
  buf1  g2440(.din(new_new_n2398__), .dout(n9033));
  buf1  g2441(.din(new_new_n1824__), .dout(n9036));
  buf1  g2442(.din(new_new_n2402__), .dout(n9039));
  buf1  g2443(.din(new_new_n1826__), .dout(n9042));
  buf1  g2444(.din(new_new_n1828__), .dout(n9045));
  buf1  g2445(.din(new_new_n1830__), .dout(n9048));
  buf1  g2446(.din(new_new_n1832__), .dout(n9051));
  buf1  g2447(.din(new_new_n2412__), .dout(n9054));
  buf1  g2448(.din(new_new_n1834__), .dout(n9057));
  buf1  g2449(.din(new_new_n1836__), .dout(n9060));
  buf1  g2450(.din(new_new_n1838__), .dout(n9063));
  buf1  g2451(.din(new_new_n2420__), .dout(n9066));
  buf1  g2452(.din(new_new_n1840__), .dout(n9069));
  buf1  g2453(.din(new_new_n2424__), .dout(n9072));
  buf1  g2454(.din(new_new_n1842__), .dout(n9075));
  buf1  g2455(.din(new_new_n2428__), .dout(n9078));
  buf1  g2456(.din(new_new_n1844__), .dout(n9081));
  buf1  g2457(.din(new_new_n2432__), .dout(n9084));
  buf1  g2458(.din(new_new_n1846__), .dout(n9087));
  buf1  g2459(.din(new_new_n2436__), .dout(n9090));
  buf1  g2460(.din(new_new_n1848__), .dout(n9093));
  buf1  g2461(.din(new_new_n2440__), .dout(n9096));
  buf1  g2462(.din(new_new_n2442__), .dout(n9099));
  buf1  g2463(.din(new_new_n2444__), .dout(n9102));
  buf1  g2464(.din(new_new_n1850__), .dout(n9105));
  buf1  g2465(.din(new_new_n1852__), .dout(n9108));
  buf1  g2466(.din(new_new_n5519__), .dout(n9111));
  buf1  g2467(.din(new_new_n1854__), .dout(n9114));
  buf1  g2468(.din(new_new_n2454__), .dout(n9117));
  buf1  g2469(.din(new_new_n5515__), .dout(n9120));
  buf1  g2470(.din(new_new_n1856__), .dout(n9123));
  buf1  g2471(.din(new_new_n5526__), .dout(n9126));
  buf1  g2472(.din(new_new_n1858__), .dout(n9129));
  buf1  g2473(.din(new_new_n5525__), .dout(n9132));
  buf1  g2474(.din(new_new_n1860__), .dout(n9135));
  buf1  g2475(.din(new_new_n2468__), .dout(n9138));
  buf1  g2476(.din(new_new_n2470__), .dout(n9141));
  buf1  g2477(.din(new_new_n5751__), .dout(n9144));
  buf1  g2478(.din(new_new_n1862__), .dout(n9147));
  buf1  g2479(.din(new_new_n2476__), .dout(n9150));
  buf1  g2480(.din(new_new_n2478__), .dout(n9153));
  buf1  g2481(.din(new_new_n5753__), .dout(n9156));
  buf1  g2482(.din(new_new_n1868__), .dout(n9159));
  buf1  g2483(.din(new_new_n2484__), .dout(n9162));
  buf1  g2484(.din(new_new_n2486__), .dout(n9165));
  buf1  g2485(.din(new_new_n2488__), .dout(n9168));
  buf1  g2486(.din(new_new_n1870__), .dout(n9171));
  buf1  g2487(.din(new_new_n2492__), .dout(n9174));
  buf1  g2488(.din(new_new_n1872__), .dout(n9177));
  buf1  g2489(.din(new_new_n2496__), .dout(n9180));
  buf1  g2490(.din(new_new_n1874__), .dout(n9183));
  buf1  g2491(.din(new_new_n2500__), .dout(n9186));
  buf1  g2492(.din(new_new_n1876__), .dout(n9189));
  buf1  g2493(.din(new_new_n2504__), .dout(n9192));
  buf1  g2494(.din(new_new_n1878__), .dout(n9195));
  buf1  g2495(.din(new_new_n2508__), .dout(n9198));
  buf1  g2496(.din(new_new_n1880__), .dout(n9201));
  buf1  g2497(.din(new_new_n2512__), .dout(n9204));
  buf1  g2498(.din(new_new_n1882__), .dout(n9207));
  buf1  g2499(.din(new_new_n2516__), .dout(n9210));
  buf1  g2500(.din(new_new_n2518__), .dout(n9213));
  buf1  g2501(.din(new_new_n1884__), .dout(n9216));
  buf1  g2502(.din(new_new_n2522__), .dout(n9219));
  buf1  g2503(.din(new_new_n2524__), .dout(n9222));
  buf1  g2504(.din(new_new_n1886__), .dout(n9225));
  buf1  g2505(.din(new_new_n2528__), .dout(n9228));
  buf1  g2506(.din(new_new_n2530__), .dout(n9231));
  buf1  g2507(.din(new_new_n1888__), .dout(n9234));
  buf1  g2508(.din(new_new_n2534__), .dout(n9237));
  buf1  g2509(.din(new_new_n2536__), .dout(n9240));
  buf1  g2510(.din(new_new_n5327__), .dout(n9243));
  buf1  g2511(.din(new_new_n5583__), .dout(n9246));
  buf1  g2512(.din(new_new_n5568__), .dout(n9249));
  buf1  g2513(.din(new_new_n5567__), .dout(n9252));
  buf1  g2514(.din(new_new_n2610__), .dout(n9255));
  buf1  g2515(.din(new_new_n2612__), .dout(n9258));
  buf1  g2516(.din(new_new_n2650__), .dout(n9261));
  buf1  g2517(.din(new_new_n2652__), .dout(n9264));
  buf1  g2518(.din(new_new_n5564__), .dout(n9267));
  buf1  g2519(.din(new_new_n5103__), .dout(n9270));
  buf1  g2520(.din(new_new_n2674__), .dout(n9273));
  buf1  g2521(.din(new_new_n2676__), .dout(n9276));
  buf1  g2522(.din(new_new_n2686__), .dout(n9279));
  buf1  g2523(.din(new_new_n5565__), .dout(n9282));
  buf1  g2524(.din(new_new_n2800__), .dout(n9285));
  buf1  g2525(.din(new_new_n5332__), .dout(n9288));
  buf1  g2526(.din(new_new_n5322__), .dout(n9291));
  buf1  g2527(.din(new_new_n5330__), .dout(n9294));
  buf1  g2528(.din(new_new_n2806__), .dout(n9297));
  buf1  g2529(.din(new_new_n5755__), .dout(n9300));
  buf1  g2530(.din(new_new_n5467__), .dout(n9303));
  buf1  g2531(.din(new_new_n5459__), .dout(n9306));
  buf1  g2532(.din(new_new_n5576__), .dout(n9309));
  buf1  g2533(.din(new_new_n5594__), .dout(n9312));
  buf1  g2534(.din(new_new_n5219__), .dout(n9315));
  buf1  g2535(.din(new_new_n5425__), .dout(n9318));
  buf1  g2536(.din(new_new_n5431__), .dout(n9321));
  buf1  g2537(.din(new_new_n5407__), .dout(n9324));
  buf1  g2538(.din(new_new_n5215__), .dout(n9327));
  buf1  g2539(.din(new_new_n5422__), .dout(n9330));
  buf1  g2540(.din(new_new_n5428__), .dout(n9333));
  buf1  g2541(.din(new_new_n5542__), .dout(n9336));
  buf1  g2542(.din(new_new_n5440__), .dout(n9339));
  buf1  g2543(.din(new_new_n5433__), .dout(n9342));
  buf1  g2544(.din(new_new_n5452__), .dout(n9345));
  buf1  g2545(.din(n9303), .dout(n9348));
  buf1  g2546(.din(n9306), .dout(n9351));
  buf1  g2547(.din(new_new_n5756__), .dout(n9354));
  buf1  g2548(.din(new_new_n5384__), .dout(n9357));
  buf1  g2549(.din(new_new_n5402__), .dout(n9360));
  buf1  g2550(.din(new_new_n5757__), .dout(n9363));
  buf1  g2551(.din(new_new_n5696__), .dout(n9366));
  buf1  g2552(.din(new_new_n5758__), .dout(n9369));
  buf1  g2553(.din(n9312), .dout(n9372));
  buf1  g2554(.din(n9315), .dout(n9375));
  buf1  g2555(.din(n9318), .dout(n9378));
  buf1  g2556(.din(n9321), .dout(n9381));
  buf1  g2557(.din(n9324), .dout(n9384));
  buf1  g2558(.din(n9327), .dout(n9387));
  buf1  g2559(.din(n9330), .dout(n9390));
  buf1  g2560(.din(n9333), .dout(n9393));
  buf1  g2561(.din(new_new_n5471__), .dout(n9396));
  buf1  g2562(.din(new_new_n5447__), .dout(n9399));
  buf1  g2563(.din(new_new_n5450__), .dout(n9402));
  buf1  g2564(.din(new_new_n5690__), .dout(n9405));
  buf1  g2565(.din(new_new_n5442__), .dout(n9408));
  buf1  g2566(.din(new_new_n5435__), .dout(n9411));
  buf1  g2567(.din(new_new_n5759__), .dout(n9414));
  buf1  g2568(.din(n9309), .dout(n9417));
  buf1  g2569(.din(n9354), .dout(n9420));
  buf1  g2570(.din(n9357), .dout(n9423));
  buf1  g2571(.din(n9360), .dout(n9426));
  buf1  g2572(.din(n9363), .dout(n9429));
  buf1  g2573(.din(n9366), .dout(n9432));
  buf1  g2574(.din(n9369), .dout(n9435));
  buf1  g2575(.din(new_new_n5762__), .dout(n9438));
  buf1  g2576(.din(new_new_n5601__), .dout(n9441));
  buf1  g2577(.din(new_new_n5472__), .dout(n9444));
  buf1  g2578(.din(n9405), .dout(n9447));
  buf1  g2579(.din(new_new_n5699__), .dout(n9450));
  buf1  g2580(.din(n9414), .dout(n9453));
  buf1  g2581(.din(new_new_n5686__), .dout(n9456));
  buf1  g2582(.din(new_new_n5693__), .dout(n9459));
  buf1  g2583(.din(n9438), .dout(n9462));
  buf1  g2584(.din(n9441), .dout(n9465));
  buf1  g2585(.din(new_new_n5691__), .dout(n9468));
  buf1  g2586(.din(new_new_n5480__), .dout(n9471));
  buf1  g2587(.din(new_new_n5489__), .dout(n9474));
  buf1  g2588(.din(n9471), .dout(n9477));
  buf1  g2589(.din(n9474), .dout(n9480));
  buf1  g2590(.din(n9144), .dout(n9483));
  buf1  g2591(.din(n9156), .dout(n9486));
  not1  g2592(.din(new_new_n5585__), .dout(n9489));
  not1  g2593(.din(new_new_n5584__), .dout(n9492));
  buf1  g2594(.din(new_new_n5764__), .dout(n9495));
  buf1  g2595(.din(new_new_n5765__), .dout(n9498));
  buf1  g2596(.din(new_new_n5335__), .dout(n9501));
  buf1  g2597(.din(new_new_n5337__), .dout(n9504));
  buf1  g2598(.din(new_new_n5766__), .dout(n9507));
  buf1  g2599(.din(new_new_n5767__), .dout(n9510));
  buf1  g2600(.din(new_new_n5768__), .dout(n9513));
  buf1  g2601(.din(new_new_n5769__), .dout(n9516));
  buf1  g2602(.din(new_new_n5770__), .dout(n9519));
  buf1  g2603(.din(new_new_n5771__), .dout(n9522));
  buf1  g2604(.din(n9450), .dout(n9525));
  not1  g2605(.din(new_new_n5603__), .dout(n9528));
  not1  g2606(.din(new_new_n5610__), .dout(n9531));
  not1  g2607(.din(new_new_n5614__), .dout(n9534));
  not1  g2608(.din(new_new_n5616__), .dout(n9537));
  not1  g2609(.din(new_new_n5620__), .dout(n9540));
  not1  g2610(.din(new_new_n5624__), .dout(n9543));
  not1  g2611(.din(new_new_n5631__), .dout(n9546));
  not1  g2612(.din(new_new_n5633__), .dout(n9549));
  buf1  g2613(.din(new_new_n5640__), .dout(n9552));
  buf1  g2614(.din(new_new_n5647__), .dout(n9555));
  buf1  g2615(.din(new_new_n5649__), .dout(n9558));
  buf1  g2616(.din(new_new_n5651__), .dout(n9561));
  not1  g2617(.din(new_new_n5655__), .dout(n9564));
  not1  g2618(.din(new_new_n5659__), .dout(n9567));
  not1  g2619(.din(new_new_n5663__), .dout(n9570));
  not1  g2620(.din(new_new_n5667__), .dout(n9573));
  not1  g2621(.din(new_new_n5608__), .dout(n9576));
  not1  g2622(.din(new_new_n5612__), .dout(n9579));
  not1  g2623(.din(new_new_n5618__), .dout(n9582));
  not1  g2624(.din(new_new_n5622__), .dout(n9585));
  buf1  g2625(.din(new_new_n5639__), .dout(n9588));
  buf1  g2626(.din(new_new_n5646__), .dout(n9591));
  not1  g2627(.din(new_new_n5630__), .dout(n9594));
  buf1  g2628(.din(n9588), .dout(n9597));
  buf1  g2629(.din(n9591), .dout(n9600));
  buf1  g2630(.din(n9594), .dout(n9603));
  buf1  g2631(.din(new_new_n5761__), .dout(n9606));
  not1  g2632(.din(new_new_n5653__), .dout(n9609));
  not1  g2633(.din(new_new_n5657__), .dout(n9612));
  not1  g2634(.din(new_new_n5661__), .dout(n9615));
  not1  g2635(.din(new_new_n5665__), .dout(n9618));
  buf1  g2636(.din(new_new_n5773__), .dout(n9621));
  buf1  g2637(.din(new_new_n5775__), .dout(n9624));
  buf1  g2638(.din(new_new_n5777__), .dout(n9627));
  buf1  g2639(.din(new_new_n5701__), .dout(n9630));
  buf1  g2640(.din(new_new_n5779__), .dout(n9633));
  not1  g2641(.din(new_new_n5782__), .dout(n9636));
  buf1  g2642(.din(n9636), .dout(n9639));
  buf1  g2643(.din(new_new_n5589__), .dout(n9642));
  not1  g2644(.din(new_new_n5586__), .dout(n9645));
  buf1  g2645(.din(new_new_n2080__), .dout(n9648));
  buf1  g2646(.din(new_new_n5738__), .dout(n9651));
  buf1  g2647(.din(new_new_n5720__), .dout(n9654));
  buf1  g2648(.din(new_new_n5588__), .dout(n9657));
  buf1  g2649(.din(new_new_n5785__), .dout(n9660));
  buf1  g2650(.din(new_new_n5786__), .dout(n9663));
  buf1  g2651(.din(new_new_n2626__), .dout(n9666));
  buf1  g2652(.din(new_new_n2628__), .dout(n9669));
  buf1  g2653(.din(new_new_n2630__), .dout(n9672));
  buf1  g2654(.din(new_new_n2632__), .dout(n9675));
  buf1  g2655(.din(new_new_n2634__), .dout(n9678));
  buf1  g2656(.din(new_new_n2636__), .dout(n9681));
  buf1  g2657(.din(new_new_n2638__), .dout(n9684));
  buf1  g2658(.din(new_new_n2640__), .dout(n9687));
  buf1  g2659(.din(new_new_n2658__), .dout(n9690));
  buf1  g2660(.din(new_new_n2660__), .dout(n9693));
  buf1  g2661(.din(new_new_n2662__), .dout(n9696));
  buf1  g2662(.din(new_new_n2664__), .dout(n9699));
  buf1  g2663(.din(new_new_n2666__), .dout(n9702));
  buf1  g2664(.din(new_new_n2668__), .dout(n9705));
  buf1  g2665(.din(new_new_n2680__), .dout(n9708));
  buf1  g2666(.din(new_new_n2728__), .dout(n9711));
  buf1  g2667(.din(n9300), .dout(n9714));
  buf1  g2668(.din(n9336), .dout(n9717));
  buf1  g2669(.din(new_new_n5460__), .dout(n9720));
  not1  g2670(.din(new_new_n4053__), .dout(n9723));
  buf1  g2671(.din(new_new_n4055__), .dout(n9726));
  not1  g2672(.din(new_new_n4072__), .dout(n9729));
  buf1  g2673(.din(new_new_n4074__), .dout(n9732));
  buf1  g2674(.din(new_new_n4076__), .dout(n9735));
  buf1  g2675(.din(new_new_n4078__), .dout(n9738));
  not1  g2676(.din(new_new_n4089__), .dout(n9741));
  buf1  g2677(.din(new_new_n4091__), .dout(n9744));
  not1  g2678(.din(new_new_n4093__), .dout(n9747));
  not1  g2679(.din(new_new_n4095__), .dout(n9750));
  not1  g2680(.din(new_new_n4097__), .dout(n9753));
  not1  g2681(.din(new_new_n4099__), .dout(n9756));
  buf1  g2682(.din(new_new_n5481__), .dout(n9759));
  buf1  g2683(.din(new_new_n5490__), .dout(n9762));
  buf1  g2684(.din(new_new_n4102__), .dout(n9765));
  buf1  g2685(.din(new_new_n4105__), .dout(n9768));
  buf1  g2686(.din(new_new_n4108__), .dout(n9771));
  buf1  g2687(.din(new_new_n4111__), .dout(n9774));
  buf1  g2688(.din(new_new_n4114__), .dout(n9777));
  buf1  g2689(.din(new_new_n4117__), .dout(n9780));
  buf1  g2690(.din(new_new_n4120__), .dout(n9783));
  buf1  g2691(.din(new_new_n4123__), .dout(n9786));
  buf1  g2692(.din(new_new_n4126__), .dout(n9789));
  buf1  g2693(.din(new_new_n4129__), .dout(n9792));
  buf1  g2694(.din(new_new_n4132__), .dout(n9795));
  buf1  g2695(.din(new_new_n4135__), .dout(n9798));
  buf1  g2696(.din(new_new_n4138__), .dout(n9801));
  buf1  g2697(.din(new_new_n4141__), .dout(n9804));
  buf1  g2698(.din(new_new_n4144__), .dout(n9807));
  buf1  g2699(.din(new_new_n4147__), .dout(n9810));
  buf1  g2700(.din(new_new_n5750__), .dout(n9813));
  buf1  g2701(.din(new_new_n5752__), .dout(n9816));
  buf1  g2702(.din(new_new_n4150__), .dout(n9819));
  not1  g2703(.din(new_new_n4151__), .dout(n9822));
  buf1  g2704(.din(n9495), .dout(n9825));
  buf1  g2705(.din(n9498), .dout(n9828));
  buf1  g2706(.din(new_new_n5334__), .dout(n9831));
  buf1  g2707(.din(new_new_n5336__), .dout(n9834));
  buf1  g2708(.din(n9507), .dout(n9837));
  buf1  g2709(.din(n9510), .dout(n9840));
  buf1  g2710(.din(n9513), .dout(n9843));
  buf1  g2711(.din(n9516), .dout(n9846));
  buf1  g2712(.din(n9519), .dout(n9849));
  buf1  g2713(.din(n9522), .dout(n9852));
  buf1  g2714(.din(new_new_n5763__), .dout(n9855));
  buf1  g2715(.din(n9621), .dout(n9858));
  buf1  g2716(.din(n9624), .dout(n9861));
  buf1  g2717(.din(n9627), .dout(n9864));
  buf1  g2718(.din(new_new_n5703__), .dout(n9867));
  buf1  g2719(.din(n9633), .dout(n9870));
  not1  g2720(.din(new_new_n5783__), .dout(n9873));
  buf1  g2721(.din(n9873), .dout(n9876));
  not1  g2722(.din(new_new_n5789__), .dout(n9879));
  buf1  g2723(.din(n9651), .dout(n9882));
  buf1  g2724(.din(n9654), .dout(n9885));
  buf1  g2725(.din(new_new_n2494__), .dout(n9888));
  buf1  g2726(.din(new_new_n2498__), .dout(n9891));
  buf1  g2727(.din(new_new_n2502__), .dout(n9894));
  buf1  g2728(.din(new_new_n2506__), .dout(n9897));
  buf1  g2729(.din(new_new_n5451__), .dout(n9900));
  buf1  g2730(.din(new_new_n5466__), .dout(n9903));
  buf1  g2731(.din(new_new_n5446__), .dout(n9906));
  buf1  g2732(.din(new_new_n5449__), .dout(n9909));
  buf1  g2733(.din(n9408), .dout(n9912));
  buf1  g2734(.din(n9411), .dout(n9915));
  buf1  g2735(.din(n9444), .dout(n9918));
  buf1  g2736(.din(new_new_n4161__), .dout(n9921));
  buf1  g2737(.din(new_new_n4168__), .dout(n9924));
  buf1  g2738(.din(new_new_n5600__), .dout(n9927));
  buf1  g2739(.din(n9468), .dout(n9930));
  buf1  g2740(.din(new_new_n5739__), .dout(n9933));
  buf1  g2741(.din(new_new_n5721__), .dout(n9936));
  not1  g2742(.din(new_new_n4169__), .dout(n9939));
  not1  g2743(.din(new_new_n4170__), .dout(n9942));
  not1  g2744(.din(new_new_n4171__), .dout(n9945));
  not1  g2745(.din(new_new_n4172__), .dout(n9948));
  not1  g2746(.din(new_new_n4173__), .dout(n9951));
  not1  g2747(.din(new_new_n4174__), .dout(n9954));
  not1  g2748(.din(new_new_n4175__), .dout(n9957));
  not1  g2749(.din(new_new_n4176__), .dout(n9960));
  buf1  g2750(.din(new_new_n4177__), .dout(n9963));
  buf1  g2751(.din(new_new_n4178__), .dout(n9966));
  buf1  g2752(.din(new_new_n4179__), .dout(n9969));
  buf1  g2753(.din(new_new_n4180__), .dout(n9972));
  not1  g2754(.din(new_new_n4181__), .dout(n9975));
  not1  g2755(.din(new_new_n4182__), .dout(n9978));
  not1  g2756(.din(new_new_n4183__), .dout(n9981));
  not1  g2757(.din(new_new_n4184__), .dout(n9984));
  not1  g2758(.din(new_new_n4185__), .dout(n9987));
  not1  g2759(.din(new_new_n4186__), .dout(n9990));
  not1  g2760(.din(new_new_n4187__), .dout(n9993));
  not1  g2761(.din(new_new_n4188__), .dout(n9996));
  buf1  g2762(.din(new_new_n4189__), .dout(n9999));
  buf1  g2763(.din(new_new_n4190__), .dout(n10002));
  not1  g2764(.din(new_new_n4191__), .dout(n10005));
  buf1  g2765(.din(new_new_n4192__), .dout(n10008));
  buf1  g2766(.din(new_new_n4193__), .dout(n10011));
  not1  g2767(.din(new_new_n4194__), .dout(n10014));
  not1  g2768(.din(new_new_n4195__), .dout(n10017));
  not1  g2769(.din(new_new_n4196__), .dout(n10020));
  not1  g2770(.din(new_new_n4197__), .dout(n10023));
  not1  g2771(.din(new_new_n4198__), .dout(n10026));
  not1  g2772(.din(new_new_n4199__), .dout(n10029));
  not1  g2773(.din(new_new_n4200__), .dout(n10032));
  buf1  g2774(.din(n9660), .dout(n10035));
  buf1  g2775(.din(n9663), .dout(n10038));
  buf1  g2776(.din(new_new_n4211__), .dout(n10041));
  buf1  g2777(.din(new_new_n4222__), .dout(n10044));
  buf1  g2778(.din(new_new_n4229__), .dout(n10047));
  buf1  g2779(.din(new_new_n5754__), .dout(n10050));
  buf1  g2780(.din(new_new_n4240__), .dout(n10053));
  buf1  g2781(.din(n9720), .dout(n10056));
  buf1  g2782(.din(n9759), .dout(n10059));
  buf1  g2783(.din(n9762), .dout(n10062));
  buf1  g2784(.din(new_new_n4243__), .dout(n10065));
  buf1  g2785(.din(new_new_n4246__), .dout(n10068));
  buf1  g2786(.din(new_new_n4249__), .dout(n10071));
  buf1  g2787(.din(new_new_n4252__), .dout(n10074));
  buf1  g2788(.din(n9855), .dout(n10077));
  buf1  g2789(.din(new_new_n4256__), .dout(n10080));
  buf1  g2790(.din(new_new_n4260__), .dout(n10083));
  buf1  g2791(.din(new_new_n5772__), .dout(n10086));
  buf1  g2792(.din(new_new_n5774__), .dout(n10089));
  buf1  g2793(.din(new_new_n5776__), .dout(n10092));
  buf1  g2794(.din(n9867), .dout(n10095));
  buf1  g2795(.din(new_new_n5778__), .dout(n10098));
  not1  g2796(.din(new_new_n5784__), .dout(n10101));
  buf1  g2797(.din(n10101), .dout(n10104));
  buf1  g2798(.din(new_new_n1940__), .dout(n10107));
  buf1  g2799(.din(new_new_n2104__), .dout(n10110));
  buf1  g2800(.din(new_new_n2108__), .dout(n10113));
  buf1  g2801(.din(new_new_n2134__), .dout(n10116));
  buf1  g2802(.din(new_new_n2138__), .dout(n10119));
  buf1  g2803(.din(new_new_n2166__), .dout(n10122));
  buf1  g2804(.din(new_new_n2170__), .dout(n10125));
  buf1  g2805(.din(new_new_n2198__), .dout(n10128));
  buf1  g2806(.din(new_new_n2202__), .dout(n10131));
  buf1  g2807(.din(new_new_n2406__), .dout(n10134));
  buf1  g2808(.din(new_new_n2410__), .dout(n10137));
  buf1  g2809(.din(new_new_n2416__), .dout(n10140));
  buf1  g2810(.din(new_new_n2418__), .dout(n10143));
  buf1  g2811(.din(new_new_n2448__), .dout(n10146));
  buf1  g2812(.din(new_new_n2450__), .dout(n10149));
  buf1  g2813(.din(new_new_n2460__), .dout(n10152));
  buf1  g2814(.din(new_new_n2464__), .dout(n10155));
  buf1  g2815(.din(new_new_n4262__), .dout(n10158));
  buf1  g2816(.din(new_new_n4264__), .dout(n10161));
  buf1  g2817(.din(new_new_n4266__), .dout(n10164));
  buf1  g2818(.din(new_new_n4268__), .dout(n10167));
  buf1  g2819(.din(new_new_n4270__), .dout(n10170));
  buf1  g2820(.din(new_new_n4271__), .dout(n10173));
  not1  g2821(.din(new_new_n5587__), .dout(n10176));
  buf1  g2822(.din(new_new_n4273__), .dout(n10179));
  buf1  g2823(.din(new_new_n4275__), .dout(n10182));
  buf1  g2824(.din(new_new_n4277__), .dout(n10185));
  buf1  g2825(.din(n9879), .dout(n10188));
  not1  g2826(.din(new_new_n5788__), .dout(n10191));
  buf1  g2827(.din(new_new_n4279__), .dout(n10194));
  buf1  g2828(.din(new_new_n4281__), .dout(n10197));
  buf1  g2829(.din(new_new_n2094__), .dout(n10200));
  buf1  g2830(.din(new_new_n2106__), .dout(n10203));
  buf1  g2831(.din(new_new_n2126__), .dout(n10206));
  buf1  g2832(.din(new_new_n2136__), .dout(n10209));
  buf1  g2833(.din(new_new_n2156__), .dout(n10212));
  buf1  g2834(.din(new_new_n2168__), .dout(n10215));
  buf1  g2835(.din(new_new_n2188__), .dout(n10218));
  buf1  g2836(.din(new_new_n2200__), .dout(n10221));
  buf1  g2837(.din(new_new_n2216__), .dout(n10224));
  buf1  g2838(.din(new_new_n2240__), .dout(n10227));
  buf1  g2839(.din(new_new_n2246__), .dout(n10230));
  buf1  g2840(.din(new_new_n2270__), .dout(n10233));
  buf1  g2841(.din(new_new_n2276__), .dout(n10236));
  buf1  g2842(.din(new_new_n2300__), .dout(n10239));
  buf1  g2843(.din(new_new_n2306__), .dout(n10242));
  buf1  g2844(.din(new_new_n2330__), .dout(n10245));
  buf1  g2845(.din(n9933), .dout(n10248));
  buf1  g2846(.din(n9936), .dout(n10251));
  buf1  g2847(.din(new_new_n4292__), .dout(n10254));
  buf1  g2848(.din(new_new_n4303__), .dout(n10257));
  buf1  g2849(.din(new_new_n4305__), .dout(n10260));
  not1  g2850(.din(new_new_n5790__), .dout(n10263));
  buf1  g2851(.din(n10263), .dout(n10266));
  buf1  g2852(.din(new_new_n1732__), .dout(n10269));
  buf1  g2853(.din(new_new_n1734__), .dout(n10272));
  buf1  g2854(.din(new_new_n1752__), .dout(n10275));
  buf1  g2855(.din(new_new_n1754__), .dout(n10278));
  buf1  g2856(.din(new_new_n1772__), .dout(n10281));
  buf1  g2857(.din(new_new_n1774__), .dout(n10284));
  buf1  g2858(.din(new_new_n1792__), .dout(n10287));
  buf1  g2859(.din(new_new_n1794__), .dout(n10290));
  buf1  g2860(.din(new_new_n1864__), .dout(n10293));
  buf1  g2861(.din(new_new_n1866__), .dout(n10296));
  buf1  g2862(.din(new_new_n2377__), .dout(new_new_n5047__));
  buf1  g2863(.din(new_new_n2343__), .dout(new_new_n5048__));
  buf1  g2864(.din(new_new_n5048__), .dout(new_new_n5049__));
  buf1  g2865(.din(new_new_n5048__), .dout(new_new_n5050__));
  buf1  g2866(.din(new_new_n3250__), .dout(new_new_n5051__));
  buf1  g2867(.din(new_new_n5051__), .dout(new_new_n5052__));
  buf1  g2868(.din(new_new_n2285__), .dout(new_new_n5053__));
  buf1  g2869(.din(new_new_n2125__), .dout(new_new_n5054__));
  buf1  g2870(.din(new_new_n2255__), .dout(new_new_n5055__));
  buf1  g2871(.din(new_new_n2155__), .dout(new_new_n5056__));
  buf1  g2872(.din(new_new_n2315__), .dout(new_new_n5057__));
  buf1  g2873(.din(new_new_n2187__), .dout(new_new_n5058__));
  buf1  g2874(.din(new_new_n2225__), .dout(new_new_n5059__));
  buf1  g2875(.din(new_new_n2093__), .dout(new_new_n5060__));
  buf1  g2876(.din(new_new_n3258__), .dout(new_new_n5061__));
  buf1  g2877(.din(new_new_n3255__), .dout(new_new_n5062__));
  buf1  g2878(.din(new_new_n2384__), .dout(new_new_n5063__));
  buf1  g2879(.din(new_new_n5063__), .dout(new_new_n5064__));
  buf1  g2880(.din(new_new_n2385__), .dout(new_new_n5065__));
  buf1  g2881(.din(new_new_n5065__), .dout(new_new_n5066__));
  buf1  g2882(.din(new_new_n3265__), .dout(new_new_n5067__));
  buf1  g2883(.din(new_new_n3262__), .dout(new_new_n5068__));
  buf1  g2884(.din(new_new_n5068__), .dout(new_new_n5069__));
  buf1  g2885(.din(new_new_n5068__), .dout(new_new_n5070__));
  buf1  g2886(.din(new_new_n2392__), .dout(new_new_n5071__));
  buf1  g2887(.din(new_new_n5071__), .dout(new_new_n5072__));
  buf1  g2888(.din(new_new_n5072__), .dout(new_new_n5073__));
  buf1  g2889(.din(new_new_n5071__), .dout(new_new_n5074__));
  buf1  g2890(.din(new_new_n2564__), .dout(new_new_n5075__));
  buf1  g2891(.din(new_new_n2393__), .dout(new_new_n5076__));
  buf1  g2892(.din(new_new_n5076__), .dout(new_new_n5077__));
  buf1  g2893(.din(new_new_n5077__), .dout(new_new_n5078__));
  buf1  g2894(.din(new_new_n5076__), .dout(new_new_n5079__));
  buf1  g2895(.din(new_new_n2562__), .dout(new_new_n5080__));
  buf1  g2896(.din(new_new_n2547__), .dout(new_new_n5081__));
  buf1  g2897(.din(new_new_n3283__), .dout(new_new_n5082__));
  buf1  g2898(.din(new_new_n2571__), .dout(new_new_n5083__));
  buf1  g2899(.din(new_new_n3287__), .dout(new_new_n5084__));
  buf1  g2900(.din(new_new_n1949__), .dout(new_new_n5085__));
  buf1  g2901(.din(new_new_n2925__), .dout(new_new_n5086__));
  buf1  g2902(.din(new_new_n2856__), .dout(new_new_n5087__));
  buf1  g2903(.din(new_new_n2924__), .dout(new_new_n5088__));
  buf1  g2904(.din(new_new_n2857__), .dout(new_new_n5089__));
  buf1  g2905(.din(new_new_n2568__), .dout(new_new_n5090__));
  buf1  g2906(.din(new_new_n5090__), .dout(new_new_n5091__));
  buf1  g2907(.din(new_new_n2079__), .dout(new_new_n5092__));
  buf1  g2908(.din(new_new_n2926__), .dout(new_new_n5093__));
  buf1  g2909(.din(new_new_n3434__), .dout(new_new_n5094__));
  buf1  g2910(.din(new_new_n3412__), .dout(new_new_n5095__));
  buf1  g2911(.din(new_new_n3310__), .dout(new_new_n5096__));
  buf1  g2912(.din(new_new_n3325__), .dout(new_new_n5097__));
  buf1  g2913(.din(new_new_n3295__), .dout(new_new_n5098__));
  buf1  g2914(.din(new_new_n3437__), .dout(new_new_n5099__));
  buf1  g2915(.din(new_new_n2673__), .dout(new_new_n5100__));
  buf1  g2916(.din(new_new_n2672__), .dout(new_new_n5101__));
  buf1  g2917(.din(new_new_n5101__), .dout(new_new_n5102__));
  buf1  g2918(.din(new_new_n5101__), .dout(new_new_n5103__));
  buf1  g2919(.din(new_new_n2966__), .dout(new_new_n5104__));
  buf1  g2920(.din(new_new_n2968__), .dout(new_new_n5105__));
  buf1  g2921(.din(new_new_n2813__), .dout(new_new_n5106__));
  buf1  g2922(.din(new_new_n2815__), .dout(new_new_n5107__));
  buf1  g2923(.din(new_new_n3084__), .dout(new_new_n5108__));
  buf1  g2924(.din(new_new_n5108__), .dout(new_new_n5109__));
  buf1  g2925(.din(new_new_n5109__), .dout(new_new_n5110__));
  buf1  g2926(.din(new_new_n5109__), .dout(new_new_n5111__));
  buf1  g2927(.din(new_new_n5108__), .dout(new_new_n5112__));
  buf1  g2928(.din(new_new_n5112__), .dout(new_new_n5113__));
  buf1  g2929(.din(new_new_n5112__), .dout(new_new_n5114__));
  buf1  g2930(.din(new_new_n3086__), .dout(new_new_n5115__));
  buf1  g2931(.din(new_new_n5115__), .dout(new_new_n5116__));
  buf1  g2932(.din(new_new_n5116__), .dout(new_new_n5117__));
  buf1  g2933(.din(new_new_n5116__), .dout(new_new_n5118__));
  buf1  g2934(.din(new_new_n5115__), .dout(new_new_n5119__));
  buf1  g2935(.din(new_new_n5119__), .dout(new_new_n5120__));
  buf1  g2936(.din(new_new_n5119__), .dout(new_new_n5121__));
  buf1  g2937(.din(new_new_n2885__), .dout(new_new_n5122__));
  buf1  g2938(.din(new_new_n5122__), .dout(new_new_n5123__));
  buf1  g2939(.din(new_new_n5123__), .dout(new_new_n5124__));
  buf1  g2940(.din(new_new_n5123__), .dout(new_new_n5125__));
  buf1  g2941(.din(new_new_n5122__), .dout(new_new_n5126__));
  buf1  g2942(.din(new_new_n5126__), .dout(new_new_n5127__));
  buf1  g2943(.din(new_new_n5126__), .dout(new_new_n5128__));
  buf1  g2944(.din(new_new_n2887__), .dout(new_new_n5129__));
  buf1  g2945(.din(new_new_n5129__), .dout(new_new_n5130__));
  buf1  g2946(.din(new_new_n5130__), .dout(new_new_n5131__));
  buf1  g2947(.din(new_new_n5130__), .dout(new_new_n5132__));
  buf1  g2948(.din(new_new_n5129__), .dout(new_new_n5133__));
  buf1  g2949(.din(new_new_n5133__), .dout(new_new_n5134__));
  buf1  g2950(.din(new_new_n5133__), .dout(new_new_n5135__));
  buf1  g2951(.din(new_new_n3210__), .dout(new_new_n5136__));
  buf1  g2952(.din(new_new_n5136__), .dout(new_new_n5137__));
  buf1  g2953(.din(new_new_n5137__), .dout(new_new_n5138__));
  buf1  g2954(.din(new_new_n5138__), .dout(new_new_n5139__));
  buf1  g2955(.din(new_new_n5138__), .dout(new_new_n5140__));
  buf1  g2956(.din(new_new_n5137__), .dout(new_new_n5141__));
  buf1  g2957(.din(new_new_n5136__), .dout(new_new_n5142__));
  buf1  g2958(.din(new_new_n5142__), .dout(new_new_n5143__));
  buf1  g2959(.din(new_new_n5142__), .dout(new_new_n5144__));
  buf1  g2960(.din(new_new_n3211__), .dout(new_new_n5145__));
  buf1  g2961(.din(new_new_n5145__), .dout(new_new_n5146__));
  buf1  g2962(.din(new_new_n5146__), .dout(new_new_n5147__));
  buf1  g2963(.din(new_new_n5146__), .dout(new_new_n5148__));
  buf1  g2964(.din(new_new_n5145__), .dout(new_new_n5149__));
  buf1  g2965(.din(new_new_n3212__), .dout(new_new_n5150__));
  buf1  g2966(.din(new_new_n5150__), .dout(new_new_n5151__));
  buf1  g2967(.din(new_new_n5151__), .dout(new_new_n5152__));
  buf1  g2968(.din(new_new_n5152__), .dout(new_new_n5153__));
  buf1  g2969(.din(new_new_n5152__), .dout(new_new_n5154__));
  buf1  g2970(.din(new_new_n5151__), .dout(new_new_n5155__));
  buf1  g2971(.din(new_new_n5150__), .dout(new_new_n5156__));
  buf1  g2972(.din(new_new_n5156__), .dout(new_new_n5157__));
  buf1  g2973(.din(new_new_n5156__), .dout(new_new_n5158__));
  buf1  g2974(.din(new_new_n3213__), .dout(new_new_n5159__));
  buf1  g2975(.din(new_new_n5159__), .dout(new_new_n5160__));
  buf1  g2976(.din(new_new_n5160__), .dout(new_new_n5161__));
  buf1  g2977(.din(new_new_n5160__), .dout(new_new_n5162__));
  buf1  g2978(.din(new_new_n5159__), .dout(new_new_n5163__));
  buf1  g2979(.din(new_new_n3001__), .dout(new_new_n5164__));
  buf1  g2980(.din(new_new_n5164__), .dout(new_new_n5165__));
  buf1  g2981(.din(new_new_n5165__), .dout(new_new_n5166__));
  buf1  g2982(.din(new_new_n5166__), .dout(new_new_n5167__));
  buf1  g2983(.din(new_new_n5166__), .dout(new_new_n5168__));
  buf1  g2984(.din(new_new_n5165__), .dout(new_new_n5169__));
  buf1  g2985(.din(new_new_n5164__), .dout(new_new_n5170__));
  buf1  g2986(.din(new_new_n5170__), .dout(new_new_n5171__));
  buf1  g2987(.din(new_new_n5170__), .dout(new_new_n5172__));
  buf1  g2988(.din(new_new_n3000__), .dout(new_new_n5173__));
  buf1  g2989(.din(new_new_n5173__), .dout(new_new_n5174__));
  buf1  g2990(.din(new_new_n5174__), .dout(new_new_n5175__));
  buf1  g2991(.din(new_new_n5174__), .dout(new_new_n5176__));
  buf1  g2992(.din(new_new_n5173__), .dout(new_new_n5177__));
  buf1  g2993(.din(new_new_n3003__), .dout(new_new_n5178__));
  buf1  g2994(.din(new_new_n5178__), .dout(new_new_n5179__));
  buf1  g2995(.din(new_new_n5179__), .dout(new_new_n5180__));
  buf1  g2996(.din(new_new_n5180__), .dout(new_new_n5181__));
  buf1  g2997(.din(new_new_n5180__), .dout(new_new_n5182__));
  buf1  g2998(.din(new_new_n5179__), .dout(new_new_n5183__));
  buf1  g2999(.din(new_new_n5178__), .dout(new_new_n5184__));
  buf1  g3000(.din(new_new_n5184__), .dout(new_new_n5185__));
  buf1  g3001(.din(new_new_n5184__), .dout(new_new_n5186__));
  buf1  g3002(.din(new_new_n3002__), .dout(new_new_n5187__));
  buf1  g3003(.din(new_new_n5187__), .dout(new_new_n5188__));
  buf1  g3004(.din(new_new_n5188__), .dout(new_new_n5189__));
  buf1  g3005(.din(new_new_n5188__), .dout(new_new_n5190__));
  buf1  g3006(.din(new_new_n5187__), .dout(new_new_n5191__));
  buf1  g3007(.din(new_new_n3220__), .dout(new_new_n5192__));
  buf1  g3008(.din(new_new_n5192__), .dout(new_new_n5193__));
  buf1  g3009(.din(new_new_n5193__), .dout(new_new_n5194__));
  buf1  g3010(.din(new_new_n5194__), .dout(new_new_n5195__));
  buf1  g3011(.din(new_new_n5194__), .dout(new_new_n5196__));
  buf1  g3012(.din(new_new_n5193__), .dout(new_new_n5197__));
  buf1  g3013(.din(new_new_n5197__), .dout(new_new_n5198__));
  buf1  g3014(.din(new_new_n5192__), .dout(new_new_n5199__));
  buf1  g3015(.din(new_new_n5199__), .dout(new_new_n5200__));
  buf1  g3016(.din(new_new_n5199__), .dout(new_new_n5201__));
  buf1  g3017(.din(new_new_n3145__), .dout(new_new_n5202__));
  buf1  g3018(.din(new_new_n3221__), .dout(new_new_n5203__));
  buf1  g3019(.din(new_new_n5203__), .dout(new_new_n5204__));
  buf1  g3020(.din(new_new_n5204__), .dout(new_new_n5205__));
  buf1  g3021(.din(new_new_n5205__), .dout(new_new_n5206__));
  buf1  g3022(.din(new_new_n5205__), .dout(new_new_n5207__));
  buf1  g3023(.din(new_new_n5204__), .dout(new_new_n5208__));
  buf1  g3024(.din(new_new_n5208__), .dout(new_new_n5209__));
  buf1  g3025(.din(new_new_n5203__), .dout(new_new_n5210__));
  buf1  g3026(.din(new_new_n5210__), .dout(new_new_n5211__));
  buf1  g3027(.din(new_new_n5210__), .dout(new_new_n5212__));
  buf1  g3028(.din(new_new_n3144__), .dout(new_new_n5213__));
  buf1  g3029(.din(new_new_n5213__), .dout(new_new_n5214__));
  buf1  g3030(.din(new_new_n5213__), .dout(new_new_n5215__));
  buf1  g3031(.din(new_new_n3137__), .dout(new_new_n5216__));
  buf1  g3032(.din(new_new_n3136__), .dout(new_new_n5217__));
  buf1  g3033(.din(new_new_n5217__), .dout(new_new_n5218__));
  buf1  g3034(.din(new_new_n5217__), .dout(new_new_n5219__));
  buf1  g3035(.din(new_new_n3222__), .dout(new_new_n5220__));
  buf1  g3036(.din(new_new_n5220__), .dout(new_new_n5221__));
  buf1  g3037(.din(new_new_n5221__), .dout(new_new_n5222__));
  buf1  g3038(.din(new_new_n5222__), .dout(new_new_n5223__));
  buf1  g3039(.din(new_new_n5222__), .dout(new_new_n5224__));
  buf1  g3040(.din(new_new_n5221__), .dout(new_new_n5225__));
  buf1  g3041(.din(new_new_n5225__), .dout(new_new_n5226__));
  buf1  g3042(.din(new_new_n5220__), .dout(new_new_n5227__));
  buf1  g3043(.din(new_new_n5227__), .dout(new_new_n5228__));
  buf1  g3044(.din(new_new_n5227__), .dout(new_new_n5229__));
  buf1  g3045(.din(new_new_n3223__), .dout(new_new_n5230__));
  buf1  g3046(.din(new_new_n5230__), .dout(new_new_n5231__));
  buf1  g3047(.din(new_new_n5231__), .dout(new_new_n5232__));
  buf1  g3048(.din(new_new_n5232__), .dout(new_new_n5233__));
  buf1  g3049(.din(new_new_n5232__), .dout(new_new_n5234__));
  buf1  g3050(.din(new_new_n5231__), .dout(new_new_n5235__));
  buf1  g3051(.din(new_new_n5235__), .dout(new_new_n5236__));
  buf1  g3052(.din(new_new_n5230__), .dout(new_new_n5237__));
  buf1  g3053(.din(new_new_n5237__), .dout(new_new_n5238__));
  buf1  g3054(.din(new_new_n5237__), .dout(new_new_n5239__));
  buf1  g3055(.din(new_new_n3567__), .dout(new_new_n5240__));
  buf1  g3056(.din(new_new_n5240__), .dout(new_new_n5241__));
  buf1  g3057(.din(new_new_n5240__), .dout(new_new_n5242__));
  buf1  g3058(.din(new_new_n3570__), .dout(new_new_n5243__));
  buf1  g3059(.din(new_new_n5243__), .dout(new_new_n5244__));
  buf1  g3060(.din(new_new_n3574__), .dout(new_new_n5245__));
  buf1  g3061(.din(new_new_n3585__), .dout(new_new_n5246__));
  buf1  g3062(.din(new_new_n5246__), .dout(new_new_n5247__));
  buf1  g3063(.din(new_new_n5247__), .dout(new_new_n5248__));
  buf1  g3064(.din(new_new_n5246__), .dout(new_new_n5249__));
  buf1  g3065(.din(new_new_n3584__), .dout(new_new_n5250__));
  buf1  g3066(.din(new_new_n5250__), .dout(new_new_n5251__));
  buf1  g3067(.din(new_new_n5251__), .dout(new_new_n5252__));
  buf1  g3068(.din(new_new_n5250__), .dout(new_new_n5253__));
  buf1  g3069(.din(new_new_n3591__), .dout(new_new_n5254__));
  buf1  g3070(.din(new_new_n5254__), .dout(new_new_n5255__));
  buf1  g3071(.din(new_new_n5254__), .dout(new_new_n5256__));
  buf1  g3072(.din(new_new_n3590__), .dout(new_new_n5257__));
  buf1  g3073(.din(new_new_n5257__), .dout(new_new_n5258__));
  buf1  g3074(.din(new_new_n5257__), .dout(new_new_n5259__));
  buf1  g3075(.din(new_new_n3599__), .dout(new_new_n5260__));
  buf1  g3076(.din(new_new_n5260__), .dout(new_new_n5261__));
  buf1  g3077(.din(new_new_n3598__), .dout(new_new_n5262__));
  buf1  g3078(.din(new_new_n5262__), .dout(new_new_n5263__));
  buf1  g3079(.din(new_new_n2782__), .dout(new_new_n5264__));
  buf1  g3080(.din(new_new_n2783__), .dout(new_new_n5265__));
  buf1  g3081(.din(new_new_n3609__), .dout(new_new_n5266__));
  buf1  g3082(.din(new_new_n3608__), .dout(new_new_n5267__));
  buf1  g3083(.din(new_new_n2690__), .dout(new_new_n5268__));
  buf1  g3084(.din(new_new_n5268__), .dout(new_new_n5269__));
  buf1  g3085(.din(new_new_n2691__), .dout(new_new_n5270__));
  buf1  g3086(.din(new_new_n5270__), .dout(new_new_n5271__));
  buf1  g3087(.din(new_new_n3091__), .dout(new_new_n5272__));
  buf1  g3088(.din(new_new_n3090__), .dout(new_new_n5273__));
  buf1  g3089(.din(new_new_n3581__), .dout(new_new_n5274__));
  buf1  g3090(.din(new_new_n3665__), .dout(new_new_n5275__));
  buf1  g3091(.din(new_new_n5275__), .dout(new_new_n5276__));
  buf1  g3092(.din(new_new_n5275__), .dout(new_new_n5277__));
  buf1  g3093(.din(new_new_n3668__), .dout(new_new_n5278__));
  buf1  g3094(.din(new_new_n5278__), .dout(new_new_n5279__));
  buf1  g3095(.din(new_new_n3672__), .dout(new_new_n5280__));
  buf1  g3096(.din(new_new_n3683__), .dout(new_new_n5281__));
  buf1  g3097(.din(new_new_n5281__), .dout(new_new_n5282__));
  buf1  g3098(.din(new_new_n5282__), .dout(new_new_n5283__));
  buf1  g3099(.din(new_new_n5281__), .dout(new_new_n5284__));
  buf1  g3100(.din(new_new_n3682__), .dout(new_new_n5285__));
  buf1  g3101(.din(new_new_n5285__), .dout(new_new_n5286__));
  buf1  g3102(.din(new_new_n5286__), .dout(new_new_n5287__));
  buf1  g3103(.din(new_new_n5285__), .dout(new_new_n5288__));
  buf1  g3104(.din(new_new_n3689__), .dout(new_new_n5289__));
  buf1  g3105(.din(new_new_n5289__), .dout(new_new_n5290__));
  buf1  g3106(.din(new_new_n5289__), .dout(new_new_n5291__));
  buf1  g3107(.din(new_new_n3688__), .dout(new_new_n5292__));
  buf1  g3108(.din(new_new_n5292__), .dout(new_new_n5293__));
  buf1  g3109(.din(new_new_n5292__), .dout(new_new_n5294__));
  buf1  g3110(.din(new_new_n3697__), .dout(new_new_n5295__));
  buf1  g3111(.din(new_new_n5295__), .dout(new_new_n5296__));
  buf1  g3112(.din(new_new_n3696__), .dout(new_new_n5297__));
  buf1  g3113(.din(new_new_n5297__), .dout(new_new_n5298__));
  buf1  g3114(.din(new_new_n3707__), .dout(new_new_n5299__));
  buf1  g3115(.din(new_new_n3706__), .dout(new_new_n5300__));
  buf1  g3116(.din(new_new_n3095__), .dout(new_new_n5301__));
  buf1  g3117(.din(new_new_n3094__), .dout(new_new_n5302__));
  buf1  g3118(.din(new_new_n3679__), .dout(new_new_n5303__));
  buf1  g3119(.din(new_new_n2988__), .dout(new_new_n5304__));
  buf1  g3120(.din(new_new_n2981__), .dout(new_new_n5305__));
  buf1  g3121(.din(new_new_n2989__), .dout(new_new_n5306__));
  buf1  g3122(.din(new_new_n2980__), .dout(new_new_n5307__));
  buf1  g3123(.din(new_new_n2990__), .dout(new_new_n5308__));
  buf1  g3124(.din(new_new_n2987__), .dout(new_new_n5309__));
  buf1  g3125(.din(new_new_n2991__), .dout(new_new_n5310__));
  buf1  g3126(.din(new_new_n2986__), .dout(new_new_n5311__));
  buf1  g3127(.din(new_new_n2526__), .dout(new_new_n5312__));
  buf1  g3128(.din(new_new_n2521__), .dout(new_new_n5313__));
  buf1  g3129(.din(new_new_n2527__), .dout(new_new_n5314__));
  buf1  g3130(.din(new_new_n2520__), .dout(new_new_n5315__));
  buf1  g3131(.din(new_new_n2679__), .dout(new_new_n5316__));
  buf1  g3132(.din(new_new_n2586__), .dout(new_new_n5317__));
  buf1  g3133(.din(new_new_n2678__), .dout(new_new_n5318__));
  buf1  g3134(.din(new_new_n2587__), .dout(new_new_n5319__));
  buf1  g3135(.din(new_new_n3074__), .dout(new_new_n5320__));
  buf1  g3136(.din(new_new_n5320__), .dout(new_new_n5321__));
  buf1  g3137(.din(new_new_n5320__), .dout(new_new_n5322__));
  buf1  g3138(.din(new_new_n2577__), .dout(new_new_n5323__));
  buf1  g3139(.din(new_new_n3075__), .dout(new_new_n5324__));
  buf1  g3140(.din(new_new_n2576__), .dout(new_new_n5325__));
  buf1  g3141(.din(new_new_n5325__), .dout(new_new_n5326__));
  buf1  g3142(.din(new_new_n5325__), .dout(new_new_n5327__));
  buf1  g3143(.din(new_new_n3077__), .dout(new_new_n5328__));
  buf1  g3144(.din(new_new_n3073__), .dout(new_new_n5329__));
  buf1  g3145(.din(new_new_n3076__), .dout(new_new_n5330__));
  buf1  g3146(.din(new_new_n5330__), .dout(new_new_n5331__));
  buf1  g3147(.din(new_new_n3072__), .dout(new_new_n5332__));
  buf1  g3148(.din(new_new_n5332__), .dout(new_new_n5333__));
  buf1  g3149(.din(new_new_n3773__), .dout(new_new_n5334__));
  buf1  g3150(.din(new_new_n5334__), .dout(new_new_n5335__));
  buf1  g3151(.din(new_new_n3779__), .dout(new_new_n5336__));
  buf1  g3152(.din(new_new_n5336__), .dout(new_new_n5337__));
  buf1  g3153(.din(new_new_n2972__), .dout(new_new_n5338__));
  buf1  g3154(.din(new_new_n2971__), .dout(new_new_n5339__));
  buf1  g3155(.din(new_new_n2973__), .dout(new_new_n5340__));
  buf1  g3156(.din(new_new_n2970__), .dout(new_new_n5341__));
  buf1  g3157(.din(new_new_n2976__), .dout(new_new_n5342__));
  buf1  g3158(.din(new_new_n2975__), .dout(new_new_n5343__));
  buf1  g3159(.din(new_new_n2977__), .dout(new_new_n5344__));
  buf1  g3160(.din(new_new_n2974__), .dout(new_new_n5345__));
  buf1  g3161(.din(new_new_n3824__), .dout(new_new_n5346__));
  buf1  g3162(.din(new_new_n3817__), .dout(new_new_n5347__));
  buf1  g3163(.din(new_new_n3829__), .dout(new_new_n5348__));
  buf1  g3164(.din(new_new_n3818__), .dout(new_new_n5349__));
  buf1  g3165(.din(new_new_n3830__), .dout(new_new_n5350__));
  buf1  g3166(.din(new_new_n3823__), .dout(new_new_n5351__));
  buf1  g3167(.din(new_new_n3080__), .dout(new_new_n5352__));
  buf1  g3168(.din(new_new_n2982__), .dout(new_new_n5353__));
  buf1  g3169(.din(new_new_n3081__), .dout(new_new_n5354__));
  buf1  g3170(.din(new_new_n2983__), .dout(new_new_n5355__));
  buf1  g3171(.din(new_new_n2985__), .dout(new_new_n5356__));
  buf1  g3172(.din(new_new_n2978__), .dout(new_new_n5357__));
  buf1  g3173(.din(new_new_n2984__), .dout(new_new_n5358__));
  buf1  g3174(.din(new_new_n2979__), .dout(new_new_n5359__));
  buf1  g3175(.din(new_new_n3852__), .dout(new_new_n5360__));
  buf1  g3176(.din(new_new_n3847__), .dout(new_new_n5361__));
  buf1  g3177(.din(new_new_n3859__), .dout(new_new_n5362__));
  buf1  g3178(.din(new_new_n3846__), .dout(new_new_n5363__));
  buf1  g3179(.din(new_new_n3858__), .dout(new_new_n5364__));
  buf1  g3180(.din(new_new_n3853__), .dout(new_new_n5365__));
  buf1  g3181(.din(new_new_n3110__), .dout(new_new_n5366__));
  buf1  g3182(.din(new_new_n3109__), .dout(new_new_n5367__));
  buf1  g3183(.din(new_new_n3111__), .dout(new_new_n5368__));
  buf1  g3184(.din(new_new_n3108__), .dout(new_new_n5369__));
  buf1  g3185(.din(new_new_n2998__), .dout(new_new_n5370__));
  buf1  g3186(.din(new_new_n2996__), .dout(new_new_n5371__));
  buf1  g3187(.din(new_new_n2999__), .dout(new_new_n5372__));
  buf1  g3188(.din(new_new_n2997__), .dout(new_new_n5373__));
  buf1  g3189(.din(new_new_n3882__), .dout(new_new_n5374__));
  buf1  g3190(.din(new_new_n3875__), .dout(new_new_n5375__));
  buf1  g3191(.din(new_new_n3887__), .dout(new_new_n5376__));
  buf1  g3192(.din(new_new_n3876__), .dout(new_new_n5377__));
  buf1  g3193(.din(new_new_n3888__), .dout(new_new_n5378__));
  buf1  g3194(.din(new_new_n3881__), .dout(new_new_n5379__));
  buf1  g3195(.din(new_new_n2457__), .dout(new_new_n5380__));
  buf1  g3196(.din(new_new_n2415__), .dout(new_new_n5381__));
  buf1  g3197(.din(new_new_n2422__), .dout(new_new_n5382__));
  buf1  g3198(.din(new_new_n5382__), .dout(new_new_n5383__));
  buf1  g3199(.din(new_new_n5382__), .dout(new_new_n5384__));
  buf1  g3200(.din(new_new_n3117__), .dout(new_new_n5385__));
  buf1  g3201(.din(new_new_n5385__), .dout(new_new_n5386__));
  buf1  g3202(.din(new_new_n5386__), .dout(new_new_n5387__));
  buf1  g3203(.din(new_new_n5387__), .dout(new_new_n5388__));
  buf1  g3204(.din(new_new_n5387__), .dout(new_new_n5389__));
  buf1  g3205(.din(new_new_n5386__), .dout(new_new_n5390__));
  buf1  g3206(.din(new_new_n5390__), .dout(new_new_n5391__));
  buf1  g3207(.din(new_new_n5390__), .dout(new_new_n5392__));
  buf1  g3208(.din(new_new_n5385__), .dout(new_new_n5393__));
  buf1  g3209(.din(new_new_n5393__), .dout(new_new_n5394__));
  buf1  g3210(.din(new_new_n5394__), .dout(new_new_n5395__));
  buf1  g3211(.din(new_new_n5394__), .dout(new_new_n5396__));
  buf1  g3212(.din(new_new_n5393__), .dout(new_new_n5397__));
  buf1  g3213(.din(new_new_n5397__), .dout(new_new_n5398__));
  buf1  g3214(.din(new_new_n5397__), .dout(new_new_n5399__));
  buf1  g3215(.din(new_new_n2426__), .dout(new_new_n5400__));
  buf1  g3216(.din(new_new_n5400__), .dout(new_new_n5401__));
  buf1  g3217(.din(new_new_n5400__), .dout(new_new_n5402__));
  buf1  g3218(.din(new_new_n3142__), .dout(new_new_n5403__));
  buf1  g3219(.din(new_new_n5403__), .dout(new_new_n5404__));
  buf1  g3220(.din(new_new_n5404__), .dout(new_new_n5405__));
  buf1  g3221(.din(new_new_n5404__), .dout(new_new_n5406__));
  buf1  g3222(.din(new_new_n5403__), .dout(new_new_n5407__));
  buf1  g3223(.din(new_new_n3918__), .dout(new_new_n5408__));
  buf1  g3224(.din(new_new_n5408__), .dout(new_new_n5409__));
  buf1  g3225(.din(new_new_n5408__), .dout(new_new_n5410__));
  buf1  g3226(.din(new_new_n2435__), .dout(new_new_n5411__));
  buf1  g3227(.din(new_new_n3917__), .dout(new_new_n5412__));
  buf1  g3228(.din(new_new_n5412__), .dout(new_new_n5413__));
  buf1  g3229(.din(new_new_n5413__), .dout(new_new_n5414__));
  buf1  g3230(.din(new_new_n5413__), .dout(new_new_n5415__));
  buf1  g3231(.din(new_new_n5412__), .dout(new_new_n5416__));
  buf1  g3232(.din(new_new_n5416__), .dout(new_new_n5417__));
  buf1  g3233(.din(new_new_n5416__), .dout(new_new_n5418__));
  buf1  g3234(.din(new_new_n2439__), .dout(new_new_n5419__));
  buf1  g3235(.din(new_new_n3146__), .dout(new_new_n5420__));
  buf1  g3236(.din(new_new_n5420__), .dout(new_new_n5421__));
  buf1  g3237(.din(new_new_n5420__), .dout(new_new_n5422__));
  buf1  g3238(.din(new_new_n3138__), .dout(new_new_n5423__));
  buf1  g3239(.din(new_new_n5423__), .dout(new_new_n5424__));
  buf1  g3240(.din(new_new_n5423__), .dout(new_new_n5425__));
  buf1  g3241(.din(new_new_n3148__), .dout(new_new_n5426__));
  buf1  g3242(.din(new_new_n5426__), .dout(new_new_n5427__));
  buf1  g3243(.din(new_new_n5426__), .dout(new_new_n5428__));
  buf1  g3244(.din(new_new_n3140__), .dout(new_new_n5429__));
  buf1  g3245(.din(new_new_n5429__), .dout(new_new_n5430__));
  buf1  g3246(.din(new_new_n5429__), .dout(new_new_n5431__));
  buf1  g3247(.din(new_new_n3451__), .dout(new_new_n5432__));
  buf1  g3248(.din(new_new_n5432__), .dout(new_new_n5433__));
  buf1  g3249(.din(new_new_n5433__), .dout(new_new_n5434__));
  buf1  g3250(.din(new_new_n5432__), .dout(new_new_n5435__));
  buf1  g3251(.din(new_new_n3171__), .dout(new_new_n5436__));
  buf1  g3252(.din(new_new_n5436__), .dout(new_new_n5437__));
  buf1  g3253(.din(new_new_n5436__), .dout(new_new_n5438__));
  buf1  g3254(.din(new_new_n3448__), .dout(new_new_n5439__));
  buf1  g3255(.din(new_new_n5439__), .dout(new_new_n5440__));
  buf1  g3256(.din(new_new_n5440__), .dout(new_new_n5441__));
  buf1  g3257(.din(new_new_n5439__), .dout(new_new_n5442__));
  buf1  g3258(.din(new_new_n3173__), .dout(new_new_n5443__));
  buf1  g3259(.din(new_new_n5443__), .dout(new_new_n5444__));
  buf1  g3260(.din(new_new_n5443__), .dout(new_new_n5445__));
  buf1  g3261(.din(new_new_n3476__), .dout(new_new_n5446__));
  buf1  g3262(.din(new_new_n5446__), .dout(new_new_n5447__));
  buf1  g3263(.din(new_new_n2965__), .dout(new_new_n5448__));
  buf1  g3264(.din(new_new_n3487__), .dout(new_new_n5449__));
  buf1  g3265(.din(new_new_n5449__), .dout(new_new_n5450__));
  buf1  g3266(.din(new_new_n3454__), .dout(new_new_n5451__));
  buf1  g3267(.din(new_new_n5451__), .dout(new_new_n5452__));
  buf1  g3268(.din(new_new_n2964__), .dout(new_new_n5453__));
  buf1  g3269(.din(new_new_n3216__), .dout(new_new_n5454__));
  buf1  g3270(.din(new_new_n5454__), .dout(new_new_n5455__));
  buf1  g3271(.din(new_new_n5455__), .dout(new_new_n5456__));
  buf1  g3272(.din(new_new_n5455__), .dout(new_new_n5457__));
  buf1  g3273(.din(new_new_n5454__), .dout(new_new_n5458__));
  buf1  g3274(.din(new_new_n5458__), .dout(new_new_n5459__));
  buf1  g3275(.din(new_new_n5458__), .dout(new_new_n5460__));
  buf1  g3276(.din(new_new_n3170__), .dout(new_new_n5461__));
  buf1  g3277(.din(new_new_n3214__), .dout(new_new_n5462__));
  buf1  g3278(.din(new_new_n5462__), .dout(new_new_n5463__));
  buf1  g3279(.din(new_new_n5463__), .dout(new_new_n5464__));
  buf1  g3280(.din(new_new_n5463__), .dout(new_new_n5465__));
  buf1  g3281(.din(new_new_n5462__), .dout(new_new_n5466__));
  buf1  g3282(.din(new_new_n5466__), .dout(new_new_n5467__));
  buf1  g3283(.din(new_new_n3172__), .dout(new_new_n5468__));
  buf1  g3284(.din(new_new_n2431__), .dout(new_new_n5469__));
  buf1  g3285(.din(new_new_n3465__), .dout(new_new_n5470__));
  buf1  g3286(.din(new_new_n5470__), .dout(new_new_n5471__));
  buf1  g3287(.din(new_new_n5470__), .dout(new_new_n5472__));
  buf1  g3288(.din(new_new_n3240__), .dout(new_new_n5473__));
  buf1  g3289(.din(new_new_n5473__), .dout(new_new_n5474__));
  buf1  g3290(.din(new_new_n5474__), .dout(new_new_n5475__));
  buf1  g3291(.din(new_new_n5475__), .dout(new_new_n5476__));
  buf1  g3292(.din(new_new_n5475__), .dout(new_new_n5477__));
  buf1  g3293(.din(new_new_n5474__), .dout(new_new_n5478__));
  buf1  g3294(.din(new_new_n5473__), .dout(new_new_n5479__));
  buf1  g3295(.din(new_new_n5479__), .dout(new_new_n5480__));
  buf1  g3296(.din(new_new_n5479__), .dout(new_new_n5481__));
  buf1  g3297(.din(new_new_n3242__), .dout(new_new_n5482__));
  buf1  g3298(.din(new_new_n5482__), .dout(new_new_n5483__));
  buf1  g3299(.din(new_new_n5483__), .dout(new_new_n5484__));
  buf1  g3300(.din(new_new_n5484__), .dout(new_new_n5485__));
  buf1  g3301(.din(new_new_n5484__), .dout(new_new_n5486__));
  buf1  g3302(.din(new_new_n5483__), .dout(new_new_n5487__));
  buf1  g3303(.din(new_new_n5482__), .dout(new_new_n5488__));
  buf1  g3304(.din(new_new_n5488__), .dout(new_new_n5489__));
  buf1  g3305(.din(new_new_n5488__), .dout(new_new_n5490__));
  buf1  g3306(.din(new_new_n3241__), .dout(new_new_n5491__));
  buf1  g3307(.din(new_new_n5491__), .dout(new_new_n5492__));
  buf1  g3308(.din(new_new_n5492__), .dout(new_new_n5493__));
  buf1  g3309(.din(new_new_n5492__), .dout(new_new_n5494__));
  buf1  g3310(.din(new_new_n5491__), .dout(new_new_n5495__));
  buf1  g3311(.din(new_new_n3243__), .dout(new_new_n5496__));
  buf1  g3312(.din(new_new_n5496__), .dout(new_new_n5497__));
  buf1  g3313(.din(new_new_n5497__), .dout(new_new_n5498__));
  buf1  g3314(.din(new_new_n5497__), .dout(new_new_n5499__));
  buf1  g3315(.din(new_new_n5496__), .dout(new_new_n5500__));
  buf1  g3316(.din(new_new_n2615__), .dout(new_new_n5501__));
  buf1  g3317(.din(new_new_n2590__), .dout(new_new_n5502__));
  buf1  g3318(.din(new_new_n2614__), .dout(new_new_n5503__));
  buf1  g3319(.din(new_new_n2591__), .dout(new_new_n5504__));
  buf1  g3320(.din(new_new_n2588__), .dout(new_new_n5505__));
  buf1  g3321(.din(new_new_n2532__), .dout(new_new_n5506__));
  buf1  g3322(.din(new_new_n2589__), .dout(new_new_n5507__));
  buf1  g3323(.din(new_new_n2533__), .dout(new_new_n5508__));
  buf1  g3324(.din(new_new_n4047__), .dout(new_new_n5509__));
  buf1  g3325(.din(new_new_n4041__), .dout(new_new_n5510__));
  buf1  g3326(.din(new_new_n4051__), .dout(new_new_n5511__));
  buf1  g3327(.din(new_new_n5511__), .dout(new_new_n5512__));
  buf1  g3328(.din(new_new_n5511__), .dout(new_new_n5513__));
  buf1  g3329(.din(new_new_n4048__), .dout(new_new_n5514__));
  buf1  g3330(.din(new_new_n2624__), .dout(new_new_n5515__));
  buf1  g3331(.din(new_new_n5515__), .dout(new_new_n5516__));
  buf1  g3332(.din(new_new_n2597__), .dout(new_new_n5517__));
  buf1  g3333(.din(new_new_n2625__), .dout(new_new_n5518__));
  buf1  g3334(.din(new_new_n2596__), .dout(new_new_n5519__));
  buf1  g3335(.din(new_new_n5519__), .dout(new_new_n5520__));
  buf1  g3336(.din(new_new_n2594__), .dout(new_new_n5521__));
  buf1  g3337(.din(new_new_n2538__), .dout(new_new_n5522__));
  buf1  g3338(.din(new_new_n2595__), .dout(new_new_n5523__));
  buf1  g3339(.din(new_new_n2539__), .dout(new_new_n5524__));
  buf1  g3340(.din(new_new_n2600__), .dout(new_new_n5525__));
  buf1  g3341(.din(new_new_n2598__), .dout(new_new_n5526__));
  buf1  g3342(.din(new_new_n4066__), .dout(new_new_n5527__));
  buf1  g3343(.din(new_new_n4060__), .dout(new_new_n5528__));
  buf1  g3344(.din(new_new_n4070__), .dout(new_new_n5529__));
  buf1  g3345(.din(new_new_n5529__), .dout(new_new_n5530__));
  buf1  g3346(.din(new_new_n5529__), .dout(new_new_n5531__));
  buf1  g3347(.din(new_new_n4067__), .dout(new_new_n5532__));
  buf1  g3348(.din(new_new_n4042__), .dout(new_new_n5533__));
  buf1  g3349(.din(new_new_n4061__), .dout(new_new_n5534__));
  buf1  g3350(.din(new_new_n2958__), .dout(new_new_n5535__));
  buf1  g3351(.din(new_new_n2957__), .dout(new_new_n5536__));
  buf1  g3352(.din(new_new_n2959__), .dout(new_new_n5537__));
  buf1  g3353(.din(new_new_n2956__), .dout(new_new_n5538__));
  buf1  g3354(.din(new_new_n4083__), .dout(new_new_n5539__));
  buf1  g3355(.din(new_new_n3445__), .dout(new_new_n5540__));
  buf1  g3356(.din(new_new_n5540__), .dout(new_new_n5541__));
  buf1  g3357(.din(new_new_n5540__), .dout(new_new_n5542__));
  buf1  g3358(.din(new_new_n4087__), .dout(new_new_n5543__));
  buf1  g3359(.din(new_new_n5543__), .dout(new_new_n5544__));
  buf1  g3360(.din(new_new_n5543__), .dout(new_new_n5545__));
  buf1  g3361(.din(new_new_n4084__), .dout(new_new_n5546__));
  buf1  g3362(.din(new_new_n3444__), .dout(new_new_n5547__));
  buf1  g3363(.din(new_new_n1970__), .dout(new_new_n5548__));
  buf1  g3364(.din(new_new_n5548__), .dout(new_new_n5549__));
  buf1  g3365(.din(new_new_n5549__), .dout(new_new_n5550__));
  buf1  g3366(.din(new_new_n5550__), .dout(new_new_n5551__));
  buf1  g3367(.din(new_new_n5549__), .dout(new_new_n5552__));
  buf1  g3368(.din(new_new_n5548__), .dout(new_new_n5553__));
  buf1  g3369(.din(new_new_n5553__), .dout(new_new_n5554__));
  buf1  g3370(.din(new_new_n5553__), .dout(new_new_n5555__));
  buf1  g3371(.din(new_new_n1971__), .dout(new_new_n5556__));
  buf1  g3372(.din(new_new_n5556__), .dout(new_new_n5557__));
  buf1  g3373(.din(new_new_n5557__), .dout(new_new_n5558__));
  buf1  g3374(.din(new_new_n5558__), .dout(new_new_n5559__));
  buf1  g3375(.din(new_new_n5557__), .dout(new_new_n5560__));
  buf1  g3376(.din(new_new_n5556__), .dout(new_new_n5561__));
  buf1  g3377(.din(new_new_n5561__), .dout(new_new_n5562__));
  buf1  g3378(.din(new_new_n5561__), .dout(new_new_n5563__));
  buf1  g3379(.din(new_new_n2670__), .dout(new_new_n5564__));
  buf1  g3380(.din(new_new_n2798__), .dout(new_new_n5565__));
  buf1  g3381(.din(new_new_n5565__), .dout(new_new_n5566__));
  buf1  g3382(.din(new_new_n2582__), .dout(new_new_n5567__));
  buf1  g3383(.din(new_new_n2580__), .dout(new_new_n5568__));
  buf1  g3384(.din(new_new_n2038__), .dout(new_new_n5569__));
  buf1  g3385(.din(new_new_n5569__), .dout(new_new_n5570__));
  buf1  g3386(.din(new_new_n5570__), .dout(new_new_n5571__));
  buf1  g3387(.din(new_new_n5571__), .dout(new_new_n5572__));
  buf1  g3388(.din(new_new_n5570__), .dout(new_new_n5573__));
  buf1  g3389(.din(new_new_n5569__), .dout(new_new_n5574__));
  buf1  g3390(.din(new_new_n5574__), .dout(new_new_n5575__));
  buf1  g3391(.din(new_new_n5574__), .dout(new_new_n5576__));
  buf1  g3392(.din(new_new_n2039__), .dout(new_new_n5577__));
  buf1  g3393(.din(new_new_n5577__), .dout(new_new_n5578__));
  buf1  g3394(.din(new_new_n5578__), .dout(new_new_n5579__));
  buf1  g3395(.din(new_new_n5578__), .dout(new_new_n5580__));
  buf1  g3396(.din(new_new_n5577__), .dout(new_new_n5581__));
  buf1  g3397(.din(new_new_n5581__), .dout(new_new_n5582__));
  buf1  g3398(.din(new_new_n2578__), .dout(new_new_n5583__));
  buf1  g3399(.din(new_new_n3761__), .dout(new_new_n5584__));
  buf1  g3400(.din(new_new_n3663__), .dout(new_new_n5585__));
  buf1  g3401(.din(new_new_n4036__), .dout(new_new_n5586__));
  buf1  g3402(.din(new_new_n4152__), .dout(new_new_n5587__));
  buf1  g3403(.din(new_new_n4025__), .dout(new_new_n5588__));
  buf1  g3404(.din(new_new_n5588__), .dout(new_new_n5589__));
  buf1  g3405(.din(new_new_n3143__), .dout(new_new_n5590__));
  buf1  g3406(.din(new_new_n3135__), .dout(new_new_n5591__));
  buf1  g3407(.din(new_new_n3134__), .dout(new_new_n5592__));
  buf1  g3408(.din(new_new_n5592__), .dout(new_new_n5593__));
  buf1  g3409(.din(new_new_n5592__), .dout(new_new_n5594__));
  buf1  g3410(.din(new_new_n4159__), .dout(new_new_n5595__));
  buf1  g3411(.din(new_new_n3553__), .dout(new_new_n5596__));
  buf1  g3412(.din(new_new_n5596__), .dout(new_new_n5597__));
  buf1  g3413(.din(new_new_n5597__), .dout(new_new_n5598__));
  buf1  g3414(.din(new_new_n5597__), .dout(new_new_n5599__));
  buf1  g3415(.din(new_new_n5596__), .dout(new_new_n5600__));
  buf1  g3416(.din(new_new_n5600__), .dout(new_new_n5601__));
  buf1  g3417(.din(new_new_n4166__), .dout(new_new_n5602__));
  buf1  g3418(.din(new_new_n3902__), .dout(new_new_n5603__));
  buf1  g3419(.din(new_new_n5603__), .dout(new_new_n5604__));
  buf1  g3420(.din(new_new_n3530__), .dout(new_new_n5605__));
  buf1  g3421(.din(new_new_n5605__), .dout(new_new_n5606__));
  buf1  g3422(.din(new_new_n5605__), .dout(new_new_n5607__));
  buf1  g3423(.din(new_new_n3947__), .dout(new_new_n5608__));
  buf1  g3424(.din(new_new_n5608__), .dout(new_new_n5609__));
  buf1  g3425(.din(new_new_n3904__), .dout(new_new_n5610__));
  buf1  g3426(.din(new_new_n5610__), .dout(new_new_n5611__));
  buf1  g3427(.din(new_new_n3949__), .dout(new_new_n5612__));
  buf1  g3428(.din(new_new_n5612__), .dout(new_new_n5613__));
  buf1  g3429(.din(new_new_n3906__), .dout(new_new_n5614__));
  buf1  g3430(.din(new_new_n5614__), .dout(new_new_n5615__));
  buf1  g3431(.din(new_new_n3909__), .dout(new_new_n5616__));
  buf1  g3432(.din(new_new_n5616__), .dout(new_new_n5617__));
  buf1  g3433(.din(new_new_n3951__), .dout(new_new_n5618__));
  buf1  g3434(.din(new_new_n5618__), .dout(new_new_n5619__));
  buf1  g3435(.din(new_new_n3911__), .dout(new_new_n5620__));
  buf1  g3436(.din(new_new_n5620__), .dout(new_new_n5621__));
  buf1  g3437(.din(new_new_n3953__), .dout(new_new_n5622__));
  buf1  g3438(.din(new_new_n5622__), .dout(new_new_n5623__));
  buf1  g3439(.din(new_new_n3913__), .dout(new_new_n5624__));
  buf1  g3440(.din(new_new_n5624__), .dout(new_new_n5625__));
  buf1  g3441(.din(new_new_n3959__), .dout(new_new_n5626__));
  buf1  g3442(.din(new_new_n5626__), .dout(new_new_n5627__));
  buf1  g3443(.din(new_new_n5627__), .dout(new_new_n5628__));
  buf1  g3444(.din(new_new_n5627__), .dout(new_new_n5629__));
  buf1  g3445(.din(new_new_n5626__), .dout(new_new_n5630__));
  buf1  g3446(.din(new_new_n3919__), .dout(new_new_n5631__));
  buf1  g3447(.din(new_new_n5631__), .dout(new_new_n5632__));
  buf1  g3448(.din(new_new_n3921__), .dout(new_new_n5633__));
  buf1  g3449(.din(new_new_n5633__), .dout(new_new_n5634__));
  buf1  g3450(.din(new_new_n3955__), .dout(new_new_n5635__));
  buf1  g3451(.din(new_new_n5635__), .dout(new_new_n5636__));
  buf1  g3452(.din(new_new_n5636__), .dout(new_new_n5637__));
  buf1  g3453(.din(new_new_n5636__), .dout(new_new_n5638__));
  buf1  g3454(.din(new_new_n5635__), .dout(new_new_n5639__));
  buf1  g3455(.din(new_new_n3923__), .dout(new_new_n5640__));
  buf1  g3456(.din(new_new_n5640__), .dout(new_new_n5641__));
  buf1  g3457(.din(new_new_n3957__), .dout(new_new_n5642__));
  buf1  g3458(.din(new_new_n5642__), .dout(new_new_n5643__));
  buf1  g3459(.din(new_new_n5643__), .dout(new_new_n5644__));
  buf1  g3460(.din(new_new_n5643__), .dout(new_new_n5645__));
  buf1  g3461(.din(new_new_n5642__), .dout(new_new_n5646__));
  buf1  g3462(.din(new_new_n3925__), .dout(new_new_n5647__));
  buf1  g3463(.din(new_new_n5647__), .dout(new_new_n5648__));
  buf1  g3464(.din(new_new_n3927__), .dout(new_new_n5649__));
  buf1  g3465(.din(new_new_n5649__), .dout(new_new_n5650__));
  buf1  g3466(.din(new_new_n3929__), .dout(new_new_n5651__));
  buf1  g3467(.din(new_new_n5651__), .dout(new_new_n5652__));
  buf1  g3468(.din(new_new_n3963__), .dout(new_new_n5653__));
  buf1  g3469(.din(new_new_n5653__), .dout(new_new_n5654__));
  buf1  g3470(.din(new_new_n3933__), .dout(new_new_n5655__));
  buf1  g3471(.din(new_new_n5655__), .dout(new_new_n5656__));
  buf1  g3472(.din(new_new_n3967__), .dout(new_new_n5657__));
  buf1  g3473(.din(new_new_n5657__), .dout(new_new_n5658__));
  buf1  g3474(.din(new_new_n3937__), .dout(new_new_n5659__));
  buf1  g3475(.din(new_new_n5659__), .dout(new_new_n5660__));
  buf1  g3476(.din(new_new_n3971__), .dout(new_new_n5661__));
  buf1  g3477(.din(new_new_n5661__), .dout(new_new_n5662__));
  buf1  g3478(.din(new_new_n3941__), .dout(new_new_n5663__));
  buf1  g3479(.din(new_new_n5663__), .dout(new_new_n5664__));
  buf1  g3480(.din(new_new_n3975__), .dout(new_new_n5665__));
  buf1  g3481(.din(new_new_n5665__), .dout(new_new_n5666__));
  buf1  g3482(.din(new_new_n3945__), .dout(new_new_n5667__));
  buf1  g3483(.din(new_new_n5667__), .dout(new_new_n5668__));
  buf1  g3484(.din(new_new_n2696__), .dout(new_new_n5669__));
  buf1  g3485(.din(new_new_n5669__), .dout(new_new_n5670__));
  buf1  g3486(.din(new_new_n5669__), .dout(new_new_n5671__));
  buf1  g3487(.din(new_new_n2698__), .dout(new_new_n5672__));
  buf1  g3488(.din(new_new_n5672__), .dout(new_new_n5673__));
  buf1  g3489(.din(new_new_n5672__), .dout(new_new_n5674__));
  buf1  g3490(.din(new_new_n2693__), .dout(new_new_n5675__));
  buf1  g3491(.din(new_new_n5675__), .dout(new_new_n5676__));
  buf1  g3492(.din(new_new_n5675__), .dout(new_new_n5677__));
  buf1  g3493(.din(new_new_n2695__), .dout(new_new_n5678__));
  buf1  g3494(.din(new_new_n5678__), .dout(new_new_n5679__));
  buf1  g3495(.din(new_new_n5678__), .dout(new_new_n5680__));
  buf1  g3496(.din(new_new_n2699__), .dout(new_new_n5681__));
  buf1  g3497(.din(new_new_n2697__), .dout(new_new_n5682__));
  buf1  g3498(.din(new_new_n2692__), .dout(new_new_n5683__));
  buf1  g3499(.din(new_new_n2694__), .dout(new_new_n5684__));
  buf1  g3500(.din(new_new_n3552__), .dout(new_new_n5685__));
  buf1  g3501(.din(new_new_n3558__), .dout(new_new_n5686__));
  buf1  g3502(.din(new_new_n3509__), .dout(new_new_n5687__));
  buf1  g3503(.din(new_new_n5687__), .dout(new_new_n5688__));
  buf1  g3504(.din(new_new_n5688__), .dout(new_new_n5689__));
  buf1  g3505(.din(new_new_n5688__), .dout(new_new_n5690__));
  buf1  g3506(.din(new_new_n5687__), .dout(new_new_n5691__));
  buf1  g3507(.din(new_new_n3508__), .dout(new_new_n5692__));
  buf1  g3508(.din(new_new_n3564__), .dout(new_new_n5693__));
  buf1  g3509(.din(new_new_n2438__), .dout(new_new_n5694__));
  buf1  g3510(.din(new_new_n5694__), .dout(new_new_n5695__));
  buf1  g3511(.din(new_new_n5694__), .dout(new_new_n5696__));
  buf1  g3512(.din(new_new_n2404__), .dout(new_new_n5697__));
  buf1  g3513(.din(new_new_n5697__), .dout(new_new_n5698__));
  buf1  g3514(.din(new_new_n5697__), .dout(new_new_n5699__));
  buf1  g3515(.din(new_new_n4001__), .dout(new_new_n5700__));
  buf1  g3516(.din(new_new_n5700__), .dout(new_new_n5701__));
  buf1  g3517(.din(new_new_n5701__), .dout(new_new_n5702__));
  buf1  g3518(.din(new_new_n5700__), .dout(new_new_n5703__));
  buf1  g3519(.din(new_new_n2353__), .dout(new_new_n5704__));
  buf1  g3520(.din(new_new_n5704__), .dout(new_new_n5705__));
  buf1  g3521(.din(new_new_n5705__), .dout(new_new_n5706__));
  buf1  g3522(.din(new_new_n5705__), .dout(new_new_n5707__));
  buf1  g3523(.din(new_new_n5704__), .dout(new_new_n5708__));
  buf1  g3524(.din(new_new_n5708__), .dout(new_new_n5709__));
  buf1  g3525(.din(new_new_n5708__), .dout(new_new_n5710__));
  buf1  g3526(.din(new_new_n2368__), .dout(new_new_n5711__));
  buf1  g3527(.din(new_new_n5711__), .dout(new_new_n5712__));
  buf1  g3528(.din(new_new_n5712__), .dout(new_new_n5713__));
  buf1  g3529(.din(new_new_n5713__), .dout(new_new_n5714__));
  buf1  g3530(.din(new_new_n5713__), .dout(new_new_n5715__));
  buf1  g3531(.din(new_new_n5712__), .dout(new_new_n5716__));
  buf1  g3532(.din(new_new_n5716__), .dout(new_new_n5717__));
  buf1  g3533(.din(new_new_n5716__), .dout(new_new_n5718__));
  buf1  g3534(.din(new_new_n5711__), .dout(new_new_n5719__));
  buf1  g3535(.din(new_new_n5719__), .dout(new_new_n5720__));
  buf1  g3536(.din(new_new_n5719__), .dout(new_new_n5721__));
  buf1  g3537(.din(new_new_n2369__), .dout(new_new_n5722__));
  buf1  g3538(.din(new_new_n5722__), .dout(new_new_n5723__));
  buf1  g3539(.din(new_new_n5723__), .dout(new_new_n5724__));
  buf1  g3540(.din(new_new_n5723__), .dout(new_new_n5725__));
  buf1  g3541(.din(new_new_n5722__), .dout(new_new_n5726__));
  buf1  g3542(.din(new_new_n5726__), .dout(new_new_n5727__));
  buf1  g3543(.din(new_new_n5726__), .dout(new_new_n5728__));
  buf1  g3544(.din(new_new_n2352__), .dout(new_new_n5729__));
  buf1  g3545(.din(new_new_n5729__), .dout(new_new_n5730__));
  buf1  g3546(.din(new_new_n5730__), .dout(new_new_n5731__));
  buf1  g3547(.din(new_new_n5731__), .dout(new_new_n5732__));
  buf1  g3548(.din(new_new_n5731__), .dout(new_new_n5733__));
  buf1  g3549(.din(new_new_n5730__), .dout(new_new_n5734__));
  buf1  g3550(.din(new_new_n5734__), .dout(new_new_n5735__));
  buf1  g3551(.din(new_new_n5734__), .dout(new_new_n5736__));
  buf1  g3552(.din(new_new_n5729__), .dout(new_new_n5737__));
  buf1  g3553(.din(new_new_n5737__), .dout(new_new_n5738__));
  buf1  g3554(.din(new_new_n5737__), .dout(new_new_n5739__));
  buf1  g3555(.din(new_new_n2401__), .dout(new_new_n5740__));
  buf1  g3556(.din(new_new_n2447__), .dout(new_new_n5741__));
  buf1  g3557(.din(new_new_n5741__), .dout(new_new_n5742__));
  buf1  g3558(.din(new_new_n3259__), .dout(new_new_n5743__));
  buf1  g3559(.din(new_new_n3273__), .dout(new_new_n5744__));
  buf1  g3560(.din(new_new_n3276__), .dout(new_new_n5745__));
  buf1  g3561(.din(new_new_n3282__), .dout(new_new_n5746__));
  buf1  g3562(.din(new_new_n3396__), .dout(new_new_n5747__));
  buf1  g3563(.din(new_new_n3430__), .dout(new_new_n5748__));
  buf1  g3564(.din(new_new_n3443__), .dout(new_new_n5749__));
  buf1  g3565(.din(new_new_n2472__), .dout(new_new_n5750__));
  buf1  g3566(.din(new_new_n5750__), .dout(new_new_n5751__));
  buf1  g3567(.din(new_new_n2480__), .dout(new_new_n5752__));
  buf1  g3568(.din(new_new_n5752__), .dout(new_new_n5753__));
  buf1  g3569(.din(new_new_n2808__), .dout(new_new_n5754__));
  buf1  g3570(.din(new_new_n5754__), .dout(new_new_n5755__));
  buf1  g3571(.din(new_new_n2414__), .dout(new_new_n5756__));
  buf1  g3572(.din(new_new_n2434__), .dout(new_new_n5757__));
  buf1  g3573(.din(new_new_n2456__), .dout(new_new_n5758__));
  buf1  g3574(.din(new_new_n2430__), .dout(new_new_n5759__));
  buf1  g3575(.din(new_new_n3531__), .dout(new_new_n5760__));
  buf1  g3576(.din(new_new_n5760__), .dout(new_new_n5761__));
  buf1  g3577(.din(new_new_n5761__), .dout(new_new_n5762__));
  buf1  g3578(.din(new_new_n5760__), .dout(new_new_n5763__));
  buf1  g3579(.din(new_new_n3764__), .dout(new_new_n5764__));
  buf1  g3580(.din(new_new_n3767__), .dout(new_new_n5765__));
  buf1  g3581(.din(new_new_n3794__), .dout(new_new_n5766__));
  buf1  g3582(.din(new_new_n3809__), .dout(new_new_n5767__));
  buf1  g3583(.din(new_new_n3812__), .dout(new_new_n5768__));
  buf1  g3584(.din(new_new_n3841__), .dout(new_new_n5769__));
  buf1  g3585(.din(new_new_n3870__), .dout(new_new_n5770__));
  buf1  g3586(.din(new_new_n3899__), .dout(new_new_n5771__));
  buf1  g3587(.din(new_new_n3977__), .dout(new_new_n5772__));
  buf1  g3588(.din(new_new_n5772__), .dout(new_new_n5773__));
  buf1  g3589(.din(new_new_n3979__), .dout(new_new_n5774__));
  buf1  g3590(.din(new_new_n5774__), .dout(new_new_n5775__));
  buf1  g3591(.din(new_new_n3990__), .dout(new_new_n5776__));
  buf1  g3592(.din(new_new_n5776__), .dout(new_new_n5777__));
  buf1  g3593(.din(new_new_n4012__), .dout(new_new_n5778__));
  buf1  g3594(.din(new_new_n5778__), .dout(new_new_n5779__));
  buf1  g3595(.din(new_new_n4014__), .dout(new_new_n5780__));
  buf1  g3596(.din(new_new_n5780__), .dout(new_new_n5781__));
  buf1  g3597(.din(new_new_n5781__), .dout(new_new_n5782__));
  buf1  g3598(.din(new_new_n5781__), .dout(new_new_n5783__));
  buf1  g3599(.din(new_new_n5780__), .dout(new_new_n5784__));
  buf1  g3600(.din(new_new_n2510__), .dout(new_new_n5785__));
  buf1  g3601(.din(new_new_n2514__), .dout(new_new_n5786__));
  buf1  g3602(.din(new_new_n4154__), .dout(new_new_n5787__));
  buf1  g3603(.din(new_new_n5787__), .dout(new_new_n5788__));
  buf1  g3604(.din(new_new_n5788__), .dout(new_new_n5789__));
  buf1  g3605(.din(new_new_n5787__), .dout(new_new_n5790__));
  always @ (posedge clock) begin
    n1416_lo <= n8268;
    n1419_lo <= n8271;
    n1422_lo <= n8274;
    n1425_lo <= n8277;
    n1428_lo <= n8280;
    n1431_lo <= n8283;
    n1434_lo <= n8286;
    n1437_lo <= n8289;
    n1440_lo <= n8292;
    n1443_lo <= n8295;
    n1446_lo <= n8298;
    n1449_lo <= n8301;
    n1452_lo <= n8304;
    n1455_lo <= n8307;
    n1458_lo <= n8310;
    n1464_lo <= n8313;
    n1467_lo <= n8316;
    n1470_lo <= n8319;
    n1476_lo <= n8322;
    n1479_lo <= n8325;
    n1482_lo <= n8328;
    n1488_lo <= n8331;
    n1491_lo <= n8334;
    n1494_lo <= n8337;
    n1497_lo <= n8340;
    n1500_lo <= n8343;
    n1512_lo <= n8346;
    n1515_lo <= n8349;
    n1518_lo <= n8352;
    n1521_lo <= n8355;
    n1524_lo <= n8358;
    n1527_lo <= n8361;
    n1530_lo <= n8364;
    n1533_lo <= n8367;
    n1536_lo <= n8370;
    n1539_lo <= n8373;
    n1542_lo <= n8376;
    n1545_lo <= n8379;
    n1548_lo <= n8382;
    n1551_lo <= n8385;
    n1554_lo <= n8388;
    n1560_lo <= n8391;
    n1563_lo <= n8394;
    n1566_lo <= n8397;
    n1572_lo <= n8400;
    n1575_lo <= n8403;
    n1578_lo <= n8406;
    n1584_lo <= n8409;
    n1587_lo <= n8412;
    n1590_lo <= n8415;
    n1596_lo <= n8418;
    n1599_lo <= n8421;
    n1602_lo <= n8424;
    n1608_lo <= n8427;
    n1611_lo <= n8430;
    n1614_lo <= n8433;
    n1620_lo <= n8436;
    n1623_lo <= n8439;
    n1626_lo <= n8442;
    n1632_lo <= n8445;
    n1635_lo <= n8448;
    n1638_lo <= n8451;
    n1644_lo <= n8454;
    n1647_lo <= n8457;
    n1650_lo <= n8460;
    n1656_lo <= n8463;
    n1659_lo <= n8466;
    n1662_lo <= n8469;
    n1668_lo <= n8472;
    n1671_lo <= n8475;
    n1674_lo <= n8478;
    n1677_lo <= n8481;
    n1680_lo <= n8484;
    n1683_lo <= n8487;
    n1686_lo <= n8490;
    n1692_lo <= n8493;
    n1695_lo <= n8496;
    n1698_lo <= n8499;
    n1704_lo <= n8502;
    n1707_lo <= n8505;
    n1710_lo <= n8508;
    n1716_lo <= n8511;
    n1719_lo <= n8514;
    n1722_lo <= n8517;
    n1728_lo <= n8520;
    n1731_lo <= n8523;
    n1734_lo <= n8526;
    n1740_lo <= n8529;
    n1743_lo <= n8532;
    n1746_lo <= n8535;
    n1749_lo <= n8538;
    n1752_lo <= n8541;
    n1755_lo <= n8544;
    n1758_lo <= n8547;
    n1761_lo <= n8550;
    n1764_lo <= n8553;
    n1776_lo <= n8556;
    n1779_lo <= n8559;
    n1788_lo <= n8562;
    n1791_lo <= n8565;
    n1794_lo <= n8568;
    n1797_lo <= n8571;
    n1800_lo <= n8574;
    n1812_lo <= n8577;
    n1824_lo <= n8580;
    n1836_lo <= n8583;
    n1848_lo <= n8586;
    n1860_lo <= n8589;
    n1872_lo <= n8592;
    n1884_lo <= n8595;
    n1896_lo <= n8598;
    n1899_lo <= n8601;
    n1908_lo <= n8604;
    n1911_lo <= n8607;
    n1920_lo <= n8610;
    n1923_lo <= n8613;
    n1926_lo <= n8616;
    n1929_lo <= n8619;
    n1932_lo <= n8622;
    n1944_lo <= n8625;
    n1956_lo <= n8628;
    n1968_lo <= n8631;
    n1980_lo <= n8634;
    n1992_lo <= n8637;
    n2004_lo <= n8640;
    n2016_lo <= n8643;
    n2019_lo <= n8646;
    n2028_lo <= n8649;
    n2031_lo <= n8652;
    n2040_lo <= n8655;
    n2043_lo <= n8658;
    n2046_lo <= n8661;
    n2049_lo <= n8664;
    n2052_lo <= n8667;
    n2064_lo <= n8670;
    n2076_lo <= n8673;
    n2088_lo <= n8676;
    n2100_lo <= n8679;
    n2112_lo <= n8682;
    n2124_lo <= n8685;
    n2136_lo <= n8688;
    n2148_lo <= n8691;
    n2151_lo <= n8694;
    n2160_lo <= n8697;
    n2163_lo <= n8700;
    n2172_lo <= n8703;
    n2175_lo <= n8706;
    n2178_lo <= n8709;
    n2181_lo <= n8712;
    n2184_lo <= n8715;
    n2196_lo <= n8718;
    n2208_lo <= n8721;
    n2220_lo <= n8724;
    n2232_lo <= n8727;
    n2244_lo <= n8730;
    n2256_lo <= n8733;
    n2268_lo <= n8736;
    n2280_lo <= n8739;
    n2283_lo <= n8742;
    n2292_lo <= n8745;
    n2295_lo <= n8748;
    n2298_lo <= n8751;
    n2301_lo <= n8754;
    n2304_lo <= n8757;
    n2316_lo <= n8760;
    n2319_lo <= n8763;
    n2322_lo <= n8766;
    n2325_lo <= n8769;
    n2328_lo <= n8772;
    n2331_lo <= n8775;
    n2340_lo <= n8778;
    n2343_lo <= n8781;
    n2376_lo <= n8784;
    n2379_lo <= n8787;
    n2388_lo <= n8790;
    n2400_lo <= n8793;
    n2412_lo <= n8796;
    n2415_lo <= n8799;
    n2424_lo <= n8802;
    n2436_lo <= n8805;
    n2439_lo <= n8808;
    n2442_lo <= n8811;
    n2445_lo <= n8814;
    n2448_lo <= n8817;
    n2451_lo <= n8820;
    n2460_lo <= n8823;
    n2463_lo <= n8826;
    n2496_lo <= n8829;
    n2499_lo <= n8832;
    n2508_lo <= n8835;
    n2520_lo <= n8838;
    n2532_lo <= n8841;
    n2535_lo <= n8844;
    n2544_lo <= n8847;
    n2556_lo <= n8850;
    n2559_lo <= n8853;
    n2562_lo <= n8856;
    n2565_lo <= n8859;
    n2568_lo <= n8862;
    n2571_lo <= n8865;
    n2580_lo <= n8868;
    n2583_lo <= n8871;
    n2616_lo <= n8874;
    n2619_lo <= n8877;
    n2628_lo <= n8880;
    n2640_lo <= n8883;
    n2652_lo <= n8886;
    n2655_lo <= n8889;
    n2664_lo <= n8892;
    n2676_lo <= n8895;
    n2679_lo <= n8898;
    n2682_lo <= n8901;
    n2685_lo <= n8904;
    n2688_lo <= n8907;
    n2691_lo <= n8910;
    n2700_lo <= n8913;
    n2703_lo <= n8916;
    n2736_lo <= n8919;
    n2739_lo <= n8922;
    n2748_lo <= n8925;
    n2760_lo <= n8928;
    n2772_lo <= n8931;
    n2775_lo <= n8934;
    n2784_lo <= n8937;
    n2787_lo <= n8940;
    n2790_lo <= n8943;
    n2793_lo <= n8946;
    n2796_lo <= n8949;
    n2799_lo <= n8952;
    n2802_lo <= n8955;
    n2805_lo <= n8958;
    n2808_lo <= n8961;
    n2820_lo <= n8964;
    n2823_lo <= n8967;
    n2826_lo <= n8970;
    n2832_lo <= n8973;
    n2835_lo <= n8976;
    n2838_lo <= n8979;
    n2841_lo <= n8982;
    n2844_lo <= n8985;
    n2856_lo <= n8988;
    n2859_lo <= n8991;
    n2862_lo <= n8994;
    n2865_lo <= n8997;
    n2868_lo <= n9000;
    n2871_lo <= n9003;
    n2874_lo <= n9006;
    n2877_lo <= n9009;
    n2880_lo <= n9012;
    n2883_lo <= n9015;
    n2886_lo <= n9018;
    n2889_lo <= n9021;
    n2892_lo <= n9024;
    n2895_lo <= n9027;
    n2898_lo <= n9030;
    n2901_lo <= n9033;
    n2904_lo <= n9036;
    n2907_lo <= n9039;
    n2916_lo <= n9042;
    n2928_lo <= n9045;
    n2940_lo <= n9048;
    n2952_lo <= n9051;
    n2955_lo <= n9054;
    n2964_lo <= n9057;
    n2976_lo <= n9060;
    n2988_lo <= n9063;
    n2991_lo <= n9066;
    n3000_lo <= n9069;
    n3003_lo <= n9072;
    n3012_lo <= n9075;
    n3015_lo <= n9078;
    n3024_lo <= n9081;
    n3027_lo <= n9084;
    n3036_lo <= n9087;
    n3039_lo <= n9090;
    n3048_lo <= n9093;
    n3051_lo <= n9096;
    n3054_lo <= n9099;
    n3057_lo <= n9102;
    n3060_lo <= n9105;
    n3072_lo <= n9108;
    n3081_lo <= n9111;
    n3084_lo <= n9114;
    n3087_lo <= n9117;
    n3093_lo <= n9120;
    n3096_lo <= n9123;
    n3105_lo <= n9126;
    n3108_lo <= n9129;
    n3117_lo <= n9132;
    n3120_lo <= n9135;
    n3123_lo <= n9138;
    n3126_lo <= n9141;
    n3129_lo <= n9144;
    n3132_lo <= n9147;
    n3135_lo <= n9150;
    n3138_lo <= n9153;
    n3141_lo <= n9156;
    n3168_lo <= n9159;
    n3171_lo <= n9162;
    n3174_lo <= n9165;
    n3177_lo <= n9168;
    n3180_lo <= n9171;
    n3183_lo <= n9174;
    n3192_lo <= n9177;
    n3195_lo <= n9180;
    n3204_lo <= n9183;
    n3207_lo <= n9186;
    n3216_lo <= n9189;
    n3219_lo <= n9192;
    n3228_lo <= n9195;
    n3231_lo <= n9198;
    n3240_lo <= n9201;
    n3243_lo <= n9204;
    n3252_lo <= n9207;
    n3255_lo <= n9210;
    n3258_lo <= n9213;
    n3264_lo <= n9216;
    n3267_lo <= n9219;
    n3270_lo <= n9222;
    n3276_lo <= n9225;
    n3279_lo <= n9228;
    n3282_lo <= n9231;
    n3288_lo <= n9234;
    n3291_lo <= n9237;
    n3294_lo <= n9240;
    n4537_o2 <= n9243;
    n4538_o2 <= n9246;
    n4710_o2 <= n9249;
    n4711_o2 <= n9252;
    n1211_inv <= n9255;
    n1214_inv <= n9258;
    n1217_inv <= n9261;
    n1220_inv <= n9264;
    n4927_o2 <= n9267;
    n4928_o2 <= n9270;
    n1229_inv <= n9273;
    n1232_inv <= n9276;
    n1235_inv <= n9279;
    n5178_o2 <= n9282;
    n5179_o2 <= n9285;
    n5477_o2 <= n9288;
    n5478_o2 <= n9291;
    n5479_o2 <= n9294;
    n5222_o2 <= n9297;
    n5223_o2 <= n9300;
    n5553_o2 <= n9303;
    n5554_o2 <= n9306;
    G491_o2 <= n9309;
    n2922_lo_buf_o2 <= n9312;
    n2946_lo_buf_o2 <= n9315;
    n2970_lo_buf_o2 <= n9318;
    n2982_lo_buf_o2 <= n9321;
    n3066_lo_buf_o2 <= n9324;
    n3078_lo_buf_o2 <= n9327;
    n3102_lo_buf_o2 <= n9330;
    n3114_lo_buf_o2 <= n9333;
    G1321_o2 <= n9336;
    G1033_o2 <= n9339;
    G1030_o2 <= n9342;
    G1072_o2 <= n9345;
    n1304_inv <= n9348;
    n1307_inv <= n9351;
    n2958_lo_buf_o2 <= n9354;
    n2994_lo_buf_o2 <= n9357;
    n3006_lo_buf_o2 <= n9360;
    n3030_lo_buf_o2 <= n9363;
    n3042_lo_buf_o2 <= n9366;
    n3090_lo_buf_o2 <= n9369;
    n1328_inv <= n9372;
    n1331_inv <= n9375;
    n1334_inv <= n9378;
    n1337_inv <= n9381;
    n1340_inv <= n9384;
    n1343_inv <= n9387;
    n1346_inv <= n9390;
    n1349_inv <= n9393;
    G1036_o2 <= n9396;
    G1062_o2 <= n9399;
    G1067_o2 <= n9402;
    G1014_o2 <= n9405;
    n1364_inv <= n9408;
    n1367_inv <= n9411;
    n3018_lo_buf_o2 <= n9414;
    G766_o2 <= n9417;
    n1376_inv <= n9420;
    n1379_inv <= n9423;
    n1382_inv <= n9426;
    n1385_inv <= n9429;
    n1388_inv <= n9432;
    n1391_inv <= n9435;
    G1017_o2 <= n9438;
    G1008_o2 <= n9441;
    n1400_inv <= n9444;
    n1403_inv <= n9447;
    n2910_lo_buf_o2 <= n9450;
    n1409_inv <= n9453;
    G2138_o2 <= n9456;
    G2147_o2 <= n9459;
    n1418_inv <= n9462;
    G1137_o2 <= n9465;
    G1329_o2 <= n9468;
    G374_o2 <= n9471;
    G386_o2 <= n9474;
    G663_o2 <= n9477;
    G674_o2 <= n9480;
    G578_o2 <= n9483;
    G575_o2 <= n9486;
    G2505_o2 <= n9489;
    n1448_inv <= n9492;
    G987_o2 <= n9495;
    G984_o2 <= n9498;
    G1862_o2 <= n9501;
    G1859_o2 <= n9504;
    G1260_o2 <= n9507;
    G1865_o2 <= n9510;
    G2073_o2 <= n9513;
    G1402_o2 <= n9516;
    G2048_o2 <= n9519;
    G2276_o2 <= n9522;
    n1481_inv <= n9525;
    G2141_o2 <= n9528;
    G2008_o2 <= n9531;
    G2011_o2 <= n9534;
    G2150_o2 <= n9537;
    G2026_o2 <= n9540;
    G2029_o2 <= n9543;
    G2023_o2 <= n9546;
    G2041_o2 <= n9549;
    G2017_o2 <= n9552;
    G2020_o2 <= n9555;
    G2035_o2 <= n9558;
    G2038_o2 <= n9561;
    G2228_o2 <= n9564;
    G2231_o2 <= n9567;
    G2234_o2 <= n9570;
    G2237_o2 <= n9573;
    G1904_o2 <= n9576;
    G1907_o2 <= n9579;
    G1928_o2 <= n9582;
    G1931_o2 <= n9585;
    G1893_o2 <= n9588;
    G1896_o2 <= n9591;
    G1899_o2 <= n9594;
    G1937_o2 <= n9597;
    G1940_o2 <= n9600;
    G1943_o2 <= n9603;
    G1336_o2 <= n9606;
    G1996_o2 <= n9609;
    G1999_o2 <= n9612;
    G2002_o2 <= n9615;
    G2005_o2 <= n9618;
    G2014_o2 <= n9621;
    G2032_o2 <= n9624;
    G1076_o2 <= n9627;
    G1002_o2 <= n9630;
    G998_o2 <= n9633;
    G1890_o2 <= n9636;
    G1934_o2 <= n9639;
    G1044_o2 <= n9642;
    G1039_o2 <= n9645;
    n1770_lo_buf_o2 <= n9648;
    G342_o2 <= n9651;
    G354_o2 <= n9654;
    G1193_o2 <= n9657;
    n3234_lo_buf_o2 <= n9660;
    n3246_lo_buf_o2 <= n9663;
    G783_o2 <= n9666;
    G786_o2 <= n9669;
    G792_o2 <= n9672;
    G795_o2 <= n9675;
    G815_o2 <= n9678;
    G818_o2 <= n9681;
    G824_o2 <= n9684;
    G827_o2 <= n9687;
    G789_o2 <= n9690;
    G798_o2 <= n9693;
    G801_o2 <= n9696;
    G807_o2 <= n9699;
    G812_o2 <= n9702;
    G821_o2 <= n9705;
    G804_o2 <= n9708;
    G780_o2 <= n9711;
    G1231_o2 <= n9714;
    G1572_o2 <= n9717;
    G1377_o2 <= n9720;
    G1253_o2 <= n9723;
    G1359_o2 <= n9726;
    G1258_o2 <= n9729;
    G1367_o2 <= n9732;
    G1358_o2 <= n9735;
    G1366_o2 <= n9738;
    G2057_o2 <= n9741;
    G2117_o2 <= n9744;
    G2118_o2 <= n9747;
    G1254_o2 <= n9750;
    G1259_o2 <= n9753;
    G2058_o2 <= n9756;
    G405_o2 <= n9759;
    G417_o2 <= n9762;
    G1269_o2 <= n9765;
    G1275_o2 <= n9768;
    G1287_o2 <= n9771;
    G1266_o2 <= n9774;
    G1272_o2 <= n9777;
    G1278_o2 <= n9780;
    G1281_o2 <= n9783;
    G1284_o2 <= n9786;
    G1290_o2 <= n9789;
    G1293_o2 <= n9792;
    G1299_o2 <= n9795;
    G1305_o2 <= n9798;
    G1296_o2 <= n9801;
    G1302_o2 <= n9804;
    G1308_o2 <= n9807;
    G1311_o2 <= n9810;
    G811_o2 <= n9813;
    G810_o2 <= n9816;
    G1728_o2 <= n9819;
    G2512_o2 <= n9822;
    G1114_o2 <= n9825;
    G1113_o2 <= n9828;
    G1992_o2 <= n9831;
    G1991_o2 <= n9834;
    G1426_o2 <= n9837;
    G1966_o2 <= n9840;
    G2211_o2 <= n9843;
    G1509_o2 <= n9846;
    G2153_o2 <= n9849;
    G2329_o2 <= n9852;
    G1540_o2 <= n9855;
    G2167_o2 <= n9858;
    G2191_o2 <= n9861;
    G1234_o2 <= n9864;
    G1132_o2 <= n9867;
    G1129_o2 <= n9870;
    G2088_o2 <= n9873;
    G2106_o2 <= n9876;
    G1314_o2 <= n9879;
    G636_o2 <= n9882;
    G647_o2 <= n9885;
    n3186_lo_buf_o2 <= n9888;
    n3198_lo_buf_o2 <= n9891;
    n3210_lo_buf_o2 <= n9894;
    n3222_lo_buf_o2 <= n9897;
    G1225_o2 <= n9900;
    G1342_o2 <= n9903;
    G1222_o2 <= n9906;
    G1228_o2 <= n9909;
    G1348_o2 <= n9912;
    G1345_o2 <= n9915;
    G1351_o2 <= n9918;
    G2242_o2 <= n9921;
    G2260_o2 <= n9924;
    G1374_o2 <= n9927;
    G1537_o2 <= n9930;
    G301_o2 <= n9933;
    G313_o2 <= n9936;
    G2365_o2 <= n9939;
    G2255_o2 <= n9942;
    G2253_o2 <= n9945;
    G2395_o2 <= n9948;
    G2272_o2 <= n9951;
    G2270_o2 <= n9954;
    G2245_o2 <= n9957;
    G2262_o2 <= n9960;
    G2249_o2 <= n9963;
    G2247_o2 <= n9966;
    G2266_o2 <= n9969;
    G2264_o2 <= n9972;
    G2403_o2 <= n9975;
    G2401_o2 <= n9978;
    G2410_o2 <= n9981;
    G2408_o2 <= n9984;
    G2306_o2 <= n9987;
    G2305_o2 <= n9990;
    G2314_o2 <= n9993;
    G2313_o2 <= n9996;
    G2303_o2 <= n9999;
    G2302_o2 <= n10002;
    G2301_o2 <= n10005;
    G2311_o2 <= n10008;
    G2310_o2 <= n10011;
    G2309_o2 <= n10014;
    G2404_o2 <= n10017;
    G2411_o2 <= n10020;
    G2420_o2 <= n10023;
    G2419_o2 <= n10026;
    G2433_o2 <= n10029;
    G2432_o2 <= n10032;
    G402_o2 <= n10035;
    G403_o2 <= n10038;
    G1053_o2 <= n10041;
    G1049_o2 <= n10044;
    n2003_inv <= n10047;
    G1364_o2 <= n10050;
    G1079_o2 <= n10053;
    G1478_o2 <= n10056;
    G707_o2 <= n10059;
    G718_o2 <= n10062;
    G2417_o2 <= n10065;
    G2414_o2 <= n10068;
    G2431_o2 <= n10071;
    G2428_o2 <= n10074;
    G1653_o2 <= n10077;
    G2213_o2 <= n10080;
    G2221_o2 <= n10083;
    G2250_o2 <= n10086;
    G2267_o2 <= n10089;
    G1365_o2 <= n10092;
    G1368_o2 <= n10095;
    G1371_o2 <= n10098;
    G2218_o2 <= n10101;
    G2225_o2 <= n10104;
    n1503_lo_buf_o2 <= n10107;
    n1863_lo_buf_o2 <= n10110;
    n1887_lo_buf_o2 <= n10113;
    n1983_lo_buf_o2 <= n10116;
    n2007_lo_buf_o2 <= n10119;
    n2115_lo_buf_o2 <= n10122;
    n2139_lo_buf_o2 <= n10125;
    n2247_lo_buf_o2 <= n10128;
    n2271_lo_buf_o2 <= n10131;
    n2919_lo_buf_o2 <= n10134;
    n2943_lo_buf_o2 <= n10137;
    n2967_lo_buf_o2 <= n10140;
    n2979_lo_buf_o2 <= n10143;
    n3063_lo_buf_o2 <= n10146;
    n3075_lo_buf_o2 <= n10149;
    n3099_lo_buf_o2 <= n10152;
    n3111_lo_buf_o2 <= n10155;
    G878_o2 <= n10158;
    G875_o2 <= n10161;
    G661_o2 <= n10164;
    G660_o2 <= n10167;
    G879_o2 <= n10170;
    G876_o2 <= n10173;
    G1320_o2 <= n10176;
    G941_o2 <= n10179;
    G732_o2 <= n10182;
    G942_o2 <= n10185;
    G1493_o2 <= n10188;
    G1498_o2 <= n10191;
    G877_o2 <= n10194;
    G874_o2 <= n10197;
    n1806_lo_buf_o2 <= n10200;
    n1878_lo_buf_o2 <= n10203;
    n1938_lo_buf_o2 <= n10206;
    n1998_lo_buf_o2 <= n10209;
    n2058_lo_buf_o2 <= n10212;
    n2130_lo_buf_o2 <= n10215;
    n2190_lo_buf_o2 <= n10218;
    n2262_lo_buf_o2 <= n10221;
    n2310_lo_buf_o2 <= n10224;
    n2406_lo_buf_o2 <= n10227;
    n2430_lo_buf_o2 <= n10230;
    n2526_lo_buf_o2 <= n10233;
    n2550_lo_buf_o2 <= n10236;
    n2646_lo_buf_o2 <= n10239;
    n2670_lo_buf_o2 <= n10242;
    n2766_lo_buf_o2 <= n10245;
    G603_o2 <= n10248;
    G614_o2 <= n10251;
    G1026_o2 <= n10254;
    G1021_o2 <= n10257;
    G940_o2 <= n10260;
    G1636_o2 <= n10263;
    G1684_o2 <= n10266;
    n2352_lo_buf_o2 <= n10269;
    n2364_lo_buf_o2 <= n10272;
    n2472_lo_buf_o2 <= n10275;
    n2484_lo_buf_o2 <= n10278;
    n2592_lo_buf_o2 <= n10281;
    n2604_lo_buf_o2 <= n10284;
    n2712_lo_buf_o2 <= n10287;
    n2724_lo_buf_o2 <= n10290;
    n3150_lo_buf_o2 <= n10293;
    n3162_lo_buf_o2 <= n10296;
  end
  initial begin
    n1416_lo <= 1'b0;
    n1419_lo <= 1'b0;
    n1422_lo <= 1'b0;
    n1425_lo <= 1'b0;
    n1428_lo <= 1'b0;
    n1431_lo <= 1'b0;
    n1434_lo <= 1'b0;
    n1437_lo <= 1'b0;
    n1440_lo <= 1'b0;
    n1443_lo <= 1'b0;
    n1446_lo <= 1'b0;
    n1449_lo <= 1'b0;
    n1452_lo <= 1'b0;
    n1455_lo <= 1'b0;
    n1458_lo <= 1'b0;
    n1464_lo <= 1'b0;
    n1467_lo <= 1'b0;
    n1470_lo <= 1'b0;
    n1476_lo <= 1'b0;
    n1479_lo <= 1'b0;
    n1482_lo <= 1'b0;
    n1488_lo <= 1'b0;
    n1491_lo <= 1'b0;
    n1494_lo <= 1'b0;
    n1497_lo <= 1'b0;
    n1500_lo <= 1'b0;
    n1512_lo <= 1'b0;
    n1515_lo <= 1'b0;
    n1518_lo <= 1'b0;
    n1521_lo <= 1'b0;
    n1524_lo <= 1'b0;
    n1527_lo <= 1'b0;
    n1530_lo <= 1'b0;
    n1533_lo <= 1'b0;
    n1536_lo <= 1'b0;
    n1539_lo <= 1'b0;
    n1542_lo <= 1'b0;
    n1545_lo <= 1'b0;
    n1548_lo <= 1'b0;
    n1551_lo <= 1'b0;
    n1554_lo <= 1'b0;
    n1560_lo <= 1'b0;
    n1563_lo <= 1'b0;
    n1566_lo <= 1'b0;
    n1572_lo <= 1'b0;
    n1575_lo <= 1'b0;
    n1578_lo <= 1'b0;
    n1584_lo <= 1'b0;
    n1587_lo <= 1'b0;
    n1590_lo <= 1'b0;
    n1596_lo <= 1'b0;
    n1599_lo <= 1'b0;
    n1602_lo <= 1'b0;
    n1608_lo <= 1'b0;
    n1611_lo <= 1'b0;
    n1614_lo <= 1'b0;
    n1620_lo <= 1'b0;
    n1623_lo <= 1'b0;
    n1626_lo <= 1'b0;
    n1632_lo <= 1'b0;
    n1635_lo <= 1'b0;
    n1638_lo <= 1'b0;
    n1644_lo <= 1'b0;
    n1647_lo <= 1'b0;
    n1650_lo <= 1'b0;
    n1656_lo <= 1'b0;
    n1659_lo <= 1'b0;
    n1662_lo <= 1'b0;
    n1668_lo <= 1'b0;
    n1671_lo <= 1'b0;
    n1674_lo <= 1'b0;
    n1677_lo <= 1'b0;
    n1680_lo <= 1'b0;
    n1683_lo <= 1'b0;
    n1686_lo <= 1'b0;
    n1692_lo <= 1'b0;
    n1695_lo <= 1'b0;
    n1698_lo <= 1'b0;
    n1704_lo <= 1'b0;
    n1707_lo <= 1'b0;
    n1710_lo <= 1'b0;
    n1716_lo <= 1'b0;
    n1719_lo <= 1'b0;
    n1722_lo <= 1'b0;
    n1728_lo <= 1'b0;
    n1731_lo <= 1'b0;
    n1734_lo <= 1'b0;
    n1740_lo <= 1'b0;
    n1743_lo <= 1'b0;
    n1746_lo <= 1'b0;
    n1749_lo <= 1'b0;
    n1752_lo <= 1'b0;
    n1755_lo <= 1'b0;
    n1758_lo <= 1'b0;
    n1761_lo <= 1'b0;
    n1764_lo <= 1'b0;
    n1776_lo <= 1'b0;
    n1779_lo <= 1'b0;
    n1788_lo <= 1'b0;
    n1791_lo <= 1'b0;
    n1794_lo <= 1'b0;
    n1797_lo <= 1'b0;
    n1800_lo <= 1'b0;
    n1812_lo <= 1'b0;
    n1824_lo <= 1'b0;
    n1836_lo <= 1'b0;
    n1848_lo <= 1'b0;
    n1860_lo <= 1'b0;
    n1872_lo <= 1'b0;
    n1884_lo <= 1'b0;
    n1896_lo <= 1'b0;
    n1899_lo <= 1'b0;
    n1908_lo <= 1'b0;
    n1911_lo <= 1'b0;
    n1920_lo <= 1'b0;
    n1923_lo <= 1'b0;
    n1926_lo <= 1'b0;
    n1929_lo <= 1'b0;
    n1932_lo <= 1'b0;
    n1944_lo <= 1'b0;
    n1956_lo <= 1'b0;
    n1968_lo <= 1'b0;
    n1980_lo <= 1'b0;
    n1992_lo <= 1'b0;
    n2004_lo <= 1'b0;
    n2016_lo <= 1'b0;
    n2019_lo <= 1'b0;
    n2028_lo <= 1'b0;
    n2031_lo <= 1'b0;
    n2040_lo <= 1'b0;
    n2043_lo <= 1'b0;
    n2046_lo <= 1'b0;
    n2049_lo <= 1'b0;
    n2052_lo <= 1'b0;
    n2064_lo <= 1'b0;
    n2076_lo <= 1'b0;
    n2088_lo <= 1'b0;
    n2100_lo <= 1'b0;
    n2112_lo <= 1'b0;
    n2124_lo <= 1'b0;
    n2136_lo <= 1'b0;
    n2148_lo <= 1'b0;
    n2151_lo <= 1'b0;
    n2160_lo <= 1'b0;
    n2163_lo <= 1'b0;
    n2172_lo <= 1'b0;
    n2175_lo <= 1'b0;
    n2178_lo <= 1'b0;
    n2181_lo <= 1'b0;
    n2184_lo <= 1'b0;
    n2196_lo <= 1'b0;
    n2208_lo <= 1'b0;
    n2220_lo <= 1'b0;
    n2232_lo <= 1'b0;
    n2244_lo <= 1'b0;
    n2256_lo <= 1'b0;
    n2268_lo <= 1'b0;
    n2280_lo <= 1'b0;
    n2283_lo <= 1'b0;
    n2292_lo <= 1'b0;
    n2295_lo <= 1'b0;
    n2298_lo <= 1'b0;
    n2301_lo <= 1'b0;
    n2304_lo <= 1'b0;
    n2316_lo <= 1'b0;
    n2319_lo <= 1'b0;
    n2322_lo <= 1'b0;
    n2325_lo <= 1'b0;
    n2328_lo <= 1'b0;
    n2331_lo <= 1'b0;
    n2340_lo <= 1'b0;
    n2343_lo <= 1'b0;
    n2376_lo <= 1'b0;
    n2379_lo <= 1'b0;
    n2388_lo <= 1'b0;
    n2400_lo <= 1'b0;
    n2412_lo <= 1'b0;
    n2415_lo <= 1'b0;
    n2424_lo <= 1'b0;
    n2436_lo <= 1'b0;
    n2439_lo <= 1'b0;
    n2442_lo <= 1'b0;
    n2445_lo <= 1'b0;
    n2448_lo <= 1'b0;
    n2451_lo <= 1'b0;
    n2460_lo <= 1'b0;
    n2463_lo <= 1'b0;
    n2496_lo <= 1'b0;
    n2499_lo <= 1'b0;
    n2508_lo <= 1'b0;
    n2520_lo <= 1'b0;
    n2532_lo <= 1'b0;
    n2535_lo <= 1'b0;
    n2544_lo <= 1'b0;
    n2556_lo <= 1'b0;
    n2559_lo <= 1'b0;
    n2562_lo <= 1'b0;
    n2565_lo <= 1'b0;
    n2568_lo <= 1'b0;
    n2571_lo <= 1'b0;
    n2580_lo <= 1'b0;
    n2583_lo <= 1'b0;
    n2616_lo <= 1'b0;
    n2619_lo <= 1'b0;
    n2628_lo <= 1'b0;
    n2640_lo <= 1'b0;
    n2652_lo <= 1'b0;
    n2655_lo <= 1'b0;
    n2664_lo <= 1'b0;
    n2676_lo <= 1'b0;
    n2679_lo <= 1'b0;
    n2682_lo <= 1'b0;
    n2685_lo <= 1'b0;
    n2688_lo <= 1'b0;
    n2691_lo <= 1'b0;
    n2700_lo <= 1'b0;
    n2703_lo <= 1'b0;
    n2736_lo <= 1'b0;
    n2739_lo <= 1'b0;
    n2748_lo <= 1'b0;
    n2760_lo <= 1'b0;
    n2772_lo <= 1'b0;
    n2775_lo <= 1'b0;
    n2784_lo <= 1'b0;
    n2787_lo <= 1'b0;
    n2790_lo <= 1'b0;
    n2793_lo <= 1'b0;
    n2796_lo <= 1'b0;
    n2799_lo <= 1'b0;
    n2802_lo <= 1'b0;
    n2805_lo <= 1'b0;
    n2808_lo <= 1'b0;
    n2820_lo <= 1'b0;
    n2823_lo <= 1'b0;
    n2826_lo <= 1'b0;
    n2832_lo <= 1'b0;
    n2835_lo <= 1'b0;
    n2838_lo <= 1'b0;
    n2841_lo <= 1'b0;
    n2844_lo <= 1'b0;
    n2856_lo <= 1'b0;
    n2859_lo <= 1'b0;
    n2862_lo <= 1'b0;
    n2865_lo <= 1'b0;
    n2868_lo <= 1'b0;
    n2871_lo <= 1'b0;
    n2874_lo <= 1'b0;
    n2877_lo <= 1'b0;
    n2880_lo <= 1'b0;
    n2883_lo <= 1'b0;
    n2886_lo <= 1'b0;
    n2889_lo <= 1'b0;
    n2892_lo <= 1'b0;
    n2895_lo <= 1'b0;
    n2898_lo <= 1'b0;
    n2901_lo <= 1'b0;
    n2904_lo <= 1'b0;
    n2907_lo <= 1'b0;
    n2916_lo <= 1'b0;
    n2928_lo <= 1'b0;
    n2940_lo <= 1'b0;
    n2952_lo <= 1'b0;
    n2955_lo <= 1'b0;
    n2964_lo <= 1'b0;
    n2976_lo <= 1'b0;
    n2988_lo <= 1'b0;
    n2991_lo <= 1'b0;
    n3000_lo <= 1'b0;
    n3003_lo <= 1'b0;
    n3012_lo <= 1'b0;
    n3015_lo <= 1'b0;
    n3024_lo <= 1'b0;
    n3027_lo <= 1'b0;
    n3036_lo <= 1'b0;
    n3039_lo <= 1'b0;
    n3048_lo <= 1'b0;
    n3051_lo <= 1'b0;
    n3054_lo <= 1'b0;
    n3057_lo <= 1'b0;
    n3060_lo <= 1'b0;
    n3072_lo <= 1'b0;
    n3081_lo <= 1'b0;
    n3084_lo <= 1'b0;
    n3087_lo <= 1'b0;
    n3093_lo <= 1'b0;
    n3096_lo <= 1'b0;
    n3105_lo <= 1'b0;
    n3108_lo <= 1'b0;
    n3117_lo <= 1'b0;
    n3120_lo <= 1'b0;
    n3123_lo <= 1'b0;
    n3126_lo <= 1'b0;
    n3129_lo <= 1'b0;
    n3132_lo <= 1'b0;
    n3135_lo <= 1'b0;
    n3138_lo <= 1'b0;
    n3141_lo <= 1'b0;
    n3168_lo <= 1'b0;
    n3171_lo <= 1'b0;
    n3174_lo <= 1'b0;
    n3177_lo <= 1'b0;
    n3180_lo <= 1'b0;
    n3183_lo <= 1'b0;
    n3192_lo <= 1'b0;
    n3195_lo <= 1'b0;
    n3204_lo <= 1'b0;
    n3207_lo <= 1'b0;
    n3216_lo <= 1'b0;
    n3219_lo <= 1'b0;
    n3228_lo <= 1'b0;
    n3231_lo <= 1'b0;
    n3240_lo <= 1'b0;
    n3243_lo <= 1'b0;
    n3252_lo <= 1'b0;
    n3255_lo <= 1'b0;
    n3258_lo <= 1'b0;
    n3264_lo <= 1'b0;
    n3267_lo <= 1'b0;
    n3270_lo <= 1'b0;
    n3276_lo <= 1'b0;
    n3279_lo <= 1'b0;
    n3282_lo <= 1'b0;
    n3288_lo <= 1'b0;
    n3291_lo <= 1'b0;
    n3294_lo <= 1'b0;
    n4537_o2 <= 1'b0;
    n4538_o2 <= 1'b0;
    n4710_o2 <= 1'b0;
    n4711_o2 <= 1'b0;
    n1211_inv <= 1'b0;
    n1214_inv <= 1'b0;
    n1217_inv <= 1'b0;
    n1220_inv <= 1'b0;
    n4927_o2 <= 1'b0;
    n4928_o2 <= 1'b0;
    n1229_inv <= 1'b0;
    n1232_inv <= 1'b0;
    n1235_inv <= 1'b0;
    n5178_o2 <= 1'b0;
    n5179_o2 <= 1'b0;
    n5477_o2 <= 1'b0;
    n5478_o2 <= 1'b0;
    n5479_o2 <= 1'b0;
    n5222_o2 <= 1'b0;
    n5223_o2 <= 1'b0;
    n5553_o2 <= 1'b0;
    n5554_o2 <= 1'b0;
    G491_o2 <= 1'b0;
    n2922_lo_buf_o2 <= 1'b0;
    n2946_lo_buf_o2 <= 1'b0;
    n2970_lo_buf_o2 <= 1'b0;
    n2982_lo_buf_o2 <= 1'b0;
    n3066_lo_buf_o2 <= 1'b0;
    n3078_lo_buf_o2 <= 1'b0;
    n3102_lo_buf_o2 <= 1'b0;
    n3114_lo_buf_o2 <= 1'b0;
    G1321_o2 <= 1'b0;
    G1033_o2 <= 1'b0;
    G1030_o2 <= 1'b0;
    G1072_o2 <= 1'b0;
    n1304_inv <= 1'b0;
    n1307_inv <= 1'b0;
    n2958_lo_buf_o2 <= 1'b0;
    n2994_lo_buf_o2 <= 1'b0;
    n3006_lo_buf_o2 <= 1'b0;
    n3030_lo_buf_o2 <= 1'b0;
    n3042_lo_buf_o2 <= 1'b0;
    n3090_lo_buf_o2 <= 1'b0;
    n1328_inv <= 1'b0;
    n1331_inv <= 1'b0;
    n1334_inv <= 1'b0;
    n1337_inv <= 1'b0;
    n1340_inv <= 1'b0;
    n1343_inv <= 1'b0;
    n1346_inv <= 1'b0;
    n1349_inv <= 1'b0;
    G1036_o2 <= 1'b0;
    G1062_o2 <= 1'b0;
    G1067_o2 <= 1'b0;
    G1014_o2 <= 1'b0;
    n1364_inv <= 1'b0;
    n1367_inv <= 1'b0;
    n3018_lo_buf_o2 <= 1'b0;
    G766_o2 <= 1'b0;
    n1376_inv <= 1'b0;
    n1379_inv <= 1'b0;
    n1382_inv <= 1'b0;
    n1385_inv <= 1'b0;
    n1388_inv <= 1'b0;
    n1391_inv <= 1'b0;
    G1017_o2 <= 1'b0;
    G1008_o2 <= 1'b0;
    n1400_inv <= 1'b0;
    n1403_inv <= 1'b0;
    n2910_lo_buf_o2 <= 1'b0;
    n1409_inv <= 1'b0;
    G2138_o2 <= 1'b0;
    G2147_o2 <= 1'b0;
    n1418_inv <= 1'b0;
    G1137_o2 <= 1'b0;
    G1329_o2 <= 1'b0;
    G374_o2 <= 1'b0;
    G386_o2 <= 1'b0;
    G663_o2 <= 1'b0;
    G674_o2 <= 1'b0;
    G578_o2 <= 1'b0;
    G575_o2 <= 1'b0;
    G2505_o2 <= 1'b0;
    n1448_inv <= 1'b0;
    G987_o2 <= 1'b0;
    G984_o2 <= 1'b0;
    G1862_o2 <= 1'b0;
    G1859_o2 <= 1'b0;
    G1260_o2 <= 1'b0;
    G1865_o2 <= 1'b0;
    G2073_o2 <= 1'b0;
    G1402_o2 <= 1'b0;
    G2048_o2 <= 1'b0;
    G2276_o2 <= 1'b0;
    n1481_inv <= 1'b0;
    G2141_o2 <= 1'b0;
    G2008_o2 <= 1'b0;
    G2011_o2 <= 1'b0;
    G2150_o2 <= 1'b0;
    G2026_o2 <= 1'b0;
    G2029_o2 <= 1'b0;
    G2023_o2 <= 1'b0;
    G2041_o2 <= 1'b0;
    G2017_o2 <= 1'b0;
    G2020_o2 <= 1'b0;
    G2035_o2 <= 1'b0;
    G2038_o2 <= 1'b0;
    G2228_o2 <= 1'b0;
    G2231_o2 <= 1'b0;
    G2234_o2 <= 1'b0;
    G2237_o2 <= 1'b0;
    G1904_o2 <= 1'b0;
    G1907_o2 <= 1'b0;
    G1928_o2 <= 1'b0;
    G1931_o2 <= 1'b0;
    G1893_o2 <= 1'b0;
    G1896_o2 <= 1'b0;
    G1899_o2 <= 1'b0;
    G1937_o2 <= 1'b0;
    G1940_o2 <= 1'b0;
    G1943_o2 <= 1'b0;
    G1336_o2 <= 1'b0;
    G1996_o2 <= 1'b0;
    G1999_o2 <= 1'b0;
    G2002_o2 <= 1'b0;
    G2005_o2 <= 1'b0;
    G2014_o2 <= 1'b0;
    G2032_o2 <= 1'b0;
    G1076_o2 <= 1'b0;
    G1002_o2 <= 1'b0;
    G998_o2 <= 1'b0;
    G1890_o2 <= 1'b0;
    G1934_o2 <= 1'b0;
    G1044_o2 <= 1'b0;
    G1039_o2 <= 1'b0;
    n1770_lo_buf_o2 <= 1'b0;
    G342_o2 <= 1'b0;
    G354_o2 <= 1'b0;
    G1193_o2 <= 1'b0;
    n3234_lo_buf_o2 <= 1'b0;
    n3246_lo_buf_o2 <= 1'b0;
    G783_o2 <= 1'b0;
    G786_o2 <= 1'b0;
    G792_o2 <= 1'b0;
    G795_o2 <= 1'b0;
    G815_o2 <= 1'b0;
    G818_o2 <= 1'b0;
    G824_o2 <= 1'b0;
    G827_o2 <= 1'b0;
    G789_o2 <= 1'b0;
    G798_o2 <= 1'b0;
    G801_o2 <= 1'b0;
    G807_o2 <= 1'b0;
    G812_o2 <= 1'b0;
    G821_o2 <= 1'b0;
    G804_o2 <= 1'b0;
    G780_o2 <= 1'b0;
    G1231_o2 <= 1'b0;
    G1572_o2 <= 1'b0;
    G1377_o2 <= 1'b0;
    G1253_o2 <= 1'b0;
    G1359_o2 <= 1'b0;
    G1258_o2 <= 1'b0;
    G1367_o2 <= 1'b0;
    G1358_o2 <= 1'b0;
    G1366_o2 <= 1'b0;
    G2057_o2 <= 1'b0;
    G2117_o2 <= 1'b0;
    G2118_o2 <= 1'b0;
    G1254_o2 <= 1'b0;
    G1259_o2 <= 1'b0;
    G2058_o2 <= 1'b0;
    G405_o2 <= 1'b0;
    G417_o2 <= 1'b0;
    G1269_o2 <= 1'b0;
    G1275_o2 <= 1'b0;
    G1287_o2 <= 1'b0;
    G1266_o2 <= 1'b0;
    G1272_o2 <= 1'b0;
    G1278_o2 <= 1'b0;
    G1281_o2 <= 1'b0;
    G1284_o2 <= 1'b0;
    G1290_o2 <= 1'b0;
    G1293_o2 <= 1'b0;
    G1299_o2 <= 1'b0;
    G1305_o2 <= 1'b0;
    G1296_o2 <= 1'b0;
    G1302_o2 <= 1'b0;
    G1308_o2 <= 1'b0;
    G1311_o2 <= 1'b0;
    G811_o2 <= 1'b0;
    G810_o2 <= 1'b0;
    G1728_o2 <= 1'b0;
    G2512_o2 <= 1'b0;
    G1114_o2 <= 1'b0;
    G1113_o2 <= 1'b0;
    G1992_o2 <= 1'b0;
    G1991_o2 <= 1'b0;
    G1426_o2 <= 1'b0;
    G1966_o2 <= 1'b0;
    G2211_o2 <= 1'b0;
    G1509_o2 <= 1'b0;
    G2153_o2 <= 1'b0;
    G2329_o2 <= 1'b0;
    G1540_o2 <= 1'b0;
    G2167_o2 <= 1'b0;
    G2191_o2 <= 1'b0;
    G1234_o2 <= 1'b0;
    G1132_o2 <= 1'b0;
    G1129_o2 <= 1'b0;
    G2088_o2 <= 1'b0;
    G2106_o2 <= 1'b0;
    G1314_o2 <= 1'b0;
    G636_o2 <= 1'b0;
    G647_o2 <= 1'b0;
    n3186_lo_buf_o2 <= 1'b0;
    n3198_lo_buf_o2 <= 1'b0;
    n3210_lo_buf_o2 <= 1'b0;
    n3222_lo_buf_o2 <= 1'b0;
    G1225_o2 <= 1'b0;
    G1342_o2 <= 1'b0;
    G1222_o2 <= 1'b0;
    G1228_o2 <= 1'b0;
    G1348_o2 <= 1'b0;
    G1345_o2 <= 1'b0;
    G1351_o2 <= 1'b0;
    G2242_o2 <= 1'b0;
    G2260_o2 <= 1'b0;
    G1374_o2 <= 1'b0;
    G1537_o2 <= 1'b0;
    G301_o2 <= 1'b0;
    G313_o2 <= 1'b0;
    G2365_o2 <= 1'b0;
    G2255_o2 <= 1'b0;
    G2253_o2 <= 1'b0;
    G2395_o2 <= 1'b0;
    G2272_o2 <= 1'b0;
    G2270_o2 <= 1'b0;
    G2245_o2 <= 1'b0;
    G2262_o2 <= 1'b0;
    G2249_o2 <= 1'b0;
    G2247_o2 <= 1'b0;
    G2266_o2 <= 1'b0;
    G2264_o2 <= 1'b0;
    G2403_o2 <= 1'b0;
    G2401_o2 <= 1'b0;
    G2410_o2 <= 1'b0;
    G2408_o2 <= 1'b0;
    G2306_o2 <= 1'b0;
    G2305_o2 <= 1'b0;
    G2314_o2 <= 1'b0;
    G2313_o2 <= 1'b0;
    G2303_o2 <= 1'b0;
    G2302_o2 <= 1'b0;
    G2301_o2 <= 1'b0;
    G2311_o2 <= 1'b0;
    G2310_o2 <= 1'b0;
    G2309_o2 <= 1'b0;
    G2404_o2 <= 1'b0;
    G2411_o2 <= 1'b0;
    G2420_o2 <= 1'b0;
    G2419_o2 <= 1'b0;
    G2433_o2 <= 1'b0;
    G2432_o2 <= 1'b0;
    G402_o2 <= 1'b0;
    G403_o2 <= 1'b0;
    G1053_o2 <= 1'b0;
    G1049_o2 <= 1'b0;
    n2003_inv <= 1'b0;
    G1364_o2 <= 1'b0;
    G1079_o2 <= 1'b0;
    G1478_o2 <= 1'b0;
    G707_o2 <= 1'b0;
    G718_o2 <= 1'b0;
    G2417_o2 <= 1'b0;
    G2414_o2 <= 1'b0;
    G2431_o2 <= 1'b0;
    G2428_o2 <= 1'b0;
    G1653_o2 <= 1'b0;
    G2213_o2 <= 1'b0;
    G2221_o2 <= 1'b0;
    G2250_o2 <= 1'b0;
    G2267_o2 <= 1'b0;
    G1365_o2 <= 1'b0;
    G1368_o2 <= 1'b0;
    G1371_o2 <= 1'b0;
    G2218_o2 <= 1'b0;
    G2225_o2 <= 1'b0;
    n1503_lo_buf_o2 <= 1'b0;
    n1863_lo_buf_o2 <= 1'b0;
    n1887_lo_buf_o2 <= 1'b0;
    n1983_lo_buf_o2 <= 1'b0;
    n2007_lo_buf_o2 <= 1'b0;
    n2115_lo_buf_o2 <= 1'b0;
    n2139_lo_buf_o2 <= 1'b0;
    n2247_lo_buf_o2 <= 1'b0;
    n2271_lo_buf_o2 <= 1'b0;
    n2919_lo_buf_o2 <= 1'b0;
    n2943_lo_buf_o2 <= 1'b0;
    n2967_lo_buf_o2 <= 1'b0;
    n2979_lo_buf_o2 <= 1'b0;
    n3063_lo_buf_o2 <= 1'b0;
    n3075_lo_buf_o2 <= 1'b0;
    n3099_lo_buf_o2 <= 1'b0;
    n3111_lo_buf_o2 <= 1'b0;
    G878_o2 <= 1'b0;
    G875_o2 <= 1'b0;
    G661_o2 <= 1'b0;
    G660_o2 <= 1'b0;
    G879_o2 <= 1'b0;
    G876_o2 <= 1'b0;
    G1320_o2 <= 1'b0;
    G941_o2 <= 1'b0;
    G732_o2 <= 1'b0;
    G942_o2 <= 1'b0;
    G1493_o2 <= 1'b0;
    G1498_o2 <= 1'b0;
    G877_o2 <= 1'b0;
    G874_o2 <= 1'b0;
    n1806_lo_buf_o2 <= 1'b0;
    n1878_lo_buf_o2 <= 1'b0;
    n1938_lo_buf_o2 <= 1'b0;
    n1998_lo_buf_o2 <= 1'b0;
    n2058_lo_buf_o2 <= 1'b0;
    n2130_lo_buf_o2 <= 1'b0;
    n2190_lo_buf_o2 <= 1'b0;
    n2262_lo_buf_o2 <= 1'b0;
    n2310_lo_buf_o2 <= 1'b0;
    n2406_lo_buf_o2 <= 1'b0;
    n2430_lo_buf_o2 <= 1'b0;
    n2526_lo_buf_o2 <= 1'b0;
    n2550_lo_buf_o2 <= 1'b0;
    n2646_lo_buf_o2 <= 1'b0;
    n2670_lo_buf_o2 <= 1'b0;
    n2766_lo_buf_o2 <= 1'b0;
    G603_o2 <= 1'b0;
    G614_o2 <= 1'b0;
    G1026_o2 <= 1'b0;
    G1021_o2 <= 1'b0;
    G940_o2 <= 1'b0;
    G1636_o2 <= 1'b0;
    G1684_o2 <= 1'b0;
    n2352_lo_buf_o2 <= 1'b0;
    n2364_lo_buf_o2 <= 1'b0;
    n2472_lo_buf_o2 <= 1'b0;
    n2484_lo_buf_o2 <= 1'b0;
    n2592_lo_buf_o2 <= 1'b0;
    n2604_lo_buf_o2 <= 1'b0;
    n2712_lo_buf_o2 <= 1'b0;
    n2724_lo_buf_o2 <= 1'b0;
    n3150_lo_buf_o2 <= 1'b0;
    n3162_lo_buf_o2 <= 1'b0;
  end
endmodule


