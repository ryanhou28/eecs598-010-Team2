
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  G42,
  G43,
  G44,
  G45,
  G46,
  G47,
  G48,
  G49,
  G50,
  G51,
  G52,
  G53,
  G54,
  G55,
  G56,
  G57,
  G58,
  G59,
  G60,
  G61,
  G62,
  G63,
  G64,
  G65,
  G66,
  G67,
  G68,
  G69,
  G70,
  G71,
  G72,
  G73,
  G74,
  G75,
  G76,
  G77,
  G78,
  G79,
  G80,
  G81,
  G82,
  G83,
  G84,
  G85,
  G86,
  G87,
  G88,
  G89,
  G90,
  G91,
  G92,
  G93,
  G94,
  G95,
  G96,
  G97,
  G98,
  G99,
  G100,
  G101,
  G102,
  G103,
  G104,
  G105,
  G106,
  G107,
  G108,
  G109,
  G110,
  G111,
  G112,
  G113,
  G114,
  G115,
  G116,
  G117,
  G118,
  G119,
  G120,
  G121,
  G122,
  G123,
  G124,
  G125,
  G126,
  G127,
  G128,
  G129,
  G130,
  G131,
  G132,
  G133,
  G134,
  G135,
  G136,
  G137,
  G138,
  G139,
  G140,
  G141,
  G142,
  G143,
  G144,
  G145,
  G146,
  G147,
  G148,
  G149,
  G150,
  G151,
  G152,
  G153,
  G154,
  G155,
  G156,
  G157,
  G158,
  G159,
  G160,
  G161,
  G162,
  G163,
  G164,
  G165,
  G166,
  G167,
  G168,
  G169,
  G170,
  G171,
  G172,
  G173,
  G174,
  G175,
  G176,
  G177,
  G178,
  n2610_lo,
  n2613_lo,
  n2616_lo,
  n2619_lo,
  n2622_lo,
  n2625_lo,
  n2628_lo,
  n2631_lo,
  n2634_lo,
  n2637_lo,
  n2640_lo,
  n2643_lo,
  n2646_lo,
  n2649_lo,
  n2652_lo,
  n2655_lo,
  n2658_lo,
  n2661_lo,
  n2664_lo,
  n2667_lo,
  n2670_lo,
  n2673_lo,
  n2676_lo,
  n2679_lo,
  n2682_lo,
  n2685_lo,
  n2688_lo,
  n2691_lo,
  n2694_lo,
  n2697_lo,
  n2700_lo,
  n2703_lo,
  n2706_lo,
  n2709_lo,
  n2712_lo,
  n2715_lo,
  n2718_lo,
  n2721_lo,
  n2724_lo,
  n2727_lo,
  n2730_lo,
  n2733_lo,
  n2736_lo,
  n2739_lo,
  n2742_lo,
  n2745_lo,
  n2748_lo,
  n2751_lo,
  n2754_lo,
  n2757_lo,
  n2760_lo,
  n2763_lo,
  n2766_lo,
  n2769_lo,
  n2772_lo,
  n2775_lo,
  n2778_lo,
  n2781_lo,
  n2784_lo,
  n2787_lo,
  n2790_lo,
  n2793_lo,
  n2796_lo,
  n2799_lo,
  n2802_lo,
  n2805_lo,
  n2808_lo,
  n2811_lo,
  n2814_lo,
  n2817_lo,
  n2820_lo,
  n2823_lo,
  n2826_lo,
  n2829_lo,
  n2832_lo,
  n2835_lo,
  n2838_lo,
  n2841_lo,
  n2844_lo,
  n2847_lo,
  n2850_lo,
  n2853_lo,
  n2856_lo,
  n2859_lo,
  n2862_lo,
  n2865_lo,
  n2868_lo,
  n2871_lo,
  n2874_lo,
  n2877_lo,
  n2880_lo,
  n2883_lo,
  n2886_lo,
  n2889_lo,
  n2892_lo,
  n2895_lo,
  n2898_lo,
  n2901_lo,
  n2904_lo,
  n2907_lo,
  n2910_lo,
  n2913_lo,
  n2916_lo,
  n2919_lo,
  n2922_lo,
  n2925_lo,
  n2928_lo,
  n2931_lo,
  n2934_lo,
  n2937_lo,
  n2940_lo,
  n2943_lo,
  n2946_lo,
  n2949_lo,
  n2952_lo,
  n2955_lo,
  n2958_lo,
  n2961_lo,
  n2964_lo,
  n2967_lo,
  n2970_lo,
  n2973_lo,
  n2976_lo,
  n2979_lo,
  n2982_lo,
  n2985_lo,
  n2988_lo,
  n2991_lo,
  n2994_lo,
  n2997_lo,
  n3000_lo,
  n3003_lo,
  n3006_lo,
  n3009_lo,
  n3012_lo,
  n3015_lo,
  n3018_lo,
  n3021_lo,
  n3024_lo,
  n3027_lo,
  n3030_lo,
  n3033_lo,
  n3036_lo,
  n3039_lo,
  n3042_lo,
  n3045_lo,
  n3048_lo,
  n3051_lo,
  n3054_lo,
  n3057_lo,
  n3060_lo,
  n3063_lo,
  n3066_lo,
  n3069_lo,
  n3072_lo,
  n3075_lo,
  n3078_lo,
  n3081_lo,
  n3084_lo,
  n3087_lo,
  n3090_lo,
  n3093_lo,
  n3096_lo,
  n3099_lo,
  n3102_lo,
  n3105_lo,
  n3108_lo,
  n3111_lo,
  n3114_lo,
  n3117_lo,
  n3120_lo,
  n3123_lo,
  n3126_lo,
  n3129_lo,
  n3132_lo,
  n3135_lo,
  n3138_lo,
  n3141_lo,
  n3144_lo,
  n3147_lo,
  n3150_lo,
  n3153_lo,
  n3156_lo,
  n3159_lo,
  n3162_lo,
  n3165_lo,
  n3168_lo,
  n3171_lo,
  n3174_lo,
  n3177_lo,
  n3180_lo,
  n3183_lo,
  n3186_lo,
  n3189_lo,
  n3192_lo,
  n3195_lo,
  n3198_lo,
  n3201_lo,
  n3204_lo,
  n3207_lo,
  n3210_lo,
  n3213_lo,
  n3216_lo,
  n3219_lo,
  n3222_lo,
  n3225_lo,
  n3228_lo,
  n3231_lo,
  n3234_lo,
  n3237_lo,
  n3240_lo,
  n3243_lo,
  n3246_lo,
  n3249_lo,
  n3252_lo,
  n3255_lo,
  n3258_lo,
  n3261_lo,
  n3264_lo,
  n3267_lo,
  n3270_lo,
  n3273_lo,
  n3276_lo,
  n3279_lo,
  n3282_lo,
  n3285_lo,
  n3288_lo,
  n3291_lo,
  n3294_lo,
  n3297_lo,
  n3300_lo,
  n3303_lo,
  n3306_lo,
  n3309_lo,
  n3312_lo,
  n3315_lo,
  n3318_lo,
  n3321_lo,
  n3324_lo,
  n3327_lo,
  n3330_lo,
  n3333_lo,
  n3336_lo,
  n3339_lo,
  n3342_lo,
  n3345_lo,
  n3348_lo,
  n3351_lo,
  n3354_lo,
  n3357_lo,
  n3360_lo,
  n3363_lo,
  n3366_lo,
  n3369_lo,
  n3372_lo,
  n3375_lo,
  n3378_lo,
  n3381_lo,
  n3384_lo,
  n3387_lo,
  n3390_lo,
  n3393_lo,
  n3396_lo,
  n3399_lo,
  n3402_lo,
  n3405_lo,
  n3408_lo,
  n3411_lo,
  n3414_lo,
  n3417_lo,
  n3420_lo,
  n3423_lo,
  n3426_lo,
  n3429_lo,
  n3432_lo,
  n3435_lo,
  n3438_lo,
  n3441_lo,
  n3444_lo,
  n3447_lo,
  n3450_lo,
  n3453_lo,
  n3456_lo,
  n3459_lo,
  n3462_lo,
  n3465_lo,
  n3468_lo,
  n3471_lo,
  n3474_lo,
  n3477_lo,
  n3480_lo,
  n3483_lo,
  n3486_lo,
  n3489_lo,
  n3492_lo,
  n3495_lo,
  n3498_lo,
  n3501_lo,
  n3504_lo,
  n3507_lo,
  n3510_lo,
  n3513_lo,
  n3516_lo,
  n3519_lo,
  n3522_lo,
  n3525_lo,
  n3528_lo,
  n3531_lo,
  n3534_lo,
  n3537_lo,
  n3540_lo,
  n3543_lo,
  n3546_lo,
  n3549_lo,
  n3552_lo,
  n3555_lo,
  n3558_lo,
  n3561_lo,
  n3564_lo,
  n3567_lo,
  n3570_lo,
  n3573_lo,
  n3576_lo,
  n3579_lo,
  n3582_lo,
  n3585_lo,
  n3588_lo,
  n3591_lo,
  n3594_lo,
  n3597_lo,
  n3600_lo,
  n3603_lo,
  n3606_lo,
  n3609_lo,
  n3612_lo,
  n3615_lo,
  n3618_lo,
  n3621_lo,
  n3624_lo,
  n3627_lo,
  n3630_lo,
  n3633_lo,
  n3636_lo,
  n3639_lo,
  n3642_lo,
  n3645_lo,
  n3648_lo,
  n3651_lo,
  n3654_lo,
  n3657_lo,
  n3666_lo,
  n3669_lo,
  n3678_lo,
  n3687_lo,
  n3690_lo,
  n3702_lo,
  n3711_lo,
  n3714_lo,
  n3726_lo,
  n3735_lo,
  n3738_lo,
  n3750_lo,
  n3753_lo,
  n3759_lo,
  n3762_lo,
  n3765_lo,
  n3774_lo,
  n3777_lo,
  n3786_lo,
  n3789_lo,
  n3792_lo,
  n3795_lo,
  n3798_lo,
  n3801_lo,
  n3810_lo,
  n3813_lo,
  n3822_lo,
  n3825_lo,
  n3834_lo,
  n3843_lo,
  n3846_lo,
  n3867_lo,
  n3891_lo,
  n3915_lo,
  n3930_lo,
  n3933_lo,
  n3936_lo,
  n3942_lo,
  n3945_lo,
  n3948_lo,
  n3954_lo,
  n3957_lo,
  n3963_lo,
  n3966_lo,
  n3969_lo,
  n3975_lo,
  n3978_lo,
  n3987_lo,
  n3990_lo,
  n4002_lo,
  n4011_lo,
  n4014_lo,
  n4026_lo,
  n4035_lo,
  n4038_lo,
  n4050_lo,
  n4053_lo,
  n4059_lo,
  n4062_lo,
  n4065_lo,
  n4098_lo,
  n4107_lo,
  n4119_lo,
  n4131_lo,
  n4143_lo,
  n4155_lo,
  n4167_lo,
  n4179_lo,
  n4182_lo,
  n4185_lo,
  n4188_lo,
  n4194_lo,
  n4197_lo,
  n4200_lo,
  n4206_lo,
  n4209_lo,
  n4212_lo,
  n4215_lo,
  n4227_lo,
  n4230_lo,
  n4233_lo,
  n4236_lo,
  n4239_lo,
  n4242_lo,
  n4251_lo,
  n4263_lo,
  n4275_lo,
  n4278_lo,
  n4287_lo,
  n4290_lo,
  n4293_lo,
  n4299_lo,
  n4302_lo,
  n4305_lo,
  n4311_lo,
  n4314_lo,
  n4323_lo,
  n4326_lo,
  n4335_lo,
  n4338_lo,
  n4347_lo,
  n4350_lo,
  n4359_lo,
  n4362_lo,
  n4365_lo,
  n4371_lo,
  n4374_lo,
  n4383_lo,
  n4395_lo,
  n4407_lo,
  n4410_lo,
  n4413_lo,
  n4416_lo,
  n4419_lo,
  n4422_lo,
  n4425_lo,
  n4428_lo,
  n4431_lo,
  n4434_lo,
  n4437_lo,
  n4440_lo,
  n4443_lo,
  n4446_lo,
  n4449_lo,
  n4452_lo,
  n4455_lo,
  n4458_lo,
  n4461_lo,
  n4464_lo,
  n4467_lo,
  n4470_lo,
  n4473_lo,
  n4476_lo,
  n4479_lo,
  n4482_lo,
  n4485_lo,
  n4488_lo,
  n4494_lo,
  n4497_lo,
  n4500_lo,
  n4503_lo,
  n4506_lo,
  n4509_lo,
  n4512_lo,
  n4515_lo,
  n4518_lo,
  n4521_lo,
  n4524_lo,
  n4527_lo,
  n4530_lo,
  n4533_lo,
  n4536_lo,
  n4539_lo,
  n4542_lo,
  n4545_lo,
  n4548_lo,
  n4554_lo,
  n4557_lo,
  n4560_lo,
  n4563_lo,
  n4566_lo,
  n4569_lo,
  n4572_lo,
  n4575_lo,
  n4578_lo,
  n4581_lo,
  n4584_lo,
  n4587_lo,
  n4590_lo,
  n4593_lo,
  n4596_lo,
  n4599_lo,
  n4602_lo,
  n4605_lo,
  n4608_lo,
  n4611_lo,
  n4614_lo,
  n4617_lo,
  n4620_lo,
  n4623_lo,
  n4626_lo,
  n4629_lo,
  n4632_lo,
  n4635_lo,
  n4638_lo,
  n4641_lo,
  n4644_lo,
  n4647_lo,
  n4650_lo,
  n4653_lo,
  n4656_lo,
  n4659_lo,
  n4662_lo,
  n4665_lo,
  n4668_lo,
  n4671_lo,
  n4674_lo,
  n4677_lo,
  n4680_lo,
  n4683_lo,
  n4686_lo,
  n4689_lo,
  n4692_lo,
  n4695_lo,
  n4698_lo,
  n4701_lo,
  n4704_lo,
  n4707_lo,
  n4710_lo,
  n4713_lo,
  n4716_lo,
  n4719_lo,
  n4722_lo,
  n4725_lo,
  n4728_lo,
  n4731_lo,
  n4734_lo,
  n4737_lo,
  n4740_lo,
  n4743_lo,
  n6382_o2,
  n6383_o2,
  n6419_o2,
  n6420_o2,
  n6435_o2,
  n6436_o2,
  n6448_o2,
  n6449_o2,
  n6613_o2,
  n6614_o2,
  n6641_o2,
  n6658_o2,
  n6757_o2,
  n6756_o2,
  n7116_o2,
  n7156_o2,
  n6549_o2,
  n6550_o2,
  n7357_o2,
  n7358_o2,
  n7359_o2,
  n7360_o2,
  n6621_o2,
  n6623_o2,
  n6625_o2,
  n6626_o2,
  n6627_o2,
  n6628_o2,
  n6629_o2,
  n6630_o2,
  n6669_o2,
  n7449_o2,
  n7450_o2,
  n7451_o2,
  n7452_o2,
  n6682_o2,
  n6683_o2,
  n6684_o2,
  n6685_o2,
  n7463_o2,
  n6686_o2,
  n6687_o2,
  n6688_o2,
  n6689_o2,
  n6772_o2,
  n6773_o2,
  n6774_o2,
  n6775_o2,
  G3467_o2,
  G2810_o2,
  n6833_o2,
  n6945_o2,
  n6947_o2,
  n6949_o2,
  n6951_o2,
  n6888_o2,
  n6889_o2,
  n6936_o2,
  n6954_o2,
  n6955_o2,
  n6956_o2,
  n6957_o2,
  n6958_o2,
  n6982_o2,
  n6984_o2,
  n6974_o2,
  n6975_o2,
  n6999_o2,
  n7015_o2,
  n7016_o2,
  n7017_o2,
  n7018_o2,
  n7005_o2,
  n7019_o2,
  n7022_o2,
  n7023_o2,
  n7132_o2,
  n7133_o2,
  n7135_o2,
  n7136_o2,
  n7175_o2,
  n7155_o2,
  G3060_o2,
  n7383_o2,
  G3802_o2,
  G3859_o2,
  n7355_o2,
  n7356_o2,
  G4054_o2,
  G4068_o2,
  n7384_o2,
  n7387_o2,
  n7388_o2,
  n7389_o2,
  n7386_o2,
  n7453_o2,
  n7431_o2,
  n7432_o2,
  n7433_o2,
  n7430_o2,
  n7485_o2,
  n7486_o2,
  G2508_o2,
  G2486_o2,
  n2326_inv,
  n2329_inv,
  n3756_lo_buf_o2,
  n4056_lo_buf_o2,
  G3474_o2,
  n2341_inv,
  n7396_o2,
  n7398_o2,
  n7400_o2,
  n7401_o2,
  n7402_o2,
  n7403_o2,
  n7404_o2,
  n7405_o2,
  G2711_o2,
  n2371_inv,
  n7490_o2,
  n7527_o2,
  n7528_o2,
  n7529_o2,
  n7530_o2,
  n7523_o2,
  n7524_o2,
  n7525_o2,
  n7526_o2,
  n4296_lo_buf_o2,
  n4368_lo_buf_o2,
  G2466_o2,
  G2404_o2,
  n7534_o2,
  n7535_o2,
  n7536_o2,
  n7533_o2,
  G1060_o2,
  G963_o2,
  G2448_o2,
  G2685_o2,
  G2679_o2,
  G2774_o2,
  G2780_o2,
  G2759_o2,
  G2737_o2,
  G2850_o2,
  G3393_o2,
  G3404_o2,
  G3559_o2,
  G2744_o2,
  n3708_lo_buf_o2,
  n3840_lo_buf_o2,
  n4008_lo_buf_o2,
  n4104_lo_buf_o2,
  G1821_o2,
  G1734_o2,
  G3517_o2,
  G3533_o2,
  G3629_o2,
  G3645_o2,
  n2497_inv,
  G2731_o2,
  G2844_o2,
  n3732_lo_buf_o2,
  n4032_lo_buf_o2,
  G3552_o2,
  G2271_o2,
  n4248_lo_buf_o2,
  n4332_lo_buf_o2,
  n4344_lo_buf_o2,
  n4380_lo_buf_o2,
  G2398_o2,
  G2480_o2,
  G2418_o2,
  G1455_o2,
  G1449_o2,
  G1452_o2,
  G1425_o2,
  G1428_o2,
  G1419_o2,
  G1422_o2,
  n4308_lo_buf_o2,
  G2675_o2,
  G3035_o2,
  G3026_o2,
  G3029_o2,
  G3032_o2,
  G2999_o2,
  G3002_o2,
  G2770_o2,
  G3008_o2,
  G2073_o2,
  G2752_o2,
  G3005_o2,
  G5108_o2,
  G5135_o2,
  G5111_o2,
  G5138_o2,
  G3415_o2,
  G3386_o2,
  G3570_o2,
  G2430_o2,
  G3495_o2,
  G3621_o2,
  n4284_lo_buf_o2,
  n4356_lo_buf_o2,
  G2472_o2,
  G2410_o2,
  n3960_lo_buf_o2,
  n3972_lo_buf_o2,
  n2647_inv,
  n2650_inv,
  n3684_lo_buf_o2,
  n4080_lo_buf_o2,
  n4092_lo_buf_o2,
  n2662_inv,
  n2665_inv,
  G1147_o2,
  G2705_o2,
  G2693_o2,
  G2696_o2,
  G2700_o2,
  G2915_o2,
  G2966_o2,
  G2540_o2,
  G2788_o2,
  G2792_o2,
  G2797_o2,
  G2804_o2,
  G1038_o2,
  G1044_o2,
  G1090_o2,
  G1096_o2,
  G1029_o2,
  G3942_o2,
  G3954_o2,
  G4011_o2,
  G4017_o2,
  G1141_o2,
  G1081_o2,
  G2146_o2,
  G2145_o2,
  G2144_o2,
  G2143_o2,
  G2142_o2,
  G2141_o2,
  G2140_o2,
  G2139_o2,
  G3769_o2,
  G3773_o2,
  G3768_o2,
  G4101_o2,
  G3161_o2,
  G4143_o2,
  G3828_o2,
  G3831_o2,
  G3334_o2,
  G3335_o2,
  G3180_o2,
  G3340_o2,
  G3339_o2,
  G3341_o2,
  G3234_o2,
  G3829_o2,
  G3338_o2,
  G3336_o2,
  G3770_o2,
  G3918_o2,
  G3774_o2,
  G3921_o2,
  G3832_o2,
  G3993_o2,
  G2076_o2,
  G2071_o2,
  G2072_o2,
  G2069_o2,
  G2070_o2,
  G2067_o2,
  G2068_o2,
  G4095_o2,
  G3272_o2,
  G3269_o2,
  G3270_o2,
  G3271_o2,
  G3265_o2,
  G3266_o2,
  G4137_o2,
  G3268_o2,
  G2361_o2,
  G3228_o2,
  G3267_o2,
  G2336_o2,
  G3459_o2,
  G3428_o2,
  G3438_o2,
  G3449_o2,
  G3421_o2,
  G3576_o2,
  G3303_o2,
  G3583_o2,
  G3594_o2,
  G3674_o2,
  G3685_o2,
  G4504_o2,
  G4180_o2,
  G5123_o2,
  G5142_o2,
  G5126_o2,
  G5144_o2,
  G3912_o2,
  G4417_o2,
  G4420_o2,
  G3969_o2,
  G4023_o2,
  G2720_o2,
  G2837_o2,
  n2965_inv,
  n2968_inv,
  n2971_inv,
  n2974_inv,
  G1876_o2,
  G4996_o2,
  G4984_o2,
  G4920_o2,
  G4923_o2,
  G4930_o2,
  G4933_o2,
  n4320_lo_buf_o2,
  G2424_o2,
  G3317_o2,
  G3503_o2,
  G3485_o2,
  G3611_o2,
  n3864_lo_buf_o2,
  n3888_lo_buf_o2,
  n4116_lo_buf_o2,
  n4128_lo_buf_o2,
  n4140_lo_buf_o2,
  n4152_lo_buf_o2,
  G1815_o2,
  G1728_o2,
  G1035_o2,
  G1041_o2,
  G1087_o2,
  G1093_o2,
  G1132_o2,
  G1108_o2,
  G1138_o2,
  G1114_o2,
  G1807_o2,
  G2108_o2,
  G1126_o2,
  G1899_o2,
  G2134_o2,
  G1852_o2,
  G2116_o2,
  G2543_o2,
  G2727_o2,
  G2715_o2,
  G2832_o2,
  G1873_o2,
  G3291_o2,
  G5025_o2,
  G5036_o2,
  G3132_o2,
  G5038_o2,
  G5039_o2,
  n3118_inv,
  n3121_inv,
  n3124_inv,
  n3127_inv,
  n3984_lo_buf_o2,
  G1802_o2,
  G1804_o2,
  G1849_o2,
  G1851_o2,
  G2492_o2,
  G1799_o2,
  G4231_o2,
  G4234_o2,
  G4245_o2,
  G4247_o2,
  G1894_o2,
  G1846_o2,
  G4238_o2,
  G4249_o2,
  G2293_o2,
  G5022_o2,
  G5006_o2,
  G4944_o2,
  G4946_o2,
  G4954_o2,
  G4956_o2,
  G3546_o2,
  G3658_o2,
  G1344_o2,
  G2921_o2,
  n3912_lo_buf_o2,
  G1835_o2,
  G3810_o2,
  G3866_o2,
  G3811_o2,
  G2269_o2,
  G3812_o2,
  G3867_o2,
  G3868_o2,
  G3809_o2,
  G3716_o2,
  G4529_o2,
  G4670_o2,
  G4493_o2,
  G4580_o2,
  G3822_o2,
  G3877_o2,
  G4131_o2,
  G4170_o2,
  G4051_o2,
  G4065_o2,
  G4697_o2,
  G4706_o2,
  G2460_o2,
  G2454_o2,
  G2392_o2,
  G2386_o2,
  n4260_lo_buf_o2,
  n4272_lo_buf_o2,
  n4392_lo_buf_o2,
  n4404_lo_buf_o2,
  G1512_o2,
  G3135_o2,
  G2379_o2,
  n4164_lo_buf_o2,
  n4176_lo_buf_o2,
  n4224_lo_buf_o2,
  G2975_o2,
  G2978_o2,
  G2933_o2,
  G2936_o2,
  G1356_o2,
  G1359_o2,
  G1398_o2,
  G1401_o2,
  G5193,
  G5194,
  G5195,
  G5196,
  G5197,
  G5198,
  G5199,
  G5200,
  G5201,
  G5202,
  G5203,
  G5204,
  G5205,
  G5206,
  G5207,
  G5208,
  G5209,
  G5210,
  G5211,
  G5212,
  G5213,
  G5214,
  G5215,
  G5216,
  G5217,
  G5218,
  G5219,
  G5220,
  G5221,
  G5222,
  G5223,
  G5224,
  G5225,
  G5226,
  G5227,
  G5228,
  G5229,
  G5230,
  G5231,
  G5232,
  G5233,
  G5234,
  G5235,
  G5236,
  G5237,
  G5238,
  G5239,
  G5240,
  G5241,
  G5242,
  G5243,
  G5244,
  G5245,
  G5246,
  G5247,
  G5248,
  G5249,
  G5250,
  G5251,
  G5252,
  G5253,
  G5254,
  G5255,
  G5256,
  G5257,
  G5258,
  G5259,
  G5260,
  G5261,
  G5262,
  G5263,
  G5264,
  G5265,
  G5266,
  G5267,
  G5268,
  G5269,
  G5270,
  G5271,
  G5272,
  G5273,
  G5274,
  G5275,
  G5276,
  G5277,
  G5278,
  G5279,
  G5280,
  G5281,
  G5282,
  G5283,
  G5284,
  G5285,
  G5286,
  G5287,
  G5288,
  G5289,
  G5290,
  G5291,
  G5292,
  G5293,
  G5294,
  G5295,
  G5296,
  G5297,
  G5298,
  G5299,
  G5300,
  G5301,
  G5302,
  G5303,
  G5304,
  G5305,
  G5306,
  G5307,
  G5308,
  G5309,
  G5310,
  G5311,
  G5312,
  G5313,
  G5314,
  G5315,
  n2610_li,
  n2613_li,
  n2616_li,
  n2619_li,
  n2622_li,
  n2625_li,
  n2628_li,
  n2631_li,
  n2634_li,
  n2637_li,
  n2640_li,
  n2643_li,
  n2646_li,
  n2649_li,
  n2652_li,
  n2655_li,
  n2658_li,
  n2661_li,
  n2664_li,
  n2667_li,
  n2670_li,
  n2673_li,
  n2676_li,
  n2679_li,
  n2682_li,
  n2685_li,
  n2688_li,
  n2691_li,
  n2694_li,
  n2697_li,
  n2700_li,
  n2703_li,
  n2706_li,
  n2709_li,
  n2712_li,
  n2715_li,
  n2718_li,
  n2721_li,
  n2724_li,
  n2727_li,
  n2730_li,
  n2733_li,
  n2736_li,
  n2739_li,
  n2742_li,
  n2745_li,
  n2748_li,
  n2751_li,
  n2754_li,
  n2757_li,
  n2760_li,
  n2763_li,
  n2766_li,
  n2769_li,
  n2772_li,
  n2775_li,
  n2778_li,
  n2781_li,
  n2784_li,
  n2787_li,
  n2790_li,
  n2793_li,
  n2796_li,
  n2799_li,
  n2802_li,
  n2805_li,
  n2808_li,
  n2811_li,
  n2814_li,
  n2817_li,
  n2820_li,
  n2823_li,
  n2826_li,
  n2829_li,
  n2832_li,
  n2835_li,
  n2838_li,
  n2841_li,
  n2844_li,
  n2847_li,
  n2850_li,
  n2853_li,
  n2856_li,
  n2859_li,
  n2862_li,
  n2865_li,
  n2868_li,
  n2871_li,
  n2874_li,
  n2877_li,
  n2880_li,
  n2883_li,
  n2886_li,
  n2889_li,
  n2892_li,
  n2895_li,
  n2898_li,
  n2901_li,
  n2904_li,
  n2907_li,
  n2910_li,
  n2913_li,
  n2916_li,
  n2919_li,
  n2922_li,
  n2925_li,
  n2928_li,
  n2931_li,
  n2934_li,
  n2937_li,
  n2940_li,
  n2943_li,
  n2946_li,
  n2949_li,
  n2952_li,
  n2955_li,
  n2958_li,
  n2961_li,
  n2964_li,
  n2967_li,
  n2970_li,
  n2973_li,
  n2976_li,
  n2979_li,
  n2982_li,
  n2985_li,
  n2988_li,
  n2991_li,
  n2994_li,
  n2997_li,
  n3000_li,
  n3003_li,
  n3006_li,
  n3009_li,
  n3012_li,
  n3015_li,
  n3018_li,
  n3021_li,
  n3024_li,
  n3027_li,
  n3030_li,
  n3033_li,
  n3036_li,
  n3039_li,
  n3042_li,
  n3045_li,
  n3048_li,
  n3051_li,
  n3054_li,
  n3057_li,
  n3060_li,
  n3063_li,
  n3066_li,
  n3069_li,
  n3072_li,
  n3075_li,
  n3078_li,
  n3081_li,
  n3084_li,
  n3087_li,
  n3090_li,
  n3093_li,
  n3096_li,
  n3099_li,
  n3102_li,
  n3105_li,
  n3108_li,
  n3111_li,
  n3114_li,
  n3117_li,
  n3120_li,
  n3123_li,
  n3126_li,
  n3129_li,
  n3132_li,
  n3135_li,
  n3138_li,
  n3141_li,
  n3144_li,
  n3147_li,
  n3150_li,
  n3153_li,
  n3156_li,
  n3159_li,
  n3162_li,
  n3165_li,
  n3168_li,
  n3171_li,
  n3174_li,
  n3177_li,
  n3180_li,
  n3183_li,
  n3186_li,
  n3189_li,
  n3192_li,
  n3195_li,
  n3198_li,
  n3201_li,
  n3204_li,
  n3207_li,
  n3210_li,
  n3213_li,
  n3216_li,
  n3219_li,
  n3222_li,
  n3225_li,
  n3228_li,
  n3231_li,
  n3234_li,
  n3237_li,
  n3240_li,
  n3243_li,
  n3246_li,
  n3249_li,
  n3252_li,
  n3255_li,
  n3258_li,
  n3261_li,
  n3264_li,
  n3267_li,
  n3270_li,
  n3273_li,
  n3276_li,
  n3279_li,
  n3282_li,
  n3285_li,
  n3288_li,
  n3291_li,
  n3294_li,
  n3297_li,
  n3300_li,
  n3303_li,
  n3306_li,
  n3309_li,
  n3312_li,
  n3315_li,
  n3318_li,
  n3321_li,
  n3324_li,
  n3327_li,
  n3330_li,
  n3333_li,
  n3336_li,
  n3339_li,
  n3342_li,
  n3345_li,
  n3348_li,
  n3351_li,
  n3354_li,
  n3357_li,
  n3360_li,
  n3363_li,
  n3366_li,
  n3369_li,
  n3372_li,
  n3375_li,
  n3378_li,
  n3381_li,
  n3384_li,
  n3387_li,
  n3390_li,
  n3393_li,
  n3396_li,
  n3399_li,
  n3402_li,
  n3405_li,
  n3408_li,
  n3411_li,
  n3414_li,
  n3417_li,
  n3420_li,
  n3423_li,
  n3426_li,
  n3429_li,
  n3432_li,
  n3435_li,
  n3438_li,
  n3441_li,
  n3444_li,
  n3447_li,
  n3450_li,
  n3453_li,
  n3456_li,
  n3459_li,
  n3462_li,
  n3465_li,
  n3468_li,
  n3471_li,
  n3474_li,
  n3477_li,
  n3480_li,
  n3483_li,
  n3486_li,
  n3489_li,
  n3492_li,
  n3495_li,
  n3498_li,
  n3501_li,
  n3504_li,
  n3507_li,
  n3510_li,
  n3513_li,
  n3516_li,
  n3519_li,
  n3522_li,
  n3525_li,
  n3528_li,
  n3531_li,
  n3534_li,
  n3537_li,
  n3540_li,
  n3543_li,
  n3546_li,
  n3549_li,
  n3552_li,
  n3555_li,
  n3558_li,
  n3561_li,
  n3564_li,
  n3567_li,
  n3570_li,
  n3573_li,
  n3576_li,
  n3579_li,
  n3582_li,
  n3585_li,
  n3588_li,
  n3591_li,
  n3594_li,
  n3597_li,
  n3600_li,
  n3603_li,
  n3606_li,
  n3609_li,
  n3612_li,
  n3615_li,
  n3618_li,
  n3621_li,
  n3624_li,
  n3627_li,
  n3630_li,
  n3633_li,
  n3636_li,
  n3639_li,
  n3642_li,
  n3645_li,
  n3648_li,
  n3651_li,
  n3654_li,
  n3657_li,
  n3666_li,
  n3669_li,
  n3678_li,
  n3687_li,
  n3690_li,
  n3702_li,
  n3711_li,
  n3714_li,
  n3726_li,
  n3735_li,
  n3738_li,
  n3750_li,
  n3753_li,
  n3759_li,
  n3762_li,
  n3765_li,
  n3774_li,
  n3777_li,
  n3786_li,
  n3789_li,
  n3792_li,
  n3795_li,
  n3798_li,
  n3801_li,
  n3810_li,
  n3813_li,
  n3822_li,
  n3825_li,
  n3834_li,
  n3843_li,
  n3846_li,
  n3867_li,
  n3891_li,
  n3915_li,
  n3930_li,
  n3933_li,
  n3936_li,
  n3942_li,
  n3945_li,
  n3948_li,
  n3954_li,
  n3957_li,
  n3963_li,
  n3966_li,
  n3969_li,
  n3975_li,
  n3978_li,
  n3987_li,
  n3990_li,
  n4002_li,
  n4011_li,
  n4014_li,
  n4026_li,
  n4035_li,
  n4038_li,
  n4050_li,
  n4053_li,
  n4059_li,
  n4062_li,
  n4065_li,
  n4098_li,
  n4107_li,
  n4119_li,
  n4131_li,
  n4143_li,
  n4155_li,
  n4167_li,
  n4179_li,
  n4182_li,
  n4185_li,
  n4188_li,
  n4194_li,
  n4197_li,
  n4200_li,
  n4206_li,
  n4209_li,
  n4212_li,
  n4215_li,
  n4227_li,
  n4230_li,
  n4233_li,
  n4236_li,
  n4239_li,
  n4242_li,
  n4251_li,
  n4263_li,
  n4275_li,
  n4278_li,
  n4287_li,
  n4290_li,
  n4293_li,
  n4299_li,
  n4302_li,
  n4305_li,
  n4311_li,
  n4314_li,
  n4323_li,
  n4326_li,
  n4335_li,
  n4338_li,
  n4347_li,
  n4350_li,
  n4359_li,
  n4362_li,
  n4365_li,
  n4371_li,
  n4374_li,
  n4383_li,
  n4395_li,
  n4407_li,
  n4410_li,
  n4413_li,
  n4416_li,
  n4419_li,
  n4422_li,
  n4425_li,
  n4428_li,
  n4431_li,
  n4434_li,
  n4437_li,
  n4440_li,
  n4443_li,
  n4446_li,
  n4449_li,
  n4452_li,
  n4455_li,
  n4458_li,
  n4461_li,
  n4464_li,
  n4467_li,
  n4470_li,
  n4473_li,
  n4476_li,
  n4479_li,
  n4482_li,
  n4485_li,
  n4488_li,
  n4494_li,
  n4497_li,
  n4500_li,
  n4503_li,
  n4506_li,
  n4509_li,
  n4512_li,
  n4515_li,
  n4518_li,
  n4521_li,
  n4524_li,
  n4527_li,
  n4530_li,
  n4533_li,
  n4536_li,
  n4539_li,
  n4542_li,
  n4545_li,
  n4548_li,
  n4554_li,
  n4557_li,
  n4560_li,
  n4563_li,
  n4566_li,
  n4569_li,
  n4572_li,
  n4575_li,
  n4578_li,
  n4581_li,
  n4584_li,
  n4587_li,
  n4590_li,
  n4593_li,
  n4596_li,
  n4599_li,
  n4602_li,
  n4605_li,
  n4608_li,
  n4611_li,
  n4614_li,
  n4617_li,
  n4620_li,
  n4623_li,
  n4626_li,
  n4629_li,
  n4632_li,
  n4635_li,
  n4638_li,
  n4641_li,
  n4644_li,
  n4647_li,
  n4650_li,
  n4653_li,
  n4656_li,
  n4659_li,
  n4662_li,
  n4665_li,
  n4668_li,
  n4671_li,
  n4674_li,
  n4677_li,
  n4680_li,
  n4683_li,
  n4686_li,
  n4689_li,
  n4692_li,
  n4695_li,
  n4698_li,
  n4701_li,
  n4704_li,
  n4707_li,
  n4710_li,
  n4713_li,
  n4716_li,
  n4719_li,
  n4722_li,
  n4725_li,
  n4728_li,
  n4731_li,
  n4734_li,
  n4737_li,
  n4740_li,
  n4743_li,
  n6382_i2,
  n6383_i2,
  n6419_i2,
  n6420_i2,
  n6435_i2,
  n6436_i2,
  n6448_i2,
  n6449_i2,
  n6613_i2,
  n6614_i2,
  n6641_i2,
  n6658_i2,
  n6757_i2,
  n6756_i2,
  n7116_i2,
  n7156_i2,
  n6549_i2,
  n6550_i2,
  n7357_i2,
  n7358_i2,
  n7359_i2,
  n7360_i2,
  n6621_i2,
  n6623_i2,
  n6625_i2,
  n6626_i2,
  n6627_i2,
  n6628_i2,
  n6629_i2,
  n6630_i2,
  n6669_i2,
  n7449_i2,
  n7450_i2,
  n7451_i2,
  n7452_i2,
  n6682_i2,
  n6683_i2,
  n6684_i2,
  n6685_i2,
  n7463_i2,
  n6686_i2,
  n6687_i2,
  n6688_i2,
  n6689_i2,
  n6772_i2,
  n6773_i2,
  n6774_i2,
  n6775_i2,
  G3467_i2,
  G2810_i2,
  n6833_i2,
  n6945_i2,
  n6947_i2,
  n6949_i2,
  n6951_i2,
  n6888_i2,
  n6889_i2,
  n6936_i2,
  n6954_i2,
  n6955_i2,
  n6956_i2,
  n6957_i2,
  n6958_i2,
  n6982_i2,
  n6984_i2,
  n6974_i2,
  n6975_i2,
  n6999_i2,
  n7015_i2,
  n7016_i2,
  n7017_i2,
  n7018_i2,
  n7005_i2,
  n7019_i2,
  n7022_i2,
  n7023_i2,
  n7132_i2,
  n7133_i2,
  n7135_i2,
  n7136_i2,
  n7175_i2,
  n7155_i2,
  G3060_i2,
  n7383_i2,
  G3802_i2,
  G3859_i2,
  n7355_i2,
  n7356_i2,
  G4054_i2,
  G4068_i2,
  n7384_i2,
  n7387_i2,
  n7388_i2,
  n7389_i2,
  n7386_i2,
  n7453_i2,
  n7431_i2,
  n7432_i2,
  n7433_i2,
  n7430_i2,
  n7485_i2,
  n7486_i2,
  G2508_i2,
  G2486_i2,
  n7245_i2,
  n7246_i2,
  n3756_lo_buf_i2,
  n4056_lo_buf_i2,
  G3474_i2,
  G2817_i2,
  n7396_i2,
  n7398_i2,
  n7400_i2,
  n7401_i2,
  n7402_i2,
  n7403_i2,
  n7404_i2,
  n7405_i2,
  G2711_i2,
  G2828_i2,
  n7490_i2,
  n7527_i2,
  n7528_i2,
  n7529_i2,
  n7530_i2,
  n7523_i2,
  n7524_i2,
  n7525_i2,
  n7526_i2,
  n4296_lo_buf_i2,
  n4368_lo_buf_i2,
  G2466_i2,
  G2404_i2,
  n7534_i2,
  n7535_i2,
  n7536_i2,
  n7533_i2,
  G1060_i2,
  G963_i2,
  G2448_i2,
  G2685_i2,
  G2679_i2,
  G2774_i2,
  G2780_i2,
  G2759_i2,
  G2737_i2,
  G2850_i2,
  G3393_i2,
  G3404_i2,
  G3559_i2,
  G2744_i2,
  n3708_lo_buf_i2,
  n3840_lo_buf_i2,
  n4008_lo_buf_i2,
  n4104_lo_buf_i2,
  G1821_i2,
  G1734_i2,
  G3517_i2,
  G3533_i2,
  G3629_i2,
  G3645_i2,
  G2857_i2,
  G2731_i2,
  G2844_i2,
  n3732_lo_buf_i2,
  n4032_lo_buf_i2,
  G3552_i2,
  G2271_i2,
  n4248_lo_buf_i2,
  n4332_lo_buf_i2,
  n4344_lo_buf_i2,
  n4380_lo_buf_i2,
  G2398_i2,
  G2480_i2,
  G2418_i2,
  G1455_i2,
  G1449_i2,
  G1452_i2,
  G1425_i2,
  G1428_i2,
  G1419_i2,
  G1422_i2,
  n4308_lo_buf_i2,
  G2675_i2,
  G3035_i2,
  G3026_i2,
  G3029_i2,
  G3032_i2,
  G2999_i2,
  G3002_i2,
  G2770_i2,
  G3008_i2,
  G2073_i2,
  G2752_i2,
  G3005_i2,
  G5108_i2,
  G5135_i2,
  G5111_i2,
  G5138_i2,
  G3415_i2,
  G3386_i2,
  G3570_i2,
  G2430_i2,
  G3495_i2,
  G3621_i2,
  n4284_lo_buf_i2,
  n4356_lo_buf_i2,
  G2472_i2,
  G2410_i2,
  n3960_lo_buf_i2,
  n3972_lo_buf_i2,
  G2865_i2,
  G970_i2,
  n3684_lo_buf_i2,
  n4080_lo_buf_i2,
  n4092_lo_buf_i2,
  G1053_i2,
  G956_i2,
  G1147_i2,
  G2705_i2,
  G2693_i2,
  G2696_i2,
  G2700_i2,
  G2915_i2,
  G2966_i2,
  G2540_i2,
  G2788_i2,
  G2792_i2,
  G2797_i2,
  G2804_i2,
  G1038_i2,
  G1044_i2,
  G1090_i2,
  G1096_i2,
  G1029_i2,
  G3942_i2,
  G3954_i2,
  G4011_i2,
  G4017_i2,
  G1141_i2,
  G1081_i2,
  G2146_i2,
  G2145_i2,
  G2144_i2,
  G2143_i2,
  G2142_i2,
  G2141_i2,
  G2140_i2,
  G2139_i2,
  G3769_i2,
  G3773_i2,
  G3768_i2,
  G4101_i2,
  G3161_i2,
  G4143_i2,
  G3828_i2,
  G3831_i2,
  G3334_i2,
  G3335_i2,
  G3180_i2,
  G3340_i2,
  G3339_i2,
  G3341_i2,
  G3234_i2,
  G3829_i2,
  G3338_i2,
  G3336_i2,
  G3770_i2,
  G3918_i2,
  G3774_i2,
  G3921_i2,
  G3832_i2,
  G3993_i2,
  G2076_i2,
  G2071_i2,
  G2072_i2,
  G2069_i2,
  G2070_i2,
  G2067_i2,
  G2068_i2,
  G4095_i2,
  G3272_i2,
  G3269_i2,
  G3270_i2,
  G3271_i2,
  G3265_i2,
  G3266_i2,
  G4137_i2,
  G3268_i2,
  G2361_i2,
  G3228_i2,
  G3267_i2,
  G2336_i2,
  G3459_i2,
  G3428_i2,
  G3438_i2,
  G3449_i2,
  G3421_i2,
  G3576_i2,
  G3303_i2,
  G3583_i2,
  G3594_i2,
  G3674_i2,
  G3685_i2,
  G4504_i2,
  G4180_i2,
  G5123_i2,
  G5142_i2,
  G5126_i2,
  G5144_i2,
  G3912_i2,
  G4417_i2,
  G4420_i2,
  G3969_i2,
  G4023_i2,
  G2720_i2,
  G2837_i2,
  G836_i2,
  G848_i2,
  G813_i2,
  G825_i2,
  G1876_i2,
  G4996_i2,
  G4984_i2,
  G4920_i2,
  G4923_i2,
  G4930_i2,
  G4933_i2,
  n4320_lo_buf_i2,
  G2424_i2,
  G3317_i2,
  G3503_i2,
  G3485_i2,
  G3611_i2,
  n3864_lo_buf_i2,
  n3888_lo_buf_i2,
  n4116_lo_buf_i2,
  n4128_lo_buf_i2,
  n4140_lo_buf_i2,
  n4152_lo_buf_i2,
  G1815_i2,
  G1728_i2,
  G1035_i2,
  G1041_i2,
  G1087_i2,
  G1093_i2,
  G1132_i2,
  G1108_i2,
  G1138_i2,
  G1114_i2,
  G1807_i2,
  G2108_i2,
  G1126_i2,
  G1899_i2,
  G2134_i2,
  G1852_i2,
  G2116_i2,
  G2543_i2,
  G2727_i2,
  G2715_i2,
  G2832_i2,
  G1873_i2,
  G3291_i2,
  G5025_i2,
  G5036_i2,
  G3132_i2,
  G5038_i2,
  G5039_i2,
  G1150_i2,
  G1162_i2,
  G804_i2,
  G1172_i2,
  n3984_lo_buf_i2,
  G1802_i2,
  G1804_i2,
  G1849_i2,
  G1851_i2,
  G2492_i2,
  G1799_i2,
  G4231_i2,
  G4234_i2,
  G4245_i2,
  G4247_i2,
  G1894_i2,
  G1846_i2,
  G4238_i2,
  G4249_i2,
  G2293_i2,
  G5022_i2,
  G5006_i2,
  G4944_i2,
  G4946_i2,
  G4954_i2,
  G4956_i2,
  G3546_i2,
  G3658_i2,
  G1344_i2,
  G2921_i2,
  n3912_lo_buf_i2,
  G1835_i2,
  G3810_i2,
  G3866_i2,
  G3811_i2,
  G2269_i2,
  G3812_i2,
  G3867_i2,
  G3868_i2,
  G3809_i2,
  G3716_i2,
  G4529_i2,
  G4670_i2,
  G4493_i2,
  G4580_i2,
  G3822_i2,
  G3877_i2,
  G4131_i2,
  G4170_i2,
  G4051_i2,
  G4065_i2,
  G4697_i2,
  G4706_i2,
  G2460_i2,
  G2454_i2,
  G2392_i2,
  G2386_i2,
  n4260_lo_buf_i2,
  n4272_lo_buf_i2,
  n4392_lo_buf_i2,
  n4404_lo_buf_i2,
  G1512_i2,
  G3135_i2,
  G2379_i2,
  n4164_lo_buf_i2,
  n4176_lo_buf_i2,
  n4224_lo_buf_i2,
  G2975_i2,
  G2978_i2,
  G2933_i2,
  G2936_i2,
  G1356_i2,
  G1359_i2,
  G1398_i2,
  G1401_i2
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input G42;input G43;input G44;input G45;input G46;input G47;input G48;input G49;input G50;input G51;input G52;input G53;input G54;input G55;input G56;input G57;input G58;input G59;input G60;input G61;input G62;input G63;input G64;input G65;input G66;input G67;input G68;input G69;input G70;input G71;input G72;input G73;input G74;input G75;input G76;input G77;input G78;input G79;input G80;input G81;input G82;input G83;input G84;input G85;input G86;input G87;input G88;input G89;input G90;input G91;input G92;input G93;input G94;input G95;input G96;input G97;input G98;input G99;input G100;input G101;input G102;input G103;input G104;input G105;input G106;input G107;input G108;input G109;input G110;input G111;input G112;input G113;input G114;input G115;input G116;input G117;input G118;input G119;input G120;input G121;input G122;input G123;input G124;input G125;input G126;input G127;input G128;input G129;input G130;input G131;input G132;input G133;input G134;input G135;input G136;input G137;input G138;input G139;input G140;input G141;input G142;input G143;input G144;input G145;input G146;input G147;input G148;input G149;input G150;input G151;input G152;input G153;input G154;input G155;input G156;input G157;input G158;input G159;input G160;input G161;input G162;input G163;input G164;input G165;input G166;input G167;input G168;input G169;input G170;input G171;input G172;input G173;input G174;input G175;input G176;input G177;input G178;input n2610_lo;input n2613_lo;input n2616_lo;input n2619_lo;input n2622_lo;input n2625_lo;input n2628_lo;input n2631_lo;input n2634_lo;input n2637_lo;input n2640_lo;input n2643_lo;input n2646_lo;input n2649_lo;input n2652_lo;input n2655_lo;input n2658_lo;input n2661_lo;input n2664_lo;input n2667_lo;input n2670_lo;input n2673_lo;input n2676_lo;input n2679_lo;input n2682_lo;input n2685_lo;input n2688_lo;input n2691_lo;input n2694_lo;input n2697_lo;input n2700_lo;input n2703_lo;input n2706_lo;input n2709_lo;input n2712_lo;input n2715_lo;input n2718_lo;input n2721_lo;input n2724_lo;input n2727_lo;input n2730_lo;input n2733_lo;input n2736_lo;input n2739_lo;input n2742_lo;input n2745_lo;input n2748_lo;input n2751_lo;input n2754_lo;input n2757_lo;input n2760_lo;input n2763_lo;input n2766_lo;input n2769_lo;input n2772_lo;input n2775_lo;input n2778_lo;input n2781_lo;input n2784_lo;input n2787_lo;input n2790_lo;input n2793_lo;input n2796_lo;input n2799_lo;input n2802_lo;input n2805_lo;input n2808_lo;input n2811_lo;input n2814_lo;input n2817_lo;input n2820_lo;input n2823_lo;input n2826_lo;input n2829_lo;input n2832_lo;input n2835_lo;input n2838_lo;input n2841_lo;input n2844_lo;input n2847_lo;input n2850_lo;input n2853_lo;input n2856_lo;input n2859_lo;input n2862_lo;input n2865_lo;input n2868_lo;input n2871_lo;input n2874_lo;input n2877_lo;input n2880_lo;input n2883_lo;input n2886_lo;input n2889_lo;input n2892_lo;input n2895_lo;input n2898_lo;input n2901_lo;input n2904_lo;input n2907_lo;input n2910_lo;input n2913_lo;input n2916_lo;input n2919_lo;input n2922_lo;input n2925_lo;input n2928_lo;input n2931_lo;input n2934_lo;input n2937_lo;input n2940_lo;input n2943_lo;input n2946_lo;input n2949_lo;input n2952_lo;input n2955_lo;input n2958_lo;input n2961_lo;input n2964_lo;input n2967_lo;input n2970_lo;input n2973_lo;input n2976_lo;input n2979_lo;input n2982_lo;input n2985_lo;input n2988_lo;input n2991_lo;input n2994_lo;input n2997_lo;input n3000_lo;input n3003_lo;input n3006_lo;input n3009_lo;input n3012_lo;input n3015_lo;input n3018_lo;input n3021_lo;input n3024_lo;input n3027_lo;input n3030_lo;input n3033_lo;input n3036_lo;input n3039_lo;input n3042_lo;input n3045_lo;input n3048_lo;input n3051_lo;input n3054_lo;input n3057_lo;input n3060_lo;input n3063_lo;input n3066_lo;input n3069_lo;input n3072_lo;input n3075_lo;input n3078_lo;input n3081_lo;input n3084_lo;input n3087_lo;input n3090_lo;input n3093_lo;input n3096_lo;input n3099_lo;input n3102_lo;input n3105_lo;input n3108_lo;input n3111_lo;input n3114_lo;input n3117_lo;input n3120_lo;input n3123_lo;input n3126_lo;input n3129_lo;input n3132_lo;input n3135_lo;input n3138_lo;input n3141_lo;input n3144_lo;input n3147_lo;input n3150_lo;input n3153_lo;input n3156_lo;input n3159_lo;input n3162_lo;input n3165_lo;input n3168_lo;input n3171_lo;input n3174_lo;input n3177_lo;input n3180_lo;input n3183_lo;input n3186_lo;input n3189_lo;input n3192_lo;input n3195_lo;input n3198_lo;input n3201_lo;input n3204_lo;input n3207_lo;input n3210_lo;input n3213_lo;input n3216_lo;input n3219_lo;input n3222_lo;input n3225_lo;input n3228_lo;input n3231_lo;input n3234_lo;input n3237_lo;input n3240_lo;input n3243_lo;input n3246_lo;input n3249_lo;input n3252_lo;input n3255_lo;input n3258_lo;input n3261_lo;input n3264_lo;input n3267_lo;input n3270_lo;input n3273_lo;input n3276_lo;input n3279_lo;input n3282_lo;input n3285_lo;input n3288_lo;input n3291_lo;input n3294_lo;input n3297_lo;input n3300_lo;input n3303_lo;input n3306_lo;input n3309_lo;input n3312_lo;input n3315_lo;input n3318_lo;input n3321_lo;input n3324_lo;input n3327_lo;input n3330_lo;input n3333_lo;input n3336_lo;input n3339_lo;input n3342_lo;input n3345_lo;input n3348_lo;input n3351_lo;input n3354_lo;input n3357_lo;input n3360_lo;input n3363_lo;input n3366_lo;input n3369_lo;input n3372_lo;input n3375_lo;input n3378_lo;input n3381_lo;input n3384_lo;input n3387_lo;input n3390_lo;input n3393_lo;input n3396_lo;input n3399_lo;input n3402_lo;input n3405_lo;input n3408_lo;input n3411_lo;input n3414_lo;input n3417_lo;input n3420_lo;input n3423_lo;input n3426_lo;input n3429_lo;input n3432_lo;input n3435_lo;input n3438_lo;input n3441_lo;input n3444_lo;input n3447_lo;input n3450_lo;input n3453_lo;input n3456_lo;input n3459_lo;input n3462_lo;input n3465_lo;input n3468_lo;input n3471_lo;input n3474_lo;input n3477_lo;input n3480_lo;input n3483_lo;input n3486_lo;input n3489_lo;input n3492_lo;input n3495_lo;input n3498_lo;input n3501_lo;input n3504_lo;input n3507_lo;input n3510_lo;input n3513_lo;input n3516_lo;input n3519_lo;input n3522_lo;input n3525_lo;input n3528_lo;input n3531_lo;input n3534_lo;input n3537_lo;input n3540_lo;input n3543_lo;input n3546_lo;input n3549_lo;input n3552_lo;input n3555_lo;input n3558_lo;input n3561_lo;input n3564_lo;input n3567_lo;input n3570_lo;input n3573_lo;input n3576_lo;input n3579_lo;input n3582_lo;input n3585_lo;input n3588_lo;input n3591_lo;input n3594_lo;input n3597_lo;input n3600_lo;input n3603_lo;input n3606_lo;input n3609_lo;input n3612_lo;input n3615_lo;input n3618_lo;input n3621_lo;input n3624_lo;input n3627_lo;input n3630_lo;input n3633_lo;input n3636_lo;input n3639_lo;input n3642_lo;input n3645_lo;input n3648_lo;input n3651_lo;input n3654_lo;input n3657_lo;input n3666_lo;input n3669_lo;input n3678_lo;input n3687_lo;input n3690_lo;input n3702_lo;input n3711_lo;input n3714_lo;input n3726_lo;input n3735_lo;input n3738_lo;input n3750_lo;input n3753_lo;input n3759_lo;input n3762_lo;input n3765_lo;input n3774_lo;input n3777_lo;input n3786_lo;input n3789_lo;input n3792_lo;input n3795_lo;input n3798_lo;input n3801_lo;input n3810_lo;input n3813_lo;input n3822_lo;input n3825_lo;input n3834_lo;input n3843_lo;input n3846_lo;input n3867_lo;input n3891_lo;input n3915_lo;input n3930_lo;input n3933_lo;input n3936_lo;input n3942_lo;input n3945_lo;input n3948_lo;input n3954_lo;input n3957_lo;input n3963_lo;input n3966_lo;input n3969_lo;input n3975_lo;input n3978_lo;input n3987_lo;input n3990_lo;input n4002_lo;input n4011_lo;input n4014_lo;input n4026_lo;input n4035_lo;input n4038_lo;input n4050_lo;input n4053_lo;input n4059_lo;input n4062_lo;input n4065_lo;input n4098_lo;input n4107_lo;input n4119_lo;input n4131_lo;input n4143_lo;input n4155_lo;input n4167_lo;input n4179_lo;input n4182_lo;input n4185_lo;input n4188_lo;input n4194_lo;input n4197_lo;input n4200_lo;input n4206_lo;input n4209_lo;input n4212_lo;input n4215_lo;input n4227_lo;input n4230_lo;input n4233_lo;input n4236_lo;input n4239_lo;input n4242_lo;input n4251_lo;input n4263_lo;input n4275_lo;input n4278_lo;input n4287_lo;input n4290_lo;input n4293_lo;input n4299_lo;input n4302_lo;input n4305_lo;input n4311_lo;input n4314_lo;input n4323_lo;input n4326_lo;input n4335_lo;input n4338_lo;input n4347_lo;input n4350_lo;input n4359_lo;input n4362_lo;input n4365_lo;input n4371_lo;input n4374_lo;input n4383_lo;input n4395_lo;input n4407_lo;input n4410_lo;input n4413_lo;input n4416_lo;input n4419_lo;input n4422_lo;input n4425_lo;input n4428_lo;input n4431_lo;input n4434_lo;input n4437_lo;input n4440_lo;input n4443_lo;input n4446_lo;input n4449_lo;input n4452_lo;input n4455_lo;input n4458_lo;input n4461_lo;input n4464_lo;input n4467_lo;input n4470_lo;input n4473_lo;input n4476_lo;input n4479_lo;input n4482_lo;input n4485_lo;input n4488_lo;input n4494_lo;input n4497_lo;input n4500_lo;input n4503_lo;input n4506_lo;input n4509_lo;input n4512_lo;input n4515_lo;input n4518_lo;input n4521_lo;input n4524_lo;input n4527_lo;input n4530_lo;input n4533_lo;input n4536_lo;input n4539_lo;input n4542_lo;input n4545_lo;input n4548_lo;input n4554_lo;input n4557_lo;input n4560_lo;input n4563_lo;input n4566_lo;input n4569_lo;input n4572_lo;input n4575_lo;input n4578_lo;input n4581_lo;input n4584_lo;input n4587_lo;input n4590_lo;input n4593_lo;input n4596_lo;input n4599_lo;input n4602_lo;input n4605_lo;input n4608_lo;input n4611_lo;input n4614_lo;input n4617_lo;input n4620_lo;input n4623_lo;input n4626_lo;input n4629_lo;input n4632_lo;input n4635_lo;input n4638_lo;input n4641_lo;input n4644_lo;input n4647_lo;input n4650_lo;input n4653_lo;input n4656_lo;input n4659_lo;input n4662_lo;input n4665_lo;input n4668_lo;input n4671_lo;input n4674_lo;input n4677_lo;input n4680_lo;input n4683_lo;input n4686_lo;input n4689_lo;input n4692_lo;input n4695_lo;input n4698_lo;input n4701_lo;input n4704_lo;input n4707_lo;input n4710_lo;input n4713_lo;input n4716_lo;input n4719_lo;input n4722_lo;input n4725_lo;input n4728_lo;input n4731_lo;input n4734_lo;input n4737_lo;input n4740_lo;input n4743_lo;input n6382_o2;input n6383_o2;input n6419_o2;input n6420_o2;input n6435_o2;input n6436_o2;input n6448_o2;input n6449_o2;input n6613_o2;input n6614_o2;input n6641_o2;input n6658_o2;input n6757_o2;input n6756_o2;input n7116_o2;input n7156_o2;input n6549_o2;input n6550_o2;input n7357_o2;input n7358_o2;input n7359_o2;input n7360_o2;input n6621_o2;input n6623_o2;input n6625_o2;input n6626_o2;input n6627_o2;input n6628_o2;input n6629_o2;input n6630_o2;input n6669_o2;input n7449_o2;input n7450_o2;input n7451_o2;input n7452_o2;input n6682_o2;input n6683_o2;input n6684_o2;input n6685_o2;input n7463_o2;input n6686_o2;input n6687_o2;input n6688_o2;input n6689_o2;input n6772_o2;input n6773_o2;input n6774_o2;input n6775_o2;input G3467_o2;input G2810_o2;input n6833_o2;input n6945_o2;input n6947_o2;input n6949_o2;input n6951_o2;input n6888_o2;input n6889_o2;input n6936_o2;input n6954_o2;input n6955_o2;input n6956_o2;input n6957_o2;input n6958_o2;input n6982_o2;input n6984_o2;input n6974_o2;input n6975_o2;input n6999_o2;input n7015_o2;input n7016_o2;input n7017_o2;input n7018_o2;input n7005_o2;input n7019_o2;input n7022_o2;input n7023_o2;input n7132_o2;input n7133_o2;input n7135_o2;input n7136_o2;input n7175_o2;input n7155_o2;input G3060_o2;input n7383_o2;input G3802_o2;input G3859_o2;input n7355_o2;input n7356_o2;input G4054_o2;input G4068_o2;input n7384_o2;input n7387_o2;input n7388_o2;input n7389_o2;input n7386_o2;input n7453_o2;input n7431_o2;input n7432_o2;input n7433_o2;input n7430_o2;input n7485_o2;input n7486_o2;input G2508_o2;input G2486_o2;input n2326_inv;input n2329_inv;input n3756_lo_buf_o2;input n4056_lo_buf_o2;input G3474_o2;input n2341_inv;input n7396_o2;input n7398_o2;input n7400_o2;input n7401_o2;input n7402_o2;input n7403_o2;input n7404_o2;input n7405_o2;input G2711_o2;input n2371_inv;input n7490_o2;input n7527_o2;input n7528_o2;input n7529_o2;input n7530_o2;input n7523_o2;input n7524_o2;input n7525_o2;input n7526_o2;input n4296_lo_buf_o2;input n4368_lo_buf_o2;input G2466_o2;input G2404_o2;input n7534_o2;input n7535_o2;input n7536_o2;input n7533_o2;input G1060_o2;input G963_o2;input G2448_o2;input G2685_o2;input G2679_o2;input G2774_o2;input G2780_o2;input G2759_o2;input G2737_o2;input G2850_o2;input G3393_o2;input G3404_o2;input G3559_o2;input G2744_o2;input n3708_lo_buf_o2;input n3840_lo_buf_o2;input n4008_lo_buf_o2;input n4104_lo_buf_o2;input G1821_o2;input G1734_o2;input G3517_o2;input G3533_o2;input G3629_o2;input G3645_o2;input n2497_inv;input G2731_o2;input G2844_o2;input n3732_lo_buf_o2;input n4032_lo_buf_o2;input G3552_o2;input G2271_o2;input n4248_lo_buf_o2;input n4332_lo_buf_o2;input n4344_lo_buf_o2;input n4380_lo_buf_o2;input G2398_o2;input G2480_o2;input G2418_o2;input G1455_o2;input G1449_o2;input G1452_o2;input G1425_o2;input G1428_o2;input G1419_o2;input G1422_o2;input n4308_lo_buf_o2;input G2675_o2;input G3035_o2;input G3026_o2;input G3029_o2;input G3032_o2;input G2999_o2;input G3002_o2;input G2770_o2;input G3008_o2;input G2073_o2;input G2752_o2;input G3005_o2;input G5108_o2;input G5135_o2;input G5111_o2;input G5138_o2;input G3415_o2;input G3386_o2;input G3570_o2;input G2430_o2;input G3495_o2;input G3621_o2;input n4284_lo_buf_o2;input n4356_lo_buf_o2;input G2472_o2;input G2410_o2;input n3960_lo_buf_o2;input n3972_lo_buf_o2;input n2647_inv;input n2650_inv;input n3684_lo_buf_o2;input n4080_lo_buf_o2;input n4092_lo_buf_o2;input n2662_inv;input n2665_inv;input G1147_o2;input G2705_o2;input G2693_o2;input G2696_o2;input G2700_o2;input G2915_o2;input G2966_o2;input G2540_o2;input G2788_o2;input G2792_o2;input G2797_o2;input G2804_o2;input G1038_o2;input G1044_o2;input G1090_o2;input G1096_o2;input G1029_o2;input G3942_o2;input G3954_o2;input G4011_o2;input G4017_o2;input G1141_o2;input G1081_o2;input G2146_o2;input G2145_o2;input G2144_o2;input G2143_o2;input G2142_o2;input G2141_o2;input G2140_o2;input G2139_o2;input G3769_o2;input G3773_o2;input G3768_o2;input G4101_o2;input G3161_o2;input G4143_o2;input G3828_o2;input G3831_o2;input G3334_o2;input G3335_o2;input G3180_o2;input G3340_o2;input G3339_o2;input G3341_o2;input G3234_o2;input G3829_o2;input G3338_o2;input G3336_o2;input G3770_o2;input G3918_o2;input G3774_o2;input G3921_o2;input G3832_o2;input G3993_o2;input G2076_o2;input G2071_o2;input G2072_o2;input G2069_o2;input G2070_o2;input G2067_o2;input G2068_o2;input G4095_o2;input G3272_o2;input G3269_o2;input G3270_o2;input G3271_o2;input G3265_o2;input G3266_o2;input G4137_o2;input G3268_o2;input G2361_o2;input G3228_o2;input G3267_o2;input G2336_o2;input G3459_o2;input G3428_o2;input G3438_o2;input G3449_o2;input G3421_o2;input G3576_o2;input G3303_o2;input G3583_o2;input G3594_o2;input G3674_o2;input G3685_o2;input G4504_o2;input G4180_o2;input G5123_o2;input G5142_o2;input G5126_o2;input G5144_o2;input G3912_o2;input G4417_o2;input G4420_o2;input G3969_o2;input G4023_o2;input G2720_o2;input G2837_o2;input n2965_inv;input n2968_inv;input n2971_inv;input n2974_inv;input G1876_o2;input G4996_o2;input G4984_o2;input G4920_o2;input G4923_o2;input G4930_o2;input G4933_o2;input n4320_lo_buf_o2;input G2424_o2;input G3317_o2;input G3503_o2;input G3485_o2;input G3611_o2;input n3864_lo_buf_o2;input n3888_lo_buf_o2;input n4116_lo_buf_o2;input n4128_lo_buf_o2;input n4140_lo_buf_o2;input n4152_lo_buf_o2;input G1815_o2;input G1728_o2;input G1035_o2;input G1041_o2;input G1087_o2;input G1093_o2;input G1132_o2;input G1108_o2;input G1138_o2;input G1114_o2;input G1807_o2;input G2108_o2;input G1126_o2;input G1899_o2;input G2134_o2;input G1852_o2;input G2116_o2;input G2543_o2;input G2727_o2;input G2715_o2;input G2832_o2;input G1873_o2;input G3291_o2;input G5025_o2;input G5036_o2;input G3132_o2;input G5038_o2;input G5039_o2;input n3118_inv;input n3121_inv;input n3124_inv;input n3127_inv;input n3984_lo_buf_o2;input G1802_o2;input G1804_o2;input G1849_o2;input G1851_o2;input G2492_o2;input G1799_o2;input G4231_o2;input G4234_o2;input G4245_o2;input G4247_o2;input G1894_o2;input G1846_o2;input G4238_o2;input G4249_o2;input G2293_o2;input G5022_o2;input G5006_o2;input G4944_o2;input G4946_o2;input G4954_o2;input G4956_o2;input G3546_o2;input G3658_o2;input G1344_o2;input G2921_o2;input n3912_lo_buf_o2;input G1835_o2;input G3810_o2;input G3866_o2;input G3811_o2;input G2269_o2;input G3812_o2;input G3867_o2;input G3868_o2;input G3809_o2;input G3716_o2;input G4529_o2;input G4670_o2;input G4493_o2;input G4580_o2;input G3822_o2;input G3877_o2;input G4131_o2;input G4170_o2;input G4051_o2;input G4065_o2;input G4697_o2;input G4706_o2;input G2460_o2;input G2454_o2;input G2392_o2;input G2386_o2;input n4260_lo_buf_o2;input n4272_lo_buf_o2;input n4392_lo_buf_o2;input n4404_lo_buf_o2;input G1512_o2;input G3135_o2;input G2379_o2;input n4164_lo_buf_o2;input n4176_lo_buf_o2;input n4224_lo_buf_o2;input G2975_o2;input G2978_o2;input G2933_o2;input G2936_o2;input G1356_o2;input G1359_o2;input G1398_o2;input G1401_o2;
  output G5193;output G5194;output G5195;output G5196;output G5197;output G5198;output G5199;output G5200;output G5201;output G5202;output G5203;output G5204;output G5205;output G5206;output G5207;output G5208;output G5209;output G5210;output G5211;output G5212;output G5213;output G5214;output G5215;output G5216;output G5217;output G5218;output G5219;output G5220;output G5221;output G5222;output G5223;output G5224;output G5225;output G5226;output G5227;output G5228;output G5229;output G5230;output G5231;output G5232;output G5233;output G5234;output G5235;output G5236;output G5237;output G5238;output G5239;output G5240;output G5241;output G5242;output G5243;output G5244;output G5245;output G5246;output G5247;output G5248;output G5249;output G5250;output G5251;output G5252;output G5253;output G5254;output G5255;output G5256;output G5257;output G5258;output G5259;output G5260;output G5261;output G5262;output G5263;output G5264;output G5265;output G5266;output G5267;output G5268;output G5269;output G5270;output G5271;output G5272;output G5273;output G5274;output G5275;output G5276;output G5277;output G5278;output G5279;output G5280;output G5281;output G5282;output G5283;output G5284;output G5285;output G5286;output G5287;output G5288;output G5289;output G5290;output G5291;output G5292;output G5293;output G5294;output G5295;output G5296;output G5297;output G5298;output G5299;output G5300;output G5301;output G5302;output G5303;output G5304;output G5305;output G5306;output G5307;output G5308;output G5309;output G5310;output G5311;output G5312;output G5313;output G5314;output G5315;output n2610_li;output n2613_li;output n2616_li;output n2619_li;output n2622_li;output n2625_li;output n2628_li;output n2631_li;output n2634_li;output n2637_li;output n2640_li;output n2643_li;output n2646_li;output n2649_li;output n2652_li;output n2655_li;output n2658_li;output n2661_li;output n2664_li;output n2667_li;output n2670_li;output n2673_li;output n2676_li;output n2679_li;output n2682_li;output n2685_li;output n2688_li;output n2691_li;output n2694_li;output n2697_li;output n2700_li;output n2703_li;output n2706_li;output n2709_li;output n2712_li;output n2715_li;output n2718_li;output n2721_li;output n2724_li;output n2727_li;output n2730_li;output n2733_li;output n2736_li;output n2739_li;output n2742_li;output n2745_li;output n2748_li;output n2751_li;output n2754_li;output n2757_li;output n2760_li;output n2763_li;output n2766_li;output n2769_li;output n2772_li;output n2775_li;output n2778_li;output n2781_li;output n2784_li;output n2787_li;output n2790_li;output n2793_li;output n2796_li;output n2799_li;output n2802_li;output n2805_li;output n2808_li;output n2811_li;output n2814_li;output n2817_li;output n2820_li;output n2823_li;output n2826_li;output n2829_li;output n2832_li;output n2835_li;output n2838_li;output n2841_li;output n2844_li;output n2847_li;output n2850_li;output n2853_li;output n2856_li;output n2859_li;output n2862_li;output n2865_li;output n2868_li;output n2871_li;output n2874_li;output n2877_li;output n2880_li;output n2883_li;output n2886_li;output n2889_li;output n2892_li;output n2895_li;output n2898_li;output n2901_li;output n2904_li;output n2907_li;output n2910_li;output n2913_li;output n2916_li;output n2919_li;output n2922_li;output n2925_li;output n2928_li;output n2931_li;output n2934_li;output n2937_li;output n2940_li;output n2943_li;output n2946_li;output n2949_li;output n2952_li;output n2955_li;output n2958_li;output n2961_li;output n2964_li;output n2967_li;output n2970_li;output n2973_li;output n2976_li;output n2979_li;output n2982_li;output n2985_li;output n2988_li;output n2991_li;output n2994_li;output n2997_li;output n3000_li;output n3003_li;output n3006_li;output n3009_li;output n3012_li;output n3015_li;output n3018_li;output n3021_li;output n3024_li;output n3027_li;output n3030_li;output n3033_li;output n3036_li;output n3039_li;output n3042_li;output n3045_li;output n3048_li;output n3051_li;output n3054_li;output n3057_li;output n3060_li;output n3063_li;output n3066_li;output n3069_li;output n3072_li;output n3075_li;output n3078_li;output n3081_li;output n3084_li;output n3087_li;output n3090_li;output n3093_li;output n3096_li;output n3099_li;output n3102_li;output n3105_li;output n3108_li;output n3111_li;output n3114_li;output n3117_li;output n3120_li;output n3123_li;output n3126_li;output n3129_li;output n3132_li;output n3135_li;output n3138_li;output n3141_li;output n3144_li;output n3147_li;output n3150_li;output n3153_li;output n3156_li;output n3159_li;output n3162_li;output n3165_li;output n3168_li;output n3171_li;output n3174_li;output n3177_li;output n3180_li;output n3183_li;output n3186_li;output n3189_li;output n3192_li;output n3195_li;output n3198_li;output n3201_li;output n3204_li;output n3207_li;output n3210_li;output n3213_li;output n3216_li;output n3219_li;output n3222_li;output n3225_li;output n3228_li;output n3231_li;output n3234_li;output n3237_li;output n3240_li;output n3243_li;output n3246_li;output n3249_li;output n3252_li;output n3255_li;output n3258_li;output n3261_li;output n3264_li;output n3267_li;output n3270_li;output n3273_li;output n3276_li;output n3279_li;output n3282_li;output n3285_li;output n3288_li;output n3291_li;output n3294_li;output n3297_li;output n3300_li;output n3303_li;output n3306_li;output n3309_li;output n3312_li;output n3315_li;output n3318_li;output n3321_li;output n3324_li;output n3327_li;output n3330_li;output n3333_li;output n3336_li;output n3339_li;output n3342_li;output n3345_li;output n3348_li;output n3351_li;output n3354_li;output n3357_li;output n3360_li;output n3363_li;output n3366_li;output n3369_li;output n3372_li;output n3375_li;output n3378_li;output n3381_li;output n3384_li;output n3387_li;output n3390_li;output n3393_li;output n3396_li;output n3399_li;output n3402_li;output n3405_li;output n3408_li;output n3411_li;output n3414_li;output n3417_li;output n3420_li;output n3423_li;output n3426_li;output n3429_li;output n3432_li;output n3435_li;output n3438_li;output n3441_li;output n3444_li;output n3447_li;output n3450_li;output n3453_li;output n3456_li;output n3459_li;output n3462_li;output n3465_li;output n3468_li;output n3471_li;output n3474_li;output n3477_li;output n3480_li;output n3483_li;output n3486_li;output n3489_li;output n3492_li;output n3495_li;output n3498_li;output n3501_li;output n3504_li;output n3507_li;output n3510_li;output n3513_li;output n3516_li;output n3519_li;output n3522_li;output n3525_li;output n3528_li;output n3531_li;output n3534_li;output n3537_li;output n3540_li;output n3543_li;output n3546_li;output n3549_li;output n3552_li;output n3555_li;output n3558_li;output n3561_li;output n3564_li;output n3567_li;output n3570_li;output n3573_li;output n3576_li;output n3579_li;output n3582_li;output n3585_li;output n3588_li;output n3591_li;output n3594_li;output n3597_li;output n3600_li;output n3603_li;output n3606_li;output n3609_li;output n3612_li;output n3615_li;output n3618_li;output n3621_li;output n3624_li;output n3627_li;output n3630_li;output n3633_li;output n3636_li;output n3639_li;output n3642_li;output n3645_li;output n3648_li;output n3651_li;output n3654_li;output n3657_li;output n3666_li;output n3669_li;output n3678_li;output n3687_li;output n3690_li;output n3702_li;output n3711_li;output n3714_li;output n3726_li;output n3735_li;output n3738_li;output n3750_li;output n3753_li;output n3759_li;output n3762_li;output n3765_li;output n3774_li;output n3777_li;output n3786_li;output n3789_li;output n3792_li;output n3795_li;output n3798_li;output n3801_li;output n3810_li;output n3813_li;output n3822_li;output n3825_li;output n3834_li;output n3843_li;output n3846_li;output n3867_li;output n3891_li;output n3915_li;output n3930_li;output n3933_li;output n3936_li;output n3942_li;output n3945_li;output n3948_li;output n3954_li;output n3957_li;output n3963_li;output n3966_li;output n3969_li;output n3975_li;output n3978_li;output n3987_li;output n3990_li;output n4002_li;output n4011_li;output n4014_li;output n4026_li;output n4035_li;output n4038_li;output n4050_li;output n4053_li;output n4059_li;output n4062_li;output n4065_li;output n4098_li;output n4107_li;output n4119_li;output n4131_li;output n4143_li;output n4155_li;output n4167_li;output n4179_li;output n4182_li;output n4185_li;output n4188_li;output n4194_li;output n4197_li;output n4200_li;output n4206_li;output n4209_li;output n4212_li;output n4215_li;output n4227_li;output n4230_li;output n4233_li;output n4236_li;output n4239_li;output n4242_li;output n4251_li;output n4263_li;output n4275_li;output n4278_li;output n4287_li;output n4290_li;output n4293_li;output n4299_li;output n4302_li;output n4305_li;output n4311_li;output n4314_li;output n4323_li;output n4326_li;output n4335_li;output n4338_li;output n4347_li;output n4350_li;output n4359_li;output n4362_li;output n4365_li;output n4371_li;output n4374_li;output n4383_li;output n4395_li;output n4407_li;output n4410_li;output n4413_li;output n4416_li;output n4419_li;output n4422_li;output n4425_li;output n4428_li;output n4431_li;output n4434_li;output n4437_li;output n4440_li;output n4443_li;output n4446_li;output n4449_li;output n4452_li;output n4455_li;output n4458_li;output n4461_li;output n4464_li;output n4467_li;output n4470_li;output n4473_li;output n4476_li;output n4479_li;output n4482_li;output n4485_li;output n4488_li;output n4494_li;output n4497_li;output n4500_li;output n4503_li;output n4506_li;output n4509_li;output n4512_li;output n4515_li;output n4518_li;output n4521_li;output n4524_li;output n4527_li;output n4530_li;output n4533_li;output n4536_li;output n4539_li;output n4542_li;output n4545_li;output n4548_li;output n4554_li;output n4557_li;output n4560_li;output n4563_li;output n4566_li;output n4569_li;output n4572_li;output n4575_li;output n4578_li;output n4581_li;output n4584_li;output n4587_li;output n4590_li;output n4593_li;output n4596_li;output n4599_li;output n4602_li;output n4605_li;output n4608_li;output n4611_li;output n4614_li;output n4617_li;output n4620_li;output n4623_li;output n4626_li;output n4629_li;output n4632_li;output n4635_li;output n4638_li;output n4641_li;output n4644_li;output n4647_li;output n4650_li;output n4653_li;output n4656_li;output n4659_li;output n4662_li;output n4665_li;output n4668_li;output n4671_li;output n4674_li;output n4677_li;output n4680_li;output n4683_li;output n4686_li;output n4689_li;output n4692_li;output n4695_li;output n4698_li;output n4701_li;output n4704_li;output n4707_li;output n4710_li;output n4713_li;output n4716_li;output n4719_li;output n4722_li;output n4725_li;output n4728_li;output n4731_li;output n4734_li;output n4737_li;output n4740_li;output n4743_li;output n6382_i2;output n6383_i2;output n6419_i2;output n6420_i2;output n6435_i2;output n6436_i2;output n6448_i2;output n6449_i2;output n6613_i2;output n6614_i2;output n6641_i2;output n6658_i2;output n6757_i2;output n6756_i2;output n7116_i2;output n7156_i2;output n6549_i2;output n6550_i2;output n7357_i2;output n7358_i2;output n7359_i2;output n7360_i2;output n6621_i2;output n6623_i2;output n6625_i2;output n6626_i2;output n6627_i2;output n6628_i2;output n6629_i2;output n6630_i2;output n6669_i2;output n7449_i2;output n7450_i2;output n7451_i2;output n7452_i2;output n6682_i2;output n6683_i2;output n6684_i2;output n6685_i2;output n7463_i2;output n6686_i2;output n6687_i2;output n6688_i2;output n6689_i2;output n6772_i2;output n6773_i2;output n6774_i2;output n6775_i2;output G3467_i2;output G2810_i2;output n6833_i2;output n6945_i2;output n6947_i2;output n6949_i2;output n6951_i2;output n6888_i2;output n6889_i2;output n6936_i2;output n6954_i2;output n6955_i2;output n6956_i2;output n6957_i2;output n6958_i2;output n6982_i2;output n6984_i2;output n6974_i2;output n6975_i2;output n6999_i2;output n7015_i2;output n7016_i2;output n7017_i2;output n7018_i2;output n7005_i2;output n7019_i2;output n7022_i2;output n7023_i2;output n7132_i2;output n7133_i2;output n7135_i2;output n7136_i2;output n7175_i2;output n7155_i2;output G3060_i2;output n7383_i2;output G3802_i2;output G3859_i2;output n7355_i2;output n7356_i2;output G4054_i2;output G4068_i2;output n7384_i2;output n7387_i2;output n7388_i2;output n7389_i2;output n7386_i2;output n7453_i2;output n7431_i2;output n7432_i2;output n7433_i2;output n7430_i2;output n7485_i2;output n7486_i2;output G2508_i2;output G2486_i2;output n7245_i2;output n7246_i2;output n3756_lo_buf_i2;output n4056_lo_buf_i2;output G3474_i2;output G2817_i2;output n7396_i2;output n7398_i2;output n7400_i2;output n7401_i2;output n7402_i2;output n7403_i2;output n7404_i2;output n7405_i2;output G2711_i2;output G2828_i2;output n7490_i2;output n7527_i2;output n7528_i2;output n7529_i2;output n7530_i2;output n7523_i2;output n7524_i2;output n7525_i2;output n7526_i2;output n4296_lo_buf_i2;output n4368_lo_buf_i2;output G2466_i2;output G2404_i2;output n7534_i2;output n7535_i2;output n7536_i2;output n7533_i2;output G1060_i2;output G963_i2;output G2448_i2;output G2685_i2;output G2679_i2;output G2774_i2;output G2780_i2;output G2759_i2;output G2737_i2;output G2850_i2;output G3393_i2;output G3404_i2;output G3559_i2;output G2744_i2;output n3708_lo_buf_i2;output n3840_lo_buf_i2;output n4008_lo_buf_i2;output n4104_lo_buf_i2;output G1821_i2;output G1734_i2;output G3517_i2;output G3533_i2;output G3629_i2;output G3645_i2;output G2857_i2;output G2731_i2;output G2844_i2;output n3732_lo_buf_i2;output n4032_lo_buf_i2;output G3552_i2;output G2271_i2;output n4248_lo_buf_i2;output n4332_lo_buf_i2;output n4344_lo_buf_i2;output n4380_lo_buf_i2;output G2398_i2;output G2480_i2;output G2418_i2;output G1455_i2;output G1449_i2;output G1452_i2;output G1425_i2;output G1428_i2;output G1419_i2;output G1422_i2;output n4308_lo_buf_i2;output G2675_i2;output G3035_i2;output G3026_i2;output G3029_i2;output G3032_i2;output G2999_i2;output G3002_i2;output G2770_i2;output G3008_i2;output G2073_i2;output G2752_i2;output G3005_i2;output G5108_i2;output G5135_i2;output G5111_i2;output G5138_i2;output G3415_i2;output G3386_i2;output G3570_i2;output G2430_i2;output G3495_i2;output G3621_i2;output n4284_lo_buf_i2;output n4356_lo_buf_i2;output G2472_i2;output G2410_i2;output n3960_lo_buf_i2;output n3972_lo_buf_i2;output G2865_i2;output G970_i2;output n3684_lo_buf_i2;output n4080_lo_buf_i2;output n4092_lo_buf_i2;output G1053_i2;output G956_i2;output G1147_i2;output G2705_i2;output G2693_i2;output G2696_i2;output G2700_i2;output G2915_i2;output G2966_i2;output G2540_i2;output G2788_i2;output G2792_i2;output G2797_i2;output G2804_i2;output G1038_i2;output G1044_i2;output G1090_i2;output G1096_i2;output G1029_i2;output G3942_i2;output G3954_i2;output G4011_i2;output G4017_i2;output G1141_i2;output G1081_i2;output G2146_i2;output G2145_i2;output G2144_i2;output G2143_i2;output G2142_i2;output G2141_i2;output G2140_i2;output G2139_i2;output G3769_i2;output G3773_i2;output G3768_i2;output G4101_i2;output G3161_i2;output G4143_i2;output G3828_i2;output G3831_i2;output G3334_i2;output G3335_i2;output G3180_i2;output G3340_i2;output G3339_i2;output G3341_i2;output G3234_i2;output G3829_i2;output G3338_i2;output G3336_i2;output G3770_i2;output G3918_i2;output G3774_i2;output G3921_i2;output G3832_i2;output G3993_i2;output G2076_i2;output G2071_i2;output G2072_i2;output G2069_i2;output G2070_i2;output G2067_i2;output G2068_i2;output G4095_i2;output G3272_i2;output G3269_i2;output G3270_i2;output G3271_i2;output G3265_i2;output G3266_i2;output G4137_i2;output G3268_i2;output G2361_i2;output G3228_i2;output G3267_i2;output G2336_i2;output G3459_i2;output G3428_i2;output G3438_i2;output G3449_i2;output G3421_i2;output G3576_i2;output G3303_i2;output G3583_i2;output G3594_i2;output G3674_i2;output G3685_i2;output G4504_i2;output G4180_i2;output G5123_i2;output G5142_i2;output G5126_i2;output G5144_i2;output G3912_i2;output G4417_i2;output G4420_i2;output G3969_i2;output G4023_i2;output G2720_i2;output G2837_i2;output G836_i2;output G848_i2;output G813_i2;output G825_i2;output G1876_i2;output G4996_i2;output G4984_i2;output G4920_i2;output G4923_i2;output G4930_i2;output G4933_i2;output n4320_lo_buf_i2;output G2424_i2;output G3317_i2;output G3503_i2;output G3485_i2;output G3611_i2;output n3864_lo_buf_i2;output n3888_lo_buf_i2;output n4116_lo_buf_i2;output n4128_lo_buf_i2;output n4140_lo_buf_i2;output n4152_lo_buf_i2;output G1815_i2;output G1728_i2;output G1035_i2;output G1041_i2;output G1087_i2;output G1093_i2;output G1132_i2;output G1108_i2;output G1138_i2;output G1114_i2;output G1807_i2;output G2108_i2;output G1126_i2;output G1899_i2;output G2134_i2;output G1852_i2;output G2116_i2;output G2543_i2;output G2727_i2;output G2715_i2;output G2832_i2;output G1873_i2;output G3291_i2;output G5025_i2;output G5036_i2;output G3132_i2;output G5038_i2;output G5039_i2;output G1150_i2;output G1162_i2;output G804_i2;output G1172_i2;output n3984_lo_buf_i2;output G1802_i2;output G1804_i2;output G1849_i2;output G1851_i2;output G2492_i2;output G1799_i2;output G4231_i2;output G4234_i2;output G4245_i2;output G4247_i2;output G1894_i2;output G1846_i2;output G4238_i2;output G4249_i2;output G2293_i2;output G5022_i2;output G5006_i2;output G4944_i2;output G4946_i2;output G4954_i2;output G4956_i2;output G3546_i2;output G3658_i2;output G1344_i2;output G2921_i2;output n3912_lo_buf_i2;output G1835_i2;output G3810_i2;output G3866_i2;output G3811_i2;output G2269_i2;output G3812_i2;output G3867_i2;output G3868_i2;output G3809_i2;output G3716_i2;output G4529_i2;output G4670_i2;output G4493_i2;output G4580_i2;output G3822_i2;output G3877_i2;output G4131_i2;output G4170_i2;output G4051_i2;output G4065_i2;output G4697_i2;output G4706_i2;output G2460_i2;output G2454_i2;output G2392_i2;output G2386_i2;output n4260_lo_buf_i2;output n4272_lo_buf_i2;output n4392_lo_buf_i2;output n4404_lo_buf_i2;output G1512_i2;output G3135_i2;output G2379_i2;output n4164_lo_buf_i2;output n4176_lo_buf_i2;output n4224_lo_buf_i2;output G2975_i2;output G2978_i2;output G2933_i2;output G2936_i2;output G1356_i2;output G1359_i2;output G1398_i2;output G1401_i2;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire G51_p;
  wire G51_n;
  wire G52_p;
  wire G52_n;
  wire G53_p;
  wire G53_n;
  wire G54_p;
  wire G54_n;
  wire G55_p;
  wire G55_n;
  wire G56_p;
  wire G56_n;
  wire G57_p;
  wire G57_n;
  wire G58_p;
  wire G58_n;
  wire G59_p;
  wire G59_n;
  wire G60_p;
  wire G60_n;
  wire G61_p;
  wire G61_n;
  wire G62_p;
  wire G62_n;
  wire G63_p;
  wire G63_n;
  wire G64_p;
  wire G64_n;
  wire G65_p;
  wire G65_n;
  wire G66_p;
  wire G66_n;
  wire G67_p;
  wire G67_n;
  wire G68_p;
  wire G68_n;
  wire G69_p;
  wire G69_n;
  wire G70_p;
  wire G70_n;
  wire G71_p;
  wire G71_n;
  wire G72_p;
  wire G72_n;
  wire G73_p;
  wire G73_n;
  wire G74_p;
  wire G74_n;
  wire G75_p;
  wire G75_n;
  wire G76_p;
  wire G76_n;
  wire G77_p;
  wire G77_n;
  wire G78_p;
  wire G78_n;
  wire G79_p;
  wire G79_n;
  wire G80_p;
  wire G80_n;
  wire G81_p;
  wire G81_n;
  wire G82_p;
  wire G82_n;
  wire G83_p;
  wire G83_n;
  wire G84_p;
  wire G84_n;
  wire G85_p;
  wire G85_n;
  wire G86_p;
  wire G86_n;
  wire G87_p;
  wire G87_n;
  wire G88_p;
  wire G88_n;
  wire G89_p;
  wire G89_n;
  wire G90_p;
  wire G90_n;
  wire G91_p;
  wire G91_n;
  wire G92_p;
  wire G92_n;
  wire G93_p;
  wire G93_n;
  wire G94_p;
  wire G94_n;
  wire G95_p;
  wire G95_n;
  wire G96_p;
  wire G96_n;
  wire G97_p;
  wire G97_n;
  wire G98_p;
  wire G98_n;
  wire G99_p;
  wire G99_n;
  wire G100_p;
  wire G100_n;
  wire G101_p;
  wire G101_n;
  wire G102_p;
  wire G102_n;
  wire G103_p;
  wire G103_n;
  wire G104_p;
  wire G104_n;
  wire G105_p;
  wire G105_n;
  wire G106_p;
  wire G106_n;
  wire G107_p;
  wire G107_n;
  wire G108_p;
  wire G108_n;
  wire G109_p;
  wire G109_n;
  wire G110_p;
  wire G110_n;
  wire G111_p;
  wire G111_n;
  wire G112_p;
  wire G112_n;
  wire G113_p;
  wire G113_n;
  wire G114_p;
  wire G114_n;
  wire G115_p;
  wire G115_n;
  wire G116_p;
  wire G116_n;
  wire G117_p;
  wire G117_n;
  wire G118_p;
  wire G118_n;
  wire G119_p;
  wire G119_n;
  wire G120_p;
  wire G120_n;
  wire G121_p;
  wire G121_n;
  wire G122_p;
  wire G122_n;
  wire G123_p;
  wire G123_n;
  wire G124_p;
  wire G124_n;
  wire G125_p;
  wire G125_n;
  wire G126_p;
  wire G126_n;
  wire G127_p;
  wire G127_n;
  wire G128_p;
  wire G128_n;
  wire G129_p;
  wire G129_n;
  wire G130_p;
  wire G130_n;
  wire G131_p;
  wire G131_n;
  wire G132_p;
  wire G132_n;
  wire G133_p;
  wire G133_n;
  wire G134_p;
  wire G134_n;
  wire G135_p;
  wire G135_n;
  wire G136_p;
  wire G136_n;
  wire G137_p;
  wire G137_n;
  wire G138_p;
  wire G138_n;
  wire G139_p;
  wire G139_n;
  wire G140_p;
  wire G140_n;
  wire G141_p;
  wire G141_n;
  wire G142_p;
  wire G142_n;
  wire G143_p;
  wire G143_n;
  wire G144_p;
  wire G144_n;
  wire G145_p;
  wire G145_n;
  wire G146_p;
  wire G146_n;
  wire G147_p;
  wire G147_n;
  wire G148_p;
  wire G148_n;
  wire G149_p;
  wire G149_n;
  wire G150_p;
  wire G150_n;
  wire G151_p;
  wire G151_n;
  wire G152_p;
  wire G152_n;
  wire G153_p;
  wire G153_n;
  wire G154_p;
  wire G154_n;
  wire G155_p;
  wire G155_n;
  wire G156_p;
  wire G156_n;
  wire G157_p;
  wire G157_n;
  wire G158_p;
  wire G158_n;
  wire G159_p;
  wire G159_n;
  wire G160_p;
  wire G160_n;
  wire G161_p;
  wire G161_n;
  wire G162_p;
  wire G162_n;
  wire G163_p;
  wire G163_n;
  wire G164_p;
  wire G164_n;
  wire G165_p;
  wire G165_n;
  wire G166_p;
  wire G166_n;
  wire G167_p;
  wire G167_n;
  wire G168_p;
  wire G168_n;
  wire G169_p;
  wire G169_n;
  wire G170_p;
  wire G170_n;
  wire G171_p;
  wire G171_n;
  wire G172_p;
  wire G172_n;
  wire G173_p;
  wire G173_n;
  wire G174_p;
  wire G174_n;
  wire G175_p;
  wire G175_n;
  wire G176_p;
  wire G176_n;
  wire G177_p;
  wire G177_n;
  wire G178_p;
  wire G178_n;
  wire n2610_lo_p;
  wire n2610_lo_n;
  wire n2613_lo_p;
  wire n2613_lo_n;
  wire n2616_lo_p;
  wire n2616_lo_n;
  wire n2619_lo_p;
  wire n2619_lo_n;
  wire n2622_lo_p;
  wire n2622_lo_n;
  wire n2625_lo_p;
  wire n2625_lo_n;
  wire n2628_lo_p;
  wire n2628_lo_n;
  wire n2631_lo_p;
  wire n2631_lo_n;
  wire n2634_lo_p;
  wire n2634_lo_n;
  wire n2637_lo_p;
  wire n2637_lo_n;
  wire n2640_lo_p;
  wire n2640_lo_n;
  wire n2643_lo_p;
  wire n2643_lo_n;
  wire n2646_lo_p;
  wire n2646_lo_n;
  wire n2649_lo_p;
  wire n2649_lo_n;
  wire n2652_lo_p;
  wire n2652_lo_n;
  wire n2655_lo_p;
  wire n2655_lo_n;
  wire n2658_lo_p;
  wire n2658_lo_n;
  wire n2661_lo_p;
  wire n2661_lo_n;
  wire n2664_lo_p;
  wire n2664_lo_n;
  wire n2667_lo_p;
  wire n2667_lo_n;
  wire n2670_lo_p;
  wire n2670_lo_n;
  wire n2673_lo_p;
  wire n2673_lo_n;
  wire n2676_lo_p;
  wire n2676_lo_n;
  wire n2679_lo_p;
  wire n2679_lo_n;
  wire n2682_lo_p;
  wire n2682_lo_n;
  wire n2685_lo_p;
  wire n2685_lo_n;
  wire n2688_lo_p;
  wire n2688_lo_n;
  wire n2691_lo_p;
  wire n2691_lo_n;
  wire n2694_lo_p;
  wire n2694_lo_n;
  wire n2697_lo_p;
  wire n2697_lo_n;
  wire n2700_lo_p;
  wire n2700_lo_n;
  wire n2703_lo_p;
  wire n2703_lo_n;
  wire n2706_lo_p;
  wire n2706_lo_n;
  wire n2709_lo_p;
  wire n2709_lo_n;
  wire n2712_lo_p;
  wire n2712_lo_n;
  wire n2715_lo_p;
  wire n2715_lo_n;
  wire n2718_lo_p;
  wire n2718_lo_n;
  wire n2721_lo_p;
  wire n2721_lo_n;
  wire n2724_lo_p;
  wire n2724_lo_n;
  wire n2727_lo_p;
  wire n2727_lo_n;
  wire n2730_lo_p;
  wire n2730_lo_n;
  wire n2733_lo_p;
  wire n2733_lo_n;
  wire n2736_lo_p;
  wire n2736_lo_n;
  wire n2739_lo_p;
  wire n2739_lo_n;
  wire n2742_lo_p;
  wire n2742_lo_n;
  wire n2745_lo_p;
  wire n2745_lo_n;
  wire n2748_lo_p;
  wire n2748_lo_n;
  wire n2751_lo_p;
  wire n2751_lo_n;
  wire n2754_lo_p;
  wire n2754_lo_n;
  wire n2757_lo_p;
  wire n2757_lo_n;
  wire n2760_lo_p;
  wire n2760_lo_n;
  wire n2763_lo_p;
  wire n2763_lo_n;
  wire n2766_lo_p;
  wire n2766_lo_n;
  wire n2769_lo_p;
  wire n2769_lo_n;
  wire n2772_lo_p;
  wire n2772_lo_n;
  wire n2775_lo_p;
  wire n2775_lo_n;
  wire n2778_lo_p;
  wire n2778_lo_n;
  wire n2781_lo_p;
  wire n2781_lo_n;
  wire n2784_lo_p;
  wire n2784_lo_n;
  wire n2787_lo_p;
  wire n2787_lo_n;
  wire n2790_lo_p;
  wire n2790_lo_n;
  wire n2793_lo_p;
  wire n2793_lo_n;
  wire n2796_lo_p;
  wire n2796_lo_n;
  wire n2799_lo_p;
  wire n2799_lo_n;
  wire n2802_lo_p;
  wire n2802_lo_n;
  wire n2805_lo_p;
  wire n2805_lo_n;
  wire n2808_lo_p;
  wire n2808_lo_n;
  wire n2811_lo_p;
  wire n2811_lo_n;
  wire n2814_lo_p;
  wire n2814_lo_n;
  wire n2817_lo_p;
  wire n2817_lo_n;
  wire n2820_lo_p;
  wire n2820_lo_n;
  wire n2823_lo_p;
  wire n2823_lo_n;
  wire n2826_lo_p;
  wire n2826_lo_n;
  wire n2829_lo_p;
  wire n2829_lo_n;
  wire n2832_lo_p;
  wire n2832_lo_n;
  wire n2835_lo_p;
  wire n2835_lo_n;
  wire n2838_lo_p;
  wire n2838_lo_n;
  wire n2841_lo_p;
  wire n2841_lo_n;
  wire n2844_lo_p;
  wire n2844_lo_n;
  wire n2847_lo_p;
  wire n2847_lo_n;
  wire n2850_lo_p;
  wire n2850_lo_n;
  wire n2853_lo_p;
  wire n2853_lo_n;
  wire n2856_lo_p;
  wire n2856_lo_n;
  wire n2859_lo_p;
  wire n2859_lo_n;
  wire n2862_lo_p;
  wire n2862_lo_n;
  wire n2865_lo_p;
  wire n2865_lo_n;
  wire n2868_lo_p;
  wire n2868_lo_n;
  wire n2871_lo_p;
  wire n2871_lo_n;
  wire n2874_lo_p;
  wire n2874_lo_n;
  wire n2877_lo_p;
  wire n2877_lo_n;
  wire n2880_lo_p;
  wire n2880_lo_n;
  wire n2883_lo_p;
  wire n2883_lo_n;
  wire n2886_lo_p;
  wire n2886_lo_n;
  wire n2889_lo_p;
  wire n2889_lo_n;
  wire n2892_lo_p;
  wire n2892_lo_n;
  wire n2895_lo_p;
  wire n2895_lo_n;
  wire n2898_lo_p;
  wire n2898_lo_n;
  wire n2901_lo_p;
  wire n2901_lo_n;
  wire n2904_lo_p;
  wire n2904_lo_n;
  wire n2907_lo_p;
  wire n2907_lo_n;
  wire n2910_lo_p;
  wire n2910_lo_n;
  wire n2913_lo_p;
  wire n2913_lo_n;
  wire n2916_lo_p;
  wire n2916_lo_n;
  wire n2919_lo_p;
  wire n2919_lo_n;
  wire n2922_lo_p;
  wire n2922_lo_n;
  wire n2925_lo_p;
  wire n2925_lo_n;
  wire n2928_lo_p;
  wire n2928_lo_n;
  wire n2931_lo_p;
  wire n2931_lo_n;
  wire n2934_lo_p;
  wire n2934_lo_n;
  wire n2937_lo_p;
  wire n2937_lo_n;
  wire n2940_lo_p;
  wire n2940_lo_n;
  wire n2943_lo_p;
  wire n2943_lo_n;
  wire n2946_lo_p;
  wire n2946_lo_n;
  wire n2949_lo_p;
  wire n2949_lo_n;
  wire n2952_lo_p;
  wire n2952_lo_n;
  wire n2955_lo_p;
  wire n2955_lo_n;
  wire n2958_lo_p;
  wire n2958_lo_n;
  wire n2961_lo_p;
  wire n2961_lo_n;
  wire n2964_lo_p;
  wire n2964_lo_n;
  wire n2967_lo_p;
  wire n2967_lo_n;
  wire n2970_lo_p;
  wire n2970_lo_n;
  wire n2973_lo_p;
  wire n2973_lo_n;
  wire n2976_lo_p;
  wire n2976_lo_n;
  wire n2979_lo_p;
  wire n2979_lo_n;
  wire n2982_lo_p;
  wire n2982_lo_n;
  wire n2985_lo_p;
  wire n2985_lo_n;
  wire n2988_lo_p;
  wire n2988_lo_n;
  wire n2991_lo_p;
  wire n2991_lo_n;
  wire n2994_lo_p;
  wire n2994_lo_n;
  wire n2997_lo_p;
  wire n2997_lo_n;
  wire n3000_lo_p;
  wire n3000_lo_n;
  wire n3003_lo_p;
  wire n3003_lo_n;
  wire n3006_lo_p;
  wire n3006_lo_n;
  wire n3009_lo_p;
  wire n3009_lo_n;
  wire n3012_lo_p;
  wire n3012_lo_n;
  wire n3015_lo_p;
  wire n3015_lo_n;
  wire n3018_lo_p;
  wire n3018_lo_n;
  wire n3021_lo_p;
  wire n3021_lo_n;
  wire n3024_lo_p;
  wire n3024_lo_n;
  wire n3027_lo_p;
  wire n3027_lo_n;
  wire n3030_lo_p;
  wire n3030_lo_n;
  wire n3033_lo_p;
  wire n3033_lo_n;
  wire n3036_lo_p;
  wire n3036_lo_n;
  wire n3039_lo_p;
  wire n3039_lo_n;
  wire n3042_lo_p;
  wire n3042_lo_n;
  wire n3045_lo_p;
  wire n3045_lo_n;
  wire n3048_lo_p;
  wire n3048_lo_n;
  wire n3051_lo_p;
  wire n3051_lo_n;
  wire n3054_lo_p;
  wire n3054_lo_n;
  wire n3057_lo_p;
  wire n3057_lo_n;
  wire n3060_lo_p;
  wire n3060_lo_n;
  wire n3063_lo_p;
  wire n3063_lo_n;
  wire n3066_lo_p;
  wire n3066_lo_n;
  wire n3069_lo_p;
  wire n3069_lo_n;
  wire n3072_lo_p;
  wire n3072_lo_n;
  wire n3075_lo_p;
  wire n3075_lo_n;
  wire n3078_lo_p;
  wire n3078_lo_n;
  wire n3081_lo_p;
  wire n3081_lo_n;
  wire n3084_lo_p;
  wire n3084_lo_n;
  wire n3087_lo_p;
  wire n3087_lo_n;
  wire n3090_lo_p;
  wire n3090_lo_n;
  wire n3093_lo_p;
  wire n3093_lo_n;
  wire n3096_lo_p;
  wire n3096_lo_n;
  wire n3099_lo_p;
  wire n3099_lo_n;
  wire n3102_lo_p;
  wire n3102_lo_n;
  wire n3105_lo_p;
  wire n3105_lo_n;
  wire n3108_lo_p;
  wire n3108_lo_n;
  wire n3111_lo_p;
  wire n3111_lo_n;
  wire n3114_lo_p;
  wire n3114_lo_n;
  wire n3117_lo_p;
  wire n3117_lo_n;
  wire n3120_lo_p;
  wire n3120_lo_n;
  wire n3123_lo_p;
  wire n3123_lo_n;
  wire n3126_lo_p;
  wire n3126_lo_n;
  wire n3129_lo_p;
  wire n3129_lo_n;
  wire n3132_lo_p;
  wire n3132_lo_n;
  wire n3135_lo_p;
  wire n3135_lo_n;
  wire n3138_lo_p;
  wire n3138_lo_n;
  wire n3141_lo_p;
  wire n3141_lo_n;
  wire n3144_lo_p;
  wire n3144_lo_n;
  wire n3147_lo_p;
  wire n3147_lo_n;
  wire n3150_lo_p;
  wire n3150_lo_n;
  wire n3153_lo_p;
  wire n3153_lo_n;
  wire n3156_lo_p;
  wire n3156_lo_n;
  wire n3159_lo_p;
  wire n3159_lo_n;
  wire n3162_lo_p;
  wire n3162_lo_n;
  wire n3165_lo_p;
  wire n3165_lo_n;
  wire n3168_lo_p;
  wire n3168_lo_n;
  wire n3171_lo_p;
  wire n3171_lo_n;
  wire n3174_lo_p;
  wire n3174_lo_n;
  wire n3177_lo_p;
  wire n3177_lo_n;
  wire n3180_lo_p;
  wire n3180_lo_n;
  wire n3183_lo_p;
  wire n3183_lo_n;
  wire n3186_lo_p;
  wire n3186_lo_n;
  wire n3189_lo_p;
  wire n3189_lo_n;
  wire n3192_lo_p;
  wire n3192_lo_n;
  wire n3195_lo_p;
  wire n3195_lo_n;
  wire n3198_lo_p;
  wire n3198_lo_n;
  wire n3201_lo_p;
  wire n3201_lo_n;
  wire n3204_lo_p;
  wire n3204_lo_n;
  wire n3207_lo_p;
  wire n3207_lo_n;
  wire n3210_lo_p;
  wire n3210_lo_n;
  wire n3213_lo_p;
  wire n3213_lo_n;
  wire n3216_lo_p;
  wire n3216_lo_n;
  wire n3219_lo_p;
  wire n3219_lo_n;
  wire n3222_lo_p;
  wire n3222_lo_n;
  wire n3225_lo_p;
  wire n3225_lo_n;
  wire n3228_lo_p;
  wire n3228_lo_n;
  wire n3231_lo_p;
  wire n3231_lo_n;
  wire n3234_lo_p;
  wire n3234_lo_n;
  wire n3237_lo_p;
  wire n3237_lo_n;
  wire n3240_lo_p;
  wire n3240_lo_n;
  wire n3243_lo_p;
  wire n3243_lo_n;
  wire n3246_lo_p;
  wire n3246_lo_n;
  wire n3249_lo_p;
  wire n3249_lo_n;
  wire n3252_lo_p;
  wire n3252_lo_n;
  wire n3255_lo_p;
  wire n3255_lo_n;
  wire n3258_lo_p;
  wire n3258_lo_n;
  wire n3261_lo_p;
  wire n3261_lo_n;
  wire n3264_lo_p;
  wire n3264_lo_n;
  wire n3267_lo_p;
  wire n3267_lo_n;
  wire n3270_lo_p;
  wire n3270_lo_n;
  wire n3273_lo_p;
  wire n3273_lo_n;
  wire n3276_lo_p;
  wire n3276_lo_n;
  wire n3279_lo_p;
  wire n3279_lo_n;
  wire n3282_lo_p;
  wire n3282_lo_n;
  wire n3285_lo_p;
  wire n3285_lo_n;
  wire n3288_lo_p;
  wire n3288_lo_n;
  wire n3291_lo_p;
  wire n3291_lo_n;
  wire n3294_lo_p;
  wire n3294_lo_n;
  wire n3297_lo_p;
  wire n3297_lo_n;
  wire n3300_lo_p;
  wire n3300_lo_n;
  wire n3303_lo_p;
  wire n3303_lo_n;
  wire n3306_lo_p;
  wire n3306_lo_n;
  wire n3309_lo_p;
  wire n3309_lo_n;
  wire n3312_lo_p;
  wire n3312_lo_n;
  wire n3315_lo_p;
  wire n3315_lo_n;
  wire n3318_lo_p;
  wire n3318_lo_n;
  wire n3321_lo_p;
  wire n3321_lo_n;
  wire n3324_lo_p;
  wire n3324_lo_n;
  wire n3327_lo_p;
  wire n3327_lo_n;
  wire n3330_lo_p;
  wire n3330_lo_n;
  wire n3333_lo_p;
  wire n3333_lo_n;
  wire n3336_lo_p;
  wire n3336_lo_n;
  wire n3339_lo_p;
  wire n3339_lo_n;
  wire n3342_lo_p;
  wire n3342_lo_n;
  wire n3345_lo_p;
  wire n3345_lo_n;
  wire n3348_lo_p;
  wire n3348_lo_n;
  wire n3351_lo_p;
  wire n3351_lo_n;
  wire n3354_lo_p;
  wire n3354_lo_n;
  wire n3357_lo_p;
  wire n3357_lo_n;
  wire n3360_lo_p;
  wire n3360_lo_n;
  wire n3363_lo_p;
  wire n3363_lo_n;
  wire n3366_lo_p;
  wire n3366_lo_n;
  wire n3369_lo_p;
  wire n3369_lo_n;
  wire n3372_lo_p;
  wire n3372_lo_n;
  wire n3375_lo_p;
  wire n3375_lo_n;
  wire n3378_lo_p;
  wire n3378_lo_n;
  wire n3381_lo_p;
  wire n3381_lo_n;
  wire n3384_lo_p;
  wire n3384_lo_n;
  wire n3387_lo_p;
  wire n3387_lo_n;
  wire n3390_lo_p;
  wire n3390_lo_n;
  wire n3393_lo_p;
  wire n3393_lo_n;
  wire n3396_lo_p;
  wire n3396_lo_n;
  wire n3399_lo_p;
  wire n3399_lo_n;
  wire n3402_lo_p;
  wire n3402_lo_n;
  wire n3405_lo_p;
  wire n3405_lo_n;
  wire n3408_lo_p;
  wire n3408_lo_n;
  wire n3411_lo_p;
  wire n3411_lo_n;
  wire n3414_lo_p;
  wire n3414_lo_n;
  wire n3417_lo_p;
  wire n3417_lo_n;
  wire n3420_lo_p;
  wire n3420_lo_n;
  wire n3423_lo_p;
  wire n3423_lo_n;
  wire n3426_lo_p;
  wire n3426_lo_n;
  wire n3429_lo_p;
  wire n3429_lo_n;
  wire n3432_lo_p;
  wire n3432_lo_n;
  wire n3435_lo_p;
  wire n3435_lo_n;
  wire n3438_lo_p;
  wire n3438_lo_n;
  wire n3441_lo_p;
  wire n3441_lo_n;
  wire n3444_lo_p;
  wire n3444_lo_n;
  wire n3447_lo_p;
  wire n3447_lo_n;
  wire n3450_lo_p;
  wire n3450_lo_n;
  wire n3453_lo_p;
  wire n3453_lo_n;
  wire n3456_lo_p;
  wire n3456_lo_n;
  wire n3459_lo_p;
  wire n3459_lo_n;
  wire n3462_lo_p;
  wire n3462_lo_n;
  wire n3465_lo_p;
  wire n3465_lo_n;
  wire n3468_lo_p;
  wire n3468_lo_n;
  wire n3471_lo_p;
  wire n3471_lo_n;
  wire n3474_lo_p;
  wire n3474_lo_n;
  wire n3477_lo_p;
  wire n3477_lo_n;
  wire n3480_lo_p;
  wire n3480_lo_n;
  wire n3483_lo_p;
  wire n3483_lo_n;
  wire n3486_lo_p;
  wire n3486_lo_n;
  wire n3489_lo_p;
  wire n3489_lo_n;
  wire n3492_lo_p;
  wire n3492_lo_n;
  wire n3495_lo_p;
  wire n3495_lo_n;
  wire n3498_lo_p;
  wire n3498_lo_n;
  wire n3501_lo_p;
  wire n3501_lo_n;
  wire n3504_lo_p;
  wire n3504_lo_n;
  wire n3507_lo_p;
  wire n3507_lo_n;
  wire n3510_lo_p;
  wire n3510_lo_n;
  wire n3513_lo_p;
  wire n3513_lo_n;
  wire n3516_lo_p;
  wire n3516_lo_n;
  wire n3519_lo_p;
  wire n3519_lo_n;
  wire n3522_lo_p;
  wire n3522_lo_n;
  wire n3525_lo_p;
  wire n3525_lo_n;
  wire n3528_lo_p;
  wire n3528_lo_n;
  wire n3531_lo_p;
  wire n3531_lo_n;
  wire n3534_lo_p;
  wire n3534_lo_n;
  wire n3537_lo_p;
  wire n3537_lo_n;
  wire n3540_lo_p;
  wire n3540_lo_n;
  wire n3543_lo_p;
  wire n3543_lo_n;
  wire n3546_lo_p;
  wire n3546_lo_n;
  wire n3549_lo_p;
  wire n3549_lo_n;
  wire n3552_lo_p;
  wire n3552_lo_n;
  wire n3555_lo_p;
  wire n3555_lo_n;
  wire n3558_lo_p;
  wire n3558_lo_n;
  wire n3561_lo_p;
  wire n3561_lo_n;
  wire n3564_lo_p;
  wire n3564_lo_n;
  wire n3567_lo_p;
  wire n3567_lo_n;
  wire n3570_lo_p;
  wire n3570_lo_n;
  wire n3573_lo_p;
  wire n3573_lo_n;
  wire n3576_lo_p;
  wire n3576_lo_n;
  wire n3579_lo_p;
  wire n3579_lo_n;
  wire n3582_lo_p;
  wire n3582_lo_n;
  wire n3585_lo_p;
  wire n3585_lo_n;
  wire n3588_lo_p;
  wire n3588_lo_n;
  wire n3591_lo_p;
  wire n3591_lo_n;
  wire n3594_lo_p;
  wire n3594_lo_n;
  wire n3597_lo_p;
  wire n3597_lo_n;
  wire n3600_lo_p;
  wire n3600_lo_n;
  wire n3603_lo_p;
  wire n3603_lo_n;
  wire n3606_lo_p;
  wire n3606_lo_n;
  wire n3609_lo_p;
  wire n3609_lo_n;
  wire n3612_lo_p;
  wire n3612_lo_n;
  wire n3615_lo_p;
  wire n3615_lo_n;
  wire n3618_lo_p;
  wire n3618_lo_n;
  wire n3621_lo_p;
  wire n3621_lo_n;
  wire n3624_lo_p;
  wire n3624_lo_n;
  wire n3627_lo_p;
  wire n3627_lo_n;
  wire n3630_lo_p;
  wire n3630_lo_n;
  wire n3633_lo_p;
  wire n3633_lo_n;
  wire n3636_lo_p;
  wire n3636_lo_n;
  wire n3639_lo_p;
  wire n3639_lo_n;
  wire n3642_lo_p;
  wire n3642_lo_n;
  wire n3645_lo_p;
  wire n3645_lo_n;
  wire n3648_lo_p;
  wire n3648_lo_n;
  wire n3651_lo_p;
  wire n3651_lo_n;
  wire n3654_lo_p;
  wire n3654_lo_n;
  wire n3657_lo_p;
  wire n3657_lo_n;
  wire n3666_lo_p;
  wire n3666_lo_n;
  wire n3669_lo_p;
  wire n3669_lo_n;
  wire n3678_lo_p;
  wire n3678_lo_n;
  wire n3687_lo_p;
  wire n3687_lo_n;
  wire n3690_lo_p;
  wire n3690_lo_n;
  wire n3702_lo_p;
  wire n3702_lo_n;
  wire n3711_lo_p;
  wire n3711_lo_n;
  wire n3714_lo_p;
  wire n3714_lo_n;
  wire n3726_lo_p;
  wire n3726_lo_n;
  wire n3735_lo_p;
  wire n3735_lo_n;
  wire n3738_lo_p;
  wire n3738_lo_n;
  wire n3750_lo_p;
  wire n3750_lo_n;
  wire n3753_lo_p;
  wire n3753_lo_n;
  wire n3759_lo_p;
  wire n3759_lo_n;
  wire n3762_lo_p;
  wire n3762_lo_n;
  wire n3765_lo_p;
  wire n3765_lo_n;
  wire n3774_lo_p;
  wire n3774_lo_n;
  wire n3777_lo_p;
  wire n3777_lo_n;
  wire n3786_lo_p;
  wire n3786_lo_n;
  wire n3789_lo_p;
  wire n3789_lo_n;
  wire n3792_lo_p;
  wire n3792_lo_n;
  wire n3795_lo_p;
  wire n3795_lo_n;
  wire n3798_lo_p;
  wire n3798_lo_n;
  wire n3801_lo_p;
  wire n3801_lo_n;
  wire n3810_lo_p;
  wire n3810_lo_n;
  wire n3813_lo_p;
  wire n3813_lo_n;
  wire n3822_lo_p;
  wire n3822_lo_n;
  wire n3825_lo_p;
  wire n3825_lo_n;
  wire n3834_lo_p;
  wire n3834_lo_n;
  wire n3843_lo_p;
  wire n3843_lo_n;
  wire n3846_lo_p;
  wire n3846_lo_n;
  wire n3867_lo_p;
  wire n3867_lo_n;
  wire n3891_lo_p;
  wire n3891_lo_n;
  wire n3915_lo_p;
  wire n3915_lo_n;
  wire n3930_lo_p;
  wire n3930_lo_n;
  wire n3933_lo_p;
  wire n3933_lo_n;
  wire n3936_lo_p;
  wire n3936_lo_n;
  wire n3942_lo_p;
  wire n3942_lo_n;
  wire n3945_lo_p;
  wire n3945_lo_n;
  wire n3948_lo_p;
  wire n3948_lo_n;
  wire n3954_lo_p;
  wire n3954_lo_n;
  wire n3957_lo_p;
  wire n3957_lo_n;
  wire n3963_lo_p;
  wire n3963_lo_n;
  wire n3966_lo_p;
  wire n3966_lo_n;
  wire n3969_lo_p;
  wire n3969_lo_n;
  wire n3975_lo_p;
  wire n3975_lo_n;
  wire n3978_lo_p;
  wire n3978_lo_n;
  wire n3987_lo_p;
  wire n3987_lo_n;
  wire n3990_lo_p;
  wire n3990_lo_n;
  wire n4002_lo_p;
  wire n4002_lo_n;
  wire n4011_lo_p;
  wire n4011_lo_n;
  wire n4014_lo_p;
  wire n4014_lo_n;
  wire n4026_lo_p;
  wire n4026_lo_n;
  wire n4035_lo_p;
  wire n4035_lo_n;
  wire n4038_lo_p;
  wire n4038_lo_n;
  wire n4050_lo_p;
  wire n4050_lo_n;
  wire n4053_lo_p;
  wire n4053_lo_n;
  wire n4059_lo_p;
  wire n4059_lo_n;
  wire n4062_lo_p;
  wire n4062_lo_n;
  wire n4065_lo_p;
  wire n4065_lo_n;
  wire n4098_lo_p;
  wire n4098_lo_n;
  wire n4107_lo_p;
  wire n4107_lo_n;
  wire n4119_lo_p;
  wire n4119_lo_n;
  wire n4131_lo_p;
  wire n4131_lo_n;
  wire n4143_lo_p;
  wire n4143_lo_n;
  wire n4155_lo_p;
  wire n4155_lo_n;
  wire n4167_lo_p;
  wire n4167_lo_n;
  wire n4179_lo_p;
  wire n4179_lo_n;
  wire n4182_lo_p;
  wire n4182_lo_n;
  wire n4185_lo_p;
  wire n4185_lo_n;
  wire n4188_lo_p;
  wire n4188_lo_n;
  wire n4194_lo_p;
  wire n4194_lo_n;
  wire n4197_lo_p;
  wire n4197_lo_n;
  wire n4200_lo_p;
  wire n4200_lo_n;
  wire n4206_lo_p;
  wire n4206_lo_n;
  wire n4209_lo_p;
  wire n4209_lo_n;
  wire n4212_lo_p;
  wire n4212_lo_n;
  wire n4215_lo_p;
  wire n4215_lo_n;
  wire n4227_lo_p;
  wire n4227_lo_n;
  wire n4230_lo_p;
  wire n4230_lo_n;
  wire n4233_lo_p;
  wire n4233_lo_n;
  wire n4236_lo_p;
  wire n4236_lo_n;
  wire n4239_lo_p;
  wire n4239_lo_n;
  wire n4242_lo_p;
  wire n4242_lo_n;
  wire n4251_lo_p;
  wire n4251_lo_n;
  wire n4263_lo_p;
  wire n4263_lo_n;
  wire n4275_lo_p;
  wire n4275_lo_n;
  wire n4278_lo_p;
  wire n4278_lo_n;
  wire n4287_lo_p;
  wire n4287_lo_n;
  wire n4290_lo_p;
  wire n4290_lo_n;
  wire n4293_lo_p;
  wire n4293_lo_n;
  wire n4299_lo_p;
  wire n4299_lo_n;
  wire n4302_lo_p;
  wire n4302_lo_n;
  wire n4305_lo_p;
  wire n4305_lo_n;
  wire n4311_lo_p;
  wire n4311_lo_n;
  wire n4314_lo_p;
  wire n4314_lo_n;
  wire n4323_lo_p;
  wire n4323_lo_n;
  wire n4326_lo_p;
  wire n4326_lo_n;
  wire n4335_lo_p;
  wire n4335_lo_n;
  wire n4338_lo_p;
  wire n4338_lo_n;
  wire n4347_lo_p;
  wire n4347_lo_n;
  wire n4350_lo_p;
  wire n4350_lo_n;
  wire n4359_lo_p;
  wire n4359_lo_n;
  wire n4362_lo_p;
  wire n4362_lo_n;
  wire n4365_lo_p;
  wire n4365_lo_n;
  wire n4371_lo_p;
  wire n4371_lo_n;
  wire n4374_lo_p;
  wire n4374_lo_n;
  wire n4383_lo_p;
  wire n4383_lo_n;
  wire n4395_lo_p;
  wire n4395_lo_n;
  wire n4407_lo_p;
  wire n4407_lo_n;
  wire n4410_lo_p;
  wire n4410_lo_n;
  wire n4413_lo_p;
  wire n4413_lo_n;
  wire n4416_lo_p;
  wire n4416_lo_n;
  wire n4419_lo_p;
  wire n4419_lo_n;
  wire n4422_lo_p;
  wire n4422_lo_n;
  wire n4425_lo_p;
  wire n4425_lo_n;
  wire n4428_lo_p;
  wire n4428_lo_n;
  wire n4431_lo_p;
  wire n4431_lo_n;
  wire n4434_lo_p;
  wire n4434_lo_n;
  wire n4437_lo_p;
  wire n4437_lo_n;
  wire n4440_lo_p;
  wire n4440_lo_n;
  wire n4443_lo_p;
  wire n4443_lo_n;
  wire n4446_lo_p;
  wire n4446_lo_n;
  wire n4449_lo_p;
  wire n4449_lo_n;
  wire n4452_lo_p;
  wire n4452_lo_n;
  wire n4455_lo_p;
  wire n4455_lo_n;
  wire n4458_lo_p;
  wire n4458_lo_n;
  wire n4461_lo_p;
  wire n4461_lo_n;
  wire n4464_lo_p;
  wire n4464_lo_n;
  wire n4467_lo_p;
  wire n4467_lo_n;
  wire n4470_lo_p;
  wire n4470_lo_n;
  wire n4473_lo_p;
  wire n4473_lo_n;
  wire n4476_lo_p;
  wire n4476_lo_n;
  wire n4479_lo_p;
  wire n4479_lo_n;
  wire n4482_lo_p;
  wire n4482_lo_n;
  wire n4485_lo_p;
  wire n4485_lo_n;
  wire n4488_lo_p;
  wire n4488_lo_n;
  wire n4494_lo_p;
  wire n4494_lo_n;
  wire n4497_lo_p;
  wire n4497_lo_n;
  wire n4500_lo_p;
  wire n4500_lo_n;
  wire n4503_lo_p;
  wire n4503_lo_n;
  wire n4506_lo_p;
  wire n4506_lo_n;
  wire n4509_lo_p;
  wire n4509_lo_n;
  wire n4512_lo_p;
  wire n4512_lo_n;
  wire n4515_lo_p;
  wire n4515_lo_n;
  wire n4518_lo_p;
  wire n4518_lo_n;
  wire n4521_lo_p;
  wire n4521_lo_n;
  wire n4524_lo_p;
  wire n4524_lo_n;
  wire n4527_lo_p;
  wire n4527_lo_n;
  wire n4530_lo_p;
  wire n4530_lo_n;
  wire n4533_lo_p;
  wire n4533_lo_n;
  wire n4536_lo_p;
  wire n4536_lo_n;
  wire n4539_lo_p;
  wire n4539_lo_n;
  wire n4542_lo_p;
  wire n4542_lo_n;
  wire n4545_lo_p;
  wire n4545_lo_n;
  wire n4548_lo_p;
  wire n4548_lo_n;
  wire n4554_lo_p;
  wire n4554_lo_n;
  wire n4557_lo_p;
  wire n4557_lo_n;
  wire n4560_lo_p;
  wire n4560_lo_n;
  wire n4563_lo_p;
  wire n4563_lo_n;
  wire n4566_lo_p;
  wire n4566_lo_n;
  wire n4569_lo_p;
  wire n4569_lo_n;
  wire n4572_lo_p;
  wire n4572_lo_n;
  wire n4575_lo_p;
  wire n4575_lo_n;
  wire n4578_lo_p;
  wire n4578_lo_n;
  wire n4581_lo_p;
  wire n4581_lo_n;
  wire n4584_lo_p;
  wire n4584_lo_n;
  wire n4587_lo_p;
  wire n4587_lo_n;
  wire n4590_lo_p;
  wire n4590_lo_n;
  wire n4593_lo_p;
  wire n4593_lo_n;
  wire n4596_lo_p;
  wire n4596_lo_n;
  wire n4599_lo_p;
  wire n4599_lo_n;
  wire n4602_lo_p;
  wire n4602_lo_n;
  wire n4605_lo_p;
  wire n4605_lo_n;
  wire n4608_lo_p;
  wire n4608_lo_n;
  wire n4611_lo_p;
  wire n4611_lo_n;
  wire n4614_lo_p;
  wire n4614_lo_n;
  wire n4617_lo_p;
  wire n4617_lo_n;
  wire n4620_lo_p;
  wire n4620_lo_n;
  wire n4623_lo_p;
  wire n4623_lo_n;
  wire n4626_lo_p;
  wire n4626_lo_n;
  wire n4629_lo_p;
  wire n4629_lo_n;
  wire n4632_lo_p;
  wire n4632_lo_n;
  wire n4635_lo_p;
  wire n4635_lo_n;
  wire n4638_lo_p;
  wire n4638_lo_n;
  wire n4641_lo_p;
  wire n4641_lo_n;
  wire n4644_lo_p;
  wire n4644_lo_n;
  wire n4647_lo_p;
  wire n4647_lo_n;
  wire n4650_lo_p;
  wire n4650_lo_n;
  wire n4653_lo_p;
  wire n4653_lo_n;
  wire n4656_lo_p;
  wire n4656_lo_n;
  wire n4659_lo_p;
  wire n4659_lo_n;
  wire n4662_lo_p;
  wire n4662_lo_n;
  wire n4665_lo_p;
  wire n4665_lo_n;
  wire n4668_lo_p;
  wire n4668_lo_n;
  wire n4671_lo_p;
  wire n4671_lo_n;
  wire n4674_lo_p;
  wire n4674_lo_n;
  wire n4677_lo_p;
  wire n4677_lo_n;
  wire n4680_lo_p;
  wire n4680_lo_n;
  wire n4683_lo_p;
  wire n4683_lo_n;
  wire n4686_lo_p;
  wire n4686_lo_n;
  wire n4689_lo_p;
  wire n4689_lo_n;
  wire n4692_lo_p;
  wire n4692_lo_n;
  wire n4695_lo_p;
  wire n4695_lo_n;
  wire n4698_lo_p;
  wire n4698_lo_n;
  wire n4701_lo_p;
  wire n4701_lo_n;
  wire n4704_lo_p;
  wire n4704_lo_n;
  wire n4707_lo_p;
  wire n4707_lo_n;
  wire n4710_lo_p;
  wire n4710_lo_n;
  wire n4713_lo_p;
  wire n4713_lo_n;
  wire n4716_lo_p;
  wire n4716_lo_n;
  wire n4719_lo_p;
  wire n4719_lo_n;
  wire n4722_lo_p;
  wire n4722_lo_n;
  wire n4725_lo_p;
  wire n4725_lo_n;
  wire n4728_lo_p;
  wire n4728_lo_n;
  wire n4731_lo_p;
  wire n4731_lo_n;
  wire n4734_lo_p;
  wire n4734_lo_n;
  wire n4737_lo_p;
  wire n4737_lo_n;
  wire n4740_lo_p;
  wire n4740_lo_n;
  wire n4743_lo_p;
  wire n4743_lo_n;
  wire n6382_o2_p;
  wire n6382_o2_n;
  wire n6383_o2_p;
  wire n6383_o2_n;
  wire n6419_o2_p;
  wire n6419_o2_n;
  wire n6420_o2_p;
  wire n6420_o2_n;
  wire n6435_o2_p;
  wire n6435_o2_n;
  wire n6436_o2_p;
  wire n6436_o2_n;
  wire n6448_o2_p;
  wire n6448_o2_n;
  wire n6449_o2_p;
  wire n6449_o2_n;
  wire n6613_o2_p;
  wire n6613_o2_n;
  wire n6614_o2_p;
  wire n6614_o2_n;
  wire n6641_o2_p;
  wire n6641_o2_n;
  wire n6658_o2_p;
  wire n6658_o2_n;
  wire n6757_o2_p;
  wire n6757_o2_n;
  wire n6756_o2_p;
  wire n6756_o2_n;
  wire n7116_o2_p;
  wire n7116_o2_n;
  wire n7156_o2_p;
  wire n7156_o2_n;
  wire n6549_o2_p;
  wire n6549_o2_n;
  wire n6550_o2_p;
  wire n6550_o2_n;
  wire n7357_o2_p;
  wire n7357_o2_n;
  wire n7358_o2_p;
  wire n7358_o2_n;
  wire n7359_o2_p;
  wire n7359_o2_n;
  wire n7360_o2_p;
  wire n7360_o2_n;
  wire n6621_o2_p;
  wire n6621_o2_n;
  wire n6623_o2_p;
  wire n6623_o2_n;
  wire n6625_o2_p;
  wire n6625_o2_n;
  wire n6626_o2_p;
  wire n6626_o2_n;
  wire n6627_o2_p;
  wire n6627_o2_n;
  wire n6628_o2_p;
  wire n6628_o2_n;
  wire n6629_o2_p;
  wire n6629_o2_n;
  wire n6630_o2_p;
  wire n6630_o2_n;
  wire n6669_o2_p;
  wire n6669_o2_n;
  wire n7449_o2_p;
  wire n7449_o2_n;
  wire n7450_o2_p;
  wire n7450_o2_n;
  wire n7451_o2_p;
  wire n7451_o2_n;
  wire n7452_o2_p;
  wire n7452_o2_n;
  wire n6682_o2_p;
  wire n6682_o2_n;
  wire n6683_o2_p;
  wire n6683_o2_n;
  wire n6684_o2_p;
  wire n6684_o2_n;
  wire n6685_o2_p;
  wire n6685_o2_n;
  wire n7463_o2_p;
  wire n7463_o2_n;
  wire n6686_o2_p;
  wire n6686_o2_n;
  wire n6687_o2_p;
  wire n6687_o2_n;
  wire n6688_o2_p;
  wire n6688_o2_n;
  wire n6689_o2_p;
  wire n6689_o2_n;
  wire n6772_o2_p;
  wire n6772_o2_n;
  wire n6773_o2_p;
  wire n6773_o2_n;
  wire n6774_o2_p;
  wire n6774_o2_n;
  wire n6775_o2_p;
  wire n6775_o2_n;
  wire G3467_o2_p;
  wire G3467_o2_n;
  wire G2810_o2_p;
  wire G2810_o2_n;
  wire n6833_o2_p;
  wire n6833_o2_n;
  wire n6945_o2_p;
  wire n6945_o2_n;
  wire n6947_o2_p;
  wire n6947_o2_n;
  wire n6949_o2_p;
  wire n6949_o2_n;
  wire n6951_o2_p;
  wire n6951_o2_n;
  wire n6888_o2_p;
  wire n6888_o2_n;
  wire n6889_o2_p;
  wire n6889_o2_n;
  wire n6936_o2_p;
  wire n6936_o2_n;
  wire n6954_o2_p;
  wire n6954_o2_n;
  wire n6955_o2_p;
  wire n6955_o2_n;
  wire n6956_o2_p;
  wire n6956_o2_n;
  wire n6957_o2_p;
  wire n6957_o2_n;
  wire n6958_o2_p;
  wire n6958_o2_n;
  wire n6982_o2_p;
  wire n6982_o2_n;
  wire n6984_o2_p;
  wire n6984_o2_n;
  wire n6974_o2_p;
  wire n6974_o2_n;
  wire n6975_o2_p;
  wire n6975_o2_n;
  wire n6999_o2_p;
  wire n6999_o2_n;
  wire n7015_o2_p;
  wire n7015_o2_n;
  wire n7016_o2_p;
  wire n7016_o2_n;
  wire n7017_o2_p;
  wire n7017_o2_n;
  wire n7018_o2_p;
  wire n7018_o2_n;
  wire n7005_o2_p;
  wire n7005_o2_n;
  wire n7019_o2_p;
  wire n7019_o2_n;
  wire n7022_o2_p;
  wire n7022_o2_n;
  wire n7023_o2_p;
  wire n7023_o2_n;
  wire n7132_o2_p;
  wire n7132_o2_n;
  wire n7133_o2_p;
  wire n7133_o2_n;
  wire n7135_o2_p;
  wire n7135_o2_n;
  wire n7136_o2_p;
  wire n7136_o2_n;
  wire n7175_o2_p;
  wire n7175_o2_n;
  wire n7155_o2_p;
  wire n7155_o2_n;
  wire G3060_o2_p;
  wire G3060_o2_n;
  wire n7383_o2_p;
  wire n7383_o2_n;
  wire G3802_o2_p;
  wire G3802_o2_n;
  wire G3859_o2_p;
  wire G3859_o2_n;
  wire n7355_o2_p;
  wire n7355_o2_n;
  wire n7356_o2_p;
  wire n7356_o2_n;
  wire G4054_o2_p;
  wire G4054_o2_n;
  wire G4068_o2_p;
  wire G4068_o2_n;
  wire n7384_o2_p;
  wire n7384_o2_n;
  wire n7387_o2_p;
  wire n7387_o2_n;
  wire n7388_o2_p;
  wire n7388_o2_n;
  wire n7389_o2_p;
  wire n7389_o2_n;
  wire n7386_o2_p;
  wire n7386_o2_n;
  wire n7453_o2_p;
  wire n7453_o2_n;
  wire n7431_o2_p;
  wire n7431_o2_n;
  wire n7432_o2_p;
  wire n7432_o2_n;
  wire n7433_o2_p;
  wire n7433_o2_n;
  wire n7430_o2_p;
  wire n7430_o2_n;
  wire n7485_o2_p;
  wire n7485_o2_n;
  wire n7486_o2_p;
  wire n7486_o2_n;
  wire G2508_o2_p;
  wire G2508_o2_n;
  wire G2486_o2_p;
  wire G2486_o2_n;
  wire n2326_inv_p;
  wire n2326_inv_n;
  wire n2329_inv_p;
  wire n2329_inv_n;
  wire n3756_lo_buf_o2_p;
  wire n3756_lo_buf_o2_n;
  wire n4056_lo_buf_o2_p;
  wire n4056_lo_buf_o2_n;
  wire G3474_o2_p;
  wire G3474_o2_n;
  wire n2341_inv_p;
  wire n2341_inv_n;
  wire n7396_o2_p;
  wire n7396_o2_n;
  wire n7398_o2_p;
  wire n7398_o2_n;
  wire n7400_o2_p;
  wire n7400_o2_n;
  wire n7401_o2_p;
  wire n7401_o2_n;
  wire n7402_o2_p;
  wire n7402_o2_n;
  wire n7403_o2_p;
  wire n7403_o2_n;
  wire n7404_o2_p;
  wire n7404_o2_n;
  wire n7405_o2_p;
  wire n7405_o2_n;
  wire G2711_o2_p;
  wire G2711_o2_n;
  wire n2371_inv_p;
  wire n2371_inv_n;
  wire n7490_o2_p;
  wire n7490_o2_n;
  wire n7527_o2_p;
  wire n7527_o2_n;
  wire n7528_o2_p;
  wire n7528_o2_n;
  wire n7529_o2_p;
  wire n7529_o2_n;
  wire n7530_o2_p;
  wire n7530_o2_n;
  wire n7523_o2_p;
  wire n7523_o2_n;
  wire n7524_o2_p;
  wire n7524_o2_n;
  wire n7525_o2_p;
  wire n7525_o2_n;
  wire n7526_o2_p;
  wire n7526_o2_n;
  wire n4296_lo_buf_o2_p;
  wire n4296_lo_buf_o2_n;
  wire n4368_lo_buf_o2_p;
  wire n4368_lo_buf_o2_n;
  wire G2466_o2_p;
  wire G2466_o2_n;
  wire G2404_o2_p;
  wire G2404_o2_n;
  wire n7534_o2_p;
  wire n7534_o2_n;
  wire n7535_o2_p;
  wire n7535_o2_n;
  wire n7536_o2_p;
  wire n7536_o2_n;
  wire n7533_o2_p;
  wire n7533_o2_n;
  wire G1060_o2_p;
  wire G1060_o2_n;
  wire G963_o2_p;
  wire G963_o2_n;
  wire G2448_o2_p;
  wire G2448_o2_n;
  wire G2685_o2_p;
  wire G2685_o2_n;
  wire G2679_o2_p;
  wire G2679_o2_n;
  wire G2774_o2_p;
  wire G2774_o2_n;
  wire G2780_o2_p;
  wire G2780_o2_n;
  wire G2759_o2_p;
  wire G2759_o2_n;
  wire G2737_o2_p;
  wire G2737_o2_n;
  wire G2850_o2_p;
  wire G2850_o2_n;
  wire G3393_o2_p;
  wire G3393_o2_n;
  wire G3404_o2_p;
  wire G3404_o2_n;
  wire G3559_o2_p;
  wire G3559_o2_n;
  wire G2744_o2_p;
  wire G2744_o2_n;
  wire n3708_lo_buf_o2_p;
  wire n3708_lo_buf_o2_n;
  wire n3840_lo_buf_o2_p;
  wire n3840_lo_buf_o2_n;
  wire n4008_lo_buf_o2_p;
  wire n4008_lo_buf_o2_n;
  wire n4104_lo_buf_o2_p;
  wire n4104_lo_buf_o2_n;
  wire G1821_o2_p;
  wire G1821_o2_n;
  wire G1734_o2_p;
  wire G1734_o2_n;
  wire G3517_o2_p;
  wire G3517_o2_n;
  wire G3533_o2_p;
  wire G3533_o2_n;
  wire G3629_o2_p;
  wire G3629_o2_n;
  wire G3645_o2_p;
  wire G3645_o2_n;
  wire n2497_inv_p;
  wire n2497_inv_n;
  wire G2731_o2_p;
  wire G2731_o2_n;
  wire G2844_o2_p;
  wire G2844_o2_n;
  wire n3732_lo_buf_o2_p;
  wire n3732_lo_buf_o2_n;
  wire n4032_lo_buf_o2_p;
  wire n4032_lo_buf_o2_n;
  wire G3552_o2_p;
  wire G3552_o2_n;
  wire G2271_o2_p;
  wire G2271_o2_n;
  wire n4248_lo_buf_o2_p;
  wire n4248_lo_buf_o2_n;
  wire n4332_lo_buf_o2_p;
  wire n4332_lo_buf_o2_n;
  wire n4344_lo_buf_o2_p;
  wire n4344_lo_buf_o2_n;
  wire n4380_lo_buf_o2_p;
  wire n4380_lo_buf_o2_n;
  wire G2398_o2_p;
  wire G2398_o2_n;
  wire G2480_o2_p;
  wire G2480_o2_n;
  wire G2418_o2_p;
  wire G2418_o2_n;
  wire G1455_o2_p;
  wire G1455_o2_n;
  wire G1449_o2_p;
  wire G1449_o2_n;
  wire G1452_o2_p;
  wire G1452_o2_n;
  wire G1425_o2_p;
  wire G1425_o2_n;
  wire G1428_o2_p;
  wire G1428_o2_n;
  wire G1419_o2_p;
  wire G1419_o2_n;
  wire G1422_o2_p;
  wire G1422_o2_n;
  wire n4308_lo_buf_o2_p;
  wire n4308_lo_buf_o2_n;
  wire G2675_o2_p;
  wire G2675_o2_n;
  wire G3035_o2_p;
  wire G3035_o2_n;
  wire G3026_o2_p;
  wire G3026_o2_n;
  wire G3029_o2_p;
  wire G3029_o2_n;
  wire G3032_o2_p;
  wire G3032_o2_n;
  wire G2999_o2_p;
  wire G2999_o2_n;
  wire G3002_o2_p;
  wire G3002_o2_n;
  wire G2770_o2_p;
  wire G2770_o2_n;
  wire G3008_o2_p;
  wire G3008_o2_n;
  wire G2073_o2_p;
  wire G2073_o2_n;
  wire G2752_o2_p;
  wire G2752_o2_n;
  wire G3005_o2_p;
  wire G3005_o2_n;
  wire G5108_o2_p;
  wire G5108_o2_n;
  wire G5135_o2_p;
  wire G5135_o2_n;
  wire G5111_o2_p;
  wire G5111_o2_n;
  wire G5138_o2_p;
  wire G5138_o2_n;
  wire G3415_o2_p;
  wire G3415_o2_n;
  wire G3386_o2_p;
  wire G3386_o2_n;
  wire G3570_o2_p;
  wire G3570_o2_n;
  wire G2430_o2_p;
  wire G2430_o2_n;
  wire G3495_o2_p;
  wire G3495_o2_n;
  wire G3621_o2_p;
  wire G3621_o2_n;
  wire n4284_lo_buf_o2_p;
  wire n4284_lo_buf_o2_n;
  wire n4356_lo_buf_o2_p;
  wire n4356_lo_buf_o2_n;
  wire G2472_o2_p;
  wire G2472_o2_n;
  wire G2410_o2_p;
  wire G2410_o2_n;
  wire n3960_lo_buf_o2_p;
  wire n3960_lo_buf_o2_n;
  wire n3972_lo_buf_o2_p;
  wire n3972_lo_buf_o2_n;
  wire n2647_inv_p;
  wire n2647_inv_n;
  wire n2650_inv_p;
  wire n2650_inv_n;
  wire n3684_lo_buf_o2_p;
  wire n3684_lo_buf_o2_n;
  wire n4080_lo_buf_o2_p;
  wire n4080_lo_buf_o2_n;
  wire n4092_lo_buf_o2_p;
  wire n4092_lo_buf_o2_n;
  wire n2662_inv_p;
  wire n2662_inv_n;
  wire n2665_inv_p;
  wire n2665_inv_n;
  wire G1147_o2_p;
  wire G1147_o2_n;
  wire G2705_o2_p;
  wire G2705_o2_n;
  wire G2693_o2_p;
  wire G2693_o2_n;
  wire G2696_o2_p;
  wire G2696_o2_n;
  wire G2700_o2_p;
  wire G2700_o2_n;
  wire G2915_o2_p;
  wire G2915_o2_n;
  wire G2966_o2_p;
  wire G2966_o2_n;
  wire G2540_o2_p;
  wire G2540_o2_n;
  wire G2788_o2_p;
  wire G2788_o2_n;
  wire G2792_o2_p;
  wire G2792_o2_n;
  wire G2797_o2_p;
  wire G2797_o2_n;
  wire G2804_o2_p;
  wire G2804_o2_n;
  wire G1038_o2_p;
  wire G1038_o2_n;
  wire G1044_o2_p;
  wire G1044_o2_n;
  wire G1090_o2_p;
  wire G1090_o2_n;
  wire G1096_o2_p;
  wire G1096_o2_n;
  wire G1029_o2_p;
  wire G1029_o2_n;
  wire G3942_o2_p;
  wire G3942_o2_n;
  wire G3954_o2_p;
  wire G3954_o2_n;
  wire G4011_o2_p;
  wire G4011_o2_n;
  wire G4017_o2_p;
  wire G4017_o2_n;
  wire G1141_o2_p;
  wire G1141_o2_n;
  wire G1081_o2_p;
  wire G1081_o2_n;
  wire G2146_o2_p;
  wire G2146_o2_n;
  wire G2145_o2_p;
  wire G2145_o2_n;
  wire G2144_o2_p;
  wire G2144_o2_n;
  wire G2143_o2_p;
  wire G2143_o2_n;
  wire G2142_o2_p;
  wire G2142_o2_n;
  wire G2141_o2_p;
  wire G2141_o2_n;
  wire G2140_o2_p;
  wire G2140_o2_n;
  wire G2139_o2_p;
  wire G2139_o2_n;
  wire G3769_o2_p;
  wire G3769_o2_n;
  wire G3773_o2_p;
  wire G3773_o2_n;
  wire G3768_o2_p;
  wire G3768_o2_n;
  wire G4101_o2_p;
  wire G4101_o2_n;
  wire G3161_o2_p;
  wire G3161_o2_n;
  wire G4143_o2_p;
  wire G4143_o2_n;
  wire G3828_o2_p;
  wire G3828_o2_n;
  wire G3831_o2_p;
  wire G3831_o2_n;
  wire G3334_o2_p;
  wire G3334_o2_n;
  wire G3335_o2_p;
  wire G3335_o2_n;
  wire G3180_o2_p;
  wire G3180_o2_n;
  wire G3340_o2_p;
  wire G3340_o2_n;
  wire G3339_o2_p;
  wire G3339_o2_n;
  wire G3341_o2_p;
  wire G3341_o2_n;
  wire G3234_o2_p;
  wire G3234_o2_n;
  wire G3829_o2_p;
  wire G3829_o2_n;
  wire G3338_o2_p;
  wire G3338_o2_n;
  wire G3336_o2_p;
  wire G3336_o2_n;
  wire G3770_o2_p;
  wire G3770_o2_n;
  wire G3918_o2_p;
  wire G3918_o2_n;
  wire G3774_o2_p;
  wire G3774_o2_n;
  wire G3921_o2_p;
  wire G3921_o2_n;
  wire G3832_o2_p;
  wire G3832_o2_n;
  wire G3993_o2_p;
  wire G3993_o2_n;
  wire G2076_o2_p;
  wire G2076_o2_n;
  wire G2071_o2_p;
  wire G2071_o2_n;
  wire G2072_o2_p;
  wire G2072_o2_n;
  wire G2069_o2_p;
  wire G2069_o2_n;
  wire G2070_o2_p;
  wire G2070_o2_n;
  wire G2067_o2_p;
  wire G2067_o2_n;
  wire G2068_o2_p;
  wire G2068_o2_n;
  wire G4095_o2_p;
  wire G4095_o2_n;
  wire G3272_o2_p;
  wire G3272_o2_n;
  wire G3269_o2_p;
  wire G3269_o2_n;
  wire G3270_o2_p;
  wire G3270_o2_n;
  wire G3271_o2_p;
  wire G3271_o2_n;
  wire G3265_o2_p;
  wire G3265_o2_n;
  wire G3266_o2_p;
  wire G3266_o2_n;
  wire G4137_o2_p;
  wire G4137_o2_n;
  wire G3268_o2_p;
  wire G3268_o2_n;
  wire G2361_o2_p;
  wire G2361_o2_n;
  wire G3228_o2_p;
  wire G3228_o2_n;
  wire G3267_o2_p;
  wire G3267_o2_n;
  wire G2336_o2_p;
  wire G2336_o2_n;
  wire G3459_o2_p;
  wire G3459_o2_n;
  wire G3428_o2_p;
  wire G3428_o2_n;
  wire G3438_o2_p;
  wire G3438_o2_n;
  wire G3449_o2_p;
  wire G3449_o2_n;
  wire G3421_o2_p;
  wire G3421_o2_n;
  wire G3576_o2_p;
  wire G3576_o2_n;
  wire G3303_o2_p;
  wire G3303_o2_n;
  wire G3583_o2_p;
  wire G3583_o2_n;
  wire G3594_o2_p;
  wire G3594_o2_n;
  wire G3674_o2_p;
  wire G3674_o2_n;
  wire G3685_o2_p;
  wire G3685_o2_n;
  wire G4504_o2_p;
  wire G4504_o2_n;
  wire G4180_o2_p;
  wire G4180_o2_n;
  wire G5123_o2_p;
  wire G5123_o2_n;
  wire G5142_o2_p;
  wire G5142_o2_n;
  wire G5126_o2_p;
  wire G5126_o2_n;
  wire G5144_o2_p;
  wire G5144_o2_n;
  wire G3912_o2_p;
  wire G3912_o2_n;
  wire G4417_o2_p;
  wire G4417_o2_n;
  wire G4420_o2_p;
  wire G4420_o2_n;
  wire G3969_o2_p;
  wire G3969_o2_n;
  wire G4023_o2_p;
  wire G4023_o2_n;
  wire G2720_o2_p;
  wire G2720_o2_n;
  wire G2837_o2_p;
  wire G2837_o2_n;
  wire n2965_inv_p;
  wire n2965_inv_n;
  wire n2968_inv_p;
  wire n2968_inv_n;
  wire n2971_inv_p;
  wire n2971_inv_n;
  wire n2974_inv_p;
  wire n2974_inv_n;
  wire G1876_o2_p;
  wire G1876_o2_n;
  wire G4996_o2_p;
  wire G4996_o2_n;
  wire G4984_o2_p;
  wire G4984_o2_n;
  wire G4920_o2_p;
  wire G4920_o2_n;
  wire G4923_o2_p;
  wire G4923_o2_n;
  wire G4930_o2_p;
  wire G4930_o2_n;
  wire G4933_o2_p;
  wire G4933_o2_n;
  wire n4320_lo_buf_o2_p;
  wire n4320_lo_buf_o2_n;
  wire G2424_o2_p;
  wire G2424_o2_n;
  wire G3317_o2_p;
  wire G3317_o2_n;
  wire G3503_o2_p;
  wire G3503_o2_n;
  wire G3485_o2_p;
  wire G3485_o2_n;
  wire G3611_o2_p;
  wire G3611_o2_n;
  wire n3864_lo_buf_o2_p;
  wire n3864_lo_buf_o2_n;
  wire n3888_lo_buf_o2_p;
  wire n3888_lo_buf_o2_n;
  wire n4116_lo_buf_o2_p;
  wire n4116_lo_buf_o2_n;
  wire n4128_lo_buf_o2_p;
  wire n4128_lo_buf_o2_n;
  wire n4140_lo_buf_o2_p;
  wire n4140_lo_buf_o2_n;
  wire n4152_lo_buf_o2_p;
  wire n4152_lo_buf_o2_n;
  wire G1815_o2_p;
  wire G1815_o2_n;
  wire G1728_o2_p;
  wire G1728_o2_n;
  wire G1035_o2_p;
  wire G1035_o2_n;
  wire G1041_o2_p;
  wire G1041_o2_n;
  wire G1087_o2_p;
  wire G1087_o2_n;
  wire G1093_o2_p;
  wire G1093_o2_n;
  wire G1132_o2_p;
  wire G1132_o2_n;
  wire G1108_o2_p;
  wire G1108_o2_n;
  wire G1138_o2_p;
  wire G1138_o2_n;
  wire G1114_o2_p;
  wire G1114_o2_n;
  wire G1807_o2_p;
  wire G1807_o2_n;
  wire G2108_o2_p;
  wire G2108_o2_n;
  wire G1126_o2_p;
  wire G1126_o2_n;
  wire G1899_o2_p;
  wire G1899_o2_n;
  wire G2134_o2_p;
  wire G2134_o2_n;
  wire G1852_o2_p;
  wire G1852_o2_n;
  wire G2116_o2_p;
  wire G2116_o2_n;
  wire G2543_o2_p;
  wire G2543_o2_n;
  wire G2727_o2_p;
  wire G2727_o2_n;
  wire G2715_o2_p;
  wire G2715_o2_n;
  wire G2832_o2_p;
  wire G2832_o2_n;
  wire G1873_o2_p;
  wire G1873_o2_n;
  wire G3291_o2_p;
  wire G3291_o2_n;
  wire G5025_o2_p;
  wire G5025_o2_n;
  wire G5036_o2_p;
  wire G5036_o2_n;
  wire G3132_o2_p;
  wire G3132_o2_n;
  wire G5038_o2_p;
  wire G5038_o2_n;
  wire G5039_o2_p;
  wire G5039_o2_n;
  wire n3118_inv_p;
  wire n3118_inv_n;
  wire n3121_inv_p;
  wire n3121_inv_n;
  wire n3124_inv_p;
  wire n3124_inv_n;
  wire n3127_inv_p;
  wire n3127_inv_n;
  wire n3984_lo_buf_o2_p;
  wire n3984_lo_buf_o2_n;
  wire G1802_o2_p;
  wire G1802_o2_n;
  wire G1804_o2_p;
  wire G1804_o2_n;
  wire G1849_o2_p;
  wire G1849_o2_n;
  wire G1851_o2_p;
  wire G1851_o2_n;
  wire G2492_o2_p;
  wire G2492_o2_n;
  wire G1799_o2_p;
  wire G1799_o2_n;
  wire G4231_o2_p;
  wire G4231_o2_n;
  wire G4234_o2_p;
  wire G4234_o2_n;
  wire G4245_o2_p;
  wire G4245_o2_n;
  wire G4247_o2_p;
  wire G4247_o2_n;
  wire G1894_o2_p;
  wire G1894_o2_n;
  wire G1846_o2_p;
  wire G1846_o2_n;
  wire G4238_o2_p;
  wire G4238_o2_n;
  wire G4249_o2_p;
  wire G4249_o2_n;
  wire G2293_o2_p;
  wire G2293_o2_n;
  wire G5022_o2_p;
  wire G5022_o2_n;
  wire G5006_o2_p;
  wire G5006_o2_n;
  wire G4944_o2_p;
  wire G4944_o2_n;
  wire G4946_o2_p;
  wire G4946_o2_n;
  wire G4954_o2_p;
  wire G4954_o2_n;
  wire G4956_o2_p;
  wire G4956_o2_n;
  wire G3546_o2_p;
  wire G3546_o2_n;
  wire G3658_o2_p;
  wire G3658_o2_n;
  wire G1344_o2_p;
  wire G1344_o2_n;
  wire G2921_o2_p;
  wire G2921_o2_n;
  wire n3912_lo_buf_o2_p;
  wire n3912_lo_buf_o2_n;
  wire G1835_o2_p;
  wire G1835_o2_n;
  wire G3810_o2_p;
  wire G3810_o2_n;
  wire G3866_o2_p;
  wire G3866_o2_n;
  wire G3811_o2_p;
  wire G3811_o2_n;
  wire G2269_o2_p;
  wire G2269_o2_n;
  wire G3812_o2_p;
  wire G3812_o2_n;
  wire G3867_o2_p;
  wire G3867_o2_n;
  wire G3868_o2_p;
  wire G3868_o2_n;
  wire G3809_o2_p;
  wire G3809_o2_n;
  wire G3716_o2_p;
  wire G3716_o2_n;
  wire G4529_o2_p;
  wire G4529_o2_n;
  wire G4670_o2_p;
  wire G4670_o2_n;
  wire G4493_o2_p;
  wire G4493_o2_n;
  wire G4580_o2_p;
  wire G4580_o2_n;
  wire G3822_o2_p;
  wire G3822_o2_n;
  wire G3877_o2_p;
  wire G3877_o2_n;
  wire G4131_o2_p;
  wire G4131_o2_n;
  wire G4170_o2_p;
  wire G4170_o2_n;
  wire G4051_o2_p;
  wire G4051_o2_n;
  wire G4065_o2_p;
  wire G4065_o2_n;
  wire G4697_o2_p;
  wire G4697_o2_n;
  wire G4706_o2_p;
  wire G4706_o2_n;
  wire G2460_o2_p;
  wire G2460_o2_n;
  wire G2454_o2_p;
  wire G2454_o2_n;
  wire G2392_o2_p;
  wire G2392_o2_n;
  wire G2386_o2_p;
  wire G2386_o2_n;
  wire n4260_lo_buf_o2_p;
  wire n4260_lo_buf_o2_n;
  wire n4272_lo_buf_o2_p;
  wire n4272_lo_buf_o2_n;
  wire n4392_lo_buf_o2_p;
  wire n4392_lo_buf_o2_n;
  wire n4404_lo_buf_o2_p;
  wire n4404_lo_buf_o2_n;
  wire G1512_o2_p;
  wire G1512_o2_n;
  wire G3135_o2_p;
  wire G3135_o2_n;
  wire G2379_o2_p;
  wire G2379_o2_n;
  wire n4164_lo_buf_o2_p;
  wire n4164_lo_buf_o2_n;
  wire n4176_lo_buf_o2_p;
  wire n4176_lo_buf_o2_n;
  wire n4224_lo_buf_o2_p;
  wire n4224_lo_buf_o2_n;
  wire G2975_o2_p;
  wire G2975_o2_n;
  wire G2978_o2_p;
  wire G2978_o2_n;
  wire G2933_o2_p;
  wire G2933_o2_n;
  wire G2936_o2_p;
  wire G2936_o2_n;
  wire G1356_o2_p;
  wire G1356_o2_n;
  wire G1359_o2_p;
  wire G1359_o2_n;
  wire G1398_o2_p;
  wire G1398_o2_n;
  wire G1401_o2_p;
  wire G1401_o2_n;
  wire g1192_p;
  wire g1192_n;
  wire g1193_p;
  wire g1193_n;
  wire g1194_p;
  wire g1194_n;
  wire g1195_p;
  wire g1195_n;
  wire g1196_p;
  wire g1196_n;
  wire g1197_p;
  wire g1197_n;
  wire g1198_p;
  wire g1198_n;
  wire g1199_p;
  wire g1199_n;
  wire g1200_p;
  wire g1200_n;
  wire g1201_p;
  wire g1201_n;
  wire g1202_p;
  wire g1202_n;
  wire g1203_p;
  wire g1203_n;
  wire g1204_p;
  wire g1204_n;
  wire g1205_p;
  wire g1205_n;
  wire g1206_p;
  wire g1206_n;
  wire g1207_p;
  wire g1207_n;
  wire g1208_p;
  wire g1208_n;
  wire g1209_p;
  wire g1209_n;
  wire g1210_p;
  wire g1210_n;
  wire g1211_p;
  wire g1211_n;
  wire g1212_p;
  wire g1212_n;
  wire g1213_p;
  wire g1213_n;
  wire g1214_p;
  wire g1214_n;
  wire g1215_p;
  wire g1215_n;
  wire g1216_p;
  wire g1216_n;
  wire g1217_p;
  wire g1217_n;
  wire g1218_p;
  wire g1218_n;
  wire g1219_p;
  wire g1219_n;
  wire g1220_p;
  wire g1220_n;
  wire g1221_p;
  wire g1221_n;
  wire g1222_p;
  wire g1222_n;
  wire g1223_p;
  wire g1223_n;
  wire g1224_p;
  wire g1224_n;
  wire g1225_p;
  wire g1225_n;
  wire g1226_p;
  wire g1226_n;
  wire g1227_p;
  wire g1227_n;
  wire g1228_p;
  wire g1228_n;
  wire g1229_p;
  wire g1229_n;
  wire g1230_p;
  wire g1230_n;
  wire g1231_p;
  wire g1231_n;
  wire g1232_p;
  wire g1232_n;
  wire g1233_p;
  wire g1233_n;
  wire g1234_p;
  wire g1234_n;
  wire g1235_p;
  wire g1235_n;
  wire g1236_p;
  wire g1236_n;
  wire g1237_p;
  wire g1237_n;
  wire g1238_p;
  wire g1238_n;
  wire g1239_p;
  wire g1239_n;
  wire g1240_p;
  wire g1240_n;
  wire g1241_p;
  wire g1241_n;
  wire g1242_p;
  wire g1242_n;
  wire g1243_p;
  wire g1243_n;
  wire g1244_p;
  wire g1244_n;
  wire g1245_p;
  wire g1245_n;
  wire g1246_p;
  wire g1246_n;
  wire g1247_p;
  wire g1247_n;
  wire g1248_p;
  wire g1248_n;
  wire g1249_p;
  wire g1249_n;
  wire g1250_p;
  wire g1250_n;
  wire g1251_p;
  wire g1251_n;
  wire g1252_p;
  wire g1252_n;
  wire g1253_p;
  wire g1253_n;
  wire g1254_p;
  wire g1254_n;
  wire g1255_p;
  wire g1255_n;
  wire g1256_p;
  wire g1256_n;
  wire g1257_p;
  wire g1257_n;
  wire g1258_p;
  wire g1258_n;
  wire g1259_p;
  wire g1259_n;
  wire g1260_p;
  wire g1260_n;
  wire g1261_p;
  wire g1261_n;
  wire g1262_p;
  wire g1262_n;
  wire g1263_p;
  wire g1263_n;
  wire g1264_p;
  wire g1264_n;
  wire g1265_p;
  wire g1265_n;
  wire g1266_p;
  wire g1266_n;
  wire g1267_p;
  wire g1267_n;
  wire g1268_p;
  wire g1268_n;
  wire g1269_p;
  wire g1269_n;
  wire g1270_p;
  wire g1270_n;
  wire g1271_p;
  wire g1271_n;
  wire g1272_p;
  wire g1272_n;
  wire g1273_p;
  wire g1273_n;
  wire g1274_p;
  wire g1274_n;
  wire g1275_p;
  wire g1275_n;
  wire g1276_p;
  wire g1276_n;
  wire g1277_p;
  wire g1277_n;
  wire g1278_p;
  wire g1278_n;
  wire g1279_p;
  wire g1279_n;
  wire g1280_p;
  wire g1280_n;
  wire g1281_p;
  wire g1281_n;
  wire g1282_p;
  wire g1282_n;
  wire g1283_p;
  wire g1283_n;
  wire g1284_p;
  wire g1284_n;
  wire g1285_p;
  wire g1285_n;
  wire g1286_p;
  wire g1286_n;
  wire g1287_p;
  wire g1287_n;
  wire g1288_p;
  wire g1288_n;
  wire g1289_p;
  wire g1289_n;
  wire g1290_p;
  wire g1290_n;
  wire g1291_p;
  wire g1291_n;
  wire g1292_p;
  wire g1292_n;
  wire g1293_p;
  wire g1293_n;
  wire g1294_p;
  wire g1294_n;
  wire g1295_p;
  wire g1295_n;
  wire g1296_p;
  wire g1296_n;
  wire g1297_p;
  wire g1297_n;
  wire g1298_p;
  wire g1298_n;
  wire g1299_p;
  wire g1299_n;
  wire g1300_p;
  wire g1300_n;
  wire g1301_p;
  wire g1301_n;
  wire g1302_p;
  wire g1302_n;
  wire g1303_p;
  wire g1303_n;
  wire g1304_p;
  wire g1304_n;
  wire g1305_p;
  wire g1305_n;
  wire g1306_p;
  wire g1306_n;
  wire g1307_p;
  wire g1307_n;
  wire g1308_p;
  wire g1308_n;
  wire g1309_p;
  wire g1309_n;
  wire g1310_p;
  wire g1310_n;
  wire g1311_p;
  wire g1311_n;
  wire g1312_p;
  wire g1312_n;
  wire g1313_p;
  wire g1313_n;
  wire g1314_p;
  wire g1314_n;
  wire g1315_p;
  wire g1315_n;
  wire g1316_p;
  wire g1316_n;
  wire g1317_p;
  wire g1317_n;
  wire g1318_p;
  wire g1318_n;
  wire g1319_p;
  wire g1319_n;
  wire g1320_p;
  wire g1320_n;
  wire g1321_p;
  wire g1321_n;
  wire g1322_p;
  wire g1322_n;
  wire g1323_p;
  wire g1323_n;
  wire g1324_p;
  wire g1324_n;
  wire g1325_p;
  wire g1325_n;
  wire g1326_p;
  wire g1326_n;
  wire g1327_p;
  wire g1327_n;
  wire g1328_p;
  wire g1328_n;
  wire g1329_p;
  wire g1329_n;
  wire g1330_p;
  wire g1330_n;
  wire g1331_p;
  wire g1331_n;
  wire g1332_p;
  wire g1332_n;
  wire g1333_p;
  wire g1333_n;
  wire g1334_p;
  wire g1334_n;
  wire g1335_p;
  wire g1335_n;
  wire g1336_p;
  wire g1336_n;
  wire g1337_p;
  wire g1337_n;
  wire g1338_p;
  wire g1338_n;
  wire g1339_p;
  wire g1339_n;
  wire g1340_p;
  wire g1340_n;
  wire g1341_p;
  wire g1341_n;
  wire g1342_p;
  wire g1342_n;
  wire g1343_p;
  wire g1343_n;
  wire g1344_p;
  wire g1344_n;
  wire g1345_p;
  wire g1345_n;
  wire g1346_p;
  wire g1346_n;
  wire g1347_p;
  wire g1347_n;
  wire g1348_p;
  wire g1348_n;
  wire g1349_p;
  wire g1349_n;
  wire g1350_p;
  wire g1350_n;
  wire g1351_p;
  wire g1351_n;
  wire g1352_p;
  wire g1352_n;
  wire g1353_p;
  wire g1353_n;
  wire g1354_p;
  wire g1354_n;
  wire g1355_p;
  wire g1355_n;
  wire g1356_p;
  wire g1356_n;
  wire g1357_p;
  wire g1357_n;
  wire g1358_p;
  wire g1358_n;
  wire g1359_p;
  wire g1359_n;
  wire g1360_p;
  wire g1360_n;
  wire g1361_p;
  wire g1361_n;
  wire g1362_p;
  wire g1362_n;
  wire g1363_p;
  wire g1363_n;
  wire g1364_p;
  wire g1364_n;
  wire g1365_p;
  wire g1365_n;
  wire g1366_p;
  wire g1366_n;
  wire g1367_p;
  wire g1367_n;
  wire g1368_p;
  wire g1368_n;
  wire g1369_p;
  wire g1369_n;
  wire g1370_p;
  wire g1370_n;
  wire g1371_p;
  wire g1371_n;
  wire g1372_p;
  wire g1372_n;
  wire g1373_p;
  wire g1373_n;
  wire g1374_p;
  wire g1374_n;
  wire g1375_p;
  wire g1375_n;
  wire g1376_p;
  wire g1376_n;
  wire g1377_p;
  wire g1377_n;
  wire g1378_p;
  wire g1378_n;
  wire g1379_p;
  wire g1379_n;
  wire g1380_p;
  wire g1380_n;
  wire g1381_p;
  wire g1381_n;
  wire g1382_p;
  wire g1382_n;
  wire g1383_p;
  wire g1383_n;
  wire g1384_p;
  wire g1384_n;
  wire g1385_p;
  wire g1385_n;
  wire g1386_p;
  wire g1386_n;
  wire g1387_p;
  wire g1387_n;
  wire g1388_p;
  wire g1388_n;
  wire g1389_p;
  wire g1389_n;
  wire g1390_p;
  wire g1390_n;
  wire g1391_p;
  wire g1391_n;
  wire g1392_p;
  wire g1392_n;
  wire g1393_p;
  wire g1393_n;
  wire g1394_p;
  wire g1394_n;
  wire g1395_p;
  wire g1395_n;
  wire g1396_p;
  wire g1396_n;
  wire g1397_p;
  wire g1397_n;
  wire g1398_p;
  wire g1398_n;
  wire g1399_p;
  wire g1399_n;
  wire g1400_p;
  wire g1400_n;
  wire g1401_p;
  wire g1401_n;
  wire g1402_p;
  wire g1402_n;
  wire g1403_p;
  wire g1403_n;
  wire g1404_p;
  wire g1404_n;
  wire g1405_p;
  wire g1405_n;
  wire g1406_p;
  wire g1406_n;
  wire g1407_p;
  wire g1407_n;
  wire g1408_p;
  wire g1408_n;
  wire g1409_p;
  wire g1409_n;
  wire g1410_p;
  wire g1410_n;
  wire g1411_p;
  wire g1411_n;
  wire g1412_p;
  wire g1412_n;
  wire g1413_p;
  wire g1413_n;
  wire g1414_p;
  wire g1414_n;
  wire g1415_p;
  wire g1415_n;
  wire g1416_p;
  wire g1416_n;
  wire g1417_p;
  wire g1417_n;
  wire g1418_p;
  wire g1418_n;
  wire g1419_p;
  wire g1419_n;
  wire g1420_p;
  wire g1420_n;
  wire g1421_p;
  wire g1421_n;
  wire g1422_p;
  wire g1422_n;
  wire g1423_p;
  wire g1423_n;
  wire g1424_p;
  wire g1424_n;
  wire g1425_p;
  wire g1425_n;
  wire g1426_p;
  wire g1426_n;
  wire g1427_p;
  wire g1427_n;
  wire g1428_p;
  wire g1428_n;
  wire g1429_p;
  wire g1429_n;
  wire g1430_p;
  wire g1430_n;
  wire g1431_p;
  wire g1431_n;
  wire g1432_p;
  wire g1432_n;
  wire g1433_p;
  wire g1433_n;
  wire g1434_p;
  wire g1434_n;
  wire g1435_p;
  wire g1435_n;
  wire g1436_p;
  wire g1436_n;
  wire g1437_p;
  wire g1437_n;
  wire g1438_p;
  wire g1438_n;
  wire g1439_p;
  wire g1439_n;
  wire g1440_p;
  wire g1440_n;
  wire g1441_p;
  wire g1441_n;
  wire g1442_p;
  wire g1442_n;
  wire g1443_p;
  wire g1443_n;
  wire g1444_p;
  wire g1444_n;
  wire g1445_p;
  wire g1445_n;
  wire g1446_p;
  wire g1446_n;
  wire g1447_p;
  wire g1447_n;
  wire g1448_p;
  wire g1448_n;
  wire g1449_p;
  wire g1449_n;
  wire g1450_p;
  wire g1450_n;
  wire g1451_p;
  wire g1451_n;
  wire g1452_p;
  wire g1452_n;
  wire g1453_p;
  wire g1453_n;
  wire g1454_p;
  wire g1454_n;
  wire g1455_p;
  wire g1455_n;
  wire g1456_p;
  wire g1456_n;
  wire g1457_p;
  wire g1457_n;
  wire g1458_p;
  wire g1458_n;
  wire g1459_p;
  wire g1459_n;
  wire g1460_p;
  wire g1460_n;
  wire g1461_p;
  wire g1461_n;
  wire g1462_p;
  wire g1462_n;
  wire g1463_p;
  wire g1463_n;
  wire g1464_p;
  wire g1464_n;
  wire g1465_p;
  wire g1465_n;
  wire g1466_p;
  wire g1466_n;
  wire g1467_p;
  wire g1467_n;
  wire g1468_p;
  wire g1468_n;
  wire g1469_p;
  wire g1469_n;
  wire g1470_p;
  wire g1470_n;
  wire g1471_p;
  wire g1471_n;
  wire g1472_p;
  wire g1472_n;
  wire g1473_p;
  wire g1473_n;
  wire g1474_p;
  wire g1474_n;
  wire g1475_p;
  wire g1475_n;
  wire g1476_p;
  wire g1476_n;
  wire g1477_p;
  wire g1477_n;
  wire g1478_p;
  wire g1478_n;
  wire g1479_p;
  wire g1479_n;
  wire g1480_p;
  wire g1480_n;
  wire g1481_p;
  wire g1481_n;
  wire g1482_p;
  wire g1482_n;
  wire g1483_p;
  wire g1483_n;
  wire g1484_p;
  wire g1484_n;
  wire g1485_p;
  wire g1485_n;
  wire g1486_p;
  wire g1486_n;
  wire g1487_p;
  wire g1487_n;
  wire g1488_p;
  wire g1488_n;
  wire g1489_p;
  wire g1489_n;
  wire g1490_p;
  wire g1490_n;
  wire g1491_p;
  wire g1491_n;
  wire g1492_p;
  wire g1492_n;
  wire g1493_p;
  wire g1493_n;
  wire g1494_p;
  wire g1494_n;
  wire g1495_p;
  wire g1495_n;
  wire g1496_p;
  wire g1496_n;
  wire g1497_p;
  wire g1497_n;
  wire g1498_p;
  wire g1498_n;
  wire g1499_p;
  wire g1499_n;
  wire g1500_p;
  wire g1500_n;
  wire g1501_p;
  wire g1501_n;
  wire g1502_p;
  wire g1502_n;
  wire g1503_p;
  wire g1503_n;
  wire g1504_p;
  wire g1504_n;
  wire g1505_p;
  wire g1505_n;
  wire g1506_p;
  wire g1506_n;
  wire g1507_p;
  wire g1507_n;
  wire g1508_p;
  wire g1508_n;
  wire g1509_p;
  wire g1509_n;
  wire g1510_p;
  wire g1510_n;
  wire g1511_p;
  wire g1511_n;
  wire g1512_p;
  wire g1512_n;
  wire g1513_p;
  wire g1513_n;
  wire g1514_p;
  wire g1514_n;
  wire g1515_p;
  wire g1515_n;
  wire g1516_p;
  wire g1516_n;
  wire g1517_p;
  wire g1517_n;
  wire g1518_p;
  wire g1518_n;
  wire g1519_p;
  wire g1519_n;
  wire g1520_p;
  wire g1520_n;
  wire g1521_p;
  wire g1521_n;
  wire g1522_p;
  wire g1522_n;
  wire g1523_p;
  wire g1523_n;
  wire g1524_p;
  wire g1524_n;
  wire g1525_p;
  wire g1525_n;
  wire g1526_p;
  wire g1526_n;
  wire g1527_p;
  wire g1527_n;
  wire g1528_p;
  wire g1528_n;
  wire g1529_p;
  wire g1529_n;
  wire g1530_p;
  wire g1530_n;
  wire g1531_p;
  wire g1531_n;
  wire g1532_p;
  wire g1532_n;
  wire g1533_p;
  wire g1533_n;
  wire g1534_p;
  wire g1534_n;
  wire g1535_p;
  wire g1535_n;
  wire g1536_p;
  wire g1536_n;
  wire g1537_p;
  wire g1537_n;
  wire g1538_p;
  wire g1538_n;
  wire g1539_p;
  wire g1539_n;
  wire g1540_p;
  wire g1540_n;
  wire g1541_p;
  wire g1541_n;
  wire g1542_p;
  wire g1542_n;
  wire g1543_p;
  wire g1543_n;
  wire g1544_p;
  wire g1544_n;
  wire g1545_p;
  wire g1545_n;
  wire g1546_p;
  wire g1546_n;
  wire g1547_p;
  wire g1547_n;
  wire g1548_p;
  wire g1548_n;
  wire g1549_p;
  wire g1549_n;
  wire g1550_p;
  wire g1550_n;
  wire g1551_p;
  wire g1551_n;
  wire g1552_p;
  wire g1552_n;
  wire g1553_p;
  wire g1553_n;
  wire g1554_p;
  wire g1554_n;
  wire g1555_p;
  wire g1555_n;
  wire g1556_p;
  wire g1556_n;
  wire g1557_p;
  wire g1557_n;
  wire g1558_p;
  wire g1558_n;
  wire g1559_p;
  wire g1559_n;
  wire g1560_p;
  wire g1560_n;
  wire g1561_p;
  wire g1561_n;
  wire g1562_p;
  wire g1562_n;
  wire g1563_p;
  wire g1563_n;
  wire g1564_p;
  wire g1564_n;
  wire g1565_p;
  wire g1565_n;
  wire g1566_p;
  wire g1566_n;
  wire g1567_p;
  wire g1567_n;
  wire g1568_p;
  wire g1568_n;
  wire g1569_p;
  wire g1569_n;
  wire g1570_p;
  wire g1570_n;
  wire g1571_p;
  wire g1571_n;
  wire g1572_p;
  wire g1572_n;
  wire g1573_p;
  wire g1573_n;
  wire g1574_p;
  wire g1574_n;
  wire g1575_p;
  wire g1575_n;
  wire g1576_p;
  wire g1576_n;
  wire g1577_p;
  wire g1577_n;
  wire g1578_p;
  wire g1578_n;
  wire g1579_p;
  wire g1579_n;
  wire g1580_p;
  wire g1580_n;
  wire g1581_p;
  wire g1581_n;
  wire g1582_p;
  wire g1582_n;
  wire g1583_p;
  wire g1583_n;
  wire g1584_p;
  wire g1584_n;
  wire g1585_p;
  wire g1585_n;
  wire g1586_p;
  wire g1586_n;
  wire g1587_p;
  wire g1587_n;
  wire g1588_p;
  wire g1588_n;
  wire g1589_p;
  wire g1589_n;
  wire g1590_p;
  wire g1590_n;
  wire g1591_p;
  wire g1591_n;
  wire g1592_p;
  wire g1592_n;
  wire g1593_p;
  wire g1593_n;
  wire g1594_p;
  wire g1594_n;
  wire g1595_p;
  wire g1595_n;
  wire g1596_p;
  wire g1596_n;
  wire g1597_p;
  wire g1597_n;
  wire g1598_p;
  wire g1598_n;
  wire g1599_p;
  wire g1599_n;
  wire g1600_p;
  wire g1600_n;
  wire g1601_p;
  wire g1601_n;
  wire g1602_p;
  wire g1602_n;
  wire g1603_p;
  wire g1603_n;
  wire g1604_p;
  wire g1604_n;
  wire g1605_p;
  wire g1605_n;
  wire g1606_p;
  wire g1606_n;
  wire g1607_p;
  wire g1607_n;
  wire g1608_p;
  wire g1608_n;
  wire g1609_p;
  wire g1609_n;
  wire g1610_p;
  wire g1610_n;
  wire g1611_p;
  wire g1611_n;
  wire g1612_p;
  wire g1612_n;
  wire g1613_p;
  wire g1613_n;
  wire g1614_p;
  wire g1614_n;
  wire g1615_p;
  wire g1615_n;
  wire g1616_p;
  wire g1616_n;
  wire g1617_p;
  wire g1617_n;
  wire g1618_p;
  wire g1618_n;
  wire g1619_p;
  wire g1619_n;
  wire g1620_p;
  wire g1620_n;
  wire g1621_p;
  wire g1621_n;
  wire g1622_p;
  wire g1622_n;
  wire g1623_p;
  wire g1623_n;
  wire g1624_p;
  wire g1624_n;
  wire g1625_p;
  wire g1625_n;
  wire g1626_p;
  wire g1626_n;
  wire g1627_p;
  wire g1627_n;
  wire g1628_p;
  wire g1628_n;
  wire g1629_p;
  wire g1629_n;
  wire g1630_p;
  wire g1630_n;
  wire g1631_p;
  wire g1631_n;
  wire g1632_p;
  wire g1632_n;
  wire g1633_p;
  wire g1633_n;
  wire g1634_p;
  wire g1634_n;
  wire g1635_p;
  wire g1635_n;
  wire g1636_p;
  wire g1636_n;
  wire g1637_p;
  wire g1637_n;
  wire g1638_p;
  wire g1638_n;
  wire g1639_p;
  wire g1639_n;
  wire g1640_p;
  wire g1640_n;
  wire g1641_p;
  wire g1641_n;
  wire g1642_p;
  wire g1642_n;
  wire g1643_p;
  wire g1643_n;
  wire g1644_p;
  wire g1644_n;
  wire g1645_p;
  wire g1645_n;
  wire g1646_p;
  wire g1646_n;
  wire g1647_p;
  wire g1647_n;
  wire g1648_p;
  wire g1648_n;
  wire g1649_p;
  wire g1649_n;
  wire g1650_p;
  wire g1650_n;
  wire g1651_p;
  wire g1651_n;
  wire g1652_p;
  wire g1652_n;
  wire g1653_p;
  wire g1653_n;
  wire g1654_p;
  wire g1654_n;
  wire g1655_p;
  wire g1655_n;
  wire g1656_p;
  wire g1656_n;
  wire g1657_p;
  wire g1657_n;
  wire g1658_p;
  wire g1658_n;
  wire g1659_p;
  wire g1659_n;
  wire g1660_p;
  wire g1660_n;
  wire g1661_p;
  wire g1661_n;
  wire g1662_p;
  wire g1662_n;
  wire g1663_p;
  wire g1663_n;
  wire g1664_p;
  wire g1664_n;
  wire g1665_p;
  wire g1665_n;
  wire g1666_p;
  wire g1666_n;
  wire g1667_p;
  wire g1667_n;
  wire g1668_p;
  wire g1668_n;
  wire g1669_p;
  wire g1669_n;
  wire g1670_p;
  wire g1670_n;
  wire g1671_p;
  wire g1671_n;
  wire g1672_p;
  wire g1672_n;
  wire g1673_p;
  wire g1673_n;
  wire g1674_p;
  wire g1674_n;
  wire g1675_p;
  wire g1675_n;
  wire g1676_p;
  wire g1676_n;
  wire g1677_p;
  wire g1677_n;
  wire g1678_p;
  wire g1678_n;
  wire g1679_p;
  wire g1679_n;
  wire g1680_p;
  wire g1680_n;
  wire g1681_p;
  wire g1681_n;
  wire g1682_p;
  wire g1682_n;
  wire g1683_p;
  wire g1683_n;
  wire g1684_p;
  wire g1684_n;
  wire g1685_p;
  wire g1685_n;
  wire g1686_p;
  wire g1686_n;
  wire g1687_p;
  wire g1687_n;
  wire g1688_p;
  wire g1688_n;
  wire g1689_p;
  wire g1689_n;
  wire g1690_p;
  wire g1690_n;
  wire g1691_p;
  wire g1691_n;
  wire g1692_p;
  wire g1692_n;
  wire g1693_p;
  wire g1693_n;
  wire g1694_p;
  wire g1694_n;
  wire g1695_p;
  wire g1695_n;
  wire g1696_p;
  wire g1696_n;
  wire g1697_p;
  wire g1697_n;
  wire g1698_p;
  wire g1698_n;
  wire g1699_p;
  wire g1699_n;
  wire g1700_p;
  wire g1700_n;
  wire g1701_p;
  wire g1701_n;
  wire g1702_p;
  wire g1702_n;
  wire g1703_p;
  wire g1703_n;
  wire g1704_p;
  wire g1704_n;
  wire g1705_p;
  wire g1705_n;
  wire g1706_p;
  wire g1706_n;
  wire g1707_p;
  wire g1707_n;
  wire g1708_p;
  wire g1708_n;
  wire g1709_p;
  wire g1709_n;
  wire g1710_p;
  wire g1710_n;
  wire g1711_p;
  wire g1711_n;
  wire g1712_p;
  wire g1712_n;
  wire g1713_p;
  wire g1713_n;
  wire g1714_p;
  wire g1714_n;
  wire g1715_p;
  wire g1715_n;
  wire g1716_p;
  wire g1716_n;
  wire g1717_p;
  wire g1717_n;
  wire g1718_p;
  wire g1718_n;
  wire g1719_p;
  wire g1719_n;
  wire g1720_p;
  wire g1720_n;
  wire g1721_p;
  wire g1721_n;
  wire g1722_p;
  wire g1722_n;
  wire g1723_p;
  wire g1723_n;
  wire g1724_p;
  wire g1724_n;
  wire g1725_p;
  wire g1725_n;
  wire g1726_p;
  wire g1726_n;
  wire g1727_p;
  wire g1727_n;
  wire g1728_p;
  wire g1728_n;
  wire g1729_p;
  wire g1729_n;
  wire g1730_p;
  wire g1730_n;
  wire g1731_p;
  wire g1731_n;
  wire g1732_p;
  wire g1732_n;
  wire g1733_p;
  wire g1733_n;
  wire g1734_p;
  wire g1734_n;
  wire g1735_p;
  wire g1735_n;
  wire g1736_p;
  wire g1736_n;
  wire g1737_p;
  wire g1737_n;
  wire g1738_p;
  wire g1738_n;
  wire g1739_p;
  wire g1739_n;
  wire g1740_p;
  wire g1740_n;
  wire g1741_p;
  wire g1741_n;
  wire g1742_p;
  wire g1742_n;
  wire g1743_p;
  wire g1743_n;
  wire g1744_p;
  wire g1744_n;
  wire g1745_p;
  wire g1745_n;
  wire g1746_p;
  wire g1746_n;
  wire g1747_p;
  wire g1747_n;
  wire g1748_p;
  wire g1748_n;
  wire g1749_p;
  wire g1749_n;
  wire g1750_p;
  wire g1750_n;
  wire g1751_p;
  wire g1751_n;
  wire g1752_p;
  wire g1752_n;
  wire g1753_p;
  wire g1753_n;
  wire g1754_p;
  wire g1754_n;
  wire g1755_p;
  wire g1755_n;
  wire g1756_p;
  wire g1756_n;
  wire g1757_p;
  wire g1757_n;
  wire g1758_p;
  wire g1758_n;
  wire g1759_p;
  wire g1759_n;
  wire g1760_p;
  wire g1760_n;
  wire g1761_p;
  wire g1761_n;
  wire g1762_p;
  wire g1762_n;
  wire g1763_p;
  wire g1763_n;
  wire g1764_p;
  wire g1764_n;
  wire g1765_p;
  wire g1765_n;
  wire g1766_p;
  wire g1766_n;
  wire g1767_p;
  wire g1767_n;
  wire g1768_p;
  wire g1768_n;
  wire g1769_p;
  wire g1769_n;
  wire g1770_p;
  wire g1770_n;
  wire g1771_p;
  wire g1771_n;
  wire g1772_p;
  wire g1772_n;
  wire g1773_p;
  wire g1773_n;
  wire g1774_p;
  wire g1774_n;
  wire g1775_p;
  wire g1775_n;
  wire g1776_p;
  wire g1776_n;
  wire g1777_p;
  wire g1777_n;
  wire g1778_p;
  wire g1778_n;
  wire g1779_p;
  wire g1779_n;
  wire g1780_p;
  wire g1780_n;
  wire g1781_p;
  wire g1781_n;
  wire g1782_p;
  wire g1782_n;
  wire g1783_p;
  wire g1783_n;
  wire g1784_p;
  wire g1784_n;
  wire g1785_p;
  wire g1785_n;
  wire g1786_p;
  wire g1786_n;
  wire g1787_p;
  wire g1787_n;
  wire g1788_p;
  wire g1788_n;
  wire g1789_p;
  wire g1789_n;
  wire g1790_p;
  wire g1790_n;
  wire g1791_p;
  wire g1791_n;
  wire g1792_p;
  wire g1792_n;
  wire g1793_p;
  wire g1793_n;
  wire g1794_p;
  wire g1794_n;
  wire g1795_p;
  wire g1795_n;
  wire g1796_p;
  wire g1796_n;
  wire g1797_p;
  wire g1797_n;
  wire g1798_p;
  wire g1798_n;
  wire g1799_p;
  wire g1799_n;
  wire g1800_p;
  wire g1800_n;
  wire g1801_p;
  wire g1801_n;
  wire g1802_p;
  wire g1802_n;
  wire g1803_p;
  wire g1803_n;
  wire g1804_p;
  wire g1804_n;
  wire g1805_p;
  wire g1805_n;
  wire g1806_p;
  wire g1806_n;
  wire g1807_p;
  wire g1807_n;
  wire g1808_p;
  wire g1808_n;
  wire g1809_p;
  wire g1809_n;
  wire g1810_p;
  wire g1810_n;
  wire g1811_p;
  wire g1811_n;
  wire g1812_p;
  wire g1812_n;
  wire g1813_p;
  wire g1813_n;
  wire g1814_p;
  wire g1814_n;
  wire g1815_p;
  wire g1815_n;
  wire g1816_p;
  wire g1816_n;
  wire g1817_p;
  wire g1817_n;
  wire g1818_p;
  wire g1818_n;
  wire g1819_p;
  wire g1819_n;
  wire g1820_p;
  wire g1820_n;
  wire g1821_p;
  wire g1821_n;
  wire g1822_p;
  wire g1822_n;
  wire g1823_p;
  wire g1823_n;
  wire g1824_p;
  wire g1824_n;
  wire g1825_p;
  wire g1825_n;
  wire g1826_p;
  wire g1826_n;
  wire g1827_p;
  wire g1827_n;
  wire g1828_p;
  wire g1828_n;
  wire g1829_p;
  wire g1829_n;
  wire g1830_p;
  wire g1830_n;
  wire g1831_p;
  wire g1831_n;
  wire g1832_p;
  wire g1832_n;
  wire g1833_p;
  wire g1833_n;
  wire g1834_p;
  wire g1834_n;
  wire g1835_p;
  wire g1835_n;
  wire g1836_p;
  wire g1836_n;
  wire g1837_p;
  wire g1837_n;
  wire g1838_p;
  wire g1838_n;
  wire g1839_p;
  wire g1839_n;
  wire g1840_p;
  wire g1840_n;
  wire g1841_p;
  wire g1841_n;
  wire g1842_p;
  wire g1842_n;
  wire g1843_p;
  wire g1843_n;
  wire g1844_p;
  wire g1844_n;
  wire g1845_p;
  wire g1845_n;
  wire g1846_p;
  wire g1846_n;
  wire g1847_p;
  wire g1847_n;
  wire g1848_p;
  wire g1848_n;
  wire g1849_p;
  wire g1849_n;
  wire g1850_p;
  wire g1850_n;
  wire g1851_p;
  wire g1851_n;
  wire g1852_p;
  wire g1852_n;
  wire g1853_p;
  wire g1853_n;
  wire g1854_p;
  wire g1854_n;
  wire g1855_p;
  wire g1855_n;
  wire g1856_p;
  wire g1856_n;
  wire g1857_p;
  wire g1857_n;
  wire g1858_p;
  wire g1858_n;
  wire g1859_p;
  wire g1859_n;
  wire g1860_p;
  wire g1860_n;
  wire g1861_p;
  wire g1861_n;
  wire g1862_p;
  wire g1862_n;
  wire g1863_p;
  wire g1863_n;
  wire g1864_p;
  wire g1864_n;
  wire g1865_p;
  wire g1865_n;
  wire g1866_p;
  wire g1866_n;
  wire g1867_p;
  wire g1867_n;
  wire g1868_p;
  wire g1868_n;
  wire g1869_p;
  wire g1869_n;
  wire g1870_p;
  wire g1870_n;
  wire g1871_p;
  wire g1871_n;
  wire g1872_p;
  wire g1872_n;
  wire g1873_p;
  wire g1873_n;
  wire g1874_p;
  wire g1874_n;
  wire g1875_p;
  wire g1875_n;
  wire g1876_p;
  wire g1876_n;
  wire g1877_p;
  wire g1877_n;
  wire g1878_p;
  wire g1878_n;
  wire g1879_p;
  wire g1879_n;
  wire g1880_p;
  wire g1880_n;
  wire g1881_p;
  wire g1881_n;
  wire g1882_p;
  wire g1882_n;
  wire g1883_p;
  wire g1883_n;
  wire g1884_p;
  wire g1884_n;
  wire g1885_p;
  wire g1885_n;
  wire g1886_p;
  wire g1886_n;
  wire g1887_p;
  wire g1887_n;
  wire g1888_p;
  wire g1888_n;
  wire g1889_p;
  wire g1889_n;
  wire g1890_p;
  wire g1890_n;
  wire g1891_p;
  wire g1891_n;
  wire g1892_p;
  wire g1892_n;
  wire g1893_p;
  wire g1893_n;
  wire g1894_p;
  wire g1894_n;
  wire g1895_p;
  wire g1895_n;
  wire g1896_p;
  wire g1896_n;
  wire g1897_p;
  wire g1897_n;
  wire g1898_p;
  wire g1898_n;
  wire g1899_p;
  wire g1899_n;
  wire g1900_p;
  wire g1900_n;
  wire g1901_p;
  wire g1901_n;
  wire g1902_p;
  wire g1902_n;
  wire g1903_p;
  wire g1903_n;
  wire g1904_p;
  wire g1904_n;
  wire g1905_p;
  wire g1905_n;
  wire g1906_p;
  wire g1906_n;
  wire g1907_p;
  wire g1907_n;
  wire g1908_p;
  wire g1908_n;
  wire g1909_p;
  wire g1909_n;
  wire g1910_p;
  wire g1910_n;
  wire g1911_p;
  wire g1911_n;
  wire g1912_p;
  wire g1912_n;
  wire g1913_p;
  wire g1913_n;
  wire g1914_p;
  wire g1914_n;
  wire g1915_p;
  wire g1915_n;
  wire g1916_p;
  wire g1916_n;
  wire g1917_p;
  wire g1917_n;
  wire g1918_p;
  wire g1918_n;
  wire g1919_p;
  wire g1919_n;
  wire g1920_p;
  wire g1920_n;
  wire g1921_p;
  wire g1921_n;
  wire g1922_p;
  wire g1922_n;
  wire g1923_p;
  wire g1923_n;
  wire g1924_p;
  wire g1924_n;
  wire g1925_p;
  wire g1925_n;
  wire g1926_p;
  wire g1926_n;
  wire g1927_p;
  wire g1927_n;
  wire g1928_p;
  wire g1928_n;
  wire g1929_p;
  wire g1929_n;
  wire g1930_p;
  wire g1930_n;
  wire g1931_p;
  wire g1931_n;
  wire g1932_p;
  wire g1932_n;
  wire g1933_p;
  wire g1933_n;
  wire g1934_p;
  wire g1934_n;
  wire g1935_p;
  wire g1935_n;
  wire g1936_p;
  wire g1936_n;
  wire g1937_p;
  wire g1937_n;
  wire g1938_p;
  wire g1938_n;
  wire g1939_p;
  wire g1939_n;
  wire g1940_p;
  wire g1940_n;
  wire g1941_p;
  wire g1941_n;
  wire g1942_p;
  wire g1942_n;
  wire g1943_p;
  wire g1943_n;
  wire g1944_p;
  wire g1944_n;
  wire g1945_p;
  wire g1945_n;
  wire g1946_p;
  wire g1946_n;
  wire g1947_p;
  wire g1947_n;
  wire g1948_p;
  wire g1948_n;
  wire g1949_p;
  wire g1949_n;
  wire g1950_p;
  wire g1950_n;
  wire g1951_p;
  wire g1951_n;
  wire g1952_p;
  wire g1952_n;
  wire g1953_p;
  wire g1953_n;
  wire g1954_p;
  wire g1954_n;
  wire g1955_p;
  wire g1955_n;
  wire g1956_p;
  wire g1956_n;
  wire g1957_p;
  wire g1957_n;
  wire g1958_p;
  wire g1958_n;
  wire g1959_p;
  wire g1959_n;
  wire g1960_p;
  wire g1960_n;
  wire g1961_p;
  wire g1961_n;
  wire g1962_p;
  wire g1962_n;
  wire g1963_p;
  wire g1963_n;
  wire g1964_p;
  wire g1964_n;
  wire g1965_p;
  wire g1965_n;
  wire g1966_p;
  wire g1966_n;
  wire g1967_p;
  wire g1967_n;
  wire g1968_p;
  wire g1968_n;
  wire g1969_p;
  wire g1969_n;
  wire g1970_p;
  wire g1970_n;
  wire g1971_p;
  wire g1971_n;
  wire g1972_p;
  wire g1972_n;
  wire g1973_p;
  wire g1973_n;
  wire g1974_p;
  wire g1974_n;
  wire g1975_p;
  wire g1975_n;
  wire g1976_p;
  wire g1976_n;
  wire g1977_p;
  wire g1977_n;
  wire g1978_p;
  wire g1978_n;
  wire g1979_p;
  wire g1979_n;
  wire g1980_p;
  wire g1980_n;
  wire g1981_p;
  wire g1981_n;
  wire g1982_p;
  wire g1982_n;
  wire g1983_p;
  wire g1983_n;
  wire g1984_p;
  wire g1984_n;
  wire g1985_p;
  wire g1985_n;
  wire g1986_p;
  wire g1986_n;
  wire g1987_p;
  wire g1987_n;
  wire g1988_p;
  wire g1988_n;
  wire g1989_p;
  wire g1989_n;
  wire g1990_p;
  wire g1990_n;
  wire g1991_p;
  wire g1991_n;
  wire g1992_p;
  wire g1992_n;
  wire g1993_p;
  wire g1993_n;
  wire g1994_p;
  wire g1994_n;
  wire g1995_p;
  wire g1995_n;
  wire g1996_p;
  wire g1996_n;
  wire g1997_p;
  wire g1997_n;
  wire g1998_p;
  wire g1998_n;
  wire g1999_p;
  wire g1999_n;
  wire g2000_p;
  wire g2000_n;
  wire g2001_p;
  wire g2001_n;
  wire g2002_p;
  wire g2002_n;
  wire g2003_p;
  wire g2003_n;
  wire g2004_p;
  wire g2004_n;
  wire g2005_p;
  wire g2005_n;
  wire g2006_p;
  wire g2006_n;
  wire g2007_p;
  wire g2007_n;
  wire g2008_p;
  wire g2008_n;
  wire g2009_p;
  wire g2009_n;
  wire g2010_p;
  wire g2010_n;
  wire g2011_p;
  wire g2011_n;
  wire g2012_p;
  wire g2012_n;
  wire g2013_p;
  wire g2013_n;
  wire g2014_p;
  wire g2014_n;
  wire g2015_p;
  wire g2015_n;
  wire g2016_p;
  wire g2016_n;
  wire g2017_p;
  wire g2017_n;
  wire g2018_p;
  wire g2018_n;
  wire g2019_p;
  wire g2019_n;
  wire g2020_p;
  wire g2020_n;
  wire g2021_p;
  wire g2021_n;
  wire g2022_p;
  wire g2022_n;
  wire g2023_p;
  wire g2023_n;
  wire g2024_p;
  wire g2024_n;
  wire g2025_p;
  wire g2025_n;
  wire g2026_p;
  wire g2026_n;
  wire g2027_p;
  wire g2027_n;
  wire g2028_p;
  wire g2028_n;
  wire g2029_p;
  wire g2029_n;
  wire g2030_p;
  wire g2030_n;
  wire g2031_p;
  wire g2031_n;
  wire g2032_p;
  wire g2032_n;
  wire g2033_p;
  wire g2033_n;
  wire g2034_p;
  wire g2034_n;
  wire g2035_p;
  wire g2035_n;
  wire g2036_p;
  wire g2036_n;
  wire g2037_p;
  wire g2037_n;
  wire g2038_p;
  wire g2038_n;
  wire g2039_p;
  wire g2039_n;
  wire g2040_p;
  wire g2040_n;
  wire g2041_p;
  wire g2041_n;
  wire g2042_p;
  wire g2042_n;
  wire g2043_p;
  wire g2043_n;
  wire g2044_p;
  wire g2044_n;
  wire g2045_p;
  wire g2045_n;
  wire g2046_p;
  wire g2046_n;
  wire g2047_p;
  wire g2047_n;
  wire g2048_p;
  wire g2048_n;
  wire g2049_p;
  wire g2049_n;
  wire g2050_p;
  wire g2050_n;
  wire g2051_p;
  wire g2051_n;
  wire g2052_p;
  wire g2052_n;
  wire g2053_p;
  wire g2053_n;
  wire g2054_p;
  wire g2054_n;
  wire g2055_p;
  wire g2055_n;
  wire g2056_p;
  wire g2056_n;
  wire g2057_p;
  wire g2057_n;
  wire g2058_p;
  wire g2058_n;
  wire g2059_p;
  wire g2059_n;
  wire g2060_p;
  wire g2060_n;
  wire g2061_p;
  wire g2061_n;
  wire g2062_p;
  wire g2062_n;
  wire g2063_p;
  wire g2063_n;
  wire g2064_p;
  wire g2064_n;
  wire g2065_p;
  wire g2065_n;
  wire g2066_p;
  wire g2066_n;
  wire g2067_p;
  wire g2067_n;
  wire g2068_p;
  wire g2068_n;
  wire g2069_p;
  wire g2069_n;
  wire g2070_p;
  wire g2070_n;
  wire g2071_p;
  wire g2071_n;
  wire g2072_p;
  wire g2072_n;
  wire g2073_p;
  wire g2073_n;
  wire g2074_p;
  wire g2074_n;
  wire g2075_p;
  wire g2075_n;
  wire g2076_p;
  wire g2076_n;
  wire g2077_p;
  wire g2077_n;
  wire g2078_p;
  wire g2078_n;
  wire g2079_p;
  wire g2079_n;
  wire g2080_p;
  wire g2080_n;
  wire g2081_p;
  wire g2081_n;
  wire g2082_p;
  wire g2082_n;
  wire g2083_p;
  wire g2083_n;
  wire g2084_p;
  wire g2084_n;
  wire g2085_p;
  wire g2085_n;
  wire g2086_p;
  wire g2086_n;
  wire g2087_p;
  wire g2087_n;
  wire g2088_p;
  wire g2088_n;
  wire g2089_p;
  wire g2089_n;
  wire g2090_p;
  wire g2090_n;
  wire g2091_p;
  wire g2091_n;
  wire g2092_p;
  wire g2092_n;
  wire g2093_p;
  wire g2093_n;
  wire g2094_p;
  wire g2094_n;
  wire g2095_p;
  wire g2095_n;
  wire g2096_p;
  wire g2096_n;
  wire g2097_p;
  wire g2097_n;
  wire g2098_p;
  wire g2098_n;
  wire g2099_p;
  wire g2099_n;
  wire g2100_p;
  wire g2100_n;
  wire g2101_p;
  wire g2101_n;
  wire g2102_p;
  wire g2102_n;
  wire g2103_p;
  wire g2103_n;
  wire g2104_p;
  wire g2104_n;
  wire g2105_p;
  wire g2105_n;
  wire g2106_p;
  wire g2106_n;
  wire g2107_p;
  wire g2107_n;
  wire g2108_p;
  wire g2108_n;
  wire g2109_p;
  wire g2109_n;
  wire g2110_p;
  wire g2110_n;
  wire g2111_p;
  wire g2111_n;
  wire g2112_p;
  wire g2112_n;
  wire g2113_p;
  wire g2113_n;
  wire g2114_p;
  wire g2114_n;
  wire g2115_p;
  wire g2115_n;
  wire g2116_p;
  wire g2116_n;
  wire g2117_p;
  wire g2117_n;
  wire g2118_p;
  wire g2118_n;
  wire g2119_p;
  wire g2119_n;
  wire g2120_p;
  wire g2120_n;
  wire g2121_p;
  wire g2121_n;
  wire g2122_p;
  wire g2122_n;
  wire g2123_p;
  wire g2123_n;
  wire g2124_p;
  wire g2124_n;
  wire g2125_p;
  wire g2125_n;
  wire g2126_p;
  wire g2126_n;
  wire g2127_p;
  wire g2127_n;
  wire g2128_p;
  wire g2128_n;
  wire g2129_p;
  wire g2129_n;
  wire g2130_p;
  wire g2130_n;
  wire g2131_p;
  wire g2131_n;
  wire g2132_p;
  wire g2132_n;
  wire g2133_p;
  wire g2133_n;
  wire g2134_p;
  wire g2134_n;
  wire g2135_p;
  wire g2135_n;
  wire g2136_p;
  wire g2136_n;
  wire g2137_p;
  wire g2137_n;
  wire g2138_p;
  wire g2138_n;
  wire g2139_p;
  wire g2139_n;
  wire g2140_p;
  wire g2140_n;
  wire g2141_p;
  wire g2141_n;
  wire g2142_p;
  wire g2142_n;
  wire g2143_p;
  wire g2143_n;
  wire g2144_p;
  wire g2144_n;
  wire g2145_p;
  wire g2145_n;
  wire g2146_p;
  wire g2146_n;
  wire g2147_p;
  wire g2147_n;
  wire g2148_p;
  wire g2148_n;
  wire g2149_p;
  wire g2149_n;
  wire g2150_p;
  wire g2150_n;
  wire g2151_p;
  wire g2151_n;
  wire g2152_p;
  wire g2152_n;
  wire g2153_p;
  wire g2153_n;
  wire g2154_p;
  wire g2154_n;
  wire g2155_p;
  wire g2155_n;
  wire g2156_p;
  wire g2156_n;
  wire g2157_p;
  wire g2157_n;
  wire g2158_p;
  wire g2158_n;
  wire g2159_p;
  wire g2159_n;
  wire g2160_p;
  wire g2160_n;
  wire g2161_p;
  wire g2161_n;
  wire g2162_p;
  wire g2162_n;
  wire g2163_p;
  wire g2163_n;
  wire g2164_p;
  wire g2164_n;
  wire g2165_p;
  wire g2165_n;
  wire g2166_p;
  wire g2166_n;
  wire g2167_p;
  wire g2167_n;
  wire g2168_p;
  wire g2168_n;
  wire g2169_p;
  wire g2169_n;
  wire g2170_p;
  wire g2170_n;
  wire g2171_p;
  wire g2171_n;
  wire g2172_p;
  wire g2172_n;
  wire g2173_p;
  wire g2173_n;
  wire g2174_p;
  wire g2174_n;
  wire g2175_p;
  wire g2175_n;
  wire g2176_p;
  wire g2176_n;
  wire g2177_p;
  wire g2177_n;
  wire g2178_p;
  wire g2178_n;
  wire g2179_p;
  wire g2179_n;
  wire g2180_p;
  wire g2180_n;
  wire g2181_p;
  wire g2181_n;
  wire g2182_p;
  wire g2182_n;
  wire g2183_p;
  wire g2183_n;
  wire g2184_p;
  wire g2184_n;
  wire g2185_p;
  wire g2185_n;
  wire g2186_p;
  wire g2186_n;
  wire g2187_p;
  wire g2187_n;
  wire g2188_p;
  wire g2188_n;
  wire g2189_p;
  wire g2189_n;
  wire g2190_p;
  wire g2190_n;
  wire g2191_p;
  wire g2191_n;
  wire g2192_p;
  wire g2192_n;
  wire g2193_p;
  wire g2193_n;
  wire g2194_p;
  wire g2194_n;
  wire g2195_p;
  wire g2195_n;
  wire g2196_p;
  wire g2196_n;
  wire g2197_p;
  wire g2197_n;
  wire g2198_p;
  wire g2198_n;
  wire g2199_p;
  wire g2199_n;
  wire g2200_p;
  wire g2200_n;
  wire g2201_p;
  wire g2201_n;
  wire g2202_p;
  wire g2202_n;
  wire g2203_p;
  wire g2203_n;
  wire g2204_p;
  wire g2204_n;
  wire g2205_p;
  wire g2205_n;
  wire g2206_p;
  wire g2206_n;
  wire g2207_p;
  wire g2207_n;
  wire g2208_p;
  wire g2208_n;
  wire g2209_p;
  wire g2209_n;
  wire g2210_p;
  wire g2210_n;
  wire g2211_p;
  wire g2211_n;
  wire g2212_p;
  wire g2212_n;
  wire g2213_p;
  wire g2213_n;
  wire g2214_p;
  wire g2214_n;
  wire g2215_p;
  wire g2215_n;
  wire g2216_p;
  wire g2216_n;
  wire g2217_p;
  wire g2217_n;
  wire g2218_p;
  wire g2218_n;
  wire g2219_p;
  wire g2219_n;
  wire g2220_p;
  wire g2220_n;
  wire g2221_p;
  wire g2221_n;
  wire g2222_p;
  wire g2222_n;
  wire g2223_p;
  wire g2223_n;
  wire g2224_p;
  wire g2224_n;
  wire g2225_p;
  wire g2225_n;
  wire g2226_p;
  wire g2226_n;
  wire g2227_p;
  wire g2227_n;
  wire g2228_p;
  wire g2228_n;
  wire g2229_p;
  wire g2229_n;
  wire g2230_p;
  wire g2230_n;
  wire g2231_p;
  wire g2231_n;
  wire g2232_p;
  wire g2232_n;
  wire g2233_p;
  wire g2233_n;
  wire g2234_p;
  wire g2234_n;
  wire g2235_p;
  wire g2235_n;
  wire g2236_p;
  wire g2236_n;
  wire g2237_p;
  wire g2237_n;
  wire g2238_p;
  wire g2238_n;
  wire g2239_p;
  wire g2239_n;
  wire g2240_p;
  wire g2240_n;
  wire g2241_p;
  wire g2241_n;
  wire g2242_p;
  wire g2242_n;
  wire g2243_p;
  wire g2243_n;
  wire g2244_p;
  wire g2244_n;
  wire g2245_p;
  wire g2245_n;
  wire g2246_p;
  wire g2246_n;
  wire g2247_p;
  wire g2247_n;
  wire g2248_p;
  wire g2248_n;
  wire g2249_p;
  wire g2249_n;
  wire g2250_p;
  wire g2250_n;
  wire g2251_p;
  wire g2251_n;
  wire g2252_p;
  wire g2252_n;
  wire g2253_p;
  wire g2253_n;
  wire g2254_p;
  wire g2254_n;
  wire g2255_p;
  wire g2255_n;
  wire g2256_p;
  wire g2256_n;
  wire g2257_p;
  wire g2257_n;
  wire g2258_p;
  wire g2258_n;
  wire g2259_p;
  wire g2259_n;
  wire g2260_p;
  wire g2260_n;
  wire g2261_p;
  wire g2261_n;
  wire g2262_p;
  wire g2262_n;
  wire g2263_p;
  wire g2263_n;
  wire g2264_p;
  wire g2264_n;
  wire g2265_p;
  wire g2265_n;
  wire g2266_p;
  wire g2266_n;
  wire g2267_p;
  wire g2267_n;
  wire g2268_p;
  wire g2268_n;
  wire g2269_p;
  wire g2269_n;
  wire g2270_p;
  wire g2270_n;
  wire g2271_p;
  wire g2271_n;
  wire g2272_p;
  wire g2272_n;
  wire g2273_p;
  wire g2273_n;
  wire g2274_p;
  wire g2274_n;
  wire g2275_p;
  wire g2275_n;
  wire g2276_p;
  wire g2276_n;
  wire g2277_p;
  wire g2277_n;
  wire g2278_p;
  wire g2278_n;
  wire g2279_p;
  wire g2279_n;
  wire g2280_p;
  wire g2280_n;
  wire g2281_p;
  wire g2281_n;
  wire g2282_p;
  wire g2282_n;
  wire g2283_p;
  wire g2283_n;
  wire g2284_p;
  wire g2284_n;
  wire g2285_p;
  wire g2285_n;
  wire g2286_p;
  wire g2286_n;
  wire g2287_p;
  wire g2287_n;
  wire g2288_p;
  wire g2288_n;
  wire g2289_p;
  wire g2289_n;
  wire g2290_p;
  wire g2290_n;
  wire g2291_p;
  wire g2291_n;
  wire g2292_p;
  wire g2292_n;
  wire g2293_p;
  wire g2293_n;
  wire g2294_p;
  wire g2294_n;
  wire g2295_p;
  wire g2295_n;
  wire g2296_p;
  wire g2296_n;
  wire g2297_p;
  wire g2297_n;
  wire g2298_p;
  wire g2298_n;
  wire g2299_p;
  wire g2299_n;
  wire g2300_p;
  wire g2300_n;
  wire g2301_p;
  wire g2301_n;
  wire g2302_p;
  wire g2302_n;
  wire g2303_p;
  wire g2303_n;
  wire g2304_p;
  wire g2304_n;
  wire g2305_p;
  wire g2305_n;
  wire g2306_p;
  wire g2306_n;
  wire g2307_p;
  wire g2307_n;
  wire g2308_p;
  wire g2308_n;
  wire g2309_p;
  wire g2309_n;
  wire g2310_p;
  wire g2310_n;
  wire g2311_p;
  wire g2311_n;
  wire g2312_p;
  wire g2312_n;
  wire g2313_p;
  wire g2313_n;
  wire g2314_p;
  wire g2314_n;
  wire g2315_p;
  wire g2315_n;
  wire g2316_p;
  wire g2316_n;
  wire g2317_p;
  wire g2317_n;
  wire g2318_p;
  wire g2318_n;
  wire g2319_p;
  wire g2319_n;
  wire g2320_p;
  wire g2320_n;
  wire g2321_p;
  wire g2321_n;
  wire g2322_p;
  wire g2322_n;
  wire g2323_p;
  wire g2323_n;
  wire g2324_p;
  wire g2324_n;
  wire g2325_p;
  wire g2325_n;
  wire g2326_p;
  wire g2326_n;
  wire g2327_p;
  wire g2327_n;
  wire g2328_p;
  wire g2328_n;
  wire g2329_p;
  wire g2329_n;
  wire g2330_p;
  wire g2330_n;
  wire g2331_p;
  wire g2331_n;
  wire g2332_p;
  wire g2332_n;
  wire g2333_p;
  wire g2333_n;
  wire g2334_p;
  wire g2334_n;
  wire g2335_p;
  wire g2335_n;
  wire g2336_p;
  wire g2336_n;
  wire g2337_p;
  wire g2337_n;
  wire g2338_p;
  wire g2338_n;
  wire g2339_p;
  wire g2339_n;
  wire g2340_p;
  wire g2340_n;
  wire g2341_p;
  wire g2341_n;
  wire g2342_p;
  wire g2342_n;
  wire g2343_p;
  wire g2343_n;
  wire g2344_p;
  wire g2344_n;
  wire g2345_p;
  wire g2345_n;
  wire g2346_p;
  wire g2346_n;
  wire g2347_p;
  wire g2347_n;
  wire g2348_p;
  wire g2348_n;
  wire g2349_p;
  wire g2349_n;
  wire g2350_p;
  wire g2350_n;
  wire g2351_p;
  wire g2351_n;
  wire g2352_p;
  wire g2352_n;
  wire g2353_p;
  wire g2353_n;
  wire g2354_p;
  wire g2354_n;
  wire g2355_p;
  wire g2355_n;
  wire g2356_p;
  wire g2356_n;
  wire g2357_p;
  wire g2357_n;
  wire g2358_p;
  wire g2358_n;
  wire g2359_p;
  wire g2359_n;
  wire g2360_p;
  wire g2360_n;
  wire g2361_p;
  wire g2361_n;
  wire g2362_p;
  wire g2362_n;
  wire g2363_p;
  wire g2363_n;
  wire g2364_p;
  wire g2364_n;
  wire g2365_p;
  wire g2365_n;
  wire g2366_p;
  wire g2366_n;
  wire g2367_p;
  wire g2367_n;
  wire g2368_p;
  wire g2368_n;
  wire g2369_p;
  wire g2369_n;
  wire g2370_p;
  wire g2370_n;
  wire g2371_p;
  wire g2371_n;
  wire g2372_p;
  wire g2372_n;
  wire g2373_p;
  wire g2373_n;
  wire g2374_p;
  wire g2374_n;
  wire g2375_p;
  wire g2375_n;
  wire g2376_p;
  wire g2376_n;
  wire g2377_p;
  wire g2377_n;
  wire g2378_p;
  wire g2378_n;
  wire g2379_p;
  wire g2379_n;
  wire g2380_p;
  wire g2380_n;
  wire g2381_p;
  wire g2381_n;
  wire g2382_p;
  wire g2382_n;
  wire g2383_p;
  wire g2383_n;
  wire g2384_p;
  wire g2384_n;
  wire g2385_p;
  wire g2385_n;
  wire g2386_p;
  wire g2386_n;
  wire g2387_p;
  wire g2387_n;
  wire g2388_p;
  wire g2388_n;
  wire g2389_p;
  wire g2389_n;
  wire g2390_p;
  wire g2390_n;
  wire g2391_p;
  wire g2391_n;
  wire g2392_p;
  wire g2392_n;
  wire g2393_p;
  wire g2393_n;
  wire g2394_p;
  wire g2394_n;
  wire g2395_p;
  wire g2395_n;
  wire g2396_p;
  wire g2396_n;
  wire g2397_p;
  wire g2397_n;
  wire g2398_p;
  wire g2398_n;
  wire g2399_p;
  wire g2399_n;
  wire g2400_p;
  wire g2400_n;
  wire g2401_p;
  wire g2401_n;
  wire g2402_p;
  wire g2402_n;
  wire g2403_p;
  wire g2403_n;
  wire g2404_p;
  wire g2404_n;
  wire g2405_p;
  wire g2405_n;
  wire g2406_p;
  wire g2406_n;
  wire g2407_p;
  wire g2407_n;
  wire g2408_p;
  wire g2408_n;
  wire g2409_p;
  wire g2409_n;
  wire g2410_p;
  wire g2410_n;
  wire g2411_p;
  wire g2411_n;
  wire g2412_p;
  wire g2412_n;
  wire g2413_p;
  wire g2413_n;
  wire g2414_p;
  wire g2414_n;
  wire g2415_p;
  wire g2415_n;
  wire g2416_p;
  wire g2416_n;
  wire g2417_p;
  wire g2417_n;
  wire g2418_p;
  wire g2418_n;
  wire g2419_p;
  wire g2419_n;
  wire g2420_p;
  wire g2420_n;
  wire g2421_p;
  wire g2421_n;
  wire g2422_p;
  wire g2422_n;
  wire g2423_p;
  wire g2423_n;
  wire g2424_p;
  wire g2424_n;
  wire g2425_p;
  wire g2425_n;
  wire g2426_p;
  wire g2426_n;
  wire g2427_p;
  wire g2427_n;
  wire g2428_p;
  wire g2428_n;
  wire g2429_p;
  wire g2429_n;
  wire g2430_p;
  wire g2430_n;
  wire g2431_p;
  wire g2431_n;
  wire g2432_p;
  wire g2432_n;
  wire g2433_p;
  wire g2433_n;
  wire g2434_p;
  wire g2434_n;
  wire g2435_p;
  wire g2435_n;
  wire g2436_p;
  wire g2436_n;
  wire g2437_p;
  wire g2437_n;
  wire g2438_p;
  wire g2438_n;
  wire g2439_p;
  wire g2439_n;
  wire g2440_p;
  wire g2440_n;
  wire g2441_p;
  wire g2441_n;
  wire g2442_p;
  wire g2442_n;
  wire g2443_p;
  wire g2443_n;
  wire g2444_p;
  wire g2444_n;
  wire g2445_p;
  wire g2445_n;
  wire g2446_p;
  wire g2446_n;
  wire g2447_p;
  wire g2447_n;
  wire g2448_p;
  wire g2448_n;
  wire g2449_p;
  wire g2449_n;
  wire g2450_p;
  wire g2450_n;
  wire g2451_p;
  wire g2451_n;
  wire g2452_p;
  wire g2452_n;
  wire g2453_p;
  wire g2453_n;
  wire g2454_p;
  wire g2454_n;
  wire g2455_p;
  wire g2455_n;
  wire g2456_p;
  wire g2456_n;
  wire g2457_p;
  wire g2457_n;
  wire g2458_p;
  wire g2458_n;
  wire g2459_p;
  wire g2459_n;
  wire g2460_p;
  wire g2460_n;
  wire g2461_p;
  wire g2461_n;
  wire g2462_p;
  wire g2462_n;
  wire g2463_p;
  wire g2463_n;
  wire g2464_p;
  wire g2464_n;
  wire g2465_p;
  wire g2465_n;
  wire g2466_p;
  wire g2466_n;
  wire g2467_p;
  wire g2467_n;
  wire g2468_p;
  wire g2468_n;
  wire g2469_p;
  wire g2469_n;
  wire g2470_p;
  wire g2470_n;
  wire g2471_p;
  wire g2471_n;
  wire g2472_p;
  wire g2472_n;
  wire g2473_p;
  wire g2473_n;
  wire g2474_p;
  wire g2474_n;
  wire g2475_p;
  wire g2475_n;
  wire g2476_p;
  wire g2476_n;
  wire g2477_p;
  wire g2477_n;
  wire g2478_p;
  wire g2478_n;
  wire g2479_p;
  wire g2479_n;
  wire g2480_p;
  wire g2480_n;
  wire g2481_p;
  wire g2481_n;
  wire g2482_p;
  wire g2482_n;
  wire g2483_p;
  wire g2483_n;
  wire g2484_p;
  wire g2484_n;
  wire g2485_p;
  wire g2485_n;
  wire g2486_p;
  wire g2486_n;
  wire g2487_p;
  wire g2487_n;
  wire g2488_p;
  wire g2488_n;
  wire g2489_p;
  wire g2489_n;
  wire g2490_p;
  wire g2490_n;
  wire g2491_p;
  wire g2491_n;
  wire g2492_p;
  wire g2492_n;
  wire g2493_p;
  wire g2493_n;
  wire g2494_p;
  wire g2494_n;
  wire g2495_p;
  wire g2495_n;
  wire g2496_p;
  wire g2496_n;
  wire g2497_p;
  wire g2497_n;
  wire g2498_p;
  wire g2498_n;
  wire g2499_p;
  wire g2499_n;
  wire g2500_p;
  wire g2500_n;
  wire g2501_p;
  wire g2501_n;
  wire g2502_p;
  wire g2502_n;
  wire g2503_p;
  wire g2503_n;
  wire g2504_p;
  wire g2504_n;
  wire g2505_p;
  wire g2505_n;
  wire g2506_p;
  wire g2506_n;
  wire g2507_p;
  wire g2507_n;
  wire g2508_p;
  wire g2508_n;
  wire g2509_p;
  wire g2509_n;
  wire g2510_p;
  wire g2510_n;
  wire g2511_p;
  wire g2511_n;
  wire g2512_p;
  wire g2512_n;
  wire g2513_p;
  wire g2513_n;
  wire g2514_p;
  wire g2514_n;
  wire g2515_p;
  wire g2515_n;
  wire g2516_p;
  wire g2516_n;
  wire g2517_p;
  wire g2517_n;
  wire g2518_p;
  wire g2518_n;
  wire g2519_p;
  wire g2519_n;
  wire g2520_p;
  wire g2520_n;
  wire g2521_p;
  wire g2521_n;
  wire g2522_p;
  wire g2522_n;
  wire g2523_p;
  wire g2523_n;
  wire g2524_p;
  wire g2524_n;
  wire g2525_p;
  wire g2525_n;
  wire g2526_p;
  wire g2526_n;
  wire g2527_p;
  wire g2527_n;
  wire g2528_p;
  wire g2528_n;
  wire g2529_p;
  wire g2529_n;
  wire g2530_p;
  wire g2530_n;
  wire g2531_p;
  wire g2531_n;
  wire g2532_p;
  wire g2532_n;
  wire g2533_p;
  wire g2533_n;
  wire g2534_p;
  wire g2534_n;
  wire g2535_p;
  wire g2535_n;
  wire g2536_p;
  wire g2536_n;
  wire g2537_p;
  wire g2537_n;
  wire g2538_p;
  wire g2538_n;
  wire g2539_p;
  wire g2539_n;
  wire g2540_p;
  wire g2540_n;
  wire g2541_p;
  wire g2541_n;
  wire g2542_p;
  wire g2542_n;
  wire g2543_p;
  wire g2543_n;
  wire g2544_p;
  wire g2544_n;
  wire g2545_p;
  wire g2545_n;
  wire g2546_p;
  wire g2546_n;
  wire g2547_p;
  wire g2547_n;
  wire g2548_p;
  wire g2548_n;
  wire g2549_p;
  wire g2549_n;
  wire g2550_p;
  wire g2550_n;
  wire g2551_p;
  wire g2551_n;
  wire g2552_p;
  wire g2552_n;
  wire g2553_p;
  wire g2553_n;
  wire g2554_p;
  wire g2554_n;
  wire g2555_p;
  wire g2555_n;
  wire g2556_p;
  wire g2556_n;
  wire g2557_p;
  wire g2557_n;
  wire g2558_p;
  wire g2558_n;
  wire g2559_p;
  wire g2559_n;
  wire g2560_p;
  wire g2560_n;
  wire g2561_p;
  wire g2561_n;
  wire g2562_p;
  wire g2562_n;
  wire g2563_p;
  wire g2563_n;
  wire g2564_p;
  wire g2564_n;
  wire g2565_p;
  wire g2565_n;
  wire g2566_p;
  wire g2566_n;
  wire g2567_p;
  wire g2567_n;
  wire g2568_p;
  wire g2568_n;
  wire g2569_p;
  wire g2569_n;
  wire g2570_p;
  wire g2570_n;
  wire g2571_p;
  wire g2571_n;
  wire g2572_p;
  wire g2572_n;
  wire g2573_p;
  wire g2573_n;
  wire g2574_p;
  wire g2574_n;
  wire g2575_p;
  wire g2575_n;
  wire g2576_p;
  wire g2576_n;
  wire g2577_p;
  wire g2577_n;
  wire g2578_p;
  wire g2578_n;
  wire g2579_p;
  wire g2579_n;
  wire g2580_p;
  wire g2580_n;
  wire g2581_p;
  wire g2581_n;
  wire g2582_p;
  wire g2582_n;
  wire g2583_p;
  wire g2583_n;
  wire g2584_p;
  wire g2584_n;
  wire g2585_p;
  wire g2585_n;
  wire g2586_p;
  wire g2586_n;
  wire g2587_p;
  wire g2587_n;
  wire g2588_p;
  wire g2588_n;
  wire g2589_p;
  wire g2589_n;
  wire g2590_p;
  wire g2590_n;
  wire g2591_p;
  wire g2591_n;
  wire g2592_p;
  wire g2592_n;
  wire g2593_p;
  wire g2593_n;
  wire g2594_p;
  wire g2594_n;
  wire g2595_p;
  wire g2595_n;
  wire g2596_p;
  wire g2596_n;
  wire g2597_p;
  wire g2597_n;
  wire g2598_p;
  wire g2598_n;
  wire g2599_p;
  wire g2599_n;
  wire g2600_p;
  wire g2600_n;
  wire g2601_p;
  wire g2601_n;
  wire g2602_p;
  wire g2602_n;
  wire g2603_p;
  wire g2603_n;
  wire g2604_p;
  wire g2604_n;
  wire g2605_p;
  wire g2605_n;
  wire g2606_p;
  wire g2606_n;
  wire g2607_p;
  wire g2607_n;
  wire g2608_p;
  wire g2608_n;
  wire g2609_p;
  wire g2609_n;
  wire g2610_p;
  wire g2610_n;
  wire g2611_p;
  wire g2611_n;
  wire g2612_p;
  wire g2612_n;
  wire g2613_p;
  wire g2613_n;
  wire g2614_p;
  wire g2614_n;
  wire g2615_p;
  wire g2615_n;
  wire g2616_p;
  wire g2616_n;
  wire g2617_p;
  wire g2617_n;
  wire g2618_p;
  wire g2618_n;
  wire g2619_p;
  wire g2619_n;
  wire g2620_p;
  wire g2620_n;
  wire g2621_p;
  wire g2621_n;
  wire g2622_p;
  wire g2622_n;
  wire g2623_p;
  wire g2623_n;
  wire g2624_p;
  wire g2624_n;
  wire g2625_p;
  wire g2625_n;
  wire g2626_p;
  wire g2626_n;
  wire g2627_p;
  wire g2627_n;
  wire g2628_p;
  wire g2628_n;
  wire g2629_p;
  wire g2629_n;
  wire g2630_p;
  wire g2630_n;
  wire g2631_p;
  wire g2631_n;
  wire g2632_p;
  wire g2632_n;
  wire g2633_p;
  wire g2633_n;
  wire g2634_p;
  wire g2634_n;
  wire g2635_p;
  wire g2635_n;
  wire g2636_p;
  wire g2636_n;
  wire g2637_p;
  wire g2637_n;
  wire g2638_p;
  wire g2638_n;
  wire g2639_p;
  wire g2639_n;
  wire g2640_p;
  wire g2640_n;
  wire g2641_p;
  wire g2641_n;
  wire g2642_p;
  wire g2642_n;
  wire g2643_p;
  wire g2643_n;
  wire g2644_p;
  wire g2644_n;
  wire g2645_p;
  wire g2645_n;
  wire g2646_p;
  wire g2646_n;
  wire g2647_p;
  wire g2647_n;
  wire g2648_p;
  wire g2648_n;
  wire g2649_p;
  wire g2649_n;
  wire g2650_p;
  wire g2650_n;
  wire g2651_p;
  wire g2651_n;
  wire g2652_p;
  wire g2652_n;
  wire g2653_p;
  wire g2653_n;
  wire g2654_p;
  wire g2654_n;
  wire g2655_p;
  wire g2655_n;
  wire g2656_p;
  wire g2656_n;
  wire g2657_p;
  wire g2657_n;
  wire g2658_p;
  wire g2658_n;
  wire g2659_p;
  wire g2659_n;
  wire g2660_p;
  wire g2660_n;
  wire g2661_p;
  wire g2661_n;
  wire g2662_p;
  wire g2662_n;
  wire g2663_p;
  wire g2663_n;
  wire g2664_p;
  wire g2664_n;
  wire g2665_p;
  wire g2665_n;
  wire g2666_p;
  wire g2666_n;
  wire g2667_p;
  wire g2667_n;
  wire g2668_p;
  wire g2668_n;
  wire g2669_p;
  wire g2669_n;
  wire g2670_p;
  wire g2670_n;
  wire g2671_p;
  wire g2671_n;
  wire g2672_p;
  wire g2672_n;
  wire g2673_p;
  wire g2673_n;
  wire g2674_p;
  wire g2674_n;
  wire g2675_p;
  wire g2675_n;
  wire g2676_p;
  wire g2676_n;
  wire g2677_p;
  wire g2677_n;
  wire g2678_p;
  wire g2678_n;
  wire g2679_p;
  wire g2679_n;
  wire g2680_p;
  wire g2680_n;
  wire g2681_p;
  wire g2681_n;
  wire g2682_p;
  wire g2682_n;
  wire g2683_p;
  wire g2683_n;
  wire g2684_p;
  wire g2684_n;
  wire g2685_p;
  wire g2685_n;
  wire g2686_p;
  wire g2686_n;
  wire g2687_p;
  wire g2687_n;
  wire g2688_p;
  wire g2688_n;
  wire g2689_p;
  wire g2689_n;
  wire g2690_p;
  wire g2690_n;
  wire g2691_p;
  wire g2691_n;
  wire g2692_p;
  wire g2692_n;
  wire g2693_p;
  wire g2693_n;
  wire g2694_p;
  wire g2694_n;
  wire g2695_p;
  wire g2695_n;
  wire g2696_p;
  wire g2696_n;
  wire g2697_p;
  wire g2697_n;
  wire g2698_p;
  wire g2698_n;
  wire g2699_p;
  wire g2699_n;
  wire g2700_p;
  wire g2700_n;
  wire g2701_p;
  wire g2701_n;
  wire g2702_p;
  wire g2702_n;
  wire g2703_p;
  wire g2703_n;
  wire g2704_p;
  wire g2704_n;
  wire g2705_p;
  wire g2705_n;
  wire g2706_p;
  wire g2706_n;
  wire g2707_p;
  wire g2707_n;
  wire g2708_p;
  wire g2708_n;
  wire g2709_p;
  wire g2709_n;
  wire g2710_p;
  wire g2710_n;
  wire g2711_p;
  wire g2711_n;
  wire g2712_p;
  wire g2712_n;
  wire g2713_p;
  wire g2713_n;
  wire g2714_p;
  wire g2714_n;
  wire g2715_p;
  wire g2715_n;
  wire g2716_p;
  wire g2716_n;
  wire g2717_p;
  wire g2717_n;
  wire g2718_p;
  wire g2718_n;
  wire g2719_p;
  wire g2719_n;
  wire g2720_p;
  wire g2720_n;
  wire g2721_p;
  wire g2721_n;
  wire g2722_p;
  wire g2722_n;
  wire g2723_p;
  wire g2723_n;
  wire g2724_p;
  wire g2724_n;
  wire g2725_p;
  wire g2725_n;
  wire g2726_p;
  wire g2726_n;
  wire g2727_p;
  wire g2727_n;
  wire g2728_p;
  wire g2728_n;
  wire g2729_p;
  wire g2729_n;
  wire g2730_p;
  wire g2730_n;
  wire g2731_p;
  wire g2731_n;
  wire g2732_p;
  wire g2732_n;
  wire g2733_p;
  wire g2733_n;
  wire g2734_p;
  wire g2734_n;
  wire g2735_p;
  wire g2735_n;
  wire g2736_p;
  wire g2736_n;
  wire g2737_p;
  wire g2737_n;
  wire g2738_p;
  wire g2738_n;
  wire g2739_p;
  wire g2739_n;
  wire g2740_p;
  wire g2740_n;
  wire g2741_p;
  wire g2741_n;
  wire g2742_p;
  wire g2742_n;
  wire g2743_p;
  wire g2743_n;
  wire g2744_p;
  wire g2744_n;
  wire g2745_p;
  wire g2745_n;
  wire g2746_p;
  wire g2746_n;
  wire g2747_p;
  wire g2747_n;
  wire g2748_p;
  wire g2748_n;
  wire g2749_p;
  wire g2749_n;
  wire g2750_p;
  wire g2750_n;
  wire g2751_p;
  wire g2751_n;
  wire g2752_p;
  wire g2752_n;
  wire g2753_p;
  wire g2753_n;
  wire g2754_p;
  wire g2754_n;
  wire g2755_p;
  wire g2755_n;
  wire g2756_p;
  wire g2756_n;
  wire g2757_p;
  wire g2757_n;
  wire g2758_p;
  wire g2758_n;
  wire g2759_p;
  wire g2759_n;
  wire g2760_p;
  wire g2760_n;
  wire g2761_p;
  wire g2761_n;
  wire g2762_p;
  wire g2762_n;
  wire g2763_p;
  wire g2763_n;
  wire g2764_p;
  wire g2764_n;
  wire g2765_p;
  wire g2765_n;
  wire g2766_p;
  wire g2766_n;
  wire g2767_p;
  wire g2767_n;
  wire g2768_p;
  wire g2768_n;
  wire g2769_p;
  wire g2769_n;
  wire g2770_p;
  wire g2770_n;
  wire g2771_p;
  wire g2771_n;
  wire g2772_p;
  wire g2772_n;
  wire g2773_p;
  wire g2773_n;
  wire g2774_p;
  wire g2774_n;
  wire g2775_p;
  wire g2775_n;
  wire g2776_p;
  wire g2776_n;
  wire g2777_p;
  wire g2777_n;
  wire g2778_p;
  wire g2778_n;
  wire g2779_p;
  wire g2779_n;
  wire g2780_p;
  wire g2780_n;
  wire g2781_p;
  wire g2781_n;
  wire g2782_p;
  wire g2782_n;
  wire g2783_p;
  wire g2783_n;
  wire g2784_p;
  wire g2784_n;
  wire g2785_p;
  wire g2785_n;
  wire g2786_p;
  wire g2786_n;
  wire g2787_p;
  wire g2787_n;
  wire g2788_p;
  wire g2788_n;
  wire g2789_p;
  wire g2789_n;
  wire g2790_p;
  wire g2790_n;
  wire g2791_p;
  wire g2791_n;
  wire g2792_p;
  wire g2792_n;
  wire g2793_p;
  wire g2793_n;
  wire g2794_p;
  wire g2794_n;
  wire g2795_p;
  wire g2795_n;
  wire g2796_p;
  wire g2796_n;
  wire g2797_p;
  wire g2797_n;
  wire g2798_p;
  wire g2798_n;
  wire g2799_p;
  wire g2799_n;
  wire g2800_p;
  wire g2800_n;
  wire g2801_p;
  wire g2801_n;
  wire g2802_p;
  wire g2802_n;
  wire g2803_p;
  wire g2803_n;
  wire g2804_p;
  wire g2804_n;
  wire g2805_p;
  wire g2805_n;
  wire g2806_p;
  wire g2806_n;
  wire g2807_p;
  wire g2807_n;
  wire g2808_p;
  wire g2808_n;
  wire g2809_p;
  wire g2809_n;
  wire g2810_p;
  wire g2810_n;
  wire g2811_p;
  wire g2811_n;
  wire g2812_p;
  wire g2812_n;
  wire g2813_p;
  wire g2813_n;
  wire g2814_p;
  wire g2814_n;
  wire g2815_p;
  wire g2815_n;
  wire g2816_p;
  wire g2816_n;
  wire g2817_p;
  wire g2817_n;
  wire g2818_p;
  wire g2818_n;
  wire g2819_p;
  wire g2819_n;
  wire g2820_p;
  wire g2820_n;
  wire g2821_p;
  wire g2821_n;
  wire g2822_p;
  wire g2822_n;
  wire g2823_p;
  wire g2823_n;
  wire g2824_p;
  wire g2824_n;
  wire g2825_p;
  wire g2825_n;
  wire g2826_p;
  wire g2826_n;
  wire g2827_p;
  wire g2827_n;
  wire g2828_p;
  wire g2828_n;
  wire g2829_p;
  wire g2829_n;
  wire g2830_p;
  wire g2830_n;
  wire g2831_p;
  wire g2831_n;
  wire g2832_p;
  wire g2832_n;
  wire g2833_p;
  wire g2833_n;
  wire g2834_p;
  wire g2834_n;
  wire g2835_p;
  wire g2835_n;
  wire g2836_p;
  wire g2836_n;
  wire g2837_p;
  wire g2837_n;
  wire g2838_p;
  wire g2838_n;
  wire g2839_p;
  wire g2839_n;
  wire g2840_p;
  wire g2840_n;
  wire g2841_p;
  wire g2841_n;
  wire g2842_p;
  wire g2842_n;
  wire g2843_p;
  wire g2843_n;
  wire g2844_p;
  wire g2844_n;
  wire g2845_p;
  wire g2845_n;
  wire g2846_p;
  wire g2846_n;
  wire g2847_p;
  wire g2847_n;
  wire g2848_p;
  wire g2848_n;
  wire g2849_p;
  wire g2849_n;
  wire g2850_p;
  wire g2850_n;
  wire g2851_p;
  wire g2851_n;
  wire g2852_p;
  wire g2852_n;
  wire g2853_p;
  wire g2853_n;
  wire g2854_p;
  wire g2854_n;
  wire g2855_p;
  wire g2855_n;
  wire g2856_p;
  wire g2856_n;
  wire g2857_p;
  wire g2857_n;
  wire g2858_p;
  wire g2858_n;
  wire g2859_p;
  wire g2859_n;
  wire g2860_p;
  wire g2860_n;
  wire g2861_p;
  wire g2861_n;
  wire g2862_p;
  wire g2862_n;
  wire g2863_p;
  wire g2863_n;
  wire g2864_p;
  wire g2864_n;
  wire g2865_p;
  wire g2865_n;
  wire g2866_p;
  wire g2866_n;
  wire g2867_p;
  wire g2867_n;
  wire g2868_p;
  wire g2868_n;
  wire g2869_p;
  wire g2869_n;
  wire g2870_p;
  wire g2870_n;
  wire g2871_p;
  wire g2871_n;
  wire g2872_p;
  wire g2872_n;
  wire g2873_p;
  wire g2873_n;
  wire g2874_p;
  wire g2874_n;
  wire g2875_p;
  wire g2875_n;
  wire g2876_p;
  wire g2876_n;
  wire g2877_p;
  wire g2877_n;
  wire g2878_p;
  wire g2878_n;
  wire g2879_p;
  wire g2879_n;
  wire g2880_p;
  wire g2880_n;
  wire g2881_p;
  wire g2881_n;
  wire g2882_p;
  wire g2882_n;
  wire g2883_p;
  wire g2883_n;
  wire g2884_p;
  wire g2884_n;
  wire g2885_p;
  wire g2885_n;
  wire g2886_p;
  wire g2886_n;
  wire g2887_p;
  wire g2887_n;
  wire g2888_p;
  wire g2888_n;
  wire g2889_p;
  wire g2889_n;
  wire g2890_p;
  wire g2890_n;
  wire g2891_p;
  wire g2891_n;
  wire g2892_p;
  wire g2892_n;
  wire g2893_p;
  wire g2893_n;
  wire g2894_p;
  wire g2894_n;
  wire g2895_p;
  wire g2895_n;
  wire g2896_p;
  wire g2896_n;
  wire g2897_p;
  wire g2897_n;
  wire g2898_p;
  wire g2898_n;
  wire g2899_p;
  wire g2899_n;
  wire g2900_p;
  wire g2900_n;
  wire g2901_p;
  wire g2901_n;
  wire g2902_p;
  wire g2902_n;
  wire g2903_p;
  wire g2903_n;
  wire g2904_p;
  wire g2904_n;
  wire g2905_p;
  wire g2905_n;
  wire g2906_p;
  wire g2906_n;
  wire g2907_p;
  wire g2907_n;
  wire g2908_p;
  wire g2908_n;
  wire g2909_p;
  wire g2909_n;
  wire g2910_p;
  wire g2910_n;
  wire g2911_p;
  wire g2911_n;
  wire g2912_p;
  wire g2912_n;
  wire g2913_p;
  wire g2913_n;
  wire g2914_p;
  wire g2914_n;
  wire g2915_p;
  wire g2915_n;
  wire g2916_p;
  wire g2916_n;
  wire g2917_p;
  wire g2917_n;
  wire g2918_p;
  wire g2918_n;
  wire g2919_p;
  wire g2919_n;
  wire g2920_p;
  wire g2920_n;
  wire g2921_p;
  wire g2921_n;
  wire g2922_p;
  wire g2922_n;
  wire g2923_p;
  wire g2923_n;
  wire g2924_p;
  wire g2924_n;
  wire g2925_p;
  wire g2925_n;
  wire g2926_p;
  wire g2926_n;
  wire g2927_p;
  wire g2927_n;
  wire g2928_p;
  wire g2928_n;
  wire g2929_p;
  wire g2929_n;
  wire g2930_p;
  wire g2930_n;
  wire g2931_p;
  wire g2931_n;
  wire g2932_p;
  wire g2932_n;
  wire g2933_p;
  wire g2933_n;
  wire g2934_p;
  wire g2934_n;
  wire g2935_p;
  wire g2935_n;
  wire g2936_p;
  wire g2936_n;
  wire g2937_p;
  wire g2937_n;
  wire g2938_p;
  wire g2938_n;
  wire g2939_p;
  wire g2939_n;
  wire g2940_p;
  wire g2940_n;
  wire g2941_p;
  wire g2941_n;
  wire g2942_p;
  wire g2942_n;
  wire g2943_p;
  wire g2943_n;
  wire g2944_p;
  wire g2944_n;
  wire g2945_p;
  wire g2945_n;
  wire g2946_p;
  wire g2946_n;
  wire g2947_p;
  wire g2947_n;
  wire g2948_p;
  wire g2948_n;
  wire g2949_p;
  wire g2949_n;
  wire g2950_p;
  wire g2950_n;
  wire g2951_p;
  wire g2951_n;
  wire g2952_p;
  wire g2952_n;
  wire g2953_p;
  wire g2953_n;
  wire g2954_p;
  wire g2954_n;
  wire g2955_p;
  wire g2955_n;
  wire g2956_p;
  wire g2956_n;
  wire g2957_p;
  wire g2957_n;
  wire g2958_p;
  wire g2958_n;
  wire g2959_p;
  wire g2959_n;
  wire g2960_p;
  wire g2960_n;
  wire g2961_p;
  wire g2961_n;
  wire g2962_p;
  wire g2962_n;
  wire g2963_p;
  wire g2963_n;
  wire g2964_p;
  wire g2964_n;
  wire g2965_p;
  wire g2965_n;
  wire g2966_p;
  wire g2966_n;
  wire g2967_p;
  wire g2967_n;
  wire g2968_p;
  wire g2968_n;
  wire g2969_p;
  wire g2969_n;
  wire g2970_p;
  wire g2970_n;
  wire g2971_p;
  wire g2971_n;
  wire g2972_p;
  wire g2972_n;
  wire g2973_p;
  wire g2973_n;
  wire g2974_p;
  wire g2974_n;
  wire g2975_p;
  wire g2975_n;
  wire g2976_p;
  wire g2976_n;
  wire g2977_p;
  wire g2977_n;
  wire g2978_p;
  wire g2978_n;
  wire g2979_p;
  wire g2979_n;
  wire g2980_p;
  wire g2980_n;
  wire g2981_p;
  wire g2981_n;
  wire g2982_p;
  wire g2982_n;
  wire g2983_p;
  wire g2983_n;
  wire g2984_p;
  wire g2984_n;
  wire g2985_p;
  wire g2985_n;
  wire g2986_p;
  wire g2986_n;
  wire g2987_p;
  wire g2987_n;
  wire g2988_p;
  wire g2988_n;
  wire g2989_p;
  wire g2989_n;
  wire g2990_p;
  wire g2990_n;
  wire g2991_p;
  wire g2991_n;
  wire g2992_p;
  wire g2992_n;
  wire g2993_p;
  wire g2993_n;
  wire g2994_p;
  wire g2994_n;
  wire g2995_p;
  wire g2995_n;
  wire g2996_p;
  wire g2996_n;
  wire g2997_p;
  wire g2997_n;
  wire g2998_p;
  wire g2998_n;
  wire g2999_p;
  wire g2999_n;
  wire g3000_p;
  wire g3000_n;
  wire g3001_p;
  wire g3001_n;
  wire g3002_p;
  wire g3002_n;
  wire g3003_p;
  wire g3003_n;
  wire g3004_p;
  wire g3004_n;
  wire g3005_p;
  wire g3005_n;
  wire g3006_p;
  wire g3006_n;
  wire g3007_p;
  wire g3007_n;
  wire g3008_p;
  wire g3008_n;
  wire g3009_p;
  wire g3009_n;
  wire g3010_p;
  wire g3010_n;
  wire g3011_p;
  wire g3011_n;
  wire g3012_p;
  wire g3012_n;
  wire g3013_p;
  wire g3013_n;
  wire g3014_p;
  wire g3014_n;
  wire g3015_p;
  wire g3015_n;
  wire g3016_p;
  wire g3016_n;
  wire g3017_p;
  wire g3017_n;
  wire g3018_p;
  wire g3018_n;
  wire g3019_p;
  wire g3019_n;
  wire g3020_p;
  wire g3020_n;
  wire g3021_p;
  wire g3021_n;
  wire g3022_p;
  wire g3022_n;
  wire g3023_p;
  wire g3023_n;
  wire g3024_p;
  wire g3024_n;
  wire g3025_p;
  wire g3025_n;
  wire g3026_p;
  wire g3026_n;
  wire g3027_p;
  wire g3027_n;
  wire g3028_p;
  wire g3028_n;
  wire g3029_p;
  wire g3029_n;
  wire g3030_p;
  wire g3030_n;
  wire g3031_p;
  wire g3031_n;
  wire g3032_p;
  wire g3032_n;
  wire g3033_p;
  wire g3033_n;
  wire g3034_p;
  wire g3034_n;
  wire g3035_p;
  wire g3035_n;
  wire g3036_p;
  wire g3036_n;
  wire g3037_p;
  wire g3037_n;
  wire g3038_p;
  wire g3038_n;
  wire g3039_p;
  wire g3039_n;
  wire g3040_p;
  wire g3040_n;
  wire g3041_p;
  wire g3041_n;
  wire g3042_p;
  wire g3042_n;
  wire g3043_p;
  wire g3043_n;
  wire g3044_p;
  wire g3044_n;
  wire g3045_p;
  wire g3045_n;
  wire g3046_p;
  wire g3046_n;
  wire g3047_p;
  wire g3047_n;
  wire g3048_p;
  wire g3048_n;
  wire g3049_p;
  wire g3049_n;
  wire g3050_p;
  wire g3050_n;
  wire g3051_p;
  wire g3051_n;
  wire g3052_p;
  wire g3052_n;
  wire g3053_p;
  wire g3053_n;
  wire g3054_p;
  wire g3054_n;
  wire g3055_p;
  wire g3055_n;
  wire g3056_p;
  wire g3056_n;
  wire g3057_p;
  wire g3057_n;
  wire g3058_p;
  wire g3058_n;
  wire g3059_p;
  wire g3059_n;
  wire g3060_p;
  wire g3060_n;
  wire g3061_p;
  wire g3061_n;
  wire g3062_p;
  wire g3062_n;
  wire g3063_p;
  wire g3063_n;
  wire g3064_p;
  wire g3064_n;
  wire g3065_p;
  wire g3065_n;
  wire g3066_p;
  wire g3066_n;
  wire g3067_p;
  wire g3067_n;
  wire g3068_p;
  wire g3068_n;
  wire g3069_p;
  wire g3069_n;
  wire g3070_p;
  wire g3070_n;
  wire g3071_p;
  wire g3071_n;
  wire g3072_p;
  wire g3072_n;
  wire g3073_p;
  wire g3073_n;
  wire g3074_p;
  wire g3074_n;
  wire g3075_p;
  wire g3075_n;
  wire g3076_p;
  wire g3076_n;
  wire g3077_p;
  wire g3077_n;
  wire g3078_p;
  wire g3078_n;
  wire g3079_p;
  wire g3079_n;
  wire g3080_p;
  wire g3080_n;
  wire g3081_p;
  wire g3081_n;
  wire g3082_p;
  wire g3082_n;
  wire g3083_p;
  wire g3083_n;
  wire g3084_p;
  wire g3084_n;
  wire g3085_p;
  wire g3085_n;
  wire g3086_p;
  wire g3086_n;
  wire g3087_p;
  wire g3087_n;
  wire g3088_p;
  wire g3088_n;
  wire g3089_p;
  wire g3089_n;
  wire g3090_p;
  wire g3090_n;
  wire g3091_p;
  wire g3091_n;
  wire g3092_p;
  wire g3092_n;
  wire g3093_p;
  wire g3093_n;
  wire g3094_p;
  wire g3094_n;
  wire g3095_p;
  wire g3095_n;
  wire g3096_p;
  wire g3096_n;
  wire g3097_p;
  wire g3097_n;
  wire g3098_p;
  wire g3098_n;
  wire g3099_p;
  wire g3099_n;
  wire g3100_p;
  wire g3100_n;
  wire g3101_p;
  wire g3101_n;
  wire g3102_p;
  wire g3102_n;
  wire g3103_p;
  wire g3103_n;
  wire g3104_p;
  wire g3104_n;
  wire g3105_p;
  wire g3105_n;
  wire g3106_p;
  wire g3106_n;
  wire g3107_p;
  wire g3107_n;
  wire g3108_p;
  wire g3108_n;
  wire g3109_p;
  wire g3109_n;
  wire g3110_p;
  wire g3110_n;
  wire g3111_p;
  wire g3111_n;
  wire g3112_p;
  wire g3112_n;
  wire g3113_p;
  wire g3113_n;
  wire g3114_p;
  wire g3114_n;
  wire g3115_p;
  wire g3115_n;
  wire g3116_p;
  wire g3116_n;
  wire g3117_p;
  wire g3117_n;
  wire g3118_p;
  wire g3118_n;
  wire g3119_p;
  wire g3119_n;
  wire g3120_p;
  wire g3120_n;
  wire g3121_p;
  wire g3121_n;
  wire g3122_p;
  wire g3122_n;
  wire g3123_p;
  wire g3123_n;
  wire g3124_p;
  wire g3124_n;
  wire g3125_p;
  wire g3125_n;
  wire g3126_p;
  wire g3126_n;
  wire g3127_p;
  wire g3127_n;
  wire g3128_p;
  wire g3128_n;
  wire g3129_p;
  wire g3129_n;
  wire g3130_p;
  wire g3130_n;
  wire g3131_p;
  wire g3131_n;
  wire g3132_p;
  wire g3132_n;
  wire g3133_p;
  wire g3133_n;
  wire g3134_p;
  wire g3134_n;
  wire g3135_p;
  wire g3135_n;
  wire g3136_p;
  wire g3136_n;
  wire g3137_p;
  wire g3137_n;
  wire g3138_p;
  wire g3138_n;
  wire g3139_p;
  wire g3139_n;
  wire g3140_p;
  wire g3140_n;
  wire g3141_p;
  wire g3141_n;
  wire g3142_p;
  wire g3142_n;
  wire g3143_p;
  wire g3143_n;
  wire g3144_p;
  wire g3144_n;
  wire g3145_p;
  wire g3145_n;
  wire g3146_p;
  wire g3146_n;
  wire g3147_p;
  wire g3147_n;
  wire g3148_p;
  wire g3148_n;
  wire g3149_p;
  wire g3149_n;
  wire g3150_p;
  wire g3150_n;
  wire g3151_p;
  wire g3151_n;
  wire g3152_p;
  wire g3152_n;
  wire g3153_p;
  wire g3153_n;
  wire g3154_p;
  wire g3154_n;
  wire g3155_p;
  wire g3155_n;
  wire g3156_p;
  wire g3156_n;
  wire g3157_p;
  wire g3157_n;
  wire g3158_p;
  wire g3158_n;
  wire g3159_p;
  wire g3159_n;
  wire g3160_p;
  wire g3160_n;
  wire g3161_p;
  wire g3161_n;
  wire g3162_p;
  wire g3162_n;
  wire g3163_p;
  wire g3163_n;
  wire g3164_p;
  wire g3164_n;
  wire g3165_p;
  wire g3165_n;
  wire g3166_p;
  wire g3166_n;
  wire g3167_p;
  wire g3167_n;
  wire g3168_p;
  wire g3168_n;
  wire g3169_p;
  wire g3169_n;
  wire g3170_p;
  wire g3170_n;
  wire g3171_p;
  wire g3171_n;
  wire g3172_p;
  wire g3172_n;
  wire g3173_p;
  wire g3173_n;
  wire g3174_p;
  wire g3174_n;
  wire g3175_p;
  wire g3175_n;
  wire g3176_p;
  wire g3176_n;
  wire g3177_p;
  wire g3177_n;
  wire g3178_p;
  wire g3178_n;
  wire n3399_lo_p_spl_;
  wire n2619_lo_p_spl_;
  wire n4587_lo_n_spl_;
  wire n2739_lo_n_spl_;
  wire n4455_lo_n_spl_;
  wire n4239_lo_n_spl_;
  wire g1198_n_spl_;
  wire g1198_n_spl_0;
  wire g1198_n_spl_00;
  wire g1198_n_spl_000;
  wire g1198_n_spl_001;
  wire g1198_n_spl_01;
  wire g1198_n_spl_010;
  wire g1198_n_spl_011;
  wire g1198_n_spl_1;
  wire g1198_n_spl_10;
  wire g1198_n_spl_100;
  wire g1198_n_spl_11;
  wire n4563_lo_n_spl_;
  wire n4563_lo_n_spl_0;
  wire n4563_lo_n_spl_00;
  wire n4563_lo_n_spl_01;
  wire n4563_lo_n_spl_1;
  wire n4563_lo_n_spl_10;
  wire n4563_lo_n_spl_11;
  wire n4563_lo_p_spl_;
  wire n4563_lo_p_spl_0;
  wire n4563_lo_p_spl_00;
  wire n4563_lo_p_spl_01;
  wire n4563_lo_p_spl_1;
  wire n4563_lo_p_spl_10;
  wire n4563_lo_p_spl_11;
  wire n2991_lo_n_spl_;
  wire g1198_p_spl_;
  wire g1216_n_spl_;
  wire g1216_n_spl_0;
  wire g1216_n_spl_1;
  wire g1217_n_spl_;
  wire g1217_n_spl_0;
  wire g1217_n_spl_1;
  wire n3399_lo_n_spl_;
  wire n3399_lo_n_spl_0;
  wire n3399_lo_n_spl_00;
  wire n3399_lo_n_spl_1;
  wire n7357_o2_p_spl_;
  wire n7357_o2_p_spl_0;
  wire n4359_lo_n_spl_;
  wire n4035_lo_p_spl_;
  wire n7359_o2_p_spl_;
  wire n7359_o2_p_spl_0;
  wire n4035_lo_n_spl_;
  wire n7449_o2_n_spl_;
  wire n7449_o2_n_spl_0;
  wire n7452_o2_n_spl_;
  wire n7452_o2_n_spl_0;
  wire n4347_lo_n_spl_;
  wire n4011_lo_p_spl_;
  wire n4011_lo_n_spl_;
  wire n3963_lo_n_spl_;
  wire n3963_lo_n_spl_0;
  wire n3963_lo_p_spl_;
  wire g1265_p_spl_;
  wire g1255_p_spl_;
  wire g1268_p_spl_;
  wire n4635_lo_p_spl_;
  wire n4635_lo_p_spl_0;
  wire n4635_lo_p_spl_00;
  wire n4635_lo_p_spl_000;
  wire n4635_lo_p_spl_001;
  wire n4635_lo_p_spl_01;
  wire n4635_lo_p_spl_010;
  wire n4635_lo_p_spl_011;
  wire n4635_lo_p_spl_1;
  wire n4635_lo_p_spl_10;
  wire n4635_lo_p_spl_11;
  wire n4407_lo_n_spl_;
  wire n4143_lo_p_spl_;
  wire n4623_lo_p_spl_;
  wire n4623_lo_p_spl_0;
  wire n4623_lo_p_spl_00;
  wire n4623_lo_p_spl_000;
  wire n4623_lo_p_spl_001;
  wire n4623_lo_p_spl_01;
  wire n4623_lo_p_spl_010;
  wire n4623_lo_p_spl_1;
  wire n4623_lo_p_spl_10;
  wire n4623_lo_p_spl_11;
  wire n4143_lo_n_spl_;
  wire n4599_lo_n_spl_;
  wire n4599_lo_n_spl_0;
  wire n4599_lo_n_spl_00;
  wire n4599_lo_n_spl_000;
  wire n4599_lo_n_spl_001;
  wire n4599_lo_n_spl_01;
  wire n4599_lo_n_spl_010;
  wire n4599_lo_n_spl_011;
  wire n4599_lo_n_spl_1;
  wire n4599_lo_n_spl_10;
  wire n4599_lo_n_spl_11;
  wire n4611_lo_n_spl_;
  wire n4611_lo_n_spl_0;
  wire n4611_lo_n_spl_00;
  wire n4611_lo_n_spl_000;
  wire n4611_lo_n_spl_001;
  wire n4611_lo_n_spl_01;
  wire n4611_lo_n_spl_010;
  wire n4611_lo_n_spl_1;
  wire n4611_lo_n_spl_10;
  wire n4611_lo_n_spl_11;
  wire n4395_lo_n_spl_;
  wire n4119_lo_p_spl_;
  wire n4119_lo_n_spl_;
  wire n4371_lo_n_spl_;
  wire n4371_lo_n_spl_0;
  wire n4059_lo_p_spl_;
  wire n4059_lo_n_spl_;
  wire n4371_lo_p_spl_;
  wire g1294_p_spl_;
  wire g1284_p_spl_;
  wire g1297_p_spl_;
  wire g1307_p_spl_;
  wire n4299_lo_n_spl_;
  wire n4299_lo_n_spl_0;
  wire n3759_lo_p_spl_;
  wire n3759_lo_n_spl_;
  wire n4299_lo_p_spl_;
  wire n4287_lo_n_spl_;
  wire n3735_lo_p_spl_;
  wire n3735_lo_n_spl_;
  wire n4335_lo_n_spl_;
  wire n3711_lo_p_spl_;
  wire n3711_lo_n_spl_;
  wire n4323_lo_n_spl_;
  wire n3687_lo_p_spl_;
  wire n3687_lo_n_spl_;
  wire g1332_p_spl_;
  wire g1322_p_spl_;
  wire g1342_p_spl_;
  wire g1352_p_spl_;
  wire n4227_lo_n_spl_;
  wire n3915_lo_p_spl_;
  wire n3915_lo_n_spl_;
  wire n4275_lo_n_spl_;
  wire n3891_lo_p_spl_;
  wire n3891_lo_n_spl_;
  wire n4263_lo_n_spl_;
  wire n3867_lo_p_spl_;
  wire n3867_lo_n_spl_;
  wire n4251_lo_n_spl_;
  wire n3843_lo_p_spl_;
  wire n3843_lo_n_spl_;
  wire g1375_p_spl_;
  wire g1365_p_spl_;
  wire g1385_p_spl_;
  wire g1395_p_spl_;
  wire n6419_o2_n_spl_;
  wire n6613_o2_n_spl_;
  wire n6613_o2_n_spl_0;
  wire G3467_o2_n_spl_;
  wire G3467_o2_n_spl_0;
  wire G3467_o2_n_spl_1;
  wire g1403_n_spl_;
  wire G3570_o2_n_spl_;
  wire G2759_o2_p_spl_;
  wire G2759_o2_p_spl_0;
  wire G2759_o2_p_spl_1;
  wire G3559_o2_n_spl_;
  wire G3559_o2_n_spl_0;
  wire G2752_o2_p_spl_;
  wire G2752_o2_p_spl_0;
  wire G2752_o2_p_spl_00;
  wire G2752_o2_p_spl_01;
  wire G2752_o2_p_spl_1;
  wire G3303_o2_p_spl_;
  wire G3303_o2_p_spl_0;
  wire G3303_o2_p_spl_00;
  wire G3303_o2_p_spl_000;
  wire G3303_o2_p_spl_01;
  wire G3303_o2_p_spl_1;
  wire G3303_o2_p_spl_10;
  wire G3303_o2_p_spl_11;
  wire G2797_o2_n_spl_;
  wire G2797_o2_n_spl_0;
  wire G3303_o2_n_spl_;
  wire G3303_o2_n_spl_0;
  wire G3303_o2_n_spl_00;
  wire G3303_o2_n_spl_000;
  wire G3303_o2_n_spl_01;
  wire G3303_o2_n_spl_1;
  wire G3303_o2_n_spl_10;
  wire G3303_o2_n_spl_11;
  wire G2797_o2_p_spl_;
  wire G2797_o2_p_spl_0;
  wire G3583_o2_p_spl_;
  wire G3583_o2_p_spl_0;
  wire G3583_o2_p_spl_00;
  wire G3583_o2_p_spl_01;
  wire G3583_o2_p_spl_1;
  wire G3583_o2_n_spl_;
  wire G3583_o2_n_spl_0;
  wire G3583_o2_n_spl_00;
  wire G3583_o2_n_spl_01;
  wire G3583_o2_n_spl_1;
  wire G3576_o2_p_spl_;
  wire G3576_o2_p_spl_0;
  wire G3576_o2_p_spl_00;
  wire G3576_o2_p_spl_01;
  wire G3576_o2_p_spl_1;
  wire G3576_o2_n_spl_;
  wire G3576_o2_n_spl_0;
  wire G3576_o2_n_spl_00;
  wire G3576_o2_n_spl_01;
  wire G3576_o2_n_spl_1;
  wire G3594_o2_p_spl_;
  wire G3594_o2_p_spl_0;
  wire G3594_o2_p_spl_00;
  wire G3594_o2_p_spl_01;
  wire G3594_o2_p_spl_1;
  wire G3594_o2_n_spl_;
  wire G3594_o2_n_spl_0;
  wire G3594_o2_n_spl_00;
  wire G3594_o2_n_spl_01;
  wire G3594_o2_n_spl_1;
  wire g1411_n_spl_;
  wire g1407_n_spl_;
  wire n6420_o2_n_spl_;
  wire n6614_o2_p_spl_;
  wire n6614_o2_p_spl_0;
  wire G2810_o2_p_spl_;
  wire G2810_o2_p_spl_0;
  wire G2810_o2_p_spl_1;
  wire g1415_n_spl_;
  wire G3415_o2_n_spl_;
  wire G3393_o2_n_spl_;
  wire G3393_o2_n_spl_0;
  wire G3393_o2_n_spl_1;
  wire G3404_o2_n_spl_;
  wire G3404_o2_n_spl_0;
  wire G3386_o2_n_spl_;
  wire G3386_o2_n_spl_0;
  wire G3386_o2_n_spl_00;
  wire G3386_o2_n_spl_1;
  wire G3428_o2_p_spl_;
  wire G3428_o2_p_spl_0;
  wire G3428_o2_p_spl_00;
  wire G3428_o2_p_spl_000;
  wire G3428_o2_p_spl_01;
  wire G3428_o2_p_spl_1;
  wire G3428_o2_p_spl_10;
  wire G3428_o2_p_spl_11;
  wire G3459_o2_p_spl_;
  wire G3459_o2_p_spl_0;
  wire G3428_o2_n_spl_;
  wire G3428_o2_n_spl_0;
  wire G3428_o2_n_spl_00;
  wire G3428_o2_n_spl_000;
  wire G3428_o2_n_spl_01;
  wire G3428_o2_n_spl_1;
  wire G3428_o2_n_spl_10;
  wire G3428_o2_n_spl_11;
  wire G3459_o2_n_spl_;
  wire G3459_o2_n_spl_0;
  wire G3438_o2_p_spl_;
  wire G3438_o2_p_spl_0;
  wire G3438_o2_p_spl_00;
  wire G3438_o2_p_spl_01;
  wire G3438_o2_p_spl_1;
  wire G3438_o2_n_spl_;
  wire G3438_o2_n_spl_0;
  wire G3438_o2_n_spl_00;
  wire G3438_o2_n_spl_01;
  wire G3438_o2_n_spl_1;
  wire G3421_o2_p_spl_;
  wire G3421_o2_p_spl_0;
  wire G3421_o2_p_spl_00;
  wire G3421_o2_p_spl_01;
  wire G3421_o2_p_spl_1;
  wire G3421_o2_n_spl_;
  wire G3421_o2_n_spl_0;
  wire G3421_o2_n_spl_00;
  wire G3421_o2_n_spl_01;
  wire G3421_o2_n_spl_1;
  wire G3449_o2_p_spl_;
  wire G3449_o2_p_spl_0;
  wire G3449_o2_p_spl_00;
  wire G3449_o2_p_spl_01;
  wire G3449_o2_p_spl_1;
  wire G3449_o2_n_spl_;
  wire G3449_o2_n_spl_0;
  wire G3449_o2_n_spl_00;
  wire G3449_o2_n_spl_01;
  wire G3449_o2_n_spl_1;
  wire g1423_n_spl_;
  wire g1419_n_spl_;
  wire g1430_p_spl_;
  wire g1427_n_spl_;
  wire g1430_n_spl_;
  wire g1427_p_spl_;
  wire g1435_p_spl_;
  wire g1435_p_spl_0;
  wire g1435_p_spl_1;
  wire g1434_n_spl_;
  wire g1434_n_spl_0;
  wire g1434_n_spl_1;
  wire g1435_n_spl_;
  wire g1435_n_spl_0;
  wire g1435_n_spl_1;
  wire g1434_p_spl_;
  wire g1434_p_spl_0;
  wire g1434_p_spl_1;
  wire G1147_o2_n_spl_;
  wire G1147_o2_n_spl_0;
  wire G1147_o2_n_spl_1;
  wire G1147_o2_p_spl_;
  wire G1147_o2_p_spl_0;
  wire G1147_o2_p_spl_1;
  wire g1455_p_spl_;
  wire g1452_n_spl_;
  wire g1455_n_spl_;
  wire g1452_p_spl_;
  wire g1460_p_spl_;
  wire g1460_p_spl_0;
  wire g1460_p_spl_1;
  wire g1459_n_spl_;
  wire g1459_n_spl_0;
  wire g1459_n_spl_1;
  wire g1460_n_spl_;
  wire g1460_n_spl_0;
  wire g1460_n_spl_1;
  wire g1459_p_spl_;
  wire g1459_p_spl_0;
  wire g1459_p_spl_1;
  wire G2336_o2_p_spl_;
  wire G2336_o2_p_spl_0;
  wire G2336_o2_p_spl_1;
  wire G2336_o2_n_spl_;
  wire G2336_o2_n_spl_0;
  wire G2336_o2_n_spl_1;
  wire n4311_lo_n_spl_;
  wire n4311_lo_n_spl_0;
  wire g1475_n_spl_;
  wire G2770_o2_p_spl_;
  wire G2774_o2_n_spl_;
  wire G2780_o2_n_spl_;
  wire n7463_o2_n_spl_;
  wire n7463_o2_n_spl_0;
  wire n7463_o2_n_spl_1;
  wire G2540_o2_p_spl_;
  wire G2540_o2_n_spl_;
  wire G2788_o2_p_spl_;
  wire G2788_o2_p_spl_0;
  wire G2788_o2_n_spl_;
  wire G2788_o2_n_spl_0;
  wire G2792_o2_p_spl_;
  wire G2792_o2_p_spl_0;
  wire G2792_o2_n_spl_;
  wire G2792_o2_n_spl_0;
  wire g1503_p_spl_;
  wire g1503_n_spl_;
  wire G2804_o2_n_spl_;
  wire G2804_o2_n_spl_0;
  wire G2804_o2_n_spl_1;
  wire G2804_o2_p_spl_;
  wire G2804_o2_p_spl_0;
  wire G2804_o2_p_spl_1;
  wire g1510_p_spl_;
  wire G2675_o2_n_spl_;
  wire G2679_o2_n_spl_;
  wire G2685_o2_n_spl_;
  wire G2693_o2_p_spl_;
  wire G2693_o2_n_spl_;
  wire G2696_o2_p_spl_;
  wire G2696_o2_p_spl_0;
  wire G2696_o2_n_spl_;
  wire G2696_o2_n_spl_0;
  wire G2700_o2_p_spl_;
  wire G2700_o2_p_spl_0;
  wire G2700_o2_n_spl_;
  wire G2700_o2_n_spl_0;
  wire g1529_p_spl_;
  wire g1529_n_spl_;
  wire G2705_o2_p_spl_;
  wire G2705_o2_p_spl_0;
  wire G2705_o2_p_spl_1;
  wire G2705_o2_n_spl_;
  wire G2705_o2_n_spl_0;
  wire G2705_o2_n_spl_1;
  wire g1536_p_spl_;
  wire n7358_o2_p_spl_;
  wire n7360_o2_p_spl_;
  wire n4719_lo_p_spl_;
  wire n4719_lo_p_spl_0;
  wire n4719_lo_p_spl_00;
  wire n4719_lo_p_spl_000;
  wire n4719_lo_p_spl_0000;
  wire n4719_lo_p_spl_00000;
  wire n4719_lo_p_spl_00001;
  wire n4719_lo_p_spl_0001;
  wire n4719_lo_p_spl_00010;
  wire n4719_lo_p_spl_00011;
  wire n4719_lo_p_spl_001;
  wire n4719_lo_p_spl_0010;
  wire n4719_lo_p_spl_00100;
  wire n4719_lo_p_spl_00101;
  wire n4719_lo_p_spl_0011;
  wire n4719_lo_p_spl_00110;
  wire n4719_lo_p_spl_00111;
  wire n4719_lo_p_spl_01;
  wire n4719_lo_p_spl_010;
  wire n4719_lo_p_spl_0100;
  wire n4719_lo_p_spl_01000;
  wire n4719_lo_p_spl_0101;
  wire n4719_lo_p_spl_011;
  wire n4719_lo_p_spl_0110;
  wire n4719_lo_p_spl_0111;
  wire n4719_lo_p_spl_1;
  wire n4719_lo_p_spl_10;
  wire n4719_lo_p_spl_100;
  wire n4719_lo_p_spl_1000;
  wire n4719_lo_p_spl_1001;
  wire n4719_lo_p_spl_101;
  wire n4719_lo_p_spl_1010;
  wire n4719_lo_p_spl_1011;
  wire n4719_lo_p_spl_11;
  wire n4719_lo_p_spl_110;
  wire n4719_lo_p_spl_1100;
  wire n4719_lo_p_spl_1101;
  wire n4719_lo_p_spl_111;
  wire n4719_lo_p_spl_1110;
  wire n4719_lo_p_spl_1111;
  wire n4731_lo_p_spl_;
  wire n4731_lo_p_spl_0;
  wire n4731_lo_p_spl_00;
  wire n4731_lo_p_spl_000;
  wire n4731_lo_p_spl_0000;
  wire n4731_lo_p_spl_00000;
  wire n4731_lo_p_spl_00001;
  wire n4731_lo_p_spl_0001;
  wire n4731_lo_p_spl_00010;
  wire n4731_lo_p_spl_00011;
  wire n4731_lo_p_spl_001;
  wire n4731_lo_p_spl_0010;
  wire n4731_lo_p_spl_00100;
  wire n4731_lo_p_spl_00101;
  wire n4731_lo_p_spl_0011;
  wire n4731_lo_p_spl_00110;
  wire n4731_lo_p_spl_00111;
  wire n4731_lo_p_spl_01;
  wire n4731_lo_p_spl_010;
  wire n4731_lo_p_spl_0100;
  wire n4731_lo_p_spl_01000;
  wire n4731_lo_p_spl_0101;
  wire n4731_lo_p_spl_011;
  wire n4731_lo_p_spl_0110;
  wire n4731_lo_p_spl_0111;
  wire n4731_lo_p_spl_1;
  wire n4731_lo_p_spl_10;
  wire n4731_lo_p_spl_100;
  wire n4731_lo_p_spl_1000;
  wire n4731_lo_p_spl_1001;
  wire n4731_lo_p_spl_101;
  wire n4731_lo_p_spl_1010;
  wire n4731_lo_p_spl_1011;
  wire n4731_lo_p_spl_11;
  wire n4731_lo_p_spl_110;
  wire n4731_lo_p_spl_1100;
  wire n4731_lo_p_spl_1101;
  wire n4731_lo_p_spl_111;
  wire n4731_lo_p_spl_1110;
  wire n4731_lo_p_spl_1111;
  wire n2859_lo_p_spl_;
  wire n2859_lo_p_spl_0;
  wire n2859_lo_n_spl_;
  wire n2859_lo_n_spl_0;
  wire g1557_n_spl_;
  wire n4719_lo_n_spl_;
  wire n4719_lo_n_spl_0;
  wire n4719_lo_n_spl_00;
  wire n4719_lo_n_spl_000;
  wire n4719_lo_n_spl_0000;
  wire n4719_lo_n_spl_0001;
  wire n4719_lo_n_spl_001;
  wire n4719_lo_n_spl_0010;
  wire n4719_lo_n_spl_0011;
  wire n4719_lo_n_spl_01;
  wire n4719_lo_n_spl_010;
  wire n4719_lo_n_spl_0100;
  wire n4719_lo_n_spl_0101;
  wire n4719_lo_n_spl_011;
  wire n4719_lo_n_spl_0110;
  wire n4719_lo_n_spl_0111;
  wire n4719_lo_n_spl_1;
  wire n4719_lo_n_spl_10;
  wire n4719_lo_n_spl_100;
  wire n4719_lo_n_spl_101;
  wire n4719_lo_n_spl_11;
  wire n4719_lo_n_spl_110;
  wire n4719_lo_n_spl_111;
  wire n4731_lo_n_spl_;
  wire n4731_lo_n_spl_0;
  wire n4731_lo_n_spl_00;
  wire n4731_lo_n_spl_000;
  wire n4731_lo_n_spl_0000;
  wire n4731_lo_n_spl_0001;
  wire n4731_lo_n_spl_001;
  wire n4731_lo_n_spl_0010;
  wire n4731_lo_n_spl_0011;
  wire n4731_lo_n_spl_01;
  wire n4731_lo_n_spl_010;
  wire n4731_lo_n_spl_0100;
  wire n4731_lo_n_spl_0101;
  wire n4731_lo_n_spl_011;
  wire n4731_lo_n_spl_0110;
  wire n4731_lo_n_spl_0111;
  wire n4731_lo_n_spl_1;
  wire n4731_lo_n_spl_10;
  wire n4731_lo_n_spl_100;
  wire n4731_lo_n_spl_101;
  wire n4731_lo_n_spl_11;
  wire n4731_lo_n_spl_110;
  wire n4731_lo_n_spl_111;
  wire g1566_n_spl_;
  wire g1566_n_spl_0;
  wire g1566_p_spl_;
  wire g1566_p_spl_0;
  wire g1570_n_spl_;
  wire n2631_lo_p_spl_;
  wire n2631_lo_p_spl_0;
  wire n2631_lo_n_spl_;
  wire n2631_lo_n_spl_0;
  wire g1581_n_spl_;
  wire G3228_o2_p_spl_;
  wire G4137_o2_n_spl_;
  wire G3228_o2_n_spl_;
  wire G4137_o2_p_spl_;
  wire g1592_p_spl_;
  wire g1592_p_spl_0;
  wire g1592_p_spl_00;
  wire g1592_p_spl_1;
  wire g1592_n_spl_;
  wire g1592_n_spl_0;
  wire g1592_n_spl_00;
  wire g1592_n_spl_1;
  wire g1596_p_spl_;
  wire g1596_n_spl_;
  wire G2752_o2_n_spl_;
  wire g1563_n_spl_;
  wire g1563_n_spl_0;
  wire g1563_n_spl_00;
  wire g1563_n_spl_1;
  wire n4683_lo_p_spl_;
  wire n4683_lo_p_spl_0;
  wire n4683_lo_p_spl_00;
  wire n4683_lo_p_spl_000;
  wire n4683_lo_p_spl_0000;
  wire n4683_lo_p_spl_0001;
  wire n4683_lo_p_spl_001;
  wire n4683_lo_p_spl_0010;
  wire n4683_lo_p_spl_0011;
  wire n4683_lo_p_spl_01;
  wire n4683_lo_p_spl_010;
  wire n4683_lo_p_spl_011;
  wire n4683_lo_p_spl_1;
  wire n4683_lo_p_spl_10;
  wire n4683_lo_p_spl_100;
  wire n4683_lo_p_spl_101;
  wire n4683_lo_p_spl_11;
  wire n4683_lo_p_spl_110;
  wire n4683_lo_p_spl_111;
  wire n4671_lo_p_spl_;
  wire n4671_lo_p_spl_0;
  wire n4671_lo_p_spl_00;
  wire n4671_lo_p_spl_000;
  wire n4671_lo_p_spl_0000;
  wire n4671_lo_p_spl_0001;
  wire n4671_lo_p_spl_001;
  wire n4671_lo_p_spl_0010;
  wire n4671_lo_p_spl_0011;
  wire n4671_lo_p_spl_01;
  wire n4671_lo_p_spl_010;
  wire n4671_lo_p_spl_011;
  wire n4671_lo_p_spl_1;
  wire n4671_lo_p_spl_10;
  wire n4671_lo_p_spl_100;
  wire n4671_lo_p_spl_101;
  wire n4671_lo_p_spl_11;
  wire n4671_lo_p_spl_110;
  wire n4671_lo_p_spl_111;
  wire g1587_n_spl_;
  wire g1587_n_spl_0;
  wire g1587_n_spl_00;
  wire g1587_n_spl_1;
  wire n4683_lo_n_spl_;
  wire n4683_lo_n_spl_0;
  wire n4683_lo_n_spl_00;
  wire n4683_lo_n_spl_000;
  wire n4683_lo_n_spl_0000;
  wire n4683_lo_n_spl_0001;
  wire n4683_lo_n_spl_001;
  wire n4683_lo_n_spl_0010;
  wire n4683_lo_n_spl_0011;
  wire n4683_lo_n_spl_01;
  wire n4683_lo_n_spl_010;
  wire n4683_lo_n_spl_011;
  wire n4683_lo_n_spl_1;
  wire n4683_lo_n_spl_10;
  wire n4683_lo_n_spl_100;
  wire n4683_lo_n_spl_101;
  wire n4683_lo_n_spl_11;
  wire n4683_lo_n_spl_110;
  wire n4683_lo_n_spl_111;
  wire n2643_lo_p_spl_;
  wire n4671_lo_n_spl_;
  wire n4671_lo_n_spl_0;
  wire n4671_lo_n_spl_00;
  wire n4671_lo_n_spl_000;
  wire n4671_lo_n_spl_0000;
  wire n4671_lo_n_spl_0001;
  wire n4671_lo_n_spl_001;
  wire n4671_lo_n_spl_0010;
  wire n4671_lo_n_spl_0011;
  wire n4671_lo_n_spl_01;
  wire n4671_lo_n_spl_010;
  wire n4671_lo_n_spl_011;
  wire n4671_lo_n_spl_1;
  wire n4671_lo_n_spl_10;
  wire n4671_lo_n_spl_100;
  wire n4671_lo_n_spl_101;
  wire n4671_lo_n_spl_11;
  wire n4671_lo_n_spl_110;
  wire n4671_lo_n_spl_111;
  wire n2871_lo_p_spl_;
  wire g1616_p_spl_;
  wire g1616_n_spl_;
  wire g1618_p_spl_;
  wire g1618_n_spl_;
  wire g1621_p_spl_;
  wire g1621_n_spl_;
  wire g1629_n_spl_;
  wire g1643_n_spl_;
  wire g1658_n_spl_;
  wire n4695_lo_p_spl_;
  wire n4695_lo_p_spl_0;
  wire n4695_lo_p_spl_00;
  wire n4695_lo_p_spl_000;
  wire n4695_lo_p_spl_0000;
  wire n4695_lo_p_spl_0001;
  wire n4695_lo_p_spl_001;
  wire n4695_lo_p_spl_0010;
  wire n4695_lo_p_spl_0011;
  wire n4695_lo_p_spl_01;
  wire n4695_lo_p_spl_010;
  wire n4695_lo_p_spl_011;
  wire n4695_lo_p_spl_1;
  wire n4695_lo_p_spl_10;
  wire n4695_lo_p_spl_100;
  wire n4695_lo_p_spl_101;
  wire n4695_lo_p_spl_11;
  wire n4695_lo_p_spl_110;
  wire n4695_lo_p_spl_111;
  wire n4707_lo_p_spl_;
  wire n4707_lo_p_spl_0;
  wire n4707_lo_p_spl_00;
  wire n4707_lo_p_spl_000;
  wire n4707_lo_p_spl_0000;
  wire n4707_lo_p_spl_0001;
  wire n4707_lo_p_spl_001;
  wire n4707_lo_p_spl_0010;
  wire n4707_lo_p_spl_0011;
  wire n4707_lo_p_spl_01;
  wire n4707_lo_p_spl_010;
  wire n4707_lo_p_spl_011;
  wire n4707_lo_p_spl_1;
  wire n4707_lo_p_spl_10;
  wire n4707_lo_p_spl_100;
  wire n4707_lo_p_spl_101;
  wire n4707_lo_p_spl_11;
  wire n4707_lo_p_spl_110;
  wire n4707_lo_p_spl_111;
  wire n4695_lo_n_spl_;
  wire n4695_lo_n_spl_0;
  wire n4695_lo_n_spl_00;
  wire n4695_lo_n_spl_000;
  wire n4695_lo_n_spl_0000;
  wire n4695_lo_n_spl_0001;
  wire n4695_lo_n_spl_001;
  wire n4695_lo_n_spl_0010;
  wire n4695_lo_n_spl_0011;
  wire n4695_lo_n_spl_01;
  wire n4695_lo_n_spl_010;
  wire n4695_lo_n_spl_011;
  wire n4695_lo_n_spl_1;
  wire n4695_lo_n_spl_10;
  wire n4695_lo_n_spl_100;
  wire n4695_lo_n_spl_101;
  wire n4695_lo_n_spl_11;
  wire n4695_lo_n_spl_110;
  wire n4695_lo_n_spl_111;
  wire n4707_lo_n_spl_;
  wire n4707_lo_n_spl_0;
  wire n4707_lo_n_spl_00;
  wire n4707_lo_n_spl_000;
  wire n4707_lo_n_spl_0000;
  wire n4707_lo_n_spl_0001;
  wire n4707_lo_n_spl_001;
  wire n4707_lo_n_spl_0010;
  wire n4707_lo_n_spl_0011;
  wire n4707_lo_n_spl_01;
  wire n4707_lo_n_spl_010;
  wire n4707_lo_n_spl_011;
  wire n4707_lo_n_spl_1;
  wire n4707_lo_n_spl_10;
  wire n4707_lo_n_spl_100;
  wire n4707_lo_n_spl_101;
  wire n4707_lo_n_spl_11;
  wire n4707_lo_n_spl_110;
  wire n4707_lo_n_spl_111;
  wire g1679_p_spl_;
  wire g1679_n_spl_;
  wire g1681_p_spl_;
  wire g1681_n_spl_;
  wire g1683_p_spl_;
  wire g1683_p_spl_0;
  wire g1683_n_spl_;
  wire g1683_n_spl_0;
  wire g1685_p_spl_;
  wire g1685_n_spl_;
  wire g1693_n_spl_;
  wire g1707_n_spl_;
  wire g1722_n_spl_;
  wire g1734_n_spl_;
  wire g1746_p_spl_;
  wire g1743_n_spl_;
  wire g1746_n_spl_;
  wire g1743_p_spl_;
  wire g1751_p_spl_;
  wire g1751_p_spl_0;
  wire g1751_p_spl_1;
  wire g1750_n_spl_;
  wire g1750_n_spl_0;
  wire g1750_n_spl_1;
  wire g1751_n_spl_;
  wire g1751_n_spl_0;
  wire g1751_n_spl_1;
  wire g1750_p_spl_;
  wire g1750_p_spl_0;
  wire g1750_p_spl_1;
  wire G3674_o2_p_spl_;
  wire G3674_o2_p_spl_0;
  wire G3674_o2_p_spl_1;
  wire G3674_o2_n_spl_;
  wire G3674_o2_n_spl_0;
  wire G3674_o2_n_spl_1;
  wire g1771_p_spl_;
  wire g1768_n_spl_;
  wire g1771_n_spl_;
  wire g1768_p_spl_;
  wire g1776_p_spl_;
  wire g1776_p_spl_0;
  wire g1776_p_spl_1;
  wire g1775_n_spl_;
  wire g1775_n_spl_0;
  wire g1775_n_spl_1;
  wire g1776_n_spl_;
  wire g1776_n_spl_0;
  wire g1776_n_spl_1;
  wire g1775_p_spl_;
  wire g1775_p_spl_0;
  wire g1775_p_spl_1;
  wire G3685_o2_n_spl_;
  wire G3685_o2_n_spl_0;
  wire G3685_o2_n_spl_1;
  wire G3685_o2_p_spl_;
  wire G3685_o2_p_spl_0;
  wire G3685_o2_p_spl_1;
  wire g1792_p_spl_;
  wire g1792_p_spl_0;
  wire g1792_p_spl_1;
  wire g1792_n_spl_;
  wire g1792_n_spl_0;
  wire g1792_n_spl_1;
  wire g1795_n_spl_;
  wire g1804_n_spl_;
  wire g1815_n_spl_;
  wire g1827_n_spl_;
  wire g1838_n_spl_;
  wire g1847_n_spl_;
  wire g1858_n_spl_;
  wire g1601_n_spl_;
  wire g1601_n_spl_0;
  wire g1601_n_spl_1;
  wire n4503_lo_p_spl_;
  wire n4503_lo_p_spl_0;
  wire n4503_lo_p_spl_00;
  wire n4503_lo_p_spl_000;
  wire n4503_lo_p_spl_0000;
  wire n4503_lo_p_spl_0001;
  wire n4503_lo_p_spl_001;
  wire n4503_lo_p_spl_0010;
  wire n4503_lo_p_spl_0011;
  wire n4503_lo_p_spl_01;
  wire n4503_lo_p_spl_010;
  wire n4503_lo_p_spl_011;
  wire n4503_lo_p_spl_1;
  wire n4503_lo_p_spl_10;
  wire n4503_lo_p_spl_100;
  wire n4503_lo_p_spl_101;
  wire n4503_lo_p_spl_11;
  wire n4503_lo_p_spl_110;
  wire n4503_lo_p_spl_111;
  wire n4515_lo_p_spl_;
  wire n4515_lo_p_spl_0;
  wire n4515_lo_p_spl_00;
  wire n4515_lo_p_spl_000;
  wire n4515_lo_p_spl_0000;
  wire n4515_lo_p_spl_0001;
  wire n4515_lo_p_spl_001;
  wire n4515_lo_p_spl_0010;
  wire n4515_lo_p_spl_0011;
  wire n4515_lo_p_spl_01;
  wire n4515_lo_p_spl_010;
  wire n4515_lo_p_spl_011;
  wire n4515_lo_p_spl_1;
  wire n4515_lo_p_spl_10;
  wire n4515_lo_p_spl_100;
  wire n4515_lo_p_spl_101;
  wire n4515_lo_p_spl_11;
  wire n4515_lo_p_spl_110;
  wire n4515_lo_p_spl_111;
  wire n4503_lo_n_spl_;
  wire n4503_lo_n_spl_0;
  wire n4503_lo_n_spl_00;
  wire n4503_lo_n_spl_000;
  wire n4503_lo_n_spl_0000;
  wire n4503_lo_n_spl_0001;
  wire n4503_lo_n_spl_001;
  wire n4503_lo_n_spl_0010;
  wire n4503_lo_n_spl_0011;
  wire n4503_lo_n_spl_01;
  wire n4503_lo_n_spl_010;
  wire n4503_lo_n_spl_011;
  wire n4503_lo_n_spl_1;
  wire n4503_lo_n_spl_10;
  wire n4503_lo_n_spl_100;
  wire n4503_lo_n_spl_101;
  wire n4503_lo_n_spl_11;
  wire n4503_lo_n_spl_110;
  wire n4503_lo_n_spl_111;
  wire n3567_lo_p_spl_;
  wire n4515_lo_n_spl_;
  wire n4515_lo_n_spl_0;
  wire n4515_lo_n_spl_00;
  wire n4515_lo_n_spl_000;
  wire n4515_lo_n_spl_0000;
  wire n4515_lo_n_spl_0001;
  wire n4515_lo_n_spl_001;
  wire n4515_lo_n_spl_0010;
  wire n4515_lo_n_spl_0011;
  wire n4515_lo_n_spl_01;
  wire n4515_lo_n_spl_010;
  wire n4515_lo_n_spl_011;
  wire n4515_lo_n_spl_1;
  wire n4515_lo_n_spl_10;
  wire n4515_lo_n_spl_100;
  wire n4515_lo_n_spl_101;
  wire n4515_lo_n_spl_11;
  wire n4515_lo_n_spl_110;
  wire n4515_lo_n_spl_111;
  wire n3579_lo_p_spl_;
  wire n3375_lo_p_spl_;
  wire n3375_lo_p_spl_0;
  wire n3375_lo_p_spl_00;
  wire n3375_lo_p_spl_000;
  wire n3375_lo_p_spl_0000;
  wire n3375_lo_p_spl_0001;
  wire n3375_lo_p_spl_001;
  wire n3375_lo_p_spl_0010;
  wire n3375_lo_p_spl_0011;
  wire n3375_lo_p_spl_01;
  wire n3375_lo_p_spl_010;
  wire n3375_lo_p_spl_0100;
  wire n3375_lo_p_spl_011;
  wire n3375_lo_p_spl_1;
  wire n3375_lo_p_spl_10;
  wire n3375_lo_p_spl_100;
  wire n3375_lo_p_spl_101;
  wire n3375_lo_p_spl_11;
  wire n3375_lo_p_spl_110;
  wire n3375_lo_p_spl_111;
  wire n4527_lo_p_spl_;
  wire n4527_lo_p_spl_0;
  wire n4527_lo_p_spl_00;
  wire n4527_lo_p_spl_000;
  wire n4527_lo_p_spl_0000;
  wire n4527_lo_p_spl_0001;
  wire n4527_lo_p_spl_001;
  wire n4527_lo_p_spl_0010;
  wire n4527_lo_p_spl_0011;
  wire n4527_lo_p_spl_01;
  wire n4527_lo_p_spl_010;
  wire n4527_lo_p_spl_011;
  wire n4527_lo_p_spl_1;
  wire n4527_lo_p_spl_10;
  wire n4527_lo_p_spl_100;
  wire n4527_lo_p_spl_101;
  wire n4527_lo_p_spl_11;
  wire n4527_lo_p_spl_110;
  wire n4527_lo_p_spl_111;
  wire n4539_lo_p_spl_;
  wire n4539_lo_p_spl_0;
  wire n4539_lo_p_spl_00;
  wire n4539_lo_p_spl_000;
  wire n4539_lo_p_spl_0000;
  wire n4539_lo_p_spl_0001;
  wire n4539_lo_p_spl_001;
  wire n4539_lo_p_spl_0010;
  wire n4539_lo_p_spl_0011;
  wire n4539_lo_p_spl_01;
  wire n4539_lo_p_spl_010;
  wire n4539_lo_p_spl_011;
  wire n4539_lo_p_spl_1;
  wire n4539_lo_p_spl_10;
  wire n4539_lo_p_spl_100;
  wire n4539_lo_p_spl_101;
  wire n4539_lo_p_spl_11;
  wire n4539_lo_p_spl_110;
  wire n4539_lo_p_spl_111;
  wire n4527_lo_n_spl_;
  wire n4527_lo_n_spl_0;
  wire n4527_lo_n_spl_00;
  wire n4527_lo_n_spl_000;
  wire n4527_lo_n_spl_0000;
  wire n4527_lo_n_spl_0001;
  wire n4527_lo_n_spl_001;
  wire n4527_lo_n_spl_0010;
  wire n4527_lo_n_spl_0011;
  wire n4527_lo_n_spl_01;
  wire n4527_lo_n_spl_010;
  wire n4527_lo_n_spl_011;
  wire n4527_lo_n_spl_1;
  wire n4527_lo_n_spl_10;
  wire n4527_lo_n_spl_100;
  wire n4527_lo_n_spl_101;
  wire n4527_lo_n_spl_11;
  wire n4527_lo_n_spl_110;
  wire n4527_lo_n_spl_111;
  wire n4539_lo_n_spl_;
  wire n4539_lo_n_spl_0;
  wire n4539_lo_n_spl_00;
  wire n4539_lo_n_spl_000;
  wire n4539_lo_n_spl_0000;
  wire n4539_lo_n_spl_0001;
  wire n4539_lo_n_spl_001;
  wire n4539_lo_n_spl_0010;
  wire n4539_lo_n_spl_0011;
  wire n4539_lo_n_spl_01;
  wire n4539_lo_n_spl_010;
  wire n4539_lo_n_spl_011;
  wire n4539_lo_n_spl_1;
  wire n4539_lo_n_spl_10;
  wire n4539_lo_n_spl_100;
  wire n4539_lo_n_spl_101;
  wire n4539_lo_n_spl_11;
  wire n4539_lo_n_spl_110;
  wire n4539_lo_n_spl_111;
  wire g1635_n_spl_;
  wire g1635_n_spl_0;
  wire g1635_n_spl_00;
  wire g1635_n_spl_1;
  wire g1699_n_spl_;
  wire g1699_n_spl_0;
  wire g1699_n_spl_00;
  wire g1699_n_spl_1;
  wire n2799_lo_p_spl_;
  wire n2775_lo_p_spl_;
  wire g1649_n_spl_;
  wire g1649_n_spl_0;
  wire g1649_n_spl_00;
  wire g1649_n_spl_1;
  wire g1713_n_spl_;
  wire g1713_n_spl_0;
  wire g1713_n_spl_00;
  wire g1713_n_spl_1;
  wire n2931_lo_p_spl_;
  wire n2679_lo_p_spl_;
  wire g1664_n_spl_;
  wire g1664_n_spl_0;
  wire g1664_n_spl_00;
  wire g1664_n_spl_1;
  wire g1728_n_spl_;
  wire g1728_n_spl_0;
  wire g1728_n_spl_00;
  wire g1728_n_spl_1;
  wire n2919_lo_p_spl_;
  wire n2667_lo_p_spl_;
  wire g1576_n_spl_;
  wire g1576_n_spl_0;
  wire g1576_n_spl_00;
  wire g1576_n_spl_1;
  wire g1740_n_spl_;
  wire g1740_n_spl_0;
  wire g1740_n_spl_00;
  wire g1740_n_spl_1;
  wire n2895_lo_p_spl_;
  wire n2907_lo_p_spl_;
  wire n3639_lo_p_spl_;
  wire n3519_lo_p_spl_;
  wire n3591_lo_p_spl_;
  wire n3471_lo_p_spl_;
  wire n3459_lo_p_spl_;
  wire n3447_lo_p_spl_;
  wire n3435_lo_p_spl_;
  wire n3423_lo_p_spl_;
  wire g1271_p_spl_;
  wire n4659_lo_n_spl_;
  wire n4647_lo_n_spl_;
  wire n7463_o2_p_spl_;
  wire n3339_lo_p_spl_;
  wire n3339_lo_n_spl_;
  wire g2078_n_spl_;
  wire g2078_p_spl_;
  wire g2081_n_spl_;
  wire n4659_lo_p_spl_;
  wire n3255_lo_p_spl_;
  wire n4647_lo_p_spl_;
  wire g1601_p_spl_;
  wire g2092_n_spl_;
  wire n4467_lo_n_spl_;
  wire n4443_lo_n_spl_;
  wire g1765_n_spl_;
  wire n4479_lo_n_spl_;
  wire g1790_n_spl_;
  wire g1449_n_spl_;
  wire g1474_n_spl_;
  wire n3795_lo_n_spl_;
  wire n7156_o2_n_spl_;
  wire n7156_o2_p_spl_;
  wire g2103_n_spl_;
  wire g2103_n_spl_0;
  wire g2103_n_spl_00;
  wire g2103_n_spl_1;
  wire g2154_n_spl_;
  wire g2154_n_spl_0;
  wire g2154_n_spl_00;
  wire g2154_n_spl_1;
  wire n3111_lo_p_spl_;
  wire n3099_lo_p_spl_;
  wire g2111_n_spl_;
  wire g2111_n_spl_0;
  wire g2111_n_spl_00;
  wire g2111_n_spl_1;
  wire g2162_n_spl_;
  wire g2162_n_spl_0;
  wire g2162_n_spl_00;
  wire g2162_n_spl_1;
  wire n2811_lo_p_spl_;
  wire n2823_lo_p_spl_;
  wire g2119_n_spl_;
  wire g2119_n_spl_0;
  wire g2119_n_spl_00;
  wire g2119_n_spl_1;
  wire g2170_n_spl_;
  wire g2170_n_spl_0;
  wire g2170_n_spl_00;
  wire g2170_n_spl_1;
  wire n3075_lo_p_spl_;
  wire n3087_lo_p_spl_;
  wire g2127_n_spl_;
  wire g2127_n_spl_0;
  wire g2127_n_spl_00;
  wire g2127_n_spl_1;
  wire g2178_n_spl_;
  wire g2178_n_spl_0;
  wire g2178_n_spl_00;
  wire g2178_n_spl_1;
  wire n3039_lo_p_spl_;
  wire n2787_lo_p_spl_;
  wire n3651_lo_p_spl_;
  wire n3531_lo_p_spl_;
  wire n3627_lo_p_spl_;
  wire n3507_lo_p_spl_;
  wire n3615_lo_p_spl_;
  wire n3495_lo_p_spl_;
  wire n3603_lo_p_spl_;
  wire n3483_lo_p_spl_;
  wire g2365_n_spl_;
  wire g2370_p_spl_;
  wire g2375_n_spl_;
  wire g2381_n_spl_;
  wire g2386_p_spl_;
  wire g2399_n_spl_;
  wire g2399_n_spl_0;
  wire g2399_n_spl_1;
  wire g2407_n_spl_;
  wire g2407_n_spl_0;
  wire g2407_n_spl_1;
  wire n2655_lo_p_spl_;
  wire n2883_lo_p_spl_;
  wire n3543_lo_p_spl_;
  wire n3555_lo_p_spl_;
  wire n2968_inv_n_spl_;
  wire n2968_inv_n_spl_0;
  wire n2968_inv_n_spl_00;
  wire n2968_inv_n_spl_01;
  wire n2968_inv_n_spl_1;
  wire n2968_inv_n_spl_10;
  wire n2968_inv_n_spl_11;
  wire n4308_lo_buf_o2_p_spl_;
  wire n4308_lo_buf_o2_p_spl_0;
  wire n4308_lo_buf_o2_p_spl_00;
  wire n4308_lo_buf_o2_p_spl_1;
  wire n2968_inv_p_spl_;
  wire n2968_inv_p_spl_0;
  wire n2968_inv_p_spl_00;
  wire n2968_inv_p_spl_000;
  wire n2968_inv_p_spl_01;
  wire n2968_inv_p_spl_1;
  wire n2968_inv_p_spl_10;
  wire n2968_inv_p_spl_11;
  wire n4308_lo_buf_o2_n_spl_;
  wire n4308_lo_buf_o2_n_spl_0;
  wire n4308_lo_buf_o2_n_spl_1;
  wire n2974_inv_n_spl_;
  wire n2974_inv_n_spl_0;
  wire n2974_inv_n_spl_00;
  wire n2974_inv_n_spl_01;
  wire n2974_inv_n_spl_1;
  wire n2974_inv_n_spl_10;
  wire n2974_inv_p_spl_;
  wire n2974_inv_p_spl_0;
  wire n2974_inv_p_spl_00;
  wire n2974_inv_p_spl_01;
  wire n2974_inv_p_spl_1;
  wire n2974_inv_p_spl_10;
  wire n2974_inv_p_spl_11;
  wire n3121_inv_n_spl_;
  wire n3121_inv_n_spl_0;
  wire n3121_inv_n_spl_00;
  wire n3121_inv_n_spl_01;
  wire n3121_inv_n_spl_1;
  wire n3121_inv_n_spl_10;
  wire n3121_inv_n_spl_11;
  wire G1873_o2_p_spl_;
  wire n3121_inv_p_spl_;
  wire n3121_inv_p_spl_0;
  wire n3121_inv_p_spl_00;
  wire n3121_inv_p_spl_000;
  wire n3121_inv_p_spl_01;
  wire n3121_inv_p_spl_1;
  wire n3121_inv_p_spl_10;
  wire n3121_inv_p_spl_11;
  wire G1873_o2_n_spl_;
  wire n3124_inv_n_spl_;
  wire n3124_inv_n_spl_0;
  wire n3124_inv_n_spl_00;
  wire n3124_inv_n_spl_01;
  wire n3124_inv_n_spl_1;
  wire n3124_inv_n_spl_10;
  wire n3124_inv_p_spl_;
  wire n3124_inv_p_spl_0;
  wire n3124_inv_p_spl_00;
  wire n3124_inv_p_spl_01;
  wire n3124_inv_p_spl_1;
  wire n3124_inv_p_spl_10;
  wire n3124_inv_p_spl_11;
  wire n6955_o2_p_spl_;
  wire n6955_o2_n_spl_;
  wire n6954_o2_p_spl_;
  wire n6954_o2_p_spl_0;
  wire n6954_o2_p_spl_00;
  wire n6954_o2_p_spl_01;
  wire n6954_o2_p_spl_1;
  wire n6954_o2_p_spl_10;
  wire n6954_o2_n_spl_;
  wire n6954_o2_n_spl_0;
  wire n6954_o2_n_spl_00;
  wire n6954_o2_n_spl_01;
  wire n6954_o2_n_spl_1;
  wire n6954_o2_n_spl_10;
  wire n7387_o2_p_spl_;
  wire n7387_o2_p_spl_0;
  wire n7387_o2_p_spl_00;
  wire n7387_o2_p_spl_01;
  wire n7387_o2_p_spl_1;
  wire n7387_o2_n_spl_;
  wire n7387_o2_n_spl_0;
  wire n7387_o2_n_spl_00;
  wire n7387_o2_n_spl_01;
  wire n7387_o2_n_spl_1;
  wire G3495_o2_p_spl_;
  wire G3495_o2_p_spl_0;
  wire G3495_o2_p_spl_00;
  wire G3495_o2_p_spl_1;
  wire G3495_o2_n_spl_;
  wire G3495_o2_n_spl_0;
  wire G3495_o2_n_spl_00;
  wire G3495_o2_n_spl_1;
  wire n6957_o2_p_spl_;
  wire n6957_o2_n_spl_;
  wire n6956_o2_p_spl_;
  wire n6956_o2_p_spl_0;
  wire n6956_o2_p_spl_00;
  wire n6956_o2_p_spl_01;
  wire n6956_o2_p_spl_1;
  wire n6956_o2_p_spl_10;
  wire n6956_o2_n_spl_;
  wire n6956_o2_n_spl_0;
  wire n6956_o2_n_spl_00;
  wire n6956_o2_n_spl_01;
  wire n6956_o2_n_spl_1;
  wire n6956_o2_n_spl_10;
  wire n7386_o2_p_spl_;
  wire n7386_o2_p_spl_0;
  wire n7386_o2_p_spl_00;
  wire n7386_o2_p_spl_01;
  wire n7386_o2_p_spl_1;
  wire n7386_o2_n_spl_;
  wire n7386_o2_n_spl_0;
  wire n7386_o2_n_spl_00;
  wire n7386_o2_n_spl_01;
  wire n7386_o2_n_spl_1;
  wire G3621_o2_p_spl_;
  wire G3621_o2_p_spl_0;
  wire G3621_o2_p_spl_00;
  wire G3621_o2_p_spl_1;
  wire G3621_o2_n_spl_;
  wire G3621_o2_n_spl_0;
  wire G3621_o2_n_spl_00;
  wire G3621_o2_n_spl_1;
  wire G2404_o2_p_spl_;
  wire G2404_o2_p_spl_0;
  wire G2404_o2_p_spl_1;
  wire n4296_lo_buf_o2_p_spl_;
  wire n4296_lo_buf_o2_p_spl_0;
  wire n4296_lo_buf_o2_p_spl_1;
  wire G2404_o2_n_spl_;
  wire G2404_o2_n_spl_0;
  wire n4296_lo_buf_o2_n_spl_;
  wire n4296_lo_buf_o2_n_spl_0;
  wire G2466_o2_p_spl_;
  wire G2466_o2_p_spl_0;
  wire G2466_o2_p_spl_1;
  wire n4368_lo_buf_o2_p_spl_;
  wire n4368_lo_buf_o2_p_spl_0;
  wire n4368_lo_buf_o2_p_spl_1;
  wire G2466_o2_n_spl_;
  wire G2466_o2_n_spl_0;
  wire n4368_lo_buf_o2_n_spl_;
  wire n4368_lo_buf_o2_n_spl_0;
  wire n6772_o2_n_spl_;
  wire n6772_o2_n_spl_0;
  wire n6772_o2_p_spl_;
  wire n6772_o2_p_spl_0;
  wire n6772_o2_p_spl_1;
  wire G2424_o2_p_spl_;
  wire n4320_lo_buf_o2_p_spl_;
  wire G1821_o2_p_spl_;
  wire n4053_lo_p_spl_;
  wire n4053_lo_p_spl_0;
  wire n4053_lo_p_spl_00;
  wire n4053_lo_p_spl_1;
  wire n4053_lo_n_spl_;
  wire G1060_o2_n_spl_;
  wire G1734_o2_p_spl_;
  wire n3753_lo_p_spl_;
  wire n3753_lo_p_spl_0;
  wire n3753_lo_p_spl_00;
  wire n3753_lo_p_spl_1;
  wire n3753_lo_n_spl_;
  wire G963_o2_n_spl_;
  wire n4164_lo_buf_o2_p_spl_;
  wire G1815_o2_p_spl_;
  wire G1815_o2_p_spl_0;
  wire G1815_o2_n_spl_;
  wire n4176_lo_buf_o2_p_spl_;
  wire n2662_inv_n_spl_;
  wire n2662_inv_p_spl_;
  wire n2662_inv_p_spl_0;
  wire n7136_o2_p_spl_;
  wire n7136_o2_p_spl_0;
  wire n7136_o2_p_spl_1;
  wire n7132_o2_p_spl_;
  wire n7132_o2_p_spl_0;
  wire n7132_o2_p_spl_00;
  wire n7132_o2_p_spl_01;
  wire n7132_o2_p_spl_1;
  wire n7132_o2_p_spl_10;
  wire n7023_o2_p_spl_;
  wire n7023_o2_p_spl_0;
  wire n7016_o2_p_spl_;
  wire n7016_o2_p_spl_0;
  wire n7016_o2_p_spl_00;
  wire n7016_o2_p_spl_01;
  wire n7016_o2_p_spl_1;
  wire n7022_o2_n_spl_;
  wire n7022_o2_n_spl_0;
  wire n7017_o2_n_spl_;
  wire n7017_o2_n_spl_0;
  wire n7017_o2_n_spl_00;
  wire n7017_o2_n_spl_01;
  wire n7017_o2_n_spl_1;
  wire n7135_o2_n_spl_;
  wire n7133_o2_n_spl_;
  wire n7133_o2_n_spl_0;
  wire n7133_o2_n_spl_00;
  wire n7133_o2_n_spl_1;
  wire n4272_lo_buf_o2_p_spl_;
  wire G2386_o2_p_spl_;
  wire n4404_lo_buf_o2_p_spl_;
  wire G2454_o2_p_spl_;
  wire n7384_o2_p_spl_;
  wire n7384_o2_p_spl_0;
  wire n7383_o2_n_spl_;
  wire n7383_o2_n_spl_0;
  wire n7383_o2_n_spl_1;
  wire n7384_o2_n_spl_;
  wire n7383_o2_p_spl_;
  wire n7383_o2_p_spl_0;
  wire n7383_o2_p_spl_00;
  wire n7383_o2_p_spl_01;
  wire n7383_o2_p_spl_1;
  wire n7016_o2_n_spl_;
  wire n7016_o2_n_spl_0;
  wire n7016_o2_n_spl_1;
  wire n7023_o2_n_spl_;
  wire n7022_o2_p_spl_;
  wire n7022_o2_p_spl_0;
  wire n7022_o2_p_spl_1;
  wire n7017_o2_p_spl_;
  wire n7017_o2_p_spl_0;
  wire n7017_o2_p_spl_00;
  wire n7017_o2_p_spl_01;
  wire n7017_o2_p_spl_1;
  wire n4224_lo_buf_o2_p_spl_;
  wire n4224_lo_buf_o2_p_spl_0;
  wire n4224_lo_buf_o2_p_spl_00;
  wire n4224_lo_buf_o2_p_spl_1;
  wire G2379_o2_p_spl_;
  wire G2379_o2_p_spl_0;
  wire G2379_o2_p_spl_00;
  wire G2379_o2_p_spl_1;
  wire n4224_lo_buf_o2_n_spl_;
  wire n4224_lo_buf_o2_n_spl_0;
  wire n4224_lo_buf_o2_n_spl_1;
  wire G2379_o2_n_spl_;
  wire G2379_o2_n_spl_0;
  wire G2379_o2_n_spl_1;
  wire G1356_o2_p_spl_;
  wire G2933_o2_n_spl_;
  wire G1356_o2_n_spl_;
  wire G2933_o2_p_spl_;
  wire G1359_o2_p_spl_;
  wire G2936_o2_n_spl_;
  wire G1359_o2_n_spl_;
  wire G2936_o2_p_spl_;
  wire G1398_o2_p_spl_;
  wire G2975_o2_n_spl_;
  wire G1398_o2_n_spl_;
  wire G2975_o2_p_spl_;
  wire G1401_o2_p_spl_;
  wire G2978_o2_n_spl_;
  wire G1401_o2_n_spl_;
  wire G2978_o2_p_spl_;
  wire n4260_lo_buf_o2_p_spl_;
  wire G2392_o2_p_spl_;
  wire n4392_lo_buf_o2_p_spl_;
  wire G2460_o2_p_spl_;
  wire n4098_lo_p_spl_;
  wire G1728_o2_p_spl_;
  wire n3834_lo_p_spl_;
  wire n2665_inv_p_spl_;
  wire n4080_lo_buf_o2_p_spl_;
  wire n4080_lo_buf_o2_p_spl_0;
  wire n4080_lo_buf_o2_p_spl_00;
  wire n4080_lo_buf_o2_p_spl_01;
  wire n4080_lo_buf_o2_p_spl_1;
  wire n4080_lo_buf_o2_p_spl_10;
  wire n4002_lo_p_spl_;
  wire n4080_lo_buf_o2_n_spl_;
  wire n4080_lo_buf_o2_n_spl_0;
  wire n4080_lo_buf_o2_n_spl_00;
  wire n4080_lo_buf_o2_n_spl_1;
  wire n4092_lo_buf_o2_p_spl_;
  wire n4092_lo_buf_o2_p_spl_0;
  wire n4092_lo_buf_o2_p_spl_00;
  wire n4092_lo_buf_o2_p_spl_01;
  wire n4092_lo_buf_o2_p_spl_1;
  wire n4092_lo_buf_o2_p_spl_10;
  wire n3702_lo_p_spl_;
  wire n4092_lo_buf_o2_n_spl_;
  wire n4092_lo_buf_o2_n_spl_0;
  wire n4092_lo_buf_o2_n_spl_00;
  wire n4092_lo_buf_o2_n_spl_1;
  wire g2565_p_spl_;
  wire g2452_p_spl_;
  wire g2452_p_spl_0;
  wire g2452_p_spl_1;
  wire g2565_n_spl_;
  wire g2452_n_spl_;
  wire g2452_n_spl_0;
  wire g2452_n_spl_00;
  wire g2452_n_spl_1;
  wire G3474_o2_p_spl_;
  wire G3474_o2_p_spl_0;
  wire G3474_o2_n_spl_;
  wire g2571_p_spl_;
  wire g2485_n_spl_;
  wire g2485_n_spl_0;
  wire n4488_lo_p_spl_;
  wire n4488_lo_p_spl_0;
  wire g2576_p_spl_;
  wire g2576_n_spl_;
  wire g2582_p_spl_;
  wire g2485_p_spl_;
  wire g2466_p_spl_;
  wire n4488_lo_n_spl_;
  wire n4488_lo_n_spl_0;
  wire g2593_p_spl_;
  wire g2593_n_spl_;
  wire g2603_p_spl_;
  wire g2603_n_spl_;
  wire g2614_p_spl_;
  wire G2492_o2_p_spl_;
  wire G2492_o2_p_spl_0;
  wire G2492_o2_p_spl_00;
  wire G2492_o2_p_spl_000;
  wire G2492_o2_p_spl_001;
  wire G2492_o2_p_spl_01;
  wire G2492_o2_p_spl_1;
  wire G2492_o2_p_spl_10;
  wire G2492_o2_p_spl_11;
  wire g2614_n_spl_;
  wire G2492_o2_n_spl_;
  wire G2492_o2_n_spl_0;
  wire G2492_o2_n_spl_1;
  wire n2341_inv_p_spl_;
  wire n2341_inv_p_spl_0;
  wire n2341_inv_n_spl_;
  wire g2620_n_spl_;
  wire g2500_p_spl_;
  wire n4548_lo_n_spl_;
  wire n4548_lo_n_spl_0;
  wire g2625_p_spl_;
  wire g2625_n_spl_;
  wire g2631_n_spl_;
  wire g2500_n_spl_;
  wire g2500_n_spl_0;
  wire g2470_p_spl_;
  wire n4548_lo_p_spl_;
  wire n4548_lo_p_spl_0;
  wire g2642_p_spl_;
  wire g2642_n_spl_;
  wire g2652_p_spl_;
  wire g2652_n_spl_;
  wire n7132_o2_n_spl_;
  wire n7132_o2_n_spl_0;
  wire n7132_o2_n_spl_1;
  wire n7136_o2_n_spl_;
  wire G2430_o2_p_spl_;
  wire G2430_o2_p_spl_0;
  wire G2430_o2_n_spl_;
  wire n7135_o2_p_spl_;
  wire n7135_o2_p_spl_0;
  wire n7135_o2_p_spl_1;
  wire n7133_o2_p_spl_;
  wire n7133_o2_p_spl_0;
  wire n7133_o2_p_spl_00;
  wire n7133_o2_p_spl_01;
  wire n7133_o2_p_spl_1;
  wire n3657_lo_p_spl_;
  wire n3657_lo_p_spl_0;
  wire n3657_lo_p_spl_00;
  wire n3657_lo_p_spl_1;
  wire n4293_lo_p_spl_;
  wire n4293_lo_p_spl_0;
  wire n4293_lo_p_spl_1;
  wire g2514_n_spl_;
  wire n4365_lo_p_spl_;
  wire n4365_lo_p_spl_0;
  wire n4365_lo_p_spl_1;
  wire g2511_n_spl_;
  wire n4026_lo_p_spl_;
  wire n3726_lo_p_spl_;
  wire n6775_o2_p_spl_;
  wire n6775_o2_p_spl_0;
  wire n6775_o2_p_spl_1;
  wire n6774_o2_p_spl_;
  wire n6774_o2_p_spl_0;
  wire n6774_o2_p_spl_00;
  wire n6774_o2_p_spl_01;
  wire n6774_o2_p_spl_1;
  wire n7019_o2_p_spl_;
  wire n7019_o2_p_spl_0;
  wire n7019_o2_p_spl_1;
  wire n7015_o2_p_spl_;
  wire n7015_o2_p_spl_0;
  wire n7015_o2_p_spl_1;
  wire n6688_o2_p_spl_;
  wire n6688_o2_p_spl_0;
  wire n6688_o2_p_spl_1;
  wire n6682_o2_p_spl_;
  wire n6682_o2_p_spl_0;
  wire n6682_o2_p_spl_00;
  wire n6682_o2_p_spl_01;
  wire n6682_o2_p_spl_1;
  wire n6689_o2_p_spl_;
  wire n6689_o2_p_spl_0;
  wire n6689_o2_p_spl_1;
  wire n6683_o2_p_spl_;
  wire n6683_o2_p_spl_0;
  wire n6683_o2_p_spl_00;
  wire n6683_o2_p_spl_01;
  wire n6683_o2_p_spl_1;
  wire n7005_o2_p_spl_;
  wire n7005_o2_p_spl_0;
  wire n7018_o2_p_spl_;
  wire n7018_o2_p_spl_0;
  wire n7018_o2_p_spl_00;
  wire n7018_o2_p_spl_1;
  wire n6686_o2_p_spl_;
  wire n6686_o2_p_spl_0;
  wire n6684_o2_p_spl_;
  wire n6684_o2_p_spl_0;
  wire n6684_o2_p_spl_00;
  wire n6684_o2_p_spl_01;
  wire n6684_o2_p_spl_1;
  wire n6687_o2_p_spl_;
  wire n6687_o2_p_spl_0;
  wire n6685_o2_p_spl_;
  wire n6685_o2_p_spl_0;
  wire n6685_o2_p_spl_00;
  wire n6685_o2_p_spl_01;
  wire n6685_o2_p_spl_1;
  wire n6623_o2_p_spl_;
  wire n6621_o2_p_spl_;
  wire n6669_o2_n_spl_;
  wire n6669_o2_n_spl_0;
  wire n6669_o2_n_spl_00;
  wire n6669_o2_n_spl_1;
  wire n3936_lo_p_spl_;
  wire n6669_o2_p_spl_;
  wire n6669_o2_p_spl_0;
  wire n6669_o2_p_spl_00;
  wire n6669_o2_p_spl_01;
  wire n6669_o2_p_spl_1;
  wire n3936_lo_n_spl_;
  wire n6627_o2_p_spl_;
  wire n6625_o2_p_spl_;
  wire n4188_lo_p_spl_;
  wire g2529_n_spl_;
  wire g2529_n_spl_0;
  wire g2529_n_spl_1;
  wire g2518_p_spl_;
  wire g2702_p_spl_;
  wire g2702_p_spl_0;
  wire g2526_n_spl_;
  wire g2526_n_spl_0;
  wire g2526_n_spl_00;
  wire g2526_n_spl_1;
  wire g2519_p_spl_;
  wire g2519_p_spl_0;
  wire g2520_n_spl_;
  wire g2520_n_spl_0;
  wire G2486_o2_p_spl_;
  wire G2486_o2_p_spl_0;
  wire G2486_o2_p_spl_00;
  wire G2486_o2_p_spl_01;
  wire G2486_o2_p_spl_1;
  wire G2486_o2_p_spl_10;
  wire G2486_o2_p_spl_11;
  wire g2521_n_spl_;
  wire g2707_n_spl_;
  wire g2707_n_spl_0;
  wire n6686_o2_n_spl_;
  wire n6687_o2_n_spl_;
  wire g2714_n_spl_;
  wire n6833_o2_p_spl_;
  wire n6833_o2_p_spl_0;
  wire n6833_o2_p_spl_1;
  wire g2669_n_spl_;
  wire g2532_n_spl_;
  wire g2532_n_spl_0;
  wire g2719_p_spl_;
  wire g2663_n_spl_;
  wire g2723_p_spl_;
  wire g2704_p_spl_;
  wire g2562_p_spl_;
  wire g2703_p_spl_;
  wire g2706_n_spl_;
  wire g2709_n_spl_;
  wire n3756_lo_buf_o2_p_spl_;
  wire n6947_o2_p_spl_;
  wire n6774_o2_n_spl_;
  wire n6774_o2_n_spl_0;
  wire n6774_o2_n_spl_1;
  wire n7015_o2_n_spl_;
  wire n6682_o2_n_spl_;
  wire n6682_o2_n_spl_0;
  wire n6682_o2_n_spl_1;
  wire n6683_o2_n_spl_;
  wire n6683_o2_n_spl_0;
  wire n6683_o2_n_spl_1;
  wire n7018_o2_n_spl_;
  wire n7018_o2_n_spl_0;
  wire n7005_o2_n_spl_;
  wire n6684_o2_n_spl_;
  wire n6684_o2_n_spl_0;
  wire n6684_o2_n_spl_1;
  wire n6685_o2_n_spl_;
  wire n6685_o2_n_spl_0;
  wire n6685_o2_n_spl_1;
  wire n2965_inv_n_spl_;
  wire n2965_inv_n_spl_0;
  wire n2965_inv_n_spl_00;
  wire n2965_inv_n_spl_01;
  wire n2965_inv_n_spl_1;
  wire n2965_inv_p_spl_;
  wire n2965_inv_p_spl_0;
  wire n2965_inv_p_spl_00;
  wire n2965_inv_p_spl_01;
  wire n2965_inv_p_spl_1;
  wire n2965_inv_p_spl_10;
  wire G1138_o2_n_spl_;
  wire G1138_o2_p_spl_;
  wire n2971_inv_n_spl_;
  wire n2971_inv_n_spl_0;
  wire n2971_inv_n_spl_00;
  wire n2971_inv_n_spl_01;
  wire n2971_inv_n_spl_1;
  wire n2971_inv_p_spl_;
  wire n2971_inv_p_spl_0;
  wire n2971_inv_p_spl_00;
  wire n2971_inv_p_spl_01;
  wire n2971_inv_p_spl_1;
  wire n2971_inv_p_spl_10;
  wire n3118_inv_n_spl_;
  wire n3118_inv_n_spl_0;
  wire n3118_inv_n_spl_00;
  wire n3118_inv_n_spl_01;
  wire n3118_inv_n_spl_1;
  wire n3118_inv_n_spl_10;
  wire n3118_inv_n_spl_11;
  wire n6982_o2_n_spl_;
  wire n3118_inv_p_spl_;
  wire n3118_inv_p_spl_0;
  wire n3118_inv_p_spl_00;
  wire n3118_inv_p_spl_000;
  wire n3118_inv_p_spl_01;
  wire n3118_inv_p_spl_1;
  wire n3118_inv_p_spl_10;
  wire n3118_inv_p_spl_11;
  wire n6982_o2_p_spl_;
  wire n6982_o2_p_spl_0;
  wire n6982_o2_p_spl_00;
  wire n6982_o2_p_spl_1;
  wire n3127_inv_n_spl_;
  wire n3127_inv_n_spl_0;
  wire n3127_inv_n_spl_00;
  wire n3127_inv_n_spl_01;
  wire n3127_inv_n_spl_1;
  wire n3127_inv_n_spl_10;
  wire n3127_inv_n_spl_11;
  wire n3127_inv_p_spl_;
  wire n3127_inv_p_spl_0;
  wire n3127_inv_p_spl_00;
  wire n3127_inv_p_spl_000;
  wire n3127_inv_p_spl_01;
  wire n3127_inv_p_spl_1;
  wire n3127_inv_p_spl_10;
  wire n3127_inv_p_spl_11;
  wire G1132_o2_n_spl_;
  wire G1132_o2_p_spl_;
  wire n6945_o2_n_spl_;
  wire n6945_o2_p_spl_;
  wire n6945_o2_p_spl_0;
  wire n6945_o2_p_spl_00;
  wire n6945_o2_p_spl_1;
  wire g2787_n_spl_;
  wire g2777_p_spl_;
  wire g2787_p_spl_;
  wire g2777_n_spl_;
  wire G1126_o2_n_spl_;
  wire G1126_o2_p_spl_;
  wire n7175_o2_n_spl_;
  wire n7175_o2_p_spl_;
  wire n7175_o2_p_spl_0;
  wire n7175_o2_p_spl_00;
  wire n7175_o2_p_spl_1;
  wire g2800_p_spl_;
  wire g2462_p_spl_;
  wire g2800_n_spl_;
  wire g2462_n_spl_;
  wire g2462_n_spl_0;
  wire G1114_o2_n_spl_;
  wire G1114_o2_p_spl_;
  wire n6984_o2_n_spl_;
  wire n6984_o2_p_spl_;
  wire n6984_o2_p_spl_0;
  wire n6984_o2_p_spl_00;
  wire n6984_o2_p_spl_1;
  wire G1108_o2_n_spl_;
  wire G1108_o2_p_spl_;
  wire n6949_o2_n_spl_;
  wire n6949_o2_p_spl_;
  wire n6949_o2_p_spl_0;
  wire n6949_o2_p_spl_00;
  wire n6949_o2_p_spl_1;
  wire g2826_n_spl_;
  wire g2816_p_spl_;
  wire g2826_p_spl_;
  wire g2816_n_spl_;
  wire n7453_o2_n_spl_;
  wire n7453_o2_p_spl_;
  wire n7453_o2_p_spl_0;
  wire n7453_o2_p_spl_00;
  wire n7453_o2_p_spl_1;
  wire n3960_lo_buf_o2_n_spl_;
  wire n3960_lo_buf_o2_p_spl_;
  wire n3960_lo_buf_o2_p_spl_0;
  wire n3960_lo_buf_o2_p_spl_00;
  wire n3960_lo_buf_o2_p_spl_1;
  wire g2835_p_spl_;
  wire g2832_p_spl_;
  wire g2835_n_spl_;
  wire g2832_n_spl_;
  wire G1041_o2_n_spl_;
  wire G1041_o2_p_spl_;
  wire G1035_o2_n_spl_;
  wire G1035_o2_p_spl_;
  wire g2871_n_spl_;
  wire g2861_p_spl_;
  wire g2871_p_spl_;
  wire g2861_n_spl_;
  wire g2886_n_spl_;
  wire g2880_p_spl_;
  wire g2886_p_spl_;
  wire g2880_n_spl_;
  wire g2874_n_spl_;
  wire g2851_p_spl_;
  wire g2889_p_spl_;
  wire g2851_n_spl_;
  wire g2889_n_spl_;
  wire g2874_p_spl_;
  wire G1093_o2_n_spl_;
  wire G1093_o2_p_spl_;
  wire G1087_o2_n_spl_;
  wire G1087_o2_p_spl_;
  wire g2920_n_spl_;
  wire g2910_p_spl_;
  wire g2920_p_spl_;
  wire g2910_n_spl_;
  wire g2932_n_spl_;
  wire g2926_p_spl_;
  wire g2932_p_spl_;
  wire g2926_n_spl_;
  wire g2923_p_spl_;
  wire g2503_n_spl_;
  wire g2935_n_spl_;
  wire g2503_p_spl_;
  wire g2503_p_spl_0;
  wire g2935_p_spl_;
  wire g2923_n_spl_;
  wire g2684_n_spl_;
  wire g2684_n_spl_0;
  wire n4278_lo_p_spl_;
  wire n4278_lo_p_spl_0;
  wire g2681_n_spl_;
  wire g2681_n_spl_0;
  wire n4350_lo_p_spl_;
  wire n4350_lo_p_spl_0;
  wire G2727_o2_p_spl_;
  wire g2953_p_spl_;
  wire g2952_n_spl_;
  wire g2953_n_spl_;
  wire g2952_p_spl_;
  wire g2956_p_spl_;
  wire G3552_o2_n_spl_;
  wire G3552_o2_n_spl_0;
  wire G3552_o2_n_spl_1;
  wire g2956_n_spl_;
  wire G3552_o2_p_spl_;
  wire G3552_o2_p_spl_0;
  wire G3552_o2_p_spl_00;
  wire G3552_o2_p_spl_1;
  wire G3533_o2_p_spl_;
  wire G3533_o2_p_spl_0;
  wire G3533_o2_n_spl_;
  wire G2543_o2_p_spl_;
  wire g2967_p_spl_;
  wire g2966_n_spl_;
  wire g2967_n_spl_;
  wire g2966_p_spl_;
  wire g2970_p_spl_;
  wire n2647_inv_p_spl_;
  wire n2647_inv_p_spl_0;
  wire n2647_inv_p_spl_00;
  wire n2647_inv_p_spl_1;
  wire g2970_n_spl_;
  wire n2647_inv_n_spl_;
  wire n2647_inv_n_spl_0;
  wire n2647_inv_n_spl_1;
  wire G3645_o2_p_spl_;
  wire G3645_o2_p_spl_0;
  wire G3645_o2_n_spl_;
  wire g2507_n_spl_;
  wire g2507_n_spl_0;
  wire g2507_n_spl_1;
  wire G2715_o2_p_spl_;
  wire g2507_p_spl_;
  wire g2507_p_spl_0;
  wire G3485_o2_p_spl_;
  wire G3485_o2_p_spl_0;
  wire G3485_o2_p_spl_00;
  wire G3485_o2_p_spl_01;
  wire G3485_o2_p_spl_1;
  wire G3485_o2_p_spl_10;
  wire G2720_o2_p_spl_;
  wire G2720_o2_p_spl_0;
  wire G2720_o2_p_spl_1;
  wire G3485_o2_n_spl_;
  wire G2720_o2_n_spl_;
  wire G2720_o2_n_spl_0;
  wire G3546_o2_p_spl_;
  wire G3546_o2_p_spl_0;
  wire G3546_o2_p_spl_1;
  wire G3546_o2_n_spl_;
  wire G3546_o2_n_spl_0;
  wire g2508_p_spl_;
  wire g2983_p_spl_;
  wire g2983_p_spl_0;
  wire g2983_n_spl_;
  wire g2983_n_spl_0;
  wire G4051_o2_n_spl_;
  wire G4051_o2_n_spl_0;
  wire G4051_o2_p_spl_;
  wire G4051_o2_p_spl_0;
  wire G2410_o2_p_spl_;
  wire n4284_lo_buf_o2_p_spl_;
  wire g2986_n_spl_;
  wire g2985_n_spl_;
  wire g2986_p_spl_;
  wire g2985_p_spl_;
  wire g2989_p_spl_;
  wire g2984_n_spl_;
  wire g2989_n_spl_;
  wire g2984_p_spl_;
  wire g2998_p_spl_;
  wire g2998_n_spl_;
  wire g2504_p_spl_;
  wire g2504_p_spl_0;
  wire g2504_p_spl_1;
  wire G2832_o2_p_spl_;
  wire g2504_n_spl_;
  wire g2504_n_spl_0;
  wire g2504_n_spl_00;
  wire g2504_n_spl_01;
  wire g2504_n_spl_1;
  wire g2504_n_spl_10;
  wire G3611_o2_p_spl_;
  wire G3611_o2_p_spl_0;
  wire G3611_o2_p_spl_00;
  wire G3611_o2_p_spl_01;
  wire G3611_o2_p_spl_1;
  wire G3611_o2_p_spl_10;
  wire G2837_o2_p_spl_;
  wire G2837_o2_p_spl_0;
  wire G2837_o2_p_spl_1;
  wire G3611_o2_n_spl_;
  wire G2837_o2_n_spl_;
  wire G2837_o2_n_spl_0;
  wire G3658_o2_p_spl_;
  wire G3658_o2_p_spl_0;
  wire G3658_o2_p_spl_1;
  wire G3658_o2_n_spl_;
  wire G3658_o2_n_spl_0;
  wire g3011_p_spl_;
  wire g3011_p_spl_0;
  wire g3011_n_spl_;
  wire g3011_n_spl_0;
  wire G4065_o2_n_spl_;
  wire G4065_o2_n_spl_0;
  wire G4065_o2_p_spl_;
  wire G4065_o2_p_spl_0;
  wire G2472_o2_p_spl_;
  wire n4356_lo_buf_o2_p_spl_;
  wire g3014_n_spl_;
  wire g3013_n_spl_;
  wire g3014_p_spl_;
  wire g3013_p_spl_;
  wire g3017_p_spl_;
  wire g3012_n_spl_;
  wire g3017_n_spl_;
  wire g3012_p_spl_;
  wire g3026_p_spl_;
  wire g3026_n_spl_;
  wire n3678_lo_p_spl_;
  wire g2552_p_spl_;
  wire g2552_p_spl_0;
  wire n4374_lo_p_spl_;
  wire n4374_lo_p_spl_0;
  wire g2552_n_spl_;
  wire g2552_n_spl_0;
  wire n4374_lo_n_spl_;
  wire n4374_lo_n_spl_0;
  wire n4242_lo_p_spl_;
  wire n4242_lo_p_spl_0;
  wire g2555_n_spl_;
  wire g2555_n_spl_0;
  wire n4326_lo_p_spl_;
  wire n4326_lo_p_spl_0;
  wire g2561_n_spl_;
  wire g2561_n_spl_0;
  wire n4338_lo_p_spl_;
  wire n4338_lo_p_spl_0;
  wire g2558_n_spl_;
  wire g2558_n_spl_0;
  wire n4248_lo_buf_o2_p_spl_;
  wire n4248_lo_buf_o2_p_spl_0;
  wire n3801_lo_n_spl_;
  wire n3801_lo_n_spl_0;
  wire n3813_lo_n_spl_;
  wire n3813_lo_n_spl_0;
  wire n3840_lo_buf_o2_p_spl_;
  wire n3840_lo_buf_o2_p_spl_0;
  wire n3840_lo_buf_o2_p_spl_1;
  wire g2672_n_spl_;
  wire g2672_n_spl_0;
  wire n4305_lo_n_spl_;
  wire G4697_o2_p_spl_;
  wire G4131_o2_n_spl_;
  wire G4697_o2_n_spl_;
  wire G4131_o2_p_spl_;
  wire g3067_p_spl_;
  wire g3067_n_spl_;
  wire g3073_n_spl_;
  wire g2675_n_spl_;
  wire g2675_n_spl_0;
  wire g2675_n_spl_00;
  wire g2675_n_spl_1;
  wire G4706_o2_n_spl_;
  wire G4170_o2_n_spl_;
  wire G4706_o2_p_spl_;
  wire G4170_o2_p_spl_;
  wire g3077_p_spl_;
  wire g3077_n_spl_;
  wire g3083_n_spl_;
  wire g2678_n_spl_;
  wire g2678_n_spl_0;
  wire g2678_n_spl_00;
  wire g2678_n_spl_1;
  wire n3957_lo_p_spl_;
  wire n3969_lo_p_spl_;
  wire g2536_n_spl_;
  wire g2536_n_spl_0;
  wire g2536_n_spl_1;
  wire g2522_p_spl_;
  wire g2522_p_spl_0;
  wire g2536_p_spl_;
  wire g2536_p_spl_0;
  wire g2522_n_spl_;
  wire g3098_p_spl_;
  wire g3041_n_spl_;
  wire g3041_n_spl_0;
  wire g3041_n_spl_00;
  wire g3041_n_spl_1;
  wire g2542_n_spl_;
  wire g2542_n_spl_0;
  wire g2523_p_spl_;
  wire g2523_p_spl_0;
  wire g2542_p_spl_;
  wire g2542_p_spl_0;
  wire g2523_n_spl_;
  wire g3100_n_spl_;
  wire g3038_p_spl_;
  wire g3038_p_spl_0;
  wire g3038_p_spl_1;
  wire g2539_n_spl_;
  wire g2539_n_spl_0;
  wire g2539_n_spl_00;
  wire g2539_n_spl_01;
  wire g2539_n_spl_1;
  wire g2539_p_spl_;
  wire g2539_p_spl_0;
  wire g2533_p_spl_;
  wire g2533_p_spl_0;
  wire g2533_p_spl_00;
  wire g2533_p_spl_1;
  wire g2533_n_spl_;
  wire g2533_n_spl_0;
  wire g2533_n_spl_1;
  wire g3103_p_spl_;
  wire n3978_lo_p_spl_;
  wire g2550_n_spl_;
  wire g2550_n_spl_0;
  wire g3106_p_spl_;
  wire g2545_n_spl_;
  wire g2545_n_spl_0;
  wire g2545_p_spl_;
  wire g2545_p_spl_0;
  wire g2545_p_spl_1;
  wire g2517_p_spl_;
  wire g2517_p_spl_0;
  wire g2517_p_spl_1;
  wire g2517_n_spl_;
  wire g2517_n_spl_0;
  wire g2517_n_spl_00;
  wire g2517_n_spl_01;
  wire g2517_n_spl_1;
  wire g2517_n_spl_10;
  wire g2517_n_spl_11;
  wire g3110_n_spl_;
  wire g3112_n_spl_;
  wire g2546_p_spl_;
  wire g2546_p_spl_0;
  wire g2547_n_spl_;
  wire g2547_p_spl_;
  wire g3119_p_spl_;
  wire g3119_p_spl_0;
  wire g3121_p_spl_;
  wire g3122_n_spl_;
  wire g3123_n_spl_;
  wire g3120_p_spl_;
  wire g3126_n_spl_;
  wire g3131_p_spl_;
  wire g3131_p_spl_0;
  wire g3131_n_spl_;
  wire g3131_n_spl_0;
  wire g3136_p_spl_;
  wire g3128_n_spl_;
  wire g3093_n_spl_;
  wire g3044_n_spl_;
  wire g3044_n_spl_0;
  wire g3096_n_spl_;
  wire g3047_n_spl_;
  wire g3047_n_spl_0;
  wire g3115_p_spl_;
  wire g3061_p_spl_;
  wire g3099_p_spl_;
  wire g3104_p_spl_;
  wire g3116_n_spl_;
  wire g3060_n_spl_;
  wire g3101_n_spl_;
  wire g3111_n_spl_;
  wire g2947_p_spl_;
  wire g3062_p_spl_;
  wire g2948_p_spl_;
  wire g3063_p_spl_;
  wire g3119_n_spl_;
  wire G126_p_spl_;
  wire G123_p_spl_;
  wire G123_p_spl_0;
  wire G123_p_spl_00;
  wire G123_p_spl_1;
  wire G127_p_spl_;
  wire G123_n_spl_;
  wire G128_p_spl_;
  wire G129_p_spl_;
  wire G124_p_spl_;
  wire G124_p_spl_0;
  wire G124_p_spl_00;
  wire G124_p_spl_01;
  wire G124_p_spl_1;
  wire G105_p_spl_;
  wire G124_n_spl_;
  wire G124_n_spl_0;
  wire G107_p_spl_;
  wire G109_p_spl_;
  wire n4419_lo_n_spl_;
  wire n4419_lo_n_spl_0;
  wire n4431_lo_p_spl_;
  wire n2619_lo_n_spl_;
  wire n2619_lo_n_spl_0;
  wire n2619_lo_n_spl_1;
  wire n3975_lo_n_spl_;
  wire g1207_n_spl_;
  wire n4056_lo_buf_o2_p_spl_;
  wire n2650_inv_p_spl_;
  wire n2650_inv_p_spl_0;
  wire n7396_o2_p_spl_;
  wire n7396_o2_p_spl_0;
  wire n7396_o2_p_spl_1;
  wire n7398_o2_p_spl_;
  wire n7398_o2_p_spl_0;
  wire n7398_o2_p_spl_1;
  wire n7400_o2_p_spl_;
  wire n7400_o2_p_spl_0;
  wire n7400_o2_p_spl_1;
  wire n7402_o2_p_spl_;
  wire n7402_o2_p_spl_0;
  wire n7402_o2_p_spl_1;
  wire n3708_lo_buf_o2_p_spl_;
  wire n4008_lo_buf_o2_p_spl_;
  wire n3732_lo_buf_o2_p_spl_;
  wire n4032_lo_buf_o2_p_spl_;
  wire n3684_lo_buf_o2_p_spl_;
  wire g2592_p_spl_;
  wire g2611_n_spl_;
  wire g2641_n_spl_;
  wire g2660_n_spl_;
  wire g2666_n_spl_;
  wire n3801_lo_p_spl_;
  wire n3813_lo_p_spl_;
  wire g2962_p_spl_;
  wire g2976_p_spl_;
  wire g2995_n_spl_;
  wire g3004_n_spl_;
  wire g3023_p_spl_;
  wire g3032_p_spl_;
  wire n4314_lo_p_spl_;
  wire n4314_lo_p_spl_0;
  wire g3035_n_spl_;
  wire g3035_n_spl_0;
  wire n3777_lo_p_spl_;
  wire n3825_lo_p_spl_;
  wire g3166_n_spl_;
  wire g3169_n_spl_;
  wire g3172_n_spl_;
  wire g3175_n_spl_;
  wire G138_p_spl_;
  wire G139_p_spl_;
  wire G149_p_spl_;
  wire G150_p_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    G37_p,
    G37
  );


  not

  (
    G37_n,
    G37
  );


  buf

  (
    G38_p,
    G38
  );


  not

  (
    G38_n,
    G38
  );


  buf

  (
    G39_p,
    G39
  );


  not

  (
    G39_n,
    G39
  );


  buf

  (
    G40_p,
    G40
  );


  not

  (
    G40_n,
    G40
  );


  buf

  (
    G41_p,
    G41
  );


  not

  (
    G41_n,
    G41
  );


  buf

  (
    G42_p,
    G42
  );


  not

  (
    G42_n,
    G42
  );


  buf

  (
    G43_p,
    G43
  );


  not

  (
    G43_n,
    G43
  );


  buf

  (
    G44_p,
    G44
  );


  not

  (
    G44_n,
    G44
  );


  buf

  (
    G45_p,
    G45
  );


  not

  (
    G45_n,
    G45
  );


  buf

  (
    G46_p,
    G46
  );


  not

  (
    G46_n,
    G46
  );


  buf

  (
    G47_p,
    G47
  );


  not

  (
    G47_n,
    G47
  );


  buf

  (
    G48_p,
    G48
  );


  not

  (
    G48_n,
    G48
  );


  buf

  (
    G49_p,
    G49
  );


  not

  (
    G49_n,
    G49
  );


  buf

  (
    G50_p,
    G50
  );


  not

  (
    G50_n,
    G50
  );


  buf

  (
    G51_p,
    G51
  );


  not

  (
    G51_n,
    G51
  );


  buf

  (
    G52_p,
    G52
  );


  not

  (
    G52_n,
    G52
  );


  buf

  (
    G53_p,
    G53
  );


  not

  (
    G53_n,
    G53
  );


  buf

  (
    G54_p,
    G54
  );


  not

  (
    G54_n,
    G54
  );


  buf

  (
    G55_p,
    G55
  );


  not

  (
    G55_n,
    G55
  );


  buf

  (
    G56_p,
    G56
  );


  not

  (
    G56_n,
    G56
  );


  buf

  (
    G57_p,
    G57
  );


  not

  (
    G57_n,
    G57
  );


  buf

  (
    G58_p,
    G58
  );


  not

  (
    G58_n,
    G58
  );


  buf

  (
    G59_p,
    G59
  );


  not

  (
    G59_n,
    G59
  );


  buf

  (
    G60_p,
    G60
  );


  not

  (
    G60_n,
    G60
  );


  buf

  (
    G61_p,
    G61
  );


  not

  (
    G61_n,
    G61
  );


  buf

  (
    G62_p,
    G62
  );


  not

  (
    G62_n,
    G62
  );


  buf

  (
    G63_p,
    G63
  );


  not

  (
    G63_n,
    G63
  );


  buf

  (
    G64_p,
    G64
  );


  not

  (
    G64_n,
    G64
  );


  buf

  (
    G65_p,
    G65
  );


  not

  (
    G65_n,
    G65
  );


  buf

  (
    G66_p,
    G66
  );


  not

  (
    G66_n,
    G66
  );


  buf

  (
    G67_p,
    G67
  );


  not

  (
    G67_n,
    G67
  );


  buf

  (
    G68_p,
    G68
  );


  not

  (
    G68_n,
    G68
  );


  buf

  (
    G69_p,
    G69
  );


  not

  (
    G69_n,
    G69
  );


  buf

  (
    G70_p,
    G70
  );


  not

  (
    G70_n,
    G70
  );


  buf

  (
    G71_p,
    G71
  );


  not

  (
    G71_n,
    G71
  );


  buf

  (
    G72_p,
    G72
  );


  not

  (
    G72_n,
    G72
  );


  buf

  (
    G73_p,
    G73
  );


  not

  (
    G73_n,
    G73
  );


  buf

  (
    G74_p,
    G74
  );


  not

  (
    G74_n,
    G74
  );


  buf

  (
    G75_p,
    G75
  );


  not

  (
    G75_n,
    G75
  );


  buf

  (
    G76_p,
    G76
  );


  not

  (
    G76_n,
    G76
  );


  buf

  (
    G77_p,
    G77
  );


  not

  (
    G77_n,
    G77
  );


  buf

  (
    G78_p,
    G78
  );


  not

  (
    G78_n,
    G78
  );


  buf

  (
    G79_p,
    G79
  );


  not

  (
    G79_n,
    G79
  );


  buf

  (
    G80_p,
    G80
  );


  not

  (
    G80_n,
    G80
  );


  buf

  (
    G81_p,
    G81
  );


  not

  (
    G81_n,
    G81
  );


  buf

  (
    G82_p,
    G82
  );


  not

  (
    G82_n,
    G82
  );


  buf

  (
    G83_p,
    G83
  );


  not

  (
    G83_n,
    G83
  );


  buf

  (
    G84_p,
    G84
  );


  not

  (
    G84_n,
    G84
  );


  buf

  (
    G85_p,
    G85
  );


  not

  (
    G85_n,
    G85
  );


  buf

  (
    G86_p,
    G86
  );


  not

  (
    G86_n,
    G86
  );


  buf

  (
    G87_p,
    G87
  );


  not

  (
    G87_n,
    G87
  );


  buf

  (
    G88_p,
    G88
  );


  not

  (
    G88_n,
    G88
  );


  buf

  (
    G89_p,
    G89
  );


  not

  (
    G89_n,
    G89
  );


  buf

  (
    G90_p,
    G90
  );


  not

  (
    G90_n,
    G90
  );


  buf

  (
    G91_p,
    G91
  );


  not

  (
    G91_n,
    G91
  );


  buf

  (
    G92_p,
    G92
  );


  not

  (
    G92_n,
    G92
  );


  buf

  (
    G93_p,
    G93
  );


  not

  (
    G93_n,
    G93
  );


  buf

  (
    G94_p,
    G94
  );


  not

  (
    G94_n,
    G94
  );


  buf

  (
    G95_p,
    G95
  );


  not

  (
    G95_n,
    G95
  );


  buf

  (
    G96_p,
    G96
  );


  not

  (
    G96_n,
    G96
  );


  buf

  (
    G97_p,
    G97
  );


  not

  (
    G97_n,
    G97
  );


  buf

  (
    G98_p,
    G98
  );


  not

  (
    G98_n,
    G98
  );


  buf

  (
    G99_p,
    G99
  );


  not

  (
    G99_n,
    G99
  );


  buf

  (
    G100_p,
    G100
  );


  not

  (
    G100_n,
    G100
  );


  buf

  (
    G101_p,
    G101
  );


  not

  (
    G101_n,
    G101
  );


  buf

  (
    G102_p,
    G102
  );


  not

  (
    G102_n,
    G102
  );


  buf

  (
    G103_p,
    G103
  );


  not

  (
    G103_n,
    G103
  );


  buf

  (
    G104_p,
    G104
  );


  not

  (
    G104_n,
    G104
  );


  buf

  (
    G105_p,
    G105
  );


  not

  (
    G105_n,
    G105
  );


  buf

  (
    G106_p,
    G106
  );


  not

  (
    G106_n,
    G106
  );


  buf

  (
    G107_p,
    G107
  );


  not

  (
    G107_n,
    G107
  );


  buf

  (
    G108_p,
    G108
  );


  not

  (
    G108_n,
    G108
  );


  buf

  (
    G109_p,
    G109
  );


  not

  (
    G109_n,
    G109
  );


  buf

  (
    G110_p,
    G110
  );


  not

  (
    G110_n,
    G110
  );


  buf

  (
    G111_p,
    G111
  );


  not

  (
    G111_n,
    G111
  );


  buf

  (
    G112_p,
    G112
  );


  not

  (
    G112_n,
    G112
  );


  buf

  (
    G113_p,
    G113
  );


  not

  (
    G113_n,
    G113
  );


  buf

  (
    G114_p,
    G114
  );


  not

  (
    G114_n,
    G114
  );


  buf

  (
    G115_p,
    G115
  );


  not

  (
    G115_n,
    G115
  );


  buf

  (
    G116_p,
    G116
  );


  not

  (
    G116_n,
    G116
  );


  buf

  (
    G117_p,
    G117
  );


  not

  (
    G117_n,
    G117
  );


  buf

  (
    G118_p,
    G118
  );


  not

  (
    G118_n,
    G118
  );


  buf

  (
    G119_p,
    G119
  );


  not

  (
    G119_n,
    G119
  );


  buf

  (
    G120_p,
    G120
  );


  not

  (
    G120_n,
    G120
  );


  buf

  (
    G121_p,
    G121
  );


  not

  (
    G121_n,
    G121
  );


  buf

  (
    G122_p,
    G122
  );


  not

  (
    G122_n,
    G122
  );


  buf

  (
    G123_p,
    G123
  );


  not

  (
    G123_n,
    G123
  );


  buf

  (
    G124_p,
    G124
  );


  not

  (
    G124_n,
    G124
  );


  buf

  (
    G125_p,
    G125
  );


  not

  (
    G125_n,
    G125
  );


  buf

  (
    G126_p,
    G126
  );


  not

  (
    G126_n,
    G126
  );


  buf

  (
    G127_p,
    G127
  );


  not

  (
    G127_n,
    G127
  );


  buf

  (
    G128_p,
    G128
  );


  not

  (
    G128_n,
    G128
  );


  buf

  (
    G129_p,
    G129
  );


  not

  (
    G129_n,
    G129
  );


  buf

  (
    G130_p,
    G130
  );


  not

  (
    G130_n,
    G130
  );


  buf

  (
    G131_p,
    G131
  );


  not

  (
    G131_n,
    G131
  );


  buf

  (
    G132_p,
    G132
  );


  not

  (
    G132_n,
    G132
  );


  buf

  (
    G133_p,
    G133
  );


  not

  (
    G133_n,
    G133
  );


  buf

  (
    G134_p,
    G134
  );


  not

  (
    G134_n,
    G134
  );


  buf

  (
    G135_p,
    G135
  );


  not

  (
    G135_n,
    G135
  );


  buf

  (
    G136_p,
    G136
  );


  not

  (
    G136_n,
    G136
  );


  buf

  (
    G137_p,
    G137
  );


  not

  (
    G137_n,
    G137
  );


  buf

  (
    G138_p,
    G138
  );


  not

  (
    G138_n,
    G138
  );


  buf

  (
    G139_p,
    G139
  );


  not

  (
    G139_n,
    G139
  );


  buf

  (
    G140_p,
    G140
  );


  not

  (
    G140_n,
    G140
  );


  buf

  (
    G141_p,
    G141
  );


  not

  (
    G141_n,
    G141
  );


  buf

  (
    G142_p,
    G142
  );


  not

  (
    G142_n,
    G142
  );


  buf

  (
    G143_p,
    G143
  );


  not

  (
    G143_n,
    G143
  );


  buf

  (
    G144_p,
    G144
  );


  not

  (
    G144_n,
    G144
  );


  buf

  (
    G145_p,
    G145
  );


  not

  (
    G145_n,
    G145
  );


  buf

  (
    G146_p,
    G146
  );


  not

  (
    G146_n,
    G146
  );


  buf

  (
    G147_p,
    G147
  );


  not

  (
    G147_n,
    G147
  );


  buf

  (
    G148_p,
    G148
  );


  not

  (
    G148_n,
    G148
  );


  buf

  (
    G149_p,
    G149
  );


  not

  (
    G149_n,
    G149
  );


  buf

  (
    G150_p,
    G150
  );


  not

  (
    G150_n,
    G150
  );


  buf

  (
    G151_p,
    G151
  );


  not

  (
    G151_n,
    G151
  );


  buf

  (
    G152_p,
    G152
  );


  not

  (
    G152_n,
    G152
  );


  buf

  (
    G153_p,
    G153
  );


  not

  (
    G153_n,
    G153
  );


  buf

  (
    G154_p,
    G154
  );


  not

  (
    G154_n,
    G154
  );


  buf

  (
    G155_p,
    G155
  );


  not

  (
    G155_n,
    G155
  );


  buf

  (
    G156_p,
    G156
  );


  not

  (
    G156_n,
    G156
  );


  buf

  (
    G157_p,
    G157
  );


  not

  (
    G157_n,
    G157
  );


  buf

  (
    G158_p,
    G158
  );


  not

  (
    G158_n,
    G158
  );


  buf

  (
    G159_p,
    G159
  );


  not

  (
    G159_n,
    G159
  );


  buf

  (
    G160_p,
    G160
  );


  not

  (
    G160_n,
    G160
  );


  buf

  (
    G161_p,
    G161
  );


  not

  (
    G161_n,
    G161
  );


  buf

  (
    G162_p,
    G162
  );


  not

  (
    G162_n,
    G162
  );


  buf

  (
    G163_p,
    G163
  );


  not

  (
    G163_n,
    G163
  );


  buf

  (
    G164_p,
    G164
  );


  not

  (
    G164_n,
    G164
  );


  buf

  (
    G165_p,
    G165
  );


  not

  (
    G165_n,
    G165
  );


  buf

  (
    G166_p,
    G166
  );


  not

  (
    G166_n,
    G166
  );


  buf

  (
    G167_p,
    G167
  );


  not

  (
    G167_n,
    G167
  );


  buf

  (
    G168_p,
    G168
  );


  not

  (
    G168_n,
    G168
  );


  buf

  (
    G169_p,
    G169
  );


  not

  (
    G169_n,
    G169
  );


  buf

  (
    G170_p,
    G170
  );


  not

  (
    G170_n,
    G170
  );


  buf

  (
    G171_p,
    G171
  );


  not

  (
    G171_n,
    G171
  );


  buf

  (
    G172_p,
    G172
  );


  not

  (
    G172_n,
    G172
  );


  buf

  (
    G173_p,
    G173
  );


  not

  (
    G173_n,
    G173
  );


  buf

  (
    G174_p,
    G174
  );


  not

  (
    G174_n,
    G174
  );


  buf

  (
    G175_p,
    G175
  );


  not

  (
    G175_n,
    G175
  );


  buf

  (
    G176_p,
    G176
  );


  not

  (
    G176_n,
    G176
  );


  buf

  (
    G177_p,
    G177
  );


  not

  (
    G177_n,
    G177
  );


  buf

  (
    G178_p,
    G178
  );


  not

  (
    G178_n,
    G178
  );


  buf

  (
    n2610_lo_p,
    n2610_lo
  );


  not

  (
    n2610_lo_n,
    n2610_lo
  );


  buf

  (
    n2613_lo_p,
    n2613_lo
  );


  not

  (
    n2613_lo_n,
    n2613_lo
  );


  buf

  (
    n2616_lo_p,
    n2616_lo
  );


  not

  (
    n2616_lo_n,
    n2616_lo
  );


  buf

  (
    n2619_lo_p,
    n2619_lo
  );


  not

  (
    n2619_lo_n,
    n2619_lo
  );


  buf

  (
    n2622_lo_p,
    n2622_lo
  );


  not

  (
    n2622_lo_n,
    n2622_lo
  );


  buf

  (
    n2625_lo_p,
    n2625_lo
  );


  not

  (
    n2625_lo_n,
    n2625_lo
  );


  buf

  (
    n2628_lo_p,
    n2628_lo
  );


  not

  (
    n2628_lo_n,
    n2628_lo
  );


  buf

  (
    n2631_lo_p,
    n2631_lo
  );


  not

  (
    n2631_lo_n,
    n2631_lo
  );


  buf

  (
    n2634_lo_p,
    n2634_lo
  );


  not

  (
    n2634_lo_n,
    n2634_lo
  );


  buf

  (
    n2637_lo_p,
    n2637_lo
  );


  not

  (
    n2637_lo_n,
    n2637_lo
  );


  buf

  (
    n2640_lo_p,
    n2640_lo
  );


  not

  (
    n2640_lo_n,
    n2640_lo
  );


  buf

  (
    n2643_lo_p,
    n2643_lo
  );


  not

  (
    n2643_lo_n,
    n2643_lo
  );


  buf

  (
    n2646_lo_p,
    n2646_lo
  );


  not

  (
    n2646_lo_n,
    n2646_lo
  );


  buf

  (
    n2649_lo_p,
    n2649_lo
  );


  not

  (
    n2649_lo_n,
    n2649_lo
  );


  buf

  (
    n2652_lo_p,
    n2652_lo
  );


  not

  (
    n2652_lo_n,
    n2652_lo
  );


  buf

  (
    n2655_lo_p,
    n2655_lo
  );


  not

  (
    n2655_lo_n,
    n2655_lo
  );


  buf

  (
    n2658_lo_p,
    n2658_lo
  );


  not

  (
    n2658_lo_n,
    n2658_lo
  );


  buf

  (
    n2661_lo_p,
    n2661_lo
  );


  not

  (
    n2661_lo_n,
    n2661_lo
  );


  buf

  (
    n2664_lo_p,
    n2664_lo
  );


  not

  (
    n2664_lo_n,
    n2664_lo
  );


  buf

  (
    n2667_lo_p,
    n2667_lo
  );


  not

  (
    n2667_lo_n,
    n2667_lo
  );


  buf

  (
    n2670_lo_p,
    n2670_lo
  );


  not

  (
    n2670_lo_n,
    n2670_lo
  );


  buf

  (
    n2673_lo_p,
    n2673_lo
  );


  not

  (
    n2673_lo_n,
    n2673_lo
  );


  buf

  (
    n2676_lo_p,
    n2676_lo
  );


  not

  (
    n2676_lo_n,
    n2676_lo
  );


  buf

  (
    n2679_lo_p,
    n2679_lo
  );


  not

  (
    n2679_lo_n,
    n2679_lo
  );


  buf

  (
    n2682_lo_p,
    n2682_lo
  );


  not

  (
    n2682_lo_n,
    n2682_lo
  );


  buf

  (
    n2685_lo_p,
    n2685_lo
  );


  not

  (
    n2685_lo_n,
    n2685_lo
  );


  buf

  (
    n2688_lo_p,
    n2688_lo
  );


  not

  (
    n2688_lo_n,
    n2688_lo
  );


  buf

  (
    n2691_lo_p,
    n2691_lo
  );


  not

  (
    n2691_lo_n,
    n2691_lo
  );


  buf

  (
    n2694_lo_p,
    n2694_lo
  );


  not

  (
    n2694_lo_n,
    n2694_lo
  );


  buf

  (
    n2697_lo_p,
    n2697_lo
  );


  not

  (
    n2697_lo_n,
    n2697_lo
  );


  buf

  (
    n2700_lo_p,
    n2700_lo
  );


  not

  (
    n2700_lo_n,
    n2700_lo
  );


  buf

  (
    n2703_lo_p,
    n2703_lo
  );


  not

  (
    n2703_lo_n,
    n2703_lo
  );


  buf

  (
    n2706_lo_p,
    n2706_lo
  );


  not

  (
    n2706_lo_n,
    n2706_lo
  );


  buf

  (
    n2709_lo_p,
    n2709_lo
  );


  not

  (
    n2709_lo_n,
    n2709_lo
  );


  buf

  (
    n2712_lo_p,
    n2712_lo
  );


  not

  (
    n2712_lo_n,
    n2712_lo
  );


  buf

  (
    n2715_lo_p,
    n2715_lo
  );


  not

  (
    n2715_lo_n,
    n2715_lo
  );


  buf

  (
    n2718_lo_p,
    n2718_lo
  );


  not

  (
    n2718_lo_n,
    n2718_lo
  );


  buf

  (
    n2721_lo_p,
    n2721_lo
  );


  not

  (
    n2721_lo_n,
    n2721_lo
  );


  buf

  (
    n2724_lo_p,
    n2724_lo
  );


  not

  (
    n2724_lo_n,
    n2724_lo
  );


  buf

  (
    n2727_lo_p,
    n2727_lo
  );


  not

  (
    n2727_lo_n,
    n2727_lo
  );


  buf

  (
    n2730_lo_p,
    n2730_lo
  );


  not

  (
    n2730_lo_n,
    n2730_lo
  );


  buf

  (
    n2733_lo_p,
    n2733_lo
  );


  not

  (
    n2733_lo_n,
    n2733_lo
  );


  buf

  (
    n2736_lo_p,
    n2736_lo
  );


  not

  (
    n2736_lo_n,
    n2736_lo
  );


  buf

  (
    n2739_lo_p,
    n2739_lo
  );


  not

  (
    n2739_lo_n,
    n2739_lo
  );


  buf

  (
    n2742_lo_p,
    n2742_lo
  );


  not

  (
    n2742_lo_n,
    n2742_lo
  );


  buf

  (
    n2745_lo_p,
    n2745_lo
  );


  not

  (
    n2745_lo_n,
    n2745_lo
  );


  buf

  (
    n2748_lo_p,
    n2748_lo
  );


  not

  (
    n2748_lo_n,
    n2748_lo
  );


  buf

  (
    n2751_lo_p,
    n2751_lo
  );


  not

  (
    n2751_lo_n,
    n2751_lo
  );


  buf

  (
    n2754_lo_p,
    n2754_lo
  );


  not

  (
    n2754_lo_n,
    n2754_lo
  );


  buf

  (
    n2757_lo_p,
    n2757_lo
  );


  not

  (
    n2757_lo_n,
    n2757_lo
  );


  buf

  (
    n2760_lo_p,
    n2760_lo
  );


  not

  (
    n2760_lo_n,
    n2760_lo
  );


  buf

  (
    n2763_lo_p,
    n2763_lo
  );


  not

  (
    n2763_lo_n,
    n2763_lo
  );


  buf

  (
    n2766_lo_p,
    n2766_lo
  );


  not

  (
    n2766_lo_n,
    n2766_lo
  );


  buf

  (
    n2769_lo_p,
    n2769_lo
  );


  not

  (
    n2769_lo_n,
    n2769_lo
  );


  buf

  (
    n2772_lo_p,
    n2772_lo
  );


  not

  (
    n2772_lo_n,
    n2772_lo
  );


  buf

  (
    n2775_lo_p,
    n2775_lo
  );


  not

  (
    n2775_lo_n,
    n2775_lo
  );


  buf

  (
    n2778_lo_p,
    n2778_lo
  );


  not

  (
    n2778_lo_n,
    n2778_lo
  );


  buf

  (
    n2781_lo_p,
    n2781_lo
  );


  not

  (
    n2781_lo_n,
    n2781_lo
  );


  buf

  (
    n2784_lo_p,
    n2784_lo
  );


  not

  (
    n2784_lo_n,
    n2784_lo
  );


  buf

  (
    n2787_lo_p,
    n2787_lo
  );


  not

  (
    n2787_lo_n,
    n2787_lo
  );


  buf

  (
    n2790_lo_p,
    n2790_lo
  );


  not

  (
    n2790_lo_n,
    n2790_lo
  );


  buf

  (
    n2793_lo_p,
    n2793_lo
  );


  not

  (
    n2793_lo_n,
    n2793_lo
  );


  buf

  (
    n2796_lo_p,
    n2796_lo
  );


  not

  (
    n2796_lo_n,
    n2796_lo
  );


  buf

  (
    n2799_lo_p,
    n2799_lo
  );


  not

  (
    n2799_lo_n,
    n2799_lo
  );


  buf

  (
    n2802_lo_p,
    n2802_lo
  );


  not

  (
    n2802_lo_n,
    n2802_lo
  );


  buf

  (
    n2805_lo_p,
    n2805_lo
  );


  not

  (
    n2805_lo_n,
    n2805_lo
  );


  buf

  (
    n2808_lo_p,
    n2808_lo
  );


  not

  (
    n2808_lo_n,
    n2808_lo
  );


  buf

  (
    n2811_lo_p,
    n2811_lo
  );


  not

  (
    n2811_lo_n,
    n2811_lo
  );


  buf

  (
    n2814_lo_p,
    n2814_lo
  );


  not

  (
    n2814_lo_n,
    n2814_lo
  );


  buf

  (
    n2817_lo_p,
    n2817_lo
  );


  not

  (
    n2817_lo_n,
    n2817_lo
  );


  buf

  (
    n2820_lo_p,
    n2820_lo
  );


  not

  (
    n2820_lo_n,
    n2820_lo
  );


  buf

  (
    n2823_lo_p,
    n2823_lo
  );


  not

  (
    n2823_lo_n,
    n2823_lo
  );


  buf

  (
    n2826_lo_p,
    n2826_lo
  );


  not

  (
    n2826_lo_n,
    n2826_lo
  );


  buf

  (
    n2829_lo_p,
    n2829_lo
  );


  not

  (
    n2829_lo_n,
    n2829_lo
  );


  buf

  (
    n2832_lo_p,
    n2832_lo
  );


  not

  (
    n2832_lo_n,
    n2832_lo
  );


  buf

  (
    n2835_lo_p,
    n2835_lo
  );


  not

  (
    n2835_lo_n,
    n2835_lo
  );


  buf

  (
    n2838_lo_p,
    n2838_lo
  );


  not

  (
    n2838_lo_n,
    n2838_lo
  );


  buf

  (
    n2841_lo_p,
    n2841_lo
  );


  not

  (
    n2841_lo_n,
    n2841_lo
  );


  buf

  (
    n2844_lo_p,
    n2844_lo
  );


  not

  (
    n2844_lo_n,
    n2844_lo
  );


  buf

  (
    n2847_lo_p,
    n2847_lo
  );


  not

  (
    n2847_lo_n,
    n2847_lo
  );


  buf

  (
    n2850_lo_p,
    n2850_lo
  );


  not

  (
    n2850_lo_n,
    n2850_lo
  );


  buf

  (
    n2853_lo_p,
    n2853_lo
  );


  not

  (
    n2853_lo_n,
    n2853_lo
  );


  buf

  (
    n2856_lo_p,
    n2856_lo
  );


  not

  (
    n2856_lo_n,
    n2856_lo
  );


  buf

  (
    n2859_lo_p,
    n2859_lo
  );


  not

  (
    n2859_lo_n,
    n2859_lo
  );


  buf

  (
    n2862_lo_p,
    n2862_lo
  );


  not

  (
    n2862_lo_n,
    n2862_lo
  );


  buf

  (
    n2865_lo_p,
    n2865_lo
  );


  not

  (
    n2865_lo_n,
    n2865_lo
  );


  buf

  (
    n2868_lo_p,
    n2868_lo
  );


  not

  (
    n2868_lo_n,
    n2868_lo
  );


  buf

  (
    n2871_lo_p,
    n2871_lo
  );


  not

  (
    n2871_lo_n,
    n2871_lo
  );


  buf

  (
    n2874_lo_p,
    n2874_lo
  );


  not

  (
    n2874_lo_n,
    n2874_lo
  );


  buf

  (
    n2877_lo_p,
    n2877_lo
  );


  not

  (
    n2877_lo_n,
    n2877_lo
  );


  buf

  (
    n2880_lo_p,
    n2880_lo
  );


  not

  (
    n2880_lo_n,
    n2880_lo
  );


  buf

  (
    n2883_lo_p,
    n2883_lo
  );


  not

  (
    n2883_lo_n,
    n2883_lo
  );


  buf

  (
    n2886_lo_p,
    n2886_lo
  );


  not

  (
    n2886_lo_n,
    n2886_lo
  );


  buf

  (
    n2889_lo_p,
    n2889_lo
  );


  not

  (
    n2889_lo_n,
    n2889_lo
  );


  buf

  (
    n2892_lo_p,
    n2892_lo
  );


  not

  (
    n2892_lo_n,
    n2892_lo
  );


  buf

  (
    n2895_lo_p,
    n2895_lo
  );


  not

  (
    n2895_lo_n,
    n2895_lo
  );


  buf

  (
    n2898_lo_p,
    n2898_lo
  );


  not

  (
    n2898_lo_n,
    n2898_lo
  );


  buf

  (
    n2901_lo_p,
    n2901_lo
  );


  not

  (
    n2901_lo_n,
    n2901_lo
  );


  buf

  (
    n2904_lo_p,
    n2904_lo
  );


  not

  (
    n2904_lo_n,
    n2904_lo
  );


  buf

  (
    n2907_lo_p,
    n2907_lo
  );


  not

  (
    n2907_lo_n,
    n2907_lo
  );


  buf

  (
    n2910_lo_p,
    n2910_lo
  );


  not

  (
    n2910_lo_n,
    n2910_lo
  );


  buf

  (
    n2913_lo_p,
    n2913_lo
  );


  not

  (
    n2913_lo_n,
    n2913_lo
  );


  buf

  (
    n2916_lo_p,
    n2916_lo
  );


  not

  (
    n2916_lo_n,
    n2916_lo
  );


  buf

  (
    n2919_lo_p,
    n2919_lo
  );


  not

  (
    n2919_lo_n,
    n2919_lo
  );


  buf

  (
    n2922_lo_p,
    n2922_lo
  );


  not

  (
    n2922_lo_n,
    n2922_lo
  );


  buf

  (
    n2925_lo_p,
    n2925_lo
  );


  not

  (
    n2925_lo_n,
    n2925_lo
  );


  buf

  (
    n2928_lo_p,
    n2928_lo
  );


  not

  (
    n2928_lo_n,
    n2928_lo
  );


  buf

  (
    n2931_lo_p,
    n2931_lo
  );


  not

  (
    n2931_lo_n,
    n2931_lo
  );


  buf

  (
    n2934_lo_p,
    n2934_lo
  );


  not

  (
    n2934_lo_n,
    n2934_lo
  );


  buf

  (
    n2937_lo_p,
    n2937_lo
  );


  not

  (
    n2937_lo_n,
    n2937_lo
  );


  buf

  (
    n2940_lo_p,
    n2940_lo
  );


  not

  (
    n2940_lo_n,
    n2940_lo
  );


  buf

  (
    n2943_lo_p,
    n2943_lo
  );


  not

  (
    n2943_lo_n,
    n2943_lo
  );


  buf

  (
    n2946_lo_p,
    n2946_lo
  );


  not

  (
    n2946_lo_n,
    n2946_lo
  );


  buf

  (
    n2949_lo_p,
    n2949_lo
  );


  not

  (
    n2949_lo_n,
    n2949_lo
  );


  buf

  (
    n2952_lo_p,
    n2952_lo
  );


  not

  (
    n2952_lo_n,
    n2952_lo
  );


  buf

  (
    n2955_lo_p,
    n2955_lo
  );


  not

  (
    n2955_lo_n,
    n2955_lo
  );


  buf

  (
    n2958_lo_p,
    n2958_lo
  );


  not

  (
    n2958_lo_n,
    n2958_lo
  );


  buf

  (
    n2961_lo_p,
    n2961_lo
  );


  not

  (
    n2961_lo_n,
    n2961_lo
  );


  buf

  (
    n2964_lo_p,
    n2964_lo
  );


  not

  (
    n2964_lo_n,
    n2964_lo
  );


  buf

  (
    n2967_lo_p,
    n2967_lo
  );


  not

  (
    n2967_lo_n,
    n2967_lo
  );


  buf

  (
    n2970_lo_p,
    n2970_lo
  );


  not

  (
    n2970_lo_n,
    n2970_lo
  );


  buf

  (
    n2973_lo_p,
    n2973_lo
  );


  not

  (
    n2973_lo_n,
    n2973_lo
  );


  buf

  (
    n2976_lo_p,
    n2976_lo
  );


  not

  (
    n2976_lo_n,
    n2976_lo
  );


  buf

  (
    n2979_lo_p,
    n2979_lo
  );


  not

  (
    n2979_lo_n,
    n2979_lo
  );


  buf

  (
    n2982_lo_p,
    n2982_lo
  );


  not

  (
    n2982_lo_n,
    n2982_lo
  );


  buf

  (
    n2985_lo_p,
    n2985_lo
  );


  not

  (
    n2985_lo_n,
    n2985_lo
  );


  buf

  (
    n2988_lo_p,
    n2988_lo
  );


  not

  (
    n2988_lo_n,
    n2988_lo
  );


  buf

  (
    n2991_lo_p,
    n2991_lo
  );


  not

  (
    n2991_lo_n,
    n2991_lo
  );


  buf

  (
    n2994_lo_p,
    n2994_lo
  );


  not

  (
    n2994_lo_n,
    n2994_lo
  );


  buf

  (
    n2997_lo_p,
    n2997_lo
  );


  not

  (
    n2997_lo_n,
    n2997_lo
  );


  buf

  (
    n3000_lo_p,
    n3000_lo
  );


  not

  (
    n3000_lo_n,
    n3000_lo
  );


  buf

  (
    n3003_lo_p,
    n3003_lo
  );


  not

  (
    n3003_lo_n,
    n3003_lo
  );


  buf

  (
    n3006_lo_p,
    n3006_lo
  );


  not

  (
    n3006_lo_n,
    n3006_lo
  );


  buf

  (
    n3009_lo_p,
    n3009_lo
  );


  not

  (
    n3009_lo_n,
    n3009_lo
  );


  buf

  (
    n3012_lo_p,
    n3012_lo
  );


  not

  (
    n3012_lo_n,
    n3012_lo
  );


  buf

  (
    n3015_lo_p,
    n3015_lo
  );


  not

  (
    n3015_lo_n,
    n3015_lo
  );


  buf

  (
    n3018_lo_p,
    n3018_lo
  );


  not

  (
    n3018_lo_n,
    n3018_lo
  );


  buf

  (
    n3021_lo_p,
    n3021_lo
  );


  not

  (
    n3021_lo_n,
    n3021_lo
  );


  buf

  (
    n3024_lo_p,
    n3024_lo
  );


  not

  (
    n3024_lo_n,
    n3024_lo
  );


  buf

  (
    n3027_lo_p,
    n3027_lo
  );


  not

  (
    n3027_lo_n,
    n3027_lo
  );


  buf

  (
    n3030_lo_p,
    n3030_lo
  );


  not

  (
    n3030_lo_n,
    n3030_lo
  );


  buf

  (
    n3033_lo_p,
    n3033_lo
  );


  not

  (
    n3033_lo_n,
    n3033_lo
  );


  buf

  (
    n3036_lo_p,
    n3036_lo
  );


  not

  (
    n3036_lo_n,
    n3036_lo
  );


  buf

  (
    n3039_lo_p,
    n3039_lo
  );


  not

  (
    n3039_lo_n,
    n3039_lo
  );


  buf

  (
    n3042_lo_p,
    n3042_lo
  );


  not

  (
    n3042_lo_n,
    n3042_lo
  );


  buf

  (
    n3045_lo_p,
    n3045_lo
  );


  not

  (
    n3045_lo_n,
    n3045_lo
  );


  buf

  (
    n3048_lo_p,
    n3048_lo
  );


  not

  (
    n3048_lo_n,
    n3048_lo
  );


  buf

  (
    n3051_lo_p,
    n3051_lo
  );


  not

  (
    n3051_lo_n,
    n3051_lo
  );


  buf

  (
    n3054_lo_p,
    n3054_lo
  );


  not

  (
    n3054_lo_n,
    n3054_lo
  );


  buf

  (
    n3057_lo_p,
    n3057_lo
  );


  not

  (
    n3057_lo_n,
    n3057_lo
  );


  buf

  (
    n3060_lo_p,
    n3060_lo
  );


  not

  (
    n3060_lo_n,
    n3060_lo
  );


  buf

  (
    n3063_lo_p,
    n3063_lo
  );


  not

  (
    n3063_lo_n,
    n3063_lo
  );


  buf

  (
    n3066_lo_p,
    n3066_lo
  );


  not

  (
    n3066_lo_n,
    n3066_lo
  );


  buf

  (
    n3069_lo_p,
    n3069_lo
  );


  not

  (
    n3069_lo_n,
    n3069_lo
  );


  buf

  (
    n3072_lo_p,
    n3072_lo
  );


  not

  (
    n3072_lo_n,
    n3072_lo
  );


  buf

  (
    n3075_lo_p,
    n3075_lo
  );


  not

  (
    n3075_lo_n,
    n3075_lo
  );


  buf

  (
    n3078_lo_p,
    n3078_lo
  );


  not

  (
    n3078_lo_n,
    n3078_lo
  );


  buf

  (
    n3081_lo_p,
    n3081_lo
  );


  not

  (
    n3081_lo_n,
    n3081_lo
  );


  buf

  (
    n3084_lo_p,
    n3084_lo
  );


  not

  (
    n3084_lo_n,
    n3084_lo
  );


  buf

  (
    n3087_lo_p,
    n3087_lo
  );


  not

  (
    n3087_lo_n,
    n3087_lo
  );


  buf

  (
    n3090_lo_p,
    n3090_lo
  );


  not

  (
    n3090_lo_n,
    n3090_lo
  );


  buf

  (
    n3093_lo_p,
    n3093_lo
  );


  not

  (
    n3093_lo_n,
    n3093_lo
  );


  buf

  (
    n3096_lo_p,
    n3096_lo
  );


  not

  (
    n3096_lo_n,
    n3096_lo
  );


  buf

  (
    n3099_lo_p,
    n3099_lo
  );


  not

  (
    n3099_lo_n,
    n3099_lo
  );


  buf

  (
    n3102_lo_p,
    n3102_lo
  );


  not

  (
    n3102_lo_n,
    n3102_lo
  );


  buf

  (
    n3105_lo_p,
    n3105_lo
  );


  not

  (
    n3105_lo_n,
    n3105_lo
  );


  buf

  (
    n3108_lo_p,
    n3108_lo
  );


  not

  (
    n3108_lo_n,
    n3108_lo
  );


  buf

  (
    n3111_lo_p,
    n3111_lo
  );


  not

  (
    n3111_lo_n,
    n3111_lo
  );


  buf

  (
    n3114_lo_p,
    n3114_lo
  );


  not

  (
    n3114_lo_n,
    n3114_lo
  );


  buf

  (
    n3117_lo_p,
    n3117_lo
  );


  not

  (
    n3117_lo_n,
    n3117_lo
  );


  buf

  (
    n3120_lo_p,
    n3120_lo
  );


  not

  (
    n3120_lo_n,
    n3120_lo
  );


  buf

  (
    n3123_lo_p,
    n3123_lo
  );


  not

  (
    n3123_lo_n,
    n3123_lo
  );


  buf

  (
    n3126_lo_p,
    n3126_lo
  );


  not

  (
    n3126_lo_n,
    n3126_lo
  );


  buf

  (
    n3129_lo_p,
    n3129_lo
  );


  not

  (
    n3129_lo_n,
    n3129_lo
  );


  buf

  (
    n3132_lo_p,
    n3132_lo
  );


  not

  (
    n3132_lo_n,
    n3132_lo
  );


  buf

  (
    n3135_lo_p,
    n3135_lo
  );


  not

  (
    n3135_lo_n,
    n3135_lo
  );


  buf

  (
    n3138_lo_p,
    n3138_lo
  );


  not

  (
    n3138_lo_n,
    n3138_lo
  );


  buf

  (
    n3141_lo_p,
    n3141_lo
  );


  not

  (
    n3141_lo_n,
    n3141_lo
  );


  buf

  (
    n3144_lo_p,
    n3144_lo
  );


  not

  (
    n3144_lo_n,
    n3144_lo
  );


  buf

  (
    n3147_lo_p,
    n3147_lo
  );


  not

  (
    n3147_lo_n,
    n3147_lo
  );


  buf

  (
    n3150_lo_p,
    n3150_lo
  );


  not

  (
    n3150_lo_n,
    n3150_lo
  );


  buf

  (
    n3153_lo_p,
    n3153_lo
  );


  not

  (
    n3153_lo_n,
    n3153_lo
  );


  buf

  (
    n3156_lo_p,
    n3156_lo
  );


  not

  (
    n3156_lo_n,
    n3156_lo
  );


  buf

  (
    n3159_lo_p,
    n3159_lo
  );


  not

  (
    n3159_lo_n,
    n3159_lo
  );


  buf

  (
    n3162_lo_p,
    n3162_lo
  );


  not

  (
    n3162_lo_n,
    n3162_lo
  );


  buf

  (
    n3165_lo_p,
    n3165_lo
  );


  not

  (
    n3165_lo_n,
    n3165_lo
  );


  buf

  (
    n3168_lo_p,
    n3168_lo
  );


  not

  (
    n3168_lo_n,
    n3168_lo
  );


  buf

  (
    n3171_lo_p,
    n3171_lo
  );


  not

  (
    n3171_lo_n,
    n3171_lo
  );


  buf

  (
    n3174_lo_p,
    n3174_lo
  );


  not

  (
    n3174_lo_n,
    n3174_lo
  );


  buf

  (
    n3177_lo_p,
    n3177_lo
  );


  not

  (
    n3177_lo_n,
    n3177_lo
  );


  buf

  (
    n3180_lo_p,
    n3180_lo
  );


  not

  (
    n3180_lo_n,
    n3180_lo
  );


  buf

  (
    n3183_lo_p,
    n3183_lo
  );


  not

  (
    n3183_lo_n,
    n3183_lo
  );


  buf

  (
    n3186_lo_p,
    n3186_lo
  );


  not

  (
    n3186_lo_n,
    n3186_lo
  );


  buf

  (
    n3189_lo_p,
    n3189_lo
  );


  not

  (
    n3189_lo_n,
    n3189_lo
  );


  buf

  (
    n3192_lo_p,
    n3192_lo
  );


  not

  (
    n3192_lo_n,
    n3192_lo
  );


  buf

  (
    n3195_lo_p,
    n3195_lo
  );


  not

  (
    n3195_lo_n,
    n3195_lo
  );


  buf

  (
    n3198_lo_p,
    n3198_lo
  );


  not

  (
    n3198_lo_n,
    n3198_lo
  );


  buf

  (
    n3201_lo_p,
    n3201_lo
  );


  not

  (
    n3201_lo_n,
    n3201_lo
  );


  buf

  (
    n3204_lo_p,
    n3204_lo
  );


  not

  (
    n3204_lo_n,
    n3204_lo
  );


  buf

  (
    n3207_lo_p,
    n3207_lo
  );


  not

  (
    n3207_lo_n,
    n3207_lo
  );


  buf

  (
    n3210_lo_p,
    n3210_lo
  );


  not

  (
    n3210_lo_n,
    n3210_lo
  );


  buf

  (
    n3213_lo_p,
    n3213_lo
  );


  not

  (
    n3213_lo_n,
    n3213_lo
  );


  buf

  (
    n3216_lo_p,
    n3216_lo
  );


  not

  (
    n3216_lo_n,
    n3216_lo
  );


  buf

  (
    n3219_lo_p,
    n3219_lo
  );


  not

  (
    n3219_lo_n,
    n3219_lo
  );


  buf

  (
    n3222_lo_p,
    n3222_lo
  );


  not

  (
    n3222_lo_n,
    n3222_lo
  );


  buf

  (
    n3225_lo_p,
    n3225_lo
  );


  not

  (
    n3225_lo_n,
    n3225_lo
  );


  buf

  (
    n3228_lo_p,
    n3228_lo
  );


  not

  (
    n3228_lo_n,
    n3228_lo
  );


  buf

  (
    n3231_lo_p,
    n3231_lo
  );


  not

  (
    n3231_lo_n,
    n3231_lo
  );


  buf

  (
    n3234_lo_p,
    n3234_lo
  );


  not

  (
    n3234_lo_n,
    n3234_lo
  );


  buf

  (
    n3237_lo_p,
    n3237_lo
  );


  not

  (
    n3237_lo_n,
    n3237_lo
  );


  buf

  (
    n3240_lo_p,
    n3240_lo
  );


  not

  (
    n3240_lo_n,
    n3240_lo
  );


  buf

  (
    n3243_lo_p,
    n3243_lo
  );


  not

  (
    n3243_lo_n,
    n3243_lo
  );


  buf

  (
    n3246_lo_p,
    n3246_lo
  );


  not

  (
    n3246_lo_n,
    n3246_lo
  );


  buf

  (
    n3249_lo_p,
    n3249_lo
  );


  not

  (
    n3249_lo_n,
    n3249_lo
  );


  buf

  (
    n3252_lo_p,
    n3252_lo
  );


  not

  (
    n3252_lo_n,
    n3252_lo
  );


  buf

  (
    n3255_lo_p,
    n3255_lo
  );


  not

  (
    n3255_lo_n,
    n3255_lo
  );


  buf

  (
    n3258_lo_p,
    n3258_lo
  );


  not

  (
    n3258_lo_n,
    n3258_lo
  );


  buf

  (
    n3261_lo_p,
    n3261_lo
  );


  not

  (
    n3261_lo_n,
    n3261_lo
  );


  buf

  (
    n3264_lo_p,
    n3264_lo
  );


  not

  (
    n3264_lo_n,
    n3264_lo
  );


  buf

  (
    n3267_lo_p,
    n3267_lo
  );


  not

  (
    n3267_lo_n,
    n3267_lo
  );


  buf

  (
    n3270_lo_p,
    n3270_lo
  );


  not

  (
    n3270_lo_n,
    n3270_lo
  );


  buf

  (
    n3273_lo_p,
    n3273_lo
  );


  not

  (
    n3273_lo_n,
    n3273_lo
  );


  buf

  (
    n3276_lo_p,
    n3276_lo
  );


  not

  (
    n3276_lo_n,
    n3276_lo
  );


  buf

  (
    n3279_lo_p,
    n3279_lo
  );


  not

  (
    n3279_lo_n,
    n3279_lo
  );


  buf

  (
    n3282_lo_p,
    n3282_lo
  );


  not

  (
    n3282_lo_n,
    n3282_lo
  );


  buf

  (
    n3285_lo_p,
    n3285_lo
  );


  not

  (
    n3285_lo_n,
    n3285_lo
  );


  buf

  (
    n3288_lo_p,
    n3288_lo
  );


  not

  (
    n3288_lo_n,
    n3288_lo
  );


  buf

  (
    n3291_lo_p,
    n3291_lo
  );


  not

  (
    n3291_lo_n,
    n3291_lo
  );


  buf

  (
    n3294_lo_p,
    n3294_lo
  );


  not

  (
    n3294_lo_n,
    n3294_lo
  );


  buf

  (
    n3297_lo_p,
    n3297_lo
  );


  not

  (
    n3297_lo_n,
    n3297_lo
  );


  buf

  (
    n3300_lo_p,
    n3300_lo
  );


  not

  (
    n3300_lo_n,
    n3300_lo
  );


  buf

  (
    n3303_lo_p,
    n3303_lo
  );


  not

  (
    n3303_lo_n,
    n3303_lo
  );


  buf

  (
    n3306_lo_p,
    n3306_lo
  );


  not

  (
    n3306_lo_n,
    n3306_lo
  );


  buf

  (
    n3309_lo_p,
    n3309_lo
  );


  not

  (
    n3309_lo_n,
    n3309_lo
  );


  buf

  (
    n3312_lo_p,
    n3312_lo
  );


  not

  (
    n3312_lo_n,
    n3312_lo
  );


  buf

  (
    n3315_lo_p,
    n3315_lo
  );


  not

  (
    n3315_lo_n,
    n3315_lo
  );


  buf

  (
    n3318_lo_p,
    n3318_lo
  );


  not

  (
    n3318_lo_n,
    n3318_lo
  );


  buf

  (
    n3321_lo_p,
    n3321_lo
  );


  not

  (
    n3321_lo_n,
    n3321_lo
  );


  buf

  (
    n3324_lo_p,
    n3324_lo
  );


  not

  (
    n3324_lo_n,
    n3324_lo
  );


  buf

  (
    n3327_lo_p,
    n3327_lo
  );


  not

  (
    n3327_lo_n,
    n3327_lo
  );


  buf

  (
    n3330_lo_p,
    n3330_lo
  );


  not

  (
    n3330_lo_n,
    n3330_lo
  );


  buf

  (
    n3333_lo_p,
    n3333_lo
  );


  not

  (
    n3333_lo_n,
    n3333_lo
  );


  buf

  (
    n3336_lo_p,
    n3336_lo
  );


  not

  (
    n3336_lo_n,
    n3336_lo
  );


  buf

  (
    n3339_lo_p,
    n3339_lo
  );


  not

  (
    n3339_lo_n,
    n3339_lo
  );


  buf

  (
    n3342_lo_p,
    n3342_lo
  );


  not

  (
    n3342_lo_n,
    n3342_lo
  );


  buf

  (
    n3345_lo_p,
    n3345_lo
  );


  not

  (
    n3345_lo_n,
    n3345_lo
  );


  buf

  (
    n3348_lo_p,
    n3348_lo
  );


  not

  (
    n3348_lo_n,
    n3348_lo
  );


  buf

  (
    n3351_lo_p,
    n3351_lo
  );


  not

  (
    n3351_lo_n,
    n3351_lo
  );


  buf

  (
    n3354_lo_p,
    n3354_lo
  );


  not

  (
    n3354_lo_n,
    n3354_lo
  );


  buf

  (
    n3357_lo_p,
    n3357_lo
  );


  not

  (
    n3357_lo_n,
    n3357_lo
  );


  buf

  (
    n3360_lo_p,
    n3360_lo
  );


  not

  (
    n3360_lo_n,
    n3360_lo
  );


  buf

  (
    n3363_lo_p,
    n3363_lo
  );


  not

  (
    n3363_lo_n,
    n3363_lo
  );


  buf

  (
    n3366_lo_p,
    n3366_lo
  );


  not

  (
    n3366_lo_n,
    n3366_lo
  );


  buf

  (
    n3369_lo_p,
    n3369_lo
  );


  not

  (
    n3369_lo_n,
    n3369_lo
  );


  buf

  (
    n3372_lo_p,
    n3372_lo
  );


  not

  (
    n3372_lo_n,
    n3372_lo
  );


  buf

  (
    n3375_lo_p,
    n3375_lo
  );


  not

  (
    n3375_lo_n,
    n3375_lo
  );


  buf

  (
    n3378_lo_p,
    n3378_lo
  );


  not

  (
    n3378_lo_n,
    n3378_lo
  );


  buf

  (
    n3381_lo_p,
    n3381_lo
  );


  not

  (
    n3381_lo_n,
    n3381_lo
  );


  buf

  (
    n3384_lo_p,
    n3384_lo
  );


  not

  (
    n3384_lo_n,
    n3384_lo
  );


  buf

  (
    n3387_lo_p,
    n3387_lo
  );


  not

  (
    n3387_lo_n,
    n3387_lo
  );


  buf

  (
    n3390_lo_p,
    n3390_lo
  );


  not

  (
    n3390_lo_n,
    n3390_lo
  );


  buf

  (
    n3393_lo_p,
    n3393_lo
  );


  not

  (
    n3393_lo_n,
    n3393_lo
  );


  buf

  (
    n3396_lo_p,
    n3396_lo
  );


  not

  (
    n3396_lo_n,
    n3396_lo
  );


  buf

  (
    n3399_lo_p,
    n3399_lo
  );


  not

  (
    n3399_lo_n,
    n3399_lo
  );


  buf

  (
    n3402_lo_p,
    n3402_lo
  );


  not

  (
    n3402_lo_n,
    n3402_lo
  );


  buf

  (
    n3405_lo_p,
    n3405_lo
  );


  not

  (
    n3405_lo_n,
    n3405_lo
  );


  buf

  (
    n3408_lo_p,
    n3408_lo
  );


  not

  (
    n3408_lo_n,
    n3408_lo
  );


  buf

  (
    n3411_lo_p,
    n3411_lo
  );


  not

  (
    n3411_lo_n,
    n3411_lo
  );


  buf

  (
    n3414_lo_p,
    n3414_lo
  );


  not

  (
    n3414_lo_n,
    n3414_lo
  );


  buf

  (
    n3417_lo_p,
    n3417_lo
  );


  not

  (
    n3417_lo_n,
    n3417_lo
  );


  buf

  (
    n3420_lo_p,
    n3420_lo
  );


  not

  (
    n3420_lo_n,
    n3420_lo
  );


  buf

  (
    n3423_lo_p,
    n3423_lo
  );


  not

  (
    n3423_lo_n,
    n3423_lo
  );


  buf

  (
    n3426_lo_p,
    n3426_lo
  );


  not

  (
    n3426_lo_n,
    n3426_lo
  );


  buf

  (
    n3429_lo_p,
    n3429_lo
  );


  not

  (
    n3429_lo_n,
    n3429_lo
  );


  buf

  (
    n3432_lo_p,
    n3432_lo
  );


  not

  (
    n3432_lo_n,
    n3432_lo
  );


  buf

  (
    n3435_lo_p,
    n3435_lo
  );


  not

  (
    n3435_lo_n,
    n3435_lo
  );


  buf

  (
    n3438_lo_p,
    n3438_lo
  );


  not

  (
    n3438_lo_n,
    n3438_lo
  );


  buf

  (
    n3441_lo_p,
    n3441_lo
  );


  not

  (
    n3441_lo_n,
    n3441_lo
  );


  buf

  (
    n3444_lo_p,
    n3444_lo
  );


  not

  (
    n3444_lo_n,
    n3444_lo
  );


  buf

  (
    n3447_lo_p,
    n3447_lo
  );


  not

  (
    n3447_lo_n,
    n3447_lo
  );


  buf

  (
    n3450_lo_p,
    n3450_lo
  );


  not

  (
    n3450_lo_n,
    n3450_lo
  );


  buf

  (
    n3453_lo_p,
    n3453_lo
  );


  not

  (
    n3453_lo_n,
    n3453_lo
  );


  buf

  (
    n3456_lo_p,
    n3456_lo
  );


  not

  (
    n3456_lo_n,
    n3456_lo
  );


  buf

  (
    n3459_lo_p,
    n3459_lo
  );


  not

  (
    n3459_lo_n,
    n3459_lo
  );


  buf

  (
    n3462_lo_p,
    n3462_lo
  );


  not

  (
    n3462_lo_n,
    n3462_lo
  );


  buf

  (
    n3465_lo_p,
    n3465_lo
  );


  not

  (
    n3465_lo_n,
    n3465_lo
  );


  buf

  (
    n3468_lo_p,
    n3468_lo
  );


  not

  (
    n3468_lo_n,
    n3468_lo
  );


  buf

  (
    n3471_lo_p,
    n3471_lo
  );


  not

  (
    n3471_lo_n,
    n3471_lo
  );


  buf

  (
    n3474_lo_p,
    n3474_lo
  );


  not

  (
    n3474_lo_n,
    n3474_lo
  );


  buf

  (
    n3477_lo_p,
    n3477_lo
  );


  not

  (
    n3477_lo_n,
    n3477_lo
  );


  buf

  (
    n3480_lo_p,
    n3480_lo
  );


  not

  (
    n3480_lo_n,
    n3480_lo
  );


  buf

  (
    n3483_lo_p,
    n3483_lo
  );


  not

  (
    n3483_lo_n,
    n3483_lo
  );


  buf

  (
    n3486_lo_p,
    n3486_lo
  );


  not

  (
    n3486_lo_n,
    n3486_lo
  );


  buf

  (
    n3489_lo_p,
    n3489_lo
  );


  not

  (
    n3489_lo_n,
    n3489_lo
  );


  buf

  (
    n3492_lo_p,
    n3492_lo
  );


  not

  (
    n3492_lo_n,
    n3492_lo
  );


  buf

  (
    n3495_lo_p,
    n3495_lo
  );


  not

  (
    n3495_lo_n,
    n3495_lo
  );


  buf

  (
    n3498_lo_p,
    n3498_lo
  );


  not

  (
    n3498_lo_n,
    n3498_lo
  );


  buf

  (
    n3501_lo_p,
    n3501_lo
  );


  not

  (
    n3501_lo_n,
    n3501_lo
  );


  buf

  (
    n3504_lo_p,
    n3504_lo
  );


  not

  (
    n3504_lo_n,
    n3504_lo
  );


  buf

  (
    n3507_lo_p,
    n3507_lo
  );


  not

  (
    n3507_lo_n,
    n3507_lo
  );


  buf

  (
    n3510_lo_p,
    n3510_lo
  );


  not

  (
    n3510_lo_n,
    n3510_lo
  );


  buf

  (
    n3513_lo_p,
    n3513_lo
  );


  not

  (
    n3513_lo_n,
    n3513_lo
  );


  buf

  (
    n3516_lo_p,
    n3516_lo
  );


  not

  (
    n3516_lo_n,
    n3516_lo
  );


  buf

  (
    n3519_lo_p,
    n3519_lo
  );


  not

  (
    n3519_lo_n,
    n3519_lo
  );


  buf

  (
    n3522_lo_p,
    n3522_lo
  );


  not

  (
    n3522_lo_n,
    n3522_lo
  );


  buf

  (
    n3525_lo_p,
    n3525_lo
  );


  not

  (
    n3525_lo_n,
    n3525_lo
  );


  buf

  (
    n3528_lo_p,
    n3528_lo
  );


  not

  (
    n3528_lo_n,
    n3528_lo
  );


  buf

  (
    n3531_lo_p,
    n3531_lo
  );


  not

  (
    n3531_lo_n,
    n3531_lo
  );


  buf

  (
    n3534_lo_p,
    n3534_lo
  );


  not

  (
    n3534_lo_n,
    n3534_lo
  );


  buf

  (
    n3537_lo_p,
    n3537_lo
  );


  not

  (
    n3537_lo_n,
    n3537_lo
  );


  buf

  (
    n3540_lo_p,
    n3540_lo
  );


  not

  (
    n3540_lo_n,
    n3540_lo
  );


  buf

  (
    n3543_lo_p,
    n3543_lo
  );


  not

  (
    n3543_lo_n,
    n3543_lo
  );


  buf

  (
    n3546_lo_p,
    n3546_lo
  );


  not

  (
    n3546_lo_n,
    n3546_lo
  );


  buf

  (
    n3549_lo_p,
    n3549_lo
  );


  not

  (
    n3549_lo_n,
    n3549_lo
  );


  buf

  (
    n3552_lo_p,
    n3552_lo
  );


  not

  (
    n3552_lo_n,
    n3552_lo
  );


  buf

  (
    n3555_lo_p,
    n3555_lo
  );


  not

  (
    n3555_lo_n,
    n3555_lo
  );


  buf

  (
    n3558_lo_p,
    n3558_lo
  );


  not

  (
    n3558_lo_n,
    n3558_lo
  );


  buf

  (
    n3561_lo_p,
    n3561_lo
  );


  not

  (
    n3561_lo_n,
    n3561_lo
  );


  buf

  (
    n3564_lo_p,
    n3564_lo
  );


  not

  (
    n3564_lo_n,
    n3564_lo
  );


  buf

  (
    n3567_lo_p,
    n3567_lo
  );


  not

  (
    n3567_lo_n,
    n3567_lo
  );


  buf

  (
    n3570_lo_p,
    n3570_lo
  );


  not

  (
    n3570_lo_n,
    n3570_lo
  );


  buf

  (
    n3573_lo_p,
    n3573_lo
  );


  not

  (
    n3573_lo_n,
    n3573_lo
  );


  buf

  (
    n3576_lo_p,
    n3576_lo
  );


  not

  (
    n3576_lo_n,
    n3576_lo
  );


  buf

  (
    n3579_lo_p,
    n3579_lo
  );


  not

  (
    n3579_lo_n,
    n3579_lo
  );


  buf

  (
    n3582_lo_p,
    n3582_lo
  );


  not

  (
    n3582_lo_n,
    n3582_lo
  );


  buf

  (
    n3585_lo_p,
    n3585_lo
  );


  not

  (
    n3585_lo_n,
    n3585_lo
  );


  buf

  (
    n3588_lo_p,
    n3588_lo
  );


  not

  (
    n3588_lo_n,
    n3588_lo
  );


  buf

  (
    n3591_lo_p,
    n3591_lo
  );


  not

  (
    n3591_lo_n,
    n3591_lo
  );


  buf

  (
    n3594_lo_p,
    n3594_lo
  );


  not

  (
    n3594_lo_n,
    n3594_lo
  );


  buf

  (
    n3597_lo_p,
    n3597_lo
  );


  not

  (
    n3597_lo_n,
    n3597_lo
  );


  buf

  (
    n3600_lo_p,
    n3600_lo
  );


  not

  (
    n3600_lo_n,
    n3600_lo
  );


  buf

  (
    n3603_lo_p,
    n3603_lo
  );


  not

  (
    n3603_lo_n,
    n3603_lo
  );


  buf

  (
    n3606_lo_p,
    n3606_lo
  );


  not

  (
    n3606_lo_n,
    n3606_lo
  );


  buf

  (
    n3609_lo_p,
    n3609_lo
  );


  not

  (
    n3609_lo_n,
    n3609_lo
  );


  buf

  (
    n3612_lo_p,
    n3612_lo
  );


  not

  (
    n3612_lo_n,
    n3612_lo
  );


  buf

  (
    n3615_lo_p,
    n3615_lo
  );


  not

  (
    n3615_lo_n,
    n3615_lo
  );


  buf

  (
    n3618_lo_p,
    n3618_lo
  );


  not

  (
    n3618_lo_n,
    n3618_lo
  );


  buf

  (
    n3621_lo_p,
    n3621_lo
  );


  not

  (
    n3621_lo_n,
    n3621_lo
  );


  buf

  (
    n3624_lo_p,
    n3624_lo
  );


  not

  (
    n3624_lo_n,
    n3624_lo
  );


  buf

  (
    n3627_lo_p,
    n3627_lo
  );


  not

  (
    n3627_lo_n,
    n3627_lo
  );


  buf

  (
    n3630_lo_p,
    n3630_lo
  );


  not

  (
    n3630_lo_n,
    n3630_lo
  );


  buf

  (
    n3633_lo_p,
    n3633_lo
  );


  not

  (
    n3633_lo_n,
    n3633_lo
  );


  buf

  (
    n3636_lo_p,
    n3636_lo
  );


  not

  (
    n3636_lo_n,
    n3636_lo
  );


  buf

  (
    n3639_lo_p,
    n3639_lo
  );


  not

  (
    n3639_lo_n,
    n3639_lo
  );


  buf

  (
    n3642_lo_p,
    n3642_lo
  );


  not

  (
    n3642_lo_n,
    n3642_lo
  );


  buf

  (
    n3645_lo_p,
    n3645_lo
  );


  not

  (
    n3645_lo_n,
    n3645_lo
  );


  buf

  (
    n3648_lo_p,
    n3648_lo
  );


  not

  (
    n3648_lo_n,
    n3648_lo
  );


  buf

  (
    n3651_lo_p,
    n3651_lo
  );


  not

  (
    n3651_lo_n,
    n3651_lo
  );


  buf

  (
    n3654_lo_p,
    n3654_lo
  );


  not

  (
    n3654_lo_n,
    n3654_lo
  );


  buf

  (
    n3657_lo_p,
    n3657_lo
  );


  not

  (
    n3657_lo_n,
    n3657_lo
  );


  buf

  (
    n3666_lo_p,
    n3666_lo
  );


  not

  (
    n3666_lo_n,
    n3666_lo
  );


  buf

  (
    n3669_lo_p,
    n3669_lo
  );


  not

  (
    n3669_lo_n,
    n3669_lo
  );


  buf

  (
    n3678_lo_p,
    n3678_lo
  );


  not

  (
    n3678_lo_n,
    n3678_lo
  );


  buf

  (
    n3687_lo_p,
    n3687_lo
  );


  not

  (
    n3687_lo_n,
    n3687_lo
  );


  buf

  (
    n3690_lo_p,
    n3690_lo
  );


  not

  (
    n3690_lo_n,
    n3690_lo
  );


  buf

  (
    n3702_lo_p,
    n3702_lo
  );


  not

  (
    n3702_lo_n,
    n3702_lo
  );


  buf

  (
    n3711_lo_p,
    n3711_lo
  );


  not

  (
    n3711_lo_n,
    n3711_lo
  );


  buf

  (
    n3714_lo_p,
    n3714_lo
  );


  not

  (
    n3714_lo_n,
    n3714_lo
  );


  buf

  (
    n3726_lo_p,
    n3726_lo
  );


  not

  (
    n3726_lo_n,
    n3726_lo
  );


  buf

  (
    n3735_lo_p,
    n3735_lo
  );


  not

  (
    n3735_lo_n,
    n3735_lo
  );


  buf

  (
    n3738_lo_p,
    n3738_lo
  );


  not

  (
    n3738_lo_n,
    n3738_lo
  );


  buf

  (
    n3750_lo_p,
    n3750_lo
  );


  not

  (
    n3750_lo_n,
    n3750_lo
  );


  buf

  (
    n3753_lo_p,
    n3753_lo
  );


  not

  (
    n3753_lo_n,
    n3753_lo
  );


  buf

  (
    n3759_lo_p,
    n3759_lo
  );


  not

  (
    n3759_lo_n,
    n3759_lo
  );


  buf

  (
    n3762_lo_p,
    n3762_lo
  );


  not

  (
    n3762_lo_n,
    n3762_lo
  );


  buf

  (
    n3765_lo_p,
    n3765_lo
  );


  not

  (
    n3765_lo_n,
    n3765_lo
  );


  buf

  (
    n3774_lo_p,
    n3774_lo
  );


  not

  (
    n3774_lo_n,
    n3774_lo
  );


  buf

  (
    n3777_lo_p,
    n3777_lo
  );


  not

  (
    n3777_lo_n,
    n3777_lo
  );


  buf

  (
    n3786_lo_p,
    n3786_lo
  );


  not

  (
    n3786_lo_n,
    n3786_lo
  );


  buf

  (
    n3789_lo_p,
    n3789_lo
  );


  not

  (
    n3789_lo_n,
    n3789_lo
  );


  buf

  (
    n3792_lo_p,
    n3792_lo
  );


  not

  (
    n3792_lo_n,
    n3792_lo
  );


  buf

  (
    n3795_lo_p,
    n3795_lo
  );


  not

  (
    n3795_lo_n,
    n3795_lo
  );


  buf

  (
    n3798_lo_p,
    n3798_lo
  );


  not

  (
    n3798_lo_n,
    n3798_lo
  );


  buf

  (
    n3801_lo_p,
    n3801_lo
  );


  not

  (
    n3801_lo_n,
    n3801_lo
  );


  buf

  (
    n3810_lo_p,
    n3810_lo
  );


  not

  (
    n3810_lo_n,
    n3810_lo
  );


  buf

  (
    n3813_lo_p,
    n3813_lo
  );


  not

  (
    n3813_lo_n,
    n3813_lo
  );


  buf

  (
    n3822_lo_p,
    n3822_lo
  );


  not

  (
    n3822_lo_n,
    n3822_lo
  );


  buf

  (
    n3825_lo_p,
    n3825_lo
  );


  not

  (
    n3825_lo_n,
    n3825_lo
  );


  buf

  (
    n3834_lo_p,
    n3834_lo
  );


  not

  (
    n3834_lo_n,
    n3834_lo
  );


  buf

  (
    n3843_lo_p,
    n3843_lo
  );


  not

  (
    n3843_lo_n,
    n3843_lo
  );


  buf

  (
    n3846_lo_p,
    n3846_lo
  );


  not

  (
    n3846_lo_n,
    n3846_lo
  );


  buf

  (
    n3867_lo_p,
    n3867_lo
  );


  not

  (
    n3867_lo_n,
    n3867_lo
  );


  buf

  (
    n3891_lo_p,
    n3891_lo
  );


  not

  (
    n3891_lo_n,
    n3891_lo
  );


  buf

  (
    n3915_lo_p,
    n3915_lo
  );


  not

  (
    n3915_lo_n,
    n3915_lo
  );


  buf

  (
    n3930_lo_p,
    n3930_lo
  );


  not

  (
    n3930_lo_n,
    n3930_lo
  );


  buf

  (
    n3933_lo_p,
    n3933_lo
  );


  not

  (
    n3933_lo_n,
    n3933_lo
  );


  buf

  (
    n3936_lo_p,
    n3936_lo
  );


  not

  (
    n3936_lo_n,
    n3936_lo
  );


  buf

  (
    n3942_lo_p,
    n3942_lo
  );


  not

  (
    n3942_lo_n,
    n3942_lo
  );


  buf

  (
    n3945_lo_p,
    n3945_lo
  );


  not

  (
    n3945_lo_n,
    n3945_lo
  );


  buf

  (
    n3948_lo_p,
    n3948_lo
  );


  not

  (
    n3948_lo_n,
    n3948_lo
  );


  buf

  (
    n3954_lo_p,
    n3954_lo
  );


  not

  (
    n3954_lo_n,
    n3954_lo
  );


  buf

  (
    n3957_lo_p,
    n3957_lo
  );


  not

  (
    n3957_lo_n,
    n3957_lo
  );


  buf

  (
    n3963_lo_p,
    n3963_lo
  );


  not

  (
    n3963_lo_n,
    n3963_lo
  );


  buf

  (
    n3966_lo_p,
    n3966_lo
  );


  not

  (
    n3966_lo_n,
    n3966_lo
  );


  buf

  (
    n3969_lo_p,
    n3969_lo
  );


  not

  (
    n3969_lo_n,
    n3969_lo
  );


  buf

  (
    n3975_lo_p,
    n3975_lo
  );


  not

  (
    n3975_lo_n,
    n3975_lo
  );


  buf

  (
    n3978_lo_p,
    n3978_lo
  );


  not

  (
    n3978_lo_n,
    n3978_lo
  );


  buf

  (
    n3987_lo_p,
    n3987_lo
  );


  not

  (
    n3987_lo_n,
    n3987_lo
  );


  buf

  (
    n3990_lo_p,
    n3990_lo
  );


  not

  (
    n3990_lo_n,
    n3990_lo
  );


  buf

  (
    n4002_lo_p,
    n4002_lo
  );


  not

  (
    n4002_lo_n,
    n4002_lo
  );


  buf

  (
    n4011_lo_p,
    n4011_lo
  );


  not

  (
    n4011_lo_n,
    n4011_lo
  );


  buf

  (
    n4014_lo_p,
    n4014_lo
  );


  not

  (
    n4014_lo_n,
    n4014_lo
  );


  buf

  (
    n4026_lo_p,
    n4026_lo
  );


  not

  (
    n4026_lo_n,
    n4026_lo
  );


  buf

  (
    n4035_lo_p,
    n4035_lo
  );


  not

  (
    n4035_lo_n,
    n4035_lo
  );


  buf

  (
    n4038_lo_p,
    n4038_lo
  );


  not

  (
    n4038_lo_n,
    n4038_lo
  );


  buf

  (
    n4050_lo_p,
    n4050_lo
  );


  not

  (
    n4050_lo_n,
    n4050_lo
  );


  buf

  (
    n4053_lo_p,
    n4053_lo
  );


  not

  (
    n4053_lo_n,
    n4053_lo
  );


  buf

  (
    n4059_lo_p,
    n4059_lo
  );


  not

  (
    n4059_lo_n,
    n4059_lo
  );


  buf

  (
    n4062_lo_p,
    n4062_lo
  );


  not

  (
    n4062_lo_n,
    n4062_lo
  );


  buf

  (
    n4065_lo_p,
    n4065_lo
  );


  not

  (
    n4065_lo_n,
    n4065_lo
  );


  buf

  (
    n4098_lo_p,
    n4098_lo
  );


  not

  (
    n4098_lo_n,
    n4098_lo
  );


  buf

  (
    n4107_lo_p,
    n4107_lo
  );


  not

  (
    n4107_lo_n,
    n4107_lo
  );


  buf

  (
    n4119_lo_p,
    n4119_lo
  );


  not

  (
    n4119_lo_n,
    n4119_lo
  );


  buf

  (
    n4131_lo_p,
    n4131_lo
  );


  not

  (
    n4131_lo_n,
    n4131_lo
  );


  buf

  (
    n4143_lo_p,
    n4143_lo
  );


  not

  (
    n4143_lo_n,
    n4143_lo
  );


  buf

  (
    n4155_lo_p,
    n4155_lo
  );


  not

  (
    n4155_lo_n,
    n4155_lo
  );


  buf

  (
    n4167_lo_p,
    n4167_lo
  );


  not

  (
    n4167_lo_n,
    n4167_lo
  );


  buf

  (
    n4179_lo_p,
    n4179_lo
  );


  not

  (
    n4179_lo_n,
    n4179_lo
  );


  buf

  (
    n4182_lo_p,
    n4182_lo
  );


  not

  (
    n4182_lo_n,
    n4182_lo
  );


  buf

  (
    n4185_lo_p,
    n4185_lo
  );


  not

  (
    n4185_lo_n,
    n4185_lo
  );


  buf

  (
    n4188_lo_p,
    n4188_lo
  );


  not

  (
    n4188_lo_n,
    n4188_lo
  );


  buf

  (
    n4194_lo_p,
    n4194_lo
  );


  not

  (
    n4194_lo_n,
    n4194_lo
  );


  buf

  (
    n4197_lo_p,
    n4197_lo
  );


  not

  (
    n4197_lo_n,
    n4197_lo
  );


  buf

  (
    n4200_lo_p,
    n4200_lo
  );


  not

  (
    n4200_lo_n,
    n4200_lo
  );


  buf

  (
    n4206_lo_p,
    n4206_lo
  );


  not

  (
    n4206_lo_n,
    n4206_lo
  );


  buf

  (
    n4209_lo_p,
    n4209_lo
  );


  not

  (
    n4209_lo_n,
    n4209_lo
  );


  buf

  (
    n4212_lo_p,
    n4212_lo
  );


  not

  (
    n4212_lo_n,
    n4212_lo
  );


  buf

  (
    n4215_lo_p,
    n4215_lo
  );


  not

  (
    n4215_lo_n,
    n4215_lo
  );


  buf

  (
    n4227_lo_p,
    n4227_lo
  );


  not

  (
    n4227_lo_n,
    n4227_lo
  );


  buf

  (
    n4230_lo_p,
    n4230_lo
  );


  not

  (
    n4230_lo_n,
    n4230_lo
  );


  buf

  (
    n4233_lo_p,
    n4233_lo
  );


  not

  (
    n4233_lo_n,
    n4233_lo
  );


  buf

  (
    n4236_lo_p,
    n4236_lo
  );


  not

  (
    n4236_lo_n,
    n4236_lo
  );


  buf

  (
    n4239_lo_p,
    n4239_lo
  );


  not

  (
    n4239_lo_n,
    n4239_lo
  );


  buf

  (
    n4242_lo_p,
    n4242_lo
  );


  not

  (
    n4242_lo_n,
    n4242_lo
  );


  buf

  (
    n4251_lo_p,
    n4251_lo
  );


  not

  (
    n4251_lo_n,
    n4251_lo
  );


  buf

  (
    n4263_lo_p,
    n4263_lo
  );


  not

  (
    n4263_lo_n,
    n4263_lo
  );


  buf

  (
    n4275_lo_p,
    n4275_lo
  );


  not

  (
    n4275_lo_n,
    n4275_lo
  );


  buf

  (
    n4278_lo_p,
    n4278_lo
  );


  not

  (
    n4278_lo_n,
    n4278_lo
  );


  buf

  (
    n4287_lo_p,
    n4287_lo
  );


  not

  (
    n4287_lo_n,
    n4287_lo
  );


  buf

  (
    n4290_lo_p,
    n4290_lo
  );


  not

  (
    n4290_lo_n,
    n4290_lo
  );


  buf

  (
    n4293_lo_p,
    n4293_lo
  );


  not

  (
    n4293_lo_n,
    n4293_lo
  );


  buf

  (
    n4299_lo_p,
    n4299_lo
  );


  not

  (
    n4299_lo_n,
    n4299_lo
  );


  buf

  (
    n4302_lo_p,
    n4302_lo
  );


  not

  (
    n4302_lo_n,
    n4302_lo
  );


  buf

  (
    n4305_lo_p,
    n4305_lo
  );


  not

  (
    n4305_lo_n,
    n4305_lo
  );


  buf

  (
    n4311_lo_p,
    n4311_lo
  );


  not

  (
    n4311_lo_n,
    n4311_lo
  );


  buf

  (
    n4314_lo_p,
    n4314_lo
  );


  not

  (
    n4314_lo_n,
    n4314_lo
  );


  buf

  (
    n4323_lo_p,
    n4323_lo
  );


  not

  (
    n4323_lo_n,
    n4323_lo
  );


  buf

  (
    n4326_lo_p,
    n4326_lo
  );


  not

  (
    n4326_lo_n,
    n4326_lo
  );


  buf

  (
    n4335_lo_p,
    n4335_lo
  );


  not

  (
    n4335_lo_n,
    n4335_lo
  );


  buf

  (
    n4338_lo_p,
    n4338_lo
  );


  not

  (
    n4338_lo_n,
    n4338_lo
  );


  buf

  (
    n4347_lo_p,
    n4347_lo
  );


  not

  (
    n4347_lo_n,
    n4347_lo
  );


  buf

  (
    n4350_lo_p,
    n4350_lo
  );


  not

  (
    n4350_lo_n,
    n4350_lo
  );


  buf

  (
    n4359_lo_p,
    n4359_lo
  );


  not

  (
    n4359_lo_n,
    n4359_lo
  );


  buf

  (
    n4362_lo_p,
    n4362_lo
  );


  not

  (
    n4362_lo_n,
    n4362_lo
  );


  buf

  (
    n4365_lo_p,
    n4365_lo
  );


  not

  (
    n4365_lo_n,
    n4365_lo
  );


  buf

  (
    n4371_lo_p,
    n4371_lo
  );


  not

  (
    n4371_lo_n,
    n4371_lo
  );


  buf

  (
    n4374_lo_p,
    n4374_lo
  );


  not

  (
    n4374_lo_n,
    n4374_lo
  );


  buf

  (
    n4383_lo_p,
    n4383_lo
  );


  not

  (
    n4383_lo_n,
    n4383_lo
  );


  buf

  (
    n4395_lo_p,
    n4395_lo
  );


  not

  (
    n4395_lo_n,
    n4395_lo
  );


  buf

  (
    n4407_lo_p,
    n4407_lo
  );


  not

  (
    n4407_lo_n,
    n4407_lo
  );


  buf

  (
    n4410_lo_p,
    n4410_lo
  );


  not

  (
    n4410_lo_n,
    n4410_lo
  );


  buf

  (
    n4413_lo_p,
    n4413_lo
  );


  not

  (
    n4413_lo_n,
    n4413_lo
  );


  buf

  (
    n4416_lo_p,
    n4416_lo
  );


  not

  (
    n4416_lo_n,
    n4416_lo
  );


  buf

  (
    n4419_lo_p,
    n4419_lo
  );


  not

  (
    n4419_lo_n,
    n4419_lo
  );


  buf

  (
    n4422_lo_p,
    n4422_lo
  );


  not

  (
    n4422_lo_n,
    n4422_lo
  );


  buf

  (
    n4425_lo_p,
    n4425_lo
  );


  not

  (
    n4425_lo_n,
    n4425_lo
  );


  buf

  (
    n4428_lo_p,
    n4428_lo
  );


  not

  (
    n4428_lo_n,
    n4428_lo
  );


  buf

  (
    n4431_lo_p,
    n4431_lo
  );


  not

  (
    n4431_lo_n,
    n4431_lo
  );


  buf

  (
    n4434_lo_p,
    n4434_lo
  );


  not

  (
    n4434_lo_n,
    n4434_lo
  );


  buf

  (
    n4437_lo_p,
    n4437_lo
  );


  not

  (
    n4437_lo_n,
    n4437_lo
  );


  buf

  (
    n4440_lo_p,
    n4440_lo
  );


  not

  (
    n4440_lo_n,
    n4440_lo
  );


  buf

  (
    n4443_lo_p,
    n4443_lo
  );


  not

  (
    n4443_lo_n,
    n4443_lo
  );


  buf

  (
    n4446_lo_p,
    n4446_lo
  );


  not

  (
    n4446_lo_n,
    n4446_lo
  );


  buf

  (
    n4449_lo_p,
    n4449_lo
  );


  not

  (
    n4449_lo_n,
    n4449_lo
  );


  buf

  (
    n4452_lo_p,
    n4452_lo
  );


  not

  (
    n4452_lo_n,
    n4452_lo
  );


  buf

  (
    n4455_lo_p,
    n4455_lo
  );


  not

  (
    n4455_lo_n,
    n4455_lo
  );


  buf

  (
    n4458_lo_p,
    n4458_lo
  );


  not

  (
    n4458_lo_n,
    n4458_lo
  );


  buf

  (
    n4461_lo_p,
    n4461_lo
  );


  not

  (
    n4461_lo_n,
    n4461_lo
  );


  buf

  (
    n4464_lo_p,
    n4464_lo
  );


  not

  (
    n4464_lo_n,
    n4464_lo
  );


  buf

  (
    n4467_lo_p,
    n4467_lo
  );


  not

  (
    n4467_lo_n,
    n4467_lo
  );


  buf

  (
    n4470_lo_p,
    n4470_lo
  );


  not

  (
    n4470_lo_n,
    n4470_lo
  );


  buf

  (
    n4473_lo_p,
    n4473_lo
  );


  not

  (
    n4473_lo_n,
    n4473_lo
  );


  buf

  (
    n4476_lo_p,
    n4476_lo
  );


  not

  (
    n4476_lo_n,
    n4476_lo
  );


  buf

  (
    n4479_lo_p,
    n4479_lo
  );


  not

  (
    n4479_lo_n,
    n4479_lo
  );


  buf

  (
    n4482_lo_p,
    n4482_lo
  );


  not

  (
    n4482_lo_n,
    n4482_lo
  );


  buf

  (
    n4485_lo_p,
    n4485_lo
  );


  not

  (
    n4485_lo_n,
    n4485_lo
  );


  buf

  (
    n4488_lo_p,
    n4488_lo
  );


  not

  (
    n4488_lo_n,
    n4488_lo
  );


  buf

  (
    n4494_lo_p,
    n4494_lo
  );


  not

  (
    n4494_lo_n,
    n4494_lo
  );


  buf

  (
    n4497_lo_p,
    n4497_lo
  );


  not

  (
    n4497_lo_n,
    n4497_lo
  );


  buf

  (
    n4500_lo_p,
    n4500_lo
  );


  not

  (
    n4500_lo_n,
    n4500_lo
  );


  buf

  (
    n4503_lo_p,
    n4503_lo
  );


  not

  (
    n4503_lo_n,
    n4503_lo
  );


  buf

  (
    n4506_lo_p,
    n4506_lo
  );


  not

  (
    n4506_lo_n,
    n4506_lo
  );


  buf

  (
    n4509_lo_p,
    n4509_lo
  );


  not

  (
    n4509_lo_n,
    n4509_lo
  );


  buf

  (
    n4512_lo_p,
    n4512_lo
  );


  not

  (
    n4512_lo_n,
    n4512_lo
  );


  buf

  (
    n4515_lo_p,
    n4515_lo
  );


  not

  (
    n4515_lo_n,
    n4515_lo
  );


  buf

  (
    n4518_lo_p,
    n4518_lo
  );


  not

  (
    n4518_lo_n,
    n4518_lo
  );


  buf

  (
    n4521_lo_p,
    n4521_lo
  );


  not

  (
    n4521_lo_n,
    n4521_lo
  );


  buf

  (
    n4524_lo_p,
    n4524_lo
  );


  not

  (
    n4524_lo_n,
    n4524_lo
  );


  buf

  (
    n4527_lo_p,
    n4527_lo
  );


  not

  (
    n4527_lo_n,
    n4527_lo
  );


  buf

  (
    n4530_lo_p,
    n4530_lo
  );


  not

  (
    n4530_lo_n,
    n4530_lo
  );


  buf

  (
    n4533_lo_p,
    n4533_lo
  );


  not

  (
    n4533_lo_n,
    n4533_lo
  );


  buf

  (
    n4536_lo_p,
    n4536_lo
  );


  not

  (
    n4536_lo_n,
    n4536_lo
  );


  buf

  (
    n4539_lo_p,
    n4539_lo
  );


  not

  (
    n4539_lo_n,
    n4539_lo
  );


  buf

  (
    n4542_lo_p,
    n4542_lo
  );


  not

  (
    n4542_lo_n,
    n4542_lo
  );


  buf

  (
    n4545_lo_p,
    n4545_lo
  );


  not

  (
    n4545_lo_n,
    n4545_lo
  );


  buf

  (
    n4548_lo_p,
    n4548_lo
  );


  not

  (
    n4548_lo_n,
    n4548_lo
  );


  buf

  (
    n4554_lo_p,
    n4554_lo
  );


  not

  (
    n4554_lo_n,
    n4554_lo
  );


  buf

  (
    n4557_lo_p,
    n4557_lo
  );


  not

  (
    n4557_lo_n,
    n4557_lo
  );


  buf

  (
    n4560_lo_p,
    n4560_lo
  );


  not

  (
    n4560_lo_n,
    n4560_lo
  );


  buf

  (
    n4563_lo_p,
    n4563_lo
  );


  not

  (
    n4563_lo_n,
    n4563_lo
  );


  buf

  (
    n4566_lo_p,
    n4566_lo
  );


  not

  (
    n4566_lo_n,
    n4566_lo
  );


  buf

  (
    n4569_lo_p,
    n4569_lo
  );


  not

  (
    n4569_lo_n,
    n4569_lo
  );


  buf

  (
    n4572_lo_p,
    n4572_lo
  );


  not

  (
    n4572_lo_n,
    n4572_lo
  );


  buf

  (
    n4575_lo_p,
    n4575_lo
  );


  not

  (
    n4575_lo_n,
    n4575_lo
  );


  buf

  (
    n4578_lo_p,
    n4578_lo
  );


  not

  (
    n4578_lo_n,
    n4578_lo
  );


  buf

  (
    n4581_lo_p,
    n4581_lo
  );


  not

  (
    n4581_lo_n,
    n4581_lo
  );


  buf

  (
    n4584_lo_p,
    n4584_lo
  );


  not

  (
    n4584_lo_n,
    n4584_lo
  );


  buf

  (
    n4587_lo_p,
    n4587_lo
  );


  not

  (
    n4587_lo_n,
    n4587_lo
  );


  buf

  (
    n4590_lo_p,
    n4590_lo
  );


  not

  (
    n4590_lo_n,
    n4590_lo
  );


  buf

  (
    n4593_lo_p,
    n4593_lo
  );


  not

  (
    n4593_lo_n,
    n4593_lo
  );


  buf

  (
    n4596_lo_p,
    n4596_lo
  );


  not

  (
    n4596_lo_n,
    n4596_lo
  );


  buf

  (
    n4599_lo_p,
    n4599_lo
  );


  not

  (
    n4599_lo_n,
    n4599_lo
  );


  buf

  (
    n4602_lo_p,
    n4602_lo
  );


  not

  (
    n4602_lo_n,
    n4602_lo
  );


  buf

  (
    n4605_lo_p,
    n4605_lo
  );


  not

  (
    n4605_lo_n,
    n4605_lo
  );


  buf

  (
    n4608_lo_p,
    n4608_lo
  );


  not

  (
    n4608_lo_n,
    n4608_lo
  );


  buf

  (
    n4611_lo_p,
    n4611_lo
  );


  not

  (
    n4611_lo_n,
    n4611_lo
  );


  buf

  (
    n4614_lo_p,
    n4614_lo
  );


  not

  (
    n4614_lo_n,
    n4614_lo
  );


  buf

  (
    n4617_lo_p,
    n4617_lo
  );


  not

  (
    n4617_lo_n,
    n4617_lo
  );


  buf

  (
    n4620_lo_p,
    n4620_lo
  );


  not

  (
    n4620_lo_n,
    n4620_lo
  );


  buf

  (
    n4623_lo_p,
    n4623_lo
  );


  not

  (
    n4623_lo_n,
    n4623_lo
  );


  buf

  (
    n4626_lo_p,
    n4626_lo
  );


  not

  (
    n4626_lo_n,
    n4626_lo
  );


  buf

  (
    n4629_lo_p,
    n4629_lo
  );


  not

  (
    n4629_lo_n,
    n4629_lo
  );


  buf

  (
    n4632_lo_p,
    n4632_lo
  );


  not

  (
    n4632_lo_n,
    n4632_lo
  );


  buf

  (
    n4635_lo_p,
    n4635_lo
  );


  not

  (
    n4635_lo_n,
    n4635_lo
  );


  buf

  (
    n4638_lo_p,
    n4638_lo
  );


  not

  (
    n4638_lo_n,
    n4638_lo
  );


  buf

  (
    n4641_lo_p,
    n4641_lo
  );


  not

  (
    n4641_lo_n,
    n4641_lo
  );


  buf

  (
    n4644_lo_p,
    n4644_lo
  );


  not

  (
    n4644_lo_n,
    n4644_lo
  );


  buf

  (
    n4647_lo_p,
    n4647_lo
  );


  not

  (
    n4647_lo_n,
    n4647_lo
  );


  buf

  (
    n4650_lo_p,
    n4650_lo
  );


  not

  (
    n4650_lo_n,
    n4650_lo
  );


  buf

  (
    n4653_lo_p,
    n4653_lo
  );


  not

  (
    n4653_lo_n,
    n4653_lo
  );


  buf

  (
    n4656_lo_p,
    n4656_lo
  );


  not

  (
    n4656_lo_n,
    n4656_lo
  );


  buf

  (
    n4659_lo_p,
    n4659_lo
  );


  not

  (
    n4659_lo_n,
    n4659_lo
  );


  buf

  (
    n4662_lo_p,
    n4662_lo
  );


  not

  (
    n4662_lo_n,
    n4662_lo
  );


  buf

  (
    n4665_lo_p,
    n4665_lo
  );


  not

  (
    n4665_lo_n,
    n4665_lo
  );


  buf

  (
    n4668_lo_p,
    n4668_lo
  );


  not

  (
    n4668_lo_n,
    n4668_lo
  );


  buf

  (
    n4671_lo_p,
    n4671_lo
  );


  not

  (
    n4671_lo_n,
    n4671_lo
  );


  buf

  (
    n4674_lo_p,
    n4674_lo
  );


  not

  (
    n4674_lo_n,
    n4674_lo
  );


  buf

  (
    n4677_lo_p,
    n4677_lo
  );


  not

  (
    n4677_lo_n,
    n4677_lo
  );


  buf

  (
    n4680_lo_p,
    n4680_lo
  );


  not

  (
    n4680_lo_n,
    n4680_lo
  );


  buf

  (
    n4683_lo_p,
    n4683_lo
  );


  not

  (
    n4683_lo_n,
    n4683_lo
  );


  buf

  (
    n4686_lo_p,
    n4686_lo
  );


  not

  (
    n4686_lo_n,
    n4686_lo
  );


  buf

  (
    n4689_lo_p,
    n4689_lo
  );


  not

  (
    n4689_lo_n,
    n4689_lo
  );


  buf

  (
    n4692_lo_p,
    n4692_lo
  );


  not

  (
    n4692_lo_n,
    n4692_lo
  );


  buf

  (
    n4695_lo_p,
    n4695_lo
  );


  not

  (
    n4695_lo_n,
    n4695_lo
  );


  buf

  (
    n4698_lo_p,
    n4698_lo
  );


  not

  (
    n4698_lo_n,
    n4698_lo
  );


  buf

  (
    n4701_lo_p,
    n4701_lo
  );


  not

  (
    n4701_lo_n,
    n4701_lo
  );


  buf

  (
    n4704_lo_p,
    n4704_lo
  );


  not

  (
    n4704_lo_n,
    n4704_lo
  );


  buf

  (
    n4707_lo_p,
    n4707_lo
  );


  not

  (
    n4707_lo_n,
    n4707_lo
  );


  buf

  (
    n4710_lo_p,
    n4710_lo
  );


  not

  (
    n4710_lo_n,
    n4710_lo
  );


  buf

  (
    n4713_lo_p,
    n4713_lo
  );


  not

  (
    n4713_lo_n,
    n4713_lo
  );


  buf

  (
    n4716_lo_p,
    n4716_lo
  );


  not

  (
    n4716_lo_n,
    n4716_lo
  );


  buf

  (
    n4719_lo_p,
    n4719_lo
  );


  not

  (
    n4719_lo_n,
    n4719_lo
  );


  buf

  (
    n4722_lo_p,
    n4722_lo
  );


  not

  (
    n4722_lo_n,
    n4722_lo
  );


  buf

  (
    n4725_lo_p,
    n4725_lo
  );


  not

  (
    n4725_lo_n,
    n4725_lo
  );


  buf

  (
    n4728_lo_p,
    n4728_lo
  );


  not

  (
    n4728_lo_n,
    n4728_lo
  );


  buf

  (
    n4731_lo_p,
    n4731_lo
  );


  not

  (
    n4731_lo_n,
    n4731_lo
  );


  buf

  (
    n4734_lo_p,
    n4734_lo
  );


  not

  (
    n4734_lo_n,
    n4734_lo
  );


  buf

  (
    n4737_lo_p,
    n4737_lo
  );


  not

  (
    n4737_lo_n,
    n4737_lo
  );


  buf

  (
    n4740_lo_p,
    n4740_lo
  );


  not

  (
    n4740_lo_n,
    n4740_lo
  );


  buf

  (
    n4743_lo_p,
    n4743_lo
  );


  not

  (
    n4743_lo_n,
    n4743_lo
  );


  buf

  (
    n6382_o2_p,
    n6382_o2
  );


  not

  (
    n6382_o2_n,
    n6382_o2
  );


  buf

  (
    n6383_o2_p,
    n6383_o2
  );


  not

  (
    n6383_o2_n,
    n6383_o2
  );


  buf

  (
    n6419_o2_p,
    n6419_o2
  );


  not

  (
    n6419_o2_n,
    n6419_o2
  );


  buf

  (
    n6420_o2_p,
    n6420_o2
  );


  not

  (
    n6420_o2_n,
    n6420_o2
  );


  buf

  (
    n6435_o2_p,
    n6435_o2
  );


  not

  (
    n6435_o2_n,
    n6435_o2
  );


  buf

  (
    n6436_o2_p,
    n6436_o2
  );


  not

  (
    n6436_o2_n,
    n6436_o2
  );


  buf

  (
    n6448_o2_p,
    n6448_o2
  );


  not

  (
    n6448_o2_n,
    n6448_o2
  );


  buf

  (
    n6449_o2_p,
    n6449_o2
  );


  not

  (
    n6449_o2_n,
    n6449_o2
  );


  buf

  (
    n6613_o2_p,
    n6613_o2
  );


  not

  (
    n6613_o2_n,
    n6613_o2
  );


  buf

  (
    n6614_o2_p,
    n6614_o2
  );


  not

  (
    n6614_o2_n,
    n6614_o2
  );


  buf

  (
    n6641_o2_p,
    n6641_o2
  );


  not

  (
    n6641_o2_n,
    n6641_o2
  );


  buf

  (
    n6658_o2_p,
    n6658_o2
  );


  not

  (
    n6658_o2_n,
    n6658_o2
  );


  buf

  (
    n6757_o2_p,
    n6757_o2
  );


  not

  (
    n6757_o2_n,
    n6757_o2
  );


  buf

  (
    n6756_o2_p,
    n6756_o2
  );


  not

  (
    n6756_o2_n,
    n6756_o2
  );


  buf

  (
    n7116_o2_p,
    n7116_o2
  );


  not

  (
    n7116_o2_n,
    n7116_o2
  );


  buf

  (
    n7156_o2_p,
    n7156_o2
  );


  not

  (
    n7156_o2_n,
    n7156_o2
  );


  buf

  (
    n6549_o2_p,
    n6549_o2
  );


  not

  (
    n6549_o2_n,
    n6549_o2
  );


  buf

  (
    n6550_o2_p,
    n6550_o2
  );


  not

  (
    n6550_o2_n,
    n6550_o2
  );


  buf

  (
    n7357_o2_p,
    n7357_o2
  );


  not

  (
    n7357_o2_n,
    n7357_o2
  );


  buf

  (
    n7358_o2_p,
    n7358_o2
  );


  not

  (
    n7358_o2_n,
    n7358_o2
  );


  buf

  (
    n7359_o2_p,
    n7359_o2
  );


  not

  (
    n7359_o2_n,
    n7359_o2
  );


  buf

  (
    n7360_o2_p,
    n7360_o2
  );


  not

  (
    n7360_o2_n,
    n7360_o2
  );


  buf

  (
    n6621_o2_p,
    n6621_o2
  );


  not

  (
    n6621_o2_n,
    n6621_o2
  );


  buf

  (
    n6623_o2_p,
    n6623_o2
  );


  not

  (
    n6623_o2_n,
    n6623_o2
  );


  buf

  (
    n6625_o2_p,
    n6625_o2
  );


  not

  (
    n6625_o2_n,
    n6625_o2
  );


  buf

  (
    n6626_o2_p,
    n6626_o2
  );


  not

  (
    n6626_o2_n,
    n6626_o2
  );


  buf

  (
    n6627_o2_p,
    n6627_o2
  );


  not

  (
    n6627_o2_n,
    n6627_o2
  );


  buf

  (
    n6628_o2_p,
    n6628_o2
  );


  not

  (
    n6628_o2_n,
    n6628_o2
  );


  buf

  (
    n6629_o2_p,
    n6629_o2
  );


  not

  (
    n6629_o2_n,
    n6629_o2
  );


  buf

  (
    n6630_o2_p,
    n6630_o2
  );


  not

  (
    n6630_o2_n,
    n6630_o2
  );


  buf

  (
    n6669_o2_p,
    n6669_o2
  );


  not

  (
    n6669_o2_n,
    n6669_o2
  );


  buf

  (
    n7449_o2_p,
    n7449_o2
  );


  not

  (
    n7449_o2_n,
    n7449_o2
  );


  buf

  (
    n7450_o2_p,
    n7450_o2
  );


  not

  (
    n7450_o2_n,
    n7450_o2
  );


  buf

  (
    n7451_o2_p,
    n7451_o2
  );


  not

  (
    n7451_o2_n,
    n7451_o2
  );


  buf

  (
    n7452_o2_p,
    n7452_o2
  );


  not

  (
    n7452_o2_n,
    n7452_o2
  );


  buf

  (
    n6682_o2_p,
    n6682_o2
  );


  not

  (
    n6682_o2_n,
    n6682_o2
  );


  buf

  (
    n6683_o2_p,
    n6683_o2
  );


  not

  (
    n6683_o2_n,
    n6683_o2
  );


  buf

  (
    n6684_o2_p,
    n6684_o2
  );


  not

  (
    n6684_o2_n,
    n6684_o2
  );


  buf

  (
    n6685_o2_p,
    n6685_o2
  );


  not

  (
    n6685_o2_n,
    n6685_o2
  );


  buf

  (
    n7463_o2_p,
    n7463_o2
  );


  not

  (
    n7463_o2_n,
    n7463_o2
  );


  buf

  (
    n6686_o2_p,
    n6686_o2
  );


  not

  (
    n6686_o2_n,
    n6686_o2
  );


  buf

  (
    n6687_o2_p,
    n6687_o2
  );


  not

  (
    n6687_o2_n,
    n6687_o2
  );


  buf

  (
    n6688_o2_p,
    n6688_o2
  );


  not

  (
    n6688_o2_n,
    n6688_o2
  );


  buf

  (
    n6689_o2_p,
    n6689_o2
  );


  not

  (
    n6689_o2_n,
    n6689_o2
  );


  buf

  (
    n6772_o2_p,
    n6772_o2
  );


  not

  (
    n6772_o2_n,
    n6772_o2
  );


  buf

  (
    n6773_o2_p,
    n6773_o2
  );


  not

  (
    n6773_o2_n,
    n6773_o2
  );


  buf

  (
    n6774_o2_p,
    n6774_o2
  );


  not

  (
    n6774_o2_n,
    n6774_o2
  );


  buf

  (
    n6775_o2_p,
    n6775_o2
  );


  not

  (
    n6775_o2_n,
    n6775_o2
  );


  buf

  (
    G3467_o2_p,
    G3467_o2
  );


  not

  (
    G3467_o2_n,
    G3467_o2
  );


  buf

  (
    G2810_o2_p,
    G2810_o2
  );


  not

  (
    G2810_o2_n,
    G2810_o2
  );


  buf

  (
    n6833_o2_p,
    n6833_o2
  );


  not

  (
    n6833_o2_n,
    n6833_o2
  );


  buf

  (
    n6945_o2_p,
    n6945_o2
  );


  not

  (
    n6945_o2_n,
    n6945_o2
  );


  buf

  (
    n6947_o2_p,
    n6947_o2
  );


  not

  (
    n6947_o2_n,
    n6947_o2
  );


  buf

  (
    n6949_o2_p,
    n6949_o2
  );


  not

  (
    n6949_o2_n,
    n6949_o2
  );


  buf

  (
    n6951_o2_p,
    n6951_o2
  );


  not

  (
    n6951_o2_n,
    n6951_o2
  );


  buf

  (
    n6888_o2_p,
    n6888_o2
  );


  not

  (
    n6888_o2_n,
    n6888_o2
  );


  buf

  (
    n6889_o2_p,
    n6889_o2
  );


  not

  (
    n6889_o2_n,
    n6889_o2
  );


  buf

  (
    n6936_o2_p,
    n6936_o2
  );


  not

  (
    n6936_o2_n,
    n6936_o2
  );


  buf

  (
    n6954_o2_p,
    n6954_o2
  );


  not

  (
    n6954_o2_n,
    n6954_o2
  );


  buf

  (
    n6955_o2_p,
    n6955_o2
  );


  not

  (
    n6955_o2_n,
    n6955_o2
  );


  buf

  (
    n6956_o2_p,
    n6956_o2
  );


  not

  (
    n6956_o2_n,
    n6956_o2
  );


  buf

  (
    n6957_o2_p,
    n6957_o2
  );


  not

  (
    n6957_o2_n,
    n6957_o2
  );


  buf

  (
    n6958_o2_p,
    n6958_o2
  );


  not

  (
    n6958_o2_n,
    n6958_o2
  );


  buf

  (
    n6982_o2_p,
    n6982_o2
  );


  not

  (
    n6982_o2_n,
    n6982_o2
  );


  buf

  (
    n6984_o2_p,
    n6984_o2
  );


  not

  (
    n6984_o2_n,
    n6984_o2
  );


  buf

  (
    n6974_o2_p,
    n6974_o2
  );


  not

  (
    n6974_o2_n,
    n6974_o2
  );


  buf

  (
    n6975_o2_p,
    n6975_o2
  );


  not

  (
    n6975_o2_n,
    n6975_o2
  );


  buf

  (
    n6999_o2_p,
    n6999_o2
  );


  not

  (
    n6999_o2_n,
    n6999_o2
  );


  buf

  (
    n7015_o2_p,
    n7015_o2
  );


  not

  (
    n7015_o2_n,
    n7015_o2
  );


  buf

  (
    n7016_o2_p,
    n7016_o2
  );


  not

  (
    n7016_o2_n,
    n7016_o2
  );


  buf

  (
    n7017_o2_p,
    n7017_o2
  );


  not

  (
    n7017_o2_n,
    n7017_o2
  );


  buf

  (
    n7018_o2_p,
    n7018_o2
  );


  not

  (
    n7018_o2_n,
    n7018_o2
  );


  buf

  (
    n7005_o2_p,
    n7005_o2
  );


  not

  (
    n7005_o2_n,
    n7005_o2
  );


  buf

  (
    n7019_o2_p,
    n7019_o2
  );


  not

  (
    n7019_o2_n,
    n7019_o2
  );


  buf

  (
    n7022_o2_p,
    n7022_o2
  );


  not

  (
    n7022_o2_n,
    n7022_o2
  );


  buf

  (
    n7023_o2_p,
    n7023_o2
  );


  not

  (
    n7023_o2_n,
    n7023_o2
  );


  buf

  (
    n7132_o2_p,
    n7132_o2
  );


  not

  (
    n7132_o2_n,
    n7132_o2
  );


  buf

  (
    n7133_o2_p,
    n7133_o2
  );


  not

  (
    n7133_o2_n,
    n7133_o2
  );


  buf

  (
    n7135_o2_p,
    n7135_o2
  );


  not

  (
    n7135_o2_n,
    n7135_o2
  );


  buf

  (
    n7136_o2_p,
    n7136_o2
  );


  not

  (
    n7136_o2_n,
    n7136_o2
  );


  buf

  (
    n7175_o2_p,
    n7175_o2
  );


  not

  (
    n7175_o2_n,
    n7175_o2
  );


  buf

  (
    n7155_o2_p,
    n7155_o2
  );


  not

  (
    n7155_o2_n,
    n7155_o2
  );


  buf

  (
    G3060_o2_p,
    G3060_o2
  );


  not

  (
    G3060_o2_n,
    G3060_o2
  );


  buf

  (
    n7383_o2_p,
    n7383_o2
  );


  not

  (
    n7383_o2_n,
    n7383_o2
  );


  buf

  (
    G3802_o2_p,
    G3802_o2
  );


  not

  (
    G3802_o2_n,
    G3802_o2
  );


  buf

  (
    G3859_o2_p,
    G3859_o2
  );


  not

  (
    G3859_o2_n,
    G3859_o2
  );


  buf

  (
    n7355_o2_p,
    n7355_o2
  );


  not

  (
    n7355_o2_n,
    n7355_o2
  );


  buf

  (
    n7356_o2_p,
    n7356_o2
  );


  not

  (
    n7356_o2_n,
    n7356_o2
  );


  buf

  (
    G4054_o2_p,
    G4054_o2
  );


  not

  (
    G4054_o2_n,
    G4054_o2
  );


  buf

  (
    G4068_o2_p,
    G4068_o2
  );


  not

  (
    G4068_o2_n,
    G4068_o2
  );


  buf

  (
    n7384_o2_p,
    n7384_o2
  );


  not

  (
    n7384_o2_n,
    n7384_o2
  );


  buf

  (
    n7387_o2_p,
    n7387_o2
  );


  not

  (
    n7387_o2_n,
    n7387_o2
  );


  buf

  (
    n7388_o2_p,
    n7388_o2
  );


  not

  (
    n7388_o2_n,
    n7388_o2
  );


  buf

  (
    n7389_o2_p,
    n7389_o2
  );


  not

  (
    n7389_o2_n,
    n7389_o2
  );


  buf

  (
    n7386_o2_p,
    n7386_o2
  );


  not

  (
    n7386_o2_n,
    n7386_o2
  );


  buf

  (
    n7453_o2_p,
    n7453_o2
  );


  not

  (
    n7453_o2_n,
    n7453_o2
  );


  buf

  (
    n7431_o2_p,
    n7431_o2
  );


  not

  (
    n7431_o2_n,
    n7431_o2
  );


  buf

  (
    n7432_o2_p,
    n7432_o2
  );


  not

  (
    n7432_o2_n,
    n7432_o2
  );


  buf

  (
    n7433_o2_p,
    n7433_o2
  );


  not

  (
    n7433_o2_n,
    n7433_o2
  );


  buf

  (
    n7430_o2_p,
    n7430_o2
  );


  not

  (
    n7430_o2_n,
    n7430_o2
  );


  buf

  (
    n7485_o2_p,
    n7485_o2
  );


  not

  (
    n7485_o2_n,
    n7485_o2
  );


  buf

  (
    n7486_o2_p,
    n7486_o2
  );


  not

  (
    n7486_o2_n,
    n7486_o2
  );


  buf

  (
    G2508_o2_p,
    G2508_o2
  );


  not

  (
    G2508_o2_n,
    G2508_o2
  );


  buf

  (
    G2486_o2_p,
    G2486_o2
  );


  not

  (
    G2486_o2_n,
    G2486_o2
  );


  buf

  (
    n2326_inv_p,
    n2326_inv
  );


  not

  (
    n2326_inv_n,
    n2326_inv
  );


  buf

  (
    n2329_inv_p,
    n2329_inv
  );


  not

  (
    n2329_inv_n,
    n2329_inv
  );


  buf

  (
    n3756_lo_buf_o2_p,
    n3756_lo_buf_o2
  );


  not

  (
    n3756_lo_buf_o2_n,
    n3756_lo_buf_o2
  );


  buf

  (
    n4056_lo_buf_o2_p,
    n4056_lo_buf_o2
  );


  not

  (
    n4056_lo_buf_o2_n,
    n4056_lo_buf_o2
  );


  buf

  (
    G3474_o2_p,
    G3474_o2
  );


  not

  (
    G3474_o2_n,
    G3474_o2
  );


  buf

  (
    n2341_inv_p,
    n2341_inv
  );


  not

  (
    n2341_inv_n,
    n2341_inv
  );


  buf

  (
    n7396_o2_p,
    n7396_o2
  );


  not

  (
    n7396_o2_n,
    n7396_o2
  );


  buf

  (
    n7398_o2_p,
    n7398_o2
  );


  not

  (
    n7398_o2_n,
    n7398_o2
  );


  buf

  (
    n7400_o2_p,
    n7400_o2
  );


  not

  (
    n7400_o2_n,
    n7400_o2
  );


  buf

  (
    n7401_o2_p,
    n7401_o2
  );


  not

  (
    n7401_o2_n,
    n7401_o2
  );


  buf

  (
    n7402_o2_p,
    n7402_o2
  );


  not

  (
    n7402_o2_n,
    n7402_o2
  );


  buf

  (
    n7403_o2_p,
    n7403_o2
  );


  not

  (
    n7403_o2_n,
    n7403_o2
  );


  buf

  (
    n7404_o2_p,
    n7404_o2
  );


  not

  (
    n7404_o2_n,
    n7404_o2
  );


  buf

  (
    n7405_o2_p,
    n7405_o2
  );


  not

  (
    n7405_o2_n,
    n7405_o2
  );


  buf

  (
    G2711_o2_p,
    G2711_o2
  );


  not

  (
    G2711_o2_n,
    G2711_o2
  );


  buf

  (
    n2371_inv_p,
    n2371_inv
  );


  not

  (
    n2371_inv_n,
    n2371_inv
  );


  buf

  (
    n7490_o2_p,
    n7490_o2
  );


  not

  (
    n7490_o2_n,
    n7490_o2
  );


  buf

  (
    n7527_o2_p,
    n7527_o2
  );


  not

  (
    n7527_o2_n,
    n7527_o2
  );


  buf

  (
    n7528_o2_p,
    n7528_o2
  );


  not

  (
    n7528_o2_n,
    n7528_o2
  );


  buf

  (
    n7529_o2_p,
    n7529_o2
  );


  not

  (
    n7529_o2_n,
    n7529_o2
  );


  buf

  (
    n7530_o2_p,
    n7530_o2
  );


  not

  (
    n7530_o2_n,
    n7530_o2
  );


  buf

  (
    n7523_o2_p,
    n7523_o2
  );


  not

  (
    n7523_o2_n,
    n7523_o2
  );


  buf

  (
    n7524_o2_p,
    n7524_o2
  );


  not

  (
    n7524_o2_n,
    n7524_o2
  );


  buf

  (
    n7525_o2_p,
    n7525_o2
  );


  not

  (
    n7525_o2_n,
    n7525_o2
  );


  buf

  (
    n7526_o2_p,
    n7526_o2
  );


  not

  (
    n7526_o2_n,
    n7526_o2
  );


  buf

  (
    n4296_lo_buf_o2_p,
    n4296_lo_buf_o2
  );


  not

  (
    n4296_lo_buf_o2_n,
    n4296_lo_buf_o2
  );


  buf

  (
    n4368_lo_buf_o2_p,
    n4368_lo_buf_o2
  );


  not

  (
    n4368_lo_buf_o2_n,
    n4368_lo_buf_o2
  );


  buf

  (
    G2466_o2_p,
    G2466_o2
  );


  not

  (
    G2466_o2_n,
    G2466_o2
  );


  buf

  (
    G2404_o2_p,
    G2404_o2
  );


  not

  (
    G2404_o2_n,
    G2404_o2
  );


  buf

  (
    n7534_o2_p,
    n7534_o2
  );


  not

  (
    n7534_o2_n,
    n7534_o2
  );


  buf

  (
    n7535_o2_p,
    n7535_o2
  );


  not

  (
    n7535_o2_n,
    n7535_o2
  );


  buf

  (
    n7536_o2_p,
    n7536_o2
  );


  not

  (
    n7536_o2_n,
    n7536_o2
  );


  buf

  (
    n7533_o2_p,
    n7533_o2
  );


  not

  (
    n7533_o2_n,
    n7533_o2
  );


  buf

  (
    G1060_o2_p,
    G1060_o2
  );


  not

  (
    G1060_o2_n,
    G1060_o2
  );


  buf

  (
    G963_o2_p,
    G963_o2
  );


  not

  (
    G963_o2_n,
    G963_o2
  );


  buf

  (
    G2448_o2_p,
    G2448_o2
  );


  not

  (
    G2448_o2_n,
    G2448_o2
  );


  buf

  (
    G2685_o2_p,
    G2685_o2
  );


  not

  (
    G2685_o2_n,
    G2685_o2
  );


  buf

  (
    G2679_o2_p,
    G2679_o2
  );


  not

  (
    G2679_o2_n,
    G2679_o2
  );


  buf

  (
    G2774_o2_p,
    G2774_o2
  );


  not

  (
    G2774_o2_n,
    G2774_o2
  );


  buf

  (
    G2780_o2_p,
    G2780_o2
  );


  not

  (
    G2780_o2_n,
    G2780_o2
  );


  buf

  (
    G2759_o2_p,
    G2759_o2
  );


  not

  (
    G2759_o2_n,
    G2759_o2
  );


  buf

  (
    G2737_o2_p,
    G2737_o2
  );


  not

  (
    G2737_o2_n,
    G2737_o2
  );


  buf

  (
    G2850_o2_p,
    G2850_o2
  );


  not

  (
    G2850_o2_n,
    G2850_o2
  );


  buf

  (
    G3393_o2_p,
    G3393_o2
  );


  not

  (
    G3393_o2_n,
    G3393_o2
  );


  buf

  (
    G3404_o2_p,
    G3404_o2
  );


  not

  (
    G3404_o2_n,
    G3404_o2
  );


  buf

  (
    G3559_o2_p,
    G3559_o2
  );


  not

  (
    G3559_o2_n,
    G3559_o2
  );


  buf

  (
    G2744_o2_p,
    G2744_o2
  );


  not

  (
    G2744_o2_n,
    G2744_o2
  );


  buf

  (
    n3708_lo_buf_o2_p,
    n3708_lo_buf_o2
  );


  not

  (
    n3708_lo_buf_o2_n,
    n3708_lo_buf_o2
  );


  buf

  (
    n3840_lo_buf_o2_p,
    n3840_lo_buf_o2
  );


  not

  (
    n3840_lo_buf_o2_n,
    n3840_lo_buf_o2
  );


  buf

  (
    n4008_lo_buf_o2_p,
    n4008_lo_buf_o2
  );


  not

  (
    n4008_lo_buf_o2_n,
    n4008_lo_buf_o2
  );


  buf

  (
    n4104_lo_buf_o2_p,
    n4104_lo_buf_o2
  );


  not

  (
    n4104_lo_buf_o2_n,
    n4104_lo_buf_o2
  );


  buf

  (
    G1821_o2_p,
    G1821_o2
  );


  not

  (
    G1821_o2_n,
    G1821_o2
  );


  buf

  (
    G1734_o2_p,
    G1734_o2
  );


  not

  (
    G1734_o2_n,
    G1734_o2
  );


  buf

  (
    G3517_o2_p,
    G3517_o2
  );


  not

  (
    G3517_o2_n,
    G3517_o2
  );


  buf

  (
    G3533_o2_p,
    G3533_o2
  );


  not

  (
    G3533_o2_n,
    G3533_o2
  );


  buf

  (
    G3629_o2_p,
    G3629_o2
  );


  not

  (
    G3629_o2_n,
    G3629_o2
  );


  buf

  (
    G3645_o2_p,
    G3645_o2
  );


  not

  (
    G3645_o2_n,
    G3645_o2
  );


  buf

  (
    n2497_inv_p,
    n2497_inv
  );


  not

  (
    n2497_inv_n,
    n2497_inv
  );


  buf

  (
    G2731_o2_p,
    G2731_o2
  );


  not

  (
    G2731_o2_n,
    G2731_o2
  );


  buf

  (
    G2844_o2_p,
    G2844_o2
  );


  not

  (
    G2844_o2_n,
    G2844_o2
  );


  buf

  (
    n3732_lo_buf_o2_p,
    n3732_lo_buf_o2
  );


  not

  (
    n3732_lo_buf_o2_n,
    n3732_lo_buf_o2
  );


  buf

  (
    n4032_lo_buf_o2_p,
    n4032_lo_buf_o2
  );


  not

  (
    n4032_lo_buf_o2_n,
    n4032_lo_buf_o2
  );


  buf

  (
    G3552_o2_p,
    G3552_o2
  );


  not

  (
    G3552_o2_n,
    G3552_o2
  );


  buf

  (
    G2271_o2_p,
    G2271_o2
  );


  not

  (
    G2271_o2_n,
    G2271_o2
  );


  buf

  (
    n4248_lo_buf_o2_p,
    n4248_lo_buf_o2
  );


  not

  (
    n4248_lo_buf_o2_n,
    n4248_lo_buf_o2
  );


  buf

  (
    n4332_lo_buf_o2_p,
    n4332_lo_buf_o2
  );


  not

  (
    n4332_lo_buf_o2_n,
    n4332_lo_buf_o2
  );


  buf

  (
    n4344_lo_buf_o2_p,
    n4344_lo_buf_o2
  );


  not

  (
    n4344_lo_buf_o2_n,
    n4344_lo_buf_o2
  );


  buf

  (
    n4380_lo_buf_o2_p,
    n4380_lo_buf_o2
  );


  not

  (
    n4380_lo_buf_o2_n,
    n4380_lo_buf_o2
  );


  buf

  (
    G2398_o2_p,
    G2398_o2
  );


  not

  (
    G2398_o2_n,
    G2398_o2
  );


  buf

  (
    G2480_o2_p,
    G2480_o2
  );


  not

  (
    G2480_o2_n,
    G2480_o2
  );


  buf

  (
    G2418_o2_p,
    G2418_o2
  );


  not

  (
    G2418_o2_n,
    G2418_o2
  );


  buf

  (
    G1455_o2_p,
    G1455_o2
  );


  not

  (
    G1455_o2_n,
    G1455_o2
  );


  buf

  (
    G1449_o2_p,
    G1449_o2
  );


  not

  (
    G1449_o2_n,
    G1449_o2
  );


  buf

  (
    G1452_o2_p,
    G1452_o2
  );


  not

  (
    G1452_o2_n,
    G1452_o2
  );


  buf

  (
    G1425_o2_p,
    G1425_o2
  );


  not

  (
    G1425_o2_n,
    G1425_o2
  );


  buf

  (
    G1428_o2_p,
    G1428_o2
  );


  not

  (
    G1428_o2_n,
    G1428_o2
  );


  buf

  (
    G1419_o2_p,
    G1419_o2
  );


  not

  (
    G1419_o2_n,
    G1419_o2
  );


  buf

  (
    G1422_o2_p,
    G1422_o2
  );


  not

  (
    G1422_o2_n,
    G1422_o2
  );


  buf

  (
    n4308_lo_buf_o2_p,
    n4308_lo_buf_o2
  );


  not

  (
    n4308_lo_buf_o2_n,
    n4308_lo_buf_o2
  );


  buf

  (
    G2675_o2_p,
    G2675_o2
  );


  not

  (
    G2675_o2_n,
    G2675_o2
  );


  buf

  (
    G3035_o2_p,
    G3035_o2
  );


  not

  (
    G3035_o2_n,
    G3035_o2
  );


  buf

  (
    G3026_o2_p,
    G3026_o2
  );


  not

  (
    G3026_o2_n,
    G3026_o2
  );


  buf

  (
    G3029_o2_p,
    G3029_o2
  );


  not

  (
    G3029_o2_n,
    G3029_o2
  );


  buf

  (
    G3032_o2_p,
    G3032_o2
  );


  not

  (
    G3032_o2_n,
    G3032_o2
  );


  buf

  (
    G2999_o2_p,
    G2999_o2
  );


  not

  (
    G2999_o2_n,
    G2999_o2
  );


  buf

  (
    G3002_o2_p,
    G3002_o2
  );


  not

  (
    G3002_o2_n,
    G3002_o2
  );


  buf

  (
    G2770_o2_p,
    G2770_o2
  );


  not

  (
    G2770_o2_n,
    G2770_o2
  );


  buf

  (
    G3008_o2_p,
    G3008_o2
  );


  not

  (
    G3008_o2_n,
    G3008_o2
  );


  buf

  (
    G2073_o2_p,
    G2073_o2
  );


  not

  (
    G2073_o2_n,
    G2073_o2
  );


  buf

  (
    G2752_o2_p,
    G2752_o2
  );


  not

  (
    G2752_o2_n,
    G2752_o2
  );


  buf

  (
    G3005_o2_p,
    G3005_o2
  );


  not

  (
    G3005_o2_n,
    G3005_o2
  );


  buf

  (
    G5108_o2_p,
    G5108_o2
  );


  not

  (
    G5108_o2_n,
    G5108_o2
  );


  buf

  (
    G5135_o2_p,
    G5135_o2
  );


  not

  (
    G5135_o2_n,
    G5135_o2
  );


  buf

  (
    G5111_o2_p,
    G5111_o2
  );


  not

  (
    G5111_o2_n,
    G5111_o2
  );


  buf

  (
    G5138_o2_p,
    G5138_o2
  );


  not

  (
    G5138_o2_n,
    G5138_o2
  );


  buf

  (
    G3415_o2_p,
    G3415_o2
  );


  not

  (
    G3415_o2_n,
    G3415_o2
  );


  buf

  (
    G3386_o2_p,
    G3386_o2
  );


  not

  (
    G3386_o2_n,
    G3386_o2
  );


  buf

  (
    G3570_o2_p,
    G3570_o2
  );


  not

  (
    G3570_o2_n,
    G3570_o2
  );


  buf

  (
    G2430_o2_p,
    G2430_o2
  );


  not

  (
    G2430_o2_n,
    G2430_o2
  );


  buf

  (
    G3495_o2_p,
    G3495_o2
  );


  not

  (
    G3495_o2_n,
    G3495_o2
  );


  buf

  (
    G3621_o2_p,
    G3621_o2
  );


  not

  (
    G3621_o2_n,
    G3621_o2
  );


  buf

  (
    n4284_lo_buf_o2_p,
    n4284_lo_buf_o2
  );


  not

  (
    n4284_lo_buf_o2_n,
    n4284_lo_buf_o2
  );


  buf

  (
    n4356_lo_buf_o2_p,
    n4356_lo_buf_o2
  );


  not

  (
    n4356_lo_buf_o2_n,
    n4356_lo_buf_o2
  );


  buf

  (
    G2472_o2_p,
    G2472_o2
  );


  not

  (
    G2472_o2_n,
    G2472_o2
  );


  buf

  (
    G2410_o2_p,
    G2410_o2
  );


  not

  (
    G2410_o2_n,
    G2410_o2
  );


  buf

  (
    n3960_lo_buf_o2_p,
    n3960_lo_buf_o2
  );


  not

  (
    n3960_lo_buf_o2_n,
    n3960_lo_buf_o2
  );


  buf

  (
    n3972_lo_buf_o2_p,
    n3972_lo_buf_o2
  );


  not

  (
    n3972_lo_buf_o2_n,
    n3972_lo_buf_o2
  );


  buf

  (
    n2647_inv_p,
    n2647_inv
  );


  not

  (
    n2647_inv_n,
    n2647_inv
  );


  buf

  (
    n2650_inv_p,
    n2650_inv
  );


  not

  (
    n2650_inv_n,
    n2650_inv
  );


  buf

  (
    n3684_lo_buf_o2_p,
    n3684_lo_buf_o2
  );


  not

  (
    n3684_lo_buf_o2_n,
    n3684_lo_buf_o2
  );


  buf

  (
    n4080_lo_buf_o2_p,
    n4080_lo_buf_o2
  );


  not

  (
    n4080_lo_buf_o2_n,
    n4080_lo_buf_o2
  );


  buf

  (
    n4092_lo_buf_o2_p,
    n4092_lo_buf_o2
  );


  not

  (
    n4092_lo_buf_o2_n,
    n4092_lo_buf_o2
  );


  buf

  (
    n2662_inv_p,
    n2662_inv
  );


  not

  (
    n2662_inv_n,
    n2662_inv
  );


  buf

  (
    n2665_inv_p,
    n2665_inv
  );


  not

  (
    n2665_inv_n,
    n2665_inv
  );


  buf

  (
    G1147_o2_p,
    G1147_o2
  );


  not

  (
    G1147_o2_n,
    G1147_o2
  );


  buf

  (
    G2705_o2_p,
    G2705_o2
  );


  not

  (
    G2705_o2_n,
    G2705_o2
  );


  buf

  (
    G2693_o2_p,
    G2693_o2
  );


  not

  (
    G2693_o2_n,
    G2693_o2
  );


  buf

  (
    G2696_o2_p,
    G2696_o2
  );


  not

  (
    G2696_o2_n,
    G2696_o2
  );


  buf

  (
    G2700_o2_p,
    G2700_o2
  );


  not

  (
    G2700_o2_n,
    G2700_o2
  );


  buf

  (
    G2915_o2_p,
    G2915_o2
  );


  not

  (
    G2915_o2_n,
    G2915_o2
  );


  buf

  (
    G2966_o2_p,
    G2966_o2
  );


  not

  (
    G2966_o2_n,
    G2966_o2
  );


  buf

  (
    G2540_o2_p,
    G2540_o2
  );


  not

  (
    G2540_o2_n,
    G2540_o2
  );


  buf

  (
    G2788_o2_p,
    G2788_o2
  );


  not

  (
    G2788_o2_n,
    G2788_o2
  );


  buf

  (
    G2792_o2_p,
    G2792_o2
  );


  not

  (
    G2792_o2_n,
    G2792_o2
  );


  buf

  (
    G2797_o2_p,
    G2797_o2
  );


  not

  (
    G2797_o2_n,
    G2797_o2
  );


  buf

  (
    G2804_o2_p,
    G2804_o2
  );


  not

  (
    G2804_o2_n,
    G2804_o2
  );


  buf

  (
    G1038_o2_p,
    G1038_o2
  );


  not

  (
    G1038_o2_n,
    G1038_o2
  );


  buf

  (
    G1044_o2_p,
    G1044_o2
  );


  not

  (
    G1044_o2_n,
    G1044_o2
  );


  buf

  (
    G1090_o2_p,
    G1090_o2
  );


  not

  (
    G1090_o2_n,
    G1090_o2
  );


  buf

  (
    G1096_o2_p,
    G1096_o2
  );


  not

  (
    G1096_o2_n,
    G1096_o2
  );


  buf

  (
    G1029_o2_p,
    G1029_o2
  );


  not

  (
    G1029_o2_n,
    G1029_o2
  );


  buf

  (
    G3942_o2_p,
    G3942_o2
  );


  not

  (
    G3942_o2_n,
    G3942_o2
  );


  buf

  (
    G3954_o2_p,
    G3954_o2
  );


  not

  (
    G3954_o2_n,
    G3954_o2
  );


  buf

  (
    G4011_o2_p,
    G4011_o2
  );


  not

  (
    G4011_o2_n,
    G4011_o2
  );


  buf

  (
    G4017_o2_p,
    G4017_o2
  );


  not

  (
    G4017_o2_n,
    G4017_o2
  );


  buf

  (
    G1141_o2_p,
    G1141_o2
  );


  not

  (
    G1141_o2_n,
    G1141_o2
  );


  buf

  (
    G1081_o2_p,
    G1081_o2
  );


  not

  (
    G1081_o2_n,
    G1081_o2
  );


  buf

  (
    G2146_o2_p,
    G2146_o2
  );


  not

  (
    G2146_o2_n,
    G2146_o2
  );


  buf

  (
    G2145_o2_p,
    G2145_o2
  );


  not

  (
    G2145_o2_n,
    G2145_o2
  );


  buf

  (
    G2144_o2_p,
    G2144_o2
  );


  not

  (
    G2144_o2_n,
    G2144_o2
  );


  buf

  (
    G2143_o2_p,
    G2143_o2
  );


  not

  (
    G2143_o2_n,
    G2143_o2
  );


  buf

  (
    G2142_o2_p,
    G2142_o2
  );


  not

  (
    G2142_o2_n,
    G2142_o2
  );


  buf

  (
    G2141_o2_p,
    G2141_o2
  );


  not

  (
    G2141_o2_n,
    G2141_o2
  );


  buf

  (
    G2140_o2_p,
    G2140_o2
  );


  not

  (
    G2140_o2_n,
    G2140_o2
  );


  buf

  (
    G2139_o2_p,
    G2139_o2
  );


  not

  (
    G2139_o2_n,
    G2139_o2
  );


  buf

  (
    G3769_o2_p,
    G3769_o2
  );


  not

  (
    G3769_o2_n,
    G3769_o2
  );


  buf

  (
    G3773_o2_p,
    G3773_o2
  );


  not

  (
    G3773_o2_n,
    G3773_o2
  );


  buf

  (
    G3768_o2_p,
    G3768_o2
  );


  not

  (
    G3768_o2_n,
    G3768_o2
  );


  buf

  (
    G4101_o2_p,
    G4101_o2
  );


  not

  (
    G4101_o2_n,
    G4101_o2
  );


  buf

  (
    G3161_o2_p,
    G3161_o2
  );


  not

  (
    G3161_o2_n,
    G3161_o2
  );


  buf

  (
    G4143_o2_p,
    G4143_o2
  );


  not

  (
    G4143_o2_n,
    G4143_o2
  );


  buf

  (
    G3828_o2_p,
    G3828_o2
  );


  not

  (
    G3828_o2_n,
    G3828_o2
  );


  buf

  (
    G3831_o2_p,
    G3831_o2
  );


  not

  (
    G3831_o2_n,
    G3831_o2
  );


  buf

  (
    G3334_o2_p,
    G3334_o2
  );


  not

  (
    G3334_o2_n,
    G3334_o2
  );


  buf

  (
    G3335_o2_p,
    G3335_o2
  );


  not

  (
    G3335_o2_n,
    G3335_o2
  );


  buf

  (
    G3180_o2_p,
    G3180_o2
  );


  not

  (
    G3180_o2_n,
    G3180_o2
  );


  buf

  (
    G3340_o2_p,
    G3340_o2
  );


  not

  (
    G3340_o2_n,
    G3340_o2
  );


  buf

  (
    G3339_o2_p,
    G3339_o2
  );


  not

  (
    G3339_o2_n,
    G3339_o2
  );


  buf

  (
    G3341_o2_p,
    G3341_o2
  );


  not

  (
    G3341_o2_n,
    G3341_o2
  );


  buf

  (
    G3234_o2_p,
    G3234_o2
  );


  not

  (
    G3234_o2_n,
    G3234_o2
  );


  buf

  (
    G3829_o2_p,
    G3829_o2
  );


  not

  (
    G3829_o2_n,
    G3829_o2
  );


  buf

  (
    G3338_o2_p,
    G3338_o2
  );


  not

  (
    G3338_o2_n,
    G3338_o2
  );


  buf

  (
    G3336_o2_p,
    G3336_o2
  );


  not

  (
    G3336_o2_n,
    G3336_o2
  );


  buf

  (
    G3770_o2_p,
    G3770_o2
  );


  not

  (
    G3770_o2_n,
    G3770_o2
  );


  buf

  (
    G3918_o2_p,
    G3918_o2
  );


  not

  (
    G3918_o2_n,
    G3918_o2
  );


  buf

  (
    G3774_o2_p,
    G3774_o2
  );


  not

  (
    G3774_o2_n,
    G3774_o2
  );


  buf

  (
    G3921_o2_p,
    G3921_o2
  );


  not

  (
    G3921_o2_n,
    G3921_o2
  );


  buf

  (
    G3832_o2_p,
    G3832_o2
  );


  not

  (
    G3832_o2_n,
    G3832_o2
  );


  buf

  (
    G3993_o2_p,
    G3993_o2
  );


  not

  (
    G3993_o2_n,
    G3993_o2
  );


  buf

  (
    G2076_o2_p,
    G2076_o2
  );


  not

  (
    G2076_o2_n,
    G2076_o2
  );


  buf

  (
    G2071_o2_p,
    G2071_o2
  );


  not

  (
    G2071_o2_n,
    G2071_o2
  );


  buf

  (
    G2072_o2_p,
    G2072_o2
  );


  not

  (
    G2072_o2_n,
    G2072_o2
  );


  buf

  (
    G2069_o2_p,
    G2069_o2
  );


  not

  (
    G2069_o2_n,
    G2069_o2
  );


  buf

  (
    G2070_o2_p,
    G2070_o2
  );


  not

  (
    G2070_o2_n,
    G2070_o2
  );


  buf

  (
    G2067_o2_p,
    G2067_o2
  );


  not

  (
    G2067_o2_n,
    G2067_o2
  );


  buf

  (
    G2068_o2_p,
    G2068_o2
  );


  not

  (
    G2068_o2_n,
    G2068_o2
  );


  buf

  (
    G4095_o2_p,
    G4095_o2
  );


  not

  (
    G4095_o2_n,
    G4095_o2
  );


  buf

  (
    G3272_o2_p,
    G3272_o2
  );


  not

  (
    G3272_o2_n,
    G3272_o2
  );


  buf

  (
    G3269_o2_p,
    G3269_o2
  );


  not

  (
    G3269_o2_n,
    G3269_o2
  );


  buf

  (
    G3270_o2_p,
    G3270_o2
  );


  not

  (
    G3270_o2_n,
    G3270_o2
  );


  buf

  (
    G3271_o2_p,
    G3271_o2
  );


  not

  (
    G3271_o2_n,
    G3271_o2
  );


  buf

  (
    G3265_o2_p,
    G3265_o2
  );


  not

  (
    G3265_o2_n,
    G3265_o2
  );


  buf

  (
    G3266_o2_p,
    G3266_o2
  );


  not

  (
    G3266_o2_n,
    G3266_o2
  );


  buf

  (
    G4137_o2_p,
    G4137_o2
  );


  not

  (
    G4137_o2_n,
    G4137_o2
  );


  buf

  (
    G3268_o2_p,
    G3268_o2
  );


  not

  (
    G3268_o2_n,
    G3268_o2
  );


  buf

  (
    G2361_o2_p,
    G2361_o2
  );


  not

  (
    G2361_o2_n,
    G2361_o2
  );


  buf

  (
    G3228_o2_p,
    G3228_o2
  );


  not

  (
    G3228_o2_n,
    G3228_o2
  );


  buf

  (
    G3267_o2_p,
    G3267_o2
  );


  not

  (
    G3267_o2_n,
    G3267_o2
  );


  buf

  (
    G2336_o2_p,
    G2336_o2
  );


  not

  (
    G2336_o2_n,
    G2336_o2
  );


  buf

  (
    G3459_o2_p,
    G3459_o2
  );


  not

  (
    G3459_o2_n,
    G3459_o2
  );


  buf

  (
    G3428_o2_p,
    G3428_o2
  );


  not

  (
    G3428_o2_n,
    G3428_o2
  );


  buf

  (
    G3438_o2_p,
    G3438_o2
  );


  not

  (
    G3438_o2_n,
    G3438_o2
  );


  buf

  (
    G3449_o2_p,
    G3449_o2
  );


  not

  (
    G3449_o2_n,
    G3449_o2
  );


  buf

  (
    G3421_o2_p,
    G3421_o2
  );


  not

  (
    G3421_o2_n,
    G3421_o2
  );


  buf

  (
    G3576_o2_p,
    G3576_o2
  );


  not

  (
    G3576_o2_n,
    G3576_o2
  );


  buf

  (
    G3303_o2_p,
    G3303_o2
  );


  not

  (
    G3303_o2_n,
    G3303_o2
  );


  buf

  (
    G3583_o2_p,
    G3583_o2
  );


  not

  (
    G3583_o2_n,
    G3583_o2
  );


  buf

  (
    G3594_o2_p,
    G3594_o2
  );


  not

  (
    G3594_o2_n,
    G3594_o2
  );


  buf

  (
    G3674_o2_p,
    G3674_o2
  );


  not

  (
    G3674_o2_n,
    G3674_o2
  );


  buf

  (
    G3685_o2_p,
    G3685_o2
  );


  not

  (
    G3685_o2_n,
    G3685_o2
  );


  buf

  (
    G4504_o2_p,
    G4504_o2
  );


  not

  (
    G4504_o2_n,
    G4504_o2
  );


  buf

  (
    G4180_o2_p,
    G4180_o2
  );


  not

  (
    G4180_o2_n,
    G4180_o2
  );


  buf

  (
    G5123_o2_p,
    G5123_o2
  );


  not

  (
    G5123_o2_n,
    G5123_o2
  );


  buf

  (
    G5142_o2_p,
    G5142_o2
  );


  not

  (
    G5142_o2_n,
    G5142_o2
  );


  buf

  (
    G5126_o2_p,
    G5126_o2
  );


  not

  (
    G5126_o2_n,
    G5126_o2
  );


  buf

  (
    G5144_o2_p,
    G5144_o2
  );


  not

  (
    G5144_o2_n,
    G5144_o2
  );


  buf

  (
    G3912_o2_p,
    G3912_o2
  );


  not

  (
    G3912_o2_n,
    G3912_o2
  );


  buf

  (
    G4417_o2_p,
    G4417_o2
  );


  not

  (
    G4417_o2_n,
    G4417_o2
  );


  buf

  (
    G4420_o2_p,
    G4420_o2
  );


  not

  (
    G4420_o2_n,
    G4420_o2
  );


  buf

  (
    G3969_o2_p,
    G3969_o2
  );


  not

  (
    G3969_o2_n,
    G3969_o2
  );


  buf

  (
    G4023_o2_p,
    G4023_o2
  );


  not

  (
    G4023_o2_n,
    G4023_o2
  );


  buf

  (
    G2720_o2_p,
    G2720_o2
  );


  not

  (
    G2720_o2_n,
    G2720_o2
  );


  buf

  (
    G2837_o2_p,
    G2837_o2
  );


  not

  (
    G2837_o2_n,
    G2837_o2
  );


  buf

  (
    n2965_inv_p,
    n2965_inv
  );


  not

  (
    n2965_inv_n,
    n2965_inv
  );


  buf

  (
    n2968_inv_p,
    n2968_inv
  );


  not

  (
    n2968_inv_n,
    n2968_inv
  );


  buf

  (
    n2971_inv_p,
    n2971_inv
  );


  not

  (
    n2971_inv_n,
    n2971_inv
  );


  buf

  (
    n2974_inv_p,
    n2974_inv
  );


  not

  (
    n2974_inv_n,
    n2974_inv
  );


  buf

  (
    G1876_o2_p,
    G1876_o2
  );


  not

  (
    G1876_o2_n,
    G1876_o2
  );


  buf

  (
    G4996_o2_p,
    G4996_o2
  );


  not

  (
    G4996_o2_n,
    G4996_o2
  );


  buf

  (
    G4984_o2_p,
    G4984_o2
  );


  not

  (
    G4984_o2_n,
    G4984_o2
  );


  buf

  (
    G4920_o2_p,
    G4920_o2
  );


  not

  (
    G4920_o2_n,
    G4920_o2
  );


  buf

  (
    G4923_o2_p,
    G4923_o2
  );


  not

  (
    G4923_o2_n,
    G4923_o2
  );


  buf

  (
    G4930_o2_p,
    G4930_o2
  );


  not

  (
    G4930_o2_n,
    G4930_o2
  );


  buf

  (
    G4933_o2_p,
    G4933_o2
  );


  not

  (
    G4933_o2_n,
    G4933_o2
  );


  buf

  (
    n4320_lo_buf_o2_p,
    n4320_lo_buf_o2
  );


  not

  (
    n4320_lo_buf_o2_n,
    n4320_lo_buf_o2
  );


  buf

  (
    G2424_o2_p,
    G2424_o2
  );


  not

  (
    G2424_o2_n,
    G2424_o2
  );


  buf

  (
    G3317_o2_p,
    G3317_o2
  );


  not

  (
    G3317_o2_n,
    G3317_o2
  );


  buf

  (
    G3503_o2_p,
    G3503_o2
  );


  not

  (
    G3503_o2_n,
    G3503_o2
  );


  buf

  (
    G3485_o2_p,
    G3485_o2
  );


  not

  (
    G3485_o2_n,
    G3485_o2
  );


  buf

  (
    G3611_o2_p,
    G3611_o2
  );


  not

  (
    G3611_o2_n,
    G3611_o2
  );


  buf

  (
    n3864_lo_buf_o2_p,
    n3864_lo_buf_o2
  );


  not

  (
    n3864_lo_buf_o2_n,
    n3864_lo_buf_o2
  );


  buf

  (
    n3888_lo_buf_o2_p,
    n3888_lo_buf_o2
  );


  not

  (
    n3888_lo_buf_o2_n,
    n3888_lo_buf_o2
  );


  buf

  (
    n4116_lo_buf_o2_p,
    n4116_lo_buf_o2
  );


  not

  (
    n4116_lo_buf_o2_n,
    n4116_lo_buf_o2
  );


  buf

  (
    n4128_lo_buf_o2_p,
    n4128_lo_buf_o2
  );


  not

  (
    n4128_lo_buf_o2_n,
    n4128_lo_buf_o2
  );


  buf

  (
    n4140_lo_buf_o2_p,
    n4140_lo_buf_o2
  );


  not

  (
    n4140_lo_buf_o2_n,
    n4140_lo_buf_o2
  );


  buf

  (
    n4152_lo_buf_o2_p,
    n4152_lo_buf_o2
  );


  not

  (
    n4152_lo_buf_o2_n,
    n4152_lo_buf_o2
  );


  buf

  (
    G1815_o2_p,
    G1815_o2
  );


  not

  (
    G1815_o2_n,
    G1815_o2
  );


  buf

  (
    G1728_o2_p,
    G1728_o2
  );


  not

  (
    G1728_o2_n,
    G1728_o2
  );


  buf

  (
    G1035_o2_p,
    G1035_o2
  );


  not

  (
    G1035_o2_n,
    G1035_o2
  );


  buf

  (
    G1041_o2_p,
    G1041_o2
  );


  not

  (
    G1041_o2_n,
    G1041_o2
  );


  buf

  (
    G1087_o2_p,
    G1087_o2
  );


  not

  (
    G1087_o2_n,
    G1087_o2
  );


  buf

  (
    G1093_o2_p,
    G1093_o2
  );


  not

  (
    G1093_o2_n,
    G1093_o2
  );


  buf

  (
    G1132_o2_p,
    G1132_o2
  );


  not

  (
    G1132_o2_n,
    G1132_o2
  );


  buf

  (
    G1108_o2_p,
    G1108_o2
  );


  not

  (
    G1108_o2_n,
    G1108_o2
  );


  buf

  (
    G1138_o2_p,
    G1138_o2
  );


  not

  (
    G1138_o2_n,
    G1138_o2
  );


  buf

  (
    G1114_o2_p,
    G1114_o2
  );


  not

  (
    G1114_o2_n,
    G1114_o2
  );


  buf

  (
    G1807_o2_p,
    G1807_o2
  );


  not

  (
    G1807_o2_n,
    G1807_o2
  );


  buf

  (
    G2108_o2_p,
    G2108_o2
  );


  not

  (
    G2108_o2_n,
    G2108_o2
  );


  buf

  (
    G1126_o2_p,
    G1126_o2
  );


  not

  (
    G1126_o2_n,
    G1126_o2
  );


  buf

  (
    G1899_o2_p,
    G1899_o2
  );


  not

  (
    G1899_o2_n,
    G1899_o2
  );


  buf

  (
    G2134_o2_p,
    G2134_o2
  );


  not

  (
    G2134_o2_n,
    G2134_o2
  );


  buf

  (
    G1852_o2_p,
    G1852_o2
  );


  not

  (
    G1852_o2_n,
    G1852_o2
  );


  buf

  (
    G2116_o2_p,
    G2116_o2
  );


  not

  (
    G2116_o2_n,
    G2116_o2
  );


  buf

  (
    G2543_o2_p,
    G2543_o2
  );


  not

  (
    G2543_o2_n,
    G2543_o2
  );


  buf

  (
    G2727_o2_p,
    G2727_o2
  );


  not

  (
    G2727_o2_n,
    G2727_o2
  );


  buf

  (
    G2715_o2_p,
    G2715_o2
  );


  not

  (
    G2715_o2_n,
    G2715_o2
  );


  buf

  (
    G2832_o2_p,
    G2832_o2
  );


  not

  (
    G2832_o2_n,
    G2832_o2
  );


  buf

  (
    G1873_o2_p,
    G1873_o2
  );


  not

  (
    G1873_o2_n,
    G1873_o2
  );


  buf

  (
    G3291_o2_p,
    G3291_o2
  );


  not

  (
    G3291_o2_n,
    G3291_o2
  );


  buf

  (
    G5025_o2_p,
    G5025_o2
  );


  not

  (
    G5025_o2_n,
    G5025_o2
  );


  buf

  (
    G5036_o2_p,
    G5036_o2
  );


  not

  (
    G5036_o2_n,
    G5036_o2
  );


  buf

  (
    G3132_o2_p,
    G3132_o2
  );


  not

  (
    G3132_o2_n,
    G3132_o2
  );


  buf

  (
    G5038_o2_p,
    G5038_o2
  );


  not

  (
    G5038_o2_n,
    G5038_o2
  );


  buf

  (
    G5039_o2_p,
    G5039_o2
  );


  not

  (
    G5039_o2_n,
    G5039_o2
  );


  buf

  (
    n3118_inv_p,
    n3118_inv
  );


  not

  (
    n3118_inv_n,
    n3118_inv
  );


  buf

  (
    n3121_inv_p,
    n3121_inv
  );


  not

  (
    n3121_inv_n,
    n3121_inv
  );


  buf

  (
    n3124_inv_p,
    n3124_inv
  );


  not

  (
    n3124_inv_n,
    n3124_inv
  );


  buf

  (
    n3127_inv_p,
    n3127_inv
  );


  not

  (
    n3127_inv_n,
    n3127_inv
  );


  buf

  (
    n3984_lo_buf_o2_p,
    n3984_lo_buf_o2
  );


  not

  (
    n3984_lo_buf_o2_n,
    n3984_lo_buf_o2
  );


  buf

  (
    G1802_o2_p,
    G1802_o2
  );


  not

  (
    G1802_o2_n,
    G1802_o2
  );


  buf

  (
    G1804_o2_p,
    G1804_o2
  );


  not

  (
    G1804_o2_n,
    G1804_o2
  );


  buf

  (
    G1849_o2_p,
    G1849_o2
  );


  not

  (
    G1849_o2_n,
    G1849_o2
  );


  buf

  (
    G1851_o2_p,
    G1851_o2
  );


  not

  (
    G1851_o2_n,
    G1851_o2
  );


  buf

  (
    G2492_o2_p,
    G2492_o2
  );


  not

  (
    G2492_o2_n,
    G2492_o2
  );


  buf

  (
    G1799_o2_p,
    G1799_o2
  );


  not

  (
    G1799_o2_n,
    G1799_o2
  );


  buf

  (
    G4231_o2_p,
    G4231_o2
  );


  not

  (
    G4231_o2_n,
    G4231_o2
  );


  buf

  (
    G4234_o2_p,
    G4234_o2
  );


  not

  (
    G4234_o2_n,
    G4234_o2
  );


  buf

  (
    G4245_o2_p,
    G4245_o2
  );


  not

  (
    G4245_o2_n,
    G4245_o2
  );


  buf

  (
    G4247_o2_p,
    G4247_o2
  );


  not

  (
    G4247_o2_n,
    G4247_o2
  );


  buf

  (
    G1894_o2_p,
    G1894_o2
  );


  not

  (
    G1894_o2_n,
    G1894_o2
  );


  buf

  (
    G1846_o2_p,
    G1846_o2
  );


  not

  (
    G1846_o2_n,
    G1846_o2
  );


  buf

  (
    G4238_o2_p,
    G4238_o2
  );


  not

  (
    G4238_o2_n,
    G4238_o2
  );


  buf

  (
    G4249_o2_p,
    G4249_o2
  );


  not

  (
    G4249_o2_n,
    G4249_o2
  );


  buf

  (
    G2293_o2_p,
    G2293_o2
  );


  not

  (
    G2293_o2_n,
    G2293_o2
  );


  buf

  (
    G5022_o2_p,
    G5022_o2
  );


  not

  (
    G5022_o2_n,
    G5022_o2
  );


  buf

  (
    G5006_o2_p,
    G5006_o2
  );


  not

  (
    G5006_o2_n,
    G5006_o2
  );


  buf

  (
    G4944_o2_p,
    G4944_o2
  );


  not

  (
    G4944_o2_n,
    G4944_o2
  );


  buf

  (
    G4946_o2_p,
    G4946_o2
  );


  not

  (
    G4946_o2_n,
    G4946_o2
  );


  buf

  (
    G4954_o2_p,
    G4954_o2
  );


  not

  (
    G4954_o2_n,
    G4954_o2
  );


  buf

  (
    G4956_o2_p,
    G4956_o2
  );


  not

  (
    G4956_o2_n,
    G4956_o2
  );


  buf

  (
    G3546_o2_p,
    G3546_o2
  );


  not

  (
    G3546_o2_n,
    G3546_o2
  );


  buf

  (
    G3658_o2_p,
    G3658_o2
  );


  not

  (
    G3658_o2_n,
    G3658_o2
  );


  buf

  (
    G1344_o2_p,
    G1344_o2
  );


  not

  (
    G1344_o2_n,
    G1344_o2
  );


  buf

  (
    G2921_o2_p,
    G2921_o2
  );


  not

  (
    G2921_o2_n,
    G2921_o2
  );


  buf

  (
    n3912_lo_buf_o2_p,
    n3912_lo_buf_o2
  );


  not

  (
    n3912_lo_buf_o2_n,
    n3912_lo_buf_o2
  );


  buf

  (
    G1835_o2_p,
    G1835_o2
  );


  not

  (
    G1835_o2_n,
    G1835_o2
  );


  buf

  (
    G3810_o2_p,
    G3810_o2
  );


  not

  (
    G3810_o2_n,
    G3810_o2
  );


  buf

  (
    G3866_o2_p,
    G3866_o2
  );


  not

  (
    G3866_o2_n,
    G3866_o2
  );


  buf

  (
    G3811_o2_p,
    G3811_o2
  );


  not

  (
    G3811_o2_n,
    G3811_o2
  );


  buf

  (
    G2269_o2_p,
    G2269_o2
  );


  not

  (
    G2269_o2_n,
    G2269_o2
  );


  buf

  (
    G3812_o2_p,
    G3812_o2
  );


  not

  (
    G3812_o2_n,
    G3812_o2
  );


  buf

  (
    G3867_o2_p,
    G3867_o2
  );


  not

  (
    G3867_o2_n,
    G3867_o2
  );


  buf

  (
    G3868_o2_p,
    G3868_o2
  );


  not

  (
    G3868_o2_n,
    G3868_o2
  );


  buf

  (
    G3809_o2_p,
    G3809_o2
  );


  not

  (
    G3809_o2_n,
    G3809_o2
  );


  buf

  (
    G3716_o2_p,
    G3716_o2
  );


  not

  (
    G3716_o2_n,
    G3716_o2
  );


  buf

  (
    G4529_o2_p,
    G4529_o2
  );


  not

  (
    G4529_o2_n,
    G4529_o2
  );


  buf

  (
    G4670_o2_p,
    G4670_o2
  );


  not

  (
    G4670_o2_n,
    G4670_o2
  );


  buf

  (
    G4493_o2_p,
    G4493_o2
  );


  not

  (
    G4493_o2_n,
    G4493_o2
  );


  buf

  (
    G4580_o2_p,
    G4580_o2
  );


  not

  (
    G4580_o2_n,
    G4580_o2
  );


  buf

  (
    G3822_o2_p,
    G3822_o2
  );


  not

  (
    G3822_o2_n,
    G3822_o2
  );


  buf

  (
    G3877_o2_p,
    G3877_o2
  );


  not

  (
    G3877_o2_n,
    G3877_o2
  );


  buf

  (
    G4131_o2_p,
    G4131_o2
  );


  not

  (
    G4131_o2_n,
    G4131_o2
  );


  buf

  (
    G4170_o2_p,
    G4170_o2
  );


  not

  (
    G4170_o2_n,
    G4170_o2
  );


  buf

  (
    G4051_o2_p,
    G4051_o2
  );


  not

  (
    G4051_o2_n,
    G4051_o2
  );


  buf

  (
    G4065_o2_p,
    G4065_o2
  );


  not

  (
    G4065_o2_n,
    G4065_o2
  );


  buf

  (
    G4697_o2_p,
    G4697_o2
  );


  not

  (
    G4697_o2_n,
    G4697_o2
  );


  buf

  (
    G4706_o2_p,
    G4706_o2
  );


  not

  (
    G4706_o2_n,
    G4706_o2
  );


  buf

  (
    G2460_o2_p,
    G2460_o2
  );


  not

  (
    G2460_o2_n,
    G2460_o2
  );


  buf

  (
    G2454_o2_p,
    G2454_o2
  );


  not

  (
    G2454_o2_n,
    G2454_o2
  );


  buf

  (
    G2392_o2_p,
    G2392_o2
  );


  not

  (
    G2392_o2_n,
    G2392_o2
  );


  buf

  (
    G2386_o2_p,
    G2386_o2
  );


  not

  (
    G2386_o2_n,
    G2386_o2
  );


  buf

  (
    n4260_lo_buf_o2_p,
    n4260_lo_buf_o2
  );


  not

  (
    n4260_lo_buf_o2_n,
    n4260_lo_buf_o2
  );


  buf

  (
    n4272_lo_buf_o2_p,
    n4272_lo_buf_o2
  );


  not

  (
    n4272_lo_buf_o2_n,
    n4272_lo_buf_o2
  );


  buf

  (
    n4392_lo_buf_o2_p,
    n4392_lo_buf_o2
  );


  not

  (
    n4392_lo_buf_o2_n,
    n4392_lo_buf_o2
  );


  buf

  (
    n4404_lo_buf_o2_p,
    n4404_lo_buf_o2
  );


  not

  (
    n4404_lo_buf_o2_n,
    n4404_lo_buf_o2
  );


  buf

  (
    G1512_o2_p,
    G1512_o2
  );


  not

  (
    G1512_o2_n,
    G1512_o2
  );


  buf

  (
    G3135_o2_p,
    G3135_o2
  );


  not

  (
    G3135_o2_n,
    G3135_o2
  );


  buf

  (
    G2379_o2_p,
    G2379_o2
  );


  not

  (
    G2379_o2_n,
    G2379_o2
  );


  buf

  (
    n4164_lo_buf_o2_p,
    n4164_lo_buf_o2
  );


  not

  (
    n4164_lo_buf_o2_n,
    n4164_lo_buf_o2
  );


  buf

  (
    n4176_lo_buf_o2_p,
    n4176_lo_buf_o2
  );


  not

  (
    n4176_lo_buf_o2_n,
    n4176_lo_buf_o2
  );


  buf

  (
    n4224_lo_buf_o2_p,
    n4224_lo_buf_o2
  );


  not

  (
    n4224_lo_buf_o2_n,
    n4224_lo_buf_o2
  );


  buf

  (
    G2975_o2_p,
    G2975_o2
  );


  not

  (
    G2975_o2_n,
    G2975_o2
  );


  buf

  (
    G2978_o2_p,
    G2978_o2
  );


  not

  (
    G2978_o2_n,
    G2978_o2
  );


  buf

  (
    G2933_o2_p,
    G2933_o2
  );


  not

  (
    G2933_o2_n,
    G2933_o2
  );


  buf

  (
    G2936_o2_p,
    G2936_o2
  );


  not

  (
    G2936_o2_n,
    G2936_o2
  );


  buf

  (
    G1356_o2_p,
    G1356_o2
  );


  not

  (
    G1356_o2_n,
    G1356_o2
  );


  buf

  (
    G1359_o2_p,
    G1359_o2
  );


  not

  (
    G1359_o2_n,
    G1359_o2
  );


  buf

  (
    G1398_o2_p,
    G1398_o2
  );


  not

  (
    G1398_o2_n,
    G1398_o2
  );


  buf

  (
    G1401_o2_p,
    G1401_o2
  );


  not

  (
    G1401_o2_n,
    G1401_o2
  );


  and

  (
    g1192_p,
    n4479_lo_p,
    n4443_lo_p
  );


  and

  (
    g1193_p,
    n3411_lo_p,
    n3399_lo_p_spl_
  );


  and

  (
    g1194_p,
    n4215_lo_p,
    n2619_lo_p_spl_
  );


  and

  (
    g1195_p,
    n4587_lo_n_spl_,
    n3363_lo_p
  );


  or

  (
    g1196_n,
    n4575_lo_p,
    n2739_lo_n_spl_
  );


  or

  (
    g1197_n,
    n4455_lo_n_spl_,
    n4239_lo_n_spl_
  );


  and

  (
    g1198_p,
    n2751_lo_p,
    n2739_lo_p
  );


  or

  (
    g1198_n,
    n2751_lo_n,
    n2739_lo_n_spl_
  );


  or

  (
    g1199_n,
    g1198_n_spl_000,
    n3387_lo_n
  );


  or

  (
    g1200_n,
    n4563_lo_n_spl_00,
    n3015_lo_n
  );


  or

  (
    g1201_n,
    n4563_lo_p_spl_00,
    n3003_lo_n
  );


  and

  (
    g1202_p,
    g1201_n,
    g1200_n
  );


  or

  (
    g1203_n,
    g1202_p,
    g1198_n_spl_000
  );


  or

  (
    g1204_n,
    n4563_lo_n_spl_00,
    n2763_lo_n
  );


  or

  (
    g1205_n,
    n4563_lo_p_spl_00,
    n3027_lo_n
  );


  and

  (
    g1206_p,
    g1205_n,
    g1204_n
  );


  or

  (
    g1207_n,
    g1206_p,
    g1198_n_spl_001
  );


  or

  (
    g1208_n,
    n4563_lo_n_spl_01,
    n2991_lo_n_spl_
  );


  or

  (
    g1209_n,
    n4563_lo_p_spl_01,
    n2991_lo_n_spl_
  );


  and

  (
    g1210_p,
    g1209_n,
    g1208_n
  );


  or

  (
    g1211_n,
    g1210_p,
    g1198_n_spl_001
  );


  or

  (
    g1212_n,
    n4563_lo_n_spl_01,
    n2703_lo_n
  );


  or

  (
    g1213_n,
    g1212_n,
    g1198_n_spl_010
  );


  or

  (
    g1214_n,
    n4563_lo_p_spl_01,
    n2715_lo_n
  );


  or

  (
    g1215_n,
    g1214_n,
    g1198_n_spl_010
  );


  or

  (
    g1216_n,
    g1198_p_spl_,
    n4563_lo_n_spl_10
  );


  or

  (
    g1217_n,
    g1198_p_spl_,
    n4563_lo_p_spl_10
  );


  and

  (
    g1218_p,
    g1215_n,
    g1213_n
  );


  and

  (
    g1219_p,
    g1218_p,
    g1216_n_spl_0
  );


  and

  (
    g1220_p,
    g1219_p,
    g1217_n_spl_0
  );


  or

  (
    g1221_n,
    g1220_p,
    n3399_lo_n_spl_00
  );


  or

  (
    g1222_n,
    n4563_lo_n_spl_10,
    n2727_lo_n
  );


  or

  (
    g1223_n,
    g1222_n,
    g1198_n_spl_011
  );


  or

  (
    g1224_n,
    n4563_lo_p_spl_10,
    n2967_lo_n
  );


  or

  (
    g1225_n,
    g1224_n,
    g1198_n_spl_011
  );


  and

  (
    g1226_p,
    g1225_n,
    g1223_n
  );


  and

  (
    g1227_p,
    g1226_p,
    g1216_n_spl_0
  );


  and

  (
    g1228_p,
    g1227_p,
    g1217_n_spl_0
  );


  or

  (
    g1229_n,
    g1228_p,
    n3399_lo_n_spl_00
  );


  or

  (
    g1230_n,
    n4563_lo_n_spl_11,
    n2943_lo_n
  );


  or

  (
    g1231_n,
    g1230_n,
    g1198_n_spl_100
  );


  or

  (
    g1232_n,
    n4563_lo_p_spl_11,
    n2691_lo_n
  );


  or

  (
    g1233_n,
    g1232_n,
    g1198_n_spl_100
  );


  and

  (
    g1234_p,
    g1233_n,
    g1231_n
  );


  and

  (
    g1235_p,
    g1234_p,
    g1216_n_spl_1
  );


  and

  (
    g1236_p,
    g1235_p,
    g1217_n_spl_1
  );


  or

  (
    g1237_n,
    g1236_p,
    n3399_lo_n_spl_0
  );


  or

  (
    g1238_n,
    n4563_lo_n_spl_11,
    n2979_lo_n
  );


  or

  (
    g1239_n,
    g1238_n,
    g1198_n_spl_10
  );


  or

  (
    g1240_n,
    n4563_lo_p_spl_11,
    n2955_lo_n
  );


  or

  (
    g1241_n,
    g1240_n,
    g1198_n_spl_11
  );


  and

  (
    g1242_p,
    g1241_n,
    g1239_n
  );


  and

  (
    g1243_p,
    g1242_p,
    g1216_n_spl_1
  );


  and

  (
    g1244_p,
    g1243_p,
    g1217_n_spl_1
  );


  or

  (
    g1245_n,
    g1244_p,
    n3399_lo_n_spl_1
  );


  or

  (
    g1246_n,
    n7357_o2_p_spl_0,
    n4359_lo_n_spl_
  );


  or

  (
    g1247_n,
    g1246_n,
    n4035_lo_p_spl_
  );


  or

  (
    g1248_n,
    n7359_o2_p_spl_0,
    n4359_lo_n_spl_
  );


  or

  (
    g1249_n,
    g1248_n,
    n4035_lo_n_spl_
  );


  and

  (
    g1250_p,
    g1249_n,
    g1247_n
  );


  and

  (
    g1251_p,
    n7449_o2_n_spl_0,
    n4035_lo_n_spl_
  );


  and

  (
    g1252_p,
    n7452_o2_n_spl_0,
    n4035_lo_p_spl_
  );


  or

  (
    g1253_n,
    g1252_p,
    g1251_p
  );


  or

  (
    g1254_n,
    g1253_n,
    n4359_lo_p
  );


  and

  (
    g1255_p,
    g1254_n,
    g1250_p
  );


  or

  (
    g1256_n,
    n7357_o2_p_spl_0,
    n4347_lo_n_spl_
  );


  or

  (
    g1257_n,
    g1256_n,
    n4011_lo_p_spl_
  );


  or

  (
    g1258_n,
    n7359_o2_p_spl_0,
    n4347_lo_n_spl_
  );


  or

  (
    g1259_n,
    g1258_n,
    n4011_lo_n_spl_
  );


  and

  (
    g1260_p,
    g1259_n,
    g1257_n
  );


  and

  (
    g1261_p,
    n7449_o2_n_spl_0,
    n4011_lo_n_spl_
  );


  and

  (
    g1262_p,
    n7452_o2_n_spl_0,
    n4011_lo_p_spl_
  );


  or

  (
    g1263_n,
    g1262_p,
    g1261_p
  );


  or

  (
    g1264_n,
    g1263_n,
    n4347_lo_p
  );


  and

  (
    g1265_p,
    g1264_n,
    g1260_p
  );


  or

  (
    g1266_n,
    n7357_o2_p_spl_,
    n3987_lo_p
  );


  or

  (
    g1267_n,
    n7359_o2_p_spl_,
    n3987_lo_n
  );


  and

  (
    g1268_p,
    g1267_n,
    g1266_n
  );


  and

  (
    g1269_p,
    n7449_o2_n_spl_,
    n3963_lo_n_spl_0
  );


  or

  (
    g1269_n,
    n7449_o2_p,
    n3963_lo_p_spl_
  );


  and

  (
    g1270_p,
    n7452_o2_n_spl_,
    n3963_lo_p_spl_
  );


  or

  (
    g1270_n,
    n7452_o2_p,
    n3963_lo_n_spl_0
  );


  and

  (
    g1271_p,
    g1270_n,
    g1269_n
  );


  or

  (
    g1271_n,
    g1270_p,
    g1269_p
  );


  or

  (
    g1272_n,
    g1265_p_spl_,
    g1255_p_spl_
  );


  or

  (
    g1273_n,
    g1272_n,
    g1268_p_spl_
  );


  or

  (
    g1274_n,
    g1273_n,
    g1271_n
  );


  or

  (
    g1275_n,
    n4635_lo_p_spl_000,
    n4407_lo_n_spl_
  );


  or

  (
    g1276_n,
    g1275_n,
    n4143_lo_p_spl_
  );


  or

  (
    g1277_n,
    n4623_lo_p_spl_000,
    n4407_lo_n_spl_
  );


  or

  (
    g1278_n,
    g1277_n,
    n4143_lo_n_spl_
  );


  and

  (
    g1279_p,
    g1278_n,
    g1276_n
  );


  and

  (
    g1280_p,
    n4599_lo_n_spl_000,
    n4143_lo_n_spl_
  );


  and

  (
    g1281_p,
    n4611_lo_n_spl_000,
    n4143_lo_p_spl_
  );


  or

  (
    g1282_n,
    g1281_p,
    g1280_p
  );


  or

  (
    g1283_n,
    g1282_n,
    n4407_lo_p
  );


  and

  (
    g1284_p,
    g1283_n,
    g1279_p
  );


  or

  (
    g1285_n,
    n4635_lo_p_spl_000,
    n4395_lo_n_spl_
  );


  or

  (
    g1286_n,
    g1285_n,
    n4119_lo_p_spl_
  );


  or

  (
    g1287_n,
    n4623_lo_p_spl_000,
    n4395_lo_n_spl_
  );


  or

  (
    g1288_n,
    g1287_n,
    n4119_lo_n_spl_
  );


  and

  (
    g1289_p,
    g1288_n,
    g1286_n
  );


  and

  (
    g1290_p,
    n4599_lo_n_spl_000,
    n4119_lo_n_spl_
  );


  and

  (
    g1291_p,
    n4611_lo_n_spl_000,
    n4119_lo_p_spl_
  );


  or

  (
    g1292_n,
    g1291_p,
    g1290_p
  );


  or

  (
    g1293_n,
    g1292_n,
    n4395_lo_p
  );


  and

  (
    g1294_p,
    g1293_n,
    g1289_p
  );


  or

  (
    g1295_n,
    n4635_lo_p_spl_001,
    n4383_lo_n
  );


  or

  (
    g1296_n,
    n4599_lo_n_spl_001,
    n4383_lo_p
  );


  and

  (
    g1297_p,
    g1296_n,
    g1295_n
  );


  or

  (
    g1298_n,
    n4635_lo_p_spl_001,
    n4371_lo_n_spl_0
  );


  or

  (
    g1299_n,
    g1298_n,
    n4059_lo_p_spl_
  );


  or

  (
    g1300_n,
    n4623_lo_p_spl_001,
    n4371_lo_n_spl_0
  );


  or

  (
    g1301_n,
    g1300_n,
    n4059_lo_n_spl_
  );


  and

  (
    g1302_p,
    g1301_n,
    g1299_n
  );


  and

  (
    g1303_p,
    n4599_lo_n_spl_001,
    n4059_lo_n_spl_
  );


  and

  (
    g1304_p,
    n4611_lo_n_spl_001,
    n4059_lo_p_spl_
  );


  or

  (
    g1305_n,
    g1304_p,
    g1303_p
  );


  or

  (
    g1306_n,
    g1305_n,
    n4371_lo_p_spl_
  );


  and

  (
    g1307_p,
    g1306_n,
    g1302_p
  );


  or

  (
    g1308_n,
    g1294_p_spl_,
    g1284_p_spl_
  );


  or

  (
    g1309_n,
    g1308_n,
    g1297_p_spl_
  );


  or

  (
    g1310_n,
    g1309_n,
    g1307_p_spl_
  );


  or

  (
    g1311_n,
    g1310_n,
    g1274_n
  );


  or

  (
    g1312_n,
    g1311_n,
    G2508_o2_p
  );


  or

  (
    g1313_n,
    n4635_lo_p_spl_010,
    n4299_lo_n_spl_0
  );


  or

  (
    g1314_n,
    g1313_n,
    n3759_lo_p_spl_
  );


  or

  (
    g1315_n,
    n4623_lo_p_spl_001,
    n4299_lo_n_spl_0
  );


  or

  (
    g1316_n,
    g1315_n,
    n3759_lo_n_spl_
  );


  and

  (
    g1317_p,
    g1316_n,
    g1314_n
  );


  and

  (
    g1318_p,
    n4599_lo_n_spl_010,
    n3759_lo_n_spl_
  );


  and

  (
    g1319_p,
    n4611_lo_n_spl_001,
    n3759_lo_p_spl_
  );


  or

  (
    g1320_n,
    g1319_p,
    g1318_p
  );


  or

  (
    g1321_n,
    g1320_n,
    n4299_lo_p_spl_
  );


  and

  (
    g1322_p,
    g1321_n,
    g1317_p
  );


  or

  (
    g1323_n,
    n4635_lo_p_spl_010,
    n4287_lo_n_spl_
  );


  or

  (
    g1324_n,
    g1323_n,
    n3735_lo_p_spl_
  );


  or

  (
    g1325_n,
    n4623_lo_p_spl_010,
    n4287_lo_n_spl_
  );


  or

  (
    g1326_n,
    g1325_n,
    n3735_lo_n_spl_
  );


  and

  (
    g1327_p,
    g1326_n,
    g1324_n
  );


  and

  (
    g1328_p,
    n4599_lo_n_spl_010,
    n3735_lo_n_spl_
  );


  and

  (
    g1329_p,
    n4611_lo_n_spl_010,
    n3735_lo_p_spl_
  );


  or

  (
    g1330_n,
    g1329_p,
    g1328_p
  );


  or

  (
    g1331_n,
    g1330_n,
    n4287_lo_p
  );


  and

  (
    g1332_p,
    g1331_n,
    g1327_p
  );


  or

  (
    g1333_n,
    n4635_lo_p_spl_011,
    n4335_lo_n_spl_
  );


  or

  (
    g1334_n,
    g1333_n,
    n3711_lo_p_spl_
  );


  or

  (
    g1335_n,
    n4623_lo_p_spl_010,
    n4335_lo_n_spl_
  );


  or

  (
    g1336_n,
    g1335_n,
    n3711_lo_n_spl_
  );


  and

  (
    g1337_p,
    g1336_n,
    g1334_n
  );


  and

  (
    g1338_p,
    n4599_lo_n_spl_011,
    n3711_lo_n_spl_
  );


  and

  (
    g1339_p,
    n4611_lo_n_spl_010,
    n3711_lo_p_spl_
  );


  or

  (
    g1340_n,
    g1339_p,
    g1338_p
  );


  or

  (
    g1341_n,
    g1340_n,
    n4335_lo_p
  );


  and

  (
    g1342_p,
    g1341_n,
    g1337_p
  );


  or

  (
    g1343_n,
    n4635_lo_p_spl_011,
    n4323_lo_n_spl_
  );


  or

  (
    g1344_n,
    g1343_n,
    n3687_lo_p_spl_
  );


  or

  (
    g1345_n,
    n4623_lo_p_spl_01,
    n4323_lo_n_spl_
  );


  or

  (
    g1346_n,
    g1345_n,
    n3687_lo_n_spl_
  );


  and

  (
    g1347_p,
    g1346_n,
    g1344_n
  );


  and

  (
    g1348_p,
    n4599_lo_n_spl_011,
    n3687_lo_n_spl_
  );


  and

  (
    g1349_p,
    n4611_lo_n_spl_01,
    n3687_lo_p_spl_
  );


  or

  (
    g1350_n,
    g1349_p,
    g1348_p
  );


  or

  (
    g1351_n,
    g1350_n,
    n4323_lo_p
  );


  and

  (
    g1352_p,
    g1351_n,
    g1347_p
  );


  or

  (
    g1353_n,
    g1332_p_spl_,
    g1322_p_spl_
  );


  or

  (
    g1354_n,
    g1353_n,
    g1342_p_spl_
  );


  or

  (
    g1355_n,
    g1354_n,
    g1352_p_spl_
  );


  or

  (
    g1356_n,
    n4635_lo_p_spl_10,
    n4227_lo_n_spl_
  );


  or

  (
    g1357_n,
    g1356_n,
    n3915_lo_p_spl_
  );


  or

  (
    g1358_n,
    n4623_lo_p_spl_10,
    n4227_lo_n_spl_
  );


  or

  (
    g1359_n,
    g1358_n,
    n3915_lo_n_spl_
  );


  and

  (
    g1360_p,
    g1359_n,
    g1357_n
  );


  and

  (
    g1361_p,
    n4599_lo_n_spl_10,
    n3915_lo_n_spl_
  );


  and

  (
    g1362_p,
    n4611_lo_n_spl_10,
    n3915_lo_p_spl_
  );


  or

  (
    g1363_n,
    g1362_p,
    g1361_p
  );


  or

  (
    g1364_n,
    g1363_n,
    n4227_lo_p
  );


  and

  (
    g1365_p,
    g1364_n,
    g1360_p
  );


  or

  (
    g1366_n,
    n4635_lo_p_spl_10,
    n4275_lo_n_spl_
  );


  or

  (
    g1367_n,
    g1366_n,
    n3891_lo_p_spl_
  );


  or

  (
    g1368_n,
    n4623_lo_p_spl_10,
    n4275_lo_n_spl_
  );


  or

  (
    g1369_n,
    g1368_n,
    n3891_lo_n_spl_
  );


  and

  (
    g1370_p,
    g1369_n,
    g1367_n
  );


  and

  (
    g1371_p,
    n4599_lo_n_spl_10,
    n3891_lo_n_spl_
  );


  and

  (
    g1372_p,
    n4611_lo_n_spl_10,
    n3891_lo_p_spl_
  );


  or

  (
    g1373_n,
    g1372_p,
    g1371_p
  );


  or

  (
    g1374_n,
    g1373_n,
    n4275_lo_p
  );


  and

  (
    g1375_p,
    g1374_n,
    g1370_p
  );


  or

  (
    g1376_n,
    n4635_lo_p_spl_11,
    n4263_lo_n_spl_
  );


  or

  (
    g1377_n,
    g1376_n,
    n3867_lo_p_spl_
  );


  or

  (
    g1378_n,
    n4623_lo_p_spl_11,
    n4263_lo_n_spl_
  );


  or

  (
    g1379_n,
    g1378_n,
    n3867_lo_n_spl_
  );


  and

  (
    g1380_p,
    g1379_n,
    g1377_n
  );


  and

  (
    g1381_p,
    n4599_lo_n_spl_11,
    n3867_lo_n_spl_
  );


  and

  (
    g1382_p,
    n4611_lo_n_spl_11,
    n3867_lo_p_spl_
  );


  or

  (
    g1383_n,
    g1382_p,
    g1381_p
  );


  or

  (
    g1384_n,
    g1383_n,
    n4263_lo_p
  );


  and

  (
    g1385_p,
    g1384_n,
    g1380_p
  );


  or

  (
    g1386_n,
    n4635_lo_p_spl_11,
    n4251_lo_n_spl_
  );


  or

  (
    g1387_n,
    g1386_n,
    n3843_lo_p_spl_
  );


  or

  (
    g1388_n,
    n4623_lo_p_spl_11,
    n4251_lo_n_spl_
  );


  or

  (
    g1389_n,
    g1388_n,
    n3843_lo_n_spl_
  );


  and

  (
    g1390_p,
    g1389_n,
    g1387_n
  );


  and

  (
    g1391_p,
    n4599_lo_n_spl_11,
    n3843_lo_n_spl_
  );


  and

  (
    g1392_p,
    n4611_lo_n_spl_11,
    n3843_lo_p_spl_
  );


  or

  (
    g1393_n,
    g1392_p,
    g1391_p
  );


  or

  (
    g1394_n,
    g1393_n,
    n4251_lo_p
  );


  and

  (
    g1395_p,
    g1394_n,
    g1390_p
  );


  or

  (
    g1396_n,
    g1375_p_spl_,
    g1365_p_spl_
  );


  or

  (
    g1397_n,
    g1396_n,
    g1385_p_spl_
  );


  or

  (
    g1398_n,
    g1397_n,
    g1395_p_spl_
  );


  or

  (
    g1399_n,
    g1398_n,
    g1355_n
  );


  or

  (
    g1400_n,
    g1399_n,
    G3060_o2_n
  );


  or

  (
    g1401_n,
    n6448_o2_n,
    n6419_o2_n_spl_
  );


  or

  (
    g1402_n,
    g1401_n,
    n6613_o2_n_spl_0
  );


  or

  (
    g1403_n,
    g1402_n,
    G3467_o2_n_spl_0
  );


  or

  (
    g1404_n,
    g1403_n_spl_,
    G3802_o2_n
  );


  or

  (
    g1405_n,
    G3570_o2_n_spl_,
    G2759_o2_p_spl_0
  );


  or

  (
    g1406_n,
    g1405_n,
    G3559_o2_n_spl_0
  );


  or

  (
    g1407_n,
    g1406_n,
    G2752_o2_p_spl_00
  );


  and

  (
    g1408_p,
    G3303_o2_p_spl_000,
    G2797_o2_n_spl_0
  );


  or

  (
    g1408_n,
    G3303_o2_n_spl_000,
    G2797_o2_p_spl_0
  );


  and

  (
    g1409_p,
    g1408_p,
    G3583_o2_p_spl_00
  );


  or

  (
    g1409_n,
    g1408_n,
    G3583_o2_n_spl_00
  );


  and

  (
    g1410_p,
    g1409_p,
    G3576_o2_p_spl_00
  );


  or

  (
    g1410_n,
    g1409_n,
    G3576_o2_n_spl_00
  );


  and

  (
    g1411_p,
    g1410_p,
    G3594_o2_p_spl_00
  );


  or

  (
    g1411_n,
    g1410_n,
    G3594_o2_n_spl_00
  );


  or

  (
    g1412_n,
    g1411_n_spl_,
    g1407_n_spl_
  );


  or

  (
    g1413_n,
    n6449_o2_n,
    n6420_o2_n_spl_
  );


  or

  (
    g1414_n,
    g1413_n,
    n6614_o2_p_spl_0
  );


  or

  (
    g1415_n,
    g1414_n,
    G2810_o2_p_spl_0
  );


  or

  (
    g1416_n,
    g1415_n_spl_,
    G3859_o2_n
  );


  or

  (
    g1417_n,
    G3415_o2_n_spl_,
    G3393_o2_n_spl_0
  );


  or

  (
    g1418_n,
    g1417_n,
    G3404_o2_n_spl_0
  );


  or

  (
    g1419_n,
    g1418_n,
    G3386_o2_n_spl_00
  );


  and

  (
    g1420_p,
    G3428_o2_p_spl_000,
    G3459_o2_p_spl_0
  );


  or

  (
    g1420_n,
    G3428_o2_n_spl_000,
    G3459_o2_n_spl_0
  );


  and

  (
    g1421_p,
    g1420_p,
    G3438_o2_p_spl_00
  );


  or

  (
    g1421_n,
    g1420_n,
    G3438_o2_n_spl_00
  );


  and

  (
    g1422_p,
    g1421_p,
    G3421_o2_p_spl_00
  );


  or

  (
    g1422_n,
    g1421_n,
    G3421_o2_n_spl_00
  );


  and

  (
    g1423_p,
    g1422_p,
    G3449_o2_p_spl_00
  );


  or

  (
    g1423_n,
    g1422_n,
    G3449_o2_n_spl_00
  );


  or

  (
    g1424_n,
    g1423_n_spl_,
    g1419_n_spl_
  );


  and

  (
    g1425_p,
    G2067_o2_p,
    G1422_o2_n
  );


  or

  (
    g1425_n,
    G2067_o2_n,
    G1422_o2_p
  );


  and

  (
    g1426_p,
    G2068_o2_p,
    G1419_o2_n
  );


  or

  (
    g1426_n,
    G2068_o2_n,
    G1419_o2_p
  );


  and

  (
    g1427_p,
    g1426_n,
    g1425_n
  );


  or

  (
    g1427_n,
    g1426_p,
    g1425_p
  );


  and

  (
    g1428_p,
    G2069_o2_p,
    G1428_o2_n
  );


  or

  (
    g1428_n,
    G2069_o2_n,
    G1428_o2_p
  );


  and

  (
    g1429_p,
    G2070_o2_p,
    G1425_o2_n
  );


  or

  (
    g1429_n,
    G2070_o2_n,
    G1425_o2_p
  );


  and

  (
    g1430_p,
    g1429_n,
    g1428_n
  );


  or

  (
    g1430_n,
    g1429_p,
    g1428_p
  );


  and

  (
    g1431_p,
    g1430_p_spl_,
    g1427_n_spl_
  );


  or

  (
    g1431_n,
    g1430_n_spl_,
    g1427_p_spl_
  );


  and

  (
    g1432_p,
    g1430_n_spl_,
    g1427_p_spl_
  );


  or

  (
    g1432_n,
    g1430_p_spl_,
    g1427_n_spl_
  );


  and

  (
    g1433_p,
    g1432_n,
    g1431_n
  );


  or

  (
    g1433_n,
    g1432_p,
    g1431_p
  );


  and

  (
    g1434_p,
    G2139_o2_n,
    G2140_o2_n
  );


  or

  (
    g1434_n,
    G2139_o2_p,
    G2140_o2_p
  );


  and

  (
    g1435_p,
    G2141_o2_n,
    G2142_o2_n
  );


  or

  (
    g1435_n,
    G2141_o2_p,
    G2142_o2_p
  );


  and

  (
    g1436_p,
    g1435_p_spl_0,
    g1434_n_spl_0
  );


  or

  (
    g1436_n,
    g1435_n_spl_0,
    g1434_p_spl_0
  );


  and

  (
    g1437_p,
    g1436_p,
    G1147_o2_n_spl_0
  );


  or

  (
    g1437_n,
    g1436_n,
    G1147_o2_p_spl_0
  );


  and

  (
    g1438_p,
    g1435_p_spl_0,
    g1434_p_spl_0
  );


  or

  (
    g1438_n,
    g1435_n_spl_0,
    g1434_n_spl_0
  );


  and

  (
    g1439_p,
    g1438_p,
    G1147_o2_p_spl_0
  );


  or

  (
    g1439_n,
    g1438_n,
    G1147_o2_n_spl_0
  );


  and

  (
    g1440_p,
    g1439_n,
    g1437_n
  );


  or

  (
    g1440_n,
    g1439_p,
    g1437_p
  );


  and

  (
    g1441_p,
    g1435_n_spl_1,
    g1434_p_spl_1
  );


  or

  (
    g1441_n,
    g1435_p_spl_1,
    g1434_n_spl_1
  );


  and

  (
    g1442_p,
    g1441_p,
    G1147_o2_n_spl_1
  );


  or

  (
    g1442_n,
    g1441_n,
    G1147_o2_p_spl_1
  );


  and

  (
    g1443_p,
    g1435_n_spl_1,
    g1434_n_spl_1
  );


  or

  (
    g1443_n,
    g1435_p_spl_1,
    g1434_p_spl_1
  );


  and

  (
    g1444_p,
    g1443_p,
    G1147_o2_p_spl_1
  );


  or

  (
    g1444_n,
    g1443_n,
    G1147_o2_n_spl_1
  );


  and

  (
    g1445_p,
    g1444_n,
    g1442_n
  );


  or

  (
    g1445_n,
    g1444_p,
    g1442_p
  );


  and

  (
    g1446_p,
    g1445_p,
    g1440_p
  );


  or

  (
    g1446_n,
    g1445_n,
    g1440_n
  );


  and

  (
    g1447_p,
    g1446_p,
    g1433_n
  );


  and

  (
    g1448_p,
    g1446_n,
    g1433_p
  );


  or

  (
    g1449_n,
    g1448_p,
    g1447_p
  );


  and

  (
    g1450_p,
    G2071_o2_p,
    G1452_o2_n
  );


  or

  (
    g1450_n,
    G2071_o2_n,
    G1452_o2_p
  );


  and

  (
    g1451_p,
    G2072_o2_p,
    G1449_o2_n
  );


  or

  (
    g1451_n,
    G2072_o2_n,
    G1449_o2_p
  );


  and

  (
    g1452_p,
    g1451_n,
    g1450_n
  );


  or

  (
    g1452_n,
    g1451_p,
    g1450_p
  );


  and

  (
    g1453_p,
    G2361_o2_n,
    G1455_o2_n
  );


  or

  (
    g1453_n,
    G2361_o2_p,
    G1455_o2_p
  );


  and

  (
    g1454_p,
    G2076_o2_p,
    G2073_o2_p
  );


  or

  (
    g1454_n,
    G2076_o2_n,
    G2073_o2_n
  );


  and

  (
    g1455_p,
    g1454_n,
    g1453_n
  );


  or

  (
    g1455_n,
    g1454_p,
    g1453_p
  );


  and

  (
    g1456_p,
    g1455_p_spl_,
    g1452_n_spl_
  );


  or

  (
    g1456_n,
    g1455_n_spl_,
    g1452_p_spl_
  );


  and

  (
    g1457_p,
    g1455_n_spl_,
    g1452_p_spl_
  );


  or

  (
    g1457_n,
    g1455_p_spl_,
    g1452_n_spl_
  );


  and

  (
    g1458_p,
    g1457_n,
    g1456_n
  );


  or

  (
    g1458_n,
    g1457_p,
    g1456_p
  );


  and

  (
    g1459_p,
    G2143_o2_n,
    G2144_o2_n
  );


  or

  (
    g1459_n,
    G2143_o2_p,
    G2144_o2_p
  );


  and

  (
    g1460_p,
    G2145_o2_n,
    G2146_o2_n
  );


  or

  (
    g1460_n,
    G2145_o2_p,
    G2146_o2_p
  );


  and

  (
    g1461_p,
    g1460_p_spl_0,
    g1459_n_spl_0
  );


  or

  (
    g1461_n,
    g1460_n_spl_0,
    g1459_p_spl_0
  );


  and

  (
    g1462_p,
    g1461_p,
    G2336_o2_p_spl_0
  );


  or

  (
    g1462_n,
    g1461_n,
    G2336_o2_n_spl_0
  );


  and

  (
    g1463_p,
    g1460_p_spl_0,
    g1459_p_spl_0
  );


  or

  (
    g1463_n,
    g1460_n_spl_0,
    g1459_n_spl_0
  );


  and

  (
    g1464_p,
    g1463_p,
    G2336_o2_n_spl_0
  );


  or

  (
    g1464_n,
    g1463_n,
    G2336_o2_p_spl_0
  );


  and

  (
    g1465_p,
    g1464_n,
    g1462_n
  );


  or

  (
    g1465_n,
    g1464_p,
    g1462_p
  );


  and

  (
    g1466_p,
    g1460_n_spl_1,
    g1459_p_spl_1
  );


  or

  (
    g1466_n,
    g1460_p_spl_1,
    g1459_n_spl_1
  );


  and

  (
    g1467_p,
    g1466_p,
    G2336_o2_p_spl_1
  );


  or

  (
    g1467_n,
    g1466_n,
    G2336_o2_n_spl_1
  );


  and

  (
    g1468_p,
    g1460_n_spl_1,
    g1459_n_spl_1
  );


  or

  (
    g1468_n,
    g1460_p_spl_1,
    g1459_p_spl_1
  );


  and

  (
    g1469_p,
    g1468_p,
    G2336_o2_n_spl_1
  );


  or

  (
    g1469_n,
    g1468_n,
    G2336_o2_p_spl_1
  );


  and

  (
    g1470_p,
    g1469_n,
    g1467_n
  );


  or

  (
    g1470_n,
    g1469_p,
    g1467_p
  );


  and

  (
    g1471_p,
    g1470_p,
    g1465_p
  );


  or

  (
    g1471_n,
    g1470_n,
    g1465_n
  );


  and

  (
    g1472_p,
    g1471_p,
    g1458_n
  );


  and

  (
    g1473_p,
    g1471_n,
    g1458_p
  );


  or

  (
    g1474_n,
    g1473_p,
    g1472_p
  );


  or

  (
    g1475_n,
    n7116_o2_n,
    n4311_lo_n_spl_0
  );


  or

  (
    g1476_n,
    G3467_o2_n_spl_0,
    n6641_o2_n
  );


  or

  (
    g1477_n,
    G3467_o2_n_spl_1,
    n6613_o2_n_spl_0
  );


  or

  (
    g1478_n,
    g1477_n,
    n6435_o2_n
  );


  or

  (
    g1479_n,
    G3467_o2_n_spl_1,
    n6419_o2_n_spl_
  );


  or

  (
    g1480_n,
    g1479_n,
    n6382_o2_n
  );


  or

  (
    g1481_n,
    g1480_n,
    n6613_o2_n_spl_
  );


  and

  (
    g1482_p,
    g1476_n,
    g1475_n_spl_
  );


  and

  (
    g1483_p,
    g1482_p,
    g1478_n
  );


  and

  (
    g1484_p,
    g1483_p,
    g1481_n
  );


  or

  (
    g1485_n,
    g1403_n_spl_,
    G4054_o2_n
  );


  and

  (
    g1486_p,
    g1485_n,
    g1484_p
  );


  or

  (
    g1487_n,
    G2752_o2_p_spl_00,
    G2770_o2_p_spl_
  );


  or

  (
    g1488_n,
    G2752_o2_p_spl_01,
    G2759_o2_p_spl_0
  );


  or

  (
    g1489_n,
    g1488_n,
    G2774_o2_n_spl_
  );


  or

  (
    g1490_n,
    G2752_o2_p_spl_01,
    G3559_o2_n_spl_0
  );


  or

  (
    g1491_n,
    g1490_n,
    G2780_o2_n_spl_
  );


  or

  (
    g1492_n,
    g1491_n,
    G2759_o2_p_spl_1
  );


  and

  (
    g1493_p,
    g1487_n,
    n7463_o2_n_spl_0
  );


  and

  (
    g1494_p,
    g1493_p,
    g1489_n
  );


  and

  (
    g1495_p,
    g1494_p,
    g1492_n
  );


  and

  (
    g1496_p,
    n6756_o2_p,
    n4371_lo_p_spl_
  );


  or

  (
    g1496_n,
    n6756_o2_n,
    n4371_lo_n_spl_
  );


  and

  (
    g1497_p,
    G3576_o2_p_spl_00,
    G2540_o2_p_spl_
  );


  or

  (
    g1497_n,
    G3576_o2_n_spl_00,
    G2540_o2_n_spl_
  );


  and

  (
    g1498_p,
    G3303_o2_p_spl_000,
    G3576_o2_p_spl_01
  );


  or

  (
    g1498_n,
    G3303_o2_n_spl_000,
    G3576_o2_n_spl_01
  );


  and

  (
    g1499_p,
    g1498_p,
    G2788_o2_p_spl_0
  );


  or

  (
    g1499_n,
    g1498_n,
    G2788_o2_n_spl_0
  );


  and

  (
    g1500_p,
    G3583_o2_p_spl_00,
    G3576_o2_p_spl_01
  );


  or

  (
    g1500_n,
    G3583_o2_n_spl_00,
    G3576_o2_n_spl_01
  );


  and

  (
    g1501_p,
    g1500_p,
    G2792_o2_p_spl_0
  );


  or

  (
    g1501_n,
    g1500_n,
    G2792_o2_n_spl_0
  );


  and

  (
    g1502_p,
    g1501_p,
    G3303_o2_p_spl_00
  );


  or

  (
    g1502_n,
    g1501_n,
    G3303_o2_n_spl_00
  );


  and

  (
    g1503_p,
    G3594_o2_p_spl_00,
    G3583_o2_p_spl_01
  );


  or

  (
    g1503_n,
    G3594_o2_n_spl_00,
    G3583_o2_n_spl_01
  );


  and

  (
    g1504_p,
    g1503_p_spl_,
    G3576_o2_p_spl_1
  );


  or

  (
    g1504_n,
    g1503_n_spl_,
    G3576_o2_n_spl_1
  );


  and

  (
    g1505_p,
    g1504_p,
    G2804_o2_n_spl_0
  );


  or

  (
    g1505_n,
    g1504_n,
    G2804_o2_p_spl_0
  );


  and

  (
    g1506_p,
    g1505_p,
    G3303_o2_p_spl_01
  );


  or

  (
    g1506_n,
    g1505_n,
    G3303_o2_n_spl_01
  );


  and

  (
    g1507_p,
    g1497_n,
    g1496_n
  );


  or

  (
    g1507_n,
    g1497_p,
    g1496_p
  );


  and

  (
    g1508_p,
    g1507_p,
    g1499_n
  );


  or

  (
    g1508_n,
    g1507_n,
    g1499_p
  );


  and

  (
    g1509_p,
    g1508_p,
    g1502_n
  );


  or

  (
    g1509_n,
    g1508_n,
    g1502_p
  );


  and

  (
    g1510_p,
    g1509_p,
    g1506_n
  );


  or

  (
    g1510_n,
    g1509_n,
    g1506_p
  );


  or

  (
    g1511_n,
    g1510_p_spl_,
    g1407_n_spl_
  );


  and

  (
    g1512_p,
    g1511_n,
    g1495_p
  );


  or

  (
    g1513_n,
    G3386_o2_n_spl_00,
    G2675_o2_n_spl_
  );


  or

  (
    g1514_n,
    G3386_o2_n_spl_0,
    G3393_o2_n_spl_0
  );


  or

  (
    g1515_n,
    g1514_n,
    G2679_o2_n_spl_
  );


  or

  (
    g1516_n,
    G3386_o2_n_spl_1,
    G3404_o2_n_spl_0
  );


  or

  (
    g1517_n,
    g1516_n,
    G2685_o2_n_spl_
  );


  or

  (
    g1518_n,
    g1517_n,
    G3393_o2_n_spl_1
  );


  and

  (
    g1519_p,
    g1513_n,
    g1475_n_spl_
  );


  and

  (
    g1520_p,
    g1519_p,
    g1515_n
  );


  and

  (
    g1521_p,
    g1520_p,
    g1518_n
  );


  and

  (
    g1522_p,
    n6757_o2_p,
    n4299_lo_p_spl_
  );


  or

  (
    g1522_n,
    n6757_o2_n,
    n4299_lo_n_spl_
  );


  and

  (
    g1523_p,
    G3421_o2_p_spl_00,
    G2693_o2_p_spl_
  );


  or

  (
    g1523_n,
    G3421_o2_n_spl_00,
    G2693_o2_n_spl_
  );


  and

  (
    g1524_p,
    G3421_o2_p_spl_01,
    G3428_o2_p_spl_000
  );


  or

  (
    g1524_n,
    G3421_o2_n_spl_01,
    G3428_o2_n_spl_000
  );


  and

  (
    g1525_p,
    g1524_p,
    G2696_o2_p_spl_0
  );


  or

  (
    g1525_n,
    g1524_n,
    G2696_o2_n_spl_0
  );


  and

  (
    g1526_p,
    G3421_o2_p_spl_01,
    G3438_o2_p_spl_00
  );


  or

  (
    g1526_n,
    G3421_o2_n_spl_01,
    G3438_o2_n_spl_00
  );


  and

  (
    g1527_p,
    g1526_p,
    G2700_o2_p_spl_0
  );


  or

  (
    g1527_n,
    g1526_n,
    G2700_o2_n_spl_0
  );


  and

  (
    g1528_p,
    g1527_p,
    G3428_o2_p_spl_00
  );


  or

  (
    g1528_n,
    g1527_n,
    G3428_o2_n_spl_00
  );


  and

  (
    g1529_p,
    G3449_o2_p_spl_00,
    G3438_o2_p_spl_01
  );


  or

  (
    g1529_n,
    G3449_o2_n_spl_00,
    G3438_o2_n_spl_01
  );


  and

  (
    g1530_p,
    g1529_p_spl_,
    G3421_o2_p_spl_1
  );


  or

  (
    g1530_n,
    g1529_n_spl_,
    G3421_o2_n_spl_1
  );


  and

  (
    g1531_p,
    g1530_p,
    G2705_o2_p_spl_0
  );


  or

  (
    g1531_n,
    g1530_n,
    G2705_o2_n_spl_0
  );


  and

  (
    g1532_p,
    g1531_p,
    G3428_o2_p_spl_01
  );


  or

  (
    g1532_n,
    g1531_n,
    G3428_o2_n_spl_01
  );


  and

  (
    g1533_p,
    g1523_n,
    g1522_n
  );


  or

  (
    g1533_n,
    g1523_p,
    g1522_p
  );


  and

  (
    g1534_p,
    g1533_p,
    g1525_n
  );


  or

  (
    g1534_n,
    g1533_n,
    g1525_p
  );


  and

  (
    g1535_p,
    g1534_p,
    g1528_n
  );


  or

  (
    g1535_n,
    g1534_n,
    g1528_p
  );


  and

  (
    g1536_p,
    g1535_p,
    g1532_n
  );


  or

  (
    g1536_n,
    g1535_n,
    g1532_p
  );


  or

  (
    g1537_n,
    g1536_p_spl_,
    g1419_n_spl_
  );


  and

  (
    g1538_p,
    g1537_n,
    g1521_p
  );


  or

  (
    g1539_n,
    G2810_o2_p_spl_0,
    n6658_o2_p
  );


  or

  (
    g1540_n,
    G2810_o2_p_spl_1,
    n6614_o2_p_spl_0
  );


  or

  (
    g1541_n,
    g1540_n,
    n6436_o2_n
  );


  or

  (
    g1542_n,
    G2810_o2_p_spl_1,
    n6420_o2_n_spl_
  );


  or

  (
    g1543_n,
    g1542_n,
    n6383_o2_n
  );


  or

  (
    g1544_n,
    g1543_n,
    n6614_o2_p_spl_
  );


  and

  (
    g1545_p,
    g1539_n,
    n7463_o2_n_spl_0
  );


  and

  (
    g1546_p,
    g1545_p,
    g1541_n
  );


  and

  (
    g1547_p,
    g1546_p,
    g1544_n
  );


  or

  (
    g1548_n,
    g1415_n_spl_,
    G4068_o2_n
  );


  and

  (
    g1549_p,
    g1548_n,
    g1547_p
  );


  or

  (
    g1550_n,
    n7358_o2_p_spl_,
    n4167_lo_p
  );


  or

  (
    g1551_n,
    n7360_o2_p_spl_,
    n4167_lo_n
  );


  and

  (
    g1552_p,
    g1551_n,
    g1550_n
  );


  and

  (
    g1553_p,
    g1552_p,
    n4719_lo_p_spl_00000
  );


  and

  (
    g1554_p,
    g1553_p,
    n4731_lo_p_spl_00000
  );


  and

  (
    g1555_p,
    G2797_o2_p_spl_0,
    n2859_lo_p_spl_0
  );


  and

  (
    g1556_p,
    G2797_o2_n_spl_0,
    n2859_lo_n_spl_0
  );


  or

  (
    g1557_n,
    g1556_p,
    g1555_p
  );


  and

  (
    g1558_p,
    g1557_n_spl_,
    n4719_lo_n_spl_0000
  );


  and

  (
    g1559_p,
    g1558_p,
    n4731_lo_p_spl_00000
  );


  and

  (
    g1560_p,
    n4719_lo_p_spl_00000,
    n3327_lo_p
  );


  and

  (
    g1561_p,
    g1560_p,
    n4731_lo_n_spl_0000
  );


  or

  (
    g1562_n,
    g1559_p,
    g1554_p
  );


  or

  (
    g1563_n,
    g1562_n,
    g1561_p
  );


  and

  (
    g1564_p,
    g1284_p_spl_,
    n4719_lo_p_spl_00001
  );


  and

  (
    g1565_p,
    g1564_p,
    n4731_lo_p_spl_00001
  );


  and

  (
    g1566_p,
    G2797_o2_n_spl_,
    n2859_lo_p_spl_0
  );


  or

  (
    g1566_n,
    G2797_o2_p_spl_,
    n2859_lo_n_spl_0
  );


  and

  (
    g1567_p,
    g1566_n_spl_0,
    G2804_o2_p_spl_0
  );


  or

  (
    g1567_n,
    g1566_p_spl_0,
    G2804_o2_n_spl_0
  );


  and

  (
    g1568_p,
    g1567_p,
    G3594_o2_n_spl_01
  );


  and

  (
    g1569_p,
    g1567_n,
    G3594_o2_p_spl_01
  );


  or

  (
    g1570_n,
    g1569_p,
    g1568_p
  );


  and

  (
    g1571_p,
    g1570_n_spl_,
    n4719_lo_n_spl_0000
  );


  and

  (
    g1572_p,
    g1571_p,
    n4731_lo_p_spl_00001
  );


  and

  (
    g1573_p,
    n4719_lo_p_spl_00001,
    n3303_lo_p
  );


  and

  (
    g1574_p,
    g1573_p,
    n4731_lo_n_spl_0000
  );


  or

  (
    g1575_n,
    g1572_p,
    g1565_p
  );


  or

  (
    g1576_n,
    g1575_n,
    g1574_p
  );


  and

  (
    g1577_p,
    g1365_p_spl_,
    n4719_lo_p_spl_00010
  );


  and

  (
    g1578_p,
    g1577_p,
    n4731_lo_p_spl_00010
  );


  and

  (
    g1579_p,
    G3459_o2_n_spl_0,
    n2631_lo_p_spl_0
  );


  and

  (
    g1580_p,
    G3459_o2_p_spl_0,
    n2631_lo_n_spl_0
  );


  or

  (
    g1581_n,
    g1580_p,
    g1579_p
  );


  and

  (
    g1582_p,
    g1581_n_spl_,
    n4719_lo_n_spl_0001
  );


  and

  (
    g1583_p,
    g1582_p,
    n4731_lo_p_spl_00010
  );


  and

  (
    g1584_p,
    n4719_lo_p_spl_00010,
    n3183_lo_p
  );


  and

  (
    g1585_p,
    g1584_p,
    n4731_lo_n_spl_0001
  );


  or

  (
    g1586_n,
    g1583_p,
    g1578_p
  );


  or

  (
    g1587_n,
    g1586_n,
    g1585_p
  );


  and

  (
    g1588_p,
    G3228_o2_p_spl_,
    G4137_o2_n_spl_
  );


  or

  (
    g1588_n,
    G3228_o2_n_spl_,
    G4137_o2_p_spl_
  );


  and

  (
    g1589_p,
    G3228_o2_n_spl_,
    G4137_o2_p_spl_
  );


  or

  (
    g1589_n,
    G3228_o2_p_spl_,
    G4137_o2_n_spl_
  );


  and

  (
    g1590_p,
    g1589_n,
    g1588_n
  );


  or

  (
    g1590_n,
    g1589_p,
    g1588_p
  );


  and

  (
    g1591_p,
    g1411_p,
    n2859_lo_p_spl_
  );


  or

  (
    g1591_n,
    g1411_n_spl_,
    n2859_lo_n_spl_
  );


  and

  (
    g1592_p,
    g1591_n,
    g1510_p_spl_
  );


  or

  (
    g1592_n,
    g1591_p,
    g1510_n
  );


  and

  (
    g1593_p,
    g1592_p_spl_00,
    g1590_p
  );


  or

  (
    g1593_n,
    g1592_n_spl_00,
    g1590_n
  );


  and

  (
    g1594_p,
    G3161_o2_n,
    G2770_o2_p_spl_
  );


  or

  (
    g1594_n,
    G3161_o2_p,
    G2770_o2_n
  );


  and

  (
    g1595_p,
    g1594_p,
    G3828_o2_n
  );


  or

  (
    g1595_n,
    g1594_n,
    G3828_o2_p
  );


  and

  (
    g1596_p,
    g1595_p,
    G3829_o2_n
  );


  or

  (
    g1596_n,
    g1595_n,
    G3829_o2_p
  );


  and

  (
    g1597_p,
    g1596_p_spl_,
    G2752_o2_p_spl_1
  );


  or

  (
    g1597_n,
    g1596_n_spl_,
    G2752_o2_n_spl_
  );


  and

  (
    g1598_p,
    g1596_n_spl_,
    G2752_o2_n_spl_
  );


  or

  (
    g1598_n,
    g1596_p_spl_,
    G2752_o2_p_spl_1
  );


  and

  (
    g1599_p,
    g1598_n,
    g1597_n
  );


  or

  (
    g1599_n,
    g1598_p,
    g1597_p
  );


  and

  (
    g1600_p,
    g1599_n,
    g1592_n_spl_00
  );


  or

  (
    g1600_n,
    g1599_p,
    g1592_p_spl_00
  );


  and

  (
    g1601_p,
    g1600_n,
    g1593_n
  );


  or

  (
    g1601_n,
    g1600_p,
    g1593_p
  );


  and

  (
    g1602_p,
    g1563_n_spl_00,
    n4683_lo_p_spl_0000
  );


  and

  (
    g1603_p,
    g1602_p,
    n4671_lo_p_spl_0000
  );


  and

  (
    g1604_p,
    g1587_n_spl_00,
    n4683_lo_n_spl_0000
  );


  and

  (
    g1605_p,
    g1604_p,
    n4671_lo_p_spl_0000
  );


  and

  (
    g1606_p,
    n4683_lo_p_spl_0000,
    n2643_lo_p_spl_
  );


  and

  (
    g1607_p,
    g1606_p,
    n4671_lo_n_spl_0000
  );


  and

  (
    g1608_p,
    n4683_lo_n_spl_0000,
    n2871_lo_p_spl_
  );


  and

  (
    g1609_p,
    g1608_p,
    n4671_lo_n_spl_0000
  );


  or

  (
    g1610_n,
    g1605_p,
    g1603_p
  );


  or

  (
    g1611_n,
    g1610_n,
    g1607_p
  );


  or

  (
    g1612_n,
    g1611_n,
    g1609_p
  );


  and

  (
    g1613_p,
    g1307_p_spl_,
    n4719_lo_p_spl_00011
  );


  and

  (
    g1614_p,
    g1613_p,
    n4731_lo_p_spl_00011
  );


  and

  (
    g1615_p,
    G3303_o2_p_spl_01,
    G2788_o2_p_spl_0
  );


  or

  (
    g1615_n,
    G3303_o2_n_spl_01,
    G2788_o2_n_spl_0
  );


  and

  (
    g1616_p,
    G3583_o2_p_spl_01,
    G2792_o2_p_spl_0
  );


  or

  (
    g1616_n,
    G3583_o2_n_spl_01,
    G2792_o2_n_spl_0
  );


  and

  (
    g1617_p,
    g1616_p_spl_,
    G3303_o2_p_spl_10
  );


  or

  (
    g1617_n,
    g1616_n_spl_,
    G3303_o2_n_spl_10
  );


  and

  (
    g1618_p,
    g1503_p_spl_,
    G2804_o2_n_spl_1
  );


  or

  (
    g1618_n,
    g1503_n_spl_,
    G2804_o2_p_spl_1
  );


  and

  (
    g1619_p,
    g1618_p_spl_,
    G3303_o2_p_spl_10
  );


  or

  (
    g1619_n,
    g1618_n_spl_,
    G3303_o2_n_spl_10
  );


  and

  (
    g1620_p,
    g1566_p_spl_0,
    G3583_o2_p_spl_1
  );


  or

  (
    g1620_n,
    g1566_n_spl_0,
    G3583_o2_n_spl_1
  );


  and

  (
    g1621_p,
    g1620_p,
    G3594_o2_p_spl_01
  );


  or

  (
    g1621_n,
    g1620_n,
    G3594_o2_n_spl_01
  );


  and

  (
    g1622_p,
    g1621_p_spl_,
    G3303_o2_p_spl_11
  );


  or

  (
    g1622_n,
    g1621_n_spl_,
    G3303_o2_n_spl_11
  );


  and

  (
    g1623_p,
    g1615_n,
    G2540_o2_n_spl_
  );


  or

  (
    g1623_n,
    g1615_p,
    G2540_o2_p_spl_
  );


  and

  (
    g1624_p,
    g1623_p,
    g1617_n
  );


  or

  (
    g1624_n,
    g1623_n,
    g1617_p
  );


  and

  (
    g1625_p,
    g1624_p,
    g1619_n
  );


  or

  (
    g1625_n,
    g1624_n,
    g1619_p
  );


  and

  (
    g1626_p,
    g1625_p,
    g1622_n
  );


  or

  (
    g1626_n,
    g1625_n,
    g1622_p
  );


  and

  (
    g1627_p,
    g1626_p,
    G3576_o2_n_spl_1
  );


  and

  (
    g1628_p,
    g1626_n,
    G3576_o2_p_spl_1
  );


  or

  (
    g1629_n,
    g1628_p,
    g1627_p
  );


  and

  (
    g1630_p,
    g1629_n_spl_,
    n4719_lo_n_spl_0001
  );


  and

  (
    g1631_p,
    g1630_p,
    n4731_lo_p_spl_00011
  );


  and

  (
    g1632_p,
    n4719_lo_p_spl_00011,
    n2835_lo_p
  );


  and

  (
    g1633_p,
    g1632_p,
    n4731_lo_n_spl_0001
  );


  or

  (
    g1634_n,
    g1631_p,
    g1614_p
  );


  or

  (
    g1635_n,
    g1634_n,
    g1633_p
  );


  and

  (
    g1636_p,
    g1297_p_spl_,
    n4719_lo_p_spl_00100
  );


  and

  (
    g1637_p,
    g1636_p,
    n4731_lo_p_spl_00100
  );


  and

  (
    g1638_p,
    g1616_n_spl_,
    G2788_o2_n_spl_
  );


  or

  (
    g1638_n,
    g1616_p_spl_,
    G2788_o2_p_spl_
  );


  and

  (
    g1639_p,
    g1638_p,
    g1618_n_spl_
  );


  or

  (
    g1639_n,
    g1638_n,
    g1618_p_spl_
  );


  and

  (
    g1640_p,
    g1639_p,
    g1621_n_spl_
  );


  or

  (
    g1640_n,
    g1639_n,
    g1621_p_spl_
  );


  and

  (
    g1641_p,
    g1640_p,
    G3303_o2_n_spl_11
  );


  and

  (
    g1642_p,
    g1640_n,
    G3303_o2_p_spl_11
  );


  or

  (
    g1643_n,
    g1642_p,
    g1641_p
  );


  and

  (
    g1644_p,
    g1643_n_spl_,
    n4719_lo_n_spl_0010
  );


  and

  (
    g1645_p,
    g1644_p,
    n4731_lo_p_spl_00100
  );


  and

  (
    g1646_p,
    n4719_lo_p_spl_00100,
    n3315_lo_p
  );


  and

  (
    g1647_p,
    g1646_p,
    n4731_lo_n_spl_0010
  );


  or

  (
    g1648_n,
    g1645_p,
    g1637_p
  );


  or

  (
    g1649_n,
    g1648_n,
    g1647_p
  );


  and

  (
    g1650_p,
    g1294_p_spl_,
    n4719_lo_p_spl_00101
  );


  and

  (
    g1651_p,
    g1650_p,
    n4731_lo_p_spl_00101
  );


  and

  (
    g1652_p,
    G3594_o2_p_spl_1,
    G2804_o2_n_spl_1
  );


  or

  (
    g1652_n,
    G3594_o2_n_spl_1,
    G2804_o2_p_spl_1
  );


  and

  (
    g1653_p,
    g1566_p_spl_,
    G3594_o2_p_spl_1
  );


  or

  (
    g1653_n,
    g1566_n_spl_,
    G3594_o2_n_spl_1
  );


  and

  (
    g1654_p,
    g1652_n,
    G2792_o2_n_spl_
  );


  or

  (
    g1654_n,
    g1652_p,
    G2792_o2_p_spl_
  );


  and

  (
    g1655_p,
    g1654_p,
    g1653_n
  );


  or

  (
    g1655_n,
    g1654_n,
    g1653_p
  );


  and

  (
    g1656_p,
    g1655_p,
    G3583_o2_n_spl_1
  );


  and

  (
    g1657_p,
    g1655_n,
    G3583_o2_p_spl_1
  );


  or

  (
    g1658_n,
    g1657_p,
    g1656_p
  );


  and

  (
    g1659_p,
    g1658_n_spl_,
    n4719_lo_n_spl_0010
  );


  and

  (
    g1660_p,
    g1659_p,
    n4731_lo_p_spl_00101
  );


  and

  (
    g1661_p,
    n4719_lo_p_spl_00101,
    n3207_lo_p
  );


  and

  (
    g1662_p,
    g1661_p,
    n4731_lo_n_spl_0010
  );


  or

  (
    g1663_n,
    g1660_p,
    g1651_p
  );


  or

  (
    g1664_n,
    g1663_n,
    g1662_p
  );


  and

  (
    g1665_p,
    g1563_n_spl_00,
    n4695_lo_p_spl_0000
  );


  and

  (
    g1666_p,
    g1665_p,
    n4707_lo_p_spl_0000
  );


  and

  (
    g1667_p,
    g1587_n_spl_00,
    n4695_lo_n_spl_0000
  );


  and

  (
    g1668_p,
    g1667_p,
    n4707_lo_p_spl_0000
  );


  and

  (
    g1669_p,
    n4695_lo_p_spl_0000,
    n2643_lo_p_spl_
  );


  and

  (
    g1670_p,
    g1669_p,
    n4707_lo_n_spl_0000
  );


  and

  (
    g1671_p,
    n4695_lo_n_spl_0000,
    n2871_lo_p_spl_
  );


  and

  (
    g1672_p,
    g1671_p,
    n4707_lo_n_spl_0000
  );


  or

  (
    g1673_n,
    g1668_p,
    g1666_p
  );


  or

  (
    g1674_n,
    g1673_n,
    g1670_p
  );


  or

  (
    g1675_n,
    g1674_n,
    g1672_p
  );


  and

  (
    g1676_p,
    g1322_p_spl_,
    n4719_lo_p_spl_00110
  );


  and

  (
    g1677_p,
    g1676_p,
    n4731_lo_p_spl_00110
  );


  and

  (
    g1678_p,
    G3428_o2_p_spl_01,
    G2696_o2_p_spl_0
  );


  or

  (
    g1678_n,
    G3428_o2_n_spl_01,
    G2696_o2_n_spl_0
  );


  and

  (
    g1679_p,
    G3438_o2_p_spl_01,
    G2700_o2_p_spl_0
  );


  or

  (
    g1679_n,
    G3438_o2_n_spl_01,
    G2700_o2_n_spl_0
  );


  and

  (
    g1680_p,
    g1679_p_spl_,
    G3428_o2_p_spl_10
  );


  or

  (
    g1680_n,
    g1679_n_spl_,
    G3428_o2_n_spl_10
  );


  and

  (
    g1681_p,
    g1529_p_spl_,
    G2705_o2_p_spl_0
  );


  or

  (
    g1681_n,
    g1529_n_spl_,
    G2705_o2_n_spl_0
  );


  and

  (
    g1682_p,
    g1681_p_spl_,
    G3428_o2_p_spl_10
  );


  or

  (
    g1682_n,
    g1681_n_spl_,
    G3428_o2_n_spl_10
  );


  and

  (
    g1683_p,
    G3459_o2_p_spl_,
    n2631_lo_p_spl_0
  );


  or

  (
    g1683_n,
    G3459_o2_n_spl_,
    n2631_lo_n_spl_0
  );


  and

  (
    g1684_p,
    g1683_p_spl_0,
    G3438_o2_p_spl_1
  );


  or

  (
    g1684_n,
    g1683_n_spl_0,
    G3438_o2_n_spl_1
  );


  and

  (
    g1685_p,
    g1684_p,
    G3449_o2_p_spl_01
  );


  or

  (
    g1685_n,
    g1684_n,
    G3449_o2_n_spl_01
  );


  and

  (
    g1686_p,
    g1685_p_spl_,
    G3428_o2_p_spl_11
  );


  or

  (
    g1686_n,
    g1685_n_spl_,
    G3428_o2_n_spl_11
  );


  and

  (
    g1687_p,
    g1678_n,
    G2693_o2_n_spl_
  );


  or

  (
    g1687_n,
    g1678_p,
    G2693_o2_p_spl_
  );


  and

  (
    g1688_p,
    g1687_p,
    g1680_n
  );


  or

  (
    g1688_n,
    g1687_n,
    g1680_p
  );


  and

  (
    g1689_p,
    g1688_p,
    g1682_n
  );


  or

  (
    g1689_n,
    g1688_n,
    g1682_p
  );


  and

  (
    g1690_p,
    g1689_p,
    g1686_n
  );


  or

  (
    g1690_n,
    g1689_n,
    g1686_p
  );


  and

  (
    g1691_p,
    g1690_p,
    G3421_o2_n_spl_1
  );


  and

  (
    g1692_p,
    g1690_n,
    G3421_o2_p_spl_1
  );


  or

  (
    g1693_n,
    g1692_p,
    g1691_p
  );


  and

  (
    g1694_p,
    g1693_n_spl_,
    n4719_lo_n_spl_0011
  );


  and

  (
    g1695_p,
    g1694_p,
    n4731_lo_p_spl_00110
  );


  and

  (
    g1696_p,
    n4719_lo_p_spl_00110,
    n3243_lo_p
  );


  and

  (
    g1697_p,
    g1696_p,
    n4731_lo_n_spl_0011
  );


  or

  (
    g1698_n,
    g1695_p,
    g1677_p
  );


  or

  (
    g1699_n,
    g1698_n,
    g1697_p
  );


  and

  (
    g1700_p,
    g1395_p_spl_,
    n4719_lo_p_spl_00111
  );


  and

  (
    g1701_p,
    g1700_p,
    n4731_lo_p_spl_00111
  );


  and

  (
    g1702_p,
    g1679_n_spl_,
    G2696_o2_n_spl_
  );


  or

  (
    g1702_n,
    g1679_p_spl_,
    G2696_o2_p_spl_
  );


  and

  (
    g1703_p,
    g1702_p,
    g1681_n_spl_
  );


  or

  (
    g1703_n,
    g1702_n,
    g1681_p_spl_
  );


  and

  (
    g1704_p,
    g1703_p,
    g1685_n_spl_
  );


  or

  (
    g1704_n,
    g1703_n,
    g1685_p_spl_
  );


  and

  (
    g1705_p,
    g1704_p,
    G3428_o2_n_spl_11
  );


  and

  (
    g1706_p,
    g1704_n,
    G3428_o2_p_spl_11
  );


  or

  (
    g1707_n,
    g1706_p,
    g1705_p
  );


  and

  (
    g1708_p,
    g1707_n_spl_,
    n4719_lo_n_spl_0011
  );


  and

  (
    g1709_p,
    g1708_p,
    n4731_lo_p_spl_00111
  );


  and

  (
    g1710_p,
    n4719_lo_p_spl_00111,
    n3291_lo_p
  );


  and

  (
    g1711_p,
    g1710_p,
    n4731_lo_n_spl_0011
  );


  or

  (
    g1712_n,
    g1709_p,
    g1701_p
  );


  or

  (
    g1713_n,
    g1712_n,
    g1711_p
  );


  and

  (
    g1714_p,
    g1385_p_spl_,
    n4719_lo_p_spl_01000
  );


  and

  (
    g1715_p,
    g1714_p,
    n4731_lo_p_spl_01000
  );


  and

  (
    g1716_p,
    G3449_o2_p_spl_01,
    G2705_o2_p_spl_1
  );


  or

  (
    g1716_n,
    G3449_o2_n_spl_01,
    G2705_o2_n_spl_1
  );


  and

  (
    g1717_p,
    g1683_p_spl_0,
    G3449_o2_p_spl_1
  );


  or

  (
    g1717_n,
    g1683_n_spl_0,
    G3449_o2_n_spl_1
  );


  and

  (
    g1718_p,
    g1716_n,
    G2700_o2_n_spl_
  );


  or

  (
    g1718_n,
    g1716_p,
    G2700_o2_p_spl_
  );


  and

  (
    g1719_p,
    g1718_p,
    g1717_n
  );


  or

  (
    g1719_n,
    g1718_n,
    g1717_p
  );


  and

  (
    g1720_p,
    g1719_p,
    G3438_o2_n_spl_1
  );


  and

  (
    g1721_p,
    g1719_n,
    G3438_o2_p_spl_1
  );


  or

  (
    g1722_n,
    g1721_p,
    g1720_p
  );


  and

  (
    g1723_p,
    g1722_n_spl_,
    n4719_lo_n_spl_0100
  );


  and

  (
    g1724_p,
    g1723_p,
    n4731_lo_p_spl_01000
  );


  and

  (
    g1725_p,
    n4719_lo_p_spl_01000,
    n3279_lo_p
  );


  and

  (
    g1726_p,
    g1725_p,
    n4731_lo_n_spl_0100
  );


  or

  (
    g1727_n,
    g1724_p,
    g1715_p
  );


  or

  (
    g1728_n,
    g1727_n,
    g1726_p
  );


  and

  (
    g1729_p,
    g1375_p_spl_,
    n4719_lo_p_spl_0100
  );


  and

  (
    g1730_p,
    g1729_p,
    n4731_lo_p_spl_0100
  );


  and

  (
    g1731_p,
    g1683_n_spl_,
    G2705_o2_n_spl_1
  );


  or

  (
    g1731_n,
    g1683_p_spl_,
    G2705_o2_p_spl_1
  );


  and

  (
    g1732_p,
    g1731_p,
    G3449_o2_n_spl_1
  );


  and

  (
    g1733_p,
    g1731_n,
    G3449_o2_p_spl_1
  );


  or

  (
    g1734_n,
    g1733_p,
    g1732_p
  );


  and

  (
    g1735_p,
    g1734_n_spl_,
    n4719_lo_n_spl_0100
  );


  and

  (
    g1736_p,
    g1735_p,
    n4731_lo_p_spl_0101
  );


  and

  (
    g1737_p,
    n4719_lo_p_spl_0101,
    n3267_lo_p
  );


  and

  (
    g1738_p,
    g1737_p,
    n4731_lo_n_spl_0100
  );


  or

  (
    g1739_n,
    g1736_p,
    g1730_p
  );


  or

  (
    g1740_n,
    g1739_n,
    g1738_p
  );


  and

  (
    g1741_p,
    G3265_o2_p,
    G3002_o2_n
  );


  or

  (
    g1741_n,
    G3265_o2_n,
    G3002_o2_p
  );


  and

  (
    g1742_p,
    G3266_o2_p,
    G2999_o2_n
  );


  or

  (
    g1742_n,
    G3266_o2_n,
    G2999_o2_p
  );


  and

  (
    g1743_p,
    g1742_n,
    g1741_n
  );


  or

  (
    g1743_n,
    g1742_p,
    g1741_p
  );


  and

  (
    g1744_p,
    G3267_o2_p,
    G3008_o2_n
  );


  or

  (
    g1744_n,
    G3267_o2_n,
    G3008_o2_p
  );


  and

  (
    g1745_p,
    G3268_o2_p,
    G3005_o2_n
  );


  or

  (
    g1745_n,
    G3268_o2_n,
    G3005_o2_p
  );


  and

  (
    g1746_p,
    g1745_n,
    g1744_n
  );


  or

  (
    g1746_n,
    g1745_p,
    g1744_p
  );


  and

  (
    g1747_p,
    g1746_p_spl_,
    g1743_n_spl_
  );


  or

  (
    g1747_n,
    g1746_n_spl_,
    g1743_p_spl_
  );


  and

  (
    g1748_p,
    g1746_n_spl_,
    g1743_p_spl_
  );


  or

  (
    g1748_n,
    g1746_p_spl_,
    g1743_n_spl_
  );


  and

  (
    g1749_p,
    g1748_n,
    g1747_n
  );


  or

  (
    g1749_n,
    g1748_p,
    g1747_p
  );


  and

  (
    g1750_p,
    G3335_o2_n,
    G3334_o2_n
  );


  or

  (
    g1750_n,
    G3335_o2_p,
    G3334_o2_p
  );


  and

  (
    g1751_p,
    G3336_o2_n,
    G3180_o2_p
  );


  or

  (
    g1751_n,
    G3336_o2_p,
    G3180_o2_n
  );


  and

  (
    g1752_p,
    g1751_p_spl_0,
    g1750_n_spl_0
  );


  or

  (
    g1752_n,
    g1751_n_spl_0,
    g1750_p_spl_0
  );


  and

  (
    g1753_p,
    g1752_p,
    G3674_o2_p_spl_0
  );


  or

  (
    g1753_n,
    g1752_n,
    G3674_o2_n_spl_0
  );


  and

  (
    g1754_p,
    g1751_p_spl_0,
    g1750_p_spl_0
  );


  or

  (
    g1754_n,
    g1751_n_spl_0,
    g1750_n_spl_0
  );


  and

  (
    g1755_p,
    g1754_p,
    G3674_o2_n_spl_0
  );


  or

  (
    g1755_n,
    g1754_n,
    G3674_o2_p_spl_0
  );


  and

  (
    g1756_p,
    g1755_n,
    g1753_n
  );


  or

  (
    g1756_n,
    g1755_p,
    g1753_p
  );


  and

  (
    g1757_p,
    g1751_n_spl_1,
    g1750_p_spl_1
  );


  or

  (
    g1757_n,
    g1751_p_spl_1,
    g1750_n_spl_1
  );


  and

  (
    g1758_p,
    g1757_p,
    G3674_o2_p_spl_1
  );


  or

  (
    g1758_n,
    g1757_n,
    G3674_o2_n_spl_1
  );


  and

  (
    g1759_p,
    g1751_n_spl_1,
    g1750_n_spl_1
  );


  or

  (
    g1759_n,
    g1751_p_spl_1,
    g1750_p_spl_1
  );


  and

  (
    g1760_p,
    g1759_p,
    G3674_o2_n_spl_1
  );


  or

  (
    g1760_n,
    g1759_n,
    G3674_o2_p_spl_1
  );


  and

  (
    g1761_p,
    g1760_n,
    g1758_n
  );


  or

  (
    g1761_n,
    g1760_p,
    g1758_p
  );


  and

  (
    g1762_p,
    g1761_p,
    g1756_p
  );


  or

  (
    g1762_n,
    g1761_n,
    g1756_n
  );


  and

  (
    g1763_p,
    g1762_p,
    g1749_n
  );


  and

  (
    g1764_p,
    g1762_n,
    g1749_p
  );


  or

  (
    g1765_n,
    g1764_p,
    g1763_p
  );


  and

  (
    g1766_p,
    G3269_o2_p,
    G3029_o2_n
  );


  or

  (
    g1766_n,
    G3269_o2_n,
    G3029_o2_p
  );


  and

  (
    g1767_p,
    G3270_o2_p,
    G3026_o2_n
  );


  or

  (
    g1767_n,
    G3270_o2_n,
    G3026_o2_p
  );


  and

  (
    g1768_p,
    g1767_n,
    g1766_n
  );


  or

  (
    g1768_n,
    g1767_p,
    g1766_p
  );


  and

  (
    g1769_p,
    G3271_o2_p,
    G3035_o2_n
  );


  or

  (
    g1769_n,
    G3271_o2_n,
    G3035_o2_p
  );


  and

  (
    g1770_p,
    G3272_o2_p,
    G3032_o2_n
  );


  or

  (
    g1770_n,
    G3272_o2_n,
    G3032_o2_p
  );


  and

  (
    g1771_p,
    g1770_n,
    g1769_n
  );


  or

  (
    g1771_n,
    g1770_p,
    g1769_p
  );


  and

  (
    g1772_p,
    g1771_p_spl_,
    g1768_n_spl_
  );


  or

  (
    g1772_n,
    g1771_n_spl_,
    g1768_p_spl_
  );


  and

  (
    g1773_p,
    g1771_n_spl_,
    g1768_p_spl_
  );


  or

  (
    g1773_n,
    g1771_p_spl_,
    g1768_n_spl_
  );


  and

  (
    g1774_p,
    g1773_n,
    g1772_n
  );


  or

  (
    g1774_n,
    g1773_p,
    g1772_p
  );


  and

  (
    g1775_p,
    G3338_o2_n,
    G3339_o2_n
  );


  or

  (
    g1775_n,
    G3338_o2_p,
    G3339_o2_p
  );


  and

  (
    g1776_p,
    G3341_o2_n,
    G3340_o2_n
  );


  or

  (
    g1776_n,
    G3341_o2_p,
    G3340_o2_p
  );


  and

  (
    g1777_p,
    g1776_p_spl_0,
    g1775_n_spl_0
  );


  or

  (
    g1777_n,
    g1776_n_spl_0,
    g1775_p_spl_0
  );


  and

  (
    g1778_p,
    g1777_p,
    G3685_o2_n_spl_0
  );


  or

  (
    g1778_n,
    g1777_n,
    G3685_o2_p_spl_0
  );


  and

  (
    g1779_p,
    g1776_p_spl_0,
    g1775_p_spl_0
  );


  or

  (
    g1779_n,
    g1776_n_spl_0,
    g1775_n_spl_0
  );


  and

  (
    g1780_p,
    g1779_p,
    G3685_o2_p_spl_0
  );


  or

  (
    g1780_n,
    g1779_n,
    G3685_o2_n_spl_0
  );


  and

  (
    g1781_p,
    g1780_n,
    g1778_n
  );


  or

  (
    g1781_n,
    g1780_p,
    g1778_p
  );


  and

  (
    g1782_p,
    g1776_n_spl_1,
    g1775_p_spl_1
  );


  or

  (
    g1782_n,
    g1776_p_spl_1,
    g1775_n_spl_1
  );


  and

  (
    g1783_p,
    g1782_p,
    G3685_o2_n_spl_1
  );


  or

  (
    g1783_n,
    g1782_n,
    G3685_o2_p_spl_1
  );


  and

  (
    g1784_p,
    g1776_n_spl_1,
    g1775_n_spl_1
  );


  or

  (
    g1784_n,
    g1776_p_spl_1,
    g1775_p_spl_1
  );


  and

  (
    g1785_p,
    g1784_p,
    G3685_o2_p_spl_1
  );


  or

  (
    g1785_n,
    g1784_n,
    G3685_o2_n_spl_1
  );


  and

  (
    g1786_p,
    g1785_n,
    g1783_n
  );


  or

  (
    g1786_n,
    g1785_p,
    g1783_p
  );


  and

  (
    g1787_p,
    g1786_p,
    g1781_p
  );


  or

  (
    g1787_n,
    g1786_n,
    g1781_n
  );


  and

  (
    g1788_p,
    g1787_p,
    g1774_n
  );


  and

  (
    g1789_p,
    g1787_n,
    g1774_p
  );


  or

  (
    g1790_n,
    g1789_p,
    g1788_p
  );


  and

  (
    g1791_p,
    g1423_p,
    n2631_lo_p_spl_
  );


  or

  (
    g1791_n,
    g1423_n_spl_,
    n2631_lo_n_spl_
  );


  and

  (
    g1792_p,
    g1791_n,
    g1536_p_spl_
  );


  or

  (
    g1792_n,
    g1791_p,
    g1536_n
  );


  and

  (
    g1793_p,
    g1792_p_spl_0,
    G3415_o2_p
  );


  and

  (
    g1794_p,
    g1792_n_spl_0,
    G3415_o2_n_spl_
  );


  or

  (
    g1795_n,
    g1794_p,
    g1793_p
  );


  and

  (
    g1796_p,
    G3404_o2_n_spl_,
    G2685_o2_p
  );


  and

  (
    g1797_p,
    G3404_o2_p,
    G2685_o2_n_spl_
  );


  or

  (
    g1798_n,
    g1797_p,
    g1796_p
  );


  and

  (
    g1799_p,
    g1798_n,
    g1792_p_spl_0
  );


  or

  (
    g1800_n,
    G3921_o2_p,
    G2915_o2_n
  );


  or

  (
    g1801_n,
    G3921_o2_n,
    G2915_o2_p
  );


  and

  (
    g1802_p,
    g1801_n,
    g1800_n
  );


  and

  (
    g1803_p,
    g1802_p,
    g1792_n_spl_0
  );


  or

  (
    g1804_n,
    g1803_p,
    g1799_p
  );


  or

  (
    g1805_n,
    G3918_o2_p,
    G4101_o2_n
  );


  or

  (
    g1806_n,
    G3918_o2_n,
    G4101_o2_p
  );


  and

  (
    g1807_p,
    g1806_n,
    g1805_n
  );


  and

  (
    g1808_p,
    g1807_p,
    g1792_p_spl_1
  );


  and

  (
    g1809_p,
    G3773_o2_n,
    G2679_o2_n_spl_
  );


  or

  (
    g1809_n,
    G3773_o2_p,
    G2679_o2_p
  );


  and

  (
    g1810_p,
    g1809_p,
    G3774_o2_n
  );


  or

  (
    g1810_n,
    g1809_n,
    G3774_o2_p
  );


  and

  (
    g1811_p,
    g1810_p,
    G3393_o2_n_spl_1
  );


  and

  (
    g1812_p,
    g1810_n,
    G3393_o2_p
  );


  or

  (
    g1813_n,
    g1812_p,
    g1811_p
  );


  and

  (
    g1814_p,
    g1813_n,
    g1792_n_spl_1
  );


  or

  (
    g1815_n,
    g1814_p,
    g1808_p
  );


  or

  (
    g1816_n,
    G3912_o2_p,
    G4095_o2_n
  );


  or

  (
    g1817_n,
    G3912_o2_n,
    G4095_o2_p
  );


  and

  (
    g1818_p,
    g1817_n,
    g1816_n
  );


  and

  (
    g1819_p,
    g1818_p,
    g1792_p_spl_1
  );


  and

  (
    g1820_p,
    G3768_o2_n,
    G2675_o2_n_spl_
  );


  or

  (
    g1820_n,
    G3768_o2_p,
    G2675_o2_p
  );


  and

  (
    g1821_p,
    g1820_p,
    G3769_o2_n
  );


  or

  (
    g1821_n,
    g1820_n,
    G3769_o2_p
  );


  and

  (
    g1822_p,
    g1821_p,
    G3770_o2_n
  );


  or

  (
    g1822_n,
    g1821_n,
    G3770_o2_p
  );


  and

  (
    g1823_p,
    g1822_p,
    G3386_o2_n_spl_1
  );


  and

  (
    g1824_p,
    g1822_n,
    G3386_o2_p
  );


  or

  (
    g1825_n,
    g1824_p,
    g1823_p
  );


  and

  (
    g1826_p,
    g1825_n,
    g1792_n_spl_1
  );


  or

  (
    g1827_n,
    g1826_p,
    g1819_p
  );


  or

  (
    g1828_n,
    g1734_n_spl_,
    g1581_n_spl_
  );


  or

  (
    g1829_n,
    g1828_n,
    g1722_n_spl_
  );


  or

  (
    g1830_n,
    g1829_n,
    g1707_n_spl_
  );


  or

  (
    g1831_n,
    g1830_n,
    g1693_n_spl_
  );


  or

  (
    g1832_n,
    g1831_n,
    g1795_n_spl_
  );


  or

  (
    g1833_n,
    g1832_n,
    g1804_n_spl_
  );


  or

  (
    g1834_n,
    g1833_n,
    g1815_n_spl_
  );


  or

  (
    g1835_n,
    g1834_n,
    g1827_n_spl_
  );


  and

  (
    g1836_p,
    g1592_p_spl_0,
    G3570_o2_p
  );


  and

  (
    g1837_p,
    g1592_n_spl_0,
    G3570_o2_n_spl_
  );


  or

  (
    g1838_n,
    g1837_p,
    g1836_p
  );


  and

  (
    g1839_p,
    G3559_o2_n_spl_,
    G2780_o2_p
  );


  and

  (
    g1840_p,
    G3559_o2_p,
    G2780_o2_n_spl_
  );


  or

  (
    g1841_n,
    g1840_p,
    g1839_p
  );


  and

  (
    g1842_p,
    g1841_n,
    g1592_p_spl_1
  );


  or

  (
    g1843_n,
    G3993_o2_p,
    G2966_o2_n
  );


  or

  (
    g1844_n,
    G3993_o2_n,
    G2966_o2_p
  );


  and

  (
    g1845_p,
    g1844_n,
    g1843_n
  );


  and

  (
    g1846_p,
    g1845_p,
    g1592_n_spl_1
  );


  or

  (
    g1847_n,
    g1846_p,
    g1842_p
  );


  or

  (
    g1848_n,
    G3234_o2_n,
    G4143_o2_n
  );


  or

  (
    g1849_n,
    G3234_o2_p,
    G4143_o2_p
  );


  and

  (
    g1850_p,
    g1849_n,
    g1848_n
  );


  and

  (
    g1851_p,
    g1850_p,
    g1592_p_spl_1
  );


  and

  (
    g1852_p,
    G3831_o2_n,
    G2774_o2_n_spl_
  );


  or

  (
    g1852_n,
    G3831_o2_p,
    G2774_o2_p
  );


  and

  (
    g1853_p,
    g1852_p,
    G3832_o2_n
  );


  or

  (
    g1853_n,
    g1852_n,
    G3832_o2_p
  );


  and

  (
    g1854_p,
    g1853_p,
    G2759_o2_p_spl_1
  );


  and

  (
    g1855_p,
    g1853_n,
    G2759_o2_n
  );


  or

  (
    g1856_n,
    g1855_p,
    g1854_p
  );


  and

  (
    g1857_p,
    g1856_n,
    g1592_n_spl_1
  );


  or

  (
    g1858_n,
    g1857_p,
    g1851_p
  );


  or

  (
    g1859_n,
    g1570_n_spl_,
    g1557_n_spl_
  );


  or

  (
    g1860_n,
    g1859_n,
    g1658_n_spl_
  );


  or

  (
    g1861_n,
    g1860_n,
    g1643_n_spl_
  );


  or

  (
    g1862_n,
    g1861_n,
    g1629_n_spl_
  );


  or

  (
    g1863_n,
    g1862_n,
    g1838_n_spl_
  );


  or

  (
    g1864_n,
    g1863_n,
    g1847_n_spl_
  );


  or

  (
    g1865_n,
    g1864_n,
    g1858_n_spl_
  );


  or

  (
    g1866_n,
    g1865_n,
    g1601_n_spl_0
  );


  and

  (
    g1867_p,
    g1563_n_spl_0,
    n4503_lo_p_spl_0000
  );


  and

  (
    g1868_p,
    g1867_p,
    n4515_lo_p_spl_0000
  );


  and

  (
    g1869_p,
    g1587_n_spl_0,
    n4503_lo_n_spl_0000
  );


  and

  (
    g1870_p,
    g1869_p,
    n4515_lo_p_spl_0000
  );


  and

  (
    g1871_p,
    n4503_lo_p_spl_0000,
    n3567_lo_p_spl_
  );


  and

  (
    g1872_p,
    g1871_p,
    n4515_lo_n_spl_0000
  );


  and

  (
    g1873_p,
    n4503_lo_n_spl_0000,
    n3579_lo_p_spl_
  );


  and

  (
    g1874_p,
    g1873_p,
    n4515_lo_n_spl_0000
  );


  or

  (
    g1875_n,
    g1870_p,
    g1868_p
  );


  or

  (
    g1876_n,
    g1875_n,
    g1872_p
  );


  or

  (
    g1877_n,
    g1876_n,
    g1874_p
  );


  and

  (
    g1878_p,
    g1877_n,
    n3375_lo_p_spl_0000
  );


  and

  (
    g1879_p,
    g1563_n_spl_1,
    n4527_lo_p_spl_0000
  );


  and

  (
    g1880_p,
    g1879_p,
    n4539_lo_p_spl_0000
  );


  and

  (
    g1881_p,
    g1587_n_spl_1,
    n4527_lo_n_spl_0000
  );


  and

  (
    g1882_p,
    g1881_p,
    n4539_lo_p_spl_0000
  );


  and

  (
    g1883_p,
    n4527_lo_p_spl_0000,
    n3567_lo_p_spl_
  );


  and

  (
    g1884_p,
    g1883_p,
    n4539_lo_n_spl_0000
  );


  and

  (
    g1885_p,
    n4527_lo_n_spl_0000,
    n3579_lo_p_spl_
  );


  and

  (
    g1886_p,
    g1885_p,
    n4539_lo_n_spl_0000
  );


  or

  (
    g1887_n,
    g1882_p,
    g1880_p
  );


  or

  (
    g1888_n,
    g1887_n,
    g1884_p
  );


  or

  (
    g1889_n,
    g1888_n,
    g1886_p
  );


  and

  (
    g1890_p,
    g1889_n,
    n3375_lo_p_spl_0000
  );


  and

  (
    g1891_p,
    g1635_n_spl_00,
    n4683_lo_p_spl_0001
  );


  and

  (
    g1892_p,
    g1891_p,
    n4671_lo_p_spl_0001
  );


  and

  (
    g1893_p,
    g1699_n_spl_00,
    n4683_lo_n_spl_0001
  );


  and

  (
    g1894_p,
    g1893_p,
    n4671_lo_p_spl_0001
  );


  and

  (
    g1895_p,
    n4683_lo_p_spl_0001,
    n2799_lo_p_spl_
  );


  and

  (
    g1896_p,
    g1895_p,
    n4671_lo_n_spl_0001
  );


  and

  (
    g1897_p,
    n4683_lo_n_spl_0001,
    n2775_lo_p_spl_
  );


  and

  (
    g1898_p,
    g1897_p,
    n4671_lo_n_spl_0001
  );


  or

  (
    g1899_n,
    g1894_p,
    g1892_p
  );


  or

  (
    g1900_n,
    g1899_n,
    g1896_p
  );


  or

  (
    g1901_n,
    g1900_n,
    g1898_p
  );


  and

  (
    g1902_p,
    g1649_n_spl_00,
    n4683_lo_p_spl_0010
  );


  and

  (
    g1903_p,
    g1902_p,
    n4671_lo_p_spl_0010
  );


  and

  (
    g1904_p,
    g1713_n_spl_00,
    n4683_lo_n_spl_0010
  );


  and

  (
    g1905_p,
    g1904_p,
    n4671_lo_p_spl_0010
  );


  and

  (
    g1906_p,
    n4683_lo_p_spl_0010,
    n2931_lo_p_spl_
  );


  and

  (
    g1907_p,
    g1906_p,
    n4671_lo_n_spl_0010
  );


  and

  (
    g1908_p,
    n4683_lo_n_spl_0010,
    n2679_lo_p_spl_
  );


  and

  (
    g1909_p,
    g1908_p,
    n4671_lo_n_spl_0010
  );


  or

  (
    g1910_n,
    g1905_p,
    g1903_p
  );


  or

  (
    g1911_n,
    g1910_n,
    g1907_p
  );


  or

  (
    g1912_n,
    g1911_n,
    g1909_p
  );


  and

  (
    g1913_p,
    g1664_n_spl_00,
    n4683_lo_p_spl_0011
  );


  and

  (
    g1914_p,
    g1913_p,
    n4671_lo_p_spl_0011
  );


  and

  (
    g1915_p,
    g1728_n_spl_00,
    n4683_lo_n_spl_0011
  );


  and

  (
    g1916_p,
    g1915_p,
    n4671_lo_p_spl_0011
  );


  and

  (
    g1917_p,
    n4683_lo_p_spl_0011,
    n2919_lo_p_spl_
  );


  and

  (
    g1918_p,
    g1917_p,
    n4671_lo_n_spl_0011
  );


  and

  (
    g1919_p,
    n4683_lo_n_spl_0011,
    n2667_lo_p_spl_
  );


  and

  (
    g1920_p,
    g1919_p,
    n4671_lo_n_spl_0011
  );


  or

  (
    g1921_n,
    g1916_p,
    g1914_p
  );


  or

  (
    g1922_n,
    g1921_n,
    g1918_p
  );


  or

  (
    g1923_n,
    g1922_n,
    g1920_p
  );


  and

  (
    g1924_p,
    g1576_n_spl_00,
    n4683_lo_p_spl_010
  );


  and

  (
    g1925_p,
    g1924_p,
    n4671_lo_p_spl_010
  );


  and

  (
    g1926_p,
    g1740_n_spl_00,
    n4683_lo_n_spl_010
  );


  and

  (
    g1927_p,
    g1926_p,
    n4671_lo_p_spl_010
  );


  and

  (
    g1928_p,
    n4683_lo_p_spl_010,
    n2895_lo_p_spl_
  );


  and

  (
    g1929_p,
    g1928_p,
    n4671_lo_n_spl_010
  );


  and

  (
    g1930_p,
    n4683_lo_n_spl_010,
    n2907_lo_p_spl_
  );


  and

  (
    g1931_p,
    g1930_p,
    n4671_lo_n_spl_010
  );


  or

  (
    g1932_n,
    g1927_p,
    g1925_p
  );


  or

  (
    g1933_n,
    g1932_n,
    g1929_p
  );


  or

  (
    g1934_n,
    g1933_n,
    g1931_p
  );


  and

  (
    g1935_p,
    g1635_n_spl_00,
    n4695_lo_p_spl_0001
  );


  and

  (
    g1936_p,
    g1935_p,
    n4707_lo_p_spl_0001
  );


  and

  (
    g1937_p,
    g1699_n_spl_00,
    n4695_lo_n_spl_0001
  );


  and

  (
    g1938_p,
    g1937_p,
    n4707_lo_p_spl_0001
  );


  and

  (
    g1939_p,
    n4695_lo_p_spl_0001,
    n2799_lo_p_spl_
  );


  and

  (
    g1940_p,
    g1939_p,
    n4707_lo_n_spl_0001
  );


  and

  (
    g1941_p,
    n4695_lo_n_spl_0001,
    n2775_lo_p_spl_
  );


  and

  (
    g1942_p,
    g1941_p,
    n4707_lo_n_spl_0001
  );


  or

  (
    g1943_n,
    g1938_p,
    g1936_p
  );


  or

  (
    g1944_n,
    g1943_n,
    g1940_p
  );


  or

  (
    g1945_n,
    g1944_n,
    g1942_p
  );


  and

  (
    g1946_p,
    g1649_n_spl_00,
    n4695_lo_p_spl_0010
  );


  and

  (
    g1947_p,
    g1946_p,
    n4707_lo_p_spl_0010
  );


  and

  (
    g1948_p,
    g1713_n_spl_00,
    n4695_lo_n_spl_0010
  );


  and

  (
    g1949_p,
    g1948_p,
    n4707_lo_p_spl_0010
  );


  and

  (
    g1950_p,
    n4695_lo_p_spl_0010,
    n2931_lo_p_spl_
  );


  and

  (
    g1951_p,
    g1950_p,
    n4707_lo_n_spl_0010
  );


  and

  (
    g1952_p,
    n4695_lo_n_spl_0010,
    n2679_lo_p_spl_
  );


  and

  (
    g1953_p,
    g1952_p,
    n4707_lo_n_spl_0010
  );


  or

  (
    g1954_n,
    g1949_p,
    g1947_p
  );


  or

  (
    g1955_n,
    g1954_n,
    g1951_p
  );


  or

  (
    g1956_n,
    g1955_n,
    g1953_p
  );


  and

  (
    g1957_p,
    g1664_n_spl_00,
    n4695_lo_p_spl_0011
  );


  and

  (
    g1958_p,
    g1957_p,
    n4707_lo_p_spl_0011
  );


  and

  (
    g1959_p,
    g1728_n_spl_00,
    n4695_lo_n_spl_0011
  );


  and

  (
    g1960_p,
    g1959_p,
    n4707_lo_p_spl_0011
  );


  and

  (
    g1961_p,
    n4695_lo_p_spl_0011,
    n2919_lo_p_spl_
  );


  and

  (
    g1962_p,
    g1961_p,
    n4707_lo_n_spl_0011
  );


  and

  (
    g1963_p,
    n4695_lo_n_spl_0011,
    n2667_lo_p_spl_
  );


  and

  (
    g1964_p,
    g1963_p,
    n4707_lo_n_spl_0011
  );


  or

  (
    g1965_n,
    g1960_p,
    g1958_p
  );


  or

  (
    g1966_n,
    g1965_n,
    g1962_p
  );


  or

  (
    g1967_n,
    g1966_n,
    g1964_p
  );


  and

  (
    g1968_p,
    g1576_n_spl_00,
    n4695_lo_p_spl_010
  );


  and

  (
    g1969_p,
    g1968_p,
    n4707_lo_p_spl_010
  );


  and

  (
    g1970_p,
    g1740_n_spl_00,
    n4695_lo_n_spl_010
  );


  and

  (
    g1971_p,
    g1970_p,
    n4707_lo_p_spl_010
  );


  and

  (
    g1972_p,
    n4695_lo_p_spl_010,
    n2895_lo_p_spl_
  );


  and

  (
    g1973_p,
    g1972_p,
    n4707_lo_n_spl_010
  );


  and

  (
    g1974_p,
    n4695_lo_n_spl_010,
    n2907_lo_p_spl_
  );


  and

  (
    g1975_p,
    g1974_p,
    n4707_lo_n_spl_010
  );


  or

  (
    g1976_n,
    g1971_p,
    g1969_p
  );


  or

  (
    g1977_n,
    g1976_n,
    g1973_p
  );


  or

  (
    g1978_n,
    g1977_n,
    g1975_p
  );


  and

  (
    g1979_p,
    g1635_n_spl_0,
    n4503_lo_p_spl_0001
  );


  and

  (
    g1980_p,
    g1979_p,
    n4515_lo_p_spl_0001
  );


  and

  (
    g1981_p,
    g1699_n_spl_0,
    n4503_lo_n_spl_0001
  );


  and

  (
    g1982_p,
    g1981_p,
    n4515_lo_p_spl_0001
  );


  and

  (
    g1983_p,
    n4503_lo_p_spl_0001,
    n3639_lo_p_spl_
  );


  and

  (
    g1984_p,
    g1983_p,
    n4515_lo_n_spl_0001
  );


  and

  (
    g1985_p,
    n4503_lo_n_spl_0001,
    n3519_lo_p_spl_
  );


  and

  (
    g1986_p,
    g1985_p,
    n4515_lo_n_spl_0001
  );


  or

  (
    g1987_n,
    g1982_p,
    g1980_p
  );


  or

  (
    g1988_n,
    g1987_n,
    g1984_p
  );


  or

  (
    g1989_n,
    g1988_n,
    g1986_p
  );


  and

  (
    g1990_p,
    g1989_n,
    n3375_lo_p_spl_0001
  );


  and

  (
    g1991_p,
    g1576_n_spl_0,
    n4503_lo_p_spl_0010
  );


  and

  (
    g1992_p,
    g1991_p,
    n4515_lo_p_spl_0010
  );


  and

  (
    g1993_p,
    g1740_n_spl_0,
    n4503_lo_n_spl_0010
  );


  and

  (
    g1994_p,
    g1993_p,
    n4515_lo_p_spl_0010
  );


  and

  (
    g1995_p,
    n4503_lo_p_spl_0010,
    n3591_lo_p_spl_
  );


  and

  (
    g1996_p,
    g1995_p,
    n4515_lo_n_spl_0010
  );


  and

  (
    g1997_p,
    n4503_lo_n_spl_0010,
    n3471_lo_p_spl_
  );


  and

  (
    g1998_p,
    g1997_p,
    n4515_lo_n_spl_0010
  );


  or

  (
    g1999_n,
    g1994_p,
    g1992_p
  );


  or

  (
    g2000_n,
    g1999_n,
    g1996_p
  );


  or

  (
    g2001_n,
    g2000_n,
    g1998_p
  );


  and

  (
    g2002_p,
    g2001_n,
    n3375_lo_p_spl_0001
  );


  and

  (
    g2003_p,
    g1664_n_spl_0,
    n4503_lo_p_spl_0011
  );


  and

  (
    g2004_p,
    g2003_p,
    n4515_lo_p_spl_0011
  );


  and

  (
    g2005_p,
    g1728_n_spl_0,
    n4503_lo_n_spl_0011
  );


  and

  (
    g2006_p,
    g2005_p,
    n4515_lo_p_spl_0011
  );


  and

  (
    g2007_p,
    n4503_lo_p_spl_0011,
    n3459_lo_p_spl_
  );


  and

  (
    g2008_p,
    g2007_p,
    n4515_lo_n_spl_0011
  );


  and

  (
    g2009_p,
    n4503_lo_n_spl_0011,
    n3447_lo_p_spl_
  );


  and

  (
    g2010_p,
    g2009_p,
    n4515_lo_n_spl_0011
  );


  or

  (
    g2011_n,
    g2006_p,
    g2004_p
  );


  or

  (
    g2012_n,
    g2011_n,
    g2008_p
  );


  or

  (
    g2013_n,
    g2012_n,
    g2010_p
  );


  and

  (
    g2014_p,
    g2013_n,
    n3375_lo_p_spl_0010
  );


  and

  (
    g2015_p,
    g1649_n_spl_0,
    n4503_lo_p_spl_010
  );


  and

  (
    g2016_p,
    g2015_p,
    n4515_lo_p_spl_010
  );


  and

  (
    g2017_p,
    g1713_n_spl_0,
    n4503_lo_n_spl_010
  );


  and

  (
    g2018_p,
    g2017_p,
    n4515_lo_p_spl_010
  );


  and

  (
    g2019_p,
    n4503_lo_p_spl_010,
    n3435_lo_p_spl_
  );


  and

  (
    g2020_p,
    g2019_p,
    n4515_lo_n_spl_010
  );


  and

  (
    g2021_p,
    n4503_lo_n_spl_010,
    n3423_lo_p_spl_
  );


  and

  (
    g2022_p,
    g2021_p,
    n4515_lo_n_spl_010
  );


  or

  (
    g2023_n,
    g2018_p,
    g2016_p
  );


  or

  (
    g2024_n,
    g2023_n,
    g2020_p
  );


  or

  (
    g2025_n,
    g2024_n,
    g2022_p
  );


  and

  (
    g2026_p,
    g2025_n,
    n3375_lo_p_spl_0010
  );


  and

  (
    g2027_p,
    g1635_n_spl_1,
    n4527_lo_p_spl_0001
  );


  and

  (
    g2028_p,
    g2027_p,
    n4539_lo_p_spl_0001
  );


  and

  (
    g2029_p,
    g1699_n_spl_1,
    n4527_lo_n_spl_0001
  );


  and

  (
    g2030_p,
    g2029_p,
    n4539_lo_p_spl_0001
  );


  and

  (
    g2031_p,
    n4527_lo_p_spl_0001,
    n3639_lo_p_spl_
  );


  and

  (
    g2032_p,
    g2031_p,
    n4539_lo_n_spl_0001
  );


  and

  (
    g2033_p,
    n4527_lo_n_spl_0001,
    n3519_lo_p_spl_
  );


  and

  (
    g2034_p,
    g2033_p,
    n4539_lo_n_spl_0001
  );


  or

  (
    g2035_n,
    g2030_p,
    g2028_p
  );


  or

  (
    g2036_n,
    g2035_n,
    g2032_p
  );


  or

  (
    g2037_n,
    g2036_n,
    g2034_p
  );


  and

  (
    g2038_p,
    g2037_n,
    n3375_lo_p_spl_0011
  );


  and

  (
    g2039_p,
    g1576_n_spl_1,
    n4527_lo_p_spl_0010
  );


  and

  (
    g2040_p,
    g2039_p,
    n4539_lo_p_spl_0010
  );


  and

  (
    g2041_p,
    g1740_n_spl_1,
    n4527_lo_n_spl_0010
  );


  and

  (
    g2042_p,
    g2041_p,
    n4539_lo_p_spl_0010
  );


  and

  (
    g2043_p,
    n4527_lo_p_spl_0010,
    n3591_lo_p_spl_
  );


  and

  (
    g2044_p,
    g2043_p,
    n4539_lo_n_spl_0010
  );


  and

  (
    g2045_p,
    n4527_lo_n_spl_0010,
    n3471_lo_p_spl_
  );


  and

  (
    g2046_p,
    g2045_p,
    n4539_lo_n_spl_0010
  );


  or

  (
    g2047_n,
    g2042_p,
    g2040_p
  );


  or

  (
    g2048_n,
    g2047_n,
    g2044_p
  );


  or

  (
    g2049_n,
    g2048_n,
    g2046_p
  );


  and

  (
    g2050_p,
    g2049_n,
    n3375_lo_p_spl_0011
  );


  and

  (
    g2051_p,
    g1664_n_spl_1,
    n4527_lo_p_spl_0011
  );


  and

  (
    g2052_p,
    g2051_p,
    n4539_lo_p_spl_0011
  );


  and

  (
    g2053_p,
    g1728_n_spl_1,
    n4527_lo_n_spl_0011
  );


  and

  (
    g2054_p,
    g2053_p,
    n4539_lo_p_spl_0011
  );


  and

  (
    g2055_p,
    n4527_lo_p_spl_0011,
    n3459_lo_p_spl_
  );


  and

  (
    g2056_p,
    g2055_p,
    n4539_lo_n_spl_0011
  );


  and

  (
    g2057_p,
    n4527_lo_n_spl_0011,
    n3447_lo_p_spl_
  );


  and

  (
    g2058_p,
    g2057_p,
    n4539_lo_n_spl_0011
  );


  or

  (
    g2059_n,
    g2054_p,
    g2052_p
  );


  or

  (
    g2060_n,
    g2059_n,
    g2056_p
  );


  or

  (
    g2061_n,
    g2060_n,
    g2058_p
  );


  and

  (
    g2062_p,
    g2061_n,
    n3375_lo_p_spl_0100
  );


  and

  (
    g2063_p,
    g1649_n_spl_1,
    n4527_lo_p_spl_010
  );


  and

  (
    g2064_p,
    g2063_p,
    n4539_lo_p_spl_010
  );


  and

  (
    g2065_p,
    g1713_n_spl_1,
    n4527_lo_n_spl_010
  );


  and

  (
    g2066_p,
    g2065_p,
    n4539_lo_p_spl_010
  );


  and

  (
    g2067_p,
    n4527_lo_p_spl_010,
    n3435_lo_p_spl_
  );


  and

  (
    g2068_p,
    g2067_p,
    n4539_lo_n_spl_010
  );


  and

  (
    g2069_p,
    n4527_lo_n_spl_010,
    n3423_lo_p_spl_
  );


  and

  (
    g2070_p,
    g2069_p,
    n4539_lo_n_spl_010
  );


  or

  (
    g2071_n,
    g2066_p,
    g2064_p
  );


  or

  (
    g2072_n,
    g2071_n,
    g2068_p
  );


  or

  (
    g2073_n,
    g2072_n,
    g2070_p
  );


  and

  (
    g2074_p,
    g2073_n,
    n3375_lo_p_spl_0100
  );


  or

  (
    g2075_n,
    n4743_lo_n,
    n3351_lo_n
  );


  and

  (
    g2076_p,
    g1271_p_spl_,
    n4659_lo_n_spl_
  );


  and

  (
    g2077_p,
    g2076_p,
    n4647_lo_n_spl_
  );


  and

  (
    g2078_p,
    n7463_o2_p_spl_,
    n3339_lo_p_spl_
  );


  or

  (
    g2078_n,
    n7463_o2_n_spl_1,
    n3339_lo_n_spl_
  );


  and

  (
    g2079_p,
    g2078_n_spl_,
    n7463_o2_p_spl_
  );


  or

  (
    g2079_n,
    g2078_p_spl_,
    n7463_o2_n_spl_1
  );


  and

  (
    g2080_p,
    g2078_n_spl_,
    n3339_lo_p_spl_
  );


  or

  (
    g2080_n,
    g2078_p_spl_,
    n3339_lo_n_spl_
  );


  and

  (
    g2081_p,
    g2080_n,
    g2079_n
  );


  or

  (
    g2081_n,
    g2080_p,
    g2079_p
  );


  and

  (
    g2082_p,
    g2081_n_spl_,
    n4659_lo_p_spl_
  );


  and

  (
    g2083_p,
    g2082_p,
    n4647_lo_n_spl_
  );


  and

  (
    g2084_p,
    n4659_lo_n_spl_,
    n3255_lo_p_spl_
  );


  and

  (
    g2085_p,
    g2084_p,
    n4647_lo_p_spl_
  );


  and

  (
    g2086_p,
    g1601_n_spl_0,
    n4659_lo_p_spl_
  );


  and

  (
    g2087_p,
    g2086_p,
    n4647_lo_p_spl_
  );


  or

  (
    g2088_n,
    g2083_p,
    g2077_p
  );


  or

  (
    g2089_n,
    g2088_n,
    g2085_p
  );


  or

  (
    g2090_n,
    g2089_n,
    g2087_p
  );


  and

  (
    g2091_p,
    g2090_n,
    g2075_n
  );


  or

  (
    g2092_n,
    g2081_p,
    g1601_p_spl_
  );


  and

  (
    g2093_p,
    g2092_n_spl_,
    g2081_n_spl_
  );


  and

  (
    g2094_p,
    g2092_n_spl_,
    g1601_n_spl_1
  );


  or

  (
    g2095_n,
    g2094_p,
    g2093_p
  );


  and

  (
    g2096_p,
    g1271_p_spl_,
    n4719_lo_p_spl_0101
  );


  and

  (
    g2097_p,
    g2096_p,
    n4731_lo_p_spl_0101
  );


  and

  (
    g2098_p,
    g1601_n_spl_1,
    n4719_lo_n_spl_0101
  );


  and

  (
    g2099_p,
    g2098_p,
    n4731_lo_p_spl_0110
  );


  and

  (
    g2100_p,
    n4719_lo_p_spl_0110,
    n3255_lo_p_spl_
  );


  and

  (
    g2101_p,
    g2100_p,
    n4731_lo_n_spl_0101
  );


  or

  (
    g2102_n,
    g2099_p,
    g2097_p
  );


  or

  (
    g2103_n,
    g2102_n,
    g2101_p
  );


  and

  (
    g2104_p,
    g1268_p_spl_,
    n4719_lo_p_spl_0110
  );


  and

  (
    g2105_p,
    g2104_p,
    n4731_lo_p_spl_0110
  );


  and

  (
    g2106_p,
    g1858_n_spl_,
    n4719_lo_n_spl_0101
  );


  and

  (
    g2107_p,
    g2106_p,
    n4731_lo_p_spl_0111
  );


  and

  (
    g2108_p,
    n4719_lo_p_spl_0111,
    n3231_lo_p
  );


  and

  (
    g2109_p,
    g2108_p,
    n4731_lo_n_spl_0101
  );


  or

  (
    g2110_n,
    g2107_p,
    g2105_p
  );


  or

  (
    g2111_n,
    g2110_n,
    g2109_p
  );


  and

  (
    g2112_p,
    g1265_p_spl_,
    n4719_lo_p_spl_0111
  );


  and

  (
    g2113_p,
    g2112_p,
    n4731_lo_p_spl_0111
  );


  and

  (
    g2114_p,
    g1847_n_spl_,
    n4719_lo_n_spl_0110
  );


  and

  (
    g2115_p,
    g2114_p,
    n4731_lo_p_spl_1000
  );


  and

  (
    g2116_p,
    n4719_lo_p_spl_1000,
    n3171_lo_p
  );


  and

  (
    g2117_p,
    g2116_p,
    n4731_lo_n_spl_0110
  );


  or

  (
    g2118_n,
    g2115_p,
    g2113_p
  );


  or

  (
    g2119_n,
    g2118_n,
    g2117_p
  );


  and

  (
    g2120_p,
    g1255_p_spl_,
    n4719_lo_p_spl_1000
  );


  and

  (
    g2121_p,
    g2120_p,
    n4731_lo_p_spl_1000
  );


  and

  (
    g2122_p,
    g1838_n_spl_,
    n4719_lo_n_spl_0110
  );


  and

  (
    g2123_p,
    g2122_p,
    n4731_lo_p_spl_1001
  );


  and

  (
    g2124_p,
    n4719_lo_p_spl_1001,
    n3123_lo_p
  );


  and

  (
    g2125_p,
    g2124_p,
    n4731_lo_n_spl_0110
  );


  or

  (
    g2126_n,
    g2123_p,
    g2121_p
  );


  or

  (
    g2127_n,
    g2126_n,
    g2125_p
  );


  or

  (
    g2128_n,
    n4467_lo_n_spl_,
    n4239_lo_n_spl_
  );


  or

  (
    g2129_n,
    g2128_n,
    n4455_lo_n_spl_
  );


  or

  (
    g2130_n,
    g2129_n,
    n4443_lo_n_spl_
  );


  or

  (
    g2131_n,
    g1765_n_spl_,
    n4479_lo_n_spl_
  );


  or

  (
    g2132_n,
    g2131_n,
    g1790_n_spl_
  );


  or

  (
    g2133_n,
    g2132_n,
    g1449_n_spl_
  );


  or

  (
    g2134_n,
    g2133_n,
    g1474_n_spl_
  );


  or

  (
    g2135_n,
    g2134_n,
    g2130_n
  );


  or

  (
    g2136_n,
    g2135_n,
    n3795_lo_n_spl_
  );


  or

  (
    g2137_n,
    n7358_o2_p_spl_,
    n4311_lo_n_spl_0
  );


  or

  (
    g2138_n,
    g2137_n,
    n7156_o2_n_spl_
  );


  or

  (
    g2139_n,
    n7360_o2_p_spl_,
    n4311_lo_n_spl_
  );


  or

  (
    g2140_n,
    g2139_n,
    n7156_o2_p_spl_
  );


  and

  (
    g2141_p,
    g2140_n,
    g2138_n
  );


  and

  (
    g2142_p,
    n7450_o2_n,
    n7156_o2_p_spl_
  );


  and

  (
    g2143_p,
    n7451_o2_n,
    n7156_o2_n_spl_
  );


  or

  (
    g2144_n,
    g2143_p,
    g2142_p
  );


  or

  (
    g2145_n,
    g2144_n,
    n4311_lo_p
  );


  and

  (
    g2146_p,
    g2145_n,
    g2141_p
  );


  and

  (
    g2147_p,
    g2146_p,
    n4719_lo_p_spl_1001
  );


  and

  (
    g2148_p,
    g2147_p,
    n4731_lo_p_spl_1001
  );


  and

  (
    g2149_p,
    g1827_n_spl_,
    n4719_lo_n_spl_0111
  );


  and

  (
    g2150_p,
    g2149_p,
    n4731_lo_p_spl_1010
  );


  and

  (
    g2151_p,
    n4719_lo_p_spl_1010,
    n3159_lo_p
  );


  and

  (
    g2152_p,
    g2151_p,
    n4731_lo_n_spl_0111
  );


  or

  (
    g2153_n,
    g2150_p,
    g2148_p
  );


  or

  (
    g2154_n,
    g2153_n,
    g2152_p
  );


  and

  (
    g2155_p,
    g1352_p_spl_,
    n4719_lo_p_spl_1010
  );


  and

  (
    g2156_p,
    g2155_p,
    n4731_lo_p_spl_1010
  );


  and

  (
    g2157_p,
    g1815_n_spl_,
    n4719_lo_n_spl_0111
  );


  and

  (
    g2158_p,
    g2157_p,
    n4731_lo_p_spl_1011
  );


  and

  (
    g2159_p,
    n4719_lo_p_spl_1011,
    n3147_lo_p
  );


  and

  (
    g2160_p,
    g2159_p,
    n4731_lo_n_spl_0111
  );


  or

  (
    g2161_n,
    g2158_p,
    g2156_p
  );


  or

  (
    g2162_n,
    g2161_n,
    g2160_p
  );


  and

  (
    g2163_p,
    g1342_p_spl_,
    n4719_lo_p_spl_1011
  );


  and

  (
    g2164_p,
    g2163_p,
    n4731_lo_p_spl_1011
  );


  and

  (
    g2165_p,
    g1804_n_spl_,
    n4719_lo_n_spl_100
  );


  and

  (
    g2166_p,
    g2165_p,
    n4731_lo_p_spl_1100
  );


  and

  (
    g2167_p,
    n4719_lo_p_spl_1100,
    n2847_lo_p
  );


  and

  (
    g2168_p,
    g2167_p,
    n4731_lo_n_spl_100
  );


  or

  (
    g2169_n,
    g2166_p,
    g2164_p
  );


  or

  (
    g2170_n,
    g2169_n,
    g2168_p
  );


  and

  (
    g2171_p,
    g1332_p_spl_,
    n4719_lo_p_spl_1100
  );


  and

  (
    g2172_p,
    g2171_p,
    n4731_lo_p_spl_1100
  );


  and

  (
    g2173_p,
    g1795_n_spl_,
    n4719_lo_n_spl_100
  );


  and

  (
    g2174_p,
    g2173_p,
    n4731_lo_p_spl_1101
  );


  and

  (
    g2175_p,
    n4719_lo_p_spl_1101,
    n3135_lo_p
  );


  and

  (
    g2176_p,
    g2175_p,
    n4731_lo_n_spl_100
  );


  or

  (
    g2177_n,
    g2174_p,
    g2172_p
  );


  or

  (
    g2178_n,
    g2177_n,
    g2176_p
  );


  and

  (
    g2179_p,
    g2103_n_spl_00,
    n4695_lo_p_spl_011
  );


  and

  (
    g2180_p,
    g2179_p,
    n4707_lo_p_spl_011
  );


  and

  (
    g2181_p,
    g2154_n_spl_00,
    n4695_lo_n_spl_011
  );


  and

  (
    g2182_p,
    g2181_p,
    n4707_lo_p_spl_011
  );


  and

  (
    g2183_p,
    n4695_lo_p_spl_011,
    n3111_lo_p_spl_
  );


  and

  (
    g2184_p,
    g2183_p,
    n4707_lo_n_spl_011
  );


  and

  (
    g2185_p,
    n4695_lo_n_spl_011,
    n3099_lo_p_spl_
  );


  and

  (
    g2186_p,
    g2185_p,
    n4707_lo_n_spl_011
  );


  or

  (
    g2187_n,
    g2182_p,
    g2180_p
  );


  or

  (
    g2188_n,
    g2187_n,
    g2184_p
  );


  or

  (
    g2189_n,
    g2188_n,
    g2186_p
  );


  and

  (
    g2190_p,
    g2103_n_spl_00,
    n4683_lo_p_spl_011
  );


  and

  (
    g2191_p,
    g2190_p,
    n4671_lo_p_spl_011
  );


  and

  (
    g2192_p,
    g2154_n_spl_00,
    n4683_lo_n_spl_011
  );


  and

  (
    g2193_p,
    g2192_p,
    n4671_lo_p_spl_011
  );


  and

  (
    g2194_p,
    n4683_lo_p_spl_011,
    n3111_lo_p_spl_
  );


  and

  (
    g2195_p,
    g2194_p,
    n4671_lo_n_spl_011
  );


  and

  (
    g2196_p,
    n4683_lo_n_spl_011,
    n3099_lo_p_spl_
  );


  and

  (
    g2197_p,
    g2196_p,
    n4671_lo_n_spl_011
  );


  or

  (
    g2198_n,
    g2193_p,
    g2191_p
  );


  or

  (
    g2199_n,
    g2198_n,
    g2195_p
  );


  or

  (
    g2200_n,
    g2199_n,
    g2197_p
  );


  and

  (
    g2201_p,
    g2111_n_spl_00,
    n4683_lo_p_spl_100
  );


  and

  (
    g2202_p,
    g2201_p,
    n4671_lo_p_spl_100
  );


  and

  (
    g2203_p,
    g2162_n_spl_00,
    n4683_lo_n_spl_100
  );


  and

  (
    g2204_p,
    g2203_p,
    n4671_lo_p_spl_100
  );


  and

  (
    g2205_p,
    n4683_lo_p_spl_100,
    n2811_lo_p_spl_
  );


  and

  (
    g2206_p,
    g2205_p,
    n4671_lo_n_spl_100
  );


  and

  (
    g2207_p,
    n4683_lo_n_spl_100,
    n2823_lo_p_spl_
  );


  and

  (
    g2208_p,
    g2207_p,
    n4671_lo_n_spl_100
  );


  or

  (
    g2209_n,
    g2204_p,
    g2202_p
  );


  or

  (
    g2210_n,
    g2209_n,
    g2206_p
  );


  or

  (
    g2211_n,
    g2210_n,
    g2208_p
  );


  and

  (
    g2212_p,
    g2119_n_spl_00,
    n4683_lo_p_spl_101
  );


  and

  (
    g2213_p,
    g2212_p,
    n4671_lo_p_spl_101
  );


  and

  (
    g2214_p,
    g2170_n_spl_00,
    n4683_lo_n_spl_101
  );


  and

  (
    g2215_p,
    g2214_p,
    n4671_lo_p_spl_101
  );


  and

  (
    g2216_p,
    n4683_lo_p_spl_101,
    n3075_lo_p_spl_
  );


  and

  (
    g2217_p,
    g2216_p,
    n4671_lo_n_spl_101
  );


  and

  (
    g2218_p,
    n4683_lo_n_spl_101,
    n3087_lo_p_spl_
  );


  and

  (
    g2219_p,
    g2218_p,
    n4671_lo_n_spl_101
  );


  or

  (
    g2220_n,
    g2215_p,
    g2213_p
  );


  or

  (
    g2221_n,
    g2220_n,
    g2217_p
  );


  or

  (
    g2222_n,
    g2221_n,
    g2219_p
  );


  and

  (
    g2223_p,
    g2127_n_spl_00,
    n4683_lo_p_spl_110
  );


  and

  (
    g2224_p,
    g2223_p,
    n4671_lo_p_spl_110
  );


  and

  (
    g2225_p,
    g2178_n_spl_00,
    n4683_lo_n_spl_110
  );


  and

  (
    g2226_p,
    g2225_p,
    n4671_lo_p_spl_110
  );


  and

  (
    g2227_p,
    n4683_lo_p_spl_110,
    n3039_lo_p_spl_
  );


  and

  (
    g2228_p,
    g2227_p,
    n4671_lo_n_spl_110
  );


  and

  (
    g2229_p,
    n4683_lo_n_spl_110,
    n2787_lo_p_spl_
  );


  and

  (
    g2230_p,
    g2229_p,
    n4671_lo_n_spl_110
  );


  or

  (
    g2231_n,
    g2226_p,
    g2224_p
  );


  or

  (
    g2232_n,
    g2231_n,
    g2228_p
  );


  or

  (
    g2233_n,
    g2232_n,
    g2230_p
  );


  and

  (
    g2234_p,
    g2111_n_spl_00,
    n4695_lo_p_spl_100
  );


  and

  (
    g2235_p,
    g2234_p,
    n4707_lo_p_spl_100
  );


  and

  (
    g2236_p,
    g2162_n_spl_00,
    n4695_lo_n_spl_100
  );


  and

  (
    g2237_p,
    g2236_p,
    n4707_lo_p_spl_100
  );


  and

  (
    g2238_p,
    n4695_lo_p_spl_100,
    n2811_lo_p_spl_
  );


  and

  (
    g2239_p,
    g2238_p,
    n4707_lo_n_spl_100
  );


  and

  (
    g2240_p,
    n4695_lo_n_spl_100,
    n2823_lo_p_spl_
  );


  and

  (
    g2241_p,
    g2240_p,
    n4707_lo_n_spl_100
  );


  or

  (
    g2242_n,
    g2237_p,
    g2235_p
  );


  or

  (
    g2243_n,
    g2242_n,
    g2239_p
  );


  or

  (
    g2244_n,
    g2243_n,
    g2241_p
  );


  and

  (
    g2245_p,
    g2119_n_spl_00,
    n4695_lo_p_spl_101
  );


  and

  (
    g2246_p,
    g2245_p,
    n4707_lo_p_spl_101
  );


  and

  (
    g2247_p,
    g2170_n_spl_00,
    n4695_lo_n_spl_101
  );


  and

  (
    g2248_p,
    g2247_p,
    n4707_lo_p_spl_101
  );


  and

  (
    g2249_p,
    n4695_lo_p_spl_101,
    n3075_lo_p_spl_
  );


  and

  (
    g2250_p,
    g2249_p,
    n4707_lo_n_spl_101
  );


  and

  (
    g2251_p,
    n4695_lo_n_spl_101,
    n3087_lo_p_spl_
  );


  and

  (
    g2252_p,
    g2251_p,
    n4707_lo_n_spl_101
  );


  or

  (
    g2253_n,
    g2248_p,
    g2246_p
  );


  or

  (
    g2254_n,
    g2253_n,
    g2250_p
  );


  or

  (
    g2255_n,
    g2254_n,
    g2252_p
  );


  and

  (
    g2256_p,
    g2127_n_spl_00,
    n4695_lo_p_spl_110
  );


  and

  (
    g2257_p,
    g2256_p,
    n4707_lo_p_spl_110
  );


  and

  (
    g2258_p,
    g2178_n_spl_00,
    n4695_lo_n_spl_110
  );


  and

  (
    g2259_p,
    g2258_p,
    n4707_lo_p_spl_110
  );


  and

  (
    g2260_p,
    n4695_lo_p_spl_110,
    n3039_lo_p_spl_
  );


  and

  (
    g2261_p,
    g2260_p,
    n4707_lo_n_spl_110
  );


  and

  (
    g2262_p,
    n4695_lo_n_spl_110,
    n2787_lo_p_spl_
  );


  and

  (
    g2263_p,
    g2262_p,
    n4707_lo_n_spl_110
  );


  or

  (
    g2264_n,
    g2259_p,
    g2257_p
  );


  or

  (
    g2265_n,
    g2264_n,
    g2261_p
  );


  or

  (
    g2266_n,
    g2265_n,
    g2263_p
  );


  and

  (
    g2267_p,
    g2127_n_spl_0,
    n4503_lo_p_spl_011
  );


  and

  (
    g2268_p,
    g2267_p,
    n4515_lo_p_spl_011
  );


  and

  (
    g2269_p,
    g2178_n_spl_0,
    n4503_lo_n_spl_011
  );


  and

  (
    g2270_p,
    g2269_p,
    n4515_lo_p_spl_011
  );


  and

  (
    g2271_p,
    n4503_lo_p_spl_011,
    n3651_lo_p_spl_
  );


  and

  (
    g2272_p,
    g2271_p,
    n4515_lo_n_spl_011
  );


  and

  (
    g2273_p,
    n4503_lo_n_spl_011,
    n3531_lo_p_spl_
  );


  and

  (
    g2274_p,
    g2273_p,
    n4515_lo_n_spl_011
  );


  or

  (
    g2275_n,
    g2270_p,
    g2268_p
  );


  or

  (
    g2276_n,
    g2275_n,
    g2272_p
  );


  or

  (
    g2277_n,
    g2276_n,
    g2274_p
  );


  and

  (
    g2278_p,
    g2277_n,
    n3375_lo_p_spl_010
  );


  and

  (
    g2279_p,
    g2119_n_spl_0,
    n4503_lo_p_spl_100
  );


  and

  (
    g2280_p,
    g2279_p,
    n4515_lo_p_spl_100
  );


  and

  (
    g2281_p,
    g2170_n_spl_0,
    n4503_lo_n_spl_100
  );


  and

  (
    g2282_p,
    g2281_p,
    n4515_lo_p_spl_100
  );


  and

  (
    g2283_p,
    n4503_lo_p_spl_100,
    n3627_lo_p_spl_
  );


  and

  (
    g2284_p,
    g2283_p,
    n4515_lo_n_spl_100
  );


  and

  (
    g2285_p,
    n4503_lo_n_spl_100,
    n3507_lo_p_spl_
  );


  and

  (
    g2286_p,
    g2285_p,
    n4515_lo_n_spl_100
  );


  or

  (
    g2287_n,
    g2282_p,
    g2280_p
  );


  or

  (
    g2288_n,
    g2287_n,
    g2284_p
  );


  or

  (
    g2289_n,
    g2288_n,
    g2286_p
  );


  and

  (
    g2290_p,
    g2289_n,
    n3375_lo_p_spl_011
  );


  and

  (
    g2291_p,
    g2111_n_spl_0,
    n4503_lo_p_spl_101
  );


  and

  (
    g2292_p,
    g2291_p,
    n4515_lo_p_spl_101
  );


  and

  (
    g2293_p,
    g2162_n_spl_0,
    n4503_lo_n_spl_101
  );


  and

  (
    g2294_p,
    g2293_p,
    n4515_lo_p_spl_101
  );


  and

  (
    g2295_p,
    n4503_lo_p_spl_101,
    n3615_lo_p_spl_
  );


  and

  (
    g2296_p,
    g2295_p,
    n4515_lo_n_spl_101
  );


  and

  (
    g2297_p,
    n4503_lo_n_spl_101,
    n3495_lo_p_spl_
  );


  and

  (
    g2298_p,
    g2297_p,
    n4515_lo_n_spl_101
  );


  or

  (
    g2299_n,
    g2294_p,
    g2292_p
  );


  or

  (
    g2300_n,
    g2299_n,
    g2296_p
  );


  or

  (
    g2301_n,
    g2300_n,
    g2298_p
  );


  and

  (
    g2302_p,
    g2301_n,
    n3375_lo_p_spl_011
  );


  and

  (
    g2303_p,
    g2103_n_spl_0,
    n4503_lo_p_spl_110
  );


  and

  (
    g2304_p,
    g2303_p,
    n4515_lo_p_spl_110
  );


  and

  (
    g2305_p,
    g2154_n_spl_0,
    n4503_lo_n_spl_110
  );


  and

  (
    g2306_p,
    g2305_p,
    n4515_lo_p_spl_110
  );


  and

  (
    g2307_p,
    n4503_lo_p_spl_110,
    n3603_lo_p_spl_
  );


  and

  (
    g2308_p,
    g2307_p,
    n4515_lo_n_spl_110
  );


  and

  (
    g2309_p,
    n4503_lo_n_spl_110,
    n3483_lo_p_spl_
  );


  and

  (
    g2310_p,
    g2309_p,
    n4515_lo_n_spl_110
  );


  or

  (
    g2311_n,
    g2306_p,
    g2304_p
  );


  or

  (
    g2312_n,
    g2311_n,
    g2308_p
  );


  or

  (
    g2313_n,
    g2312_n,
    g2310_p
  );


  and

  (
    g2314_p,
    g2313_n,
    n3375_lo_p_spl_100
  );


  and

  (
    g2315_p,
    g2127_n_spl_1,
    n4527_lo_p_spl_011
  );


  and

  (
    g2316_p,
    g2315_p,
    n4539_lo_p_spl_011
  );


  and

  (
    g2317_p,
    g2178_n_spl_1,
    n4527_lo_n_spl_011
  );


  and

  (
    g2318_p,
    g2317_p,
    n4539_lo_p_spl_011
  );


  and

  (
    g2319_p,
    n4527_lo_p_spl_011,
    n3651_lo_p_spl_
  );


  and

  (
    g2320_p,
    g2319_p,
    n4539_lo_n_spl_011
  );


  and

  (
    g2321_p,
    n4527_lo_n_spl_011,
    n3531_lo_p_spl_
  );


  and

  (
    g2322_p,
    g2321_p,
    n4539_lo_n_spl_011
  );


  or

  (
    g2323_n,
    g2318_p,
    g2316_p
  );


  or

  (
    g2324_n,
    g2323_n,
    g2320_p
  );


  or

  (
    g2325_n,
    g2324_n,
    g2322_p
  );


  and

  (
    g2326_p,
    g2325_n,
    n3375_lo_p_spl_100
  );


  and

  (
    g2327_p,
    g2119_n_spl_1,
    n4527_lo_p_spl_100
  );


  and

  (
    g2328_p,
    g2327_p,
    n4539_lo_p_spl_100
  );


  and

  (
    g2329_p,
    g2170_n_spl_1,
    n4527_lo_n_spl_100
  );


  and

  (
    g2330_p,
    g2329_p,
    n4539_lo_p_spl_100
  );


  and

  (
    g2331_p,
    n4527_lo_p_spl_100,
    n3627_lo_p_spl_
  );


  and

  (
    g2332_p,
    g2331_p,
    n4539_lo_n_spl_100
  );


  and

  (
    g2333_p,
    n4527_lo_n_spl_100,
    n3507_lo_p_spl_
  );


  and

  (
    g2334_p,
    g2333_p,
    n4539_lo_n_spl_100
  );


  or

  (
    g2335_n,
    g2330_p,
    g2328_p
  );


  or

  (
    g2336_n,
    g2335_n,
    g2332_p
  );


  or

  (
    g2337_n,
    g2336_n,
    g2334_p
  );


  and

  (
    g2338_p,
    g2337_n,
    n3375_lo_p_spl_101
  );


  and

  (
    g2339_p,
    g2111_n_spl_1,
    n4527_lo_p_spl_101
  );


  and

  (
    g2340_p,
    g2339_p,
    n4539_lo_p_spl_101
  );


  and

  (
    g2341_p,
    g2162_n_spl_1,
    n4527_lo_n_spl_101
  );


  and

  (
    g2342_p,
    g2341_p,
    n4539_lo_p_spl_101
  );


  and

  (
    g2343_p,
    n4527_lo_p_spl_101,
    n3615_lo_p_spl_
  );


  and

  (
    g2344_p,
    g2343_p,
    n4539_lo_n_spl_101
  );


  and

  (
    g2345_p,
    n4527_lo_n_spl_101,
    n3495_lo_p_spl_
  );


  and

  (
    g2346_p,
    g2345_p,
    n4539_lo_n_spl_101
  );


  or

  (
    g2347_n,
    g2342_p,
    g2340_p
  );


  or

  (
    g2348_n,
    g2347_n,
    g2344_p
  );


  or

  (
    g2349_n,
    g2348_n,
    g2346_p
  );


  and

  (
    g2350_p,
    g2349_n,
    n3375_lo_p_spl_101
  );


  and

  (
    g2351_p,
    g2103_n_spl_1,
    n4527_lo_p_spl_110
  );


  and

  (
    g2352_p,
    g2351_p,
    n4539_lo_p_spl_110
  );


  and

  (
    g2353_p,
    g2154_n_spl_1,
    n4527_lo_n_spl_110
  );


  and

  (
    g2354_p,
    g2353_p,
    n4539_lo_p_spl_110
  );


  and

  (
    g2355_p,
    n4527_lo_p_spl_110,
    n3603_lo_p_spl_
  );


  and

  (
    g2356_p,
    g2355_p,
    n4539_lo_n_spl_110
  );


  and

  (
    g2357_p,
    n4527_lo_n_spl_110,
    n3483_lo_p_spl_
  );


  and

  (
    g2358_p,
    g2357_p,
    n4539_lo_n_spl_110
  );


  or

  (
    g2359_n,
    g2354_p,
    g2352_p
  );


  or

  (
    g2360_n,
    g2359_n,
    g2356_p
  );


  or

  (
    g2361_n,
    g2360_n,
    g2358_p
  );


  and

  (
    g2362_p,
    g2361_n,
    n3375_lo_p_spl_110
  );


  and

  (
    g2363_p,
    G4420_o2_n,
    G4180_o2_n
  );


  and

  (
    g2364_p,
    G4420_o2_p,
    G4180_o2_p
  );


  or

  (
    g2365_n,
    g2364_p,
    g2363_p
  );


  or

  (
    g2366_n,
    g2365_n_spl_,
    n4719_lo_n_spl_101
  );


  or

  (
    g2367_n,
    g2366_n,
    n4731_lo_n_spl_101
  );


  or

  (
    g2368_n,
    G5126_o2_p,
    G5138_o2_n
  );


  or

  (
    g2369_n,
    G5144_o2_p,
    G5111_o2_n
  );


  and

  (
    g2370_p,
    g2369_n,
    g2368_n
  );


  or

  (
    g2371_n,
    g2370_p_spl_,
    n4719_lo_p_spl_1101
  );


  or

  (
    g2372_n,
    g2371_n,
    n4731_lo_n_spl_101
  );


  or

  (
    g2373_n,
    n4719_lo_n_spl_101,
    n3219_lo_n
  );


  or

  (
    g2374_n,
    g2373_n,
    n4731_lo_p_spl_1101
  );


  or

  (
    g2375_n,
    n4731_lo_p_spl_1110,
    n4719_lo_p_spl_1110
  );


  and

  (
    g2376_p,
    g2372_n,
    g2367_n
  );


  and

  (
    g2377_p,
    g2376_p,
    g2374_n
  );


  and

  (
    g2378_p,
    g2377_p,
    g2375_n_spl_
  );


  and

  (
    g2379_p,
    G4417_o2_p,
    G4504_o2_n
  );


  and

  (
    g2380_p,
    G4417_o2_n,
    G4504_o2_p
  );


  or

  (
    g2381_n,
    g2380_p,
    g2379_p
  );


  or

  (
    g2382_n,
    g2381_n_spl_,
    n4719_lo_n_spl_110
  );


  or

  (
    g2383_n,
    g2382_n,
    n4731_lo_n_spl_110
  );


  or

  (
    g2384_n,
    G5123_o2_n,
    G5135_o2_n
  );


  or

  (
    g2385_n,
    G5142_o2_p,
    G5108_o2_p
  );


  and

  (
    g2386_p,
    g2385_n,
    g2384_n
  );


  or

  (
    g2387_n,
    g2386_p_spl_,
    n4719_lo_p_spl_1110
  );


  or

  (
    g2388_n,
    g2387_n,
    n4731_lo_n_spl_110
  );


  or

  (
    g2389_n,
    n4719_lo_n_spl_110,
    n3195_lo_n
  );


  or

  (
    g2390_n,
    g2389_n,
    n4731_lo_p_spl_1110
  );


  and

  (
    g2391_p,
    g2388_n,
    g2383_n
  );


  and

  (
    g2392_p,
    g2391_p,
    g2390_n
  );


  and

  (
    g2393_p,
    g2392_p,
    g2375_n_spl_
  );


  and

  (
    g2394_p,
    g2365_n_spl_,
    n4719_lo_p_spl_1111
  );


  and

  (
    g2395_p,
    g2370_p_spl_,
    n4719_lo_n_spl_111
  );


  or

  (
    g2396_n,
    g2395_p,
    g2394_p
  );


  and

  (
    g2397_p,
    g2396_n,
    n4731_lo_p_spl_1111
  );


  and

  (
    g2398_p,
    n4731_lo_n_spl_111,
    n3051_lo_p
  );


  or

  (
    g2399_n,
    g2398_p,
    g2397_p
  );


  and

  (
    g2400_p,
    g2399_n_spl_0,
    n4683_lo_p_spl_111
  );


  and

  (
    g2401_p,
    g2400_p,
    n4671_lo_p_spl_111
  );


  and

  (
    g2402_p,
    g2381_n_spl_,
    n4719_lo_p_spl_1111
  );


  and

  (
    g2403_p,
    g2386_p_spl_,
    n4719_lo_n_spl_111
  );


  or

  (
    g2404_n,
    g2403_p,
    g2402_p
  );


  and

  (
    g2405_p,
    g2404_n,
    n4731_lo_p_spl_1111
  );


  and

  (
    g2406_p,
    n4731_lo_n_spl_111,
    n3063_lo_p
  );


  or

  (
    g2407_n,
    g2406_p,
    g2405_p
  );


  and

  (
    g2408_p,
    g2407_n_spl_0,
    n4683_lo_n_spl_111
  );


  and

  (
    g2409_p,
    g2408_p,
    n4671_lo_p_spl_111
  );


  and

  (
    g2410_p,
    n4683_lo_p_spl_111,
    n2655_lo_p_spl_
  );


  and

  (
    g2411_p,
    g2410_p,
    n4671_lo_n_spl_111
  );


  and

  (
    g2412_p,
    n4683_lo_n_spl_111,
    n2883_lo_p_spl_
  );


  and

  (
    g2413_p,
    g2412_p,
    n4671_lo_n_spl_111
  );


  or

  (
    g2414_n,
    g2409_p,
    g2401_p
  );


  or

  (
    g2415_n,
    g2414_n,
    g2411_p
  );


  or

  (
    g2416_n,
    g2415_n,
    g2413_p
  );


  and

  (
    g2417_p,
    g2399_n_spl_0,
    n4695_lo_p_spl_111
  );


  and

  (
    g2418_p,
    g2417_p,
    n4707_lo_p_spl_111
  );


  and

  (
    g2419_p,
    g2407_n_spl_0,
    n4695_lo_n_spl_111
  );


  and

  (
    g2420_p,
    g2419_p,
    n4707_lo_p_spl_111
  );


  and

  (
    g2421_p,
    n4695_lo_p_spl_111,
    n2655_lo_p_spl_
  );


  and

  (
    g2422_p,
    g2421_p,
    n4707_lo_n_spl_111
  );


  and

  (
    g2423_p,
    n4695_lo_n_spl_111,
    n2883_lo_p_spl_
  );


  and

  (
    g2424_p,
    g2423_p,
    n4707_lo_n_spl_111
  );


  or

  (
    g2425_n,
    g2420_p,
    g2418_p
  );


  or

  (
    g2426_n,
    g2425_n,
    g2422_p
  );


  or

  (
    g2427_n,
    g2426_n,
    g2424_p
  );


  and

  (
    g2428_p,
    g2399_n_spl_1,
    n4503_lo_p_spl_111
  );


  and

  (
    g2429_p,
    g2428_p,
    n4515_lo_p_spl_111
  );


  and

  (
    g2430_p,
    g2407_n_spl_1,
    n4503_lo_n_spl_111
  );


  and

  (
    g2431_p,
    g2430_p,
    n4515_lo_p_spl_111
  );


  and

  (
    g2432_p,
    n4503_lo_p_spl_111,
    n3543_lo_p_spl_
  );


  and

  (
    g2433_p,
    g2432_p,
    n4515_lo_n_spl_111
  );


  and

  (
    g2434_p,
    n4503_lo_n_spl_111,
    n3555_lo_p_spl_
  );


  and

  (
    g2435_p,
    g2434_p,
    n4515_lo_n_spl_111
  );


  or

  (
    g2436_n,
    g2431_p,
    g2429_p
  );


  or

  (
    g2437_n,
    g2436_n,
    g2433_p
  );


  or

  (
    g2438_n,
    g2437_n,
    g2435_p
  );


  and

  (
    g2439_p,
    g2438_n,
    n3375_lo_p_spl_110
  );


  and

  (
    g2440_p,
    g2399_n_spl_1,
    n4527_lo_p_spl_111
  );


  and

  (
    g2441_p,
    g2440_p,
    n4539_lo_p_spl_111
  );


  and

  (
    g2442_p,
    g2407_n_spl_1,
    n4527_lo_n_spl_111
  );


  and

  (
    g2443_p,
    g2442_p,
    n4539_lo_p_spl_111
  );


  and

  (
    g2444_p,
    n4527_lo_p_spl_111,
    n3543_lo_p_spl_
  );


  and

  (
    g2445_p,
    g2444_p,
    n4539_lo_n_spl_111
  );


  and

  (
    g2446_p,
    n4527_lo_n_spl_111,
    n3555_lo_p_spl_
  );


  and

  (
    g2447_p,
    g2446_p,
    n4539_lo_n_spl_111
  );


  or

  (
    g2448_n,
    g2443_p,
    g2441_p
  );


  or

  (
    g2449_n,
    g2448_n,
    g2445_p
  );


  or

  (
    g2450_n,
    g2449_n,
    g2447_p
  );


  and

  (
    g2451_p,
    g2450_n,
    n3375_lo_p_spl_111
  );


  and

  (
    g2452_p,
    G3132_o2_n,
    G3291_o2_n
  );


  or

  (
    g2452_n,
    G3132_o2_p,
    G3291_o2_p
  );


  and

  (
    g2453_p,
    n2968_inv_n_spl_00,
    n4308_lo_buf_o2_p_spl_00
  );


  or

  (
    g2453_n,
    n2968_inv_p_spl_000,
    n4308_lo_buf_o2_n_spl_0
  );


  and

  (
    g2454_p,
    g2453_p,
    G1876_o2_p
  );


  or

  (
    g2454_n,
    g2453_n,
    G1876_o2_n
  );


  and

  (
    g2455_p,
    n2974_inv_n_spl_00,
    n4308_lo_buf_o2_p_spl_00
  );


  or

  (
    g2455_n,
    n2974_inv_p_spl_00,
    n4308_lo_buf_o2_n_spl_0
  );


  and

  (
    g2456_p,
    g2455_p,
    G2293_o2_n
  );


  or

  (
    g2456_n,
    g2455_n,
    G2293_o2_p
  );


  and

  (
    g2457_p,
    g2456_n,
    g2454_n
  );


  or

  (
    g2457_n,
    g2456_p,
    g2454_p
  );


  and

  (
    g2458_p,
    n3121_inv_n_spl_00,
    G1873_o2_p_spl_
  );


  or

  (
    g2458_n,
    n3121_inv_p_spl_000,
    G1873_o2_n_spl_
  );


  and

  (
    g2459_p,
    n3124_inv_n_spl_00,
    G1873_o2_n_spl_
  );


  or

  (
    g2459_n,
    n3124_inv_p_spl_00,
    G1873_o2_p_spl_
  );


  and

  (
    g2460_p,
    g2459_n,
    g2458_n
  );


  or

  (
    g2460_n,
    g2459_p,
    g2458_p
  );


  and

  (
    g2461_p,
    g2460_p,
    n4308_lo_buf_o2_n_spl_1
  );


  or

  (
    g2461_n,
    g2460_n,
    n4308_lo_buf_o2_p_spl_0
  );


  and

  (
    g2462_p,
    g2461_n,
    g2457_p
  );


  or

  (
    g2462_n,
    g2461_p,
    g2457_n
  );


  and

  (
    g2463_p,
    n6999_o2_p,
    n6955_o2_p_spl_
  );


  or

  (
    g2463_n,
    n6999_o2_n,
    n6955_o2_n_spl_
  );


  and

  (
    g2464_p,
    g2463_p,
    n6954_o2_p_spl_00
  );


  or

  (
    g2464_n,
    g2463_n,
    n6954_o2_n_spl_00
  );


  and

  (
    g2465_p,
    g2464_p,
    n7387_o2_p_spl_00
  );


  or

  (
    g2465_n,
    g2464_n,
    n7387_o2_n_spl_00
  );


  and

  (
    g2466_p,
    g2465_p,
    G3495_o2_p_spl_00
  );


  or

  (
    g2466_n,
    g2465_n,
    G3495_o2_n_spl_00
  );


  and

  (
    g2467_p,
    n7155_o2_n,
    n6957_o2_p_spl_
  );


  or

  (
    g2467_n,
    n7155_o2_p,
    n6957_o2_n_spl_
  );


  and

  (
    g2468_p,
    g2467_p,
    n6956_o2_p_spl_00
  );


  or

  (
    g2468_n,
    g2467_n,
    n6956_o2_n_spl_00
  );


  and

  (
    g2469_p,
    g2468_p,
    n7386_o2_p_spl_00
  );


  or

  (
    g2469_n,
    g2468_n,
    n7386_o2_n_spl_00
  );


  and

  (
    g2470_p,
    g2469_p,
    G3621_o2_p_spl_00
  );


  or

  (
    g2470_n,
    g2469_n,
    G3621_o2_n_spl_00
  );


  and

  (
    g2471_p,
    G2404_o2_p_spl_0,
    n4296_lo_buf_o2_p_spl_0
  );


  or

  (
    g2471_n,
    G2404_o2_n_spl_0,
    n4296_lo_buf_o2_n_spl_0
  );


  and

  (
    g2472_p,
    G3495_o2_p_spl_00,
    n7431_o2_p
  );


  or

  (
    g2472_n,
    G3495_o2_n_spl_00,
    n7431_o2_n
  );


  and

  (
    g2473_p,
    G3495_o2_p_spl_0,
    n7387_o2_p_spl_00
  );


  or

  (
    g2473_n,
    G3495_o2_n_spl_0,
    n7387_o2_n_spl_00
  );


  and

  (
    g2474_p,
    g2473_p,
    n6974_o2_p
  );


  or

  (
    g2474_n,
    g2473_n,
    n6974_o2_n
  );


  and

  (
    g2475_p,
    G3495_o2_p_spl_1,
    n6954_o2_p_spl_00
  );


  or

  (
    g2475_n,
    G3495_o2_n_spl_1,
    n6954_o2_n_spl_00
  );


  and

  (
    g2476_p,
    g2475_p,
    n6888_o2_p
  );


  or

  (
    g2476_n,
    g2475_n,
    n6888_o2_n
  );


  and

  (
    g2477_p,
    g2476_p,
    n7387_o2_p_spl_01
  );


  or

  (
    g2477_n,
    g2476_n,
    n7387_o2_n_spl_01
  );


  and

  (
    g2478_p,
    n6955_o2_p_spl_,
    n6954_o2_p_spl_01
  );


  or

  (
    g2478_n,
    n6955_o2_n_spl_,
    n6954_o2_n_spl_01
  );


  and

  (
    g2479_p,
    g2478_p,
    G3495_o2_p_spl_1
  );


  or

  (
    g2479_n,
    g2478_n,
    G3495_o2_n_spl_1
  );


  and

  (
    g2480_p,
    g2479_p,
    n6936_o2_p
  );


  or

  (
    g2480_n,
    g2479_n,
    n6936_o2_n
  );


  and

  (
    g2481_p,
    g2480_p,
    n7387_o2_p_spl_01
  );


  or

  (
    g2481_n,
    g2480_n,
    n7387_o2_n_spl_01
  );


  and

  (
    g2482_p,
    g2472_n,
    g2471_n
  );


  or

  (
    g2482_n,
    g2472_p,
    g2471_p
  );


  and

  (
    g2483_p,
    g2482_p,
    g2474_n
  );


  or

  (
    g2483_n,
    g2482_n,
    g2474_p
  );


  and

  (
    g2484_p,
    g2483_p,
    g2477_n
  );


  or

  (
    g2484_n,
    g2483_n,
    g2477_p
  );


  and

  (
    g2485_p,
    g2484_p,
    g2481_n
  );


  or

  (
    g2485_n,
    g2484_n,
    g2481_p
  );


  and

  (
    g2486_p,
    G2466_o2_p_spl_0,
    n4368_lo_buf_o2_p_spl_0
  );


  or

  (
    g2486_n,
    G2466_o2_n_spl_0,
    n4368_lo_buf_o2_n_spl_0
  );


  and

  (
    g2487_p,
    G3621_o2_p_spl_00,
    n7430_o2_p
  );


  or

  (
    g2487_n,
    G3621_o2_n_spl_00,
    n7430_o2_n
  );


  and

  (
    g2488_p,
    G3621_o2_p_spl_0,
    n7386_o2_p_spl_00
  );


  or

  (
    g2488_n,
    G3621_o2_n_spl_0,
    n7386_o2_n_spl_00
  );


  and

  (
    g2489_p,
    g2488_p,
    n6975_o2_p
  );


  or

  (
    g2489_n,
    g2488_n,
    n6975_o2_n
  );


  and

  (
    g2490_p,
    G3621_o2_p_spl_1,
    n6956_o2_p_spl_00
  );


  or

  (
    g2490_n,
    G3621_o2_n_spl_1,
    n6956_o2_n_spl_00
  );


  and

  (
    g2491_p,
    g2490_p,
    n6889_o2_p
  );


  or

  (
    g2491_n,
    g2490_n,
    n6889_o2_n
  );


  and

  (
    g2492_p,
    g2491_p,
    n7386_o2_p_spl_01
  );


  or

  (
    g2492_n,
    g2491_n,
    n7386_o2_n_spl_01
  );


  and

  (
    g2493_p,
    n6957_o2_p_spl_,
    n6956_o2_p_spl_01
  );


  or

  (
    g2493_n,
    n6957_o2_n_spl_,
    n6956_o2_n_spl_01
  );


  and

  (
    g2494_p,
    g2493_p,
    G3621_o2_p_spl_1
  );


  or

  (
    g2494_n,
    g2493_n,
    G3621_o2_n_spl_1
  );


  and

  (
    g2495_p,
    g2494_p,
    n6958_o2_n
  );


  or

  (
    g2495_n,
    g2494_n,
    n6958_o2_p
  );


  and

  (
    g2496_p,
    g2495_p,
    n7386_o2_p_spl_01
  );


  or

  (
    g2496_n,
    g2495_n,
    n7386_o2_n_spl_01
  );


  and

  (
    g2497_p,
    g2487_n,
    g2486_n
  );


  or

  (
    g2497_n,
    g2487_p,
    g2486_p
  );


  and

  (
    g2498_p,
    g2497_p,
    g2489_n
  );


  or

  (
    g2498_n,
    g2497_n,
    g2489_p
  );


  and

  (
    g2499_p,
    g2498_p,
    g2492_n
  );


  or

  (
    g2499_n,
    g2498_n,
    g2492_p
  );


  and

  (
    g2500_p,
    g2499_p,
    g2496_n
  );


  or

  (
    g2500_n,
    g2499_n,
    g2496_p
  );


  and

  (
    g2501_p,
    n2968_inv_n_spl_00,
    n6772_o2_n_spl_0
  );


  or

  (
    g2501_n,
    n2968_inv_p_spl_000,
    n6772_o2_p_spl_0
  );


  and

  (
    g2502_p,
    n2974_inv_n_spl_00,
    n6772_o2_p_spl_0
  );


  or

  (
    g2502_n,
    n2974_inv_p_spl_00,
    n6772_o2_n_spl_0
  );


  and

  (
    g2503_p,
    g2502_n,
    g2501_n
  );


  or

  (
    g2503_n,
    g2502_p,
    g2501_p
  );


  and

  (
    g2504_p,
    G2269_o2_n,
    G1835_o2_n
  );


  or

  (
    g2504_n,
    G2269_o2_p,
    G1835_o2_p
  );


  and

  (
    g2505_p,
    G1512_o2_p,
    G2921_o2_n
  );


  or

  (
    g2505_n,
    G1512_o2_n,
    G2921_o2_p
  );


  and

  (
    g2506_p,
    G3135_o2_p,
    G1344_o2_n
  );


  or

  (
    g2506_n,
    G3135_o2_n,
    G1344_o2_p
  );


  and

  (
    g2507_p,
    g2506_n,
    g2505_n
  );


  or

  (
    g2507_n,
    g2506_p,
    g2505_p
  );


  and

  (
    g2508_p,
    G2424_o2_p_spl_,
    n4320_lo_buf_o2_p_spl_
  );


  or

  (
    g2508_n,
    G2424_o2_n,
    n4320_lo_buf_o2_n
  );


  and

  (
    g2509_p,
    G1821_o2_p_spl_,
    n4053_lo_p_spl_00
  );


  or

  (
    g2509_n,
    G1821_o2_n,
    n4053_lo_n_spl_
  );


  and

  (
    g2510_p,
    G1060_o2_n_spl_,
    n4065_lo_p
  );


  or

  (
    g2510_n,
    G1060_o2_p,
    n4065_lo_n
  );


  and

  (
    g2511_p,
    g2510_n,
    g2509_n
  );


  or

  (
    g2511_n,
    g2510_p,
    g2509_p
  );


  and

  (
    g2512_p,
    G1734_o2_p_spl_,
    n3753_lo_p_spl_00
  );


  or

  (
    g2512_n,
    G1734_o2_n,
    n3753_lo_n_spl_
  );


  and

  (
    g2513_p,
    G963_o2_n_spl_,
    n3765_lo_p
  );


  or

  (
    g2513_n,
    G963_o2_p,
    n3765_lo_n
  );


  and

  (
    g2514_p,
    g2513_n,
    g2512_n
  );


  or

  (
    g2514_n,
    g2513_p,
    g2512_p
  );


  and

  (
    g2515_p,
    n4164_lo_buf_o2_p_spl_,
    G1815_o2_p_spl_0
  );


  or

  (
    g2515_n,
    n4164_lo_buf_o2_n,
    G1815_o2_n_spl_
  );


  and

  (
    g2516_p,
    n4176_lo_buf_o2_p_spl_,
    n2662_inv_n_spl_
  );


  or

  (
    g2516_n,
    n4176_lo_buf_o2_n,
    n2662_inv_p_spl_0
  );


  and

  (
    g2517_p,
    g2516_n,
    g2515_n
  );


  or

  (
    g2517_n,
    g2516_p,
    g2515_p
  );


  and

  (
    g2518_p,
    n7136_o2_p_spl_0,
    n7132_o2_p_spl_00
  );


  and

  (
    g2519_p,
    n7023_o2_p_spl_0,
    n7016_o2_p_spl_00
  );


  or

  (
    g2520_n,
    n7022_o2_n_spl_0,
    n7017_o2_n_spl_00
  );


  or

  (
    g2521_n,
    n7135_o2_n_spl_,
    n7133_o2_n_spl_00
  );


  and

  (
    g2522_p,
    n4272_lo_buf_o2_p_spl_,
    G2386_o2_p_spl_
  );


  or

  (
    g2522_n,
    n4272_lo_buf_o2_n,
    G2386_o2_n
  );


  and

  (
    g2523_p,
    n4404_lo_buf_o2_p_spl_,
    G2454_o2_p_spl_
  );


  or

  (
    g2523_n,
    n4404_lo_buf_o2_n,
    G2454_o2_n
  );


  and

  (
    g2524_p,
    n7384_o2_p_spl_0,
    n7383_o2_n_spl_0
  );


  and

  (
    g2525_p,
    n7384_o2_n_spl_,
    n7383_o2_p_spl_00
  );


  or

  (
    g2526_n,
    g2525_p,
    g2524_p
  );


  and

  (
    g2527_p,
    n7023_o2_p_spl_0,
    n7016_o2_n_spl_0
  );


  and

  (
    g2528_p,
    n7023_o2_n_spl_,
    n7016_o2_p_spl_00
  );


  or

  (
    g2529_n,
    g2528_p,
    g2527_p
  );


  and

  (
    g2530_p,
    n7022_o2_p_spl_0,
    n7017_o2_n_spl_00
  );


  or

  (
    g2530_n,
    n7022_o2_n_spl_0,
    n7017_o2_p_spl_00
  );


  and

  (
    g2531_p,
    n7022_o2_n_spl_,
    n7017_o2_p_spl_00
  );


  or

  (
    g2531_n,
    n7022_o2_p_spl_0,
    n7017_o2_n_spl_01
  );


  and

  (
    g2532_p,
    g2531_n,
    g2530_n
  );


  or

  (
    g2532_n,
    g2531_p,
    g2530_p
  );


  and

  (
    g2533_p,
    n4224_lo_buf_o2_p_spl_00,
    G2379_o2_p_spl_00
  );


  or

  (
    g2533_n,
    n4224_lo_buf_o2_n_spl_0,
    G2379_o2_n_spl_0
  );


  and

  (
    g2534_p,
    G1356_o2_p_spl_,
    G2933_o2_n_spl_
  );


  or

  (
    g2534_n,
    G1356_o2_n_spl_,
    G2933_o2_p_spl_
  );


  and

  (
    g2535_p,
    G1356_o2_n_spl_,
    G2933_o2_p_spl_
  );


  or

  (
    g2535_n,
    G1356_o2_p_spl_,
    G2933_o2_n_spl_
  );


  and

  (
    g2536_p,
    g2535_n,
    g2534_n
  );


  or

  (
    g2536_n,
    g2535_p,
    g2534_p
  );


  and

  (
    g2537_p,
    G1359_o2_p_spl_,
    G2936_o2_n_spl_
  );


  or

  (
    g2537_n,
    G1359_o2_n_spl_,
    G2936_o2_p_spl_
  );


  and

  (
    g2538_p,
    G1359_o2_n_spl_,
    G2936_o2_p_spl_
  );


  or

  (
    g2538_n,
    G1359_o2_p_spl_,
    G2936_o2_n_spl_
  );


  and

  (
    g2539_p,
    g2538_n,
    g2537_n
  );


  or

  (
    g2539_n,
    g2538_p,
    g2537_p
  );


  and

  (
    g2540_p,
    G1398_o2_p_spl_,
    G2975_o2_n_spl_
  );


  or

  (
    g2540_n,
    G1398_o2_n_spl_,
    G2975_o2_p_spl_
  );


  and

  (
    g2541_p,
    G1398_o2_n_spl_,
    G2975_o2_p_spl_
  );


  or

  (
    g2541_n,
    G1398_o2_p_spl_,
    G2975_o2_n_spl_
  );


  and

  (
    g2542_p,
    g2541_n,
    g2540_n
  );


  or

  (
    g2542_n,
    g2541_p,
    g2540_p
  );


  and

  (
    g2543_p,
    G1401_o2_p_spl_,
    G2978_o2_n_spl_
  );


  or

  (
    g2543_n,
    G1401_o2_n_spl_,
    G2978_o2_p_spl_
  );


  and

  (
    g2544_p,
    G1401_o2_n_spl_,
    G2978_o2_p_spl_
  );


  or

  (
    g2544_n,
    G1401_o2_p_spl_,
    G2978_o2_n_spl_
  );


  and

  (
    g2545_p,
    g2544_n,
    g2543_n
  );


  or

  (
    g2545_n,
    g2544_p,
    g2543_p
  );


  and

  (
    g2546_p,
    n4260_lo_buf_o2_p_spl_,
    G2392_o2_p_spl_
  );


  or

  (
    g2546_n,
    n4260_lo_buf_o2_n,
    G2392_o2_n
  );


  and

  (
    g2547_p,
    n4392_lo_buf_o2_p_spl_,
    G2460_o2_p_spl_
  );


  or

  (
    g2547_n,
    n4392_lo_buf_o2_n,
    G2460_o2_n
  );


  and

  (
    g2548_p,
    n4224_lo_buf_o2_p_spl_00,
    G2379_o2_n_spl_0
  );


  or

  (
    g2548_n,
    n4224_lo_buf_o2_n_spl_0,
    G2379_o2_p_spl_00
  );


  and

  (
    g2549_p,
    n4224_lo_buf_o2_n_spl_1,
    G2379_o2_p_spl_0
  );


  or

  (
    g2549_n,
    n4224_lo_buf_o2_p_spl_0,
    G2379_o2_n_spl_1
  );


  and

  (
    g2550_p,
    g2549_n,
    g2548_n
  );


  or

  (
    g2550_n,
    g2549_p,
    g2548_p
  );


  and

  (
    g2551_p,
    n2662_inv_n_spl_,
    n4098_lo_p_spl_
  );


  or

  (
    g2551_n,
    n2662_inv_p_spl_0,
    n4098_lo_n
  );


  and

  (
    g2552_p,
    g2551_n,
    G1815_o2_n_spl_
  );


  or

  (
    g2552_n,
    g2551_p,
    G1815_o2_p_spl_0
  );


  and

  (
    g2553_p,
    G1728_o2_p_spl_,
    n3834_lo_p_spl_
  );


  or

  (
    g2553_n,
    G1728_o2_n,
    n3834_lo_n
  );


  and

  (
    g2554_p,
    n2665_inv_n,
    n3846_lo_p
  );


  or

  (
    g2554_n,
    n2665_inv_p_spl_,
    n3846_lo_n
  );


  and

  (
    g2555_p,
    g2554_n,
    g2553_n
  );


  or

  (
    g2555_n,
    g2554_p,
    g2553_p
  );


  and

  (
    g2556_p,
    n4080_lo_buf_o2_p_spl_00,
    n4002_lo_p_spl_
  );


  or

  (
    g2556_n,
    n4080_lo_buf_o2_n_spl_00,
    n4002_lo_n
  );


  and

  (
    g2557_p,
    n4080_lo_buf_o2_n_spl_00,
    n4014_lo_p
  );


  or

  (
    g2557_n,
    n4080_lo_buf_o2_p_spl_00,
    n4014_lo_n
  );


  and

  (
    g2558_p,
    g2557_n,
    g2556_n
  );


  or

  (
    g2558_n,
    g2557_p,
    g2556_p
  );


  and

  (
    g2559_p,
    n4092_lo_buf_o2_p_spl_00,
    n3702_lo_p_spl_
  );


  or

  (
    g2559_n,
    n4092_lo_buf_o2_n_spl_00,
    n3702_lo_n
  );


  and

  (
    g2560_p,
    n4092_lo_buf_o2_n_spl_00,
    n3714_lo_p
  );


  or

  (
    g2560_n,
    n4092_lo_buf_o2_p_spl_00,
    n3714_lo_n
  );


  and

  (
    g2561_p,
    g2560_n,
    g2559_n
  );


  or

  (
    g2561_n,
    g2560_p,
    g2559_p
  );


  and

  (
    g2562_p,
    n7384_o2_p_spl_0,
    n7383_o2_p_spl_00
  );


  and

  (
    g2563_p,
    G4946_o2_n,
    G3954_o2_n
  );


  or

  (
    g2563_n,
    G4946_o2_p,
    G3954_o2_p
  );


  and

  (
    g2564_p,
    G4234_o2_p,
    G4923_o2_p
  );


  or

  (
    g2564_n,
    G4234_o2_n,
    G4923_o2_n
  );


  and

  (
    g2565_p,
    g2564_n,
    g2563_n
  );


  or

  (
    g2565_n,
    g2564_p,
    g2563_p
  );


  and

  (
    g2566_p,
    g2565_p_spl_,
    g2452_p_spl_0
  );


  or

  (
    g2566_n,
    g2565_n_spl_,
    g2452_n_spl_00
  );


  and

  (
    g2567_p,
    g2565_n_spl_,
    g2452_n_spl_00
  );


  or

  (
    g2567_n,
    g2565_p_spl_,
    g2452_p_spl_0
  );


  and

  (
    g2568_p,
    g2567_n,
    g2566_n
  );


  or

  (
    g2568_n,
    g2567_p,
    g2566_p
  );


  or

  (
    g2569_n,
    g2568_n,
    G3474_o2_p_spl_0
  );


  or

  (
    g2570_n,
    g2568_p,
    G3474_o2_n_spl_
  );


  and

  (
    g2571_p,
    g2570_n,
    g2569_n
  );


  or

  (
    g2572_n,
    g2571_p_spl_,
    g2485_n_spl_0
  );


  or

  (
    g2573_n,
    g2572_n,
    n4488_lo_p_spl_0
  );


  and

  (
    g2574_p,
    G4944_o2_n,
    G3942_o2_n
  );


  or

  (
    g2574_n,
    G4944_o2_p,
    G3942_o2_p
  );


  and

  (
    g2575_p,
    G4231_o2_p,
    G4920_o2_p
  );


  or

  (
    g2575_n,
    G4231_o2_n,
    G4920_o2_n
  );


  and

  (
    g2576_p,
    g2575_n,
    g2574_n
  );


  or

  (
    g2576_n,
    g2575_p,
    g2574_p
  );


  and

  (
    g2577_p,
    g2576_p_spl_,
    g2452_p_spl_1
  );


  or

  (
    g2577_n,
    g2576_n_spl_,
    g2452_n_spl_0
  );


  and

  (
    g2578_p,
    g2576_n_spl_,
    g2452_n_spl_1
  );


  or

  (
    g2578_n,
    g2576_p_spl_,
    g2452_p_spl_1
  );


  and

  (
    g2579_p,
    g2578_n,
    g2577_n
  );


  or

  (
    g2579_n,
    g2578_p,
    g2577_p
  );


  or

  (
    g2580_n,
    g2579_n,
    G3474_o2_p_spl_0
  );


  or

  (
    g2581_n,
    g2579_p,
    G3474_o2_n_spl_
  );


  and

  (
    g2582_p,
    g2581_n,
    g2580_n
  );


  or

  (
    g2583_n,
    g2582_p_spl_,
    g2485_p_spl_
  );


  or

  (
    g2584_n,
    g2583_n,
    n4488_lo_p_spl_0
  );


  and

  (
    g2585_p,
    g2485_p_spl_,
    g2466_n
  );


  or

  (
    g2585_n,
    g2485_n_spl_0,
    g2466_p_spl_
  );


  or

  (
    g2586_n,
    g2585_n,
    g2571_p_spl_
  );


  or

  (
    g2587_n,
    g2586_n,
    n4488_lo_n_spl_0
  );


  or

  (
    g2588_n,
    g2585_p,
    g2582_p_spl_
  );


  or

  (
    g2589_n,
    g2588_n,
    n4488_lo_n_spl_0
  );


  and

  (
    g2590_p,
    g2584_n,
    g2573_n
  );


  and

  (
    g2591_p,
    g2590_p,
    g2587_n
  );


  and

  (
    g2592_p,
    g2591_p,
    g2589_n
  );


  and

  (
    g2593_p,
    G5038_o2_p,
    G5025_o2_n
  );


  or

  (
    g2593_n,
    G5038_o2_n,
    G5025_o2_p
  );


  and

  (
    g2594_p,
    g2593_p_spl_,
    n6954_o2_n_spl_01
  );


  or

  (
    g2594_n,
    g2593_n_spl_,
    n6954_o2_p_spl_01
  );


  and

  (
    g2595_p,
    g2593_n_spl_,
    n6954_o2_p_spl_10
  );


  or

  (
    g2595_n,
    g2593_p_spl_,
    n6954_o2_n_spl_10
  );


  and

  (
    g2596_p,
    g2595_n,
    g2594_n
  );


  or

  (
    g2596_n,
    g2595_p,
    g2594_p
  );


  or

  (
    g2597_n,
    g2596_n,
    n7387_o2_p_spl_1
  );


  or

  (
    g2598_n,
    g2596_p,
    n7387_o2_n_spl_1
  );


  and

  (
    g2599_p,
    g2598_n,
    g2597_n
  );


  and

  (
    g2600_p,
    g2599_p,
    n4488_lo_n_spl_
  );


  and

  (
    g2601_p,
    G5022_o2_p,
    G3969_o2_n
  );


  or

  (
    g2601_n,
    G5022_o2_n,
    G3969_o2_p
  );


  and

  (
    g2602_p,
    G4238_o2_p,
    G4996_o2_n
  );


  or

  (
    g2602_n,
    G4238_o2_n,
    G4996_o2_p
  );


  and

  (
    g2603_p,
    g2602_n,
    g2601_n
  );


  or

  (
    g2603_n,
    g2602_p,
    g2601_p
  );


  and

  (
    g2604_p,
    g2603_p_spl_,
    n6954_o2_n_spl_10
  );


  or

  (
    g2604_n,
    g2603_n_spl_,
    n6954_o2_p_spl_10
  );


  and

  (
    g2605_p,
    g2603_n_spl_,
    n6954_o2_p_spl_1
  );


  or

  (
    g2605_n,
    g2603_p_spl_,
    n6954_o2_n_spl_1
  );


  and

  (
    g2606_p,
    g2605_n,
    g2604_n
  );


  or

  (
    g2606_n,
    g2605_p,
    g2604_p
  );


  and

  (
    g2607_p,
    g2606_p,
    n7387_o2_n_spl_1
  );


  and

  (
    g2608_p,
    g2606_n,
    n7387_o2_p_spl_1
  );


  or

  (
    g2609_n,
    g2608_p,
    g2607_p
  );


  and

  (
    g2610_p,
    g2609_n,
    n4488_lo_p_spl_
  );


  or

  (
    g2611_n,
    g2610_p,
    g2600_p
  );


  and

  (
    g2612_p,
    G4956_o2_p,
    G4017_o2_n
  );


  or

  (
    g2612_n,
    G4956_o2_n,
    G4017_o2_p
  );


  and

  (
    g2613_p,
    G4247_o2_p,
    G4933_o2_n
  );


  or

  (
    g2613_n,
    G4247_o2_n,
    G4933_o2_p
  );


  and

  (
    g2614_p,
    g2613_n,
    g2612_n
  );


  or

  (
    g2614_n,
    g2613_p,
    g2612_p
  );


  and

  (
    g2615_p,
    g2614_p_spl_,
    G2492_o2_p_spl_000
  );


  or

  (
    g2615_n,
    g2614_n_spl_,
    G2492_o2_n_spl_0
  );


  and

  (
    g2616_p,
    g2614_n_spl_,
    G2492_o2_n_spl_0
  );


  or

  (
    g2616_n,
    g2614_p_spl_,
    G2492_o2_p_spl_000
  );


  and

  (
    g2617_p,
    g2616_n,
    g2615_n
  );


  or

  (
    g2617_n,
    g2616_p,
    g2615_p
  );


  and

  (
    g2618_p,
    g2617_p,
    n2341_inv_p_spl_0
  );


  and

  (
    g2619_p,
    g2617_n,
    n2341_inv_n_spl_
  );


  or

  (
    g2620_n,
    g2619_p,
    g2618_p
  );


  and

  (
    g2621_p,
    g2620_n_spl_,
    g2500_p_spl_
  );


  and

  (
    g2622_p,
    g2621_p,
    n4548_lo_n_spl_0
  );


  and

  (
    g2623_p,
    G4954_o2_p,
    G4011_o2_n
  );


  or

  (
    g2623_n,
    G4954_o2_n,
    G4011_o2_p
  );


  and

  (
    g2624_p,
    G4245_o2_p,
    G4930_o2_n
  );


  or

  (
    g2624_n,
    G4245_o2_n,
    G4930_o2_p
  );


  and

  (
    g2625_p,
    g2624_n,
    g2623_n
  );


  or

  (
    g2625_n,
    g2624_p,
    g2623_p
  );


  and

  (
    g2626_p,
    g2625_p_spl_,
    G2492_o2_p_spl_001
  );


  or

  (
    g2626_n,
    g2625_n_spl_,
    G2492_o2_n_spl_1
  );


  and

  (
    g2627_p,
    g2625_n_spl_,
    G2492_o2_n_spl_1
  );


  or

  (
    g2627_n,
    g2625_p_spl_,
    G2492_o2_p_spl_001
  );


  and

  (
    g2628_p,
    g2627_n,
    g2626_n
  );


  or

  (
    g2628_n,
    g2627_p,
    g2626_p
  );


  and

  (
    g2629_p,
    g2628_p,
    n2341_inv_p_spl_0
  );


  and

  (
    g2630_p,
    g2628_n,
    n2341_inv_n_spl_
  );


  or

  (
    g2631_n,
    g2630_p,
    g2629_p
  );


  and

  (
    g2632_p,
    g2631_n_spl_,
    g2500_n_spl_0
  );


  and

  (
    g2633_p,
    g2632_p,
    n4548_lo_n_spl_0
  );


  and

  (
    g2634_p,
    g2500_p_spl_,
    g2470_n
  );


  or

  (
    g2634_n,
    g2500_n_spl_0,
    g2470_p_spl_
  );


  and

  (
    g2635_p,
    g2634_p,
    g2620_n_spl_
  );


  and

  (
    g2636_p,
    g2635_p,
    n4548_lo_p_spl_0
  );


  and

  (
    g2637_p,
    g2634_n,
    g2631_n_spl_
  );


  and

  (
    g2638_p,
    g2637_p,
    n4548_lo_p_spl_0
  );


  or

  (
    g2639_n,
    g2633_p,
    g2622_p
  );


  or

  (
    g2640_n,
    g2639_n,
    g2636_p
  );


  or

  (
    g2641_n,
    g2640_n,
    g2638_p
  );


  and

  (
    g2642_p,
    G5039_o2_p,
    G5036_o2_n
  );


  or

  (
    g2642_n,
    G5039_o2_n,
    G5036_o2_p
  );


  and

  (
    g2643_p,
    g2642_p_spl_,
    n6956_o2_n_spl_01
  );


  or

  (
    g2643_n,
    g2642_n_spl_,
    n6956_o2_p_spl_01
  );


  and

  (
    g2644_p,
    g2642_n_spl_,
    n6956_o2_p_spl_10
  );


  or

  (
    g2644_n,
    g2642_p_spl_,
    n6956_o2_n_spl_10
  );


  and

  (
    g2645_p,
    g2644_n,
    g2643_n
  );


  or

  (
    g2645_n,
    g2644_p,
    g2643_p
  );


  or

  (
    g2646_n,
    g2645_n,
    n7386_o2_p_spl_1
  );


  or

  (
    g2647_n,
    g2645_p,
    n7386_o2_n_spl_1
  );


  and

  (
    g2648_p,
    g2647_n,
    g2646_n
  );


  and

  (
    g2649_p,
    g2648_p,
    n4548_lo_n_spl_
  );


  and

  (
    g2650_p,
    G5006_o2_p,
    G4023_o2_n
  );


  or

  (
    g2650_n,
    G5006_o2_n,
    G4023_o2_p
  );


  and

  (
    g2651_p,
    G4249_o2_p,
    G4984_o2_n
  );


  or

  (
    g2651_n,
    G4249_o2_n,
    G4984_o2_p
  );


  and

  (
    g2652_p,
    g2651_n,
    g2650_n
  );


  or

  (
    g2652_n,
    g2651_p,
    g2650_p
  );


  and

  (
    g2653_p,
    g2652_p_spl_,
    n6956_o2_n_spl_10
  );


  or

  (
    g2653_n,
    g2652_n_spl_,
    n6956_o2_p_spl_10
  );


  and

  (
    g2654_p,
    g2652_n_spl_,
    n6956_o2_p_spl_1
  );


  or

  (
    g2654_n,
    g2652_p_spl_,
    n6956_o2_n_spl_1
  );


  and

  (
    g2655_p,
    g2654_n,
    g2653_n
  );


  or

  (
    g2655_n,
    g2654_p,
    g2653_p
  );


  and

  (
    g2656_p,
    g2655_p,
    n7386_o2_n_spl_1
  );


  and

  (
    g2657_p,
    g2655_n,
    n7386_o2_p_spl_1
  );


  or

  (
    g2658_n,
    g2657_p,
    g2656_p
  );


  and

  (
    g2659_p,
    g2658_n,
    n4548_lo_p_spl_
  );


  or

  (
    g2660_n,
    g2659_p,
    g2649_p
  );


  and

  (
    g2661_p,
    n7136_o2_p_spl_0,
    n7132_o2_n_spl_0
  );


  and

  (
    g2662_p,
    n7136_o2_n_spl_,
    n7132_o2_p_spl_00
  );


  or

  (
    g2663_n,
    g2662_p,
    g2661_p
  );


  and

  (
    g2664_p,
    G2430_o2_p_spl_0,
    n4308_lo_buf_o2_n_spl_1
  );


  and

  (
    g2665_p,
    G2430_o2_n_spl_,
    n4308_lo_buf_o2_p_spl_1
  );


  or

  (
    g2666_n,
    g2665_p,
    g2664_p
  );


  and

  (
    g2667_p,
    n7135_o2_p_spl_0,
    n7133_o2_n_spl_00
  );


  and

  (
    g2668_p,
    n7135_o2_n_spl_,
    n7133_o2_p_spl_00
  );


  or

  (
    g2669_n,
    g2668_p,
    g2667_p
  );


  and

  (
    g2670_p,
    G1734_o2_p_spl_,
    n3657_lo_p_spl_00
  );


  and

  (
    g2671_p,
    G963_o2_n_spl_,
    n3669_lo_p
  );


  or

  (
    g2672_n,
    g2671_p,
    g2670_p
  );


  and

  (
    g2673_p,
    g2514_p,
    n4293_lo_p_spl_0
  );


  and

  (
    g2674_p,
    g2514_n_spl_,
    n4293_lo_n
  );


  or

  (
    g2675_n,
    g2674_p,
    g2673_p
  );


  and

  (
    g2676_p,
    g2511_p,
    n4365_lo_p_spl_0
  );


  and

  (
    g2677_p,
    g2511_n_spl_,
    n4365_lo_n
  );


  or

  (
    g2678_n,
    g2677_p,
    g2676_p
  );


  and

  (
    g2679_p,
    n4080_lo_buf_o2_p_spl_01,
    n4026_lo_p_spl_
  );


  or

  (
    g2679_n,
    n4080_lo_buf_o2_n_spl_0,
    n4026_lo_n
  );


  and

  (
    g2680_p,
    n4080_lo_buf_o2_n_spl_1,
    n4038_lo_p
  );


  or

  (
    g2680_n,
    n4080_lo_buf_o2_p_spl_01,
    n4038_lo_n
  );


  and

  (
    g2681_p,
    g2680_n,
    g2679_n
  );


  or

  (
    g2681_n,
    g2680_p,
    g2679_p
  );


  and

  (
    g2682_p,
    n4092_lo_buf_o2_p_spl_01,
    n3726_lo_p_spl_
  );


  or

  (
    g2682_n,
    n4092_lo_buf_o2_n_spl_0,
    n3726_lo_n
  );


  and

  (
    g2683_p,
    n4092_lo_buf_o2_n_spl_1,
    n3738_lo_p
  );


  or

  (
    g2683_n,
    n4092_lo_buf_o2_p_spl_01,
    n3738_lo_n
  );


  and

  (
    g2684_p,
    g2683_n,
    g2682_n
  );


  or

  (
    g2684_n,
    g2683_p,
    g2682_p
  );


  and

  (
    g2685_p,
    n6775_o2_p_spl_0,
    n6774_o2_p_spl_00
  );


  and

  (
    g2686_p,
    n7019_o2_p_spl_0,
    n7015_o2_p_spl_0
  );


  and

  (
    g2687_p,
    n6688_o2_p_spl_0,
    n6682_o2_p_spl_00
  );


  and

  (
    g2688_p,
    n6689_o2_p_spl_0,
    n6683_o2_p_spl_00
  );


  or

  (
    g2689_n,
    n7136_o2_p_spl_1,
    n7132_o2_p_spl_01
  );


  or

  (
    g2690_n,
    n7135_o2_p_spl_0,
    n7133_o2_p_spl_00
  );


  and

  (
    g2691_p,
    n7005_o2_p_spl_0,
    n7018_o2_p_spl_00
  );


  and

  (
    g2692_p,
    n6686_o2_p_spl_0,
    n6684_o2_p_spl_00
  );


  and

  (
    g2693_p,
    n6687_o2_p_spl_0,
    n6685_o2_p_spl_00
  );


  and

  (
    g2694_p,
    n6623_o2_p_spl_,
    n6621_o2_n
  );


  and

  (
    g2695_p,
    n6623_o2_n,
    n6621_o2_p_spl_
  );


  and

  (
    g2696_p,
    n6669_o2_n_spl_00,
    n3936_lo_p_spl_
  );


  and

  (
    g2697_p,
    n6669_o2_p_spl_00,
    n3936_lo_n_spl_
  );


  and

  (
    g2698_p,
    n6627_o2_p_spl_,
    n6625_o2_n
  );


  and

  (
    g2699_p,
    n6627_o2_n,
    n6625_o2_p_spl_
  );


  and

  (
    g2700_p,
    n6772_o2_n_spl_,
    n4188_lo_p_spl_
  );


  and

  (
    g2701_p,
    n6772_o2_p_spl_1,
    n4188_lo_n
  );


  and

  (
    g2702_p,
    g2529_n_spl_0,
    g2518_p_spl_
  );


  and

  (
    g2703_p,
    g2702_p_spl_0,
    g2526_n_spl_00
  );


  and

  (
    g2704_p,
    g2526_n_spl_00,
    g2519_p_spl_0
  );


  or

  (
    g2705_n,
    g2702_p_spl_0,
    g2519_p_spl_0
  );


  or

  (
    g2706_n,
    g2520_n_spl_0,
    G2486_o2_p_spl_00
  );


  or

  (
    g2707_n,
    g2532_p,
    g2521_n_spl_
  );


  and

  (
    g2708_p,
    g2707_n_spl_0,
    g2520_n_spl_0
  );


  or

  (
    g2709_n,
    g2707_n_spl_0,
    G2486_o2_p_spl_00
  );


  and

  (
    g2710_p,
    n6687_o2_p_spl_0,
    n6686_o2_n_spl_
  );


  and

  (
    g2711_p,
    n6687_o2_n_spl_,
    n6686_o2_p_spl_0
  );


  and

  (
    g2712_p,
    n6629_o2_p,
    n4188_lo_p_spl_
  );


  and

  (
    g2713_p,
    n6549_o2_n,
    n4200_lo_p
  );


  or

  (
    g2714_n,
    g2713_p,
    g2712_p
  );


  or

  (
    g2715_n,
    g2714_n_spl_,
    n6833_o2_p_spl_0
  );


  and

  (
    g2716_p,
    n7384_o2_p_spl_,
    n7023_o2_n_spl_
  );


  and

  (
    g2717_p,
    G2404_o2_p_spl_0,
    n7136_o2_n_spl_
  );


  and

  (
    g2718_p,
    n7384_o2_n_spl_,
    n7023_o2_p_spl_
  );


  and

  (
    g2719_p,
    g2669_n_spl_,
    g2532_n_spl_0
  );


  and

  (
    g2720_p,
    g2719_p_spl_,
    G2486_o2_n
  );


  and

  (
    g2721_p,
    G2404_o2_n_spl_0,
    n7136_o2_p_spl_1
  );


  and

  (
    g2722_p,
    g2714_n_spl_,
    n6833_o2_p_spl_0
  );


  and

  (
    g2723_p,
    g2663_n_spl_,
    g2529_n_spl_0
  );


  and

  (
    g2724_p,
    g2723_p_spl_,
    g2526_n_spl_0
  );


  or

  (
    g2725_n,
    g2704_p_spl_,
    g2562_p_spl_
  );


  or

  (
    g2726_n,
    g2725_n,
    g2703_p_spl_
  );


  and

  (
    g2727_p,
    g2706_n_spl_,
    G2486_o2_p_spl_01
  );


  and

  (
    g2728_p,
    g2727_p,
    g2709_n_spl_
  );


  and

  (
    g2729_p,
    n3756_lo_buf_o2_p_spl_,
    n6947_o2_n
  );


  and

  (
    g2730_p,
    n3756_lo_buf_o2_n,
    n6947_o2_p_spl_
  );


  or

  (
    g2731_n,
    g2730_p,
    g2729_p
  );


  and

  (
    g2732_p,
    n6775_o2_p_spl_0,
    n6774_o2_n_spl_0
  );


  and

  (
    g2733_p,
    n6775_o2_n,
    n6774_o2_p_spl_00
  );


  or

  (
    g2734_n,
    g2733_p,
    g2732_p
  );


  and

  (
    g2735_p,
    n7019_o2_p_spl_0,
    n7015_o2_n_spl_
  );


  and

  (
    g2736_p,
    n7019_o2_n,
    n7015_o2_p_spl_0
  );


  or

  (
    g2737_n,
    g2736_p,
    g2735_p
  );


  and

  (
    g2738_p,
    n6688_o2_p_spl_0,
    n6682_o2_n_spl_0
  );


  and

  (
    g2739_p,
    n6688_o2_n,
    n6682_o2_p_spl_00
  );


  or

  (
    g2740_n,
    g2739_p,
    g2738_p
  );


  and

  (
    g2741_p,
    n6689_o2_p_spl_0,
    n6683_o2_n_spl_0
  );


  and

  (
    g2742_p,
    n6689_o2_n,
    n6683_o2_p_spl_00
  );


  or

  (
    g2743_n,
    g2742_p,
    g2741_p
  );


  and

  (
    g2744_p,
    G2404_o2_p_spl_1,
    n4296_lo_buf_o2_n_spl_0
  );


  and

  (
    g2745_p,
    G2404_o2_n_spl_,
    n4296_lo_buf_o2_p_spl_0
  );


  or

  (
    g2746_n,
    g2745_p,
    g2744_p
  );


  and

  (
    g2747_p,
    G2466_o2_p_spl_0,
    n4368_lo_buf_o2_n_spl_0
  );


  and

  (
    g2748_p,
    G2466_o2_n_spl_0,
    n4368_lo_buf_o2_p_spl_0
  );


  or

  (
    g2749_n,
    g2748_p,
    g2747_p
  );


  and

  (
    g2750_p,
    n7005_o2_p_spl_0,
    n7018_o2_n_spl_0
  );


  and

  (
    g2751_p,
    n7005_o2_n_spl_,
    n7018_o2_p_spl_00
  );


  or

  (
    g2752_n,
    g2751_p,
    g2750_p
  );


  and

  (
    g2753_p,
    n6686_o2_p_spl_,
    n6684_o2_n_spl_0
  );


  and

  (
    g2754_p,
    n6686_o2_n_spl_,
    n6684_o2_p_spl_00
  );


  or

  (
    g2755_n,
    g2754_p,
    g2753_p
  );


  and

  (
    g2756_p,
    n6687_o2_p_spl_,
    n6685_o2_n_spl_0
  );


  and

  (
    g2757_p,
    n6687_o2_n_spl_,
    n6685_o2_p_spl_00
  );


  or

  (
    g2758_n,
    g2757_p,
    g2756_p
  );


  and

  (
    g2759_p,
    G2466_o2_p_spl_1,
    n7005_o2_n_spl_
  );


  and

  (
    g2760_p,
    G2466_o2_n_spl_,
    n7005_o2_p_spl_
  );


  or

  (
    g2761_n,
    g2760_p,
    g2759_p
  );


  and

  (
    g2762_p,
    n6630_o2_p,
    n3936_lo_p_spl_
  );


  or

  (
    g2762_n,
    n6630_o2_n,
    n3936_lo_n_spl_
  );


  and

  (
    g2763_p,
    n6550_o2_n,
    n3948_lo_p
  );


  or

  (
    g2763_n,
    n6550_o2_p,
    n3948_lo_n
  );


  and

  (
    g2764_p,
    g2763_n,
    g2762_n
  );


  or

  (
    g2764_n,
    g2763_p,
    g2762_p
  );


  or

  (
    g2765_n,
    g2764_n,
    G2430_o2_p_spl_0
  );


  or

  (
    g2766_n,
    g2764_p,
    G2430_o2_n_spl_
  );


  and

  (
    g2767_p,
    g2766_n,
    g2765_n
  );


  and

  (
    g2768_p,
    n2965_inv_n_spl_00,
    n7132_o2_p_spl_01
  );


  or

  (
    g2768_n,
    n2965_inv_p_spl_00,
    n7132_o2_n_spl_0
  );


  and

  (
    g2769_p,
    g2768_p,
    G1138_o2_n_spl_
  );


  or

  (
    g2769_n,
    g2768_n,
    G1138_o2_p_spl_
  );


  and

  (
    g2770_p,
    n2971_inv_n_spl_00,
    n7132_o2_p_spl_10
  );


  or

  (
    g2770_n,
    n2971_inv_p_spl_00,
    n7132_o2_n_spl_1
  );


  and

  (
    g2771_p,
    g2770_p,
    G1138_o2_p_spl_
  );


  or

  (
    g2771_n,
    g2770_n,
    G1138_o2_n_spl_
  );


  and

  (
    g2772_p,
    g2771_n,
    g2769_n
  );


  or

  (
    g2772_n,
    g2771_p,
    g2769_p
  );


  and

  (
    g2773_p,
    n3118_inv_n_spl_00,
    n6982_o2_n_spl_
  );


  or

  (
    g2773_n,
    n3118_inv_p_spl_000,
    n6982_o2_p_spl_00
  );


  and

  (
    g2774_p,
    n3127_inv_n_spl_00,
    n6982_o2_p_spl_00
  );


  or

  (
    g2774_n,
    n3127_inv_p_spl_000,
    n6982_o2_n_spl_
  );


  and

  (
    g2775_p,
    g2774_n,
    g2773_n
  );


  or

  (
    g2775_n,
    g2774_p,
    g2773_p
  );


  and

  (
    g2776_p,
    g2775_p,
    n7132_o2_n_spl_1
  );


  or

  (
    g2776_n,
    g2775_n,
    n7132_o2_p_spl_10
  );


  and

  (
    g2777_p,
    g2776_n,
    g2772_p
  );


  or

  (
    g2777_n,
    g2776_p,
    g2772_n
  );


  and

  (
    g2778_p,
    n2965_inv_n_spl_00,
    n7016_o2_p_spl_01
  );


  or

  (
    g2778_n,
    n2965_inv_p_spl_00,
    n7016_o2_n_spl_0
  );


  and

  (
    g2779_p,
    g2778_p,
    G1132_o2_n_spl_
  );


  or

  (
    g2779_n,
    g2778_n,
    G1132_o2_p_spl_
  );


  and

  (
    g2780_p,
    n2971_inv_n_spl_00,
    n7016_o2_p_spl_01
  );


  or

  (
    g2780_n,
    n2971_inv_p_spl_00,
    n7016_o2_n_spl_1
  );


  and

  (
    g2781_p,
    g2780_p,
    G1132_o2_p_spl_
  );


  or

  (
    g2781_n,
    g2780_n,
    G1132_o2_n_spl_
  );


  and

  (
    g2782_p,
    g2781_n,
    g2779_n
  );


  or

  (
    g2782_n,
    g2781_p,
    g2779_p
  );


  and

  (
    g2783_p,
    n3118_inv_n_spl_00,
    n6945_o2_n_spl_
  );


  or

  (
    g2783_n,
    n3118_inv_p_spl_000,
    n6945_o2_p_spl_00
  );


  and

  (
    g2784_p,
    n3127_inv_n_spl_00,
    n6945_o2_p_spl_00
  );


  or

  (
    g2784_n,
    n3127_inv_p_spl_000,
    n6945_o2_n_spl_
  );


  and

  (
    g2785_p,
    g2784_n,
    g2783_n
  );


  or

  (
    g2785_n,
    g2784_p,
    g2783_p
  );


  and

  (
    g2786_p,
    g2785_p,
    n7016_o2_n_spl_1
  );


  or

  (
    g2786_n,
    g2785_n,
    n7016_o2_p_spl_1
  );


  and

  (
    g2787_p,
    g2786_n,
    g2782_p
  );


  or

  (
    g2787_n,
    g2786_p,
    g2782_n
  );


  and

  (
    g2788_p,
    g2787_n_spl_,
    g2777_p_spl_
  );


  or

  (
    g2788_n,
    g2787_p_spl_,
    g2777_n_spl_
  );


  and

  (
    g2789_p,
    g2787_p_spl_,
    g2777_n_spl_
  );


  or

  (
    g2789_n,
    g2787_n_spl_,
    g2777_p_spl_
  );


  and

  (
    g2790_p,
    g2789_n,
    g2788_n
  );


  or

  (
    g2790_n,
    g2789_p,
    g2788_p
  );


  and

  (
    g2791_p,
    n2965_inv_n_spl_01,
    n7383_o2_p_spl_01
  );


  or

  (
    g2791_n,
    n2965_inv_p_spl_01,
    n7383_o2_n_spl_0
  );


  and

  (
    g2792_p,
    g2791_p,
    G1126_o2_n_spl_
  );


  or

  (
    g2792_n,
    g2791_n,
    G1126_o2_p_spl_
  );


  and

  (
    g2793_p,
    n2971_inv_n_spl_01,
    n7383_o2_p_spl_01
  );


  or

  (
    g2793_n,
    n2971_inv_p_spl_01,
    n7383_o2_n_spl_1
  );


  and

  (
    g2794_p,
    g2793_p,
    G1126_o2_p_spl_
  );


  or

  (
    g2794_n,
    g2793_n,
    G1126_o2_n_spl_
  );


  and

  (
    g2795_p,
    g2794_n,
    g2792_n
  );


  or

  (
    g2795_n,
    g2794_p,
    g2792_p
  );


  and

  (
    g2796_p,
    n3118_inv_n_spl_01,
    n7175_o2_n_spl_
  );


  or

  (
    g2796_n,
    n3118_inv_p_spl_00,
    n7175_o2_p_spl_00
  );


  and

  (
    g2797_p,
    n3127_inv_n_spl_01,
    n7175_o2_p_spl_00
  );


  or

  (
    g2797_n,
    n3127_inv_p_spl_00,
    n7175_o2_n_spl_
  );


  and

  (
    g2798_p,
    g2797_n,
    g2796_n
  );


  or

  (
    g2798_n,
    g2797_p,
    g2796_p
  );


  and

  (
    g2799_p,
    g2798_p,
    n7383_o2_n_spl_1
  );


  or

  (
    g2799_n,
    g2798_n,
    n7383_o2_p_spl_1
  );


  and

  (
    g2800_p,
    g2799_n,
    g2795_p
  );


  or

  (
    g2800_n,
    g2799_p,
    g2795_n
  );


  and

  (
    g2801_p,
    g2800_p_spl_,
    g2462_p_spl_
  );


  or

  (
    g2801_n,
    g2800_n_spl_,
    g2462_n_spl_0
  );


  and

  (
    g2802_p,
    g2800_n_spl_,
    g2462_n_spl_0
  );


  or

  (
    g2802_n,
    g2800_p_spl_,
    g2462_p_spl_
  );


  and

  (
    g2803_p,
    g2802_n,
    g2801_n
  );


  or

  (
    g2803_n,
    g2802_p,
    g2801_p
  );


  or

  (
    g2804_n,
    g2803_n,
    g2790_p
  );


  or

  (
    g2805_n,
    g2803_p,
    g2790_n
  );


  and

  (
    g2806_p,
    g2805_n,
    g2804_n
  );


  and

  (
    g2807_p,
    n2968_inv_n_spl_01,
    n7133_o2_p_spl_01
  );


  or

  (
    g2807_n,
    n2968_inv_p_spl_00,
    n7133_o2_n_spl_0
  );


  and

  (
    g2808_p,
    g2807_p,
    G1114_o2_n_spl_
  );


  or

  (
    g2808_n,
    g2807_n,
    G1114_o2_p_spl_
  );


  and

  (
    g2809_p,
    n2974_inv_n_spl_01,
    n7133_o2_p_spl_01
  );


  or

  (
    g2809_n,
    n2974_inv_p_spl_01,
    n7133_o2_n_spl_1
  );


  and

  (
    g2810_p,
    g2809_p,
    G1114_o2_p_spl_
  );


  or

  (
    g2810_n,
    g2809_n,
    G1114_o2_n_spl_
  );


  and

  (
    g2811_p,
    g2810_n,
    g2808_n
  );


  or

  (
    g2811_n,
    g2810_p,
    g2808_p
  );


  and

  (
    g2812_p,
    n3121_inv_n_spl_00,
    n6984_o2_n_spl_
  );


  or

  (
    g2812_n,
    n3121_inv_p_spl_000,
    n6984_o2_p_spl_00
  );


  and

  (
    g2813_p,
    n3124_inv_n_spl_00,
    n6984_o2_p_spl_00
  );


  or

  (
    g2813_n,
    n3124_inv_p_spl_00,
    n6984_o2_n_spl_
  );


  and

  (
    g2814_p,
    g2813_n,
    g2812_n
  );


  or

  (
    g2814_n,
    g2813_p,
    g2812_p
  );


  and

  (
    g2815_p,
    g2814_p,
    n7133_o2_n_spl_1
  );


  or

  (
    g2815_n,
    g2814_n,
    n7133_o2_p_spl_1
  );


  and

  (
    g2816_p,
    g2815_n,
    g2811_p
  );


  or

  (
    g2816_n,
    g2815_p,
    g2811_n
  );


  and

  (
    g2817_p,
    n2968_inv_n_spl_01,
    n7017_o2_p_spl_01
  );


  or

  (
    g2817_n,
    n2968_inv_p_spl_01,
    n7017_o2_n_spl_01
  );


  and

  (
    g2818_p,
    g2817_p,
    G1108_o2_n_spl_
  );


  or

  (
    g2818_n,
    g2817_n,
    G1108_o2_p_spl_
  );


  and

  (
    g2819_p,
    n2974_inv_n_spl_01,
    n7017_o2_p_spl_01
  );


  or

  (
    g2819_n,
    n2974_inv_p_spl_01,
    n7017_o2_n_spl_1
  );


  and

  (
    g2820_p,
    g2819_p,
    G1108_o2_p_spl_
  );


  or

  (
    g2820_n,
    g2819_n,
    G1108_o2_n_spl_
  );


  and

  (
    g2821_p,
    g2820_n,
    g2818_n
  );


  or

  (
    g2821_n,
    g2820_p,
    g2818_p
  );


  and

  (
    g2822_p,
    n3121_inv_n_spl_01,
    n6949_o2_n_spl_
  );


  or

  (
    g2822_n,
    n3121_inv_p_spl_00,
    n6949_o2_p_spl_00
  );


  and

  (
    g2823_p,
    n3124_inv_n_spl_01,
    n6949_o2_p_spl_00
  );


  or

  (
    g2823_n,
    n3124_inv_p_spl_01,
    n6949_o2_n_spl_
  );


  and

  (
    g2824_p,
    g2823_n,
    g2822_n
  );


  or

  (
    g2824_n,
    g2823_p,
    g2822_p
  );


  and

  (
    g2825_p,
    g2824_p,
    n7017_o2_n_spl_1
  );


  or

  (
    g2825_n,
    g2824_n,
    n7017_o2_p_spl_1
  );


  and

  (
    g2826_p,
    g2825_n,
    g2821_p
  );


  or

  (
    g2826_n,
    g2825_p,
    g2821_n
  );


  and

  (
    g2827_p,
    g2826_n_spl_,
    g2816_p_spl_
  );


  or

  (
    g2827_n,
    g2826_p_spl_,
    g2816_n_spl_
  );


  and

  (
    g2828_p,
    g2826_p_spl_,
    g2816_n_spl_
  );


  or

  (
    g2828_n,
    g2826_n_spl_,
    g2816_p_spl_
  );


  and

  (
    g2829_p,
    g2828_n,
    g2827_n
  );


  or

  (
    g2829_n,
    g2828_p,
    g2827_p
  );


  and

  (
    g2830_p,
    n2968_inv_n_spl_10,
    n7453_o2_n_spl_
  );


  or

  (
    g2830_n,
    n2968_inv_p_spl_01,
    n7453_o2_p_spl_00
  );


  and

  (
    g2831_p,
    n2974_inv_n_spl_10,
    n7453_o2_p_spl_00
  );


  or

  (
    g2831_n,
    n2974_inv_p_spl_10,
    n7453_o2_n_spl_
  );


  and

  (
    g2832_p,
    g2831_n,
    g2830_n
  );


  or

  (
    g2832_n,
    g2831_p,
    g2830_p
  );


  and

  (
    g2833_p,
    n3121_inv_n_spl_01,
    n3960_lo_buf_o2_n_spl_
  );


  or

  (
    g2833_n,
    n3121_inv_p_spl_01,
    n3960_lo_buf_o2_p_spl_00
  );


  and

  (
    g2834_p,
    n3124_inv_n_spl_01,
    n3960_lo_buf_o2_p_spl_00
  );


  or

  (
    g2834_n,
    n3124_inv_p_spl_01,
    n3960_lo_buf_o2_n_spl_
  );


  and

  (
    g2835_p,
    g2834_n,
    g2833_n
  );


  or

  (
    g2835_n,
    g2834_p,
    g2833_p
  );


  and

  (
    g2836_p,
    g2835_p_spl_,
    g2832_p_spl_
  );


  or

  (
    g2836_n,
    g2835_n_spl_,
    g2832_n_spl_
  );


  and

  (
    g2837_p,
    g2835_n_spl_,
    g2832_n_spl_
  );


  or

  (
    g2837_n,
    g2835_p_spl_,
    g2832_p_spl_
  );


  and

  (
    g2838_p,
    g2837_n,
    g2836_n
  );


  or

  (
    g2838_n,
    g2837_p,
    g2836_p
  );


  or

  (
    g2839_n,
    g2838_n,
    g2829_p
  );


  or

  (
    g2840_n,
    g2838_p,
    g2829_n
  );


  and

  (
    g2841_p,
    g2840_n,
    g2839_n
  );


  and

  (
    g2842_p,
    n2965_inv_n_spl_01,
    n6774_o2_p_spl_01
  );


  or

  (
    g2842_n,
    n2965_inv_p_spl_01,
    n6774_o2_n_spl_0
  );


  and

  (
    g2843_p,
    g2842_p,
    n6669_o2_n_spl_00
  );


  or

  (
    g2843_n,
    g2842_n,
    n6669_o2_p_spl_00
  );


  and

  (
    g2844_p,
    n2971_inv_n_spl_01,
    n6774_o2_p_spl_01
  );


  or

  (
    g2844_n,
    n2971_inv_p_spl_01,
    n6774_o2_n_spl_1
  );


  and

  (
    g2845_p,
    g2844_p,
    n6669_o2_p_spl_01
  );


  or

  (
    g2845_n,
    g2844_n,
    n6669_o2_n_spl_0
  );


  and

  (
    g2846_p,
    g2845_n,
    g2843_n
  );


  or

  (
    g2846_n,
    g2845_p,
    g2843_p
  );


  and

  (
    g2847_p,
    n3118_inv_n_spl_01,
    n6669_o2_n_spl_1
  );


  or

  (
    g2847_n,
    n3118_inv_p_spl_01,
    n6669_o2_p_spl_01
  );


  and

  (
    g2848_p,
    n3127_inv_n_spl_01,
    n6669_o2_p_spl_1
  );


  or

  (
    g2848_n,
    n3127_inv_p_spl_01,
    n6669_o2_n_spl_1
  );


  and

  (
    g2849_p,
    g2848_n,
    g2847_n
  );


  or

  (
    g2849_n,
    g2848_p,
    g2847_p
  );


  and

  (
    g2850_p,
    g2849_p,
    n6774_o2_n_spl_1
  );


  or

  (
    g2850_n,
    g2849_n,
    n6774_o2_p_spl_1
  );


  and

  (
    g2851_p,
    g2850_n,
    g2846_p
  );


  or

  (
    g2851_n,
    g2850_p,
    g2846_n
  );


  and

  (
    g2852_p,
    n2965_inv_n_spl_1,
    n6683_o2_p_spl_01
  );


  or

  (
    g2852_n,
    n2965_inv_p_spl_10,
    n6683_o2_n_spl_0
  );


  and

  (
    g2853_p,
    g2852_p,
    G1044_o2_n
  );


  or

  (
    g2853_n,
    g2852_n,
    G1044_o2_p
  );


  and

  (
    g2854_p,
    n2971_inv_n_spl_1,
    n6683_o2_p_spl_01
  );


  or

  (
    g2854_n,
    n2971_inv_p_spl_10,
    n6683_o2_n_spl_1
  );


  and

  (
    g2855_p,
    g2854_p,
    G1804_o2_p
  );


  or

  (
    g2855_n,
    g2854_n,
    G1804_o2_n
  );


  and

  (
    g2856_p,
    g2855_n,
    g2853_n
  );


  or

  (
    g2856_n,
    g2855_p,
    g2853_p
  );


  and

  (
    g2857_p,
    n3118_inv_n_spl_10,
    G1041_o2_n_spl_
  );


  or

  (
    g2857_n,
    n3118_inv_p_spl_01,
    G1041_o2_p_spl_
  );


  and

  (
    g2858_p,
    n3127_inv_n_spl_10,
    G1041_o2_p_spl_
  );


  or

  (
    g2858_n,
    n3127_inv_p_spl_01,
    G1041_o2_n_spl_
  );


  and

  (
    g2859_p,
    g2858_n,
    g2857_n
  );


  or

  (
    g2859_n,
    g2858_p,
    g2857_p
  );


  and

  (
    g2860_p,
    g2859_p,
    n6683_o2_n_spl_1
  );


  or

  (
    g2860_n,
    g2859_n,
    n6683_o2_p_spl_1
  );


  and

  (
    g2861_p,
    g2860_n,
    g2856_p
  );


  or

  (
    g2861_n,
    g2860_p,
    g2856_n
  );


  and

  (
    g2862_p,
    n2965_inv_n_spl_1,
    n6682_o2_p_spl_01
  );


  or

  (
    g2862_n,
    n2965_inv_p_spl_10,
    n6682_o2_n_spl_0
  );


  and

  (
    g2863_p,
    g2862_p,
    G1038_o2_n
  );


  or

  (
    g2863_n,
    g2862_n,
    G1038_o2_p
  );


  and

  (
    g2864_p,
    n2971_inv_n_spl_1,
    n6682_o2_p_spl_01
  );


  or

  (
    g2864_n,
    n2971_inv_p_spl_10,
    n6682_o2_n_spl_1
  );


  and

  (
    g2865_p,
    g2864_p,
    G1802_o2_p
  );


  or

  (
    g2865_n,
    g2864_n,
    G1802_o2_n
  );


  and

  (
    g2866_p,
    g2865_n,
    g2863_n
  );


  or

  (
    g2866_n,
    g2865_p,
    g2863_p
  );


  and

  (
    g2867_p,
    n3118_inv_n_spl_10,
    G1035_o2_n_spl_
  );


  or

  (
    g2867_n,
    n3118_inv_p_spl_10,
    G1035_o2_p_spl_
  );


  and

  (
    g2868_p,
    n3127_inv_n_spl_10,
    G1035_o2_p_spl_
  );


  or

  (
    g2868_n,
    n3127_inv_p_spl_10,
    G1035_o2_n_spl_
  );


  and

  (
    g2869_p,
    g2868_n,
    g2867_n
  );


  or

  (
    g2869_n,
    g2868_p,
    g2867_p
  );


  and

  (
    g2870_p,
    g2869_p,
    n6682_o2_n_spl_1
  );


  or

  (
    g2870_n,
    g2869_n,
    n6682_o2_p_spl_1
  );


  and

  (
    g2871_p,
    g2870_n,
    g2866_p
  );


  or

  (
    g2871_n,
    g2870_p,
    g2866_n
  );


  and

  (
    g2872_p,
    g2871_n_spl_,
    g2861_p_spl_
  );


  or

  (
    g2872_n,
    g2871_p_spl_,
    g2861_n_spl_
  );


  and

  (
    g2873_p,
    g2871_p_spl_,
    g2861_n_spl_
  );


  or

  (
    g2873_n,
    g2871_n_spl_,
    g2861_p_spl_
  );


  and

  (
    g2874_p,
    g2873_n,
    g2872_n
  );


  or

  (
    g2874_n,
    g2873_p,
    g2872_p
  );


  and

  (
    g2875_p,
    G2108_o2_n,
    G1807_o2_n
  );


  or

  (
    g2875_n,
    G2108_o2_p,
    G1807_o2_p
  );


  and

  (
    g2876_p,
    n3118_inv_n_spl_11,
    G1029_o2_n
  );


  or

  (
    g2876_n,
    n3118_inv_p_spl_10,
    G1029_o2_p
  );


  and

  (
    g2877_p,
    G1799_o2_p,
    n3127_inv_n_spl_11
  );


  or

  (
    g2877_n,
    G1799_o2_n,
    n3127_inv_p_spl_10
  );


  and

  (
    g2878_p,
    g2877_n,
    g2876_n
  );


  or

  (
    g2878_n,
    g2877_p,
    g2876_p
  );


  and

  (
    g2879_p,
    g2878_p,
    n7015_o2_n_spl_
  );


  or

  (
    g2879_n,
    g2878_n,
    n7015_o2_p_spl_1
  );


  and

  (
    g2880_p,
    g2879_n,
    g2875_p
  );


  or

  (
    g2880_n,
    g2879_p,
    g2875_n
  );


  and

  (
    g2881_p,
    G2134_o2_n,
    G1899_o2_n
  );


  or

  (
    g2881_n,
    G2134_o2_p,
    G1899_o2_p
  );


  and

  (
    g2882_p,
    n3118_inv_n_spl_11,
    G1141_o2_n
  );


  or

  (
    g2882_n,
    n3118_inv_p_spl_11,
    G1141_o2_p
  );


  and

  (
    g2883_p,
    G1894_o2_p,
    n3127_inv_n_spl_11
  );


  or

  (
    g2883_n,
    G1894_o2_n,
    n3127_inv_p_spl_11
  );


  and

  (
    g2884_p,
    g2883_n,
    g2882_n
  );


  or

  (
    g2884_n,
    g2883_p,
    g2882_p
  );


  and

  (
    g2885_p,
    g2884_p,
    n4296_lo_buf_o2_n_spl_
  );


  or

  (
    g2885_n,
    g2884_n,
    n4296_lo_buf_o2_p_spl_1
  );


  and

  (
    g2886_p,
    g2885_n,
    g2881_p
  );


  or

  (
    g2886_n,
    g2885_p,
    g2881_n
  );


  and

  (
    g2887_p,
    g2886_n_spl_,
    g2880_p_spl_
  );


  or

  (
    g2887_n,
    g2886_p_spl_,
    g2880_n_spl_
  );


  and

  (
    g2888_p,
    g2886_p_spl_,
    g2880_n_spl_
  );


  or

  (
    g2888_n,
    g2886_n_spl_,
    g2880_p_spl_
  );


  and

  (
    g2889_p,
    g2888_n,
    g2887_n
  );


  or

  (
    g2889_n,
    g2888_p,
    g2887_p
  );


  or

  (
    g2890_n,
    g2874_n_spl_,
    g2851_p_spl_
  );


  or

  (
    g2891_n,
    g2890_n,
    g2889_p_spl_
  );


  or

  (
    g2892_n,
    g2874_n_spl_,
    g2851_n_spl_
  );


  or

  (
    g2893_n,
    g2892_n,
    g2889_n_spl_
  );


  and

  (
    g2894_p,
    g2893_n,
    g2891_n
  );


  or

  (
    g2895_n,
    g2874_p_spl_,
    g2851_n_spl_
  );


  or

  (
    g2896_n,
    g2895_n,
    g2889_p_spl_
  );


  or

  (
    g2897_n,
    g2874_p_spl_,
    g2851_p_spl_
  );


  or

  (
    g2898_n,
    g2897_n,
    g2889_n_spl_
  );


  and

  (
    g2899_p,
    g2898_n,
    g2896_n
  );


  and

  (
    g2900_p,
    g2899_p,
    g2894_p
  );


  and

  (
    g2901_p,
    n2968_inv_n_spl_10,
    n6685_o2_p_spl_01
  );


  or

  (
    g2901_n,
    n2968_inv_p_spl_10,
    n6685_o2_n_spl_0
  );


  and

  (
    g2902_p,
    g2901_p,
    G1096_o2_n
  );


  or

  (
    g2902_n,
    g2901_n,
    G1096_o2_p
  );


  and

  (
    g2903_p,
    n2974_inv_n_spl_10,
    n6685_o2_p_spl_01
  );


  or

  (
    g2903_n,
    n2974_inv_p_spl_10,
    n6685_o2_n_spl_1
  );


  and

  (
    g2904_p,
    g2903_p,
    G1851_o2_p
  );


  or

  (
    g2904_n,
    g2903_n,
    G1851_o2_n
  );


  and

  (
    g2905_p,
    g2904_n,
    g2902_n
  );


  or

  (
    g2905_n,
    g2904_p,
    g2902_p
  );


  and

  (
    g2906_p,
    n3121_inv_n_spl_10,
    G1093_o2_n_spl_
  );


  or

  (
    g2906_n,
    n3121_inv_p_spl_01,
    G1093_o2_p_spl_
  );


  and

  (
    g2907_p,
    n3124_inv_n_spl_10,
    G1093_o2_p_spl_
  );


  or

  (
    g2907_n,
    n3124_inv_p_spl_10,
    G1093_o2_n_spl_
  );


  and

  (
    g2908_p,
    g2907_n,
    g2906_n
  );


  or

  (
    g2908_n,
    g2907_p,
    g2906_p
  );


  and

  (
    g2909_p,
    g2908_p,
    n6685_o2_n_spl_1
  );


  or

  (
    g2909_n,
    g2908_n,
    n6685_o2_p_spl_1
  );


  and

  (
    g2910_p,
    g2909_n,
    g2905_p
  );


  or

  (
    g2910_n,
    g2909_p,
    g2905_n
  );


  and

  (
    g2911_p,
    n2968_inv_n_spl_11,
    n6684_o2_p_spl_01
  );


  or

  (
    g2911_n,
    n2968_inv_p_spl_10,
    n6684_o2_n_spl_0
  );


  and

  (
    g2912_p,
    g2911_p,
    G1090_o2_n
  );


  or

  (
    g2912_n,
    g2911_n,
    G1090_o2_p
  );


  and

  (
    g2913_p,
    n2974_inv_n_spl_1,
    n6684_o2_p_spl_01
  );


  or

  (
    g2913_n,
    n2974_inv_p_spl_11,
    n6684_o2_n_spl_1
  );


  and

  (
    g2914_p,
    g2913_p,
    G1849_o2_p
  );


  or

  (
    g2914_n,
    g2913_n,
    G1849_o2_n
  );


  and

  (
    g2915_p,
    g2914_n,
    g2912_n
  );


  or

  (
    g2915_n,
    g2914_p,
    g2912_p
  );


  and

  (
    g2916_p,
    n3121_inv_n_spl_10,
    G1087_o2_n_spl_
  );


  or

  (
    g2916_n,
    n3121_inv_p_spl_10,
    G1087_o2_p_spl_
  );


  and

  (
    g2917_p,
    n3124_inv_n_spl_10,
    G1087_o2_p_spl_
  );


  or

  (
    g2917_n,
    n3124_inv_p_spl_10,
    G1087_o2_n_spl_
  );


  and

  (
    g2918_p,
    g2917_n,
    g2916_n
  );


  or

  (
    g2918_n,
    g2917_p,
    g2916_p
  );


  and

  (
    g2919_p,
    g2918_p,
    n6684_o2_n_spl_1
  );


  or

  (
    g2919_n,
    g2918_n,
    n6684_o2_p_spl_1
  );


  and

  (
    g2920_p,
    g2919_n,
    g2915_p
  );


  or

  (
    g2920_n,
    g2919_p,
    g2915_n
  );


  and

  (
    g2921_p,
    g2920_n_spl_,
    g2910_p_spl_
  );


  or

  (
    g2921_n,
    g2920_p_spl_,
    g2910_n_spl_
  );


  and

  (
    g2922_p,
    g2920_p_spl_,
    g2910_n_spl_
  );


  or

  (
    g2922_n,
    g2920_n_spl_,
    g2910_p_spl_
  );


  and

  (
    g2923_p,
    g2922_n,
    g2921_n
  );


  or

  (
    g2923_n,
    g2922_p,
    g2921_p
  );


  and

  (
    g2924_p,
    n2968_inv_n_spl_11,
    n7018_o2_p_spl_0
  );


  or

  (
    g2924_n,
    n2968_inv_p_spl_11,
    n7018_o2_n_spl_0
  );


  and

  (
    g2925_p,
    n3121_inv_p_spl_10,
    n7018_o2_n_spl_
  );


  or

  (
    g2925_n,
    n3121_inv_n_spl_11,
    n7018_o2_p_spl_1
  );


  and

  (
    g2926_p,
    g2925_n,
    g2924_n
  );


  or

  (
    g2926_n,
    g2925_p,
    g2924_p
  );


  and

  (
    g2927_p,
    G2116_o2_n,
    G1852_o2_n
  );


  or

  (
    g2927_n,
    G2116_o2_p,
    G1852_o2_p
  );


  and

  (
    g2928_p,
    n3121_inv_n_spl_11,
    G1081_o2_n
  );


  or

  (
    g2928_n,
    n3121_inv_p_spl_11,
    G1081_o2_p
  );


  and

  (
    g2929_p,
    G1846_o2_p,
    n3124_inv_n_spl_1
  );


  or

  (
    g2929_n,
    G1846_o2_n,
    n3124_inv_p_spl_11
  );


  and

  (
    g2930_p,
    g2929_n,
    g2928_n
  );


  or

  (
    g2930_n,
    g2929_p,
    g2928_p
  );


  and

  (
    g2931_p,
    g2930_p,
    n4368_lo_buf_o2_n_spl_
  );


  or

  (
    g2931_n,
    g2930_n,
    n4368_lo_buf_o2_p_spl_1
  );


  and

  (
    g2932_p,
    g2931_n,
    g2927_p
  );


  or

  (
    g2932_n,
    g2931_p,
    g2927_n
  );


  and

  (
    g2933_p,
    g2932_n_spl_,
    g2926_p_spl_
  );


  or

  (
    g2933_n,
    g2932_p_spl_,
    g2926_n_spl_
  );


  and

  (
    g2934_p,
    g2932_p_spl_,
    g2926_n_spl_
  );


  or

  (
    g2934_n,
    g2932_n_spl_,
    g2926_p_spl_
  );


  and

  (
    g2935_p,
    g2934_n,
    g2933_n
  );


  or

  (
    g2935_n,
    g2934_p,
    g2933_p
  );


  and

  (
    g2936_p,
    g2923_p_spl_,
    g2503_n_spl_
  );


  and

  (
    g2937_p,
    g2936_p,
    g2935_n_spl_
  );


  and

  (
    g2938_p,
    g2923_p_spl_,
    g2503_p_spl_0
  );


  and

  (
    g2939_p,
    g2938_p,
    g2935_p_spl_
  );


  or

  (
    g2940_n,
    g2939_p,
    g2937_p
  );


  and

  (
    g2941_p,
    g2923_n_spl_,
    g2503_p_spl_0
  );


  and

  (
    g2942_p,
    g2941_p,
    g2935_n_spl_
  );


  and

  (
    g2943_p,
    g2923_n_spl_,
    g2503_n_spl_
  );


  and

  (
    g2944_p,
    g2943_p,
    g2935_p_spl_
  );


  or

  (
    g2945_n,
    g2944_p,
    g2942_p
  );


  or

  (
    g2946_n,
    g2945_n,
    g2940_n
  );


  and

  (
    g2947_p,
    g2684_n_spl_0,
    n4278_lo_p_spl_0
  );


  and

  (
    g2948_p,
    g2681_n_spl_0,
    n4350_lo_p_spl_0
  );


  and

  (
    g2949_p,
    G3809_o2_n,
    G2727_o2_n
  );


  or

  (
    g2949_n,
    G3809_o2_p,
    G2727_o2_p_spl_
  );


  and

  (
    g2950_p,
    g2949_p,
    G3810_o2_n
  );


  or

  (
    g2950_n,
    g2949_n,
    G3810_o2_p
  );


  and

  (
    g2951_p,
    g2950_p,
    G3811_o2_n
  );


  or

  (
    g2951_n,
    g2950_n,
    G3811_o2_p
  );


  and

  (
    g2952_p,
    g2951_p,
    G3812_o2_n
  );


  or

  (
    g2952_n,
    g2951_n,
    G3812_o2_p
  );


  and

  (
    g2953_p,
    G4580_o2_p,
    G4670_o2_n
  );


  or

  (
    g2953_n,
    G4580_o2_n,
    G4670_o2_p
  );


  and

  (
    g2954_p,
    g2953_p_spl_,
    g2952_n_spl_
  );


  or

  (
    g2954_n,
    g2953_n_spl_,
    g2952_p_spl_
  );


  and

  (
    g2955_p,
    g2953_n_spl_,
    g2952_p_spl_
  );


  or

  (
    g2955_n,
    g2953_p_spl_,
    g2952_n_spl_
  );


  and

  (
    g2956_p,
    g2955_n,
    g2954_n
  );


  or

  (
    g2956_n,
    g2955_p,
    g2954_p
  );


  and

  (
    g2957_p,
    g2956_p_spl_,
    G3552_o2_n_spl_0
  );


  or

  (
    g2957_n,
    g2956_n_spl_,
    G3552_o2_p_spl_00
  );


  and

  (
    g2958_p,
    g2956_n_spl_,
    G3552_o2_p_spl_00
  );


  or

  (
    g2958_n,
    g2956_p_spl_,
    G3552_o2_n_spl_0
  );


  and

  (
    g2959_p,
    g2958_n,
    g2957_n
  );


  or

  (
    g2959_n,
    g2958_p,
    g2957_p
  );


  or

  (
    g2960_n,
    g2959_n,
    G3533_o2_p_spl_0
  );


  or

  (
    g2961_n,
    g2959_p,
    G3533_o2_n_spl_
  );


  and

  (
    g2962_p,
    g2961_n,
    g2960_n
  );


  and

  (
    g2963_p,
    G3716_o2_n,
    G2543_o2_n
  );


  or

  (
    g2963_n,
    G3716_o2_p,
    G2543_o2_p_spl_
  );


  and

  (
    g2964_p,
    g2963_p,
    G3866_o2_n
  );


  or

  (
    g2964_n,
    g2963_n,
    G3866_o2_p
  );


  and

  (
    g2965_p,
    g2964_p,
    G3867_o2_n
  );


  or

  (
    g2965_n,
    g2964_n,
    G3867_o2_p
  );


  and

  (
    g2966_p,
    g2965_p,
    G3868_o2_n
  );


  or

  (
    g2966_n,
    g2965_n,
    G3868_o2_p
  );


  and

  (
    g2967_p,
    G4493_o2_n,
    G4529_o2_n
  );


  or

  (
    g2967_n,
    G4493_o2_p,
    G4529_o2_p
  );


  and

  (
    g2968_p,
    g2967_p_spl_,
    g2966_n_spl_
  );


  or

  (
    g2968_n,
    g2967_n_spl_,
    g2966_p_spl_
  );


  and

  (
    g2969_p,
    g2967_n_spl_,
    g2966_p_spl_
  );


  or

  (
    g2969_n,
    g2967_p_spl_,
    g2966_n_spl_
  );


  and

  (
    g2970_p,
    g2969_n,
    g2968_n
  );


  or

  (
    g2970_n,
    g2969_p,
    g2968_p
  );


  and

  (
    g2971_p,
    g2970_p_spl_,
    n2647_inv_p_spl_00
  );


  or

  (
    g2971_n,
    g2970_n_spl_,
    n2647_inv_n_spl_0
  );


  and

  (
    g2972_p,
    g2970_n_spl_,
    n2647_inv_n_spl_0
  );


  or

  (
    g2972_n,
    g2970_p_spl_,
    n2647_inv_p_spl_00
  );


  and

  (
    g2973_p,
    g2972_n,
    g2971_n
  );


  or

  (
    g2973_n,
    g2972_p,
    g2971_p
  );


  or

  (
    g2974_n,
    g2973_n,
    G3645_o2_p_spl_0
  );


  or

  (
    g2975_n,
    g2973_p,
    G3645_o2_n_spl_
  );


  and

  (
    g2976_p,
    g2975_n,
    g2974_n
  );


  and

  (
    g2977_p,
    g2507_n_spl_0,
    G2715_o2_p_spl_
  );


  or

  (
    g2977_n,
    g2507_p_spl_0,
    G2715_o2_n
  );


  and

  (
    g2978_p,
    G3485_o2_p_spl_00,
    G2720_o2_p_spl_0
  );


  or

  (
    g2978_n,
    G3485_o2_n_spl_,
    G2720_o2_n_spl_0
  );


  and

  (
    g2979_p,
    g2978_p,
    g2507_n_spl_0
  );


  or

  (
    g2979_n,
    g2978_n,
    g2507_p_spl_0
  );


  and

  (
    g2980_p,
    G3546_o2_p_spl_0,
    G3485_o2_p_spl_00
  );


  or

  (
    g2980_n,
    G3546_o2_n_spl_0,
    G3485_o2_n_spl_
  );


  and

  (
    g2981_p,
    g2980_p,
    g2507_n_spl_1
  );


  or

  (
    g2981_n,
    g2980_n,
    g2507_p_spl_
  );


  and

  (
    g2982_p,
    g2977_n,
    g2508_n
  );


  or

  (
    g2982_n,
    g2977_p,
    g2508_p_spl_
  );


  and

  (
    g2983_p,
    g2982_p,
    g2979_n
  );


  or

  (
    g2983_n,
    g2982_n,
    g2979_p
  );


  and

  (
    g2984_p,
    g2983_p_spl_0,
    g2981_n
  );


  or

  (
    g2984_n,
    g2983_n_spl_0,
    g2981_p
  );


  and

  (
    g2985_p,
    G4051_o2_n_spl_0,
    G3822_o2_n
  );


  or

  (
    g2985_n,
    G4051_o2_p_spl_0,
    G3822_o2_p
  );


  and

  (
    g2986_p,
    G2410_o2_n,
    n4284_lo_buf_o2_n
  );


  or

  (
    g2986_n,
    G2410_o2_p_spl_,
    n4284_lo_buf_o2_p_spl_
  );


  and

  (
    g2987_p,
    g2986_n_spl_,
    g2985_n_spl_
  );


  or

  (
    g2987_n,
    g2986_p_spl_,
    g2985_p_spl_
  );


  and

  (
    g2988_p,
    g2986_p_spl_,
    g2985_p_spl_
  );


  or

  (
    g2988_n,
    g2986_n_spl_,
    g2985_n_spl_
  );


  and

  (
    g2989_p,
    g2988_n,
    g2987_n
  );


  or

  (
    g2989_n,
    g2988_p,
    g2987_p
  );


  and

  (
    g2990_p,
    g2989_p_spl_,
    g2984_n_spl_
  );


  or

  (
    g2990_n,
    g2989_n_spl_,
    g2984_p_spl_
  );


  and

  (
    g2991_p,
    g2989_n_spl_,
    g2984_p_spl_
  );


  or

  (
    g2991_n,
    g2989_p_spl_,
    g2984_n_spl_
  );


  and

  (
    g2992_p,
    g2991_n,
    g2990_n
  );


  or

  (
    g2992_n,
    g2991_p,
    g2990_p
  );


  and

  (
    g2993_p,
    g2992_p,
    G3546_o2_n_spl_0
  );


  and

  (
    g2994_p,
    g2992_n,
    G3546_o2_p_spl_0
  );


  or

  (
    g2995_n,
    g2994_p,
    g2993_p
  );


  and

  (
    g2996_p,
    G4051_o2_n_spl_0,
    G2720_o2_p_spl_0
  );


  or

  (
    g2996_n,
    G4051_o2_p_spl_0,
    G2720_o2_n_spl_0
  );


  and

  (
    g2997_p,
    G4051_o2_p_spl_,
    G2720_o2_n_spl_
  );


  or

  (
    g2997_n,
    G4051_o2_n_spl_,
    G2720_o2_p_spl_1
  );


  and

  (
    g2998_p,
    g2997_n,
    g2996_n
  );


  or

  (
    g2998_n,
    g2997_p,
    g2996_p
  );


  and

  (
    g2999_p,
    g2998_p_spl_,
    g2983_p_spl_0
  );


  or

  (
    g2999_n,
    g2998_n_spl_,
    g2983_n_spl_0
  );


  and

  (
    g3000_p,
    g2998_n_spl_,
    g2983_n_spl_
  );


  or

  (
    g3000_n,
    g2998_p_spl_,
    g2983_p_spl_
  );


  and

  (
    g3001_p,
    g3000_n,
    g2999_n
  );


  or

  (
    g3001_n,
    g3000_p,
    g2999_p
  );


  and

  (
    g3002_p,
    g3001_p,
    G3546_o2_n_spl_
  );


  and

  (
    g3003_p,
    g3001_n,
    G3546_o2_p_spl_1
  );


  or

  (
    g3004_n,
    g3003_p,
    g3002_p
  );


  and

  (
    g3005_p,
    g2504_p_spl_0,
    G2832_o2_p_spl_
  );


  or

  (
    g3005_n,
    g2504_n_spl_00,
    G2832_o2_n
  );


  and

  (
    g3006_p,
    G3611_o2_p_spl_00,
    G2837_o2_p_spl_0
  );


  or

  (
    g3006_n,
    G3611_o2_n_spl_,
    G2837_o2_n_spl_0
  );


  and

  (
    g3007_p,
    g3006_p,
    g2504_p_spl_0
  );


  or

  (
    g3007_n,
    g3006_n,
    g2504_n_spl_00
  );


  and

  (
    g3008_p,
    G3658_o2_p_spl_0,
    G3611_o2_p_spl_00
  );


  or

  (
    g3008_n,
    G3658_o2_n_spl_0,
    G3611_o2_n_spl_
  );


  and

  (
    g3009_p,
    g3008_p,
    g2504_p_spl_1
  );


  or

  (
    g3009_n,
    g3008_n,
    g2504_n_spl_01
  );


  and

  (
    g3010_p,
    g3005_n,
    g2504_n_spl_01
  );


  or

  (
    g3010_n,
    g3005_p,
    g2504_p_spl_1
  );


  and

  (
    g3011_p,
    g3010_p,
    g3007_n
  );


  or

  (
    g3011_n,
    g3010_n,
    g3007_p
  );


  and

  (
    g3012_p,
    g3011_p_spl_0,
    g3009_n
  );


  or

  (
    g3012_n,
    g3011_n_spl_0,
    g3009_p
  );


  and

  (
    g3013_p,
    G4065_o2_n_spl_0,
    G3877_o2_n
  );


  or

  (
    g3013_n,
    G4065_o2_p_spl_0,
    G3877_o2_p
  );


  and

  (
    g3014_p,
    G2472_o2_n,
    n4356_lo_buf_o2_n
  );


  or

  (
    g3014_n,
    G2472_o2_p_spl_,
    n4356_lo_buf_o2_p_spl_
  );


  and

  (
    g3015_p,
    g3014_n_spl_,
    g3013_n_spl_
  );


  or

  (
    g3015_n,
    g3014_p_spl_,
    g3013_p_spl_
  );


  and

  (
    g3016_p,
    g3014_p_spl_,
    g3013_p_spl_
  );


  or

  (
    g3016_n,
    g3014_n_spl_,
    g3013_n_spl_
  );


  and

  (
    g3017_p,
    g3016_n,
    g3015_n
  );


  or

  (
    g3017_n,
    g3016_p,
    g3015_p
  );


  and

  (
    g3018_p,
    g3017_p_spl_,
    g3012_n_spl_
  );


  or

  (
    g3018_n,
    g3017_n_spl_,
    g3012_p_spl_
  );


  and

  (
    g3019_p,
    g3017_n_spl_,
    g3012_p_spl_
  );


  or

  (
    g3019_n,
    g3017_p_spl_,
    g3012_n_spl_
  );


  and

  (
    g3020_p,
    g3019_n,
    g3018_n
  );


  or

  (
    g3020_n,
    g3019_p,
    g3018_p
  );


  or

  (
    g3021_n,
    g3020_n,
    G3658_o2_p_spl_0
  );


  or

  (
    g3022_n,
    g3020_p,
    G3658_o2_n_spl_0
  );


  and

  (
    g3023_p,
    g3022_n,
    g3021_n
  );


  and

  (
    g3024_p,
    G4065_o2_n_spl_0,
    G2837_o2_p_spl_0
  );


  or

  (
    g3024_n,
    G4065_o2_p_spl_0,
    G2837_o2_n_spl_0
  );


  and

  (
    g3025_p,
    G4065_o2_p_spl_,
    G2837_o2_n_spl_
  );


  or

  (
    g3025_n,
    G4065_o2_n_spl_,
    G2837_o2_p_spl_1
  );


  and

  (
    g3026_p,
    g3025_n,
    g3024_n
  );


  or

  (
    g3026_n,
    g3025_p,
    g3024_p
  );


  and

  (
    g3027_p,
    g3026_p_spl_,
    g3011_p_spl_0
  );


  or

  (
    g3027_n,
    g3026_n_spl_,
    g3011_n_spl_0
  );


  and

  (
    g3028_p,
    g3026_n_spl_,
    g3011_n_spl_
  );


  or

  (
    g3028_n,
    g3026_p_spl_,
    g3011_p_spl_
  );


  and

  (
    g3029_p,
    g3028_n,
    g3027_n
  );


  or

  (
    g3029_n,
    g3028_p,
    g3027_p
  );


  or

  (
    g3030_n,
    g3029_n,
    G3658_o2_p_spl_1
  );


  or

  (
    g3031_n,
    g3029_p,
    G3658_o2_n_spl_
  );


  and

  (
    g3032_p,
    g3031_n,
    g3030_n
  );


  and

  (
    g3033_p,
    n4092_lo_buf_o2_p_spl_10,
    n3678_lo_p_spl_
  );


  and

  (
    g3034_p,
    n4092_lo_buf_o2_n_spl_1,
    n3690_lo_p
  );


  or

  (
    g3035_n,
    g3034_p,
    g3033_p
  );


  and

  (
    g3036_p,
    g2552_p_spl_0,
    n4374_lo_p_spl_0
  );


  or

  (
    g3036_n,
    g2552_n_spl_0,
    n4374_lo_n_spl_0
  );


  and

  (
    g3037_p,
    g2552_n_spl_0,
    n4374_lo_n_spl_0
  );


  or

  (
    g3037_n,
    g2552_p_spl_0,
    n4374_lo_p_spl_0
  );


  and

  (
    g3038_p,
    g3037_n,
    g3036_n
  );


  or

  (
    g3038_n,
    g3037_p,
    g3036_p
  );


  and

  (
    g3039_p,
    g2555_p,
    n4242_lo_p_spl_0
  );


  and

  (
    g3040_p,
    g2555_n_spl_0,
    n4242_lo_n
  );


  or

  (
    g3041_n,
    g3040_p,
    g3039_p
  );


  and

  (
    g3042_p,
    g2561_p,
    n4326_lo_p_spl_0
  );


  and

  (
    g3043_p,
    g2561_n_spl_0,
    n4326_lo_n
  );


  or

  (
    g3044_n,
    g3043_p,
    g3042_p
  );


  and

  (
    g3045_p,
    g2558_p,
    n4338_lo_p_spl_0
  );


  and

  (
    g3046_p,
    g2558_n_spl_0,
    n4338_lo_n
  );


  or

  (
    g3047_n,
    g3046_p,
    g3045_p
  );


  and

  (
    g3048_p,
    n4248_lo_buf_o2_p_spl_0,
    n3801_lo_n_spl_0
  );


  and

  (
    g3049_p,
    g3048_p,
    n3840_lo_buf_o2_n
  );


  and

  (
    g3050_p,
    n4248_lo_buf_o2_p_spl_0,
    n3813_lo_n_spl_0
  );


  and

  (
    g3051_p,
    g3050_p,
    n3840_lo_buf_o2_p_spl_0
  );


  and

  (
    g3052_p,
    n4293_lo_p_spl_0,
    n3801_lo_n_spl_0
  );


  and

  (
    g3053_p,
    g3052_p,
    n3753_lo_n_spl_
  );


  and

  (
    g3054_p,
    n4293_lo_p_spl_1,
    n3813_lo_n_spl_0
  );


  and

  (
    g3055_p,
    g3054_p,
    n3753_lo_p_spl_00
  );


  and

  (
    g3056_p,
    n4365_lo_p_spl_0,
    n3801_lo_n_spl_
  );


  and

  (
    g3057_p,
    g3056_p,
    n4053_lo_n_spl_
  );


  and

  (
    g3058_p,
    n4365_lo_p_spl_1,
    n3813_lo_n_spl_
  );


  and

  (
    g3059_p,
    g3058_p,
    n4053_lo_p_spl_00
  );


  or

  (
    g3060_n,
    g2552_p_spl_,
    n4374_lo_n_spl_
  );


  and

  (
    g3061_p,
    g2555_n_spl_0,
    n4242_lo_p_spl_0
  );


  and

  (
    g3062_p,
    g2561_n_spl_0,
    n4326_lo_p_spl_0
  );


  and

  (
    g3063_p,
    g2558_n_spl_0,
    n4338_lo_p_spl_0
  );


  and

  (
    g3064_p,
    g2672_n_spl_0,
    n4305_lo_n_spl_
  );


  and

  (
    g3065_p,
    G4697_o2_p_spl_,
    G4131_o2_n_spl_
  );


  or

  (
    g3065_n,
    G4697_o2_n_spl_,
    G4131_o2_p_spl_
  );


  and

  (
    g3066_p,
    G4697_o2_n_spl_,
    G4131_o2_p_spl_
  );


  or

  (
    g3066_n,
    G4697_o2_p_spl_,
    G4131_o2_n_spl_
  );


  and

  (
    g3067_p,
    g3066_n,
    g3065_n
  );


  or

  (
    g3067_n,
    g3066_p,
    g3065_p
  );


  and

  (
    g3068_p,
    g3067_p_spl_,
    G3552_o2_n_spl_1
  );


  or

  (
    g3068_n,
    g3067_n_spl_,
    G3552_o2_p_spl_0
  );


  and

  (
    g3069_p,
    g3067_n_spl_,
    G3552_o2_p_spl_1
  );


  or

  (
    g3069_n,
    g3067_p_spl_,
    G3552_o2_n_spl_1
  );


  and

  (
    g3070_p,
    g3069_n,
    g3068_n
  );


  or

  (
    g3070_n,
    g3069_p,
    g3068_p
  );


  and

  (
    g3071_p,
    g3070_p,
    G3533_o2_n_spl_
  );


  and

  (
    g3072_p,
    g3070_n,
    G3533_o2_p_spl_0
  );


  or

  (
    g3073_n,
    g3072_p,
    g3071_p
  );


  and

  (
    g3074_p,
    g3073_n_spl_,
    g2675_n_spl_00
  );


  and

  (
    g3075_p,
    G4706_o2_n_spl_,
    G4170_o2_n_spl_
  );


  or

  (
    g3075_n,
    G4706_o2_p_spl_,
    G4170_o2_p_spl_
  );


  and

  (
    g3076_p,
    G4706_o2_p_spl_,
    G4170_o2_p_spl_
  );


  or

  (
    g3076_n,
    G4706_o2_n_spl_,
    G4170_o2_n_spl_
  );


  and

  (
    g3077_p,
    g3076_n,
    g3075_n
  );


  or

  (
    g3077_n,
    g3076_p,
    g3075_p
  );


  and

  (
    g3078_p,
    g3077_p_spl_,
    n2647_inv_p_spl_0
  );


  or

  (
    g3078_n,
    g3077_n_spl_,
    n2647_inv_n_spl_1
  );


  and

  (
    g3079_p,
    g3077_n_spl_,
    n2647_inv_n_spl_1
  );


  or

  (
    g3079_n,
    g3077_p_spl_,
    n2647_inv_p_spl_1
  );


  and

  (
    g3080_p,
    g3079_n,
    g3078_n
  );


  or

  (
    g3080_n,
    g3079_p,
    g3078_p
  );


  and

  (
    g3081_p,
    g3080_p,
    G3645_o2_n_spl_
  );


  and

  (
    g3082_p,
    g3080_n,
    G3645_o2_p_spl_0
  );


  or

  (
    g3083_n,
    g3082_p,
    g3081_p
  );


  and

  (
    g3084_p,
    g3083_n_spl_,
    g2678_n_spl_00
  );


  or

  (
    g3085_n,
    g2672_n_spl_0,
    n4305_lo_n_spl_
  );


  or

  (
    g3086_n,
    g3073_n_spl_,
    g2675_n_spl_00
  );


  or

  (
    g3087_n,
    g3083_n_spl_,
    g2678_n_spl_00
  );


  and

  (
    g3088_p,
    G1821_o2_p_spl_,
    n3957_lo_p_spl_
  );


  and

  (
    g3089_p,
    G1060_o2_n_spl_,
    n3969_lo_p_spl_
  );


  or

  (
    g3090_n,
    g3089_p,
    g3088_p
  );


  and

  (
    g3091_p,
    g2684_p,
    n4278_lo_p_spl_0
  );


  and

  (
    g3092_p,
    g2684_n_spl_0,
    n4278_lo_n
  );


  or

  (
    g3093_n,
    g3092_p,
    g3091_p
  );


  and

  (
    g3094_p,
    g2681_p,
    n4350_lo_p_spl_0
  );


  and

  (
    g3095_p,
    g2681_n_spl_0,
    n4350_lo_n
  );


  or

  (
    g3096_n,
    g3095_p,
    g3094_p
  );


  and

  (
    g3097_p,
    n4080_lo_buf_o2_n_spl_1,
    n3990_lo_p
  );


  and

  (
    g3098_p,
    g2536_n_spl_0,
    g2522_p_spl_0
  );


  or

  (
    g3098_n,
    g2536_p_spl_0,
    g2522_n_spl_
  );


  and

  (
    g3099_p,
    g3098_p_spl_,
    g3041_n_spl_00
  );


  and

  (
    g3100_p,
    g2542_n_spl_0,
    g2523_p_spl_0
  );


  or

  (
    g3100_n,
    g2542_p_spl_0,
    g2523_n_spl_
  );


  or

  (
    g3101_n,
    g3100_n_spl_,
    g3038_p_spl_0
  );


  and

  (
    g3102_p,
    g2539_n_spl_00,
    g2536_n_spl_0
  );


  or

  (
    g3102_n,
    g2539_p_spl_0,
    g2536_p_spl_0
  );


  and

  (
    g3103_p,
    g3102_p,
    g2533_p_spl_00
  );


  or

  (
    g3103_n,
    g3102_n,
    g2533_n_spl_0
  );


  and

  (
    g3104_p,
    g3103_p_spl_,
    g3041_n_spl_00
  );


  and

  (
    g3105_p,
    n4080_lo_buf_o2_p_spl_10,
    n3978_lo_p_spl_
  );


  and

  (
    g3106_p,
    g2550_n_spl_0,
    g2536_n_spl_1
  );


  or

  (
    g3106_n,
    g2550_p,
    g2536_p_spl_
  );


  and

  (
    g3107_p,
    g3106_p_spl_,
    g3041_n_spl_0
  );


  and

  (
    g3108_p,
    g3107_p,
    g2539_n_spl_00
  );


  and

  (
    g3109_p,
    g2545_n_spl_0,
    g2542_n_spl_0
  );


  or

  (
    g3109_n,
    g2545_p_spl_0,
    g2542_p_spl_0
  );


  and

  (
    g3110_p,
    g3109_p,
    g2517_p_spl_0
  );


  or

  (
    g3110_n,
    g3109_n,
    g2517_n_spl_00
  );


  or

  (
    g3111_n,
    g3110_n_spl_,
    g3038_p_spl_0
  );


  or

  (
    g3112_n,
    g2542_p_spl_,
    g2517_n_spl_00
  );


  or

  (
    g3113_n,
    g3112_n_spl_,
    g3038_p_spl_1
  );


  or

  (
    g3114_n,
    g3113_n,
    g2545_p_spl_0
  );


  and

  (
    g3115_p,
    g3041_n_spl_1,
    g2546_p_spl_0
  );


  or

  (
    g3116_n,
    g3038_p_spl_1,
    g2547_n_spl_
  );


  or

  (
    g3117_n,
    g3112_n_spl_,
    g2545_p_spl_1
  );


  and

  (
    g3118_p,
    g3100_n_spl_,
    g2547_n_spl_
  );


  or

  (
    g3118_n,
    g3100_p,
    g2547_p_spl_
  );


  and

  (
    g3119_p,
    g3118_p,
    g3110_n_spl_
  );


  or

  (
    g3119_n,
    g3118_n,
    g3110_p
  );


  and

  (
    g3120_p,
    g3119_p_spl_0,
    g3117_n
  );


  and

  (
    g3121_p,
    g2545_n_spl_0,
    g2517_p_spl_0
  );


  or

  (
    g3121_n,
    g2545_p_spl_1,
    g2517_n_spl_01
  );


  and

  (
    g3122_p,
    g3121_n,
    g2523_n_spl_
  );


  or

  (
    g3122_n,
    g3121_p_spl_,
    g2523_p_spl_0
  );


  or

  (
    g3123_n,
    g3122_n_spl_,
    g3121_p_spl_
  );


  or

  (
    g3124_n,
    g3123_n_spl_,
    g3120_p_spl_
  );


  and

  (
    g3125_p,
    g2539_n_spl_01,
    g2533_p_spl_00
  );


  or

  (
    g3125_n,
    g2539_p_spl_0,
    g2533_n_spl_0
  );


  and

  (
    g3126_p,
    g3125_n,
    g2522_n_spl_
  );


  or

  (
    g3126_n,
    g3125_p,
    g2522_p_spl_0
  );


  and

  (
    g3127_p,
    g2550_n_spl_0,
    g2539_n_spl_01
  );


  or

  (
    g3128_n,
    g3127_p,
    g3126_n_spl_
  );


  and

  (
    g3129_p,
    g3106_p_spl_,
    g2539_n_spl_1
  );


  or

  (
    g3129_n,
    g3106_n,
    g2539_p_spl_
  );


  and

  (
    g3130_p,
    g3098_n,
    g2546_n
  );


  or

  (
    g3130_n,
    g3098_p_spl_,
    g2546_p_spl_0
  );


  and

  (
    g3131_p,
    g3130_p,
    g3103_n
  );


  or

  (
    g3131_n,
    g3130_n,
    g3103_p_spl_
  );


  and

  (
    g3132_p,
    g3131_p_spl_0,
    g3129_n
  );


  or

  (
    g3132_n,
    g3131_n_spl_0,
    g3129_p
  );


  and

  (
    g3133_p,
    n4224_lo_buf_o2_n_spl_1,
    G2379_o2_n_spl_1
  );


  or

  (
    g3133_n,
    n4224_lo_buf_o2_p_spl_1,
    G2379_o2_p_spl_1
  );


  or

  (
    g3134_n,
    g3133_p,
    g3132_p
  );


  or

  (
    g3135_n,
    g3133_n,
    g3132_n
  );


  and

  (
    g3136_p,
    g3135_n,
    g3134_n
  );


  and

  (
    g3137_p,
    g3136_p_spl_,
    g3128_n_spl_
  );


  and

  (
    g3138_p,
    g3123_n_spl_,
    g3120_p_spl_
  );


  or

  (
    g3139_n,
    g3136_p_spl_,
    g3128_n_spl_
  );


  and

  (
    g3140_p,
    g3093_n_spl_,
    g3044_n_spl_0
  );


  and

  (
    g3141_p,
    g3096_n_spl_,
    g3047_n_spl_0
  );


  or

  (
    g3142_n,
    g3115_p_spl_,
    g3061_p_spl_
  );


  or

  (
    g3143_n,
    g3142_n,
    g3099_p_spl_
  );


  or

  (
    g3144_n,
    g3143_n,
    g3104_p_spl_
  );


  and

  (
    g3145_p,
    g3116_n_spl_,
    g3060_n_spl_
  );


  and

  (
    g3146_p,
    g3145_p,
    g3101_n_spl_
  );


  and

  (
    g3147_p,
    g3146_p,
    g3111_n_spl_
  );


  and

  (
    g3148_p,
    g3044_n_spl_0,
    g2947_p_spl_
  );


  or

  (
    g3149_n,
    g3148_p,
    g3062_p_spl_
  );


  and

  (
    g3150_p,
    g3047_n_spl_0,
    g2948_p_spl_
  );


  or

  (
    g3151_n,
    g3150_p,
    g3063_p_spl_
  );


  and

  (
    g3152_p,
    g3131_p_spl_0,
    g2533_p_spl_0
  );


  or

  (
    g3152_n,
    g3131_n_spl_0,
    g2533_n_spl_1
  );


  and

  (
    g3153_p,
    g3131_n_spl_,
    g2533_n_spl_1
  );


  or

  (
    g3153_n,
    g3131_p_spl_,
    g2533_p_spl_1
  );


  and

  (
    g3154_p,
    g3153_n,
    g3152_n
  );


  or

  (
    g3154_n,
    g3153_p,
    g3152_p
  );


  or

  (
    g3155_n,
    g3154_n,
    g3126_n_spl_
  );


  or

  (
    g3156_n,
    g3154_p,
    g3126_p
  );


  and

  (
    g3157_p,
    g3156_n,
    g3155_n
  );


  and

  (
    g3158_p,
    g3119_p_spl_0,
    g2517_p_spl_1
  );


  or

  (
    g3158_n,
    g3119_n_spl_,
    g2517_n_spl_01
  );


  and

  (
    g3159_p,
    g3119_n_spl_,
    g2517_n_spl_10
  );


  or

  (
    g3159_n,
    g3119_p_spl_,
    g2517_p_spl_1
  );


  and

  (
    g3160_p,
    g3159_n,
    g3158_n
  );


  or

  (
    g3160_n,
    g3159_p,
    g3158_p
  );


  and

  (
    g3161_p,
    g3160_p,
    g3122_p
  );


  and

  (
    g3162_p,
    g3160_n,
    g3122_n_spl_
  );


  or

  (
    g3163_n,
    g3162_p,
    g3161_p
  );


  and

  (
    g3164_p,
    G126_p_spl_,
    G123_p_spl_00
  );


  and

  (
    g3165_p,
    G127_p_spl_,
    G123_n_spl_
  );


  or

  (
    g3166_n,
    g3165_p,
    g3164_p
  );


  and

  (
    g3167_p,
    G128_p_spl_,
    G123_p_spl_00
  );


  and

  (
    g3168_p,
    G129_p_spl_,
    G123_n_spl_
  );


  or

  (
    g3169_n,
    g3168_p,
    g3167_p
  );


  and

  (
    g3170_p,
    G124_p_spl_00,
    G105_p_spl_
  );


  and

  (
    g3171_p,
    G124_n_spl_0,
    G106_p
  );


  or

  (
    g3172_n,
    g3171_p,
    g3170_p
  );


  and

  (
    g3173_p,
    G124_p_spl_00,
    G107_p_spl_
  );


  and

  (
    g3174_p,
    G124_n_spl_0,
    G108_p
  );


  or

  (
    g3175_n,
    g3174_p,
    g3173_p
  );


  and

  (
    g3176_p,
    G124_p_spl_01,
    G109_p_spl_
  );


  and

  (
    g3177_p,
    G124_n_spl_,
    G110_p
  );


  or

  (
    g3178_n,
    g3177_p,
    g3176_p
  );


  buf

  (
    G5193,
    n3399_lo_n_spl_1
  );


  buf

  (
    G5194,
    n3963_lo_n_spl_
  );


  buf

  (
    G5195,
    n4587_lo_n_spl_
  );


  buf

  (
    G5196,
    n4419_lo_n_spl_0
  );


  buf

  (
    G5197,
    n4131_lo_n
  );


  buf

  (
    G5198,
    n4179_lo_n
  );


  buf

  (
    G5199,
    g1192_p
  );


  buf

  (
    G5200,
    n4431_lo_n
  );


  buf

  (
    G5201,
    n4419_lo_n_spl_0
  );


  buf

  (
    G5202,
    n4419_lo_n_spl_
  );


  buf

  (
    G5203,
    n4107_lo_n
  );


  buf

  (
    G5204,
    n4155_lo_n
  );


  buf

  (
    G5205,
    g1193_p
  );


  buf

  (
    G5206,
    n3795_lo_n_spl_
  );


  buf

  (
    G5207,
    n4443_lo_n_spl_
  );


  buf

  (
    G5208,
    n4479_lo_n_spl_
  );


  buf

  (
    G5209,
    n4467_lo_n_spl_
  );


  buf

  (
    G5210,
    g1194_p
  );


  buf

  (
    G5211,
    g1195_p
  );


  buf

  (
    G5212,
    g1196_n
  );


  buf

  (
    G5213,
    g1197_n
  );


  buf

  (
    G5214,
    n3375_lo_p_spl_111
  );


  buf

  (
    G5215,
    n3399_lo_p_spl_
  );


  buf

  (
    G5216,
    n2619_lo_p_spl_
  );


  buf

  (
    G5217,
    n4431_lo_p_spl_
  );


  buf

  (
    G5218,
    n3975_lo_p
  );


  buf

  (
    G5219,
    n4431_lo_p_spl_
  );


  buf

  (
    G5220,
    g1199_n
  );


  buf

  (
    G5221,
    g1198_n_spl_11
  );


  buf

  (
    G5222,
    n2619_lo_n_spl_0
  );


  buf

  (
    G5223,
    n2619_lo_n_spl_0
  );


  buf

  (
    G5224,
    n2619_lo_n_spl_1
  );


  buf

  (
    G5225,
    n2619_lo_n_spl_1
  );


  buf

  (
    G5226,
    n3975_lo_n_spl_
  );


  buf

  (
    G5227,
    n3975_lo_n_spl_
  );


  buf

  (
    G5228,
    g1203_n
  );


  buf

  (
    G5229,
    g1207_n_spl_
  );


  buf

  (
    G5230,
    g1207_n_spl_
  );


  buf

  (
    G5231,
    g1211_n
  );


  not

  (
    G5232,
    g1221_n
  );


  not

  (
    G5233,
    g1229_n
  );


  not

  (
    G5234,
    g1237_n
  );


  not

  (
    G5235,
    g1245_n
  );


  not

  (
    G5236,
    g1312_n
  );


  not

  (
    G5237,
    g1400_n
  );


  not

  (
    G5238,
    g1404_n
  );


  not

  (
    G5239,
    g1412_n
  );


  not

  (
    G5240,
    g1416_n
  );


  not

  (
    G5241,
    g1424_n
  );


  not

  (
    G5242,
    g1449_n_spl_
  );


  not

  (
    G5243,
    g1474_n_spl_
  );


  not

  (
    G5244,
    g1486_p
  );


  not

  (
    G5245,
    g1512_p
  );


  not

  (
    G5246,
    g1538_p
  );


  not

  (
    G5247,
    g1549_p
  );


  not

  (
    G5248,
    g1563_n_spl_1
  );


  not

  (
    G5249,
    g1576_n_spl_1
  );


  not

  (
    G5250,
    g1587_n_spl_1
  );


  buf

  (
    G5251,
    g1601_p_spl_
  );


  buf

  (
    G5252,
    g1612_n
  );


  not

  (
    G5253,
    g1635_n_spl_1
  );


  not

  (
    G5254,
    g1649_n_spl_1
  );


  not

  (
    G5255,
    g1664_n_spl_1
  );


  buf

  (
    G5256,
    g1675_n
  );


  not

  (
    G5257,
    g1699_n_spl_1
  );


  not

  (
    G5258,
    g1713_n_spl_1
  );


  not

  (
    G5259,
    g1728_n_spl_1
  );


  not

  (
    G5260,
    g1740_n_spl_1
  );


  not

  (
    G5261,
    g1765_n_spl_
  );


  not

  (
    G5262,
    g1790_n_spl_
  );


  not

  (
    G5263,
    g1835_n
  );


  not

  (
    G5264,
    g1866_n
  );


  buf

  (
    G5265,
    g1878_p
  );


  buf

  (
    G5266,
    g1890_p
  );


  buf

  (
    G5267,
    g1901_n
  );


  buf

  (
    G5268,
    g1912_n
  );


  buf

  (
    G5269,
    g1923_n
  );


  buf

  (
    G5270,
    g1934_n
  );


  buf

  (
    G5271,
    g1945_n
  );


  buf

  (
    G5272,
    g1956_n
  );


  buf

  (
    G5273,
    g1967_n
  );


  buf

  (
    G5274,
    g1978_n
  );


  buf

  (
    G5275,
    g1990_p
  );


  buf

  (
    G5276,
    g2002_p
  );


  buf

  (
    G5277,
    g2014_p
  );


  buf

  (
    G5278,
    g2026_p
  );


  buf

  (
    G5279,
    g2038_p
  );


  buf

  (
    G5280,
    g2050_p
  );


  buf

  (
    G5281,
    g2062_p
  );


  buf

  (
    G5282,
    g2074_p
  );


  buf

  (
    G5283,
    g2091_p
  );


  buf

  (
    G5284,
    g2095_n
  );


  not

  (
    G5285,
    g2103_n_spl_1
  );


  not

  (
    G5286,
    g2111_n_spl_1
  );


  not

  (
    G5287,
    g2119_n_spl_1
  );


  not

  (
    G5288,
    g2127_n_spl_1
  );


  not

  (
    G5289,
    g2136_n
  );


  not

  (
    G5290,
    g2154_n_spl_1
  );


  not

  (
    G5291,
    g2162_n_spl_1
  );


  not

  (
    G5292,
    g2170_n_spl_1
  );


  not

  (
    G5293,
    g2178_n_spl_1
  );


  buf

  (
    G5294,
    g2189_n
  );


  buf

  (
    G5295,
    g2200_n
  );


  buf

  (
    G5296,
    g2211_n
  );


  buf

  (
    G5297,
    g2222_n
  );


  buf

  (
    G5298,
    g2233_n
  );


  buf

  (
    G5299,
    g2244_n
  );


  buf

  (
    G5300,
    g2255_n
  );


  buf

  (
    G5301,
    g2266_n
  );


  buf

  (
    G5302,
    g2278_p
  );


  buf

  (
    G5303,
    g2290_p
  );


  buf

  (
    G5304,
    g2302_p
  );


  buf

  (
    G5305,
    g2314_p
  );


  buf

  (
    G5306,
    g2326_p
  );


  buf

  (
    G5307,
    g2338_p
  );


  buf

  (
    G5308,
    g2350_p
  );


  buf

  (
    G5309,
    g2362_p
  );


  not

  (
    G5310,
    g2378_p
  );


  not

  (
    G5311,
    g2393_p
  );


  buf

  (
    G5312,
    g2416_n
  );


  buf

  (
    G5313,
    g2427_n
  );


  not

  (
    G5314,
    g2439_p
  );


  not

  (
    G5315,
    g2451_p
  );


  buf

  (
    n2610_li,
    G1_p
  );


  buf

  (
    n2613_li,
    n2610_lo_p
  );


  buf

  (
    n2616_li,
    n2613_lo_p
  );


  buf

  (
    n2619_li,
    n2616_lo_p
  );


  buf

  (
    n2622_li,
    G2_p
  );


  buf

  (
    n2625_li,
    n2622_lo_p
  );


  buf

  (
    n2628_li,
    n2625_lo_p
  );


  buf

  (
    n2631_li,
    n2628_lo_p
  );


  buf

  (
    n2634_li,
    G3_p
  );


  buf

  (
    n2637_li,
    n2634_lo_p
  );


  buf

  (
    n2640_li,
    n2637_lo_p
  );


  buf

  (
    n2643_li,
    n2640_lo_p
  );


  buf

  (
    n2646_li,
    G4_p
  );


  buf

  (
    n2649_li,
    n2646_lo_p
  );


  buf

  (
    n2652_li,
    n2649_lo_p
  );


  buf

  (
    n2655_li,
    n2652_lo_p
  );


  buf

  (
    n2658_li,
    G5_p
  );


  buf

  (
    n2661_li,
    n2658_lo_p
  );


  buf

  (
    n2664_li,
    n2661_lo_p
  );


  buf

  (
    n2667_li,
    n2664_lo_p
  );


  buf

  (
    n2670_li,
    G6_p
  );


  buf

  (
    n2673_li,
    n2670_lo_p
  );


  buf

  (
    n2676_li,
    n2673_lo_p
  );


  buf

  (
    n2679_li,
    n2676_lo_p
  );


  buf

  (
    n2682_li,
    G7_p
  );


  buf

  (
    n2685_li,
    n2682_lo_p
  );


  buf

  (
    n2688_li,
    n2685_lo_p
  );


  buf

  (
    n2691_li,
    n2688_lo_p
  );


  buf

  (
    n2694_li,
    G8_p
  );


  buf

  (
    n2697_li,
    n2694_lo_p
  );


  buf

  (
    n2700_li,
    n2697_lo_p
  );


  buf

  (
    n2703_li,
    n2700_lo_p
  );


  buf

  (
    n2706_li,
    G9_p
  );


  buf

  (
    n2709_li,
    n2706_lo_p
  );


  buf

  (
    n2712_li,
    n2709_lo_p
  );


  buf

  (
    n2715_li,
    n2712_lo_p
  );


  buf

  (
    n2718_li,
    G10_p
  );


  buf

  (
    n2721_li,
    n2718_lo_p
  );


  buf

  (
    n2724_li,
    n2721_lo_p
  );


  buf

  (
    n2727_li,
    n2724_lo_p
  );


  buf

  (
    n2730_li,
    G11_p
  );


  buf

  (
    n2733_li,
    n2730_lo_p
  );


  buf

  (
    n2736_li,
    n2733_lo_p
  );


  buf

  (
    n2739_li,
    n2736_lo_p
  );


  buf

  (
    n2742_li,
    G12_p
  );


  buf

  (
    n2745_li,
    n2742_lo_p
  );


  buf

  (
    n2748_li,
    n2745_lo_p
  );


  buf

  (
    n2751_li,
    n2748_lo_p
  );


  buf

  (
    n2754_li,
    G13_p
  );


  buf

  (
    n2757_li,
    n2754_lo_p
  );


  buf

  (
    n2760_li,
    n2757_lo_p
  );


  buf

  (
    n2763_li,
    n2760_lo_p
  );


  buf

  (
    n2766_li,
    G14_p
  );


  buf

  (
    n2769_li,
    n2766_lo_p
  );


  buf

  (
    n2772_li,
    n2769_lo_p
  );


  buf

  (
    n2775_li,
    n2772_lo_p
  );


  buf

  (
    n2778_li,
    G15_p
  );


  buf

  (
    n2781_li,
    n2778_lo_p
  );


  buf

  (
    n2784_li,
    n2781_lo_p
  );


  buf

  (
    n2787_li,
    n2784_lo_p
  );


  buf

  (
    n2790_li,
    G16_p
  );


  buf

  (
    n2793_li,
    n2790_lo_p
  );


  buf

  (
    n2796_li,
    n2793_lo_p
  );


  buf

  (
    n2799_li,
    n2796_lo_p
  );


  buf

  (
    n2802_li,
    G17_p
  );


  buf

  (
    n2805_li,
    n2802_lo_p
  );


  buf

  (
    n2808_li,
    n2805_lo_p
  );


  buf

  (
    n2811_li,
    n2808_lo_p
  );


  buf

  (
    n2814_li,
    G18_p
  );


  buf

  (
    n2817_li,
    n2814_lo_p
  );


  buf

  (
    n2820_li,
    n2817_lo_p
  );


  buf

  (
    n2823_li,
    n2820_lo_p
  );


  buf

  (
    n2826_li,
    G19_p
  );


  buf

  (
    n2829_li,
    n2826_lo_p
  );


  buf

  (
    n2832_li,
    n2829_lo_p
  );


  buf

  (
    n2835_li,
    n2832_lo_p
  );


  buf

  (
    n2838_li,
    G20_p
  );


  buf

  (
    n2841_li,
    n2838_lo_p
  );


  buf

  (
    n2844_li,
    n2841_lo_p
  );


  buf

  (
    n2847_li,
    n2844_lo_p
  );


  buf

  (
    n2850_li,
    G21_p
  );


  buf

  (
    n2853_li,
    n2850_lo_p
  );


  buf

  (
    n2856_li,
    n2853_lo_p
  );


  buf

  (
    n2859_li,
    n2856_lo_p
  );


  buf

  (
    n2862_li,
    G22_p
  );


  buf

  (
    n2865_li,
    n2862_lo_p
  );


  buf

  (
    n2868_li,
    n2865_lo_p
  );


  buf

  (
    n2871_li,
    n2868_lo_p
  );


  buf

  (
    n2874_li,
    G23_p
  );


  buf

  (
    n2877_li,
    n2874_lo_p
  );


  buf

  (
    n2880_li,
    n2877_lo_p
  );


  buf

  (
    n2883_li,
    n2880_lo_p
  );


  buf

  (
    n2886_li,
    G24_p
  );


  buf

  (
    n2889_li,
    n2886_lo_p
  );


  buf

  (
    n2892_li,
    n2889_lo_p
  );


  buf

  (
    n2895_li,
    n2892_lo_p
  );


  buf

  (
    n2898_li,
    G25_p
  );


  buf

  (
    n2901_li,
    n2898_lo_p
  );


  buf

  (
    n2904_li,
    n2901_lo_p
  );


  buf

  (
    n2907_li,
    n2904_lo_p
  );


  buf

  (
    n2910_li,
    G26_p
  );


  buf

  (
    n2913_li,
    n2910_lo_p
  );


  buf

  (
    n2916_li,
    n2913_lo_p
  );


  buf

  (
    n2919_li,
    n2916_lo_p
  );


  buf

  (
    n2922_li,
    G27_p
  );


  buf

  (
    n2925_li,
    n2922_lo_p
  );


  buf

  (
    n2928_li,
    n2925_lo_p
  );


  buf

  (
    n2931_li,
    n2928_lo_p
  );


  buf

  (
    n2934_li,
    G28_p
  );


  buf

  (
    n2937_li,
    n2934_lo_p
  );


  buf

  (
    n2940_li,
    n2937_lo_p
  );


  buf

  (
    n2943_li,
    n2940_lo_p
  );


  buf

  (
    n2946_li,
    G29_p
  );


  buf

  (
    n2949_li,
    n2946_lo_p
  );


  buf

  (
    n2952_li,
    n2949_lo_p
  );


  buf

  (
    n2955_li,
    n2952_lo_p
  );


  buf

  (
    n2958_li,
    G30_p
  );


  buf

  (
    n2961_li,
    n2958_lo_p
  );


  buf

  (
    n2964_li,
    n2961_lo_p
  );


  buf

  (
    n2967_li,
    n2964_lo_p
  );


  buf

  (
    n2970_li,
    G31_p
  );


  buf

  (
    n2973_li,
    n2970_lo_p
  );


  buf

  (
    n2976_li,
    n2973_lo_p
  );


  buf

  (
    n2979_li,
    n2976_lo_p
  );


  buf

  (
    n2982_li,
    G32_p
  );


  buf

  (
    n2985_li,
    n2982_lo_p
  );


  buf

  (
    n2988_li,
    n2985_lo_p
  );


  buf

  (
    n2991_li,
    n2988_lo_p
  );


  buf

  (
    n2994_li,
    G33_p
  );


  buf

  (
    n2997_li,
    n2994_lo_p
  );


  buf

  (
    n3000_li,
    n2997_lo_p
  );


  buf

  (
    n3003_li,
    n3000_lo_p
  );


  buf

  (
    n3006_li,
    G34_p
  );


  buf

  (
    n3009_li,
    n3006_lo_p
  );


  buf

  (
    n3012_li,
    n3009_lo_p
  );


  buf

  (
    n3015_li,
    n3012_lo_p
  );


  buf

  (
    n3018_li,
    G35_p
  );


  buf

  (
    n3021_li,
    n3018_lo_p
  );


  buf

  (
    n3024_li,
    n3021_lo_p
  );


  buf

  (
    n3027_li,
    n3024_lo_p
  );


  buf

  (
    n3030_li,
    G36_p
  );


  buf

  (
    n3033_li,
    n3030_lo_p
  );


  buf

  (
    n3036_li,
    n3033_lo_p
  );


  buf

  (
    n3039_li,
    n3036_lo_p
  );


  buf

  (
    n3042_li,
    G37_p
  );


  buf

  (
    n3045_li,
    n3042_lo_p
  );


  buf

  (
    n3048_li,
    n3045_lo_p
  );


  buf

  (
    n3051_li,
    n3048_lo_p
  );


  buf

  (
    n3054_li,
    G38_p
  );


  buf

  (
    n3057_li,
    n3054_lo_p
  );


  buf

  (
    n3060_li,
    n3057_lo_p
  );


  buf

  (
    n3063_li,
    n3060_lo_p
  );


  buf

  (
    n3066_li,
    G39_p
  );


  buf

  (
    n3069_li,
    n3066_lo_p
  );


  buf

  (
    n3072_li,
    n3069_lo_p
  );


  buf

  (
    n3075_li,
    n3072_lo_p
  );


  buf

  (
    n3078_li,
    G40_p
  );


  buf

  (
    n3081_li,
    n3078_lo_p
  );


  buf

  (
    n3084_li,
    n3081_lo_p
  );


  buf

  (
    n3087_li,
    n3084_lo_p
  );


  buf

  (
    n3090_li,
    G41_p
  );


  buf

  (
    n3093_li,
    n3090_lo_p
  );


  buf

  (
    n3096_li,
    n3093_lo_p
  );


  buf

  (
    n3099_li,
    n3096_lo_p
  );


  buf

  (
    n3102_li,
    G42_p
  );


  buf

  (
    n3105_li,
    n3102_lo_p
  );


  buf

  (
    n3108_li,
    n3105_lo_p
  );


  buf

  (
    n3111_li,
    n3108_lo_p
  );


  buf

  (
    n3114_li,
    G43_p
  );


  buf

  (
    n3117_li,
    n3114_lo_p
  );


  buf

  (
    n3120_li,
    n3117_lo_p
  );


  buf

  (
    n3123_li,
    n3120_lo_p
  );


  buf

  (
    n3126_li,
    G44_p
  );


  buf

  (
    n3129_li,
    n3126_lo_p
  );


  buf

  (
    n3132_li,
    n3129_lo_p
  );


  buf

  (
    n3135_li,
    n3132_lo_p
  );


  buf

  (
    n3138_li,
    G45_p
  );


  buf

  (
    n3141_li,
    n3138_lo_p
  );


  buf

  (
    n3144_li,
    n3141_lo_p
  );


  buf

  (
    n3147_li,
    n3144_lo_p
  );


  buf

  (
    n3150_li,
    G46_p
  );


  buf

  (
    n3153_li,
    n3150_lo_p
  );


  buf

  (
    n3156_li,
    n3153_lo_p
  );


  buf

  (
    n3159_li,
    n3156_lo_p
  );


  buf

  (
    n3162_li,
    G47_p
  );


  buf

  (
    n3165_li,
    n3162_lo_p
  );


  buf

  (
    n3168_li,
    n3165_lo_p
  );


  buf

  (
    n3171_li,
    n3168_lo_p
  );


  buf

  (
    n3174_li,
    G48_p
  );


  buf

  (
    n3177_li,
    n3174_lo_p
  );


  buf

  (
    n3180_li,
    n3177_lo_p
  );


  buf

  (
    n3183_li,
    n3180_lo_p
  );


  buf

  (
    n3186_li,
    G49_p
  );


  buf

  (
    n3189_li,
    n3186_lo_p
  );


  buf

  (
    n3192_li,
    n3189_lo_p
  );


  buf

  (
    n3195_li,
    n3192_lo_p
  );


  buf

  (
    n3198_li,
    G50_p
  );


  buf

  (
    n3201_li,
    n3198_lo_p
  );


  buf

  (
    n3204_li,
    n3201_lo_p
  );


  buf

  (
    n3207_li,
    n3204_lo_p
  );


  buf

  (
    n3210_li,
    G51_p
  );


  buf

  (
    n3213_li,
    n3210_lo_p
  );


  buf

  (
    n3216_li,
    n3213_lo_p
  );


  buf

  (
    n3219_li,
    n3216_lo_p
  );


  buf

  (
    n3222_li,
    G52_p
  );


  buf

  (
    n3225_li,
    n3222_lo_p
  );


  buf

  (
    n3228_li,
    n3225_lo_p
  );


  buf

  (
    n3231_li,
    n3228_lo_p
  );


  buf

  (
    n3234_li,
    G53_p
  );


  buf

  (
    n3237_li,
    n3234_lo_p
  );


  buf

  (
    n3240_li,
    n3237_lo_p
  );


  buf

  (
    n3243_li,
    n3240_lo_p
  );


  buf

  (
    n3246_li,
    G54_p
  );


  buf

  (
    n3249_li,
    n3246_lo_p
  );


  buf

  (
    n3252_li,
    n3249_lo_p
  );


  buf

  (
    n3255_li,
    n3252_lo_p
  );


  buf

  (
    n3258_li,
    G55_p
  );


  buf

  (
    n3261_li,
    n3258_lo_p
  );


  buf

  (
    n3264_li,
    n3261_lo_p
  );


  buf

  (
    n3267_li,
    n3264_lo_p
  );


  buf

  (
    n3270_li,
    G56_p
  );


  buf

  (
    n3273_li,
    n3270_lo_p
  );


  buf

  (
    n3276_li,
    n3273_lo_p
  );


  buf

  (
    n3279_li,
    n3276_lo_p
  );


  buf

  (
    n3282_li,
    G57_p
  );


  buf

  (
    n3285_li,
    n3282_lo_p
  );


  buf

  (
    n3288_li,
    n3285_lo_p
  );


  buf

  (
    n3291_li,
    n3288_lo_p
  );


  buf

  (
    n3294_li,
    G58_p
  );


  buf

  (
    n3297_li,
    n3294_lo_p
  );


  buf

  (
    n3300_li,
    n3297_lo_p
  );


  buf

  (
    n3303_li,
    n3300_lo_p
  );


  buf

  (
    n3306_li,
    G59_p
  );


  buf

  (
    n3309_li,
    n3306_lo_p
  );


  buf

  (
    n3312_li,
    n3309_lo_p
  );


  buf

  (
    n3315_li,
    n3312_lo_p
  );


  buf

  (
    n3318_li,
    G60_p
  );


  buf

  (
    n3321_li,
    n3318_lo_p
  );


  buf

  (
    n3324_li,
    n3321_lo_p
  );


  buf

  (
    n3327_li,
    n3324_lo_p
  );


  buf

  (
    n3330_li,
    G61_p
  );


  buf

  (
    n3333_li,
    n3330_lo_p
  );


  buf

  (
    n3336_li,
    n3333_lo_p
  );


  buf

  (
    n3339_li,
    n3336_lo_p
  );


  buf

  (
    n3342_li,
    G62_p
  );


  buf

  (
    n3345_li,
    n3342_lo_p
  );


  buf

  (
    n3348_li,
    n3345_lo_p
  );


  buf

  (
    n3351_li,
    n3348_lo_p
  );


  buf

  (
    n3354_li,
    G63_p
  );


  buf

  (
    n3357_li,
    n3354_lo_p
  );


  buf

  (
    n3360_li,
    n3357_lo_p
  );


  buf

  (
    n3363_li,
    n3360_lo_p
  );


  buf

  (
    n3366_li,
    G64_p
  );


  buf

  (
    n3369_li,
    n3366_lo_p
  );


  buf

  (
    n3372_li,
    n3369_lo_p
  );


  buf

  (
    n3375_li,
    n3372_lo_p
  );


  buf

  (
    n3378_li,
    G65_p
  );


  buf

  (
    n3381_li,
    n3378_lo_p
  );


  buf

  (
    n3384_li,
    n3381_lo_p
  );


  buf

  (
    n3387_li,
    n3384_lo_p
  );


  buf

  (
    n3390_li,
    G66_p
  );


  buf

  (
    n3393_li,
    n3390_lo_p
  );


  buf

  (
    n3396_li,
    n3393_lo_p
  );


  buf

  (
    n3399_li,
    n3396_lo_p
  );


  buf

  (
    n3402_li,
    G67_p
  );


  buf

  (
    n3405_li,
    n3402_lo_p
  );


  buf

  (
    n3408_li,
    n3405_lo_p
  );


  buf

  (
    n3411_li,
    n3408_lo_p
  );


  buf

  (
    n3414_li,
    G68_p
  );


  buf

  (
    n3417_li,
    n3414_lo_p
  );


  buf

  (
    n3420_li,
    n3417_lo_p
  );


  buf

  (
    n3423_li,
    n3420_lo_p
  );


  buf

  (
    n3426_li,
    G69_p
  );


  buf

  (
    n3429_li,
    n3426_lo_p
  );


  buf

  (
    n3432_li,
    n3429_lo_p
  );


  buf

  (
    n3435_li,
    n3432_lo_p
  );


  buf

  (
    n3438_li,
    G70_p
  );


  buf

  (
    n3441_li,
    n3438_lo_p
  );


  buf

  (
    n3444_li,
    n3441_lo_p
  );


  buf

  (
    n3447_li,
    n3444_lo_p
  );


  buf

  (
    n3450_li,
    G71_p
  );


  buf

  (
    n3453_li,
    n3450_lo_p
  );


  buf

  (
    n3456_li,
    n3453_lo_p
  );


  buf

  (
    n3459_li,
    n3456_lo_p
  );


  buf

  (
    n3462_li,
    G72_p
  );


  buf

  (
    n3465_li,
    n3462_lo_p
  );


  buf

  (
    n3468_li,
    n3465_lo_p
  );


  buf

  (
    n3471_li,
    n3468_lo_p
  );


  buf

  (
    n3474_li,
    G73_p
  );


  buf

  (
    n3477_li,
    n3474_lo_p
  );


  buf

  (
    n3480_li,
    n3477_lo_p
  );


  buf

  (
    n3483_li,
    n3480_lo_p
  );


  buf

  (
    n3486_li,
    G74_p
  );


  buf

  (
    n3489_li,
    n3486_lo_p
  );


  buf

  (
    n3492_li,
    n3489_lo_p
  );


  buf

  (
    n3495_li,
    n3492_lo_p
  );


  buf

  (
    n3498_li,
    G75_p
  );


  buf

  (
    n3501_li,
    n3498_lo_p
  );


  buf

  (
    n3504_li,
    n3501_lo_p
  );


  buf

  (
    n3507_li,
    n3504_lo_p
  );


  buf

  (
    n3510_li,
    G76_p
  );


  buf

  (
    n3513_li,
    n3510_lo_p
  );


  buf

  (
    n3516_li,
    n3513_lo_p
  );


  buf

  (
    n3519_li,
    n3516_lo_p
  );


  buf

  (
    n3522_li,
    G77_p
  );


  buf

  (
    n3525_li,
    n3522_lo_p
  );


  buf

  (
    n3528_li,
    n3525_lo_p
  );


  buf

  (
    n3531_li,
    n3528_lo_p
  );


  buf

  (
    n3534_li,
    G78_p
  );


  buf

  (
    n3537_li,
    n3534_lo_p
  );


  buf

  (
    n3540_li,
    n3537_lo_p
  );


  buf

  (
    n3543_li,
    n3540_lo_p
  );


  buf

  (
    n3546_li,
    G79_p
  );


  buf

  (
    n3549_li,
    n3546_lo_p
  );


  buf

  (
    n3552_li,
    n3549_lo_p
  );


  buf

  (
    n3555_li,
    n3552_lo_p
  );


  buf

  (
    n3558_li,
    G80_p
  );


  buf

  (
    n3561_li,
    n3558_lo_p
  );


  buf

  (
    n3564_li,
    n3561_lo_p
  );


  buf

  (
    n3567_li,
    n3564_lo_p
  );


  buf

  (
    n3570_li,
    G81_p
  );


  buf

  (
    n3573_li,
    n3570_lo_p
  );


  buf

  (
    n3576_li,
    n3573_lo_p
  );


  buf

  (
    n3579_li,
    n3576_lo_p
  );


  buf

  (
    n3582_li,
    G82_p
  );


  buf

  (
    n3585_li,
    n3582_lo_p
  );


  buf

  (
    n3588_li,
    n3585_lo_p
  );


  buf

  (
    n3591_li,
    n3588_lo_p
  );


  buf

  (
    n3594_li,
    G83_p
  );


  buf

  (
    n3597_li,
    n3594_lo_p
  );


  buf

  (
    n3600_li,
    n3597_lo_p
  );


  buf

  (
    n3603_li,
    n3600_lo_p
  );


  buf

  (
    n3606_li,
    G84_p
  );


  buf

  (
    n3609_li,
    n3606_lo_p
  );


  buf

  (
    n3612_li,
    n3609_lo_p
  );


  buf

  (
    n3615_li,
    n3612_lo_p
  );


  buf

  (
    n3618_li,
    G85_p
  );


  buf

  (
    n3621_li,
    n3618_lo_p
  );


  buf

  (
    n3624_li,
    n3621_lo_p
  );


  buf

  (
    n3627_li,
    n3624_lo_p
  );


  buf

  (
    n3630_li,
    G86_p
  );


  buf

  (
    n3633_li,
    n3630_lo_p
  );


  buf

  (
    n3636_li,
    n3633_lo_p
  );


  buf

  (
    n3639_li,
    n3636_lo_p
  );


  buf

  (
    n3642_li,
    G87_p
  );


  buf

  (
    n3645_li,
    n3642_lo_p
  );


  buf

  (
    n3648_li,
    n3645_lo_p
  );


  buf

  (
    n3651_li,
    n3648_lo_p
  );


  buf

  (
    n3654_li,
    G88_p
  );


  buf

  (
    n3657_li,
    n3654_lo_p
  );


  buf

  (
    n3666_li,
    G89_p
  );


  buf

  (
    n3669_li,
    n3666_lo_p
  );


  buf

  (
    n3678_li,
    G90_p
  );


  buf

  (
    n3687_li,
    n7175_o2_p_spl_0
  );


  buf

  (
    n3690_li,
    G91_p
  );


  buf

  (
    n3702_li,
    G92_p
  );


  buf

  (
    n3711_li,
    n6945_o2_p_spl_0
  );


  buf

  (
    n3714_li,
    G93_p
  );


  buf

  (
    n3726_li,
    G94_p
  );


  buf

  (
    n3735_li,
    n6982_o2_p_spl_0
  );


  buf

  (
    n3738_li,
    G95_p
  );


  buf

  (
    n3750_li,
    G96_p
  );


  buf

  (
    n3753_li,
    n3750_lo_p
  );


  buf

  (
    n3759_li,
    n3756_lo_buf_o2_p_spl_
  );


  buf

  (
    n3762_li,
    G97_p
  );


  buf

  (
    n3765_li,
    n3762_lo_p
  );


  buf

  (
    n3774_li,
    G98_p
  );


  buf

  (
    n3777_li,
    n3774_lo_p
  );


  buf

  (
    n3786_li,
    G99_p
  );


  buf

  (
    n3789_li,
    n3786_lo_p
  );


  buf

  (
    n3792_li,
    n3789_lo_p
  );


  buf

  (
    n3795_li,
    n3792_lo_p
  );


  buf

  (
    n3798_li,
    G100_p
  );


  buf

  (
    n3801_li,
    n3798_lo_p
  );


  buf

  (
    n3810_li,
    G101_p
  );


  buf

  (
    n3813_li,
    n3810_lo_p
  );


  buf

  (
    n3822_li,
    G102_p
  );


  buf

  (
    n3825_li,
    n3822_lo_p
  );


  buf

  (
    n3834_li,
    G103_p
  );


  buf

  (
    n3843_li,
    n6947_o2_p_spl_
  );


  buf

  (
    n3846_li,
    G104_p
  );


  buf

  (
    n3867_li,
    n6621_o2_p_spl_
  );


  buf

  (
    n3891_li,
    n6623_o2_p_spl_
  );


  buf

  (
    n3915_li,
    n6669_o2_p_spl_1
  );


  buf

  (
    n3930_li,
    G111_p
  );


  buf

  (
    n3933_li,
    n3930_lo_p
  );


  buf

  (
    n3936_li,
    n3933_lo_p
  );


  buf

  (
    n3942_li,
    G112_p
  );


  buf

  (
    n3945_li,
    n3942_lo_p
  );


  buf

  (
    n3948_li,
    n3945_lo_p
  );


  buf

  (
    n3954_li,
    G113_p
  );


  buf

  (
    n3957_li,
    n3954_lo_p
  );


  buf

  (
    n3963_li,
    n3960_lo_buf_o2_p_spl_0
  );


  buf

  (
    n3966_li,
    G114_p
  );


  buf

  (
    n3969_li,
    n3966_lo_p
  );


  buf

  (
    n3975_li,
    n3972_lo_buf_o2_p
  );


  buf

  (
    n3978_li,
    G115_p
  );


  buf

  (
    n3987_li,
    n7453_o2_p_spl_0
  );


  buf

  (
    n3990_li,
    G116_p
  );


  buf

  (
    n4002_li,
    G117_p
  );


  buf

  (
    n4011_li,
    n6949_o2_p_spl_0
  );


  buf

  (
    n4014_li,
    G118_p
  );


  buf

  (
    n4026_li,
    G119_p
  );


  buf

  (
    n4035_li,
    n6984_o2_p_spl_0
  );


  buf

  (
    n4038_li,
    G120_p
  );


  buf

  (
    n4050_li,
    G121_p
  );


  buf

  (
    n4053_li,
    n4050_lo_p
  );


  buf

  (
    n4059_li,
    n4056_lo_buf_o2_p_spl_
  );


  buf

  (
    n4062_li,
    G122_p
  );


  buf

  (
    n4065_li,
    n4062_lo_p
  );


  buf

  (
    n4098_li,
    G125_p
  );


  buf

  (
    n4107_li,
    n6951_o2_p
  );


  buf

  (
    n4119_li,
    n6625_o2_p_spl_
  );


  buf

  (
    n4131_li,
    n6626_o2_p
  );


  buf

  (
    n4143_li,
    n6627_o2_p_spl_
  );


  buf

  (
    n4155_li,
    n6628_o2_p
  );


  buf

  (
    n4167_li,
    n6772_o2_p_spl_1
  );


  buf

  (
    n4179_li,
    n6773_o2_p
  );


  buf

  (
    n4182_li,
    G132_p
  );


  buf

  (
    n4185_li,
    n4182_lo_p
  );


  buf

  (
    n4188_li,
    n4185_lo_p
  );


  buf

  (
    n4194_li,
    G133_p
  );


  buf

  (
    n4197_li,
    n4194_lo_p
  );


  buf

  (
    n4200_li,
    n4197_lo_p
  );


  buf

  (
    n4206_li,
    G134_p
  );


  buf

  (
    n4209_li,
    n4206_lo_p
  );


  buf

  (
    n4212_li,
    n4209_lo_p
  );


  buf

  (
    n4215_li,
    n4212_lo_p
  );


  buf

  (
    n4227_li,
    n6774_o2_p_spl_1
  );


  buf

  (
    n4230_li,
    G136_p
  );


  buf

  (
    n4233_li,
    n4230_lo_p
  );


  buf

  (
    n4236_li,
    n4233_lo_p
  );


  buf

  (
    n4239_li,
    n4236_lo_p
  );


  buf

  (
    n4242_li,
    G137_p
  );


  buf

  (
    n4251_li,
    n7015_o2_p_spl_1
  );


  buf

  (
    n4263_li,
    n6682_o2_p_spl_1
  );


  buf

  (
    n4275_li,
    n6683_o2_p_spl_1
  );


  buf

  (
    n4278_li,
    G140_p
  );


  buf

  (
    n4287_li,
    n7132_o2_p_spl_1
  );


  buf

  (
    n4290_li,
    G141_p
  );


  buf

  (
    n4293_li,
    n4290_lo_p
  );


  buf

  (
    n4299_li,
    n4296_lo_buf_o2_p_spl_1
  );


  buf

  (
    n4302_li,
    G142_p
  );


  buf

  (
    n4305_li,
    n4302_lo_p
  );


  buf

  (
    n4311_li,
    n4308_lo_buf_o2_p_spl_1
  );


  buf

  (
    n4314_li,
    G143_p
  );


  buf

  (
    n4323_li,
    n7383_o2_p_spl_1
  );


  buf

  (
    n4326_li,
    G144_p
  );


  buf

  (
    n4335_li,
    n7016_o2_p_spl_1
  );


  buf

  (
    n4338_li,
    G145_p
  );


  buf

  (
    n4347_li,
    n7017_o2_p_spl_1
  );


  buf

  (
    n4350_li,
    G146_p
  );


  buf

  (
    n4359_li,
    n7133_o2_p_spl_1
  );


  buf

  (
    n4362_li,
    G147_p
  );


  buf

  (
    n4365_li,
    n4362_lo_p
  );


  buf

  (
    n4371_li,
    n4368_lo_buf_o2_p_spl_1
  );


  buf

  (
    n4374_li,
    G148_p
  );


  buf

  (
    n4383_li,
    n7018_o2_p_spl_1
  );


  buf

  (
    n4395_li,
    n6684_o2_p_spl_1
  );


  buf

  (
    n4407_li,
    n6685_o2_p_spl_1
  );


  buf

  (
    n4410_li,
    G151_p
  );


  buf

  (
    n4413_li,
    n4410_lo_p
  );


  buf

  (
    n4416_li,
    n4413_lo_p
  );


  buf

  (
    n4419_li,
    n4416_lo_p
  );


  buf

  (
    n4422_li,
    G152_p
  );


  buf

  (
    n4425_li,
    n4422_lo_p
  );


  buf

  (
    n4428_li,
    n4425_lo_p
  );


  buf

  (
    n4431_li,
    n4428_lo_p
  );


  buf

  (
    n4434_li,
    G153_p
  );


  buf

  (
    n4437_li,
    n4434_lo_p
  );


  buf

  (
    n4440_li,
    n4437_lo_p
  );


  buf

  (
    n4443_li,
    n4440_lo_p
  );


  buf

  (
    n4446_li,
    G154_p
  );


  buf

  (
    n4449_li,
    n4446_lo_p
  );


  buf

  (
    n4452_li,
    n4449_lo_p
  );


  buf

  (
    n4455_li,
    n4452_lo_p
  );


  buf

  (
    n4458_li,
    G155_p
  );


  buf

  (
    n4461_li,
    n4458_lo_p
  );


  buf

  (
    n4464_li,
    n4461_lo_p
  );


  buf

  (
    n4467_li,
    n4464_lo_p
  );


  buf

  (
    n4470_li,
    G156_p
  );


  buf

  (
    n4473_li,
    n4470_lo_p
  );


  buf

  (
    n4476_li,
    n4473_lo_p
  );


  buf

  (
    n4479_li,
    n4476_lo_p
  );


  buf

  (
    n4482_li,
    G157_p
  );


  buf

  (
    n4485_li,
    n4482_lo_p
  );


  buf

  (
    n4488_li,
    n4485_lo_p
  );


  buf

  (
    n4494_li,
    G158_p
  );


  buf

  (
    n4497_li,
    n4494_lo_p
  );


  buf

  (
    n4500_li,
    n4497_lo_p
  );


  buf

  (
    n4503_li,
    n4500_lo_p
  );


  buf

  (
    n4506_li,
    G159_p
  );


  buf

  (
    n4509_li,
    n4506_lo_p
  );


  buf

  (
    n4512_li,
    n4509_lo_p
  );


  buf

  (
    n4515_li,
    n4512_lo_p
  );


  buf

  (
    n4518_li,
    G160_p
  );


  buf

  (
    n4521_li,
    n4518_lo_p
  );


  buf

  (
    n4524_li,
    n4521_lo_p
  );


  buf

  (
    n4527_li,
    n4524_lo_p
  );


  buf

  (
    n4530_li,
    G161_p
  );


  buf

  (
    n4533_li,
    n4530_lo_p
  );


  buf

  (
    n4536_li,
    n4533_lo_p
  );


  buf

  (
    n4539_li,
    n4536_lo_p
  );


  buf

  (
    n4542_li,
    G162_p
  );


  buf

  (
    n4545_li,
    n4542_lo_p
  );


  buf

  (
    n4548_li,
    n4545_lo_p
  );


  buf

  (
    n4554_li,
    G163_p
  );


  buf

  (
    n4557_li,
    n4554_lo_p
  );


  buf

  (
    n4560_li,
    n4557_lo_p
  );


  buf

  (
    n4563_li,
    n4560_lo_p
  );


  buf

  (
    n4566_li,
    G164_p
  );


  buf

  (
    n4569_li,
    n4566_lo_p
  );


  buf

  (
    n4572_li,
    n4569_lo_p
  );


  buf

  (
    n4575_li,
    n4572_lo_p
  );


  buf

  (
    n4578_li,
    G165_p
  );


  buf

  (
    n4581_li,
    n4578_lo_p
  );


  buf

  (
    n4584_li,
    n4581_lo_p
  );


  buf

  (
    n4587_li,
    n4584_lo_p
  );


  buf

  (
    n4590_li,
    G166_p
  );


  buf

  (
    n4593_li,
    n4590_lo_p
  );


  buf

  (
    n4596_li,
    n4593_lo_p
  );


  buf

  (
    n4599_li,
    n4596_lo_p
  );


  buf

  (
    n4602_li,
    G167_p
  );


  buf

  (
    n4605_li,
    n4602_lo_p
  );


  buf

  (
    n4608_li,
    n4605_lo_p
  );


  buf

  (
    n4611_li,
    n4608_lo_p
  );


  buf

  (
    n4614_li,
    G168_p
  );


  buf

  (
    n4617_li,
    n4614_lo_p
  );


  buf

  (
    n4620_li,
    n4617_lo_p
  );


  buf

  (
    n4623_li,
    n4620_lo_p
  );


  buf

  (
    n4626_li,
    G169_p
  );


  buf

  (
    n4629_li,
    n4626_lo_p
  );


  buf

  (
    n4632_li,
    n4629_lo_p
  );


  buf

  (
    n4635_li,
    n4632_lo_p
  );


  buf

  (
    n4638_li,
    G170_p
  );


  buf

  (
    n4641_li,
    n4638_lo_p
  );


  buf

  (
    n4644_li,
    n4641_lo_p
  );


  buf

  (
    n4647_li,
    n4644_lo_p
  );


  buf

  (
    n4650_li,
    G171_p
  );


  buf

  (
    n4653_li,
    n4650_lo_p
  );


  buf

  (
    n4656_li,
    n4653_lo_p
  );


  buf

  (
    n4659_li,
    n4656_lo_p
  );


  buf

  (
    n4662_li,
    G172_p
  );


  buf

  (
    n4665_li,
    n4662_lo_p
  );


  buf

  (
    n4668_li,
    n4665_lo_p
  );


  buf

  (
    n4671_li,
    n4668_lo_p
  );


  buf

  (
    n4674_li,
    G173_p
  );


  buf

  (
    n4677_li,
    n4674_lo_p
  );


  buf

  (
    n4680_li,
    n4677_lo_p
  );


  buf

  (
    n4683_li,
    n4680_lo_p
  );


  buf

  (
    n4686_li,
    G174_p
  );


  buf

  (
    n4689_li,
    n4686_lo_p
  );


  buf

  (
    n4692_li,
    n4689_lo_p
  );


  buf

  (
    n4695_li,
    n4692_lo_p
  );


  buf

  (
    n4698_li,
    G175_p
  );


  buf

  (
    n4701_li,
    n4698_lo_p
  );


  buf

  (
    n4704_li,
    n4701_lo_p
  );


  buf

  (
    n4707_li,
    n4704_lo_p
  );


  buf

  (
    n4710_li,
    G176_p
  );


  buf

  (
    n4713_li,
    n4710_lo_p
  );


  buf

  (
    n4716_li,
    n4713_lo_p
  );


  buf

  (
    n4719_li,
    n4716_lo_p
  );


  buf

  (
    n4722_li,
    G177_p
  );


  buf

  (
    n4725_li,
    n4722_lo_p
  );


  buf

  (
    n4728_li,
    n4725_lo_p
  );


  buf

  (
    n4731_li,
    n4728_lo_p
  );


  buf

  (
    n4734_li,
    G178_p
  );


  buf

  (
    n4737_li,
    n4734_lo_p
  );


  buf

  (
    n4740_li,
    n4737_lo_p
  );


  buf

  (
    n4743_li,
    n4740_lo_p
  );


  buf

  (
    n6382_i2,
    n7355_o2_p
  );


  buf

  (
    n6383_i2,
    n7356_o2_p
  );


  buf

  (
    n6419_i2,
    n7388_o2_p
  );


  buf

  (
    n6420_i2,
    n7389_o2_p
  );


  buf

  (
    n6435_i2,
    n7432_o2_p
  );


  buf

  (
    n6436_i2,
    n7433_o2_p
  );


  buf

  (
    n6448_i2,
    n7485_o2_p
  );


  buf

  (
    n6449_i2,
    n7486_o2_p
  );


  buf

  (
    n6613_i2,
    G3474_o2_p_spl_
  );


  buf

  (
    n6614_i2,
    n2341_inv_p_spl_
  );


  buf

  (
    n6641_i2,
    G2711_o2_p
  );


  buf

  (
    n6658_i2,
    n2371_inv_p
  );


  buf

  (
    n6757_i2,
    G2404_o2_p_spl_1
  );


  buf

  (
    n6756_i2,
    G2466_o2_p_spl_1
  );


  buf

  (
    n7116_i2,
    G2430_o2_p_spl_
  );


  buf

  (
    n7156_i2,
    n2650_inv_p_spl_0
  );


  buf

  (
    n6549_i2,
    n2326_inv_p
  );


  buf

  (
    n6550_i2,
    n2329_inv_p
  );


  buf

  (
    n7357_i2,
    n2965_inv_p_spl_1
  );


  buf

  (
    n7358_i2,
    n2968_inv_p_spl_11
  );


  buf

  (
    n7359_i2,
    n2971_inv_p_spl_1
  );


  buf

  (
    n7360_i2,
    n2974_inv_p_spl_11
  );


  buf

  (
    n6621_i2,
    n7396_o2_p_spl_0
  );


  buf

  (
    n6623_i2,
    n7398_o2_p_spl_0
  );


  buf

  (
    n6625_i2,
    n7400_o2_p_spl_0
  );


  buf

  (
    n6626_i2,
    n7401_o2_p
  );


  buf

  (
    n6627_i2,
    n7402_o2_p_spl_0
  );


  buf

  (
    n6628_i2,
    n7403_o2_p
  );


  buf

  (
    n6629_i2,
    n7404_o2_p
  );


  buf

  (
    n6630_i2,
    n7405_o2_p
  );


  buf

  (
    n6669_i2,
    n7490_o2_p
  );


  buf

  (
    n7449_i2,
    n3118_inv_p_spl_11
  );


  buf

  (
    n7450_i2,
    n3121_inv_p_spl_11
  );


  buf

  (
    n7451_i2,
    n3124_inv_p_spl_11
  );


  buf

  (
    n7452_i2,
    n3127_inv_p_spl_11
  );


  buf

  (
    n6682_i2,
    n7527_o2_p
  );


  buf

  (
    n6683_i2,
    n7528_o2_p
  );


  buf

  (
    n6684_i2,
    n7529_o2_p
  );


  buf

  (
    n6685_i2,
    n7530_o2_p
  );


  buf

  (
    n7463_i2,
    G2492_o2_p_spl_01
  );


  buf

  (
    n6686_i2,
    n7523_o2_p
  );


  buf

  (
    n6687_i2,
    n7524_o2_p
  );


  buf

  (
    n6688_i2,
    n7525_o2_p
  );


  buf

  (
    n6689_i2,
    n7526_o2_p
  );


  buf

  (
    n6772_i2,
    n7534_o2_p
  );


  buf

  (
    n6773_i2,
    n7535_o2_p
  );


  buf

  (
    n6774_i2,
    n7536_o2_p
  );


  buf

  (
    n6775_i2,
    n7533_o2_p
  );


  buf

  (
    G3467_i2,
    g2452_n_spl_1
  );


  buf

  (
    G2810_i2,
    G2492_o2_p_spl_01
  );


  buf

  (
    n6833_i2,
    G2448_o2_p
  );


  buf

  (
    n6945_i2,
    n3708_lo_buf_o2_p_spl_
  );


  buf

  (
    n6947_i2,
    n3840_lo_buf_o2_p_spl_0
  );


  buf

  (
    n6949_i2,
    n4008_lo_buf_o2_p_spl_
  );


  buf

  (
    n6951_i2,
    n4104_lo_buf_o2_p
  );


  buf

  (
    n6888_i2,
    G2737_o2_p
  );


  buf

  (
    n6889_i2,
    G2850_o2_p
  );


  buf

  (
    n6936_i2,
    G2744_o2_p
  );


  buf

  (
    n6954_i2,
    G3517_o2_p
  );


  buf

  (
    n6955_i2,
    G3533_o2_p_spl_
  );


  buf

  (
    n6956_i2,
    G3629_o2_p
  );


  buf

  (
    n6957_i2,
    G3645_o2_p_spl_
  );


  buf

  (
    n6958_i2,
    n2497_inv_p
  );


  buf

  (
    n6982_i2,
    n3732_lo_buf_o2_p_spl_
  );


  buf

  (
    n6984_i2,
    n4032_lo_buf_o2_p_spl_
  );


  buf

  (
    n6974_i2,
    G2731_o2_p
  );


  buf

  (
    n6975_i2,
    G2844_o2_p
  );


  buf

  (
    n6999_i2,
    G3552_o2_p_spl_1
  );


  buf

  (
    n7015_i2,
    n4248_lo_buf_o2_p_spl_
  );


  buf

  (
    n7016_i2,
    n4332_lo_buf_o2_p
  );


  buf

  (
    n7017_i2,
    n4344_lo_buf_o2_p
  );


  buf

  (
    n7018_i2,
    n4380_lo_buf_o2_p
  );


  buf

  (
    n7005_i2,
    G2271_o2_p
  );


  buf

  (
    n7019_i2,
    G2398_o2_p
  );


  buf

  (
    n7022_i2,
    G2480_o2_p
  );


  buf

  (
    n7023_i2,
    G2418_o2_p
  );


  buf

  (
    n7132_i2,
    n4284_lo_buf_o2_p_spl_
  );


  buf

  (
    n7133_i2,
    n4356_lo_buf_o2_p_spl_
  );


  buf

  (
    n7135_i2,
    G2472_o2_p_spl_
  );


  buf

  (
    n7136_i2,
    G2410_o2_p_spl_
  );


  buf

  (
    n7175_i2,
    n3684_lo_buf_o2_p_spl_
  );


  buf

  (
    n7155_i2,
    n2647_inv_p_spl_1
  );


  buf

  (
    G3060_i2,
    g2462_n_spl_
  );


  buf

  (
    n7383_i2,
    n4320_lo_buf_o2_p_spl_
  );


  buf

  (
    G3802_i2,
    g2466_p_spl_
  );


  buf

  (
    G3859_i2,
    g2470_p_spl_
  );


  buf

  (
    n7355_i2,
    G2720_o2_p_spl_1
  );


  buf

  (
    n7356_i2,
    G2837_o2_p_spl_1
  );


  buf

  (
    G4054_i2,
    g2485_n_spl_
  );


  buf

  (
    G4068_i2,
    g2500_n_spl_
  );


  buf

  (
    n7384_i2,
    G2424_o2_p_spl_
  );


  buf

  (
    n7387_i2,
    G3503_o2_p
  );


  buf

  (
    n7388_i2,
    G3485_o2_p_spl_01
  );


  buf

  (
    n7389_i2,
    G3611_o2_p_spl_01
  );


  buf

  (
    n7386_i2,
    G3317_o2_p
  );


  buf

  (
    n7453_i2,
    n3984_lo_buf_o2_p
  );


  buf

  (
    n7431_i2,
    G2727_o2_p_spl_
  );


  buf

  (
    n7432_i2,
    G2715_o2_p_spl_
  );


  buf

  (
    n7433_i2,
    G2832_o2_p_spl_
  );


  buf

  (
    n7430_i2,
    G2543_o2_p_spl_
  );


  buf

  (
    n7485_i2,
    G3546_o2_p_spl_1
  );


  buf

  (
    n7486_i2,
    G3658_o2_p_spl_1
  );


  buf

  (
    G2508_i2,
    g2503_p_spl_
  );


  buf

  (
    G2486_i2,
    g2504_n_spl_10
  );


  buf

  (
    n7245_i2,
    n2662_inv_p_spl_
  );


  buf

  (
    n7246_i2,
    n2665_inv_p_spl_
  );


  buf

  (
    n3756_lo_buf_i2,
    n3753_lo_p_spl_0
  );


  buf

  (
    n4056_lo_buf_i2,
    n4053_lo_p_spl_0
  );


  buf

  (
    G3474_i2,
    g2507_n_spl_1
  );


  buf

  (
    G2817_i2,
    g2504_n_spl_10
  );


  buf

  (
    n7396_i2,
    n3864_lo_buf_o2_p
  );


  buf

  (
    n7398_i2,
    n3888_lo_buf_o2_p
  );


  buf

  (
    n7400_i2,
    n4116_lo_buf_o2_p
  );


  buf

  (
    n7401_i2,
    n4128_lo_buf_o2_p
  );


  buf

  (
    n7402_i2,
    n4140_lo_buf_o2_p
  );


  buf

  (
    n7403_i2,
    n4152_lo_buf_o2_p
  );


  buf

  (
    n7404_i2,
    G1815_o2_p_spl_
  );


  buf

  (
    n7405_i2,
    G1728_o2_p_spl_
  );


  buf

  (
    G2711_i2,
    g2508_p_spl_
  );


  buf

  (
    G2828_i2,
    g2504_n_spl_1
  );


  buf

  (
    n7490_i2,
    n3912_lo_buf_o2_p
  );


  buf

  (
    n7527_i2,
    n4260_lo_buf_o2_p_spl_
  );


  buf

  (
    n7528_i2,
    n4272_lo_buf_o2_p_spl_
  );


  buf

  (
    n7529_i2,
    n4392_lo_buf_o2_p_spl_
  );


  buf

  (
    n7530_i2,
    n4404_lo_buf_o2_p_spl_
  );


  buf

  (
    n7523_i2,
    G2460_o2_p_spl_
  );


  buf

  (
    n7524_i2,
    G2454_o2_p_spl_
  );


  buf

  (
    n7525_i2,
    G2392_o2_p_spl_
  );


  buf

  (
    n7526_i2,
    G2386_o2_p_spl_
  );


  buf

  (
    n4296_lo_buf_i2,
    n4293_lo_p_spl_1
  );


  buf

  (
    n4368_lo_buf_i2,
    n4365_lo_p_spl_1
  );


  buf

  (
    G2466_i2,
    g2511_n_spl_
  );


  buf

  (
    G2404_i2,
    g2514_n_spl_
  );


  buf

  (
    n7534_i2,
    n4164_lo_buf_o2_p_spl_
  );


  buf

  (
    n7535_i2,
    n4176_lo_buf_o2_p_spl_
  );


  buf

  (
    n7536_i2,
    n4224_lo_buf_o2_p_spl_1
  );


  buf

  (
    n7533_i2,
    G2379_o2_p_spl_1
  );


  buf

  (
    G1060_i2,
    n4080_lo_buf_o2_p_spl_10
  );


  buf

  (
    G963_i2,
    n4092_lo_buf_o2_p_spl_10
  );


  buf

  (
    G2448_i2,
    g2517_n_spl_10
  );


  buf

  (
    G2685_i2,
    g2518_p_spl_
  );


  buf

  (
    G2679_i2,
    g2519_p_spl_
  );


  not

  (
    G2774_i2,
    g2520_n_spl_
  );


  not

  (
    G2780_i2,
    g2521_n_spl_
  );


  buf

  (
    G2759_i2,
    G2486_o2_p_spl_01
  );


  buf

  (
    G2737_i2,
    g2522_p_spl_
  );


  buf

  (
    G2850_i2,
    g2523_p_spl_
  );


  buf

  (
    G3393_i2,
    g2526_n_spl_1
  );


  buf

  (
    G3404_i2,
    g2529_n_spl_1
  );


  buf

  (
    G3559_i2,
    g2532_n_spl_0
  );


  buf

  (
    G2744_i2,
    g2533_p_spl_1
  );


  buf

  (
    n3708_lo_buf_i2,
    n3702_lo_p_spl_
  );


  buf

  (
    n3840_lo_buf_i2,
    n3834_lo_p_spl_
  );


  buf

  (
    n4008_lo_buf_i2,
    n4002_lo_p_spl_
  );


  buf

  (
    n4104_lo_buf_i2,
    n4098_lo_p_spl_
  );


  buf

  (
    G1821_i2,
    n4080_lo_buf_o2_p_spl_1
  );


  buf

  (
    G1734_i2,
    n4092_lo_buf_o2_p_spl_1
  );


  buf

  (
    G3517_i2,
    g2536_n_spl_1
  );


  buf

  (
    G3533_i2,
    g2539_n_spl_1
  );


  buf

  (
    G3629_i2,
    g2542_n_spl_
  );


  buf

  (
    G3645_i2,
    g2545_n_spl_
  );


  buf

  (
    G2857_i2,
    g2517_n_spl_11
  );


  buf

  (
    G2731_i2,
    g2546_p_spl_
  );


  buf

  (
    G2844_i2,
    g2547_p_spl_
  );


  buf

  (
    n3732_lo_buf_i2,
    n3726_lo_p_spl_
  );


  buf

  (
    n4032_lo_buf_i2,
    n4026_lo_p_spl_
  );


  buf

  (
    G3552_i2,
    g2550_n_spl_
  );


  buf

  (
    G2271_i2,
    g2552_n_spl_
  );


  buf

  (
    n4248_lo_buf_i2,
    n4242_lo_p_spl_
  );


  buf

  (
    n4332_lo_buf_i2,
    n4326_lo_p_spl_
  );


  buf

  (
    n4344_lo_buf_i2,
    n4338_lo_p_spl_
  );


  buf

  (
    n4380_lo_buf_i2,
    n4374_lo_p_spl_
  );


  buf

  (
    G2398_i2,
    g2555_n_spl_
  );


  buf

  (
    G2480_i2,
    g2558_n_spl_
  );


  buf

  (
    G2418_i2,
    g2561_n_spl_
  );


  buf

  (
    G1455_i2,
    n7175_o2_p_spl_1
  );


  buf

  (
    G1449_i2,
    n6945_o2_p_spl_1
  );


  buf

  (
    G1452_i2,
    n6982_o2_p_spl_1
  );


  buf

  (
    G1425_i2,
    n3960_lo_buf_o2_p_spl_1
  );


  buf

  (
    G1428_i2,
    n7453_o2_p_spl_1
  );


  buf

  (
    G1419_i2,
    n6949_o2_p_spl_1
  );


  buf

  (
    G1422_i2,
    n6984_o2_p_spl_1
  );


  buf

  (
    n4308_lo_buf_i2,
    n4305_lo_p
  );


  buf

  (
    G2675_i2,
    g2562_p_spl_
  );


  buf

  (
    G3035_i2,
    n6688_o2_p_spl_1
  );


  buf

  (
    G3026_i2,
    n6689_o2_p_spl_1
  );


  buf

  (
    G3029_i2,
    n6775_o2_p_spl_1
  );


  buf

  (
    G3032_i2,
    n7019_o2_p_spl_1
  );


  buf

  (
    G2999_i2,
    n7022_o2_p_spl_1
  );


  buf

  (
    G3002_i2,
    n7135_o2_p_spl_1
  );


  buf

  (
    G2770_i2,
    G2486_o2_p_spl_10
  );


  buf

  (
    G3008_i2,
    G2486_o2_p_spl_10
  );


  buf

  (
    G2073_i2,
    n2650_inv_p_spl_0
  );


  buf

  (
    G2752_i2,
    G2492_o2_p_spl_10
  );


  buf

  (
    G3005_i2,
    G2492_o2_p_spl_10
  );


  buf

  (
    G5108_i2,
    g2592_p_spl_
  );


  buf

  (
    G5135_i2,
    g2611_n_spl_
  );


  buf

  (
    G5111_i2,
    g2641_n_spl_
  );


  buf

  (
    G5138_i2,
    g2660_n_spl_
  );


  buf

  (
    G3415_i2,
    g2663_n_spl_
  );


  buf

  (
    G3386_i2,
    g2666_n_spl_
  );


  buf

  (
    G3570_i2,
    g2669_n_spl_
  );


  buf

  (
    G2430_i2,
    g2672_n_spl_
  );


  buf

  (
    G3495_i2,
    g2675_n_spl_0
  );


  buf

  (
    G3621_i2,
    g2678_n_spl_0
  );


  buf

  (
    n4284_lo_buf_i2,
    n4278_lo_p_spl_
  );


  buf

  (
    n4356_lo_buf_i2,
    n4350_lo_p_spl_
  );


  buf

  (
    G2472_i2,
    g2681_n_spl_
  );


  buf

  (
    G2410_i2,
    g2684_n_spl_
  );


  buf

  (
    n3960_lo_buf_i2,
    n3957_lo_p_spl_
  );


  buf

  (
    n3972_lo_buf_i2,
    n3969_lo_p_spl_
  );


  buf

  (
    G2865_i2,
    g2517_n_spl_11
  );


  buf

  (
    G970_i2,
    n3657_lo_p_spl_00
  );


  buf

  (
    n3684_lo_buf_i2,
    n3678_lo_p_spl_
  );


  buf

  (
    n4080_lo_buf_i2,
    G123_p_spl_0
  );


  buf

  (
    n4092_lo_buf_i2,
    G124_p_spl_01
  );


  buf

  (
    G1053_i2,
    G123_p_spl_1
  );


  buf

  (
    G956_i2,
    G124_p_spl_1
  );


  buf

  (
    G1147_i2,
    n4056_lo_buf_o2_p_spl_
  );


  buf

  (
    G2705_i2,
    g2685_p
  );


  buf

  (
    G2693_i2,
    g2686_p
  );


  buf

  (
    G2696_i2,
    g2687_p
  );


  buf

  (
    G2700_i2,
    g2688_p
  );


  buf

  (
    G2915_i2,
    g2689_n
  );


  buf

  (
    G2966_i2,
    g2690_n
  );


  buf

  (
    G2540_i2,
    g2691_p
  );


  buf

  (
    G2788_i2,
    g2692_p
  );


  buf

  (
    G2792_i2,
    g2693_p
  );


  buf

  (
    G2797_i2,
    n6833_o2_p_spl_1
  );


  buf

  (
    G2804_i2,
    n6833_o2_p_spl_1
  );


  buf

  (
    G1038_i2,
    n7396_o2_p_spl_0
  );


  buf

  (
    G1044_i2,
    n7398_o2_p_spl_0
  );


  buf

  (
    G1090_i2,
    n7400_o2_p_spl_0
  );


  buf

  (
    G1096_i2,
    n7402_o2_p_spl_0
  );


  buf

  (
    G1029_i2,
    n3840_lo_buf_o2_p_spl_1
  );


  buf

  (
    G3942_i2,
    G3485_o2_p_spl_01
  );


  buf

  (
    G3954_i2,
    G3485_o2_p_spl_10
  );


  buf

  (
    G4011_i2,
    G3611_o2_p_spl_01
  );


  buf

  (
    G4017_i2,
    G3611_o2_p_spl_10
  );


  buf

  (
    G1141_i2,
    n3753_lo_p_spl_1
  );


  buf

  (
    G1081_i2,
    n4053_lo_p_spl_1
  );


  buf

  (
    G2146_i2,
    g2694_p
  );


  buf

  (
    G2145_i2,
    g2695_p
  );


  buf

  (
    G2144_i2,
    g2696_p
  );


  buf

  (
    G2143_i2,
    g2697_p
  );


  buf

  (
    G2142_i2,
    g2698_p
  );


  buf

  (
    G2141_i2,
    g2699_p
  );


  buf

  (
    G2140_i2,
    g2700_p
  );


  buf

  (
    G2139_i2,
    g2701_p
  );


  buf

  (
    G3769_i2,
    g2703_p_spl_
  );


  buf

  (
    G3773_i2,
    g2702_p_spl_
  );


  buf

  (
    G3768_i2,
    g2704_p_spl_
  );


  buf

  (
    G4101_i2,
    g2705_n
  );


  not

  (
    G3161_i2,
    g2706_n_spl_
  );


  not

  (
    G4143_i2,
    g2708_p
  );


  not

  (
    G3828_i2,
    g2709_n_spl_
  );


  not

  (
    G3831_i2,
    g2707_n_spl_
  );


  buf

  (
    G3334_i2,
    g2710_p
  );


  buf

  (
    G3335_i2,
    g2711_p
  );


  buf

  (
    G3180_i2,
    g2715_n
  );


  buf

  (
    G3340_i2,
    g2716_p
  );


  buf

  (
    G3339_i2,
    g2717_p
  );


  buf

  (
    G3341_i2,
    g2718_p
  );


  buf

  (
    G3234_i2,
    G2486_o2_p_spl_11
  );


  buf

  (
    G3829_i2,
    g2720_p
  );


  buf

  (
    G3338_i2,
    g2721_p
  );


  buf

  (
    G3336_i2,
    g2722_p
  );


  buf

  (
    G3770_i2,
    g2724_p
  );


  buf

  (
    G3918_i2,
    g2526_n_spl_1
  );


  buf

  (
    G3774_i2,
    g2723_p_spl_
  );


  buf

  (
    G3921_i2,
    g2529_n_spl_1
  );


  buf

  (
    G3832_i2,
    g2719_p_spl_
  );


  buf

  (
    G3993_i2,
    g2532_n_spl_
  );


  buf

  (
    G2076_i2,
    n7175_o2_p_spl_1
  );


  buf

  (
    G2071_i2,
    n6945_o2_p_spl_1
  );


  buf

  (
    G2072_i2,
    n6982_o2_p_spl_1
  );


  buf

  (
    G2069_i2,
    n3960_lo_buf_o2_p_spl_1
  );


  buf

  (
    G2070_i2,
    n7453_o2_p_spl_1
  );


  buf

  (
    G2067_i2,
    n6949_o2_p_spl_1
  );


  buf

  (
    G2068_i2,
    n6984_o2_p_spl_1
  );


  buf

  (
    G4095_i2,
    g2726_n
  );


  buf

  (
    G3272_i2,
    n6688_o2_p_spl_1
  );


  buf

  (
    G3269_i2,
    n6689_o2_p_spl_1
  );


  buf

  (
    G3270_i2,
    n6775_o2_p_spl_1
  );


  buf

  (
    G3271_i2,
    n7019_o2_p_spl_1
  );


  buf

  (
    G3265_i2,
    n7022_o2_p_spl_1
  );


  buf

  (
    G3266_i2,
    n7135_o2_p_spl_1
  );


  buf

  (
    G4137_i2,
    g2728_p
  );


  buf

  (
    G3268_i2,
    G2486_o2_p_spl_11
  );


  buf

  (
    G2361_i2,
    n2650_inv_p_spl_
  );


  buf

  (
    G3228_i2,
    G2492_o2_p_spl_11
  );


  buf

  (
    G3267_i2,
    G2492_o2_p_spl_11
  );


  buf

  (
    G2336_i2,
    g2731_n
  );


  buf

  (
    G3459_i2,
    g2734_n
  );


  buf

  (
    G3428_i2,
    g2737_n
  );


  buf

  (
    G3438_i2,
    g2740_n
  );


  buf

  (
    G3449_i2,
    g2743_n
  );


  buf

  (
    G3421_i2,
    g2746_n
  );


  buf

  (
    G3576_i2,
    g2749_n
  );


  buf

  (
    G3303_i2,
    g2752_n
  );


  buf

  (
    G3583_i2,
    g2755_n
  );


  buf

  (
    G3594_i2,
    g2758_n
  );


  buf

  (
    G3674_i2,
    g2761_n
  );


  buf

  (
    G3685_i2,
    g2767_p
  );


  buf

  (
    G4504_i2,
    g2806_p
  );


  buf

  (
    G4180_i2,
    g2841_p
  );


  buf

  (
    G5123_i2,
    g2592_p_spl_
  );


  buf

  (
    G5142_i2,
    g2611_n_spl_
  );


  buf

  (
    G5126_i2,
    g2641_n_spl_
  );


  buf

  (
    G5144_i2,
    g2660_n_spl_
  );


  buf

  (
    G3912_i2,
    g2666_n_spl_
  );


  buf

  (
    G4417_i2,
    g2900_p
  );


  buf

  (
    G4420_i2,
    g2946_n
  );


  buf

  (
    G3969_i2,
    g2675_n_spl_1
  );


  buf

  (
    G4023_i2,
    g2678_n_spl_1
  );


  buf

  (
    G2720_i2,
    g2947_p_spl_
  );


  buf

  (
    G2837_i2,
    g2948_p_spl_
  );


  buf

  (
    G836_i2,
    n3801_lo_p_spl_
  );


  buf

  (
    G848_i2,
    n3801_lo_p_spl_
  );


  buf

  (
    G813_i2,
    n3813_lo_p_spl_
  );


  buf

  (
    G825_i2,
    n3813_lo_p_spl_
  );


  buf

  (
    G1876_i2,
    n3657_lo_p_spl_0
  );


  buf

  (
    G4996_i2,
    g2962_p_spl_
  );


  buf

  (
    G4984_i2,
    g2976_p_spl_
  );


  buf

  (
    G4920_i2,
    g2995_n_spl_
  );


  buf

  (
    G4923_i2,
    g3004_n_spl_
  );


  buf

  (
    G4930_i2,
    g3023_p_spl_
  );


  buf

  (
    G4933_i2,
    g3032_p_spl_
  );


  buf

  (
    n4320_lo_buf_i2,
    n4314_lo_p_spl_0
  );


  buf

  (
    G2424_i2,
    g3035_n_spl_0
  );


  buf

  (
    G3317_i2,
    g3038_n
  );


  buf

  (
    G3503_i2,
    g3041_n_spl_1
  );


  buf

  (
    G3485_i2,
    g3044_n_spl_
  );


  buf

  (
    G3611_i2,
    g3047_n_spl_
  );


  buf

  (
    n3864_lo_buf_i2,
    G105_p_spl_
  );


  buf

  (
    n3888_lo_buf_i2,
    G107_p_spl_
  );


  buf

  (
    n4116_lo_buf_i2,
    G126_p_spl_
  );


  buf

  (
    n4128_lo_buf_i2,
    G127_p_spl_
  );


  buf

  (
    n4140_lo_buf_i2,
    G128_p_spl_
  );


  buf

  (
    n4152_lo_buf_i2,
    G129_p_spl_
  );


  buf

  (
    G1815_i2,
    G123_p_spl_1
  );


  buf

  (
    G1728_i2,
    G124_p_spl_1
  );


  buf

  (
    G1035_i2,
    n7396_o2_p_spl_1
  );


  buf

  (
    G1041_i2,
    n7398_o2_p_spl_1
  );


  buf

  (
    G1087_i2,
    n7400_o2_p_spl_1
  );


  buf

  (
    G1093_i2,
    n7402_o2_p_spl_1
  );


  buf

  (
    G1132_i2,
    n3708_lo_buf_o2_p_spl_
  );


  buf

  (
    G1108_i2,
    n4008_lo_buf_o2_p_spl_
  );


  buf

  (
    G1138_i2,
    n3732_lo_buf_o2_p_spl_
  );


  buf

  (
    G1114_i2,
    n4032_lo_buf_o2_p_spl_
  );


  buf

  (
    G1807_i2,
    g3049_p
  );


  buf

  (
    G2108_i2,
    g3051_p
  );


  buf

  (
    G1126_i2,
    n3684_lo_buf_o2_p_spl_
  );


  buf

  (
    G1899_i2,
    g3053_p
  );


  buf

  (
    G2134_i2,
    g3055_p
  );


  buf

  (
    G1852_i2,
    g3057_p
  );


  buf

  (
    G2116_i2,
    g3059_p
  );


  not

  (
    G2543_i2,
    g3060_n_spl_
  );


  buf

  (
    G2727_i2,
    g3061_p_spl_
  );


  buf

  (
    G2715_i2,
    g3062_p_spl_
  );


  buf

  (
    G2832_i2,
    g3063_p_spl_
  );


  buf

  (
    G1873_i2,
    n3657_lo_p_spl_1
  );


  buf

  (
    G3291_i2,
    g3064_p
  );


  buf

  (
    G5025_i2,
    g3074_p
  );


  buf

  (
    G5036_i2,
    g3084_p
  );


  not

  (
    G3132_i2,
    g3085_n
  );


  buf

  (
    G5038_i2,
    g3086_n
  );


  buf

  (
    G5039_i2,
    g3087_n
  );


  buf

  (
    G1150_i2,
    n3777_lo_p_spl_
  );


  buf

  (
    G1162_i2,
    n3777_lo_p_spl_
  );


  buf

  (
    G804_i2,
    n3825_lo_p_spl_
  );


  buf

  (
    G1172_i2,
    n3825_lo_p_spl_
  );


  buf

  (
    n3984_lo_buf_i2,
    n3978_lo_p_spl_
  );


  buf

  (
    G1802_i2,
    n7396_o2_p_spl_1
  );


  buf

  (
    G1804_i2,
    n7398_o2_p_spl_1
  );


  buf

  (
    G1849_i2,
    n7400_o2_p_spl_1
  );


  buf

  (
    G1851_i2,
    n7402_o2_p_spl_1
  );


  buf

  (
    G2492_i2,
    g3090_n
  );


  buf

  (
    G1799_i2,
    n3840_lo_buf_o2_p_spl_1
  );


  buf

  (
    G4231_i2,
    G3485_o2_p_spl_10
  );


  buf

  (
    G4234_i2,
    G3485_o2_p_spl_1
  );


  buf

  (
    G4245_i2,
    G3611_o2_p_spl_10
  );


  buf

  (
    G4247_i2,
    G3611_o2_p_spl_1
  );


  buf

  (
    G1894_i2,
    n3753_lo_p_spl_1
  );


  buf

  (
    G1846_i2,
    n4053_lo_p_spl_1
  );


  buf

  (
    G4238_i2,
    g2675_n_spl_1
  );


  buf

  (
    G4249_i2,
    g2678_n_spl_1
  );


  buf

  (
    G2293_i2,
    n3657_lo_p_spl_1
  );


  buf

  (
    G5022_i2,
    g2962_p_spl_
  );


  buf

  (
    G5006_i2,
    g2976_p_spl_
  );


  buf

  (
    G4944_i2,
    g2995_n_spl_
  );


  buf

  (
    G4946_i2,
    g3004_n_spl_
  );


  buf

  (
    G4954_i2,
    g3023_p_spl_
  );


  buf

  (
    G4956_i2,
    g3032_p_spl_
  );


  buf

  (
    G3546_i2,
    g3093_n_spl_
  );


  buf

  (
    G3658_i2,
    g3096_n_spl_
  );


  buf

  (
    G1344_i2,
    n4314_lo_p_spl_0
  );


  buf

  (
    G2921_i2,
    g3035_n_spl_0
  );


  buf

  (
    n3912_lo_buf_i2,
    G109_p_spl_
  );


  buf

  (
    G1835_i2,
    g3097_p
  );


  buf

  (
    G3810_i2,
    g3099_p_spl_
  );


  not

  (
    G3866_i2,
    g3101_n_spl_
  );


  buf

  (
    G3811_i2,
    g3104_p_spl_
  );


  buf

  (
    G2269_i2,
    g3105_p
  );


  buf

  (
    G3812_i2,
    g3108_p
  );


  not

  (
    G3867_i2,
    g3111_n_spl_
  );


  not

  (
    G3868_i2,
    g3114_n
  );


  buf

  (
    G3809_i2,
    g3115_p_spl_
  );


  not

  (
    G3716_i2,
    g3116_n_spl_
  );


  not

  (
    G4529_i2,
    g3124_n
  );


  buf

  (
    G4670_i2,
    g3137_p
  );


  buf

  (
    G4493_i2,
    g3138_p
  );


  buf

  (
    G4580_i2,
    g3139_n
  );


  buf

  (
    G3822_i2,
    g3140_p
  );


  buf

  (
    G3877_i2,
    g3141_p
  );


  buf

  (
    G4131_i2,
    g3144_n
  );


  not

  (
    G4170_i2,
    g3147_p
  );


  buf

  (
    G4051_i2,
    g3149_n
  );


  buf

  (
    G4065_i2,
    g3151_n
  );


  buf

  (
    G4697_i2,
    g3157_p
  );


  buf

  (
    G4706_i2,
    g3163_n
  );


  buf

  (
    G2460_i2,
    g3166_n_spl_
  );


  buf

  (
    G2454_i2,
    g3169_n_spl_
  );


  buf

  (
    G2392_i2,
    g3172_n_spl_
  );


  buf

  (
    G2386_i2,
    g3175_n_spl_
  );


  buf

  (
    n4260_lo_buf_i2,
    G138_p_spl_
  );


  buf

  (
    n4272_lo_buf_i2,
    G139_p_spl_
  );


  buf

  (
    n4392_lo_buf_i2,
    G149_p_spl_
  );


  buf

  (
    n4404_lo_buf_i2,
    G150_p_spl_
  );


  buf

  (
    G1512_i2,
    n4314_lo_p_spl_
  );


  buf

  (
    G3135_i2,
    g3035_n_spl_
  );


  buf

  (
    G2379_i2,
    g3178_n
  );


  buf

  (
    n4164_lo_buf_i2,
    G130_p
  );


  buf

  (
    n4176_lo_buf_i2,
    G131_p
  );


  buf

  (
    n4224_lo_buf_i2,
    G135_p
  );


  buf

  (
    G2975_i2,
    g3166_n_spl_
  );


  buf

  (
    G2978_i2,
    g3169_n_spl_
  );


  buf

  (
    G2933_i2,
    g3172_n_spl_
  );


  buf

  (
    G2936_i2,
    g3175_n_spl_
  );


  buf

  (
    G1356_i2,
    G138_p_spl_
  );


  buf

  (
    G1359_i2,
    G139_p_spl_
  );


  buf

  (
    G1398_i2,
    G149_p_spl_
  );


  buf

  (
    G1401_i2,
    G150_p_spl_
  );


  buf

  (
    n3399_lo_p_spl_,
    n3399_lo_p
  );


  buf

  (
    n2619_lo_p_spl_,
    n2619_lo_p
  );


  buf

  (
    n4587_lo_n_spl_,
    n4587_lo_n
  );


  buf

  (
    n2739_lo_n_spl_,
    n2739_lo_n
  );


  buf

  (
    n4455_lo_n_spl_,
    n4455_lo_n
  );


  buf

  (
    n4239_lo_n_spl_,
    n4239_lo_n
  );


  buf

  (
    g1198_n_spl_,
    g1198_n
  );


  buf

  (
    g1198_n_spl_0,
    g1198_n_spl_
  );


  buf

  (
    g1198_n_spl_00,
    g1198_n_spl_0
  );


  buf

  (
    g1198_n_spl_000,
    g1198_n_spl_00
  );


  buf

  (
    g1198_n_spl_001,
    g1198_n_spl_00
  );


  buf

  (
    g1198_n_spl_01,
    g1198_n_spl_0
  );


  buf

  (
    g1198_n_spl_010,
    g1198_n_spl_01
  );


  buf

  (
    g1198_n_spl_011,
    g1198_n_spl_01
  );


  buf

  (
    g1198_n_spl_1,
    g1198_n_spl_
  );


  buf

  (
    g1198_n_spl_10,
    g1198_n_spl_1
  );


  buf

  (
    g1198_n_spl_100,
    g1198_n_spl_10
  );


  buf

  (
    g1198_n_spl_11,
    g1198_n_spl_1
  );


  buf

  (
    n4563_lo_n_spl_,
    n4563_lo_n
  );


  buf

  (
    n4563_lo_n_spl_0,
    n4563_lo_n_spl_
  );


  buf

  (
    n4563_lo_n_spl_00,
    n4563_lo_n_spl_0
  );


  buf

  (
    n4563_lo_n_spl_01,
    n4563_lo_n_spl_0
  );


  buf

  (
    n4563_lo_n_spl_1,
    n4563_lo_n_spl_
  );


  buf

  (
    n4563_lo_n_spl_10,
    n4563_lo_n_spl_1
  );


  buf

  (
    n4563_lo_n_spl_11,
    n4563_lo_n_spl_1
  );


  buf

  (
    n4563_lo_p_spl_,
    n4563_lo_p
  );


  buf

  (
    n4563_lo_p_spl_0,
    n4563_lo_p_spl_
  );


  buf

  (
    n4563_lo_p_spl_00,
    n4563_lo_p_spl_0
  );


  buf

  (
    n4563_lo_p_spl_01,
    n4563_lo_p_spl_0
  );


  buf

  (
    n4563_lo_p_spl_1,
    n4563_lo_p_spl_
  );


  buf

  (
    n4563_lo_p_spl_10,
    n4563_lo_p_spl_1
  );


  buf

  (
    n4563_lo_p_spl_11,
    n4563_lo_p_spl_1
  );


  buf

  (
    n2991_lo_n_spl_,
    n2991_lo_n
  );


  buf

  (
    g1198_p_spl_,
    g1198_p
  );


  buf

  (
    g1216_n_spl_,
    g1216_n
  );


  buf

  (
    g1216_n_spl_0,
    g1216_n_spl_
  );


  buf

  (
    g1216_n_spl_1,
    g1216_n_spl_
  );


  buf

  (
    g1217_n_spl_,
    g1217_n
  );


  buf

  (
    g1217_n_spl_0,
    g1217_n_spl_
  );


  buf

  (
    g1217_n_spl_1,
    g1217_n_spl_
  );


  buf

  (
    n3399_lo_n_spl_,
    n3399_lo_n
  );


  buf

  (
    n3399_lo_n_spl_0,
    n3399_lo_n_spl_
  );


  buf

  (
    n3399_lo_n_spl_00,
    n3399_lo_n_spl_0
  );


  buf

  (
    n3399_lo_n_spl_1,
    n3399_lo_n_spl_
  );


  buf

  (
    n7357_o2_p_spl_,
    n7357_o2_p
  );


  buf

  (
    n7357_o2_p_spl_0,
    n7357_o2_p_spl_
  );


  buf

  (
    n4359_lo_n_spl_,
    n4359_lo_n
  );


  buf

  (
    n4035_lo_p_spl_,
    n4035_lo_p
  );


  buf

  (
    n7359_o2_p_spl_,
    n7359_o2_p
  );


  buf

  (
    n7359_o2_p_spl_0,
    n7359_o2_p_spl_
  );


  buf

  (
    n4035_lo_n_spl_,
    n4035_lo_n
  );


  buf

  (
    n7449_o2_n_spl_,
    n7449_o2_n
  );


  buf

  (
    n7449_o2_n_spl_0,
    n7449_o2_n_spl_
  );


  buf

  (
    n7452_o2_n_spl_,
    n7452_o2_n
  );


  buf

  (
    n7452_o2_n_spl_0,
    n7452_o2_n_spl_
  );


  buf

  (
    n4347_lo_n_spl_,
    n4347_lo_n
  );


  buf

  (
    n4011_lo_p_spl_,
    n4011_lo_p
  );


  buf

  (
    n4011_lo_n_spl_,
    n4011_lo_n
  );


  buf

  (
    n3963_lo_n_spl_,
    n3963_lo_n
  );


  buf

  (
    n3963_lo_n_spl_0,
    n3963_lo_n_spl_
  );


  buf

  (
    n3963_lo_p_spl_,
    n3963_lo_p
  );


  buf

  (
    g1265_p_spl_,
    g1265_p
  );


  buf

  (
    g1255_p_spl_,
    g1255_p
  );


  buf

  (
    g1268_p_spl_,
    g1268_p
  );


  buf

  (
    n4635_lo_p_spl_,
    n4635_lo_p
  );


  buf

  (
    n4635_lo_p_spl_0,
    n4635_lo_p_spl_
  );


  buf

  (
    n4635_lo_p_spl_00,
    n4635_lo_p_spl_0
  );


  buf

  (
    n4635_lo_p_spl_000,
    n4635_lo_p_spl_00
  );


  buf

  (
    n4635_lo_p_spl_001,
    n4635_lo_p_spl_00
  );


  buf

  (
    n4635_lo_p_spl_01,
    n4635_lo_p_spl_0
  );


  buf

  (
    n4635_lo_p_spl_010,
    n4635_lo_p_spl_01
  );


  buf

  (
    n4635_lo_p_spl_011,
    n4635_lo_p_spl_01
  );


  buf

  (
    n4635_lo_p_spl_1,
    n4635_lo_p_spl_
  );


  buf

  (
    n4635_lo_p_spl_10,
    n4635_lo_p_spl_1
  );


  buf

  (
    n4635_lo_p_spl_11,
    n4635_lo_p_spl_1
  );


  buf

  (
    n4407_lo_n_spl_,
    n4407_lo_n
  );


  buf

  (
    n4143_lo_p_spl_,
    n4143_lo_p
  );


  buf

  (
    n4623_lo_p_spl_,
    n4623_lo_p
  );


  buf

  (
    n4623_lo_p_spl_0,
    n4623_lo_p_spl_
  );


  buf

  (
    n4623_lo_p_spl_00,
    n4623_lo_p_spl_0
  );


  buf

  (
    n4623_lo_p_spl_000,
    n4623_lo_p_spl_00
  );


  buf

  (
    n4623_lo_p_spl_001,
    n4623_lo_p_spl_00
  );


  buf

  (
    n4623_lo_p_spl_01,
    n4623_lo_p_spl_0
  );


  buf

  (
    n4623_lo_p_spl_010,
    n4623_lo_p_spl_01
  );


  buf

  (
    n4623_lo_p_spl_1,
    n4623_lo_p_spl_
  );


  buf

  (
    n4623_lo_p_spl_10,
    n4623_lo_p_spl_1
  );


  buf

  (
    n4623_lo_p_spl_11,
    n4623_lo_p_spl_1
  );


  buf

  (
    n4143_lo_n_spl_,
    n4143_lo_n
  );


  buf

  (
    n4599_lo_n_spl_,
    n4599_lo_n
  );


  buf

  (
    n4599_lo_n_spl_0,
    n4599_lo_n_spl_
  );


  buf

  (
    n4599_lo_n_spl_00,
    n4599_lo_n_spl_0
  );


  buf

  (
    n4599_lo_n_spl_000,
    n4599_lo_n_spl_00
  );


  buf

  (
    n4599_lo_n_spl_001,
    n4599_lo_n_spl_00
  );


  buf

  (
    n4599_lo_n_spl_01,
    n4599_lo_n_spl_0
  );


  buf

  (
    n4599_lo_n_spl_010,
    n4599_lo_n_spl_01
  );


  buf

  (
    n4599_lo_n_spl_011,
    n4599_lo_n_spl_01
  );


  buf

  (
    n4599_lo_n_spl_1,
    n4599_lo_n_spl_
  );


  buf

  (
    n4599_lo_n_spl_10,
    n4599_lo_n_spl_1
  );


  buf

  (
    n4599_lo_n_spl_11,
    n4599_lo_n_spl_1
  );


  buf

  (
    n4611_lo_n_spl_,
    n4611_lo_n
  );


  buf

  (
    n4611_lo_n_spl_0,
    n4611_lo_n_spl_
  );


  buf

  (
    n4611_lo_n_spl_00,
    n4611_lo_n_spl_0
  );


  buf

  (
    n4611_lo_n_spl_000,
    n4611_lo_n_spl_00
  );


  buf

  (
    n4611_lo_n_spl_001,
    n4611_lo_n_spl_00
  );


  buf

  (
    n4611_lo_n_spl_01,
    n4611_lo_n_spl_0
  );


  buf

  (
    n4611_lo_n_spl_010,
    n4611_lo_n_spl_01
  );


  buf

  (
    n4611_lo_n_spl_1,
    n4611_lo_n_spl_
  );


  buf

  (
    n4611_lo_n_spl_10,
    n4611_lo_n_spl_1
  );


  buf

  (
    n4611_lo_n_spl_11,
    n4611_lo_n_spl_1
  );


  buf

  (
    n4395_lo_n_spl_,
    n4395_lo_n
  );


  buf

  (
    n4119_lo_p_spl_,
    n4119_lo_p
  );


  buf

  (
    n4119_lo_n_spl_,
    n4119_lo_n
  );


  buf

  (
    n4371_lo_n_spl_,
    n4371_lo_n
  );


  buf

  (
    n4371_lo_n_spl_0,
    n4371_lo_n_spl_
  );


  buf

  (
    n4059_lo_p_spl_,
    n4059_lo_p
  );


  buf

  (
    n4059_lo_n_spl_,
    n4059_lo_n
  );


  buf

  (
    n4371_lo_p_spl_,
    n4371_lo_p
  );


  buf

  (
    g1294_p_spl_,
    g1294_p
  );


  buf

  (
    g1284_p_spl_,
    g1284_p
  );


  buf

  (
    g1297_p_spl_,
    g1297_p
  );


  buf

  (
    g1307_p_spl_,
    g1307_p
  );


  buf

  (
    n4299_lo_n_spl_,
    n4299_lo_n
  );


  buf

  (
    n4299_lo_n_spl_0,
    n4299_lo_n_spl_
  );


  buf

  (
    n3759_lo_p_spl_,
    n3759_lo_p
  );


  buf

  (
    n3759_lo_n_spl_,
    n3759_lo_n
  );


  buf

  (
    n4299_lo_p_spl_,
    n4299_lo_p
  );


  buf

  (
    n4287_lo_n_spl_,
    n4287_lo_n
  );


  buf

  (
    n3735_lo_p_spl_,
    n3735_lo_p
  );


  buf

  (
    n3735_lo_n_spl_,
    n3735_lo_n
  );


  buf

  (
    n4335_lo_n_spl_,
    n4335_lo_n
  );


  buf

  (
    n3711_lo_p_spl_,
    n3711_lo_p
  );


  buf

  (
    n3711_lo_n_spl_,
    n3711_lo_n
  );


  buf

  (
    n4323_lo_n_spl_,
    n4323_lo_n
  );


  buf

  (
    n3687_lo_p_spl_,
    n3687_lo_p
  );


  buf

  (
    n3687_lo_n_spl_,
    n3687_lo_n
  );


  buf

  (
    g1332_p_spl_,
    g1332_p
  );


  buf

  (
    g1322_p_spl_,
    g1322_p
  );


  buf

  (
    g1342_p_spl_,
    g1342_p
  );


  buf

  (
    g1352_p_spl_,
    g1352_p
  );


  buf

  (
    n4227_lo_n_spl_,
    n4227_lo_n
  );


  buf

  (
    n3915_lo_p_spl_,
    n3915_lo_p
  );


  buf

  (
    n3915_lo_n_spl_,
    n3915_lo_n
  );


  buf

  (
    n4275_lo_n_spl_,
    n4275_lo_n
  );


  buf

  (
    n3891_lo_p_spl_,
    n3891_lo_p
  );


  buf

  (
    n3891_lo_n_spl_,
    n3891_lo_n
  );


  buf

  (
    n4263_lo_n_spl_,
    n4263_lo_n
  );


  buf

  (
    n3867_lo_p_spl_,
    n3867_lo_p
  );


  buf

  (
    n3867_lo_n_spl_,
    n3867_lo_n
  );


  buf

  (
    n4251_lo_n_spl_,
    n4251_lo_n
  );


  buf

  (
    n3843_lo_p_spl_,
    n3843_lo_p
  );


  buf

  (
    n3843_lo_n_spl_,
    n3843_lo_n
  );


  buf

  (
    g1375_p_spl_,
    g1375_p
  );


  buf

  (
    g1365_p_spl_,
    g1365_p
  );


  buf

  (
    g1385_p_spl_,
    g1385_p
  );


  buf

  (
    g1395_p_spl_,
    g1395_p
  );


  buf

  (
    n6419_o2_n_spl_,
    n6419_o2_n
  );


  buf

  (
    n6613_o2_n_spl_,
    n6613_o2_n
  );


  buf

  (
    n6613_o2_n_spl_0,
    n6613_o2_n_spl_
  );


  buf

  (
    G3467_o2_n_spl_,
    G3467_o2_n
  );


  buf

  (
    G3467_o2_n_spl_0,
    G3467_o2_n_spl_
  );


  buf

  (
    G3467_o2_n_spl_1,
    G3467_o2_n_spl_
  );


  buf

  (
    g1403_n_spl_,
    g1403_n
  );


  buf

  (
    G3570_o2_n_spl_,
    G3570_o2_n
  );


  buf

  (
    G2759_o2_p_spl_,
    G2759_o2_p
  );


  buf

  (
    G2759_o2_p_spl_0,
    G2759_o2_p_spl_
  );


  buf

  (
    G2759_o2_p_spl_1,
    G2759_o2_p_spl_
  );


  buf

  (
    G3559_o2_n_spl_,
    G3559_o2_n
  );


  buf

  (
    G3559_o2_n_spl_0,
    G3559_o2_n_spl_
  );


  buf

  (
    G2752_o2_p_spl_,
    G2752_o2_p
  );


  buf

  (
    G2752_o2_p_spl_0,
    G2752_o2_p_spl_
  );


  buf

  (
    G2752_o2_p_spl_00,
    G2752_o2_p_spl_0
  );


  buf

  (
    G2752_o2_p_spl_01,
    G2752_o2_p_spl_0
  );


  buf

  (
    G2752_o2_p_spl_1,
    G2752_o2_p_spl_
  );


  buf

  (
    G3303_o2_p_spl_,
    G3303_o2_p
  );


  buf

  (
    G3303_o2_p_spl_0,
    G3303_o2_p_spl_
  );


  buf

  (
    G3303_o2_p_spl_00,
    G3303_o2_p_spl_0
  );


  buf

  (
    G3303_o2_p_spl_000,
    G3303_o2_p_spl_00
  );


  buf

  (
    G3303_o2_p_spl_01,
    G3303_o2_p_spl_0
  );


  buf

  (
    G3303_o2_p_spl_1,
    G3303_o2_p_spl_
  );


  buf

  (
    G3303_o2_p_spl_10,
    G3303_o2_p_spl_1
  );


  buf

  (
    G3303_o2_p_spl_11,
    G3303_o2_p_spl_1
  );


  buf

  (
    G2797_o2_n_spl_,
    G2797_o2_n
  );


  buf

  (
    G2797_o2_n_spl_0,
    G2797_o2_n_spl_
  );


  buf

  (
    G3303_o2_n_spl_,
    G3303_o2_n
  );


  buf

  (
    G3303_o2_n_spl_0,
    G3303_o2_n_spl_
  );


  buf

  (
    G3303_o2_n_spl_00,
    G3303_o2_n_spl_0
  );


  buf

  (
    G3303_o2_n_spl_000,
    G3303_o2_n_spl_00
  );


  buf

  (
    G3303_o2_n_spl_01,
    G3303_o2_n_spl_0
  );


  buf

  (
    G3303_o2_n_spl_1,
    G3303_o2_n_spl_
  );


  buf

  (
    G3303_o2_n_spl_10,
    G3303_o2_n_spl_1
  );


  buf

  (
    G3303_o2_n_spl_11,
    G3303_o2_n_spl_1
  );


  buf

  (
    G2797_o2_p_spl_,
    G2797_o2_p
  );


  buf

  (
    G2797_o2_p_spl_0,
    G2797_o2_p_spl_
  );


  buf

  (
    G3583_o2_p_spl_,
    G3583_o2_p
  );


  buf

  (
    G3583_o2_p_spl_0,
    G3583_o2_p_spl_
  );


  buf

  (
    G3583_o2_p_spl_00,
    G3583_o2_p_spl_0
  );


  buf

  (
    G3583_o2_p_spl_01,
    G3583_o2_p_spl_0
  );


  buf

  (
    G3583_o2_p_spl_1,
    G3583_o2_p_spl_
  );


  buf

  (
    G3583_o2_n_spl_,
    G3583_o2_n
  );


  buf

  (
    G3583_o2_n_spl_0,
    G3583_o2_n_spl_
  );


  buf

  (
    G3583_o2_n_spl_00,
    G3583_o2_n_spl_0
  );


  buf

  (
    G3583_o2_n_spl_01,
    G3583_o2_n_spl_0
  );


  buf

  (
    G3583_o2_n_spl_1,
    G3583_o2_n_spl_
  );


  buf

  (
    G3576_o2_p_spl_,
    G3576_o2_p
  );


  buf

  (
    G3576_o2_p_spl_0,
    G3576_o2_p_spl_
  );


  buf

  (
    G3576_o2_p_spl_00,
    G3576_o2_p_spl_0
  );


  buf

  (
    G3576_o2_p_spl_01,
    G3576_o2_p_spl_0
  );


  buf

  (
    G3576_o2_p_spl_1,
    G3576_o2_p_spl_
  );


  buf

  (
    G3576_o2_n_spl_,
    G3576_o2_n
  );


  buf

  (
    G3576_o2_n_spl_0,
    G3576_o2_n_spl_
  );


  buf

  (
    G3576_o2_n_spl_00,
    G3576_o2_n_spl_0
  );


  buf

  (
    G3576_o2_n_spl_01,
    G3576_o2_n_spl_0
  );


  buf

  (
    G3576_o2_n_spl_1,
    G3576_o2_n_spl_
  );


  buf

  (
    G3594_o2_p_spl_,
    G3594_o2_p
  );


  buf

  (
    G3594_o2_p_spl_0,
    G3594_o2_p_spl_
  );


  buf

  (
    G3594_o2_p_spl_00,
    G3594_o2_p_spl_0
  );


  buf

  (
    G3594_o2_p_spl_01,
    G3594_o2_p_spl_0
  );


  buf

  (
    G3594_o2_p_spl_1,
    G3594_o2_p_spl_
  );


  buf

  (
    G3594_o2_n_spl_,
    G3594_o2_n
  );


  buf

  (
    G3594_o2_n_spl_0,
    G3594_o2_n_spl_
  );


  buf

  (
    G3594_o2_n_spl_00,
    G3594_o2_n_spl_0
  );


  buf

  (
    G3594_o2_n_spl_01,
    G3594_o2_n_spl_0
  );


  buf

  (
    G3594_o2_n_spl_1,
    G3594_o2_n_spl_
  );


  buf

  (
    g1411_n_spl_,
    g1411_n
  );


  buf

  (
    g1407_n_spl_,
    g1407_n
  );


  buf

  (
    n6420_o2_n_spl_,
    n6420_o2_n
  );


  buf

  (
    n6614_o2_p_spl_,
    n6614_o2_p
  );


  buf

  (
    n6614_o2_p_spl_0,
    n6614_o2_p_spl_
  );


  buf

  (
    G2810_o2_p_spl_,
    G2810_o2_p
  );


  buf

  (
    G2810_o2_p_spl_0,
    G2810_o2_p_spl_
  );


  buf

  (
    G2810_o2_p_spl_1,
    G2810_o2_p_spl_
  );


  buf

  (
    g1415_n_spl_,
    g1415_n
  );


  buf

  (
    G3415_o2_n_spl_,
    G3415_o2_n
  );


  buf

  (
    G3393_o2_n_spl_,
    G3393_o2_n
  );


  buf

  (
    G3393_o2_n_spl_0,
    G3393_o2_n_spl_
  );


  buf

  (
    G3393_o2_n_spl_1,
    G3393_o2_n_spl_
  );


  buf

  (
    G3404_o2_n_spl_,
    G3404_o2_n
  );


  buf

  (
    G3404_o2_n_spl_0,
    G3404_o2_n_spl_
  );


  buf

  (
    G3386_o2_n_spl_,
    G3386_o2_n
  );


  buf

  (
    G3386_o2_n_spl_0,
    G3386_o2_n_spl_
  );


  buf

  (
    G3386_o2_n_spl_00,
    G3386_o2_n_spl_0
  );


  buf

  (
    G3386_o2_n_spl_1,
    G3386_o2_n_spl_
  );


  buf

  (
    G3428_o2_p_spl_,
    G3428_o2_p
  );


  buf

  (
    G3428_o2_p_spl_0,
    G3428_o2_p_spl_
  );


  buf

  (
    G3428_o2_p_spl_00,
    G3428_o2_p_spl_0
  );


  buf

  (
    G3428_o2_p_spl_000,
    G3428_o2_p_spl_00
  );


  buf

  (
    G3428_o2_p_spl_01,
    G3428_o2_p_spl_0
  );


  buf

  (
    G3428_o2_p_spl_1,
    G3428_o2_p_spl_
  );


  buf

  (
    G3428_o2_p_spl_10,
    G3428_o2_p_spl_1
  );


  buf

  (
    G3428_o2_p_spl_11,
    G3428_o2_p_spl_1
  );


  buf

  (
    G3459_o2_p_spl_,
    G3459_o2_p
  );


  buf

  (
    G3459_o2_p_spl_0,
    G3459_o2_p_spl_
  );


  buf

  (
    G3428_o2_n_spl_,
    G3428_o2_n
  );


  buf

  (
    G3428_o2_n_spl_0,
    G3428_o2_n_spl_
  );


  buf

  (
    G3428_o2_n_spl_00,
    G3428_o2_n_spl_0
  );


  buf

  (
    G3428_o2_n_spl_000,
    G3428_o2_n_spl_00
  );


  buf

  (
    G3428_o2_n_spl_01,
    G3428_o2_n_spl_0
  );


  buf

  (
    G3428_o2_n_spl_1,
    G3428_o2_n_spl_
  );


  buf

  (
    G3428_o2_n_spl_10,
    G3428_o2_n_spl_1
  );


  buf

  (
    G3428_o2_n_spl_11,
    G3428_o2_n_spl_1
  );


  buf

  (
    G3459_o2_n_spl_,
    G3459_o2_n
  );


  buf

  (
    G3459_o2_n_spl_0,
    G3459_o2_n_spl_
  );


  buf

  (
    G3438_o2_p_spl_,
    G3438_o2_p
  );


  buf

  (
    G3438_o2_p_spl_0,
    G3438_o2_p_spl_
  );


  buf

  (
    G3438_o2_p_spl_00,
    G3438_o2_p_spl_0
  );


  buf

  (
    G3438_o2_p_spl_01,
    G3438_o2_p_spl_0
  );


  buf

  (
    G3438_o2_p_spl_1,
    G3438_o2_p_spl_
  );


  buf

  (
    G3438_o2_n_spl_,
    G3438_o2_n
  );


  buf

  (
    G3438_o2_n_spl_0,
    G3438_o2_n_spl_
  );


  buf

  (
    G3438_o2_n_spl_00,
    G3438_o2_n_spl_0
  );


  buf

  (
    G3438_o2_n_spl_01,
    G3438_o2_n_spl_0
  );


  buf

  (
    G3438_o2_n_spl_1,
    G3438_o2_n_spl_
  );


  buf

  (
    G3421_o2_p_spl_,
    G3421_o2_p
  );


  buf

  (
    G3421_o2_p_spl_0,
    G3421_o2_p_spl_
  );


  buf

  (
    G3421_o2_p_spl_00,
    G3421_o2_p_spl_0
  );


  buf

  (
    G3421_o2_p_spl_01,
    G3421_o2_p_spl_0
  );


  buf

  (
    G3421_o2_p_spl_1,
    G3421_o2_p_spl_
  );


  buf

  (
    G3421_o2_n_spl_,
    G3421_o2_n
  );


  buf

  (
    G3421_o2_n_spl_0,
    G3421_o2_n_spl_
  );


  buf

  (
    G3421_o2_n_spl_00,
    G3421_o2_n_spl_0
  );


  buf

  (
    G3421_o2_n_spl_01,
    G3421_o2_n_spl_0
  );


  buf

  (
    G3421_o2_n_spl_1,
    G3421_o2_n_spl_
  );


  buf

  (
    G3449_o2_p_spl_,
    G3449_o2_p
  );


  buf

  (
    G3449_o2_p_spl_0,
    G3449_o2_p_spl_
  );


  buf

  (
    G3449_o2_p_spl_00,
    G3449_o2_p_spl_0
  );


  buf

  (
    G3449_o2_p_spl_01,
    G3449_o2_p_spl_0
  );


  buf

  (
    G3449_o2_p_spl_1,
    G3449_o2_p_spl_
  );


  buf

  (
    G3449_o2_n_spl_,
    G3449_o2_n
  );


  buf

  (
    G3449_o2_n_spl_0,
    G3449_o2_n_spl_
  );


  buf

  (
    G3449_o2_n_spl_00,
    G3449_o2_n_spl_0
  );


  buf

  (
    G3449_o2_n_spl_01,
    G3449_o2_n_spl_0
  );


  buf

  (
    G3449_o2_n_spl_1,
    G3449_o2_n_spl_
  );


  buf

  (
    g1423_n_spl_,
    g1423_n
  );


  buf

  (
    g1419_n_spl_,
    g1419_n
  );


  buf

  (
    g1430_p_spl_,
    g1430_p
  );


  buf

  (
    g1427_n_spl_,
    g1427_n
  );


  buf

  (
    g1430_n_spl_,
    g1430_n
  );


  buf

  (
    g1427_p_spl_,
    g1427_p
  );


  buf

  (
    g1435_p_spl_,
    g1435_p
  );


  buf

  (
    g1435_p_spl_0,
    g1435_p_spl_
  );


  buf

  (
    g1435_p_spl_1,
    g1435_p_spl_
  );


  buf

  (
    g1434_n_spl_,
    g1434_n
  );


  buf

  (
    g1434_n_spl_0,
    g1434_n_spl_
  );


  buf

  (
    g1434_n_spl_1,
    g1434_n_spl_
  );


  buf

  (
    g1435_n_spl_,
    g1435_n
  );


  buf

  (
    g1435_n_spl_0,
    g1435_n_spl_
  );


  buf

  (
    g1435_n_spl_1,
    g1435_n_spl_
  );


  buf

  (
    g1434_p_spl_,
    g1434_p
  );


  buf

  (
    g1434_p_spl_0,
    g1434_p_spl_
  );


  buf

  (
    g1434_p_spl_1,
    g1434_p_spl_
  );


  buf

  (
    G1147_o2_n_spl_,
    G1147_o2_n
  );


  buf

  (
    G1147_o2_n_spl_0,
    G1147_o2_n_spl_
  );


  buf

  (
    G1147_o2_n_spl_1,
    G1147_o2_n_spl_
  );


  buf

  (
    G1147_o2_p_spl_,
    G1147_o2_p
  );


  buf

  (
    G1147_o2_p_spl_0,
    G1147_o2_p_spl_
  );


  buf

  (
    G1147_o2_p_spl_1,
    G1147_o2_p_spl_
  );


  buf

  (
    g1455_p_spl_,
    g1455_p
  );


  buf

  (
    g1452_n_spl_,
    g1452_n
  );


  buf

  (
    g1455_n_spl_,
    g1455_n
  );


  buf

  (
    g1452_p_spl_,
    g1452_p
  );


  buf

  (
    g1460_p_spl_,
    g1460_p
  );


  buf

  (
    g1460_p_spl_0,
    g1460_p_spl_
  );


  buf

  (
    g1460_p_spl_1,
    g1460_p_spl_
  );


  buf

  (
    g1459_n_spl_,
    g1459_n
  );


  buf

  (
    g1459_n_spl_0,
    g1459_n_spl_
  );


  buf

  (
    g1459_n_spl_1,
    g1459_n_spl_
  );


  buf

  (
    g1460_n_spl_,
    g1460_n
  );


  buf

  (
    g1460_n_spl_0,
    g1460_n_spl_
  );


  buf

  (
    g1460_n_spl_1,
    g1460_n_spl_
  );


  buf

  (
    g1459_p_spl_,
    g1459_p
  );


  buf

  (
    g1459_p_spl_0,
    g1459_p_spl_
  );


  buf

  (
    g1459_p_spl_1,
    g1459_p_spl_
  );


  buf

  (
    G2336_o2_p_spl_,
    G2336_o2_p
  );


  buf

  (
    G2336_o2_p_spl_0,
    G2336_o2_p_spl_
  );


  buf

  (
    G2336_o2_p_spl_1,
    G2336_o2_p_spl_
  );


  buf

  (
    G2336_o2_n_spl_,
    G2336_o2_n
  );


  buf

  (
    G2336_o2_n_spl_0,
    G2336_o2_n_spl_
  );


  buf

  (
    G2336_o2_n_spl_1,
    G2336_o2_n_spl_
  );


  buf

  (
    n4311_lo_n_spl_,
    n4311_lo_n
  );


  buf

  (
    n4311_lo_n_spl_0,
    n4311_lo_n_spl_
  );


  buf

  (
    g1475_n_spl_,
    g1475_n
  );


  buf

  (
    G2770_o2_p_spl_,
    G2770_o2_p
  );


  buf

  (
    G2774_o2_n_spl_,
    G2774_o2_n
  );


  buf

  (
    G2780_o2_n_spl_,
    G2780_o2_n
  );


  buf

  (
    n7463_o2_n_spl_,
    n7463_o2_n
  );


  buf

  (
    n7463_o2_n_spl_0,
    n7463_o2_n_spl_
  );


  buf

  (
    n7463_o2_n_spl_1,
    n7463_o2_n_spl_
  );


  buf

  (
    G2540_o2_p_spl_,
    G2540_o2_p
  );


  buf

  (
    G2540_o2_n_spl_,
    G2540_o2_n
  );


  buf

  (
    G2788_o2_p_spl_,
    G2788_o2_p
  );


  buf

  (
    G2788_o2_p_spl_0,
    G2788_o2_p_spl_
  );


  buf

  (
    G2788_o2_n_spl_,
    G2788_o2_n
  );


  buf

  (
    G2788_o2_n_spl_0,
    G2788_o2_n_spl_
  );


  buf

  (
    G2792_o2_p_spl_,
    G2792_o2_p
  );


  buf

  (
    G2792_o2_p_spl_0,
    G2792_o2_p_spl_
  );


  buf

  (
    G2792_o2_n_spl_,
    G2792_o2_n
  );


  buf

  (
    G2792_o2_n_spl_0,
    G2792_o2_n_spl_
  );


  buf

  (
    g1503_p_spl_,
    g1503_p
  );


  buf

  (
    g1503_n_spl_,
    g1503_n
  );


  buf

  (
    G2804_o2_n_spl_,
    G2804_o2_n
  );


  buf

  (
    G2804_o2_n_spl_0,
    G2804_o2_n_spl_
  );


  buf

  (
    G2804_o2_n_spl_1,
    G2804_o2_n_spl_
  );


  buf

  (
    G2804_o2_p_spl_,
    G2804_o2_p
  );


  buf

  (
    G2804_o2_p_spl_0,
    G2804_o2_p_spl_
  );


  buf

  (
    G2804_o2_p_spl_1,
    G2804_o2_p_spl_
  );


  buf

  (
    g1510_p_spl_,
    g1510_p
  );


  buf

  (
    G2675_o2_n_spl_,
    G2675_o2_n
  );


  buf

  (
    G2679_o2_n_spl_,
    G2679_o2_n
  );


  buf

  (
    G2685_o2_n_spl_,
    G2685_o2_n
  );


  buf

  (
    G2693_o2_p_spl_,
    G2693_o2_p
  );


  buf

  (
    G2693_o2_n_spl_,
    G2693_o2_n
  );


  buf

  (
    G2696_o2_p_spl_,
    G2696_o2_p
  );


  buf

  (
    G2696_o2_p_spl_0,
    G2696_o2_p_spl_
  );


  buf

  (
    G2696_o2_n_spl_,
    G2696_o2_n
  );


  buf

  (
    G2696_o2_n_spl_0,
    G2696_o2_n_spl_
  );


  buf

  (
    G2700_o2_p_spl_,
    G2700_o2_p
  );


  buf

  (
    G2700_o2_p_spl_0,
    G2700_o2_p_spl_
  );


  buf

  (
    G2700_o2_n_spl_,
    G2700_o2_n
  );


  buf

  (
    G2700_o2_n_spl_0,
    G2700_o2_n_spl_
  );


  buf

  (
    g1529_p_spl_,
    g1529_p
  );


  buf

  (
    g1529_n_spl_,
    g1529_n
  );


  buf

  (
    G2705_o2_p_spl_,
    G2705_o2_p
  );


  buf

  (
    G2705_o2_p_spl_0,
    G2705_o2_p_spl_
  );


  buf

  (
    G2705_o2_p_spl_1,
    G2705_o2_p_spl_
  );


  buf

  (
    G2705_o2_n_spl_,
    G2705_o2_n
  );


  buf

  (
    G2705_o2_n_spl_0,
    G2705_o2_n_spl_
  );


  buf

  (
    G2705_o2_n_spl_1,
    G2705_o2_n_spl_
  );


  buf

  (
    g1536_p_spl_,
    g1536_p
  );


  buf

  (
    n7358_o2_p_spl_,
    n7358_o2_p
  );


  buf

  (
    n7360_o2_p_spl_,
    n7360_o2_p
  );


  buf

  (
    n4719_lo_p_spl_,
    n4719_lo_p
  );


  buf

  (
    n4719_lo_p_spl_0,
    n4719_lo_p_spl_
  );


  buf

  (
    n4719_lo_p_spl_00,
    n4719_lo_p_spl_0
  );


  buf

  (
    n4719_lo_p_spl_000,
    n4719_lo_p_spl_00
  );


  buf

  (
    n4719_lo_p_spl_0000,
    n4719_lo_p_spl_000
  );


  buf

  (
    n4719_lo_p_spl_00000,
    n4719_lo_p_spl_0000
  );


  buf

  (
    n4719_lo_p_spl_00001,
    n4719_lo_p_spl_0000
  );


  buf

  (
    n4719_lo_p_spl_0001,
    n4719_lo_p_spl_000
  );


  buf

  (
    n4719_lo_p_spl_00010,
    n4719_lo_p_spl_0001
  );


  buf

  (
    n4719_lo_p_spl_00011,
    n4719_lo_p_spl_0001
  );


  buf

  (
    n4719_lo_p_spl_001,
    n4719_lo_p_spl_00
  );


  buf

  (
    n4719_lo_p_spl_0010,
    n4719_lo_p_spl_001
  );


  buf

  (
    n4719_lo_p_spl_00100,
    n4719_lo_p_spl_0010
  );


  buf

  (
    n4719_lo_p_spl_00101,
    n4719_lo_p_spl_0010
  );


  buf

  (
    n4719_lo_p_spl_0011,
    n4719_lo_p_spl_001
  );


  buf

  (
    n4719_lo_p_spl_00110,
    n4719_lo_p_spl_0011
  );


  buf

  (
    n4719_lo_p_spl_00111,
    n4719_lo_p_spl_0011
  );


  buf

  (
    n4719_lo_p_spl_01,
    n4719_lo_p_spl_0
  );


  buf

  (
    n4719_lo_p_spl_010,
    n4719_lo_p_spl_01
  );


  buf

  (
    n4719_lo_p_spl_0100,
    n4719_lo_p_spl_010
  );


  buf

  (
    n4719_lo_p_spl_01000,
    n4719_lo_p_spl_0100
  );


  buf

  (
    n4719_lo_p_spl_0101,
    n4719_lo_p_spl_010
  );


  buf

  (
    n4719_lo_p_spl_011,
    n4719_lo_p_spl_01
  );


  buf

  (
    n4719_lo_p_spl_0110,
    n4719_lo_p_spl_011
  );


  buf

  (
    n4719_lo_p_spl_0111,
    n4719_lo_p_spl_011
  );


  buf

  (
    n4719_lo_p_spl_1,
    n4719_lo_p_spl_
  );


  buf

  (
    n4719_lo_p_spl_10,
    n4719_lo_p_spl_1
  );


  buf

  (
    n4719_lo_p_spl_100,
    n4719_lo_p_spl_10
  );


  buf

  (
    n4719_lo_p_spl_1000,
    n4719_lo_p_spl_100
  );


  buf

  (
    n4719_lo_p_spl_1001,
    n4719_lo_p_spl_100
  );


  buf

  (
    n4719_lo_p_spl_101,
    n4719_lo_p_spl_10
  );


  buf

  (
    n4719_lo_p_spl_1010,
    n4719_lo_p_spl_101
  );


  buf

  (
    n4719_lo_p_spl_1011,
    n4719_lo_p_spl_101
  );


  buf

  (
    n4719_lo_p_spl_11,
    n4719_lo_p_spl_1
  );


  buf

  (
    n4719_lo_p_spl_110,
    n4719_lo_p_spl_11
  );


  buf

  (
    n4719_lo_p_spl_1100,
    n4719_lo_p_spl_110
  );


  buf

  (
    n4719_lo_p_spl_1101,
    n4719_lo_p_spl_110
  );


  buf

  (
    n4719_lo_p_spl_111,
    n4719_lo_p_spl_11
  );


  buf

  (
    n4719_lo_p_spl_1110,
    n4719_lo_p_spl_111
  );


  buf

  (
    n4719_lo_p_spl_1111,
    n4719_lo_p_spl_111
  );


  buf

  (
    n4731_lo_p_spl_,
    n4731_lo_p
  );


  buf

  (
    n4731_lo_p_spl_0,
    n4731_lo_p_spl_
  );


  buf

  (
    n4731_lo_p_spl_00,
    n4731_lo_p_spl_0
  );


  buf

  (
    n4731_lo_p_spl_000,
    n4731_lo_p_spl_00
  );


  buf

  (
    n4731_lo_p_spl_0000,
    n4731_lo_p_spl_000
  );


  buf

  (
    n4731_lo_p_spl_00000,
    n4731_lo_p_spl_0000
  );


  buf

  (
    n4731_lo_p_spl_00001,
    n4731_lo_p_spl_0000
  );


  buf

  (
    n4731_lo_p_spl_0001,
    n4731_lo_p_spl_000
  );


  buf

  (
    n4731_lo_p_spl_00010,
    n4731_lo_p_spl_0001
  );


  buf

  (
    n4731_lo_p_spl_00011,
    n4731_lo_p_spl_0001
  );


  buf

  (
    n4731_lo_p_spl_001,
    n4731_lo_p_spl_00
  );


  buf

  (
    n4731_lo_p_spl_0010,
    n4731_lo_p_spl_001
  );


  buf

  (
    n4731_lo_p_spl_00100,
    n4731_lo_p_spl_0010
  );


  buf

  (
    n4731_lo_p_spl_00101,
    n4731_lo_p_spl_0010
  );


  buf

  (
    n4731_lo_p_spl_0011,
    n4731_lo_p_spl_001
  );


  buf

  (
    n4731_lo_p_spl_00110,
    n4731_lo_p_spl_0011
  );


  buf

  (
    n4731_lo_p_spl_00111,
    n4731_lo_p_spl_0011
  );


  buf

  (
    n4731_lo_p_spl_01,
    n4731_lo_p_spl_0
  );


  buf

  (
    n4731_lo_p_spl_010,
    n4731_lo_p_spl_01
  );


  buf

  (
    n4731_lo_p_spl_0100,
    n4731_lo_p_spl_010
  );


  buf

  (
    n4731_lo_p_spl_01000,
    n4731_lo_p_spl_0100
  );


  buf

  (
    n4731_lo_p_spl_0101,
    n4731_lo_p_spl_010
  );


  buf

  (
    n4731_lo_p_spl_011,
    n4731_lo_p_spl_01
  );


  buf

  (
    n4731_lo_p_spl_0110,
    n4731_lo_p_spl_011
  );


  buf

  (
    n4731_lo_p_spl_0111,
    n4731_lo_p_spl_011
  );


  buf

  (
    n4731_lo_p_spl_1,
    n4731_lo_p_spl_
  );


  buf

  (
    n4731_lo_p_spl_10,
    n4731_lo_p_spl_1
  );


  buf

  (
    n4731_lo_p_spl_100,
    n4731_lo_p_spl_10
  );


  buf

  (
    n4731_lo_p_spl_1000,
    n4731_lo_p_spl_100
  );


  buf

  (
    n4731_lo_p_spl_1001,
    n4731_lo_p_spl_100
  );


  buf

  (
    n4731_lo_p_spl_101,
    n4731_lo_p_spl_10
  );


  buf

  (
    n4731_lo_p_spl_1010,
    n4731_lo_p_spl_101
  );


  buf

  (
    n4731_lo_p_spl_1011,
    n4731_lo_p_spl_101
  );


  buf

  (
    n4731_lo_p_spl_11,
    n4731_lo_p_spl_1
  );


  buf

  (
    n4731_lo_p_spl_110,
    n4731_lo_p_spl_11
  );


  buf

  (
    n4731_lo_p_spl_1100,
    n4731_lo_p_spl_110
  );


  buf

  (
    n4731_lo_p_spl_1101,
    n4731_lo_p_spl_110
  );


  buf

  (
    n4731_lo_p_spl_111,
    n4731_lo_p_spl_11
  );


  buf

  (
    n4731_lo_p_spl_1110,
    n4731_lo_p_spl_111
  );


  buf

  (
    n4731_lo_p_spl_1111,
    n4731_lo_p_spl_111
  );


  buf

  (
    n2859_lo_p_spl_,
    n2859_lo_p
  );


  buf

  (
    n2859_lo_p_spl_0,
    n2859_lo_p_spl_
  );


  buf

  (
    n2859_lo_n_spl_,
    n2859_lo_n
  );


  buf

  (
    n2859_lo_n_spl_0,
    n2859_lo_n_spl_
  );


  buf

  (
    g1557_n_spl_,
    g1557_n
  );


  buf

  (
    n4719_lo_n_spl_,
    n4719_lo_n
  );


  buf

  (
    n4719_lo_n_spl_0,
    n4719_lo_n_spl_
  );


  buf

  (
    n4719_lo_n_spl_00,
    n4719_lo_n_spl_0
  );


  buf

  (
    n4719_lo_n_spl_000,
    n4719_lo_n_spl_00
  );


  buf

  (
    n4719_lo_n_spl_0000,
    n4719_lo_n_spl_000
  );


  buf

  (
    n4719_lo_n_spl_0001,
    n4719_lo_n_spl_000
  );


  buf

  (
    n4719_lo_n_spl_001,
    n4719_lo_n_spl_00
  );


  buf

  (
    n4719_lo_n_spl_0010,
    n4719_lo_n_spl_001
  );


  buf

  (
    n4719_lo_n_spl_0011,
    n4719_lo_n_spl_001
  );


  buf

  (
    n4719_lo_n_spl_01,
    n4719_lo_n_spl_0
  );


  buf

  (
    n4719_lo_n_spl_010,
    n4719_lo_n_spl_01
  );


  buf

  (
    n4719_lo_n_spl_0100,
    n4719_lo_n_spl_010
  );


  buf

  (
    n4719_lo_n_spl_0101,
    n4719_lo_n_spl_010
  );


  buf

  (
    n4719_lo_n_spl_011,
    n4719_lo_n_spl_01
  );


  buf

  (
    n4719_lo_n_spl_0110,
    n4719_lo_n_spl_011
  );


  buf

  (
    n4719_lo_n_spl_0111,
    n4719_lo_n_spl_011
  );


  buf

  (
    n4719_lo_n_spl_1,
    n4719_lo_n_spl_
  );


  buf

  (
    n4719_lo_n_spl_10,
    n4719_lo_n_spl_1
  );


  buf

  (
    n4719_lo_n_spl_100,
    n4719_lo_n_spl_10
  );


  buf

  (
    n4719_lo_n_spl_101,
    n4719_lo_n_spl_10
  );


  buf

  (
    n4719_lo_n_spl_11,
    n4719_lo_n_spl_1
  );


  buf

  (
    n4719_lo_n_spl_110,
    n4719_lo_n_spl_11
  );


  buf

  (
    n4719_lo_n_spl_111,
    n4719_lo_n_spl_11
  );


  buf

  (
    n4731_lo_n_spl_,
    n4731_lo_n
  );


  buf

  (
    n4731_lo_n_spl_0,
    n4731_lo_n_spl_
  );


  buf

  (
    n4731_lo_n_spl_00,
    n4731_lo_n_spl_0
  );


  buf

  (
    n4731_lo_n_spl_000,
    n4731_lo_n_spl_00
  );


  buf

  (
    n4731_lo_n_spl_0000,
    n4731_lo_n_spl_000
  );


  buf

  (
    n4731_lo_n_spl_0001,
    n4731_lo_n_spl_000
  );


  buf

  (
    n4731_lo_n_spl_001,
    n4731_lo_n_spl_00
  );


  buf

  (
    n4731_lo_n_spl_0010,
    n4731_lo_n_spl_001
  );


  buf

  (
    n4731_lo_n_spl_0011,
    n4731_lo_n_spl_001
  );


  buf

  (
    n4731_lo_n_spl_01,
    n4731_lo_n_spl_0
  );


  buf

  (
    n4731_lo_n_spl_010,
    n4731_lo_n_spl_01
  );


  buf

  (
    n4731_lo_n_spl_0100,
    n4731_lo_n_spl_010
  );


  buf

  (
    n4731_lo_n_spl_0101,
    n4731_lo_n_spl_010
  );


  buf

  (
    n4731_lo_n_spl_011,
    n4731_lo_n_spl_01
  );


  buf

  (
    n4731_lo_n_spl_0110,
    n4731_lo_n_spl_011
  );


  buf

  (
    n4731_lo_n_spl_0111,
    n4731_lo_n_spl_011
  );


  buf

  (
    n4731_lo_n_spl_1,
    n4731_lo_n_spl_
  );


  buf

  (
    n4731_lo_n_spl_10,
    n4731_lo_n_spl_1
  );


  buf

  (
    n4731_lo_n_spl_100,
    n4731_lo_n_spl_10
  );


  buf

  (
    n4731_lo_n_spl_101,
    n4731_lo_n_spl_10
  );


  buf

  (
    n4731_lo_n_spl_11,
    n4731_lo_n_spl_1
  );


  buf

  (
    n4731_lo_n_spl_110,
    n4731_lo_n_spl_11
  );


  buf

  (
    n4731_lo_n_spl_111,
    n4731_lo_n_spl_11
  );


  buf

  (
    g1566_n_spl_,
    g1566_n
  );


  buf

  (
    g1566_n_spl_0,
    g1566_n_spl_
  );


  buf

  (
    g1566_p_spl_,
    g1566_p
  );


  buf

  (
    g1566_p_spl_0,
    g1566_p_spl_
  );


  buf

  (
    g1570_n_spl_,
    g1570_n
  );


  buf

  (
    n2631_lo_p_spl_,
    n2631_lo_p
  );


  buf

  (
    n2631_lo_p_spl_0,
    n2631_lo_p_spl_
  );


  buf

  (
    n2631_lo_n_spl_,
    n2631_lo_n
  );


  buf

  (
    n2631_lo_n_spl_0,
    n2631_lo_n_spl_
  );


  buf

  (
    g1581_n_spl_,
    g1581_n
  );


  buf

  (
    G3228_o2_p_spl_,
    G3228_o2_p
  );


  buf

  (
    G4137_o2_n_spl_,
    G4137_o2_n
  );


  buf

  (
    G3228_o2_n_spl_,
    G3228_o2_n
  );


  buf

  (
    G4137_o2_p_spl_,
    G4137_o2_p
  );


  buf

  (
    g1592_p_spl_,
    g1592_p
  );


  buf

  (
    g1592_p_spl_0,
    g1592_p_spl_
  );


  buf

  (
    g1592_p_spl_00,
    g1592_p_spl_0
  );


  buf

  (
    g1592_p_spl_1,
    g1592_p_spl_
  );


  buf

  (
    g1592_n_spl_,
    g1592_n
  );


  buf

  (
    g1592_n_spl_0,
    g1592_n_spl_
  );


  buf

  (
    g1592_n_spl_00,
    g1592_n_spl_0
  );


  buf

  (
    g1592_n_spl_1,
    g1592_n_spl_
  );


  buf

  (
    g1596_p_spl_,
    g1596_p
  );


  buf

  (
    g1596_n_spl_,
    g1596_n
  );


  buf

  (
    G2752_o2_n_spl_,
    G2752_o2_n
  );


  buf

  (
    g1563_n_spl_,
    g1563_n
  );


  buf

  (
    g1563_n_spl_0,
    g1563_n_spl_
  );


  buf

  (
    g1563_n_spl_00,
    g1563_n_spl_0
  );


  buf

  (
    g1563_n_spl_1,
    g1563_n_spl_
  );


  buf

  (
    n4683_lo_p_spl_,
    n4683_lo_p
  );


  buf

  (
    n4683_lo_p_spl_0,
    n4683_lo_p_spl_
  );


  buf

  (
    n4683_lo_p_spl_00,
    n4683_lo_p_spl_0
  );


  buf

  (
    n4683_lo_p_spl_000,
    n4683_lo_p_spl_00
  );


  buf

  (
    n4683_lo_p_spl_0000,
    n4683_lo_p_spl_000
  );


  buf

  (
    n4683_lo_p_spl_0001,
    n4683_lo_p_spl_000
  );


  buf

  (
    n4683_lo_p_spl_001,
    n4683_lo_p_spl_00
  );


  buf

  (
    n4683_lo_p_spl_0010,
    n4683_lo_p_spl_001
  );


  buf

  (
    n4683_lo_p_spl_0011,
    n4683_lo_p_spl_001
  );


  buf

  (
    n4683_lo_p_spl_01,
    n4683_lo_p_spl_0
  );


  buf

  (
    n4683_lo_p_spl_010,
    n4683_lo_p_spl_01
  );


  buf

  (
    n4683_lo_p_spl_011,
    n4683_lo_p_spl_01
  );


  buf

  (
    n4683_lo_p_spl_1,
    n4683_lo_p_spl_
  );


  buf

  (
    n4683_lo_p_spl_10,
    n4683_lo_p_spl_1
  );


  buf

  (
    n4683_lo_p_spl_100,
    n4683_lo_p_spl_10
  );


  buf

  (
    n4683_lo_p_spl_101,
    n4683_lo_p_spl_10
  );


  buf

  (
    n4683_lo_p_spl_11,
    n4683_lo_p_spl_1
  );


  buf

  (
    n4683_lo_p_spl_110,
    n4683_lo_p_spl_11
  );


  buf

  (
    n4683_lo_p_spl_111,
    n4683_lo_p_spl_11
  );


  buf

  (
    n4671_lo_p_spl_,
    n4671_lo_p
  );


  buf

  (
    n4671_lo_p_spl_0,
    n4671_lo_p_spl_
  );


  buf

  (
    n4671_lo_p_spl_00,
    n4671_lo_p_spl_0
  );


  buf

  (
    n4671_lo_p_spl_000,
    n4671_lo_p_spl_00
  );


  buf

  (
    n4671_lo_p_spl_0000,
    n4671_lo_p_spl_000
  );


  buf

  (
    n4671_lo_p_spl_0001,
    n4671_lo_p_spl_000
  );


  buf

  (
    n4671_lo_p_spl_001,
    n4671_lo_p_spl_00
  );


  buf

  (
    n4671_lo_p_spl_0010,
    n4671_lo_p_spl_001
  );


  buf

  (
    n4671_lo_p_spl_0011,
    n4671_lo_p_spl_001
  );


  buf

  (
    n4671_lo_p_spl_01,
    n4671_lo_p_spl_0
  );


  buf

  (
    n4671_lo_p_spl_010,
    n4671_lo_p_spl_01
  );


  buf

  (
    n4671_lo_p_spl_011,
    n4671_lo_p_spl_01
  );


  buf

  (
    n4671_lo_p_spl_1,
    n4671_lo_p_spl_
  );


  buf

  (
    n4671_lo_p_spl_10,
    n4671_lo_p_spl_1
  );


  buf

  (
    n4671_lo_p_spl_100,
    n4671_lo_p_spl_10
  );


  buf

  (
    n4671_lo_p_spl_101,
    n4671_lo_p_spl_10
  );


  buf

  (
    n4671_lo_p_spl_11,
    n4671_lo_p_spl_1
  );


  buf

  (
    n4671_lo_p_spl_110,
    n4671_lo_p_spl_11
  );


  buf

  (
    n4671_lo_p_spl_111,
    n4671_lo_p_spl_11
  );


  buf

  (
    g1587_n_spl_,
    g1587_n
  );


  buf

  (
    g1587_n_spl_0,
    g1587_n_spl_
  );


  buf

  (
    g1587_n_spl_00,
    g1587_n_spl_0
  );


  buf

  (
    g1587_n_spl_1,
    g1587_n_spl_
  );


  buf

  (
    n4683_lo_n_spl_,
    n4683_lo_n
  );


  buf

  (
    n4683_lo_n_spl_0,
    n4683_lo_n_spl_
  );


  buf

  (
    n4683_lo_n_spl_00,
    n4683_lo_n_spl_0
  );


  buf

  (
    n4683_lo_n_spl_000,
    n4683_lo_n_spl_00
  );


  buf

  (
    n4683_lo_n_spl_0000,
    n4683_lo_n_spl_000
  );


  buf

  (
    n4683_lo_n_spl_0001,
    n4683_lo_n_spl_000
  );


  buf

  (
    n4683_lo_n_spl_001,
    n4683_lo_n_spl_00
  );


  buf

  (
    n4683_lo_n_spl_0010,
    n4683_lo_n_spl_001
  );


  buf

  (
    n4683_lo_n_spl_0011,
    n4683_lo_n_spl_001
  );


  buf

  (
    n4683_lo_n_spl_01,
    n4683_lo_n_spl_0
  );


  buf

  (
    n4683_lo_n_spl_010,
    n4683_lo_n_spl_01
  );


  buf

  (
    n4683_lo_n_spl_011,
    n4683_lo_n_spl_01
  );


  buf

  (
    n4683_lo_n_spl_1,
    n4683_lo_n_spl_
  );


  buf

  (
    n4683_lo_n_spl_10,
    n4683_lo_n_spl_1
  );


  buf

  (
    n4683_lo_n_spl_100,
    n4683_lo_n_spl_10
  );


  buf

  (
    n4683_lo_n_spl_101,
    n4683_lo_n_spl_10
  );


  buf

  (
    n4683_lo_n_spl_11,
    n4683_lo_n_spl_1
  );


  buf

  (
    n4683_lo_n_spl_110,
    n4683_lo_n_spl_11
  );


  buf

  (
    n4683_lo_n_spl_111,
    n4683_lo_n_spl_11
  );


  buf

  (
    n2643_lo_p_spl_,
    n2643_lo_p
  );


  buf

  (
    n4671_lo_n_spl_,
    n4671_lo_n
  );


  buf

  (
    n4671_lo_n_spl_0,
    n4671_lo_n_spl_
  );


  buf

  (
    n4671_lo_n_spl_00,
    n4671_lo_n_spl_0
  );


  buf

  (
    n4671_lo_n_spl_000,
    n4671_lo_n_spl_00
  );


  buf

  (
    n4671_lo_n_spl_0000,
    n4671_lo_n_spl_000
  );


  buf

  (
    n4671_lo_n_spl_0001,
    n4671_lo_n_spl_000
  );


  buf

  (
    n4671_lo_n_spl_001,
    n4671_lo_n_spl_00
  );


  buf

  (
    n4671_lo_n_spl_0010,
    n4671_lo_n_spl_001
  );


  buf

  (
    n4671_lo_n_spl_0011,
    n4671_lo_n_spl_001
  );


  buf

  (
    n4671_lo_n_spl_01,
    n4671_lo_n_spl_0
  );


  buf

  (
    n4671_lo_n_spl_010,
    n4671_lo_n_spl_01
  );


  buf

  (
    n4671_lo_n_spl_011,
    n4671_lo_n_spl_01
  );


  buf

  (
    n4671_lo_n_spl_1,
    n4671_lo_n_spl_
  );


  buf

  (
    n4671_lo_n_spl_10,
    n4671_lo_n_spl_1
  );


  buf

  (
    n4671_lo_n_spl_100,
    n4671_lo_n_spl_10
  );


  buf

  (
    n4671_lo_n_spl_101,
    n4671_lo_n_spl_10
  );


  buf

  (
    n4671_lo_n_spl_11,
    n4671_lo_n_spl_1
  );


  buf

  (
    n4671_lo_n_spl_110,
    n4671_lo_n_spl_11
  );


  buf

  (
    n4671_lo_n_spl_111,
    n4671_lo_n_spl_11
  );


  buf

  (
    n2871_lo_p_spl_,
    n2871_lo_p
  );


  buf

  (
    g1616_p_spl_,
    g1616_p
  );


  buf

  (
    g1616_n_spl_,
    g1616_n
  );


  buf

  (
    g1618_p_spl_,
    g1618_p
  );


  buf

  (
    g1618_n_spl_,
    g1618_n
  );


  buf

  (
    g1621_p_spl_,
    g1621_p
  );


  buf

  (
    g1621_n_spl_,
    g1621_n
  );


  buf

  (
    g1629_n_spl_,
    g1629_n
  );


  buf

  (
    g1643_n_spl_,
    g1643_n
  );


  buf

  (
    g1658_n_spl_,
    g1658_n
  );


  buf

  (
    n4695_lo_p_spl_,
    n4695_lo_p
  );


  buf

  (
    n4695_lo_p_spl_0,
    n4695_lo_p_spl_
  );


  buf

  (
    n4695_lo_p_spl_00,
    n4695_lo_p_spl_0
  );


  buf

  (
    n4695_lo_p_spl_000,
    n4695_lo_p_spl_00
  );


  buf

  (
    n4695_lo_p_spl_0000,
    n4695_lo_p_spl_000
  );


  buf

  (
    n4695_lo_p_spl_0001,
    n4695_lo_p_spl_000
  );


  buf

  (
    n4695_lo_p_spl_001,
    n4695_lo_p_spl_00
  );


  buf

  (
    n4695_lo_p_spl_0010,
    n4695_lo_p_spl_001
  );


  buf

  (
    n4695_lo_p_spl_0011,
    n4695_lo_p_spl_001
  );


  buf

  (
    n4695_lo_p_spl_01,
    n4695_lo_p_spl_0
  );


  buf

  (
    n4695_lo_p_spl_010,
    n4695_lo_p_spl_01
  );


  buf

  (
    n4695_lo_p_spl_011,
    n4695_lo_p_spl_01
  );


  buf

  (
    n4695_lo_p_spl_1,
    n4695_lo_p_spl_
  );


  buf

  (
    n4695_lo_p_spl_10,
    n4695_lo_p_spl_1
  );


  buf

  (
    n4695_lo_p_spl_100,
    n4695_lo_p_spl_10
  );


  buf

  (
    n4695_lo_p_spl_101,
    n4695_lo_p_spl_10
  );


  buf

  (
    n4695_lo_p_spl_11,
    n4695_lo_p_spl_1
  );


  buf

  (
    n4695_lo_p_spl_110,
    n4695_lo_p_spl_11
  );


  buf

  (
    n4695_lo_p_spl_111,
    n4695_lo_p_spl_11
  );


  buf

  (
    n4707_lo_p_spl_,
    n4707_lo_p
  );


  buf

  (
    n4707_lo_p_spl_0,
    n4707_lo_p_spl_
  );


  buf

  (
    n4707_lo_p_spl_00,
    n4707_lo_p_spl_0
  );


  buf

  (
    n4707_lo_p_spl_000,
    n4707_lo_p_spl_00
  );


  buf

  (
    n4707_lo_p_spl_0000,
    n4707_lo_p_spl_000
  );


  buf

  (
    n4707_lo_p_spl_0001,
    n4707_lo_p_spl_000
  );


  buf

  (
    n4707_lo_p_spl_001,
    n4707_lo_p_spl_00
  );


  buf

  (
    n4707_lo_p_spl_0010,
    n4707_lo_p_spl_001
  );


  buf

  (
    n4707_lo_p_spl_0011,
    n4707_lo_p_spl_001
  );


  buf

  (
    n4707_lo_p_spl_01,
    n4707_lo_p_spl_0
  );


  buf

  (
    n4707_lo_p_spl_010,
    n4707_lo_p_spl_01
  );


  buf

  (
    n4707_lo_p_spl_011,
    n4707_lo_p_spl_01
  );


  buf

  (
    n4707_lo_p_spl_1,
    n4707_lo_p_spl_
  );


  buf

  (
    n4707_lo_p_spl_10,
    n4707_lo_p_spl_1
  );


  buf

  (
    n4707_lo_p_spl_100,
    n4707_lo_p_spl_10
  );


  buf

  (
    n4707_lo_p_spl_101,
    n4707_lo_p_spl_10
  );


  buf

  (
    n4707_lo_p_spl_11,
    n4707_lo_p_spl_1
  );


  buf

  (
    n4707_lo_p_spl_110,
    n4707_lo_p_spl_11
  );


  buf

  (
    n4707_lo_p_spl_111,
    n4707_lo_p_spl_11
  );


  buf

  (
    n4695_lo_n_spl_,
    n4695_lo_n
  );


  buf

  (
    n4695_lo_n_spl_0,
    n4695_lo_n_spl_
  );


  buf

  (
    n4695_lo_n_spl_00,
    n4695_lo_n_spl_0
  );


  buf

  (
    n4695_lo_n_spl_000,
    n4695_lo_n_spl_00
  );


  buf

  (
    n4695_lo_n_spl_0000,
    n4695_lo_n_spl_000
  );


  buf

  (
    n4695_lo_n_spl_0001,
    n4695_lo_n_spl_000
  );


  buf

  (
    n4695_lo_n_spl_001,
    n4695_lo_n_spl_00
  );


  buf

  (
    n4695_lo_n_spl_0010,
    n4695_lo_n_spl_001
  );


  buf

  (
    n4695_lo_n_spl_0011,
    n4695_lo_n_spl_001
  );


  buf

  (
    n4695_lo_n_spl_01,
    n4695_lo_n_spl_0
  );


  buf

  (
    n4695_lo_n_spl_010,
    n4695_lo_n_spl_01
  );


  buf

  (
    n4695_lo_n_spl_011,
    n4695_lo_n_spl_01
  );


  buf

  (
    n4695_lo_n_spl_1,
    n4695_lo_n_spl_
  );


  buf

  (
    n4695_lo_n_spl_10,
    n4695_lo_n_spl_1
  );


  buf

  (
    n4695_lo_n_spl_100,
    n4695_lo_n_spl_10
  );


  buf

  (
    n4695_lo_n_spl_101,
    n4695_lo_n_spl_10
  );


  buf

  (
    n4695_lo_n_spl_11,
    n4695_lo_n_spl_1
  );


  buf

  (
    n4695_lo_n_spl_110,
    n4695_lo_n_spl_11
  );


  buf

  (
    n4695_lo_n_spl_111,
    n4695_lo_n_spl_11
  );


  buf

  (
    n4707_lo_n_spl_,
    n4707_lo_n
  );


  buf

  (
    n4707_lo_n_spl_0,
    n4707_lo_n_spl_
  );


  buf

  (
    n4707_lo_n_spl_00,
    n4707_lo_n_spl_0
  );


  buf

  (
    n4707_lo_n_spl_000,
    n4707_lo_n_spl_00
  );


  buf

  (
    n4707_lo_n_spl_0000,
    n4707_lo_n_spl_000
  );


  buf

  (
    n4707_lo_n_spl_0001,
    n4707_lo_n_spl_000
  );


  buf

  (
    n4707_lo_n_spl_001,
    n4707_lo_n_spl_00
  );


  buf

  (
    n4707_lo_n_spl_0010,
    n4707_lo_n_spl_001
  );


  buf

  (
    n4707_lo_n_spl_0011,
    n4707_lo_n_spl_001
  );


  buf

  (
    n4707_lo_n_spl_01,
    n4707_lo_n_spl_0
  );


  buf

  (
    n4707_lo_n_spl_010,
    n4707_lo_n_spl_01
  );


  buf

  (
    n4707_lo_n_spl_011,
    n4707_lo_n_spl_01
  );


  buf

  (
    n4707_lo_n_spl_1,
    n4707_lo_n_spl_
  );


  buf

  (
    n4707_lo_n_spl_10,
    n4707_lo_n_spl_1
  );


  buf

  (
    n4707_lo_n_spl_100,
    n4707_lo_n_spl_10
  );


  buf

  (
    n4707_lo_n_spl_101,
    n4707_lo_n_spl_10
  );


  buf

  (
    n4707_lo_n_spl_11,
    n4707_lo_n_spl_1
  );


  buf

  (
    n4707_lo_n_spl_110,
    n4707_lo_n_spl_11
  );


  buf

  (
    n4707_lo_n_spl_111,
    n4707_lo_n_spl_11
  );


  buf

  (
    g1679_p_spl_,
    g1679_p
  );


  buf

  (
    g1679_n_spl_,
    g1679_n
  );


  buf

  (
    g1681_p_spl_,
    g1681_p
  );


  buf

  (
    g1681_n_spl_,
    g1681_n
  );


  buf

  (
    g1683_p_spl_,
    g1683_p
  );


  buf

  (
    g1683_p_spl_0,
    g1683_p_spl_
  );


  buf

  (
    g1683_n_spl_,
    g1683_n
  );


  buf

  (
    g1683_n_spl_0,
    g1683_n_spl_
  );


  buf

  (
    g1685_p_spl_,
    g1685_p
  );


  buf

  (
    g1685_n_spl_,
    g1685_n
  );


  buf

  (
    g1693_n_spl_,
    g1693_n
  );


  buf

  (
    g1707_n_spl_,
    g1707_n
  );


  buf

  (
    g1722_n_spl_,
    g1722_n
  );


  buf

  (
    g1734_n_spl_,
    g1734_n
  );


  buf

  (
    g1746_p_spl_,
    g1746_p
  );


  buf

  (
    g1743_n_spl_,
    g1743_n
  );


  buf

  (
    g1746_n_spl_,
    g1746_n
  );


  buf

  (
    g1743_p_spl_,
    g1743_p
  );


  buf

  (
    g1751_p_spl_,
    g1751_p
  );


  buf

  (
    g1751_p_spl_0,
    g1751_p_spl_
  );


  buf

  (
    g1751_p_spl_1,
    g1751_p_spl_
  );


  buf

  (
    g1750_n_spl_,
    g1750_n
  );


  buf

  (
    g1750_n_spl_0,
    g1750_n_spl_
  );


  buf

  (
    g1750_n_spl_1,
    g1750_n_spl_
  );


  buf

  (
    g1751_n_spl_,
    g1751_n
  );


  buf

  (
    g1751_n_spl_0,
    g1751_n_spl_
  );


  buf

  (
    g1751_n_spl_1,
    g1751_n_spl_
  );


  buf

  (
    g1750_p_spl_,
    g1750_p
  );


  buf

  (
    g1750_p_spl_0,
    g1750_p_spl_
  );


  buf

  (
    g1750_p_spl_1,
    g1750_p_spl_
  );


  buf

  (
    G3674_o2_p_spl_,
    G3674_o2_p
  );


  buf

  (
    G3674_o2_p_spl_0,
    G3674_o2_p_spl_
  );


  buf

  (
    G3674_o2_p_spl_1,
    G3674_o2_p_spl_
  );


  buf

  (
    G3674_o2_n_spl_,
    G3674_o2_n
  );


  buf

  (
    G3674_o2_n_spl_0,
    G3674_o2_n_spl_
  );


  buf

  (
    G3674_o2_n_spl_1,
    G3674_o2_n_spl_
  );


  buf

  (
    g1771_p_spl_,
    g1771_p
  );


  buf

  (
    g1768_n_spl_,
    g1768_n
  );


  buf

  (
    g1771_n_spl_,
    g1771_n
  );


  buf

  (
    g1768_p_spl_,
    g1768_p
  );


  buf

  (
    g1776_p_spl_,
    g1776_p
  );


  buf

  (
    g1776_p_spl_0,
    g1776_p_spl_
  );


  buf

  (
    g1776_p_spl_1,
    g1776_p_spl_
  );


  buf

  (
    g1775_n_spl_,
    g1775_n
  );


  buf

  (
    g1775_n_spl_0,
    g1775_n_spl_
  );


  buf

  (
    g1775_n_spl_1,
    g1775_n_spl_
  );


  buf

  (
    g1776_n_spl_,
    g1776_n
  );


  buf

  (
    g1776_n_spl_0,
    g1776_n_spl_
  );


  buf

  (
    g1776_n_spl_1,
    g1776_n_spl_
  );


  buf

  (
    g1775_p_spl_,
    g1775_p
  );


  buf

  (
    g1775_p_spl_0,
    g1775_p_spl_
  );


  buf

  (
    g1775_p_spl_1,
    g1775_p_spl_
  );


  buf

  (
    G3685_o2_n_spl_,
    G3685_o2_n
  );


  buf

  (
    G3685_o2_n_spl_0,
    G3685_o2_n_spl_
  );


  buf

  (
    G3685_o2_n_spl_1,
    G3685_o2_n_spl_
  );


  buf

  (
    G3685_o2_p_spl_,
    G3685_o2_p
  );


  buf

  (
    G3685_o2_p_spl_0,
    G3685_o2_p_spl_
  );


  buf

  (
    G3685_o2_p_spl_1,
    G3685_o2_p_spl_
  );


  buf

  (
    g1792_p_spl_,
    g1792_p
  );


  buf

  (
    g1792_p_spl_0,
    g1792_p_spl_
  );


  buf

  (
    g1792_p_spl_1,
    g1792_p_spl_
  );


  buf

  (
    g1792_n_spl_,
    g1792_n
  );


  buf

  (
    g1792_n_spl_0,
    g1792_n_spl_
  );


  buf

  (
    g1792_n_spl_1,
    g1792_n_spl_
  );


  buf

  (
    g1795_n_spl_,
    g1795_n
  );


  buf

  (
    g1804_n_spl_,
    g1804_n
  );


  buf

  (
    g1815_n_spl_,
    g1815_n
  );


  buf

  (
    g1827_n_spl_,
    g1827_n
  );


  buf

  (
    g1838_n_spl_,
    g1838_n
  );


  buf

  (
    g1847_n_spl_,
    g1847_n
  );


  buf

  (
    g1858_n_spl_,
    g1858_n
  );


  buf

  (
    g1601_n_spl_,
    g1601_n
  );


  buf

  (
    g1601_n_spl_0,
    g1601_n_spl_
  );


  buf

  (
    g1601_n_spl_1,
    g1601_n_spl_
  );


  buf

  (
    n4503_lo_p_spl_,
    n4503_lo_p
  );


  buf

  (
    n4503_lo_p_spl_0,
    n4503_lo_p_spl_
  );


  buf

  (
    n4503_lo_p_spl_00,
    n4503_lo_p_spl_0
  );


  buf

  (
    n4503_lo_p_spl_000,
    n4503_lo_p_spl_00
  );


  buf

  (
    n4503_lo_p_spl_0000,
    n4503_lo_p_spl_000
  );


  buf

  (
    n4503_lo_p_spl_0001,
    n4503_lo_p_spl_000
  );


  buf

  (
    n4503_lo_p_spl_001,
    n4503_lo_p_spl_00
  );


  buf

  (
    n4503_lo_p_spl_0010,
    n4503_lo_p_spl_001
  );


  buf

  (
    n4503_lo_p_spl_0011,
    n4503_lo_p_spl_001
  );


  buf

  (
    n4503_lo_p_spl_01,
    n4503_lo_p_spl_0
  );


  buf

  (
    n4503_lo_p_spl_010,
    n4503_lo_p_spl_01
  );


  buf

  (
    n4503_lo_p_spl_011,
    n4503_lo_p_spl_01
  );


  buf

  (
    n4503_lo_p_spl_1,
    n4503_lo_p_spl_
  );


  buf

  (
    n4503_lo_p_spl_10,
    n4503_lo_p_spl_1
  );


  buf

  (
    n4503_lo_p_spl_100,
    n4503_lo_p_spl_10
  );


  buf

  (
    n4503_lo_p_spl_101,
    n4503_lo_p_spl_10
  );


  buf

  (
    n4503_lo_p_spl_11,
    n4503_lo_p_spl_1
  );


  buf

  (
    n4503_lo_p_spl_110,
    n4503_lo_p_spl_11
  );


  buf

  (
    n4503_lo_p_spl_111,
    n4503_lo_p_spl_11
  );


  buf

  (
    n4515_lo_p_spl_,
    n4515_lo_p
  );


  buf

  (
    n4515_lo_p_spl_0,
    n4515_lo_p_spl_
  );


  buf

  (
    n4515_lo_p_spl_00,
    n4515_lo_p_spl_0
  );


  buf

  (
    n4515_lo_p_spl_000,
    n4515_lo_p_spl_00
  );


  buf

  (
    n4515_lo_p_spl_0000,
    n4515_lo_p_spl_000
  );


  buf

  (
    n4515_lo_p_spl_0001,
    n4515_lo_p_spl_000
  );


  buf

  (
    n4515_lo_p_spl_001,
    n4515_lo_p_spl_00
  );


  buf

  (
    n4515_lo_p_spl_0010,
    n4515_lo_p_spl_001
  );


  buf

  (
    n4515_lo_p_spl_0011,
    n4515_lo_p_spl_001
  );


  buf

  (
    n4515_lo_p_spl_01,
    n4515_lo_p_spl_0
  );


  buf

  (
    n4515_lo_p_spl_010,
    n4515_lo_p_spl_01
  );


  buf

  (
    n4515_lo_p_spl_011,
    n4515_lo_p_spl_01
  );


  buf

  (
    n4515_lo_p_spl_1,
    n4515_lo_p_spl_
  );


  buf

  (
    n4515_lo_p_spl_10,
    n4515_lo_p_spl_1
  );


  buf

  (
    n4515_lo_p_spl_100,
    n4515_lo_p_spl_10
  );


  buf

  (
    n4515_lo_p_spl_101,
    n4515_lo_p_spl_10
  );


  buf

  (
    n4515_lo_p_spl_11,
    n4515_lo_p_spl_1
  );


  buf

  (
    n4515_lo_p_spl_110,
    n4515_lo_p_spl_11
  );


  buf

  (
    n4515_lo_p_spl_111,
    n4515_lo_p_spl_11
  );


  buf

  (
    n4503_lo_n_spl_,
    n4503_lo_n
  );


  buf

  (
    n4503_lo_n_spl_0,
    n4503_lo_n_spl_
  );


  buf

  (
    n4503_lo_n_spl_00,
    n4503_lo_n_spl_0
  );


  buf

  (
    n4503_lo_n_spl_000,
    n4503_lo_n_spl_00
  );


  buf

  (
    n4503_lo_n_spl_0000,
    n4503_lo_n_spl_000
  );


  buf

  (
    n4503_lo_n_spl_0001,
    n4503_lo_n_spl_000
  );


  buf

  (
    n4503_lo_n_spl_001,
    n4503_lo_n_spl_00
  );


  buf

  (
    n4503_lo_n_spl_0010,
    n4503_lo_n_spl_001
  );


  buf

  (
    n4503_lo_n_spl_0011,
    n4503_lo_n_spl_001
  );


  buf

  (
    n4503_lo_n_spl_01,
    n4503_lo_n_spl_0
  );


  buf

  (
    n4503_lo_n_spl_010,
    n4503_lo_n_spl_01
  );


  buf

  (
    n4503_lo_n_spl_011,
    n4503_lo_n_spl_01
  );


  buf

  (
    n4503_lo_n_spl_1,
    n4503_lo_n_spl_
  );


  buf

  (
    n4503_lo_n_spl_10,
    n4503_lo_n_spl_1
  );


  buf

  (
    n4503_lo_n_spl_100,
    n4503_lo_n_spl_10
  );


  buf

  (
    n4503_lo_n_spl_101,
    n4503_lo_n_spl_10
  );


  buf

  (
    n4503_lo_n_spl_11,
    n4503_lo_n_spl_1
  );


  buf

  (
    n4503_lo_n_spl_110,
    n4503_lo_n_spl_11
  );


  buf

  (
    n4503_lo_n_spl_111,
    n4503_lo_n_spl_11
  );


  buf

  (
    n3567_lo_p_spl_,
    n3567_lo_p
  );


  buf

  (
    n4515_lo_n_spl_,
    n4515_lo_n
  );


  buf

  (
    n4515_lo_n_spl_0,
    n4515_lo_n_spl_
  );


  buf

  (
    n4515_lo_n_spl_00,
    n4515_lo_n_spl_0
  );


  buf

  (
    n4515_lo_n_spl_000,
    n4515_lo_n_spl_00
  );


  buf

  (
    n4515_lo_n_spl_0000,
    n4515_lo_n_spl_000
  );


  buf

  (
    n4515_lo_n_spl_0001,
    n4515_lo_n_spl_000
  );


  buf

  (
    n4515_lo_n_spl_001,
    n4515_lo_n_spl_00
  );


  buf

  (
    n4515_lo_n_spl_0010,
    n4515_lo_n_spl_001
  );


  buf

  (
    n4515_lo_n_spl_0011,
    n4515_lo_n_spl_001
  );


  buf

  (
    n4515_lo_n_spl_01,
    n4515_lo_n_spl_0
  );


  buf

  (
    n4515_lo_n_spl_010,
    n4515_lo_n_spl_01
  );


  buf

  (
    n4515_lo_n_spl_011,
    n4515_lo_n_spl_01
  );


  buf

  (
    n4515_lo_n_spl_1,
    n4515_lo_n_spl_
  );


  buf

  (
    n4515_lo_n_spl_10,
    n4515_lo_n_spl_1
  );


  buf

  (
    n4515_lo_n_spl_100,
    n4515_lo_n_spl_10
  );


  buf

  (
    n4515_lo_n_spl_101,
    n4515_lo_n_spl_10
  );


  buf

  (
    n4515_lo_n_spl_11,
    n4515_lo_n_spl_1
  );


  buf

  (
    n4515_lo_n_spl_110,
    n4515_lo_n_spl_11
  );


  buf

  (
    n4515_lo_n_spl_111,
    n4515_lo_n_spl_11
  );


  buf

  (
    n3579_lo_p_spl_,
    n3579_lo_p
  );


  buf

  (
    n3375_lo_p_spl_,
    n3375_lo_p
  );


  buf

  (
    n3375_lo_p_spl_0,
    n3375_lo_p_spl_
  );


  buf

  (
    n3375_lo_p_spl_00,
    n3375_lo_p_spl_0
  );


  buf

  (
    n3375_lo_p_spl_000,
    n3375_lo_p_spl_00
  );


  buf

  (
    n3375_lo_p_spl_0000,
    n3375_lo_p_spl_000
  );


  buf

  (
    n3375_lo_p_spl_0001,
    n3375_lo_p_spl_000
  );


  buf

  (
    n3375_lo_p_spl_001,
    n3375_lo_p_spl_00
  );


  buf

  (
    n3375_lo_p_spl_0010,
    n3375_lo_p_spl_001
  );


  buf

  (
    n3375_lo_p_spl_0011,
    n3375_lo_p_spl_001
  );


  buf

  (
    n3375_lo_p_spl_01,
    n3375_lo_p_spl_0
  );


  buf

  (
    n3375_lo_p_spl_010,
    n3375_lo_p_spl_01
  );


  buf

  (
    n3375_lo_p_spl_0100,
    n3375_lo_p_spl_010
  );


  buf

  (
    n3375_lo_p_spl_011,
    n3375_lo_p_spl_01
  );


  buf

  (
    n3375_lo_p_spl_1,
    n3375_lo_p_spl_
  );


  buf

  (
    n3375_lo_p_spl_10,
    n3375_lo_p_spl_1
  );


  buf

  (
    n3375_lo_p_spl_100,
    n3375_lo_p_spl_10
  );


  buf

  (
    n3375_lo_p_spl_101,
    n3375_lo_p_spl_10
  );


  buf

  (
    n3375_lo_p_spl_11,
    n3375_lo_p_spl_1
  );


  buf

  (
    n3375_lo_p_spl_110,
    n3375_lo_p_spl_11
  );


  buf

  (
    n3375_lo_p_spl_111,
    n3375_lo_p_spl_11
  );


  buf

  (
    n4527_lo_p_spl_,
    n4527_lo_p
  );


  buf

  (
    n4527_lo_p_spl_0,
    n4527_lo_p_spl_
  );


  buf

  (
    n4527_lo_p_spl_00,
    n4527_lo_p_spl_0
  );


  buf

  (
    n4527_lo_p_spl_000,
    n4527_lo_p_spl_00
  );


  buf

  (
    n4527_lo_p_spl_0000,
    n4527_lo_p_spl_000
  );


  buf

  (
    n4527_lo_p_spl_0001,
    n4527_lo_p_spl_000
  );


  buf

  (
    n4527_lo_p_spl_001,
    n4527_lo_p_spl_00
  );


  buf

  (
    n4527_lo_p_spl_0010,
    n4527_lo_p_spl_001
  );


  buf

  (
    n4527_lo_p_spl_0011,
    n4527_lo_p_spl_001
  );


  buf

  (
    n4527_lo_p_spl_01,
    n4527_lo_p_spl_0
  );


  buf

  (
    n4527_lo_p_spl_010,
    n4527_lo_p_spl_01
  );


  buf

  (
    n4527_lo_p_spl_011,
    n4527_lo_p_spl_01
  );


  buf

  (
    n4527_lo_p_spl_1,
    n4527_lo_p_spl_
  );


  buf

  (
    n4527_lo_p_spl_10,
    n4527_lo_p_spl_1
  );


  buf

  (
    n4527_lo_p_spl_100,
    n4527_lo_p_spl_10
  );


  buf

  (
    n4527_lo_p_spl_101,
    n4527_lo_p_spl_10
  );


  buf

  (
    n4527_lo_p_spl_11,
    n4527_lo_p_spl_1
  );


  buf

  (
    n4527_lo_p_spl_110,
    n4527_lo_p_spl_11
  );


  buf

  (
    n4527_lo_p_spl_111,
    n4527_lo_p_spl_11
  );


  buf

  (
    n4539_lo_p_spl_,
    n4539_lo_p
  );


  buf

  (
    n4539_lo_p_spl_0,
    n4539_lo_p_spl_
  );


  buf

  (
    n4539_lo_p_spl_00,
    n4539_lo_p_spl_0
  );


  buf

  (
    n4539_lo_p_spl_000,
    n4539_lo_p_spl_00
  );


  buf

  (
    n4539_lo_p_spl_0000,
    n4539_lo_p_spl_000
  );


  buf

  (
    n4539_lo_p_spl_0001,
    n4539_lo_p_spl_000
  );


  buf

  (
    n4539_lo_p_spl_001,
    n4539_lo_p_spl_00
  );


  buf

  (
    n4539_lo_p_spl_0010,
    n4539_lo_p_spl_001
  );


  buf

  (
    n4539_lo_p_spl_0011,
    n4539_lo_p_spl_001
  );


  buf

  (
    n4539_lo_p_spl_01,
    n4539_lo_p_spl_0
  );


  buf

  (
    n4539_lo_p_spl_010,
    n4539_lo_p_spl_01
  );


  buf

  (
    n4539_lo_p_spl_011,
    n4539_lo_p_spl_01
  );


  buf

  (
    n4539_lo_p_spl_1,
    n4539_lo_p_spl_
  );


  buf

  (
    n4539_lo_p_spl_10,
    n4539_lo_p_spl_1
  );


  buf

  (
    n4539_lo_p_spl_100,
    n4539_lo_p_spl_10
  );


  buf

  (
    n4539_lo_p_spl_101,
    n4539_lo_p_spl_10
  );


  buf

  (
    n4539_lo_p_spl_11,
    n4539_lo_p_spl_1
  );


  buf

  (
    n4539_lo_p_spl_110,
    n4539_lo_p_spl_11
  );


  buf

  (
    n4539_lo_p_spl_111,
    n4539_lo_p_spl_11
  );


  buf

  (
    n4527_lo_n_spl_,
    n4527_lo_n
  );


  buf

  (
    n4527_lo_n_spl_0,
    n4527_lo_n_spl_
  );


  buf

  (
    n4527_lo_n_spl_00,
    n4527_lo_n_spl_0
  );


  buf

  (
    n4527_lo_n_spl_000,
    n4527_lo_n_spl_00
  );


  buf

  (
    n4527_lo_n_spl_0000,
    n4527_lo_n_spl_000
  );


  buf

  (
    n4527_lo_n_spl_0001,
    n4527_lo_n_spl_000
  );


  buf

  (
    n4527_lo_n_spl_001,
    n4527_lo_n_spl_00
  );


  buf

  (
    n4527_lo_n_spl_0010,
    n4527_lo_n_spl_001
  );


  buf

  (
    n4527_lo_n_spl_0011,
    n4527_lo_n_spl_001
  );


  buf

  (
    n4527_lo_n_spl_01,
    n4527_lo_n_spl_0
  );


  buf

  (
    n4527_lo_n_spl_010,
    n4527_lo_n_spl_01
  );


  buf

  (
    n4527_lo_n_spl_011,
    n4527_lo_n_spl_01
  );


  buf

  (
    n4527_lo_n_spl_1,
    n4527_lo_n_spl_
  );


  buf

  (
    n4527_lo_n_spl_10,
    n4527_lo_n_spl_1
  );


  buf

  (
    n4527_lo_n_spl_100,
    n4527_lo_n_spl_10
  );


  buf

  (
    n4527_lo_n_spl_101,
    n4527_lo_n_spl_10
  );


  buf

  (
    n4527_lo_n_spl_11,
    n4527_lo_n_spl_1
  );


  buf

  (
    n4527_lo_n_spl_110,
    n4527_lo_n_spl_11
  );


  buf

  (
    n4527_lo_n_spl_111,
    n4527_lo_n_spl_11
  );


  buf

  (
    n4539_lo_n_spl_,
    n4539_lo_n
  );


  buf

  (
    n4539_lo_n_spl_0,
    n4539_lo_n_spl_
  );


  buf

  (
    n4539_lo_n_spl_00,
    n4539_lo_n_spl_0
  );


  buf

  (
    n4539_lo_n_spl_000,
    n4539_lo_n_spl_00
  );


  buf

  (
    n4539_lo_n_spl_0000,
    n4539_lo_n_spl_000
  );


  buf

  (
    n4539_lo_n_spl_0001,
    n4539_lo_n_spl_000
  );


  buf

  (
    n4539_lo_n_spl_001,
    n4539_lo_n_spl_00
  );


  buf

  (
    n4539_lo_n_spl_0010,
    n4539_lo_n_spl_001
  );


  buf

  (
    n4539_lo_n_spl_0011,
    n4539_lo_n_spl_001
  );


  buf

  (
    n4539_lo_n_spl_01,
    n4539_lo_n_spl_0
  );


  buf

  (
    n4539_lo_n_spl_010,
    n4539_lo_n_spl_01
  );


  buf

  (
    n4539_lo_n_spl_011,
    n4539_lo_n_spl_01
  );


  buf

  (
    n4539_lo_n_spl_1,
    n4539_lo_n_spl_
  );


  buf

  (
    n4539_lo_n_spl_10,
    n4539_lo_n_spl_1
  );


  buf

  (
    n4539_lo_n_spl_100,
    n4539_lo_n_spl_10
  );


  buf

  (
    n4539_lo_n_spl_101,
    n4539_lo_n_spl_10
  );


  buf

  (
    n4539_lo_n_spl_11,
    n4539_lo_n_spl_1
  );


  buf

  (
    n4539_lo_n_spl_110,
    n4539_lo_n_spl_11
  );


  buf

  (
    n4539_lo_n_spl_111,
    n4539_lo_n_spl_11
  );


  buf

  (
    g1635_n_spl_,
    g1635_n
  );


  buf

  (
    g1635_n_spl_0,
    g1635_n_spl_
  );


  buf

  (
    g1635_n_spl_00,
    g1635_n_spl_0
  );


  buf

  (
    g1635_n_spl_1,
    g1635_n_spl_
  );


  buf

  (
    g1699_n_spl_,
    g1699_n
  );


  buf

  (
    g1699_n_spl_0,
    g1699_n_spl_
  );


  buf

  (
    g1699_n_spl_00,
    g1699_n_spl_0
  );


  buf

  (
    g1699_n_spl_1,
    g1699_n_spl_
  );


  buf

  (
    n2799_lo_p_spl_,
    n2799_lo_p
  );


  buf

  (
    n2775_lo_p_spl_,
    n2775_lo_p
  );


  buf

  (
    g1649_n_spl_,
    g1649_n
  );


  buf

  (
    g1649_n_spl_0,
    g1649_n_spl_
  );


  buf

  (
    g1649_n_spl_00,
    g1649_n_spl_0
  );


  buf

  (
    g1649_n_spl_1,
    g1649_n_spl_
  );


  buf

  (
    g1713_n_spl_,
    g1713_n
  );


  buf

  (
    g1713_n_spl_0,
    g1713_n_spl_
  );


  buf

  (
    g1713_n_spl_00,
    g1713_n_spl_0
  );


  buf

  (
    g1713_n_spl_1,
    g1713_n_spl_
  );


  buf

  (
    n2931_lo_p_spl_,
    n2931_lo_p
  );


  buf

  (
    n2679_lo_p_spl_,
    n2679_lo_p
  );


  buf

  (
    g1664_n_spl_,
    g1664_n
  );


  buf

  (
    g1664_n_spl_0,
    g1664_n_spl_
  );


  buf

  (
    g1664_n_spl_00,
    g1664_n_spl_0
  );


  buf

  (
    g1664_n_spl_1,
    g1664_n_spl_
  );


  buf

  (
    g1728_n_spl_,
    g1728_n
  );


  buf

  (
    g1728_n_spl_0,
    g1728_n_spl_
  );


  buf

  (
    g1728_n_spl_00,
    g1728_n_spl_0
  );


  buf

  (
    g1728_n_spl_1,
    g1728_n_spl_
  );


  buf

  (
    n2919_lo_p_spl_,
    n2919_lo_p
  );


  buf

  (
    n2667_lo_p_spl_,
    n2667_lo_p
  );


  buf

  (
    g1576_n_spl_,
    g1576_n
  );


  buf

  (
    g1576_n_spl_0,
    g1576_n_spl_
  );


  buf

  (
    g1576_n_spl_00,
    g1576_n_spl_0
  );


  buf

  (
    g1576_n_spl_1,
    g1576_n_spl_
  );


  buf

  (
    g1740_n_spl_,
    g1740_n
  );


  buf

  (
    g1740_n_spl_0,
    g1740_n_spl_
  );


  buf

  (
    g1740_n_spl_00,
    g1740_n_spl_0
  );


  buf

  (
    g1740_n_spl_1,
    g1740_n_spl_
  );


  buf

  (
    n2895_lo_p_spl_,
    n2895_lo_p
  );


  buf

  (
    n2907_lo_p_spl_,
    n2907_lo_p
  );


  buf

  (
    n3639_lo_p_spl_,
    n3639_lo_p
  );


  buf

  (
    n3519_lo_p_spl_,
    n3519_lo_p
  );


  buf

  (
    n3591_lo_p_spl_,
    n3591_lo_p
  );


  buf

  (
    n3471_lo_p_spl_,
    n3471_lo_p
  );


  buf

  (
    n3459_lo_p_spl_,
    n3459_lo_p
  );


  buf

  (
    n3447_lo_p_spl_,
    n3447_lo_p
  );


  buf

  (
    n3435_lo_p_spl_,
    n3435_lo_p
  );


  buf

  (
    n3423_lo_p_spl_,
    n3423_lo_p
  );


  buf

  (
    g1271_p_spl_,
    g1271_p
  );


  buf

  (
    n4659_lo_n_spl_,
    n4659_lo_n
  );


  buf

  (
    n4647_lo_n_spl_,
    n4647_lo_n
  );


  buf

  (
    n7463_o2_p_spl_,
    n7463_o2_p
  );


  buf

  (
    n3339_lo_p_spl_,
    n3339_lo_p
  );


  buf

  (
    n3339_lo_n_spl_,
    n3339_lo_n
  );


  buf

  (
    g2078_n_spl_,
    g2078_n
  );


  buf

  (
    g2078_p_spl_,
    g2078_p
  );


  buf

  (
    g2081_n_spl_,
    g2081_n
  );


  buf

  (
    n4659_lo_p_spl_,
    n4659_lo_p
  );


  buf

  (
    n3255_lo_p_spl_,
    n3255_lo_p
  );


  buf

  (
    n4647_lo_p_spl_,
    n4647_lo_p
  );


  buf

  (
    g1601_p_spl_,
    g1601_p
  );


  buf

  (
    g2092_n_spl_,
    g2092_n
  );


  buf

  (
    n4467_lo_n_spl_,
    n4467_lo_n
  );


  buf

  (
    n4443_lo_n_spl_,
    n4443_lo_n
  );


  buf

  (
    g1765_n_spl_,
    g1765_n
  );


  buf

  (
    n4479_lo_n_spl_,
    n4479_lo_n
  );


  buf

  (
    g1790_n_spl_,
    g1790_n
  );


  buf

  (
    g1449_n_spl_,
    g1449_n
  );


  buf

  (
    g1474_n_spl_,
    g1474_n
  );


  buf

  (
    n3795_lo_n_spl_,
    n3795_lo_n
  );


  buf

  (
    n7156_o2_n_spl_,
    n7156_o2_n
  );


  buf

  (
    n7156_o2_p_spl_,
    n7156_o2_p
  );


  buf

  (
    g2103_n_spl_,
    g2103_n
  );


  buf

  (
    g2103_n_spl_0,
    g2103_n_spl_
  );


  buf

  (
    g2103_n_spl_00,
    g2103_n_spl_0
  );


  buf

  (
    g2103_n_spl_1,
    g2103_n_spl_
  );


  buf

  (
    g2154_n_spl_,
    g2154_n
  );


  buf

  (
    g2154_n_spl_0,
    g2154_n_spl_
  );


  buf

  (
    g2154_n_spl_00,
    g2154_n_spl_0
  );


  buf

  (
    g2154_n_spl_1,
    g2154_n_spl_
  );


  buf

  (
    n3111_lo_p_spl_,
    n3111_lo_p
  );


  buf

  (
    n3099_lo_p_spl_,
    n3099_lo_p
  );


  buf

  (
    g2111_n_spl_,
    g2111_n
  );


  buf

  (
    g2111_n_spl_0,
    g2111_n_spl_
  );


  buf

  (
    g2111_n_spl_00,
    g2111_n_spl_0
  );


  buf

  (
    g2111_n_spl_1,
    g2111_n_spl_
  );


  buf

  (
    g2162_n_spl_,
    g2162_n
  );


  buf

  (
    g2162_n_spl_0,
    g2162_n_spl_
  );


  buf

  (
    g2162_n_spl_00,
    g2162_n_spl_0
  );


  buf

  (
    g2162_n_spl_1,
    g2162_n_spl_
  );


  buf

  (
    n2811_lo_p_spl_,
    n2811_lo_p
  );


  buf

  (
    n2823_lo_p_spl_,
    n2823_lo_p
  );


  buf

  (
    g2119_n_spl_,
    g2119_n
  );


  buf

  (
    g2119_n_spl_0,
    g2119_n_spl_
  );


  buf

  (
    g2119_n_spl_00,
    g2119_n_spl_0
  );


  buf

  (
    g2119_n_spl_1,
    g2119_n_spl_
  );


  buf

  (
    g2170_n_spl_,
    g2170_n
  );


  buf

  (
    g2170_n_spl_0,
    g2170_n_spl_
  );


  buf

  (
    g2170_n_spl_00,
    g2170_n_spl_0
  );


  buf

  (
    g2170_n_spl_1,
    g2170_n_spl_
  );


  buf

  (
    n3075_lo_p_spl_,
    n3075_lo_p
  );


  buf

  (
    n3087_lo_p_spl_,
    n3087_lo_p
  );


  buf

  (
    g2127_n_spl_,
    g2127_n
  );


  buf

  (
    g2127_n_spl_0,
    g2127_n_spl_
  );


  buf

  (
    g2127_n_spl_00,
    g2127_n_spl_0
  );


  buf

  (
    g2127_n_spl_1,
    g2127_n_spl_
  );


  buf

  (
    g2178_n_spl_,
    g2178_n
  );


  buf

  (
    g2178_n_spl_0,
    g2178_n_spl_
  );


  buf

  (
    g2178_n_spl_00,
    g2178_n_spl_0
  );


  buf

  (
    g2178_n_spl_1,
    g2178_n_spl_
  );


  buf

  (
    n3039_lo_p_spl_,
    n3039_lo_p
  );


  buf

  (
    n2787_lo_p_spl_,
    n2787_lo_p
  );


  buf

  (
    n3651_lo_p_spl_,
    n3651_lo_p
  );


  buf

  (
    n3531_lo_p_spl_,
    n3531_lo_p
  );


  buf

  (
    n3627_lo_p_spl_,
    n3627_lo_p
  );


  buf

  (
    n3507_lo_p_spl_,
    n3507_lo_p
  );


  buf

  (
    n3615_lo_p_spl_,
    n3615_lo_p
  );


  buf

  (
    n3495_lo_p_spl_,
    n3495_lo_p
  );


  buf

  (
    n3603_lo_p_spl_,
    n3603_lo_p
  );


  buf

  (
    n3483_lo_p_spl_,
    n3483_lo_p
  );


  buf

  (
    g2365_n_spl_,
    g2365_n
  );


  buf

  (
    g2370_p_spl_,
    g2370_p
  );


  buf

  (
    g2375_n_spl_,
    g2375_n
  );


  buf

  (
    g2381_n_spl_,
    g2381_n
  );


  buf

  (
    g2386_p_spl_,
    g2386_p
  );


  buf

  (
    g2399_n_spl_,
    g2399_n
  );


  buf

  (
    g2399_n_spl_0,
    g2399_n_spl_
  );


  buf

  (
    g2399_n_spl_1,
    g2399_n_spl_
  );


  buf

  (
    g2407_n_spl_,
    g2407_n
  );


  buf

  (
    g2407_n_spl_0,
    g2407_n_spl_
  );


  buf

  (
    g2407_n_spl_1,
    g2407_n_spl_
  );


  buf

  (
    n2655_lo_p_spl_,
    n2655_lo_p
  );


  buf

  (
    n2883_lo_p_spl_,
    n2883_lo_p
  );


  buf

  (
    n3543_lo_p_spl_,
    n3543_lo_p
  );


  buf

  (
    n3555_lo_p_spl_,
    n3555_lo_p
  );


  buf

  (
    n2968_inv_n_spl_,
    n2968_inv_n
  );


  buf

  (
    n2968_inv_n_spl_0,
    n2968_inv_n_spl_
  );


  buf

  (
    n2968_inv_n_spl_00,
    n2968_inv_n_spl_0
  );


  buf

  (
    n2968_inv_n_spl_01,
    n2968_inv_n_spl_0
  );


  buf

  (
    n2968_inv_n_spl_1,
    n2968_inv_n_spl_
  );


  buf

  (
    n2968_inv_n_spl_10,
    n2968_inv_n_spl_1
  );


  buf

  (
    n2968_inv_n_spl_11,
    n2968_inv_n_spl_1
  );


  buf

  (
    n4308_lo_buf_o2_p_spl_,
    n4308_lo_buf_o2_p
  );


  buf

  (
    n4308_lo_buf_o2_p_spl_0,
    n4308_lo_buf_o2_p_spl_
  );


  buf

  (
    n4308_lo_buf_o2_p_spl_00,
    n4308_lo_buf_o2_p_spl_0
  );


  buf

  (
    n4308_lo_buf_o2_p_spl_1,
    n4308_lo_buf_o2_p_spl_
  );


  buf

  (
    n2968_inv_p_spl_,
    n2968_inv_p
  );


  buf

  (
    n2968_inv_p_spl_0,
    n2968_inv_p_spl_
  );


  buf

  (
    n2968_inv_p_spl_00,
    n2968_inv_p_spl_0
  );


  buf

  (
    n2968_inv_p_spl_000,
    n2968_inv_p_spl_00
  );


  buf

  (
    n2968_inv_p_spl_01,
    n2968_inv_p_spl_0
  );


  buf

  (
    n2968_inv_p_spl_1,
    n2968_inv_p_spl_
  );


  buf

  (
    n2968_inv_p_spl_10,
    n2968_inv_p_spl_1
  );


  buf

  (
    n2968_inv_p_spl_11,
    n2968_inv_p_spl_1
  );


  buf

  (
    n4308_lo_buf_o2_n_spl_,
    n4308_lo_buf_o2_n
  );


  buf

  (
    n4308_lo_buf_o2_n_spl_0,
    n4308_lo_buf_o2_n_spl_
  );


  buf

  (
    n4308_lo_buf_o2_n_spl_1,
    n4308_lo_buf_o2_n_spl_
  );


  buf

  (
    n2974_inv_n_spl_,
    n2974_inv_n
  );


  buf

  (
    n2974_inv_n_spl_0,
    n2974_inv_n_spl_
  );


  buf

  (
    n2974_inv_n_spl_00,
    n2974_inv_n_spl_0
  );


  buf

  (
    n2974_inv_n_spl_01,
    n2974_inv_n_spl_0
  );


  buf

  (
    n2974_inv_n_spl_1,
    n2974_inv_n_spl_
  );


  buf

  (
    n2974_inv_n_spl_10,
    n2974_inv_n_spl_1
  );


  buf

  (
    n2974_inv_p_spl_,
    n2974_inv_p
  );


  buf

  (
    n2974_inv_p_spl_0,
    n2974_inv_p_spl_
  );


  buf

  (
    n2974_inv_p_spl_00,
    n2974_inv_p_spl_0
  );


  buf

  (
    n2974_inv_p_spl_01,
    n2974_inv_p_spl_0
  );


  buf

  (
    n2974_inv_p_spl_1,
    n2974_inv_p_spl_
  );


  buf

  (
    n2974_inv_p_spl_10,
    n2974_inv_p_spl_1
  );


  buf

  (
    n2974_inv_p_spl_11,
    n2974_inv_p_spl_1
  );


  buf

  (
    n3121_inv_n_spl_,
    n3121_inv_n
  );


  buf

  (
    n3121_inv_n_spl_0,
    n3121_inv_n_spl_
  );


  buf

  (
    n3121_inv_n_spl_00,
    n3121_inv_n_spl_0
  );


  buf

  (
    n3121_inv_n_spl_01,
    n3121_inv_n_spl_0
  );


  buf

  (
    n3121_inv_n_spl_1,
    n3121_inv_n_spl_
  );


  buf

  (
    n3121_inv_n_spl_10,
    n3121_inv_n_spl_1
  );


  buf

  (
    n3121_inv_n_spl_11,
    n3121_inv_n_spl_1
  );


  buf

  (
    G1873_o2_p_spl_,
    G1873_o2_p
  );


  buf

  (
    n3121_inv_p_spl_,
    n3121_inv_p
  );


  buf

  (
    n3121_inv_p_spl_0,
    n3121_inv_p_spl_
  );


  buf

  (
    n3121_inv_p_spl_00,
    n3121_inv_p_spl_0
  );


  buf

  (
    n3121_inv_p_spl_000,
    n3121_inv_p_spl_00
  );


  buf

  (
    n3121_inv_p_spl_01,
    n3121_inv_p_spl_0
  );


  buf

  (
    n3121_inv_p_spl_1,
    n3121_inv_p_spl_
  );


  buf

  (
    n3121_inv_p_spl_10,
    n3121_inv_p_spl_1
  );


  buf

  (
    n3121_inv_p_spl_11,
    n3121_inv_p_spl_1
  );


  buf

  (
    G1873_o2_n_spl_,
    G1873_o2_n
  );


  buf

  (
    n3124_inv_n_spl_,
    n3124_inv_n
  );


  buf

  (
    n3124_inv_n_spl_0,
    n3124_inv_n_spl_
  );


  buf

  (
    n3124_inv_n_spl_00,
    n3124_inv_n_spl_0
  );


  buf

  (
    n3124_inv_n_spl_01,
    n3124_inv_n_spl_0
  );


  buf

  (
    n3124_inv_n_spl_1,
    n3124_inv_n_spl_
  );


  buf

  (
    n3124_inv_n_spl_10,
    n3124_inv_n_spl_1
  );


  buf

  (
    n3124_inv_p_spl_,
    n3124_inv_p
  );


  buf

  (
    n3124_inv_p_spl_0,
    n3124_inv_p_spl_
  );


  buf

  (
    n3124_inv_p_spl_00,
    n3124_inv_p_spl_0
  );


  buf

  (
    n3124_inv_p_spl_01,
    n3124_inv_p_spl_0
  );


  buf

  (
    n3124_inv_p_spl_1,
    n3124_inv_p_spl_
  );


  buf

  (
    n3124_inv_p_spl_10,
    n3124_inv_p_spl_1
  );


  buf

  (
    n3124_inv_p_spl_11,
    n3124_inv_p_spl_1
  );


  buf

  (
    n6955_o2_p_spl_,
    n6955_o2_p
  );


  buf

  (
    n6955_o2_n_spl_,
    n6955_o2_n
  );


  buf

  (
    n6954_o2_p_spl_,
    n6954_o2_p
  );


  buf

  (
    n6954_o2_p_spl_0,
    n6954_o2_p_spl_
  );


  buf

  (
    n6954_o2_p_spl_00,
    n6954_o2_p_spl_0
  );


  buf

  (
    n6954_o2_p_spl_01,
    n6954_o2_p_spl_0
  );


  buf

  (
    n6954_o2_p_spl_1,
    n6954_o2_p_spl_
  );


  buf

  (
    n6954_o2_p_spl_10,
    n6954_o2_p_spl_1
  );


  buf

  (
    n6954_o2_n_spl_,
    n6954_o2_n
  );


  buf

  (
    n6954_o2_n_spl_0,
    n6954_o2_n_spl_
  );


  buf

  (
    n6954_o2_n_spl_00,
    n6954_o2_n_spl_0
  );


  buf

  (
    n6954_o2_n_spl_01,
    n6954_o2_n_spl_0
  );


  buf

  (
    n6954_o2_n_spl_1,
    n6954_o2_n_spl_
  );


  buf

  (
    n6954_o2_n_spl_10,
    n6954_o2_n_spl_1
  );


  buf

  (
    n7387_o2_p_spl_,
    n7387_o2_p
  );


  buf

  (
    n7387_o2_p_spl_0,
    n7387_o2_p_spl_
  );


  buf

  (
    n7387_o2_p_spl_00,
    n7387_o2_p_spl_0
  );


  buf

  (
    n7387_o2_p_spl_01,
    n7387_o2_p_spl_0
  );


  buf

  (
    n7387_o2_p_spl_1,
    n7387_o2_p_spl_
  );


  buf

  (
    n7387_o2_n_spl_,
    n7387_o2_n
  );


  buf

  (
    n7387_o2_n_spl_0,
    n7387_o2_n_spl_
  );


  buf

  (
    n7387_o2_n_spl_00,
    n7387_o2_n_spl_0
  );


  buf

  (
    n7387_o2_n_spl_01,
    n7387_o2_n_spl_0
  );


  buf

  (
    n7387_o2_n_spl_1,
    n7387_o2_n_spl_
  );


  buf

  (
    G3495_o2_p_spl_,
    G3495_o2_p
  );


  buf

  (
    G3495_o2_p_spl_0,
    G3495_o2_p_spl_
  );


  buf

  (
    G3495_o2_p_spl_00,
    G3495_o2_p_spl_0
  );


  buf

  (
    G3495_o2_p_spl_1,
    G3495_o2_p_spl_
  );


  buf

  (
    G3495_o2_n_spl_,
    G3495_o2_n
  );


  buf

  (
    G3495_o2_n_spl_0,
    G3495_o2_n_spl_
  );


  buf

  (
    G3495_o2_n_spl_00,
    G3495_o2_n_spl_0
  );


  buf

  (
    G3495_o2_n_spl_1,
    G3495_o2_n_spl_
  );


  buf

  (
    n6957_o2_p_spl_,
    n6957_o2_p
  );


  buf

  (
    n6957_o2_n_spl_,
    n6957_o2_n
  );


  buf

  (
    n6956_o2_p_spl_,
    n6956_o2_p
  );


  buf

  (
    n6956_o2_p_spl_0,
    n6956_o2_p_spl_
  );


  buf

  (
    n6956_o2_p_spl_00,
    n6956_o2_p_spl_0
  );


  buf

  (
    n6956_o2_p_spl_01,
    n6956_o2_p_spl_0
  );


  buf

  (
    n6956_o2_p_spl_1,
    n6956_o2_p_spl_
  );


  buf

  (
    n6956_o2_p_spl_10,
    n6956_o2_p_spl_1
  );


  buf

  (
    n6956_o2_n_spl_,
    n6956_o2_n
  );


  buf

  (
    n6956_o2_n_spl_0,
    n6956_o2_n_spl_
  );


  buf

  (
    n6956_o2_n_spl_00,
    n6956_o2_n_spl_0
  );


  buf

  (
    n6956_o2_n_spl_01,
    n6956_o2_n_spl_0
  );


  buf

  (
    n6956_o2_n_spl_1,
    n6956_o2_n_spl_
  );


  buf

  (
    n6956_o2_n_spl_10,
    n6956_o2_n_spl_1
  );


  buf

  (
    n7386_o2_p_spl_,
    n7386_o2_p
  );


  buf

  (
    n7386_o2_p_spl_0,
    n7386_o2_p_spl_
  );


  buf

  (
    n7386_o2_p_spl_00,
    n7386_o2_p_spl_0
  );


  buf

  (
    n7386_o2_p_spl_01,
    n7386_o2_p_spl_0
  );


  buf

  (
    n7386_o2_p_spl_1,
    n7386_o2_p_spl_
  );


  buf

  (
    n7386_o2_n_spl_,
    n7386_o2_n
  );


  buf

  (
    n7386_o2_n_spl_0,
    n7386_o2_n_spl_
  );


  buf

  (
    n7386_o2_n_spl_00,
    n7386_o2_n_spl_0
  );


  buf

  (
    n7386_o2_n_spl_01,
    n7386_o2_n_spl_0
  );


  buf

  (
    n7386_o2_n_spl_1,
    n7386_o2_n_spl_
  );


  buf

  (
    G3621_o2_p_spl_,
    G3621_o2_p
  );


  buf

  (
    G3621_o2_p_spl_0,
    G3621_o2_p_spl_
  );


  buf

  (
    G3621_o2_p_spl_00,
    G3621_o2_p_spl_0
  );


  buf

  (
    G3621_o2_p_spl_1,
    G3621_o2_p_spl_
  );


  buf

  (
    G3621_o2_n_spl_,
    G3621_o2_n
  );


  buf

  (
    G3621_o2_n_spl_0,
    G3621_o2_n_spl_
  );


  buf

  (
    G3621_o2_n_spl_00,
    G3621_o2_n_spl_0
  );


  buf

  (
    G3621_o2_n_spl_1,
    G3621_o2_n_spl_
  );


  buf

  (
    G2404_o2_p_spl_,
    G2404_o2_p
  );


  buf

  (
    G2404_o2_p_spl_0,
    G2404_o2_p_spl_
  );


  buf

  (
    G2404_o2_p_spl_1,
    G2404_o2_p_spl_
  );


  buf

  (
    n4296_lo_buf_o2_p_spl_,
    n4296_lo_buf_o2_p
  );


  buf

  (
    n4296_lo_buf_o2_p_spl_0,
    n4296_lo_buf_o2_p_spl_
  );


  buf

  (
    n4296_lo_buf_o2_p_spl_1,
    n4296_lo_buf_o2_p_spl_
  );


  buf

  (
    G2404_o2_n_spl_,
    G2404_o2_n
  );


  buf

  (
    G2404_o2_n_spl_0,
    G2404_o2_n_spl_
  );


  buf

  (
    n4296_lo_buf_o2_n_spl_,
    n4296_lo_buf_o2_n
  );


  buf

  (
    n4296_lo_buf_o2_n_spl_0,
    n4296_lo_buf_o2_n_spl_
  );


  buf

  (
    G2466_o2_p_spl_,
    G2466_o2_p
  );


  buf

  (
    G2466_o2_p_spl_0,
    G2466_o2_p_spl_
  );


  buf

  (
    G2466_o2_p_spl_1,
    G2466_o2_p_spl_
  );


  buf

  (
    n4368_lo_buf_o2_p_spl_,
    n4368_lo_buf_o2_p
  );


  buf

  (
    n4368_lo_buf_o2_p_spl_0,
    n4368_lo_buf_o2_p_spl_
  );


  buf

  (
    n4368_lo_buf_o2_p_spl_1,
    n4368_lo_buf_o2_p_spl_
  );


  buf

  (
    G2466_o2_n_spl_,
    G2466_o2_n
  );


  buf

  (
    G2466_o2_n_spl_0,
    G2466_o2_n_spl_
  );


  buf

  (
    n4368_lo_buf_o2_n_spl_,
    n4368_lo_buf_o2_n
  );


  buf

  (
    n4368_lo_buf_o2_n_spl_0,
    n4368_lo_buf_o2_n_spl_
  );


  buf

  (
    n6772_o2_n_spl_,
    n6772_o2_n
  );


  buf

  (
    n6772_o2_n_spl_0,
    n6772_o2_n_spl_
  );


  buf

  (
    n6772_o2_p_spl_,
    n6772_o2_p
  );


  buf

  (
    n6772_o2_p_spl_0,
    n6772_o2_p_spl_
  );


  buf

  (
    n6772_o2_p_spl_1,
    n6772_o2_p_spl_
  );


  buf

  (
    G2424_o2_p_spl_,
    G2424_o2_p
  );


  buf

  (
    n4320_lo_buf_o2_p_spl_,
    n4320_lo_buf_o2_p
  );


  buf

  (
    G1821_o2_p_spl_,
    G1821_o2_p
  );


  buf

  (
    n4053_lo_p_spl_,
    n4053_lo_p
  );


  buf

  (
    n4053_lo_p_spl_0,
    n4053_lo_p_spl_
  );


  buf

  (
    n4053_lo_p_spl_00,
    n4053_lo_p_spl_0
  );


  buf

  (
    n4053_lo_p_spl_1,
    n4053_lo_p_spl_
  );


  buf

  (
    n4053_lo_n_spl_,
    n4053_lo_n
  );


  buf

  (
    G1060_o2_n_spl_,
    G1060_o2_n
  );


  buf

  (
    G1734_o2_p_spl_,
    G1734_o2_p
  );


  buf

  (
    n3753_lo_p_spl_,
    n3753_lo_p
  );


  buf

  (
    n3753_lo_p_spl_0,
    n3753_lo_p_spl_
  );


  buf

  (
    n3753_lo_p_spl_00,
    n3753_lo_p_spl_0
  );


  buf

  (
    n3753_lo_p_spl_1,
    n3753_lo_p_spl_
  );


  buf

  (
    n3753_lo_n_spl_,
    n3753_lo_n
  );


  buf

  (
    G963_o2_n_spl_,
    G963_o2_n
  );


  buf

  (
    n4164_lo_buf_o2_p_spl_,
    n4164_lo_buf_o2_p
  );


  buf

  (
    G1815_o2_p_spl_,
    G1815_o2_p
  );


  buf

  (
    G1815_o2_p_spl_0,
    G1815_o2_p_spl_
  );


  buf

  (
    G1815_o2_n_spl_,
    G1815_o2_n
  );


  buf

  (
    n4176_lo_buf_o2_p_spl_,
    n4176_lo_buf_o2_p
  );


  buf

  (
    n2662_inv_n_spl_,
    n2662_inv_n
  );


  buf

  (
    n2662_inv_p_spl_,
    n2662_inv_p
  );


  buf

  (
    n2662_inv_p_spl_0,
    n2662_inv_p_spl_
  );


  buf

  (
    n7136_o2_p_spl_,
    n7136_o2_p
  );


  buf

  (
    n7136_o2_p_spl_0,
    n7136_o2_p_spl_
  );


  buf

  (
    n7136_o2_p_spl_1,
    n7136_o2_p_spl_
  );


  buf

  (
    n7132_o2_p_spl_,
    n7132_o2_p
  );


  buf

  (
    n7132_o2_p_spl_0,
    n7132_o2_p_spl_
  );


  buf

  (
    n7132_o2_p_spl_00,
    n7132_o2_p_spl_0
  );


  buf

  (
    n7132_o2_p_spl_01,
    n7132_o2_p_spl_0
  );


  buf

  (
    n7132_o2_p_spl_1,
    n7132_o2_p_spl_
  );


  buf

  (
    n7132_o2_p_spl_10,
    n7132_o2_p_spl_1
  );


  buf

  (
    n7023_o2_p_spl_,
    n7023_o2_p
  );


  buf

  (
    n7023_o2_p_spl_0,
    n7023_o2_p_spl_
  );


  buf

  (
    n7016_o2_p_spl_,
    n7016_o2_p
  );


  buf

  (
    n7016_o2_p_spl_0,
    n7016_o2_p_spl_
  );


  buf

  (
    n7016_o2_p_spl_00,
    n7016_o2_p_spl_0
  );


  buf

  (
    n7016_o2_p_spl_01,
    n7016_o2_p_spl_0
  );


  buf

  (
    n7016_o2_p_spl_1,
    n7016_o2_p_spl_
  );


  buf

  (
    n7022_o2_n_spl_,
    n7022_o2_n
  );


  buf

  (
    n7022_o2_n_spl_0,
    n7022_o2_n_spl_
  );


  buf

  (
    n7017_o2_n_spl_,
    n7017_o2_n
  );


  buf

  (
    n7017_o2_n_spl_0,
    n7017_o2_n_spl_
  );


  buf

  (
    n7017_o2_n_spl_00,
    n7017_o2_n_spl_0
  );


  buf

  (
    n7017_o2_n_spl_01,
    n7017_o2_n_spl_0
  );


  buf

  (
    n7017_o2_n_spl_1,
    n7017_o2_n_spl_
  );


  buf

  (
    n7135_o2_n_spl_,
    n7135_o2_n
  );


  buf

  (
    n7133_o2_n_spl_,
    n7133_o2_n
  );


  buf

  (
    n7133_o2_n_spl_0,
    n7133_o2_n_spl_
  );


  buf

  (
    n7133_o2_n_spl_00,
    n7133_o2_n_spl_0
  );


  buf

  (
    n7133_o2_n_spl_1,
    n7133_o2_n_spl_
  );


  buf

  (
    n4272_lo_buf_o2_p_spl_,
    n4272_lo_buf_o2_p
  );


  buf

  (
    G2386_o2_p_spl_,
    G2386_o2_p
  );


  buf

  (
    n4404_lo_buf_o2_p_spl_,
    n4404_lo_buf_o2_p
  );


  buf

  (
    G2454_o2_p_spl_,
    G2454_o2_p
  );


  buf

  (
    n7384_o2_p_spl_,
    n7384_o2_p
  );


  buf

  (
    n7384_o2_p_spl_0,
    n7384_o2_p_spl_
  );


  buf

  (
    n7383_o2_n_spl_,
    n7383_o2_n
  );


  buf

  (
    n7383_o2_n_spl_0,
    n7383_o2_n_spl_
  );


  buf

  (
    n7383_o2_n_spl_1,
    n7383_o2_n_spl_
  );


  buf

  (
    n7384_o2_n_spl_,
    n7384_o2_n
  );


  buf

  (
    n7383_o2_p_spl_,
    n7383_o2_p
  );


  buf

  (
    n7383_o2_p_spl_0,
    n7383_o2_p_spl_
  );


  buf

  (
    n7383_o2_p_spl_00,
    n7383_o2_p_spl_0
  );


  buf

  (
    n7383_o2_p_spl_01,
    n7383_o2_p_spl_0
  );


  buf

  (
    n7383_o2_p_spl_1,
    n7383_o2_p_spl_
  );


  buf

  (
    n7016_o2_n_spl_,
    n7016_o2_n
  );


  buf

  (
    n7016_o2_n_spl_0,
    n7016_o2_n_spl_
  );


  buf

  (
    n7016_o2_n_spl_1,
    n7016_o2_n_spl_
  );


  buf

  (
    n7023_o2_n_spl_,
    n7023_o2_n
  );


  buf

  (
    n7022_o2_p_spl_,
    n7022_o2_p
  );


  buf

  (
    n7022_o2_p_spl_0,
    n7022_o2_p_spl_
  );


  buf

  (
    n7022_o2_p_spl_1,
    n7022_o2_p_spl_
  );


  buf

  (
    n7017_o2_p_spl_,
    n7017_o2_p
  );


  buf

  (
    n7017_o2_p_spl_0,
    n7017_o2_p_spl_
  );


  buf

  (
    n7017_o2_p_spl_00,
    n7017_o2_p_spl_0
  );


  buf

  (
    n7017_o2_p_spl_01,
    n7017_o2_p_spl_0
  );


  buf

  (
    n7017_o2_p_spl_1,
    n7017_o2_p_spl_
  );


  buf

  (
    n4224_lo_buf_o2_p_spl_,
    n4224_lo_buf_o2_p
  );


  buf

  (
    n4224_lo_buf_o2_p_spl_0,
    n4224_lo_buf_o2_p_spl_
  );


  buf

  (
    n4224_lo_buf_o2_p_spl_00,
    n4224_lo_buf_o2_p_spl_0
  );


  buf

  (
    n4224_lo_buf_o2_p_spl_1,
    n4224_lo_buf_o2_p_spl_
  );


  buf

  (
    G2379_o2_p_spl_,
    G2379_o2_p
  );


  buf

  (
    G2379_o2_p_spl_0,
    G2379_o2_p_spl_
  );


  buf

  (
    G2379_o2_p_spl_00,
    G2379_o2_p_spl_0
  );


  buf

  (
    G2379_o2_p_spl_1,
    G2379_o2_p_spl_
  );


  buf

  (
    n4224_lo_buf_o2_n_spl_,
    n4224_lo_buf_o2_n
  );


  buf

  (
    n4224_lo_buf_o2_n_spl_0,
    n4224_lo_buf_o2_n_spl_
  );


  buf

  (
    n4224_lo_buf_o2_n_spl_1,
    n4224_lo_buf_o2_n_spl_
  );


  buf

  (
    G2379_o2_n_spl_,
    G2379_o2_n
  );


  buf

  (
    G2379_o2_n_spl_0,
    G2379_o2_n_spl_
  );


  buf

  (
    G2379_o2_n_spl_1,
    G2379_o2_n_spl_
  );


  buf

  (
    G1356_o2_p_spl_,
    G1356_o2_p
  );


  buf

  (
    G2933_o2_n_spl_,
    G2933_o2_n
  );


  buf

  (
    G1356_o2_n_spl_,
    G1356_o2_n
  );


  buf

  (
    G2933_o2_p_spl_,
    G2933_o2_p
  );


  buf

  (
    G1359_o2_p_spl_,
    G1359_o2_p
  );


  buf

  (
    G2936_o2_n_spl_,
    G2936_o2_n
  );


  buf

  (
    G1359_o2_n_spl_,
    G1359_o2_n
  );


  buf

  (
    G2936_o2_p_spl_,
    G2936_o2_p
  );


  buf

  (
    G1398_o2_p_spl_,
    G1398_o2_p
  );


  buf

  (
    G2975_o2_n_spl_,
    G2975_o2_n
  );


  buf

  (
    G1398_o2_n_spl_,
    G1398_o2_n
  );


  buf

  (
    G2975_o2_p_spl_,
    G2975_o2_p
  );


  buf

  (
    G1401_o2_p_spl_,
    G1401_o2_p
  );


  buf

  (
    G2978_o2_n_spl_,
    G2978_o2_n
  );


  buf

  (
    G1401_o2_n_spl_,
    G1401_o2_n
  );


  buf

  (
    G2978_o2_p_spl_,
    G2978_o2_p
  );


  buf

  (
    n4260_lo_buf_o2_p_spl_,
    n4260_lo_buf_o2_p
  );


  buf

  (
    G2392_o2_p_spl_,
    G2392_o2_p
  );


  buf

  (
    n4392_lo_buf_o2_p_spl_,
    n4392_lo_buf_o2_p
  );


  buf

  (
    G2460_o2_p_spl_,
    G2460_o2_p
  );


  buf

  (
    n4098_lo_p_spl_,
    n4098_lo_p
  );


  buf

  (
    G1728_o2_p_spl_,
    G1728_o2_p
  );


  buf

  (
    n3834_lo_p_spl_,
    n3834_lo_p
  );


  buf

  (
    n2665_inv_p_spl_,
    n2665_inv_p
  );


  buf

  (
    n4080_lo_buf_o2_p_spl_,
    n4080_lo_buf_o2_p
  );


  buf

  (
    n4080_lo_buf_o2_p_spl_0,
    n4080_lo_buf_o2_p_spl_
  );


  buf

  (
    n4080_lo_buf_o2_p_spl_00,
    n4080_lo_buf_o2_p_spl_0
  );


  buf

  (
    n4080_lo_buf_o2_p_spl_01,
    n4080_lo_buf_o2_p_spl_0
  );


  buf

  (
    n4080_lo_buf_o2_p_spl_1,
    n4080_lo_buf_o2_p_spl_
  );


  buf

  (
    n4080_lo_buf_o2_p_spl_10,
    n4080_lo_buf_o2_p_spl_1
  );


  buf

  (
    n4002_lo_p_spl_,
    n4002_lo_p
  );


  buf

  (
    n4080_lo_buf_o2_n_spl_,
    n4080_lo_buf_o2_n
  );


  buf

  (
    n4080_lo_buf_o2_n_spl_0,
    n4080_lo_buf_o2_n_spl_
  );


  buf

  (
    n4080_lo_buf_o2_n_spl_00,
    n4080_lo_buf_o2_n_spl_0
  );


  buf

  (
    n4080_lo_buf_o2_n_spl_1,
    n4080_lo_buf_o2_n_spl_
  );


  buf

  (
    n4092_lo_buf_o2_p_spl_,
    n4092_lo_buf_o2_p
  );


  buf

  (
    n4092_lo_buf_o2_p_spl_0,
    n4092_lo_buf_o2_p_spl_
  );


  buf

  (
    n4092_lo_buf_o2_p_spl_00,
    n4092_lo_buf_o2_p_spl_0
  );


  buf

  (
    n4092_lo_buf_o2_p_spl_01,
    n4092_lo_buf_o2_p_spl_0
  );


  buf

  (
    n4092_lo_buf_o2_p_spl_1,
    n4092_lo_buf_o2_p_spl_
  );


  buf

  (
    n4092_lo_buf_o2_p_spl_10,
    n4092_lo_buf_o2_p_spl_1
  );


  buf

  (
    n3702_lo_p_spl_,
    n3702_lo_p
  );


  buf

  (
    n4092_lo_buf_o2_n_spl_,
    n4092_lo_buf_o2_n
  );


  buf

  (
    n4092_lo_buf_o2_n_spl_0,
    n4092_lo_buf_o2_n_spl_
  );


  buf

  (
    n4092_lo_buf_o2_n_spl_00,
    n4092_lo_buf_o2_n_spl_0
  );


  buf

  (
    n4092_lo_buf_o2_n_spl_1,
    n4092_lo_buf_o2_n_spl_
  );


  buf

  (
    g2565_p_spl_,
    g2565_p
  );


  buf

  (
    g2452_p_spl_,
    g2452_p
  );


  buf

  (
    g2452_p_spl_0,
    g2452_p_spl_
  );


  buf

  (
    g2452_p_spl_1,
    g2452_p_spl_
  );


  buf

  (
    g2565_n_spl_,
    g2565_n
  );


  buf

  (
    g2452_n_spl_,
    g2452_n
  );


  buf

  (
    g2452_n_spl_0,
    g2452_n_spl_
  );


  buf

  (
    g2452_n_spl_00,
    g2452_n_spl_0
  );


  buf

  (
    g2452_n_spl_1,
    g2452_n_spl_
  );


  buf

  (
    G3474_o2_p_spl_,
    G3474_o2_p
  );


  buf

  (
    G3474_o2_p_spl_0,
    G3474_o2_p_spl_
  );


  buf

  (
    G3474_o2_n_spl_,
    G3474_o2_n
  );


  buf

  (
    g2571_p_spl_,
    g2571_p
  );


  buf

  (
    g2485_n_spl_,
    g2485_n
  );


  buf

  (
    g2485_n_spl_0,
    g2485_n_spl_
  );


  buf

  (
    n4488_lo_p_spl_,
    n4488_lo_p
  );


  buf

  (
    n4488_lo_p_spl_0,
    n4488_lo_p_spl_
  );


  buf

  (
    g2576_p_spl_,
    g2576_p
  );


  buf

  (
    g2576_n_spl_,
    g2576_n
  );


  buf

  (
    g2582_p_spl_,
    g2582_p
  );


  buf

  (
    g2485_p_spl_,
    g2485_p
  );


  buf

  (
    g2466_p_spl_,
    g2466_p
  );


  buf

  (
    n4488_lo_n_spl_,
    n4488_lo_n
  );


  buf

  (
    n4488_lo_n_spl_0,
    n4488_lo_n_spl_
  );


  buf

  (
    g2593_p_spl_,
    g2593_p
  );


  buf

  (
    g2593_n_spl_,
    g2593_n
  );


  buf

  (
    g2603_p_spl_,
    g2603_p
  );


  buf

  (
    g2603_n_spl_,
    g2603_n
  );


  buf

  (
    g2614_p_spl_,
    g2614_p
  );


  buf

  (
    G2492_o2_p_spl_,
    G2492_o2_p
  );


  buf

  (
    G2492_o2_p_spl_0,
    G2492_o2_p_spl_
  );


  buf

  (
    G2492_o2_p_spl_00,
    G2492_o2_p_spl_0
  );


  buf

  (
    G2492_o2_p_spl_000,
    G2492_o2_p_spl_00
  );


  buf

  (
    G2492_o2_p_spl_001,
    G2492_o2_p_spl_00
  );


  buf

  (
    G2492_o2_p_spl_01,
    G2492_o2_p_spl_0
  );


  buf

  (
    G2492_o2_p_spl_1,
    G2492_o2_p_spl_
  );


  buf

  (
    G2492_o2_p_spl_10,
    G2492_o2_p_spl_1
  );


  buf

  (
    G2492_o2_p_spl_11,
    G2492_o2_p_spl_1
  );


  buf

  (
    g2614_n_spl_,
    g2614_n
  );


  buf

  (
    G2492_o2_n_spl_,
    G2492_o2_n
  );


  buf

  (
    G2492_o2_n_spl_0,
    G2492_o2_n_spl_
  );


  buf

  (
    G2492_o2_n_spl_1,
    G2492_o2_n_spl_
  );


  buf

  (
    n2341_inv_p_spl_,
    n2341_inv_p
  );


  buf

  (
    n2341_inv_p_spl_0,
    n2341_inv_p_spl_
  );


  buf

  (
    n2341_inv_n_spl_,
    n2341_inv_n
  );


  buf

  (
    g2620_n_spl_,
    g2620_n
  );


  buf

  (
    g2500_p_spl_,
    g2500_p
  );


  buf

  (
    n4548_lo_n_spl_,
    n4548_lo_n
  );


  buf

  (
    n4548_lo_n_spl_0,
    n4548_lo_n_spl_
  );


  buf

  (
    g2625_p_spl_,
    g2625_p
  );


  buf

  (
    g2625_n_spl_,
    g2625_n
  );


  buf

  (
    g2631_n_spl_,
    g2631_n
  );


  buf

  (
    g2500_n_spl_,
    g2500_n
  );


  buf

  (
    g2500_n_spl_0,
    g2500_n_spl_
  );


  buf

  (
    g2470_p_spl_,
    g2470_p
  );


  buf

  (
    n4548_lo_p_spl_,
    n4548_lo_p
  );


  buf

  (
    n4548_lo_p_spl_0,
    n4548_lo_p_spl_
  );


  buf

  (
    g2642_p_spl_,
    g2642_p
  );


  buf

  (
    g2642_n_spl_,
    g2642_n
  );


  buf

  (
    g2652_p_spl_,
    g2652_p
  );


  buf

  (
    g2652_n_spl_,
    g2652_n
  );


  buf

  (
    n7132_o2_n_spl_,
    n7132_o2_n
  );


  buf

  (
    n7132_o2_n_spl_0,
    n7132_o2_n_spl_
  );


  buf

  (
    n7132_o2_n_spl_1,
    n7132_o2_n_spl_
  );


  buf

  (
    n7136_o2_n_spl_,
    n7136_o2_n
  );


  buf

  (
    G2430_o2_p_spl_,
    G2430_o2_p
  );


  buf

  (
    G2430_o2_p_spl_0,
    G2430_o2_p_spl_
  );


  buf

  (
    G2430_o2_n_spl_,
    G2430_o2_n
  );


  buf

  (
    n7135_o2_p_spl_,
    n7135_o2_p
  );


  buf

  (
    n7135_o2_p_spl_0,
    n7135_o2_p_spl_
  );


  buf

  (
    n7135_o2_p_spl_1,
    n7135_o2_p_spl_
  );


  buf

  (
    n7133_o2_p_spl_,
    n7133_o2_p
  );


  buf

  (
    n7133_o2_p_spl_0,
    n7133_o2_p_spl_
  );


  buf

  (
    n7133_o2_p_spl_00,
    n7133_o2_p_spl_0
  );


  buf

  (
    n7133_o2_p_spl_01,
    n7133_o2_p_spl_0
  );


  buf

  (
    n7133_o2_p_spl_1,
    n7133_o2_p_spl_
  );


  buf

  (
    n3657_lo_p_spl_,
    n3657_lo_p
  );


  buf

  (
    n3657_lo_p_spl_0,
    n3657_lo_p_spl_
  );


  buf

  (
    n3657_lo_p_spl_00,
    n3657_lo_p_spl_0
  );


  buf

  (
    n3657_lo_p_spl_1,
    n3657_lo_p_spl_
  );


  buf

  (
    n4293_lo_p_spl_,
    n4293_lo_p
  );


  buf

  (
    n4293_lo_p_spl_0,
    n4293_lo_p_spl_
  );


  buf

  (
    n4293_lo_p_spl_1,
    n4293_lo_p_spl_
  );


  buf

  (
    g2514_n_spl_,
    g2514_n
  );


  buf

  (
    n4365_lo_p_spl_,
    n4365_lo_p
  );


  buf

  (
    n4365_lo_p_spl_0,
    n4365_lo_p_spl_
  );


  buf

  (
    n4365_lo_p_spl_1,
    n4365_lo_p_spl_
  );


  buf

  (
    g2511_n_spl_,
    g2511_n
  );


  buf

  (
    n4026_lo_p_spl_,
    n4026_lo_p
  );


  buf

  (
    n3726_lo_p_spl_,
    n3726_lo_p
  );


  buf

  (
    n6775_o2_p_spl_,
    n6775_o2_p
  );


  buf

  (
    n6775_o2_p_spl_0,
    n6775_o2_p_spl_
  );


  buf

  (
    n6775_o2_p_spl_1,
    n6775_o2_p_spl_
  );


  buf

  (
    n6774_o2_p_spl_,
    n6774_o2_p
  );


  buf

  (
    n6774_o2_p_spl_0,
    n6774_o2_p_spl_
  );


  buf

  (
    n6774_o2_p_spl_00,
    n6774_o2_p_spl_0
  );


  buf

  (
    n6774_o2_p_spl_01,
    n6774_o2_p_spl_0
  );


  buf

  (
    n6774_o2_p_spl_1,
    n6774_o2_p_spl_
  );


  buf

  (
    n7019_o2_p_spl_,
    n7019_o2_p
  );


  buf

  (
    n7019_o2_p_spl_0,
    n7019_o2_p_spl_
  );


  buf

  (
    n7019_o2_p_spl_1,
    n7019_o2_p_spl_
  );


  buf

  (
    n7015_o2_p_spl_,
    n7015_o2_p
  );


  buf

  (
    n7015_o2_p_spl_0,
    n7015_o2_p_spl_
  );


  buf

  (
    n7015_o2_p_spl_1,
    n7015_o2_p_spl_
  );


  buf

  (
    n6688_o2_p_spl_,
    n6688_o2_p
  );


  buf

  (
    n6688_o2_p_spl_0,
    n6688_o2_p_spl_
  );


  buf

  (
    n6688_o2_p_spl_1,
    n6688_o2_p_spl_
  );


  buf

  (
    n6682_o2_p_spl_,
    n6682_o2_p
  );


  buf

  (
    n6682_o2_p_spl_0,
    n6682_o2_p_spl_
  );


  buf

  (
    n6682_o2_p_spl_00,
    n6682_o2_p_spl_0
  );


  buf

  (
    n6682_o2_p_spl_01,
    n6682_o2_p_spl_0
  );


  buf

  (
    n6682_o2_p_spl_1,
    n6682_o2_p_spl_
  );


  buf

  (
    n6689_o2_p_spl_,
    n6689_o2_p
  );


  buf

  (
    n6689_o2_p_spl_0,
    n6689_o2_p_spl_
  );


  buf

  (
    n6689_o2_p_spl_1,
    n6689_o2_p_spl_
  );


  buf

  (
    n6683_o2_p_spl_,
    n6683_o2_p
  );


  buf

  (
    n6683_o2_p_spl_0,
    n6683_o2_p_spl_
  );


  buf

  (
    n6683_o2_p_spl_00,
    n6683_o2_p_spl_0
  );


  buf

  (
    n6683_o2_p_spl_01,
    n6683_o2_p_spl_0
  );


  buf

  (
    n6683_o2_p_spl_1,
    n6683_o2_p_spl_
  );


  buf

  (
    n7005_o2_p_spl_,
    n7005_o2_p
  );


  buf

  (
    n7005_o2_p_spl_0,
    n7005_o2_p_spl_
  );


  buf

  (
    n7018_o2_p_spl_,
    n7018_o2_p
  );


  buf

  (
    n7018_o2_p_spl_0,
    n7018_o2_p_spl_
  );


  buf

  (
    n7018_o2_p_spl_00,
    n7018_o2_p_spl_0
  );


  buf

  (
    n7018_o2_p_spl_1,
    n7018_o2_p_spl_
  );


  buf

  (
    n6686_o2_p_spl_,
    n6686_o2_p
  );


  buf

  (
    n6686_o2_p_spl_0,
    n6686_o2_p_spl_
  );


  buf

  (
    n6684_o2_p_spl_,
    n6684_o2_p
  );


  buf

  (
    n6684_o2_p_spl_0,
    n6684_o2_p_spl_
  );


  buf

  (
    n6684_o2_p_spl_00,
    n6684_o2_p_spl_0
  );


  buf

  (
    n6684_o2_p_spl_01,
    n6684_o2_p_spl_0
  );


  buf

  (
    n6684_o2_p_spl_1,
    n6684_o2_p_spl_
  );


  buf

  (
    n6687_o2_p_spl_,
    n6687_o2_p
  );


  buf

  (
    n6687_o2_p_spl_0,
    n6687_o2_p_spl_
  );


  buf

  (
    n6685_o2_p_spl_,
    n6685_o2_p
  );


  buf

  (
    n6685_o2_p_spl_0,
    n6685_o2_p_spl_
  );


  buf

  (
    n6685_o2_p_spl_00,
    n6685_o2_p_spl_0
  );


  buf

  (
    n6685_o2_p_spl_01,
    n6685_o2_p_spl_0
  );


  buf

  (
    n6685_o2_p_spl_1,
    n6685_o2_p_spl_
  );


  buf

  (
    n6623_o2_p_spl_,
    n6623_o2_p
  );


  buf

  (
    n6621_o2_p_spl_,
    n6621_o2_p
  );


  buf

  (
    n6669_o2_n_spl_,
    n6669_o2_n
  );


  buf

  (
    n6669_o2_n_spl_0,
    n6669_o2_n_spl_
  );


  buf

  (
    n6669_o2_n_spl_00,
    n6669_o2_n_spl_0
  );


  buf

  (
    n6669_o2_n_spl_1,
    n6669_o2_n_spl_
  );


  buf

  (
    n3936_lo_p_spl_,
    n3936_lo_p
  );


  buf

  (
    n6669_o2_p_spl_,
    n6669_o2_p
  );


  buf

  (
    n6669_o2_p_spl_0,
    n6669_o2_p_spl_
  );


  buf

  (
    n6669_o2_p_spl_00,
    n6669_o2_p_spl_0
  );


  buf

  (
    n6669_o2_p_spl_01,
    n6669_o2_p_spl_0
  );


  buf

  (
    n6669_o2_p_spl_1,
    n6669_o2_p_spl_
  );


  buf

  (
    n3936_lo_n_spl_,
    n3936_lo_n
  );


  buf

  (
    n6627_o2_p_spl_,
    n6627_o2_p
  );


  buf

  (
    n6625_o2_p_spl_,
    n6625_o2_p
  );


  buf

  (
    n4188_lo_p_spl_,
    n4188_lo_p
  );


  buf

  (
    g2529_n_spl_,
    g2529_n
  );


  buf

  (
    g2529_n_spl_0,
    g2529_n_spl_
  );


  buf

  (
    g2529_n_spl_1,
    g2529_n_spl_
  );


  buf

  (
    g2518_p_spl_,
    g2518_p
  );


  buf

  (
    g2702_p_spl_,
    g2702_p
  );


  buf

  (
    g2702_p_spl_0,
    g2702_p_spl_
  );


  buf

  (
    g2526_n_spl_,
    g2526_n
  );


  buf

  (
    g2526_n_spl_0,
    g2526_n_spl_
  );


  buf

  (
    g2526_n_spl_00,
    g2526_n_spl_0
  );


  buf

  (
    g2526_n_spl_1,
    g2526_n_spl_
  );


  buf

  (
    g2519_p_spl_,
    g2519_p
  );


  buf

  (
    g2519_p_spl_0,
    g2519_p_spl_
  );


  buf

  (
    g2520_n_spl_,
    g2520_n
  );


  buf

  (
    g2520_n_spl_0,
    g2520_n_spl_
  );


  buf

  (
    G2486_o2_p_spl_,
    G2486_o2_p
  );


  buf

  (
    G2486_o2_p_spl_0,
    G2486_o2_p_spl_
  );


  buf

  (
    G2486_o2_p_spl_00,
    G2486_o2_p_spl_0
  );


  buf

  (
    G2486_o2_p_spl_01,
    G2486_o2_p_spl_0
  );


  buf

  (
    G2486_o2_p_spl_1,
    G2486_o2_p_spl_
  );


  buf

  (
    G2486_o2_p_spl_10,
    G2486_o2_p_spl_1
  );


  buf

  (
    G2486_o2_p_spl_11,
    G2486_o2_p_spl_1
  );


  buf

  (
    g2521_n_spl_,
    g2521_n
  );


  buf

  (
    g2707_n_spl_,
    g2707_n
  );


  buf

  (
    g2707_n_spl_0,
    g2707_n_spl_
  );


  buf

  (
    n6686_o2_n_spl_,
    n6686_o2_n
  );


  buf

  (
    n6687_o2_n_spl_,
    n6687_o2_n
  );


  buf

  (
    g2714_n_spl_,
    g2714_n
  );


  buf

  (
    n6833_o2_p_spl_,
    n6833_o2_p
  );


  buf

  (
    n6833_o2_p_spl_0,
    n6833_o2_p_spl_
  );


  buf

  (
    n6833_o2_p_spl_1,
    n6833_o2_p_spl_
  );


  buf

  (
    g2669_n_spl_,
    g2669_n
  );


  buf

  (
    g2532_n_spl_,
    g2532_n
  );


  buf

  (
    g2532_n_spl_0,
    g2532_n_spl_
  );


  buf

  (
    g2719_p_spl_,
    g2719_p
  );


  buf

  (
    g2663_n_spl_,
    g2663_n
  );


  buf

  (
    g2723_p_spl_,
    g2723_p
  );


  buf

  (
    g2704_p_spl_,
    g2704_p
  );


  buf

  (
    g2562_p_spl_,
    g2562_p
  );


  buf

  (
    g2703_p_spl_,
    g2703_p
  );


  buf

  (
    g2706_n_spl_,
    g2706_n
  );


  buf

  (
    g2709_n_spl_,
    g2709_n
  );


  buf

  (
    n3756_lo_buf_o2_p_spl_,
    n3756_lo_buf_o2_p
  );


  buf

  (
    n6947_o2_p_spl_,
    n6947_o2_p
  );


  buf

  (
    n6774_o2_n_spl_,
    n6774_o2_n
  );


  buf

  (
    n6774_o2_n_spl_0,
    n6774_o2_n_spl_
  );


  buf

  (
    n6774_o2_n_spl_1,
    n6774_o2_n_spl_
  );


  buf

  (
    n7015_o2_n_spl_,
    n7015_o2_n
  );


  buf

  (
    n6682_o2_n_spl_,
    n6682_o2_n
  );


  buf

  (
    n6682_o2_n_spl_0,
    n6682_o2_n_spl_
  );


  buf

  (
    n6682_o2_n_spl_1,
    n6682_o2_n_spl_
  );


  buf

  (
    n6683_o2_n_spl_,
    n6683_o2_n
  );


  buf

  (
    n6683_o2_n_spl_0,
    n6683_o2_n_spl_
  );


  buf

  (
    n6683_o2_n_spl_1,
    n6683_o2_n_spl_
  );


  buf

  (
    n7018_o2_n_spl_,
    n7018_o2_n
  );


  buf

  (
    n7018_o2_n_spl_0,
    n7018_o2_n_spl_
  );


  buf

  (
    n7005_o2_n_spl_,
    n7005_o2_n
  );


  buf

  (
    n6684_o2_n_spl_,
    n6684_o2_n
  );


  buf

  (
    n6684_o2_n_spl_0,
    n6684_o2_n_spl_
  );


  buf

  (
    n6684_o2_n_spl_1,
    n6684_o2_n_spl_
  );


  buf

  (
    n6685_o2_n_spl_,
    n6685_o2_n
  );


  buf

  (
    n6685_o2_n_spl_0,
    n6685_o2_n_spl_
  );


  buf

  (
    n6685_o2_n_spl_1,
    n6685_o2_n_spl_
  );


  buf

  (
    n2965_inv_n_spl_,
    n2965_inv_n
  );


  buf

  (
    n2965_inv_n_spl_0,
    n2965_inv_n_spl_
  );


  buf

  (
    n2965_inv_n_spl_00,
    n2965_inv_n_spl_0
  );


  buf

  (
    n2965_inv_n_spl_01,
    n2965_inv_n_spl_0
  );


  buf

  (
    n2965_inv_n_spl_1,
    n2965_inv_n_spl_
  );


  buf

  (
    n2965_inv_p_spl_,
    n2965_inv_p
  );


  buf

  (
    n2965_inv_p_spl_0,
    n2965_inv_p_spl_
  );


  buf

  (
    n2965_inv_p_spl_00,
    n2965_inv_p_spl_0
  );


  buf

  (
    n2965_inv_p_spl_01,
    n2965_inv_p_spl_0
  );


  buf

  (
    n2965_inv_p_spl_1,
    n2965_inv_p_spl_
  );


  buf

  (
    n2965_inv_p_spl_10,
    n2965_inv_p_spl_1
  );


  buf

  (
    G1138_o2_n_spl_,
    G1138_o2_n
  );


  buf

  (
    G1138_o2_p_spl_,
    G1138_o2_p
  );


  buf

  (
    n2971_inv_n_spl_,
    n2971_inv_n
  );


  buf

  (
    n2971_inv_n_spl_0,
    n2971_inv_n_spl_
  );


  buf

  (
    n2971_inv_n_spl_00,
    n2971_inv_n_spl_0
  );


  buf

  (
    n2971_inv_n_spl_01,
    n2971_inv_n_spl_0
  );


  buf

  (
    n2971_inv_n_spl_1,
    n2971_inv_n_spl_
  );


  buf

  (
    n2971_inv_p_spl_,
    n2971_inv_p
  );


  buf

  (
    n2971_inv_p_spl_0,
    n2971_inv_p_spl_
  );


  buf

  (
    n2971_inv_p_spl_00,
    n2971_inv_p_spl_0
  );


  buf

  (
    n2971_inv_p_spl_01,
    n2971_inv_p_spl_0
  );


  buf

  (
    n2971_inv_p_spl_1,
    n2971_inv_p_spl_
  );


  buf

  (
    n2971_inv_p_spl_10,
    n2971_inv_p_spl_1
  );


  buf

  (
    n3118_inv_n_spl_,
    n3118_inv_n
  );


  buf

  (
    n3118_inv_n_spl_0,
    n3118_inv_n_spl_
  );


  buf

  (
    n3118_inv_n_spl_00,
    n3118_inv_n_spl_0
  );


  buf

  (
    n3118_inv_n_spl_01,
    n3118_inv_n_spl_0
  );


  buf

  (
    n3118_inv_n_spl_1,
    n3118_inv_n_spl_
  );


  buf

  (
    n3118_inv_n_spl_10,
    n3118_inv_n_spl_1
  );


  buf

  (
    n3118_inv_n_spl_11,
    n3118_inv_n_spl_1
  );


  buf

  (
    n6982_o2_n_spl_,
    n6982_o2_n
  );


  buf

  (
    n3118_inv_p_spl_,
    n3118_inv_p
  );


  buf

  (
    n3118_inv_p_spl_0,
    n3118_inv_p_spl_
  );


  buf

  (
    n3118_inv_p_spl_00,
    n3118_inv_p_spl_0
  );


  buf

  (
    n3118_inv_p_spl_000,
    n3118_inv_p_spl_00
  );


  buf

  (
    n3118_inv_p_spl_01,
    n3118_inv_p_spl_0
  );


  buf

  (
    n3118_inv_p_spl_1,
    n3118_inv_p_spl_
  );


  buf

  (
    n3118_inv_p_spl_10,
    n3118_inv_p_spl_1
  );


  buf

  (
    n3118_inv_p_spl_11,
    n3118_inv_p_spl_1
  );


  buf

  (
    n6982_o2_p_spl_,
    n6982_o2_p
  );


  buf

  (
    n6982_o2_p_spl_0,
    n6982_o2_p_spl_
  );


  buf

  (
    n6982_o2_p_spl_00,
    n6982_o2_p_spl_0
  );


  buf

  (
    n6982_o2_p_spl_1,
    n6982_o2_p_spl_
  );


  buf

  (
    n3127_inv_n_spl_,
    n3127_inv_n
  );


  buf

  (
    n3127_inv_n_spl_0,
    n3127_inv_n_spl_
  );


  buf

  (
    n3127_inv_n_spl_00,
    n3127_inv_n_spl_0
  );


  buf

  (
    n3127_inv_n_spl_01,
    n3127_inv_n_spl_0
  );


  buf

  (
    n3127_inv_n_spl_1,
    n3127_inv_n_spl_
  );


  buf

  (
    n3127_inv_n_spl_10,
    n3127_inv_n_spl_1
  );


  buf

  (
    n3127_inv_n_spl_11,
    n3127_inv_n_spl_1
  );


  buf

  (
    n3127_inv_p_spl_,
    n3127_inv_p
  );


  buf

  (
    n3127_inv_p_spl_0,
    n3127_inv_p_spl_
  );


  buf

  (
    n3127_inv_p_spl_00,
    n3127_inv_p_spl_0
  );


  buf

  (
    n3127_inv_p_spl_000,
    n3127_inv_p_spl_00
  );


  buf

  (
    n3127_inv_p_spl_01,
    n3127_inv_p_spl_0
  );


  buf

  (
    n3127_inv_p_spl_1,
    n3127_inv_p_spl_
  );


  buf

  (
    n3127_inv_p_spl_10,
    n3127_inv_p_spl_1
  );


  buf

  (
    n3127_inv_p_spl_11,
    n3127_inv_p_spl_1
  );


  buf

  (
    G1132_o2_n_spl_,
    G1132_o2_n
  );


  buf

  (
    G1132_o2_p_spl_,
    G1132_o2_p
  );


  buf

  (
    n6945_o2_n_spl_,
    n6945_o2_n
  );


  buf

  (
    n6945_o2_p_spl_,
    n6945_o2_p
  );


  buf

  (
    n6945_o2_p_spl_0,
    n6945_o2_p_spl_
  );


  buf

  (
    n6945_o2_p_spl_00,
    n6945_o2_p_spl_0
  );


  buf

  (
    n6945_o2_p_spl_1,
    n6945_o2_p_spl_
  );


  buf

  (
    g2787_n_spl_,
    g2787_n
  );


  buf

  (
    g2777_p_spl_,
    g2777_p
  );


  buf

  (
    g2787_p_spl_,
    g2787_p
  );


  buf

  (
    g2777_n_spl_,
    g2777_n
  );


  buf

  (
    G1126_o2_n_spl_,
    G1126_o2_n
  );


  buf

  (
    G1126_o2_p_spl_,
    G1126_o2_p
  );


  buf

  (
    n7175_o2_n_spl_,
    n7175_o2_n
  );


  buf

  (
    n7175_o2_p_spl_,
    n7175_o2_p
  );


  buf

  (
    n7175_o2_p_spl_0,
    n7175_o2_p_spl_
  );


  buf

  (
    n7175_o2_p_spl_00,
    n7175_o2_p_spl_0
  );


  buf

  (
    n7175_o2_p_spl_1,
    n7175_o2_p_spl_
  );


  buf

  (
    g2800_p_spl_,
    g2800_p
  );


  buf

  (
    g2462_p_spl_,
    g2462_p
  );


  buf

  (
    g2800_n_spl_,
    g2800_n
  );


  buf

  (
    g2462_n_spl_,
    g2462_n
  );


  buf

  (
    g2462_n_spl_0,
    g2462_n_spl_
  );


  buf

  (
    G1114_o2_n_spl_,
    G1114_o2_n
  );


  buf

  (
    G1114_o2_p_spl_,
    G1114_o2_p
  );


  buf

  (
    n6984_o2_n_spl_,
    n6984_o2_n
  );


  buf

  (
    n6984_o2_p_spl_,
    n6984_o2_p
  );


  buf

  (
    n6984_o2_p_spl_0,
    n6984_o2_p_spl_
  );


  buf

  (
    n6984_o2_p_spl_00,
    n6984_o2_p_spl_0
  );


  buf

  (
    n6984_o2_p_spl_1,
    n6984_o2_p_spl_
  );


  buf

  (
    G1108_o2_n_spl_,
    G1108_o2_n
  );


  buf

  (
    G1108_o2_p_spl_,
    G1108_o2_p
  );


  buf

  (
    n6949_o2_n_spl_,
    n6949_o2_n
  );


  buf

  (
    n6949_o2_p_spl_,
    n6949_o2_p
  );


  buf

  (
    n6949_o2_p_spl_0,
    n6949_o2_p_spl_
  );


  buf

  (
    n6949_o2_p_spl_00,
    n6949_o2_p_spl_0
  );


  buf

  (
    n6949_o2_p_spl_1,
    n6949_o2_p_spl_
  );


  buf

  (
    g2826_n_spl_,
    g2826_n
  );


  buf

  (
    g2816_p_spl_,
    g2816_p
  );


  buf

  (
    g2826_p_spl_,
    g2826_p
  );


  buf

  (
    g2816_n_spl_,
    g2816_n
  );


  buf

  (
    n7453_o2_n_spl_,
    n7453_o2_n
  );


  buf

  (
    n7453_o2_p_spl_,
    n7453_o2_p
  );


  buf

  (
    n7453_o2_p_spl_0,
    n7453_o2_p_spl_
  );


  buf

  (
    n7453_o2_p_spl_00,
    n7453_o2_p_spl_0
  );


  buf

  (
    n7453_o2_p_spl_1,
    n7453_o2_p_spl_
  );


  buf

  (
    n3960_lo_buf_o2_n_spl_,
    n3960_lo_buf_o2_n
  );


  buf

  (
    n3960_lo_buf_o2_p_spl_,
    n3960_lo_buf_o2_p
  );


  buf

  (
    n3960_lo_buf_o2_p_spl_0,
    n3960_lo_buf_o2_p_spl_
  );


  buf

  (
    n3960_lo_buf_o2_p_spl_00,
    n3960_lo_buf_o2_p_spl_0
  );


  buf

  (
    n3960_lo_buf_o2_p_spl_1,
    n3960_lo_buf_o2_p_spl_
  );


  buf

  (
    g2835_p_spl_,
    g2835_p
  );


  buf

  (
    g2832_p_spl_,
    g2832_p
  );


  buf

  (
    g2835_n_spl_,
    g2835_n
  );


  buf

  (
    g2832_n_spl_,
    g2832_n
  );


  buf

  (
    G1041_o2_n_spl_,
    G1041_o2_n
  );


  buf

  (
    G1041_o2_p_spl_,
    G1041_o2_p
  );


  buf

  (
    G1035_o2_n_spl_,
    G1035_o2_n
  );


  buf

  (
    G1035_o2_p_spl_,
    G1035_o2_p
  );


  buf

  (
    g2871_n_spl_,
    g2871_n
  );


  buf

  (
    g2861_p_spl_,
    g2861_p
  );


  buf

  (
    g2871_p_spl_,
    g2871_p
  );


  buf

  (
    g2861_n_spl_,
    g2861_n
  );


  buf

  (
    g2886_n_spl_,
    g2886_n
  );


  buf

  (
    g2880_p_spl_,
    g2880_p
  );


  buf

  (
    g2886_p_spl_,
    g2886_p
  );


  buf

  (
    g2880_n_spl_,
    g2880_n
  );


  buf

  (
    g2874_n_spl_,
    g2874_n
  );


  buf

  (
    g2851_p_spl_,
    g2851_p
  );


  buf

  (
    g2889_p_spl_,
    g2889_p
  );


  buf

  (
    g2851_n_spl_,
    g2851_n
  );


  buf

  (
    g2889_n_spl_,
    g2889_n
  );


  buf

  (
    g2874_p_spl_,
    g2874_p
  );


  buf

  (
    G1093_o2_n_spl_,
    G1093_o2_n
  );


  buf

  (
    G1093_o2_p_spl_,
    G1093_o2_p
  );


  buf

  (
    G1087_o2_n_spl_,
    G1087_o2_n
  );


  buf

  (
    G1087_o2_p_spl_,
    G1087_o2_p
  );


  buf

  (
    g2920_n_spl_,
    g2920_n
  );


  buf

  (
    g2910_p_spl_,
    g2910_p
  );


  buf

  (
    g2920_p_spl_,
    g2920_p
  );


  buf

  (
    g2910_n_spl_,
    g2910_n
  );


  buf

  (
    g2932_n_spl_,
    g2932_n
  );


  buf

  (
    g2926_p_spl_,
    g2926_p
  );


  buf

  (
    g2932_p_spl_,
    g2932_p
  );


  buf

  (
    g2926_n_spl_,
    g2926_n
  );


  buf

  (
    g2923_p_spl_,
    g2923_p
  );


  buf

  (
    g2503_n_spl_,
    g2503_n
  );


  buf

  (
    g2935_n_spl_,
    g2935_n
  );


  buf

  (
    g2503_p_spl_,
    g2503_p
  );


  buf

  (
    g2503_p_spl_0,
    g2503_p_spl_
  );


  buf

  (
    g2935_p_spl_,
    g2935_p
  );


  buf

  (
    g2923_n_spl_,
    g2923_n
  );


  buf

  (
    g2684_n_spl_,
    g2684_n
  );


  buf

  (
    g2684_n_spl_0,
    g2684_n_spl_
  );


  buf

  (
    n4278_lo_p_spl_,
    n4278_lo_p
  );


  buf

  (
    n4278_lo_p_spl_0,
    n4278_lo_p_spl_
  );


  buf

  (
    g2681_n_spl_,
    g2681_n
  );


  buf

  (
    g2681_n_spl_0,
    g2681_n_spl_
  );


  buf

  (
    n4350_lo_p_spl_,
    n4350_lo_p
  );


  buf

  (
    n4350_lo_p_spl_0,
    n4350_lo_p_spl_
  );


  buf

  (
    G2727_o2_p_spl_,
    G2727_o2_p
  );


  buf

  (
    g2953_p_spl_,
    g2953_p
  );


  buf

  (
    g2952_n_spl_,
    g2952_n
  );


  buf

  (
    g2953_n_spl_,
    g2953_n
  );


  buf

  (
    g2952_p_spl_,
    g2952_p
  );


  buf

  (
    g2956_p_spl_,
    g2956_p
  );


  buf

  (
    G3552_o2_n_spl_,
    G3552_o2_n
  );


  buf

  (
    G3552_o2_n_spl_0,
    G3552_o2_n_spl_
  );


  buf

  (
    G3552_o2_n_spl_1,
    G3552_o2_n_spl_
  );


  buf

  (
    g2956_n_spl_,
    g2956_n
  );


  buf

  (
    G3552_o2_p_spl_,
    G3552_o2_p
  );


  buf

  (
    G3552_o2_p_spl_0,
    G3552_o2_p_spl_
  );


  buf

  (
    G3552_o2_p_spl_00,
    G3552_o2_p_spl_0
  );


  buf

  (
    G3552_o2_p_spl_1,
    G3552_o2_p_spl_
  );


  buf

  (
    G3533_o2_p_spl_,
    G3533_o2_p
  );


  buf

  (
    G3533_o2_p_spl_0,
    G3533_o2_p_spl_
  );


  buf

  (
    G3533_o2_n_spl_,
    G3533_o2_n
  );


  buf

  (
    G2543_o2_p_spl_,
    G2543_o2_p
  );


  buf

  (
    g2967_p_spl_,
    g2967_p
  );


  buf

  (
    g2966_n_spl_,
    g2966_n
  );


  buf

  (
    g2967_n_spl_,
    g2967_n
  );


  buf

  (
    g2966_p_spl_,
    g2966_p
  );


  buf

  (
    g2970_p_spl_,
    g2970_p
  );


  buf

  (
    n2647_inv_p_spl_,
    n2647_inv_p
  );


  buf

  (
    n2647_inv_p_spl_0,
    n2647_inv_p_spl_
  );


  buf

  (
    n2647_inv_p_spl_00,
    n2647_inv_p_spl_0
  );


  buf

  (
    n2647_inv_p_spl_1,
    n2647_inv_p_spl_
  );


  buf

  (
    g2970_n_spl_,
    g2970_n
  );


  buf

  (
    n2647_inv_n_spl_,
    n2647_inv_n
  );


  buf

  (
    n2647_inv_n_spl_0,
    n2647_inv_n_spl_
  );


  buf

  (
    n2647_inv_n_spl_1,
    n2647_inv_n_spl_
  );


  buf

  (
    G3645_o2_p_spl_,
    G3645_o2_p
  );


  buf

  (
    G3645_o2_p_spl_0,
    G3645_o2_p_spl_
  );


  buf

  (
    G3645_o2_n_spl_,
    G3645_o2_n
  );


  buf

  (
    g2507_n_spl_,
    g2507_n
  );


  buf

  (
    g2507_n_spl_0,
    g2507_n_spl_
  );


  buf

  (
    g2507_n_spl_1,
    g2507_n_spl_
  );


  buf

  (
    G2715_o2_p_spl_,
    G2715_o2_p
  );


  buf

  (
    g2507_p_spl_,
    g2507_p
  );


  buf

  (
    g2507_p_spl_0,
    g2507_p_spl_
  );


  buf

  (
    G3485_o2_p_spl_,
    G3485_o2_p
  );


  buf

  (
    G3485_o2_p_spl_0,
    G3485_o2_p_spl_
  );


  buf

  (
    G3485_o2_p_spl_00,
    G3485_o2_p_spl_0
  );


  buf

  (
    G3485_o2_p_spl_01,
    G3485_o2_p_spl_0
  );


  buf

  (
    G3485_o2_p_spl_1,
    G3485_o2_p_spl_
  );


  buf

  (
    G3485_o2_p_spl_10,
    G3485_o2_p_spl_1
  );


  buf

  (
    G2720_o2_p_spl_,
    G2720_o2_p
  );


  buf

  (
    G2720_o2_p_spl_0,
    G2720_o2_p_spl_
  );


  buf

  (
    G2720_o2_p_spl_1,
    G2720_o2_p_spl_
  );


  buf

  (
    G3485_o2_n_spl_,
    G3485_o2_n
  );


  buf

  (
    G2720_o2_n_spl_,
    G2720_o2_n
  );


  buf

  (
    G2720_o2_n_spl_0,
    G2720_o2_n_spl_
  );


  buf

  (
    G3546_o2_p_spl_,
    G3546_o2_p
  );


  buf

  (
    G3546_o2_p_spl_0,
    G3546_o2_p_spl_
  );


  buf

  (
    G3546_o2_p_spl_1,
    G3546_o2_p_spl_
  );


  buf

  (
    G3546_o2_n_spl_,
    G3546_o2_n
  );


  buf

  (
    G3546_o2_n_spl_0,
    G3546_o2_n_spl_
  );


  buf

  (
    g2508_p_spl_,
    g2508_p
  );


  buf

  (
    g2983_p_spl_,
    g2983_p
  );


  buf

  (
    g2983_p_spl_0,
    g2983_p_spl_
  );


  buf

  (
    g2983_n_spl_,
    g2983_n
  );


  buf

  (
    g2983_n_spl_0,
    g2983_n_spl_
  );


  buf

  (
    G4051_o2_n_spl_,
    G4051_o2_n
  );


  buf

  (
    G4051_o2_n_spl_0,
    G4051_o2_n_spl_
  );


  buf

  (
    G4051_o2_p_spl_,
    G4051_o2_p
  );


  buf

  (
    G4051_o2_p_spl_0,
    G4051_o2_p_spl_
  );


  buf

  (
    G2410_o2_p_spl_,
    G2410_o2_p
  );


  buf

  (
    n4284_lo_buf_o2_p_spl_,
    n4284_lo_buf_o2_p
  );


  buf

  (
    g2986_n_spl_,
    g2986_n
  );


  buf

  (
    g2985_n_spl_,
    g2985_n
  );


  buf

  (
    g2986_p_spl_,
    g2986_p
  );


  buf

  (
    g2985_p_spl_,
    g2985_p
  );


  buf

  (
    g2989_p_spl_,
    g2989_p
  );


  buf

  (
    g2984_n_spl_,
    g2984_n
  );


  buf

  (
    g2989_n_spl_,
    g2989_n
  );


  buf

  (
    g2984_p_spl_,
    g2984_p
  );


  buf

  (
    g2998_p_spl_,
    g2998_p
  );


  buf

  (
    g2998_n_spl_,
    g2998_n
  );


  buf

  (
    g2504_p_spl_,
    g2504_p
  );


  buf

  (
    g2504_p_spl_0,
    g2504_p_spl_
  );


  buf

  (
    g2504_p_spl_1,
    g2504_p_spl_
  );


  buf

  (
    G2832_o2_p_spl_,
    G2832_o2_p
  );


  buf

  (
    g2504_n_spl_,
    g2504_n
  );


  buf

  (
    g2504_n_spl_0,
    g2504_n_spl_
  );


  buf

  (
    g2504_n_spl_00,
    g2504_n_spl_0
  );


  buf

  (
    g2504_n_spl_01,
    g2504_n_spl_0
  );


  buf

  (
    g2504_n_spl_1,
    g2504_n_spl_
  );


  buf

  (
    g2504_n_spl_10,
    g2504_n_spl_1
  );


  buf

  (
    G3611_o2_p_spl_,
    G3611_o2_p
  );


  buf

  (
    G3611_o2_p_spl_0,
    G3611_o2_p_spl_
  );


  buf

  (
    G3611_o2_p_spl_00,
    G3611_o2_p_spl_0
  );


  buf

  (
    G3611_o2_p_spl_01,
    G3611_o2_p_spl_0
  );


  buf

  (
    G3611_o2_p_spl_1,
    G3611_o2_p_spl_
  );


  buf

  (
    G3611_o2_p_spl_10,
    G3611_o2_p_spl_1
  );


  buf

  (
    G2837_o2_p_spl_,
    G2837_o2_p
  );


  buf

  (
    G2837_o2_p_spl_0,
    G2837_o2_p_spl_
  );


  buf

  (
    G2837_o2_p_spl_1,
    G2837_o2_p_spl_
  );


  buf

  (
    G3611_o2_n_spl_,
    G3611_o2_n
  );


  buf

  (
    G2837_o2_n_spl_,
    G2837_o2_n
  );


  buf

  (
    G2837_o2_n_spl_0,
    G2837_o2_n_spl_
  );


  buf

  (
    G3658_o2_p_spl_,
    G3658_o2_p
  );


  buf

  (
    G3658_o2_p_spl_0,
    G3658_o2_p_spl_
  );


  buf

  (
    G3658_o2_p_spl_1,
    G3658_o2_p_spl_
  );


  buf

  (
    G3658_o2_n_spl_,
    G3658_o2_n
  );


  buf

  (
    G3658_o2_n_spl_0,
    G3658_o2_n_spl_
  );


  buf

  (
    g3011_p_spl_,
    g3011_p
  );


  buf

  (
    g3011_p_spl_0,
    g3011_p_spl_
  );


  buf

  (
    g3011_n_spl_,
    g3011_n
  );


  buf

  (
    g3011_n_spl_0,
    g3011_n_spl_
  );


  buf

  (
    G4065_o2_n_spl_,
    G4065_o2_n
  );


  buf

  (
    G4065_o2_n_spl_0,
    G4065_o2_n_spl_
  );


  buf

  (
    G4065_o2_p_spl_,
    G4065_o2_p
  );


  buf

  (
    G4065_o2_p_spl_0,
    G4065_o2_p_spl_
  );


  buf

  (
    G2472_o2_p_spl_,
    G2472_o2_p
  );


  buf

  (
    n4356_lo_buf_o2_p_spl_,
    n4356_lo_buf_o2_p
  );


  buf

  (
    g3014_n_spl_,
    g3014_n
  );


  buf

  (
    g3013_n_spl_,
    g3013_n
  );


  buf

  (
    g3014_p_spl_,
    g3014_p
  );


  buf

  (
    g3013_p_spl_,
    g3013_p
  );


  buf

  (
    g3017_p_spl_,
    g3017_p
  );


  buf

  (
    g3012_n_spl_,
    g3012_n
  );


  buf

  (
    g3017_n_spl_,
    g3017_n
  );


  buf

  (
    g3012_p_spl_,
    g3012_p
  );


  buf

  (
    g3026_p_spl_,
    g3026_p
  );


  buf

  (
    g3026_n_spl_,
    g3026_n
  );


  buf

  (
    n3678_lo_p_spl_,
    n3678_lo_p
  );


  buf

  (
    g2552_p_spl_,
    g2552_p
  );


  buf

  (
    g2552_p_spl_0,
    g2552_p_spl_
  );


  buf

  (
    n4374_lo_p_spl_,
    n4374_lo_p
  );


  buf

  (
    n4374_lo_p_spl_0,
    n4374_lo_p_spl_
  );


  buf

  (
    g2552_n_spl_,
    g2552_n
  );


  buf

  (
    g2552_n_spl_0,
    g2552_n_spl_
  );


  buf

  (
    n4374_lo_n_spl_,
    n4374_lo_n
  );


  buf

  (
    n4374_lo_n_spl_0,
    n4374_lo_n_spl_
  );


  buf

  (
    n4242_lo_p_spl_,
    n4242_lo_p
  );


  buf

  (
    n4242_lo_p_spl_0,
    n4242_lo_p_spl_
  );


  buf

  (
    g2555_n_spl_,
    g2555_n
  );


  buf

  (
    g2555_n_spl_0,
    g2555_n_spl_
  );


  buf

  (
    n4326_lo_p_spl_,
    n4326_lo_p
  );


  buf

  (
    n4326_lo_p_spl_0,
    n4326_lo_p_spl_
  );


  buf

  (
    g2561_n_spl_,
    g2561_n
  );


  buf

  (
    g2561_n_spl_0,
    g2561_n_spl_
  );


  buf

  (
    n4338_lo_p_spl_,
    n4338_lo_p
  );


  buf

  (
    n4338_lo_p_spl_0,
    n4338_lo_p_spl_
  );


  buf

  (
    g2558_n_spl_,
    g2558_n
  );


  buf

  (
    g2558_n_spl_0,
    g2558_n_spl_
  );


  buf

  (
    n4248_lo_buf_o2_p_spl_,
    n4248_lo_buf_o2_p
  );


  buf

  (
    n4248_lo_buf_o2_p_spl_0,
    n4248_lo_buf_o2_p_spl_
  );


  buf

  (
    n3801_lo_n_spl_,
    n3801_lo_n
  );


  buf

  (
    n3801_lo_n_spl_0,
    n3801_lo_n_spl_
  );


  buf

  (
    n3813_lo_n_spl_,
    n3813_lo_n
  );


  buf

  (
    n3813_lo_n_spl_0,
    n3813_lo_n_spl_
  );


  buf

  (
    n3840_lo_buf_o2_p_spl_,
    n3840_lo_buf_o2_p
  );


  buf

  (
    n3840_lo_buf_o2_p_spl_0,
    n3840_lo_buf_o2_p_spl_
  );


  buf

  (
    n3840_lo_buf_o2_p_spl_1,
    n3840_lo_buf_o2_p_spl_
  );


  buf

  (
    g2672_n_spl_,
    g2672_n
  );


  buf

  (
    g2672_n_spl_0,
    g2672_n_spl_
  );


  buf

  (
    n4305_lo_n_spl_,
    n4305_lo_n
  );


  buf

  (
    G4697_o2_p_spl_,
    G4697_o2_p
  );


  buf

  (
    G4131_o2_n_spl_,
    G4131_o2_n
  );


  buf

  (
    G4697_o2_n_spl_,
    G4697_o2_n
  );


  buf

  (
    G4131_o2_p_spl_,
    G4131_o2_p
  );


  buf

  (
    g3067_p_spl_,
    g3067_p
  );


  buf

  (
    g3067_n_spl_,
    g3067_n
  );


  buf

  (
    g3073_n_spl_,
    g3073_n
  );


  buf

  (
    g2675_n_spl_,
    g2675_n
  );


  buf

  (
    g2675_n_spl_0,
    g2675_n_spl_
  );


  buf

  (
    g2675_n_spl_00,
    g2675_n_spl_0
  );


  buf

  (
    g2675_n_spl_1,
    g2675_n_spl_
  );


  buf

  (
    G4706_o2_n_spl_,
    G4706_o2_n
  );


  buf

  (
    G4170_o2_n_spl_,
    G4170_o2_n
  );


  buf

  (
    G4706_o2_p_spl_,
    G4706_o2_p
  );


  buf

  (
    G4170_o2_p_spl_,
    G4170_o2_p
  );


  buf

  (
    g3077_p_spl_,
    g3077_p
  );


  buf

  (
    g3077_n_spl_,
    g3077_n
  );


  buf

  (
    g3083_n_spl_,
    g3083_n
  );


  buf

  (
    g2678_n_spl_,
    g2678_n
  );


  buf

  (
    g2678_n_spl_0,
    g2678_n_spl_
  );


  buf

  (
    g2678_n_spl_00,
    g2678_n_spl_0
  );


  buf

  (
    g2678_n_spl_1,
    g2678_n_spl_
  );


  buf

  (
    n3957_lo_p_spl_,
    n3957_lo_p
  );


  buf

  (
    n3969_lo_p_spl_,
    n3969_lo_p
  );


  buf

  (
    g2536_n_spl_,
    g2536_n
  );


  buf

  (
    g2536_n_spl_0,
    g2536_n_spl_
  );


  buf

  (
    g2536_n_spl_1,
    g2536_n_spl_
  );


  buf

  (
    g2522_p_spl_,
    g2522_p
  );


  buf

  (
    g2522_p_spl_0,
    g2522_p_spl_
  );


  buf

  (
    g2536_p_spl_,
    g2536_p
  );


  buf

  (
    g2536_p_spl_0,
    g2536_p_spl_
  );


  buf

  (
    g2522_n_spl_,
    g2522_n
  );


  buf

  (
    g3098_p_spl_,
    g3098_p
  );


  buf

  (
    g3041_n_spl_,
    g3041_n
  );


  buf

  (
    g3041_n_spl_0,
    g3041_n_spl_
  );


  buf

  (
    g3041_n_spl_00,
    g3041_n_spl_0
  );


  buf

  (
    g3041_n_spl_1,
    g3041_n_spl_
  );


  buf

  (
    g2542_n_spl_,
    g2542_n
  );


  buf

  (
    g2542_n_spl_0,
    g2542_n_spl_
  );


  buf

  (
    g2523_p_spl_,
    g2523_p
  );


  buf

  (
    g2523_p_spl_0,
    g2523_p_spl_
  );


  buf

  (
    g2542_p_spl_,
    g2542_p
  );


  buf

  (
    g2542_p_spl_0,
    g2542_p_spl_
  );


  buf

  (
    g2523_n_spl_,
    g2523_n
  );


  buf

  (
    g3100_n_spl_,
    g3100_n
  );


  buf

  (
    g3038_p_spl_,
    g3038_p
  );


  buf

  (
    g3038_p_spl_0,
    g3038_p_spl_
  );


  buf

  (
    g3038_p_spl_1,
    g3038_p_spl_
  );


  buf

  (
    g2539_n_spl_,
    g2539_n
  );


  buf

  (
    g2539_n_spl_0,
    g2539_n_spl_
  );


  buf

  (
    g2539_n_spl_00,
    g2539_n_spl_0
  );


  buf

  (
    g2539_n_spl_01,
    g2539_n_spl_0
  );


  buf

  (
    g2539_n_spl_1,
    g2539_n_spl_
  );


  buf

  (
    g2539_p_spl_,
    g2539_p
  );


  buf

  (
    g2539_p_spl_0,
    g2539_p_spl_
  );


  buf

  (
    g2533_p_spl_,
    g2533_p
  );


  buf

  (
    g2533_p_spl_0,
    g2533_p_spl_
  );


  buf

  (
    g2533_p_spl_00,
    g2533_p_spl_0
  );


  buf

  (
    g2533_p_spl_1,
    g2533_p_spl_
  );


  buf

  (
    g2533_n_spl_,
    g2533_n
  );


  buf

  (
    g2533_n_spl_0,
    g2533_n_spl_
  );


  buf

  (
    g2533_n_spl_1,
    g2533_n_spl_
  );


  buf

  (
    g3103_p_spl_,
    g3103_p
  );


  buf

  (
    n3978_lo_p_spl_,
    n3978_lo_p
  );


  buf

  (
    g2550_n_spl_,
    g2550_n
  );


  buf

  (
    g2550_n_spl_0,
    g2550_n_spl_
  );


  buf

  (
    g3106_p_spl_,
    g3106_p
  );


  buf

  (
    g2545_n_spl_,
    g2545_n
  );


  buf

  (
    g2545_n_spl_0,
    g2545_n_spl_
  );


  buf

  (
    g2545_p_spl_,
    g2545_p
  );


  buf

  (
    g2545_p_spl_0,
    g2545_p_spl_
  );


  buf

  (
    g2545_p_spl_1,
    g2545_p_spl_
  );


  buf

  (
    g2517_p_spl_,
    g2517_p
  );


  buf

  (
    g2517_p_spl_0,
    g2517_p_spl_
  );


  buf

  (
    g2517_p_spl_1,
    g2517_p_spl_
  );


  buf

  (
    g2517_n_spl_,
    g2517_n
  );


  buf

  (
    g2517_n_spl_0,
    g2517_n_spl_
  );


  buf

  (
    g2517_n_spl_00,
    g2517_n_spl_0
  );


  buf

  (
    g2517_n_spl_01,
    g2517_n_spl_0
  );


  buf

  (
    g2517_n_spl_1,
    g2517_n_spl_
  );


  buf

  (
    g2517_n_spl_10,
    g2517_n_spl_1
  );


  buf

  (
    g2517_n_spl_11,
    g2517_n_spl_1
  );


  buf

  (
    g3110_n_spl_,
    g3110_n
  );


  buf

  (
    g3112_n_spl_,
    g3112_n
  );


  buf

  (
    g2546_p_spl_,
    g2546_p
  );


  buf

  (
    g2546_p_spl_0,
    g2546_p_spl_
  );


  buf

  (
    g2547_n_spl_,
    g2547_n
  );


  buf

  (
    g2547_p_spl_,
    g2547_p
  );


  buf

  (
    g3119_p_spl_,
    g3119_p
  );


  buf

  (
    g3119_p_spl_0,
    g3119_p_spl_
  );


  buf

  (
    g3121_p_spl_,
    g3121_p
  );


  buf

  (
    g3122_n_spl_,
    g3122_n
  );


  buf

  (
    g3123_n_spl_,
    g3123_n
  );


  buf

  (
    g3120_p_spl_,
    g3120_p
  );


  buf

  (
    g3126_n_spl_,
    g3126_n
  );


  buf

  (
    g3131_p_spl_,
    g3131_p
  );


  buf

  (
    g3131_p_spl_0,
    g3131_p_spl_
  );


  buf

  (
    g3131_n_spl_,
    g3131_n
  );


  buf

  (
    g3131_n_spl_0,
    g3131_n_spl_
  );


  buf

  (
    g3136_p_spl_,
    g3136_p
  );


  buf

  (
    g3128_n_spl_,
    g3128_n
  );


  buf

  (
    g3093_n_spl_,
    g3093_n
  );


  buf

  (
    g3044_n_spl_,
    g3044_n
  );


  buf

  (
    g3044_n_spl_0,
    g3044_n_spl_
  );


  buf

  (
    g3096_n_spl_,
    g3096_n
  );


  buf

  (
    g3047_n_spl_,
    g3047_n
  );


  buf

  (
    g3047_n_spl_0,
    g3047_n_spl_
  );


  buf

  (
    g3115_p_spl_,
    g3115_p
  );


  buf

  (
    g3061_p_spl_,
    g3061_p
  );


  buf

  (
    g3099_p_spl_,
    g3099_p
  );


  buf

  (
    g3104_p_spl_,
    g3104_p
  );


  buf

  (
    g3116_n_spl_,
    g3116_n
  );


  buf

  (
    g3060_n_spl_,
    g3060_n
  );


  buf

  (
    g3101_n_spl_,
    g3101_n
  );


  buf

  (
    g3111_n_spl_,
    g3111_n
  );


  buf

  (
    g2947_p_spl_,
    g2947_p
  );


  buf

  (
    g3062_p_spl_,
    g3062_p
  );


  buf

  (
    g2948_p_spl_,
    g2948_p
  );


  buf

  (
    g3063_p_spl_,
    g3063_p
  );


  buf

  (
    g3119_n_spl_,
    g3119_n
  );


  buf

  (
    G126_p_spl_,
    G126_p
  );


  buf

  (
    G123_p_spl_,
    G123_p
  );


  buf

  (
    G123_p_spl_0,
    G123_p_spl_
  );


  buf

  (
    G123_p_spl_00,
    G123_p_spl_0
  );


  buf

  (
    G123_p_spl_1,
    G123_p_spl_
  );


  buf

  (
    G127_p_spl_,
    G127_p
  );


  buf

  (
    G123_n_spl_,
    G123_n
  );


  buf

  (
    G128_p_spl_,
    G128_p
  );


  buf

  (
    G129_p_spl_,
    G129_p
  );


  buf

  (
    G124_p_spl_,
    G124_p
  );


  buf

  (
    G124_p_spl_0,
    G124_p_spl_
  );


  buf

  (
    G124_p_spl_00,
    G124_p_spl_0
  );


  buf

  (
    G124_p_spl_01,
    G124_p_spl_0
  );


  buf

  (
    G124_p_spl_1,
    G124_p_spl_
  );


  buf

  (
    G105_p_spl_,
    G105_p
  );


  buf

  (
    G124_n_spl_,
    G124_n
  );


  buf

  (
    G124_n_spl_0,
    G124_n_spl_
  );


  buf

  (
    G107_p_spl_,
    G107_p
  );


  buf

  (
    G109_p_spl_,
    G109_p
  );


  buf

  (
    n4419_lo_n_spl_,
    n4419_lo_n
  );


  buf

  (
    n4419_lo_n_spl_0,
    n4419_lo_n_spl_
  );


  buf

  (
    n4431_lo_p_spl_,
    n4431_lo_p
  );


  buf

  (
    n2619_lo_n_spl_,
    n2619_lo_n
  );


  buf

  (
    n2619_lo_n_spl_0,
    n2619_lo_n_spl_
  );


  buf

  (
    n2619_lo_n_spl_1,
    n2619_lo_n_spl_
  );


  buf

  (
    n3975_lo_n_spl_,
    n3975_lo_n
  );


  buf

  (
    g1207_n_spl_,
    g1207_n
  );


  buf

  (
    n4056_lo_buf_o2_p_spl_,
    n4056_lo_buf_o2_p
  );


  buf

  (
    n2650_inv_p_spl_,
    n2650_inv_p
  );


  buf

  (
    n2650_inv_p_spl_0,
    n2650_inv_p_spl_
  );


  buf

  (
    n7396_o2_p_spl_,
    n7396_o2_p
  );


  buf

  (
    n7396_o2_p_spl_0,
    n7396_o2_p_spl_
  );


  buf

  (
    n7396_o2_p_spl_1,
    n7396_o2_p_spl_
  );


  buf

  (
    n7398_o2_p_spl_,
    n7398_o2_p
  );


  buf

  (
    n7398_o2_p_spl_0,
    n7398_o2_p_spl_
  );


  buf

  (
    n7398_o2_p_spl_1,
    n7398_o2_p_spl_
  );


  buf

  (
    n7400_o2_p_spl_,
    n7400_o2_p
  );


  buf

  (
    n7400_o2_p_spl_0,
    n7400_o2_p_spl_
  );


  buf

  (
    n7400_o2_p_spl_1,
    n7400_o2_p_spl_
  );


  buf

  (
    n7402_o2_p_spl_,
    n7402_o2_p
  );


  buf

  (
    n7402_o2_p_spl_0,
    n7402_o2_p_spl_
  );


  buf

  (
    n7402_o2_p_spl_1,
    n7402_o2_p_spl_
  );


  buf

  (
    n3708_lo_buf_o2_p_spl_,
    n3708_lo_buf_o2_p
  );


  buf

  (
    n4008_lo_buf_o2_p_spl_,
    n4008_lo_buf_o2_p
  );


  buf

  (
    n3732_lo_buf_o2_p_spl_,
    n3732_lo_buf_o2_p
  );


  buf

  (
    n4032_lo_buf_o2_p_spl_,
    n4032_lo_buf_o2_p
  );


  buf

  (
    n3684_lo_buf_o2_p_spl_,
    n3684_lo_buf_o2_p
  );


  buf

  (
    g2592_p_spl_,
    g2592_p
  );


  buf

  (
    g2611_n_spl_,
    g2611_n
  );


  buf

  (
    g2641_n_spl_,
    g2641_n
  );


  buf

  (
    g2660_n_spl_,
    g2660_n
  );


  buf

  (
    g2666_n_spl_,
    g2666_n
  );


  buf

  (
    n3801_lo_p_spl_,
    n3801_lo_p
  );


  buf

  (
    n3813_lo_p_spl_,
    n3813_lo_p
  );


  buf

  (
    g2962_p_spl_,
    g2962_p
  );


  buf

  (
    g2976_p_spl_,
    g2976_p
  );


  buf

  (
    g2995_n_spl_,
    g2995_n
  );


  buf

  (
    g3004_n_spl_,
    g3004_n
  );


  buf

  (
    g3023_p_spl_,
    g3023_p
  );


  buf

  (
    g3032_p_spl_,
    g3032_p
  );


  buf

  (
    n4314_lo_p_spl_,
    n4314_lo_p
  );


  buf

  (
    n4314_lo_p_spl_0,
    n4314_lo_p_spl_
  );


  buf

  (
    g3035_n_spl_,
    g3035_n
  );


  buf

  (
    g3035_n_spl_0,
    g3035_n_spl_
  );


  buf

  (
    n3777_lo_p_spl_,
    n3777_lo_p
  );


  buf

  (
    n3825_lo_p_spl_,
    n3825_lo_p
  );


  buf

  (
    g3166_n_spl_,
    g3166_n
  );


  buf

  (
    g3169_n_spl_,
    g3169_n
  );


  buf

  (
    g3172_n_spl_,
    g3172_n
  );


  buf

  (
    g3175_n_spl_,
    g3175_n
  );


  buf

  (
    G138_p_spl_,
    G138_p
  );


  buf

  (
    G139_p_spl_,
    G139_p
  );


  buf

  (
    G149_p_spl_,
    G149_p
  );


  buf

  (
    G150_p_spl_,
    G150_p
  );


endmodule
