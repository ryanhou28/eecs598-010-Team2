



module mult(a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, product_0_, product_1_, product_2_, product_3_, product_4_, product_5_, product_6_, product_7_);input a_0_;
  input a_1_;
  input a_2_;
  input a_3_;
  input a_4_;
  input a_5_;
  input a_6_;
  input a_7_;
  input b_0_;
  input b_1_;
  input b_2_;
  input b_3_;
  input b_4_;
  input b_5_;
  input b_6_;
  input b_7_;
  output product_0_;
  output product_1_;
  output product_2_;
  output product_3_;
  output product_4_;
  output product_5_;
  output product_6_;
  output product_7_;
  
  wire wire_zeros;
  assign wire_zeros = 1'b0;
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  
  
  
  
  
  
  
  
  
  wire a_0_;
  wire a_1_;
  wire a_2_;
  wire a_3_;
  wire a_4_;
  wire a_5_;
  wire a_6_;
  wire a_7_;
  
  
  
  
  
  
  
  
  
  wire b_0_;
  wire b_1_;
  wire b_2_;
  wire b_3_;
  wire b_4_;
  wire b_5_;
  wire b_6_;
  wire b_7_;
  
  
  
  
  
  
  
  
  
  wire product_0_;
  wire product_1_;
  wire product_2_;
  wire product_3_;
  wire product_4_;
  wire product_5_;
  wire product_6_;
  wire product_7_;
  
  
  nand (_0160_, a_0_, a_0_);
  
  
  nand (_0171_, a_1_, a_1_);
  
  
  nand (_0182_, a_2_, a_2_);
  
  
  nand (_0193_, a_3_, a_3_);
  
  
  nand (_0204_, a_4_, a_4_);
  
  
  nand (_0215_, a_5_, a_5_);
  
  
  nand (_0226_, a_6_, a_6_);
  
  
  nand (_0237_, a_7_, a_7_);
  
  
  nand (_0248_, b_7_, b_7_);
  nand (_0259_, a_7_, b_3_);
  nand (_0270_, a_7_, b_4_);
  
  
  nand (_0281_, _0270_, _0270_);
  nand (_0292_, b_3_, _0281_);
  nand (_0303_, _0259_, _0270_);
  nand (_0314_, _0292_, _0303_);
  
  
  nand (_0325_, _0314_, _0314_);
  nand (_0336_, a_7_, b_5_);
  
  
  nand (_0347_, _0336_, _0336_);
  nand (_0358_, _0325_, _0347_);
  nand (_0369_, _0314_, _0336_);
  nand (_0380_, _0358_, _0369_);
  
  
  nand (_0391_, _0380_, _0380_);
  nand (_0402_, a_7_, b_1_);
  nand (_0413_, a_7_, b_0_);
  
  
  nand (_0424_, _0413_, _0413_);
  nand (_0435_, b_1_, _0424_);
  
  
  nand (_0446_, _0435_, _0435_);
  nand (_0457_, a_7_, b_2_);
  
  
  nand (_0468_, _0457_, _0457_);
  nand (_0479_, _0402_, _0413_);
  
  
  nand (_0490_, _0479_, _0479_);
  nand (_0501_, _0435_, _0479_);
  
  
  nand (_0512_, _0501_, _0501_);
  nand (_0523_, _0457_, _0501_);
  nand (_0534_, _0468_, _0512_);
  nand (_0545_, _0523_, _0534_);
  nand (_0556_, b_2_, _0446_);
  
  
  nand (_0567_, _0556_, _0556_);
  nand (_0578_, _0457_, _0490_);
  nand (_0589_, _0556_, _0578_);
  
  
  nand (_0600_, _0589_, _0589_);
  nand (_0611_, _0391_, _0600_);
  nand (_0622_, _0380_, _0589_);
  
  
  nand (_0633_, _0622_, _0622_);
  nand (_0644_, _0611_, _0622_);
  
  
  nand (_0655_, _0644_, _0644_);
  nand (_0666_, a_6_, b_5_);
  
  
  nand (_0677_, _0666_, _0666_);
  nand (_0688_, _0325_, _0677_);
  nand (_0699_, _0314_, _0666_);
  nand (_0710_, _0688_, _0699_);
  
  
  nand (_0721_, _0710_, _0710_);
  nand (_0731_, _0600_, _0721_);
  nand (_0742_, _0556_, _0731_);
  
  
  nand (_0753_, _0742_, _0742_);
  nand (_0764_, _0655_, _0742_);
  nand (_0775_, a_5_, b_6_);
  
  
  nand (_0786_, _0775_, _0775_);
  nand (_0795_, _0204_, b_7_);
  
  
  nand (_0804_, _0795_, _0795_);
  nand (_0813_, _0786_, _0804_);
  
  
  nand (_0817_, _0813_, _0813_);
  nand (_0818_, _0292_, _0688_);
  
  
  nand (_0819_, _0818_, _0818_);
  nand (_0820_, a_6_, b_6_);
  
  
  nand (_0821_, _0820_, _0820_);
  nand (_0822_, _0215_, b_7_);
  
  
  nand (_0823_, _0822_, _0822_);
  nand (_0824_, _0821_, _0823_);
  
  
  nand (_0825_, _0824_, _0824_);
  nand (_0826_, _0820_, _0822_);
  nand (_0827_, _0824_, _0826_);
  
  
  nand (_0828_, _0827_, _0827_);
  nand (_0829_, _0818_, _0828_);
  nand (_0830_, _0819_, _0827_);
  nand (_0000_, _0829_, _0830_);
  
  
  nand (_0001_, _0000_, _0000_);
  nand (_0002_, _0817_, _0001_);
  nand (_0003_, _0813_, _0000_);
  nand (_0004_, _0002_, _0003_);
  
  
  nand (_0005_, _0004_, _0004_);
  nand (_0006_, _0644_, _0753_);
  nand (_0007_, _0764_, _0006_);
  
  
  nand (_0008_, _0007_, _0007_);
  nand (_0009_, _0005_, _0008_);
  nand (_0010_, _0764_, _0009_);
  
  
  nand (_0011_, _0010_, _0010_);
  nand (_0012_, _0391_, _0567_);
  nand (_0013_, _0556_, _0633_);
  nand (_0014_, _0012_, _0013_);
  
  
  nand (_0015_, _0014_, _0014_);
  nand (_0016_, _0292_, _0358_);
  
  
  nand (_0017_, _0016_, _0016_);
  nand (_0018_, a_7_, b_6_);
  
  
  nand (_0019_, _0018_, _0018_);
  nand (_0020_, _0226_, b_7_);
  
  
  nand (_0021_, _0020_, _0020_);
  nand (_0022_, _0019_, _0020_);
  nand (_0023_, _0019_, _0021_);
  nand (_0024_, _0018_, _0020_);
  nand (_0025_, _0023_, _0024_);
  
  
  nand (_0026_, _0025_, _0025_);
  nand (_0027_, _0016_, _0026_);
  nand (_0028_, _0017_, _0025_);
  nand (_0029_, _0027_, _0028_);
  
  
  nand (_0030_, _0029_, _0029_);
  nand (_0031_, _0825_, _0030_);
  nand (_0032_, _0824_, _0029_);
  nand (_0033_, _0031_, _0032_);
  
  
  nand (_0034_, _0033_, _0033_);
  nand (_0035_, _0015_, _0034_);
  nand (_0036_, _0014_, _0033_);
  nand (_0037_, _0035_, _0036_);
  
  
  nand (_0038_, _0037_, _0037_);
  nand (_0039_, _0010_, _0038_);
  nand (_0040_, _0829_, _0002_);
  
  
  nand (_0041_, _0040_, _0040_);
  nand (_0042_, _0011_, _0037_);
  nand (_0043_, _0039_, _0042_);
  
  
  nand (_0044_, _0043_, _0043_);
  nand (_0045_, _0040_, _0044_);
  nand (_0046_, _0039_, _0045_);
  
  
  nand (_0047_, _0046_, _0046_);
  nand (_0048_, _0027_, _0031_);
  
  
  nand (_0049_, _0048_, _0048_);
  nand (_0050_, _0237_, b_7_);
  nand (_0051_, _0018_, _0050_);
  nand (_0052_, _0023_, _0051_);
  nand (_0053_, _0022_, _0050_);
  nand (_0054_, _0017_, _0052_);
  
  
  nand (_0055_, _0054_, _0054_);
  nand (_0056_, _0016_, _0053_);
  nand (_0057_, _0054_, _0056_);
  
  
  nand (_0058_, _0057_, _0057_);
  nand (_0059_, _0015_, _0057_);
  nand (_0060_, _0014_, _0058_);
  nand (_0061_, _0059_, _0060_);
  
  
  nand (_0062_, _0061_, _0061_);
  nand (_0063_, _0012_, _0035_);
  
  
  nand (_0064_, _0063_, _0063_);
  nand (_0065_, _0061_, _0063_);
  nand (_0066_, _0062_, _0064_);
  nand (_0067_, _0065_, _0066_);
  
  
  nand (_0068_, _0067_, _0067_);
  nand (_0069_, _0048_, _0068_);
  nand (_0070_, _0049_, _0067_);
  nand (_0071_, _0069_, _0070_);
  
  
  nand (_0072_, _0071_, _0071_);
  nand (_0073_, _0046_, _0072_);
  nand (_0074_, _0047_, _0071_);
  nand (_0075_, _0073_, _0074_);
  
  
  nand (_0076_, _0075_, _0075_);
  nand (_0077_, a_5_, b_5_);
  
  
  nand (_0078_, _0077_, _0077_);
  nand (_0079_, a_6_, b_4_);
  
  
  nand (_0080_, _0079_, _0079_);
  nand (_0081_, a_6_, b_3_);
  
  
  nand (_0082_, _0081_, _0081_);
  nand (_0083_, _0281_, _0082_);
  nand (_0084_, _0259_, _0079_);
  nand (_0085_, _0083_, _0084_);
  
  
  nand (_0086_, _0085_, _0085_);
  nand (_0087_, _0078_, _0086_);
  nand (_0088_, _0077_, _0085_);
  nand (_0089_, _0087_, _0088_);
  
  
  nand (_0090_, _0089_, _0089_);
  nand (_0091_, _0600_, _0090_);
  nand (_0092_, _0556_, _0091_);
  
  
  nand (_0093_, _0092_, _0092_);
  nand (_0094_, _0589_, _0710_);
  nand (_0095_, _0731_, _0094_);
  
  
  nand (_0096_, _0095_, _0095_);
  nand (_0097_, _0092_, _0096_);
  nand (_0098_, a_4_, b_6_);
  
  
  nand (_0099_, _0098_, _0098_);
  nand (_0100_, _0193_, b_7_);
  
  
  nand (_0101_, _0100_, _0100_);
  nand (_0102_, _0099_, _0101_);
  
  
  nand (_0103_, _0102_, _0102_);
  nand (_0104_, _0083_, _0087_);
  
  
  nand (_0105_, _0104_, _0104_);
  nand (_0106_, _0775_, _0795_);
  nand (_0107_, _0813_, _0106_);
  
  
  nand (_0108_, _0107_, _0107_);
  nand (_0109_, _0104_, _0108_);
  nand (_0110_, _0105_, _0107_);
  nand (_0111_, _0109_, _0110_);
  
  
  nand (_0112_, _0111_, _0111_);
  nand (_0113_, _0103_, _0112_);
  nand (_0114_, _0102_, _0111_);
  nand (_0115_, _0113_, _0114_);
  
  
  nand (_0116_, _0115_, _0115_);
  nand (_0117_, _0093_, _0095_);
  nand (_0118_, _0097_, _0117_);
  
  
  nand (_0119_, _0118_, _0118_);
  nand (_0120_, _0116_, _0119_);
  nand (_0121_, _0097_, _0120_);
  
  
  nand (_0122_, _0121_, _0121_);
  nand (_0123_, _0004_, _0007_);
  nand (_0124_, _0009_, _0123_);
  
  
  nand (_0125_, _0124_, _0124_);
  nand (_0126_, _0121_, _0125_);
  nand (_0127_, _0109_, _0113_);
  
  
  nand (_0128_, _0127_, _0127_);
  nand (_0129_, _0122_, _0124_);
  nand (_0130_, _0126_, _0129_);
  
  
  nand (_0131_, _0130_, _0130_);
  nand (_0132_, _0127_, _0131_);
  nand (_0133_, _0126_, _0132_);
  
  
  nand (_0134_, _0133_, _0133_);
  nand (_0135_, _0041_, _0043_);
  nand (_0136_, _0045_, _0135_);
  
  
  nand (_0137_, _0136_, _0136_);
  nand (_0138_, _0133_, _0137_);
  nand (_0139_, _0134_, _0136_);
  nand (_0140_, a_4_, b_5_);
  
  
  nand (_0141_, _0140_, _0140_);
  nand (_0142_, a_5_, b_4_);
  nand (_0143_, a_5_, b_3_);
  
  
  nand (_0144_, _0143_, _0143_);
  nand (_0145_, _0080_, _0144_);
  nand (_0146_, _0081_, _0142_);
  nand (_0147_, _0145_, _0146_);
  
  
  nand (_0148_, _0147_, _0147_);
  nand (_0149_, _0141_, _0148_);
  nand (_0150_, _0140_, _0147_);
  nand (_0151_, _0149_, _0150_);
  
  
  nand (_0152_, _0151_, _0151_);
  nand (_0153_, a_6_, b_2_);
  
  
  nand (_0154_, _0153_, _0153_);
  nand (_0155_, _0512_, _0154_);
  nand (_0156_, _0435_, _0155_);
  
  
  nand (_0157_, _0156_, _0156_);
  nand (_0158_, _0545_, _0157_);
  nand (_0159_, _0556_, _0158_);
  
  
  nand (_0161_, _0159_, _0159_);
  nand (_0162_, _0152_, _0161_);
  nand (_0163_, _0556_, _0162_);
  
  
  nand (_0164_, _0163_, _0163_);
  nand (_0165_, _0589_, _0089_);
  nand (_0166_, _0091_, _0165_);
  
  
  nand (_0167_, _0166_, _0166_);
  nand (_0168_, _0163_, _0167_);
  nand (_0169_, a_3_, b_6_);
  
  
  nand (_0170_, _0169_, _0169_);
  nand (_0172_, _0182_, b_7_);
  
  
  nand (_0173_, _0172_, _0172_);
  nand (_0174_, _0170_, _0173_);
  
  
  nand (_0175_, _0174_, _0174_);
  nand (_0176_, _0145_, _0149_);
  
  
  nand (_0177_, _0176_, _0176_);
  nand (_0178_, _0098_, _0100_);
  nand (_0179_, _0102_, _0178_);
  
  
  nand (_0180_, _0179_, _0179_);
  nand (_0181_, _0176_, _0180_);
  nand (_0183_, _0177_, _0179_);
  nand (_0184_, _0181_, _0183_);
  
  
  nand (_0185_, _0184_, _0184_);
  nand (_0186_, _0175_, _0185_);
  nand (_0187_, _0174_, _0184_);
  nand (_0188_, _0186_, _0187_);
  
  
  nand (_0189_, _0188_, _0188_);
  nand (_0190_, _0164_, _0166_);
  nand (_0191_, _0168_, _0190_);
  
  
  nand (_0192_, _0191_, _0191_);
  nand (_0194_, _0189_, _0192_);
  nand (_0195_, _0168_, _0194_);
  
  
  nand (_0196_, _0195_, _0195_);
  nand (_0197_, _0115_, _0118_);
  nand (_0198_, _0120_, _0197_);
  
  
  nand (_0199_, _0198_, _0198_);
  nand (_0200_, _0195_, _0199_);
  nand (_0201_, _0181_, _0186_);
  
  
  nand (_0202_, _0201_, _0201_);
  nand (_0203_, _0196_, _0198_);
  nand (_0205_, _0200_, _0203_);
  
  
  nand (_0206_, _0205_, _0205_);
  nand (_0207_, _0201_, _0206_);
  nand (_0208_, _0200_, _0207_);
  
  
  nand (_0209_, _0208_, _0208_);
  nand (_0210_, _0128_, _0130_);
  nand (_0211_, _0132_, _0210_);
  
  
  nand (_0212_, _0211_, _0211_);
  nand (_0213_, _0208_, _0212_);
  nand (_0214_, b_7_, _0424_);
  nand (_0216_, a_6_, b_1_);
  
  
  nand (_0217_, _0216_, _0216_);
  nand (_0218_, _0248_, _0413_);
  nand (_0219_, _0214_, _0218_);
  
  
  nand (_0220_, _0219_, _0219_);
  nand (_0221_, _0217_, _0220_);
  nand (_0222_, _0214_, _0221_);
  
  
  nand (_0223_, _0222_, _0222_);
  nand (_0224_, _0501_, _0153_);
  nand (_0225_, _0155_, _0224_);
  
  
  nand (_0227_, _0225_, _0225_);
  nand (_0228_, _0222_, _0227_);
  nand (_0229_, a_3_, b_5_);
  
  
  nand (_0230_, _0229_, _0229_);
  nand (_0231_, a_4_, b_4_);
  
  
  nand (_0232_, _0231_, _0231_);
  nand (_0233_, a_4_, b_3_);
  nand (_0234_, _0144_, _0232_);
  nand (_0235_, _0143_, _0231_);
  nand (_0236_, _0234_, _0235_);
  
  
  nand (_0238_, _0236_, _0236_);
  nand (_0239_, _0230_, _0238_);
  nand (_0240_, _0229_, _0236_);
  nand (_0241_, _0239_, _0240_);
  
  
  nand (_0242_, _0241_, _0241_);
  nand (_0243_, _0223_, _0225_);
  nand (_0244_, _0228_, _0243_);
  
  
  nand (_0245_, _0244_, _0244_);
  nand (_0246_, _0242_, _0245_);
  nand (_0247_, _0228_, _0246_);
  
  
  nand (_0249_, _0247_, _0247_);
  nand (_0250_, _0151_, _0159_);
  nand (_0251_, _0162_, _0250_);
  
  
  nand (_0252_, _0251_, _0251_);
  nand (_0253_, _0247_, _0252_);
  nand (_0254_, a_2_, b_6_);
  
  
  nand (_0255_, _0254_, _0254_);
  nand (_0256_, _0171_, b_7_);
  
  
  nand (_0257_, _0256_, _0256_);
  nand (_0258_, _0255_, _0257_);
  
  
  nand (_0260_, _0258_, _0258_);
  nand (_0261_, _0234_, _0239_);
  
  
  nand (_0262_, _0261_, _0261_);
  nand (_0263_, _0169_, _0172_);
  nand (_0264_, _0174_, _0263_);
  
  
  nand (_0265_, _0264_, _0264_);
  nand (_0266_, _0261_, _0265_);
  nand (_0267_, _0262_, _0264_);
  nand (_0268_, _0266_, _0267_);
  
  
  nand (_0269_, _0268_, _0268_);
  nand (_0271_, _0260_, _0269_);
  nand (_0272_, _0258_, _0268_);
  nand (_0273_, _0271_, _0272_);
  
  
  nand (_0274_, _0273_, _0273_);
  nand (_0275_, _0249_, _0251_);
  nand (_0276_, _0253_, _0275_);
  
  
  nand (_0277_, _0276_, _0276_);
  nand (_0278_, _0274_, _0277_);
  nand (_0279_, _0253_, _0278_);
  
  
  nand (_0280_, _0279_, _0279_);
  nand (_0282_, _0188_, _0191_);
  nand (_0283_, _0194_, _0282_);
  
  
  nand (_0284_, _0283_, _0283_);
  nand (_0285_, _0279_, _0284_);
  nand (_0286_, _0266_, _0271_);
  
  
  nand (_0287_, _0286_, _0286_);
  nand (_0288_, _0280_, _0283_);
  nand (_0289_, _0285_, _0288_);
  
  
  nand (_0290_, _0289_, _0289_);
  nand (_0291_, _0286_, _0290_);
  nand (_0293_, _0285_, _0291_);
  
  
  nand (_0294_, _0293_, _0293_);
  nand (_0295_, _0202_, _0205_);
  nand (_0296_, _0207_, _0295_);
  
  
  nand (_0297_, _0296_, _0296_);
  nand (_0298_, _0293_, _0297_);
  nand (_0299_, _0294_, _0296_);
  nand (_0300_, _0298_, _0299_);
  
  
  nand (_0301_, _0300_, _0300_);
  nand (_0302_, a_6_, b_0_);
  nand (_0304_, a_5_, b_1_);
  nand (_0305_, a_5_, b_0_);
  
  
  nand (_0306_, _0305_, _0305_);
  nand (_0307_, _0217_, _0306_);
  nand (_0308_, a_4_, b_2_);
  
  
  nand (_0309_, _0308_, _0308_);
  nand (_0310_, _0302_, _0304_);
  nand (_0311_, _0307_, _0310_);
  
  
  nand (_0312_, _0311_, _0311_);
  nand (_0313_, _0309_, _0312_);
  nand (_0315_, _0307_, _0313_);
  
  
  nand (_0316_, _0315_, _0315_);
  nand (_0317_, _0216_, _0219_);
  nand (_0318_, _0221_, _0317_);
  
  
  nand (_0319_, _0318_, _0318_);
  nand (_0320_, _0315_, _0319_);
  nand (_0321_, a_3_, b_4_);
  
  
  nand (_0322_, _0321_, _0321_);
  nand (_0323_, a_5_, b_2_);
  nand (_0324_, _0144_, _0309_);
  nand (_0326_, _0233_, _0323_);
  nand (_0327_, _0324_, _0326_);
  
  
  nand (_0328_, _0327_, _0327_);
  nand (_0329_, _0322_, _0328_);
  nand (_0330_, _0321_, _0327_);
  nand (_0331_, _0329_, _0330_);
  
  
  nand (_0332_, _0331_, _0331_);
  nand (_0333_, _0316_, _0318_);
  nand (_0334_, _0320_, _0333_);
  
  
  nand (_0335_, _0334_, _0334_);
  nand (_0337_, _0332_, _0335_);
  nand (_0338_, _0320_, _0337_);
  
  
  nand (_0339_, _0338_, _0338_);
  nand (_0340_, _0241_, _0244_);
  nand (_0341_, _0246_, _0340_);
  
  
  nand (_0342_, _0341_, _0341_);
  nand (_0343_, _0338_, _0342_);
  nand (_0344_, a_2_, b_5_);
  nand (_0345_, a_1_, b_6_);
  nand (_0346_, a_1_, b_5_);
  
  
  nand (_0348_, _0346_, _0346_);
  nand (_0349_, _0255_, _0348_);
  nand (_0350_, _0160_, b_7_);
  
  
  nand (_0351_, _0350_, _0350_);
  nand (_0352_, _0344_, _0345_);
  nand (_0353_, _0349_, _0352_);
  
  
  nand (_0354_, _0353_, _0353_);
  nand (_0355_, _0351_, _0354_);
  nand (_0356_, _0349_, _0355_);
  
  
  nand (_0357_, _0356_, _0356_);
  nand (_0359_, _0324_, _0329_);
  
  
  nand (_0360_, _0359_, _0359_);
  nand (_0361_, _0254_, _0256_);
  nand (_0362_, _0258_, _0361_);
  
  
  nand (_0363_, _0362_, _0362_);
  nand (_0364_, _0359_, _0363_);
  nand (_0365_, _0360_, _0362_);
  nand (_0366_, _0364_, _0365_);
  
  
  nand (_0367_, _0366_, _0366_);
  nand (_0368_, _0356_, _0367_);
  nand (_0370_, _0357_, _0366_);
  nand (_0371_, _0368_, _0370_);
  
  
  nand (_0372_, _0371_, _0371_);
  nand (_0373_, _0339_, _0341_);
  nand (_0374_, _0343_, _0373_);
  
  
  nand (_0375_, _0374_, _0374_);
  nand (_0376_, _0372_, _0375_);
  nand (_0377_, _0343_, _0376_);
  
  
  nand (_0378_, _0377_, _0377_);
  nand (_0379_, _0273_, _0276_);
  nand (_0381_, _0278_, _0379_);
  
  
  nand (_0382_, _0381_, _0381_);
  nand (_0383_, _0377_, _0382_);
  nand (_0384_, _0364_, _0368_);
  
  
  nand (_0385_, _0384_, _0384_);
  nand (_0386_, _0378_, _0381_);
  nand (_0387_, _0383_, _0386_);
  
  
  nand (_0388_, _0387_, _0387_);
  nand (_0389_, _0384_, _0388_);
  nand (_0390_, _0383_, _0389_);
  
  
  nand (_0392_, _0390_, _0390_);
  nand (_0393_, _0287_, _0289_);
  nand (_0394_, _0291_, _0393_);
  
  
  nand (_0395_, _0394_, _0394_);
  nand (_0396_, _0390_, _0395_);
  nand (_0397_, _0392_, _0394_);
  nand (_0398_, _0396_, _0397_);
  
  
  nand (_0399_, _0398_, _0398_);
  nand (_0400_, a_4_, b_1_);
  
  
  nand (_0401_, _0400_, _0400_);
  nand (_0403_, a_4_, b_0_);
  
  
  nand (_0404_, _0403_, _0403_);
  nand (_0405_, _0306_, _0401_);
  nand (_0406_, a_3_, b_2_);
  
  
  nand (_0407_, _0406_, _0406_);
  nand (_0408_, _0305_, _0400_);
  nand (_0409_, _0405_, _0408_);
  
  
  nand (_0410_, _0409_, _0409_);
  nand (_0411_, _0407_, _0410_);
  nand (_0412_, _0405_, _0411_);
  
  
  nand (_0414_, _0412_, _0412_);
  nand (_0415_, _0308_, _0311_);
  nand (_0416_, _0313_, _0415_);
  
  
  nand (_0417_, _0416_, _0416_);
  nand (_0418_, _0412_, _0417_);
  nand (_0419_, a_3_, b_3_);
  nand (_0420_, a_2_, b_4_);
  nand (_0421_, a_2_, b_3_);
  
  
  nand (_0422_, _0421_, _0421_);
  nand (_0423_, _0322_, _0422_);
  nand (_0425_, _0419_, _0420_);
  nand (_0426_, _0423_, _0425_);
  
  
  nand (_0427_, _0426_, _0426_);
  nand (_0428_, _0348_, _0427_);
  nand (_0429_, _0346_, _0426_);
  nand (_0430_, _0428_, _0429_);
  
  
  nand (_0431_, _0430_, _0430_);
  nand (_0432_, _0414_, _0416_);
  nand (_0433_, _0418_, _0432_);
  
  
  nand (_0434_, _0433_, _0433_);
  nand (_0436_, _0431_, _0434_);
  nand (_0437_, _0418_, _0436_);
  
  
  nand (_0438_, _0437_, _0437_);
  nand (_0439_, _0331_, _0334_);
  nand (_0440_, _0337_, _0439_);
  
  
  nand (_0441_, _0440_, _0440_);
  nand (_0442_, _0437_, _0441_);
  nand (_0443_, _0423_, _0428_);
  
  
  nand (_0444_, _0443_, _0443_);
  nand (_0445_, _0350_, _0353_);
  nand (_0447_, _0355_, _0445_);
  
  
  nand (_0448_, _0447_, _0447_);
  nand (_0449_, _0443_, _0448_);
  
  
  nand (_0450_, _0449_, _0449_);
  nand (_0451_, _0444_, _0447_);
  nand (_0452_, _0449_, _0451_);
  
  
  nand (_0453_, _0452_, _0452_);
  nand (_0454_, _0438_, _0440_);
  nand (_0455_, _0442_, _0454_);
  
  
  nand (_0456_, _0455_, _0455_);
  nand (_0458_, _0453_, _0456_);
  nand (_0459_, _0442_, _0458_);
  
  
  nand (_0460_, _0459_, _0459_);
  nand (_0461_, _0371_, _0374_);
  nand (_0462_, _0376_, _0461_);
  
  
  nand (_0463_, _0462_, _0462_);
  nand (_0464_, _0459_, _0463_);
  nand (_0465_, _0460_, _0462_);
  nand (_0466_, _0464_, _0465_);
  
  
  nand (_0467_, _0466_, _0466_);
  nand (_0469_, _0450_, _0467_);
  nand (_0470_, _0464_, _0469_);
  
  
  nand (_0471_, _0470_, _0470_);
  nand (_0472_, _0385_, _0387_);
  nand (_0473_, _0389_, _0472_);
  
  
  nand (_0474_, _0473_, _0473_);
  nand (_0475_, _0470_, _0474_);
  nand (_0476_, a_3_, b_1_);
  
  
  nand (_0477_, _0476_, _0476_);
  nand (_0478_, a_3_, b_0_);
  nand (_0480_, _0404_, _0477_);
  nand (_0481_, a_2_, b_2_);
  
  
  nand (_0482_, _0481_, _0481_);
  nand (_0483_, _0403_, _0476_);
  nand (_0484_, _0480_, _0483_);
  
  
  nand (_0485_, _0484_, _0484_);
  nand (_0486_, _0482_, _0485_);
  nand (_0487_, _0480_, _0486_);
  
  
  nand (_0488_, _0487_, _0487_);
  nand (_0489_, _0406_, _0409_);
  nand (_0491_, _0411_, _0489_);
  
  
  nand (_0492_, _0491_, _0491_);
  nand (_0493_, _0487_, _0492_);
  nand (_0494_, a_0_, b_5_);
  
  
  nand (_0495_, _0494_, _0494_);
  nand (_0496_, a_1_, b_4_);
  
  
  nand (_0497_, _0496_, _0496_);
  nand (_0498_, a_1_, b_3_);
  nand (_0499_, _0422_, _0497_);
  nand (_0500_, _0421_, _0496_);
  nand (_0502_, _0499_, _0500_);
  
  
  nand (_0503_, _0502_, _0502_);
  nand (_0504_, _0495_, _0503_);
  nand (_0505_, _0494_, _0502_);
  nand (_0506_, _0504_, _0505_);
  
  
  nand (_0507_, _0506_, _0506_);
  nand (_0508_, _0488_, _0491_);
  nand (_0509_, _0493_, _0508_);
  
  
  nand (_0510_, _0509_, _0509_);
  nand (_0511_, _0507_, _0510_);
  nand (_0513_, _0493_, _0511_);
  
  
  nand (_0514_, _0513_, _0513_);
  nand (_0515_, _0430_, _0433_);
  nand (_0516_, _0436_, _0515_);
  
  
  nand (_0517_, _0516_, _0516_);
  nand (_0518_, _0513_, _0517_);
  nand (_0519_, _0499_, _0504_);
  
  
  nand (_0520_, _0519_, _0519_);
  nand (_0521_, a_0_, b_6_);
  
  
  nand (_0522_, _0521_, _0521_);
  nand (_0524_, _0519_, _0522_);
  
  
  nand (_0525_, _0524_, _0524_);
  nand (_0526_, _0520_, _0521_);
  nand (_0527_, _0524_, _0526_);
  
  
  nand (_0528_, _0527_, _0527_);
  nand (_0529_, _0514_, _0516_);
  nand (_0530_, _0518_, _0529_);
  
  
  nand (_0531_, _0530_, _0530_);
  nand (_0532_, _0528_, _0531_);
  nand (_0533_, _0518_, _0532_);
  
  
  nand (_0535_, _0533_, _0533_);
  nand (_0536_, _0452_, _0455_);
  nand (_0537_, _0458_, _0536_);
  
  
  nand (_0538_, _0537_, _0537_);
  nand (_0539_, _0533_, _0538_);
  nand (_0540_, _0535_, _0537_);
  nand (_0541_, _0539_, _0540_);
  
  
  nand (_0542_, _0541_, _0541_);
  nand (_0543_, _0525_, _0542_);
  nand (_0544_, _0539_, _0543_);
  
  
  nand (_0546_, _0544_, _0544_);
  nand (_0547_, _0449_, _0466_);
  nand (_0548_, _0469_, _0547_);
  
  
  nand (_0549_, _0548_, _0548_);
  nand (_0550_, _0544_, _0549_);
  nand (_0551_, a_2_, b_1_);
  nand (_0552_, a_2_, b_0_);
  
  
  nand (_0553_, _0552_, _0552_);
  nand (_0554_, _0477_, _0553_);
  nand (_0555_, a_1_, b_2_);
  
  
  nand (_0557_, _0555_, _0555_);
  nand (_0558_, _0478_, _0551_);
  nand (_0559_, _0554_, _0558_);
  
  
  nand (_0560_, _0559_, _0559_);
  nand (_0561_, _0557_, _0560_);
  nand (_0562_, _0554_, _0561_);
  
  
  nand (_0563_, _0562_, _0562_);
  nand (_0564_, _0481_, _0484_);
  nand (_0565_, _0486_, _0564_);
  
  
  nand (_0566_, _0565_, _0565_);
  nand (_0568_, _0562_, _0566_);
  nand (_0569_, a_0_, b_4_);
  nand (_0570_, a_0_, b_3_);
  
  
  nand (_0571_, _0570_, _0570_);
  nand (_0572_, _0497_, _0571_);
  
  
  nand (_0573_, _0572_, _0572_);
  nand (_0574_, _0498_, _0569_);
  nand (_0575_, _0572_, _0574_);
  
  
  nand (_0576_, _0575_, _0575_);
  nand (_0577_, _0563_, _0565_);
  nand (_0579_, _0568_, _0577_);
  
  
  nand (_0580_, _0579_, _0579_);
  nand (_0581_, _0576_, _0580_);
  nand (_0582_, _0568_, _0581_);
  
  
  nand (_0583_, _0582_, _0582_);
  nand (_0584_, _0506_, _0509_);
  nand (_0585_, _0511_, _0584_);
  
  
  nand (_0586_, _0585_, _0585_);
  nand (_0587_, _0582_, _0586_);
  nand (_0588_, _0583_, _0585_);
  nand (_0590_, _0587_, _0588_);
  
  
  nand (_0591_, _0590_, _0590_);
  nand (_0592_, _0573_, _0591_);
  nand (_0593_, _0587_, _0592_);
  
  
  nand (_0594_, _0593_, _0593_);
  nand (_0595_, _0527_, _0530_);
  nand (_0596_, _0532_, _0595_);
  
  
  nand (_0597_, _0596_, _0596_);
  nand (_0598_, _0593_, _0597_);
  
  
  nand (_0599_, _0598_, _0598_);
  nand (_0601_, _0524_, _0541_);
  nand (_0602_, _0543_, _0601_);
  
  
  nand (_0603_, _0602_, _0602_);
  nand (_0604_, _0599_, _0603_);
  nand (_0605_, _0598_, _0602_);
  nand (_0606_, _0604_, _0605_);
  
  
  nand (_0607_, _0606_, _0606_);
  nand (_0608_, a_1_, b_1_);
  
  
  nand (_0609_, _0608_, _0608_);
  nand (_0610_, a_1_, b_0_);
  nand (_0612_, _0553_, _0609_);
  nand (_0613_, a_0_, b_2_);
  
  
  nand (_0614_, _0613_, _0613_);
  nand (_0615_, _0552_, _0608_);
  nand (_0616_, _0612_, _0615_);
  
  
  nand (_0617_, _0616_, _0616_);
  nand (_0618_, _0614_, _0617_);
  nand (_0619_, _0612_, _0618_);
  
  
  nand (_0620_, _0619_, _0619_);
  nand (_0621_, _0555_, _0559_);
  nand (_0623_, _0561_, _0621_);
  
  
  nand (_0624_, _0623_, _0623_);
  nand (_0625_, _0619_, _0624_);
  nand (_0626_, _0620_, _0623_);
  nand (_0627_, _0625_, _0626_);
  
  
  nand (_0628_, _0627_, _0627_);
  nand (_0629_, _0571_, _0628_);
  nand (_0630_, _0625_, _0629_);
  
  
  nand (_0631_, _0630_, _0630_);
  nand (_0632_, _0575_, _0579_);
  nand (_0634_, _0581_, _0632_);
  
  
  nand (_0635_, _0634_, _0634_);
  nand (_0636_, _0630_, _0635_);
  
  
  nand (_0637_, _0636_, _0636_);
  nand (_0638_, _0572_, _0590_);
  nand (_0639_, _0592_, _0638_);
  
  
  nand (_0640_, _0639_, _0639_);
  nand (_0641_, _0637_, _0640_);
  
  
  nand (_0642_, _0641_, _0641_);
  nand (_0643_, _0594_, _0596_);
  nand (_0645_, _0598_, _0643_);
  
  
  nand (_0646_, _0645_, _0645_);
  nand (_0647_, _0642_, _0646_);
  nand (_0648_, a_0_, b_1_);
  nand (_0649_, a_0_, b_0_);
  
  
  nand (_0650_, _0649_, _0649_);
  nand (_0651_, _0609_, _0650_);
  
  
  nand (_0652_, _0651_, _0651_);
  nand (_0653_, _0613_, _0616_);
  nand (_0654_, _0618_, _0653_);
  
  
  nand (_0656_, _0654_, _0654_);
  nand (_0657_, _0652_, _0656_);
  
  
  nand (_0658_, _0657_, _0657_);
  nand (_0659_, _0570_, _0627_);
  nand (_0660_, _0629_, _0659_);
  
  
  nand (_0661_, _0660_, _0660_);
  nand (_0662_, _0658_, _0661_);
  
  
  nand (_0663_, _0662_, _0662_);
  nand (_0664_, _0631_, _0634_);
  nand (_0665_, _0636_, _0664_);
  
  
  nand (_0667_, _0665_, _0665_);
  nand (_0668_, _0663_, _0667_);
  
  
  nand (_0669_, _0668_, _0668_);
  nand (_0670_, _0636_, _0639_);
  nand (_0671_, _0641_, _0670_);
  
  
  nand (_0672_, _0671_, _0671_);
  nand (_0673_, _0669_, _0672_);
  
  
  nand (_0674_, _0673_, _0673_);
  nand (_0675_, _0641_, _0645_);
  nand (_0676_, _0647_, _0675_);
  
  
  nand (_0678_, _0676_, _0676_);
  nand (_0679_, _0674_, _0678_);
  nand (_0680_, _0647_, _0679_);
  
  
  nand (_0681_, _0680_, _0680_);
  nand (_0682_, _0607_, _0680_);
  nand (_0683_, _0604_, _0682_);
  
  
  nand (_0684_, _0683_, _0683_);
  nand (_0685_, _0546_, _0548_);
  nand (_0686_, _0550_, _0685_);
  
  
  nand (_0687_, _0686_, _0686_);
  nand (_0689_, _0683_, _0687_);
  nand (_0690_, _0550_, _0689_);
  
  
  nand (_0691_, _0690_, _0690_);
  nand (_0692_, _0471_, _0473_);
  nand (_0693_, _0475_, _0692_);
  
  
  nand (_0694_, _0693_, _0693_);
  nand (_0695_, _0690_, _0694_);
  nand (_0696_, _0475_, _0695_);
  
  
  nand (_0697_, _0696_, _0696_);
  nand (_0698_, _0399_, _0696_);
  nand (_0700_, _0396_, _0698_);
  
  
  nand (_0701_, _0700_, _0700_);
  nand (_0702_, _0301_, _0700_);
  nand (_0703_, _0298_, _0702_);
  
  
  nand (_0704_, _0703_, _0703_);
  nand (_0705_, _0209_, _0211_);
  nand (_0706_, _0213_, _0705_);
  
  
  nand (_0707_, _0706_, _0706_);
  nand (_0708_, _0703_, _0707_);
  nand (_0709_, _0213_, _0708_);
  
  
  nand (_0711_, _0709_, _0709_);
  nand (_0712_, _0139_, _0709_);
  nand (_0713_, _0138_, _0711_);
  nand (_0714_, _0139_, _0713_);
  nand (_0715_, _0138_, _0712_);
  nand (_0716_, _0076_, _0715_);
  nand (_0717_, _0065_, _0069_);
  
  
  nand (_0718_, _0717_, _0717_);
  nand (_0719_, _0012_, _0059_);
  
  
  nand (_0720_, _0719_, _0719_);
  nand (_0722_, _0054_, _0720_);
  nand (_0723_, _0055_, _0719_);
  nand (_0724_, _0722_, _0723_);
  nand (_0725_, _0054_, _0719_);
  nand (_0726_, _0718_, _0724_);
  nand (_0727_, _0725_, _0726_);
  nand (_0728_, _0073_, _0727_);
  
  
  nand (_0729_, _0728_, _0728_);
  nand (_0730_, _0716_, _0729_);
  
  
  nand (product_7_, _0730_, _0730_);
  nand (_0732_, _0075_, _0714_);
  nand (_0733_, _0716_, _0732_);
  nand (_0734_, _0138_, _0139_);
  
  
  nand (_0735_, _0734_, _0734_);
  nand (_0736_, _0709_, _0734_);
  nand (_0737_, _0711_, _0735_);
  nand (_0738_, _0736_, _0737_);
  
  
  nand (_0739_, _0738_, _0738_);
  nand (_0740_, _0704_, _0706_);
  nand (_0741_, _0708_, _0740_);
  
  
  nand (_0743_, _0741_, _0741_);
  nand (_0744_, _0300_, _0701_);
  nand (_0745_, _0702_, _0744_);
  
  
  nand (_0746_, _0745_, _0745_);
  nand (_0747_, _0398_, _0697_);
  nand (_0748_, _0698_, _0747_);
  
  
  nand (_0749_, _0748_, _0748_);
  nand (_0750_, _0691_, _0693_);
  nand (_0751_, _0695_, _0750_);
  
  
  nand (_0752_, _0751_, _0751_);
  nand (_0754_, _0684_, _0686_);
  nand (_0755_, _0689_, _0754_);
  
  
  nand (_0756_, _0755_, _0755_);
  nand (_0757_, _0606_, _0681_);
  nand (_0758_, _0682_, _0757_);
  
  
  nand (_0759_, _0758_, _0758_);
  nand (_0760_, _0755_, _0758_);
  
  
  nand (_0761_, _0760_, _0760_);
  nand (_0762_, _0751_, _0761_);
  
  
  nand (_0763_, _0762_, _0762_);
  nand (_0765_, _0748_, _0763_);
  
  
  nand (_0766_, _0765_, _0765_);
  nand (_0767_, _0745_, _0766_);
  
  
  nand (_0768_, _0767_, _0767_);
  nand (_0769_, _0741_, _0768_);
  
  
  nand (_0770_, _0769_, _0769_);
  nand (_0771_, _0739_, _0770_);
  
  
  nand (_0772_, _0771_, _0771_);
  nand (_0773_, _0733_, _0772_);
  nand (_0774_, _0730_, _0773_);
  nand (_0776_, _0756_, _0759_);
  
  
  nand (_0777_, _0776_, _0776_);
  nand (_0778_, _0752_, _0777_);
  
  
  nand (_0779_, _0778_, _0778_);
  nand (_0780_, _0749_, _0779_);
  
  
  nand (_0781_, _0780_, _0780_);
  nand (_0782_, _0746_, _0781_);
  
  
  nand (_0783_, _0782_, _0782_);
  nand (_0784_, _0743_, _0783_);
  
  
  nand (_0785_, _0784_, _0784_);
  nand (_0787_, _0738_, _0785_);
  nand (_0788_, product_7_, _0787_);
  nand (_0789_, _0650_, _0788_);
  nand (product_0_, _0774_, _0789_);
  nand (_0790_, _0610_, _0648_);
  nand (_0791_, _0651_, _0790_);
  
  
  nand (_0792_, _0791_, _0791_);
  nand (_0793_, _0788_, _0792_);
  nand (product_1_, _0774_, _0793_);
  nand (_0794_, _0651_, _0654_);
  nand (_0796_, _0657_, _0794_);
  
  
  nand (_0797_, _0796_, _0796_);
  nand (_0798_, _0788_, _0797_);
  nand (product_2_, _0774_, _0798_);
  nand (_0799_, _0657_, _0660_);
  nand (_0800_, _0662_, _0799_);
  
  
  nand (_0801_, _0800_, _0800_);
  nand (_0802_, _0788_, _0801_);
  nand (product_3_, _0774_, _0802_);
  nand (_0803_, _0662_, _0665_);
  nand (_0805_, _0668_, _0803_);
  
  
  nand (_0806_, _0805_, _0805_);
  nand (_0807_, _0788_, _0806_);
  nand (product_4_, _0774_, _0807_);
  nand (_0808_, _0668_, _0671_);
  nand (_0809_, _0673_, _0808_);
  
  
  nand (_0810_, _0809_, _0809_);
  nand (_0811_, _0788_, _0810_);
  nand (product_5_, _0774_, _0811_);
  nand (_0812_, _0673_, _0676_);
  nand (_0814_, _0679_, _0812_);
  
  
  nand (_0815_, _0814_, _0814_);
  nand (_0816_, _0788_, _0815_);
  nand (product_6_, _0774_, _0816_);
endmodule
