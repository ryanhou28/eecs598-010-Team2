// Benchmark "c1355" written by ABC on Sun Oct 29 19:31:50 2023

module c1355 (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41,
    G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
    G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
    G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
    G1354, G1355  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
    G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
    G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
    G1354, G1355;
  reg n621_lo, n624_lo, n627_lo, n630_lo, n633_lo, n636_lo, n639_lo,
    n642_lo, n645_lo, n648_lo, n651_lo, n654_lo, n657_lo, n660_lo, n663_lo,
    n666_lo, n669_lo, n672_lo, n675_lo, n678_lo, n681_lo, n684_lo, n687_lo,
    n690_lo, n693_lo, n696_lo, n699_lo, n702_lo, n705_lo, n708_lo, n711_lo,
    n714_lo, n717_lo, n720_lo, n723_lo, n726_lo, n729_lo, n732_lo, n735_lo,
    n738_lo, n741_lo, n744_lo, n747_lo, n750_lo, n753_lo, n756_lo, n759_lo,
    n762_lo, n765_lo, n768_lo, n771_lo, n774_lo, n777_lo, n780_lo, n783_lo,
    n786_lo, n789_lo, n792_lo, n795_lo, n798_lo, n801_lo, n804_lo, n807_lo,
    n810_lo, n813_lo, n816_lo, n819_lo, n822_lo, n825_lo, n828_lo, n831_lo,
    n834_lo, n837_lo, n840_lo, n843_lo, n846_lo, n849_lo, n852_lo, n855_lo,
    n858_lo, n861_lo, n864_lo, n867_lo, n870_lo, n873_lo, n876_lo, n879_lo,
    n882_lo, n885_lo, n888_lo, n891_lo, n894_lo, n897_lo, n900_lo, n903_lo,
    n906_lo, n909_lo, n912_lo, n915_lo, n918_lo, n921_lo, n924_lo, n927_lo,
    n930_lo, n933_lo, n936_lo, n939_lo, n942_lo, n945_lo, n948_lo, n951_lo,
    n954_lo, n957_lo, n960_lo, n963_lo, n966_lo, n969_lo, n972_lo, n975_lo,
    n978_lo, n981_lo, n984_lo, n987_lo, n990_lo, n993_lo, n996_lo, n999_lo,
    n1002_lo, n1005_lo, n1008_lo, n1011_lo, n1014_lo, n1017_lo, n1020_lo,
    n1023_lo, n1026_lo, n1029_lo, n1032_lo, n1035_lo, n1038_lo, n1041_lo,
    n1044_lo, n1047_lo, n1050_lo, n1053_lo, n1056_lo, n1059_lo, n1062_lo,
    n1065_lo, n1068_lo, n1071_lo, n1074_lo, n1077_lo, n1080_lo, n1083_lo,
    n1086_lo, n1089_lo, n1092_lo, n1095_lo, n1098_lo, n1101_lo, n1104_lo,
    n1107_lo, n1110_lo;
  wire new_G242_, new_G245_, new_G248_, new_G251_, new_G254_, new_G257_,
    new_G260_, new_G263_, new_G266_, new_G269_, new_G272_, new_G275_,
    new_G278_, new_G281_, new_G284_, new_G287_, new_G290_, new_G293_,
    new_G296_, new_G299_, new_G302_, new_G305_, new_G308_, new_G311_,
    new_G314_, new_G317_, new_G320_, new_G323_, new_G326_, new_G329_,
    new_G332_, new_G335_, new_G338_, new_G341_, new_G344_, new_G347_,
    new_G350_, new_G353_, new_G356_, new_G359_, new_G362_, new_G363_,
    new_G364_, new_G365_, new_G366_, new_G367_, new_G368_, new_G369_,
    new_G370_, new_G371_, new_G372_, new_G373_, new_G374_, new_G375_,
    new_G376_, new_G377_, new_G378_, new_G379_, new_G380_, new_G381_,
    new_G382_, new_G383_, new_G384_, new_G385_, new_G386_, new_G387_,
    new_G388_, new_G389_, new_G390_, new_G391_, new_G392_, new_G393_,
    new_G394_, new_G395_, new_G396_, new_G397_, new_G398_, new_G399_,
    new_G400_, new_G401_, new_G402_, new_G403_, new_G404_, new_G405_,
    new_G406_, new_G407_, new_G408_, new_G409_, new_G410_, new_G411_,
    new_G412_, new_G413_, new_G414_, new_G415_, new_G416_, new_G417_,
    new_G418_, new_G419_, new_G420_, new_G421_, new_G422_, new_G423_,
    new_G424_, new_G425_, new_G426_, new_G429_, new_G432_, new_G435_,
    new_G438_, new_G441_, new_G444_, new_G447_, new_G450_, new_G453_,
    new_G456_, new_G459_, new_G462_, new_G465_, new_G468_, new_G471_,
    new_G474_, new_G477_, new_G480_, new_G483_, new_G486_, new_G489_,
    new_G492_, new_G495_, new_G498_, new_G501_, new_G504_, new_G507_,
    new_G510_, new_G513_, new_G516_, new_G519_, new_G522_, new_G525_,
    new_G528_, new_G531_, new_G534_, new_G537_, new_G540_, new_G543_,
    new_G546_, new_G549_, new_G552_, new_G555_, new_G558_, new_G561_,
    new_G564_, new_G567_, new_G570_, new_G571_, new_G572_, new_G573_,
    new_G574_, new_G575_, new_G576_, new_G577_, new_G578_, new_G579_,
    new_G580_, new_G581_, new_G582_, new_G583_, new_G584_, new_G585_,
    new_G586_, new_G587_, new_G588_, new_G589_, new_G590_, new_G591_,
    new_G592_, new_G593_, new_G594_, new_G595_, new_G596_, new_G597_,
    new_G598_, new_G599_, new_G600_, new_G601_, new_G602_, new_G607_,
    new_G612_, new_G617_, new_G622_, new_G627_, new_G632_, new_G637_,
    new_G642_, new_G645_, new_G648_, new_G651_, new_G654_, new_G657_,
    new_G660_, new_G663_, new_G666_, new_G669_, new_G672_, new_G675_,
    new_G678_, new_G681_, new_G684_, new_G687_, new_G690_, new_G691_,
    new_G692_, new_G693_, new_G694_, new_G695_, new_G696_, new_G697_,
    new_G698_, new_G699_, new_G700_, new_G701_, new_G702_, new_G703_,
    new_G704_, new_G705_, new_G706_, new_G709_, new_G712_, new_G715_,
    new_G718_, new_G721_, new_G724_, new_G727_, new_G730_, new_G733_,
    new_G736_, new_G739_, new_G742_, new_G745_, new_G748_, new_G751_,
    new_G754_, new_G755_, new_G756_, new_G757_, new_G758_, new_G759_,
    new_G760_, new_G761_, new_G762_, new_G763_, new_G764_, new_G765_,
    new_G766_, new_G767_, new_G768_, new_G769_, new_G770_, new_G773_,
    new_G776_, new_G779_, new_G782_, new_G785_, new_G788_, new_G791_,
    new_G794_, new_G797_, new_G800_, new_G803_, new_G806_, new_G809_,
    new_G812_, new_G815_, new_G818_, new_G819_, new_G820_, new_G821_,
    new_G822_, new_G823_, new_G824_, new_G825_, new_G826_, new_G827_,
    new_G828_, new_G829_, new_G830_, new_G831_, new_G832_, new_G833_,
    new_G834_, new_G847_, new_G860_, new_G873_, new_G886_, new_G899_,
    new_G912_, new_G925_, new_G938_, new_G939_, new_G940_, new_G941_,
    new_G942_, new_G943_, new_G944_, new_G945_, new_G946_, new_G947_,
    new_G948_, new_G949_, new_G950_, new_G951_, new_G952_, new_G953_,
    new_G954_, new_G955_, new_G956_, new_G957_, new_G958_, new_G959_,
    new_G960_, new_G961_, new_G962_, new_G963_, new_G964_, new_G965_,
    new_G966_, new_G967_, new_G968_, new_G969_, new_G970_, new_G971_,
    new_G972_, new_G973_, new_G974_, new_G975_, new_G976_, new_G977_,
    new_G978_, new_G979_, new_G980_, new_G981_, new_G982_, new_G983_,
    new_G984_, new_G985_, new_G986_, new_G991_, new_G996_, new_G1001_,
    new_G1006_, new_G1011_, new_G1016_, new_G1021_, new_G1026_, new_G1031_,
    new_G1036_, new_G1039_, new_G1042_, new_G1045_, new_G1048_, new_G1051_,
    new_G1054_, new_G1057_, new_G1060_, new_G1063_, new_G1066_, new_G1069_,
    new_G1072_, new_G1075_, new_G1078_, new_G1081_, new_G1084_, new_G1087_,
    new_G1090_, new_G1093_, new_G1096_, new_G1099_, new_G1102_, new_G1105_,
    new_G1108_, new_G1111_, new_G1114_, new_G1117_, new_G1120_, new_G1123_,
    new_G1126_, new_G1129_, new_G1132_, new_G1135_, new_G1138_, new_G1141_,
    new_G1144_, new_G1147_, new_G1150_, new_G1153_, new_G1156_, new_G1159_,
    new_G1162_, new_G1165_, new_G1168_, new_G1171_, new_G1174_, new_G1177_,
    new_G1180_, new_G1183_, new_G1186_, new_G1189_, new_G1192_, new_G1195_,
    new_G1198_, new_G1201_, new_G1204_, new_G1207_, new_G1210_, new_G1213_,
    new_G1216_, new_G1219_, new_G1222_, new_G1225_, new_G1228_, new_G1229_,
    new_G1230_, new_G1231_, new_G1232_, new_G1233_, new_G1234_, new_G1235_,
    new_G1236_, new_G1237_, new_G1238_, new_G1239_, new_G1240_, new_G1241_,
    new_G1242_, new_G1243_, new_G1244_, new_G1245_, new_G1246_, new_G1247_,
    new_G1248_, new_G1249_, new_G1250_, new_G1251_, new_G1252_, new_G1253_,
    new_G1254_, new_G1255_, new_G1256_, new_G1257_, new_G1258_, new_G1259_,
    new_G1260_, new_G1261_, new_G1262_, new_G1263_, new_G1264_, new_G1265_,
    new_G1266_, new_G1267_, new_G1268_, new_G1269_, new_G1270_, new_G1271_,
    new_G1272_, new_G1273_, new_G1274_, new_G1275_, new_G1276_, new_G1277_,
    new_G1278_, new_G1279_, new_G1280_, new_G1281_, new_G1282_, new_G1283_,
    new_G1284_, new_G1285_, new_G1286_, new_G1287_, new_G1288_, new_G1289_,
    new_G1290_, new_G1291_, new_G1292_, new_G1293_, new_G1294_, new_G1295_,
    new_G1296_, new_G1297_, new_G1298_, new_G1299_, new_G1300_, new_G1301_,
    new_G1302_, new_G1303_, new_G1304_, new_G1305_, new_G1306_, new_G1307_,
    new_G1308_, new_G1309_, new_G1310_, new_G1311_, new_G1312_, new_G1313_,
    new_G1314_, new_G1315_, new_G1316_, new_G1317_, new_G1318_, new_G1319_,
    new_G1320_, new_G1321_, new_G1322_, new_G1323_, n621_li, n624_li,
    n627_li, n630_li, n633_li, n636_li, n639_li, n642_li, n645_li, n648_li,
    n651_li, n654_li, n657_li, n660_li, n663_li, n666_li, n669_li, n672_li,
    n675_li, n678_li, n681_li, n684_li, n687_li, n690_li, n693_li, n696_li,
    n699_li, n702_li, n705_li, n708_li, n711_li, n714_li, n717_li, n720_li,
    n723_li, n726_li, n729_li, n732_li, n735_li, n738_li, n741_li, n744_li,
    n747_li, n750_li, n753_li, n756_li, n759_li, n762_li, n765_li, n768_li,
    n771_li, n774_li, n777_li, n780_li, n783_li, n786_li, n789_li, n792_li,
    n795_li, n798_li, n801_li, n804_li, n807_li, n810_li, n813_li, n816_li,
    n819_li, n822_li, n825_li, n828_li, n831_li, n834_li, n837_li, n840_li,
    n843_li, n846_li, n849_li, n852_li, n855_li, n858_li, n861_li, n864_li,
    n867_li, n870_li, n873_li, n876_li, n879_li, n882_li, n885_li, n888_li,
    n891_li, n894_li, n897_li, n900_li, n903_li, n906_li, n909_li, n912_li,
    n915_li, n918_li, n921_li, n924_li, n927_li, n930_li, n933_li, n936_li,
    n939_li, n942_li, n945_li, n948_li, n951_li, n954_li, n957_li, n960_li,
    n963_li, n966_li, n969_li, n972_li, n975_li, n978_li, n981_li, n984_li,
    n987_li, n990_li, n993_li, n996_li, n999_li, n1002_li, n1005_li,
    n1008_li, n1011_li, n1014_li, n1017_li, n1020_li, n1023_li, n1026_li,
    n1029_li, n1032_li, n1035_li, n1038_li, n1041_li, n1044_li, n1047_li,
    n1050_li, n1053_li, n1056_li, n1059_li, n1062_li, n1065_li, n1068_li,
    n1071_li, n1074_li, n1077_li, n1080_li, n1083_li, n1086_li, n1089_li,
    n1092_li, n1095_li, n1098_li, n1101_li, n1104_li, n1107_li, n1110_li;
  assign new_G242_ = n1014_lo & n1110_lo;
  assign new_G245_ = n1026_lo & n1110_lo;
  assign new_G248_ = n1038_lo & n1110_lo;
  assign new_G251_ = n1050_lo & n1110_lo;
  assign new_G254_ = n1062_lo & n1110_lo;
  assign new_G257_ = n1074_lo & n1110_lo;
  assign new_G260_ = n1086_lo & n1110_lo;
  assign new_G263_ = n1098_lo & n1110_lo;
  assign new_G266_ = ~n630_lo | ~n642_lo;
  assign new_G269_ = ~n654_lo | ~n666_lo;
  assign new_G272_ = ~n678_lo | ~n690_lo;
  assign new_G275_ = ~n702_lo | ~n714_lo;
  assign new_G278_ = ~n726_lo | ~n738_lo;
  assign new_G281_ = ~n750_lo | ~n762_lo;
  assign new_G284_ = ~n774_lo | ~n786_lo;
  assign new_G287_ = ~n798_lo | ~n810_lo;
  assign new_G290_ = ~n822_lo | ~n834_lo;
  assign new_G293_ = ~n846_lo | ~n858_lo;
  assign new_G296_ = ~n870_lo | ~n882_lo;
  assign new_G299_ = ~n894_lo | ~n906_lo;
  assign new_G302_ = ~n918_lo | ~n930_lo;
  assign new_G305_ = ~n942_lo | ~n954_lo;
  assign new_G308_ = ~n966_lo | ~n978_lo;
  assign new_G311_ = ~n990_lo | ~n1002_lo;
  assign new_G314_ = ~n630_lo | ~n678_lo;
  assign new_G317_ = ~n726_lo | ~n774_lo;
  assign new_G320_ = ~n642_lo | ~n690_lo;
  assign new_G323_ = ~n738_lo | ~n786_lo;
  assign new_G326_ = ~n654_lo | ~n702_lo;
  assign new_G329_ = ~n750_lo | ~n798_lo;
  assign new_G332_ = ~n666_lo | ~n714_lo;
  assign new_G335_ = ~n762_lo | ~n810_lo;
  assign new_G338_ = ~n822_lo | ~n870_lo;
  assign new_G341_ = ~n918_lo | ~n966_lo;
  assign new_G344_ = ~n834_lo | ~n882_lo;
  assign new_G347_ = ~n930_lo | ~n978_lo;
  assign new_G350_ = ~n846_lo | ~n894_lo;
  assign new_G353_ = ~n942_lo | ~n990_lo;
  assign new_G356_ = ~n858_lo | ~n906_lo;
  assign new_G359_ = ~n954_lo | ~n1002_lo;
  assign new_G362_ = ~n630_lo | ~new_G266_;
  assign new_G363_ = ~n642_lo | ~new_G266_;
  assign new_G364_ = ~n654_lo | ~new_G269_;
  assign new_G365_ = ~n666_lo | ~new_G269_;
  assign new_G366_ = ~n678_lo | ~new_G272_;
  assign new_G367_ = ~n690_lo | ~new_G272_;
  assign new_G368_ = ~n702_lo | ~new_G275_;
  assign new_G369_ = ~n714_lo | ~new_G275_;
  assign new_G370_ = ~n726_lo | ~new_G278_;
  assign new_G371_ = ~n738_lo | ~new_G278_;
  assign new_G372_ = ~n750_lo | ~new_G281_;
  assign new_G373_ = ~n762_lo | ~new_G281_;
  assign new_G374_ = ~n774_lo | ~new_G284_;
  assign new_G375_ = ~n786_lo | ~new_G284_;
  assign new_G376_ = ~n798_lo | ~new_G287_;
  assign new_G377_ = ~n810_lo | ~new_G287_;
  assign new_G378_ = ~n822_lo | ~new_G290_;
  assign new_G379_ = ~n834_lo | ~new_G290_;
  assign new_G380_ = ~n846_lo | ~new_G293_;
  assign new_G381_ = ~n858_lo | ~new_G293_;
  assign new_G382_ = ~n870_lo | ~new_G296_;
  assign new_G383_ = ~n882_lo | ~new_G296_;
  assign new_G384_ = ~n894_lo | ~new_G299_;
  assign new_G385_ = ~n906_lo | ~new_G299_;
  assign new_G386_ = ~n918_lo | ~new_G302_;
  assign new_G387_ = ~n930_lo | ~new_G302_;
  assign new_G388_ = ~n942_lo | ~new_G305_;
  assign new_G389_ = ~n954_lo | ~new_G305_;
  assign new_G390_ = ~n966_lo | ~new_G308_;
  assign new_G391_ = ~n978_lo | ~new_G308_;
  assign new_G392_ = ~n990_lo | ~new_G311_;
  assign new_G393_ = ~n1002_lo | ~new_G311_;
  assign new_G394_ = ~n630_lo | ~new_G314_;
  assign new_G395_ = ~n678_lo | ~new_G314_;
  assign new_G396_ = ~n726_lo | ~new_G317_;
  assign new_G397_ = ~n774_lo | ~new_G317_;
  assign new_G398_ = ~n642_lo | ~new_G320_;
  assign new_G399_ = ~n690_lo | ~new_G320_;
  assign new_G400_ = ~n738_lo | ~new_G323_;
  assign new_G401_ = ~n786_lo | ~new_G323_;
  assign new_G402_ = ~n654_lo | ~new_G326_;
  assign new_G403_ = ~n702_lo | ~new_G326_;
  assign new_G404_ = ~n750_lo | ~new_G329_;
  assign new_G405_ = ~n798_lo | ~new_G329_;
  assign new_G406_ = ~n666_lo | ~new_G332_;
  assign new_G407_ = ~n714_lo | ~new_G332_;
  assign new_G408_ = ~n762_lo | ~new_G335_;
  assign new_G409_ = ~n810_lo | ~new_G335_;
  assign new_G410_ = ~n822_lo | ~new_G338_;
  assign new_G411_ = ~n870_lo | ~new_G338_;
  assign new_G412_ = ~n918_lo | ~new_G341_;
  assign new_G413_ = ~n966_lo | ~new_G341_;
  assign new_G414_ = ~n834_lo | ~new_G344_;
  assign new_G415_ = ~n882_lo | ~new_G344_;
  assign new_G416_ = ~n930_lo | ~new_G347_;
  assign new_G417_ = ~n978_lo | ~new_G347_;
  assign new_G418_ = ~n846_lo | ~new_G350_;
  assign new_G419_ = ~n894_lo | ~new_G350_;
  assign new_G420_ = ~n942_lo | ~new_G353_;
  assign new_G421_ = ~n990_lo | ~new_G353_;
  assign new_G422_ = ~n858_lo | ~new_G356_;
  assign new_G423_ = ~n906_lo | ~new_G356_;
  assign new_G424_ = ~n954_lo | ~new_G359_;
  assign new_G425_ = ~n1002_lo | ~new_G359_;
  assign new_G426_ = ~new_G362_ | ~new_G363_;
  assign new_G429_ = ~new_G364_ | ~new_G365_;
  assign new_G432_ = ~new_G366_ | ~new_G367_;
  assign new_G435_ = ~new_G368_ | ~new_G369_;
  assign new_G438_ = ~new_G370_ | ~new_G371_;
  assign new_G441_ = ~new_G372_ | ~new_G373_;
  assign new_G444_ = ~new_G374_ | ~new_G375_;
  assign new_G447_ = ~new_G376_ | ~new_G377_;
  assign new_G450_ = ~new_G378_ | ~new_G379_;
  assign new_G453_ = ~new_G380_ | ~new_G381_;
  assign new_G456_ = ~new_G382_ | ~new_G383_;
  assign new_G459_ = ~new_G384_ | ~new_G385_;
  assign new_G462_ = ~new_G386_ | ~new_G387_;
  assign new_G465_ = ~new_G388_ | ~new_G389_;
  assign new_G468_ = ~new_G390_ | ~new_G391_;
  assign new_G471_ = ~new_G392_ | ~new_G393_;
  assign new_G474_ = ~new_G394_ | ~new_G395_;
  assign new_G477_ = ~new_G396_ | ~new_G397_;
  assign new_G480_ = ~new_G398_ | ~new_G399_;
  assign new_G483_ = ~new_G400_ | ~new_G401_;
  assign new_G486_ = ~new_G402_ | ~new_G403_;
  assign new_G489_ = ~new_G404_ | ~new_G405_;
  assign new_G492_ = ~new_G406_ | ~new_G407_;
  assign new_G495_ = ~new_G408_ | ~new_G409_;
  assign new_G498_ = ~new_G410_ | ~new_G411_;
  assign new_G501_ = ~new_G412_ | ~new_G413_;
  assign new_G504_ = ~new_G414_ | ~new_G415_;
  assign new_G507_ = ~new_G416_ | ~new_G417_;
  assign new_G510_ = ~new_G418_ | ~new_G419_;
  assign new_G513_ = ~new_G420_ | ~new_G421_;
  assign new_G516_ = ~new_G422_ | ~new_G423_;
  assign new_G519_ = ~new_G424_ | ~new_G425_;
  assign new_G522_ = ~new_G426_ | ~new_G429_;
  assign new_G525_ = ~new_G432_ | ~new_G435_;
  assign new_G528_ = ~new_G438_ | ~new_G441_;
  assign new_G531_ = ~new_G444_ | ~new_G447_;
  assign new_G534_ = ~new_G450_ | ~new_G453_;
  assign new_G537_ = ~new_G456_ | ~new_G459_;
  assign new_G540_ = ~new_G462_ | ~new_G465_;
  assign new_G543_ = ~new_G468_ | ~new_G471_;
  assign new_G546_ = ~new_G474_ | ~new_G477_;
  assign new_G549_ = ~new_G480_ | ~new_G483_;
  assign new_G552_ = ~new_G486_ | ~new_G489_;
  assign new_G555_ = ~new_G492_ | ~new_G495_;
  assign new_G558_ = ~new_G498_ | ~new_G501_;
  assign new_G561_ = ~new_G504_ | ~new_G507_;
  assign new_G564_ = ~new_G510_ | ~new_G513_;
  assign new_G567_ = ~new_G516_ | ~new_G519_;
  assign new_G570_ = ~new_G426_ | ~new_G522_;
  assign new_G571_ = ~new_G429_ | ~new_G522_;
  assign new_G572_ = ~new_G432_ | ~new_G525_;
  assign new_G573_ = ~new_G435_ | ~new_G525_;
  assign new_G574_ = ~new_G438_ | ~new_G528_;
  assign new_G575_ = ~new_G441_ | ~new_G528_;
  assign new_G576_ = ~new_G444_ | ~new_G531_;
  assign new_G577_ = ~new_G447_ | ~new_G531_;
  assign new_G578_ = ~new_G450_ | ~new_G534_;
  assign new_G579_ = ~new_G453_ | ~new_G534_;
  assign new_G580_ = ~new_G456_ | ~new_G537_;
  assign new_G581_ = ~new_G459_ | ~new_G537_;
  assign new_G582_ = ~new_G462_ | ~new_G540_;
  assign new_G583_ = ~new_G465_ | ~new_G540_;
  assign new_G584_ = ~new_G468_ | ~new_G543_;
  assign new_G585_ = ~new_G471_ | ~new_G543_;
  assign new_G586_ = ~new_G474_ | ~new_G546_;
  assign new_G587_ = ~new_G477_ | ~new_G546_;
  assign new_G588_ = ~new_G480_ | ~new_G549_;
  assign new_G589_ = ~new_G483_ | ~new_G549_;
  assign new_G590_ = ~new_G486_ | ~new_G552_;
  assign new_G591_ = ~new_G489_ | ~new_G552_;
  assign new_G592_ = ~new_G492_ | ~new_G555_;
  assign new_G593_ = ~new_G495_ | ~new_G555_;
  assign new_G594_ = ~new_G498_ | ~new_G558_;
  assign new_G595_ = ~new_G501_ | ~new_G558_;
  assign new_G596_ = ~new_G504_ | ~new_G561_;
  assign new_G597_ = ~new_G507_ | ~new_G561_;
  assign new_G598_ = ~new_G510_ | ~new_G564_;
  assign new_G599_ = ~new_G513_ | ~new_G564_;
  assign new_G600_ = ~new_G516_ | ~new_G567_;
  assign new_G601_ = ~new_G519_ | ~new_G567_;
  assign new_G602_ = ~new_G570_ | ~new_G571_;
  assign new_G607_ = ~new_G572_ | ~new_G573_;
  assign new_G612_ = ~new_G574_ | ~new_G575_;
  assign new_G617_ = ~new_G576_ | ~new_G577_;
  assign new_G622_ = ~new_G578_ | ~new_G579_;
  assign new_G627_ = ~new_G580_ | ~new_G581_;
  assign new_G632_ = ~new_G582_ | ~new_G583_;
  assign new_G637_ = ~new_G584_ | ~new_G585_;
  assign new_G642_ = ~new_G586_ | ~new_G587_;
  assign new_G645_ = ~new_G588_ | ~new_G589_;
  assign new_G648_ = ~new_G590_ | ~new_G591_;
  assign new_G651_ = ~new_G592_ | ~new_G593_;
  assign new_G654_ = ~new_G594_ | ~new_G595_;
  assign new_G657_ = ~new_G596_ | ~new_G597_;
  assign new_G660_ = ~new_G598_ | ~new_G599_;
  assign new_G663_ = ~new_G600_ | ~new_G601_;
  assign new_G666_ = ~new_G602_ | ~new_G607_;
  assign new_G669_ = ~new_G612_ | ~new_G617_;
  assign new_G672_ = ~new_G602_ | ~new_G612_;
  assign new_G675_ = ~new_G607_ | ~new_G617_;
  assign new_G678_ = ~new_G622_ | ~new_G627_;
  assign new_G681_ = ~new_G632_ | ~new_G637_;
  assign new_G684_ = ~new_G622_ | ~new_G632_;
  assign new_G687_ = ~new_G627_ | ~new_G637_;
  assign new_G690_ = ~new_G602_ | ~new_G666_;
  assign new_G691_ = ~new_G607_ | ~new_G666_;
  assign new_G692_ = ~new_G612_ | ~new_G669_;
  assign new_G693_ = ~new_G617_ | ~new_G669_;
  assign new_G694_ = ~new_G602_ | ~new_G672_;
  assign new_G695_ = ~new_G612_ | ~new_G672_;
  assign new_G696_ = ~new_G607_ | ~new_G675_;
  assign new_G697_ = ~new_G617_ | ~new_G675_;
  assign new_G698_ = ~new_G622_ | ~new_G678_;
  assign new_G699_ = ~new_G627_ | ~new_G678_;
  assign new_G700_ = ~new_G632_ | ~new_G681_;
  assign new_G701_ = ~new_G637_ | ~new_G681_;
  assign new_G702_ = ~new_G622_ | ~new_G684_;
  assign new_G703_ = ~new_G632_ | ~new_G684_;
  assign new_G704_ = ~new_G627_ | ~new_G687_;
  assign new_G705_ = ~new_G637_ | ~new_G687_;
  assign new_G706_ = ~new_G690_ | ~new_G691_;
  assign new_G709_ = ~new_G692_ | ~new_G693_;
  assign new_G712_ = ~new_G694_ | ~new_G695_;
  assign new_G715_ = ~new_G696_ | ~new_G697_;
  assign new_G718_ = ~new_G698_ | ~new_G699_;
  assign new_G721_ = ~new_G700_ | ~new_G701_;
  assign new_G724_ = ~new_G702_ | ~new_G703_;
  assign new_G727_ = ~new_G704_ | ~new_G705_;
  assign new_G730_ = ~new_G242_ | ~new_G718_;
  assign new_G733_ = ~new_G245_ | ~new_G721_;
  assign new_G736_ = ~new_G248_ | ~new_G724_;
  assign new_G739_ = ~new_G251_ | ~new_G727_;
  assign new_G742_ = ~new_G254_ | ~new_G706_;
  assign new_G745_ = ~new_G257_ | ~new_G709_;
  assign new_G748_ = ~new_G260_ | ~new_G712_;
  assign new_G751_ = ~new_G263_ | ~new_G715_;
  assign new_G754_ = ~new_G242_ | ~new_G730_;
  assign new_G755_ = ~new_G718_ | ~new_G730_;
  assign new_G756_ = ~new_G245_ | ~new_G733_;
  assign new_G757_ = ~new_G721_ | ~new_G733_;
  assign new_G758_ = ~new_G248_ | ~new_G736_;
  assign new_G759_ = ~new_G724_ | ~new_G736_;
  assign new_G760_ = ~new_G251_ | ~new_G739_;
  assign new_G761_ = ~new_G727_ | ~new_G739_;
  assign new_G762_ = ~new_G254_ | ~new_G742_;
  assign new_G763_ = ~new_G706_ | ~new_G742_;
  assign new_G764_ = ~new_G257_ | ~new_G745_;
  assign new_G765_ = ~new_G709_ | ~new_G745_;
  assign new_G766_ = ~new_G260_ | ~new_G748_;
  assign new_G767_ = ~new_G712_ | ~new_G748_;
  assign new_G768_ = ~new_G263_ | ~new_G751_;
  assign new_G769_ = ~new_G715_ | ~new_G751_;
  assign new_G770_ = ~new_G754_ | ~new_G755_;
  assign new_G773_ = ~new_G756_ | ~new_G757_;
  assign new_G776_ = ~new_G758_ | ~new_G759_;
  assign new_G779_ = ~new_G760_ | ~new_G761_;
  assign new_G782_ = ~new_G762_ | ~new_G763_;
  assign new_G785_ = ~new_G764_ | ~new_G765_;
  assign new_G788_ = ~new_G766_ | ~new_G767_;
  assign new_G791_ = ~new_G768_ | ~new_G769_;
  assign new_G794_ = ~new_G642_ | ~new_G770_;
  assign new_G797_ = ~new_G645_ | ~new_G773_;
  assign new_G800_ = ~new_G648_ | ~new_G776_;
  assign new_G803_ = ~new_G651_ | ~new_G779_;
  assign new_G806_ = ~new_G654_ | ~new_G782_;
  assign new_G809_ = ~new_G657_ | ~new_G785_;
  assign new_G812_ = ~new_G660_ | ~new_G788_;
  assign new_G815_ = ~new_G663_ | ~new_G791_;
  assign new_G818_ = ~new_G642_ | ~new_G794_;
  assign new_G819_ = ~new_G770_ | ~new_G794_;
  assign new_G820_ = ~new_G645_ | ~new_G797_;
  assign new_G821_ = ~new_G773_ | ~new_G797_;
  assign new_G822_ = ~new_G648_ | ~new_G800_;
  assign new_G823_ = ~new_G776_ | ~new_G800_;
  assign new_G824_ = ~new_G651_ | ~new_G803_;
  assign new_G825_ = ~new_G779_ | ~new_G803_;
  assign new_G826_ = ~new_G654_ | ~new_G806_;
  assign new_G827_ = ~new_G782_ | ~new_G806_;
  assign new_G828_ = ~new_G657_ | ~new_G809_;
  assign new_G829_ = ~new_G785_ | ~new_G809_;
  assign new_G830_ = ~new_G660_ | ~new_G812_;
  assign new_G831_ = ~new_G788_ | ~new_G812_;
  assign new_G832_ = ~new_G663_ | ~new_G815_;
  assign new_G833_ = ~new_G791_ | ~new_G815_;
  assign new_G834_ = ~new_G818_ | ~new_G819_;
  assign new_G847_ = ~new_G820_ | ~new_G821_;
  assign new_G860_ = ~new_G822_ | ~new_G823_;
  assign new_G873_ = ~new_G824_ | ~new_G825_;
  assign new_G886_ = ~new_G828_ | ~new_G829_;
  assign new_G899_ = ~new_G832_ | ~new_G833_;
  assign new_G912_ = ~new_G830_ | ~new_G831_;
  assign new_G925_ = ~new_G826_ | ~new_G827_;
  assign new_G938_ = ~new_G834_;
  assign new_G939_ = ~new_G847_;
  assign new_G940_ = ~new_G860_;
  assign new_G941_ = ~new_G834_;
  assign new_G942_ = ~new_G847_;
  assign new_G943_ = ~new_G873_;
  assign new_G944_ = ~new_G834_;
  assign new_G945_ = ~new_G860_;
  assign new_G946_ = ~new_G873_;
  assign new_G947_ = ~new_G847_;
  assign new_G948_ = ~new_G860_;
  assign new_G949_ = ~new_G873_;
  assign new_G950_ = ~new_G886_;
  assign new_G951_ = ~new_G899_;
  assign new_G952_ = ~new_G886_;
  assign new_G953_ = ~new_G912_;
  assign new_G954_ = ~new_G925_;
  assign new_G955_ = ~new_G899_;
  assign new_G956_ = ~new_G925_;
  assign new_G957_ = ~new_G912_;
  assign new_G958_ = ~new_G925_;
  assign new_G959_ = ~new_G886_;
  assign new_G960_ = ~new_G912_;
  assign new_G961_ = ~new_G925_;
  assign new_G962_ = ~new_G886_;
  assign new_G963_ = ~new_G899_;
  assign new_G964_ = ~new_G925_;
  assign new_G965_ = ~new_G912_;
  assign new_G966_ = ~new_G899_;
  assign new_G967_ = ~new_G886_;
  assign new_G968_ = ~new_G912_;
  assign new_G969_ = ~new_G899_;
  assign new_G970_ = ~new_G847_;
  assign new_G971_ = ~new_G873_;
  assign new_G972_ = ~new_G847_;
  assign new_G973_ = ~new_G860_;
  assign new_G974_ = ~new_G834_;
  assign new_G975_ = ~new_G873_;
  assign new_G976_ = ~new_G834_;
  assign new_G977_ = ~new_G860_;
  assign new_G978_ = new_G873_ & new_G938_ & new_G939_ & new_G940_;
  assign new_G979_ = new_G943_ & new_G941_ & new_G942_ & new_G860_;
  assign new_G980_ = new_G946_ & new_G944_ & new_G847_ & new_G945_;
  assign new_G981_ = new_G949_ & new_G834_ & new_G947_ & new_G948_;
  assign new_G982_ = new_G899_ & new_G958_ & new_G959_ & new_G960_;
  assign new_G983_ = new_G963_ & new_G961_ & new_G962_ & new_G912_;
  assign new_G984_ = new_G966_ & new_G964_ & new_G886_ & new_G965_;
  assign new_G985_ = new_G969_ & new_G925_ & new_G967_ & new_G968_;
  assign new_G986_ = new_G981_ | new_G980_ | new_G978_ | new_G979_;
  assign new_G991_ = new_G985_ | new_G984_ | new_G982_ | new_G983_;
  assign new_G996_ = new_G951_ & new_G925_ & new_G950_ & new_G912_ & new_G986_;
  assign new_G1001_ = new_G899_ & new_G925_ & new_G952_ & new_G953_ & new_G986_;
  assign new_G1006_ = new_G955_ & new_G954_ & new_G886_ & new_G912_ & new_G986_;
  assign new_G1011_ = new_G899_ & new_G956_ & new_G886_ & new_G957_ & new_G986_;
  assign new_G1016_ = new_G971_ & new_G834_ & new_G970_ & new_G860_ & new_G991_;
  assign new_G1021_ = new_G873_ & new_G834_ & new_G972_ & new_G973_ & new_G991_;
  assign new_G1026_ = new_G975_ & new_G974_ & new_G847_ & new_G860_ & new_G991_;
  assign new_G1031_ = new_G873_ & new_G976_ & new_G847_ & new_G977_ & new_G991_;
  assign new_G1036_ = new_G834_ & new_G996_;
  assign new_G1039_ = new_G847_ & new_G996_;
  assign new_G1042_ = new_G860_ & new_G996_;
  assign new_G1045_ = new_G873_ & new_G996_;
  assign new_G1048_ = new_G834_ & new_G1001_;
  assign new_G1051_ = new_G847_ & new_G1001_;
  assign new_G1054_ = new_G860_ & new_G1001_;
  assign new_G1057_ = new_G873_ & new_G1001_;
  assign new_G1060_ = new_G834_ & new_G1006_;
  assign new_G1063_ = new_G847_ & new_G1006_;
  assign new_G1066_ = new_G860_ & new_G1006_;
  assign new_G1069_ = new_G873_ & new_G1006_;
  assign new_G1072_ = new_G834_ & new_G1011_;
  assign new_G1075_ = new_G847_ & new_G1011_;
  assign new_G1078_ = new_G860_ & new_G1011_;
  assign new_G1081_ = new_G873_ & new_G1011_;
  assign new_G1084_ = new_G925_ & new_G1016_;
  assign new_G1087_ = new_G886_ & new_G1016_;
  assign new_G1090_ = new_G912_ & new_G1016_;
  assign new_G1093_ = new_G899_ & new_G1016_;
  assign new_G1096_ = new_G925_ & new_G1021_;
  assign new_G1099_ = new_G886_ & new_G1021_;
  assign new_G1102_ = new_G912_ & new_G1021_;
  assign new_G1105_ = new_G899_ & new_G1021_;
  assign new_G1108_ = new_G925_ & new_G1026_;
  assign new_G1111_ = new_G886_ & new_G1026_;
  assign new_G1114_ = new_G912_ & new_G1026_;
  assign new_G1117_ = new_G899_ & new_G1026_;
  assign new_G1120_ = new_G925_ & new_G1031_;
  assign new_G1123_ = new_G886_ & new_G1031_;
  assign new_G1126_ = new_G912_ & new_G1031_;
  assign new_G1129_ = new_G899_ & new_G1031_;
  assign new_G1132_ = ~n630_lo | ~new_G1036_;
  assign new_G1135_ = ~n642_lo | ~new_G1039_;
  assign new_G1138_ = ~n654_lo | ~new_G1042_;
  assign new_G1141_ = ~n666_lo | ~new_G1045_;
  assign new_G1144_ = ~n678_lo | ~new_G1048_;
  assign new_G1147_ = ~n690_lo | ~new_G1051_;
  assign new_G1150_ = ~n702_lo | ~new_G1054_;
  assign new_G1153_ = ~n714_lo | ~new_G1057_;
  assign new_G1156_ = ~n726_lo | ~new_G1060_;
  assign new_G1159_ = ~n738_lo | ~new_G1063_;
  assign new_G1162_ = ~n750_lo | ~new_G1066_;
  assign new_G1165_ = ~n762_lo | ~new_G1069_;
  assign new_G1168_ = ~n774_lo | ~new_G1072_;
  assign new_G1171_ = ~n786_lo | ~new_G1075_;
  assign new_G1174_ = ~n798_lo | ~new_G1078_;
  assign new_G1177_ = ~n810_lo | ~new_G1081_;
  assign new_G1180_ = ~n822_lo | ~new_G1084_;
  assign new_G1183_ = ~n834_lo | ~new_G1087_;
  assign new_G1186_ = ~n846_lo | ~new_G1090_;
  assign new_G1189_ = ~n858_lo | ~new_G1093_;
  assign new_G1192_ = ~n870_lo | ~new_G1096_;
  assign new_G1195_ = ~n882_lo | ~new_G1099_;
  assign new_G1198_ = ~n894_lo | ~new_G1102_;
  assign new_G1201_ = ~n906_lo | ~new_G1105_;
  assign new_G1204_ = ~n918_lo | ~new_G1108_;
  assign new_G1207_ = ~n930_lo | ~new_G1111_;
  assign new_G1210_ = ~n942_lo | ~new_G1114_;
  assign new_G1213_ = ~n954_lo | ~new_G1117_;
  assign new_G1216_ = ~n966_lo | ~new_G1120_;
  assign new_G1219_ = ~n978_lo | ~new_G1123_;
  assign new_G1222_ = ~n990_lo | ~new_G1126_;
  assign new_G1225_ = ~n1002_lo | ~new_G1129_;
  assign new_G1228_ = ~n630_lo | ~new_G1132_;
  assign new_G1229_ = ~new_G1036_ | ~new_G1132_;
  assign new_G1230_ = ~n642_lo | ~new_G1135_;
  assign new_G1231_ = ~new_G1039_ | ~new_G1135_;
  assign new_G1232_ = ~n654_lo | ~new_G1138_;
  assign new_G1233_ = ~new_G1042_ | ~new_G1138_;
  assign new_G1234_ = ~n666_lo | ~new_G1141_;
  assign new_G1235_ = ~new_G1045_ | ~new_G1141_;
  assign new_G1236_ = ~n678_lo | ~new_G1144_;
  assign new_G1237_ = ~new_G1048_ | ~new_G1144_;
  assign new_G1238_ = ~n690_lo | ~new_G1147_;
  assign new_G1239_ = ~new_G1051_ | ~new_G1147_;
  assign new_G1240_ = ~n702_lo | ~new_G1150_;
  assign new_G1241_ = ~new_G1054_ | ~new_G1150_;
  assign new_G1242_ = ~n714_lo | ~new_G1153_;
  assign new_G1243_ = ~new_G1057_ | ~new_G1153_;
  assign new_G1244_ = ~n726_lo | ~new_G1156_;
  assign new_G1245_ = ~new_G1060_ | ~new_G1156_;
  assign new_G1246_ = ~n738_lo | ~new_G1159_;
  assign new_G1247_ = ~new_G1063_ | ~new_G1159_;
  assign new_G1248_ = ~n750_lo | ~new_G1162_;
  assign new_G1249_ = ~new_G1066_ | ~new_G1162_;
  assign new_G1250_ = ~n762_lo | ~new_G1165_;
  assign new_G1251_ = ~new_G1069_ | ~new_G1165_;
  assign new_G1252_ = ~n774_lo | ~new_G1168_;
  assign new_G1253_ = ~new_G1072_ | ~new_G1168_;
  assign new_G1254_ = ~n786_lo | ~new_G1171_;
  assign new_G1255_ = ~new_G1075_ | ~new_G1171_;
  assign new_G1256_ = ~n798_lo | ~new_G1174_;
  assign new_G1257_ = ~new_G1078_ | ~new_G1174_;
  assign new_G1258_ = ~n810_lo | ~new_G1177_;
  assign new_G1259_ = ~new_G1081_ | ~new_G1177_;
  assign new_G1260_ = ~n822_lo | ~new_G1180_;
  assign new_G1261_ = ~new_G1084_ | ~new_G1180_;
  assign new_G1262_ = ~n834_lo | ~new_G1183_;
  assign new_G1263_ = ~new_G1087_ | ~new_G1183_;
  assign new_G1264_ = ~n846_lo | ~new_G1186_;
  assign new_G1265_ = ~new_G1090_ | ~new_G1186_;
  assign new_G1266_ = ~n858_lo | ~new_G1189_;
  assign new_G1267_ = ~new_G1093_ | ~new_G1189_;
  assign new_G1268_ = ~n870_lo | ~new_G1192_;
  assign new_G1269_ = ~new_G1096_ | ~new_G1192_;
  assign new_G1270_ = ~n882_lo | ~new_G1195_;
  assign new_G1271_ = ~new_G1099_ | ~new_G1195_;
  assign new_G1272_ = ~n894_lo | ~new_G1198_;
  assign new_G1273_ = ~new_G1102_ | ~new_G1198_;
  assign new_G1274_ = ~n906_lo | ~new_G1201_;
  assign new_G1275_ = ~new_G1105_ | ~new_G1201_;
  assign new_G1276_ = ~n918_lo | ~new_G1204_;
  assign new_G1277_ = ~new_G1108_ | ~new_G1204_;
  assign new_G1278_ = ~n930_lo | ~new_G1207_;
  assign new_G1279_ = ~new_G1111_ | ~new_G1207_;
  assign new_G1280_ = ~n942_lo | ~new_G1210_;
  assign new_G1281_ = ~new_G1114_ | ~new_G1210_;
  assign new_G1282_ = ~n954_lo | ~new_G1213_;
  assign new_G1283_ = ~new_G1117_ | ~new_G1213_;
  assign new_G1284_ = ~n966_lo | ~new_G1216_;
  assign new_G1285_ = ~new_G1120_ | ~new_G1216_;
  assign new_G1286_ = ~n978_lo | ~new_G1219_;
  assign new_G1287_ = ~new_G1123_ | ~new_G1219_;
  assign new_G1288_ = ~n990_lo | ~new_G1222_;
  assign new_G1289_ = ~new_G1126_ | ~new_G1222_;
  assign new_G1290_ = ~n1002_lo | ~new_G1225_;
  assign new_G1291_ = ~new_G1129_ | ~new_G1225_;
  assign new_G1292_ = ~new_G1228_ | ~new_G1229_;
  assign new_G1293_ = ~new_G1230_ | ~new_G1231_;
  assign new_G1294_ = ~new_G1232_ | ~new_G1233_;
  assign new_G1295_ = ~new_G1234_ | ~new_G1235_;
  assign new_G1296_ = ~new_G1236_ | ~new_G1237_;
  assign new_G1297_ = ~new_G1238_ | ~new_G1239_;
  assign new_G1298_ = ~new_G1240_ | ~new_G1241_;
  assign new_G1299_ = ~new_G1242_ | ~new_G1243_;
  assign new_G1300_ = ~new_G1244_ | ~new_G1245_;
  assign new_G1301_ = ~new_G1246_ | ~new_G1247_;
  assign new_G1302_ = ~new_G1248_ | ~new_G1249_;
  assign new_G1303_ = ~new_G1250_ | ~new_G1251_;
  assign new_G1304_ = ~new_G1252_ | ~new_G1253_;
  assign new_G1305_ = ~new_G1254_ | ~new_G1255_;
  assign new_G1306_ = ~new_G1256_ | ~new_G1257_;
  assign new_G1307_ = ~new_G1258_ | ~new_G1259_;
  assign new_G1308_ = ~new_G1260_ | ~new_G1261_;
  assign new_G1309_ = ~new_G1262_ | ~new_G1263_;
  assign new_G1310_ = ~new_G1264_ | ~new_G1265_;
  assign new_G1311_ = ~new_G1266_ | ~new_G1267_;
  assign new_G1312_ = ~new_G1268_ | ~new_G1269_;
  assign new_G1313_ = ~new_G1270_ | ~new_G1271_;
  assign new_G1314_ = ~new_G1272_ | ~new_G1273_;
  assign new_G1315_ = ~new_G1274_ | ~new_G1275_;
  assign new_G1316_ = ~new_G1276_ | ~new_G1277_;
  assign new_G1317_ = ~new_G1278_ | ~new_G1279_;
  assign new_G1318_ = ~new_G1280_ | ~new_G1281_;
  assign new_G1319_ = ~new_G1282_ | ~new_G1283_;
  assign new_G1320_ = ~new_G1284_ | ~new_G1285_;
  assign new_G1321_ = ~new_G1286_ | ~new_G1287_;
  assign new_G1322_ = ~new_G1288_ | ~new_G1289_;
  assign new_G1323_ = ~new_G1290_ | ~new_G1291_;
  assign G1324 = ~new_G1292_;
  assign G1325 = ~new_G1293_;
  assign G1326 = ~new_G1294_;
  assign G1327 = ~new_G1295_;
  assign G1328 = ~new_G1296_;
  assign G1329 = ~new_G1297_;
  assign G1330 = ~new_G1298_;
  assign G1331 = ~new_G1299_;
  assign G1332 = ~new_G1300_;
  assign G1333 = ~new_G1301_;
  assign G1334 = ~new_G1302_;
  assign G1335 = ~new_G1303_;
  assign G1336 = ~new_G1304_;
  assign G1337 = ~new_G1305_;
  assign G1338 = ~new_G1306_;
  assign G1339 = ~new_G1307_;
  assign G1340 = ~new_G1308_;
  assign G1341 = ~new_G1309_;
  assign G1342 = ~new_G1310_;
  assign G1343 = ~new_G1311_;
  assign G1344 = ~new_G1312_;
  assign G1345 = ~new_G1313_;
  assign G1346 = ~new_G1314_;
  assign G1347 = ~new_G1315_;
  assign G1348 = ~new_G1316_;
  assign G1349 = ~new_G1317_;
  assign G1350 = ~new_G1318_;
  assign G1351 = ~new_G1319_;
  assign G1352 = ~new_G1320_;
  assign G1353 = ~new_G1321_;
  assign G1354 = ~new_G1322_;
  assign G1355 = ~new_G1323_;
  assign n621_li = G1;
  assign n624_li = n621_lo;
  assign n627_li = n624_lo;
  assign n630_li = n627_lo;
  assign n633_li = G2;
  assign n636_li = n633_lo;
  assign n639_li = n636_lo;
  assign n642_li = n639_lo;
  assign n645_li = G3;
  assign n648_li = n645_lo;
  assign n651_li = n648_lo;
  assign n654_li = n651_lo;
  assign n657_li = G4;
  assign n660_li = n657_lo;
  assign n663_li = n660_lo;
  assign n666_li = n663_lo;
  assign n669_li = G5;
  assign n672_li = n669_lo;
  assign n675_li = n672_lo;
  assign n678_li = n675_lo;
  assign n681_li = G6;
  assign n684_li = n681_lo;
  assign n687_li = n684_lo;
  assign n690_li = n687_lo;
  assign n693_li = G7;
  assign n696_li = n693_lo;
  assign n699_li = n696_lo;
  assign n702_li = n699_lo;
  assign n705_li = G8;
  assign n708_li = n705_lo;
  assign n711_li = n708_lo;
  assign n714_li = n711_lo;
  assign n717_li = G9;
  assign n720_li = n717_lo;
  assign n723_li = n720_lo;
  assign n726_li = n723_lo;
  assign n729_li = G10;
  assign n732_li = n729_lo;
  assign n735_li = n732_lo;
  assign n738_li = n735_lo;
  assign n741_li = G11;
  assign n744_li = n741_lo;
  assign n747_li = n744_lo;
  assign n750_li = n747_lo;
  assign n753_li = G12;
  assign n756_li = n753_lo;
  assign n759_li = n756_lo;
  assign n762_li = n759_lo;
  assign n765_li = G13;
  assign n768_li = n765_lo;
  assign n771_li = n768_lo;
  assign n774_li = n771_lo;
  assign n777_li = G14;
  assign n780_li = n777_lo;
  assign n783_li = n780_lo;
  assign n786_li = n783_lo;
  assign n789_li = G15;
  assign n792_li = n789_lo;
  assign n795_li = n792_lo;
  assign n798_li = n795_lo;
  assign n801_li = G16;
  assign n804_li = n801_lo;
  assign n807_li = n804_lo;
  assign n810_li = n807_lo;
  assign n813_li = G17;
  assign n816_li = n813_lo;
  assign n819_li = n816_lo;
  assign n822_li = n819_lo;
  assign n825_li = G18;
  assign n828_li = n825_lo;
  assign n831_li = n828_lo;
  assign n834_li = n831_lo;
  assign n837_li = G19;
  assign n840_li = n837_lo;
  assign n843_li = n840_lo;
  assign n846_li = n843_lo;
  assign n849_li = G20;
  assign n852_li = n849_lo;
  assign n855_li = n852_lo;
  assign n858_li = n855_lo;
  assign n861_li = G21;
  assign n864_li = n861_lo;
  assign n867_li = n864_lo;
  assign n870_li = n867_lo;
  assign n873_li = G22;
  assign n876_li = n873_lo;
  assign n879_li = n876_lo;
  assign n882_li = n879_lo;
  assign n885_li = G23;
  assign n888_li = n885_lo;
  assign n891_li = n888_lo;
  assign n894_li = n891_lo;
  assign n897_li = G24;
  assign n900_li = n897_lo;
  assign n903_li = n900_lo;
  assign n906_li = n903_lo;
  assign n909_li = G25;
  assign n912_li = n909_lo;
  assign n915_li = n912_lo;
  assign n918_li = n915_lo;
  assign n921_li = G26;
  assign n924_li = n921_lo;
  assign n927_li = n924_lo;
  assign n930_li = n927_lo;
  assign n933_li = G27;
  assign n936_li = n933_lo;
  assign n939_li = n936_lo;
  assign n942_li = n939_lo;
  assign n945_li = G28;
  assign n948_li = n945_lo;
  assign n951_li = n948_lo;
  assign n954_li = n951_lo;
  assign n957_li = G29;
  assign n960_li = n957_lo;
  assign n963_li = n960_lo;
  assign n966_li = n963_lo;
  assign n969_li = G30;
  assign n972_li = n969_lo;
  assign n975_li = n972_lo;
  assign n978_li = n975_lo;
  assign n981_li = G31;
  assign n984_li = n981_lo;
  assign n987_li = n984_lo;
  assign n990_li = n987_lo;
  assign n993_li = G32;
  assign n996_li = n993_lo;
  assign n999_li = n996_lo;
  assign n1002_li = n999_lo;
  assign n1005_li = G33;
  assign n1008_li = n1005_lo;
  assign n1011_li = n1008_lo;
  assign n1014_li = n1011_lo;
  assign n1017_li = G34;
  assign n1020_li = n1017_lo;
  assign n1023_li = n1020_lo;
  assign n1026_li = n1023_lo;
  assign n1029_li = G35;
  assign n1032_li = n1029_lo;
  assign n1035_li = n1032_lo;
  assign n1038_li = n1035_lo;
  assign n1041_li = G36;
  assign n1044_li = n1041_lo;
  assign n1047_li = n1044_lo;
  assign n1050_li = n1047_lo;
  assign n1053_li = G37;
  assign n1056_li = n1053_lo;
  assign n1059_li = n1056_lo;
  assign n1062_li = n1059_lo;
  assign n1065_li = G38;
  assign n1068_li = n1065_lo;
  assign n1071_li = n1068_lo;
  assign n1074_li = n1071_lo;
  assign n1077_li = G39;
  assign n1080_li = n1077_lo;
  assign n1083_li = n1080_lo;
  assign n1086_li = n1083_lo;
  assign n1089_li = G40;
  assign n1092_li = n1089_lo;
  assign n1095_li = n1092_lo;
  assign n1098_li = n1095_lo;
  assign n1101_li = G41;
  assign n1104_li = n1101_lo;
  assign n1107_li = n1104_lo;
  assign n1110_li = n1107_lo;
  always @ (posedge clock) begin
    n621_lo <= n621_li;
    n624_lo <= n624_li;
    n627_lo <= n627_li;
    n630_lo <= n630_li;
    n633_lo <= n633_li;
    n636_lo <= n636_li;
    n639_lo <= n639_li;
    n642_lo <= n642_li;
    n645_lo <= n645_li;
    n648_lo <= n648_li;
    n651_lo <= n651_li;
    n654_lo <= n654_li;
    n657_lo <= n657_li;
    n660_lo <= n660_li;
    n663_lo <= n663_li;
    n666_lo <= n666_li;
    n669_lo <= n669_li;
    n672_lo <= n672_li;
    n675_lo <= n675_li;
    n678_lo <= n678_li;
    n681_lo <= n681_li;
    n684_lo <= n684_li;
    n687_lo <= n687_li;
    n690_lo <= n690_li;
    n693_lo <= n693_li;
    n696_lo <= n696_li;
    n699_lo <= n699_li;
    n702_lo <= n702_li;
    n705_lo <= n705_li;
    n708_lo <= n708_li;
    n711_lo <= n711_li;
    n714_lo <= n714_li;
    n717_lo <= n717_li;
    n720_lo <= n720_li;
    n723_lo <= n723_li;
    n726_lo <= n726_li;
    n729_lo <= n729_li;
    n732_lo <= n732_li;
    n735_lo <= n735_li;
    n738_lo <= n738_li;
    n741_lo <= n741_li;
    n744_lo <= n744_li;
    n747_lo <= n747_li;
    n750_lo <= n750_li;
    n753_lo <= n753_li;
    n756_lo <= n756_li;
    n759_lo <= n759_li;
    n762_lo <= n762_li;
    n765_lo <= n765_li;
    n768_lo <= n768_li;
    n771_lo <= n771_li;
    n774_lo <= n774_li;
    n777_lo <= n777_li;
    n780_lo <= n780_li;
    n783_lo <= n783_li;
    n786_lo <= n786_li;
    n789_lo <= n789_li;
    n792_lo <= n792_li;
    n795_lo <= n795_li;
    n798_lo <= n798_li;
    n801_lo <= n801_li;
    n804_lo <= n804_li;
    n807_lo <= n807_li;
    n810_lo <= n810_li;
    n813_lo <= n813_li;
    n816_lo <= n816_li;
    n819_lo <= n819_li;
    n822_lo <= n822_li;
    n825_lo <= n825_li;
    n828_lo <= n828_li;
    n831_lo <= n831_li;
    n834_lo <= n834_li;
    n837_lo <= n837_li;
    n840_lo <= n840_li;
    n843_lo <= n843_li;
    n846_lo <= n846_li;
    n849_lo <= n849_li;
    n852_lo <= n852_li;
    n855_lo <= n855_li;
    n858_lo <= n858_li;
    n861_lo <= n861_li;
    n864_lo <= n864_li;
    n867_lo <= n867_li;
    n870_lo <= n870_li;
    n873_lo <= n873_li;
    n876_lo <= n876_li;
    n879_lo <= n879_li;
    n882_lo <= n882_li;
    n885_lo <= n885_li;
    n888_lo <= n888_li;
    n891_lo <= n891_li;
    n894_lo <= n894_li;
    n897_lo <= n897_li;
    n900_lo <= n900_li;
    n903_lo <= n903_li;
    n906_lo <= n906_li;
    n909_lo <= n909_li;
    n912_lo <= n912_li;
    n915_lo <= n915_li;
    n918_lo <= n918_li;
    n921_lo <= n921_li;
    n924_lo <= n924_li;
    n927_lo <= n927_li;
    n930_lo <= n930_li;
    n933_lo <= n933_li;
    n936_lo <= n936_li;
    n939_lo <= n939_li;
    n942_lo <= n942_li;
    n945_lo <= n945_li;
    n948_lo <= n948_li;
    n951_lo <= n951_li;
    n954_lo <= n954_li;
    n957_lo <= n957_li;
    n960_lo <= n960_li;
    n963_lo <= n963_li;
    n966_lo <= n966_li;
    n969_lo <= n969_li;
    n972_lo <= n972_li;
    n975_lo <= n975_li;
    n978_lo <= n978_li;
    n981_lo <= n981_li;
    n984_lo <= n984_li;
    n987_lo <= n987_li;
    n990_lo <= n990_li;
    n993_lo <= n993_li;
    n996_lo <= n996_li;
    n999_lo <= n999_li;
    n1002_lo <= n1002_li;
    n1005_lo <= n1005_li;
    n1008_lo <= n1008_li;
    n1011_lo <= n1011_li;
    n1014_lo <= n1014_li;
    n1017_lo <= n1017_li;
    n1020_lo <= n1020_li;
    n1023_lo <= n1023_li;
    n1026_lo <= n1026_li;
    n1029_lo <= n1029_li;
    n1032_lo <= n1032_li;
    n1035_lo <= n1035_li;
    n1038_lo <= n1038_li;
    n1041_lo <= n1041_li;
    n1044_lo <= n1044_li;
    n1047_lo <= n1047_li;
    n1050_lo <= n1050_li;
    n1053_lo <= n1053_li;
    n1056_lo <= n1056_li;
    n1059_lo <= n1059_li;
    n1062_lo <= n1062_li;
    n1065_lo <= n1065_li;
    n1068_lo <= n1068_li;
    n1071_lo <= n1071_li;
    n1074_lo <= n1074_li;
    n1077_lo <= n1077_li;
    n1080_lo <= n1080_li;
    n1083_lo <= n1083_li;
    n1086_lo <= n1086_li;
    n1089_lo <= n1089_li;
    n1092_lo <= n1092_li;
    n1095_lo <= n1095_li;
    n1098_lo <= n1098_li;
    n1101_lo <= n1101_li;
    n1104_lo <= n1104_li;
    n1107_lo <= n1107_li;
    n1110_lo <= n1110_li;
  end
  initial begin
    n621_lo <= 1'b0;
    n624_lo <= 1'b0;
    n627_lo <= 1'b0;
    n630_lo <= 1'b0;
    n633_lo <= 1'b0;
    n636_lo <= 1'b0;
    n639_lo <= 1'b0;
    n642_lo <= 1'b0;
    n645_lo <= 1'b0;
    n648_lo <= 1'b0;
    n651_lo <= 1'b0;
    n654_lo <= 1'b0;
    n657_lo <= 1'b0;
    n660_lo <= 1'b0;
    n663_lo <= 1'b0;
    n666_lo <= 1'b0;
    n669_lo <= 1'b0;
    n672_lo <= 1'b0;
    n675_lo <= 1'b0;
    n678_lo <= 1'b0;
    n681_lo <= 1'b0;
    n684_lo <= 1'b0;
    n687_lo <= 1'b0;
    n690_lo <= 1'b0;
    n693_lo <= 1'b0;
    n696_lo <= 1'b0;
    n699_lo <= 1'b0;
    n702_lo <= 1'b0;
    n705_lo <= 1'b0;
    n708_lo <= 1'b0;
    n711_lo <= 1'b0;
    n714_lo <= 1'b0;
    n717_lo <= 1'b0;
    n720_lo <= 1'b0;
    n723_lo <= 1'b0;
    n726_lo <= 1'b0;
    n729_lo <= 1'b0;
    n732_lo <= 1'b0;
    n735_lo <= 1'b0;
    n738_lo <= 1'b0;
    n741_lo <= 1'b0;
    n744_lo <= 1'b0;
    n747_lo <= 1'b0;
    n750_lo <= 1'b0;
    n753_lo <= 1'b0;
    n756_lo <= 1'b0;
    n759_lo <= 1'b0;
    n762_lo <= 1'b0;
    n765_lo <= 1'b0;
    n768_lo <= 1'b0;
    n771_lo <= 1'b0;
    n774_lo <= 1'b0;
    n777_lo <= 1'b0;
    n780_lo <= 1'b0;
    n783_lo <= 1'b0;
    n786_lo <= 1'b0;
    n789_lo <= 1'b0;
    n792_lo <= 1'b0;
    n795_lo <= 1'b0;
    n798_lo <= 1'b0;
    n801_lo <= 1'b0;
    n804_lo <= 1'b0;
    n807_lo <= 1'b0;
    n810_lo <= 1'b0;
    n813_lo <= 1'b0;
    n816_lo <= 1'b0;
    n819_lo <= 1'b0;
    n822_lo <= 1'b0;
    n825_lo <= 1'b0;
    n828_lo <= 1'b0;
    n831_lo <= 1'b0;
    n834_lo <= 1'b0;
    n837_lo <= 1'b0;
    n840_lo <= 1'b0;
    n843_lo <= 1'b0;
    n846_lo <= 1'b0;
    n849_lo <= 1'b0;
    n852_lo <= 1'b0;
    n855_lo <= 1'b0;
    n858_lo <= 1'b0;
    n861_lo <= 1'b0;
    n864_lo <= 1'b0;
    n867_lo <= 1'b0;
    n870_lo <= 1'b0;
    n873_lo <= 1'b0;
    n876_lo <= 1'b0;
    n879_lo <= 1'b0;
    n882_lo <= 1'b0;
    n885_lo <= 1'b0;
    n888_lo <= 1'b0;
    n891_lo <= 1'b0;
    n894_lo <= 1'b0;
    n897_lo <= 1'b0;
    n900_lo <= 1'b0;
    n903_lo <= 1'b0;
    n906_lo <= 1'b0;
    n909_lo <= 1'b0;
    n912_lo <= 1'b0;
    n915_lo <= 1'b0;
    n918_lo <= 1'b0;
    n921_lo <= 1'b0;
    n924_lo <= 1'b0;
    n927_lo <= 1'b0;
    n930_lo <= 1'b0;
    n933_lo <= 1'b0;
    n936_lo <= 1'b0;
    n939_lo <= 1'b0;
    n942_lo <= 1'b0;
    n945_lo <= 1'b0;
    n948_lo <= 1'b0;
    n951_lo <= 1'b0;
    n954_lo <= 1'b0;
    n957_lo <= 1'b0;
    n960_lo <= 1'b0;
    n963_lo <= 1'b0;
    n966_lo <= 1'b0;
    n969_lo <= 1'b0;
    n972_lo <= 1'b0;
    n975_lo <= 1'b0;
    n978_lo <= 1'b0;
    n981_lo <= 1'b0;
    n984_lo <= 1'b0;
    n987_lo <= 1'b0;
    n990_lo <= 1'b0;
    n993_lo <= 1'b0;
    n996_lo <= 1'b0;
    n999_lo <= 1'b0;
    n1002_lo <= 1'b0;
    n1005_lo <= 1'b0;
    n1008_lo <= 1'b0;
    n1011_lo <= 1'b0;
    n1014_lo <= 1'b0;
    n1017_lo <= 1'b0;
    n1020_lo <= 1'b0;
    n1023_lo <= 1'b0;
    n1026_lo <= 1'b0;
    n1029_lo <= 1'b0;
    n1032_lo <= 1'b0;
    n1035_lo <= 1'b0;
    n1038_lo <= 1'b0;
    n1041_lo <= 1'b0;
    n1044_lo <= 1'b0;
    n1047_lo <= 1'b0;
    n1050_lo <= 1'b0;
    n1053_lo <= 1'b0;
    n1056_lo <= 1'b0;
    n1059_lo <= 1'b0;
    n1062_lo <= 1'b0;
    n1065_lo <= 1'b0;
    n1068_lo <= 1'b0;
    n1071_lo <= 1'b0;
    n1074_lo <= 1'b0;
    n1077_lo <= 1'b0;
    n1080_lo <= 1'b0;
    n1083_lo <= 1'b0;
    n1086_lo <= 1'b0;
    n1089_lo <= 1'b0;
    n1092_lo <= 1'b0;
    n1095_lo <= 1'b0;
    n1098_lo <= 1'b0;
    n1101_lo <= 1'b0;
    n1104_lo <= 1'b0;
    n1107_lo <= 1'b0;
    n1110_lo <= 1'b0;
  end
endmodule


