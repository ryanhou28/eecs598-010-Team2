`include "shift_reg_mem.sv"


module testbench;

    // Clock
    logic clock;

    // Define inputs
    logic signed [7:0] input_fmap;
    logic [4:0] mem_addr;
    logic signed [7:0] input_weights [31:0];
    logic enable;
    logic acc_reset;

    // Define outputs
    logic signed [7:0] output_fmap [31:0];

    // --- MEM ---
    // Define inputs to the ifmap buffer
    logic signed [7:0] ifmap_write_data [31:0];
    logic ifmap_write_enable;

    logic signed [7:0] mem_write_data [31:0];
    logic mem_write_enable;
    logic mem_reset;

    // Choose which data to write to the memory
    assign mem_write_data = (ifmap_write_enable) ? ifmap_write_data : output_fmap;

    // Instantiate the shift register memories
    shift_reg_mem shiftmem(
        .write_data(mem_write_data),
        .write_enable(mem_write_enable),
        .clk(clock),
        .reset(mem_reset),
        .read_data(input_fmap),
        .addr(mem_addr)
    );

    // Instantiate the accelerator
    accelerator accelerator1(
        .input_fmap(input_fmap),
        .input_weights(input_weights),
        .enable(enable),
        .reset(acc_reset),
        .clk(clock),
        .output_fmap(output_fmap)
    );
    
    
    always begin
        #5;
        clock=~clock;
    end

    // Define the input feature map
    localparam signed [7:0] input_nums [31:0] = '{-8, -5, 8, 0, 8, 7, -2, 7, 9, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0};

    // Define the NN Weights
    localparam signed [7:0] layer1_weights [31:0][31:0] = '{
        {2,-1,-2,1,2,-5,0,2,-1,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-4,0,-1,-4,4,3,-1,-3,-3,4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{2,-2,-5,1,-2,-2,2,-5,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{4,1,-4,-1,-3,-2,0,-5,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,-1,4,-4,-4,-3,0,-2,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-5,4,2,-1,-1,-2,2,-3,-4,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-4,0,-1,-2,-2,-2,-4,2,3,-5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-5,2,0,-4,3,4,1,0,-4,-3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-4,-4,-5,-1,3,3,-1,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{2,4,-1,-1,2,-4,3,-1,-3,-3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
    };

    localparam signed [7:0] layer2_weights [31:0][31:0] = '{
        {-2,3,1,-3,0,-4,1,1,3,-5,-2,-3,4,-5,-1,-2,-3,4,2,1,0,0,0,0,0,0,0,0,0,0,0,0},{1,3,-5,4,-2,1,-1,-5,-1,-3,-4,-1,1,-1,-4,0,-3,0,3,-2,0,0,0,0,0,0,0,0,0,0,0,0},{-3,2,-2,4,-5,4,-2,-1,-2,3,0,4,-3,-4,-4,-3,-3,-4,4,-2,0,0,0,0,0,0,0,0,0,0,0,0},{-1,2,1,0,0,-5,1,1,4,-5,-3,3,2,3,3,-4,0,4,4,0,0,0,0,0,0,0,0,0,0,0,0,0},{3,-2,4,0,-2,-2,-4,-4,3,-5,0,-2,-5,1,4,0,-2,2,0,1,0,0,0,0,0,0,0,0,0,0,0,0},{-4,-4,4,-4,3,4,4,-4,-2,-3,-2,-5,-5,-1,2,3,0,1,-5,-1,0,0,0,0,0,0,0,0,0,0,0,0},{-5,-3,-4,2,4,-2,3,-1,-1,-2,4,2,4,-2,-4,0,-1,0,2,4,0,0,0,0,0,0,0,0,0,0,0,0},{-4,2,3,3,-5,-4,3,0,-2,4,1,2,-4,0,-5,0,3,-2,-2,4,0,0,0,0,0,0,0,0,0,0,0,0},{-3,-1,-5,-1,-3,4,-4,-2,1,-1,3,-5,-1,2,1,-3,4,-1,-1,2,0,0,0,0,0,0,0,0,0,0,0,0},{-3,4,3,-2,2,-2,1,-4,1,-3,1,-5,2,0,-2,-2,2,-4,4,-4,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
    };

    localparam signed [7:0] layer3_weights [31:0][31:0] = '{
        {0,-1,0,1,1,-4,1,1,4,1,0,-4,1,4,4,-4,-3,1,4,3,3,-2,1,1,4,4,2,-5,2,-4,3,1},{1,-4,2,2,-5,-1,2,4,-1,3,1,-4,-3,0,-1,4,3,4,-4,-1,-5,2,2,2,0,2,1,-5,-2,4,0,-2},{4,4,-3,3,2,-2,-2,-5,2,-4,-3,-2,3,-3,1,-4,-5,3,4,1,4,2,1,4,-1,-4,-1,-2,-3,2,-1,2},{-3,3,-2,-1,-5,-1,4,-3,0,-1,-5,0,-1,-1,4,-4,-1,0,4,-5,-4,-5,3,2,-3,0,0,-2,3,0,2,-1},{-5,3,0,-3,-1,-5,2,0,3,-3,-1,1,2,3,3,1,2,-3,-5,-1,2,2,3,4,-4,4,-3,0,-1,1,-4,-5},{-5,-3,3,-1,-2,-4,3,-3,1,-5,-4,4,1,3,-3,2,-1,1,1,3,2,-4,-2,4,2,4,-5,-2,2,4,0,0},{3,0,-1,-1,4,-1,2,4,1,0,0,-3,-1,0,2,2,-5,4,-2,2,-1,-3,0,1,-1,3,-4,-1,-5,2,2,-5},{-5,-2,3,-4,-4,-2,-4,-2,-3,2,4,1,-2,-1,-5,0,4,-2,-1,-5,4,3,-5,-2,4,-4,2,-1,3,2,-2,3},{0,-5,2,0,-2,4,-3,-4,1,4,2,-2,-1,-2,3,-3,4,-3,4,2,4,3,-2,-2,-4,3,0,1,4,3,-4,4},{-3,4,4,3,-4,4,4,-1,2,1,1,3,2,-3,3,-1,1,-2,-3,3,0,1,3,-3,3,2,-3,-4,3,-4,3,-5},{0,-5,2,4,1,1,1,-3,-5,3,-5,1,-4,-1,0,-1,4,1,2,2,-5,0,3,-1,-5,-3,3,2,0,-3,-1,-4},{-5,4,-3,-1,-4,4,-3,-4,-1,-5,2,0,-5,-4,0,3,-4,4,2,-2,4,4,4,-2,2,4,-1,-2,-5,1,-1,-2},{0,3,-1,-3,2,0,0,-3,-5,4,4,2,0,1,3,-4,0,0,-2,-3,2,-2,-2,3,-1,-5,2,4,-4,-5,-2,-4},{-3,-4,-1,2,-4,0,1,0,2,3,-4,4,4,-5,-5,-1,-3,1,-2,1,2,3,3,1,3,-1,-4,-4,-5,3,3,-1},{-3,2,-3,-4,-2,-4,1,-5,0,-1,-5,-3,-3,-3,-4,1,0,-2,-3,-1,2,-4,-2,2,4,-1,-2,-4,3,-2,-5,-4},{3,-1,-5,3,1,2,-3,-2,-3,-5,-5,4,-2,-3,-3,0,1,1,3,3,1,0,-4,-2,4,-2,3,-2,-4,-5,2,-3},{0,2,0,-5,-3,4,3,-1,2,3,4,0,0,0,4,4,-2,3,4,1,-2,-4,-3,1,-1,-1,-2,1,-4,-4,-4,-4},{0,-5,2,-1,4,1,-5,4,2,4,0,-2,2,-4,-3,-1,2,0,0,1,1,-3,-2,2,-5,-2,1,-1,-1,-3,0,-4},{-3,-5,2,2,-2,2,-3,1,-4,3,3,0,-4,2,-3,-2,-5,-4,4,-5,1,-5,2,4,-2,-3,3,-2,-5,-1,0,-2},{-1,1,3,3,3,0,-1,4,1,1,-4,-2,-5,4,4,0,-1,4,0,-3,-5,-4,-1,4,-1,1,0,0,4,-5,-1,1},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
    };

    localparam signed [7:0] layer4_weights [31:0][31:0] = '{
        {-2,-2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-2,-2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{3,-4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-3,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,-5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-3,-3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{1,-4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{4,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-4,-2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{4,-2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-3,-4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{2,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{2,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-2,4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{4,-4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-4,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-1,-5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-5,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{2,-2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-1,-2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{0,-3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-4,-4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{3,-3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{3,4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{-3,-4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{1,-5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},{1,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
    };

    // Define a function for running the weights
    task run_nn ();
        $display("Setting input fmap");
        acc_reset = 0;
        mem_reset = 0;
        ifmap_write_enable = 1;
        mem_write_enable = 1;
        ifmap_write_data = input_nums;
        @(negedge clock);
        set_ifmap_zero();
        mem_write_enable = 0;
        ifmap_write_enable = 0;
        // Run layer 1
        // Enable the accelerator
        enable = 1;
        $display("Running layer 1");
        for (int i = 0; i < 32; i = i + 1) begin
            input_weights = layer1_weights[i];
            if (i == 31) begin
                mem_write_enable = 1;
            end
            @(negedge clock); 
        end
        // Run layer 2
        acc_reset = 1;
        mem_write_enable = 0;
        $display("Running layer 2");
        for (int i = 0; i < 32; i = i + 1) begin
            input_weights = layer2_weights[i];
            if (i == 31) begin
                mem_write_enable = 1;
            end
            @(negedge clock);
            acc_reset = 0;
        end
        // Run layer 3
        acc_reset = 1;
        mem_write_enable = 0;
        $display("Running layer 3");
        for (int i = 0; i < 32; i = i + 1) begin
            input_weights = layer3_weights[i];
            if (i == 31) begin
                mem_write_enable = 1;
            end
            @(negedge clock);
            acc_reset = 0;
        end
        // Run layer 4
        acc_reset = 1;
        mem_write_enable = 0;
        $display("Running layer 4");
        for (int i = 0; i < 32; i = i + 1) begin
            input_weights = layer4_weights[i];
            if (i == 31) begin
                mem_write_enable = 1;
            end
            @(negedge clock);
            acc_reset = 0;
        end
        mem_write_enable = 1;
        // Disable the accelerator
        $display("Inference Complete");
        // Display every output fmap
        for (int i = 0; i < 32; i = i + 1) begin
            $display("Output fmap [%d]: %d", i, output_fmap[i]);
        end
        @(negedge clock);
        mem_write_enable = 0;
        enable = 0;
        set_weights_zero();
        @(negedge clock);
    endtask

    task set_ifmap_zero();
        for (int i = 0; i < 32; i = i + 1) begin
            ifmap_write_data[0] = 0;
        end
    endtask

    task set_weights_zero();
        for (int i = 0; i < 32; i = i + 1) begin
            input_weights[0] = 0;
        end
    endtask

    initial begin
        $monitor("Time:%4.0f clock:%b enable:%b || mem_reset: %b mem_write_enable: %b | mem_write_data: [31]:%d, [30]: %d| mem_read_data: %d | mem_addr: %d || acc_reset: %b input_weights: [31]: %d, [30]: %d| output_fmap: [31]: %d, [30]: %d |",
                $time, clock, enable, mem_reset, mem_write_enable, mem_write_data[31], mem_write_data[30], input_fmap, mem_addr, acc_reset, input_weights[31], input_weights[30], output_fmap[31], output_fmap[30]);
        clock = 0;
        enable = 0;
        mem_reset = 1;
        acc_reset = 1;
        mem_write_enable = 0;
        ifmap_write_enable = 0;
        set_ifmap_zero();
        @(negedge clock);
        @(negedge clock);
        run_nn();
        @(negedge clock);
        @(negedge clock);
        @(negedge clock)

        // Run the test for some clock cycles
        for (int i = 0; i < 5; i = i + 1) begin
            @(negedge clock);
        end


        $finish;
    end

endmodule