module c1908(G1,G10,G11,G12,G13,G14,G15,G16,G17,G18,G1884,G1885,G1886,G1887,
  G1888,G1889,G1890,G1891,G1892,G1893,G1894,G1895,G1896,G1897,G1898,G1899,G19,
  G1900,G1901,G1902,G1903,G1904,G1905,G1906,G1907,G1908,G2,G20,G21,G22,G23,G24,
  G25,G26,G27,G28,G29,G3,G30,G31,G32,G33,G4,G5,G6,G7,G8,G9);
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
  G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33;
output G1884,G1885,G1886,G1887,G1888,G1889,G1890,G1891,G1892,G1893,G1894,G1895,
  G1896,G1897,G1898,G1899,G1900,G1901,G1902,G1903,G1904,G1905,G1906,G1907,
  G1908;

  wire G112,G116,G119,G123,G128,G131,G134,G138,G142,G147,G151,G154,G157,G161,
    G165,G169,G173,G174,G175,G178,G179,G182,G185,G188,G191,G194,G197,G198,G199,
    G202,G205,G212,G219,G222,G225,G228,G235,G238,G241,G248,G253,G260,G265,G268,
    G271,G274,G277,G280,G283,G286,G289,G292,G295,G298,G301,G304,G307,G310,G313,
    G314,G315,G316,G317,G318,G319,G320,G321,G322,G323,G324,G325,G326,G327,G328,
    G329,G330,G331,G332,G333,G334,G335,G338,G341,G344,G347,G350,G353,G356,G359,
    G362,G365,G368,G371,G374,G377,G380,G381,G382,G387,G391,G395,G398,G401,G404,
    G407,G410,G413,G416,G419,G422,G425,G428,G431,G434,G437,G440,G443,G446,G449,
    G452,G455,G458,G461,G464,G467,G470,G473,G476,G479,G482,G485,G488,G491,G494,
    G497,G500,G503,G506,G509,G512,G515,G518,G521,G524,G527,G530,G533,G534,G535,
    G536,G537,G538,G539,G540,G541,G542,G543,G544,G545,G546,G550,G554,G557,G560,
    G561,G562,G563,G564,G565,G566,G567,G568,G569,G570,G573,G582,G585,G586,G589,
    G590,G593,G594,G597,G598,G601,G602,G605,G606,G609,G612,G615,G616,G619,G620,
    G623,G624,G627,G628,G631,G632,G635,G636,G637,G638,G639,G640,G641,G644,G645,
    G648,G649,G650,G651,G652,G653,G654,G655,G656,G657,G660,G663,G666,G669,G672,
    G675,G678,G681,G684,G687,G690,G693,G696,G699,G700,G701,G702,G703,G704,G705,
    G706,G707,G708,G709,G710,G711,G712,G713,G714,G715,G716,G717,G718,G719,G720,
    G721,G722,G723,G724,G725,G726,G727,G728,G729,G730,G731,G734,G735,G738,G755,
    G772,G773,G774,G775,G776,G777,G778,G779,G780,G781,G782,G783,G784,G785,G786,
    G787,G788,G789,G790,G791,G792,G793,G794,G795,G796,G797,G798,G799,G802,G805,
    G806,G807,G808,G809,G810,G813,G816,G819,G822,G825,G828,G831,G834,G835,G836,
    G837,G838,G839,G840,G841,G842,G843,G844,G845,G848,G849,G850,G851,G854,G855,
    G856,G857,G858,G859,G860,G861,G864,G867,G870,G873,G876,G879,G882,G885,G888,
    G891,G894,G895,G896,G897,G898,G901,G904,G905,G906,G907,G908,G909,G910,G911,
    G914,G917,G918,G919,G920,G921,G924,G925,G926,G927,G928,G929,G930,G931,G932,
    G933,G934,G935,G936,G937,G938,G939,G940,G941,G942,G943,G944,G945,G946,G947,
    G948,G951,G952,G953,G956,G959,G962,G963,G964,G965,G966,G967,G968,G969,G970,
    G971,G972,G973,G974,G975,G976,G977,G980,G981,G984,G987,G988,G989,G993,G994,
    G995,G996,G997,G998,G999,G1000,G1003,G1006,G1009,G1012,G1015,G1019,G1022,
    G1023,G1024,G1025,G1028,G1031,G1034,G1035,G1036,G1037,G1038,G1041,G1044,
    G1047,G1050,G1053,G1056,G1059,G1062,G1065,G1066,G1067,G1068,G1069,G1072,
    G1075,G1078,G1081,G1084,G1087,G1090,G1091,G1092,G1093,G1094,G1095,G1096,
    G1097,G1098,G1099,G1100,G1103,G1104,G1107,G1110,G1111,G1112,G1113,G1114,
    G1115,G1116,G1117,G1118,G1121,G1124,G1125,G1126,G1129,G1130,G1131,G1132,
    G1135,G1138,G1139,G1140,G1143,G1144,G1145,G1148,G1151,G1152,G1153,G1154,
    G1155,G1156,G1157,G1158,G1159,G1160,G1163,G1166,G1167,G1168,G1169,G1170,
    G1171,G1174,G1175,G1176,G1177,G1178,G1181,G1182,G1185,G1186,G1187,G1188,
    G1189,G1192,G1195,G1198,G1199,G1200,G1201,G1202,G1203,G1204,G1205,G1208,
    G1209,G1212,G1215,G1216,G1217,G1218,G1219,G1220,G1221,G1222,G1225,G1226,
    G1227,G1230,G1233,G1236,G1239,G1240,G1243,G1244,G1245,G1246,G1247,G1250,
    G1251,G1252,G1253,G1256,G1259,G1260,G1261,G1262,G1263,G1264,G1265,G1266,
    G1267,G1268,G1269,G1270,G1273,G1276,G1279,G1280,G1281,G1282,G1283,G1284,
    G1287,G1290,G1293,G1296,G1299,G1302,G1305,G1308,G1309,G1310,G1311,G1312,
    G1313,G1316,G1317,G1320,G1321,G1322,G1323,G1324,G1325,G1326,G1327,G1328,
    G1329,G1330,G1331,G1332,G1333,G1334,G1335,G1336,G1337,G1338,G1339,G1340,
    G1341,G1342,G1343,G1344,G1347,G1350,G1353,G1354,G1355,G1356,G1357,G1358,
    G1359,G1362,G1363,G1366,G1369,G1370,G1371,G1374,G1375,G1378,G1381,G1382,
    G1383,G1386,G1389,G1392,G1395,G1410,G1420,G1434,G1439,G1442,G1445,G1448,
    G1451,G1454,G1457,G1458,G1459,G1460,G1461,G1462,G1463,G1464,G1465,G1466,
    G1467,G1468,G1469,G1470,G1471,G1472,G1473,G1474,G1475,G1476,G1479,G1480,
    G1483,G1484,G1487,G1488,G1489,G1490,G1493,G1496,G1499,G1502,G1505,G1508,
    G1511,G1522,G1538,G1549,G1563,G1576,G1584,G1598,G1607,G1608,G1609,G1624,
    G1625,G1642,G1645,G1648,G1651,G1654,G1657,G1660,G1663,G1666,G1669,G1672,
    G1675,G1678,G1681,G1684,G1687,G1690,G1693,G1696,G1699,G1702,G1705,G1708,
    G1711,G1712,G1713,G1714,G1715,G1716,G1717,G1718,G1719,G1722,G1725,G1728,
    G1731,G1734,G1737,G1740,G1743,G1746,G1747,G1748,G1749,G1750,G1751,G1752,
    G1753,G1754,G1755,G1756,G1757,G1758,G1759,G1760,G1761,G1762,G1763,G1764,
    G1765,G1766,G1767,G1768,G1769,G1770,G1771,G1772,G1773,G1774,G1775,G1776,
    G1777,G1778,G1779,G1780,G1781,G1782,G1783,G1784,G1785,G1786,G1787,G1788,
    G1791,G1794,G1795,G1796,G1797,G1798,G1799,G1800,G1801,G1802,G1803,G1806,
    G1809,G1810,G1817,G1818,G1819,G1820,G1821,G1822,G1825,G1828,G1831,G1834,
    G1837,G1838,G1839,G1842,G1845,G1848,G1849,G1850,G1851,G1852,G1853,G1854,
    G1855,G1856,G1857,G1858,G1859,G1860,G1861,G1862,G1863,G1864,G1865,G1866,
    G1867,G1868,G1869,G1870,G1871,G1872,G1873,G1874,G1875,G1876,G1877,G1880,
    G1881,G1882,G1883;

  not (G112,G1);
  not (G116,G2);
  not (G119,G3);
  not (G123,G4);
  not (G128,G5);
  not (G131,G6);
  not (G134,G7);
  not (G138,G8);
  not (G142,G9);
  not (G147,G10);
  not (G151,G11);
  not (G154,G12);
  not (G157,G13);
  not (G161,G14);
  not (G165,G15);
  not (G169,G16);
  nand (G173,G21,G29);
  nand (G174,G22,G30);
  not (G175,G24);
  not (G178,G24);
  not (G179,G23);
  not (G182,G23);
  not (G185,G25);
  not (G188,G26);
  not (G191,G27);
  not (G194,G28);
  not (G197,G33);
  not (G198,G33);
  not (G199,G29);
  not (G202,G30);
  not (G205,G31);
  not (G212,G31);
  not (G219,G31);
  not (G222,G31);
  not (G225,G32);
  not (G228,G32);
  not (G235,G32);
  not (G238,G33);
  not (G241,G33);
  not (G248,G33);
  not (G253,G33);
  not (G260,G33);
  not (G265,G1);
  not (G268,G2);
  not (G271,G3);
  not (G274,G4);
  not (G277,G5);
  not (G280,G6);
  not (G283,G7);
  not (G286,G8);
  not (G289,G9);
  not (G292,G10);
  not (G295,G11);
  not (G298,G12);
  not (G301,G13);
  not (G304,G14);
  not (G307,G15);
  not (G310,G16);
  not (G313,G265);
  not (G314,G268);
  not (G315,G271);
  not (G316,G274);
  not (G317,G277);
  not (G318,G280);
  not (G319,G283);
  not (G320,G286);
  not (G321,G289);
  not (G322,G292);
  not (G323,G295);
  not (G324,G298);
  not (G325,G301);
  not (G326,G304);
  not (G327,G307);
  not (G328,G310);
  nand (G329,G228,G253);
  nand (G330,G228,G253);
  nand (G331,G228,G253);
  nand (G332,G228,G253);
  nand (G333,G228,G253);
  nand (G334,G228,G253);
  not (G335,G112);
  not (G338,G116);
  not (G341,G128);
  not (G344,G131);
  not (G347,G147);
  not (G350,G165);
  and (G353,G21,G241);
  not (G356,G142);
  not (G359,G151);
  not (G362,G154);
  and (G365,G22,G241);
  not (G368,G161);
  and (G371,G17,G175,G241);
  not (G374,G169);
  not (G377,G161);
  nand (G380,G248,G199);
  nand (G381,G248,G202);
  nand (G382,G182,G24);
  nand (G387,G182,G222);
  nand (G391,G178,G222);
  not (G395,G123);
  not (G398,G138);
  not (G401,G142);
  not (G404,G161);
  not (G407,G112);
  not (G410,G112);
  not (G413,G116);
  not (G416,G151);
  not (G419,G119);
  and (G422,G19,G179,G241);
  not (G425,G154);
  not (G428,G123);
  not (G431,G157);
  and (G434,G20,G179,G241);
  not (G437,G185);
  not (G440,G185);
  not (G443,G188);
  not (G446,G188);
  not (G449,G191);
  not (G452,G191);
  not (G455,G194);
  not (G458,G194);
  and (G461,G173,G238);
  and (G464,G174,G238);
  not (G467,G119);
  not (G470,G119);
  not (G473,G134);
  not (G476,G134);
  not (G479,G169);
  not (G482,G169);
  not (G485,G157);
  not (G488,G157);
  not (G491,G123);
  not (G494,G123);
  not (G497,G128);
  not (G500,G138);
  and (G503,G18,G175,G241);
  not (G506,G165);
  not (G509,G142);
  not (G512,G142);
  not (G515,G131);
  not (G518,G138);
  not (G521,G147);
  not (G524,G165);
  not (G527,G134);
  not (G530,G147);
  not (G533,G461);
  not (G534,G464);
  not (G535,G395);
  not (G536,G398);
  not (G537,G401);
  not (G538,G404);
  not (G539,G410);
  not (G540,G422);
  not (G541,G428);
  not (G542,G431);
  not (G543,G434);
  and (G544,G17,G391);
  and (G545,G19,G387);
  nand (G546,G18,G391);
  nand (G550,G20,G387);
  nand (G554,G17,G391);
  nand (G557,G19,G387);
  not (G560,G440);
  not (G561,G437);
  not (G562,G446);
  not (G563,G443);
  not (G564,G452);
  not (G565,G449);
  not (G566,G458);
  not (G567,G455);
  nand (G568,G199,G219,G248,G382);
  nand (G569,G202,G219,G248,G382);
  nand (G570,G225,G260,G382);
  and (G573,G225,G260,G382);
  not (G582,G335);
  not (G585,G467);
  not (G586,G335);
  not (G589,G470);
  not (G590,G341);
  not (G593,G473);
  not (G594,G341);
  not (G597,G476);
  not (G598,G347);
  not (G601,G479);
  not (G602,G347);
  not (G605,G482);
  not (G606,G353);
  not (G609,G353);
  not (G612,G359);
  not (G615,G485);
  not (G616,G359);
  not (G619,G488);
  not (G620,G365);
  not (G623,G491);
  not (G624,G365);
  not (G627,G494);
  not (G628,G371);
  not (G631,G407);
  not (G632,G371);
  not (G635,G497);
  not (G636,G500);
  not (G637,G413);
  not (G638,G503);
  not (G639,G506);
  not (G640,G416);
  not (G641,G374);
  not (G644,G509);
  not (G645,G374);
  not (G648,G512);
  not (G649,G515);
  not (G650,G518);
  not (G651,G419);
  not (G652,G521);
  not (G653,G524);
  not (G654,G425);
  not (G655,G527);
  not (G656,G530);
  not (G657,G338);
  not (G660,G338);
  not (G663,G344);
  not (G666,G344);
  not (G669,G350);
  not (G672,G350);
  not (G675,G356);
  not (G678,G356);
  not (G681,G362);
  not (G684,G362);
  not (G687,G368);
  not (G690,G368);
  not (G693,G377);
  not (G696,G377);
  nand (G699,G398,G535);
  nand (G700,G395,G536);
  nand (G701,G404,G537);
  nand (G702,G401,G538);
  nand (G703,G434,G542);
  nand (G704,G431,G543);
  nand (G705,G500,G635);
  nand (G706,G497,G636);
  nand (G707,G506,G638);
  nand (G708,G503,G639);
  nand (G709,G518,G649);
  nand (G710,G515,G650);
  nand (G711,G524,G652);
  nand (G712,G521,G653);
  nand (G713,G530,G655);
  nand (G714,G527,G656);
  not (G715,G586);
  not (G716,G582);
  nand (G717,G699,G700);
  not (G718,G590);
  not (G719,G594);
  not (G720,G602);
  not (G721,G598);
  not (G722,G609);
  not (G723,G616);
  not (G724,G624);
  nand (G725,G701,G702);
  not (G726,G632);
  nand (G727,G632,G539);
  not (G728,G645);
  nand (G729,G703,G704);
  not (G730,G546);
  not (G731,G546);
  not (G734,G550);
  not (G735,G550);
  nand (G738,G568,G570);
  nand (G755,G569,G570);
  not (G772,G657);
  nand (G773,G657,G585);
  not (G774,G660);
  nand (G775,G660,G589);
  not (G776,G663);
  nand (G777,G663,G593);
  not (G778,G666);
  nand (G779,G666,G597);
  not (G780,G669);
  nand (G781,G669,G601);
  not (G782,G672);
  nand (G783,G672,G605);
  not (G784,G675);
  not (G785,G606);
  not (G786,G678);
  not (G787,G681);
  nand (G788,G681,G615);
  not (G789,G612);
  not (G790,G684);
  nand (G791,G684,G619);
  not (G792,G687);
  nand (G793,G687,G623);
  not (G794,G620);
  not (G795,G690);
  nand (G796,G690,G627);
  not (G797,G628);
  nand (G798,G628,G631);
  nand (G799,G705,G706);
  nand (G802,G707,G708);
  not (G805,G693);
  nand (G806,G693,G644);
  not (G807,G641);
  not (G808,G696);
  nand (G809,G696,G648);
  nand (G810,G709,G710);
  nand (G813,G711,G712);
  nand (G816,G713,G714);
  not (G819,G554);
  not (G822,G554);
  not (G825,G557);
  not (G828,G557);
  not (G831,G717);
  nand (G834,G410,G726);
  nand (G835,G467,G772);
  nand (G836,G470,G774);
  nand (G837,G473,G776);
  nand (G838,G476,G778);
  nand (G839,G479,G780);
  nand (G840,G482,G782);
  nand (G841,G485,G787);
  nand (G842,G488,G790);
  nand (G843,G491,G792);
  nand (G844,G494,G795);
  not (G845,G725);
  nand (G848,G407,G797);
  nand (G849,G509,G805);
  nand (G850,G512,G808);
  not (G851,G729);
  nand (G854,G834,G727);
  nand (G855,G816,G541);
  not (G856,G816);
  not (G857,G822);
  not (G858,G819);
  not (G859,G828);
  not (G860,G825);
  nand (G861,G835,G773);
  nand (G864,G836,G775);
  nand (G867,G837,G777);
  nand (G870,G838,G779);
  nand (G873,G839,G781);
  nand (G876,G840,G783);
  nand (G879,G841,G788);
  nand (G882,G842,G791);
  nand (G885,G843,G793);
  nand (G888,G844,G796);
  nand (G891,G848,G798);
  not (G894,G799);
  nand (G895,G799,G637);
  not (G896,G802);
  nand (G897,G802,G640);
  nand (G898,G849,G806);
  nand (G901,G850,G809);
  not (G904,G810);
  nand (G905,G810,G651);
  not (G906,G813);
  nand (G907,G813,G654);
  not (G908,G845);
  nand (G909,G428,G856);
  not (G910,G851);
  not (G911,G831);
  not (G914,G831);
  nand (G917,G413,G894);
  nand (G918,G416,G896);
  nand (G919,G419,G904);
  nand (G920,G425,G906);
  not (G921,G854);
  nand (G924,G864,G715);
  not (G925,G864);
  nand (G926,G861,G716);
  not (G927,G861);
  nand (G928,G867,G718);
  not (G929,G867);
  nand (G930,G870,G719);
  not (G931,G870);
  nand (G932,G876,G720);
  not (G933,G876);
  nand (G934,G873,G721);
  not (G935,G873);
  nand (G936,G882,G723);
  not (G937,G882);
  nand (G938,G888,G724);
  not (G939,G888);
  not (G940,G891);
  nand (G941,G901,G728);
  not (G942,G901);
  nand (G943,G855,G909);
  not (G944,G879);
  nand (G945,G879,G789);
  not (G946,G885);
  nand (G947,G885,G794);
  nand (G948,G895,G917);
  not (G951,G898);
  nand (G952,G898,G807);
  nand (G953,G897,G918);
  nand (G956,G907,G920);
  nand (G959,G905,G919);
  nand (G962,G586,G925);
  nand (G963,G582,G927);
  nand (G964,G590,G929);
  not (G965,G914);
  not (G966,G911);
  nand (G967,G594,G931);
  nand (G968,G602,G933);
  nand (G969,G598,G935);
  nand (G970,G616,G937);
  nand (G971,G624,G939);
  nand (G972,G645,G942);
  not (G973,G921);
  nand (G974,G612,G944);
  nand (G975,G620,G946);
  nand (G976,G641,G951);
  not (G977,G943);
  nand (G980,G924,G962);
  nand (G981,G926,G963);
  nand (G984,G928,G964);
  nand (G987,G930,G967);
  nand (G988,G932,G968);
  nand (G989,G934,G969);
  nand (G993,G936,G970);
  nand (G994,G938,G971);
  not (G995,G948);
  nand (G996,G941,G972);
  not (G997,G953);
  not (G998,G956);
  not (G999,G959);
  nand (G1000,G947,G975);
  nand (G1003,G945,G974);
  nand (G1006,G952,G976);
  not (G1009,G980);
  not (G1012,G988);
  not (G1015,G993);
  not (G1019,G987);
  nand (G1022,G959,G998);
  nand (G1023,G956,G999);
  not (G1024,G977);
  not (G1025,G994);
  not (G1028,G996);
  not (G1031,G989);
  not (G1034,G1000);
  not (G1035,G1003);
  nand (G1036,G1006,G997);
  not (G1037,G1006);
  nand (G1038,G1022,G1023);
  not (G1041,G984);
  not (G1044,G984);
  not (G1047,G989);
  not (G1050,G989);
  not (G1053,G981);
  not (G1056,G981);
  not (G1059,G1015);
  not (G1062,G1012);
  not (G1065,G1025);
  nand (G1066,G953,G1037);
  nand (G1067,G1028,G1024);
  not (G1068,G1028);
  not (G1069,G1019);
  not (G1072,G1019);
  not (G1075,G1009);
  not (G1078,G1009);
  not (G1081,G1012);
  not (G1084,G1015);
  not (G1087,G1015);
  nand (G1090,G1038,G540);
  not (G1091,G1038);
  not (G1092,G1041);
  not (G1093,G1044);
  nand (G1094,G1047,G784);
  not (G1095,G1047);
  nand (G1096,G1050,G786);
  not (G1097,G1050);
  not (G1098,G1053);
  not (G1099,G1056);
  nand (G1100,G1036,G1066);
  nand (G1103,G977,G1068);
  not (G1104,G1031);
  not (G1107,G1031);
  nand (G1110,G422,G1091);
  not (G1111,G1072);
  nand (G1112,G1075,G1092);
  not (G1113,G1075);
  nand (G1114,G1078,G1093);
  not (G1115,G1078);
  nand (G1116,G675,G1095);
  nand (G1117,G678,G1097);
  not (G1118,G1059);
  not (G1121,G1059);
  nand (G1124,G1081,G1035);
  not (G1125,G1081);
  nand (G1126,G1067,G1103);
  not (G1129,G1084);
  not (G1130,G1069);
  not (G1131,G1087);
  not (G1132,G1062);
  not (G1135,G1062);
  nand (G1138,G1100,G995);
  not (G1139,G1100);
  nand (G1140,G1090,G1110);
  nand (G1143,G1041,G1113);
  nand (G1144,G1044,G1115);
  nand (G1145,G1094,G1116);
  nand (G1148,G1096,G1117);
  nand (G1151,G1003,G1125);
  not (G1152,G1104);
  nand (G1153,G1104,G1129);
  not (G1154,G1107);
  nand (G1155,G1107,G1131);
  not (G1156,G1121);
  nand (G1157,G948,G1139);
  nand (G1158,G1126,G910);
  not (G1159,G1126);
  nand (G1160,G1112,G1143);
  nand (G1163,G1114,G1144);
  not (G1166,G1132);
  nand (G1167,G1132,G1098);
  not (G1168,G1118);
  not (G1169,G1135);
  nand (G1170,G1135,G1099);
  nand (G1171,G1124,G1151);
  nand (G1174,G1084,G1152);
  nand (G1175,G1087,G1154);
  nand (G1176,G1148,G722);
  not (G1177,G1148);
  nand (G1178,G1138,G1157);
  nand (G1181,G851,G1159);
  nand (G1182,G1140,G212);
  not (G1185,G1145);
  nand (G1186,G1145,G785);
  nand (G1187,G1053,G1166);
  nand (G1188,G1056,G1169);
  nand (G1189,G1174,G1153);
  nand (G1192,G1175,G1155);
  not (G1195,G1140);
  nand (G1198,G1163,G965);
  not (G1199,G1163);
  nand (G1200,G1160,G966);
  not (G1201,G1160);
  nand (G1202,G609,G1177);
  nand (G1203,G1171,G908);
  not (G1204,G1171);
  nand (G1205,G1158,G1181);
  nand (G1208,G606,G1185);
  nand (G1209,G1187,G1167);
  nand (G1212,G1188,G1170);
  nand (G1215,G914,G1199);
  nand (G1216,G911,G1201);
  nand (G1217,G1176,G1202);
  nand (G1218,G845,G1204);
  nand (G1219,G1192,G1111);
  not (G1220,G1192);
  not (G1221,G1195);
  nand (G1222,G1178,G212);
  not (G1225,G1189);
  nand (G1226,G1189,G1130);
  not (G1227,G1178);
  not (G1230,G1182);
  not (G1233,G1182);
  nand (G1236,G1186,G1208);
  nand (G1239,G1198,G1215);
  nand (G1240,G1200,G1216);
  nand (G1243,G1212,G1156);
  not (G1244,G1212);
  nand (G1245,G1203,G1218);
  nand (G1246,G1072,G1220);
  nand (G1247,G1205,G212);
  not (G1250,G1209);
  nand (G1251,G1209,G1168);
  nand (G1252,G1069,G1225);
  not (G1253,G1217);
  not (G1256,G1205);
  not (G1259,G1239);
  nand (G1260,G1121,G1244);
  not (G1261,G1245);
  nand (G1262,G1219,G1246);
  not (G1263,G1227);
  nand (G1264,G1233,G566);
  not (G1265,G1233);
  nand (G1266,G1230,G567);
  not (G1267,G1230);
  not (G1268,G1236);
  nand (G1269,G1118,G1250);
  not (G1270,G1222);
  not (G1273,G1222);
  nand (G1276,G1226,G1252);
  nand (G1279,G1243,G1260);
  not (G1280,G1253);
  not (G1281,G1256);
  nand (G1282,G458,G1265);
  nand (G1283,G455,G1267);
  not (G1284,G1240);
  not (G1287,G1262);
  not (G1290,G1247);
  not (G1293,G1247);
  not (G1296,G1240);
  nand (G1299,G1251,G1269);
  and (G1302,G1259,G380);
  and (G1305,G381,G1261);
  nand (G1308,G1273,G564);
  not (G1309,G1273);
  nand (G1310,G1270,G565);
  not (G1311,G1270);
  nand (G1312,G1264,G1282);
  nand (G1313,G1266,G1283);
  not (G1316,G1276);
  not (G1317,G1279);
  not (G1320,G1284);
  nand (G1321,G1284,G1280);
  not (G1322,G1287);
  nand (G1323,G1287,G973);
  nand (G1324,G1293,G859);
  not (G1325,G1293);
  nand (G1326,G1290,G860);
  not (G1327,G1290);
  nand (G1328,G452,G1309);
  nand (G1329,G449,G1311);
  not (G1330,G1312);
  not (G1331,G1296);
  nand (G1332,G1296,G1268);
  not (G1333,G1299);
  nand (G1334,G1299,G1065);
  not (G1335,G1302);
  not (G1336,G1305);
  nand (G1337,G1253,G1320);
  not (G1338,G1317);
  nand (G1339,G1317,G1034);
  nand (G1340,G921,G1322);
  nand (G1341,G828,G1325);
  nand (G1342,G825,G1327);
  nand (G1343,G1308,G1328);
  nand (G1344,G1310,G1329);
  not (G1347,G1313);
  not (G1350,G1313);
  nand (G1353,G1236,G1331);
  nand (G1354,G1025,G1333);
  nand (G1355,G1337,G1321);
  nand (G1356,G1000,G1338);
  nand (G1357,G1340,G1323);
  nand (G1358,G1324,G1341);
  nand (G1359,G1326,G1342);
  not (G1362,G1343);
  nand (G1363,G1353,G1332);
  nand (G1366,G1354,G1334);
  not (G1369,G1355);
  nand (G1370,G1356,G1339);
  nand (G1371,G1357,G212);
  not (G1374,G1358);
  not (G1375,G1344);
  not (G1378,G1344);
  not (G1381,G1363);
  not (G1382,G1366);
  nand (G1383,G1369,G212);
  nand (G1386,G1370,G212);
  not (G1389,G1359);
  not (G1392,G1359);
  and (G1395,G1347,G1375);
  and (G1410,G1350,G1375);
  and (G1420,G1347,G1378);
  and (G1434,G1350,G1378);
  not (G1439,G1371);
  not (G1442,G1371);
  not (G1445,G1383);
  not (G1448,G1383);
  not (G1451,G1386);
  not (G1454,G1386);
  nand (G1457,G1442,G562);
  not (G1458,G1442);
  nand (G1459,G1439,G563);
  not (G1460,G1439);
  nand (G1461,G1448,G857);
  not (G1462,G1448);
  nand (G1463,G1445,G858);
  not (G1464,G1445);
  nand (G1465,G1454,G560);
  not (G1466,G1454);
  nand (G1467,G1451,G561);
  not (G1468,G1451);
  nand (G1469,G446,G1458);
  nand (G1470,G443,G1460);
  nand (G1471,G822,G1462);
  nand (G1472,G819,G1464);
  nand (G1473,G440,G1466);
  nand (G1474,G437,G1468);
  nand (G1475,G1457,G1469);
  nand (G1476,G1459,G1470);
  nand (G1479,G1461,G1471);
  nand (G1480,G1463,G1472);
  nand (G1483,G1465,G1473);
  nand (G1484,G1467,G1474);
  not (G1487,G1475);
  not (G1488,G1479);
  not (G1489,G1483);
  not (G1490,G1476);
  not (G1493,G1476);
  not (G1496,G1480);
  and (G1499,G731,G1480);
  not (G1502,G1484);
  and (G1505,G735,G1484);
  nand (G1508,G1374,G1330,G1362,G1487,G546,G1489,G1488,G550);
  not (G1511,G1499);
  not (G1522,G1499);
  not (G1538,G1505);
  not (G1549,G1505);
  and (G1563,G1389,G1490);
  and (G1576,G1392,G1490);
  and (G1584,G1389,G1493);
  and (G1598,G1392,G1493);
  and (G1607,G260,G1508,G235,G235);
  and (G1608,G730,G1496);
  and (G1609,G731,G1496);
  and (G1624,G734,G1502);
  and (G1625,G735,G1502);
  nand (G1642,G1511,G1538,G1584,G1395,G738);
  nand (G1645,G1511,G1538,G1563,G1420,G738);
  nand (G1648,G1511,G1538,G1563,G1410,G738);
  nand (G1651,G1511,G1538,G1576,G1395,G738);
  nand (G1654,G1522,G1538,G1598,G1410,G755);
  nand (G1657,G1522,G1549,G1584,G1434,G755);
  nand (G1660,G1522,G1549,G1598,G1420,G755);
  and (G1663,G1511,G1538,G1584,G1395,G738);
  and (G1666,G1511,G1538,G1563,G1420,G738);
  and (G1669,G1511,G1538,G1563,G1410,G738);
  and (G1672,G1511,G1538,G1576,G1395,G738);
  and (G1675,G1522,G1538,G1598,G1410,G755);
  and (G1678,G1522,G1549,G1584,G1434,G755);
  and (G1681,G1522,G1549,G1598,G1420,G755);
  nand (G1684,G1511,G1625,G1584,G1420,G738);
  nand (G1687,G1522,G1625,G1584,G1410,G738);
  nand (G1690,G1522,G1625,G1598,G1395,G738);
  nand (G1693,G1522,G1625,G1563,G1434,G738);
  nand (G1696,G1522,G1625,G1576,G1420,G755);
  nand (G1699,G1609,G1549,G1584,G1420,G755);
  nand (G1702,G1609,G1549,G1584,G1410,G755);
  nand (G1705,G1609,G1549,G1598,G1395,G755);
  nand (G1708,G1609,G1549,G1576,G1420,G755);
  nand (G1711,G1522,G1625,G1563,G1395,G573);
  nand (G1712,G1609,G1549,G1563,G1395,G573);
  nand (G1713,G1609,G1625,G1584,G1395,G573);
  nand (G1714,G1609,G1625,G1563,G1420,G573);
  nand (G1715,G1609,G1625,G1563,G1410,G573);
  nand (G1716,G1609,G1625,G1576,G1395,G573);
  nand (G1717,G1609,G1624,G1563,G1395,G573);
  nand (G1718,G1608,G1625,G1563,G1395,G573);
  and (G1719,G1511,G1625,G1584,G1420,G738);
  and (G1722,G1522,G1625,G1584,G1410,G738);
  and (G1725,G1522,G1625,G1598,G1395,G738);
  and (G1728,G1522,G1625,G1563,G1434,G738);
  and (G1731,G1522,G1625,G1576,G1420,G755);
  and (G1734,G1609,G1549,G1584,G1420,G755);
  and (G1737,G1609,G1549,G1584,G1410,G755);
  and (G1740,G1609,G1549,G1598,G1395,G755);
  and (G1743,G1609,G1549,G1576,G1420,G755);
  nand (G1746,G1663,G313);
  not (G1747,G1663);
  nand (G1748,G1666,G314);
  not (G1749,G1666);
  nand (G1750,G1669,G315);
  not (G1751,G1669);
  nand (G1752,G1672,G316);
  not (G1753,G1672);
  nand (G1754,G1675,G322);
  not (G1755,G1675);
  nand (G1756,G1678,G327);
  not (G1757,G1678);
  nand (G1758,G1681,G328);
  not (G1759,G1681);
  and (G1760,G1711,G1712,G1713,G1714,G1715,G1716,G1717,G1718);
  nand (G1761,G265,G1747);
  nand (G1762,G268,G1749);
  nand (G1763,G271,G1751);
  nand (G1764,G274,G1753);
  nand (G1765,G1719,G317);
  not (G1766,G1719);
  nand (G1767,G1722,G318);
  not (G1768,G1722);
  nand (G1769,G1725,G319);
  not (G1770,G1725);
  nand (G1771,G1728,G320);
  not (G1772,G1728);
  nand (G1773,G1731,G321);
  not (G1774,G1731);
  nand (G1775,G292,G1755);
  nand (G1776,G1734,G323);
  not (G1777,G1734);
  nand (G1778,G1737,G324);
  not (G1779,G1737);
  nand (G1780,G1740,G325);
  not (G1781,G1740);
  nand (G1782,G1743,G326);
  not (G1783,G1743);
  nand (G1784,G307,G1757);
  nand (G1785,G310,G1759);
  nand (G1786,G1642,G1645,G1648,G1651,G1684,G1687,G1690,G1693);
  nand (G1787,G1696,G1654,G1699,G1702,G1705,G1708,G1657,G1660);
  and (G1788,G1642,G1645,G1648,G1651,G1684,G1687,G1690,G1693);
  and (G1791,G1696,G1654,G1699,G1702,G1705,G1708,G1657,G1660);
  nand (G1794,G277,G1766);
  nand (G1795,G280,G1768);
  nand (G1796,G283,G1770);
  nand (G1797,G286,G1772);
  nand (G1798,G289,G1774);
  nand (G1799,G295,G1777);
  nand (G1800,G298,G1779);
  nand (G1801,G301,G1781);
  nand (G1802,G304,G1783);
  and (G1803,G1786,G197);
  and (G1806,G1787,G198);
  and (G1809,G1788,G1791,G1760);
  nand (G1810,G1788,G1791);
  and (G1817,G260,G1508,G32,G1809);
  nand (G1818,G1803,G1335);
  not (G1819,G1803);
  nand (G1820,G1806,G1336);
  not (G1821,G1806);
  and (G1822,G544,G205,G1810);
  and (G1825,G25,G205,G1810);
  and (G1828,G27,G205,G1810);
  and (G1831,G28,G205,G1810);
  and (G1834,G545,G205,G1810);
  nand (G1837,G1302,G1819);
  nand (G1838,G1305,G1821);
  and (G1839,G26,G205,G1810);
  nand (G1842,G1818,G1837);
  nand (G1845,G1820,G1838);
  nand (G1848,G1822,G1381);
  nand (G1849,G1825,G1382);
  nand (G1850,G1828,G1263);
  nand (G1851,G1831,G1221);
  nand (G1852,G1834,G1281);
  not (G1853,G1822);
  not (G1854,G1825);
  not (G1855,G1828);
  not (G1856,G1831);
  not (G1857,G1834);
  not (G1858,G1839);
  nand (G1859,G1839,G1316);
  nand (G1860,G1363,G1853);
  nand (G1861,G1366,G1854);
  nand (G1862,G1227,G1855);
  nand (G1863,G1195,G1856);
  nand (G1864,G1256,G1857);
  nand (G1865,G1842,G533);
  not (G1866,G1842);
  nand (G1867,G1845,G534);
  not (G1868,G1845);
  nand (G1869,G1276,G1858);
  nand (G1870,G1860,G1848);
  nand (G1871,G1861,G1849);
  nand (G1872,G1862,G1850);
  nand (G1873,G1863,G1851);
  nand (G1874,G1864,G1852);
  nand (G1875,G461,G1866);
  nand (G1876,G464,G1868);
  nand (G1877,G1869,G1859);
  nand (G1880,G1877,G940);
  not (G1881,G1877);
  nand (G1882,G891,G1881);
  nand (G1883,G1880,G1882);
  nand (G1884,G1746,G1761);
  nand (G1885,G1748,G1762);
  nand (G1886,G1750,G1763);
  nand (G1887,G1752,G1764);
  nand (G1888,G1754,G1775);
  nand (G1889,G1756,G1784);
  nand (G1890,G1758,G1785);
  nand (G1891,G1765,G1794);
  nand (G1892,G1767,G1795);
  nand (G1893,G1769,G1796);
  nand (G1894,G1771,G1797);
  nand (G1895,G1773,G1798);
  nand (G1896,G1776,G1799);
  nand (G1897,G1778,G1800);
  nand (G1898,G1780,G1801);
  nand (G1899,G1782,G1802);
  nor (G1900,G1607,G1817);
  and (G1901,G1870,G329);
  and (G1902,G330,G1871);
  and (G1903,G332,G1872);
  and (G1904,G1873,G333);
  and (G1905,G334,G1874);
  nand (G1906,G1865,G1875);
  nand (G1907,G1867,G1876);
  and (G1908,G1883,G331);

endmodule
