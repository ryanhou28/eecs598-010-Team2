// Benchmark "mymod" written by ABC on Wed Nov  1 23:37:58 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58,
    G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70, G71, G72,
    G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86,
    G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G109, G110, G111, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G124,
    G125, G126, G127, G128, G129, G130, G131, G132, G133, G134, G135, G136,
    G137, G138, G139, G140, G141, G142, G143, G144, G145, G146, G147, G148,
    G149, G150, G151, G152, G153, G154, G155, G156, G157, G158, G159, G160,
    G161, G162, G163, G164, G165, G166, G167, G168, G169, G170, G171, G172,
    G173, G174, G175, G176, G177, G178,
    G5193, G5194, G5195, G5196, G5197, G5198, G5199, G5200, G5201, G5202,
    G5203, G5204, G5205, G5206, G5207, G5208, G5209, G5210, G5211, G5212,
    G5213, G5214, G5215, G5216, G5217, G5218, G5219, G5220, G5221, G5222,
    G5223, G5224, G5225, G5226, G5227, G5228, G5229, G5230, G5231, G5232,
    G5233, G5234, G5235, G5236, G5237, G5238, G5239, G5240, G5241, G5242,
    G5243, G5244, G5245, G5246, G5247, G5248, G5249, G5250, G5251, G5252,
    G5253, G5254, G5255, G5256, G5257, G5258, G5259, G5260, G5261, G5262,
    G5263, G5264, G5265, G5266, G5267, G5268, G5269, G5270, G5271, G5272,
    G5273, G5274, G5275, G5276, G5277, G5278, G5279, G5280, G5281, G5282,
    G5283, G5284, G5285, G5286, G5287, G5288, G5289, G5290, G5291, G5292,
    G5293, G5294, G5295, G5296, G5297, G5298, G5299, G5300, G5301, G5302,
    G5303, G5304, G5305, G5306, G5307, G5308, G5309, G5310, G5311, G5312,
    G5313, G5314, G5315  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70,
    G71, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98,
    G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G110,
    G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G133, G134,
    G135, G136, G137, G138, G139, G140, G141, G142, G143, G144, G145, G146,
    G147, G148, G149, G150, G151, G152, G153, G154, G155, G156, G157, G158,
    G159, G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G170,
    G171, G172, G173, G174, G175, G176, G177, G178;
  output G5193, G5194, G5195, G5196, G5197, G5198, G5199, G5200, G5201, G5202,
    G5203, G5204, G5205, G5206, G5207, G5208, G5209, G5210, G5211, G5212,
    G5213, G5214, G5215, G5216, G5217, G5218, G5219, G5220, G5221, G5222,
    G5223, G5224, G5225, G5226, G5227, G5228, G5229, G5230, G5231, G5232,
    G5233, G5234, G5235, G5236, G5237, G5238, G5239, G5240, G5241, G5242,
    G5243, G5244, G5245, G5246, G5247, G5248, G5249, G5250, G5251, G5252,
    G5253, G5254, G5255, G5256, G5257, G5258, G5259, G5260, G5261, G5262,
    G5263, G5264, G5265, G5266, G5267, G5268, G5269, G5270, G5271, G5272,
    G5273, G5274, G5275, G5276, G5277, G5278, G5279, G5280, G5281, G5282,
    G5283, G5284, G5285, G5286, G5287, G5288, G5289, G5290, G5291, G5292,
    G5293, G5294, G5295, G5296, G5297, G5298, G5299, G5300, G5301, G5302,
    G5303, G5304, G5305, G5306, G5307, G5308, G5309, G5310, G5311, G5312,
    G5313, G5314, G5315;
  reg n2610_lo, n2613_lo, n2616_lo, n2619_lo, n2622_lo, n2625_lo, n2628_lo,
    n2634_lo, n2637_lo, n2640_lo, n2643_lo, n2646_lo, n2649_lo, n2652_lo,
    n2655_lo, n2658_lo, n2661_lo, n2664_lo, n2667_lo, n2670_lo, n2673_lo,
    n2676_lo, n2679_lo, n2682_lo, n2685_lo, n2688_lo, n2691_lo, n2694_lo,
    n2697_lo, n2700_lo, n2703_lo, n2706_lo, n2709_lo, n2712_lo, n2715_lo,
    n2718_lo, n2721_lo, n2724_lo, n2727_lo, n2730_lo, n2733_lo, n2736_lo,
    n2739_lo, n2742_lo, n2745_lo, n2748_lo, n2751_lo, n2754_lo, n2757_lo,
    n2760_lo, n2763_lo, n2766_lo, n2769_lo, n2772_lo, n2775_lo, n2778_lo,
    n2781_lo, n2784_lo, n2787_lo, n2790_lo, n2793_lo, n2796_lo, n2799_lo,
    n2802_lo, n2805_lo, n2808_lo, n2811_lo, n2814_lo, n2817_lo, n2820_lo,
    n2823_lo, n2826_lo, n2829_lo, n2832_lo, n2838_lo, n2841_lo, n2844_lo,
    n2847_lo, n2850_lo, n2853_lo, n2856_lo, n2862_lo, n2865_lo, n2868_lo,
    n2871_lo, n2874_lo, n2877_lo, n2880_lo, n2883_lo, n2886_lo, n2889_lo,
    n2892_lo, n2895_lo, n2898_lo, n2901_lo, n2904_lo, n2907_lo, n2910_lo,
    n2913_lo, n2916_lo, n2919_lo, n2922_lo, n2925_lo, n2928_lo, n2931_lo,
    n2934_lo, n2937_lo, n2940_lo, n2943_lo, n2946_lo, n2949_lo, n2952_lo,
    n2955_lo, n2958_lo, n2961_lo, n2964_lo, n2967_lo, n2970_lo, n2973_lo,
    n2976_lo, n2979_lo, n2982_lo, n2985_lo, n2988_lo, n2991_lo, n2994_lo,
    n2997_lo, n3000_lo, n3003_lo, n3006_lo, n3009_lo, n3012_lo, n3015_lo,
    n3018_lo, n3021_lo, n3024_lo, n3027_lo, n3030_lo, n3033_lo, n3036_lo,
    n3039_lo, n3042_lo, n3045_lo, n3048_lo, n3051_lo, n3054_lo, n3057_lo,
    n3060_lo, n3063_lo, n3066_lo, n3069_lo, n3072_lo, n3075_lo, n3078_lo,
    n3081_lo, n3084_lo, n3087_lo, n3090_lo, n3093_lo, n3096_lo, n3099_lo,
    n3102_lo, n3105_lo, n3108_lo, n3111_lo, n3114_lo, n3117_lo, n3120_lo,
    n3126_lo, n3129_lo, n3132_lo, n3138_lo, n3141_lo, n3144_lo, n3147_lo,
    n3150_lo, n3153_lo, n3156_lo, n3162_lo, n3165_lo, n3168_lo, n3174_lo,
    n3177_lo, n3180_lo, n3186_lo, n3189_lo, n3192_lo, n3195_lo, n3198_lo,
    n3201_lo, n3204_lo, n3210_lo, n3213_lo, n3216_lo, n3219_lo, n3222_lo,
    n3225_lo, n3228_lo, n3234_lo, n3237_lo, n3240_lo, n3243_lo, n3246_lo,
    n3249_lo, n3252_lo, n3255_lo, n3258_lo, n3261_lo, n3264_lo, n3267_lo,
    n3270_lo, n3273_lo, n3276_lo, n3279_lo, n3282_lo, n3285_lo, n3288_lo,
    n3294_lo, n3297_lo, n3300_lo, n3306_lo, n3309_lo, n3312_lo, n3318_lo,
    n3321_lo, n3324_lo, n3330_lo, n3333_lo, n3336_lo, n3339_lo, n3342_lo,
    n3345_lo, n3348_lo, n3351_lo, n3354_lo, n3357_lo, n3360_lo, n3363_lo,
    n3366_lo, n3369_lo, n3372_lo, n3375_lo, n3378_lo, n3381_lo, n3384_lo,
    n3387_lo, n3390_lo, n3393_lo, n3396_lo, n3399_lo, n3402_lo, n3405_lo,
    n3408_lo, n3411_lo, n3414_lo, n3417_lo, n3420_lo, n3423_lo, n3426_lo,
    n3429_lo, n3432_lo, n3435_lo, n3438_lo, n3441_lo, n3444_lo, n3447_lo,
    n3450_lo, n3453_lo, n3456_lo, n3459_lo, n3462_lo, n3465_lo, n3468_lo,
    n3471_lo, n3474_lo, n3477_lo, n3480_lo, n3483_lo, n3486_lo, n3489_lo,
    n3492_lo, n3495_lo, n3498_lo, n3501_lo, n3504_lo, n3507_lo, n3510_lo,
    n3513_lo, n3516_lo, n3519_lo, n3522_lo, n3525_lo, n3528_lo, n3531_lo,
    n3534_lo, n3537_lo, n3540_lo, n3543_lo, n3546_lo, n3549_lo, n3552_lo,
    n3555_lo, n3558_lo, n3561_lo, n3564_lo, n3567_lo, n3570_lo, n3573_lo,
    n3576_lo, n3579_lo, n3582_lo, n3585_lo, n3588_lo, n3591_lo, n3594_lo,
    n3597_lo, n3600_lo, n3603_lo, n3606_lo, n3609_lo, n3612_lo, n3615_lo,
    n3618_lo, n3621_lo, n3624_lo, n3627_lo, n3630_lo, n3633_lo, n3636_lo,
    n3639_lo, n3642_lo, n3645_lo, n3648_lo, n3651_lo, n3654_lo, n3666_lo,
    n3750_lo, n3762_lo, n3774_lo, n3786_lo, n3789_lo, n3792_lo, n3795_lo,
    n3798_lo, n3810_lo, n3822_lo, n3834_lo, n3846_lo, n3930_lo, n3933_lo,
    n3936_lo, n3942_lo, n3945_lo, n3948_lo, n3954_lo, n3957_lo, n3963_lo,
    n3966_lo, n3969_lo, n3975_lo, n3978_lo, n3990_lo, n4050_lo, n4062_lo,
    n4098_lo, n4107_lo, n4110_lo, n4122_lo, n4131_lo, n4155_lo, n4158_lo,
    n4170_lo, n4179_lo, n4182_lo, n4185_lo, n4188_lo, n4194_lo, n4197_lo,
    n4200_lo, n4206_lo, n4209_lo, n4212_lo, n4215_lo, n4230_lo, n4233_lo,
    n4236_lo, n4239_lo, n4242_lo, n4254_lo, n4290_lo, n4293_lo, n4302_lo,
    n4314_lo, n4350_lo, n4362_lo, n4374_lo, n4386_lo, n4398_lo, n4410_lo,
    n4413_lo, n4416_lo, n4419_lo, n4422_lo, n4425_lo, n4428_lo, n4431_lo,
    n4434_lo, n4437_lo, n4440_lo, n4443_lo, n4446_lo, n4449_lo, n4452_lo,
    n4455_lo, n4458_lo, n4461_lo, n4464_lo, n4467_lo, n4470_lo, n4473_lo,
    n4476_lo, n4479_lo, n4482_lo, n4485_lo, n4488_lo, n4494_lo, n4497_lo,
    n4500_lo, n4503_lo, n4506_lo, n4509_lo, n4512_lo, n4515_lo, n4518_lo,
    n4521_lo, n4524_lo, n4527_lo, n4530_lo, n4533_lo, n4536_lo, n4539_lo,
    n4542_lo, n4545_lo, n4554_lo, n4557_lo, n4560_lo, n4563_lo, n4566_lo,
    n4569_lo, n4572_lo, n4575_lo, n4578_lo, n4581_lo, n4584_lo, n4587_lo,
    n4590_lo, n4593_lo, n4596_lo, n4602_lo, n4605_lo, n4608_lo, n4614_lo,
    n4617_lo, n4620_lo, n4626_lo, n4629_lo, n4632_lo, n4638_lo, n4641_lo,
    n4644_lo, n4647_lo, n4650_lo, n4653_lo, n4656_lo, n4659_lo, n4662_lo,
    n4665_lo, n4668_lo, n4671_lo, n4674_lo, n4677_lo, n4680_lo, n4683_lo,
    n4686_lo, n4689_lo, n4692_lo, n4695_lo, n4698_lo, n4701_lo, n4704_lo,
    n4707_lo, n4710_lo, n4713_lo, n4716_lo, n4719_lo, n4722_lo, n4725_lo,
    n4728_lo, n4731_lo, n4734_lo, n4737_lo, n4740_lo, n4743_lo, n4970_o2,
    n4972_o2, n4989_o2, n5024_o2, n5025_o2, n5029_o2, n5042_o2, n5048_o2,
    n5093_o2, n5096_o2, n5193_o2, n5199_o2, n5203_o2, n5214_o2, n5221_o2,
    n5222_o2, n5273_o2, n5365_o2, n5385_o2, n5553_o2, n5636_o2, n5782_o2,
    n5778_o2, n5323_o2, n5325_o2, n5327_o2, n5329_o2, n5816_o2, n5817_o2,
    n5837_o2, n5844_o2, n5859_o2, n5857_o2, n5369_o2, n5371_o2, n5373_o2,
    n5400_o2, n5402_o2, n5404_o2, n5406_o2, n5407_o2, n5408_o2, n2722_o2,
    n1942_inv, n5412_o2, n1948_inv, n5557_o2, n5558_o2, n5559_o2, n5564_o2,
    n5565_o2, n1966_inv, n5568_o2, n5598_o2, n5600_o2, n5601_o2, n5602_o2,
    n5603_o2, n2853_o2, n5637_o2, n1993_inv, n1996_inv, n5635_o2, n5640_o2,
    n5641_o2, n5642_o2, n5650_o2, n5652_o2, n5653_o2, n5654_o2, n5655_o2,
    n5657_o2, n2029_inv, n5661_o2, n5656_o2, n5663_o2, n2041_inv, n5795_o2,
    n5796_o2, n5797_o2, n5739_o2, n5773_o2, n2059_inv, n5799_o2, n5802_o2,
    n2068_inv, n5831_o2, n5833_o2, n5820_o2, n5823_o2, n5824_o2, n5869_o2,
    n5848_o2, n5849_o2, n5856_o2, n5896_o2, n2754_o2, n2908_o2, n5892_o2,
    n5915_o2, n5919_o2, n5918_o2, n5920_o2, n5917_o2, lo586_buf_o2,
    n2818_o2, n2863_o2, n2134_inv, n2725_o2, n3016_o2, n3013_o2, n2655_o2,
    n2149_inv, lo562_buf_o2, n2155_inv, n2531_o2, n2700_o2, n5908_o2,
    n5910_o2, n5912_o2, n5914_o2, n2753_o2, n2878_o2, n2182_inv, n5934_o2,
    n5936_o2, n5938_o2, n2728_o2, lo358_buf_o2, lo418_buf_o2, lo474_buf_o2,
    lo554_buf_o2, lo558_buf_o2, lo574_buf_o2, n2215_inv, n2218_inv,
    n2221_inv, lo450_buf_o2, n2910_o2, n2683_o2, n2828_o2, n2582_o2,
    n2600_o2, n2542_o2, n2703_o2, lo510_buf_o2, lo514_buf_o2, lo538_buf_o2,
    lo578_buf_o2, n2260_inv, n2666_o2, n2667_o2, n2660_o2, n2272_inv,
    lo454_buf_o2, n3593_o2, n3048_o2, lo410_buf_o2, lo502_buf_o2,
    lo506_buf_o2, lo550_buf_o2, lo570_buf_o2, lo582_buf_o2, n2302_inv,
    n2305_inv, n3499_o2, n2311_inv, n2870_o2, n2317_inv, n2689_o2,
    n2323_inv, n2662_o2, lo350_buf_o2, lo498_buf_o2, lo518_buf_o2,
    lo522_buf_o2, lo598_buf_o2, n2344_inv, n2347_inv, n2350_inv, n2353_inv,
    n2356_inv, n2359_inv, n2872_o2, n3313_o2, n3273_o2, n2848_o2, n2893_o2,
    n3267_o2, n2925_o2, n2839_o2, n2831_o2, n2558_o2, n2562_o2, n2825_o2,
    n3263_o2, n3517_o2, n2873_o2, n2926_o2, n3261_o2, n3268_o2, n3274_o2,
    n3314_o2, n3571_o2, n2950_o2, n2951_o2, n3022_o2, n3023_o2, n3057_o2,
    n3058_o2, n2931_o2, n2911_o2, n2959_o2, n2960_o2, n2922_o2, n2888_o2,
    n2889_o2, n3051_o2, n3052_o2, n3063_o2, n2845_o2, n2476_inv, n3281_o2,
    n3294_o2, n2885_o2, n2786_o2, n2783_o2, n2801_o2, n2572_o2, n2628_o2,
    n2609_o2, n2618_o2, n2637_o2, n2525_o2, n2551_o2, n3759_o2, n2994_o2,
    n3040_o2, n2943_o2, n2991_o2, n3034_o2, n2881_o2, n3021_o2, n3062_o2,
    n2763_o2, n2764_o2, n2775_o2, n2776_o2, n2968_o2, n2969_o2, n2798_o2,
    n3661_o2, n2694_o2, n2572_inv, n2817_o2, n2514_o2, n2501_o2, n2584_inv,
    n2505_o2, n2492_o2, lo546_buf_o2, lo590_buf_o2, lo594_buf_o2,
    n2602_inv, n2605_inv, n2709_o2, n2611_inv, n2614_inv, n2617_inv,
    n2620_inv, n3590_o2, n3591_o2, n2629_inv, n3638_o2, n3639_o2,
    n2638_inv, n2641_inv, lo458_buf_o2, lo482_buf_o2, lo566_buf_o2,
    n2718_o2, n3707_o2, n3671_o2, n3680_o2, n3749_o2, n3716_o2, n3692_o2,
    n2591_o2, n3478_o2, n3610_o2, n3611_o2, n2686_inv, n2689_inv, n2738_o2,
    n3616_o2, n3617_o2, n3031_o2, n2704_inv, n3562_o2, n2502_o2, n3560_o2,
    n3554_o2, n3555_o2, n3536_o2, n3537_o2, n3508_o2, n3650_o2, n3740_o2,
    n3484_o2, n2740_inv, n2734_o2, n2735_o2, n2711_o2, lo585_buf_o2,
    n2719_o2, n2720_o2, n2723_o2, n2724_o2, n3624_o2, n3625_o2, n3015_o2,
    n3491_o2, n2779_inv, n2811_o2, n3010_o2, n3012_o2, lo382_buf_o2,
    lo386_buf_o2, lo390_buf_o2, lo398_buf_o2, lo402_buf_o2, lo406_buf_o2,
    n3492_o2, lo366_buf_o2, lo374_buf_o2, lo426_buf_o2, lo494_buf_o2,
    n2653_o2, n2654_o2, n2715_o2, n2740_o2, n2682_o2, n2736_o2,
    lo508_buf_o2, lo512_buf_o2, lo536_buf_o2, lo576_buf_o2, lo357_buf_o2,
    lo361_buf_o2, lo417_buf_o2, lo421_buf_o2, lo473_buf_o2, lo477_buf_o2,
    lo553_buf_o2, lo557_buf_o2, lo573_buf_o2, lo434_buf_o2, lo438_buf_o2,
    lo466_buf_o2, lo470_buf_o2, lo490_buf_o2, n2657_o2, n2658_o2, n2663_o2,
    n2664_o2, n2684_o2, n2685_o2;
  wire new_new_n2042__, new_new_n2044__, new_new_n2046__, new_new_n2048__,
    new_new_n2050__, new_new_n2052__, new_new_n2054__, new_new_n2056__,
    new_new_n2058__, new_new_n2060__, new_new_n2062__, new_new_n2064__,
    new_new_n2066__, new_new_n2068__, new_new_n2070__, new_new_n2072__,
    new_new_n2074__, new_new_n2076__, new_new_n2078__, new_new_n2080__,
    new_new_n2082__, new_new_n2084__, new_new_n2086__, new_new_n2088__,
    new_new_n2090__, new_new_n2092__, new_new_n2094__, new_new_n2096__,
    new_new_n2098__, new_new_n2100__, new_new_n2102__, new_new_n2104__,
    new_new_n2106__, new_new_n2108__, new_new_n2110__, new_new_n2112__,
    new_new_n2114__, new_new_n2116__, new_new_n2118__, new_new_n2120__,
    new_new_n2122__, new_new_n2124__, new_new_n2126__, new_new_n2128__,
    new_new_n2130__, new_new_n2132__, new_new_n2134__, new_new_n2136__,
    new_new_n2138__, new_new_n2140__, new_new_n2142__, new_new_n2144__,
    new_new_n2146__, new_new_n2148__, new_new_n2150__, new_new_n2152__,
    new_new_n2154__, new_new_n2156__, new_new_n2158__, new_new_n2160__,
    new_new_n2162__, new_new_n2164__, new_new_n2166__, new_new_n2168__,
    new_new_n2170__, new_new_n2172__, new_new_n2174__, new_new_n2176__,
    new_new_n2178__, new_new_n2180__, new_new_n2182__, new_new_n2184__,
    new_new_n2186__, new_new_n2188__, new_new_n2190__, new_new_n2192__,
    new_new_n2194__, new_new_n2196__, new_new_n2198__, new_new_n2200__,
    new_new_n2202__, new_new_n2204__, new_new_n2206__, new_new_n2208__,
    new_new_n2210__, new_new_n2212__, new_new_n2214__, new_new_n2216__,
    new_new_n2218__, new_new_n2220__, new_new_n2222__, new_new_n2224__,
    new_new_n2226__, new_new_n2228__, new_new_n2230__, new_new_n2232__,
    new_new_n2234__, new_new_n2236__, new_new_n2238__, new_new_n2240__,
    new_new_n2242__, new_new_n2244__, new_new_n2246__, new_new_n2248__,
    new_new_n2250__, new_new_n2252__, new_new_n2254__, new_new_n2256__,
    new_new_n2258__, new_new_n2260__, new_new_n2262__, new_new_n2264__,
    new_new_n2266__, new_new_n2268__, new_new_n2270__, new_new_n2272__,
    new_new_n2274__, new_new_n2276__, new_new_n2278__, new_new_n2280__,
    new_new_n2282__, new_new_n2284__, new_new_n2286__, new_new_n2288__,
    new_new_n2289__, new_new_n2290__, new_new_n2292__, new_new_n2294__,
    new_new_n2296__, new_new_n2298__, new_new_n2300__, new_new_n2302__,
    new_new_n2304__, new_new_n2306__, new_new_n2308__, new_new_n2310__,
    new_new_n2312__, new_new_n2314__, new_new_n2316__, new_new_n2318__,
    new_new_n2320__, new_new_n2322__, new_new_n2324__, new_new_n2326__,
    new_new_n2328__, new_new_n2330__, new_new_n2332__, new_new_n2334__,
    new_new_n2336__, new_new_n2338__, new_new_n2340__, new_new_n2342__,
    new_new_n2344__, new_new_n2346__, new_new_n2348__, new_new_n2350__,
    new_new_n2352__, new_new_n2354__, new_new_n2356__, new_new_n2358__,
    new_new_n2360__, new_new_n2362__, new_new_n2364__, new_new_n2366__,
    new_new_n2368__, new_new_n2370__, new_new_n2372__, new_new_n2374__,
    new_new_n2376__, new_new_n2378__, new_new_n2380__, new_new_n2382__,
    new_new_n2384__, new_new_n2386__, new_new_n2388__, new_new_n2390__,
    new_new_n2392__, new_new_n2394__, new_new_n2396__, new_new_n2398__,
    new_new_n2400__, new_new_n2402__, new_new_n2404__, new_new_n2405__,
    new_new_n2406__, new_new_n2408__, new_new_n2410__, new_new_n2411__,
    new_new_n2412__, new_new_n2414__, new_new_n2416__, new_new_n2418__,
    new_new_n2420__, new_new_n2422__, new_new_n2424__, new_new_n2427__,
    new_new_n2428__, new_new_n2430__, new_new_n2432__, new_new_n2434__,
    new_new_n2436__, new_new_n2438__, new_new_n2440__, new_new_n2442__,
    new_new_n2444__, new_new_n2446__, new_new_n2448__, new_new_n2450__,
    new_new_n2452__, new_new_n2454__, new_new_n2456__, new_new_n2458__,
    new_new_n2460__, new_new_n2462__, new_new_n2464__, new_new_n2466__,
    new_new_n2468__, new_new_n2470__, new_new_n2472__, new_new_n2474__,
    new_new_n2476__, new_new_n2478__, new_new_n2480__, new_new_n2483__,
    new_new_n2484__, new_new_n2486__, new_new_n2488__, new_new_n2491__,
    new_new_n2492__, new_new_n2494__, new_new_n2496__, new_new_n2499__,
    new_new_n2500__, new_new_n2502__, new_new_n2504__, new_new_n2506__,
    new_new_n2508__, new_new_n2510__, new_new_n2512__, new_new_n2514__,
    new_new_n2516__, new_new_n2518__, new_new_n2520__, new_new_n2522__,
    new_new_n2524__, new_new_n2526__, new_new_n2528__, new_new_n2530__,
    new_new_n2532__, new_new_n2534__, new_new_n2536__, new_new_n2538__,
    new_new_n2540__, new_new_n2542__, new_new_n2544__, new_new_n2546__,
    new_new_n2548__, new_new_n2550__, new_new_n2552__, new_new_n2554__,
    new_new_n2556__, new_new_n2558__, new_new_n2559__, new_new_n2560__,
    new_new_n2562__, new_new_n2564__, new_new_n2566__, new_new_n2568__,
    new_new_n2570__, new_new_n2572__, new_new_n2575__, new_new_n2576__,
    new_new_n2578__, new_new_n2580__, new_new_n2583__, new_new_n2584__,
    new_new_n2586__, new_new_n2588__, new_new_n2591__, new_new_n2592__,
    new_new_n2594__, new_new_n2596__, new_new_n2598__, new_new_n2600__,
    new_new_n2602__, new_new_n2604__, new_new_n2606__, new_new_n2608__,
    new_new_n2610__, new_new_n2612__, new_new_n2614__, new_new_n2616__,
    new_new_n2618__, new_new_n2620__, new_new_n2622__, new_new_n2624__,
    new_new_n2626__, new_new_n2628__, new_new_n2630__, new_new_n2632__,
    new_new_n2634__, new_new_n2636__, new_new_n2638__, new_new_n2640__,
    new_new_n2642__, new_new_n2644__, new_new_n2647__, new_new_n2648__,
    new_new_n2650__, new_new_n2652__, new_new_n2655__, new_new_n2656__,
    new_new_n2658__, new_new_n2660__, new_new_n2663__, new_new_n2664__,
    new_new_n2666__, new_new_n2668__, new_new_n2671__, new_new_n2672__,
    new_new_n2674__, new_new_n2676__, new_new_n2678__, new_new_n2680__,
    new_new_n2682__, new_new_n2684__, new_new_n2687__, new_new_n2688__,
    new_new_n2690__, new_new_n2692__, new_new_n2695__, new_new_n2696__,
    new_new_n2698__, new_new_n2700__, new_new_n2702__, new_new_n2704__,
    new_new_n2706__, new_new_n2708__, new_new_n2710__, new_new_n2712__,
    new_new_n2714__, new_new_n2716__, new_new_n2718__, new_new_n2720__,
    new_new_n2722__, new_new_n2724__, new_new_n2726__, new_new_n2728__,
    new_new_n2730__, new_new_n2732__, new_new_n2734__, new_new_n2736__,
    new_new_n2738__, new_new_n2740__, new_new_n2742__, new_new_n2744__,
    new_new_n2746__, new_new_n2748__, new_new_n2750__, new_new_n2752__,
    new_new_n2754__, new_new_n2756__, new_new_n2758__, new_new_n2760__,
    new_new_n2762__, new_new_n2764__, new_new_n2766__, new_new_n2768__,
    new_new_n2770__, new_new_n2772__, new_new_n2774__, new_new_n2776__,
    new_new_n2778__, new_new_n2780__, new_new_n2782__, new_new_n2784__,
    new_new_n2786__, new_new_n2788__, new_new_n2790__, new_new_n2792__,
    new_new_n2794__, new_new_n2796__, new_new_n2798__, new_new_n2800__,
    new_new_n2802__, new_new_n2804__, new_new_n2806__, new_new_n2808__,
    new_new_n2810__, new_new_n2812__, new_new_n2814__, new_new_n2817__,
    new_new_n2818__, new_new_n2820__, new_new_n2822__, new_new_n2824__,
    new_new_n2826__, new_new_n2828__, new_new_n2830__, new_new_n2832__,
    new_new_n2834__, new_new_n2836__, new_new_n2838__, new_new_n2840__,
    new_new_n2843__, new_new_n2844__, new_new_n2846__, new_new_n2848__,
    new_new_n2850__, new_new_n2852__, new_new_n2854__, new_new_n2856__,
    new_new_n2857__, new_new_n2858__, new_new_n2860__, new_new_n2862__,
    new_new_n2865__, new_new_n2866__, new_new_n2868__, new_new_n2870__,
    new_new_n2872__, new_new_n2874__, new_new_n2876__, new_new_n2878__,
    new_new_n2880__, new_new_n2881__, new_new_n2882__, new_new_n2884__,
    new_new_n2886__, new_new_n2889__, new_new_n2890__, new_new_n2892__,
    new_new_n2894__, new_new_n2896__, new_new_n2897__, new_new_n2898__,
    new_new_n2900__, new_new_n2902__, new_new_n2904__, new_new_n2906__,
    new_new_n2908__, new_new_n2910__, new_new_n2912__, new_new_n2914__,
    new_new_n2916__, new_new_n2918__, new_new_n2920__, new_new_n2922__,
    new_new_n2924__, new_new_n2926__, new_new_n2928__, new_new_n2930__,
    new_new_n2932__, new_new_n2934__, new_new_n2936__, new_new_n2938__,
    new_new_n2940__, new_new_n2942__, new_new_n2945__, new_new_n2946__,
    new_new_n2948__, new_new_n2950__, new_new_n2952__, new_new_n2954__,
    new_new_n2956__, new_new_n2958__, new_new_n2960__, new_new_n2962__,
    new_new_n2964__, new_new_n2966__, new_new_n2968__, new_new_n2970__,
    new_new_n2972__, new_new_n2974__, new_new_n2976__, new_new_n2978__,
    new_new_n2980__, new_new_n2982__, new_new_n2984__, new_new_n2986__,
    new_new_n2988__, new_new_n2990__, new_new_n2993__, new_new_n2994__,
    new_new_n2996__, new_new_n2998__, new_new_n3001__, new_new_n3002__,
    new_new_n3004__, new_new_n3006__, new_new_n3008__, new_new_n3010__,
    new_new_n3012__, new_new_n3014__, new_new_n3016__, new_new_n3018__,
    new_new_n3020__, new_new_n3022__, new_new_n3025__, new_new_n3026__,
    new_new_n3028__, new_new_n3030__, new_new_n3032__, new_new_n3034__,
    new_new_n3036__, new_new_n3038__, new_new_n3040__, new_new_n3042__,
    new_new_n3044__, new_new_n3046__, new_new_n3048__, new_new_n3050__,
    new_new_n3052__, new_new_n3054__, new_new_n3056__, new_new_n3058__,
    new_new_n3060__, new_new_n3062__, new_new_n3064__, new_new_n3066__,
    new_new_n3068__, new_new_n3070__, new_new_n3072__, new_new_n3074__,
    new_new_n3076__, new_new_n3078__, new_new_n3080__, new_new_n3083__,
    new_new_n3084__, new_new_n3086__, new_new_n3088__, new_new_n3090__,
    new_new_n3091__, new_new_n3092__, new_new_n3093__, new_new_n3094__,
    new_new_n3096__, new_new_n3098__, new_new_n3099__, new_new_n3100__,
    new_new_n3102__, new_new_n3104__, new_new_n3105__, new_new_n3106__,
    new_new_n3108__, new_new_n3109__, new_new_n3111__, new_new_n3112__,
    new_new_n3114__, new_new_n3116__, new_new_n3117__, new_new_n3118__,
    new_new_n3120__, new_new_n3122__, new_new_n3124__, new_new_n3126__,
    new_new_n3127__, new_new_n3129__, new_new_n3130__, new_new_n3131__,
    new_new_n3132__, new_new_n3133__, new_new_n3135__, new_new_n3137__,
    new_new_n3138__, new_new_n3139__, new_new_n3140__, new_new_n3141__,
    new_new_n3143__, new_new_n3144__, new_new_n3146__, new_new_n3148__,
    new_new_n3149__, new_new_n3150__, new_new_n3152__, new_new_n3154__,
    new_new_n3156__, new_new_n3158__, new_new_n3160__, new_new_n3162__,
    new_new_n3164__, new_new_n3166__, new_new_n3168__, new_new_n3171__,
    new_new_n3172__, new_new_n3173__, new_new_n3174__, new_new_n3175__,
    new_new_n3176__, new_new_n3178__, new_new_n3179__, new_new_n3180__,
    new_new_n3182__, new_new_n3183__, new_new_n3184__, new_new_n3186__,
    new_new_n3188__, new_new_n3189__, new_new_n3190__, new_new_n3191__,
    new_new_n3192__, new_new_n3193__, new_new_n3194__, new_new_n3196__,
    new_new_n3198__, new_new_n3201__, new_new_n3202__, new_new_n3204__,
    new_new_n3206__, new_new_n3208__, new_new_n3209__, new_new_n3210__,
    new_new_n3212__, new_new_n3214__, new_new_n3217__, new_new_n3218__,
    new_new_n3220__, new_new_n3222__, new_new_n3225__, new_new_n3226__,
    new_new_n3228__, new_new_n3230__, new_new_n3233__, new_new_n3234__,
    new_new_n3236__, new_new_n3238__, new_new_n3241__, new_new_n3242__,
    new_new_n3244__, new_new_n3246__, new_new_n3247__, new_new_n3248__,
    new_new_n3250__, new_new_n3252__, new_new_n3254__, new_new_n3255__,
    new_new_n3256__, new_new_n3258__, new_new_n3260__, new_new_n3262__,
    new_new_n3263__, new_new_n3264__, new_new_n3266__, new_new_n3268__,
    new_new_n3270__, new_new_n3271__, new_new_n3272__, new_new_n3274__,
    new_new_n3276__, new_new_n3278__, new_new_n3279__, new_new_n3280__,
    new_new_n3282__, new_new_n3283__, new_new_n3284__, new_new_n3286__,
    new_new_n3288__, new_new_n3290__, new_new_n3291__, new_new_n3292__,
    new_new_n3294__, new_new_n3296__, new_new_n3298__, new_new_n3300__,
    new_new_n3302__, new_new_n3304__, new_new_n3307__, new_new_n3308__,
    new_new_n3310__, new_new_n3312__, new_new_n3314__, new_new_n3316__,
    new_new_n3318__, new_new_n3320__, new_new_n3322__, new_new_n3325__,
    new_new_n3326__, new_new_n3328__, new_new_n3331__, new_new_n3332__,
    new_new_n3334__, new_new_n3336__, new_new_n3338__, new_new_n3339__,
    new_new_n3340__, new_new_n3342__, new_new_n3344__, new_new_n3346__,
    new_new_n3347__, new_new_n3348__, new_new_n3350__, new_new_n3352__,
    new_new_n3354__, new_new_n3355__, new_new_n3356__, new_new_n3358__,
    new_new_n3360__, new_new_n3362__, new_new_n3363__, new_new_n3364__,
    new_new_n3366__, new_new_n3368__, new_new_n3370__, new_new_n3371__,
    new_new_n3372__, new_new_n3374__, new_new_n3376__, new_new_n3378__,
    new_new_n3379__, new_new_n3380__, new_new_n3382__, new_new_n3384__,
    new_new_n3385__, new_new_n3386__, new_new_n3387__, new_new_n3388__,
    new_new_n3390__, new_new_n3392__, new_new_n3393__, new_new_n3394__,
    new_new_n3395__, new_new_n3396__, new_new_n3398__, new_new_n3400__,
    new_new_n3403__, new_new_n3404__, new_new_n3405__, new_new_n3406__,
    new_new_n3407__, new_new_n3408__, new_new_n3409__, new_new_n3410__,
    new_new_n3411__, new_new_n3412__, new_new_n3413__, new_new_n3414__,
    new_new_n3415__, new_new_n3417__, new_new_n3419__, new_new_n3420__,
    new_new_n3421__, new_new_n3422__, new_new_n3423__, new_new_n3425__,
    new_new_n3426__, new_new_n3429__, new_new_n3431__, new_new_n3433__,
    new_new_n3434__, new_new_n3437__, new_new_n3438__, new_new_n3439__,
    new_new_n3440__, new_new_n3442__, new_new_n3443__, new_new_n3445__,
    new_new_n3446__, new_new_n3448__, new_new_n3449__, new_new_n3450__,
    new_new_n3451__, new_new_n3452__, new_new_n3453__, new_new_n3454__,
    new_new_n3455__, new_new_n3456__, new_new_n3457__, new_new_n3459__,
    new_new_n3461__, new_new_n3462__, new_new_n3463__, new_new_n3464__,
    new_new_n3466__, new_new_n3468__, new_new_n3470__, new_new_n3471__,
    new_new_n3472__, new_new_n3473__, new_new_n3474__, new_new_n3475__,
    new_new_n3476__, new_new_n3477__, new_new_n3478__, new_new_n3479__,
    new_new_n3480__, new_new_n3481__, new_new_n3482__, new_new_n3483__,
    new_new_n3484__, new_new_n3485__, new_new_n3486__, new_new_n3487__,
    new_new_n3489__, new_new_n3490__, new_new_n3492__, new_new_n3493__,
    new_new_n3494__, new_new_n3496__, new_new_n3497__, new_new_n3498__,
    new_new_n3500__, new_new_n3501__, new_new_n3502__, new_new_n3505__,
    new_new_n3506__, new_new_n3508__, new_new_n3509__, new_new_n3510__,
    new_new_n3511__, new_new_n3512__, new_new_n3513__, new_new_n3514__,
    new_new_n3516__, new_new_n3517__, new_new_n3518__, new_new_n3519__,
    new_new_n3520__, new_new_n3521__, new_new_n3522__, new_new_n3523__,
    new_new_n3524__, new_new_n3526__, new_new_n3528__, new_new_n3529__,
    new_new_n3530__, new_new_n3531__, new_new_n3532__, new_new_n3533__,
    new_new_n3534__, new_new_n3536__, new_new_n3537__, new_new_n3538__,
    new_new_n3540__, new_new_n3541__, new_new_n3542__, new_new_n3544__,
    new_new_n3545__, new_new_n3546__, new_new_n3548__, new_new_n3551__,
    new_new_n3552__, new_new_n3553__, new_new_n3554__, new_new_n3555__,
    new_new_n3556__, new_new_n3558__, new_new_n3559__, new_new_n3560__,
    new_new_n3561__, new_new_n3562__, new_new_n3563__, new_new_n3564__,
    new_new_n3565__, new_new_n3566__, new_new_n3568__, new_new_n3570__,
    new_new_n3571__, new_new_n3572__, new_new_n3574__, new_new_n3576__,
    new_new_n3577__, new_new_n3578__, new_new_n3579__, new_new_n3580__,
    new_new_n3582__, new_new_n3583__, new_new_n3585__, new_new_n3586__,
    new_new_n3588__, new_new_n3589__, new_new_n3590__, new_new_n3591__,
    new_new_n3592__, new_new_n3594__, new_new_n3595__, new_new_n3596__,
    new_new_n3598__, new_new_n3600__, new_new_n3602__, new_new_n3604__,
    new_new_n3606__, new_new_n3607__, new_new_n3608__, new_new_n3609__,
    new_new_n3610__, new_new_n3612__, new_new_n3613__, new_new_n3614__,
    new_new_n3616__, new_new_n3618__, new_new_n3619__, new_new_n3620__,
    new_new_n3621__, new_new_n3622__, new_new_n3623__, new_new_n3624__,
    new_new_n3625__, new_new_n3626__, new_new_n3627__, new_new_n3628__,
    new_new_n3629__, new_new_n3630__, new_new_n3631__, new_new_n3632__,
    new_new_n3634__, new_new_n3636__, new_new_n3637__, new_new_n3638__,
    new_new_n3639__, new_new_n3640__, new_new_n3641__, new_new_n3642__,
    new_new_n3643__, new_new_n3644__, new_new_n3645__, new_new_n3646__,
    new_new_n3647__, new_new_n3648__, new_new_n3649__, new_new_n3650__,
    new_new_n3652__, new_new_n3653__, new_new_n3654__, new_new_n3655__,
    new_new_n3656__, new_new_n3657__, new_new_n3658__, new_new_n3660__,
    new_new_n3661__, new_new_n3662__, new_new_n3663__, new_new_n3664__,
    new_new_n3665__, new_new_n3666__, new_new_n3667__, new_new_n3668__,
    new_new_n3669__, new_new_n3670__, new_new_n3671__, new_new_n3672__,
    new_new_n3674__, new_new_n3676__, new_new_n3678__, new_new_n3679__,
    new_new_n3680__, new_new_n3682__, new_new_n3683__, new_new_n3685__,
    new_new_n3686__, new_new_n3688__, new_new_n3690__, new_new_n3692__,
    new_new_n3694__, new_new_n3695__, new_new_n3696__, new_new_n3698__,
    new_new_n3699__, new_new_n3700__, new_new_n3701__, new_new_n3702__,
    new_new_n3704__, new_new_n3706__, new_new_n3708__, new_new_n3709__,
    new_new_n3710__, new_new_n3712__, new_new_n3714__, new_new_n3715__,
    new_new_n3716__, new_new_n3717__, new_new_n3718__, new_new_n3719__,
    new_new_n3720__, new_new_n3721__, new_new_n3722__, new_new_n3724__,
    new_new_n3725__, new_new_n3726__, new_new_n3727__, new_new_n3728__,
    new_new_n3729__, new_new_n3730__, new_new_n3732__, new_new_n3734__,
    new_new_n3735__, new_new_n3736__, new_new_n3738__, new_new_n3740__,
    new_new_n3741__, new_new_n3742__, new_new_n3743__, new_new_n3744__,
    new_new_n3745__, new_new_n3746__, new_new_n3747__, new_new_n3748__,
    new_new_n3749__, new_new_n3750__, new_new_n3752__, new_new_n3753__,
    new_new_n3754__, new_new_n3756__, new_new_n3757__, new_new_n3758__,
    new_new_n3760__, new_new_n3762__, new_new_n3764__, new_new_n3765__,
    new_new_n3766__, new_new_n3768__, new_new_n3770__, new_new_n3772__,
    new_new_n3774__, new_new_n3776__, new_new_n3778__, new_new_n3780__,
    new_new_n3782__, new_new_n3785__, new_new_n3786__, new_new_n3788__,
    new_new_n3790__, new_new_n3792__, new_new_n3793__, new_new_n3794__,
    new_new_n3796__, new_new_n3798__, new_new_n3800__, new_new_n3803__,
    new_new_n3804__, new_new_n3806__, new_new_n3808__, new_new_n3811__,
    new_new_n3812__, new_new_n3813__, new_new_n3814__, new_new_n3815__,
    new_new_n3816__, new_new_n3818__, new_new_n3821__, new_new_n3822__,
    new_new_n3825__, new_new_n3826__, new_new_n3827__, new_new_n3828__,
    new_new_n3829__, new_new_n3830__, new_new_n3831__, new_new_n3833__,
    new_new_n3834__, new_new_n3837__, new_new_n3838__, new_new_n3841__,
    new_new_n3843__, new_new_n3844__, new_new_n3846__, new_new_n3848__,
    new_new_n3850__, new_new_n3852__, new_new_n3854__, new_new_n3855__,
    new_new_n3856__, new_new_n3857__, new_new_n3858__, new_new_n3859__,
    new_new_n3860__, new_new_n3861__, new_new_n3862__, new_new_n3863__,
    new_new_n3864__, new_new_n3865__, new_new_n3866__, new_new_n3867__,
    new_new_n3868__, new_new_n3869__, new_new_n3870__, new_new_n3871__,
    new_new_n3872__, new_new_n3874__, new_new_n3876__, new_new_n3877__,
    new_new_n3878__, new_new_n3879__, new_new_n3880__, new_new_n3881__,
    new_new_n3882__, new_new_n3883__, new_new_n3884__, new_new_n3885__,
    new_new_n3887__, new_new_n3889__, new_new_n3890__, new_new_n3892__,
    new_new_n3893__, new_new_n3894__, new_new_n3895__, new_new_n3896__,
    new_new_n3897__, new_new_n3898__, new_new_n3899__, new_new_n3900__,
    new_new_n3901__, new_new_n3902__, new_new_n3903__, new_new_n3904__,
    new_new_n3905__, new_new_n3907__, new_new_n3908__, new_new_n3909__,
    new_new_n3910__, new_new_n3911__, new_new_n3912__, new_new_n3913__,
    new_new_n3915__, new_new_n3917__, new_new_n3918__, new_new_n3920__,
    new_new_n3922__, new_new_n3923__, new_new_n3924__, new_new_n3925__,
    new_new_n3926__, new_new_n3927__, new_new_n3928__, new_new_n3929__,
    new_new_n3930__, new_new_n3932__, new_new_n3934__, new_new_n3935__,
    new_new_n3936__, new_new_n3937__, new_new_n3938__, new_new_n3939__,
    new_new_n3940__, new_new_n3941__, new_new_n3942__, new_new_n3943__,
    new_new_n3944__, new_new_n3945__, new_new_n3946__, new_new_n3947__,
    new_new_n3948__, new_new_n3949__, new_new_n3950__, new_new_n3951__,
    new_new_n3952__, new_new_n3953__, new_new_n3954__, new_new_n3955__,
    new_new_n3956__, new_new_n3957__, new_new_n3958__, new_new_n3959__,
    new_new_n3960__, new_new_n3961__, new_new_n3962__, new_new_n3963__,
    new_new_n3964__, new_new_n3965__, new_new_n3966__, new_new_n3967__,
    new_new_n3968__, new_new_n3969__, new_new_n3970__, new_new_n3971__,
    new_new_n3972__, new_new_n3973__, new_new_n3974__, new_new_n3975__,
    new_new_n3976__, new_new_n3977__, new_new_n3978__, new_new_n3979__,
    new_new_n3980__, new_new_n3981__, new_new_n3982__, new_new_n3983__,
    new_new_n3984__, new_new_n3985__, new_new_n3986__, new_new_n3988__,
    new_new_n3989__, new_new_n3990__, new_new_n3991__, new_new_n3992__,
    new_new_n3993__, new_new_n3994__, new_new_n3995__, new_new_n3996__,
    new_new_n3998__, new_new_n3999__, new_new_n4000__, new_new_n4001__,
    new_new_n4002__, new_new_n4003__, new_new_n4004__, new_new_n4005__,
    new_new_n4006__, new_new_n4007__, new_new_n4008__, new_new_n4009__,
    new_new_n4010__, new_new_n4011__, new_new_n4012__, new_new_n4013__,
    new_new_n4014__, new_new_n4015__, new_new_n4016__, new_new_n4017__,
    new_new_n4018__, new_new_n4019__, new_new_n4020__, new_new_n4021__,
    new_new_n4022__, new_new_n4023__, new_new_n4024__, new_new_n4025__,
    new_new_n4026__, new_new_n4027__, new_new_n4028__, new_new_n4029__,
    new_new_n4030__, new_new_n4031__, new_new_n4032__, new_new_n4033__,
    new_new_n4034__, new_new_n4035__, new_new_n4036__, new_new_n4037__,
    new_new_n4038__, new_new_n4039__, new_new_n4040__, new_new_n4041__,
    new_new_n4042__, new_new_n4043__, new_new_n4044__, new_new_n4045__,
    new_new_n4046__, new_new_n4047__, new_new_n4048__, new_new_n4049__,
    new_new_n4050__, new_new_n4051__, new_new_n4052__, new_new_n4053__,
    new_new_n4054__, new_new_n4055__, new_new_n4056__, new_new_n4057__,
    new_new_n4058__, new_new_n4059__, new_new_n4060__, new_new_n4061__,
    new_new_n4062__, new_new_n4063__, new_new_n4064__, new_new_n4065__,
    new_new_n4066__, new_new_n4067__, new_new_n4068__, new_new_n4069__,
    new_new_n4070__, new_new_n4072__, new_new_n4074__, new_new_n4076__,
    new_new_n4077__, new_new_n4078__, new_new_n4079__, new_new_n4080__,
    new_new_n4081__, new_new_n4082__, new_new_n4083__, new_new_n4084__,
    new_new_n4085__, new_new_n4086__, new_new_n4087__, new_new_n4088__,
    new_new_n4089__, new_new_n4090__, new_new_n4091__, new_new_n4092__,
    new_new_n4093__, new_new_n4094__, new_new_n4095__, new_new_n4096__,
    new_new_n4097__, new_new_n4098__, new_new_n4099__, new_new_n4100__,
    new_new_n4101__, new_new_n4102__, new_new_n4103__, new_new_n4104__,
    new_new_n4105__, new_new_n4106__, new_new_n4108__, new_new_n4110__,
    new_new_n4111__, new_new_n4112__, new_new_n4113__, new_new_n4114__,
    new_new_n4115__, new_new_n4116__, new_new_n4117__, new_new_n4118__,
    new_new_n4119__, new_new_n4120__, new_new_n4121__, new_new_n4122__,
    new_new_n4123__, new_new_n4124__, new_new_n4125__, new_new_n4126__,
    new_new_n4127__, new_new_n4128__, new_new_n4129__, new_new_n4130__,
    new_new_n4131__, new_new_n4132__, new_new_n4133__, new_new_n4134__,
    new_new_n4135__, new_new_n4136__, new_new_n4137__, new_new_n4138__,
    new_new_n4139__, new_new_n4140__, new_new_n4141__, new_new_n4142__,
    new_new_n4143__, new_new_n4144__, new_new_n4145__, new_new_n4146__,
    new_new_n4147__, new_new_n4148__, new_new_n4149__, new_new_n4150__,
    new_new_n4151__, new_new_n4152__, new_new_n4153__, new_new_n4154__,
    new_new_n4155__, new_new_n4156__, new_new_n4157__, new_new_n4158__,
    new_new_n4159__, new_new_n4160__, new_new_n4161__, new_new_n4162__,
    new_new_n4163__, new_new_n4164__, new_new_n4165__, new_new_n4166__,
    new_new_n4167__, new_new_n4168__, new_new_n4169__, new_new_n4170__,
    new_new_n4171__, new_new_n4172__, new_new_n4173__, new_new_n4174__,
    new_new_n4175__, new_new_n4176__, new_new_n4177__, new_new_n4178__,
    new_new_n4179__, new_new_n4180__, new_new_n4181__, new_new_n4182__,
    new_new_n4183__, new_new_n4184__, new_new_n4185__, new_new_n4186__,
    new_new_n4187__, new_new_n4188__, new_new_n4189__, new_new_n4190__,
    new_new_n4191__, new_new_n4192__, new_new_n4193__, new_new_n4194__,
    new_new_n4195__, new_new_n4196__, new_new_n4197__, new_new_n4198__,
    new_new_n4199__, new_new_n4200__, new_new_n4201__, new_new_n4202__,
    new_new_n4203__, new_new_n4204__, new_new_n4205__, new_new_n4206__,
    new_new_n4207__, new_new_n4208__, new_new_n4209__, new_new_n4210__,
    new_new_n4211__, new_new_n4212__, new_new_n4213__, new_new_n4214__,
    new_new_n4215__, new_new_n4216__, new_new_n4217__, new_new_n4218__,
    new_new_n4219__, new_new_n4220__, new_new_n4221__, new_new_n4222__,
    new_new_n4223__, new_new_n4224__, new_new_n4225__, new_new_n4226__,
    new_new_n4227__, new_new_n4228__, new_new_n4229__, new_new_n4230__,
    new_new_n4231__, new_new_n4232__, new_new_n4233__, new_new_n4234__,
    new_new_n4235__, new_new_n4236__, new_new_n4237__, new_new_n4238__,
    new_new_n4239__, new_new_n4240__, new_new_n4241__, new_new_n4242__,
    new_new_n4243__, new_new_n4244__, new_new_n4245__, new_new_n4246__,
    new_new_n4247__, new_new_n4248__, new_new_n4249__, new_new_n4250__,
    new_new_n4251__, new_new_n4252__, new_new_n4253__, new_new_n4254__,
    new_new_n4255__, new_new_n4256__, new_new_n4257__, new_new_n4258__,
    new_new_n4259__, new_new_n4260__, new_new_n4261__, new_new_n4262__,
    new_new_n4263__, new_new_n4264__, new_new_n4265__, new_new_n4266__,
    new_new_n4267__, new_new_n4268__, new_new_n4269__, new_new_n4270__,
    new_new_n4271__, new_new_n4272__, new_new_n4273__, new_new_n4274__,
    new_new_n4275__, new_new_n4276__, new_new_n4277__, new_new_n4278__,
    new_new_n4279__, new_new_n4280__, new_new_n4281__, new_new_n4282__,
    new_new_n4283__, new_new_n4284__, new_new_n4285__, new_new_n4286__,
    new_new_n4287__, new_new_n4288__, new_new_n4289__, new_new_n4290__,
    new_new_n4291__, new_new_n4292__, new_new_n4293__, new_new_n4294__,
    new_new_n4295__, new_new_n4296__, new_new_n4297__, new_new_n4298__,
    new_new_n4299__, new_new_n4300__, new_new_n4301__, new_new_n4302__,
    new_new_n4303__, new_new_n4304__, new_new_n4305__, new_new_n4306__,
    new_new_n4307__, new_new_n4308__, new_new_n4309__, new_new_n4310__,
    new_new_n4311__, new_new_n4312__, new_new_n4313__, new_new_n4314__,
    new_new_n4315__, new_new_n4316__, new_new_n4317__, new_new_n4318__,
    new_new_n4319__, new_new_n4320__, new_new_n4321__, new_new_n4322__,
    new_new_n4323__, new_new_n4324__, new_new_n4325__, new_new_n4326__,
    new_new_n4327__, new_new_n4328__, new_new_n4329__, new_new_n4330__,
    new_new_n4331__, new_new_n4332__, new_new_n4333__, new_new_n4334__,
    new_new_n4335__, new_new_n4336__, new_new_n4337__, new_new_n4338__,
    new_new_n4339__, new_new_n4340__, new_new_n4341__, new_new_n4342__,
    new_new_n4343__, new_new_n4344__, new_new_n4345__, new_new_n4346__,
    new_new_n4347__, new_new_n4348__, new_new_n4349__, new_new_n4350__,
    new_new_n4351__, new_new_n4352__, new_new_n4353__, new_new_n4354__,
    new_new_n4355__, new_new_n4356__, new_new_n4357__, new_new_n4358__,
    new_new_n4359__, new_new_n4360__, new_new_n4361__, new_new_n4362__,
    new_new_n4363__, new_new_n4364__, new_new_n4365__, new_new_n4366__,
    new_new_n4367__, new_new_n4368__, new_new_n4369__, new_new_n4370__,
    new_new_n4371__, new_new_n4372__, new_new_n4373__, new_new_n4374__,
    new_new_n4375__, new_new_n4376__, new_new_n4377__, new_new_n4378__,
    new_new_n4379__, new_new_n4380__, new_new_n4381__, new_new_n4382__,
    new_new_n4383__, new_new_n4384__, new_new_n4385__, new_new_n4386__,
    new_new_n4387__, new_new_n4388__, new_new_n4389__, new_new_n4390__,
    new_new_n4391__, new_new_n4392__, new_new_n4393__, new_new_n4394__,
    new_new_n4395__, new_new_n4396__, new_new_n4397__, new_new_n4398__,
    new_new_n4399__, new_new_n4400__, new_new_n4401__, new_new_n4402__,
    new_new_n4403__, new_new_n4404__, new_new_n4405__, new_new_n4406__,
    new_new_n4407__, new_new_n4408__, new_new_n4409__, new_new_n4410__,
    new_new_n4411__, new_new_n4412__, new_new_n4413__, new_new_n4414__,
    new_new_n4415__, new_new_n4416__, new_new_n4417__, new_new_n4418__,
    new_new_n4419__, new_new_n4420__, new_new_n4421__, new_new_n4422__,
    new_new_n4423__, new_new_n4424__, new_new_n4425__, new_new_n4426__,
    new_new_n4427__, new_new_n4428__, new_new_n4429__, new_new_n4430__,
    new_new_n4431__, new_new_n4432__, new_new_n4433__, new_new_n4434__,
    new_new_n4435__, new_new_n4436__, new_new_n4437__, new_new_n4438__,
    new_new_n4439__, new_new_n4440__, new_new_n4441__, new_new_n4442__,
    new_new_n4443__, new_new_n4444__, new_new_n4445__, new_new_n4446__,
    new_new_n4447__, new_new_n4448__, new_new_n4449__, new_new_n4450__,
    new_new_n4451__, new_new_n4452__, new_new_n4453__, new_new_n4454__,
    new_new_n4455__, new_new_n4456__, new_new_n4457__, new_new_n4458__,
    new_new_n4459__, new_new_n4460__, new_new_n4461__, new_new_n4462__,
    new_new_n4463__, new_new_n4464__, new_new_n4465__, new_new_n4466__,
    new_new_n4467__, new_new_n4468__, new_new_n4469__, new_new_n4470__,
    new_new_n4471__, new_new_n4472__, new_new_n4473__, new_new_n4474__,
    new_new_n4475__, new_new_n4476__, new_new_n4477__, new_new_n4478__,
    new_new_n4479__, new_new_n4480__, new_new_n4481__, new_new_n4482__,
    new_new_n4483__, new_new_n4484__, new_new_n4485__, new_new_n4486__,
    new_new_n4487__, new_new_n4488__, new_new_n4489__, new_new_n4490__,
    new_new_n4491__, new_new_n4492__, new_new_n4493__, new_new_n4494__,
    new_new_n4495__, new_new_n4496__, new_new_n4497__, new_new_n4498__,
    new_new_n4499__, new_new_n4500__, new_new_n4501__, new_new_n4502__,
    new_new_n4503__, new_new_n4504__, new_new_n4505__, new_new_n4506__,
    new_new_n4507__, new_new_n4508__, new_new_n4509__, new_new_n4510__,
    new_new_n4511__, new_new_n4512__, new_new_n4513__, new_new_n4514__,
    new_new_n4515__, new_new_n4516__, new_new_n4517__, new_new_n4518__,
    new_new_n4519__, new_new_n4520__, new_new_n4521__, new_new_n4522__,
    new_new_n4523__, new_new_n4524__, new_new_n4525__, new_new_n4526__,
    new_new_n4527__, new_new_n4528__, new_new_n4529__, new_new_n4530__,
    new_new_n4531__, new_new_n4532__, new_new_n4533__, new_new_n4534__,
    new_new_n4535__, new_new_n4536__, new_new_n4537__, new_new_n4538__,
    new_new_n4539__, new_new_n4540__, new_new_n4541__, new_new_n4542__,
    new_new_n4543__, new_new_n4544__, new_new_n4545__, new_new_n4546__,
    new_new_n4547__, new_new_n4548__, new_new_n4549__, new_new_n4550__,
    new_new_n4551__, new_new_n4552__, new_new_n4553__, new_new_n4554__,
    new_new_n4555__, new_new_n4556__, new_new_n4557__, new_new_n4558__,
    new_new_n4559__, new_new_n4560__, new_new_n4561__, new_new_n4562__,
    new_new_n4563__, new_new_n4564__, new_new_n4565__, new_new_n4566__,
    new_new_n4567__, new_new_n4568__, new_new_n4569__, new_new_n4570__,
    new_new_n4571__, new_new_n4572__, new_new_n4573__, new_new_n4574__,
    new_new_n4575__, new_new_n4576__, new_new_n4577__, new_new_n4578__,
    new_new_n4579__, new_new_n4580__, new_new_n4581__, new_new_n4582__,
    new_new_n4583__, new_new_n4584__, new_new_n4585__, new_new_n4586__,
    new_new_n4587__, new_new_n4588__, new_new_n4589__, new_new_n4590__,
    new_new_n4591__, new_new_n4592__, new_new_n4593__, new_new_n4594__,
    new_new_n4595__, new_new_n4596__, new_new_n4597__, new_new_n4598__,
    new_new_n4599__, new_new_n4600__, new_new_n4601__, new_new_n4602__,
    new_new_n4603__, new_new_n4604__, new_new_n4605__, new_new_n4606__,
    new_new_n4607__, new_new_n4608__, new_new_n4609__, new_new_n4610__,
    new_new_n4611__, new_new_n4612__, new_new_n4613__, new_new_n4614__,
    new_new_n4615__, new_new_n4616__, new_new_n4617__, new_new_n4618__,
    new_new_n4619__, new_new_n4620__, new_new_n4621__, new_new_n4622__,
    new_new_n4623__, new_new_n4624__, new_new_n4625__, new_new_n4626__,
    new_new_n4627__, new_new_n4628__, new_new_n4629__, new_new_n4630__,
    new_new_n4631__, new_new_n4632__, new_new_n4633__, new_new_n4634__,
    new_new_n4635__, new_new_n4636__, new_new_n4637__, new_new_n4638__,
    new_new_n4639__, new_new_n4640__, new_new_n4641__, new_new_n4642__,
    new_new_n4643__, new_new_n4644__, new_new_n4645__, new_new_n4646__,
    new_new_n4647__, new_new_n4648__, new_new_n4649__, new_new_n4650__,
    new_new_n4651__, new_new_n4652__, new_new_n4653__, new_new_n4654__,
    new_new_n4655__, new_new_n4656__, new_new_n4657__, new_new_n4658__,
    new_new_n4659__, new_new_n4660__, new_new_n4661__, new_new_n4662__,
    new_new_n4663__, new_new_n4664__, new_new_n4665__, new_new_n4666__,
    new_new_n4667__, new_new_n4668__, new_new_n4669__, new_new_n4670__,
    new_new_n4671__, new_new_n4672__, new_new_n4673__, new_new_n4674__,
    new_new_n4675__, new_new_n4676__, new_new_n4677__, new_new_n4678__,
    new_new_n4679__, new_new_n4680__, new_new_n4681__, new_new_n4682__,
    new_new_n4683__, new_new_n4684__, new_new_n4685__, new_new_n4686__,
    new_new_n4687__, new_new_n4688__, new_new_n4689__, new_new_n4690__,
    new_new_n4691__, new_new_n4692__, new_new_n4693__, new_new_n4694__,
    new_new_n4695__, new_new_n4696__, new_new_n4697__, new_new_n4698__,
    new_new_n4699__, new_new_n4700__, new_new_n4701__, new_new_n4702__,
    new_new_n4703__, new_new_n4704__, new_new_n4705__, new_new_n4706__,
    new_new_n4707__, new_new_n4708__, new_new_n4709__, new_new_n4710__,
    new_new_n4711__, new_new_n4712__, new_new_n4713__, new_new_n4714__,
    new_new_n4715__, new_new_n4716__, new_new_n4717__, new_new_n4718__,
    new_new_n4719__, new_new_n4720__, new_new_n4721__, new_new_n4722__,
    new_new_n4723__, new_new_n4724__, new_new_n4725__, new_new_n4726__,
    new_new_n4727__, new_new_n4728__, new_new_n4729__, new_new_n4730__,
    new_new_n4731__, new_new_n4732__, new_new_n4733__, new_new_n4734__,
    new_new_n4735__, new_new_n4736__, new_new_n4737__, new_new_n4738__,
    new_new_n4739__, new_new_n4740__, new_new_n4741__, new_new_n4742__,
    new_new_n4743__, new_new_n4744__, new_new_n4745__, new_new_n4746__,
    new_new_n4747__, new_new_n4748__, new_new_n4749__, new_new_n4750__,
    new_new_n4751__, new_new_n4752__, new_new_n4753__, new_new_n4754__,
    new_new_n4755__, new_new_n4756__, new_new_n4757__, new_new_n4758__,
    new_new_n4759__, new_new_n4760__, new_new_n4761__, new_new_n4762__,
    new_new_n4763__, new_new_n4764__, new_new_n4765__, new_new_n4766__,
    new_new_n4767__, new_new_n4768__, new_new_n4769__, new_new_n4770__,
    new_new_n4771__, new_new_n4772__, new_new_n4773__, new_new_n4774__,
    new_new_n4775__, new_new_n4776__, new_new_n4777__, new_new_n4778__,
    new_new_n4779__, new_new_n4780__, new_new_n4781__, new_new_n4782__,
    new_new_n4783__, new_new_n4784__, new_new_n4785__, new_new_n4786__,
    new_new_n4787__, new_new_n4788__, new_new_n4789__, new_new_n4790__,
    new_new_n4791__, new_new_n4792__, new_new_n4793__, new_new_n4794__,
    new_new_n4795__, new_new_n4796__, new_new_n4797__, new_new_n4798__,
    new_new_n4799__, new_new_n4800__, new_new_n4801__, new_new_n4802__,
    new_new_n4803__, new_new_n4804__, new_new_n4805__, new_new_n4806__,
    new_new_n4807__, new_new_n4808__, new_new_n4809__, new_new_n4810__,
    new_new_n4811__, new_new_n4812__, new_new_n4813__, new_new_n4814__,
    new_new_n4815__, new_new_n4816__, new_new_n4817__, new_new_n4818__,
    new_new_n4819__, new_new_n4820__, new_new_n4821__, new_new_n4822__,
    new_new_n4823__, new_new_n4824__, new_new_n4825__, new_new_n4826__,
    new_new_n4827__, new_new_n4828__, new_new_n4829__, new_new_n4830__,
    new_new_n4831__, new_new_n4832__, new_new_n4833__, new_new_n4834__,
    new_new_n4835__, new_new_n4836__, new_new_n4837__, new_new_n4838__,
    new_new_n4839__, new_new_n4840__, new_new_n4841__, new_new_n4842__,
    new_new_n4843__, new_new_n4844__, new_new_n4845__, new_new_n4846__,
    new_new_n4847__, new_new_n4848__, new_new_n4849__, new_new_n4850__,
    new_new_n4851__, new_new_n4852__, new_new_n4853__, new_new_n4854__,
    new_new_n4855__, new_new_n4856__, new_new_n4857__, new_new_n4858__,
    new_new_n4859__, new_new_n4860__, new_new_n4861__, new_new_n4862__,
    new_new_n4863__, new_new_n4864__, new_new_n4865__, new_new_n4866__,
    new_new_n4867__, new_new_n4868__, new_new_n4869__, new_new_n4870__,
    new_new_n4871__, new_new_n4872__, new_new_n4873__, new_new_n4874__,
    new_new_n4875__, new_new_n4876__, new_new_n4877__, new_new_n4878__,
    new_new_n4879__, new_new_n4880__, new_new_n4881__, new_new_n4882__,
    new_new_n4883__, new_new_n4884__, new_new_n4885__, new_new_n4886__,
    new_new_n4887__, new_new_n4888__, new_new_n4889__, new_new_n4890__,
    new_new_n4891__, new_new_n4892__, new_new_n4893__, new_new_n4894__,
    new_new_n4895__, new_new_n4896__, new_new_n4897__, new_new_n4898__,
    new_new_n4899__, new_new_n4900__, new_new_n4901__, new_new_n4902__,
    new_new_n4903__, new_new_n4904__, new_new_n4905__, new_new_n4906__,
    new_new_n4907__, new_new_n4908__, new_new_n4909__, new_new_n4910__,
    new_new_n4911__, new_new_n4912__, new_new_n4913__, new_new_n4914__,
    new_new_n4915__, new_new_n4916__, new_new_n4917__, new_new_n4918__,
    new_new_n4919__, new_new_n4920__, new_new_n4921__, new_new_n4922__,
    new_new_n4923__, new_new_n4924__, new_new_n4925__, new_new_n4926__,
    new_new_n4927__, new_new_n4928__, new_new_n4929__, new_new_n4930__,
    new_new_n4931__, new_new_n4932__, new_new_n4933__, new_new_n4934__,
    new_new_n4935__, new_new_n4936__, new_new_n4937__, new_new_n4938__,
    new_new_n4939__, new_new_n4940__, new_new_n4941__, new_new_n4942__,
    new_new_n4943__, new_new_n4944__, new_new_n4945__, new_new_n4946__,
    new_new_n4947__, new_new_n4948__, new_new_n4949__, new_new_n4950__,
    new_new_n4951__, new_new_n4952__, new_new_n4953__, new_new_n4954__,
    new_new_n4955__, new_new_n4956__, new_new_n4957__, new_new_n4958__,
    new_new_n4959__, new_new_n4960__, new_new_n4961__, new_new_n4962__,
    new_new_n4963__, new_new_n4964__, new_new_n4965__, new_new_n4966__,
    new_new_n4967__, new_new_n4968__, new_new_n4969__, new_new_n4970__,
    new_new_n4971__, new_new_n4972__, new_new_n4973__, new_new_n4974__,
    new_new_n4975__, new_new_n4976__, new_new_n4977__, new_new_n4978__,
    new_new_n4979__, new_new_n4980__, new_new_n4981__, new_new_n4982__,
    new_new_n4983__, new_new_n4984__, new_new_n4985__, new_new_n4986__,
    new_new_n4987__, new_new_n4988__, new_new_n4989__, new_new_n4990__,
    new_new_n4991__, new_new_n4992__, new_new_n4993__, new_new_n4994__,
    new_new_n4995__, new_new_n4996__, new_new_n4997__, new_new_n4998__,
    new_new_n4999__, new_new_n5000__, new_new_n5001__, new_new_n5002__,
    new_new_n5003__, new_new_n5004__, new_new_n5005__, new_new_n5006__,
    new_new_n5007__, new_new_n5008__, new_new_n5009__, new_new_n5010__,
    new_new_n5011__, new_new_n5012__, new_new_n5013__, new_new_n5014__,
    new_new_n5015__, new_new_n5016__, new_new_n5017__, new_new_n5018__,
    new_new_n5019__, new_new_n5020__, new_new_n5021__, new_new_n5022__,
    new_new_n5023__, new_new_n5024__, new_new_n5025__, new_new_n5026__,
    new_new_n5027__, new_new_n5028__, new_new_n5029__, new_new_n5030__,
    new_new_n5031__, new_new_n5032__, new_new_n5033__, new_new_n5034__,
    new_new_n5035__, new_new_n5036__, new_new_n5037__, new_new_n5038__,
    new_new_n5039__, new_new_n5040__, new_new_n5041__, new_new_n5042__,
    new_new_n5043__, new_new_n5044__, new_new_n5045__, new_new_n5046__,
    new_new_n5047__, new_new_n5048__, new_new_n5049__, new_new_n5050__,
    new_new_n5051__, new_new_n5052__, new_new_n5053__, new_new_n5054__,
    new_new_n5055__, new_new_n5056__, new_new_n5057__, new_new_n5058__,
    new_new_n5059__, new_new_n5060__, new_new_n5061__, new_new_n5062__,
    new_new_n5063__, new_new_n5064__, new_new_n5065__, new_new_n5066__,
    new_new_n5067__, new_new_n5068__, new_new_n5069__, new_new_n5070__,
    new_new_n5071__, new_new_n5072__, new_new_n5073__, new_new_n5074__,
    new_new_n5075__, new_new_n5076__, new_new_n5077__, new_new_n5078__,
    new_new_n5079__, new_new_n5080__, new_new_n5081__, new_new_n5082__,
    new_new_n5083__, new_new_n5084__, new_new_n5085__, new_new_n5086__,
    new_new_n5087__, new_new_n5088__, new_new_n5089__, new_new_n5090__,
    new_new_n5091__, new_new_n5092__, new_new_n5093__, new_new_n5094__,
    new_new_n5095__, new_new_n5096__, new_new_n5097__, new_new_n5098__,
    new_new_n5099__, new_new_n5100__, new_new_n5101__, new_new_n5102__,
    new_new_n5103__, new_new_n5104__, new_new_n5105__, new_new_n5106__,
    new_new_n5107__, new_new_n5108__, new_new_n5109__, new_new_n5110__,
    new_new_n5111__, new_new_n5112__, new_new_n5113__, new_new_n5114__,
    new_new_n5115__, new_new_n5116__, new_new_n5117__, new_new_n5118__,
    new_new_n5119__, new_new_n5120__, new_new_n5121__, new_new_n5122__,
    new_new_n5123__, new_new_n5124__, new_new_n5125__, new_new_n5126__,
    new_new_n5127__, new_new_n5128__, new_new_n5129__, new_new_n5130__,
    new_new_n5131__, new_new_n5132__, new_new_n5133__, new_new_n5134__,
    new_new_n5135__, new_new_n5136__, new_new_n5137__, new_new_n5138__,
    new_new_n5139__, new_new_n5140__, new_new_n5141__, new_new_n5142__,
    new_new_n5143__, new_new_n5144__, new_new_n5145__, new_new_n5146__,
    new_new_n5147__, new_new_n5148__, new_new_n5149__, new_new_n5150__,
    new_new_n5151__, new_new_n5152__, new_new_n5153__, new_new_n5154__,
    new_new_n5155__, new_new_n5156__, new_new_n5157__, new_new_n5158__,
    new_new_n5159__, new_new_n5160__, new_new_n5161__, new_new_n5162__,
    new_new_n5163__, new_new_n5164__, new_new_n5165__, new_new_n5166__,
    new_new_n5167__, new_new_n5168__, new_new_n5169__, new_new_n5170__,
    new_new_n5171__, new_new_n5172__, new_new_n5173__, new_new_n5174__,
    new_new_n5175__, new_new_n5176__, new_new_n5177__, new_new_n5178__,
    new_new_n5179__, new_new_n5180__, new_new_n5181__, new_new_n5182__,
    new_new_n5183__, new_new_n5184__, new_new_n5185__, new_new_n5186__,
    new_new_n5187__, new_new_n5188__, new_new_n5189__, new_new_n5190__,
    new_new_n5191__, new_new_n5192__, new_new_n5193__, new_new_n5194__,
    new_new_n5195__, new_new_n5196__, new_new_n5197__, new_new_n5198__,
    new_new_n5199__, new_new_n5200__, new_new_n5201__, new_new_n5202__,
    new_new_n5203__, new_new_n5204__, new_new_n5205__, new_new_n5206__,
    new_new_n5207__, new_new_n5208__, new_new_n5209__, new_new_n5210__,
    new_new_n5211__, new_new_n5212__, new_new_n5213__, new_new_n5214__,
    new_new_n5215__, new_new_n5216__, new_new_n5217__, new_new_n5218__,
    new_new_n5219__, new_new_n5220__, new_new_n5221__, new_new_n5222__,
    new_new_n5223__, new_new_n5224__, new_new_n5225__, new_new_n5226__,
    new_new_n5227__, new_new_n5228__, new_new_n5229__, new_new_n5230__,
    new_new_n5231__, new_new_n5232__, new_new_n5233__, new_new_n5234__,
    new_new_n5235__, new_new_n5236__, new_new_n5237__, new_new_n5238__,
    new_new_n5239__, new_new_n5240__, new_new_n5241__, new_new_n5242__,
    new_new_n5243__, new_new_n5244__, new_new_n5245__, new_new_n5246__,
    new_new_n5247__, new_new_n5248__, new_new_n5249__, new_new_n5250__,
    new_new_n5251__, new_new_n5252__, new_new_n5253__, new_new_n5254__,
    new_new_n5255__, new_new_n5256__, new_new_n5257__, new_new_n5258__,
    new_new_n5259__, new_new_n5260__, new_new_n5261__, new_new_n5262__,
    new_new_n5263__, new_new_n5264__, new_new_n5265__, new_new_n5266__,
    new_new_n5267__, new_new_n5268__, new_new_n5269__, new_new_n5270__,
    new_new_n5271__, new_new_n5272__, new_new_n5273__, new_new_n5274__,
    new_new_n5275__, new_new_n5276__, new_new_n5277__, new_new_n5278__,
    new_new_n5279__, new_new_n5280__, new_new_n5281__, new_new_n5282__,
    new_new_n5283__, new_new_n5284__, new_new_n5285__, new_new_n5286__,
    new_new_n5287__, new_new_n5288__, new_new_n5289__, new_new_n5290__,
    new_new_n5291__, new_new_n5292__, new_new_n5293__, new_new_n5294__,
    new_new_n5295__, new_new_n5296__, new_new_n5297__, new_new_n5298__,
    new_new_n5299__, new_new_n5300__, new_new_n5301__, new_new_n5302__,
    new_new_n5303__, new_new_n5304__, new_new_n5305__, new_new_n5306__,
    new_new_n5307__, new_new_n5308__, new_new_n5309__, new_new_n5310__,
    new_new_n5311__, new_new_n5312__, new_new_n5313__, new_new_n5314__,
    new_new_n5315__, new_new_n5316__, new_new_n5317__, new_new_n5318__,
    new_new_n5319__, new_new_n5320__, new_new_n5321__, new_new_n5322__,
    new_new_n5323__, new_new_n5324__, new_new_n5325__, new_new_n5326__,
    new_new_n5327__, new_new_n5328__, new_new_n5329__, new_new_n5330__,
    new_new_n5331__, new_new_n5332__, new_new_n5333__, new_new_n5334__,
    new_new_n5335__, new_new_n5336__, new_new_n5337__, new_new_n5338__,
    new_new_n5339__, new_new_n5340__, new_new_n5341__, new_new_n5342__,
    new_new_n5343__, new_new_n5344__, new_new_n5345__, new_new_n5346__,
    new_new_n5347__, new_new_n5348__, new_new_n5349__, new_new_n5350__,
    new_new_n5351__, new_new_n5352__, new_new_n5353__, new_new_n5354__,
    new_new_n5355__, new_new_n5356__, new_new_n5357__, new_new_n5358__,
    new_new_n5359__, new_new_n5360__, new_new_n5361__, new_new_n5362__,
    new_new_n5363__, new_new_n5364__, new_new_n5365__, new_new_n5366__,
    new_new_n5367__, new_new_n5368__, new_new_n5369__, new_new_n5370__,
    new_new_n5371__, new_new_n5372__, new_new_n5373__, new_new_n5374__,
    new_new_n5375__, new_new_n5376__, new_new_n5377__, new_new_n5378__,
    new_new_n5379__, new_new_n5380__, new_new_n5381__, new_new_n5382__,
    new_new_n5383__, new_new_n5384__, new_new_n5385__, new_new_n5386__,
    new_new_n5387__, new_new_n5388__, new_new_n5389__, new_new_n5390__,
    new_new_n5391__, new_new_n5392__, new_new_n5393__, new_new_n5394__,
    new_new_n5395__, new_new_n5396__, new_new_n5397__, new_new_n5398__,
    new_new_n5399__, new_new_n5400__, new_new_n5401__, new_new_n5402__,
    new_new_n5403__, new_new_n5404__, new_new_n5405__, new_new_n5406__,
    new_new_n5407__, new_new_n5408__, new_new_n5409__, new_new_n5410__,
    new_new_n5411__, new_new_n5412__, new_new_n5413__, new_new_n5414__,
    new_new_n5415__, new_new_n5416__, new_new_n5417__, new_new_n5418__,
    new_new_n5419__, new_new_n5420__, new_new_n5421__, new_new_n5422__,
    new_new_n5423__, new_new_n5424__, new_new_n5425__, new_new_n5426__,
    new_new_n5427__, new_new_n5428__, new_new_n5429__, new_new_n5430__,
    new_new_n5431__, new_new_n5432__, new_new_n5433__, new_new_n5434__,
    new_new_n5435__, new_new_n5436__, new_new_n5437__, new_new_n5438__,
    new_new_n5439__, new_new_n5440__, new_new_n5441__, new_new_n5442__,
    new_new_n5443__, new_new_n5444__, new_new_n5445__, new_new_n5446__,
    new_new_n5447__, new_new_n5448__, new_new_n5449__, new_new_n5450__,
    new_new_n5451__, new_new_n5452__, new_new_n5453__, new_new_n5454__,
    new_new_n5455__, new_new_n5456__, new_new_n5457__, new_new_n5458__,
    new_new_n5459__, new_new_n5460__, new_new_n5461__, new_new_n5462__,
    new_new_n5463__, new_new_n5464__, new_new_n5465__, new_new_n5466__,
    new_new_n5467__, new_new_n5468__, new_new_n5469__, new_new_n5470__,
    new_new_n5471__, new_new_n5472__, new_new_n5473__, new_new_n5474__,
    new_new_n5475__, new_new_n5476__, new_new_n5477__, new_new_n5478__,
    new_new_n5479__, new_new_n5480__, new_new_n5481__, new_new_n5482__,
    new_new_n5483__, new_new_n5484__, new_new_n5485__, new_new_n5486__,
    new_new_n5487__, new_new_n5488__, new_new_n5489__, new_new_n5490__,
    new_new_n5491__, new_new_n5492__, new_new_n5493__, new_new_n5494__,
    new_new_n5495__, new_new_n5496__, new_new_n5497__, new_new_n5498__,
    new_new_n5499__, new_new_n5500__, new_new_n5501__, new_new_n5502__,
    new_new_n5503__, new_new_n5504__, new_new_n5505__, new_new_n5506__,
    new_new_n5507__, new_new_n5508__, new_new_n5509__, new_new_n5510__,
    new_new_n5511__, new_new_n5512__, new_new_n5513__, new_new_n5514__,
    new_new_n5515__, new_new_n5516__, new_new_n5517__, new_new_n5518__,
    new_new_n5519__, new_new_n5520__, new_new_n5521__, new_new_n5522__,
    new_new_n5523__, new_new_n5524__, new_new_n5525__, new_new_n5526__,
    new_new_n5527__, new_new_n5528__, new_new_n5529__, new_new_n5530__,
    new_new_n5531__, new_new_n5532__, new_new_n5533__, new_new_n5534__,
    new_new_n5535__, new_new_n5536__, new_new_n5537__, new_new_n5538__,
    new_new_n5539__, new_new_n5540__, new_new_n5541__, new_new_n5542__,
    new_new_n5543__, new_new_n5544__, new_new_n5545__, new_new_n5546__,
    new_new_n5547__, new_new_n5548__, new_new_n5549__, new_new_n5550__,
    new_new_n5551__, new_new_n5552__, new_new_n5553__, new_new_n5554__,
    new_new_n5555__, new_new_n5556__, new_new_n5557__, new_new_n5558__,
    new_new_n5559__, new_new_n5560__, new_new_n5561__, new_new_n5562__,
    new_new_n5563__, new_new_n5564__, new_new_n5565__, new_new_n5566__,
    new_new_n5567__, new_new_n5568__, new_new_n5569__, new_new_n5570__,
    new_new_n5571__, new_new_n5572__, new_new_n5573__, new_new_n5574__,
    new_new_n5575__, new_new_n5576__, new_new_n5577__, new_new_n5578__,
    new_new_n5579__, new_new_n5580__, new_new_n5581__, new_new_n5582__,
    new_new_n5583__, new_new_n5584__, new_new_n5585__, new_new_n5586__,
    new_new_n5587__, new_new_n5588__, new_new_n5589__, new_new_n5590__,
    new_new_n5591__, new_new_n5592__, new_new_n5593__, new_new_n5594__,
    new_new_n5595__, new_new_n5596__, new_new_n5597__, new_new_n5598__,
    new_new_n5599__, new_new_n5600__, new_new_n5601__, new_new_n5602__,
    new_new_n5603__, new_new_n5604__, new_new_n5605__, new_new_n5606__,
    new_new_n5607__, new_new_n5608__, new_new_n5609__, new_new_n5610__,
    new_new_n5611__, new_new_n5612__, new_new_n5613__, new_new_n5614__,
    new_new_n5615__, new_new_n5616__, new_new_n5617__, new_new_n5618__,
    new_new_n5619__, new_new_n5620__, new_new_n5621__, new_new_n5622__,
    new_new_n5623__, new_new_n5624__, new_new_n5625__, new_new_n5626__,
    new_new_n5627__, new_new_n5628__, new_new_n5629__, new_new_n5630__,
    new_new_n5631__, new_new_n5632__, new_new_n5633__, new_new_n5634__,
    new_new_n5635__, new_new_n5636__, new_new_n5637__, new_new_n5638__,
    new_new_n5639__, new_new_n5640__, new_new_n5641__, new_new_n5642__,
    new_new_n5643__, new_new_n5644__, new_new_n5645__, new_new_n5646__,
    new_new_n5647__, new_new_n5648__, new_new_n5649__, new_new_n5650__,
    new_new_n5651__, new_new_n5652__, new_new_n5653__, new_new_n5654__,
    new_new_n5655__, new_new_n5656__, new_new_n5657__, new_new_n5658__,
    new_new_n5659__, new_new_n5660__, new_new_n5661__, new_new_n5662__,
    new_new_n5663__, new_new_n5664__, new_new_n5665__, new_new_n5666__,
    new_new_n5667__, new_new_n5668__, new_new_n5669__, new_new_n5670__,
    new_new_n5671__, new_new_n5672__, new_new_n5673__, new_new_n5674__,
    new_new_n5675__, new_new_n5676__, new_new_n5677__, new_new_n5678__,
    new_new_n5679__, new_new_n5680__, new_new_n5681__, new_new_n5682__,
    new_new_n5683__, new_new_n5684__, new_new_n5685__, new_new_n5686__,
    new_new_n5687__, new_new_n5688__, new_new_n5689__, new_new_n5690__,
    new_new_n5691__, new_new_n5692__, new_new_n5693__, new_new_n5694__,
    new_new_n5695__, new_new_n5696__, new_new_n5697__, new_new_n5698__,
    new_new_n5699__, new_new_n5700__, new_new_n5701__, new_new_n5702__,
    new_new_n5703__, new_new_n5704__, new_new_n5705__, new_new_n5706__,
    new_new_n5707__, new_new_n5708__, new_new_n5709__, new_new_n5710__,
    new_new_n5711__, new_new_n5712__, new_new_n5713__, new_new_n5714__,
    new_new_n5715__, new_new_n5716__, new_new_n5717__, new_new_n5718__,
    new_new_n5719__, new_new_n5720__, new_new_n5721__, new_new_n5722__,
    new_new_n5723__, new_new_n5724__, new_new_n5725__, new_new_n5726__,
    new_new_n5727__, new_new_n5728__, new_new_n5729__, new_new_n5730__,
    new_new_n5731__, new_new_n5732__, new_new_n5733__, new_new_n5734__,
    new_new_n5735__, new_new_n5736__, new_new_n5737__, new_new_n5738__,
    new_new_n5739__, new_new_n5740__, new_new_n5741__, new_new_n5742__,
    new_new_n5743__, new_new_n5744__, new_new_n5745__, new_new_n5746__,
    new_new_n5747__, new_new_n6741__, new_new_n6742__, new_new_n6743__,
    new_new_n6744__, new_new_n6745__, new_new_n6746__, new_new_n6747__,
    new_new_n6748__, new_new_n6749__, new_new_n6750__, new_new_n6751__,
    new_new_n6752__, new_new_n6753__, new_new_n6754__, new_new_n6755__,
    new_new_n6756__, new_new_n6757__, new_new_n6758__, new_new_n6759__,
    new_new_n6760__, new_new_n6761__, new_new_n6762__, new_new_n6763__,
    new_new_n6764__, new_new_n6765__, new_new_n6766__, new_new_n6767__,
    new_new_n6768__, new_new_n6769__, new_new_n6770__, new_new_n6771__,
    new_new_n6772__, new_new_n6773__, new_new_n6774__, new_new_n6775__,
    new_new_n6776__, new_new_n6777__, new_new_n6778__, new_new_n6779__,
    new_new_n6780__, new_new_n6781__, new_new_n6782__, new_new_n6783__,
    new_new_n6784__, new_new_n6785__, new_new_n6786__, new_new_n6787__,
    new_new_n6788__, new_new_n6789__, new_new_n6790__, new_new_n6791__,
    new_new_n6792__, new_new_n6793__, new_new_n6794__, new_new_n6795__,
    new_new_n6796__, new_new_n6797__, new_new_n6798__, new_new_n6799__,
    new_new_n6800__, new_new_n6801__, new_new_n6802__, new_new_n6803__,
    new_new_n6804__, new_new_n6805__, new_new_n6806__, new_new_n6807__,
    new_new_n6808__, new_new_n6809__, new_new_n6810__, new_new_n6811__,
    new_new_n6812__, new_new_n6813__, new_new_n6814__, new_new_n6815__,
    new_new_n6816__, new_new_n6817__, new_new_n6818__, new_new_n6819__,
    new_new_n6820__, new_new_n6821__, new_new_n6822__, new_new_n6823__,
    new_new_n6824__, new_new_n6825__, new_new_n6826__, new_new_n6827__,
    new_new_n6828__, new_new_n6829__, new_new_n6830__, new_new_n6831__,
    new_new_n6832__, new_new_n6833__, new_new_n6834__, new_new_n6835__,
    new_new_n6836__, new_new_n6837__, new_new_n6838__, new_new_n6839__,
    new_new_n6840__, new_new_n6841__, new_new_n6842__, new_new_n6843__,
    new_new_n6844__, new_new_n6845__, new_new_n6846__, new_new_n6847__,
    new_new_n6848__, new_new_n6849__, new_new_n6850__, new_new_n6851__,
    new_new_n6852__, new_new_n6853__, new_new_n6854__, new_new_n6855__,
    new_new_n6856__, new_new_n6857__, new_new_n6858__, new_new_n6859__,
    new_new_n6860__, new_new_n6861__, new_new_n6862__, new_new_n6863__,
    new_new_n6864__, new_new_n6865__, new_new_n6866__, new_new_n6867__,
    new_new_n6868__, new_new_n6869__, new_new_n6870__, new_new_n6871__,
    new_new_n6872__, new_new_n6873__, new_new_n6874__, new_new_n6875__,
    new_new_n6876__, new_new_n6877__, new_new_n6878__, new_new_n6879__,
    new_new_n6880__, new_new_n6881__, new_new_n6882__, new_new_n6883__,
    new_new_n6884__, new_new_n6885__, new_new_n6886__, new_new_n6887__,
    new_new_n6888__, new_new_n6889__, new_new_n6890__, new_new_n6891__,
    new_new_n6892__, new_new_n6893__, new_new_n6894__, new_new_n6895__,
    new_new_n6896__, new_new_n6897__, new_new_n6898__, new_new_n6899__,
    new_new_n6900__, new_new_n6901__, new_new_n6902__, new_new_n6903__,
    new_new_n6904__, new_new_n6905__, new_new_n6906__, new_new_n6907__,
    new_new_n6908__, new_new_n6909__, new_new_n6910__, new_new_n6911__,
    new_new_n6912__, new_new_n6913__, new_new_n6914__, new_new_n6915__,
    new_new_n6916__, new_new_n6917__, new_new_n6918__, new_new_n6919__,
    new_new_n6920__, new_new_n6921__, new_new_n6922__, new_new_n6923__,
    new_new_n6924__, new_new_n6925__, new_new_n6926__, new_new_n6927__,
    new_new_n6928__, new_new_n6929__, new_new_n6930__, new_new_n6931__,
    new_new_n6932__, new_new_n6933__, new_new_n6934__, new_new_n6935__,
    new_new_n6936__, new_new_n6937__, new_new_n6938__, new_new_n6939__,
    new_new_n6940__, new_new_n6941__, new_new_n6942__, new_new_n6943__,
    new_new_n6944__, new_new_n6945__, new_new_n6946__, new_new_n6947__,
    new_new_n6948__, new_new_n6949__, new_new_n6950__, new_new_n6951__,
    new_new_n6952__, new_new_n6953__, new_new_n6954__, new_new_n6955__,
    new_new_n6956__, new_new_n6957__, new_new_n6958__, new_new_n6959__,
    new_new_n6960__, new_new_n6961__, new_new_n6962__, new_new_n6963__,
    new_new_n6964__, new_new_n6965__, new_new_n6966__, new_new_n6967__,
    new_new_n6968__, new_new_n6969__, new_new_n6970__, new_new_n6971__,
    new_new_n6972__, new_new_n6973__, new_new_n6974__, new_new_n6975__,
    new_new_n6976__, new_new_n6977__, new_new_n6978__, new_new_n6979__,
    new_new_n6980__, new_new_n6981__, new_new_n6982__, new_new_n6983__,
    new_new_n6984__, new_new_n6985__, new_new_n6986__, new_new_n6987__,
    new_new_n6988__, new_new_n6989__, new_new_n6990__, new_new_n6991__,
    new_new_n6992__, new_new_n6993__, new_new_n6994__, new_new_n6995__,
    new_new_n6996__, new_new_n6997__, new_new_n6998__, new_new_n6999__,
    new_new_n7000__, new_new_n7001__, new_new_n7002__, new_new_n7003__,
    new_new_n7004__, new_new_n7005__, new_new_n7006__, new_new_n7007__,
    new_new_n7008__, new_new_n7009__, new_new_n7010__, new_new_n7011__,
    new_new_n7012__, new_new_n7013__, new_new_n7014__, new_new_n7015__,
    new_new_n7016__, new_new_n7017__, new_new_n7018__, new_new_n7019__,
    new_new_n7020__, new_new_n7021__, new_new_n7022__, new_new_n7023__,
    new_new_n7024__, new_new_n7025__, new_new_n7026__, new_new_n7027__,
    new_new_n7028__, new_new_n7029__, new_new_n7030__, new_new_n7031__,
    new_new_n7032__, new_new_n7033__, new_new_n7034__, new_new_n7035__,
    new_new_n7036__, new_new_n7037__, new_new_n7038__, new_new_n7039__,
    new_new_n7040__, new_new_n7041__, new_new_n7042__, new_new_n7043__,
    new_new_n7044__, new_new_n7045__, new_new_n7046__, new_new_n7047__,
    new_new_n7048__, new_new_n7049__, new_new_n7050__, new_new_n7051__,
    new_new_n7052__, new_new_n7053__, new_new_n7054__, new_new_n7055__,
    new_new_n7056__, new_new_n7057__, new_new_n7058__, new_new_n7059__,
    new_new_n7060__, new_new_n7061__, new_new_n7062__, new_new_n7063__,
    new_new_n7064__, new_new_n7065__, new_new_n7066__, new_new_n7067__,
    new_new_n7068__, new_new_n7069__, new_new_n7070__, new_new_n7071__,
    new_new_n7072__, new_new_n7073__, new_new_n7074__, new_new_n7075__,
    new_new_n7076__, new_new_n7077__, new_new_n7078__, new_new_n7079__,
    new_new_n7080__, new_new_n7081__, new_new_n7082__, new_new_n7083__,
    new_new_n7084__, new_new_n7085__, new_new_n7086__, new_new_n7087__,
    new_new_n7088__, new_new_n7089__, new_new_n7090__, new_new_n7091__,
    new_new_n7092__, new_new_n7093__, new_new_n7094__, new_new_n7095__,
    new_new_n7096__, new_new_n7097__, new_new_n7098__, new_new_n7099__,
    new_new_n7100__, new_new_n7101__, new_new_n7102__, new_new_n7103__,
    new_new_n7104__, new_new_n7105__, new_new_n7106__, new_new_n7107__,
    new_new_n7108__, new_new_n7109__, new_new_n7110__, new_new_n7111__,
    new_new_n7112__, new_new_n7113__, new_new_n7114__, new_new_n7115__,
    new_new_n7116__, new_new_n7117__, new_new_n7118__, new_new_n7119__,
    new_new_n7120__, new_new_n7121__, new_new_n7122__, new_new_n7123__,
    new_new_n7124__, new_new_n7125__, new_new_n7126__, new_new_n7127__,
    new_new_n7128__, new_new_n7129__, new_new_n7130__, new_new_n7131__,
    new_new_n7132__, new_new_n7133__, new_new_n7134__, new_new_n7135__,
    new_new_n7136__, new_new_n7137__, new_new_n7138__, new_new_n7139__,
    new_new_n7140__, new_new_n7141__, new_new_n7142__, new_new_n7143__,
    new_new_n7144__, new_new_n7145__, new_new_n7146__, new_new_n7147__,
    new_new_n7148__, new_new_n7149__, new_new_n7150__, new_new_n7151__,
    new_new_n7152__, new_new_n7153__, new_new_n7154__, new_new_n7155__,
    new_new_n7156__, new_new_n7157__, new_new_n7158__, new_new_n7159__,
    new_new_n7160__, new_new_n7161__, new_new_n7162__, new_new_n7163__,
    new_new_n7164__, new_new_n7165__, new_new_n7166__, new_new_n7167__,
    new_new_n7168__, new_new_n7169__, new_new_n7170__, new_new_n7171__,
    new_new_n7172__, new_new_n7173__, new_new_n7174__, new_new_n7175__,
    new_new_n7176__, new_new_n7177__, new_new_n7178__, new_new_n7179__,
    new_new_n7180__, new_new_n7181__, new_new_n7182__, new_new_n7183__,
    new_new_n7184__, new_new_n7185__, new_new_n7186__, new_new_n7187__,
    new_new_n7188__, new_new_n7189__, new_new_n7190__, new_new_n7191__,
    new_new_n7192__, new_new_n7193__, new_new_n7194__, new_new_n7195__,
    new_new_n7196__, new_new_n7197__, new_new_n7198__, new_new_n7199__,
    new_new_n7200__, new_new_n7201__, new_new_n7202__, new_new_n7203__,
    new_new_n7204__, new_new_n7205__, new_new_n7206__, new_new_n7207__,
    new_new_n7208__, new_new_n7209__, new_new_n7210__, new_new_n7211__,
    new_new_n7212__, new_new_n7213__, new_new_n7214__, new_new_n7215__,
    new_new_n7216__, new_new_n7217__, new_new_n7218__, new_new_n7219__,
    new_new_n7220__, new_new_n7221__, new_new_n7222__, new_new_n7223__,
    new_new_n7224__, new_new_n7225__, new_new_n7226__, new_new_n7227__,
    new_new_n7228__, new_new_n7229__, new_new_n7230__, new_new_n7231__,
    new_new_n7232__, new_new_n7233__, new_new_n7234__, new_new_n7235__,
    new_new_n7236__, new_new_n7237__, new_new_n7238__, new_new_n7239__,
    new_new_n7240__, new_new_n7241__, new_new_n7242__, new_new_n7243__,
    new_new_n7244__, new_new_n7245__, new_new_n7246__, new_new_n7247__,
    new_new_n7248__, new_new_n7249__, new_new_n7250__, new_new_n7251__,
    new_new_n7252__, new_new_n7253__, new_new_n7254__, new_new_n7255__,
    new_new_n7256__, new_new_n7257__, new_new_n7258__, new_new_n7259__,
    new_new_n7260__, new_new_n7261__, new_new_n7262__, new_new_n7263__,
    new_new_n7264__, new_new_n7265__, new_new_n7266__, new_new_n7267__,
    new_new_n7268__, new_new_n7269__, new_new_n7270__, new_new_n7271__,
    new_new_n7272__, new_new_n7273__, new_new_n7274__, new_new_n7275__,
    new_new_n7276__, new_new_n7277__, new_new_n7278__, new_new_n7279__,
    new_new_n7280__, new_new_n7281__, new_new_n7282__, new_new_n7283__,
    new_new_n7284__, new_new_n7285__, new_new_n7286__, new_new_n7287__,
    new_new_n7288__, new_new_n7289__, new_new_n7290__, new_new_n7291__,
    new_new_n7292__, new_new_n7293__, new_new_n7294__, new_new_n7295__,
    new_new_n7296__, new_new_n7297__, new_new_n7298__, new_new_n7299__,
    new_new_n7300__, new_new_n7301__, new_new_n7302__, new_new_n7303__,
    new_new_n7304__, new_new_n7305__, new_new_n7306__, new_new_n7307__,
    new_new_n7308__, new_new_n7309__, new_new_n7310__, new_new_n7311__,
    new_new_n7312__, new_new_n7313__, new_new_n7314__, new_new_n7315__,
    new_new_n7316__, new_new_n7317__, new_new_n7318__, new_new_n7319__,
    new_new_n7320__, new_new_n7321__, new_new_n7322__, new_new_n7323__,
    new_new_n7324__, new_new_n7325__, new_new_n7326__, new_new_n7327__,
    new_new_n7328__, new_new_n7329__, new_new_n7330__, new_new_n7331__,
    new_new_n7332__, new_new_n7333__, new_new_n7334__, new_new_n7335__,
    new_new_n7336__, new_new_n7337__, new_new_n7338__, new_new_n7339__,
    new_new_n7340__, new_new_n7341__, new_new_n7342__, new_new_n7343__,
    new_new_n7344__, new_new_n7345__, new_new_n7346__, new_new_n7347__,
    new_new_n7348__, new_new_n7349__, new_new_n7350__, new_new_n7351__,
    new_new_n7352__, new_new_n7353__, new_new_n7354__, new_new_n7355__,
    new_new_n7356__, new_new_n7357__, new_new_n7358__, new_new_n7359__,
    new_new_n7360__, new_new_n7361__, new_new_n7362__, new_new_n7363__,
    new_new_n7364__, new_new_n7365__, new_new_n7366__, new_new_n7367__,
    new_new_n7368__, new_new_n7369__, new_new_n7370__, new_new_n7371__,
    new_new_n7372__, new_new_n7373__, new_new_n7374__, new_new_n7375__,
    new_new_n7376__, new_new_n7377__, new_new_n7378__, new_new_n7379__,
    new_new_n7380__, new_new_n7381__, new_new_n7382__, new_new_n7383__,
    new_new_n7384__, new_new_n7385__, new_new_n7386__, new_new_n7387__,
    new_new_n7388__, new_new_n7389__, new_new_n7390__, new_new_n7391__,
    new_new_n7392__, new_new_n7393__, new_new_n7394__, new_new_n7395__,
    new_new_n7396__, new_new_n7397__, new_new_n7398__, new_new_n7399__,
    new_new_n7400__, new_new_n7401__, new_new_n7402__, new_new_n7403__,
    new_new_n7404__, new_new_n7405__, new_new_n7406__, new_new_n7407__,
    new_new_n7408__, new_new_n7409__, new_new_n7410__, new_new_n7411__,
    new_new_n7412__, new_new_n7413__, new_new_n7414__, new_new_n7415__,
    new_new_n7416__, new_new_n7417__, new_new_n7418__, new_new_n7419__,
    new_new_n7420__, new_new_n7421__, new_new_n7422__, new_new_n7423__,
    new_new_n7424__, new_new_n7425__, new_new_n7426__, new_new_n7427__,
    new_new_n7428__, new_new_n7429__, new_new_n7430__, new_new_n7431__,
    new_new_n7432__, new_new_n7433__, new_new_n7434__, new_new_n7435__,
    new_new_n7436__, new_new_n7437__, new_new_n7438__, new_new_n7439__,
    new_new_n7440__, new_new_n7441__, new_new_n7442__, new_new_n7443__,
    new_new_n7444__, new_new_n7445__, new_new_n7446__, new_new_n7447__,
    new_new_n7448__, new_new_n7449__, new_new_n7450__, new_new_n7451__,
    new_new_n7452__, new_new_n7453__, new_new_n7454__, new_new_n7455__,
    new_new_n7456__, new_new_n7457__, new_new_n7458__, new_new_n7459__,
    new_new_n7460__, new_new_n7461__, new_new_n7462__, new_new_n7463__,
    new_new_n7464__, new_new_n7465__, new_new_n7466__, new_new_n7467__,
    new_new_n7468__, new_new_n7469__, new_new_n7470__, new_new_n7471__,
    new_new_n7472__, new_new_n7473__, new_new_n7474__, new_new_n7475__,
    new_new_n7476__, new_new_n7477__, new_new_n7478__, new_new_n7479__,
    new_new_n7480__, new_new_n7481__, new_new_n7482__, new_new_n7483__,
    new_new_n7484__, new_new_n7485__, new_new_n7486__, new_new_n7487__,
    new_new_n7488__, new_new_n7489__, new_new_n7490__, new_new_n7491__,
    new_new_n7492__, new_new_n7493__, new_new_n7494__, new_new_n7495__,
    new_new_n7496__, new_new_n7497__, new_new_n7498__, new_new_n7499__,
    new_new_n7500__, new_new_n7501__, new_new_n7502__, new_new_n7503__,
    new_new_n7504__, new_new_n7505__, new_new_n7506__, new_new_n7507__,
    new_new_n7508__, new_new_n7509__, new_new_n7510__, new_new_n7511__,
    new_new_n7512__, new_new_n7513__, new_new_n7514__, new_new_n7515__,
    new_new_n7516__, new_new_n7517__, new_new_n7518__, new_new_n7519__,
    new_new_n7520__, new_new_n7521__, new_new_n7522__, new_new_n7523__,
    new_new_n7524__, new_new_n7525__, new_new_n7526__, new_new_n7527__,
    new_new_n7528__, new_new_n7529__, new_new_n7530__, new_new_n7531__,
    new_new_n7532__, new_new_n7533__, new_new_n7534__, new_new_n7535__,
    new_new_n7536__, new_new_n7537__, new_new_n7538__, new_new_n7539__,
    new_new_n7540__, new_new_n7541__, new_new_n7542__, new_new_n7543__,
    new_new_n7544__, new_new_n7545__, new_new_n7546__, new_new_n7547__,
    new_new_n7548__, new_new_n7549__, new_new_n7550__, new_new_n7551__,
    new_new_n7552__, new_new_n7553__, new_new_n7554__, new_new_n7555__,
    new_new_n7556__, new_new_n7557__, new_new_n7558__, new_new_n7559__,
    new_new_n7560__, new_new_n7561__, new_new_n7562__, new_new_n7563__,
    new_new_n7564__, new_new_n7565__, new_new_n7566__, new_new_n7567__,
    new_new_n7568__, new_new_n7569__, new_new_n7570__, new_new_n7571__,
    new_new_n7572__, new_new_n7573__, new_new_n7574__, new_new_n7575__,
    new_new_n7576__, new_new_n7577__, new_new_n7578__, new_new_n7579__,
    new_new_n7580__, new_new_n7581__, new_new_n7582__, new_new_n7583__,
    new_new_n7584__, new_new_n7585__, new_new_n7586__, new_new_n7587__,
    new_new_n7588__, new_new_n7589__, new_new_n7590__, new_new_n7591__,
    new_new_n7592__, new_new_n7593__, new_new_n7594__, new_new_n7595__,
    new_new_n7596__, new_new_n7597__, new_new_n7598__, new_new_n7599__,
    new_new_n7600__, new_new_n7601__, new_new_n7602__, new_new_n7603__,
    new_new_n7604__, new_new_n7605__, new_new_n7606__, new_new_n7607__,
    new_new_n7608__, new_new_n7609__, new_new_n7610__, new_new_n7611__,
    new_new_n7612__, new_new_n7613__, new_new_n7614__, new_new_n7615__,
    new_new_n7616__, new_new_n7617__, new_new_n7618__, new_new_n7619__,
    new_new_n7620__, new_new_n7621__, new_new_n7622__, new_new_n7623__,
    new_new_n7624__, new_new_n7625__, new_new_n7626__, new_new_n7627__,
    new_new_n7628__, new_new_n7629__, new_new_n7630__, new_new_n7631__,
    new_new_n7632__, new_new_n7633__, new_new_n7634__, new_new_n7635__,
    new_new_n7636__, new_new_n7637__, new_new_n7638__, new_new_n7639__,
    new_new_n7640__, new_new_n7641__, new_new_n7642__, new_new_n7643__,
    new_new_n7644__, new_new_n7645__, new_new_n7646__, new_new_n7647__,
    new_new_n7648__, new_new_n7649__, new_new_n7650__, new_new_n7651__,
    new_new_n7652__, new_new_n7653__, new_new_n7654__, new_new_n7655__,
    new_new_n7656__, new_new_n7657__, new_new_n7658__, new_new_n7659__,
    new_new_n7660__, new_new_n7661__, new_new_n7662__, new_new_n7663__,
    new_new_n7664__, new_new_n7665__, new_new_n7666__, new_new_n7667__,
    new_new_n7668__, new_new_n7669__, new_new_n7670__, new_new_n7671__,
    new_new_n7672__, new_new_n7673__, new_new_n7674__, new_new_n7675__,
    new_new_n7676__, new_new_n7677__, new_new_n7678__, new_new_n7679__,
    new_new_n7680__, new_new_n7681__, new_new_n7682__, new_new_n7683__,
    new_new_n7684__, new_new_n7685__, new_new_n7686__, new_new_n7687__,
    new_new_n7688__, new_new_n7689__, new_new_n7690__, new_new_n7691__,
    new_new_n7692__, new_new_n7693__, new_new_n7694__, new_new_n7695__,
    new_new_n7696__, new_new_n7697__, new_new_n7698__, new_new_n7699__,
    new_new_n7700__, new_new_n7701__, new_new_n7702__, new_new_n7703__,
    new_new_n7704__, new_new_n7705__, new_new_n7706__, new_new_n7707__,
    new_new_n7708__, new_new_n7709__, new_new_n7710__, new_new_n7711__,
    new_new_n7712__, new_new_n7713__, new_new_n7714__, new_new_n7715__,
    new_new_n7716__, new_new_n7717__, new_new_n7718__, new_new_n7719__,
    new_new_n7720__, new_new_n7721__, new_new_n7722__, new_new_n7723__,
    new_new_n7724__, new_new_n7725__, new_new_n7726__, new_new_n7727__,
    new_new_n7728__, new_new_n7729__, new_new_n7730__, new_new_n7731__,
    new_new_n7732__, new_new_n7733__, new_new_n7734__, new_new_n7735__,
    new_new_n7736__, new_new_n7737__, new_new_n7738__, new_new_n7739__,
    new_new_n7740__, new_new_n7741__, new_new_n7742__, new_new_n7743__,
    new_new_n7744__, new_new_n7745__, new_new_n7746__, new_new_n7747__,
    new_new_n7748__, new_new_n7749__, new_new_n7750__, new_new_n7751__,
    new_new_n7752__, new_new_n7753__, new_new_n7754__, new_new_n7755__,
    new_new_n7756__, new_new_n7757__, new_new_n7758__, new_new_n7759__,
    new_new_n7760__, new_new_n7761__, new_new_n7762__, new_new_n7763__,
    new_new_n7764__, new_new_n7765__, new_new_n7766__, new_new_n7767__,
    new_new_n7768__, new_new_n7769__, new_new_n7770__, new_new_n7771__,
    new_new_n7772__, new_new_n7773__, new_new_n7774__, new_new_n7775__,
    new_new_n7776__, new_new_n7777__, new_new_n7778__, new_new_n7779__,
    new_new_n7780__, new_new_n7781__, new_new_n7782__, new_new_n7783__,
    new_new_n7784__, new_new_n7785__, new_new_n7786__, new_new_n7787__,
    new_new_n7788__, new_new_n7789__, new_new_n7790__, new_new_n7791__,
    new_new_n7792__, new_new_n7793__, new_new_n7794__, new_new_n7795__,
    new_new_n7796__, new_new_n7797__, new_new_n7798__, new_new_n7799__,
    new_new_n7800__, new_new_n7801__, new_new_n7802__, new_new_n7803__,
    new_new_n7804__, new_new_n7805__, new_new_n7806__, new_new_n7807__,
    new_new_n7808__, new_new_n7809__, new_new_n7810__, new_new_n7811__,
    new_new_n7812__, new_new_n7813__, new_new_n7814__, new_new_n7815__,
    new_new_n7816__, new_new_n7817__, new_new_n7818__, new_new_n7819__,
    new_new_n7820__, new_new_n7821__, new_new_n7822__, new_new_n7823__,
    new_new_n7824__, new_new_n7825__, new_new_n7826__, new_new_n7827__,
    new_new_n7828__, new_new_n7829__, new_new_n7830__, new_new_n7831__,
    new_new_n7832__, new_new_n7833__, new_new_n7834__, new_new_n7835__,
    new_new_n7836__, new_new_n7837__, new_new_n7838__, new_new_n7839__,
    new_new_n7840__, new_new_n7841__, new_new_n7842__, new_new_n7843__,
    new_new_n7844__, new_new_n7845__, new_new_n7846__, new_new_n7847__,
    new_new_n7848__, new_new_n7849__, new_new_n7850__, new_new_n7851__,
    new_new_n7852__, new_new_n7853__, new_new_n7854__, new_new_n7855__,
    new_new_n7856__, new_new_n7857__, new_new_n7858__, new_new_n7859__,
    new_new_n7860__, new_new_n7861__, new_new_n7862__, new_new_n7863__,
    new_new_n7864__, new_new_n7865__, new_new_n7866__, new_new_n7867__,
    new_new_n7868__, new_new_n7869__, new_new_n7870__, new_new_n7871__,
    new_new_n7872__, new_new_n7873__, new_new_n7874__, new_new_n7875__,
    new_new_n7876__, new_new_n7877__, new_new_n7878__, new_new_n7879__,
    new_new_n7880__, new_new_n7881__, new_new_n7882__, new_new_n7883__,
    new_new_n7884__, new_new_n7885__, new_new_n7886__, new_new_n7887__,
    new_new_n7888__, new_new_n7889__, new_new_n7890__, new_new_n7891__,
    new_new_n7892__, new_new_n7893__, new_new_n7894__, new_new_n7895__,
    new_new_n7896__, new_new_n7897__, new_new_n7898__, new_new_n7899__,
    new_new_n7900__, new_new_n7901__, new_new_n7902__, new_new_n7903__,
    new_new_n7904__, new_new_n7905__, new_new_n7906__, new_new_n7907__,
    new_new_n7908__, new_new_n7909__, new_new_n7910__, new_new_n7911__,
    new_new_n7912__, new_new_n7913__, new_new_n7914__, new_new_n7915__,
    new_new_n7916__, new_new_n7917__, new_new_n7918__, new_new_n7919__,
    new_new_n7920__, new_new_n7921__, new_new_n7922__, new_new_n7923__,
    new_new_n7924__, new_new_n7925__, new_new_n7926__, new_new_n7927__,
    new_new_n7928__, new_new_n7929__, new_new_n7930__, new_new_n7931__,
    new_new_n7932__, new_new_n7933__, new_new_n7934__, new_new_n7935__,
    new_new_n7936__, new_new_n7937__, new_new_n7938__, new_new_n7939__,
    new_new_n7940__, new_new_n7941__, new_new_n7942__, new_new_n7943__,
    new_new_n7944__, new_new_n7945__, new_new_n7946__, new_new_n7947__,
    new_new_n7948__, new_new_n7949__, new_new_n7950__, new_new_n7951__,
    new_new_n7952__, new_new_n7953__, new_new_n7954__, new_new_n7955__,
    new_new_n7956__, new_new_n7957__, new_new_n7958__, new_new_n7959__,
    new_new_n7960__, new_new_n7961__, new_new_n7962__, new_new_n7963__,
    new_new_n7964__, new_new_n7965__, new_new_n7966__, new_new_n7967__,
    new_new_n7968__, new_new_n7969__, new_new_n7970__, new_new_n7971__,
    new_new_n7972__, new_new_n7973__, new_new_n7974__, new_new_n7975__,
    new_new_n7976__, new_new_n7977__, new_new_n7978__, new_new_n7979__,
    new_new_n7980__, new_new_n7981__, new_new_n7982__, new_new_n7983__,
    new_new_n7984__, new_new_n7985__, new_new_n7986__, new_new_n7987__,
    new_new_n7988__, new_new_n7989__, new_new_n7990__, new_new_n7991__,
    new_new_n7992__, new_new_n7993__, new_new_n7994__, new_new_n7995__,
    new_new_n7996__, new_new_n7997__, new_new_n7998__, new_new_n7999__,
    new_new_n8000__, new_new_n8001__, new_new_n8002__, new_new_n8003__,
    new_new_n8004__, new_new_n8005__, new_new_n8006__, new_new_n8007__,
    new_new_n8008__, new_new_n8009__, new_new_n8010__, new_new_n8011__,
    new_new_n8012__, new_new_n8013__, new_new_n8014__, new_new_n8015__,
    new_new_n8016__, new_new_n8017__, new_new_n8018__, new_new_n8019__,
    new_new_n8020__, n11762, n11765, n11768, n11771, n11774, n11777,
    n11780, n11783, n11786, n11789, n11792, n11795, n11798, n11801, n11804,
    n11807, n11810, n11813, n11816, n11819, n11822, n11825, n11828, n11831,
    n11834, n11837, n11840, n11843, n11846, n11849, n11852, n11855, n11858,
    n11861, n11864, n11867, n11870, n11873, n11876, n11879, n11882, n11885,
    n11888, n11891, n11894, n11897, n11900, n11903, n11906, n11909, n11912,
    n11915, n11918, n11921, n11924, n11927, n11930, n11933, n11936, n11939,
    n11942, n11945, n11948, n11951, n11954, n11957, n11960, n11963, n11966,
    n11969, n11972, n11975, n11978, n11981, n11984, n11987, n11990, n11993,
    n11996, n11999, n12002, n12005, n12008, n12011, n12014, n12017, n12020,
    n12023, n12026, n12029, n12032, n12035, n12038, n12041, n12044, n12047,
    n12050, n12053, n12056, n12059, n12062, n12065, n12068, n12071, n12074,
    n12077, n12080, n12083, n12086, n12089, n12092, n12095, n12098, n12101,
    n12104, n12107, n12110, n12113, n12116, n12119, n12122, n12125, n12128,
    n12131, n12134, n12137, n12140, n12143, n12146, n12149, n12152, n12155,
    n12158, n12161, n12164, n12167, n12170, n12173, n12176, n12179, n12182,
    n12185, n12188, n12191, n12194, n12197, n12200, n12203, n12206, n12209,
    n12212, n12215, n12218, n12221, n12224, n12227, n12230, n12233, n12236,
    n12239, n12242, n12245, n12248, n12251, n12254, n12257, n12260, n12263,
    n12266, n12269, n12272, n12275, n12278, n12281, n12284, n12287, n12290,
    n12293, n12296, n12299, n12302, n12305, n12308, n12311, n12314, n12317,
    n12320, n12323, n12326, n12329, n12332, n12335, n12338, n12341, n12344,
    n12347, n12350, n12353, n12356, n12359, n12362, n12365, n12368, n12371,
    n12374, n12377, n12380, n12383, n12386, n12389, n12392, n12395, n12398,
    n12401, n12404, n12407, n12410, n12413, n12416, n12419, n12422, n12425,
    n12428, n12431, n12434, n12437, n12440, n12443, n12446, n12449, n12452,
    n12455, n12458, n12461, n12464, n12467, n12470, n12473, n12476, n12479,
    n12482, n12485, n12488, n12491, n12494, n12497, n12500, n12503, n12506,
    n12509, n12512, n12515, n12518, n12521, n12524, n12527, n12530, n12533,
    n12536, n12539, n12542, n12545, n12548, n12551, n12554, n12557, n12560,
    n12563, n12566, n12569, n12572, n12575, n12578, n12581, n12584, n12587,
    n12590, n12593, n12596, n12599, n12602, n12605, n12608, n12611, n12614,
    n12617, n12620, n12623, n12626, n12629, n12632, n12635, n12638, n12641,
    n12644, n12647, n12650, n12653, n12656, n12659, n12662, n12665, n12668,
    n12671, n12674, n12677, n12680, n12683, n12686, n12689, n12692, n12695,
    n12698, n12701, n12704, n12707, n12710, n12713, n12716, n12719, n12722,
    n12725, n12728, n12731, n12734, n12737, n12740, n12743, n12746, n12749,
    n12752, n12755, n12758, n12761, n12764, n12767, n12770, n12773, n12776,
    n12779, n12782, n12785, n12788, n12791, n12794, n12797, n12800, n12803,
    n12806, n12809, n12812, n12815, n12818, n12821, n12824, n12827, n12830,
    n12833, n12836, n12839, n12842, n12845, n12848, n12851, n12854, n12857,
    n12860, n12863, n12866, n12869, n12872, n12875, n12878, n12881, n12884,
    n12887, n12890, n12893, n12896, n12899, n12902, n12905, n12908, n12911,
    n12914, n12917, n12920, n12923, n12926, n12929, n12932, n12935, n12938,
    n12941, n12944, n12947, n12950, n12953, n12956, n12959, n12962, n12965,
    n12968, n12971, n12974, n12977, n12980, n12983, n12986, n12989, n12992,
    n12995, n12998, n13001, n13004, n13007, n13010, n13013, n13016, n13019,
    n13022, n13025, n13028, n13031, n13034, n13037, n13040, n13043, n13046,
    n13049, n13052, n13055, n13058, n13061, n13064, n13067, n13070, n13073,
    n13076, n13079, n13082, n13085, n13088, n13091, n13094, n13097, n13100,
    n13103, n13106, n13109, n13112, n13115, n13118, n13121, n13124, n13127,
    n13130, n13133, n13136, n13139, n13142, n13145, n13148, n13151, n13154,
    n13157, n13160, n13163, n13166, n13169, n13172, n13175, n13178, n13181,
    n13184, n13187, n13190, n13193, n13196, n13199, n13202, n13205, n13208,
    n13211, n13214, n13217, n13220, n13223, n13226, n13229, n13232, n13235,
    n13238, n13241, n13244, n13247, n13250, n13253, n13256, n13259, n13262,
    n13265, n13268, n13271, n13274, n13277, n13280, n13283, n13286, n13289,
    n13292, n13295, n13298, n13301, n13304, n13307, n13310, n13313, n13316,
    n13319, n13322, n13325, n13328, n13331, n13334, n13337, n13340, n13343,
    n13346, n13349, n13352, n13355, n13358, n13361, n13364, n13367, n13370,
    n13373, n13376, n13379, n13382, n13385, n13388, n13391, n13394, n13397,
    n13400, n13403, n13406, n13409, n13412, n13415, n13418, n13421, n13424,
    n13427, n13430, n13433, n13436, n13439, n13442, n13445, n13448, n13451,
    n13454, n13457, n13460, n13463, n13466, n13469, n13472, n13475, n13478,
    n13481, n13484, n13487, n13490, n13493, n13496, n13499, n13502, n13505,
    n13508, n13511, n13514, n13517, n13520, n13523, n13526, n13529, n13532,
    n13535, n13538, n13541, n13544, n13547, n13550, n13553, n13556, n13559,
    n13562, n13565, n13568, n13571, n13574, n13577, n13580, n13583, n13586,
    n13589, n13592, n13595, n13598, n13601, n13604, n13607, n13610, n13613,
    n13616, n13619, n13622, n13625, n13628, n13631, n13634, n13637, n13640,
    n13643, n13646, n13649, n13652, n13655, n13658, n13661, n13664, n13667,
    n13670, n13673, n13676, n13679, n13682, n13685, n13688, n13691, n13694,
    n13697, n13700, n13703, n13706, n13709, n13712, n13715, n13718, n13721,
    n13724, n13727, n13730, n13733, n13736, n13739, n13742, n13745, n13748,
    n13751, n13754, n13757, n13760, n13763, n13766, n13769, n13772, n13775,
    n13778, n13781, n13784, n13787, n13790, n13793, n13796, n13799, n13802,
    n13805, n13808, n13811, n13814, n13817, n13820, n13823, n13826, n13829,
    n13832, n13835, n13838, n13841, n13844, n13847, n13850, n13853, n13856,
    n13859, n13862, n13865, n13868, n13871, n13874, n13877, n13880, n13883,
    n13886, n13889, n13892, n13895, n13898, n13901, n13904, n13907, n13910,
    n13913, n13916, n13919, n13922, n13925, n13928, n13931, n13934, n13937,
    n13940, n13943, n13946, n13949, n13952, n13955, n13958, n13961, n13964,
    n13967, n13970, n13973, n13976, n13979, n13982, n13985, n13988, n13991,
    n13994, n13997, n14000, n14003, n14006, n14009, n14012, n14015, n14018,
    n14021, n14024, n14027, n14030, n14033, n14036, n14039, n14042, n14045,
    n14048, n14051, n14054, n14057, n14060, n14063, n14066, n14069, n14072,
    n14075, n14078, n14081, n14084, n14087, n14090, n14093, n14096, n14099,
    n14102, n14105, n14108, n14111, n14114, n14117, n14120, n14123, n14126,
    n14129, n14132, n14135, n14138, n14141, n14144, n14147, n14150, n14153,
    n14156, n14159, n14162, n14165, n14168, n14171, n14174, n14177, n14180,
    n14183, n14186, n14189, n14192, n14195, n14198, n14201, n14204, n14207,
    n14210, n14213, n14216, n14219, n14222, n14225, n14228, n14231, n14234,
    n14237, n14240, n14243, n14246, n14249, n14252, n14255, n14258, n14261,
    n14264, n14267, n14270, n14273, n14276, n14279, n14282, n14285, n14288,
    n14291, n14294, n14297, n14300, n14303, n14306, n14309, n14312, n14315,
    n14318, n14321, n14324, n14327, n14330, n14333, n14336, n14339, n14342,
    n14345, n14348, n14351, n14354, n14357, n14360, n14363, n14366, n14369;
  buf1  g0000(.din(G1), .dout(new_new_n2042__));
  buf1  g0001(.din(G2), .dout(new_new_n2044__));
  buf1  g0002(.din(G3), .dout(new_new_n2046__));
  buf1  g0003(.din(G4), .dout(new_new_n2048__));
  buf1  g0004(.din(G5), .dout(new_new_n2050__));
  buf1  g0005(.din(G6), .dout(new_new_n2052__));
  buf1  g0006(.din(G7), .dout(new_new_n2054__));
  buf1  g0007(.din(G8), .dout(new_new_n2056__));
  buf1  g0008(.din(G9), .dout(new_new_n2058__));
  buf1  g0009(.din(G10), .dout(new_new_n2060__));
  buf1  g0010(.din(G11), .dout(new_new_n2062__));
  buf1  g0011(.din(G12), .dout(new_new_n2064__));
  buf1  g0012(.din(G13), .dout(new_new_n2066__));
  buf1  g0013(.din(G14), .dout(new_new_n2068__));
  buf1  g0014(.din(G15), .dout(new_new_n2070__));
  buf1  g0015(.din(G16), .dout(new_new_n2072__));
  buf1  g0016(.din(G17), .dout(new_new_n2074__));
  buf1  g0017(.din(G18), .dout(new_new_n2076__));
  buf1  g0018(.din(G19), .dout(new_new_n2078__));
  buf1  g0019(.din(G20), .dout(new_new_n2080__));
  buf1  g0020(.din(G21), .dout(new_new_n2082__));
  buf1  g0021(.din(G22), .dout(new_new_n2084__));
  buf1  g0022(.din(G23), .dout(new_new_n2086__));
  buf1  g0023(.din(G24), .dout(new_new_n2088__));
  buf1  g0024(.din(G25), .dout(new_new_n2090__));
  buf1  g0025(.din(G26), .dout(new_new_n2092__));
  buf1  g0026(.din(G27), .dout(new_new_n2094__));
  buf1  g0027(.din(G28), .dout(new_new_n2096__));
  buf1  g0028(.din(G29), .dout(new_new_n2098__));
  buf1  g0029(.din(G30), .dout(new_new_n2100__));
  buf1  g0030(.din(G31), .dout(new_new_n2102__));
  buf1  g0031(.din(G32), .dout(new_new_n2104__));
  buf1  g0032(.din(G33), .dout(new_new_n2106__));
  buf1  g0033(.din(G34), .dout(new_new_n2108__));
  buf1  g0034(.din(G35), .dout(new_new_n2110__));
  buf1  g0035(.din(G36), .dout(new_new_n2112__));
  buf1  g0036(.din(G37), .dout(new_new_n2114__));
  buf1  g0037(.din(G38), .dout(new_new_n2116__));
  buf1  g0038(.din(G39), .dout(new_new_n2118__));
  buf1  g0039(.din(G40), .dout(new_new_n2120__));
  buf1  g0040(.din(G41), .dout(new_new_n2122__));
  buf1  g0041(.din(G42), .dout(new_new_n2124__));
  buf1  g0042(.din(G43), .dout(new_new_n2126__));
  buf1  g0043(.din(G44), .dout(new_new_n2128__));
  buf1  g0044(.din(G45), .dout(new_new_n2130__));
  buf1  g0045(.din(G46), .dout(new_new_n2132__));
  buf1  g0046(.din(G47), .dout(new_new_n2134__));
  buf1  g0047(.din(G48), .dout(new_new_n2136__));
  buf1  g0048(.din(G49), .dout(new_new_n2138__));
  buf1  g0049(.din(G50), .dout(new_new_n2140__));
  buf1  g0050(.din(G51), .dout(new_new_n2142__));
  buf1  g0051(.din(G52), .dout(new_new_n2144__));
  buf1  g0052(.din(G53), .dout(new_new_n2146__));
  buf1  g0053(.din(G54), .dout(new_new_n2148__));
  buf1  g0054(.din(G55), .dout(new_new_n2150__));
  buf1  g0055(.din(G56), .dout(new_new_n2152__));
  buf1  g0056(.din(G57), .dout(new_new_n2154__));
  buf1  g0057(.din(G58), .dout(new_new_n2156__));
  buf1  g0058(.din(G59), .dout(new_new_n2158__));
  buf1  g0059(.din(G60), .dout(new_new_n2160__));
  buf1  g0060(.din(G61), .dout(new_new_n2162__));
  buf1  g0061(.din(G62), .dout(new_new_n2164__));
  buf1  g0062(.din(G63), .dout(new_new_n2166__));
  buf1  g0063(.din(G64), .dout(new_new_n2168__));
  buf1  g0064(.din(G65), .dout(new_new_n2170__));
  buf1  g0065(.din(G66), .dout(new_new_n2172__));
  buf1  g0066(.din(G67), .dout(new_new_n2174__));
  buf1  g0067(.din(G68), .dout(new_new_n2176__));
  buf1  g0068(.din(G69), .dout(new_new_n2178__));
  buf1  g0069(.din(G70), .dout(new_new_n2180__));
  buf1  g0070(.din(G71), .dout(new_new_n2182__));
  buf1  g0071(.din(G72), .dout(new_new_n2184__));
  buf1  g0072(.din(G73), .dout(new_new_n2186__));
  buf1  g0073(.din(G74), .dout(new_new_n2188__));
  buf1  g0074(.din(G75), .dout(new_new_n2190__));
  buf1  g0075(.din(G76), .dout(new_new_n2192__));
  buf1  g0076(.din(G77), .dout(new_new_n2194__));
  buf1  g0077(.din(G78), .dout(new_new_n2196__));
  buf1  g0078(.din(G79), .dout(new_new_n2198__));
  buf1  g0079(.din(G80), .dout(new_new_n2200__));
  buf1  g0080(.din(G81), .dout(new_new_n2202__));
  buf1  g0081(.din(G82), .dout(new_new_n2204__));
  buf1  g0082(.din(G83), .dout(new_new_n2206__));
  buf1  g0083(.din(G84), .dout(new_new_n2208__));
  buf1  g0084(.din(G85), .dout(new_new_n2210__));
  buf1  g0085(.din(G86), .dout(new_new_n2212__));
  buf1  g0086(.din(G87), .dout(new_new_n2214__));
  buf1  g0087(.din(G88), .dout(new_new_n2216__));
  buf1  g0088(.din(G89), .dout(new_new_n2218__));
  buf1  g0089(.din(G90), .dout(new_new_n2220__));
  buf1  g0090(.din(G91), .dout(new_new_n2222__));
  buf1  g0091(.din(G92), .dout(new_new_n2224__));
  buf1  g0092(.din(G93), .dout(new_new_n2226__));
  buf1  g0093(.din(G94), .dout(new_new_n2228__));
  buf1  g0094(.din(G95), .dout(new_new_n2230__));
  buf1  g0095(.din(G96), .dout(new_new_n2232__));
  buf1  g0096(.din(G97), .dout(new_new_n2234__));
  buf1  g0097(.din(G98), .dout(new_new_n2236__));
  buf1  g0098(.din(G99), .dout(new_new_n2238__));
  buf1  g0099(.din(G100), .dout(new_new_n2240__));
  buf1  g0100(.din(G101), .dout(new_new_n2242__));
  buf1  g0101(.din(G102), .dout(new_new_n2244__));
  buf1  g0102(.din(G103), .dout(new_new_n2246__));
  buf1  g0103(.din(G104), .dout(new_new_n2248__));
  buf1  g0104(.din(G105), .dout(new_new_n2250__));
  buf1  g0105(.din(G106), .dout(new_new_n2252__));
  buf1  g0106(.din(G107), .dout(new_new_n2254__));
  buf1  g0107(.din(G108), .dout(new_new_n2256__));
  buf1  g0108(.din(G109), .dout(new_new_n2258__));
  buf1  g0109(.din(G110), .dout(new_new_n2260__));
  buf1  g0110(.din(G111), .dout(new_new_n2262__));
  buf1  g0111(.din(G112), .dout(new_new_n2264__));
  buf1  g0112(.din(G113), .dout(new_new_n2266__));
  buf1  g0113(.din(G114), .dout(new_new_n2268__));
  buf1  g0114(.din(G115), .dout(new_new_n2270__));
  buf1  g0115(.din(G116), .dout(new_new_n2272__));
  buf1  g0116(.din(G117), .dout(new_new_n2274__));
  buf1  g0117(.din(G118), .dout(new_new_n2276__));
  buf1  g0118(.din(G119), .dout(new_new_n2278__));
  buf1  g0119(.din(G120), .dout(new_new_n2280__));
  buf1  g0120(.din(G121), .dout(new_new_n2282__));
  buf1  g0121(.din(G122), .dout(new_new_n2284__));
  buf1  g0122(.din(G123), .dout(new_new_n2286__));
  buf1  g0123(.din(G124), .dout(new_new_n2288__));
  not1  g0124(.din(G124), .dout(new_new_n2289__));
  buf1  g0125(.din(G125), .dout(new_new_n2290__));
  buf1  g0126(.din(G126), .dout(new_new_n2292__));
  buf1  g0127(.din(G127), .dout(new_new_n2294__));
  buf1  g0128(.din(G128), .dout(new_new_n2296__));
  buf1  g0129(.din(G129), .dout(new_new_n2298__));
  buf1  g0130(.din(G130), .dout(new_new_n2300__));
  buf1  g0131(.din(G131), .dout(new_new_n2302__));
  buf1  g0132(.din(G132), .dout(new_new_n2304__));
  buf1  g0133(.din(G133), .dout(new_new_n2306__));
  buf1  g0134(.din(G134), .dout(new_new_n2308__));
  buf1  g0135(.din(G135), .dout(new_new_n2310__));
  buf1  g0136(.din(G136), .dout(new_new_n2312__));
  buf1  g0137(.din(G137), .dout(new_new_n2314__));
  buf1  g0138(.din(G138), .dout(new_new_n2316__));
  buf1  g0139(.din(G139), .dout(new_new_n2318__));
  buf1  g0140(.din(G140), .dout(new_new_n2320__));
  buf1  g0141(.din(G141), .dout(new_new_n2322__));
  buf1  g0142(.din(G142), .dout(new_new_n2324__));
  buf1  g0143(.din(G143), .dout(new_new_n2326__));
  buf1  g0144(.din(G144), .dout(new_new_n2328__));
  buf1  g0145(.din(G145), .dout(new_new_n2330__));
  buf1  g0146(.din(G146), .dout(new_new_n2332__));
  buf1  g0147(.din(G147), .dout(new_new_n2334__));
  buf1  g0148(.din(G148), .dout(new_new_n2336__));
  buf1  g0149(.din(G149), .dout(new_new_n2338__));
  buf1  g0150(.din(G150), .dout(new_new_n2340__));
  buf1  g0151(.din(G151), .dout(new_new_n2342__));
  buf1  g0152(.din(G152), .dout(new_new_n2344__));
  buf1  g0153(.din(G153), .dout(new_new_n2346__));
  buf1  g0154(.din(G154), .dout(new_new_n2348__));
  buf1  g0155(.din(G155), .dout(new_new_n2350__));
  buf1  g0156(.din(G156), .dout(new_new_n2352__));
  buf1  g0157(.din(G157), .dout(new_new_n2354__));
  buf1  g0158(.din(G158), .dout(new_new_n2356__));
  buf1  g0159(.din(G159), .dout(new_new_n2358__));
  buf1  g0160(.din(G160), .dout(new_new_n2360__));
  buf1  g0161(.din(G161), .dout(new_new_n2362__));
  buf1  g0162(.din(G162), .dout(new_new_n2364__));
  buf1  g0163(.din(G163), .dout(new_new_n2366__));
  buf1  g0164(.din(G164), .dout(new_new_n2368__));
  buf1  g0165(.din(G165), .dout(new_new_n2370__));
  buf1  g0166(.din(G166), .dout(new_new_n2372__));
  buf1  g0167(.din(G167), .dout(new_new_n2374__));
  buf1  g0168(.din(G168), .dout(new_new_n2376__));
  buf1  g0169(.din(G169), .dout(new_new_n2378__));
  buf1  g0170(.din(G170), .dout(new_new_n2380__));
  buf1  g0171(.din(G171), .dout(new_new_n2382__));
  buf1  g0172(.din(G172), .dout(new_new_n2384__));
  buf1  g0173(.din(G173), .dout(new_new_n2386__));
  buf1  g0174(.din(G174), .dout(new_new_n2388__));
  buf1  g0175(.din(G175), .dout(new_new_n2390__));
  buf1  g0176(.din(G176), .dout(new_new_n2392__));
  buf1  g0177(.din(G177), .dout(new_new_n2394__));
  buf1  g0178(.din(G178), .dout(new_new_n2396__));
  buf1  g0179(.din(n2610_lo), .dout(new_new_n2398__));
  buf1  g0180(.din(n2613_lo), .dout(new_new_n2400__));
  buf1  g0181(.din(n2616_lo), .dout(new_new_n2402__));
  buf1  g0182(.din(n2619_lo), .dout(new_new_n2404__));
  not1  g0183(.din(n2619_lo), .dout(new_new_n2405__));
  buf1  g0184(.din(n2622_lo), .dout(new_new_n2406__));
  buf1  g0185(.din(n2625_lo), .dout(new_new_n2408__));
  buf1  g0186(.din(n2628_lo), .dout(new_new_n2410__));
  not1  g0187(.din(n2628_lo), .dout(new_new_n2411__));
  buf1  g0188(.din(n2634_lo), .dout(new_new_n2412__));
  buf1  g0189(.din(n2637_lo), .dout(new_new_n2414__));
  buf1  g0190(.din(n2640_lo), .dout(new_new_n2416__));
  buf1  g0191(.din(n2643_lo), .dout(new_new_n2418__));
  buf1  g0192(.din(n2646_lo), .dout(new_new_n2420__));
  buf1  g0193(.din(n2649_lo), .dout(new_new_n2422__));
  buf1  g0194(.din(n2652_lo), .dout(new_new_n2424__));
  not1  g0195(.din(n2655_lo), .dout(new_new_n2427__));
  buf1  g0196(.din(n2658_lo), .dout(new_new_n2428__));
  buf1  g0197(.din(n2661_lo), .dout(new_new_n2430__));
  buf1  g0198(.din(n2664_lo), .dout(new_new_n2432__));
  buf1  g0199(.din(n2667_lo), .dout(new_new_n2434__));
  buf1  g0200(.din(n2670_lo), .dout(new_new_n2436__));
  buf1  g0201(.din(n2673_lo), .dout(new_new_n2438__));
  buf1  g0202(.din(n2676_lo), .dout(new_new_n2440__));
  buf1  g0203(.din(n2679_lo), .dout(new_new_n2442__));
  buf1  g0204(.din(n2682_lo), .dout(new_new_n2444__));
  buf1  g0205(.din(n2685_lo), .dout(new_new_n2446__));
  buf1  g0206(.din(n2688_lo), .dout(new_new_n2448__));
  buf1  g0207(.din(n2691_lo), .dout(new_new_n2450__));
  buf1  g0208(.din(n2694_lo), .dout(new_new_n2452__));
  buf1  g0209(.din(n2697_lo), .dout(new_new_n2454__));
  buf1  g0210(.din(n2700_lo), .dout(new_new_n2456__));
  buf1  g0211(.din(n2703_lo), .dout(new_new_n2458__));
  buf1  g0212(.din(n2706_lo), .dout(new_new_n2460__));
  buf1  g0213(.din(n2709_lo), .dout(new_new_n2462__));
  buf1  g0214(.din(n2712_lo), .dout(new_new_n2464__));
  buf1  g0215(.din(n2715_lo), .dout(new_new_n2466__));
  buf1  g0216(.din(n2718_lo), .dout(new_new_n2468__));
  buf1  g0217(.din(n2721_lo), .dout(new_new_n2470__));
  buf1  g0218(.din(n2724_lo), .dout(new_new_n2472__));
  buf1  g0219(.din(n2727_lo), .dout(new_new_n2474__));
  buf1  g0220(.din(n2730_lo), .dout(new_new_n2476__));
  buf1  g0221(.din(n2733_lo), .dout(new_new_n2478__));
  buf1  g0222(.din(n2736_lo), .dout(new_new_n2480__));
  not1  g0223(.din(n2739_lo), .dout(new_new_n2483__));
  buf1  g0224(.din(n2742_lo), .dout(new_new_n2484__));
  buf1  g0225(.din(n2745_lo), .dout(new_new_n2486__));
  buf1  g0226(.din(n2748_lo), .dout(new_new_n2488__));
  not1  g0227(.din(n2751_lo), .dout(new_new_n2491__));
  buf1  g0228(.din(n2754_lo), .dout(new_new_n2492__));
  buf1  g0229(.din(n2757_lo), .dout(new_new_n2494__));
  buf1  g0230(.din(n2760_lo), .dout(new_new_n2496__));
  not1  g0231(.din(n2763_lo), .dout(new_new_n2499__));
  buf1  g0232(.din(n2766_lo), .dout(new_new_n2500__));
  buf1  g0233(.din(n2769_lo), .dout(new_new_n2502__));
  buf1  g0234(.din(n2772_lo), .dout(new_new_n2504__));
  buf1  g0235(.din(n2775_lo), .dout(new_new_n2506__));
  buf1  g0236(.din(n2778_lo), .dout(new_new_n2508__));
  buf1  g0237(.din(n2781_lo), .dout(new_new_n2510__));
  buf1  g0238(.din(n2784_lo), .dout(new_new_n2512__));
  buf1  g0239(.din(n2787_lo), .dout(new_new_n2514__));
  buf1  g0240(.din(n2790_lo), .dout(new_new_n2516__));
  buf1  g0241(.din(n2793_lo), .dout(new_new_n2518__));
  buf1  g0242(.din(n2796_lo), .dout(new_new_n2520__));
  buf1  g0243(.din(n2799_lo), .dout(new_new_n2522__));
  buf1  g0244(.din(n2802_lo), .dout(new_new_n2524__));
  buf1  g0245(.din(n2805_lo), .dout(new_new_n2526__));
  buf1  g0246(.din(n2808_lo), .dout(new_new_n2528__));
  buf1  g0247(.din(n2811_lo), .dout(new_new_n2530__));
  buf1  g0248(.din(n2814_lo), .dout(new_new_n2532__));
  buf1  g0249(.din(n2817_lo), .dout(new_new_n2534__));
  buf1  g0250(.din(n2820_lo), .dout(new_new_n2536__));
  buf1  g0251(.din(n2823_lo), .dout(new_new_n2538__));
  buf1  g0252(.din(n2826_lo), .dout(new_new_n2540__));
  buf1  g0253(.din(n2829_lo), .dout(new_new_n2542__));
  buf1  g0254(.din(n2832_lo), .dout(new_new_n2544__));
  buf1  g0255(.din(n2838_lo), .dout(new_new_n2546__));
  buf1  g0256(.din(n2841_lo), .dout(new_new_n2548__));
  buf1  g0257(.din(n2844_lo), .dout(new_new_n2550__));
  buf1  g0258(.din(n2847_lo), .dout(new_new_n2552__));
  buf1  g0259(.din(n2850_lo), .dout(new_new_n2554__));
  buf1  g0260(.din(n2853_lo), .dout(new_new_n2556__));
  buf1  g0261(.din(n2856_lo), .dout(new_new_n2558__));
  not1  g0262(.din(n2856_lo), .dout(new_new_n2559__));
  buf1  g0263(.din(n2862_lo), .dout(new_new_n2560__));
  buf1  g0264(.din(n2865_lo), .dout(new_new_n2562__));
  buf1  g0265(.din(n2868_lo), .dout(new_new_n2564__));
  buf1  g0266(.din(n2871_lo), .dout(new_new_n2566__));
  buf1  g0267(.din(n2874_lo), .dout(new_new_n2568__));
  buf1  g0268(.din(n2877_lo), .dout(new_new_n2570__));
  buf1  g0269(.din(n2880_lo), .dout(new_new_n2572__));
  not1  g0270(.din(n2883_lo), .dout(new_new_n2575__));
  buf1  g0271(.din(n2886_lo), .dout(new_new_n2576__));
  buf1  g0272(.din(n2889_lo), .dout(new_new_n2578__));
  buf1  g0273(.din(n2892_lo), .dout(new_new_n2580__));
  not1  g0274(.din(n2895_lo), .dout(new_new_n2583__));
  buf1  g0275(.din(n2898_lo), .dout(new_new_n2584__));
  buf1  g0276(.din(n2901_lo), .dout(new_new_n2586__));
  buf1  g0277(.din(n2904_lo), .dout(new_new_n2588__));
  not1  g0278(.din(n2907_lo), .dout(new_new_n2591__));
  buf1  g0279(.din(n2910_lo), .dout(new_new_n2592__));
  buf1  g0280(.din(n2913_lo), .dout(new_new_n2594__));
  buf1  g0281(.din(n2916_lo), .dout(new_new_n2596__));
  buf1  g0282(.din(n2919_lo), .dout(new_new_n2598__));
  buf1  g0283(.din(n2922_lo), .dout(new_new_n2600__));
  buf1  g0284(.din(n2925_lo), .dout(new_new_n2602__));
  buf1  g0285(.din(n2928_lo), .dout(new_new_n2604__));
  buf1  g0286(.din(n2931_lo), .dout(new_new_n2606__));
  buf1  g0287(.din(n2934_lo), .dout(new_new_n2608__));
  buf1  g0288(.din(n2937_lo), .dout(new_new_n2610__));
  buf1  g0289(.din(n2940_lo), .dout(new_new_n2612__));
  buf1  g0290(.din(n2943_lo), .dout(new_new_n2614__));
  buf1  g0291(.din(n2946_lo), .dout(new_new_n2616__));
  buf1  g0292(.din(n2949_lo), .dout(new_new_n2618__));
  buf1  g0293(.din(n2952_lo), .dout(new_new_n2620__));
  buf1  g0294(.din(n2955_lo), .dout(new_new_n2622__));
  buf1  g0295(.din(n2958_lo), .dout(new_new_n2624__));
  buf1  g0296(.din(n2961_lo), .dout(new_new_n2626__));
  buf1  g0297(.din(n2964_lo), .dout(new_new_n2628__));
  buf1  g0298(.din(n2967_lo), .dout(new_new_n2630__));
  buf1  g0299(.din(n2970_lo), .dout(new_new_n2632__));
  buf1  g0300(.din(n2973_lo), .dout(new_new_n2634__));
  buf1  g0301(.din(n2976_lo), .dout(new_new_n2636__));
  buf1  g0302(.din(n2979_lo), .dout(new_new_n2638__));
  buf1  g0303(.din(n2982_lo), .dout(new_new_n2640__));
  buf1  g0304(.din(n2985_lo), .dout(new_new_n2642__));
  buf1  g0305(.din(n2988_lo), .dout(new_new_n2644__));
  not1  g0306(.din(n2991_lo), .dout(new_new_n2647__));
  buf1  g0307(.din(n2994_lo), .dout(new_new_n2648__));
  buf1  g0308(.din(n2997_lo), .dout(new_new_n2650__));
  buf1  g0309(.din(n3000_lo), .dout(new_new_n2652__));
  not1  g0310(.din(n3003_lo), .dout(new_new_n2655__));
  buf1  g0311(.din(n3006_lo), .dout(new_new_n2656__));
  buf1  g0312(.din(n3009_lo), .dout(new_new_n2658__));
  buf1  g0313(.din(n3012_lo), .dout(new_new_n2660__));
  not1  g0314(.din(n3015_lo), .dout(new_new_n2663__));
  buf1  g0315(.din(n3018_lo), .dout(new_new_n2664__));
  buf1  g0316(.din(n3021_lo), .dout(new_new_n2666__));
  buf1  g0317(.din(n3024_lo), .dout(new_new_n2668__));
  not1  g0318(.din(n3027_lo), .dout(new_new_n2671__));
  buf1  g0319(.din(n3030_lo), .dout(new_new_n2672__));
  buf1  g0320(.din(n3033_lo), .dout(new_new_n2674__));
  buf1  g0321(.din(n3036_lo), .dout(new_new_n2676__));
  buf1  g0322(.din(n3039_lo), .dout(new_new_n2678__));
  buf1  g0323(.din(n3042_lo), .dout(new_new_n2680__));
  buf1  g0324(.din(n3045_lo), .dout(new_new_n2682__));
  buf1  g0325(.din(n3048_lo), .dout(new_new_n2684__));
  not1  g0326(.din(n3051_lo), .dout(new_new_n2687__));
  buf1  g0327(.din(n3054_lo), .dout(new_new_n2688__));
  buf1  g0328(.din(n3057_lo), .dout(new_new_n2690__));
  buf1  g0329(.din(n3060_lo), .dout(new_new_n2692__));
  not1  g0330(.din(n3063_lo), .dout(new_new_n2695__));
  buf1  g0331(.din(n3066_lo), .dout(new_new_n2696__));
  buf1  g0332(.din(n3069_lo), .dout(new_new_n2698__));
  buf1  g0333(.din(n3072_lo), .dout(new_new_n2700__));
  buf1  g0334(.din(n3075_lo), .dout(new_new_n2702__));
  buf1  g0335(.din(n3078_lo), .dout(new_new_n2704__));
  buf1  g0336(.din(n3081_lo), .dout(new_new_n2706__));
  buf1  g0337(.din(n3084_lo), .dout(new_new_n2708__));
  buf1  g0338(.din(n3087_lo), .dout(new_new_n2710__));
  buf1  g0339(.din(n3090_lo), .dout(new_new_n2712__));
  buf1  g0340(.din(n3093_lo), .dout(new_new_n2714__));
  buf1  g0341(.din(n3096_lo), .dout(new_new_n2716__));
  buf1  g0342(.din(n3099_lo), .dout(new_new_n2718__));
  buf1  g0343(.din(n3102_lo), .dout(new_new_n2720__));
  buf1  g0344(.din(n3105_lo), .dout(new_new_n2722__));
  buf1  g0345(.din(n3108_lo), .dout(new_new_n2724__));
  buf1  g0346(.din(n3111_lo), .dout(new_new_n2726__));
  buf1  g0347(.din(n3114_lo), .dout(new_new_n2728__));
  buf1  g0348(.din(n3117_lo), .dout(new_new_n2730__));
  buf1  g0349(.din(n3120_lo), .dout(new_new_n2732__));
  buf1  g0350(.din(n3126_lo), .dout(new_new_n2734__));
  buf1  g0351(.din(n3129_lo), .dout(new_new_n2736__));
  buf1  g0352(.din(n3132_lo), .dout(new_new_n2738__));
  buf1  g0353(.din(n3138_lo), .dout(new_new_n2740__));
  buf1  g0354(.din(n3141_lo), .dout(new_new_n2742__));
  buf1  g0355(.din(n3144_lo), .dout(new_new_n2744__));
  buf1  g0356(.din(n3147_lo), .dout(new_new_n2746__));
  buf1  g0357(.din(n3150_lo), .dout(new_new_n2748__));
  buf1  g0358(.din(n3153_lo), .dout(new_new_n2750__));
  buf1  g0359(.din(n3156_lo), .dout(new_new_n2752__));
  buf1  g0360(.din(n3162_lo), .dout(new_new_n2754__));
  buf1  g0361(.din(n3165_lo), .dout(new_new_n2756__));
  buf1  g0362(.din(n3168_lo), .dout(new_new_n2758__));
  buf1  g0363(.din(n3174_lo), .dout(new_new_n2760__));
  buf1  g0364(.din(n3177_lo), .dout(new_new_n2762__));
  buf1  g0365(.din(n3180_lo), .dout(new_new_n2764__));
  buf1  g0366(.din(n3186_lo), .dout(new_new_n2766__));
  buf1  g0367(.din(n3189_lo), .dout(new_new_n2768__));
  buf1  g0368(.din(n3192_lo), .dout(new_new_n2770__));
  buf1  g0369(.din(n3195_lo), .dout(new_new_n2772__));
  buf1  g0370(.din(n3198_lo), .dout(new_new_n2774__));
  buf1  g0371(.din(n3201_lo), .dout(new_new_n2776__));
  buf1  g0372(.din(n3204_lo), .dout(new_new_n2778__));
  buf1  g0373(.din(n3210_lo), .dout(new_new_n2780__));
  buf1  g0374(.din(n3213_lo), .dout(new_new_n2782__));
  buf1  g0375(.din(n3216_lo), .dout(new_new_n2784__));
  buf1  g0376(.din(n3219_lo), .dout(new_new_n2786__));
  buf1  g0377(.din(n3222_lo), .dout(new_new_n2788__));
  buf1  g0378(.din(n3225_lo), .dout(new_new_n2790__));
  buf1  g0379(.din(n3228_lo), .dout(new_new_n2792__));
  buf1  g0380(.din(n3234_lo), .dout(new_new_n2794__));
  buf1  g0381(.din(n3237_lo), .dout(new_new_n2796__));
  buf1  g0382(.din(n3240_lo), .dout(new_new_n2798__));
  buf1  g0383(.din(n3243_lo), .dout(new_new_n2800__));
  buf1  g0384(.din(n3246_lo), .dout(new_new_n2802__));
  buf1  g0385(.din(n3249_lo), .dout(new_new_n2804__));
  buf1  g0386(.din(n3252_lo), .dout(new_new_n2806__));
  buf1  g0387(.din(n3255_lo), .dout(new_new_n2808__));
  buf1  g0388(.din(n3258_lo), .dout(new_new_n2810__));
  buf1  g0389(.din(n3261_lo), .dout(new_new_n2812__));
  buf1  g0390(.din(n3264_lo), .dout(new_new_n2814__));
  not1  g0391(.din(n3267_lo), .dout(new_new_n2817__));
  buf1  g0392(.din(n3270_lo), .dout(new_new_n2818__));
  buf1  g0393(.din(n3273_lo), .dout(new_new_n2820__));
  buf1  g0394(.din(n3276_lo), .dout(new_new_n2822__));
  buf1  g0395(.din(n3279_lo), .dout(new_new_n2824__));
  buf1  g0396(.din(n3282_lo), .dout(new_new_n2826__));
  buf1  g0397(.din(n3285_lo), .dout(new_new_n2828__));
  buf1  g0398(.din(n3288_lo), .dout(new_new_n2830__));
  buf1  g0399(.din(n3294_lo), .dout(new_new_n2832__));
  buf1  g0400(.din(n3297_lo), .dout(new_new_n2834__));
  buf1  g0401(.din(n3300_lo), .dout(new_new_n2836__));
  buf1  g0402(.din(n3306_lo), .dout(new_new_n2838__));
  buf1  g0403(.din(n3309_lo), .dout(new_new_n2840__));
  not1  g0404(.din(n3312_lo), .dout(new_new_n2843__));
  buf1  g0405(.din(n3318_lo), .dout(new_new_n2844__));
  buf1  g0406(.din(n3321_lo), .dout(new_new_n2846__));
  buf1  g0407(.din(n3324_lo), .dout(new_new_n2848__));
  buf1  g0408(.din(n3330_lo), .dout(new_new_n2850__));
  buf1  g0409(.din(n3333_lo), .dout(new_new_n2852__));
  buf1  g0410(.din(n3336_lo), .dout(new_new_n2854__));
  buf1  g0411(.din(n3339_lo), .dout(new_new_n2856__));
  not1  g0412(.din(n3339_lo), .dout(new_new_n2857__));
  buf1  g0413(.din(n3342_lo), .dout(new_new_n2858__));
  buf1  g0414(.din(n3345_lo), .dout(new_new_n2860__));
  buf1  g0415(.din(n3348_lo), .dout(new_new_n2862__));
  not1  g0416(.din(n3351_lo), .dout(new_new_n2865__));
  buf1  g0417(.din(n3354_lo), .dout(new_new_n2866__));
  buf1  g0418(.din(n3357_lo), .dout(new_new_n2868__));
  buf1  g0419(.din(n3360_lo), .dout(new_new_n2870__));
  buf1  g0420(.din(n3363_lo), .dout(new_new_n2872__));
  buf1  g0421(.din(n3366_lo), .dout(new_new_n2874__));
  buf1  g0422(.din(n3369_lo), .dout(new_new_n2876__));
  buf1  g0423(.din(n3372_lo), .dout(new_new_n2878__));
  buf1  g0424(.din(n3375_lo), .dout(new_new_n2880__));
  not1  g0425(.din(n3375_lo), .dout(new_new_n2881__));
  buf1  g0426(.din(n3378_lo), .dout(new_new_n2882__));
  buf1  g0427(.din(n3381_lo), .dout(new_new_n2884__));
  buf1  g0428(.din(n3384_lo), .dout(new_new_n2886__));
  not1  g0429(.din(n3387_lo), .dout(new_new_n2889__));
  buf1  g0430(.din(n3390_lo), .dout(new_new_n2890__));
  buf1  g0431(.din(n3393_lo), .dout(new_new_n2892__));
  buf1  g0432(.din(n3396_lo), .dout(new_new_n2894__));
  buf1  g0433(.din(n3399_lo), .dout(new_new_n2896__));
  not1  g0434(.din(n3399_lo), .dout(new_new_n2897__));
  buf1  g0435(.din(n3402_lo), .dout(new_new_n2898__));
  buf1  g0436(.din(n3405_lo), .dout(new_new_n2900__));
  buf1  g0437(.din(n3408_lo), .dout(new_new_n2902__));
  buf1  g0438(.din(n3411_lo), .dout(new_new_n2904__));
  buf1  g0439(.din(n3414_lo), .dout(new_new_n2906__));
  buf1  g0440(.din(n3417_lo), .dout(new_new_n2908__));
  buf1  g0441(.din(n3420_lo), .dout(new_new_n2910__));
  buf1  g0442(.din(n3423_lo), .dout(new_new_n2912__));
  buf1  g0443(.din(n3426_lo), .dout(new_new_n2914__));
  buf1  g0444(.din(n3429_lo), .dout(new_new_n2916__));
  buf1  g0445(.din(n3432_lo), .dout(new_new_n2918__));
  buf1  g0446(.din(n3435_lo), .dout(new_new_n2920__));
  buf1  g0447(.din(n3438_lo), .dout(new_new_n2922__));
  buf1  g0448(.din(n3441_lo), .dout(new_new_n2924__));
  buf1  g0449(.din(n3444_lo), .dout(new_new_n2926__));
  buf1  g0450(.din(n3447_lo), .dout(new_new_n2928__));
  buf1  g0451(.din(n3450_lo), .dout(new_new_n2930__));
  buf1  g0452(.din(n3453_lo), .dout(new_new_n2932__));
  buf1  g0453(.din(n3456_lo), .dout(new_new_n2934__));
  buf1  g0454(.din(n3459_lo), .dout(new_new_n2936__));
  buf1  g0455(.din(n3462_lo), .dout(new_new_n2938__));
  buf1  g0456(.din(n3465_lo), .dout(new_new_n2940__));
  buf1  g0457(.din(n3468_lo), .dout(new_new_n2942__));
  not1  g0458(.din(n3471_lo), .dout(new_new_n2945__));
  buf1  g0459(.din(n3474_lo), .dout(new_new_n2946__));
  buf1  g0460(.din(n3477_lo), .dout(new_new_n2948__));
  buf1  g0461(.din(n3480_lo), .dout(new_new_n2950__));
  buf1  g0462(.din(n3483_lo), .dout(new_new_n2952__));
  buf1  g0463(.din(n3486_lo), .dout(new_new_n2954__));
  buf1  g0464(.din(n3489_lo), .dout(new_new_n2956__));
  buf1  g0465(.din(n3492_lo), .dout(new_new_n2958__));
  buf1  g0466(.din(n3495_lo), .dout(new_new_n2960__));
  buf1  g0467(.din(n3498_lo), .dout(new_new_n2962__));
  buf1  g0468(.din(n3501_lo), .dout(new_new_n2964__));
  buf1  g0469(.din(n3504_lo), .dout(new_new_n2966__));
  buf1  g0470(.din(n3507_lo), .dout(new_new_n2968__));
  buf1  g0471(.din(n3510_lo), .dout(new_new_n2970__));
  buf1  g0472(.din(n3513_lo), .dout(new_new_n2972__));
  buf1  g0473(.din(n3516_lo), .dout(new_new_n2974__));
  buf1  g0474(.din(n3519_lo), .dout(new_new_n2976__));
  buf1  g0475(.din(n3522_lo), .dout(new_new_n2978__));
  buf1  g0476(.din(n3525_lo), .dout(new_new_n2980__));
  buf1  g0477(.din(n3528_lo), .dout(new_new_n2982__));
  buf1  g0478(.din(n3531_lo), .dout(new_new_n2984__));
  buf1  g0479(.din(n3534_lo), .dout(new_new_n2986__));
  buf1  g0480(.din(n3537_lo), .dout(new_new_n2988__));
  buf1  g0481(.din(n3540_lo), .dout(new_new_n2990__));
  not1  g0482(.din(n3543_lo), .dout(new_new_n2993__));
  buf1  g0483(.din(n3546_lo), .dout(new_new_n2994__));
  buf1  g0484(.din(n3549_lo), .dout(new_new_n2996__));
  buf1  g0485(.din(n3552_lo), .dout(new_new_n2998__));
  not1  g0486(.din(n3555_lo), .dout(new_new_n3001__));
  buf1  g0487(.din(n3558_lo), .dout(new_new_n3002__));
  buf1  g0488(.din(n3561_lo), .dout(new_new_n3004__));
  buf1  g0489(.din(n3564_lo), .dout(new_new_n3006__));
  buf1  g0490(.din(n3567_lo), .dout(new_new_n3008__));
  buf1  g0491(.din(n3570_lo), .dout(new_new_n3010__));
  buf1  g0492(.din(n3573_lo), .dout(new_new_n3012__));
  buf1  g0493(.din(n3576_lo), .dout(new_new_n3014__));
  buf1  g0494(.din(n3579_lo), .dout(new_new_n3016__));
  buf1  g0495(.din(n3582_lo), .dout(new_new_n3018__));
  buf1  g0496(.din(n3585_lo), .dout(new_new_n3020__));
  buf1  g0497(.din(n3588_lo), .dout(new_new_n3022__));
  not1  g0498(.din(n3591_lo), .dout(new_new_n3025__));
  buf1  g0499(.din(n3594_lo), .dout(new_new_n3026__));
  buf1  g0500(.din(n3597_lo), .dout(new_new_n3028__));
  buf1  g0501(.din(n3600_lo), .dout(new_new_n3030__));
  buf1  g0502(.din(n3603_lo), .dout(new_new_n3032__));
  buf1  g0503(.din(n3606_lo), .dout(new_new_n3034__));
  buf1  g0504(.din(n3609_lo), .dout(new_new_n3036__));
  buf1  g0505(.din(n3612_lo), .dout(new_new_n3038__));
  buf1  g0506(.din(n3615_lo), .dout(new_new_n3040__));
  buf1  g0507(.din(n3618_lo), .dout(new_new_n3042__));
  buf1  g0508(.din(n3621_lo), .dout(new_new_n3044__));
  buf1  g0509(.din(n3624_lo), .dout(new_new_n3046__));
  buf1  g0510(.din(n3627_lo), .dout(new_new_n3048__));
  buf1  g0511(.din(n3630_lo), .dout(new_new_n3050__));
  buf1  g0512(.din(n3633_lo), .dout(new_new_n3052__));
  buf1  g0513(.din(n3636_lo), .dout(new_new_n3054__));
  buf1  g0514(.din(n3639_lo), .dout(new_new_n3056__));
  buf1  g0515(.din(n3642_lo), .dout(new_new_n3058__));
  buf1  g0516(.din(n3645_lo), .dout(new_new_n3060__));
  buf1  g0517(.din(n3648_lo), .dout(new_new_n3062__));
  buf1  g0518(.din(n3651_lo), .dout(new_new_n3064__));
  buf1  g0519(.din(n3654_lo), .dout(new_new_n3066__));
  buf1  g0520(.din(n3666_lo), .dout(new_new_n3068__));
  buf1  g0521(.din(n3750_lo), .dout(new_new_n3070__));
  buf1  g0522(.din(n3762_lo), .dout(new_new_n3072__));
  buf1  g0523(.din(n3774_lo), .dout(new_new_n3074__));
  buf1  g0524(.din(n3786_lo), .dout(new_new_n3076__));
  buf1  g0525(.din(n3789_lo), .dout(new_new_n3078__));
  buf1  g0526(.din(n3792_lo), .dout(new_new_n3080__));
  not1  g0527(.din(n3795_lo), .dout(new_new_n3083__));
  buf1  g0528(.din(n3798_lo), .dout(new_new_n3084__));
  buf1  g0529(.din(n3810_lo), .dout(new_new_n3086__));
  buf1  g0530(.din(n3822_lo), .dout(new_new_n3088__));
  buf1  g0531(.din(n3834_lo), .dout(new_new_n3090__));
  not1  g0532(.din(n3834_lo), .dout(new_new_n3091__));
  buf1  g0533(.din(n3846_lo), .dout(new_new_n3092__));
  not1  g0534(.din(n3846_lo), .dout(new_new_n3093__));
  buf1  g0535(.din(n3930_lo), .dout(new_new_n3094__));
  buf1  g0536(.din(n3933_lo), .dout(new_new_n3096__));
  buf1  g0537(.din(n3936_lo), .dout(new_new_n3098__));
  not1  g0538(.din(n3936_lo), .dout(new_new_n3099__));
  buf1  g0539(.din(n3942_lo), .dout(new_new_n3100__));
  buf1  g0540(.din(n3945_lo), .dout(new_new_n3102__));
  buf1  g0541(.din(n3948_lo), .dout(new_new_n3104__));
  not1  g0542(.din(n3948_lo), .dout(new_new_n3105__));
  buf1  g0543(.din(n3954_lo), .dout(new_new_n3106__));
  buf1  g0544(.din(n3957_lo), .dout(new_new_n3108__));
  not1  g0545(.din(n3957_lo), .dout(new_new_n3109__));
  not1  g0546(.din(n3963_lo), .dout(new_new_n3111__));
  buf1  g0547(.din(n3966_lo), .dout(new_new_n3112__));
  buf1  g0548(.din(n3969_lo), .dout(new_new_n3114__));
  buf1  g0549(.din(n3975_lo), .dout(new_new_n3116__));
  not1  g0550(.din(n3975_lo), .dout(new_new_n3117__));
  buf1  g0551(.din(n3978_lo), .dout(new_new_n3118__));
  buf1  g0552(.din(n3990_lo), .dout(new_new_n3120__));
  buf1  g0553(.din(n4050_lo), .dout(new_new_n3122__));
  buf1  g0554(.din(n4062_lo), .dout(new_new_n3124__));
  buf1  g0555(.din(n4098_lo), .dout(new_new_n3126__));
  not1  g0556(.din(n4098_lo), .dout(new_new_n3127__));
  not1  g0557(.din(n4107_lo), .dout(new_new_n3129__));
  buf1  g0558(.din(n4110_lo), .dout(new_new_n3130__));
  not1  g0559(.din(n4110_lo), .dout(new_new_n3131__));
  buf1  g0560(.din(n4122_lo), .dout(new_new_n3132__));
  not1  g0561(.din(n4122_lo), .dout(new_new_n3133__));
  not1  g0562(.din(n4131_lo), .dout(new_new_n3135__));
  not1  g0563(.din(n4155_lo), .dout(new_new_n3137__));
  buf1  g0564(.din(n4158_lo), .dout(new_new_n3138__));
  not1  g0565(.din(n4158_lo), .dout(new_new_n3139__));
  buf1  g0566(.din(n4170_lo), .dout(new_new_n3140__));
  not1  g0567(.din(n4170_lo), .dout(new_new_n3141__));
  not1  g0568(.din(n4179_lo), .dout(new_new_n3143__));
  buf1  g0569(.din(n4182_lo), .dout(new_new_n3144__));
  buf1  g0570(.din(n4185_lo), .dout(new_new_n3146__));
  buf1  g0571(.din(n4188_lo), .dout(new_new_n3148__));
  not1  g0572(.din(n4188_lo), .dout(new_new_n3149__));
  buf1  g0573(.din(n4194_lo), .dout(new_new_n3150__));
  buf1  g0574(.din(n4197_lo), .dout(new_new_n3152__));
  buf1  g0575(.din(n4200_lo), .dout(new_new_n3154__));
  buf1  g0576(.din(n4206_lo), .dout(new_new_n3156__));
  buf1  g0577(.din(n4209_lo), .dout(new_new_n3158__));
  buf1  g0578(.din(n4212_lo), .dout(new_new_n3160__));
  buf1  g0579(.din(n4215_lo), .dout(new_new_n3162__));
  buf1  g0580(.din(n4230_lo), .dout(new_new_n3164__));
  buf1  g0581(.din(n4233_lo), .dout(new_new_n3166__));
  buf1  g0582(.din(n4236_lo), .dout(new_new_n3168__));
  not1  g0583(.din(n4239_lo), .dout(new_new_n3171__));
  buf1  g0584(.din(n4242_lo), .dout(new_new_n3172__));
  not1  g0585(.din(n4242_lo), .dout(new_new_n3173__));
  buf1  g0586(.din(n4254_lo), .dout(new_new_n3174__));
  not1  g0587(.din(n4254_lo), .dout(new_new_n3175__));
  buf1  g0588(.din(n4290_lo), .dout(new_new_n3176__));
  buf1  g0589(.din(n4293_lo), .dout(new_new_n3178__));
  not1  g0590(.din(n4293_lo), .dout(new_new_n3179__));
  buf1  g0591(.din(n4302_lo), .dout(new_new_n3180__));
  buf1  g0592(.din(n4314_lo), .dout(new_new_n3182__));
  not1  g0593(.din(n4314_lo), .dout(new_new_n3183__));
  buf1  g0594(.din(n4350_lo), .dout(new_new_n3184__));
  buf1  g0595(.din(n4362_lo), .dout(new_new_n3186__));
  buf1  g0596(.din(n4374_lo), .dout(new_new_n3188__));
  not1  g0597(.din(n4374_lo), .dout(new_new_n3189__));
  buf1  g0598(.din(n4386_lo), .dout(new_new_n3190__));
  not1  g0599(.din(n4386_lo), .dout(new_new_n3191__));
  buf1  g0600(.din(n4398_lo), .dout(new_new_n3192__));
  not1  g0601(.din(n4398_lo), .dout(new_new_n3193__));
  buf1  g0602(.din(n4410_lo), .dout(new_new_n3194__));
  buf1  g0603(.din(n4413_lo), .dout(new_new_n3196__));
  buf1  g0604(.din(n4416_lo), .dout(new_new_n3198__));
  not1  g0605(.din(n4419_lo), .dout(new_new_n3201__));
  buf1  g0606(.din(n4422_lo), .dout(new_new_n3202__));
  buf1  g0607(.din(n4425_lo), .dout(new_new_n3204__));
  buf1  g0608(.din(n4428_lo), .dout(new_new_n3206__));
  buf1  g0609(.din(n4431_lo), .dout(new_new_n3208__));
  not1  g0610(.din(n4431_lo), .dout(new_new_n3209__));
  buf1  g0611(.din(n4434_lo), .dout(new_new_n3210__));
  buf1  g0612(.din(n4437_lo), .dout(new_new_n3212__));
  buf1  g0613(.din(n4440_lo), .dout(new_new_n3214__));
  not1  g0614(.din(n4443_lo), .dout(new_new_n3217__));
  buf1  g0615(.din(n4446_lo), .dout(new_new_n3218__));
  buf1  g0616(.din(n4449_lo), .dout(new_new_n3220__));
  buf1  g0617(.din(n4452_lo), .dout(new_new_n3222__));
  not1  g0618(.din(n4455_lo), .dout(new_new_n3225__));
  buf1  g0619(.din(n4458_lo), .dout(new_new_n3226__));
  buf1  g0620(.din(n4461_lo), .dout(new_new_n3228__));
  buf1  g0621(.din(n4464_lo), .dout(new_new_n3230__));
  not1  g0622(.din(n4467_lo), .dout(new_new_n3233__));
  buf1  g0623(.din(n4470_lo), .dout(new_new_n3234__));
  buf1  g0624(.din(n4473_lo), .dout(new_new_n3236__));
  buf1  g0625(.din(n4476_lo), .dout(new_new_n3238__));
  not1  g0626(.din(n4479_lo), .dout(new_new_n3241__));
  buf1  g0627(.din(n4482_lo), .dout(new_new_n3242__));
  buf1  g0628(.din(n4485_lo), .dout(new_new_n3244__));
  buf1  g0629(.din(n4488_lo), .dout(new_new_n3246__));
  not1  g0630(.din(n4488_lo), .dout(new_new_n3247__));
  buf1  g0631(.din(n4494_lo), .dout(new_new_n3248__));
  buf1  g0632(.din(n4497_lo), .dout(new_new_n3250__));
  buf1  g0633(.din(n4500_lo), .dout(new_new_n3252__));
  buf1  g0634(.din(n4503_lo), .dout(new_new_n3254__));
  not1  g0635(.din(n4503_lo), .dout(new_new_n3255__));
  buf1  g0636(.din(n4506_lo), .dout(new_new_n3256__));
  buf1  g0637(.din(n4509_lo), .dout(new_new_n3258__));
  buf1  g0638(.din(n4512_lo), .dout(new_new_n3260__));
  buf1  g0639(.din(n4515_lo), .dout(new_new_n3262__));
  not1  g0640(.din(n4515_lo), .dout(new_new_n3263__));
  buf1  g0641(.din(n4518_lo), .dout(new_new_n3264__));
  buf1  g0642(.din(n4521_lo), .dout(new_new_n3266__));
  buf1  g0643(.din(n4524_lo), .dout(new_new_n3268__));
  buf1  g0644(.din(n4527_lo), .dout(new_new_n3270__));
  not1  g0645(.din(n4527_lo), .dout(new_new_n3271__));
  buf1  g0646(.din(n4530_lo), .dout(new_new_n3272__));
  buf1  g0647(.din(n4533_lo), .dout(new_new_n3274__));
  buf1  g0648(.din(n4536_lo), .dout(new_new_n3276__));
  buf1  g0649(.din(n4539_lo), .dout(new_new_n3278__));
  not1  g0650(.din(n4539_lo), .dout(new_new_n3279__));
  buf1  g0651(.din(n4542_lo), .dout(new_new_n3280__));
  buf1  g0652(.din(n4545_lo), .dout(new_new_n3282__));
  not1  g0653(.din(n4545_lo), .dout(new_new_n3283__));
  buf1  g0654(.din(n4554_lo), .dout(new_new_n3284__));
  buf1  g0655(.din(n4557_lo), .dout(new_new_n3286__));
  buf1  g0656(.din(n4560_lo), .dout(new_new_n3288__));
  buf1  g0657(.din(n4563_lo), .dout(new_new_n3290__));
  not1  g0658(.din(n4563_lo), .dout(new_new_n3291__));
  buf1  g0659(.din(n4566_lo), .dout(new_new_n3292__));
  buf1  g0660(.din(n4569_lo), .dout(new_new_n3294__));
  buf1  g0661(.din(n4572_lo), .dout(new_new_n3296__));
  buf1  g0662(.din(n4575_lo), .dout(new_new_n3298__));
  buf1  g0663(.din(n4578_lo), .dout(new_new_n3300__));
  buf1  g0664(.din(n4581_lo), .dout(new_new_n3302__));
  buf1  g0665(.din(n4584_lo), .dout(new_new_n3304__));
  not1  g0666(.din(n4587_lo), .dout(new_new_n3307__));
  buf1  g0667(.din(n4590_lo), .dout(new_new_n3308__));
  buf1  g0668(.din(n4593_lo), .dout(new_new_n3310__));
  buf1  g0669(.din(n4596_lo), .dout(new_new_n3312__));
  buf1  g0670(.din(n4602_lo), .dout(new_new_n3314__));
  buf1  g0671(.din(n4605_lo), .dout(new_new_n3316__));
  buf1  g0672(.din(n4608_lo), .dout(new_new_n3318__));
  buf1  g0673(.din(n4614_lo), .dout(new_new_n3320__));
  buf1  g0674(.din(n4617_lo), .dout(new_new_n3322__));
  not1  g0675(.din(n4620_lo), .dout(new_new_n3325__));
  buf1  g0676(.din(n4626_lo), .dout(new_new_n3326__));
  buf1  g0677(.din(n4629_lo), .dout(new_new_n3328__));
  not1  g0678(.din(n4632_lo), .dout(new_new_n3331__));
  buf1  g0679(.din(n4638_lo), .dout(new_new_n3332__));
  buf1  g0680(.din(n4641_lo), .dout(new_new_n3334__));
  buf1  g0681(.din(n4644_lo), .dout(new_new_n3336__));
  buf1  g0682(.din(n4647_lo), .dout(new_new_n3338__));
  not1  g0683(.din(n4647_lo), .dout(new_new_n3339__));
  buf1  g0684(.din(n4650_lo), .dout(new_new_n3340__));
  buf1  g0685(.din(n4653_lo), .dout(new_new_n3342__));
  buf1  g0686(.din(n4656_lo), .dout(new_new_n3344__));
  buf1  g0687(.din(n4659_lo), .dout(new_new_n3346__));
  not1  g0688(.din(n4659_lo), .dout(new_new_n3347__));
  buf1  g0689(.din(n4662_lo), .dout(new_new_n3348__));
  buf1  g0690(.din(n4665_lo), .dout(new_new_n3350__));
  buf1  g0691(.din(n4668_lo), .dout(new_new_n3352__));
  buf1  g0692(.din(n4671_lo), .dout(new_new_n3354__));
  not1  g0693(.din(n4671_lo), .dout(new_new_n3355__));
  buf1  g0694(.din(n4674_lo), .dout(new_new_n3356__));
  buf1  g0695(.din(n4677_lo), .dout(new_new_n3358__));
  buf1  g0696(.din(n4680_lo), .dout(new_new_n3360__));
  buf1  g0697(.din(n4683_lo), .dout(new_new_n3362__));
  not1  g0698(.din(n4683_lo), .dout(new_new_n3363__));
  buf1  g0699(.din(n4686_lo), .dout(new_new_n3364__));
  buf1  g0700(.din(n4689_lo), .dout(new_new_n3366__));
  buf1  g0701(.din(n4692_lo), .dout(new_new_n3368__));
  buf1  g0702(.din(n4695_lo), .dout(new_new_n3370__));
  not1  g0703(.din(n4695_lo), .dout(new_new_n3371__));
  buf1  g0704(.din(n4698_lo), .dout(new_new_n3372__));
  buf1  g0705(.din(n4701_lo), .dout(new_new_n3374__));
  buf1  g0706(.din(n4704_lo), .dout(new_new_n3376__));
  buf1  g0707(.din(n4707_lo), .dout(new_new_n3378__));
  not1  g0708(.din(n4707_lo), .dout(new_new_n3379__));
  buf1  g0709(.din(n4710_lo), .dout(new_new_n3380__));
  buf1  g0710(.din(n4713_lo), .dout(new_new_n3382__));
  buf1  g0711(.din(n4716_lo), .dout(new_new_n3384__));
  not1  g0712(.din(n4716_lo), .dout(new_new_n3385__));
  buf1  g0713(.din(n4719_lo), .dout(new_new_n3386__));
  not1  g0714(.din(n4719_lo), .dout(new_new_n3387__));
  buf1  g0715(.din(n4722_lo), .dout(new_new_n3388__));
  buf1  g0716(.din(n4725_lo), .dout(new_new_n3390__));
  buf1  g0717(.din(n4728_lo), .dout(new_new_n3392__));
  not1  g0718(.din(n4728_lo), .dout(new_new_n3393__));
  buf1  g0719(.din(n4731_lo), .dout(new_new_n3394__));
  not1  g0720(.din(n4731_lo), .dout(new_new_n3395__));
  buf1  g0721(.din(n4734_lo), .dout(new_new_n3396__));
  buf1  g0722(.din(n4737_lo), .dout(new_new_n3398__));
  buf1  g0723(.din(n4740_lo), .dout(new_new_n3400__));
  not1  g0724(.din(n4743_lo), .dout(new_new_n3403__));
  buf1  g0725(.din(n4970_o2), .dout(new_new_n3404__));
  not1  g0726(.din(n4970_o2), .dout(new_new_n3405__));
  buf1  g0727(.din(n4972_o2), .dout(new_new_n3406__));
  not1  g0728(.din(n4972_o2), .dout(new_new_n3407__));
  buf1  g0729(.din(n4989_o2), .dout(new_new_n3408__));
  not1  g0730(.din(n4989_o2), .dout(new_new_n3409__));
  buf1  g0731(.din(n5024_o2), .dout(new_new_n3410__));
  not1  g0732(.din(n5024_o2), .dout(new_new_n3411__));
  buf1  g0733(.din(n5025_o2), .dout(new_new_n3412__));
  not1  g0734(.din(n5025_o2), .dout(new_new_n3413__));
  buf1  g0735(.din(n5029_o2), .dout(new_new_n3414__));
  not1  g0736(.din(n5029_o2), .dout(new_new_n3415__));
  not1  g0737(.din(n5042_o2), .dout(new_new_n3417__));
  not1  g0738(.din(n5048_o2), .dout(new_new_n3419__));
  buf1  g0739(.din(n5093_o2), .dout(new_new_n3420__));
  not1  g0740(.din(n5093_o2), .dout(new_new_n3421__));
  buf1  g0741(.din(n5096_o2), .dout(new_new_n3422__));
  not1  g0742(.din(n5096_o2), .dout(new_new_n3423__));
  not1  g0743(.din(n5193_o2), .dout(new_new_n3425__));
  buf1  g0744(.din(n5199_o2), .dout(new_new_n3426__));
  not1  g0745(.din(n5203_o2), .dout(new_new_n3429__));
  not1  g0746(.din(n5214_o2), .dout(new_new_n3431__));
  not1  g0747(.din(n5221_o2), .dout(new_new_n3433__));
  buf1  g0748(.din(n5222_o2), .dout(new_new_n3434__));
  not1  g0749(.din(n5273_o2), .dout(new_new_n3437__));
  buf1  g0750(.din(n5365_o2), .dout(new_new_n3438__));
  not1  g0751(.din(n5365_o2), .dout(new_new_n3439__));
  buf1  g0752(.din(n5385_o2), .dout(new_new_n3440__));
  buf1  g0753(.din(n5553_o2), .dout(new_new_n3442__));
  not1  g0754(.din(n5553_o2), .dout(new_new_n3443__));
  not1  g0755(.din(n5636_o2), .dout(new_new_n3445__));
  buf1  g0756(.din(n5782_o2), .dout(new_new_n3446__));
  buf1  g0757(.din(n5778_o2), .dout(new_new_n3448__));
  not1  g0758(.din(n5778_o2), .dout(new_new_n3449__));
  buf1  g0759(.din(n5323_o2), .dout(new_new_n3450__));
  not1  g0760(.din(n5323_o2), .dout(new_new_n3451__));
  buf1  g0761(.din(n5325_o2), .dout(new_new_n3452__));
  not1  g0762(.din(n5325_o2), .dout(new_new_n3453__));
  buf1  g0763(.din(n5327_o2), .dout(new_new_n3454__));
  not1  g0764(.din(n5327_o2), .dout(new_new_n3455__));
  buf1  g0765(.din(n5329_o2), .dout(new_new_n3456__));
  not1  g0766(.din(n5329_o2), .dout(new_new_n3457__));
  not1  g0767(.din(n5816_o2), .dout(new_new_n3459__));
  not1  g0768(.din(n5817_o2), .dout(new_new_n3461__));
  buf1  g0769(.din(n5837_o2), .dout(new_new_n3462__));
  not1  g0770(.din(n5837_o2), .dout(new_new_n3463__));
  buf1  g0771(.din(n5844_o2), .dout(new_new_n3464__));
  buf1  g0772(.din(n5859_o2), .dout(new_new_n3466__));
  buf1  g0773(.din(n5857_o2), .dout(new_new_n3468__));
  buf1  g0774(.din(n5369_o2), .dout(new_new_n3470__));
  not1  g0775(.din(n5369_o2), .dout(new_new_n3471__));
  buf1  g0776(.din(n5371_o2), .dout(new_new_n3472__));
  not1  g0777(.din(n5371_o2), .dout(new_new_n3473__));
  buf1  g0778(.din(n5373_o2), .dout(new_new_n3474__));
  not1  g0779(.din(n5373_o2), .dout(new_new_n3475__));
  buf1  g0780(.din(n5400_o2), .dout(new_new_n3476__));
  not1  g0781(.din(n5400_o2), .dout(new_new_n3477__));
  buf1  g0782(.din(n5402_o2), .dout(new_new_n3478__));
  not1  g0783(.din(n5402_o2), .dout(new_new_n3479__));
  buf1  g0784(.din(n5404_o2), .dout(new_new_n3480__));
  not1  g0785(.din(n5404_o2), .dout(new_new_n3481__));
  buf1  g0786(.din(n5406_o2), .dout(new_new_n3482__));
  not1  g0787(.din(n5406_o2), .dout(new_new_n3483__));
  buf1  g0788(.din(n5407_o2), .dout(new_new_n3484__));
  not1  g0789(.din(n5407_o2), .dout(new_new_n3485__));
  buf1  g0790(.din(n5408_o2), .dout(new_new_n3486__));
  not1  g0791(.din(n5408_o2), .dout(new_new_n3487__));
  not1  g0792(.din(n2722_o2), .dout(new_new_n3489__));
  buf1  g0793(.din(n1942_inv), .dout(new_new_n3490__));
  buf1  g0794(.din(n5412_o2), .dout(new_new_n3492__));
  not1  g0795(.din(n5412_o2), .dout(new_new_n3493__));
  buf1  g0796(.din(n1948_inv), .dout(new_new_n3494__));
  buf1  g0797(.din(n5557_o2), .dout(new_new_n3496__));
  not1  g0798(.din(n5557_o2), .dout(new_new_n3497__));
  buf1  g0799(.din(n5558_o2), .dout(new_new_n3498__));
  buf1  g0800(.din(n5559_o2), .dout(new_new_n3500__));
  not1  g0801(.din(n5559_o2), .dout(new_new_n3501__));
  buf1  g0802(.din(n5564_o2), .dout(new_new_n3502__));
  not1  g0803(.din(n5565_o2), .dout(new_new_n3505__));
  buf1  g0804(.din(n1966_inv), .dout(new_new_n3506__));
  buf1  g0805(.din(n5568_o2), .dout(new_new_n3508__));
  not1  g0806(.din(n5568_o2), .dout(new_new_n3509__));
  buf1  g0807(.din(n5598_o2), .dout(new_new_n3510__));
  not1  g0808(.din(n5598_o2), .dout(new_new_n3511__));
  buf1  g0809(.din(n5600_o2), .dout(new_new_n3512__));
  not1  g0810(.din(n5600_o2), .dout(new_new_n3513__));
  buf1  g0811(.din(n5601_o2), .dout(new_new_n3514__));
  buf1  g0812(.din(n5602_o2), .dout(new_new_n3516__));
  not1  g0813(.din(n5602_o2), .dout(new_new_n3517__));
  buf1  g0814(.din(n5603_o2), .dout(new_new_n3518__));
  not1  g0815(.din(n5603_o2), .dout(new_new_n3519__));
  buf1  g0816(.din(n2853_o2), .dout(new_new_n3520__));
  not1  g0817(.din(n2853_o2), .dout(new_new_n3521__));
  buf1  g0818(.din(n5637_o2), .dout(new_new_n3522__));
  not1  g0819(.din(n5637_o2), .dout(new_new_n3523__));
  buf1  g0820(.din(n1993_inv), .dout(new_new_n3524__));
  buf1  g0821(.din(n1996_inv), .dout(new_new_n3526__));
  buf1  g0822(.din(n5635_o2), .dout(new_new_n3528__));
  not1  g0823(.din(n5635_o2), .dout(new_new_n3529__));
  buf1  g0824(.din(n5640_o2), .dout(new_new_n3530__));
  not1  g0825(.din(n5640_o2), .dout(new_new_n3531__));
  buf1  g0826(.din(n5641_o2), .dout(new_new_n3532__));
  not1  g0827(.din(n5641_o2), .dout(new_new_n3533__));
  buf1  g0828(.din(n5642_o2), .dout(new_new_n3534__));
  buf1  g0829(.din(n5650_o2), .dout(new_new_n3536__));
  not1  g0830(.din(n5650_o2), .dout(new_new_n3537__));
  buf1  g0831(.din(n5652_o2), .dout(new_new_n3538__));
  buf1  g0832(.din(n5653_o2), .dout(new_new_n3540__));
  not1  g0833(.din(n5653_o2), .dout(new_new_n3541__));
  buf1  g0834(.din(n5654_o2), .dout(new_new_n3542__));
  buf1  g0835(.din(n5655_o2), .dout(new_new_n3544__));
  not1  g0836(.din(n5655_o2), .dout(new_new_n3545__));
  buf1  g0837(.din(n5657_o2), .dout(new_new_n3546__));
  buf1  g0838(.din(n2029_inv), .dout(new_new_n3548__));
  not1  g0839(.din(n5661_o2), .dout(new_new_n3551__));
  buf1  g0840(.din(n5656_o2), .dout(new_new_n3552__));
  not1  g0841(.din(n5656_o2), .dout(new_new_n3553__));
  buf1  g0842(.din(n5663_o2), .dout(new_new_n3554__));
  not1  g0843(.din(n5663_o2), .dout(new_new_n3555__));
  buf1  g0844(.din(n2041_inv), .dout(new_new_n3556__));
  buf1  g0845(.din(n5795_o2), .dout(new_new_n3558__));
  not1  g0846(.din(n5795_o2), .dout(new_new_n3559__));
  buf1  g0847(.din(n5796_o2), .dout(new_new_n3560__));
  not1  g0848(.din(n5796_o2), .dout(new_new_n3561__));
  buf1  g0849(.din(n5797_o2), .dout(new_new_n3562__));
  not1  g0850(.din(n5797_o2), .dout(new_new_n3563__));
  buf1  g0851(.din(n5739_o2), .dout(new_new_n3564__));
  not1  g0852(.din(n5739_o2), .dout(new_new_n3565__));
  buf1  g0853(.din(n5773_o2), .dout(new_new_n3566__));
  buf1  g0854(.din(n2059_inv), .dout(new_new_n3568__));
  buf1  g0855(.din(n5799_o2), .dout(new_new_n3570__));
  not1  g0856(.din(n5799_o2), .dout(new_new_n3571__));
  buf1  g0857(.din(n5802_o2), .dout(new_new_n3572__));
  buf1  g0858(.din(n2068_inv), .dout(new_new_n3574__));
  buf1  g0859(.din(n5831_o2), .dout(new_new_n3576__));
  not1  g0860(.din(n5831_o2), .dout(new_new_n3577__));
  buf1  g0861(.din(n5833_o2), .dout(new_new_n3578__));
  not1  g0862(.din(n5833_o2), .dout(new_new_n3579__));
  buf1  g0863(.din(n5820_o2), .dout(new_new_n3580__));
  buf1  g0864(.din(n5823_o2), .dout(new_new_n3582__));
  not1  g0865(.din(n5823_o2), .dout(new_new_n3583__));
  not1  g0866(.din(n5824_o2), .dout(new_new_n3585__));
  buf1  g0867(.din(n5869_o2), .dout(new_new_n3586__));
  buf1  g0868(.din(n5848_o2), .dout(new_new_n3588__));
  not1  g0869(.din(n5848_o2), .dout(new_new_n3589__));
  buf1  g0870(.din(n5849_o2), .dout(new_new_n3590__));
  not1  g0871(.din(n5849_o2), .dout(new_new_n3591__));
  buf1  g0872(.din(n5856_o2), .dout(new_new_n3592__));
  buf1  g0873(.din(n5896_o2), .dout(new_new_n3594__));
  not1  g0874(.din(n5896_o2), .dout(new_new_n3595__));
  buf1  g0875(.din(n2754_o2), .dout(new_new_n3596__));
  buf1  g0876(.din(n2908_o2), .dout(new_new_n3598__));
  buf1  g0877(.din(n5892_o2), .dout(new_new_n3600__));
  buf1  g0878(.din(n5915_o2), .dout(new_new_n3602__));
  buf1  g0879(.din(n5919_o2), .dout(new_new_n3604__));
  buf1  g0880(.din(n5918_o2), .dout(new_new_n3606__));
  not1  g0881(.din(n5918_o2), .dout(new_new_n3607__));
  buf1  g0882(.din(n5920_o2), .dout(new_new_n3608__));
  not1  g0883(.din(n5920_o2), .dout(new_new_n3609__));
  buf1  g0884(.din(n5917_o2), .dout(new_new_n3610__));
  buf1  g0885(.din(lo586_buf_o2), .dout(new_new_n3612__));
  not1  g0886(.din(lo586_buf_o2), .dout(new_new_n3613__));
  buf1  g0887(.din(n2818_o2), .dout(new_new_n3614__));
  buf1  g0888(.din(n2863_o2), .dout(new_new_n3616__));
  buf1  g0889(.din(n2134_inv), .dout(new_new_n3618__));
  not1  g0890(.din(n2134_inv), .dout(new_new_n3619__));
  buf1  g0891(.din(n2725_o2), .dout(new_new_n3620__));
  not1  g0892(.din(n2725_o2), .dout(new_new_n3621__));
  buf1  g0893(.din(n3016_o2), .dout(new_new_n3622__));
  not1  g0894(.din(n3016_o2), .dout(new_new_n3623__));
  buf1  g0895(.din(n3013_o2), .dout(new_new_n3624__));
  not1  g0896(.din(n3013_o2), .dout(new_new_n3625__));
  buf1  g0897(.din(n2655_o2), .dout(new_new_n3626__));
  not1  g0898(.din(n2655_o2), .dout(new_new_n3627__));
  buf1  g0899(.din(n2149_inv), .dout(new_new_n3628__));
  not1  g0900(.din(n2149_inv), .dout(new_new_n3629__));
  buf1  g0901(.din(lo562_buf_o2), .dout(new_new_n3630__));
  not1  g0902(.din(lo562_buf_o2), .dout(new_new_n3631__));
  buf1  g0903(.din(n2155_inv), .dout(new_new_n3632__));
  buf1  g0904(.din(n2531_o2), .dout(new_new_n3634__));
  buf1  g0905(.din(n2700_o2), .dout(new_new_n3636__));
  not1  g0906(.din(n2700_o2), .dout(new_new_n3637__));
  buf1  g0907(.din(n5908_o2), .dout(new_new_n3638__));
  not1  g0908(.din(n5908_o2), .dout(new_new_n3639__));
  buf1  g0909(.din(n5910_o2), .dout(new_new_n3640__));
  not1  g0910(.din(n5910_o2), .dout(new_new_n3641__));
  buf1  g0911(.din(n5912_o2), .dout(new_new_n3642__));
  not1  g0912(.din(n5912_o2), .dout(new_new_n3643__));
  buf1  g0913(.din(n5914_o2), .dout(new_new_n3644__));
  not1  g0914(.din(n5914_o2), .dout(new_new_n3645__));
  buf1  g0915(.din(n2753_o2), .dout(new_new_n3646__));
  not1  g0916(.din(n2753_o2), .dout(new_new_n3647__));
  buf1  g0917(.din(n2878_o2), .dout(new_new_n3648__));
  not1  g0918(.din(n2878_o2), .dout(new_new_n3649__));
  buf1  g0919(.din(n2182_inv), .dout(new_new_n3650__));
  buf1  g0920(.din(n5934_o2), .dout(new_new_n3652__));
  not1  g0921(.din(n5934_o2), .dout(new_new_n3653__));
  buf1  g0922(.din(n5936_o2), .dout(new_new_n3654__));
  not1  g0923(.din(n5936_o2), .dout(new_new_n3655__));
  buf1  g0924(.din(n5938_o2), .dout(new_new_n3656__));
  not1  g0925(.din(n5938_o2), .dout(new_new_n3657__));
  buf1  g0926(.din(n2728_o2), .dout(new_new_n3658__));
  buf1  g0927(.din(lo358_buf_o2), .dout(new_new_n3660__));
  not1  g0928(.din(lo358_buf_o2), .dout(new_new_n3661__));
  buf1  g0929(.din(lo418_buf_o2), .dout(new_new_n3662__));
  not1  g0930(.din(lo418_buf_o2), .dout(new_new_n3663__));
  buf1  g0931(.din(lo474_buf_o2), .dout(new_new_n3664__));
  not1  g0932(.din(lo474_buf_o2), .dout(new_new_n3665__));
  buf1  g0933(.din(lo554_buf_o2), .dout(new_new_n3666__));
  not1  g0934(.din(lo554_buf_o2), .dout(new_new_n3667__));
  buf1  g0935(.din(lo558_buf_o2), .dout(new_new_n3668__));
  not1  g0936(.din(lo558_buf_o2), .dout(new_new_n3669__));
  buf1  g0937(.din(lo574_buf_o2), .dout(new_new_n3670__));
  not1  g0938(.din(lo574_buf_o2), .dout(new_new_n3671__));
  buf1  g0939(.din(n2215_inv), .dout(new_new_n3672__));
  buf1  g0940(.din(n2218_inv), .dout(new_new_n3674__));
  buf1  g0941(.din(n2221_inv), .dout(new_new_n3676__));
  buf1  g0942(.din(lo450_buf_o2), .dout(new_new_n3678__));
  not1  g0943(.din(lo450_buf_o2), .dout(new_new_n3679__));
  buf1  g0944(.din(n2910_o2), .dout(new_new_n3680__));
  buf1  g0945(.din(n2683_o2), .dout(new_new_n3682__));
  not1  g0946(.din(n2683_o2), .dout(new_new_n3683__));
  not1  g0947(.din(n2828_o2), .dout(new_new_n3685__));
  buf1  g0948(.din(n2582_o2), .dout(new_new_n3686__));
  buf1  g0949(.din(n2600_o2), .dout(new_new_n3688__));
  buf1  g0950(.din(n2542_o2), .dout(new_new_n3690__));
  buf1  g0951(.din(n2703_o2), .dout(new_new_n3692__));
  buf1  g0952(.din(lo510_buf_o2), .dout(new_new_n3694__));
  not1  g0953(.din(lo510_buf_o2), .dout(new_new_n3695__));
  buf1  g0954(.din(lo514_buf_o2), .dout(new_new_n3696__));
  buf1  g0955(.din(lo538_buf_o2), .dout(new_new_n3698__));
  not1  g0956(.din(lo538_buf_o2), .dout(new_new_n3699__));
  buf1  g0957(.din(lo578_buf_o2), .dout(new_new_n3700__));
  not1  g0958(.din(lo578_buf_o2), .dout(new_new_n3701__));
  buf1  g0959(.din(n2260_inv), .dout(new_new_n3702__));
  buf1  g0960(.din(n2666_o2), .dout(new_new_n3704__));
  buf1  g0961(.din(n2667_o2), .dout(new_new_n3706__));
  buf1  g0962(.din(n2660_o2), .dout(new_new_n3708__));
  not1  g0963(.din(n2660_o2), .dout(new_new_n3709__));
  buf1  g0964(.din(n2272_inv), .dout(new_new_n3710__));
  buf1  g0965(.din(lo454_buf_o2), .dout(new_new_n3712__));
  buf1  g0966(.din(n3593_o2), .dout(new_new_n3714__));
  not1  g0967(.din(n3593_o2), .dout(new_new_n3715__));
  buf1  g0968(.din(n3048_o2), .dout(new_new_n3716__));
  not1  g0969(.din(n3048_o2), .dout(new_new_n3717__));
  buf1  g0970(.din(lo410_buf_o2), .dout(new_new_n3718__));
  not1  g0971(.din(lo410_buf_o2), .dout(new_new_n3719__));
  buf1  g0972(.din(lo502_buf_o2), .dout(new_new_n3720__));
  not1  g0973(.din(lo502_buf_o2), .dout(new_new_n3721__));
  buf1  g0974(.din(lo506_buf_o2), .dout(new_new_n3722__));
  buf1  g0975(.din(lo550_buf_o2), .dout(new_new_n3724__));
  not1  g0976(.din(lo550_buf_o2), .dout(new_new_n3725__));
  buf1  g0977(.din(lo570_buf_o2), .dout(new_new_n3726__));
  not1  g0978(.din(lo570_buf_o2), .dout(new_new_n3727__));
  buf1  g0979(.din(lo582_buf_o2), .dout(new_new_n3728__));
  not1  g0980(.din(lo582_buf_o2), .dout(new_new_n3729__));
  buf1  g0981(.din(n2302_inv), .dout(new_new_n3730__));
  buf1  g0982(.din(n2305_inv), .dout(new_new_n3732__));
  buf1  g0983(.din(n3499_o2), .dout(new_new_n3734__));
  not1  g0984(.din(n3499_o2), .dout(new_new_n3735__));
  buf1  g0985(.din(n2311_inv), .dout(new_new_n3736__));
  buf1  g0986(.din(n2870_o2), .dout(new_new_n3738__));
  buf1  g0987(.din(n2317_inv), .dout(new_new_n3740__));
  not1  g0988(.din(n2317_inv), .dout(new_new_n3741__));
  buf1  g0989(.din(n2689_o2), .dout(new_new_n3742__));
  not1  g0990(.din(n2689_o2), .dout(new_new_n3743__));
  buf1  g0991(.din(n2323_inv), .dout(new_new_n3744__));
  not1  g0992(.din(n2323_inv), .dout(new_new_n3745__));
  buf1  g0993(.din(n2662_o2), .dout(new_new_n3746__));
  not1  g0994(.din(n2662_o2), .dout(new_new_n3747__));
  buf1  g0995(.din(lo350_buf_o2), .dout(new_new_n3748__));
  not1  g0996(.din(lo350_buf_o2), .dout(new_new_n3749__));
  buf1  g0997(.din(lo498_buf_o2), .dout(new_new_n3750__));
  buf1  g0998(.din(lo518_buf_o2), .dout(new_new_n3752__));
  not1  g0999(.din(lo518_buf_o2), .dout(new_new_n3753__));
  buf1  g1000(.din(lo522_buf_o2), .dout(new_new_n3754__));
  buf1  g1001(.din(lo598_buf_o2), .dout(new_new_n3756__));
  not1  g1002(.din(lo598_buf_o2), .dout(new_new_n3757__));
  buf1  g1003(.din(n2344_inv), .dout(new_new_n3758__));
  buf1  g1004(.din(n2347_inv), .dout(new_new_n3760__));
  buf1  g1005(.din(n2350_inv), .dout(new_new_n3762__));
  buf1  g1006(.din(n2353_inv), .dout(new_new_n3764__));
  not1  g1007(.din(n2353_inv), .dout(new_new_n3765__));
  buf1  g1008(.din(n2356_inv), .dout(new_new_n3766__));
  buf1  g1009(.din(n2359_inv), .dout(new_new_n3768__));
  buf1  g1010(.din(n2872_o2), .dout(new_new_n3770__));
  buf1  g1011(.din(n3313_o2), .dout(new_new_n3772__));
  buf1  g1012(.din(n3273_o2), .dout(new_new_n3774__));
  buf1  g1013(.din(n2848_o2), .dout(new_new_n3776__));
  buf1  g1014(.din(n2893_o2), .dout(new_new_n3778__));
  buf1  g1015(.din(n3267_o2), .dout(new_new_n3780__));
  buf1  g1016(.din(n2925_o2), .dout(new_new_n3782__));
  not1  g1017(.din(n2839_o2), .dout(new_new_n3785__));
  buf1  g1018(.din(n2831_o2), .dout(new_new_n3786__));
  buf1  g1019(.din(n2558_o2), .dout(new_new_n3788__));
  buf1  g1020(.din(n2562_o2), .dout(new_new_n3790__));
  buf1  g1021(.din(n2825_o2), .dout(new_new_n3792__));
  not1  g1022(.din(n2825_o2), .dout(new_new_n3793__));
  buf1  g1023(.din(n3263_o2), .dout(new_new_n3794__));
  buf1  g1024(.din(n3517_o2), .dout(new_new_n3796__));
  buf1  g1025(.din(n2873_o2), .dout(new_new_n3798__));
  buf1  g1026(.din(n2926_o2), .dout(new_new_n3800__));
  not1  g1027(.din(n3261_o2), .dout(new_new_n3803__));
  buf1  g1028(.din(n3268_o2), .dout(new_new_n3804__));
  buf1  g1029(.din(n3274_o2), .dout(new_new_n3806__));
  buf1  g1030(.din(n3314_o2), .dout(new_new_n3808__));
  not1  g1031(.din(n3571_o2), .dout(new_new_n3811__));
  buf1  g1032(.din(n2950_o2), .dout(new_new_n3812__));
  not1  g1033(.din(n2950_o2), .dout(new_new_n3813__));
  buf1  g1034(.din(n2951_o2), .dout(new_new_n3814__));
  not1  g1035(.din(n2951_o2), .dout(new_new_n3815__));
  buf1  g1036(.din(n3022_o2), .dout(new_new_n3816__));
  buf1  g1037(.din(n3023_o2), .dout(new_new_n3818__));
  not1  g1038(.din(n3057_o2), .dout(new_new_n3821__));
  buf1  g1039(.din(n3058_o2), .dout(new_new_n3822__));
  not1  g1040(.din(n2931_o2), .dout(new_new_n3825__));
  buf1  g1041(.din(n2911_o2), .dout(new_new_n3826__));
  not1  g1042(.din(n2911_o2), .dout(new_new_n3827__));
  buf1  g1043(.din(n2959_o2), .dout(new_new_n3828__));
  not1  g1044(.din(n2959_o2), .dout(new_new_n3829__));
  buf1  g1045(.din(n2960_o2), .dout(new_new_n3830__));
  not1  g1046(.din(n2960_o2), .dout(new_new_n3831__));
  not1  g1047(.din(n2922_o2), .dout(new_new_n3833__));
  buf1  g1048(.din(n2888_o2), .dout(new_new_n3834__));
  not1  g1049(.din(n2889_o2), .dout(new_new_n3837__));
  buf1  g1050(.din(n3051_o2), .dout(new_new_n3838__));
  not1  g1051(.din(n3052_o2), .dout(new_new_n3841__));
  not1  g1052(.din(n3063_o2), .dout(new_new_n3843__));
  buf1  g1053(.din(n2845_o2), .dout(new_new_n3844__));
  buf1  g1054(.din(n2476_inv), .dout(new_new_n3846__));
  buf1  g1055(.din(n3281_o2), .dout(new_new_n3848__));
  buf1  g1056(.din(n3294_o2), .dout(new_new_n3850__));
  buf1  g1057(.din(n2885_o2), .dout(new_new_n3852__));
  buf1  g1058(.din(n2786_o2), .dout(new_new_n3854__));
  not1  g1059(.din(n2786_o2), .dout(new_new_n3855__));
  buf1  g1060(.din(n2783_o2), .dout(new_new_n3856__));
  not1  g1061(.din(n2783_o2), .dout(new_new_n3857__));
  buf1  g1062(.din(n2801_o2), .dout(new_new_n3858__));
  not1  g1063(.din(n2801_o2), .dout(new_new_n3859__));
  buf1  g1064(.din(n2572_o2), .dout(new_new_n3860__));
  not1  g1065(.din(n2572_o2), .dout(new_new_n3861__));
  buf1  g1066(.din(n2628_o2), .dout(new_new_n3862__));
  not1  g1067(.din(n2628_o2), .dout(new_new_n3863__));
  buf1  g1068(.din(n2609_o2), .dout(new_new_n3864__));
  not1  g1069(.din(n2609_o2), .dout(new_new_n3865__));
  buf1  g1070(.din(n2618_o2), .dout(new_new_n3866__));
  not1  g1071(.din(n2618_o2), .dout(new_new_n3867__));
  buf1  g1072(.din(n2637_o2), .dout(new_new_n3868__));
  not1  g1073(.din(n2637_o2), .dout(new_new_n3869__));
  buf1  g1074(.din(n2525_o2), .dout(new_new_n3870__));
  not1  g1075(.din(n2525_o2), .dout(new_new_n3871__));
  buf1  g1076(.din(n2551_o2), .dout(new_new_n3872__));
  buf1  g1077(.din(n3759_o2), .dout(new_new_n3874__));
  buf1  g1078(.din(n2994_o2), .dout(new_new_n3876__));
  not1  g1079(.din(n2994_o2), .dout(new_new_n3877__));
  buf1  g1080(.din(n3040_o2), .dout(new_new_n3878__));
  not1  g1081(.din(n3040_o2), .dout(new_new_n3879__));
  buf1  g1082(.din(n2943_o2), .dout(new_new_n3880__));
  not1  g1083(.din(n2943_o2), .dout(new_new_n3881__));
  buf1  g1084(.din(n2991_o2), .dout(new_new_n3882__));
  not1  g1085(.din(n2991_o2), .dout(new_new_n3883__));
  buf1  g1086(.din(n3034_o2), .dout(new_new_n3884__));
  not1  g1087(.din(n3034_o2), .dout(new_new_n3885__));
  not1  g1088(.din(n2881_o2), .dout(new_new_n3887__));
  not1  g1089(.din(n3021_o2), .dout(new_new_n3889__));
  buf1  g1090(.din(n3062_o2), .dout(new_new_n3890__));
  buf1  g1091(.din(n2763_o2), .dout(new_new_n3892__));
  not1  g1092(.din(n2763_o2), .dout(new_new_n3893__));
  buf1  g1093(.din(n2764_o2), .dout(new_new_n3894__));
  not1  g1094(.din(n2764_o2), .dout(new_new_n3895__));
  buf1  g1095(.din(n2775_o2), .dout(new_new_n3896__));
  not1  g1096(.din(n2775_o2), .dout(new_new_n3897__));
  buf1  g1097(.din(n2776_o2), .dout(new_new_n3898__));
  not1  g1098(.din(n2776_o2), .dout(new_new_n3899__));
  buf1  g1099(.din(n2968_o2), .dout(new_new_n3900__));
  not1  g1100(.din(n2968_o2), .dout(new_new_n3901__));
  buf1  g1101(.din(n2969_o2), .dout(new_new_n3902__));
  not1  g1102(.din(n2969_o2), .dout(new_new_n3903__));
  buf1  g1103(.din(n2798_o2), .dout(new_new_n3904__));
  not1  g1104(.din(n2798_o2), .dout(new_new_n3905__));
  not1  g1105(.din(n3661_o2), .dout(new_new_n3907__));
  buf1  g1106(.din(n2694_o2), .dout(new_new_n3908__));
  not1  g1107(.din(n2694_o2), .dout(new_new_n3909__));
  buf1  g1108(.din(n2572_inv), .dout(new_new_n3910__));
  not1  g1109(.din(n2572_inv), .dout(new_new_n3911__));
  buf1  g1110(.din(n2817_o2), .dout(new_new_n3912__));
  not1  g1111(.din(n2817_o2), .dout(new_new_n3913__));
  not1  g1112(.din(n2514_o2), .dout(new_new_n3915__));
  not1  g1113(.din(n2501_o2), .dout(new_new_n3917__));
  buf1  g1114(.din(n2584_inv), .dout(new_new_n3918__));
  buf1  g1115(.din(n2505_o2), .dout(new_new_n3920__));
  buf1  g1116(.din(n2492_o2), .dout(new_new_n3922__));
  not1  g1117(.din(n2492_o2), .dout(new_new_n3923__));
  buf1  g1118(.din(lo546_buf_o2), .dout(new_new_n3924__));
  not1  g1119(.din(lo546_buf_o2), .dout(new_new_n3925__));
  buf1  g1120(.din(lo590_buf_o2), .dout(new_new_n3926__));
  not1  g1121(.din(lo590_buf_o2), .dout(new_new_n3927__));
  buf1  g1122(.din(lo594_buf_o2), .dout(new_new_n3928__));
  not1  g1123(.din(lo594_buf_o2), .dout(new_new_n3929__));
  buf1  g1124(.din(n2602_inv), .dout(new_new_n3930__));
  buf1  g1125(.din(n2605_inv), .dout(new_new_n3932__));
  buf1  g1126(.din(n2709_o2), .dout(new_new_n3934__));
  not1  g1127(.din(n2709_o2), .dout(new_new_n3935__));
  buf1  g1128(.din(n2611_inv), .dout(new_new_n3936__));
  not1  g1129(.din(n2611_inv), .dout(new_new_n3937__));
  buf1  g1130(.din(n2614_inv), .dout(new_new_n3938__));
  not1  g1131(.din(n2614_inv), .dout(new_new_n3939__));
  buf1  g1132(.din(n2617_inv), .dout(new_new_n3940__));
  not1  g1133(.din(n2617_inv), .dout(new_new_n3941__));
  buf1  g1134(.din(n2620_inv), .dout(new_new_n3942__));
  not1  g1135(.din(n2620_inv), .dout(new_new_n3943__));
  buf1  g1136(.din(n3590_o2), .dout(new_new_n3944__));
  not1  g1137(.din(n3590_o2), .dout(new_new_n3945__));
  buf1  g1138(.din(n3591_o2), .dout(new_new_n3946__));
  not1  g1139(.din(n3591_o2), .dout(new_new_n3947__));
  buf1  g1140(.din(n2629_inv), .dout(new_new_n3948__));
  not1  g1141(.din(n2629_inv), .dout(new_new_n3949__));
  buf1  g1142(.din(n3638_o2), .dout(new_new_n3950__));
  not1  g1143(.din(n3638_o2), .dout(new_new_n3951__));
  buf1  g1144(.din(n3639_o2), .dout(new_new_n3952__));
  not1  g1145(.din(n3639_o2), .dout(new_new_n3953__));
  buf1  g1146(.din(n2638_inv), .dout(new_new_n3954__));
  not1  g1147(.din(n2638_inv), .dout(new_new_n3955__));
  buf1  g1148(.din(n2641_inv), .dout(new_new_n3956__));
  not1  g1149(.din(n2641_inv), .dout(new_new_n3957__));
  buf1  g1150(.din(lo458_buf_o2), .dout(new_new_n3958__));
  not1  g1151(.din(lo458_buf_o2), .dout(new_new_n3959__));
  buf1  g1152(.din(lo482_buf_o2), .dout(new_new_n3960__));
  not1  g1153(.din(lo482_buf_o2), .dout(new_new_n3961__));
  buf1  g1154(.din(lo566_buf_o2), .dout(new_new_n3962__));
  not1  g1155(.din(lo566_buf_o2), .dout(new_new_n3963__));
  buf1  g1156(.din(n2718_o2), .dout(new_new_n3964__));
  not1  g1157(.din(n2718_o2), .dout(new_new_n3965__));
  buf1  g1158(.din(n3707_o2), .dout(new_new_n3966__));
  not1  g1159(.din(n3707_o2), .dout(new_new_n3967__));
  buf1  g1160(.din(n3671_o2), .dout(new_new_n3968__));
  not1  g1161(.din(n3671_o2), .dout(new_new_n3969__));
  buf1  g1162(.din(n3680_o2), .dout(new_new_n3970__));
  not1  g1163(.din(n3680_o2), .dout(new_new_n3971__));
  buf1  g1164(.din(n3749_o2), .dout(new_new_n3972__));
  not1  g1165(.din(n3749_o2), .dout(new_new_n3973__));
  buf1  g1166(.din(n3716_o2), .dout(new_new_n3974__));
  not1  g1167(.din(n3716_o2), .dout(new_new_n3975__));
  buf1  g1168(.din(n3692_o2), .dout(new_new_n3976__));
  not1  g1169(.din(n3692_o2), .dout(new_new_n3977__));
  buf1  g1170(.din(n2591_o2), .dout(new_new_n3978__));
  not1  g1171(.din(n2591_o2), .dout(new_new_n3979__));
  buf1  g1172(.din(n3478_o2), .dout(new_new_n3980__));
  not1  g1173(.din(n3478_o2), .dout(new_new_n3981__));
  buf1  g1174(.din(n3610_o2), .dout(new_new_n3982__));
  not1  g1175(.din(n3610_o2), .dout(new_new_n3983__));
  buf1  g1176(.din(n3611_o2), .dout(new_new_n3984__));
  not1  g1177(.din(n3611_o2), .dout(new_new_n3985__));
  buf1  g1178(.din(n2686_inv), .dout(new_new_n3986__));
  buf1  g1179(.din(n2689_inv), .dout(new_new_n3988__));
  not1  g1180(.din(n2689_inv), .dout(new_new_n3989__));
  buf1  g1181(.din(n2738_o2), .dout(new_new_n3990__));
  not1  g1182(.din(n2738_o2), .dout(new_new_n3991__));
  buf1  g1183(.din(n3616_o2), .dout(new_new_n3992__));
  not1  g1184(.din(n3616_o2), .dout(new_new_n3993__));
  buf1  g1185(.din(n3617_o2), .dout(new_new_n3994__));
  not1  g1186(.din(n3617_o2), .dout(new_new_n3995__));
  buf1  g1187(.din(n3031_o2), .dout(new_new_n3996__));
  buf1  g1188(.din(n2704_inv), .dout(new_new_n3998__));
  not1  g1189(.din(n2704_inv), .dout(new_new_n3999__));
  buf1  g1190(.din(n3562_o2), .dout(new_new_n4000__));
  not1  g1191(.din(n3562_o2), .dout(new_new_n4001__));
  buf1  g1192(.din(n2502_o2), .dout(new_new_n4002__));
  not1  g1193(.din(n2502_o2), .dout(new_new_n4003__));
  buf1  g1194(.din(n3560_o2), .dout(new_new_n4004__));
  not1  g1195(.din(n3560_o2), .dout(new_new_n4005__));
  buf1  g1196(.din(n3554_o2), .dout(new_new_n4006__));
  not1  g1197(.din(n3554_o2), .dout(new_new_n4007__));
  buf1  g1198(.din(n3555_o2), .dout(new_new_n4008__));
  not1  g1199(.din(n3555_o2), .dout(new_new_n4009__));
  buf1  g1200(.din(n3536_o2), .dout(new_new_n4010__));
  not1  g1201(.din(n3536_o2), .dout(new_new_n4011__));
  buf1  g1202(.din(n3537_o2), .dout(new_new_n4012__));
  not1  g1203(.din(n3537_o2), .dout(new_new_n4013__));
  buf1  g1204(.din(n3508_o2), .dout(new_new_n4014__));
  not1  g1205(.din(n3508_o2), .dout(new_new_n4015__));
  buf1  g1206(.din(n3650_o2), .dout(new_new_n4016__));
  not1  g1207(.din(n3650_o2), .dout(new_new_n4017__));
  buf1  g1208(.din(n3740_o2), .dout(new_new_n4018__));
  not1  g1209(.din(n3740_o2), .dout(new_new_n4019__));
  buf1  g1210(.din(n3484_o2), .dout(new_new_n4020__));
  not1  g1211(.din(n3484_o2), .dout(new_new_n4021__));
  buf1  g1212(.din(n2740_inv), .dout(new_new_n4022__));
  not1  g1213(.din(n2740_inv), .dout(new_new_n4023__));
  buf1  g1214(.din(n2734_o2), .dout(new_new_n4024__));
  not1  g1215(.din(n2734_o2), .dout(new_new_n4025__));
  buf1  g1216(.din(n2735_o2), .dout(new_new_n4026__));
  not1  g1217(.din(n2735_o2), .dout(new_new_n4027__));
  buf1  g1218(.din(n2711_o2), .dout(new_new_n4028__));
  not1  g1219(.din(n2711_o2), .dout(new_new_n4029__));
  buf1  g1220(.din(lo585_buf_o2), .dout(new_new_n4030__));
  not1  g1221(.din(lo585_buf_o2), .dout(new_new_n4031__));
  buf1  g1222(.din(n2719_o2), .dout(new_new_n4032__));
  not1  g1223(.din(n2719_o2), .dout(new_new_n4033__));
  buf1  g1224(.din(n2720_o2), .dout(new_new_n4034__));
  not1  g1225(.din(n2720_o2), .dout(new_new_n4035__));
  buf1  g1226(.din(n2723_o2), .dout(new_new_n4036__));
  not1  g1227(.din(n2723_o2), .dout(new_new_n4037__));
  buf1  g1228(.din(n2724_o2), .dout(new_new_n4038__));
  not1  g1229(.din(n2724_o2), .dout(new_new_n4039__));
  buf1  g1230(.din(n3624_o2), .dout(new_new_n4040__));
  not1  g1231(.din(n3624_o2), .dout(new_new_n4041__));
  buf1  g1232(.din(n3625_o2), .dout(new_new_n4042__));
  not1  g1233(.din(n3625_o2), .dout(new_new_n4043__));
  buf1  g1234(.din(n3015_o2), .dout(new_new_n4044__));
  not1  g1235(.din(n3015_o2), .dout(new_new_n4045__));
  buf1  g1236(.din(n3491_o2), .dout(new_new_n4046__));
  not1  g1237(.din(n3491_o2), .dout(new_new_n4047__));
  buf1  g1238(.din(n2779_inv), .dout(new_new_n4048__));
  not1  g1239(.din(n2779_inv), .dout(new_new_n4049__));
  buf1  g1240(.din(n2811_o2), .dout(new_new_n4050__));
  not1  g1241(.din(n2811_o2), .dout(new_new_n4051__));
  buf1  g1242(.din(n3010_o2), .dout(new_new_n4052__));
  not1  g1243(.din(n3010_o2), .dout(new_new_n4053__));
  buf1  g1244(.din(n3012_o2), .dout(new_new_n4054__));
  not1  g1245(.din(n3012_o2), .dout(new_new_n4055__));
  buf1  g1246(.din(lo382_buf_o2), .dout(new_new_n4056__));
  not1  g1247(.din(lo382_buf_o2), .dout(new_new_n4057__));
  buf1  g1248(.din(lo386_buf_o2), .dout(new_new_n4058__));
  not1  g1249(.din(lo386_buf_o2), .dout(new_new_n4059__));
  buf1  g1250(.din(lo390_buf_o2), .dout(new_new_n4060__));
  not1  g1251(.din(lo390_buf_o2), .dout(new_new_n4061__));
  buf1  g1252(.din(lo398_buf_o2), .dout(new_new_n4062__));
  not1  g1253(.din(lo398_buf_o2), .dout(new_new_n4063__));
  buf1  g1254(.din(lo402_buf_o2), .dout(new_new_n4064__));
  not1  g1255(.din(lo402_buf_o2), .dout(new_new_n4065__));
  buf1  g1256(.din(lo406_buf_o2), .dout(new_new_n4066__));
  not1  g1257(.din(lo406_buf_o2), .dout(new_new_n4067__));
  buf1  g1258(.din(n3492_o2), .dout(new_new_n4068__));
  not1  g1259(.din(n3492_o2), .dout(new_new_n4069__));
  buf1  g1260(.din(lo366_buf_o2), .dout(new_new_n4070__));
  buf1  g1261(.din(lo374_buf_o2), .dout(new_new_n4072__));
  buf1  g1262(.din(lo426_buf_o2), .dout(new_new_n4074__));
  buf1  g1263(.din(lo494_buf_o2), .dout(new_new_n4076__));
  not1  g1264(.din(lo494_buf_o2), .dout(new_new_n4077__));
  buf1  g1265(.din(n2653_o2), .dout(new_new_n4078__));
  not1  g1266(.din(n2653_o2), .dout(new_new_n4079__));
  buf1  g1267(.din(n2654_o2), .dout(new_new_n4080__));
  not1  g1268(.din(n2654_o2), .dout(new_new_n4081__));
  buf1  g1269(.din(n2715_o2), .dout(new_new_n4082__));
  not1  g1270(.din(n2715_o2), .dout(new_new_n4083__));
  buf1  g1271(.din(n2740_o2), .dout(new_new_n4084__));
  not1  g1272(.din(n2740_o2), .dout(new_new_n4085__));
  buf1  g1273(.din(n2682_o2), .dout(new_new_n4086__));
  not1  g1274(.din(n2682_o2), .dout(new_new_n4087__));
  buf1  g1275(.din(n2736_o2), .dout(new_new_n4088__));
  not1  g1276(.din(n2736_o2), .dout(new_new_n4089__));
  buf1  g1277(.din(lo508_buf_o2), .dout(new_new_n4090__));
  not1  g1278(.din(lo508_buf_o2), .dout(new_new_n4091__));
  buf1  g1279(.din(lo512_buf_o2), .dout(new_new_n4092__));
  not1  g1280(.din(lo512_buf_o2), .dout(new_new_n4093__));
  buf1  g1281(.din(lo536_buf_o2), .dout(new_new_n4094__));
  not1  g1282(.din(lo536_buf_o2), .dout(new_new_n4095__));
  buf1  g1283(.din(lo576_buf_o2), .dout(new_new_n4096__));
  not1  g1284(.din(lo576_buf_o2), .dout(new_new_n4097__));
  buf1  g1285(.din(lo357_buf_o2), .dout(new_new_n4098__));
  not1  g1286(.din(lo357_buf_o2), .dout(new_new_n4099__));
  buf1  g1287(.din(lo361_buf_o2), .dout(new_new_n4100__));
  not1  g1288(.din(lo361_buf_o2), .dout(new_new_n4101__));
  buf1  g1289(.din(lo417_buf_o2), .dout(new_new_n4102__));
  not1  g1290(.din(lo417_buf_o2), .dout(new_new_n4103__));
  buf1  g1291(.din(lo421_buf_o2), .dout(new_new_n4104__));
  not1  g1292(.din(lo421_buf_o2), .dout(new_new_n4105__));
  buf1  g1293(.din(lo473_buf_o2), .dout(new_new_n4106__));
  buf1  g1294(.din(lo477_buf_o2), .dout(new_new_n4108__));
  buf1  g1295(.din(lo553_buf_o2), .dout(new_new_n4110__));
  not1  g1296(.din(lo553_buf_o2), .dout(new_new_n4111__));
  buf1  g1297(.din(lo557_buf_o2), .dout(new_new_n4112__));
  not1  g1298(.din(lo557_buf_o2), .dout(new_new_n4113__));
  buf1  g1299(.din(lo573_buf_o2), .dout(new_new_n4114__));
  not1  g1300(.din(lo573_buf_o2), .dout(new_new_n4115__));
  buf1  g1301(.din(lo434_buf_o2), .dout(new_new_n4116__));
  not1  g1302(.din(lo434_buf_o2), .dout(new_new_n4117__));
  buf1  g1303(.din(lo438_buf_o2), .dout(new_new_n4118__));
  not1  g1304(.din(lo438_buf_o2), .dout(new_new_n4119__));
  buf1  g1305(.din(lo466_buf_o2), .dout(new_new_n4120__));
  not1  g1306(.din(lo466_buf_o2), .dout(new_new_n4121__));
  buf1  g1307(.din(lo470_buf_o2), .dout(new_new_n4122__));
  not1  g1308(.din(lo470_buf_o2), .dout(new_new_n4123__));
  buf1  g1309(.din(lo490_buf_o2), .dout(new_new_n4124__));
  not1  g1310(.din(lo490_buf_o2), .dout(new_new_n4125__));
  buf1  g1311(.din(n2657_o2), .dout(new_new_n4126__));
  not1  g1312(.din(n2657_o2), .dout(new_new_n4127__));
  buf1  g1313(.din(n2658_o2), .dout(new_new_n4128__));
  not1  g1314(.din(n2658_o2), .dout(new_new_n4129__));
  buf1  g1315(.din(n2663_o2), .dout(new_new_n4130__));
  not1  g1316(.din(n2663_o2), .dout(new_new_n4131__));
  buf1  g1317(.din(n2664_o2), .dout(new_new_n4132__));
  not1  g1318(.din(n2664_o2), .dout(new_new_n4133__));
  buf1  g1319(.din(n2684_o2), .dout(new_new_n4134__));
  not1  g1320(.din(n2684_o2), .dout(new_new_n4135__));
  buf1  g1321(.din(n2685_o2), .dout(new_new_n4136__));
  not1  g1322(.din(n2685_o2), .dout(new_new_n4137__));
  or1   g1323(.dina(new_new_n6741__), .dinb(new_new_n6742__), .dout(new_new_n4138__));
  and1  g1324(.dina(new_new_n6745__), .dinb(new_new_n2904__), .dout(new_new_n4139__));
  and1  g1325(.dina(new_new_n6748__), .dinb(new_new_n3162__), .dout(new_new_n4140__));
  and1  g1326(.dina(new_new_n2872__), .dinb(new_new_n6749__), .dout(new_new_n4141__));
  or1   g1327(.dina(new_new_n6750__), .dinb(new_new_n3298__), .dout(new_new_n4142__));
  or1   g1328(.dina(new_new_n3171__), .dinb(new_new_n3225__), .dout(new_new_n4143__));
  or1   g1329(.dina(new_new_n6750__), .dinb(new_new_n2491__), .dout(new_new_n4144__));
  or1   g1330(.dina(new_new_n2889__), .dinb(new_new_n6754__), .dout(new_new_n4145__));
  or1   g1331(.dina(new_new_n2663__), .dinb(new_new_n6761__), .dout(new_new_n4146__));
  or1   g1332(.dina(new_new_n2655__), .dinb(new_new_n6766__), .dout(new_new_n4147__));
  and1  g1333(.dina(new_new_n4146__), .dinb(new_new_n4147__), .dout(new_new_n4148__));
  or1   g1334(.dina(new_new_n6754__), .dinb(new_new_n4148__), .dout(new_new_n4149__));
  or1   g1335(.dina(new_new_n2499__), .dinb(new_new_n6761__), .dout(new_new_n4150__));
  or1   g1336(.dina(new_new_n2671__), .dinb(new_new_n6766__), .dout(new_new_n4151__));
  and1  g1337(.dina(new_new_n4150__), .dinb(new_new_n4151__), .dout(new_new_n4152__));
  or1   g1338(.dina(new_new_n6753__), .dinb(new_new_n4152__), .dout(new_new_n4153__));
  or1   g1339(.dina(new_new_n2647__), .dinb(new_new_n6755__), .dout(new_new_n4154__));
  and1  g1340(.dina(new_new_n2466__), .dinb(new_new_n6762__), .dout(new_new_n4155__));
  and1  g1341(.dina(new_new_n2458__), .dinb(new_new_n6767__), .dout(new_new_n4156__));
  or1   g1342(.dina(new_new_n6755__), .dinb(new_new_n4156__), .dout(new_new_n4157__));
  or1   g1343(.dina(new_new_n4155__), .dinb(new_new_n4157__), .dout(new_new_n4158__));
  and1  g1344(.dina(new_new_n6745__), .dinb(new_new_n4158__), .dout(new_new_n4159__));
  and1  g1345(.dina(new_new_n2630__), .dinb(new_new_n6762__), .dout(new_new_n4160__));
  and1  g1346(.dina(new_new_n2474__), .dinb(new_new_n6767__), .dout(new_new_n4161__));
  or1   g1347(.dina(new_new_n6757__), .dinb(new_new_n4161__), .dout(new_new_n4162__));
  or1   g1348(.dina(new_new_n4160__), .dinb(new_new_n4162__), .dout(new_new_n4163__));
  and1  g1349(.dina(new_new_n6746__), .dinb(new_new_n4163__), .dout(new_new_n4164__));
  and1  g1350(.dina(new_new_n2450__), .dinb(new_new_n6763__), .dout(new_new_n4165__));
  and1  g1351(.dina(new_new_n2614__), .dinb(new_new_n6768__), .dout(new_new_n4166__));
  or1   g1352(.dina(new_new_n6757__), .dinb(new_new_n4166__), .dout(new_new_n4167__));
  or1   g1353(.dina(new_new_n4165__), .dinb(new_new_n4167__), .dout(new_new_n4168__));
  and1  g1354(.dina(new_new_n6746__), .dinb(new_new_n4168__), .dout(new_new_n4169__));
  and1  g1355(.dina(new_new_n2622__), .dinb(new_new_n6763__), .dout(new_new_n4170__));
  and1  g1356(.dina(new_new_n2638__), .dinb(new_new_n6768__), .dout(new_new_n4171__));
  or1   g1357(.dina(new_new_n6758__), .dinb(new_new_n4171__), .dout(new_new_n4172__));
  or1   g1358(.dina(new_new_n4170__), .dinb(new_new_n4172__), .dout(new_new_n4173__));
  and1  g1359(.dina(new_new_n6747__), .dinb(new_new_n4173__), .dout(new_new_n4174__));
  and1  g1360(.dina(new_new_n3466__), .dinb(new_new_n3468__), .dout(new_new_n4175__));
  and1  g1361(.dina(new_new_n3449__), .dinb(new_new_n3634__), .dout(new_new_n4176__));
  and1  g1362(.dina(new_new_n3870__), .dinb(new_new_n4176__), .dout(new_new_n4177__));
  and1  g1363(.dina(new_new_n3690__), .dinb(new_new_n6769__), .dout(new_new_n4178__));
  and1  g1364(.dina(new_new_n4177__), .dinb(new_new_n4178__), .dout(new_new_n4179__));
  and1  g1365(.dina(new_new_n4175__), .dinb(new_new_n4179__), .dout(new_new_n4180__));
  and1  g1366(.dina(new_new_n3864__), .dinb(new_new_n3866__), .dout(new_new_n4181__));
  and1  g1367(.dina(new_new_n3862__), .dinb(new_new_n4181__), .dout(new_new_n4182__));
  or1   g1368(.dina(new_new_n3788__), .dinb(new_new_n3790__), .dout(new_new_n4183__));
  and1  g1369(.dina(new_new_n3860__), .dinb(new_new_n6770__), .dout(new_new_n4184__));
  and1  g1370(.dina(new_new_n3464__), .dinb(new_new_n3686__), .dout(new_new_n4185__));
  and1  g1371(.dina(new_new_n3688__), .dinb(new_new_n3868__), .dout(new_new_n4186__));
  and1  g1372(.dina(new_new_n4185__), .dinb(new_new_n4186__), .dout(new_new_n4187__));
  and1  g1373(.dina(new_new_n4184__), .dinb(new_new_n4187__), .dout(new_new_n4188__));
  and1  g1374(.dina(new_new_n4182__), .dinb(new_new_n4188__), .dout(new_new_n4189__));
  or1   g1375(.dina(new_new_n3419__), .dinb(new_new_n6771__), .dout(new_new_n4190__));
  or1   g1376(.dina(new_new_n3461__), .dinb(new_new_n6772__), .dout(new_new_n4191__));
  and1  g1377(.dina(new_new_n3440__), .dinb(new_new_n3489__), .dout(new_new_n4192__));
  and1  g1378(.dina(new_new_n3426__), .dinb(new_new_n4192__), .dout(new_new_n4193__));
  and1  g1379(.dina(new_new_n3434__), .dinb(new_new_n3596__), .dout(new_new_n4194__));
  and1  g1380(.dina(new_new_n4193__), .dinb(new_new_n4194__), .dout(new_new_n4195__));
  and1  g1381(.dina(new_new_n3893__), .dinb(new_new_n3895__), .dout(new_new_n4196__));
  or1   g1382(.dina(new_new_n3892__), .dinb(new_new_n3894__), .dout(new_new_n4197__));
  and1  g1383(.dina(new_new_n3897__), .dinb(new_new_n3899__), .dout(new_new_n4198__));
  or1   g1384(.dina(new_new_n3896__), .dinb(new_new_n3898__), .dout(new_new_n4199__));
  and1  g1385(.dina(new_new_n4197__), .dinb(new_new_n4198__), .dout(new_new_n4200__));
  and1  g1386(.dina(new_new_n4196__), .dinb(new_new_n4199__), .dout(new_new_n4201__));
  or1   g1387(.dina(new_new_n4200__), .dinb(new_new_n4201__), .dout(new_new_n4202__));
  and1  g1388(.dina(new_new_n6773__), .dinb(new_new_n6774__), .dout(new_new_n4203__));
  or1   g1389(.dina(new_new_n6775__), .dinb(new_new_n6776__), .dout(new_new_n4204__));
  and1  g1390(.dina(new_new_n6775__), .dinb(new_new_n6776__), .dout(new_new_n4205__));
  or1   g1391(.dina(new_new_n6773__), .dinb(new_new_n6774__), .dout(new_new_n4206__));
  and1  g1392(.dina(new_new_n4204__), .dinb(new_new_n4206__), .dout(new_new_n4207__));
  or1   g1393(.dina(new_new_n4203__), .dinb(new_new_n4205__), .dout(new_new_n4208__));
  and1  g1394(.dina(new_new_n6777__), .dinb(new_new_n6778__), .dout(new_new_n4209__));
  or1   g1395(.dina(new_new_n6779__), .dinb(new_new_n6780__), .dout(new_new_n4210__));
  and1  g1396(.dina(new_new_n6779__), .dinb(new_new_n6780__), .dout(new_new_n4211__));
  or1   g1397(.dina(new_new_n6777__), .dinb(new_new_n6778__), .dout(new_new_n4212__));
  and1  g1398(.dina(new_new_n4210__), .dinb(new_new_n4212__), .dout(new_new_n4213__));
  or1   g1399(.dina(new_new_n4209__), .dinb(new_new_n4211__), .dout(new_new_n4214__));
  and1  g1400(.dina(new_new_n4208__), .dinb(new_new_n4213__), .dout(new_new_n4215__));
  and1  g1401(.dina(new_new_n4207__), .dinb(new_new_n4214__), .dout(new_new_n4216__));
  or1   g1402(.dina(new_new_n4215__), .dinb(new_new_n4216__), .dout(new_new_n4217__));
  or1   g1403(.dina(new_new_n3459__), .dinb(new_new_n6772__), .dout(new_new_n4218__));
  or1   g1404(.dina(new_new_n3429__), .dinb(new_new_n6771__), .dout(new_new_n4219__));
  or1   g1405(.dina(new_new_n3417__), .dinb(new_new_n3433__), .dout(new_new_n4220__));
  and1  g1406(.dina(new_new_n3425__), .dinb(new_new_n4220__), .dout(new_new_n4221__));
  and1  g1407(.dina(new_new_n4219__), .dinb(new_new_n4221__), .dout(new_new_n4222__));
  and1  g1408(.dina(new_new_n4218__), .dinb(new_new_n4222__), .dout(new_new_n4223__));
  or1   g1409(.dina(new_new_n3431__), .dinb(new_new_n6782__), .dout(new_new_n4224__));
  and1  g1410(.dina(new_new_n3685__), .dinb(new_new_n6786__), .dout(new_new_n4225__));
  or1   g1411(.dina(new_new_n6801__), .dinb(new_new_n3448__), .dout(new_new_n4226__));
  and1  g1412(.dina(new_new_n6809__), .dinb(new_new_n3786__), .dout(new_new_n4227__));
  and1  g1413(.dina(new_new_n4226__), .dinb(new_new_n4227__), .dout(new_new_n4228__));
  or1   g1414(.dina(new_new_n4225__), .dinb(new_new_n4228__), .dout(new_new_n4229__));
  or1   g1415(.dina(new_new_n3439__), .dinb(new_new_n6820__), .dout(new_new_n4230__));
  and1  g1416(.dina(new_new_n6824__), .dinb(new_new_n6769__), .dout(new_new_n4231__));
  or1   g1417(.dina(new_new_n6830__), .dinb(new_new_n3785__), .dout(new_new_n4232__));
  or1   g1418(.dina(new_new_n4231__), .dinb(new_new_n4232__), .dout(new_new_n4233__));
  and1  g1419(.dina(new_new_n4230__), .dinb(new_new_n4233__), .dout(new_new_n4234__));
  and1  g1420(.dina(new_new_n6786__), .dinb(new_new_n6832__), .dout(new_new_n4235__));
  or1   g1421(.dina(new_new_n6801__), .dinb(new_new_n3861__), .dout(new_new_n4236__));
  and1  g1422(.dina(new_new_n6809__), .dinb(new_new_n3776__), .dout(new_new_n4237__));
  and1  g1423(.dina(new_new_n4236__), .dinb(new_new_n4237__), .dout(new_new_n4238__));
  or1   g1424(.dina(new_new_n4235__), .dinb(new_new_n4238__), .dout(new_new_n4239__));
  or1   g1425(.dina(new_new_n6837__), .dinb(new_new_n6854__), .dout(new_new_n4240__));
  or1   g1426(.dina(new_new_n6860__), .dinb(new_new_n6877__), .dout(new_new_n4241__));
  and1  g1427(.dina(new_new_n4240__), .dinb(new_new_n4241__), .dout(new_new_n4242__));
  and1  g1428(.dina(new_new_n6882__), .dinb(new_new_n4242__), .dout(new_new_n4243__));
  or1   g1429(.dina(new_new_n6888__), .dinb(new_new_n6837__), .dout(new_new_n4244__));
  or1   g1430(.dina(new_new_n6889__), .dinb(new_new_n6860__), .dout(new_new_n4245__));
  and1  g1431(.dina(new_new_n4244__), .dinb(new_new_n4245__), .dout(new_new_n4246__));
  and1  g1432(.dina(new_new_n6893__), .dinb(new_new_n4246__), .dout(new_new_n4247__));
  or1   g1433(.dina(new_new_n4243__), .dinb(new_new_n4247__), .dout(new_new_n4248__));
  and1  g1434(.dina(new_new_n6899__), .dinb(new_new_n6787__), .dout(new_new_n4249__));
  or1   g1435(.dina(new_new_n3770__), .dinb(new_new_n3798__), .dout(new_new_n4250__));
  and1  g1436(.dina(new_new_n6810__), .dinb(new_new_n4250__), .dout(new_new_n4251__));
  or1   g1437(.dina(new_new_n4249__), .dinb(new_new_n4251__), .dout(new_new_n4252__));
  and1  g1438(.dina(new_new_n6787__), .dinb(new_new_n6900__), .dout(new_new_n4253__));
  and1  g1439(.dina(new_new_n6810__), .dinb(new_new_n3852__), .dout(new_new_n4254__));
  or1   g1440(.dina(new_new_n4253__), .dinb(new_new_n4254__), .dout(new_new_n4255__));
  or1   g1441(.dina(new_new_n3834__), .dinb(new_new_n3837__), .dout(new_new_n4256__));
  and1  g1442(.dina(new_new_n6789__), .dinb(new_new_n6901__), .dout(new_new_n4257__));
  or1   g1443(.dina(new_new_n6800__), .dinb(new_new_n3871__), .dout(new_new_n4258__));
  and1  g1444(.dina(new_new_n6812__), .dinb(new_new_n3778__), .dout(new_new_n4259__));
  and1  g1445(.dina(new_new_n4258__), .dinb(new_new_n4259__), .dout(new_new_n4260__));
  or1   g1446(.dina(new_new_n4257__), .dinb(new_new_n4260__), .dout(new_new_n4261__));
  or1   g1447(.dina(new_new_n6906__), .dinb(new_new_n6854__), .dout(new_new_n4262__));
  or1   g1448(.dina(new_new_n6925__), .dinb(new_new_n6877__), .dout(new_new_n4263__));
  and1  g1449(.dina(new_new_n4262__), .dinb(new_new_n4263__), .dout(new_new_n4264__));
  and1  g1450(.dina(new_new_n6943__), .dinb(new_new_n4264__), .dout(new_new_n4265__));
  or1   g1451(.dina(new_new_n6888__), .dinb(new_new_n6906__), .dout(new_new_n4266__));
  or1   g1452(.dina(new_new_n6889__), .dinb(new_new_n6925__), .dout(new_new_n4267__));
  and1  g1453(.dina(new_new_n4266__), .dinb(new_new_n4267__), .dout(new_new_n4268__));
  and1  g1454(.dina(new_new_n6952__), .dinb(new_new_n4268__), .dout(new_new_n4269__));
  or1   g1455(.dina(new_new_n4265__), .dinb(new_new_n4269__), .dout(new_new_n4270__));
  and1  g1456(.dina(new_new_n3443__), .dinb(new_new_n3827__), .dout(new_new_n4271__));
  and1  g1457(.dina(new_new_n3442__), .dinb(new_new_n3826__), .dout(new_new_n4272__));
  or1   g1458(.dina(new_new_n4271__), .dinb(new_new_n4272__), .dout(new_new_n4273__));
  and1  g1459(.dina(new_new_n6789__), .dinb(new_new_n6958__), .dout(new_new_n4274__));
  and1  g1460(.dina(new_new_n2800__), .dinb(new_new_n6802__), .dout(new_new_n4275__));
  and1  g1461(.dina(new_new_n6824__), .dinb(new_new_n3865__), .dout(new_new_n4276__));
  or1   g1462(.dina(new_new_n4275__), .dinb(new_new_n4276__), .dout(new_new_n4277__));
  and1  g1463(.dina(new_new_n6812__), .dinb(new_new_n4277__), .dout(new_new_n4278__));
  or1   g1464(.dina(new_new_n4274__), .dinb(new_new_n4278__), .dout(new_new_n4279__));
  or1   g1465(.dina(new_new_n3680__), .dinb(new_new_n3833__), .dout(new_new_n4280__));
  and1  g1466(.dina(new_new_n6790__), .dinb(new_new_n6959__), .dout(new_new_n4281__));
  or1   g1467(.dina(new_new_n3782__), .dinb(new_new_n3800__), .dout(new_new_n4282__));
  and1  g1468(.dina(new_new_n6813__), .dinb(new_new_n4282__), .dout(new_new_n4283__));
  or1   g1469(.dina(new_new_n4281__), .dinb(new_new_n4283__), .dout(new_new_n4284__));
  or1   g1470(.dina(new_new_n3598__), .dinb(new_new_n3825__), .dout(new_new_n4285__));
  and1  g1471(.dina(new_new_n6790__), .dinb(new_new_n6960__), .dout(new_new_n4286__));
  and1  g1472(.dina(new_new_n2824__), .dinb(new_new_n6802__), .dout(new_new_n4287__));
  and1  g1473(.dina(new_new_n6823__), .dinb(new_new_n3863__), .dout(new_new_n4288__));
  or1   g1474(.dina(new_new_n4287__), .dinb(new_new_n4288__), .dout(new_new_n4289__));
  and1  g1475(.dina(new_new_n6813__), .dinb(new_new_n4289__), .dout(new_new_n4290__));
  or1   g1476(.dina(new_new_n4286__), .dinb(new_new_n4290__), .dout(new_new_n4291__));
  or1   g1477(.dina(new_new_n6820__), .dinb(new_new_n3880__), .dout(new_new_n4292__));
  and1  g1478(.dina(new_new_n6825__), .dinb(new_new_n6770__), .dout(new_new_n4293__));
  and1  g1479(.dina(new_new_n2817__), .dinb(new_new_n6804__), .dout(new_new_n4294__));
  or1   g1480(.dina(new_new_n6830__), .dinb(new_new_n4294__), .dout(new_new_n4295__));
  or1   g1481(.dina(new_new_n4293__), .dinb(new_new_n4295__), .dout(new_new_n4296__));
  and1  g1482(.dina(new_new_n4292__), .dinb(new_new_n4296__), .dout(new_new_n4297__));
  and1  g1483(.dina(new_new_n3813__), .dinb(new_new_n3815__), .dout(new_new_n4298__));
  or1   g1484(.dina(new_new_n3812__), .dinb(new_new_n3814__), .dout(new_new_n4299__));
  and1  g1485(.dina(new_new_n6963__), .dinb(new_new_n6965__), .dout(new_new_n4300__));
  or1   g1486(.dina(new_new_n6967__), .dinb(new_new_n6969__), .dout(new_new_n4301__));
  and1  g1487(.dina(new_new_n6967__), .dinb(new_new_n6969__), .dout(new_new_n4302__));
  or1   g1488(.dina(new_new_n6963__), .dinb(new_new_n6965__), .dout(new_new_n4303__));
  and1  g1489(.dina(new_new_n4301__), .dinb(new_new_n4303__), .dout(new_new_n4304__));
  or1   g1490(.dina(new_new_n4300__), .dinb(new_new_n4302__), .dout(new_new_n4305__));
  and1  g1491(.dina(new_new_n3828__), .dinb(new_new_n3831__), .dout(new_new_n4306__));
  or1   g1492(.dina(new_new_n3829__), .dinb(new_new_n3830__), .dout(new_new_n4307__));
  and1  g1493(.dina(new_new_n3900__), .dinb(new_new_n3903__), .dout(new_new_n4308__));
  or1   g1494(.dina(new_new_n3901__), .dinb(new_new_n3902__), .dout(new_new_n4309__));
  and1  g1495(.dina(new_new_n6970__), .dinb(new_new_n6971__), .dout(new_new_n4310__));
  or1   g1496(.dina(new_new_n6972__), .dinb(new_new_n6973__), .dout(new_new_n4311__));
  and1  g1497(.dina(new_new_n6972__), .dinb(new_new_n6973__), .dout(new_new_n4312__));
  or1   g1498(.dina(new_new_n6970__), .dinb(new_new_n6971__), .dout(new_new_n4313__));
  and1  g1499(.dina(new_new_n4311__), .dinb(new_new_n4313__), .dout(new_new_n4314__));
  or1   g1500(.dina(new_new_n4310__), .dinb(new_new_n4312__), .dout(new_new_n4315__));
  and1  g1501(.dina(new_new_n4305__), .dinb(new_new_n4314__), .dout(new_new_n4316__));
  and1  g1502(.dina(new_new_n4304__), .dinb(new_new_n4315__), .dout(new_new_n4317__));
  or1   g1503(.dina(new_new_n4316__), .dinb(new_new_n4317__), .dout(new_new_n4318__));
  and1  g1504(.dina(new_new_n6974__), .dinb(new_new_n6975__), .dout(new_new_n4319__));
  or1   g1505(.dina(new_new_n6976__), .dinb(new_new_n6977__), .dout(new_new_n4320__));
  and1  g1506(.dina(new_new_n6976__), .dinb(new_new_n6977__), .dout(new_new_n4321__));
  or1   g1507(.dina(new_new_n6974__), .dinb(new_new_n6975__), .dout(new_new_n4322__));
  and1  g1508(.dina(new_new_n4320__), .dinb(new_new_n4322__), .dout(new_new_n4323__));
  or1   g1509(.dina(new_new_n4319__), .dinb(new_new_n4321__), .dout(new_new_n4324__));
  and1  g1510(.dina(new_new_n6978__), .dinb(new_new_n6979__), .dout(new_new_n4325__));
  or1   g1511(.dina(new_new_n6980__), .dinb(new_new_n6981__), .dout(new_new_n4326__));
  and1  g1512(.dina(new_new_n6980__), .dinb(new_new_n6981__), .dout(new_new_n4327__));
  or1   g1513(.dina(new_new_n6978__), .dinb(new_new_n6979__), .dout(new_new_n4328__));
  and1  g1514(.dina(new_new_n4326__), .dinb(new_new_n4328__), .dout(new_new_n4329__));
  or1   g1515(.dina(new_new_n4325__), .dinb(new_new_n4327__), .dout(new_new_n4330__));
  and1  g1516(.dina(new_new_n6982__), .dinb(new_new_n6983__), .dout(new_new_n4331__));
  or1   g1517(.dina(new_new_n6984__), .dinb(new_new_n6985__), .dout(new_new_n4332__));
  and1  g1518(.dina(new_new_n6984__), .dinb(new_new_n6985__), .dout(new_new_n4333__));
  or1   g1519(.dina(new_new_n6982__), .dinb(new_new_n6983__), .dout(new_new_n4334__));
  and1  g1520(.dina(new_new_n4332__), .dinb(new_new_n4334__), .dout(new_new_n4335__));
  or1   g1521(.dina(new_new_n4331__), .dinb(new_new_n4333__), .dout(new_new_n4336__));
  and1  g1522(.dina(new_new_n6986__), .dinb(new_new_n6987__), .dout(new_new_n4337__));
  or1   g1523(.dina(new_new_n6988__), .dinb(new_new_n6989__), .dout(new_new_n4338__));
  and1  g1524(.dina(new_new_n6988__), .dinb(new_new_n6989__), .dout(new_new_n4339__));
  or1   g1525(.dina(new_new_n6986__), .dinb(new_new_n6987__), .dout(new_new_n4340__));
  and1  g1526(.dina(new_new_n4338__), .dinb(new_new_n4340__), .dout(new_new_n4341__));
  or1   g1527(.dina(new_new_n4337__), .dinb(new_new_n4339__), .dout(new_new_n4342__));
  and1  g1528(.dina(new_new_n6990__), .dinb(new_new_n6991__), .dout(new_new_n4343__));
  or1   g1529(.dina(new_new_n6992__), .dinb(new_new_n6993__), .dout(new_new_n4344__));
  and1  g1530(.dina(new_new_n6992__), .dinb(new_new_n6993__), .dout(new_new_n4345__));
  or1   g1531(.dina(new_new_n6990__), .dinb(new_new_n6991__), .dout(new_new_n4346__));
  and1  g1532(.dina(new_new_n4344__), .dinb(new_new_n4346__), .dout(new_new_n4347__));
  or1   g1533(.dina(new_new_n4343__), .dinb(new_new_n4345__), .dout(new_new_n4348__));
  and1  g1534(.dina(new_new_n6994__), .dinb(new_new_n6995__), .dout(new_new_n4349__));
  or1   g1535(.dina(new_new_n6996__), .dinb(new_new_n6997__), .dout(new_new_n4350__));
  and1  g1536(.dina(new_new_n6996__), .dinb(new_new_n6997__), .dout(new_new_n4351__));
  or1   g1537(.dina(new_new_n6994__), .dinb(new_new_n6995__), .dout(new_new_n4352__));
  and1  g1538(.dina(new_new_n4350__), .dinb(new_new_n4352__), .dout(new_new_n4353__));
  or1   g1539(.dina(new_new_n4349__), .dinb(new_new_n4351__), .dout(new_new_n4354__));
  and1  g1540(.dina(new_new_n4336__), .dinb(new_new_n4353__), .dout(new_new_n4355__));
  and1  g1541(.dina(new_new_n4335__), .dinb(new_new_n4354__), .dout(new_new_n4356__));
  or1   g1542(.dina(new_new_n4355__), .dinb(new_new_n4356__), .dout(new_new_n4357__));
  or1   g1543(.dina(new_new_n3816__), .dinb(new_new_n3818__), .dout(new_new_n4358__));
  or1   g1544(.dina(new_new_n6832__), .dinb(new_new_n3881__), .dout(new_new_n4359__));
  or1   g1545(.dina(new_new_n6960__), .dinb(new_new_n4359__), .dout(new_new_n4360__));
  or1   g1546(.dina(new_new_n6959__), .dinb(new_new_n4360__), .dout(new_new_n4361__));
  or1   g1547(.dina(new_new_n6958__), .dinb(new_new_n4361__), .dout(new_new_n4362__));
  or1   g1548(.dina(new_new_n6998__), .dinb(new_new_n4362__), .dout(new_new_n4363__));
  or1   g1549(.dina(new_new_n6999__), .dinb(new_new_n4363__), .dout(new_new_n4364__));
  or1   g1550(.dina(new_new_n3423__), .dinb(new_new_n3884__), .dout(new_new_n4365__));
  or1   g1551(.dina(new_new_n3422__), .dinb(new_new_n3885__), .dout(new_new_n4366__));
  and1  g1552(.dina(new_new_n4365__), .dinb(new_new_n4366__), .dout(new_new_n4367__));
  or1   g1553(.dina(new_new_n3415__), .dinb(new_new_n3879__), .dout(new_new_n4368__));
  or1   g1554(.dina(new_new_n3414__), .dinb(new_new_n3878__), .dout(new_new_n4369__));
  and1  g1555(.dina(new_new_n4368__), .dinb(new_new_n4369__), .dout(new_new_n4370__));
  or1   g1556(.dina(new_new_n7000__), .dinb(new_new_n7001__), .dout(new_new_n4371__));
  or1   g1557(.dina(new_new_n4364__), .dinb(new_new_n4371__), .dout(new_new_n4372__));
  and1  g1558(.dina(new_new_n3838__), .dinb(new_new_n3841__), .dout(new_new_n4373__));
  and1  g1559(.dina(new_new_n3821__), .dinb(new_new_n3822__), .dout(new_new_n4374__));
  or1   g1560(.dina(new_new_n3438__), .dinb(new_new_n3843__), .dout(new_new_n4375__));
  or1   g1561(.dina(new_new_n6901__), .dinb(new_new_n4375__), .dout(new_new_n4376__));
  or1   g1562(.dina(new_new_n6899__), .dinb(new_new_n4376__), .dout(new_new_n4377__));
  or1   g1563(.dina(new_new_n6900__), .dinb(new_new_n4377__), .dout(new_new_n4378__));
  or1   g1564(.dina(new_new_n7002__), .dinb(new_new_n4378__), .dout(new_new_n4379__));
  or1   g1565(.dina(new_new_n7003__), .dinb(new_new_n4379__), .dout(new_new_n4380__));
  or1   g1566(.dina(new_new_n7004__), .dinb(new_new_n4380__), .dout(new_new_n4381__));
  and1  g1567(.dina(new_new_n7009__), .dinb(new_new_n6876__), .dout(new_new_n4382__));
  and1  g1568(.dina(new_new_n7028__), .dinb(new_new_n6853__), .dout(new_new_n4383__));
  or1   g1569(.dina(new_new_n7046__), .dinb(new_new_n4383__), .dout(new_new_n4384__));
  or1   g1570(.dina(new_new_n4382__), .dinb(new_new_n4384__), .dout(new_new_n4385__));
  and1  g1571(.dina(new_new_n7052__), .dinb(new_new_n7009__), .dout(new_new_n4386__));
  and1  g1572(.dina(new_new_n7053__), .dinb(new_new_n7028__), .dout(new_new_n4387__));
  or1   g1573(.dina(new_new_n7057__), .dinb(new_new_n4387__), .dout(new_new_n4388__));
  or1   g1574(.dina(new_new_n4386__), .dinb(new_new_n4388__), .dout(new_new_n4389__));
  and1  g1575(.dina(new_new_n7067__), .dinb(new_new_n4389__), .dout(new_new_n4390__));
  and1  g1576(.dina(new_new_n4385__), .dinb(new_new_n4390__), .dout(new_new_n4391__));
  and1  g1577(.dina(new_new_n7083__), .dinb(new_new_n6878__), .dout(new_new_n4392__));
  and1  g1578(.dina(new_new_n7102__), .dinb(new_new_n6855__), .dout(new_new_n4393__));
  or1   g1579(.dina(new_new_n7120__), .dinb(new_new_n4393__), .dout(new_new_n4394__));
  or1   g1580(.dina(new_new_n4392__), .dinb(new_new_n4394__), .dout(new_new_n4395__));
  and1  g1581(.dina(new_new_n7052__), .dinb(new_new_n7083__), .dout(new_new_n4396__));
  and1  g1582(.dina(new_new_n7053__), .dinb(new_new_n7102__), .dout(new_new_n4397__));
  or1   g1583(.dina(new_new_n7129__), .dinb(new_new_n4397__), .dout(new_new_n4398__));
  or1   g1584(.dina(new_new_n4396__), .dinb(new_new_n4398__), .dout(new_new_n4399__));
  and1  g1585(.dina(new_new_n7067__), .dinb(new_new_n4399__), .dout(new_new_n4400__));
  and1  g1586(.dina(new_new_n4395__), .dinb(new_new_n4400__), .dout(new_new_n4401__));
  or1   g1587(.dina(new_new_n7135__), .dinb(new_new_n6861__), .dout(new_new_n4402__));
  or1   g1588(.dina(new_new_n7136__), .dinb(new_new_n6838__), .dout(new_new_n4403__));
  and1  g1589(.dina(new_new_n4402__), .dinb(new_new_n4403__), .dout(new_new_n4404__));
  or1   g1590(.dina(new_new_n6882__), .dinb(new_new_n4404__), .dout(new_new_n4405__));
  and1  g1591(.dina(new_new_n6838__), .dinb(new_new_n7139__), .dout(new_new_n4406__));
  and1  g1592(.dina(new_new_n6861__), .dinb(new_new_n7143__), .dout(new_new_n4407__));
  or1   g1593(.dina(new_new_n6893__), .dinb(new_new_n4407__), .dout(new_new_n4408__));
  or1   g1594(.dina(new_new_n4406__), .dinb(new_new_n4408__), .dout(new_new_n4409__));
  and1  g1595(.dina(new_new_n4405__), .dinb(new_new_n4409__), .dout(new_new_n4410__));
  or1   g1596(.dina(new_new_n7145__), .dinb(new_new_n6863__), .dout(new_new_n4411__));
  or1   g1597(.dina(new_new_n7146__), .dinb(new_new_n6840__), .dout(new_new_n4412__));
  and1  g1598(.dina(new_new_n4411__), .dinb(new_new_n4412__), .dout(new_new_n4413__));
  or1   g1599(.dina(new_new_n6883__), .dinb(new_new_n4413__), .dout(new_new_n4414__));
  and1  g1600(.dina(new_new_n6840__), .dinb(new_new_n7149__), .dout(new_new_n4415__));
  and1  g1601(.dina(new_new_n6863__), .dinb(new_new_n7153__), .dout(new_new_n4416__));
  or1   g1602(.dina(new_new_n6894__), .dinb(new_new_n4416__), .dout(new_new_n4417__));
  or1   g1603(.dina(new_new_n4415__), .dinb(new_new_n4417__), .dout(new_new_n4418__));
  and1  g1604(.dina(new_new_n4414__), .dinb(new_new_n4418__), .dout(new_new_n4419__));
  or1   g1605(.dina(new_new_n7155__), .dinb(new_new_n6864__), .dout(new_new_n4420__));
  or1   g1606(.dina(new_new_n7156__), .dinb(new_new_n6841__), .dout(new_new_n4421__));
  and1  g1607(.dina(new_new_n4420__), .dinb(new_new_n4421__), .dout(new_new_n4422__));
  or1   g1608(.dina(new_new_n6883__), .dinb(new_new_n4422__), .dout(new_new_n4423__));
  and1  g1609(.dina(new_new_n6841__), .dinb(new_new_n7159__), .dout(new_new_n4424__));
  and1  g1610(.dina(new_new_n6864__), .dinb(new_new_n7163__), .dout(new_new_n4425__));
  or1   g1611(.dina(new_new_n6894__), .dinb(new_new_n4425__), .dout(new_new_n4426__));
  or1   g1612(.dina(new_new_n4424__), .dinb(new_new_n4426__), .dout(new_new_n4427__));
  and1  g1613(.dina(new_new_n4423__), .dinb(new_new_n4427__), .dout(new_new_n4428__));
  or1   g1614(.dina(new_new_n7165__), .dinb(new_new_n6866__), .dout(new_new_n4429__));
  or1   g1615(.dina(new_new_n7166__), .dinb(new_new_n6843__), .dout(new_new_n4430__));
  and1  g1616(.dina(new_new_n4429__), .dinb(new_new_n4430__), .dout(new_new_n4431__));
  or1   g1617(.dina(new_new_n6884__), .dinb(new_new_n4431__), .dout(new_new_n4432__));
  and1  g1618(.dina(new_new_n6843__), .dinb(new_new_n7169__), .dout(new_new_n4433__));
  and1  g1619(.dina(new_new_n6866__), .dinb(new_new_n7173__), .dout(new_new_n4434__));
  or1   g1620(.dina(new_new_n6895__), .dinb(new_new_n4434__), .dout(new_new_n4435__));
  or1   g1621(.dina(new_new_n4433__), .dinb(new_new_n4435__), .dout(new_new_n4436__));
  and1  g1622(.dina(new_new_n4432__), .dinb(new_new_n4436__), .dout(new_new_n4437__));
  or1   g1623(.dina(new_new_n7135__), .dinb(new_new_n6926__), .dout(new_new_n4438__));
  or1   g1624(.dina(new_new_n7136__), .dinb(new_new_n6907__), .dout(new_new_n4439__));
  and1  g1625(.dina(new_new_n4438__), .dinb(new_new_n4439__), .dout(new_new_n4440__));
  or1   g1626(.dina(new_new_n6943__), .dinb(new_new_n4440__), .dout(new_new_n4441__));
  and1  g1627(.dina(new_new_n6907__), .dinb(new_new_n7139__), .dout(new_new_n4442__));
  and1  g1628(.dina(new_new_n6926__), .dinb(new_new_n7143__), .dout(new_new_n4443__));
  or1   g1629(.dina(new_new_n6952__), .dinb(new_new_n4443__), .dout(new_new_n4444__));
  or1   g1630(.dina(new_new_n4442__), .dinb(new_new_n4444__), .dout(new_new_n4445__));
  and1  g1631(.dina(new_new_n4441__), .dinb(new_new_n4445__), .dout(new_new_n4446__));
  or1   g1632(.dina(new_new_n7145__), .dinb(new_new_n6928__), .dout(new_new_n4447__));
  or1   g1633(.dina(new_new_n7146__), .dinb(new_new_n6909__), .dout(new_new_n4448__));
  and1  g1634(.dina(new_new_n4447__), .dinb(new_new_n4448__), .dout(new_new_n4449__));
  or1   g1635(.dina(new_new_n6944__), .dinb(new_new_n4449__), .dout(new_new_n4450__));
  and1  g1636(.dina(new_new_n6909__), .dinb(new_new_n7149__), .dout(new_new_n4451__));
  and1  g1637(.dina(new_new_n6928__), .dinb(new_new_n7153__), .dout(new_new_n4452__));
  or1   g1638(.dina(new_new_n6953__), .dinb(new_new_n4452__), .dout(new_new_n4453__));
  or1   g1639(.dina(new_new_n4451__), .dinb(new_new_n4453__), .dout(new_new_n4454__));
  and1  g1640(.dina(new_new_n4450__), .dinb(new_new_n4454__), .dout(new_new_n4455__));
  or1   g1641(.dina(new_new_n7155__), .dinb(new_new_n6929__), .dout(new_new_n4456__));
  or1   g1642(.dina(new_new_n7156__), .dinb(new_new_n6910__), .dout(new_new_n4457__));
  and1  g1643(.dina(new_new_n4456__), .dinb(new_new_n4457__), .dout(new_new_n4458__));
  or1   g1644(.dina(new_new_n6944__), .dinb(new_new_n4458__), .dout(new_new_n4459__));
  and1  g1645(.dina(new_new_n6910__), .dinb(new_new_n7159__), .dout(new_new_n4460__));
  and1  g1646(.dina(new_new_n6929__), .dinb(new_new_n7163__), .dout(new_new_n4461__));
  or1   g1647(.dina(new_new_n6953__), .dinb(new_new_n4461__), .dout(new_new_n4462__));
  or1   g1648(.dina(new_new_n4460__), .dinb(new_new_n4462__), .dout(new_new_n4463__));
  and1  g1649(.dina(new_new_n4459__), .dinb(new_new_n4463__), .dout(new_new_n4464__));
  or1   g1650(.dina(new_new_n7165__), .dinb(new_new_n6931__), .dout(new_new_n4465__));
  or1   g1651(.dina(new_new_n7166__), .dinb(new_new_n6912__), .dout(new_new_n4466__));
  and1  g1652(.dina(new_new_n4465__), .dinb(new_new_n4466__), .dout(new_new_n4467__));
  or1   g1653(.dina(new_new_n6945__), .dinb(new_new_n4467__), .dout(new_new_n4468__));
  and1  g1654(.dina(new_new_n6912__), .dinb(new_new_n7169__), .dout(new_new_n4469__));
  and1  g1655(.dina(new_new_n6931__), .dinb(new_new_n7173__), .dout(new_new_n4470__));
  or1   g1656(.dina(new_new_n6954__), .dinb(new_new_n4470__), .dout(new_new_n4471__));
  or1   g1657(.dina(new_new_n4469__), .dinb(new_new_n4471__), .dout(new_new_n4472__));
  and1  g1658(.dina(new_new_n4468__), .dinb(new_new_n4472__), .dout(new_new_n4473__));
  and1  g1659(.dina(new_new_n7010__), .dinb(new_new_n7138__), .dout(new_new_n4474__));
  and1  g1660(.dina(new_new_n7029__), .dinb(new_new_n7142__), .dout(new_new_n4475__));
  or1   g1661(.dina(new_new_n7046__), .dinb(new_new_n4475__), .dout(new_new_n4476__));
  or1   g1662(.dina(new_new_n4474__), .dinb(new_new_n4476__), .dout(new_new_n4477__));
  and1  g1663(.dina(new_new_n7175__), .dinb(new_new_n7010__), .dout(new_new_n4478__));
  and1  g1664(.dina(new_new_n7176__), .dinb(new_new_n7029__), .dout(new_new_n4479__));
  or1   g1665(.dina(new_new_n7057__), .dinb(new_new_n4479__), .dout(new_new_n4480__));
  or1   g1666(.dina(new_new_n4478__), .dinb(new_new_n4480__), .dout(new_new_n4481__));
  and1  g1667(.dina(new_new_n7066__), .dinb(new_new_n4481__), .dout(new_new_n4482__));
  and1  g1668(.dina(new_new_n4477__), .dinb(new_new_n4482__), .dout(new_new_n4483__));
  or1   g1669(.dina(new_new_n7031__), .dinb(new_new_n7168__), .dout(new_new_n4484__));
  or1   g1670(.dina(new_new_n7012__), .dinb(new_new_n7172__), .dout(new_new_n4485__));
  and1  g1671(.dina(new_new_n7058__), .dinb(new_new_n4485__), .dout(new_new_n4486__));
  and1  g1672(.dina(new_new_n4484__), .dinb(new_new_n4486__), .dout(new_new_n4487__));
  or1   g1673(.dina(new_new_n7177__), .dinb(new_new_n7031__), .dout(new_new_n4488__));
  or1   g1674(.dina(new_new_n7178__), .dinb(new_new_n7012__), .dout(new_new_n4489__));
  and1  g1675(.dina(new_new_n7047__), .dinb(new_new_n4489__), .dout(new_new_n4490__));
  and1  g1676(.dina(new_new_n4488__), .dinb(new_new_n4490__), .dout(new_new_n4491__));
  or1   g1677(.dina(new_new_n7180__), .dinb(new_new_n4491__), .dout(new_new_n4492__));
  or1   g1678(.dina(new_new_n4487__), .dinb(new_new_n4492__), .dout(new_new_n4493__));
  and1  g1679(.dina(new_new_n7013__), .dinb(new_new_n7158__), .dout(new_new_n4494__));
  and1  g1680(.dina(new_new_n7032__), .dinb(new_new_n7162__), .dout(new_new_n4495__));
  or1   g1681(.dina(new_new_n7047__), .dinb(new_new_n4495__), .dout(new_new_n4496__));
  or1   g1682(.dina(new_new_n4494__), .dinb(new_new_n4496__), .dout(new_new_n4497__));
  and1  g1683(.dina(new_new_n7182__), .dinb(new_new_n7013__), .dout(new_new_n4498__));
  and1  g1684(.dina(new_new_n7183__), .dinb(new_new_n7032__), .dout(new_new_n4499__));
  or1   g1685(.dina(new_new_n7058__), .dinb(new_new_n4499__), .dout(new_new_n4500__));
  or1   g1686(.dina(new_new_n4498__), .dinb(new_new_n4500__), .dout(new_new_n4501__));
  and1  g1687(.dina(new_new_n7068__), .dinb(new_new_n4501__), .dout(new_new_n4502__));
  and1  g1688(.dina(new_new_n4497__), .dinb(new_new_n4502__), .dout(new_new_n4503__));
  and1  g1689(.dina(new_new_n7015__), .dinb(new_new_n7148__), .dout(new_new_n4504__));
  and1  g1690(.dina(new_new_n7034__), .dinb(new_new_n7152__), .dout(new_new_n4505__));
  or1   g1691(.dina(new_new_n7048__), .dinb(new_new_n4505__), .dout(new_new_n4506__));
  or1   g1692(.dina(new_new_n4504__), .dinb(new_new_n4506__), .dout(new_new_n4507__));
  and1  g1693(.dina(new_new_n7184__), .dinb(new_new_n7015__), .dout(new_new_n4508__));
  and1  g1694(.dina(new_new_n7185__), .dinb(new_new_n7034__), .dout(new_new_n4509__));
  or1   g1695(.dina(new_new_n7059__), .dinb(new_new_n4509__), .dout(new_new_n4510__));
  or1   g1696(.dina(new_new_n4508__), .dinb(new_new_n4510__), .dout(new_new_n4511__));
  and1  g1697(.dina(new_new_n7068__), .dinb(new_new_n4511__), .dout(new_new_n4512__));
  and1  g1698(.dina(new_new_n4507__), .dinb(new_new_n4512__), .dout(new_new_n4513__));
  and1  g1699(.dina(new_new_n7084__), .dinb(new_new_n7140__), .dout(new_new_n4514__));
  and1  g1700(.dina(new_new_n7103__), .dinb(new_new_n7144__), .dout(new_new_n4515__));
  or1   g1701(.dina(new_new_n7120__), .dinb(new_new_n4515__), .dout(new_new_n4516__));
  or1   g1702(.dina(new_new_n4514__), .dinb(new_new_n4516__), .dout(new_new_n4517__));
  and1  g1703(.dina(new_new_n7175__), .dinb(new_new_n7084__), .dout(new_new_n4518__));
  and1  g1704(.dina(new_new_n7176__), .dinb(new_new_n7103__), .dout(new_new_n4519__));
  or1   g1705(.dina(new_new_n7129__), .dinb(new_new_n4519__), .dout(new_new_n4520__));
  or1   g1706(.dina(new_new_n4518__), .dinb(new_new_n4520__), .dout(new_new_n4521__));
  and1  g1707(.dina(new_new_n7070__), .dinb(new_new_n4521__), .dout(new_new_n4522__));
  and1  g1708(.dina(new_new_n4517__), .dinb(new_new_n4522__), .dout(new_new_n4523__));
  or1   g1709(.dina(new_new_n7105__), .dinb(new_new_n7170__), .dout(new_new_n4524__));
  or1   g1710(.dina(new_new_n7086__), .dinb(new_new_n7174__), .dout(new_new_n4525__));
  and1  g1711(.dina(new_new_n7130__), .dinb(new_new_n4525__), .dout(new_new_n4526__));
  and1  g1712(.dina(new_new_n4524__), .dinb(new_new_n4526__), .dout(new_new_n4527__));
  or1   g1713(.dina(new_new_n7177__), .dinb(new_new_n7105__), .dout(new_new_n4528__));
  or1   g1714(.dina(new_new_n7178__), .dinb(new_new_n7086__), .dout(new_new_n4529__));
  and1  g1715(.dina(new_new_n7121__), .dinb(new_new_n4529__), .dout(new_new_n4530__));
  and1  g1716(.dina(new_new_n4528__), .dinb(new_new_n4530__), .dout(new_new_n4531__));
  or1   g1717(.dina(new_new_n7180__), .dinb(new_new_n4531__), .dout(new_new_n4532__));
  or1   g1718(.dina(new_new_n4527__), .dinb(new_new_n4532__), .dout(new_new_n4533__));
  and1  g1719(.dina(new_new_n7087__), .dinb(new_new_n7160__), .dout(new_new_n4534__));
  and1  g1720(.dina(new_new_n7106__), .dinb(new_new_n7164__), .dout(new_new_n4535__));
  or1   g1721(.dina(new_new_n7121__), .dinb(new_new_n4535__), .dout(new_new_n4536__));
  or1   g1722(.dina(new_new_n4534__), .dinb(new_new_n4536__), .dout(new_new_n4537__));
  and1  g1723(.dina(new_new_n7182__), .dinb(new_new_n7087__), .dout(new_new_n4538__));
  and1  g1724(.dina(new_new_n7183__), .dinb(new_new_n7106__), .dout(new_new_n4539__));
  or1   g1725(.dina(new_new_n7130__), .dinb(new_new_n4539__), .dout(new_new_n4540__));
  or1   g1726(.dina(new_new_n4538__), .dinb(new_new_n4540__), .dout(new_new_n4541__));
  and1  g1727(.dina(new_new_n7070__), .dinb(new_new_n4541__), .dout(new_new_n4542__));
  and1  g1728(.dina(new_new_n4537__), .dinb(new_new_n4542__), .dout(new_new_n4543__));
  and1  g1729(.dina(new_new_n7184__), .dinb(new_new_n7089__), .dout(new_new_n4544__));
  and1  g1730(.dina(new_new_n7185__), .dinb(new_new_n7108__), .dout(new_new_n4545__));
  or1   g1731(.dina(new_new_n4544__), .dinb(new_new_n4545__), .dout(new_new_n4546__));
  and1  g1732(.dina(new_new_n7122__), .dinb(new_new_n4546__), .dout(new_new_n4547__));
  or1   g1733(.dina(new_new_n7108__), .dinb(new_new_n7150__), .dout(new_new_n4548__));
  or1   g1734(.dina(new_new_n7089__), .dinb(new_new_n7154__), .dout(new_new_n4549__));
  and1  g1735(.dina(new_new_n7131__), .dinb(new_new_n4549__), .dout(new_new_n4550__));
  and1  g1736(.dina(new_new_n4548__), .dinb(new_new_n4550__), .dout(new_new_n4551__));
  or1   g1737(.dina(new_new_n4547__), .dinb(new_new_n4551__), .dout(new_new_n4552__));
  and1  g1738(.dina(new_new_n7071__), .dinb(new_new_n4552__), .dout(new_new_n4553__));
  or1   g1739(.dina(new_new_n2865__), .dinb(new_new_n3403__), .dout(new_new_n4554__));
  and1  g1740(.dina(new_new_n2808__), .dinb(new_new_n7186__), .dout(new_new_n4555__));
  and1  g1741(.dina(new_new_n7187__), .dinb(new_new_n6962__), .dout(new_new_n4556__));
  or1   g1742(.dina(new_new_n4555__), .dinb(new_new_n4556__), .dout(new_new_n4557__));
  and1  g1743(.dina(new_new_n3338__), .dinb(new_new_n4557__), .dout(new_new_n4558__));
  and1  g1744(.dina(new_new_n7188__), .dinb(new_new_n6782__), .dout(new_new_n4559__));
  or1   g1745(.dina(new_new_n7189__), .dinb(new_new_n7190__), .dout(new_new_n4560__));
  and1  g1746(.dina(new_new_n7189__), .dinb(new_new_n7190__), .dout(new_new_n4561__));
  or1   g1747(.dina(new_new_n7188__), .dinb(new_new_n6781__), .dout(new_new_n4562__));
  and1  g1748(.dina(new_new_n4560__), .dinb(new_new_n4562__), .dout(new_new_n4563__));
  or1   g1749(.dina(new_new_n4559__), .dinb(new_new_n4561__), .dout(new_new_n4564__));
  and1  g1750(.dina(new_new_n7187__), .dinb(new_new_n7191__), .dout(new_new_n4565__));
  and1  g1751(.dina(new_new_n7186__), .dinb(new_new_n3446__), .dout(new_new_n4566__));
  or1   g1752(.dina(new_new_n4565__), .dinb(new_new_n4566__), .dout(new_new_n4567__));
  and1  g1753(.dina(new_new_n3339__), .dinb(new_new_n4567__), .dout(new_new_n4568__));
  or1   g1754(.dina(new_new_n4558__), .dinb(new_new_n4568__), .dout(new_new_n4569__));
  and1  g1755(.dina(new_new_n4554__), .dinb(new_new_n4569__), .dout(new_new_n4570__));
  or1   g1756(.dina(new_new_n6968__), .dinb(new_new_n4563__), .dout(new_new_n4571__));
  or1   g1757(.dina(new_new_n6964__), .dinb(new_new_n7191__), .dout(new_new_n4572__));
  and1  g1758(.dina(new_new_n4571__), .dinb(new_new_n4572__), .dout(new_new_n4573__));
  and1  g1759(.dina(new_new_n6964__), .dinb(new_new_n6793__), .dout(new_new_n4574__));
  and1  g1760(.dina(new_new_n3794__), .dinb(new_new_n3803__), .dout(new_new_n4575__));
  or1   g1761(.dina(new_new_n4574__), .dinb(new_new_n4575__), .dout(new_new_n4576__));
  and1  g1762(.dina(new_new_n6793__), .dinb(new_new_n7004__), .dout(new_new_n4577__));
  or1   g1763(.dina(new_new_n3780__), .dinb(new_new_n3804__), .dout(new_new_n4578__));
  and1  g1764(.dina(new_new_n6816__), .dinb(new_new_n4578__), .dout(new_new_n4579__));
  or1   g1765(.dina(new_new_n4577__), .dinb(new_new_n4579__), .dout(new_new_n4580__));
  and1  g1766(.dina(new_new_n6794__), .dinb(new_new_n7003__), .dout(new_new_n4581__));
  or1   g1767(.dina(new_new_n3774__), .dinb(new_new_n3806__), .dout(new_new_n4582__));
  and1  g1768(.dina(new_new_n6816__), .dinb(new_new_n4582__), .dout(new_new_n4583__));
  or1   g1769(.dina(new_new_n4581__), .dinb(new_new_n4583__), .dout(new_new_n4584__));
  and1  g1770(.dina(new_new_n6794__), .dinb(new_new_n7002__), .dout(new_new_n4585__));
  and1  g1771(.dina(new_new_n6817__), .dinb(new_new_n3848__), .dout(new_new_n4586__));
  or1   g1772(.dina(new_new_n4585__), .dinb(new_new_n4586__), .dout(new_new_n4587__));
  or1   g1773(.dina(new_new_n7192__), .dinb(new_new_n7193__), .dout(new_new_n4588__));
  or1   g1774(.dina(new_new_n7194__), .dinb(new_new_n4588__), .dout(new_new_n4589__));
  or1   g1775(.dina(new_new_n7195__), .dinb(new_new_n4589__), .dout(new_new_n4590__));
  or1   g1776(.dina(new_new_n7196__), .dinb(new_new_n4590__), .dout(new_new_n4591__));
  or1   g1777(.dina(new_new_n7197__), .dinb(new_new_n4591__), .dout(new_new_n4592__));
  or1   g1778(.dina(new_new_n7198__), .dinb(new_new_n4592__), .dout(new_new_n4593__));
  or1   g1779(.dina(new_new_n7199__), .dinb(new_new_n4593__), .dout(new_new_n4594__));
  and1  g1780(.dina(new_new_n6796__), .dinb(new_new_n6999__), .dout(new_new_n4595__));
  and1  g1781(.dina(new_new_n6817__), .dinb(new_new_n3850__), .dout(new_new_n4596__));
  or1   g1782(.dina(new_new_n4595__), .dinb(new_new_n4596__), .dout(new_new_n4597__));
  and1  g1783(.dina(new_new_n6796__), .dinb(new_new_n7000__), .dout(new_new_n4598__));
  and1  g1784(.dina(new_new_n2746__), .dinb(new_new_n6804__), .dout(new_new_n4599__));
  and1  g1785(.dina(new_new_n6825__), .dinb(new_new_n3867__), .dout(new_new_n4600__));
  or1   g1786(.dina(new_new_n4599__), .dinb(new_new_n4600__), .dout(new_new_n4601__));
  and1  g1787(.dina(new_new_n6819__), .dinb(new_new_n4601__), .dout(new_new_n4602__));
  or1   g1788(.dina(new_new_n4598__), .dinb(new_new_n4602__), .dout(new_new_n4603__));
  and1  g1789(.dina(new_new_n6797__), .dinb(new_new_n7001__), .dout(new_new_n4604__));
  and1  g1790(.dina(new_new_n2552__), .dinb(new_new_n6805__), .dout(new_new_n4605__));
  and1  g1791(.dina(new_new_n6827__), .dinb(new_new_n3869__), .dout(new_new_n4606__));
  or1   g1792(.dina(new_new_n4605__), .dinb(new_new_n4606__), .dout(new_new_n4607__));
  and1  g1793(.dina(new_new_n6819__), .dinb(new_new_n4607__), .dout(new_new_n4608__));
  or1   g1794(.dina(new_new_n4604__), .dinb(new_new_n4608__), .dout(new_new_n4609__));
  and1  g1795(.dina(new_new_n6797__), .dinb(new_new_n6998__), .dout(new_new_n4610__));
  or1   g1796(.dina(new_new_n3772__), .dinb(new_new_n3808__), .dout(new_new_n4611__));
  and1  g1797(.dina(new_new_n6818__), .dinb(new_new_n4611__), .dout(new_new_n4612__));
  or1   g1798(.dina(new_new_n4610__), .dinb(new_new_n4612__), .dout(new_new_n4613__));
  and1  g1799(.dina(new_new_n7200__), .dinb(new_new_n6913__), .dout(new_new_n4614__));
  and1  g1800(.dina(new_new_n7201__), .dinb(new_new_n6932__), .dout(new_new_n4615__));
  or1   g1801(.dina(new_new_n4614__), .dinb(new_new_n4615__), .dout(new_new_n4616__));
  and1  g1802(.dina(new_new_n6954__), .dinb(new_new_n4616__), .dout(new_new_n4617__));
  and1  g1803(.dina(new_new_n6913__), .dinb(new_new_n7204__), .dout(new_new_n4618__));
  and1  g1804(.dina(new_new_n6932__), .dinb(new_new_n7208__), .dout(new_new_n4619__));
  or1   g1805(.dina(new_new_n4618__), .dinb(new_new_n4619__), .dout(new_new_n4620__));
  and1  g1806(.dina(new_new_n6945__), .dinb(new_new_n4620__), .dout(new_new_n4621__));
  or1   g1807(.dina(new_new_n4617__), .dinb(new_new_n4621__), .dout(new_new_n4622__));
  and1  g1808(.dina(new_new_n6844__), .dinb(new_new_n7204__), .dout(new_new_n4623__));
  and1  g1809(.dina(new_new_n6867__), .dinb(new_new_n7208__), .dout(new_new_n4624__));
  or1   g1810(.dina(new_new_n6895__), .dinb(new_new_n4624__), .dout(new_new_n4625__));
  or1   g1811(.dina(new_new_n4623__), .dinb(new_new_n4625__), .dout(new_new_n4626__));
  or1   g1812(.dina(new_new_n7200__), .dinb(new_new_n6867__), .dout(new_new_n4627__));
  or1   g1813(.dina(new_new_n7201__), .dinb(new_new_n6844__), .dout(new_new_n4628__));
  and1  g1814(.dina(new_new_n4627__), .dinb(new_new_n4628__), .dout(new_new_n4629__));
  or1   g1815(.dina(new_new_n6884__), .dinb(new_new_n4629__), .dout(new_new_n4630__));
  and1  g1816(.dina(new_new_n4626__), .dinb(new_new_n4630__), .dout(new_new_n4631__));
  or1   g1817(.dina(new_new_n7210__), .dinb(new_new_n6870__), .dout(new_new_n4632__));
  or1   g1818(.dina(new_new_n7211__), .dinb(new_new_n6847__), .dout(new_new_n4633__));
  and1  g1819(.dina(new_new_n4632__), .dinb(new_new_n4633__), .dout(new_new_n4634__));
  or1   g1820(.dina(new_new_n6886__), .dinb(new_new_n4634__), .dout(new_new_n4635__));
  and1  g1821(.dina(new_new_n6847__), .dinb(new_new_n7214__), .dout(new_new_n4636__));
  and1  g1822(.dina(new_new_n6870__), .dinb(new_new_n7218__), .dout(new_new_n4637__));
  or1   g1823(.dina(new_new_n6897__), .dinb(new_new_n4637__), .dout(new_new_n4638__));
  or1   g1824(.dina(new_new_n4636__), .dinb(new_new_n4638__), .dout(new_new_n4639__));
  and1  g1825(.dina(new_new_n4635__), .dinb(new_new_n4639__), .dout(new_new_n4640__));
  or1   g1826(.dina(new_new_n7220__), .dinb(new_new_n6871__), .dout(new_new_n4641__));
  or1   g1827(.dina(new_new_n7221__), .dinb(new_new_n6848__), .dout(new_new_n4642__));
  and1  g1828(.dina(new_new_n4641__), .dinb(new_new_n4642__), .dout(new_new_n4643__));
  or1   g1829(.dina(new_new_n6886__), .dinb(new_new_n4643__), .dout(new_new_n4644__));
  and1  g1830(.dina(new_new_n6848__), .dinb(new_new_n7224__), .dout(new_new_n4645__));
  and1  g1831(.dina(new_new_n6871__), .dinb(new_new_n7228__), .dout(new_new_n4646__));
  or1   g1832(.dina(new_new_n6897__), .dinb(new_new_n4646__), .dout(new_new_n4647__));
  or1   g1833(.dina(new_new_n4645__), .dinb(new_new_n4647__), .dout(new_new_n4648__));
  and1  g1834(.dina(new_new_n4644__), .dinb(new_new_n4648__), .dout(new_new_n4649__));
  or1   g1835(.dina(new_new_n7230__), .dinb(new_new_n6873__), .dout(new_new_n4650__));
  or1   g1836(.dina(new_new_n7231__), .dinb(new_new_n6850__), .dout(new_new_n4651__));
  and1  g1837(.dina(new_new_n4650__), .dinb(new_new_n4651__), .dout(new_new_n4652__));
  or1   g1838(.dina(new_new_n6887__), .dinb(new_new_n4652__), .dout(new_new_n4653__));
  and1  g1839(.dina(new_new_n6850__), .dinb(new_new_n7234__), .dout(new_new_n4654__));
  and1  g1840(.dina(new_new_n6873__), .dinb(new_new_n7238__), .dout(new_new_n4655__));
  or1   g1841(.dina(new_new_n6898__), .dinb(new_new_n4655__), .dout(new_new_n4656__));
  or1   g1842(.dina(new_new_n4654__), .dinb(new_new_n4656__), .dout(new_new_n4657__));
  and1  g1843(.dina(new_new_n4653__), .dinb(new_new_n4657__), .dout(new_new_n4658__));
  or1   g1844(.dina(new_new_n7210__), .dinb(new_new_n6935__), .dout(new_new_n4659__));
  or1   g1845(.dina(new_new_n7211__), .dinb(new_new_n6916__), .dout(new_new_n4660__));
  and1  g1846(.dina(new_new_n4659__), .dinb(new_new_n4660__), .dout(new_new_n4661__));
  or1   g1847(.dina(new_new_n6947__), .dinb(new_new_n4661__), .dout(new_new_n4662__));
  and1  g1848(.dina(new_new_n6916__), .dinb(new_new_n7214__), .dout(new_new_n4663__));
  and1  g1849(.dina(new_new_n6935__), .dinb(new_new_n7218__), .dout(new_new_n4664__));
  or1   g1850(.dina(new_new_n6956__), .dinb(new_new_n4664__), .dout(new_new_n4665__));
  or1   g1851(.dina(new_new_n4663__), .dinb(new_new_n4665__), .dout(new_new_n4666__));
  and1  g1852(.dina(new_new_n4662__), .dinb(new_new_n4666__), .dout(new_new_n4667__));
  or1   g1853(.dina(new_new_n7220__), .dinb(new_new_n6936__), .dout(new_new_n4668__));
  or1   g1854(.dina(new_new_n7221__), .dinb(new_new_n6917__), .dout(new_new_n4669__));
  and1  g1855(.dina(new_new_n4668__), .dinb(new_new_n4669__), .dout(new_new_n4670__));
  or1   g1856(.dina(new_new_n6947__), .dinb(new_new_n4670__), .dout(new_new_n4671__));
  and1  g1857(.dina(new_new_n6917__), .dinb(new_new_n7224__), .dout(new_new_n4672__));
  and1  g1858(.dina(new_new_n6936__), .dinb(new_new_n7228__), .dout(new_new_n4673__));
  or1   g1859(.dina(new_new_n6956__), .dinb(new_new_n4673__), .dout(new_new_n4674__));
  or1   g1860(.dina(new_new_n4672__), .dinb(new_new_n4674__), .dout(new_new_n4675__));
  and1  g1861(.dina(new_new_n4671__), .dinb(new_new_n4675__), .dout(new_new_n4676__));
  or1   g1862(.dina(new_new_n7230__), .dinb(new_new_n6938__), .dout(new_new_n4677__));
  or1   g1863(.dina(new_new_n7231__), .dinb(new_new_n6919__), .dout(new_new_n4678__));
  and1  g1864(.dina(new_new_n4677__), .dinb(new_new_n4678__), .dout(new_new_n4679__));
  or1   g1865(.dina(new_new_n6948__), .dinb(new_new_n4679__), .dout(new_new_n4680__));
  and1  g1866(.dina(new_new_n6919__), .dinb(new_new_n7234__), .dout(new_new_n4681__));
  and1  g1867(.dina(new_new_n6938__), .dinb(new_new_n7238__), .dout(new_new_n4682__));
  or1   g1868(.dina(new_new_n6957__), .dinb(new_new_n4682__), .dout(new_new_n4683__));
  or1   g1869(.dina(new_new_n4681__), .dinb(new_new_n4683__), .dout(new_new_n4684__));
  and1  g1870(.dina(new_new_n4680__), .dinb(new_new_n4684__), .dout(new_new_n4685__));
  and1  g1871(.dina(new_new_n7016__), .dinb(new_new_n7233__), .dout(new_new_n4686__));
  and1  g1872(.dina(new_new_n7035__), .dinb(new_new_n7237__), .dout(new_new_n4687__));
  or1   g1873(.dina(new_new_n7048__), .dinb(new_new_n4687__), .dout(new_new_n4688__));
  or1   g1874(.dina(new_new_n4686__), .dinb(new_new_n4688__), .dout(new_new_n4689__));
  and1  g1875(.dina(new_new_n7240__), .dinb(new_new_n7016__), .dout(new_new_n4690__));
  and1  g1876(.dina(new_new_n7241__), .dinb(new_new_n7035__), .dout(new_new_n4691__));
  or1   g1877(.dina(new_new_n7059__), .dinb(new_new_n4691__), .dout(new_new_n4692__));
  or1   g1878(.dina(new_new_n4690__), .dinb(new_new_n4692__), .dout(new_new_n4693__));
  and1  g1879(.dina(new_new_n7071__), .dinb(new_new_n4693__), .dout(new_new_n4694__));
  and1  g1880(.dina(new_new_n4689__), .dinb(new_new_n4694__), .dout(new_new_n4695__));
  and1  g1881(.dina(new_new_n7019__), .dinb(new_new_n7223__), .dout(new_new_n4696__));
  and1  g1882(.dina(new_new_n7038__), .dinb(new_new_n7227__), .dout(new_new_n4697__));
  or1   g1883(.dina(new_new_n7050__), .dinb(new_new_n4697__), .dout(new_new_n4698__));
  or1   g1884(.dina(new_new_n4696__), .dinb(new_new_n4698__), .dout(new_new_n4699__));
  and1  g1885(.dina(new_new_n7242__), .dinb(new_new_n7019__), .dout(new_new_n4700__));
  and1  g1886(.dina(new_new_n7243__), .dinb(new_new_n7038__), .dout(new_new_n4701__));
  or1   g1887(.dina(new_new_n7061__), .dinb(new_new_n4701__), .dout(new_new_n4702__));
  or1   g1888(.dina(new_new_n4700__), .dinb(new_new_n4702__), .dout(new_new_n4703__));
  and1  g1889(.dina(new_new_n7074__), .dinb(new_new_n4703__), .dout(new_new_n4704__));
  and1  g1890(.dina(new_new_n4699__), .dinb(new_new_n4704__), .dout(new_new_n4705__));
  and1  g1891(.dina(new_new_n7020__), .dinb(new_new_n7213__), .dout(new_new_n4706__));
  and1  g1892(.dina(new_new_n7039__), .dinb(new_new_n7217__), .dout(new_new_n4707__));
  or1   g1893(.dina(new_new_n7050__), .dinb(new_new_n4707__), .dout(new_new_n4708__));
  or1   g1894(.dina(new_new_n4706__), .dinb(new_new_n4708__), .dout(new_new_n4709__));
  and1  g1895(.dina(new_new_n7244__), .dinb(new_new_n7020__), .dout(new_new_n4710__));
  and1  g1896(.dina(new_new_n7245__), .dinb(new_new_n7039__), .dout(new_new_n4711__));
  or1   g1897(.dina(new_new_n7061__), .dinb(new_new_n4711__), .dout(new_new_n4712__));
  or1   g1898(.dina(new_new_n4710__), .dinb(new_new_n4712__), .dout(new_new_n4713__));
  and1  g1899(.dina(new_new_n7074__), .dinb(new_new_n4713__), .dout(new_new_n4714__));
  and1  g1900(.dina(new_new_n4709__), .dinb(new_new_n4714__), .dout(new_new_n4715__));
  and1  g1901(.dina(new_new_n7246__), .dinb(new_new_n7022__), .dout(new_new_n4716__));
  and1  g1902(.dina(new_new_n7247__), .dinb(new_new_n7041__), .dout(new_new_n4717__));
  or1   g1903(.dina(new_new_n4716__), .dinb(new_new_n4717__), .dout(new_new_n4718__));
  and1  g1904(.dina(new_new_n7051__), .dinb(new_new_n4718__), .dout(new_new_n4719__));
  and1  g1905(.dina(new_new_n7022__), .dinb(new_new_n7203__), .dout(new_new_n4720__));
  and1  g1906(.dina(new_new_n7041__), .dinb(new_new_n7207__), .dout(new_new_n4721__));
  or1   g1907(.dina(new_new_n4720__), .dinb(new_new_n4721__), .dout(new_new_n4722__));
  and1  g1908(.dina(new_new_n7062__), .dinb(new_new_n4722__), .dout(new_new_n4723__));
  or1   g1909(.dina(new_new_n4719__), .dinb(new_new_n4723__), .dout(new_new_n4724__));
  and1  g1910(.dina(new_new_n7075__), .dinb(new_new_n4724__), .dout(new_new_n4725__));
  and1  g1911(.dina(new_new_n7240__), .dinb(new_new_n7090__), .dout(new_new_n4726__));
  and1  g1912(.dina(new_new_n7241__), .dinb(new_new_n7109__), .dout(new_new_n4727__));
  or1   g1913(.dina(new_new_n4726__), .dinb(new_new_n4727__), .dout(new_new_n4728__));
  and1  g1914(.dina(new_new_n7122__), .dinb(new_new_n4728__), .dout(new_new_n4729__));
  or1   g1915(.dina(new_new_n7109__), .dinb(new_new_n7235__), .dout(new_new_n4730__));
  or1   g1916(.dina(new_new_n7090__), .dinb(new_new_n7239__), .dout(new_new_n4731__));
  and1  g1917(.dina(new_new_n7131__), .dinb(new_new_n4731__), .dout(new_new_n4732__));
  and1  g1918(.dina(new_new_n4730__), .dinb(new_new_n4732__), .dout(new_new_n4733__));
  or1   g1919(.dina(new_new_n4729__), .dinb(new_new_n4733__), .dout(new_new_n4734__));
  and1  g1920(.dina(new_new_n7075__), .dinb(new_new_n4734__), .dout(new_new_n4735__));
  and1  g1921(.dina(new_new_n7093__), .dinb(new_new_n7225__), .dout(new_new_n4736__));
  and1  g1922(.dina(new_new_n7112__), .dinb(new_new_n7229__), .dout(new_new_n4737__));
  or1   g1923(.dina(new_new_n7124__), .dinb(new_new_n4737__), .dout(new_new_n4738__));
  or1   g1924(.dina(new_new_n4736__), .dinb(new_new_n4738__), .dout(new_new_n4739__));
  and1  g1925(.dina(new_new_n7242__), .dinb(new_new_n7093__), .dout(new_new_n4740__));
  and1  g1926(.dina(new_new_n7243__), .dinb(new_new_n7112__), .dout(new_new_n4741__));
  or1   g1927(.dina(new_new_n7133__), .dinb(new_new_n4741__), .dout(new_new_n4742__));
  or1   g1928(.dina(new_new_n4740__), .dinb(new_new_n4742__), .dout(new_new_n4743__));
  and1  g1929(.dina(new_new_n7077__), .dinb(new_new_n4743__), .dout(new_new_n4744__));
  and1  g1930(.dina(new_new_n4739__), .dinb(new_new_n4744__), .dout(new_new_n4745__));
  and1  g1931(.dina(new_new_n7094__), .dinb(new_new_n7215__), .dout(new_new_n4746__));
  and1  g1932(.dina(new_new_n7113__), .dinb(new_new_n7219__), .dout(new_new_n4747__));
  or1   g1933(.dina(new_new_n7124__), .dinb(new_new_n4747__), .dout(new_new_n4748__));
  or1   g1934(.dina(new_new_n4746__), .dinb(new_new_n4748__), .dout(new_new_n4749__));
  and1  g1935(.dina(new_new_n7244__), .dinb(new_new_n7094__), .dout(new_new_n4750__));
  and1  g1936(.dina(new_new_n7245__), .dinb(new_new_n7113__), .dout(new_new_n4751__));
  or1   g1937(.dina(new_new_n7133__), .dinb(new_new_n4751__), .dout(new_new_n4752__));
  or1   g1938(.dina(new_new_n4750__), .dinb(new_new_n4752__), .dout(new_new_n4753__));
  and1  g1939(.dina(new_new_n7077__), .dinb(new_new_n4753__), .dout(new_new_n4754__));
  and1  g1940(.dina(new_new_n4749__), .dinb(new_new_n4754__), .dout(new_new_n4755__));
  and1  g1941(.dina(new_new_n7096__), .dinb(new_new_n7205__), .dout(new_new_n4756__));
  and1  g1942(.dina(new_new_n7115__), .dinb(new_new_n7209__), .dout(new_new_n4757__));
  or1   g1943(.dina(new_new_n7125__), .dinb(new_new_n4757__), .dout(new_new_n4758__));
  or1   g1944(.dina(new_new_n4756__), .dinb(new_new_n4758__), .dout(new_new_n4759__));
  and1  g1945(.dina(new_new_n7246__), .dinb(new_new_n7096__), .dout(new_new_n4760__));
  and1  g1946(.dina(new_new_n7247__), .dinb(new_new_n7115__), .dout(new_new_n4761__));
  or1   g1947(.dina(new_new_n7134__), .dinb(new_new_n4761__), .dout(new_new_n4762__));
  or1   g1948(.dina(new_new_n4760__), .dinb(new_new_n4762__), .dout(new_new_n4763__));
  and1  g1949(.dina(new_new_n7078__), .dinb(new_new_n4763__), .dout(new_new_n4764__));
  and1  g1950(.dina(new_new_n4759__), .dinb(new_new_n4764__), .dout(new_new_n4765__));
  or1   g1951(.dina(new_new_n3796__), .dinb(new_new_n3811__), .dout(new_new_n4766__));
  or1   g1952(.dina(new_new_n6831__), .dinb(new_new_n6827__), .dout(new_new_n4767__));
  or1   g1953(.dina(new_new_n2786__), .dinb(new_new_n7248__), .dout(new_new_n4768__));
  and1  g1954(.dina(new_new_n7249__), .dinb(new_new_n4768__), .dout(new_new_n4769__));
  and1  g1955(.dina(new_new_n6831__), .dinb(new_new_n3907__), .dout(new_new_n4770__));
  or1   g1956(.dina(new_new_n6805__), .dinb(new_new_n3874__), .dout(new_new_n4771__));
  or1   g1957(.dina(new_new_n4770__), .dinb(new_new_n4771__), .dout(new_new_n4772__));
  or1   g1958(.dina(new_new_n2772__), .dinb(new_new_n7248__), .dout(new_new_n4773__));
  and1  g1959(.dina(new_new_n7250__), .dinb(new_new_n4773__), .dout(new_new_n4774__));
  and1  g1960(.dina(new_new_n7251__), .dinb(new_new_n6851__), .dout(new_new_n4775__));
  and1  g1961(.dina(new_new_n7252__), .dinb(new_new_n6874__), .dout(new_new_n4776__));
  or1   g1962(.dina(new_new_n4775__), .dinb(new_new_n4776__), .dout(new_new_n4777__));
  and1  g1963(.dina(new_new_n6898__), .dinb(new_new_n4777__), .dout(new_new_n4778__));
  or1   g1964(.dina(new_new_n2695__), .dinb(new_new_n6828__), .dout(new_new_n4779__));
  and1  g1965(.dina(new_new_n7250__), .dinb(new_new_n4779__), .dout(new_new_n4780__));
  or1   g1966(.dina(new_new_n6874__), .dinb(new_new_n7254__), .dout(new_new_n4781__));
  or1   g1967(.dina(new_new_n2687__), .dinb(new_new_n6828__), .dout(new_new_n4782__));
  and1  g1968(.dina(new_new_n7249__), .dinb(new_new_n4782__), .dout(new_new_n4783__));
  or1   g1969(.dina(new_new_n6851__), .dinb(new_new_n7257__), .dout(new_new_n4784__));
  and1  g1970(.dina(new_new_n6887__), .dinb(new_new_n4784__), .dout(new_new_n4785__));
  and1  g1971(.dina(new_new_n4781__), .dinb(new_new_n4785__), .dout(new_new_n4786__));
  or1   g1972(.dina(new_new_n4778__), .dinb(new_new_n4786__), .dout(new_new_n4787__));
  and1  g1973(.dina(new_new_n7251__), .dinb(new_new_n6920__), .dout(new_new_n4788__));
  and1  g1974(.dina(new_new_n7252__), .dinb(new_new_n6939__), .dout(new_new_n4789__));
  or1   g1975(.dina(new_new_n4788__), .dinb(new_new_n4789__), .dout(new_new_n4790__));
  and1  g1976(.dina(new_new_n6957__), .dinb(new_new_n4790__), .dout(new_new_n4791__));
  or1   g1977(.dina(new_new_n6939__), .dinb(new_new_n7254__), .dout(new_new_n4792__));
  or1   g1978(.dina(new_new_n6920__), .dinb(new_new_n7257__), .dout(new_new_n4793__));
  and1  g1979(.dina(new_new_n6948__), .dinb(new_new_n4793__), .dout(new_new_n4794__));
  and1  g1980(.dina(new_new_n4792__), .dinb(new_new_n4794__), .dout(new_new_n4795__));
  or1   g1981(.dina(new_new_n4791__), .dinb(new_new_n4795__), .dout(new_new_n4796__));
  or1   g1982(.dina(new_new_n7042__), .dinb(new_new_n7255__), .dout(new_new_n4797__));
  or1   g1983(.dina(new_new_n7023__), .dinb(new_new_n7258__), .dout(new_new_n4798__));
  and1  g1984(.dina(new_new_n7062__), .dinb(new_new_n4798__), .dout(new_new_n4799__));
  and1  g1985(.dina(new_new_n4797__), .dinb(new_new_n4799__), .dout(new_new_n4800__));
  or1   g1986(.dina(new_new_n7259__), .dinb(new_new_n7042__), .dout(new_new_n4801__));
  or1   g1987(.dina(new_new_n7260__), .dinb(new_new_n7023__), .dout(new_new_n4802__));
  and1  g1988(.dina(new_new_n7051__), .dinb(new_new_n4802__), .dout(new_new_n4803__));
  and1  g1989(.dina(new_new_n4801__), .dinb(new_new_n4803__), .dout(new_new_n4804__));
  or1   g1990(.dina(new_new_n7181__), .dinb(new_new_n4804__), .dout(new_new_n4805__));
  or1   g1991(.dina(new_new_n4800__), .dinb(new_new_n4805__), .dout(new_new_n4806__));
  or1   g1992(.dina(new_new_n7259__), .dinb(new_new_n7116__), .dout(new_new_n4807__));
  or1   g1993(.dina(new_new_n7260__), .dinb(new_new_n7097__), .dout(new_new_n4808__));
  and1  g1994(.dina(new_new_n4807__), .dinb(new_new_n4808__), .dout(new_new_n4809__));
  or1   g1995(.dina(new_new_n7134__), .dinb(new_new_n4809__), .dout(new_new_n4810__));
  and1  g1996(.dina(new_new_n7097__), .dinb(new_new_n7255__), .dout(new_new_n4811__));
  and1  g1997(.dina(new_new_n7116__), .dinb(new_new_n7258__), .dout(new_new_n4812__));
  or1   g1998(.dina(new_new_n7125__), .dinb(new_new_n4812__), .dout(new_new_n4813__));
  or1   g1999(.dina(new_new_n4811__), .dinb(new_new_n4813__), .dout(new_new_n4814__));
  and1  g2000(.dina(new_new_n4810__), .dinb(new_new_n4814__), .dout(new_new_n4815__));
  or1   g2001(.dina(new_new_n7181__), .dinb(new_new_n4815__), .dout(new_new_n4816__));
  and1  g2002(.dina(new_new_n7262__), .dinb(new_new_n7264__), .dout(new_new_n4817__));
  or1   g2003(.dina(new_new_n7266__), .dinb(new_new_n7268__), .dout(new_new_n4818__));
  and1  g2004(.dina(new_new_n7266__), .dinb(new_new_n7268__), .dout(new_new_n4819__));
  or1   g2005(.dina(new_new_n7262__), .dinb(new_new_n7264__), .dout(new_new_n4820__));
  and1  g2006(.dina(new_new_n7269__), .dinb(new_new_n4820__), .dout(new_new_n4821__));
  or1   g2007(.dina(new_new_n4817__), .dinb(new_new_n4819__), .dout(new_new_n4822__));
  or1   g2008(.dina(new_new_n7272__), .dinb(new_new_n7274__), .dout(new_new_n4823__));
  and1  g2009(.dina(new_new_n7276__), .dinb(new_new_n3600__), .dout(new_new_n4824__));
  or1   g2010(.dina(new_new_n3566__), .dinb(new_new_n4824__), .dout(new_new_n4825__));
  and1  g2011(.dina(new_new_n7278__), .dinb(new_new_n7279__), .dout(new_new_n4826__));
  and1  g2012(.dina(new_new_n3709__), .dinb(new_new_n3913__), .dout(new_new_n4827__));
  or1   g2013(.dina(new_new_n3708__), .dinb(new_new_n3912__), .dout(new_new_n4828__));
  and1  g2014(.dina(new_new_n3935__), .dinb(new_new_n7280__), .dout(new_new_n4829__));
  or1   g2015(.dina(new_new_n3934__), .dinb(new_new_n7282__), .dout(new_new_n4830__));
  and1  g2016(.dina(new_new_n4033__), .dinb(new_new_n4035__), .dout(new_new_n4831__));
  or1   g2017(.dina(new_new_n4032__), .dinb(new_new_n4034__), .dout(new_new_n4832__));
  and1  g2018(.dina(new_new_n4037__), .dinb(new_new_n4039__), .dout(new_new_n4833__));
  or1   g2019(.dina(new_new_n4036__), .dinb(new_new_n4038__), .dout(new_new_n4834__));
  and1  g2020(.dina(new_new_n4045__), .dinb(new_new_n7283__), .dout(new_new_n4835__));
  or1   g2021(.dina(new_new_n4044__), .dinb(new_new_n7284__), .dout(new_new_n4836__));
  and1  g2022(.dina(new_new_n7283__), .dinb(new_new_n4055__), .dout(new_new_n4837__));
  or1   g2023(.dina(new_new_n7284__), .dinb(new_new_n4054__), .dout(new_new_n4838__));
  and1  g2024(.dina(new_new_n4079__), .dinb(new_new_n4080__), .dout(new_new_n4839__));
  or1   g2025(.dina(new_new_n7285__), .dinb(new_new_n4081__), .dout(new_new_n4840__));
  and1  g2026(.dina(new_new_n7287__), .dinb(new_new_n7288__), .dout(new_new_n4841__));
  or1   g2027(.dina(new_new_n7289__), .dinb(new_new_n4089__), .dout(new_new_n4842__));
  and1  g2028(.dina(new_new_n7291__), .dinb(new_new_n7293__), .dout(new_new_n4843__));
  or1   g2029(.dina(new_new_n7294__), .dinb(new_new_n7295__), .dout(new_new_n4844__));
  and1  g2030(.dina(new_new_n7299__), .dinb(new_new_n3560__), .dout(new_new_n4845__));
  and1  g2031(.dina(new_new_n7310__), .dinb(new_new_n3561__), .dout(new_new_n4846__));
  or1   g2032(.dina(new_new_n4845__), .dinb(new_new_n4846__), .dout(new_new_n4847__));
  and1  g2033(.dina(new_new_n7319__), .dinb(new_new_n7322__), .dout(new_new_n4848__));
  or1   g2034(.dina(new_new_n7325__), .dinb(new_new_n7328__), .dout(new_new_n4849__));
  and1  g2035(.dina(new_new_n7325__), .dinb(new_new_n4058__), .dout(new_new_n4850__));
  or1   g2036(.dina(new_new_n7319__), .dinb(new_new_n4059__), .dout(new_new_n4851__));
  and1  g2037(.dina(new_new_n4849__), .dinb(new_new_n4851__), .dout(new_new_n4852__));
  or1   g2038(.dina(new_new_n4848__), .dinb(new_new_n4850__), .dout(new_new_n4853__));
  and1  g2039(.dina(new_new_n3765__), .dinb(new_new_n7330__), .dout(new_new_n4854__));
  or1   g2040(.dina(new_new_n7331__), .dinb(new_new_n3949__), .dout(new_new_n4855__));
  and1  g2041(.dina(new_new_n4026__), .dinb(new_new_n7333__), .dout(new_new_n4856__));
  or1   g2042(.dina(new_new_n4027__), .dinb(new_new_n7336__), .dout(new_new_n4857__));
  and1  g2043(.dina(new_new_n7337__), .dinb(new_new_n4857__), .dout(new_new_n4858__));
  or1   g2044(.dina(new_new_n7338__), .dinb(new_new_n4856__), .dout(new_new_n4859__));
  and1  g2045(.dina(new_new_n7340__), .dinb(new_new_n7342__), .dout(new_new_n4860__));
  or1   g2046(.dina(new_new_n7344__), .dinb(new_new_n7345__), .dout(new_new_n4861__));
  and1  g2047(.dina(new_new_n7280__), .dinb(new_new_n4861__), .dout(new_new_n4862__));
  or1   g2048(.dina(new_new_n7282__), .dinb(new_new_n4860__), .dout(new_new_n4863__));
  and1  g2049(.dina(new_new_n7348__), .dinb(new_new_n7351__), .dout(new_new_n4864__));
  or1   g2050(.dina(new_new_n7353__), .dinb(new_new_n7355__), .dout(new_new_n4865__));
  and1  g2051(.dina(new_new_n7353__), .dinb(new_new_n7355__), .dout(new_new_n4866__));
  or1   g2052(.dina(new_new_n7348__), .dinb(new_new_n7351__), .dout(new_new_n4867__));
  and1  g2053(.dina(new_new_n7356__), .dinb(new_new_n4867__), .dout(new_new_n4868__));
  or1   g2054(.dina(new_new_n7357__), .dinb(new_new_n4866__), .dout(new_new_n4869__));
  and1  g2055(.dina(new_new_n4127__), .dinb(new_new_n4129__), .dout(new_new_n4870__));
  or1   g2056(.dina(new_new_n4126__), .dinb(new_new_n4128__), .dout(new_new_n4871__));
  and1  g2057(.dina(new_new_n4131__), .dinb(new_new_n4133__), .dout(new_new_n4872__));
  or1   g2058(.dina(new_new_n4130__), .dinb(new_new_n4132__), .dout(new_new_n4873__));
  and1  g2059(.dina(new_new_n4135__), .dinb(new_new_n4137__), .dout(new_new_n4874__));
  or1   g2060(.dina(new_new_n4134__), .dinb(new_new_n4136__), .dout(new_new_n4875__));
  or1   g2061(.dina(new_new_n3546__), .dinb(new_new_n7358__), .dout(new_new_n4876__));
  and1  g2062(.dina(new_new_n7359__), .dinb(new_new_n7360__), .dout(new_new_n4877__));
  and1  g2063(.dina(new_new_n7362__), .dinb(new_new_n7365__), .dout(new_new_n4878__));
  or1   g2064(.dina(new_new_n7367__), .dinb(new_new_n7368__), .dout(new_new_n4879__));
  and1  g2065(.dina(new_new_n2558__), .dinb(new_new_n7370__), .dout(new_new_n4880__));
  and1  g2066(.dina(new_new_n2559__), .dinb(new_new_n3591__), .dout(new_new_n4881__));
  or1   g2067(.dina(new_new_n4880__), .dinb(new_new_n4881__), .dout(new_new_n4882__));
  and1  g2068(.dina(new_new_n7299__), .dinb(new_new_n7372__), .dout(new_new_n4883__));
  and1  g2069(.dina(new_new_n7377__), .dinb(new_new_n7385__), .dout(new_new_n4884__));
  or1   g2070(.dina(new_new_n4883__), .dinb(new_new_n4884__), .dout(new_new_n4885__));
  and1  g2071(.dina(new_new_n3558__), .dinb(new_new_n4885__), .dout(new_new_n4886__));
  and1  g2072(.dina(new_new_n7390__), .dinb(new_new_n7385__), .dout(new_new_n4887__));
  and1  g2073(.dina(new_new_n7310__), .dinb(new_new_n7372__), .dout(new_new_n4888__));
  or1   g2074(.dina(new_new_n4887__), .dinb(new_new_n4888__), .dout(new_new_n4889__));
  and1  g2075(.dina(new_new_n3559__), .dinb(new_new_n4889__), .dout(new_new_n4890__));
  or1   g2076(.dina(new_new_n4886__), .dinb(new_new_n4890__), .dout(new_new_n4891__));
  and1  g2077(.dina(new_new_n7300__), .dinb(new_new_n7398__), .dout(new_new_n4892__));
  and1  g2078(.dina(new_new_n7377__), .dinb(new_new_n7400__), .dout(new_new_n4893__));
  or1   g2079(.dina(new_new_n4892__), .dinb(new_new_n4893__), .dout(new_new_n4894__));
  and1  g2080(.dina(new_new_n3484__), .dinb(new_new_n4894__), .dout(new_new_n4895__));
  and1  g2081(.dina(new_new_n7390__), .dinb(new_new_n7400__), .dout(new_new_n4896__));
  and1  g2082(.dina(new_new_n7311__), .dinb(new_new_n7398__), .dout(new_new_n4897__));
  or1   g2083(.dina(new_new_n4896__), .dinb(new_new_n4897__), .dout(new_new_n4898__));
  and1  g2084(.dina(new_new_n3485__), .dinb(new_new_n4898__), .dout(new_new_n4899__));
  or1   g2085(.dina(new_new_n4895__), .dinb(new_new_n4899__), .dout(new_new_n4900__));
  and1  g2086(.dina(new_new_n7300__), .dinb(new_new_n7402__), .dout(new_new_n4901__));
  and1  g2087(.dina(new_new_n7378__), .dinb(new_new_n7404__), .dout(new_new_n4902__));
  or1   g2088(.dina(new_new_n4901__), .dinb(new_new_n4902__), .dout(new_new_n4903__));
  and1  g2089(.dina(new_new_n3612__), .dinb(new_new_n4903__), .dout(new_new_n4904__));
  and1  g2090(.dina(new_new_n7391__), .dinb(new_new_n7404__), .dout(new_new_n4905__));
  and1  g2091(.dina(new_new_n7311__), .dinb(new_new_n7402__), .dout(new_new_n4906__));
  or1   g2092(.dina(new_new_n4905__), .dinb(new_new_n4906__), .dout(new_new_n4907__));
  and1  g2093(.dina(new_new_n3613__), .dinb(new_new_n4907__), .dout(new_new_n4908__));
  or1   g2094(.dina(new_new_n4904__), .dinb(new_new_n4908__), .dout(new_new_n4909__));
  and1  g2095(.dina(new_new_n7407__), .dinb(new_new_n7410__), .dout(new_new_n4910__));
  or1   g2096(.dina(new_new_n7412__), .dinb(new_new_n7414__), .dout(new_new_n4911__));
  and1  g2097(.dina(new_new_n7412__), .dinb(new_new_n7414__), .dout(new_new_n4912__));
  or1   g2098(.dina(new_new_n7407__), .dinb(new_new_n7410__), .dout(new_new_n4913__));
  and1  g2099(.dina(new_new_n4911__), .dinb(new_new_n4913__), .dout(new_new_n4914__));
  or1   g2100(.dina(new_new_n7415__), .dinb(new_new_n4912__), .dout(new_new_n4915__));
  and1  g2101(.dina(new_new_n7419__), .dinb(new_new_n7425__), .dout(new_new_n4916__));
  or1   g2102(.dina(new_new_n7429__), .dinb(new_new_n4117__), .dout(new_new_n4917__));
  and1  g2103(.dina(new_new_n7429__), .dinb(new_new_n4118__), .dout(new_new_n4918__));
  or1   g2104(.dina(new_new_n7419__), .dinb(new_new_n4119__), .dout(new_new_n4919__));
  and1  g2105(.dina(new_new_n4917__), .dinb(new_new_n4919__), .dout(new_new_n4920__));
  or1   g2106(.dina(new_new_n4916__), .dinb(new_new_n4918__), .dout(new_new_n4921__));
  and1  g2107(.dina(new_new_n7435__), .dinb(new_new_n7437__), .dout(new_new_n4922__));
  or1   g2108(.dina(new_new_n4113__), .dinb(new_new_n4872__), .dout(new_new_n4923__));
  or1   g2109(.dina(new_new_n7435__), .dinb(new_new_n7437__), .dout(new_new_n4924__));
  and1  g2110(.dina(new_new_n7439__), .dinb(new_new_n7441__), .dout(new_new_n4925__));
  or1   g2111(.dina(new_new_n4115__), .dinb(new_new_n4870__), .dout(new_new_n4926__));
  and1  g2112(.dina(new_new_n7442__), .dinb(new_new_n7446__), .dout(new_new_n4927__));
  or1   g2113(.dina(new_new_n4121__), .dinb(new_new_n7457__), .dout(new_new_n4928__));
  and1  g2114(.dina(new_new_n4122__), .dinb(new_new_n7457__), .dout(new_new_n4929__));
  or1   g2115(.dina(new_new_n4123__), .dinb(new_new_n7446__), .dout(new_new_n4930__));
  and1  g2116(.dina(new_new_n4928__), .dinb(new_new_n4930__), .dout(new_new_n4931__));
  or1   g2117(.dina(new_new_n4927__), .dinb(new_new_n4929__), .dout(new_new_n4932__));
  or1   g2118(.dina(new_new_n7362__), .dinb(new_new_n7365__), .dout(new_new_n4933__));
  and1  g2119(.dina(new_new_n7333__), .dinb(new_new_n7464__), .dout(new_new_n4934__));
  or1   g2120(.dina(new_new_n7336__), .dinb(new_new_n4842__), .dout(new_new_n4935__));
  and1  g2121(.dina(new_new_n7338__), .dinb(new_new_n7287__), .dout(new_new_n4936__));
  or1   g2122(.dina(new_new_n7337__), .dinb(new_new_n7289__), .dout(new_new_n4937__));
  and1  g2123(.dina(new_new_n3991__), .dinb(new_new_n4937__), .dout(new_new_n4938__));
  or1   g2124(.dina(new_new_n3990__), .dinb(new_new_n4936__), .dout(new_new_n4939__));
  and1  g2125(.dina(new_new_n4935__), .dinb(new_new_n4938__), .dout(new_new_n4940__));
  or1   g2126(.dina(new_new_n4934__), .dinb(new_new_n4939__), .dout(new_new_n4941__));
  and1  g2127(.dina(new_new_n7466__), .dinb(new_new_n7467__), .dout(new_new_n4942__));
  or1   g2128(.dina(new_new_n7468__), .dinb(new_new_n7469__), .dout(new_new_n4943__));
  and1  g2129(.dina(new_new_n7356__), .dinb(new_new_n7470__), .dout(new_new_n4944__));
  or1   g2130(.dina(new_new_n7357__), .dinb(new_new_n7471__), .dout(new_new_n4945__));
  and1  g2131(.dina(new_new_n7420__), .dinb(new_new_n7472__), .dout(new_new_n4946__));
  or1   g2132(.dina(new_new_n7428__), .dinb(new_new_n4099__), .dout(new_new_n4947__));
  and1  g2133(.dina(new_new_n7430__), .dinb(new_new_n4100__), .dout(new_new_n4948__));
  or1   g2134(.dina(new_new_n7420__), .dinb(new_new_n4101__), .dout(new_new_n4949__));
  and1  g2135(.dina(new_new_n4947__), .dinb(new_new_n4949__), .dout(new_new_n4950__));
  or1   g2136(.dina(new_new_n4946__), .dinb(new_new_n4948__), .dout(new_new_n4951__));
  and1  g2137(.dina(new_new_n7421__), .dinb(new_new_n7473__), .dout(new_new_n4952__));
  or1   g2138(.dina(new_new_n7430__), .dinb(new_new_n4103__), .dout(new_new_n4953__));
  and1  g2139(.dina(new_new_n7432__), .dinb(new_new_n4104__), .dout(new_new_n4954__));
  or1   g2140(.dina(new_new_n7421__), .dinb(new_new_n4105__), .dout(new_new_n4955__));
  and1  g2141(.dina(new_new_n4953__), .dinb(new_new_n4955__), .dout(new_new_n4956__));
  or1   g2142(.dina(new_new_n4952__), .dinb(new_new_n4954__), .dout(new_new_n4957__));
  and1  g2143(.dina(new_new_n4047__), .dinb(new_new_n4068__), .dout(new_new_n4958__));
  or1   g2144(.dina(new_new_n4046__), .dinb(new_new_n4069__), .dout(new_new_n4959__));
  and1  g2145(.dina(new_new_n7475__), .dinb(new_new_n7476__), .dout(new_new_n4960__));
  or1   g2146(.dina(new_new_n7478__), .dinb(new_new_n7480__), .dout(new_new_n4961__));
  and1  g2147(.dina(new_new_n7478__), .dinb(new_new_n7480__), .dout(new_new_n4962__));
  or1   g2148(.dina(new_new_n7475__), .dinb(new_new_n7476__), .dout(new_new_n4963__));
  and1  g2149(.dina(new_new_n4961__), .dinb(new_new_n4963__), .dout(new_new_n4964__));
  or1   g2150(.dina(new_new_n4960__), .dinb(new_new_n4962__), .dout(new_new_n4965__));
  and1  g2151(.dina(new_new_n4855__), .dinb(new_new_n4964__), .dout(new_new_n4966__));
  and1  g2152(.dina(new_new_n7482__), .dinb(new_new_n4965__), .dout(new_new_n4967__));
  or1   g2153(.dina(new_new_n7483__), .dinb(new_new_n4967__), .dout(new_new_n4968__));
  and1  g2154(.dina(new_new_n7484__), .dinb(new_new_n7447__), .dout(new_new_n4969__));
  and1  g2155(.dina(new_new_n4108__), .dinb(new_new_n7458__), .dout(new_new_n4970__));
  or1   g2156(.dina(new_new_n4969__), .dinb(new_new_n4970__), .dout(new_new_n4971__));
  and1  g2157(.dina(new_new_n7468__), .dinb(new_new_n7469__), .dout(new_new_n4972__));
  or1   g2158(.dina(new_new_n7466__), .dinb(new_new_n7467__), .dout(new_new_n4973__));
  and1  g2159(.dina(new_new_n7470__), .dinb(new_new_n4973__), .dout(new_new_n4974__));
  or1   g2160(.dina(new_new_n7471__), .dinb(new_new_n4972__), .dout(new_new_n4975__));
  and1  g2161(.dina(new_new_n7486__), .dinb(new_new_n7488__), .dout(new_new_n4976__));
  or1   g2162(.dina(new_new_n4095__), .dinb(new_new_n4920__), .dout(new_new_n4977__));
  and1  g2163(.dina(new_new_n7490__), .dinb(new_new_n7492__), .dout(new_new_n4978__));
  or1   g2164(.dina(new_new_n4111__), .dinb(new_new_n4874__), .dout(new_new_n4979__));
  or1   g2165(.dina(new_new_n7490__), .dinb(new_new_n7492__), .dout(new_new_n4980__));
  and1  g2166(.dina(new_new_n4979__), .dinb(new_new_n4980__), .dout(new_new_n4981__));
  and1  g2167(.dina(new_new_n4923__), .dinb(new_new_n7494__), .dout(new_new_n4982__));
  or1   g2168(.dina(new_new_n7439__), .dinb(new_new_n7441__), .dout(new_new_n4983__));
  and1  g2169(.dina(new_new_n4926__), .dinb(new_new_n4983__), .dout(new_new_n4984__));
  and1  g2170(.dina(new_new_n7496__), .dinb(new_new_n7447__), .dout(new_new_n4985__));
  or1   g2171(.dina(new_new_n4091__), .dinb(new_new_n7458__), .dout(new_new_n4986__));
  and1  g2172(.dina(new_new_n7497__), .dinb(new_new_n7460__), .dout(new_new_n4987__));
  or1   g2173(.dina(new_new_n4093__), .dinb(new_new_n7449__), .dout(new_new_n4988__));
  and1  g2174(.dina(new_new_n4986__), .dinb(new_new_n4988__), .dout(new_new_n4989__));
  or1   g2175(.dina(new_new_n4985__), .dinb(new_new_n4987__), .dout(new_new_n4990__));
  and1  g2176(.dina(new_new_n7499__), .dinb(new_new_n7501__), .dout(new_new_n4991__));
  or1   g2177(.dina(new_new_n3175__), .dinb(new_new_n4956__), .dout(new_new_n4992__));
  and1  g2178(.dina(new_new_n7503__), .dinb(new_new_n7505__), .dout(new_new_n4993__));
  or1   g2179(.dina(new_new_n3183__), .dinb(new_new_n4950__), .dout(new_new_n4994__));
  and1  g2180(.dina(new_new_n7507__), .dinb(new_new_n7509__), .dout(new_new_n4995__));
  and1  g2181(.dina(new_new_n7511__), .dinb(new_new_n7513__), .dout(new_new_n4996__));
  or1   g2182(.dina(new_new_n4097__), .dinb(new_new_n4931__), .dout(new_new_n4997__));
  or1   g2183(.dina(new_new_n7511__), .dinb(new_new_n7513__), .dout(new_new_n4998__));
  and1  g2184(.dina(new_new_n4997__), .dinb(new_new_n7514__), .dout(new_new_n4999__));
  and1  g2185(.dina(new_new_n7515__), .dinb(new_new_n7517__), .dout(new_new_n5000__));
  and1  g2186(.dina(new_new_n2544__), .dinb(new_new_n7521__), .dout(new_new_n5001__));
  and1  g2187(.dina(new_new_n2738__), .dinb(new_new_n7521__), .dout(new_new_n5002__));
  and1  g2188(.dina(new_new_n2758__), .dinb(new_new_n7522__), .dout(new_new_n5003__));
  or1   g2189(.dina(new_new_n2764__), .dinb(new_new_n7531__), .dout(new_new_n5004__));
  or1   g2190(.dina(new_new_n2778__), .dinb(new_new_n7531__), .dout(new_new_n5005__));
  and1  g2191(.dina(new_new_n2792__), .dinb(new_new_n7522__), .dout(new_new_n5006__));
  and1  g2192(.dina(new_new_n2830__), .dinb(new_new_n7524__), .dout(new_new_n5007__));
  or1   g2193(.dina(new_new_n2836__), .dinb(new_new_n7532__), .dout(new_new_n5008__));
  or1   g2194(.dina(new_new_n2848__), .dinb(new_new_n7532__), .dout(new_new_n5009__));
  and1  g2195(.dina(new_new_n7302__), .dinb(new_new_n7542__), .dout(new_new_n5010__));
  and1  g2196(.dina(new_new_n7378__), .dinb(new_new_n7544__), .dout(new_new_n5011__));
  or1   g2197(.dina(new_new_n5010__), .dinb(new_new_n5011__), .dout(new_new_n5012__));
  and1  g2198(.dina(new_new_n3482__), .dinb(new_new_n5012__), .dout(new_new_n5013__));
  and1  g2199(.dina(new_new_n7391__), .dinb(new_new_n7544__), .dout(new_new_n5014__));
  and1  g2200(.dina(new_new_n7313__), .dinb(new_new_n7542__), .dout(new_new_n5015__));
  or1   g2201(.dina(new_new_n5014__), .dinb(new_new_n5015__), .dout(new_new_n5016__));
  and1  g2202(.dina(new_new_n3483__), .dinb(new_new_n5016__), .dout(new_new_n5017__));
  and1  g2203(.dina(new_new_n7546__), .dinb(new_new_n7534__), .dout(new_new_n5018__));
  or1   g2204(.dina(new_new_n7547__), .dinb(new_new_n7534__), .dout(new_new_n5019__));
  and1  g2205(.dina(new_new_n7549__), .dinb(new_new_n5019__), .dout(new_new_n5020__));
  and1  g2206(.dina(new_new_n7550__), .dinb(new_new_n3609__), .dout(new_new_n5021__));
  or1   g2207(.dina(new_new_n7551__), .dinb(new_new_n7553__), .dout(new_new_n5022__));
  and1  g2208(.dina(new_new_n3629__), .dinb(new_new_n5022__), .dout(new_new_n5023__));
  or1   g2209(.dina(new_new_n7554__), .dinb(new_new_n5021__), .dout(new_new_n5024__));
  and1  g2210(.dina(new_new_n7555__), .dinb(new_new_n7556__), .dout(new_new_n5025__));
  or1   g2211(.dina(new_new_n7557__), .dinb(new_new_n7558__), .dout(new_new_n5026__));
  and1  g2212(.dina(new_new_n7557__), .dinb(new_new_n7558__), .dout(new_new_n5027__));
  or1   g2213(.dina(new_new_n7555__), .dinb(new_new_n7556__), .dout(new_new_n5028__));
  and1  g2214(.dina(new_new_n5026__), .dinb(new_new_n5028__), .dout(new_new_n5029__));
  or1   g2215(.dina(new_new_n5025__), .dinb(new_new_n5027__), .dout(new_new_n5030__));
  and1  g2216(.dina(new_new_n7559__), .dinb(new_new_n7560__), .dout(new_new_n5031__));
  or1   g2217(.dina(new_new_n7561__), .dinb(new_new_n7562__), .dout(new_new_n5032__));
  and1  g2218(.dina(new_new_n7561__), .dinb(new_new_n7562__), .dout(new_new_n5033__));
  or1   g2219(.dina(new_new_n7559__), .dinb(new_new_n7560__), .dout(new_new_n5034__));
  and1  g2220(.dina(new_new_n5032__), .dinb(new_new_n5034__), .dout(new_new_n5035__));
  or1   g2221(.dina(new_new_n5031__), .dinb(new_new_n5033__), .dout(new_new_n5036__));
  and1  g2222(.dina(new_new_n7563__), .dinb(new_new_n3734__), .dout(new_new_n5037__));
  or1   g2223(.dina(new_new_n7272__), .dinb(new_new_n3735__), .dout(new_new_n5038__));
  and1  g2224(.dina(new_new_n7271__), .dinb(new_new_n4015__), .dout(new_new_n5039__));
  or1   g2225(.dina(new_new_n7563__), .dinb(new_new_n4014__), .dout(new_new_n5040__));
  and1  g2226(.dina(new_new_n5038__), .dinb(new_new_n5040__), .dout(new_new_n5041__));
  or1   g2227(.dina(new_new_n5037__), .dinb(new_new_n5039__), .dout(new_new_n5042__));
  and1  g2228(.dina(new_new_n7565__), .dinb(new_new_n7566__), .dout(new_new_n5043__));
  or1   g2229(.dina(new_new_n7568__), .dinb(new_new_n7569__), .dout(new_new_n5044__));
  and1  g2230(.dina(new_new_n7568__), .dinb(new_new_n7569__), .dout(new_new_n5045__));
  or1   g2231(.dina(new_new_n7565__), .dinb(new_new_n7566__), .dout(new_new_n5046__));
  and1  g2232(.dina(new_new_n5044__), .dinb(new_new_n5046__), .dout(new_new_n5047__));
  or1   g2233(.dina(new_new_n5043__), .dinb(new_new_n5045__), .dout(new_new_n5048__));
  and1  g2234(.dina(new_new_n5036__), .dinb(new_new_n5047__), .dout(new_new_n5049__));
  and1  g2235(.dina(new_new_n5035__), .dinb(new_new_n5048__), .dout(new_new_n5050__));
  or1   g2236(.dina(new_new_n5049__), .dinb(new_new_n5050__), .dout(new_new_n5051__));
  and1  g2237(.dina(new_new_n7546__), .dinb(new_new_n5051__), .dout(new_new_n5052__));
  or1   g2238(.dina(new_new_n7524__), .dinb(new_new_n7570__), .dout(new_new_n5053__));
  or1   g2239(.dina(new_new_n7523__), .dinb(new_new_n7571__), .dout(new_new_n5054__));
  and1  g2240(.dina(new_new_n7535__), .dinb(new_new_n3923__), .dout(new_new_n5055__));
  and1  g2241(.dina(new_new_n7535__), .dinb(new_new_n3920__), .dout(new_new_n5056__));
  and1  g2242(.dina(new_new_n7538__), .dinb(new_new_n3915__), .dout(new_new_n5057__));
  or1   g2243(.dina(new_new_n7526__), .dinb(new_new_n7572__), .dout(new_new_n5058__));
  and1  g2244(.dina(new_new_n4011__), .dinb(new_new_n4013__), .dout(new_new_n5059__));
  or1   g2245(.dina(new_new_n4010__), .dinb(new_new_n4012__), .dout(new_new_n5060__));
  and1  g2246(.dina(new_new_n4007__), .dinb(new_new_n4009__), .dout(new_new_n5061__));
  or1   g2247(.dina(new_new_n4006__), .dinb(new_new_n4008__), .dout(new_new_n5062__));
  and1  g2248(.dina(new_new_n7573__), .dinb(new_new_n7574__), .dout(new_new_n5063__));
  or1   g2249(.dina(new_new_n7575__), .dinb(new_new_n7576__), .dout(new_new_n5064__));
  and1  g2250(.dina(new_new_n7575__), .dinb(new_new_n7576__), .dout(new_new_n5065__));
  or1   g2251(.dina(new_new_n7573__), .dinb(new_new_n7574__), .dout(new_new_n5066__));
  and1  g2252(.dina(new_new_n5064__), .dinb(new_new_n5066__), .dout(new_new_n5067__));
  or1   g2253(.dina(new_new_n5063__), .dinb(new_new_n5065__), .dout(new_new_n5068__));
  and1  g2254(.dina(new_new_n4003__), .dinb(new_new_n4004__), .dout(new_new_n5069__));
  or1   g2255(.dina(new_new_n7577__), .dinb(new_new_n4005__), .dout(new_new_n5070__));
  and1  g2256(.dina(new_new_n3999__), .dinb(new_new_n4001__), .dout(new_new_n5071__));
  or1   g2257(.dina(new_new_n7578__), .dinb(new_new_n4000__), .dout(new_new_n5072__));
  and1  g2258(.dina(new_new_n7579__), .dinb(new_new_n7580__), .dout(new_new_n5073__));
  or1   g2259(.dina(new_new_n7581__), .dinb(new_new_n7582__), .dout(new_new_n5074__));
  and1  g2260(.dina(new_new_n7581__), .dinb(new_new_n7582__), .dout(new_new_n5075__));
  or1   g2261(.dina(new_new_n7579__), .dinb(new_new_n7580__), .dout(new_new_n5076__));
  and1  g2262(.dina(new_new_n5074__), .dinb(new_new_n5076__), .dout(new_new_n5077__));
  or1   g2263(.dina(new_new_n5073__), .dinb(new_new_n5075__), .dout(new_new_n5078__));
  and1  g2264(.dina(new_new_n5067__), .dinb(new_new_n5077__), .dout(new_new_n5079__));
  and1  g2265(.dina(new_new_n5068__), .dinb(new_new_n5078__), .dout(new_new_n5080__));
  or1   g2266(.dina(new_new_n7545__), .dinb(new_new_n5080__), .dout(new_new_n5081__));
  or1   g2267(.dina(new_new_n5079__), .dinb(new_new_n5081__), .dout(new_new_n5082__));
  and1  g2268(.dina(new_new_n7538__), .dinb(new_new_n5082__), .dout(new_new_n5083__));
  and1  g2269(.dina(new_new_n3509__), .dinb(new_new_n3528__), .dout(new_new_n5084__));
  and1  g2270(.dina(new_new_n3508__), .dinb(new_new_n3529__), .dout(new_new_n5085__));
  and1  g2271(.dina(new_new_n7276__), .dinb(new_new_n7584__), .dout(new_new_n5086__));
  or1   g2272(.dina(new_new_n7586__), .dinb(new_new_n7588__), .dout(new_new_n5087__));
  and1  g2273(.dina(new_new_n7590__), .dinb(new_new_n5087__), .dout(new_new_n5088__));
  or1   g2274(.dina(new_new_n7594__), .dinb(new_new_n5086__), .dout(new_new_n5089__));
  and1  g2275(.dina(new_new_n3533__), .dinb(new_new_n7598__), .dout(new_new_n5090__));
  and1  g2276(.dina(new_new_n3532__), .dinb(new_new_n7602__), .dout(new_new_n5091__));
  and1  g2277(.dina(new_new_n3580__), .dinb(new_new_n7604__), .dout(new_new_n5092__));
  and1  g2278(.dina(new_new_n3551__), .dinb(new_new_n7606__), .dout(new_new_n5093__));
  or1   g2279(.dina(new_new_n5092__), .dinb(new_new_n5093__), .dout(new_new_n5094__));
  or1   g2280(.dina(new_new_n7273__), .dinb(new_new_n7607__), .dout(new_new_n5095__));
  and1  g2281(.dina(new_new_n7273__), .dinb(new_new_n7607__), .dout(new_new_n5096__));
  or1   g2282(.dina(new_new_n7278__), .dinb(new_new_n7279__), .dout(new_new_n5097__));
  or1   g2283(.dina(new_new_n3586__), .dinb(new_new_n7608__), .dout(new_new_n5098__));
  and1  g2284(.dina(new_new_n7610__), .dinb(new_new_n3474__), .dout(new_new_n5099__));
  and1  g2285(.dina(new_new_n3154__), .dinb(new_new_n3475__), .dout(new_new_n5100__));
  or1   g2286(.dina(new_new_n5099__), .dinb(new_new_n5100__), .dout(new_new_n5101__));
  or1   g2287(.dina(new_new_n7370__), .dinb(new_new_n7611__), .dout(new_new_n5102__));
  and1  g2288(.dina(new_new_n7369__), .dinb(new_new_n7611__), .dout(new_new_n5103__));
  or1   g2289(.dina(new_new_n7359__), .dinb(new_new_n7360__), .dout(new_new_n5104__));
  and1  g2290(.dina(new_new_n7553__), .dinb(new_new_n7612__), .dout(new_new_n5105__));
  or1   g2291(.dina(new_new_n7552__), .dinb(new_new_n7612__), .dout(new_new_n5106__));
  or1   g2292(.dina(new_new_n7606__), .dinb(new_new_n7613__), .dout(new_new_n5107__));
  and1  g2293(.dina(new_new_n3585__), .dinb(new_new_n5107__), .dout(new_new_n5108__));
  and1  g2294(.dina(new_new_n7263__), .dinb(new_new_n7614__), .dout(new_new_n5109__));
  or1   g2295(.dina(new_new_n7263__), .dinb(new_new_n7614__), .dout(new_new_n5110__));
  or1   g2296(.dina(new_new_n7567__), .dinb(new_new_n7615__), .dout(new_new_n5111__));
  and1  g2297(.dina(new_new_n7277__), .dinb(new_new_n7616__), .dout(new_new_n5112__));
  or1   g2298(.dina(new_new_n7586__), .dinb(new_new_n3583__), .dout(new_new_n5113__));
  or1   g2299(.dina(new_new_n7277__), .dinb(new_new_n7616__), .dout(new_new_n5114__));
  and1  g2300(.dina(new_new_n7617__), .dinb(new_new_n5114__), .dout(new_new_n5115__));
  and1  g2301(.dina(new_new_n3127__), .dinb(new_new_n7460__), .dout(new_new_n5116__));
  or1   g2302(.dina(new_new_n7618__), .dinb(new_new_n7449__), .dout(new_new_n5117__));
  and1  g2303(.dina(new_new_n2732__), .dinb(new_new_n7526__), .dout(new_new_n5118__));
  and1  g2304(.dina(new_new_n7539__), .dinb(new_new_n3917__), .dout(new_new_n5119__));
  or1   g2305(.dina(new_new_n5118__), .dinb(new_new_n5119__), .dout(new_new_n5120__));
  and1  g2306(.dina(new_new_n2752__), .dinb(new_new_n7527__), .dout(new_new_n5121__));
  and1  g2307(.dina(new_new_n7539__), .dinb(new_new_n7620__), .dout(new_new_n5122__));
  or1   g2308(.dina(new_new_n5121__), .dinb(new_new_n5122__), .dout(new_new_n5123__));
  or1   g2309(.dina(new_new_n2843__), .dinb(new_new_n7540__), .dout(new_new_n5124__));
  or1   g2310(.dina(new_new_n7527__), .dinb(new_new_n7621__), .dout(new_new_n5125__));
  and1  g2311(.dina(new_new_n5124__), .dinb(new_new_n5125__), .dout(new_new_n5126__));
  or1   g2312(.dina(new_new_n7623__), .dinb(new_new_n3536__), .dout(new_new_n5127__));
  or1   g2313(.dina(new_new_n7625__), .dinb(new_new_n3537__), .dout(new_new_n5128__));
  and1  g2314(.dina(new_new_n5127__), .dinb(new_new_n5128__), .dout(new_new_n5129__));
  and1  g2315(.dina(new_new_n7627__), .dinb(new_new_n7397__), .dout(new_new_n5130__));
  and1  g2316(.dina(new_new_n7629__), .dinb(new_new_n7399__), .dout(new_new_n5131__));
  or1   g2317(.dina(new_new_n5130__), .dinb(new_new_n5131__), .dout(new_new_n5132__));
  and1  g2318(.dina(new_new_n7541__), .dinb(new_new_n7631__), .dout(new_new_n5133__));
  and1  g2319(.dina(new_new_n7543__), .dinb(new_new_n7633__), .dout(new_new_n5134__));
  or1   g2320(.dina(new_new_n5133__), .dinb(new_new_n5134__), .dout(new_new_n5135__));
  and1  g2321(.dina(new_new_n7302__), .dinb(new_new_n7635__), .dout(new_new_n5136__));
  and1  g2322(.dina(new_new_n7380__), .dinb(new_new_n7638__), .dout(new_new_n5137__));
  or1   g2323(.dina(new_new_n5136__), .dinb(new_new_n5137__), .dout(new_new_n5138__));
  and1  g2324(.dina(new_new_n3500__), .dinb(new_new_n5138__), .dout(new_new_n5139__));
  and1  g2325(.dina(new_new_n7393__), .dinb(new_new_n7638__), .dout(new_new_n5140__));
  and1  g2326(.dina(new_new_n7313__), .dinb(new_new_n7635__), .dout(new_new_n5141__));
  or1   g2327(.dina(new_new_n5140__), .dinb(new_new_n5141__), .dout(new_new_n5142__));
  and1  g2328(.dina(new_new_n3501__), .dinb(new_new_n5142__), .dout(new_new_n5143__));
  or1   g2329(.dina(new_new_n5139__), .dinb(new_new_n5143__), .dout(new_new_n5144__));
  and1  g2330(.dina(new_new_n7303__), .dinb(new_new_n7633__), .dout(new_new_n5145__));
  and1  g2331(.dina(new_new_n7380__), .dinb(new_new_n7631__), .dout(new_new_n5146__));
  or1   g2332(.dina(new_new_n5145__), .dinb(new_new_n5146__), .dout(new_new_n5147__));
  and1  g2333(.dina(new_new_n3516__), .dinb(new_new_n5147__), .dout(new_new_n5148__));
  and1  g2334(.dina(new_new_n7393__), .dinb(new_new_n7630__), .dout(new_new_n5149__));
  and1  g2335(.dina(new_new_n7314__), .dinb(new_new_n7632__), .dout(new_new_n5150__));
  or1   g2336(.dina(new_new_n5149__), .dinb(new_new_n5150__), .dout(new_new_n5151__));
  and1  g2337(.dina(new_new_n3517__), .dinb(new_new_n5151__), .dout(new_new_n5152__));
  or1   g2338(.dina(new_new_n5148__), .dinb(new_new_n5152__), .dout(new_new_n5153__));
  and1  g2339(.dina(new_new_n7303__), .dinb(new_new_n7641__), .dout(new_new_n5154__));
  and1  g2340(.dina(new_new_n7379__), .dinb(new_new_n7644__), .dout(new_new_n5155__));
  or1   g2341(.dina(new_new_n5154__), .dinb(new_new_n5155__), .dout(new_new_n5156__));
  and1  g2342(.dina(new_new_n3630__), .dinb(new_new_n5156__), .dout(new_new_n5157__));
  and1  g2343(.dina(new_new_n7392__), .dinb(new_new_n7644__), .dout(new_new_n5158__));
  and1  g2344(.dina(new_new_n7314__), .dinb(new_new_n7641__), .dout(new_new_n5159__));
  or1   g2345(.dina(new_new_n5158__), .dinb(new_new_n5159__), .dout(new_new_n5160__));
  and1  g2346(.dina(new_new_n3631__), .dinb(new_new_n5160__), .dout(new_new_n5161__));
  or1   g2347(.dina(new_new_n5157__), .dinb(new_new_n5161__), .dout(new_new_n5162__));
  and1  g2348(.dina(new_new_n7305__), .dinb(new_new_n7625__), .dout(new_new_n5163__));
  and1  g2349(.dina(new_new_n7382__), .dinb(new_new_n7623__), .dout(new_new_n5164__));
  or1   g2350(.dina(new_new_n5163__), .dinb(new_new_n5164__), .dout(new_new_n5165__));
  and1  g2351(.dina(new_new_n3518__), .dinb(new_new_n5165__), .dout(new_new_n5166__));
  and1  g2352(.dina(new_new_n7395__), .dinb(new_new_n7622__), .dout(new_new_n5167__));
  and1  g2353(.dina(new_new_n7316__), .dinb(new_new_n7624__), .dout(new_new_n5168__));
  or1   g2354(.dina(new_new_n5167__), .dinb(new_new_n5168__), .dout(new_new_n5169__));
  and1  g2355(.dina(new_new_n3519__), .dinb(new_new_n5169__), .dout(new_new_n5170__));
  or1   g2356(.dina(new_new_n5166__), .dinb(new_new_n5170__), .dout(new_new_n5171__));
  and1  g2357(.dina(new_new_n7305__), .dinb(new_new_n7629__), .dout(new_new_n5172__));
  and1  g2358(.dina(new_new_n7382__), .dinb(new_new_n7627__), .dout(new_new_n5173__));
  or1   g2359(.dina(new_new_n5172__), .dinb(new_new_n5173__), .dout(new_new_n5174__));
  and1  g2360(.dina(new_new_n3486__), .dinb(new_new_n5174__), .dout(new_new_n5175__));
  and1  g2361(.dina(new_new_n7395__), .dinb(new_new_n7626__), .dout(new_new_n5176__));
  and1  g2362(.dina(new_new_n7316__), .dinb(new_new_n7628__), .dout(new_new_n5177__));
  or1   g2363(.dina(new_new_n5176__), .dinb(new_new_n5177__), .dout(new_new_n5178__));
  and1  g2364(.dina(new_new_n3487__), .dinb(new_new_n5178__), .dout(new_new_n5179__));
  or1   g2365(.dina(new_new_n5175__), .dinb(new_new_n5179__), .dout(new_new_n5180__));
  and1  g2366(.dina(new_new_n7306__), .dinb(new_new_n7647__), .dout(new_new_n5181__));
  and1  g2367(.dina(new_new_n7383__), .dinb(new_new_n7649__), .dout(new_new_n5182__));
  or1   g2368(.dina(new_new_n5181__), .dinb(new_new_n5182__), .dout(new_new_n5183__));
  and1  g2369(.dina(new_new_n3562__), .dinb(new_new_n5183__), .dout(new_new_n5184__));
  and1  g2370(.dina(new_new_n7396__), .dinb(new_new_n7649__), .dout(new_new_n5185__));
  and1  g2371(.dina(new_new_n7317__), .dinb(new_new_n7647__), .dout(new_new_n5186__));
  or1   g2372(.dina(new_new_n5185__), .dinb(new_new_n5186__), .dout(new_new_n5187__));
  and1  g2373(.dina(new_new_n3563__), .dinb(new_new_n5187__), .dout(new_new_n5188__));
  or1   g2374(.dina(new_new_n5184__), .dinb(new_new_n5188__), .dout(new_new_n5189__));
  and1  g2375(.dina(new_new_n7306__), .dinb(new_new_n7651__), .dout(new_new_n5190__));
  and1  g2376(.dina(new_new_n7383__), .dinb(new_new_n7653__), .dout(new_new_n5191__));
  or1   g2377(.dina(new_new_n5190__), .dinb(new_new_n5191__), .dout(new_new_n5192__));
  and1  g2378(.dina(new_new_n3544__), .dinb(new_new_n5192__), .dout(new_new_n5193__));
  and1  g2379(.dina(new_new_n7396__), .dinb(new_new_n7653__), .dout(new_new_n5194__));
  and1  g2380(.dina(new_new_n7317__), .dinb(new_new_n7651__), .dout(new_new_n5195__));
  or1   g2381(.dina(new_new_n5194__), .dinb(new_new_n5195__), .dout(new_new_n5196__));
  and1  g2382(.dina(new_new_n3545__), .dinb(new_new_n5196__), .dout(new_new_n5197__));
  or1   g2383(.dina(new_new_n5193__), .dinb(new_new_n5197__), .dout(new_new_n5198__));
  and1  g2384(.dina(new_new_n7654__), .dinb(new_new_n7655__), .dout(new_new_n5199__));
  or1   g2385(.dina(new_new_n7656__), .dinb(new_new_n7657__), .dout(new_new_n5200__));
  and1  g2386(.dina(new_new_n7656__), .dinb(new_new_n7657__), .dout(new_new_n5201__));
  or1   g2387(.dina(new_new_n7654__), .dinb(new_new_n7655__), .dout(new_new_n5202__));
  and1  g2388(.dina(new_new_n5200__), .dinb(new_new_n5202__), .dout(new_new_n5203__));
  or1   g2389(.dina(new_new_n5199__), .dinb(new_new_n5201__), .dout(new_new_n5204__));
  and1  g2390(.dina(new_new_n7658__), .dinb(new_new_n7620__), .dout(new_new_n5205__));
  or1   g2391(.dina(new_new_n7659__), .dinb(new_new_n7661__), .dout(new_new_n5206__));
  and1  g2392(.dina(new_new_n7659__), .dinb(new_new_n7661__), .dout(new_new_n5207__));
  or1   g2393(.dina(new_new_n7658__), .dinb(new_new_n7619__), .dout(new_new_n5208__));
  and1  g2394(.dina(new_new_n5206__), .dinb(new_new_n5208__), .dout(new_new_n5209__));
  or1   g2395(.dina(new_new_n5205__), .dinb(new_new_n5207__), .dout(new_new_n5210__));
  and1  g2396(.dina(new_new_n7662__), .dinb(new_new_n7663__), .dout(new_new_n5211__));
  or1   g2397(.dina(new_new_n7664__), .dinb(new_new_n7665__), .dout(new_new_n5212__));
  and1  g2398(.dina(new_new_n7664__), .dinb(new_new_n7665__), .dout(new_new_n5213__));
  or1   g2399(.dina(new_new_n7662__), .dinb(new_new_n7663__), .dout(new_new_n5214__));
  and1  g2400(.dina(new_new_n5212__), .dinb(new_new_n5214__), .dout(new_new_n5215__));
  or1   g2401(.dina(new_new_n5211__), .dinb(new_new_n5213__), .dout(new_new_n5216__));
  and1  g2402(.dina(new_new_n7666__), .dinb(new_new_n7667__), .dout(new_new_n5217__));
  or1   g2403(.dina(new_new_n7668__), .dinb(new_new_n7669__), .dout(new_new_n5218__));
  and1  g2404(.dina(new_new_n7668__), .dinb(new_new_n7669__), .dout(new_new_n5219__));
  or1   g2405(.dina(new_new_n7666__), .dinb(new_new_n7667__), .dout(new_new_n5220__));
  and1  g2406(.dina(new_new_n5218__), .dinb(new_new_n5220__), .dout(new_new_n5221__));
  or1   g2407(.dina(new_new_n5217__), .dinb(new_new_n5219__), .dout(new_new_n5222__));
  and1  g2408(.dina(new_new_n7670__), .dinb(new_new_n7671__), .dout(new_new_n5223__));
  or1   g2409(.dina(new_new_n7672__), .dinb(new_new_n7673__), .dout(new_new_n5224__));
  and1  g2410(.dina(new_new_n7672__), .dinb(new_new_n7673__), .dout(new_new_n5225__));
  or1   g2411(.dina(new_new_n7670__), .dinb(new_new_n7671__), .dout(new_new_n5226__));
  and1  g2412(.dina(new_new_n5224__), .dinb(new_new_n5226__), .dout(new_new_n5227__));
  or1   g2413(.dina(new_new_n5223__), .dinb(new_new_n5225__), .dout(new_new_n5228__));
  and1  g2414(.dina(new_new_n7674__), .dinb(new_new_n7675__), .dout(new_new_n5229__));
  or1   g2415(.dina(new_new_n7676__), .dinb(new_new_n7677__), .dout(new_new_n5230__));
  and1  g2416(.dina(new_new_n7676__), .dinb(new_new_n7677__), .dout(new_new_n5231__));
  or1   g2417(.dina(new_new_n7674__), .dinb(new_new_n7675__), .dout(new_new_n5232__));
  and1  g2418(.dina(new_new_n5230__), .dinb(new_new_n5232__), .dout(new_new_n5233__));
  or1   g2419(.dina(new_new_n5229__), .dinb(new_new_n5231__), .dout(new_new_n5234__));
  or1   g2420(.dina(new_new_n5215__), .dinb(new_new_n5234__), .dout(new_new_n5235__));
  or1   g2421(.dina(new_new_n5216__), .dinb(new_new_n5233__), .dout(new_new_n5236__));
  and1  g2422(.dina(new_new_n7549__), .dinb(new_new_n5236__), .dout(new_new_n5237__));
  and1  g2423(.dina(new_new_n5235__), .dinb(new_new_n5237__), .dout(new_new_n5238__));
  and1  g2424(.dina(new_new_n3493__), .dinb(new_new_n3636__), .dout(new_new_n5239__));
  and1  g2425(.dina(new_new_n3492__), .dinb(new_new_n3637__), .dout(new_new_n5240__));
  or1   g2426(.dina(new_new_n5239__), .dinb(new_new_n5240__), .dout(new_new_n5241__));
  or1   g2427(.dina(new_new_n3505__), .dinb(new_new_n7602__), .dout(new_new_n5242__));
  or1   g2428(.dina(new_new_n3502__), .dinb(new_new_n7598__), .dout(new_new_n5243__));
  and1  g2429(.dina(new_new_n5242__), .dinb(new_new_n5243__), .dout(new_new_n5244__));
  and1  g2430(.dina(new_new_n3523__), .dinb(new_new_n7617__), .dout(new_new_n5245__));
  or1   g2431(.dina(new_new_n3522__), .dinb(new_new_n5112__), .dout(new_new_n5246__));
  or1   g2432(.dina(new_new_n3530__), .dinb(new_new_n5246__), .dout(new_new_n5247__));
  or1   g2433(.dina(new_new_n3531__), .dinb(new_new_n5245__), .dout(new_new_n5248__));
  and1  g2434(.dina(new_new_n5247__), .dinb(new_new_n5248__), .dout(new_new_n5249__));
  and1  g2435(.dina(new_new_n7679__), .dinb(new_new_n7680__), .dout(new_new_n5250__));
  or1   g2436(.dina(new_new_n7682__), .dinb(new_new_n7683__), .dout(new_new_n5251__));
  and1  g2437(.dina(new_new_n3104__), .dinb(new_new_n7683__), .dout(new_new_n5252__));
  or1   g2438(.dina(new_new_n3105__), .dinb(new_new_n7680__), .dout(new_new_n5253__));
  and1  g2439(.dina(new_new_n5251__), .dinb(new_new_n5253__), .dout(new_new_n5254__));
  or1   g2440(.dina(new_new_n5250__), .dinb(new_new_n5252__), .dout(new_new_n5255__));
  or1   g2441(.dina(new_new_n3588__), .dinb(new_new_n5255__), .dout(new_new_n5256__));
  or1   g2442(.dina(new_new_n3589__), .dinb(new_new_n5254__), .dout(new_new_n5257__));
  and1  g2443(.dina(new_new_n5256__), .dinb(new_new_n5257__), .dout(new_new_n5258__));
  and1  g2444(.dina(new_new_n3592__), .dinb(new_new_n7597__), .dout(new_new_n5259__));
  and1  g2445(.dina(new_new_n7684__), .dinb(new_new_n7601__), .dout(new_new_n5260__));
  or1   g2446(.dina(new_new_n5259__), .dinb(new_new_n5260__), .dout(new_new_n5261__));
  or1   g2447(.dina(new_new_n7550__), .dinb(new_new_n3649__), .dout(new_new_n5262__));
  or1   g2448(.dina(new_new_n7551__), .dinb(new_new_n3648__), .dout(new_new_n5263__));
  and1  g2449(.dina(new_new_n5262__), .dinb(new_new_n5263__), .dout(new_new_n5264__));
  and1  g2450(.dina(new_new_n3624__), .dinb(new_new_n7599__), .dout(new_new_n5265__));
  or1   g2451(.dina(new_new_n3625__), .dinb(new_new_n7603__), .dout(new_new_n5266__));
  and1  g2452(.dina(new_new_n3622__), .dinb(new_new_n7603__), .dout(new_new_n5267__));
  or1   g2453(.dina(new_new_n3623__), .dinb(new_new_n7599__), .dout(new_new_n5268__));
  and1  g2454(.dina(new_new_n5266__), .dinb(new_new_n5268__), .dout(new_new_n5269__));
  or1   g2455(.dina(new_new_n5265__), .dinb(new_new_n5267__), .dout(new_new_n5270__));
  and1  g2456(.dina(new_new_n7685__), .dinb(new_new_n5269__), .dout(new_new_n5271__));
  and1  g2457(.dina(new_new_n3627__), .dinb(new_new_n5270__), .dout(new_new_n5272__));
  or1   g2458(.dina(new_new_n5271__), .dinb(new_new_n5272__), .dout(new_new_n5273__));
  and1  g2459(.dina(new_new_n7274__), .dinb(new_new_n7604__), .dout(new_new_n5274__));
  and1  g2460(.dina(new_new_n3646__), .dinb(new_new_n7605__), .dout(new_new_n5275__));
  or1   g2461(.dina(new_new_n5274__), .dinb(new_new_n5275__), .dout(new_new_n5276__));
  and1  g2462(.dina(new_new_n3472__), .dinb(new_new_n3481__), .dout(new_new_n5277__));
  and1  g2463(.dina(new_new_n3473__), .dinb(new_new_n3480__), .dout(new_new_n5278__));
  or1   g2464(.dina(new_new_n5277__), .dinb(new_new_n5278__), .dout(new_new_n5279__));
  or1   g2465(.dina(new_new_n3576__), .dinb(new_new_n3679__), .dout(new_new_n5280__));
  or1   g2466(.dina(new_new_n3577__), .dinb(new_new_n7686__), .dout(new_new_n5281__));
  and1  g2467(.dina(new_new_n5280__), .dinb(new_new_n5281__), .dout(new_new_n5282__));
  and1  g2468(.dina(new_new_n7687__), .dinb(new_new_n7688__), .dout(new_new_n5283__));
  or1   g2469(.dina(new_new_n7687__), .dinb(new_new_n7688__), .dout(new_new_n5284__));
  and1  g2470(.dina(new_new_n7689__), .dinb(new_new_n7690__), .dout(new_new_n5285__));
  or1   g2471(.dina(new_new_n7610__), .dinb(new_new_n7691__), .dout(new_new_n5286__));
  and1  g2472(.dina(new_new_n7609__), .dinb(new_new_n7691__), .dout(new_new_n5287__));
  or1   g2473(.dina(new_new_n7689__), .dinb(new_new_n7690__), .dout(new_new_n5288__));
  and1  g2474(.dina(new_new_n5286__), .dinb(new_new_n5288__), .dout(new_new_n5289__));
  or1   g2475(.dina(new_new_n5285__), .dinb(new_new_n5287__), .dout(new_new_n5290__));
  and1  g2476(.dina(new_new_n7403__), .dinb(new_new_n5289__), .dout(new_new_n5291__));
  and1  g2477(.dina(new_new_n7401__), .dinb(new_new_n5290__), .dout(new_new_n5292__));
  or1   g2478(.dina(new_new_n5291__), .dinb(new_new_n5292__), .dout(new_new_n5293__));
  or1   g2479(.dina(new_new_n7652__), .dinb(new_new_n7646__), .dout(new_new_n5294__));
  or1   g2480(.dina(new_new_n7650__), .dinb(new_new_n7648__), .dout(new_new_n5295__));
  and1  g2481(.dina(new_new_n5294__), .dinb(new_new_n5295__), .dout(new_new_n5296__));
  and1  g2482(.dina(new_new_n7692__), .dinb(new_new_n7693__), .dout(new_new_n5297__));
  or1   g2483(.dina(new_new_n7692__), .dinb(new_new_n7693__), .dout(new_new_n5298__));
  and1  g2484(.dina(new_new_n3565__), .dinb(new_new_n3620__), .dout(new_new_n5299__));
  and1  g2485(.dina(new_new_n3564__), .dinb(new_new_n3621__), .dout(new_new_n5300__));
  or1   g2486(.dina(new_new_n5299__), .dinb(new_new_n5300__), .dout(new_new_n5301__));
  and1  g2487(.dina(new_new_n3553__), .dinb(new_new_n3570__), .dout(new_new_n5302__));
  and1  g2488(.dina(new_new_n3552__), .dinb(new_new_n3571__), .dout(new_new_n5303__));
  or1   g2489(.dina(new_new_n5302__), .dinb(new_new_n5303__), .dout(new_new_n5304__));
  or1   g2490(.dina(new_new_n7694__), .dinb(new_new_n7695__), .dout(new_new_n5305__));
  and1  g2491(.dina(new_new_n7694__), .dinb(new_new_n7695__), .dout(new_new_n5306__));
  and1  g2492(.dina(new_new_n7373__), .dinb(new_new_n7645__), .dout(new_new_n5307__));
  or1   g2493(.dina(new_new_n7386__), .dinb(new_new_n7642__), .dout(new_new_n5308__));
  and1  g2494(.dina(new_new_n7386__), .dinb(new_new_n7642__), .dout(new_new_n5309__));
  or1   g2495(.dina(new_new_n7373__), .dinb(new_new_n7645__), .dout(new_new_n5310__));
  and1  g2496(.dina(new_new_n5308__), .dinb(new_new_n5310__), .dout(new_new_n5311__));
  or1   g2497(.dina(new_new_n5307__), .dinb(new_new_n5309__), .dout(new_new_n5312__));
  and1  g2498(.dina(new_new_n7682__), .dinb(new_new_n7639__), .dout(new_new_n5313__));
  or1   g2499(.dina(new_new_n7679__), .dinb(new_new_n7636__), .dout(new_new_n5314__));
  and1  g2500(.dina(new_new_n7678__), .dinb(new_new_n7636__), .dout(new_new_n5315__));
  or1   g2501(.dina(new_new_n7681__), .dinb(new_new_n7639__), .dout(new_new_n5316__));
  and1  g2502(.dina(new_new_n5314__), .dinb(new_new_n5316__), .dout(new_new_n5317__));
  or1   g2503(.dina(new_new_n5313__), .dinb(new_new_n5315__), .dout(new_new_n5318__));
  or1   g2504(.dina(new_new_n5312__), .dinb(new_new_n5318__), .dout(new_new_n5319__));
  or1   g2505(.dina(new_new_n5311__), .dinb(new_new_n5317__), .dout(new_new_n5320__));
  and1  g2506(.dina(new_new_n5319__), .dinb(new_new_n5320__), .dout(new_new_n5321__));
  and1  g2507(.dina(new_new_n3944__), .dinb(new_new_n3947__), .dout(new_new_n5322__));
  or1   g2508(.dina(new_new_n3945__), .dinb(new_new_n3946__), .dout(new_new_n5323__));
  and1  g2509(.dina(new_new_n3683__), .dinb(new_new_n3714__), .dout(new_new_n5324__));
  or1   g2510(.dina(new_new_n3682__), .dinb(new_new_n3715__), .dout(new_new_n5325__));
  and1  g2511(.dina(new_new_n7696__), .dinb(new_new_n7697__), .dout(new_new_n5326__));
  or1   g2512(.dina(new_new_n7698__), .dinb(new_new_n7699__), .dout(new_new_n5327__));
  and1  g2513(.dina(new_new_n7698__), .dinb(new_new_n7699__), .dout(new_new_n5328__));
  or1   g2514(.dina(new_new_n7696__), .dinb(new_new_n7697__), .dout(new_new_n5329__));
  and1  g2515(.dina(new_new_n5327__), .dinb(new_new_n5329__), .dout(new_new_n5330__));
  or1   g2516(.dina(new_new_n5326__), .dinb(new_new_n5328__), .dout(new_new_n5331__));
  and1  g2517(.dina(new_new_n7701__), .dinb(new_new_n5331__), .dout(new_new_n5332__));
  or1   g2518(.dina(new_new_n7704__), .dinb(new_new_n5330__), .dout(new_new_n5333__));
  and1  g2519(.dina(new_new_n3983__), .dinb(new_new_n3984__), .dout(new_new_n5334__));
  or1   g2520(.dina(new_new_n3982__), .dinb(new_new_n3985__), .dout(new_new_n5335__));
  and1  g2521(.dina(new_new_n3992__), .dinb(new_new_n3995__), .dout(new_new_n5336__));
  or1   g2522(.dina(new_new_n3993__), .dinb(new_new_n3994__), .dout(new_new_n5337__));
  and1  g2523(.dina(new_new_n7706__), .dinb(new_new_n7707__), .dout(new_new_n5338__));
  or1   g2524(.dina(new_new_n7708__), .dinb(new_new_n7709__), .dout(new_new_n5339__));
  and1  g2525(.dina(new_new_n7708__), .dinb(new_new_n7709__), .dout(new_new_n5340__));
  or1   g2526(.dina(new_new_n7706__), .dinb(new_new_n7707__), .dout(new_new_n5341__));
  and1  g2527(.dina(new_new_n5339__), .dinb(new_new_n5341__), .dout(new_new_n5342__));
  or1   g2528(.dina(new_new_n5338__), .dinb(new_new_n5340__), .dout(new_new_n5343__));
  and1  g2529(.dina(new_new_n7704__), .dinb(new_new_n5342__), .dout(new_new_n5344__));
  or1   g2530(.dina(new_new_n7701__), .dinb(new_new_n5343__), .dout(new_new_n5345__));
  and1  g2531(.dina(new_new_n5333__), .dinb(new_new_n5345__), .dout(new_new_n5346__));
  or1   g2532(.dina(new_new_n5332__), .dinb(new_new_n5344__), .dout(new_new_n5347__));
  and1  g2533(.dina(new_new_n3951__), .dinb(new_new_n3952__), .dout(new_new_n5348__));
  or1   g2534(.dina(new_new_n3950__), .dinb(new_new_n3953__), .dout(new_new_n5349__));
  and1  g2535(.dina(new_new_n7590__), .dinb(new_new_n7588__), .dout(new_new_n5350__));
  or1   g2536(.dina(new_new_n7594__), .dinb(new_new_n7584__), .dout(new_new_n5351__));
  and1  g2537(.dina(new_new_n7710__), .dinb(new_new_n5351__), .dout(new_new_n5352__));
  or1   g2538(.dina(new_new_n7711__), .dinb(new_new_n5350__), .dout(new_new_n5353__));
  and1  g2539(.dina(new_new_n7591__), .dinb(new_new_n4017__), .dout(new_new_n5354__));
  or1   g2540(.dina(new_new_n7593__), .dinb(new_new_n4016__), .dout(new_new_n5355__));
  and1  g2541(.dina(new_new_n7587__), .dinb(new_new_n7712__), .dout(new_new_n5356__));
  or1   g2542(.dina(new_new_n7585__), .dinb(new_new_n7713__), .dout(new_new_n5357__));
  and1  g2543(.dina(new_new_n5353__), .dinb(new_new_n5357__), .dout(new_new_n5358__));
  or1   g2544(.dina(new_new_n5352__), .dinb(new_new_n5356__), .dout(new_new_n5359__));
  and1  g2545(.dina(new_new_n7705__), .dinb(new_new_n5359__), .dout(new_new_n5360__));
  or1   g2546(.dina(new_new_n7702__), .dinb(new_new_n5358__), .dout(new_new_n5361__));
  and1  g2547(.dina(new_new_n7595__), .dinb(new_new_n7710__), .dout(new_new_n5362__));
  or1   g2548(.dina(new_new_n7591__), .dinb(new_new_n7711__), .dout(new_new_n5363__));
  and1  g2549(.dina(new_new_n7713__), .dinb(new_new_n5363__), .dout(new_new_n5364__));
  or1   g2550(.dina(new_new_n7712__), .dinb(new_new_n5362__), .dout(new_new_n5365__));
  and1  g2551(.dina(new_new_n7702__), .dinb(new_new_n5365__), .dout(new_new_n5366__));
  or1   g2552(.dina(new_new_n7705__), .dinb(new_new_n5364__), .dout(new_new_n5367__));
  and1  g2553(.dina(new_new_n5361__), .dinb(new_new_n5367__), .dout(new_new_n5368__));
  or1   g2554(.dina(new_new_n5360__), .dinb(new_new_n5366__), .dout(new_new_n5369__));
  or1   g2555(.dina(new_new_n5346__), .dinb(new_new_n5369__), .dout(new_new_n5370__));
  or1   g2556(.dina(new_new_n5347__), .dinb(new_new_n5368__), .dout(new_new_n5371__));
  and1  g2557(.dina(new_new_n5370__), .dinb(new_new_n5371__), .dout(new_new_n5372__));
  or1   g2558(.dina(new_new_n7486__), .dinb(new_new_n7488__), .dout(new_new_n5373__));
  and1  g2559(.dina(new_new_n7714__), .dinb(new_new_n7716__), .dout(new_new_n5374__));
  or1   g2560(.dina(new_new_n4978__), .dinb(new_new_n5374__), .dout(new_new_n5375__));
  and1  g2561(.dina(new_new_n7717__), .dinb(new_new_n7517__), .dout(new_new_n5376__));
  and1  g2562(.dina(new_new_n7718__), .dinb(new_new_n7722__), .dout(new_new_n5377__));
  and1  g2563(.dina(new_new_n7735__), .dinb(new_new_n7739__), .dout(new_new_n5378__));
  or1   g2564(.dina(new_new_n5377__), .dinb(new_new_n5378__), .dout(new_new_n5379__));
  and1  g2565(.dina(new_new_n3700__), .dinb(new_new_n5379__), .dout(new_new_n5380__));
  and1  g2566(.dina(new_new_n7735__), .dinb(new_new_n7753__), .dout(new_new_n5381__));
  and1  g2567(.dina(new_new_n7718__), .dinb(new_new_n7766__), .dout(new_new_n5382__));
  or1   g2568(.dina(new_new_n5381__), .dinb(new_new_n5382__), .dout(new_new_n5383__));
  and1  g2569(.dina(new_new_n3701__), .dinb(new_new_n5383__), .dout(new_new_n5384__));
  or1   g2570(.dina(new_new_n5380__), .dinb(new_new_n5384__), .dout(new_new_n5385__));
  and1  g2571(.dina(new_new_n7777__), .dinb(new_new_n7722__), .dout(new_new_n5386__));
  and1  g2572(.dina(new_new_n7779__), .dinb(new_new_n7739__), .dout(new_new_n5387__));
  or1   g2573(.dina(new_new_n5386__), .dinb(new_new_n5387__), .dout(new_new_n5388__));
  and1  g2574(.dina(new_new_n3728__), .dinb(new_new_n5388__), .dout(new_new_n5389__));
  and1  g2575(.dina(new_new_n7779__), .dinb(new_new_n7753__), .dout(new_new_n5390__));
  and1  g2576(.dina(new_new_n7777__), .dinb(new_new_n7766__), .dout(new_new_n5391__));
  or1   g2577(.dina(new_new_n5390__), .dinb(new_new_n5391__), .dout(new_new_n5392__));
  and1  g2578(.dina(new_new_n3729__), .dinb(new_new_n5392__), .dout(new_new_n5393__));
  or1   g2579(.dina(new_new_n5389__), .dinb(new_new_n5393__), .dout(new_new_n5394__));
  and1  g2580(.dina(new_new_n3753__), .dinb(new_new_n7723__), .dout(new_new_n5395__));
  and1  g2581(.dina(new_new_n7780__), .dinb(new_new_n7740__), .dout(new_new_n5396__));
  or1   g2582(.dina(new_new_n5395__), .dinb(new_new_n5396__), .dout(new_new_n5397__));
  and1  g2583(.dina(new_new_n3959__), .dinb(new_new_n7723__), .dout(new_new_n5398__));
  and1  g2584(.dina(new_new_n7781__), .dinb(new_new_n7740__), .dout(new_new_n5399__));
  or1   g2585(.dina(new_new_n5398__), .dinb(new_new_n5399__), .dout(new_new_n5400__));
  or1   g2586(.dina(new_new_n7783__), .dinb(new_new_n7767__), .dout(new_new_n5401__));
  or1   g2587(.dina(new_new_n3109__), .dinb(new_new_n7754__), .dout(new_new_n5402__));
  and1  g2588(.dina(new_new_n5401__), .dinb(new_new_n5402__), .dout(new_new_n5403__));
  and1  g2589(.dina(new_new_n7784__), .dinb(new_new_n7423__), .dout(new_new_n5404__));
  or1   g2590(.dina(new_new_n3091__), .dinb(new_new_n7432__), .dout(new_new_n5405__));
  and1  g2591(.dina(new_new_n3092__), .dinb(new_new_n7433__), .dout(new_new_n5406__));
  or1   g2592(.dina(new_new_n3093__), .dinb(new_new_n7423__), .dout(new_new_n5407__));
  and1  g2593(.dina(new_new_n5405__), .dinb(new_new_n5407__), .dout(new_new_n5408__));
  or1   g2594(.dina(new_new_n5404__), .dinb(new_new_n5406__), .dout(new_new_n5409__));
  and1  g2595(.dina(new_new_n7785__), .dinb(new_new_n7450__), .dout(new_new_n5410__));
  or1   g2596(.dina(new_new_n3131__), .dinb(new_new_n7459__), .dout(new_new_n5411__));
  and1  g2597(.dina(new_new_n7786__), .dinb(new_new_n7462__), .dout(new_new_n5412__));
  or1   g2598(.dina(new_new_n3133__), .dinb(new_new_n7450__), .dout(new_new_n5413__));
  and1  g2599(.dina(new_new_n5411__), .dinb(new_new_n5413__), .dout(new_new_n5414__));
  or1   g2600(.dina(new_new_n5410__), .dinb(new_new_n5412__), .dout(new_new_n5415__));
  or1   g2601(.dina(new_new_n3193__), .dinb(new_new_n4989__), .dout(new_new_n5416__));
  or1   g2602(.dina(new_new_n7499__), .dinb(new_new_n7501__), .dout(new_new_n5417__));
  and1  g2603(.dina(new_new_n4992__), .dinb(new_new_n5417__), .dout(new_new_n5418__));
  or1   g2604(.dina(new_new_n7503__), .dinb(new_new_n7505__), .dout(new_new_n5419__));
  and1  g2605(.dina(new_new_n4994__), .dinb(new_new_n5419__), .dout(new_new_n5420__));
  and1  g2606(.dina(new_new_n7788__), .dinb(new_new_n7366__), .dout(new_new_n5421__));
  or1   g2607(.dina(new_new_n7791__), .dinb(new_new_n7368__), .dout(new_new_n5422__));
  and1  g2608(.dina(new_new_n4023__), .dinb(new_new_n5422__), .dout(new_new_n5423__));
  or1   g2609(.dina(new_new_n7793__), .dinb(new_new_n5421__), .dout(new_new_n5424__));
  and1  g2610(.dina(new_new_n7795__), .dinb(new_new_n7797__), .dout(new_new_n5425__));
  or1   g2611(.dina(new_new_n7415__), .dinb(new_new_n5425__), .dout(new_new_n5426__));
  or1   g2612(.dina(new_new_n7799__), .dinb(new_new_n7801__), .dout(new_new_n5427__));
  or1   g2613(.dina(new_new_n7803__), .dinb(new_new_n7805__), .dout(new_new_n5428__));
  and1  g2614(.dina(new_new_n7806__), .dinb(new_new_n7788__), .dout(new_new_n5429__));
  or1   g2615(.dina(new_new_n7808__), .dinb(new_new_n7791__), .dout(new_new_n5430__));
  and1  g2616(.dina(new_new_n7808__), .dinb(new_new_n7792__), .dout(new_new_n5431__));
  or1   g2617(.dina(new_new_n7806__), .dinb(new_new_n7789__), .dout(new_new_n5432__));
  and1  g2618(.dina(new_new_n5430__), .dinb(new_new_n5432__), .dout(new_new_n5433__));
  or1   g2619(.dina(new_new_n5429__), .dinb(new_new_n5431__), .dout(new_new_n5434__));
  and1  g2620(.dina(new_new_n7810__), .dinb(new_new_n7811__), .dout(new_new_n5435__));
  or1   g2621(.dina(new_new_n7813__), .dinb(new_new_n7815__), .dout(new_new_n5436__));
  and1  g2622(.dina(new_new_n7813__), .dinb(new_new_n7815__), .dout(new_new_n5437__));
  or1   g2623(.dina(new_new_n7810__), .dinb(new_new_n7811__), .dout(new_new_n5438__));
  and1  g2624(.dina(new_new_n5436__), .dinb(new_new_n5438__), .dout(new_new_n5439__));
  or1   g2625(.dina(new_new_n5435__), .dinb(new_new_n5437__), .dout(new_new_n5440__));
  and1  g2626(.dina(new_new_n3743__), .dinb(new_new_n3955__), .dout(new_new_n5441__));
  or1   g2627(.dina(new_new_n7816__), .dinb(new_new_n7817__), .dout(new_new_n5442__));
  and1  g2628(.dina(new_new_n7799__), .dinb(new_new_n5442__), .dout(new_new_n5443__));
  or1   g2629(.dina(new_new_n7819__), .dinb(new_new_n5441__), .dout(new_new_n5444__));
  and1  g2630(.dina(new_new_n7822__), .dinb(new_new_n7824__), .dout(new_new_n5445__));
  or1   g2631(.dina(new_new_n7797__), .dinb(new_new_n7826__), .dout(new_new_n5446__));
  and1  g2632(.dina(new_new_n7796__), .dinb(new_new_n7826__), .dout(new_new_n5447__));
  or1   g2633(.dina(new_new_n7822__), .dinb(new_new_n7824__), .dout(new_new_n5448__));
  and1  g2634(.dina(new_new_n5446__), .dinb(new_new_n5448__), .dout(new_new_n5449__));
  or1   g2635(.dina(new_new_n5445__), .dinb(new_new_n5447__), .dout(new_new_n5450__));
  and1  g2636(.dina(new_new_n5440__), .dinb(new_new_n5450__), .dout(new_new_n5451__));
  and1  g2637(.dina(new_new_n5439__), .dinb(new_new_n5449__), .dout(new_new_n5452__));
  or1   g2638(.dina(new_new_n5451__), .dinb(new_new_n5452__), .dout(new_new_n5453__));
  and1  g2639(.dina(new_new_n7803__), .dinb(new_new_n7827__), .dout(new_new_n5454__));
  or1   g2640(.dina(new_new_n7804__), .dinb(new_new_n7827__), .dout(new_new_n5455__));
  or1   g2641(.dina(new_new_n7507__), .dinb(new_new_n7509__), .dout(new_new_n5456__));
  and1  g2642(.dina(new_new_n4041__), .dinb(new_new_n4042__), .dout(new_new_n5457__));
  or1   g2643(.dina(new_new_n4040__), .dinb(new_new_n4043__), .dout(new_new_n5458__));
  and1  g2644(.dina(new_new_n7829__), .dinb(new_new_n7830__), .dout(new_new_n5459__));
  or1   g2645(.dina(new_new_n7831__), .dinb(new_new_n7832__), .dout(new_new_n5460__));
  and1  g2646(.dina(new_new_n7831__), .dinb(new_new_n7832__), .dout(new_new_n5461__));
  or1   g2647(.dina(new_new_n7829__), .dinb(new_new_n7830__), .dout(new_new_n5462__));
  and1  g2648(.dina(new_new_n5460__), .dinb(new_new_n5462__), .dout(new_new_n5463__));
  or1   g2649(.dina(new_new_n5459__), .dinb(new_new_n5461__), .dout(new_new_n5464__));
  and1  g2650(.dina(new_new_n7833__), .dinb(new_new_n5463__), .dout(new_new_n5465__));
  or1   g2651(.dina(new_new_n7835__), .dinb(new_new_n7837__), .dout(new_new_n5466__));
  and1  g2652(.dina(new_new_n7835__), .dinb(new_new_n7837__), .dout(new_new_n5467__));
  or1   g2653(.dina(new_new_n7838__), .dinb(new_new_n5467__), .dout(new_new_n5468__));
  and1  g2654(.dina(new_new_n7294__), .dinb(new_new_n7295__), .dout(new_new_n5469__));
  or1   g2655(.dina(new_new_n7291__), .dinb(new_new_n7293__), .dout(new_new_n5470__));
  and1  g2656(.dina(new_new_n4844__), .dinb(new_new_n5470__), .dout(new_new_n5471__));
  or1   g2657(.dina(new_new_n7839__), .dinb(new_new_n5469__), .dout(new_new_n5472__));
  and1  g2658(.dina(new_new_n7841__), .dinb(new_new_n7842__), .dout(new_new_n5473__));
  or1   g2659(.dina(new_new_n7843__), .dinb(new_new_n7844__), .dout(new_new_n5474__));
  and1  g2660(.dina(new_new_n7843__), .dinb(new_new_n7844__), .dout(new_new_n5475__));
  or1   g2661(.dina(new_new_n7841__), .dinb(new_new_n7842__), .dout(new_new_n5476__));
  and1  g2662(.dina(new_new_n5474__), .dinb(new_new_n5476__), .dout(new_new_n5477__));
  or1   g2663(.dina(new_new_n5473__), .dinb(new_new_n5475__), .dout(new_new_n5478__));
  and1  g2664(.dina(new_new_n7845__), .dinb(new_new_n7847__), .dout(new_new_n5479__));
  or1   g2665(.dina(new_new_n7845__), .dinb(new_new_n7847__), .dout(new_new_n5480__));
  and1  g2666(.dina(new_new_n4977__), .dinb(new_new_n7848__), .dout(new_new_n5481__));
  and1  g2667(.dina(new_new_n7849__), .dinb(new_new_n7850__), .dout(new_new_n5482__));
  or1   g2668(.dina(new_new_n4996__), .dinb(new_new_n5482__), .dout(new_new_n5483__));
  and1  g2669(.dina(new_new_n7783__), .dinb(new_new_n7851__), .dout(new_new_n5484__));
  and1  g2670(.dina(new_new_n7852__), .dinb(new_new_n3657__), .dout(new_new_n5485__));
  or1   g2671(.dina(new_new_n5484__), .dinb(new_new_n5485__), .dout(new_new_n5486__));
  and1  g2672(.dina(new_new_n7853__), .dinb(new_new_n7725__), .dout(new_new_n5487__));
  and1  g2673(.dina(new_new_n7855__), .dinb(new_new_n7742__), .dout(new_new_n5488__));
  or1   g2674(.dina(new_new_n5487__), .dinb(new_new_n5488__), .dout(new_new_n5489__));
  and1  g2675(.dina(new_new_n7856__), .dinb(new_new_n5489__), .dout(new_new_n5490__));
  and1  g2676(.dina(new_new_n7855__), .dinb(new_new_n7754__), .dout(new_new_n5491__));
  and1  g2677(.dina(new_new_n7853__), .dinb(new_new_n7767__), .dout(new_new_n5492__));
  or1   g2678(.dina(new_new_n5491__), .dinb(new_new_n5492__), .dout(new_new_n5493__));
  and1  g2679(.dina(new_new_n3667__), .dinb(new_new_n5493__), .dout(new_new_n5494__));
  or1   g2680(.dina(new_new_n5490__), .dinb(new_new_n5494__), .dout(new_new_n5495__));
  and1  g2681(.dina(new_new_n7857__), .dinb(new_new_n7725__), .dout(new_new_n5496__));
  and1  g2682(.dina(new_new_n7859__), .dinb(new_new_n7742__), .dout(new_new_n5497__));
  or1   g2683(.dina(new_new_n5496__), .dinb(new_new_n5497__), .dout(new_new_n5498__));
  and1  g2684(.dina(new_new_n7860__), .dinb(new_new_n5498__), .dout(new_new_n5499__));
  and1  g2685(.dina(new_new_n7859__), .dinb(new_new_n7756__), .dout(new_new_n5500__));
  and1  g2686(.dina(new_new_n7857__), .dinb(new_new_n7769__), .dout(new_new_n5501__));
  or1   g2687(.dina(new_new_n5500__), .dinb(new_new_n5501__), .dout(new_new_n5502__));
  and1  g2688(.dina(new_new_n3669__), .dinb(new_new_n5502__), .dout(new_new_n5503__));
  or1   g2689(.dina(new_new_n5499__), .dinb(new_new_n5503__), .dout(new_new_n5504__));
  and1  g2690(.dina(new_new_n7861__), .dinb(new_new_n7726__), .dout(new_new_n5505__));
  and1  g2691(.dina(new_new_n7863__), .dinb(new_new_n7743__), .dout(new_new_n5506__));
  or1   g2692(.dina(new_new_n5505__), .dinb(new_new_n5506__), .dout(new_new_n5507__));
  and1  g2693(.dina(new_new_n7864__), .dinb(new_new_n5507__), .dout(new_new_n5508__));
  and1  g2694(.dina(new_new_n7863__), .dinb(new_new_n7756__), .dout(new_new_n5509__));
  and1  g2695(.dina(new_new_n7861__), .dinb(new_new_n7769__), .dout(new_new_n5510__));
  or1   g2696(.dina(new_new_n5509__), .dinb(new_new_n5510__), .dout(new_new_n5511__));
  and1  g2697(.dina(new_new_n3671__), .dinb(new_new_n5511__), .dout(new_new_n5512__));
  or1   g2698(.dina(new_new_n5508__), .dinb(new_new_n5512__), .dout(new_new_n5513__));
  and1  g2699(.dina(new_new_n7865__), .dinb(new_new_n7726__), .dout(new_new_n5514__));
  and1  g2700(.dina(new_new_n7867__), .dinb(new_new_n7743__), .dout(new_new_n5515__));
  or1   g2701(.dina(new_new_n5514__), .dinb(new_new_n5515__), .dout(new_new_n5516__));
  and1  g2702(.dina(new_new_n7868__), .dinb(new_new_n5516__), .dout(new_new_n5517__));
  and1  g2703(.dina(new_new_n7867__), .dinb(new_new_n7757__), .dout(new_new_n5518__));
  and1  g2704(.dina(new_new_n7865__), .dinb(new_new_n7770__), .dout(new_new_n5519__));
  or1   g2705(.dina(new_new_n5518__), .dinb(new_new_n5519__), .dout(new_new_n5520__));
  and1  g2706(.dina(new_new_n3699__), .dinb(new_new_n5520__), .dout(new_new_n5521__));
  or1   g2707(.dina(new_new_n5517__), .dinb(new_new_n5521__), .dout(new_new_n5522__));
  and1  g2708(.dina(new_new_n7869__), .dinb(new_new_n7729__), .dout(new_new_n5523__));
  and1  g2709(.dina(new_new_n7871__), .dinb(new_new_n7746__), .dout(new_new_n5524__));
  or1   g2710(.dina(new_new_n5523__), .dinb(new_new_n5524__), .dout(new_new_n5525__));
  and1  g2711(.dina(new_new_n7872__), .dinb(new_new_n5525__), .dout(new_new_n5526__));
  and1  g2712(.dina(new_new_n7871__), .dinb(new_new_n7757__), .dout(new_new_n5527__));
  and1  g2713(.dina(new_new_n7869__), .dinb(new_new_n7770__), .dout(new_new_n5528__));
  or1   g2714(.dina(new_new_n5527__), .dinb(new_new_n5528__), .dout(new_new_n5529__));
  and1  g2715(.dina(new_new_n3725__), .dinb(new_new_n5529__), .dout(new_new_n5530__));
  or1   g2716(.dina(new_new_n5526__), .dinb(new_new_n5530__), .dout(new_new_n5531__));
  and1  g2717(.dina(new_new_n7873__), .dinb(new_new_n7729__), .dout(new_new_n5532__));
  and1  g2718(.dina(new_new_n7875__), .dinb(new_new_n7746__), .dout(new_new_n5533__));
  or1   g2719(.dina(new_new_n5532__), .dinb(new_new_n5533__), .dout(new_new_n5534__));
  and1  g2720(.dina(new_new_n7876__), .dinb(new_new_n5534__), .dout(new_new_n5535__));
  and1  g2721(.dina(new_new_n7875__), .dinb(new_new_n7760__), .dout(new_new_n5536__));
  and1  g2722(.dina(new_new_n7873__), .dinb(new_new_n7773__), .dout(new_new_n5537__));
  or1   g2723(.dina(new_new_n5536__), .dinb(new_new_n5537__), .dout(new_new_n5538__));
  and1  g2724(.dina(new_new_n3727__), .dinb(new_new_n5538__), .dout(new_new_n5539__));
  or1   g2725(.dina(new_new_n5535__), .dinb(new_new_n5539__), .dout(new_new_n5540__));
  and1  g2726(.dina(new_new_n7877__), .dinb(new_new_n7747__), .dout(new_new_n5541__));
  and1  g2727(.dina(new_new_n7879__), .dinb(new_new_n7730__), .dout(new_new_n5542__));
  or1   g2728(.dina(new_new_n5541__), .dinb(new_new_n5542__), .dout(new_new_n5543__));
  and1  g2729(.dina(new_new_n3962__), .dinb(new_new_n5543__), .dout(new_new_n5544__));
  and1  g2730(.dina(new_new_n7877__), .dinb(new_new_n7760__), .dout(new_new_n5545__));
  and1  g2731(.dina(new_new_n7879__), .dinb(new_new_n7773__), .dout(new_new_n5546__));
  or1   g2732(.dina(new_new_n5545__), .dinb(new_new_n5546__), .dout(new_new_n5547__));
  and1  g2733(.dina(new_new_n3963__), .dinb(new_new_n5547__), .dout(new_new_n5548__));
  or1   g2734(.dina(new_new_n5544__), .dinb(new_new_n5548__), .dout(new_new_n5549__));
  and1  g2735(.dina(new_new_n7344__), .dinb(new_new_n7881__), .dout(new_new_n5550__));
  or1   g2736(.dina(new_new_n7340__), .dinb(new_new_n7882__), .dout(new_new_n5551__));
  and1  g2737(.dina(new_new_n7341__), .dinb(new_new_n7882__), .dout(new_new_n5552__));
  or1   g2738(.dina(new_new_n7343__), .dinb(new_new_n7881__), .dout(new_new_n5553__));
  and1  g2739(.dina(new_new_n5551__), .dinb(new_new_n5553__), .dout(new_new_n5554__));
  or1   g2740(.dina(new_new_n5550__), .dinb(new_new_n5552__), .dout(new_new_n5555__));
  and1  g2741(.dina(new_new_n7335__), .dinb(new_new_n5555__), .dout(new_new_n5556__));
  and1  g2742(.dina(new_new_n7334__), .dinb(new_new_n5554__), .dout(new_new_n5557__));
  or1   g2743(.dina(new_new_n5556__), .dinb(new_new_n5557__), .dout(new_new_n5558__));
  and1  g2744(.dina(new_new_n7821__), .dinb(new_new_n7805__), .dout(new_new_n5559__));
  and1  g2745(.dina(new_new_n7809__), .dinb(new_new_n7800__), .dout(new_new_n5560__));
  or1   g2746(.dina(new_new_n7814__), .dinb(new_new_n7819__), .dout(new_new_n5561__));
  and1  g2747(.dina(new_new_n7363__), .dinb(new_new_n7820__), .dout(new_new_n5562__));
  or1   g2748(.dina(new_new_n7367__), .dinb(new_new_n7800__), .dout(new_new_n5563__));
  and1  g2749(.dina(new_new_n7792__), .dinb(new_new_n5563__), .dout(new_new_n5564__));
  or1   g2750(.dina(new_new_n7789__), .dinb(new_new_n5562__), .dout(new_new_n5565__));
  and1  g2751(.dina(new_new_n7883__), .dinb(new_new_n7884__), .dout(new_new_n5566__));
  or1   g2752(.dina(new_new_n7885__), .dinb(new_new_n7886__), .dout(new_new_n5567__));
  and1  g2753(.dina(new_new_n7885__), .dinb(new_new_n7886__), .dout(new_new_n5568__));
  or1   g2754(.dina(new_new_n7883__), .dinb(new_new_n7884__), .dout(new_new_n5569__));
  and1  g2755(.dina(new_new_n5567__), .dinb(new_new_n5569__), .dout(new_new_n5570__));
  or1   g2756(.dina(new_new_n5566__), .dinb(new_new_n5568__), .dout(new_new_n5571__));
  and1  g2757(.dina(new_new_n5561__), .dinb(new_new_n5570__), .dout(new_new_n5572__));
  and1  g2758(.dina(new_new_n5560__), .dinb(new_new_n5571__), .dout(new_new_n5573__));
  or1   g2759(.dina(new_new_n5572__), .dinb(new_new_n5573__), .dout(new_new_n5574__));
  or1   g2760(.dina(new_new_n7887__), .dinb(new_new_n7888__), .dout(new_new_n5575__));
  and1  g2761(.dina(new_new_n7887__), .dinb(new_new_n7888__), .dout(new_new_n5576__));
  and1  g2762(.dina(new_new_n7889__), .dinb(new_new_n7424__), .dout(new_new_n5577__));
  and1  g2763(.dina(new_new_n3068__), .dinb(new_new_n7433__), .dout(new_new_n5578__));
  or1   g2764(.dina(new_new_n5577__), .dinb(new_new_n5578__), .dout(new_new_n5579__));
  or1   g2765(.dina(new_new_n3139__), .dinb(new_new_n7462__), .dout(new_new_n5580__));
  or1   g2766(.dina(new_new_n3141__), .dinb(new_new_n7452__), .dout(new_new_n5581__));
  and1  g2767(.dina(new_new_n5580__), .dinb(new_new_n5581__), .dout(new_new_n5582__));
  or1   g2768(.dina(new_new_n3189__), .dinb(new_new_n5116__), .dout(new_new_n5583__));
  and1  g2769(.dina(new_new_n7801__), .dinb(new_new_n7890__), .dout(new_new_n5584__));
  or1   g2770(.dina(new_new_n7795__), .dinb(new_new_n7825__), .dout(new_new_n5585__));
  or1   g2771(.dina(new_new_n7804__), .dinb(new_new_n7823__), .dout(new_new_n5586__));
  and1  g2772(.dina(new_new_n5585__), .dinb(new_new_n5586__), .dout(new_new_n5587__));
  or1   g2773(.dina(new_new_n7891__), .dinb(new_new_n7892__), .dout(new_new_n5588__));
  and1  g2774(.dina(new_new_n7891__), .dinb(new_new_n7892__), .dout(new_new_n5589__));
  or1   g2775(.dina(new_new_n7894__), .dinb(new_new_n7895__), .dout(new_new_n5590__));
  or1   g2776(.dina(new_new_n7897__), .dinb(new_new_n7898__), .dout(new_new_n5591__));
  and1  g2777(.dina(new_new_n7900__), .dinb(new_new_n7902__), .dout(new_new_n5592__));
  or1   g2778(.dina(new_new_n7900__), .dinb(new_new_n7902__), .dout(new_new_n5593__));
  and1  g2779(.dina(new_new_n7904__), .dinb(new_new_n7906__), .dout(new_new_n5594__));
  or1   g2780(.dina(new_new_n7904__), .dinb(new_new_n7906__), .dout(new_new_n5595__));
  and1  g2781(.dina(new_new_n7908__), .dinb(new_new_n7730__), .dout(new_new_n5596__));
  or1   g2782(.dina(new_new_n7909__), .dinb(new_new_n7912__), .dout(new_new_n5597__));
  and1  g2783(.dina(new_new_n7909__), .dinb(new_new_n7774__), .dout(new_new_n5598__));
  or1   g2784(.dina(new_new_n7908__), .dinb(new_new_n7916__), .dout(new_new_n5599__));
  and1  g2785(.dina(new_new_n5597__), .dinb(new_new_n5599__), .dout(new_new_n5600__));
  or1   g2786(.dina(new_new_n5596__), .dinb(new_new_n5598__), .dout(new_new_n5601__));
  and1  g2787(.dina(new_new_n7919__), .dinb(new_new_n7732__), .dout(new_new_n5602__));
  or1   g2788(.dina(new_new_n7923__), .dinb(new_new_n7912__), .dout(new_new_n5603__));
  and1  g2789(.dina(new_new_n7923__), .dinb(new_new_n7747__), .dout(new_new_n5604__));
  or1   g2790(.dina(new_new_n7919__), .dinb(new_new_n7926__), .dout(new_new_n5605__));
  and1  g2791(.dina(new_new_n5603__), .dinb(new_new_n5605__), .dout(new_new_n5606__));
  or1   g2792(.dina(new_new_n5602__), .dinb(new_new_n5604__), .dout(new_new_n5607__));
  and1  g2793(.dina(new_new_n7347__), .dinb(new_new_n5607__), .dout(new_new_n5608__));
  or1   g2794(.dina(new_new_n7354__), .dinb(new_new_n5606__), .dout(new_new_n5609__));
  and1  g2795(.dina(new_new_n7922__), .dinb(new_new_n7761__), .dout(new_new_n5610__));
  or1   g2796(.dina(new_new_n7920__), .dinb(new_new_n7929__), .dout(new_new_n5611__));
  and1  g2797(.dina(new_new_n7920__), .dinb(new_new_n7774__), .dout(new_new_n5612__));
  or1   g2798(.dina(new_new_n7924__), .dinb(new_new_n7916__), .dout(new_new_n5613__));
  and1  g2799(.dina(new_new_n5611__), .dinb(new_new_n5613__), .dout(new_new_n5614__));
  or1   g2800(.dina(new_new_n5610__), .dinb(new_new_n5612__), .dout(new_new_n5615__));
  and1  g2801(.dina(new_new_n7354__), .dinb(new_new_n5615__), .dout(new_new_n5616__));
  or1   g2802(.dina(new_new_n7349__), .dinb(new_new_n5614__), .dout(new_new_n5617__));
  and1  g2803(.dina(new_new_n5609__), .dinb(new_new_n5617__), .dout(new_new_n5618__));
  or1   g2804(.dina(new_new_n5608__), .dinb(new_new_n5616__), .dout(new_new_n5619__));
  and1  g2805(.dina(new_new_n5600__), .dinb(new_new_n5619__), .dout(new_new_n5620__));
  and1  g2806(.dina(new_new_n5601__), .dinb(new_new_n5618__), .dout(new_new_n5621__));
  or1   g2807(.dina(new_new_n5620__), .dinb(new_new_n5621__), .dout(new_new_n5622__));
  or1   g2808(.dina(new_new_n7932__), .dinb(new_new_n7933__), .dout(new_new_n5623__));
  and1  g2809(.dina(new_new_n7932__), .dinb(new_new_n7933__), .dout(new_new_n5624__));
  and1  g2810(.dina(new_new_n7934__), .dinb(new_new_n7732__), .dout(new_new_n5625__));
  and1  g2811(.dina(new_new_n7936__), .dinb(new_new_n7749__), .dout(new_new_n5626__));
  or1   g2812(.dina(new_new_n5625__), .dinb(new_new_n5626__), .dout(new_new_n5627__));
  and1  g2813(.dina(new_new_n7937__), .dinb(new_new_n5627__), .dout(new_new_n5628__));
  and1  g2814(.dina(new_new_n7936__), .dinb(new_new_n7761__), .dout(new_new_n5629__));
  and1  g2815(.dina(new_new_n7934__), .dinb(new_new_n7776__), .dout(new_new_n5630__));
  or1   g2816(.dina(new_new_n5629__), .dinb(new_new_n5630__), .dout(new_new_n5631__));
  and1  g2817(.dina(new_new_n3757__), .dinb(new_new_n5631__), .dout(new_new_n5632__));
  or1   g2818(.dina(new_new_n5628__), .dinb(new_new_n5632__), .dout(new_new_n5633__));
  or1   g2819(.dina(new_new_n7939__), .dinb(new_new_n7911__), .dout(new_new_n5634__));
  or1   g2820(.dina(new_new_n7940__), .dinb(new_new_n7926__), .dout(new_new_n5635__));
  and1  g2821(.dina(new_new_n5634__), .dinb(new_new_n5635__), .dout(new_new_n5636__));
  or1   g2822(.dina(new_new_n3929__), .dinb(new_new_n5636__), .dout(new_new_n5637__));
  or1   g2823(.dina(new_new_n7940__), .dinb(new_new_n7929__), .dout(new_new_n5638__));
  or1   g2824(.dina(new_new_n7939__), .dinb(new_new_n7915__), .dout(new_new_n5639__));
  and1  g2825(.dina(new_new_n5638__), .dinb(new_new_n5639__), .dout(new_new_n5640__));
  or1   g2826(.dina(new_new_n7941__), .dinb(new_new_n5640__), .dout(new_new_n5641__));
  and1  g2827(.dina(new_new_n5637__), .dinb(new_new_n5641__), .dout(new_new_n5642__));
  or1   g2828(.dina(new_new_n7942__), .dinb(new_new_n7943__), .dout(new_new_n5643__));
  and1  g2829(.dina(new_new_n7942__), .dinb(new_new_n7943__), .dout(new_new_n5644__));
  and1  g2830(.dina(new_new_n3957__), .dinb(new_new_n7479__), .dout(new_new_n5645__));
  and1  g2831(.dina(new_new_n7944__), .dinb(new_new_n7474__), .dout(new_new_n5646__));
  or1   g2832(.dina(new_new_n5645__), .dinb(new_new_n5646__), .dout(new_new_n5647__));
  and1  g2833(.dina(new_new_n7482__), .dinb(new_new_n5647__), .dout(new_new_n5648__));
  or1   g2834(.dina(new_new_n7483__), .dinb(new_new_n5648__), .dout(new_new_n5649__));
  and1  g2835(.dina(new_new_n4944__), .dinb(new_new_n5649__), .dout(new_new_n5650__));
  and1  g2836(.dina(new_new_n7945__), .dinb(new_new_n7946__), .dout(new_new_n5651__));
  or1   g2837(.dina(new_new_n5650__), .dinb(new_new_n5651__), .dout(new_new_n5652__));
  and1  g2838(.dina(new_new_n7948__), .dinb(new_new_n7949__), .dout(new_new_n5653__));
  or1   g2839(.dina(new_new_n7950__), .dinb(new_new_n7952__), .dout(new_new_n5654__));
  and1  g2840(.dina(new_new_n7950__), .dinb(new_new_n7952__), .dout(new_new_n5655__));
  or1   g2841(.dina(new_new_n7948__), .dinb(new_new_n7949__), .dout(new_new_n5656__));
  and1  g2842(.dina(new_new_n7836__), .dinb(new_new_n5656__), .dout(new_new_n5657__));
  or1   g2843(.dina(new_new_n7833__), .dinb(new_new_n5655__), .dout(new_new_n5658__));
  and1  g2844(.dina(new_new_n5654__), .dinb(new_new_n5657__), .dout(new_new_n5659__));
  or1   g2845(.dina(new_new_n5653__), .dinb(new_new_n5658__), .dout(new_new_n5660__));
  and1  g2846(.dina(new_new_n5466__), .dinb(new_new_n5660__), .dout(new_new_n5661__));
  or1   g2847(.dina(new_new_n7838__), .dinb(new_new_n5659__), .dout(new_new_n5662__));
  or1   g2848(.dina(new_new_n5477__), .dinb(new_new_n5661__), .dout(new_new_n5663__));
  or1   g2849(.dina(new_new_n7846__), .dinb(new_new_n5662__), .dout(new_new_n5664__));
  and1  g2850(.dina(new_new_n5663__), .dinb(new_new_n5664__), .dout(new_new_n5665__));
  and1  g2851(.dina(new_new_n7954__), .dinb(new_new_n7733__), .dout(new_new_n5666__));
  or1   g2852(.dina(new_new_n7958__), .dinb(new_new_n7913__), .dout(new_new_n5667__));
  and1  g2853(.dina(new_new_n7958__), .dinb(new_new_n7749__), .dout(new_new_n5668__));
  or1   g2854(.dina(new_new_n7954__), .dinb(new_new_n7927__), .dout(new_new_n5669__));
  and1  g2855(.dina(new_new_n5667__), .dinb(new_new_n5669__), .dout(new_new_n5670__));
  or1   g2856(.dina(new_new_n5666__), .dinb(new_new_n5668__), .dout(new_new_n5671__));
  and1  g2857(.dina(new_new_n7961__), .dinb(new_new_n5671__), .dout(new_new_n5672__));
  or1   g2858(.dina(new_new_n7962__), .dinb(new_new_n5670__), .dout(new_new_n5673__));
  and1  g2859(.dina(new_new_n7957__), .dinb(new_new_n7762__), .dout(new_new_n5674__));
  or1   g2860(.dina(new_new_n7955__), .dinb(new_new_n7930__), .dout(new_new_n5675__));
  and1  g2861(.dina(new_new_n7955__), .dinb(new_new_n7776__), .dout(new_new_n5676__));
  or1   g2862(.dina(new_new_n7959__), .dinb(new_new_n7917__), .dout(new_new_n5677__));
  and1  g2863(.dina(new_new_n5675__), .dinb(new_new_n5677__), .dout(new_new_n5678__));
  or1   g2864(.dina(new_new_n5674__), .dinb(new_new_n5676__), .dout(new_new_n5679__));
  and1  g2865(.dina(new_new_n7962__), .dinb(new_new_n5679__), .dout(new_new_n5680__));
  or1   g2866(.dina(new_new_n7961__), .dinb(new_new_n5678__), .dout(new_new_n5681__));
  and1  g2867(.dina(new_new_n5673__), .dinb(new_new_n5681__), .dout(new_new_n5682__));
  or1   g2868(.dina(new_new_n5672__), .dinb(new_new_n5680__), .dout(new_new_n5683__));
  and1  g2869(.dina(new_new_n7328__), .dinb(new_new_n7733__), .dout(new_new_n5684__));
  or1   g2870(.dina(new_new_n7322__), .dinb(new_new_n7913__), .dout(new_new_n5685__));
  and1  g2871(.dina(new_new_n7323__), .dinb(new_new_n7748__), .dout(new_new_n5686__));
  or1   g2872(.dina(new_new_n7327__), .dinb(new_new_n7927__), .dout(new_new_n5687__));
  and1  g2873(.dina(new_new_n5685__), .dinb(new_new_n5687__), .dout(new_new_n5688__));
  or1   g2874(.dina(new_new_n5684__), .dinb(new_new_n5686__), .dout(new_new_n5689__));
  and1  g2875(.dina(new_new_n7406__), .dinb(new_new_n5689__), .dout(new_new_n5690__));
  or1   g2876(.dina(new_new_n7413__), .dinb(new_new_n5688__), .dout(new_new_n5691__));
  and1  g2877(.dina(new_new_n7323__), .dinb(new_new_n7762__), .dout(new_new_n5692__));
  or1   g2878(.dina(new_new_n7329__), .dinb(new_new_n7930__), .dout(new_new_n5693__));
  and1  g2879(.dina(new_new_n7329__), .dinb(new_new_n7775__), .dout(new_new_n5694__));
  or1   g2880(.dina(new_new_n7324__), .dinb(new_new_n7917__), .dout(new_new_n5695__));
  and1  g2881(.dina(new_new_n5693__), .dinb(new_new_n5695__), .dout(new_new_n5696__));
  or1   g2882(.dina(new_new_n5692__), .dinb(new_new_n5694__), .dout(new_new_n5697__));
  and1  g2883(.dina(new_new_n7413__), .dinb(new_new_n5697__), .dout(new_new_n5698__));
  or1   g2884(.dina(new_new_n7408__), .dinb(new_new_n5696__), .dout(new_new_n5699__));
  and1  g2885(.dina(new_new_n5691__), .dinb(new_new_n5699__), .dout(new_new_n5700__));
  or1   g2886(.dina(new_new_n5690__), .dinb(new_new_n5698__), .dout(new_new_n5701__));
  and1  g2887(.dina(new_new_n5682__), .dinb(new_new_n5701__), .dout(new_new_n5702__));
  and1  g2888(.dina(new_new_n5683__), .dinb(new_new_n5700__), .dout(new_new_n5703__));
  or1   g2889(.dina(new_new_n5702__), .dinb(new_new_n5703__), .dout(new_new_n5704__));
  and1  g2890(.dina(new_new_n7963__), .dinb(new_new_n4862__), .dout(new_new_n5705__));
  or1   g2891(.dina(new_new_n7964__), .dinb(new_new_n7965__), .dout(new_new_n5706__));
  and1  g2892(.dina(new_new_n7964__), .dinb(new_new_n7342__), .dout(new_new_n5707__));
  or1   g2893(.dina(new_new_n7963__), .dinb(new_new_n7345__), .dout(new_new_n5708__));
  and1  g2894(.dina(new_new_n5706__), .dinb(new_new_n5708__), .dout(new_new_n5709__));
  or1   g2895(.dina(new_new_n5705__), .dinb(new_new_n5707__), .dout(new_new_n5710__));
  and1  g2896(.dina(new_new_n7966__), .dinb(new_new_n5710__), .dout(new_new_n5711__));
  and1  g2897(.dina(new_new_n4975__), .dinb(new_new_n5709__), .dout(new_new_n5712__));
  or1   g2898(.dina(new_new_n5711__), .dinb(new_new_n5712__), .dout(new_new_n5713__));
  or1   g2899(.dina(new_new_n3173__), .dinb(new_new_n5408__), .dout(new_new_n5714__));
  or1   g2900(.dina(new_new_n3191__), .dinb(new_new_n5414__), .dout(new_new_n5715__));
  or1   g2901(.dina(new_new_n7967__), .dinb(new_new_n7968__), .dout(new_new_n5716__));
  or1   g2902(.dina(new_new_n7969__), .dinb(new_new_n7970__), .dout(new_new_n5717__));
  and1  g2903(.dina(new_new_n7971__), .dinb(new_new_n5717__), .dout(new_new_n5718__));
  and1  g2904(.dina(new_new_n7972__), .dinb(new_new_n7452__), .dout(new_new_n5719__));
  and1  g2905(.dina(new_new_n3120__), .dinb(new_new_n7463__), .dout(new_new_n5720__));
  and1  g2906(.dina(new_new_n7973__), .dinb(new_new_n7453__), .dout(new_new_n5721__));
  and1  g2907(.dina(new_new_n3124__), .dinb(new_new_n7463__), .dout(new_new_n5722__));
  and1  g2908(.dina(new_new_n7494__), .dinb(new_new_n7975__), .dout(new_new_n5723__));
  or1   g2909(.dina(new_new_n7495__), .dinb(new_new_n7975__), .dout(new_new_n5724__));
  and1  g2910(.dina(new_new_n7894__), .dinb(new_new_n7977__), .dout(new_new_n5725__));
  and1  g2911(.dina(new_new_n7514__), .dinb(new_new_n7980__), .dout(new_new_n5726__));
  and1  g2912(.dina(new_new_n7716__), .dinb(new_new_n7981__), .dout(new_new_n5727__));
  and1  g2913(.dina(new_new_n7982__), .dinb(new_new_n7983__), .dout(new_new_n5728__));
  or1   g2914(.dina(new_new_n7984__), .dinb(new_new_n5728__), .dout(new_new_n5729__));
  and1  g2915(.dina(new_new_n7897__), .dinb(new_new_n7977__), .dout(new_new_n5730__));
  or1   g2916(.dina(new_new_n7985__), .dinb(new_new_n5730__), .dout(new_new_n5731__));
  and1  g2917(.dina(new_new_n7978__), .dinb(new_new_n7898__), .dout(new_new_n5732__));
  or1   g2918(.dina(new_new_n7980__), .dinb(new_new_n7986__), .dout(new_new_n5733__));
  and1  g2919(.dina(new_new_n7988__), .dinb(new_new_n7990__), .dout(new_new_n5734__));
  or1   g2920(.dina(new_new_n7988__), .dinb(new_new_n7990__), .dout(new_new_n5735__));
  and1  g2921(.dina(new_new_n7991__), .dinb(new_new_n7992__), .dout(new_new_n5736__));
  or1   g2922(.dina(new_new_n7993__), .dinb(new_new_n7994__), .dout(new_new_n5737__));
  and1  g2923(.dina(new_new_n7995__), .dinb(new_new_n5737__), .dout(new_new_n5738__));
  or1   g2924(.dina(new_new_n7996__), .dinb(new_new_n7997__), .dout(new_new_n5739__));
  and1  g2925(.dina(new_new_n7998__), .dinb(new_new_n5739__), .dout(new_new_n5740__));
  and1  g2926(.dina(new_new_n7999__), .dinb(new_new_n8000__), .dout(new_new_n5741__));
  and1  g2927(.dina(new_new_n8001__), .dinb(new_new_n8003__), .dout(new_new_n5742__));
  and1  g2928(.dina(new_new_n2226__), .dinb(new_new_n8006__), .dout(new_new_n5743__));
  and1  g2929(.dina(new_new_n8007__), .dinb(new_new_n8003__), .dout(new_new_n5744__));
  and1  g2930(.dina(new_new_n2230__), .dinb(new_new_n8006__), .dout(new_new_n5745__));
  and1  g2931(.dina(new_new_n8008__), .dinb(new_new_n8004__), .dout(new_new_n5746__));
  and1  g2932(.dina(new_new_n2256__), .dinb(new_new_n8005__), .dout(new_new_n5747__));
  buf1  g2933(.din(new_new_n2897__), .dout(G5193));
  buf1  g2934(.din(new_new_n3111__), .dout(G5194));
  buf1  g2935(.din(new_new_n6749__), .dout(G5195));
  buf1  g2936(.din(new_new_n8010__), .dout(G5196));
  buf1  g2937(.din(new_new_n3135__), .dout(G5197));
  buf1  g2938(.din(new_new_n3143__), .dout(G5198));
  not1  g2939(.din(new_new_n7194__), .dout(G5199));
  buf1  g2940(.din(new_new_n3209__), .dout(G5200));
  buf1  g2941(.din(G5196), .dout(G5201));
  buf1  g2942(.din(new_new_n8009__), .dout(G5202));
  buf1  g2943(.din(new_new_n3129__), .dout(G5203));
  buf1  g2944(.din(new_new_n3137__), .dout(G5204));
  buf1  g2945(.din(new_new_n4139__), .dout(G5205));
  buf1  g2946(.din(new_new_n7192__), .dout(G5206));
  buf1  g2947(.din(new_new_n6741__), .dout(G5207));
  buf1  g2948(.din(new_new_n6742__), .dout(G5208));
  buf1  g2949(.din(new_new_n7193__), .dout(G5209));
  buf1  g2950(.din(new_new_n4140__), .dout(G5210));
  buf1  g2951(.din(new_new_n4141__), .dout(G5211));
  buf1  g2952(.din(new_new_n4142__), .dout(G5212));
  buf1  g2953(.din(new_new_n7195__), .dout(G5213));
  buf1  g2954(.din(new_new_n7078__), .dout(G5214));
  buf1  g2955(.din(new_new_n6747__), .dout(G5215));
  buf1  g2956(.din(new_new_n6748__), .dout(G5216));
  buf1  g2957(.din(new_new_n8011__), .dout(G5217));
  buf1  g2958(.din(new_new_n3116__), .dout(G5218));
  buf1  g2959(.din(G5217), .dout(G5219));
  buf1  g2960(.din(new_new_n4145__), .dout(G5220));
  buf1  g2961(.din(new_new_n6758__), .dout(G5221));
  buf1  g2962(.din(new_new_n8013__), .dout(G5222));
  buf1  g2963(.din(G5222), .dout(G5223));
  buf1  g2964(.din(new_new_n8014__), .dout(G5224));
  buf1  g2965(.din(G5224), .dout(G5225));
  buf1  g2966(.din(new_new_n8015__), .dout(G5226));
  buf1  g2967(.din(G5226), .dout(G5227));
  buf1  g2968(.din(new_new_n4149__), .dout(G5228));
  buf1  g2969(.din(new_new_n8016__), .dout(G5229));
  buf1  g2970(.din(G5229), .dout(G5230));
  buf1  g2971(.din(new_new_n4154__), .dout(G5231));
  buf1  g2972(.din(new_new_n4159__), .dout(G5232));
  buf1  g2973(.din(new_new_n4164__), .dout(G5233));
  buf1  g2974(.din(new_new_n4169__), .dout(G5234));
  buf1  g2975(.din(new_new_n4174__), .dout(G5235));
  buf1  g2976(.din(new_new_n4180__), .dout(G5236));
  buf1  g2977(.din(new_new_n4189__), .dout(G5237));
  not1  g2978(.din(new_new_n8017__), .dout(G5238));
  buf1  g2979(.din(new_new_n8018__), .dout(G5239));
  buf1  g2980(.din(G5239), .dout(G5240));
  buf1  g2981(.din(G5238), .dout(G5241));
  not1  g2982(.din(new_new_n7196__), .dout(G5242));
  not1  g2983(.din(new_new_n7197__), .dout(G5243));
  not1  g2984(.din(new_new_n8019__), .dout(G5244));
  buf1  g2985(.din(new_new_n8020__), .dout(G5245));
  buf1  g2986(.din(G5244), .dout(G5246));
  buf1  g2987(.din(G5245), .dout(G5247));
  not1  g2988(.din(new_new_n6855__), .dout(G5248));
  buf1  g2989(.din(new_new_n7174__), .dout(G5249));
  not1  g2990(.din(new_new_n6878__), .dout(G5250));
  buf1  g2991(.din(new_new_n6968__), .dout(G5251));
  buf1  g2992(.din(new_new_n4248__), .dout(G5252));
  not1  g2993(.din(new_new_n7144__), .dout(G5253));
  not1  g2994(.din(new_new_n7154__), .dout(G5254));
  not1  g2995(.din(new_new_n7164__), .dout(G5255));
  buf1  g2996(.din(new_new_n4270__), .dout(G5256));
  not1  g2997(.din(new_new_n7140__), .dout(G5257));
  not1  g2998(.din(new_new_n7150__), .dout(G5258));
  not1  g2999(.din(new_new_n7160__), .dout(G5259));
  buf1  g3000(.din(new_new_n7170__), .dout(G5260));
  not1  g3001(.din(new_new_n7198__), .dout(G5261));
  not1  g3002(.din(new_new_n7199__), .dout(G5262));
  not1  g3003(.din(new_new_n4372__), .dout(G5263));
  not1  g3004(.din(new_new_n4381__), .dout(G5264));
  buf1  g3005(.din(new_new_n4391__), .dout(G5265));
  buf1  g3006(.din(new_new_n4401__), .dout(G5266));
  buf1  g3007(.din(new_new_n4410__), .dout(G5267));
  buf1  g3008(.din(new_new_n4419__), .dout(G5268));
  buf1  g3009(.din(new_new_n4428__), .dout(G5269));
  not1  g3010(.din(new_new_n4437__), .dout(G5270));
  buf1  g3011(.din(new_new_n4446__), .dout(G5271));
  buf1  g3012(.din(new_new_n4455__), .dout(G5272));
  buf1  g3013(.din(new_new_n4464__), .dout(G5273));
  not1  g3014(.din(new_new_n4473__), .dout(G5274));
  buf1  g3015(.din(new_new_n4483__), .dout(G5275));
  not1  g3016(.din(new_new_n4493__), .dout(G5276));
  buf1  g3017(.din(new_new_n4503__), .dout(G5277));
  buf1  g3018(.din(new_new_n4513__), .dout(G5278));
  buf1  g3019(.din(new_new_n4523__), .dout(G5279));
  not1  g3020(.din(new_new_n4533__), .dout(G5280));
  buf1  g3021(.din(new_new_n4543__), .dout(G5281));
  buf1  g3022(.din(new_new_n4553__), .dout(G5282));
  buf1  g3023(.din(new_new_n4570__), .dout(G5283));
  buf1  g3024(.din(new_new_n4573__), .dout(G5284));
  not1  g3025(.din(new_new_n7209__), .dout(G5285));
  not1  g3026(.din(new_new_n7219__), .dout(G5286));
  not1  g3027(.din(new_new_n7229__), .dout(G5287));
  not1  g3028(.din(new_new_n7239__), .dout(G5288));
  not1  g3029(.din(new_new_n4594__), .dout(G5289));
  not1  g3030(.din(new_new_n7205__), .dout(G5290));
  not1  g3031(.din(new_new_n7215__), .dout(G5291));
  not1  g3032(.din(new_new_n7225__), .dout(G5292));
  not1  g3033(.din(new_new_n7235__), .dout(G5293));
  buf1  g3034(.din(new_new_n4622__), .dout(G5294));
  buf1  g3035(.din(new_new_n4631__), .dout(G5295));
  buf1  g3036(.din(new_new_n4640__), .dout(G5296));
  buf1  g3037(.din(new_new_n4649__), .dout(G5297));
  buf1  g3038(.din(new_new_n4658__), .dout(G5298));
  buf1  g3039(.din(new_new_n4667__), .dout(G5299));
  buf1  g3040(.din(new_new_n4676__), .dout(G5300));
  buf1  g3041(.din(new_new_n4685__), .dout(G5301));
  buf1  g3042(.din(new_new_n4695__), .dout(G5302));
  buf1  g3043(.din(new_new_n4705__), .dout(G5303));
  buf1  g3044(.din(new_new_n4715__), .dout(G5304));
  buf1  g3045(.din(new_new_n4725__), .dout(G5305));
  buf1  g3046(.din(new_new_n4735__), .dout(G5306));
  buf1  g3047(.din(new_new_n4745__), .dout(G5307));
  buf1  g3048(.din(new_new_n4755__), .dout(G5308));
  buf1  g3049(.din(new_new_n4765__), .dout(G5309));
  buf1  g3050(.din(new_new_n4769__), .dout(G5310));
  buf1  g3051(.din(new_new_n4774__), .dout(G5311));
  not1  g3052(.din(new_new_n4787__), .dout(G5312));
  not1  g3053(.din(new_new_n4796__), .dout(G5313));
  buf1  g3054(.din(new_new_n4806__), .dout(G5314));
  buf1  g3055(.din(new_new_n4816__), .dout(G5315));
  buf1  g3056(.din(new_new_n2042__), .dout(n11762));
  buf1  g3057(.din(new_new_n2398__), .dout(n11765));
  buf1  g3058(.din(new_new_n2400__), .dout(n11768));
  buf1  g3059(.din(new_new_n2402__), .dout(n11771));
  buf1  g3060(.din(new_new_n2044__), .dout(n11774));
  buf1  g3061(.din(new_new_n2406__), .dout(n11777));
  buf1  g3062(.din(new_new_n2408__), .dout(n11780));
  buf1  g3063(.din(new_new_n2046__), .dout(n11783));
  buf1  g3064(.din(new_new_n2412__), .dout(n11786));
  buf1  g3065(.din(new_new_n2414__), .dout(n11789));
  buf1  g3066(.din(new_new_n2416__), .dout(n11792));
  buf1  g3067(.din(new_new_n2048__), .dout(n11795));
  buf1  g3068(.din(new_new_n2420__), .dout(n11798));
  buf1  g3069(.din(new_new_n2422__), .dout(n11801));
  buf1  g3070(.din(new_new_n2424__), .dout(n11804));
  buf1  g3071(.din(new_new_n2050__), .dout(n11807));
  buf1  g3072(.din(new_new_n2428__), .dout(n11810));
  buf1  g3073(.din(new_new_n2430__), .dout(n11813));
  buf1  g3074(.din(new_new_n2432__), .dout(n11816));
  buf1  g3075(.din(new_new_n2052__), .dout(n11819));
  buf1  g3076(.din(new_new_n2436__), .dout(n11822));
  buf1  g3077(.din(new_new_n2438__), .dout(n11825));
  buf1  g3078(.din(new_new_n2440__), .dout(n11828));
  buf1  g3079(.din(new_new_n2054__), .dout(n11831));
  buf1  g3080(.din(new_new_n2444__), .dout(n11834));
  buf1  g3081(.din(new_new_n2446__), .dout(n11837));
  buf1  g3082(.din(new_new_n2448__), .dout(n11840));
  buf1  g3083(.din(new_new_n2056__), .dout(n11843));
  buf1  g3084(.din(new_new_n2452__), .dout(n11846));
  buf1  g3085(.din(new_new_n2454__), .dout(n11849));
  buf1  g3086(.din(new_new_n2456__), .dout(n11852));
  buf1  g3087(.din(new_new_n2058__), .dout(n11855));
  buf1  g3088(.din(new_new_n2460__), .dout(n11858));
  buf1  g3089(.din(new_new_n2462__), .dout(n11861));
  buf1  g3090(.din(new_new_n2464__), .dout(n11864));
  buf1  g3091(.din(new_new_n2060__), .dout(n11867));
  buf1  g3092(.din(new_new_n2468__), .dout(n11870));
  buf1  g3093(.din(new_new_n2470__), .dout(n11873));
  buf1  g3094(.din(new_new_n2472__), .dout(n11876));
  buf1  g3095(.din(new_new_n2062__), .dout(n11879));
  buf1  g3096(.din(new_new_n2476__), .dout(n11882));
  buf1  g3097(.din(new_new_n2478__), .dout(n11885));
  buf1  g3098(.din(new_new_n2480__), .dout(n11888));
  buf1  g3099(.din(new_new_n2064__), .dout(n11891));
  buf1  g3100(.din(new_new_n2484__), .dout(n11894));
  buf1  g3101(.din(new_new_n2486__), .dout(n11897));
  buf1  g3102(.din(new_new_n2488__), .dout(n11900));
  buf1  g3103(.din(new_new_n2066__), .dout(n11903));
  buf1  g3104(.din(new_new_n2492__), .dout(n11906));
  buf1  g3105(.din(new_new_n2494__), .dout(n11909));
  buf1  g3106(.din(new_new_n2496__), .dout(n11912));
  buf1  g3107(.din(new_new_n2068__), .dout(n11915));
  buf1  g3108(.din(new_new_n2500__), .dout(n11918));
  buf1  g3109(.din(new_new_n2502__), .dout(n11921));
  buf1  g3110(.din(new_new_n2504__), .dout(n11924));
  buf1  g3111(.din(new_new_n2070__), .dout(n11927));
  buf1  g3112(.din(new_new_n2508__), .dout(n11930));
  buf1  g3113(.din(new_new_n2510__), .dout(n11933));
  buf1  g3114(.din(new_new_n2512__), .dout(n11936));
  buf1  g3115(.din(new_new_n2072__), .dout(n11939));
  buf1  g3116(.din(new_new_n2516__), .dout(n11942));
  buf1  g3117(.din(new_new_n2518__), .dout(n11945));
  buf1  g3118(.din(new_new_n2520__), .dout(n11948));
  buf1  g3119(.din(new_new_n2074__), .dout(n11951));
  buf1  g3120(.din(new_new_n2524__), .dout(n11954));
  buf1  g3121(.din(new_new_n2526__), .dout(n11957));
  buf1  g3122(.din(new_new_n2528__), .dout(n11960));
  buf1  g3123(.din(new_new_n2076__), .dout(n11963));
  buf1  g3124(.din(new_new_n2532__), .dout(n11966));
  buf1  g3125(.din(new_new_n2534__), .dout(n11969));
  buf1  g3126(.din(new_new_n2536__), .dout(n11972));
  buf1  g3127(.din(new_new_n2078__), .dout(n11975));
  buf1  g3128(.din(new_new_n2540__), .dout(n11978));
  buf1  g3129(.din(new_new_n2542__), .dout(n11981));
  buf1  g3130(.din(new_new_n2080__), .dout(n11984));
  buf1  g3131(.din(new_new_n2546__), .dout(n11987));
  buf1  g3132(.din(new_new_n2548__), .dout(n11990));
  buf1  g3133(.din(new_new_n2550__), .dout(n11993));
  buf1  g3134(.din(new_new_n2082__), .dout(n11996));
  buf1  g3135(.din(new_new_n2554__), .dout(n11999));
  buf1  g3136(.din(new_new_n2556__), .dout(n12002));
  buf1  g3137(.din(new_new_n2084__), .dout(n12005));
  buf1  g3138(.din(new_new_n2560__), .dout(n12008));
  buf1  g3139(.din(new_new_n2562__), .dout(n12011));
  buf1  g3140(.din(new_new_n2564__), .dout(n12014));
  buf1  g3141(.din(new_new_n2086__), .dout(n12017));
  buf1  g3142(.din(new_new_n2568__), .dout(n12020));
  buf1  g3143(.din(new_new_n2570__), .dout(n12023));
  buf1  g3144(.din(new_new_n2572__), .dout(n12026));
  buf1  g3145(.din(new_new_n2088__), .dout(n12029));
  buf1  g3146(.din(new_new_n2576__), .dout(n12032));
  buf1  g3147(.din(new_new_n2578__), .dout(n12035));
  buf1  g3148(.din(new_new_n2580__), .dout(n12038));
  buf1  g3149(.din(new_new_n2090__), .dout(n12041));
  buf1  g3150(.din(new_new_n2584__), .dout(n12044));
  buf1  g3151(.din(new_new_n2586__), .dout(n12047));
  buf1  g3152(.din(new_new_n2588__), .dout(n12050));
  buf1  g3153(.din(new_new_n2092__), .dout(n12053));
  buf1  g3154(.din(new_new_n2592__), .dout(n12056));
  buf1  g3155(.din(new_new_n2594__), .dout(n12059));
  buf1  g3156(.din(new_new_n2596__), .dout(n12062));
  buf1  g3157(.din(new_new_n2094__), .dout(n12065));
  buf1  g3158(.din(new_new_n2600__), .dout(n12068));
  buf1  g3159(.din(new_new_n2602__), .dout(n12071));
  buf1  g3160(.din(new_new_n2604__), .dout(n12074));
  buf1  g3161(.din(new_new_n2096__), .dout(n12077));
  buf1  g3162(.din(new_new_n2608__), .dout(n12080));
  buf1  g3163(.din(new_new_n2610__), .dout(n12083));
  buf1  g3164(.din(new_new_n2612__), .dout(n12086));
  buf1  g3165(.din(new_new_n2098__), .dout(n12089));
  buf1  g3166(.din(new_new_n2616__), .dout(n12092));
  buf1  g3167(.din(new_new_n2618__), .dout(n12095));
  buf1  g3168(.din(new_new_n2620__), .dout(n12098));
  buf1  g3169(.din(new_new_n2100__), .dout(n12101));
  buf1  g3170(.din(new_new_n2624__), .dout(n12104));
  buf1  g3171(.din(new_new_n2626__), .dout(n12107));
  buf1  g3172(.din(new_new_n2628__), .dout(n12110));
  buf1  g3173(.din(new_new_n2102__), .dout(n12113));
  buf1  g3174(.din(new_new_n2632__), .dout(n12116));
  buf1  g3175(.din(new_new_n2634__), .dout(n12119));
  buf1  g3176(.din(new_new_n2636__), .dout(n12122));
  buf1  g3177(.din(new_new_n2104__), .dout(n12125));
  buf1  g3178(.din(new_new_n2640__), .dout(n12128));
  buf1  g3179(.din(new_new_n2642__), .dout(n12131));
  buf1  g3180(.din(new_new_n2644__), .dout(n12134));
  buf1  g3181(.din(new_new_n2106__), .dout(n12137));
  buf1  g3182(.din(new_new_n2648__), .dout(n12140));
  buf1  g3183(.din(new_new_n2650__), .dout(n12143));
  buf1  g3184(.din(new_new_n2652__), .dout(n12146));
  buf1  g3185(.din(new_new_n2108__), .dout(n12149));
  buf1  g3186(.din(new_new_n2656__), .dout(n12152));
  buf1  g3187(.din(new_new_n2658__), .dout(n12155));
  buf1  g3188(.din(new_new_n2660__), .dout(n12158));
  buf1  g3189(.din(new_new_n2110__), .dout(n12161));
  buf1  g3190(.din(new_new_n2664__), .dout(n12164));
  buf1  g3191(.din(new_new_n2666__), .dout(n12167));
  buf1  g3192(.din(new_new_n2668__), .dout(n12170));
  buf1  g3193(.din(new_new_n2112__), .dout(n12173));
  buf1  g3194(.din(new_new_n2672__), .dout(n12176));
  buf1  g3195(.din(new_new_n2674__), .dout(n12179));
  buf1  g3196(.din(new_new_n2676__), .dout(n12182));
  buf1  g3197(.din(new_new_n2114__), .dout(n12185));
  buf1  g3198(.din(new_new_n2680__), .dout(n12188));
  buf1  g3199(.din(new_new_n2682__), .dout(n12191));
  buf1  g3200(.din(new_new_n2684__), .dout(n12194));
  buf1  g3201(.din(new_new_n2116__), .dout(n12197));
  buf1  g3202(.din(new_new_n2688__), .dout(n12200));
  buf1  g3203(.din(new_new_n2690__), .dout(n12203));
  buf1  g3204(.din(new_new_n2692__), .dout(n12206));
  buf1  g3205(.din(new_new_n2118__), .dout(n12209));
  buf1  g3206(.din(new_new_n2696__), .dout(n12212));
  buf1  g3207(.din(new_new_n2698__), .dout(n12215));
  buf1  g3208(.din(new_new_n2700__), .dout(n12218));
  buf1  g3209(.din(new_new_n2120__), .dout(n12221));
  buf1  g3210(.din(new_new_n2704__), .dout(n12224));
  buf1  g3211(.din(new_new_n2706__), .dout(n12227));
  buf1  g3212(.din(new_new_n2708__), .dout(n12230));
  buf1  g3213(.din(new_new_n2122__), .dout(n12233));
  buf1  g3214(.din(new_new_n2712__), .dout(n12236));
  buf1  g3215(.din(new_new_n2714__), .dout(n12239));
  buf1  g3216(.din(new_new_n2716__), .dout(n12242));
  buf1  g3217(.din(new_new_n2124__), .dout(n12245));
  buf1  g3218(.din(new_new_n2720__), .dout(n12248));
  buf1  g3219(.din(new_new_n2722__), .dout(n12251));
  buf1  g3220(.din(new_new_n2724__), .dout(n12254));
  buf1  g3221(.din(new_new_n2126__), .dout(n12257));
  buf1  g3222(.din(new_new_n2728__), .dout(n12260));
  buf1  g3223(.din(new_new_n2730__), .dout(n12263));
  buf1  g3224(.din(new_new_n2128__), .dout(n12266));
  buf1  g3225(.din(new_new_n2734__), .dout(n12269));
  buf1  g3226(.din(new_new_n2736__), .dout(n12272));
  buf1  g3227(.din(new_new_n2130__), .dout(n12275));
  buf1  g3228(.din(new_new_n2740__), .dout(n12278));
  buf1  g3229(.din(new_new_n2742__), .dout(n12281));
  buf1  g3230(.din(new_new_n2744__), .dout(n12284));
  buf1  g3231(.din(new_new_n2132__), .dout(n12287));
  buf1  g3232(.din(new_new_n2748__), .dout(n12290));
  buf1  g3233(.din(new_new_n2750__), .dout(n12293));
  buf1  g3234(.din(new_new_n2134__), .dout(n12296));
  buf1  g3235(.din(new_new_n2754__), .dout(n12299));
  buf1  g3236(.din(new_new_n2756__), .dout(n12302));
  buf1  g3237(.din(new_new_n2136__), .dout(n12305));
  buf1  g3238(.din(new_new_n2760__), .dout(n12308));
  buf1  g3239(.din(new_new_n2762__), .dout(n12311));
  buf1  g3240(.din(new_new_n2138__), .dout(n12314));
  buf1  g3241(.din(new_new_n2766__), .dout(n12317));
  buf1  g3242(.din(new_new_n2768__), .dout(n12320));
  buf1  g3243(.din(new_new_n2770__), .dout(n12323));
  buf1  g3244(.din(new_new_n2140__), .dout(n12326));
  buf1  g3245(.din(new_new_n2774__), .dout(n12329));
  buf1  g3246(.din(new_new_n2776__), .dout(n12332));
  buf1  g3247(.din(new_new_n2142__), .dout(n12335));
  buf1  g3248(.din(new_new_n2780__), .dout(n12338));
  buf1  g3249(.din(new_new_n2782__), .dout(n12341));
  buf1  g3250(.din(new_new_n2784__), .dout(n12344));
  buf1  g3251(.din(new_new_n2144__), .dout(n12347));
  buf1  g3252(.din(new_new_n2788__), .dout(n12350));
  buf1  g3253(.din(new_new_n2790__), .dout(n12353));
  buf1  g3254(.din(new_new_n2146__), .dout(n12356));
  buf1  g3255(.din(new_new_n2794__), .dout(n12359));
  buf1  g3256(.din(new_new_n2796__), .dout(n12362));
  buf1  g3257(.din(new_new_n2798__), .dout(n12365));
  buf1  g3258(.din(new_new_n2148__), .dout(n12368));
  buf1  g3259(.din(new_new_n2802__), .dout(n12371));
  buf1  g3260(.din(new_new_n2804__), .dout(n12374));
  buf1  g3261(.din(new_new_n7547__), .dout(n12377));
  buf1  g3262(.din(new_new_n2150__), .dout(n12380));
  buf1  g3263(.din(new_new_n2810__), .dout(n12383));
  buf1  g3264(.din(new_new_n2812__), .dout(n12386));
  buf1  g3265(.din(new_new_n2814__), .dout(n12389));
  buf1  g3266(.din(new_new_n2152__), .dout(n12392));
  buf1  g3267(.din(new_new_n2818__), .dout(n12395));
  buf1  g3268(.din(new_new_n2820__), .dout(n12398));
  buf1  g3269(.din(new_new_n2822__), .dout(n12401));
  buf1  g3270(.din(new_new_n2154__), .dout(n12404));
  buf1  g3271(.din(new_new_n2826__), .dout(n12407));
  buf1  g3272(.din(new_new_n2828__), .dout(n12410));
  buf1  g3273(.din(new_new_n2156__), .dout(n12413));
  buf1  g3274(.din(new_new_n2832__), .dout(n12416));
  buf1  g3275(.din(new_new_n2834__), .dout(n12419));
  buf1  g3276(.din(new_new_n2158__), .dout(n12422));
  buf1  g3277(.din(new_new_n2838__), .dout(n12425));
  buf1  g3278(.din(new_new_n2840__), .dout(n12428));
  buf1  g3279(.din(new_new_n2160__), .dout(n12431));
  buf1  g3280(.din(new_new_n2844__), .dout(n12434));
  buf1  g3281(.din(new_new_n2846__), .dout(n12437));
  buf1  g3282(.din(new_new_n2162__), .dout(n12440));
  buf1  g3283(.din(new_new_n2850__), .dout(n12443));
  buf1  g3284(.din(new_new_n2852__), .dout(n12446));
  buf1  g3285(.din(new_new_n2854__), .dout(n12449));
  buf1  g3286(.din(new_new_n2164__), .dout(n12452));
  buf1  g3287(.din(new_new_n2858__), .dout(n12455));
  buf1  g3288(.din(new_new_n2860__), .dout(n12458));
  buf1  g3289(.din(new_new_n2862__), .dout(n12461));
  buf1  g3290(.din(new_new_n2166__), .dout(n12464));
  buf1  g3291(.din(new_new_n2866__), .dout(n12467));
  buf1  g3292(.din(new_new_n2868__), .dout(n12470));
  buf1  g3293(.din(new_new_n2870__), .dout(n12473));
  buf1  g3294(.din(new_new_n2168__), .dout(n12476));
  buf1  g3295(.din(new_new_n2874__), .dout(n12479));
  buf1  g3296(.din(new_new_n2876__), .dout(n12482));
  buf1  g3297(.din(new_new_n2878__), .dout(n12485));
  buf1  g3298(.din(new_new_n2170__), .dout(n12488));
  buf1  g3299(.din(new_new_n2882__), .dout(n12491));
  buf1  g3300(.din(new_new_n2884__), .dout(n12494));
  buf1  g3301(.din(new_new_n2886__), .dout(n12497));
  buf1  g3302(.din(new_new_n2172__), .dout(n12500));
  buf1  g3303(.din(new_new_n2890__), .dout(n12503));
  buf1  g3304(.din(new_new_n2892__), .dout(n12506));
  buf1  g3305(.din(new_new_n2894__), .dout(n12509));
  buf1  g3306(.din(new_new_n2174__), .dout(n12512));
  buf1  g3307(.din(new_new_n2898__), .dout(n12515));
  buf1  g3308(.din(new_new_n2900__), .dout(n12518));
  buf1  g3309(.din(new_new_n2902__), .dout(n12521));
  buf1  g3310(.din(new_new_n2176__), .dout(n12524));
  buf1  g3311(.din(new_new_n2906__), .dout(n12527));
  buf1  g3312(.din(new_new_n2908__), .dout(n12530));
  buf1  g3313(.din(new_new_n2910__), .dout(n12533));
  buf1  g3314(.din(new_new_n2178__), .dout(n12536));
  buf1  g3315(.din(new_new_n2914__), .dout(n12539));
  buf1  g3316(.din(new_new_n2916__), .dout(n12542));
  buf1  g3317(.din(new_new_n2918__), .dout(n12545));
  buf1  g3318(.din(new_new_n2180__), .dout(n12548));
  buf1  g3319(.din(new_new_n2922__), .dout(n12551));
  buf1  g3320(.din(new_new_n2924__), .dout(n12554));
  buf1  g3321(.din(new_new_n2926__), .dout(n12557));
  buf1  g3322(.din(new_new_n2182__), .dout(n12560));
  buf1  g3323(.din(new_new_n2930__), .dout(n12563));
  buf1  g3324(.din(new_new_n2932__), .dout(n12566));
  buf1  g3325(.din(new_new_n2934__), .dout(n12569));
  buf1  g3326(.din(new_new_n2184__), .dout(n12572));
  buf1  g3327(.din(new_new_n2938__), .dout(n12575));
  buf1  g3328(.din(new_new_n2940__), .dout(n12578));
  buf1  g3329(.din(new_new_n2942__), .dout(n12581));
  buf1  g3330(.din(new_new_n2186__), .dout(n12584));
  buf1  g3331(.din(new_new_n2946__), .dout(n12587));
  buf1  g3332(.din(new_new_n2948__), .dout(n12590));
  buf1  g3333(.din(new_new_n2950__), .dout(n12593));
  buf1  g3334(.din(new_new_n2188__), .dout(n12596));
  buf1  g3335(.din(new_new_n2954__), .dout(n12599));
  buf1  g3336(.din(new_new_n2956__), .dout(n12602));
  buf1  g3337(.din(new_new_n2958__), .dout(n12605));
  buf1  g3338(.din(new_new_n2190__), .dout(n12608));
  buf1  g3339(.din(new_new_n2962__), .dout(n12611));
  buf1  g3340(.din(new_new_n2964__), .dout(n12614));
  buf1  g3341(.din(new_new_n2966__), .dout(n12617));
  buf1  g3342(.din(new_new_n2192__), .dout(n12620));
  buf1  g3343(.din(new_new_n2970__), .dout(n12623));
  buf1  g3344(.din(new_new_n2972__), .dout(n12626));
  buf1  g3345(.din(new_new_n2974__), .dout(n12629));
  buf1  g3346(.din(new_new_n2194__), .dout(n12632));
  buf1  g3347(.din(new_new_n2978__), .dout(n12635));
  buf1  g3348(.din(new_new_n2980__), .dout(n12638));
  buf1  g3349(.din(new_new_n2982__), .dout(n12641));
  buf1  g3350(.din(new_new_n2196__), .dout(n12644));
  buf1  g3351(.din(new_new_n2986__), .dout(n12647));
  buf1  g3352(.din(new_new_n2988__), .dout(n12650));
  buf1  g3353(.din(new_new_n2990__), .dout(n12653));
  buf1  g3354(.din(new_new_n2198__), .dout(n12656));
  buf1  g3355(.din(new_new_n2994__), .dout(n12659));
  buf1  g3356(.din(new_new_n2996__), .dout(n12662));
  buf1  g3357(.din(new_new_n2998__), .dout(n12665));
  buf1  g3358(.din(new_new_n2200__), .dout(n12668));
  buf1  g3359(.din(new_new_n3002__), .dout(n12671));
  buf1  g3360(.din(new_new_n3004__), .dout(n12674));
  buf1  g3361(.din(new_new_n3006__), .dout(n12677));
  buf1  g3362(.din(new_new_n2202__), .dout(n12680));
  buf1  g3363(.din(new_new_n3010__), .dout(n12683));
  buf1  g3364(.din(new_new_n3012__), .dout(n12686));
  buf1  g3365(.din(new_new_n3014__), .dout(n12689));
  buf1  g3366(.din(new_new_n2204__), .dout(n12692));
  buf1  g3367(.din(new_new_n3018__), .dout(n12695));
  buf1  g3368(.din(new_new_n3020__), .dout(n12698));
  buf1  g3369(.din(new_new_n3022__), .dout(n12701));
  buf1  g3370(.din(new_new_n2206__), .dout(n12704));
  buf1  g3371(.din(new_new_n3026__), .dout(n12707));
  buf1  g3372(.din(new_new_n3028__), .dout(n12710));
  buf1  g3373(.din(new_new_n3030__), .dout(n12713));
  buf1  g3374(.din(new_new_n2208__), .dout(n12716));
  buf1  g3375(.din(new_new_n3034__), .dout(n12719));
  buf1  g3376(.din(new_new_n3036__), .dout(n12722));
  buf1  g3377(.din(new_new_n3038__), .dout(n12725));
  buf1  g3378(.din(new_new_n2210__), .dout(n12728));
  buf1  g3379(.din(new_new_n3042__), .dout(n12731));
  buf1  g3380(.din(new_new_n3044__), .dout(n12734));
  buf1  g3381(.din(new_new_n3046__), .dout(n12737));
  buf1  g3382(.din(new_new_n2212__), .dout(n12740));
  buf1  g3383(.din(new_new_n3050__), .dout(n12743));
  buf1  g3384(.din(new_new_n3052__), .dout(n12746));
  buf1  g3385(.din(new_new_n3054__), .dout(n12749));
  buf1  g3386(.din(new_new_n2214__), .dout(n12752));
  buf1  g3387(.din(new_new_n3058__), .dout(n12755));
  buf1  g3388(.din(new_new_n3060__), .dout(n12758));
  buf1  g3389(.din(new_new_n3062__), .dout(n12761));
  buf1  g3390(.din(new_new_n2216__), .dout(n12764));
  buf1  g3391(.din(new_new_n2218__), .dout(n12767));
  buf1  g3392(.din(new_new_n2232__), .dout(n12770));
  buf1  g3393(.din(new_new_n2234__), .dout(n12773));
  buf1  g3394(.din(new_new_n2236__), .dout(n12776));
  buf1  g3395(.din(new_new_n2238__), .dout(n12779));
  buf1  g3396(.din(new_new_n3076__), .dout(n12782));
  buf1  g3397(.din(new_new_n3078__), .dout(n12785));
  buf1  g3398(.din(new_new_n3080__), .dout(n12788));
  buf1  g3399(.din(new_new_n2240__), .dout(n12791));
  buf1  g3400(.din(new_new_n2242__), .dout(n12794));
  buf1  g3401(.din(new_new_n2244__), .dout(n12797));
  buf1  g3402(.din(new_new_n2246__), .dout(n12800));
  buf1  g3403(.din(new_new_n2248__), .dout(n12803));
  buf1  g3404(.din(new_new_n2262__), .dout(n12806));
  buf1  g3405(.din(new_new_n3094__), .dout(n12809));
  buf1  g3406(.din(new_new_n3096__), .dout(n12812));
  buf1  g3407(.din(new_new_n2264__), .dout(n12815));
  buf1  g3408(.din(new_new_n3100__), .dout(n12818));
  buf1  g3409(.din(new_new_n3102__), .dout(n12821));
  buf1  g3410(.din(new_new_n2266__), .dout(n12824));
  buf1  g3411(.din(new_new_n3106__), .dout(n12827));
  buf1  g3412(.din(new_new_n7686__), .dout(n12830));
  buf1  g3413(.din(new_new_n2268__), .dout(n12833));
  buf1  g3414(.din(new_new_n3112__), .dout(n12836));
  buf1  g3415(.din(new_new_n3712__), .dout(n12839));
  buf1  g3416(.din(new_new_n2270__), .dout(n12842));
  buf1  g3417(.din(new_new_n2272__), .dout(n12845));
  buf1  g3418(.din(new_new_n2282__), .dout(n12848));
  buf1  g3419(.din(new_new_n2284__), .dout(n12851));
  buf1  g3420(.din(new_new_n2290__), .dout(n12854));
  buf1  g3421(.din(new_new_n3538__), .dout(n12857));
  buf1  g3422(.din(new_new_n2292__), .dout(n12860));
  buf1  g3423(.din(new_new_n2294__), .dout(n12863));
  buf1  g3424(.din(new_new_n3514__), .dout(n12866));
  buf1  g3425(.din(new_new_n3498__), .dout(n12869));
  buf1  g3426(.din(new_new_n2300__), .dout(n12872));
  buf1  g3427(.din(new_new_n2302__), .dout(n12875));
  buf1  g3428(.din(new_new_n3542__), .dout(n12878));
  buf1  g3429(.din(new_new_n2304__), .dout(n12881));
  buf1  g3430(.din(new_new_n3144__), .dout(n12884));
  buf1  g3431(.din(new_new_n3146__), .dout(n12887));
  buf1  g3432(.din(new_new_n2306__), .dout(n12890));
  buf1  g3433(.din(new_new_n3150__), .dout(n12893));
  buf1  g3434(.din(new_new_n3152__), .dout(n12896));
  buf1  g3435(.din(new_new_n2308__), .dout(n12899));
  buf1  g3436(.din(new_new_n3156__), .dout(n12902));
  buf1  g3437(.din(new_new_n3158__), .dout(n12905));
  buf1  g3438(.din(new_new_n3160__), .dout(n12908));
  buf1  g3439(.din(new_new_n2312__), .dout(n12911));
  buf1  g3440(.din(new_new_n3164__), .dout(n12914));
  buf1  g3441(.din(new_new_n3166__), .dout(n12917));
  buf1  g3442(.din(new_new_n3168__), .dout(n12920));
  buf1  g3443(.din(new_new_n2314__), .dout(n12923));
  buf1  g3444(.din(new_new_n2316__), .dout(n12926));
  buf1  g3445(.din(new_new_n2322__), .dout(n12929));
  buf1  g3446(.din(new_new_n3176__), .dout(n12932));
  buf1  g3447(.din(new_new_n2324__), .dout(n12935));
  buf1  g3448(.din(new_new_n2326__), .dout(n12938));
  buf1  g3449(.din(new_new_n2332__), .dout(n12941));
  buf1  g3450(.din(new_new_n2334__), .dout(n12944));
  buf1  g3451(.din(new_new_n2336__), .dout(n12947));
  buf1  g3452(.din(new_new_n2338__), .dout(n12950));
  buf1  g3453(.din(new_new_n2340__), .dout(n12953));
  buf1  g3454(.din(new_new_n2342__), .dout(n12956));
  buf1  g3455(.din(new_new_n3194__), .dout(n12959));
  buf1  g3456(.din(new_new_n3196__), .dout(n12962));
  buf1  g3457(.din(new_new_n3198__), .dout(n12965));
  buf1  g3458(.din(new_new_n2344__), .dout(n12968));
  buf1  g3459(.din(new_new_n3202__), .dout(n12971));
  buf1  g3460(.din(new_new_n3204__), .dout(n12974));
  buf1  g3461(.din(new_new_n3206__), .dout(n12977));
  buf1  g3462(.din(new_new_n2346__), .dout(n12980));
  buf1  g3463(.din(new_new_n3210__), .dout(n12983));
  buf1  g3464(.din(new_new_n3212__), .dout(n12986));
  buf1  g3465(.din(new_new_n3214__), .dout(n12989));
  buf1  g3466(.din(new_new_n2348__), .dout(n12992));
  buf1  g3467(.din(new_new_n3218__), .dout(n12995));
  buf1  g3468(.din(new_new_n3220__), .dout(n12998));
  buf1  g3469(.din(new_new_n3222__), .dout(n13001));
  buf1  g3470(.din(new_new_n2350__), .dout(n13004));
  buf1  g3471(.din(new_new_n3226__), .dout(n13007));
  buf1  g3472(.din(new_new_n3228__), .dout(n13010));
  buf1  g3473(.din(new_new_n3230__), .dout(n13013));
  buf1  g3474(.din(new_new_n2352__), .dout(n13016));
  buf1  g3475(.din(new_new_n3234__), .dout(n13019));
  buf1  g3476(.din(new_new_n3236__), .dout(n13022));
  buf1  g3477(.din(new_new_n3238__), .dout(n13025));
  buf1  g3478(.din(new_new_n2354__), .dout(n13028));
  buf1  g3479(.din(new_new_n3242__), .dout(n13031));
  buf1  g3480(.din(new_new_n3244__), .dout(n13034));
  buf1  g3481(.din(new_new_n2356__), .dout(n13037));
  buf1  g3482(.din(new_new_n3248__), .dout(n13040));
  buf1  g3483(.din(new_new_n3250__), .dout(n13043));
  buf1  g3484(.din(new_new_n3252__), .dout(n13046));
  buf1  g3485(.din(new_new_n2358__), .dout(n13049));
  buf1  g3486(.din(new_new_n3256__), .dout(n13052));
  buf1  g3487(.din(new_new_n3258__), .dout(n13055));
  buf1  g3488(.din(new_new_n3260__), .dout(n13058));
  buf1  g3489(.din(new_new_n2360__), .dout(n13061));
  buf1  g3490(.din(new_new_n3264__), .dout(n13064));
  buf1  g3491(.din(new_new_n3266__), .dout(n13067));
  buf1  g3492(.din(new_new_n3268__), .dout(n13070));
  buf1  g3493(.din(new_new_n2362__), .dout(n13073));
  buf1  g3494(.din(new_new_n3272__), .dout(n13076));
  buf1  g3495(.din(new_new_n3274__), .dout(n13079));
  buf1  g3496(.din(new_new_n3276__), .dout(n13082));
  buf1  g3497(.din(new_new_n2364__), .dout(n13085));
  buf1  g3498(.din(new_new_n3280__), .dout(n13088));
  buf1  g3499(.din(new_new_n2366__), .dout(n13091));
  buf1  g3500(.din(new_new_n3284__), .dout(n13094));
  buf1  g3501(.din(new_new_n3286__), .dout(n13097));
  buf1  g3502(.din(new_new_n3288__), .dout(n13100));
  buf1  g3503(.din(new_new_n2368__), .dout(n13103));
  buf1  g3504(.din(new_new_n3292__), .dout(n13106));
  buf1  g3505(.din(new_new_n3294__), .dout(n13109));
  buf1  g3506(.din(new_new_n3296__), .dout(n13112));
  buf1  g3507(.din(new_new_n2370__), .dout(n13115));
  buf1  g3508(.din(new_new_n3300__), .dout(n13118));
  buf1  g3509(.din(new_new_n3302__), .dout(n13121));
  buf1  g3510(.din(new_new_n3304__), .dout(n13124));
  buf1  g3511(.din(new_new_n2372__), .dout(n13127));
  buf1  g3512(.din(new_new_n3308__), .dout(n13130));
  buf1  g3513(.din(new_new_n3310__), .dout(n13133));
  buf1  g3514(.din(new_new_n2374__), .dout(n13136));
  buf1  g3515(.din(new_new_n3314__), .dout(n13139));
  buf1  g3516(.din(new_new_n3316__), .dout(n13142));
  buf1  g3517(.din(new_new_n2376__), .dout(n13145));
  buf1  g3518(.din(new_new_n3320__), .dout(n13148));
  buf1  g3519(.din(new_new_n3322__), .dout(n13151));
  buf1  g3520(.din(new_new_n2378__), .dout(n13154));
  buf1  g3521(.din(new_new_n3326__), .dout(n13157));
  buf1  g3522(.din(new_new_n3328__), .dout(n13160));
  buf1  g3523(.din(new_new_n2380__), .dout(n13163));
  buf1  g3524(.din(new_new_n3332__), .dout(n13166));
  buf1  g3525(.din(new_new_n3334__), .dout(n13169));
  buf1  g3526(.din(new_new_n3336__), .dout(n13172));
  buf1  g3527(.din(new_new_n2382__), .dout(n13175));
  buf1  g3528(.din(new_new_n3340__), .dout(n13178));
  buf1  g3529(.din(new_new_n3342__), .dout(n13181));
  buf1  g3530(.din(new_new_n3344__), .dout(n13184));
  buf1  g3531(.din(new_new_n2384__), .dout(n13187));
  buf1  g3532(.din(new_new_n3348__), .dout(n13190));
  buf1  g3533(.din(new_new_n3350__), .dout(n13193));
  buf1  g3534(.din(new_new_n3352__), .dout(n13196));
  buf1  g3535(.din(new_new_n2386__), .dout(n13199));
  buf1  g3536(.din(new_new_n3356__), .dout(n13202));
  buf1  g3537(.din(new_new_n3358__), .dout(n13205));
  buf1  g3538(.din(new_new_n3360__), .dout(n13208));
  buf1  g3539(.din(new_new_n2388__), .dout(n13211));
  buf1  g3540(.din(new_new_n3364__), .dout(n13214));
  buf1  g3541(.din(new_new_n3366__), .dout(n13217));
  buf1  g3542(.din(new_new_n3368__), .dout(n13220));
  buf1  g3543(.din(new_new_n2390__), .dout(n13223));
  buf1  g3544(.din(new_new_n3372__), .dout(n13226));
  buf1  g3545(.din(new_new_n3374__), .dout(n13229));
  buf1  g3546(.din(new_new_n3376__), .dout(n13232));
  buf1  g3547(.din(new_new_n2392__), .dout(n13235));
  buf1  g3548(.din(new_new_n3380__), .dout(n13238));
  buf1  g3549(.din(new_new_n3382__), .dout(n13241));
  buf1  g3550(.din(new_new_n7548__), .dout(n13244));
  buf1  g3551(.din(new_new_n2394__), .dout(n13247));
  buf1  g3552(.din(new_new_n3388__), .dout(n13250));
  buf1  g3553(.din(new_new_n3390__), .dout(n13253));
  buf1  g3554(.din(new_new_n7540__), .dout(n13256));
  buf1  g3555(.din(new_new_n2396__), .dout(n13259));
  buf1  g3556(.din(new_new_n3396__), .dout(n13262));
  buf1  g3557(.din(new_new_n3398__), .dout(n13265));
  buf1  g3558(.din(new_new_n3400__), .dout(n13268));
  buf1  g3559(.din(new_new_n3490__), .dout(n13271));
  buf1  g3560(.din(new_new_n3494__), .dout(n13274));
  buf1  g3561(.din(new_new_n3506__), .dout(n13277));
  buf1  g3562(.din(new_new_n3524__), .dout(n13280));
  buf1  g3563(.din(new_new_n3526__), .dout(n13283));
  buf1  g3564(.din(new_new_n3534__), .dout(n13286));
  buf1  g3565(.din(new_new_n3548__), .dout(n13289));
  buf1  g3566(.din(new_new_n3556__), .dout(n13292));
  buf1  g3567(.din(new_new_n3568__), .dout(n13295));
  buf1  g3568(.din(new_new_n3574__), .dout(n13298));
  buf1  g3569(.din(new_new_n3602__), .dout(n13301));
  buf1  g3570(.din(new_new_n3610__), .dout(n13304));
  buf1  g3571(.din(new_new_n7684__), .dout(n13307));
  buf1  g3572(.din(new_new_n7265__), .dout(n13310));
  buf1  g3573(.din(new_new_n7685__), .dout(n13313));
  buf1  g3574(.din(new_new_n7554__), .dout(n13316));
  buf1  g3575(.din(new_new_n3632__), .dout(n13319));
  buf1  g3576(.din(new_new_n3650__), .dout(n13322));
  buf1  g3577(.din(new_new_n3658__), .dout(n13325));
  buf1  g3578(.din(new_new_n3692__), .dout(n13328));
  buf1  g3579(.din(new_new_n3738__), .dout(n13331));
  buf1  g3580(.din(new_new_n3922__), .dout(n13334));
  buf1  g3581(.din(new_new_n3918__), .dout(n13337));
  buf1  g3582(.din(new_new_n7862__), .dout(n13340));
  buf1  g3583(.din(new_new_n7858__), .dout(n13343));
  buf1  g3584(.din(new_new_n7854__), .dout(n13346));
  buf1  g3585(.din(new_new_n7318__), .dout(n13349));
  buf1  g3586(.din(new_new_n7595__), .dout(n13352));
  buf1  g3587(.din(new_new_n7585__), .dout(n13355));
  buf1  g3588(.din(new_new_n7267__), .dout(n13358));
  buf1  g3589(.din(new_new_n7660__), .dout(n13361));
  buf1  g3590(.din(new_new_n7577__), .dout(n13364));
  buf1  g3591(.din(new_new_n7578__), .dout(n13367));
  buf1  g3592(.din(new_new_n7866__), .dout(n13370));
  buf1  g3593(.din(new_new_n7734__), .dout(n13373));
  buf1  g3594(.din(new_new_n7851__), .dout(n13376));
  buf1  g3595(.din(new_new_n7874__), .dout(n13379));
  buf1  g3596(.din(new_new_n7870__), .dout(n13382));
  buf1  g3597(.din(new_new_n7778__), .dout(n13385));
  buf1  g3598(.din(new_new_n7856__), .dout(n13388));
  buf1  g3599(.din(new_new_n7860__), .dout(n13391));
  buf1  g3600(.din(new_new_n7864__), .dout(n13394));
  buf1  g3601(.din(new_new_n7269__), .dout(n13397));
  buf1  g3602(.din(new_new_n3672__), .dout(n13400));
  buf1  g3603(.din(new_new_n3674__), .dout(n13403));
  buf1  g3604(.din(new_new_n3676__), .dout(n13406));
  buf1  g3605(.din(new_new_n7935__), .dout(n13409));
  buf1  g3606(.din(new_new_n3696__), .dout(n13412));
  buf1  g3607(.din(new_new_n7868__), .dout(n13415));
  buf1  g3608(.din(new_new_n3704__), .dout(n13418));
  buf1  g3609(.din(new_new_n3706__), .dout(n13421));
  buf1  g3610(.din(new_new_n3702__), .dout(n13424));
  buf1  g3611(.din(new_new_n3710__), .dout(n13427));
  buf1  g3612(.din(new_new_n7959__), .dout(n13430));
  buf1  g3613(.din(new_new_n7938__), .dout(n13433));
  buf1  g3614(.din(new_new_n3722__), .dout(n13436));
  buf1  g3615(.din(new_new_n7872__), .dout(n13439));
  buf1  g3616(.din(new_new_n7876__), .dout(n13442));
  buf1  g3617(.din(new_new_n7564__), .dout(n13445));
  buf1  g3618(.din(new_new_n7807__), .dout(n13448));
  buf1  g3619(.din(new_new_n3730__), .dout(n13451));
  buf1  g3620(.din(new_new_n3732__), .dout(n13454));
  buf1  g3621(.din(new_new_n3736__), .dout(n13457));
  buf1  g3622(.din(new_new_n7816__), .dout(n13460));
  buf1  g3623(.din(new_new_n7836__), .dout(n13463));
  buf1  g3624(.din(new_new_n7840__), .dout(n13466));
  buf1  g3625(.din(new_new_n7878__), .dout(n13469));
  buf1  g3626(.din(new_new_n3750__), .dout(n13472));
  buf1  g3627(.din(new_new_n7780__), .dout(n13475));
  buf1  g3628(.din(new_new_n3754__), .dout(n13478));
  buf1  g3629(.din(new_new_n7937__), .dout(n13481));
  buf1  g3630(.din(new_new_n3760__), .dout(n13484));
  buf1  g3631(.din(new_new_n3762__), .dout(n13487));
  buf1  g3632(.din(new_new_n7331__), .dout(n13490));
  buf1  g3633(.din(new_new_n3758__), .dout(n13493));
  buf1  g3634(.din(new_new_n3766__), .dout(n13496));
  buf1  g3635(.din(new_new_n3768__), .dout(n13499));
  buf1  g3636(.din(new_new_n7960__), .dout(n13502));
  buf1  g3637(.din(new_new_n7907__), .dout(n13505));
  buf1  g3638(.din(new_new_n7941__), .dout(n13508));
  buf1  g3639(.din(new_new_n3846__), .dout(n13511));
  buf1  g3640(.din(new_new_n7814__), .dout(n13514));
  buf1  g3641(.din(new_new_n3930__), .dout(n13517));
  buf1  g3642(.din(new_new_n3932__), .dout(n13520));
  buf1  g3643(.din(new_new_n7363__), .dout(n13523));
  buf1  g3644(.din(new_new_n7290__), .dout(n13526));
  buf1  g3645(.din(new_new_n7781__), .dout(n13529));
  buf1  g3646(.din(new_new_n7924__), .dout(n13532));
  buf1  g3647(.din(new_new_n7330__), .dout(n13535));
  buf1  g3648(.din(new_new_n7817__), .dout(n13538));
  buf1  g3649(.din(new_new_n7944__), .dout(n13541));
  buf1  g3650(.din(new_new_n7793__), .dout(n13544));
  buf1  g3651(.din(new_new_n3986__), .dout(n13547));
  buf1  g3652(.din(new_new_n7341__), .dout(n13550));
  buf1  g3653(.din(new_new_n3996__), .dout(n13553));
  buf1  g3654(.din(new_new_n7324__), .dout(n13556));
  not1  g3655(.din(new_new_n7613__), .dout(n13559));
  buf1  g3656(.din(new_new_n7358__), .dout(n13562));
  buf1  g3657(.din(new_new_n7820__), .dout(n13565));
  buf1  g3658(.din(new_new_n7285__), .dout(n13568));
  buf1  g3659(.din(new_new_n7366__), .dout(n13571));
  buf1  g3660(.din(new_new_n7286__), .dout(n13574));
  buf1  g3661(.din(new_new_n7288__), .dout(n13577));
  buf1  g3662(.din(new_new_n7281__), .dout(n13580));
  buf1  g3663(.din(new_new_n7349__), .dout(n13583));
  buf1  g3664(.din(new_new_n7947__), .dout(n13586));
  buf1  g3665(.din(new_new_n7334__), .dout(n13589));
  buf1  g3666(.din(new_new_n7479__), .dout(n13592));
  buf1  g3667(.din(new_new_n7350__), .dout(n13595));
  buf1  g3668(.din(new_new_n7951__), .dout(n13598));
  buf1  g3669(.din(new_new_n7828__), .dout(n13601));
  buf1  g3670(.din(new_new_n7292__), .dout(n13604));
  buf1  g3671(.din(new_new_n7464__), .dout(n13607));
  buf1  g3672(.din(new_new_n7408__), .dout(n13610));
  buf1  g3673(.din(new_new_n7839__), .dout(n13613));
  buf1  g3674(.din(new_new_n7621__), .dout(n13616));
  buf1  g3675(.din(new_new_n7409__), .dout(n13619));
  buf1  g3676(.din(new_new_n4070__), .dout(n13622));
  buf1  g3677(.din(new_new_n4072__), .dout(n13625));
  buf1  g3678(.din(new_new_n4074__), .dout(n13628));
  buf1  g3679(.din(new_new_n7424__), .dout(n13631));
  buf1  g3680(.din(new_new_n7481__), .dout(n13634));
  buf1  g3681(.din(new_new_n7880__), .dout(n13637));
  buf1  g3682(.din(new_new_n7965__), .dout(n13640));
  buf1  g3683(.din(new_new_n7425__), .dout(n13643));
  buf1  g3684(.din(new_new_n7442__), .dout(n13646));
  buf1  g3685(.din(new_new_n7453__), .dout(n13649));
  buf1  g3686(.din(new_new_n7465__), .dout(n13652));
  buf1  g3687(.din(new_new_n7472__), .dout(n13655));
  buf1  g3688(.din(new_new_n7473__), .dout(n13658));
  buf1  g3689(.din(new_new_n7484__), .dout(n13661));
  buf1  g3690(.din(new_new_n7489__), .dout(n13664));
  buf1  g3691(.din(new_new_n7434__), .dout(n13667));
  buf1  g3692(.din(new_new_n7438__), .dout(n13670));
  buf1  g3693(.din(new_new_n7440__), .dout(n13673));
  buf1  g3694(.din(new_new_n7436__), .dout(n13676));
  buf1  g3695(.din(new_new_n7491__), .dout(n13679));
  buf1  g3696(.din(new_new_n7782__), .dout(n13682));
  buf1  g3697(.din(new_new_n7608__), .dout(n13685));
  buf1  g3698(.din(new_new_n4878__), .dout(n13688));
  not1  g3699(.din(new_new_n7615__), .dout(n13691));
  buf1  g3700(.din(new_new_n7571__), .dout(n13694));
  buf1  g3701(.din(new_new_n7572__), .dout(n13697));
  buf1  g3702(.din(new_new_n7570__), .dout(n13700));
  buf1  g3703(.din(new_new_n7794__), .dout(n13703));
  buf1  g3704(.din(new_new_n7496__), .dout(n13706));
  buf1  g3705(.din(new_new_n7497__), .dout(n13709));
  buf1  g3706(.din(new_new_n7485__), .dout(n13712));
  buf1  g3707(.din(new_new_n7510__), .dout(n13715));
  buf1  g3708(.din(new_new_n7487__), .dout(n13718));
  buf1  g3709(.din(new_new_n7717__), .dout(n13721));
  buf1  g3710(.din(new_new_n7495__), .dout(n13724));
  buf1  g3711(.din(new_new_n7893__), .dout(n13727));
  buf1  g3712(.din(new_new_n7512__), .dout(n13730));
  buf1  g3713(.din(new_new_n7852__), .dout(n13733));
  buf1  g3714(.din(new_new_n7890__), .dout(n13736));
  buf1  g3715(.din(new_new_n7945__), .dout(n13739));
  buf1  g3716(.din(new_new_n7784__), .dout(n13742));
  buf1  g3717(.din(new_new_n7785__), .dout(n13745));
  buf1  g3718(.din(new_new_n7786__), .dout(n13748));
  buf1  g3719(.din(new_new_n7498__), .dout(n13751));
  buf1  g3720(.din(new_new_n7502__), .dout(n13754));
  buf1  g3721(.din(new_new_n7506__), .dout(n13757));
  buf1  g3722(.din(new_new_n7504__), .dout(n13760));
  buf1  g3723(.din(new_new_n7500__), .dout(n13763));
  not1  g3724(.din(new_new_n7946__), .dout(n13766));
  buf1  g3725(.din(new_new_n7508__), .dout(n13769));
  buf1  g3726(.din(new_new_n7966__), .dout(n13772));
  buf1  g3727(.din(new_new_n7714__), .dout(n13775));
  buf1  g3728(.din(new_new_n7715__), .dout(n13778));
  buf1  g3729(.din(new_new_n7515__), .dout(n13781));
  buf1  g3730(.din(new_new_n7516__), .dout(n13784));
  buf1  g3731(.din(new_new_n7889__), .dout(n13787));
  buf1  g3732(.din(new_new_n7618__), .dout(n13790));
  buf1  g3733(.din(new_new_n3138__), .dout(n13793));
  buf1  g3734(.din(new_new_n3140__), .dout(n13796));
  buf1  g3735(.din(new_new_n7969__), .dout(n13799));
  buf1  g3736(.din(new_new_n7970__), .dout(n13802));
  buf1  g3737(.din(new_new_n7984__), .dout(n13805));
  buf1  g3738(.din(new_new_n7985__), .dout(n13808));
  buf1  g3739(.din(new_new_n7849__), .dout(n13811));
  buf1  g3740(.din(new_new_n7850__), .dout(n13814));
  buf1  g3741(.din(new_new_n7895__), .dout(n13817));
  buf1  g3742(.din(new_new_n5001__), .dout(n13820));
  buf1  g3743(.din(new_new_n5002__), .dout(n13823));
  buf1  g3744(.din(new_new_n5003__), .dout(n13826));
  buf1  g3745(.din(new_new_n5004__), .dout(n13829));
  buf1  g3746(.din(new_new_n5005__), .dout(n13832));
  buf1  g3747(.din(new_new_n5006__), .dout(n13835));
  buf1  g3748(.din(new_new_n5007__), .dout(n13838));
  buf1  g3749(.din(new_new_n5008__), .dout(n13841));
  buf1  g3750(.din(new_new_n5009__), .dout(n13844));
  buf1  g3751(.din(new_new_n5013__), .dout(n13847));
  buf1  g3752(.din(new_new_n5017__), .dout(n13850));
  buf1  g3753(.din(new_new_n5018__), .dout(n13853));
  buf1  g3754(.din(new_new_n5020__), .dout(n13856));
  buf1  g3755(.din(new_new_n5052__), .dout(n13859));
  not1  g3756(.din(new_new_n5053__), .dout(n13862));
  not1  g3757(.din(new_new_n5054__), .dout(n13865));
  buf1  g3758(.din(new_new_n5055__), .dout(n13868));
  buf1  g3759(.din(new_new_n5056__), .dout(n13871));
  buf1  g3760(.din(new_new_n5057__), .dout(n13874));
  not1  g3761(.din(new_new_n5058__), .dout(n13877));
  buf1  g3762(.din(new_new_n5083__), .dout(n13880));
  buf1  g3763(.din(new_new_n5084__), .dout(n13883));
  buf1  g3764(.din(new_new_n5085__), .dout(n13886));
  buf1  g3765(.din(new_new_n5090__), .dout(n13889));
  buf1  g3766(.din(new_new_n5091__), .dout(n13892));
  not1  g3767(.din(new_new_n5095__), .dout(n13895));
  not1  g3768(.din(new_new_n5096__), .dout(n13898));
  buf1  g3769(.din(new_new_n5097__), .dout(n13901));
  buf1  g3770(.din(new_new_n5098__), .dout(n13904));
  buf1  g3771(.din(new_new_n5102__), .dout(n13907));
  buf1  g3772(.din(new_new_n5103__), .dout(n13910));
  buf1  g3773(.din(new_new_n5104__), .dout(n13913));
  buf1  g3774(.din(new_new_n5105__), .dout(n13916));
  buf1  g3775(.din(new_new_n5106__), .dout(n13919));
  not1  g3776(.din(new_new_n5109__), .dout(n13922));
  not1  g3777(.din(new_new_n5110__), .dout(n13925));
  not1  g3778(.din(new_new_n5111__), .dout(n13928));
  buf1  g3779(.din(new_new_n5115__), .dout(n13931));
  buf1  g3780(.din(new_new_n7994__), .dout(n13934));
  buf1  g3781(.din(new_new_n5120__), .dout(n13937));
  buf1  g3782(.din(new_new_n5123__), .dout(n13940));
  not1  g3783(.din(new_new_n5126__), .dout(n13943));
  buf1  g3784(.din(new_new_n5129__), .dout(n13946));
  buf1  g3785(.din(new_new_n5132__), .dout(n13949));
  buf1  g3786(.din(new_new_n5135__), .dout(n13952));
  buf1  g3787(.din(new_new_n5144__), .dout(n13955));
  buf1  g3788(.din(new_new_n5153__), .dout(n13958));
  buf1  g3789(.din(new_new_n5162__), .dout(n13961));
  buf1  g3790(.din(new_new_n5171__), .dout(n13964));
  buf1  g3791(.din(new_new_n5180__), .dout(n13967));
  buf1  g3792(.din(new_new_n5189__), .dout(n13970));
  buf1  g3793(.din(new_new_n5198__), .dout(n13973));
  buf1  g3794(.din(new_new_n5238__), .dout(n13976));
  buf1  g3795(.din(new_new_n5241__), .dout(n13979));
  buf1  g3796(.din(new_new_n5244__), .dout(n13982));
  buf1  g3797(.din(new_new_n5249__), .dout(n13985));
  buf1  g3798(.din(new_new_n5258__), .dout(n13988));
  buf1  g3799(.din(new_new_n5261__), .dout(n13991));
  buf1  g3800(.din(new_new_n5264__), .dout(n13994));
  buf1  g3801(.din(new_new_n5273__), .dout(n13997));
  buf1  g3802(.din(new_new_n5276__), .dout(n14000));
  buf1  g3803(.din(new_new_n5283__), .dout(n14003));
  not1  g3804(.din(new_new_n5284__), .dout(n14006));
  buf1  g3805(.din(new_new_n5297__), .dout(n14009));
  not1  g3806(.din(new_new_n5298__), .dout(n14012));
  buf1  g3807(.din(new_new_n5305__), .dout(n14015));
  buf1  g3808(.din(new_new_n5306__), .dout(n14018));
  buf1  g3809(.din(new_new_n5321__), .dout(n14021));
  buf1  g3810(.din(new_new_n5372__), .dout(n14024));
  buf1  g3811(.din(new_new_n7848__), .dout(n14027));
  buf1  g3812(.din(new_new_n7982__), .dout(n14030));
  buf1  g3813(.din(new_new_n7896__), .dout(n14033));
  buf1  g3814(.din(new_new_n7899__), .dout(n14036));
  buf1  g3815(.din(new_new_n7903__), .dout(n14039));
  not1  g3816(.din(new_new_n7931__), .dout(n14042));
  not1  g3817(.din(new_new_n7901__), .dout(n14045));
  buf1  g3818(.din(new_new_n7905__), .dout(n14048));
  buf1  g3819(.din(new_new_n7996__), .dout(n14051));
  buf1  g3820(.din(new_new_n7993__), .dout(n14054));
  buf1  g3821(.din(new_new_n7967__), .dout(n14057));
  buf1  g3822(.din(new_new_n7997__), .dout(n14060));
  buf1  g3823(.din(new_new_n7968__), .dout(n14063));
  not1  g3824(.din(new_new_n7971__), .dout(n14066));
  buf1  g3825(.din(new_new_n7983__), .dout(n14069));
  buf1  g3826(.din(new_new_n7978__), .dout(n14072));
  buf1  g3827(.din(new_new_n5426__), .dout(n14075));
  not1  g3828(.din(new_new_n5428__), .dout(n14078));
  not1  g3829(.din(new_new_n5454__), .dout(n14081));
  not1  g3830(.din(new_new_n5455__), .dout(n14084));
  buf1  g3831(.din(new_new_n7979__), .dout(n14087));
  buf1  g3832(.din(new_new_n5479__), .dout(n14090));
  buf1  g3833(.din(new_new_n5480__), .dout(n14093));
  buf1  g3834(.din(new_new_n7981__), .dout(n14096));
  buf1  g3835(.din(new_new_n7986__), .dout(n14099));
  buf1  g3836(.din(new_new_n7972__), .dout(n14102));
  buf1  g3837(.din(new_new_n7973__), .dout(n14105));
  buf1  g3838(.din(new_new_n7987__), .dout(n14108));
  buf1  g3839(.din(new_new_n5486__), .dout(n14111));
  buf1  g3840(.din(new_new_n5495__), .dout(n14114));
  buf1  g3841(.din(new_new_n5504__), .dout(n14117));
  buf1  g3842(.din(new_new_n5513__), .dout(n14120));
  buf1  g3843(.din(new_new_n5522__), .dout(n14123));
  buf1  g3844(.din(new_new_n5531__), .dout(n14126));
  buf1  g3845(.din(new_new_n5540__), .dout(n14129));
  buf1  g3846(.din(new_new_n5549__), .dout(n14132));
  buf1  g3847(.din(new_new_n5558__), .dout(n14135));
  not1  g3848(.din(new_new_n5575__), .dout(n14138));
  not1  g3849(.din(new_new_n5576__), .dout(n14141));
  buf1  g3850(.din(new_new_n7989__), .dout(n14144));
  not1  g3851(.din(new_new_n7991__), .dout(n14147));
  not1  g3852(.din(new_new_n7995__), .dout(n14150));
  buf1  g3853(.din(new_new_n5588__), .dout(n14153));
  buf1  g3854(.din(new_new_n5589__), .dout(n14156));
  buf1  g3855(.din(new_new_n7974__), .dout(n14159));
  buf1  g3856(.din(new_new_n5592__), .dout(n14162));
  not1  g3857(.din(new_new_n5593__), .dout(n14165));
  buf1  g3858(.din(new_new_n5594__), .dout(n14168));
  buf1  g3859(.din(new_new_n5595__), .dout(n14171));
  not1  g3860(.din(new_new_n5623__), .dout(n14174));
  buf1  g3861(.din(new_new_n5624__), .dout(n14177));
  not1  g3862(.din(new_new_n5643__), .dout(n14180));
  buf1  g3863(.din(new_new_n5644__), .dout(n14183));
  not1  g3864(.din(new_new_n5652__), .dout(n14186));
  buf1  g3865(.din(new_new_n5665__), .dout(n14189));
  buf1  g3866(.din(new_new_n5704__), .dout(n14192));
  buf1  g3867(.din(new_new_n5713__), .dout(n14195));
  not1  g3868(.din(new_new_n7998__), .dout(n14198));
  not1  g3869(.din(new_new_n7999__), .dout(n14201));
  buf1  g3870(.din(new_new_n8000__), .dout(n14204));
  buf1  g3871(.din(new_new_n7992__), .dout(n14207));
  buf1  g3872(.din(new_new_n3186__), .dout(n14210));
  buf1  g3873(.din(new_new_n5719__), .dout(n14213));
  buf1  g3874(.din(new_new_n5720__), .dout(n14216));
  buf1  g3875(.din(new_new_n5721__), .dout(n14219));
  buf1  g3876(.din(new_new_n5722__), .dout(n14222));
  buf1  g3877(.din(new_new_n5723__), .dout(n14225));
  buf1  g3878(.din(new_new_n5724__), .dout(n14228));
  buf1  g3879(.din(new_new_n5725__), .dout(n14231));
  buf1  g3880(.din(new_new_n5726__), .dout(n14234));
  buf1  g3881(.din(new_new_n5727__), .dout(n14237));
  buf1  g3882(.din(new_new_n5729__), .dout(n14240));
  buf1  g3883(.din(new_new_n5731__), .dout(n14243));
  buf1  g3884(.din(new_new_n5732__), .dout(n14246));
  buf1  g3885(.din(new_new_n3070__), .dout(n14249));
  buf1  g3886(.din(new_new_n3072__), .dout(n14252));
  buf1  g3887(.din(new_new_n3074__), .dout(n14255));
  buf1  g3888(.din(new_new_n3084__), .dout(n14258));
  buf1  g3889(.din(new_new_n3086__), .dout(n14261));
  buf1  g3890(.din(new_new_n3088__), .dout(n14264));
  buf1  g3891(.din(new_new_n5733__), .dout(n14267));
  buf1  g3892(.din(new_new_n8001__), .dout(n14270));
  buf1  g3893(.din(new_new_n8007__), .dout(n14273));
  buf1  g3894(.din(new_new_n8008__), .dout(n14276));
  buf1  g3895(.din(new_new_n8004__), .dout(n14279));
  buf1  g3896(.din(new_new_n5734__), .dout(n14282));
  buf1  g3897(.din(new_new_n5735__), .dout(n14285));
  buf1  g3898(.din(new_new_n5736__), .dout(n14288));
  buf1  g3899(.din(new_new_n5738__), .dout(n14291));
  buf1  g3900(.din(new_new_n5740__), .dout(n14294));
  buf1  g3901(.din(new_new_n5741__), .dout(n14297));
  buf1  g3902(.din(new_new_n2296__), .dout(n14300));
  buf1  g3903(.din(new_new_n2298__), .dout(n14303));
  buf1  g3904(.din(new_new_n2310__), .dout(n14306));
  buf1  g3905(.din(new_new_n2330__), .dout(n14309));
  buf1  g3906(.din(new_new_n2220__), .dout(n14312));
  buf1  g3907(.din(new_new_n2222__), .dout(n14315));
  buf1  g3908(.din(new_new_n2250__), .dout(n14318));
  buf1  g3909(.din(new_new_n2252__), .dout(n14321));
  buf1  g3910(.din(new_new_n2278__), .dout(n14324));
  buf1  g3911(.din(new_new_n2280__), .dout(n14327));
  buf1  g3912(.din(new_new_n2318__), .dout(n14330));
  buf1  g3913(.din(new_new_n2320__), .dout(n14333));
  buf1  g3914(.din(new_new_n2328__), .dout(n14336));
  buf1  g3915(.din(new_new_n2258__), .dout(n14339));
  buf1  g3916(.din(new_new_n2260__), .dout(n14342));
  buf1  g3917(.din(new_new_n2274__), .dout(n14345));
  buf1  g3918(.din(new_new_n2276__), .dout(n14348));
  buf1  g3919(.din(new_new_n2286__), .dout(n14351));
  buf1  g3920(.din(new_new_n5742__), .dout(n14354));
  buf1  g3921(.din(new_new_n5743__), .dout(n14357));
  buf1  g3922(.din(new_new_n5744__), .dout(n14360));
  buf1  g3923(.din(new_new_n5745__), .dout(n14363));
  buf1  g3924(.din(new_new_n5746__), .dout(n14366));
  buf1  g3925(.din(new_new_n5747__), .dout(n14369));
  buf1  g3926(.din(new_new_n3217__), .dout(new_new_n6741__));
  buf1  g3927(.din(new_new_n3241__), .dout(new_new_n6742__));
  buf1  g3928(.din(new_new_n2896__), .dout(new_new_n6743__));
  buf1  g3929(.din(new_new_n6743__), .dout(new_new_n6744__));
  buf1  g3930(.din(new_new_n6744__), .dout(new_new_n6745__));
  buf1  g3931(.din(new_new_n6744__), .dout(new_new_n6746__));
  buf1  g3932(.din(new_new_n6743__), .dout(new_new_n6747__));
  buf1  g3933(.din(new_new_n2404__), .dout(new_new_n6748__));
  buf1  g3934(.din(new_new_n3307__), .dout(new_new_n6749__));
  buf1  g3935(.din(new_new_n2483__), .dout(new_new_n6750__));
  buf1  g3936(.din(new_new_n4144__), .dout(new_new_n6751__));
  buf1  g3937(.din(new_new_n6751__), .dout(new_new_n6752__));
  buf1  g3938(.din(new_new_n6752__), .dout(new_new_n6753__));
  buf1  g3939(.din(new_new_n6753__), .dout(new_new_n6754__));
  buf1  g3940(.din(new_new_n6752__), .dout(new_new_n6755__));
  buf1  g3941(.din(new_new_n6751__), .dout(new_new_n6756__));
  buf1  g3942(.din(new_new_n6756__), .dout(new_new_n6757__));
  buf1  g3943(.din(new_new_n6756__), .dout(new_new_n6758__));
  buf1  g3944(.din(new_new_n3291__), .dout(new_new_n6759__));
  buf1  g3945(.din(new_new_n6759__), .dout(new_new_n6760__));
  buf1  g3946(.din(new_new_n6760__), .dout(new_new_n6761__));
  buf1  g3947(.din(new_new_n6760__), .dout(new_new_n6762__));
  buf1  g3948(.din(new_new_n6759__), .dout(new_new_n6763__));
  buf1  g3949(.din(new_new_n3290__), .dout(new_new_n6764__));
  buf1  g3950(.din(new_new_n6764__), .dout(new_new_n6765__));
  buf1  g3951(.din(new_new_n6765__), .dout(new_new_n6766__));
  buf1  g3952(.din(new_new_n6765__), .dout(new_new_n6767__));
  buf1  g3953(.din(new_new_n6764__), .dout(new_new_n6768__));
  buf1  g3954(.din(new_new_n3872__), .dout(new_new_n6769__));
  buf1  g3955(.din(new_new_n4183__), .dout(new_new_n6770__));
  buf1  g3956(.din(new_new_n3437__), .dout(new_new_n6771__));
  buf1  g3957(.din(new_new_n4190__), .dout(new_new_n6772__));
  buf1  g3958(.din(new_new_n3854__), .dout(new_new_n6773__));
  buf1  g3959(.din(new_new_n3856__), .dout(new_new_n6774__));
  buf1  g3960(.din(new_new_n3855__), .dout(new_new_n6775__));
  buf1  g3961(.din(new_new_n3857__), .dout(new_new_n6776__));
  buf1  g3962(.din(new_new_n3859__), .dout(new_new_n6777__));
  buf1  g3963(.din(new_new_n3905__), .dout(new_new_n6778__));
  buf1  g3964(.din(new_new_n3858__), .dout(new_new_n6779__));
  buf1  g3965(.din(new_new_n3904__), .dout(new_new_n6780__));
  buf1  g3966(.din(new_new_n3462__), .dout(new_new_n6781__));
  buf1  g3967(.din(new_new_n6781__), .dout(new_new_n6782__));
  buf1  g3968(.din(new_new_n3792__), .dout(new_new_n6783__));
  buf1  g3969(.din(new_new_n6783__), .dout(new_new_n6784__));
  buf1  g3970(.din(new_new_n6784__), .dout(new_new_n6785__));
  buf1  g3971(.din(new_new_n6785__), .dout(new_new_n6786__));
  buf1  g3972(.din(new_new_n6785__), .dout(new_new_n6787__));
  buf1  g3973(.din(new_new_n6784__), .dout(new_new_n6788__));
  buf1  g3974(.din(new_new_n6788__), .dout(new_new_n6789__));
  buf1  g3975(.din(new_new_n6788__), .dout(new_new_n6790__));
  buf1  g3976(.din(new_new_n6783__), .dout(new_new_n6791__));
  buf1  g3977(.din(new_new_n6791__), .dout(new_new_n6792__));
  buf1  g3978(.din(new_new_n6792__), .dout(new_new_n6793__));
  buf1  g3979(.din(new_new_n6792__), .dout(new_new_n6794__));
  buf1  g3980(.din(new_new_n6791__), .dout(new_new_n6795__));
  buf1  g3981(.din(new_new_n6795__), .dout(new_new_n6796__));
  buf1  g3982(.din(new_new_n6795__), .dout(new_new_n6797__));
  buf1  g3983(.din(new_new_n3395__), .dout(new_new_n6798__));
  buf1  g3984(.din(new_new_n6798__), .dout(new_new_n6799__));
  buf1  g3985(.din(new_new_n6799__), .dout(new_new_n6800__));
  buf1  g3986(.din(new_new_n6800__), .dout(new_new_n6801__));
  buf1  g3987(.din(new_new_n6799__), .dout(new_new_n6802__));
  buf1  g3988(.din(new_new_n6798__), .dout(new_new_n6803__));
  buf1  g3989(.din(new_new_n6803__), .dout(new_new_n6804__));
  buf1  g3990(.din(new_new_n6803__), .dout(new_new_n6805__));
  buf1  g3991(.din(new_new_n3386__), .dout(new_new_n6806__));
  buf1  g3992(.din(new_new_n6806__), .dout(new_new_n6807__));
  buf1  g3993(.din(new_new_n6807__), .dout(new_new_n6808__));
  buf1  g3994(.din(new_new_n6808__), .dout(new_new_n6809__));
  buf1  g3995(.din(new_new_n6808__), .dout(new_new_n6810__));
  buf1  g3996(.din(new_new_n6807__), .dout(new_new_n6811__));
  buf1  g3997(.din(new_new_n6811__), .dout(new_new_n6812__));
  buf1  g3998(.din(new_new_n6811__), .dout(new_new_n6813__));
  buf1  g3999(.din(new_new_n6806__), .dout(new_new_n6814__));
  buf1  g4000(.din(new_new_n6814__), .dout(new_new_n6815__));
  buf1  g4001(.din(new_new_n6815__), .dout(new_new_n6816__));
  buf1  g4002(.din(new_new_n6815__), .dout(new_new_n6817__));
  buf1  g4003(.din(new_new_n6814__), .dout(new_new_n6818__));
  buf1  g4004(.din(new_new_n6818__), .dout(new_new_n6819__));
  buf1  g4005(.din(new_new_n3793__), .dout(new_new_n6820__));
  buf1  g4006(.din(new_new_n3394__), .dout(new_new_n6821__));
  buf1  g4007(.din(new_new_n6821__), .dout(new_new_n6822__));
  buf1  g4008(.din(new_new_n6822__), .dout(new_new_n6823__));
  buf1  g4009(.din(new_new_n6823__), .dout(new_new_n6824__));
  buf1  g4010(.din(new_new_n6822__), .dout(new_new_n6825__));
  buf1  g4011(.din(new_new_n6821__), .dout(new_new_n6826__));
  buf1  g4012(.din(new_new_n6826__), .dout(new_new_n6827__));
  buf1  g4013(.din(new_new_n6826__), .dout(new_new_n6828__));
  buf1  g4014(.din(new_new_n3387__), .dout(new_new_n6829__));
  buf1  g4015(.din(new_new_n6829__), .dout(new_new_n6830__));
  buf1  g4016(.din(new_new_n6829__), .dout(new_new_n6831__));
  buf1  g4017(.din(new_new_n3844__), .dout(new_new_n6832__));
  buf1  g4018(.din(new_new_n3363__), .dout(new_new_n6833__));
  buf1  g4019(.din(new_new_n6833__), .dout(new_new_n6834__));
  buf1  g4020(.din(new_new_n6834__), .dout(new_new_n6835__));
  buf1  g4021(.din(new_new_n6835__), .dout(new_new_n6836__));
  buf1  g4022(.din(new_new_n6836__), .dout(new_new_n6837__));
  buf1  g4023(.din(new_new_n6836__), .dout(new_new_n6838__));
  buf1  g4024(.din(new_new_n6835__), .dout(new_new_n6839__));
  buf1  g4025(.din(new_new_n6839__), .dout(new_new_n6840__));
  buf1  g4026(.din(new_new_n6839__), .dout(new_new_n6841__));
  buf1  g4027(.din(new_new_n6834__), .dout(new_new_n6842__));
  buf1  g4028(.din(new_new_n6842__), .dout(new_new_n6843__));
  buf1  g4029(.din(new_new_n6842__), .dout(new_new_n6844__));
  buf1  g4030(.din(new_new_n6833__), .dout(new_new_n6845__));
  buf1  g4031(.din(new_new_n6845__), .dout(new_new_n6846__));
  buf1  g4032(.din(new_new_n6846__), .dout(new_new_n6847__));
  buf1  g4033(.din(new_new_n6846__), .dout(new_new_n6848__));
  buf1  g4034(.din(new_new_n6845__), .dout(new_new_n6849__));
  buf1  g4035(.din(new_new_n6849__), .dout(new_new_n6850__));
  buf1  g4036(.din(new_new_n6849__), .dout(new_new_n6851__));
  buf1  g4037(.din(new_new_n4229__), .dout(new_new_n6852__));
  buf1  g4038(.din(new_new_n6852__), .dout(new_new_n6853__));
  buf1  g4039(.din(new_new_n6853__), .dout(new_new_n6854__));
  buf1  g4040(.din(new_new_n6852__), .dout(new_new_n6855__));
  buf1  g4041(.din(new_new_n3362__), .dout(new_new_n6856__));
  buf1  g4042(.din(new_new_n6856__), .dout(new_new_n6857__));
  buf1  g4043(.din(new_new_n6857__), .dout(new_new_n6858__));
  buf1  g4044(.din(new_new_n6858__), .dout(new_new_n6859__));
  buf1  g4045(.din(new_new_n6859__), .dout(new_new_n6860__));
  buf1  g4046(.din(new_new_n6859__), .dout(new_new_n6861__));
  buf1  g4047(.din(new_new_n6858__), .dout(new_new_n6862__));
  buf1  g4048(.din(new_new_n6862__), .dout(new_new_n6863__));
  buf1  g4049(.din(new_new_n6862__), .dout(new_new_n6864__));
  buf1  g4050(.din(new_new_n6857__), .dout(new_new_n6865__));
  buf1  g4051(.din(new_new_n6865__), .dout(new_new_n6866__));
  buf1  g4052(.din(new_new_n6865__), .dout(new_new_n6867__));
  buf1  g4053(.din(new_new_n6856__), .dout(new_new_n6868__));
  buf1  g4054(.din(new_new_n6868__), .dout(new_new_n6869__));
  buf1  g4055(.din(new_new_n6869__), .dout(new_new_n6870__));
  buf1  g4056(.din(new_new_n6869__), .dout(new_new_n6871__));
  buf1  g4057(.din(new_new_n6868__), .dout(new_new_n6872__));
  buf1  g4058(.din(new_new_n6872__), .dout(new_new_n6873__));
  buf1  g4059(.din(new_new_n6872__), .dout(new_new_n6874__));
  buf1  g4060(.din(new_new_n4239__), .dout(new_new_n6875__));
  buf1  g4061(.din(new_new_n6875__), .dout(new_new_n6876__));
  buf1  g4062(.din(new_new_n6876__), .dout(new_new_n6877__));
  buf1  g4063(.din(new_new_n6875__), .dout(new_new_n6878__));
  buf1  g4064(.din(new_new_n3354__), .dout(new_new_n6879__));
  buf1  g4065(.din(new_new_n6879__), .dout(new_new_n6880__));
  buf1  g4066(.din(new_new_n6880__), .dout(new_new_n6881__));
  buf1  g4067(.din(new_new_n6881__), .dout(new_new_n6882__));
  buf1  g4068(.din(new_new_n6881__), .dout(new_new_n6883__));
  buf1  g4069(.din(new_new_n6880__), .dout(new_new_n6884__));
  buf1  g4070(.din(new_new_n6879__), .dout(new_new_n6885__));
  buf1  g4071(.din(new_new_n6885__), .dout(new_new_n6886__));
  buf1  g4072(.din(new_new_n6885__), .dout(new_new_n6887__));
  buf1  g4073(.din(new_new_n2418__), .dout(new_new_n6888__));
  buf1  g4074(.din(new_new_n2566__), .dout(new_new_n6889__));
  buf1  g4075(.din(new_new_n3355__), .dout(new_new_n6890__));
  buf1  g4076(.din(new_new_n6890__), .dout(new_new_n6891__));
  buf1  g4077(.din(new_new_n6891__), .dout(new_new_n6892__));
  buf1  g4078(.din(new_new_n6892__), .dout(new_new_n6893__));
  buf1  g4079(.din(new_new_n6892__), .dout(new_new_n6894__));
  buf1  g4080(.din(new_new_n6891__), .dout(new_new_n6895__));
  buf1  g4081(.din(new_new_n6890__), .dout(new_new_n6896__));
  buf1  g4082(.din(new_new_n6896__), .dout(new_new_n6897__));
  buf1  g4083(.din(new_new_n6896__), .dout(new_new_n6898__));
  buf1  g4084(.din(new_new_n3445__), .dout(new_new_n6899__));
  buf1  g4085(.din(new_new_n3887__), .dout(new_new_n6900__));
  buf1  g4086(.din(new_new_n4256__), .dout(new_new_n6901__));
  buf1  g4087(.din(new_new_n3371__), .dout(new_new_n6902__));
  buf1  g4088(.din(new_new_n6902__), .dout(new_new_n6903__));
  buf1  g4089(.din(new_new_n6903__), .dout(new_new_n6904__));
  buf1  g4090(.din(new_new_n6904__), .dout(new_new_n6905__));
  buf1  g4091(.din(new_new_n6905__), .dout(new_new_n6906__));
  buf1  g4092(.din(new_new_n6905__), .dout(new_new_n6907__));
  buf1  g4093(.din(new_new_n6904__), .dout(new_new_n6908__));
  buf1  g4094(.din(new_new_n6908__), .dout(new_new_n6909__));
  buf1  g4095(.din(new_new_n6908__), .dout(new_new_n6910__));
  buf1  g4096(.din(new_new_n6903__), .dout(new_new_n6911__));
  buf1  g4097(.din(new_new_n6911__), .dout(new_new_n6912__));
  buf1  g4098(.din(new_new_n6911__), .dout(new_new_n6913__));
  buf1  g4099(.din(new_new_n6902__), .dout(new_new_n6914__));
  buf1  g4100(.din(new_new_n6914__), .dout(new_new_n6915__));
  buf1  g4101(.din(new_new_n6915__), .dout(new_new_n6916__));
  buf1  g4102(.din(new_new_n6915__), .dout(new_new_n6917__));
  buf1  g4103(.din(new_new_n6914__), .dout(new_new_n6918__));
  buf1  g4104(.din(new_new_n6918__), .dout(new_new_n6919__));
  buf1  g4105(.din(new_new_n6918__), .dout(new_new_n6920__));
  buf1  g4106(.din(new_new_n3370__), .dout(new_new_n6921__));
  buf1  g4107(.din(new_new_n6921__), .dout(new_new_n6922__));
  buf1  g4108(.din(new_new_n6922__), .dout(new_new_n6923__));
  buf1  g4109(.din(new_new_n6923__), .dout(new_new_n6924__));
  buf1  g4110(.din(new_new_n6924__), .dout(new_new_n6925__));
  buf1  g4111(.din(new_new_n6924__), .dout(new_new_n6926__));
  buf1  g4112(.din(new_new_n6923__), .dout(new_new_n6927__));
  buf1  g4113(.din(new_new_n6927__), .dout(new_new_n6928__));
  buf1  g4114(.din(new_new_n6927__), .dout(new_new_n6929__));
  buf1  g4115(.din(new_new_n6922__), .dout(new_new_n6930__));
  buf1  g4116(.din(new_new_n6930__), .dout(new_new_n6931__));
  buf1  g4117(.din(new_new_n6930__), .dout(new_new_n6932__));
  buf1  g4118(.din(new_new_n6921__), .dout(new_new_n6933__));
  buf1  g4119(.din(new_new_n6933__), .dout(new_new_n6934__));
  buf1  g4120(.din(new_new_n6934__), .dout(new_new_n6935__));
  buf1  g4121(.din(new_new_n6934__), .dout(new_new_n6936__));
  buf1  g4122(.din(new_new_n6933__), .dout(new_new_n6937__));
  buf1  g4123(.din(new_new_n6937__), .dout(new_new_n6938__));
  buf1  g4124(.din(new_new_n6937__), .dout(new_new_n6939__));
  buf1  g4125(.din(new_new_n3378__), .dout(new_new_n6940__));
  buf1  g4126(.din(new_new_n6940__), .dout(new_new_n6941__));
  buf1  g4127(.din(new_new_n6941__), .dout(new_new_n6942__));
  buf1  g4128(.din(new_new_n6942__), .dout(new_new_n6943__));
  buf1  g4129(.din(new_new_n6942__), .dout(new_new_n6944__));
  buf1  g4130(.din(new_new_n6941__), .dout(new_new_n6945__));
  buf1  g4131(.din(new_new_n6940__), .dout(new_new_n6946__));
  buf1  g4132(.din(new_new_n6946__), .dout(new_new_n6947__));
  buf1  g4133(.din(new_new_n6946__), .dout(new_new_n6948__));
  buf1  g4134(.din(new_new_n3379__), .dout(new_new_n6949__));
  buf1  g4135(.din(new_new_n6949__), .dout(new_new_n6950__));
  buf1  g4136(.din(new_new_n6950__), .dout(new_new_n6951__));
  buf1  g4137(.din(new_new_n6951__), .dout(new_new_n6952__));
  buf1  g4138(.din(new_new_n6951__), .dout(new_new_n6953__));
  buf1  g4139(.din(new_new_n6950__), .dout(new_new_n6954__));
  buf1  g4140(.din(new_new_n6949__), .dout(new_new_n6955__));
  buf1  g4141(.din(new_new_n6955__), .dout(new_new_n6956__));
  buf1  g4142(.din(new_new_n6955__), .dout(new_new_n6957__));
  buf1  g4143(.din(new_new_n4273__), .dout(new_new_n6958__));
  buf1  g4144(.din(new_new_n4280__), .dout(new_new_n6959__));
  buf1  g4145(.din(new_new_n4285__), .dout(new_new_n6960__));
  buf1  g4146(.din(new_new_n3521__), .dout(new_new_n6961__));
  buf1  g4147(.din(new_new_n6961__), .dout(new_new_n6962__));
  buf1  g4148(.din(new_new_n6962__), .dout(new_new_n6963__));
  buf1  g4149(.din(new_new_n6961__), .dout(new_new_n6964__));
  buf1  g4150(.din(new_new_n4299__), .dout(new_new_n6965__));
  buf1  g4151(.din(new_new_n3520__), .dout(new_new_n6966__));
  buf1  g4152(.din(new_new_n6966__), .dout(new_new_n6967__));
  buf1  g4153(.din(new_new_n6966__), .dout(new_new_n6968__));
  buf1  g4154(.din(new_new_n4298__), .dout(new_new_n6969__));
  buf1  g4155(.din(new_new_n4306__), .dout(new_new_n6970__));
  buf1  g4156(.din(new_new_n4309__), .dout(new_new_n6971__));
  buf1  g4157(.din(new_new_n4307__), .dout(new_new_n6972__));
  buf1  g4158(.din(new_new_n4308__), .dout(new_new_n6973__));
  buf1  g4159(.din(new_new_n3407__), .dout(new_new_n6974__));
  buf1  g4160(.din(new_new_n3408__), .dout(new_new_n6975__));
  buf1  g4161(.din(new_new_n3406__), .dout(new_new_n6976__));
  buf1  g4162(.din(new_new_n3409__), .dout(new_new_n6977__));
  buf1  g4163(.din(new_new_n3413__), .dout(new_new_n6978__));
  buf1  g4164(.din(new_new_n3420__), .dout(new_new_n6979__));
  buf1  g4165(.din(new_new_n3412__), .dout(new_new_n6980__));
  buf1  g4166(.din(new_new_n3421__), .dout(new_new_n6981__));
  buf1  g4167(.din(new_new_n4324__), .dout(new_new_n6982__));
  buf1  g4168(.din(new_new_n4329__), .dout(new_new_n6983__));
  buf1  g4169(.din(new_new_n4323__), .dout(new_new_n6984__));
  buf1  g4170(.din(new_new_n4330__), .dout(new_new_n6985__));
  buf1  g4171(.din(new_new_n3877__), .dout(new_new_n6986__));
  buf1  g4172(.din(new_new_n3882__), .dout(new_new_n6987__));
  buf1  g4173(.din(new_new_n3876__), .dout(new_new_n6988__));
  buf1  g4174(.din(new_new_n3883__), .dout(new_new_n6989__));
  buf1  g4175(.din(new_new_n3404__), .dout(new_new_n6990__));
  buf1  g4176(.din(new_new_n3411__), .dout(new_new_n6991__));
  buf1  g4177(.din(new_new_n3405__), .dout(new_new_n6992__));
  buf1  g4178(.din(new_new_n3410__), .dout(new_new_n6993__));
  buf1  g4179(.din(new_new_n4342__), .dout(new_new_n6994__));
  buf1  g4180(.din(new_new_n4347__), .dout(new_new_n6995__));
  buf1  g4181(.din(new_new_n4341__), .dout(new_new_n6996__));
  buf1  g4182(.din(new_new_n4348__), .dout(new_new_n6997__));
  buf1  g4183(.din(new_new_n4358__), .dout(new_new_n6998__));
  buf1  g4184(.din(new_new_n3889__), .dout(new_new_n6999__));
  buf1  g4185(.din(new_new_n4367__), .dout(new_new_n7000__));
  buf1  g4186(.din(new_new_n4370__), .dout(new_new_n7001__));
  buf1  g4187(.din(new_new_n3890__), .dout(new_new_n7002__));
  buf1  g4188(.din(new_new_n4374__), .dout(new_new_n7003__));
  buf1  g4189(.din(new_new_n4373__), .dout(new_new_n7004__));
  buf1  g4190(.din(new_new_n3255__), .dout(new_new_n7005__));
  buf1  g4191(.din(new_new_n7005__), .dout(new_new_n7006__));
  buf1  g4192(.din(new_new_n7006__), .dout(new_new_n7007__));
  buf1  g4193(.din(new_new_n7007__), .dout(new_new_n7008__));
  buf1  g4194(.din(new_new_n7008__), .dout(new_new_n7009__));
  buf1  g4195(.din(new_new_n7008__), .dout(new_new_n7010__));
  buf1  g4196(.din(new_new_n7007__), .dout(new_new_n7011__));
  buf1  g4197(.din(new_new_n7011__), .dout(new_new_n7012__));
  buf1  g4198(.din(new_new_n7011__), .dout(new_new_n7013__));
  buf1  g4199(.din(new_new_n7006__), .dout(new_new_n7014__));
  buf1  g4200(.din(new_new_n7014__), .dout(new_new_n7015__));
  buf1  g4201(.din(new_new_n7014__), .dout(new_new_n7016__));
  buf1  g4202(.din(new_new_n7005__), .dout(new_new_n7017__));
  buf1  g4203(.din(new_new_n7017__), .dout(new_new_n7018__));
  buf1  g4204(.din(new_new_n7018__), .dout(new_new_n7019__));
  buf1  g4205(.din(new_new_n7018__), .dout(new_new_n7020__));
  buf1  g4206(.din(new_new_n7017__), .dout(new_new_n7021__));
  buf1  g4207(.din(new_new_n7021__), .dout(new_new_n7022__));
  buf1  g4208(.din(new_new_n7021__), .dout(new_new_n7023__));
  buf1  g4209(.din(new_new_n3254__), .dout(new_new_n7024__));
  buf1  g4210(.din(new_new_n7024__), .dout(new_new_n7025__));
  buf1  g4211(.din(new_new_n7025__), .dout(new_new_n7026__));
  buf1  g4212(.din(new_new_n7026__), .dout(new_new_n7027__));
  buf1  g4213(.din(new_new_n7027__), .dout(new_new_n7028__));
  buf1  g4214(.din(new_new_n7027__), .dout(new_new_n7029__));
  buf1  g4215(.din(new_new_n7026__), .dout(new_new_n7030__));
  buf1  g4216(.din(new_new_n7030__), .dout(new_new_n7031__));
  buf1  g4217(.din(new_new_n7030__), .dout(new_new_n7032__));
  buf1  g4218(.din(new_new_n7025__), .dout(new_new_n7033__));
  buf1  g4219(.din(new_new_n7033__), .dout(new_new_n7034__));
  buf1  g4220(.din(new_new_n7033__), .dout(new_new_n7035__));
  buf1  g4221(.din(new_new_n7024__), .dout(new_new_n7036__));
  buf1  g4222(.din(new_new_n7036__), .dout(new_new_n7037__));
  buf1  g4223(.din(new_new_n7037__), .dout(new_new_n7038__));
  buf1  g4224(.din(new_new_n7037__), .dout(new_new_n7039__));
  buf1  g4225(.din(new_new_n7036__), .dout(new_new_n7040__));
  buf1  g4226(.din(new_new_n7040__), .dout(new_new_n7041__));
  buf1  g4227(.din(new_new_n7040__), .dout(new_new_n7042__));
  buf1  g4228(.din(new_new_n3263__), .dout(new_new_n7043__));
  buf1  g4229(.din(new_new_n7043__), .dout(new_new_n7044__));
  buf1  g4230(.din(new_new_n7044__), .dout(new_new_n7045__));
  buf1  g4231(.din(new_new_n7045__), .dout(new_new_n7046__));
  buf1  g4232(.din(new_new_n7045__), .dout(new_new_n7047__));
  buf1  g4233(.din(new_new_n7044__), .dout(new_new_n7048__));
  buf1  g4234(.din(new_new_n7043__), .dout(new_new_n7049__));
  buf1  g4235(.din(new_new_n7049__), .dout(new_new_n7050__));
  buf1  g4236(.din(new_new_n7049__), .dout(new_new_n7051__));
  buf1  g4237(.din(new_new_n3016__), .dout(new_new_n7052__));
  buf1  g4238(.din(new_new_n3008__), .dout(new_new_n7053__));
  buf1  g4239(.din(new_new_n3262__), .dout(new_new_n7054__));
  buf1  g4240(.din(new_new_n7054__), .dout(new_new_n7055__));
  buf1  g4241(.din(new_new_n7055__), .dout(new_new_n7056__));
  buf1  g4242(.din(new_new_n7056__), .dout(new_new_n7057__));
  buf1  g4243(.din(new_new_n7056__), .dout(new_new_n7058__));
  buf1  g4244(.din(new_new_n7055__), .dout(new_new_n7059__));
  buf1  g4245(.din(new_new_n7054__), .dout(new_new_n7060__));
  buf1  g4246(.din(new_new_n7060__), .dout(new_new_n7061__));
  buf1  g4247(.din(new_new_n7060__), .dout(new_new_n7062__));
  buf1  g4248(.din(new_new_n2880__), .dout(new_new_n7063__));
  buf1  g4249(.din(new_new_n7063__), .dout(new_new_n7064__));
  buf1  g4250(.din(new_new_n7064__), .dout(new_new_n7065__));
  buf1  g4251(.din(new_new_n7065__), .dout(new_new_n7066__));
  buf1  g4252(.din(new_new_n7066__), .dout(new_new_n7067__));
  buf1  g4253(.din(new_new_n7065__), .dout(new_new_n7068__));
  buf1  g4254(.din(new_new_n7064__), .dout(new_new_n7069__));
  buf1  g4255(.din(new_new_n7069__), .dout(new_new_n7070__));
  buf1  g4256(.din(new_new_n7069__), .dout(new_new_n7071__));
  buf1  g4257(.din(new_new_n7063__), .dout(new_new_n7072__));
  buf1  g4258(.din(new_new_n7072__), .dout(new_new_n7073__));
  buf1  g4259(.din(new_new_n7073__), .dout(new_new_n7074__));
  buf1  g4260(.din(new_new_n7073__), .dout(new_new_n7075__));
  buf1  g4261(.din(new_new_n7072__), .dout(new_new_n7076__));
  buf1  g4262(.din(new_new_n7076__), .dout(new_new_n7077__));
  buf1  g4263(.din(new_new_n7076__), .dout(new_new_n7078__));
  buf1  g4264(.din(new_new_n3271__), .dout(new_new_n7079__));
  buf1  g4265(.din(new_new_n7079__), .dout(new_new_n7080__));
  buf1  g4266(.din(new_new_n7080__), .dout(new_new_n7081__));
  buf1  g4267(.din(new_new_n7081__), .dout(new_new_n7082__));
  buf1  g4268(.din(new_new_n7082__), .dout(new_new_n7083__));
  buf1  g4269(.din(new_new_n7082__), .dout(new_new_n7084__));
  buf1  g4270(.din(new_new_n7081__), .dout(new_new_n7085__));
  buf1  g4271(.din(new_new_n7085__), .dout(new_new_n7086__));
  buf1  g4272(.din(new_new_n7085__), .dout(new_new_n7087__));
  buf1  g4273(.din(new_new_n7080__), .dout(new_new_n7088__));
  buf1  g4274(.din(new_new_n7088__), .dout(new_new_n7089__));
  buf1  g4275(.din(new_new_n7088__), .dout(new_new_n7090__));
  buf1  g4276(.din(new_new_n7079__), .dout(new_new_n7091__));
  buf1  g4277(.din(new_new_n7091__), .dout(new_new_n7092__));
  buf1  g4278(.din(new_new_n7092__), .dout(new_new_n7093__));
  buf1  g4279(.din(new_new_n7092__), .dout(new_new_n7094__));
  buf1  g4280(.din(new_new_n7091__), .dout(new_new_n7095__));
  buf1  g4281(.din(new_new_n7095__), .dout(new_new_n7096__));
  buf1  g4282(.din(new_new_n7095__), .dout(new_new_n7097__));
  buf1  g4283(.din(new_new_n3270__), .dout(new_new_n7098__));
  buf1  g4284(.din(new_new_n7098__), .dout(new_new_n7099__));
  buf1  g4285(.din(new_new_n7099__), .dout(new_new_n7100__));
  buf1  g4286(.din(new_new_n7100__), .dout(new_new_n7101__));
  buf1  g4287(.din(new_new_n7101__), .dout(new_new_n7102__));
  buf1  g4288(.din(new_new_n7101__), .dout(new_new_n7103__));
  buf1  g4289(.din(new_new_n7100__), .dout(new_new_n7104__));
  buf1  g4290(.din(new_new_n7104__), .dout(new_new_n7105__));
  buf1  g4291(.din(new_new_n7104__), .dout(new_new_n7106__));
  buf1  g4292(.din(new_new_n7099__), .dout(new_new_n7107__));
  buf1  g4293(.din(new_new_n7107__), .dout(new_new_n7108__));
  buf1  g4294(.din(new_new_n7107__), .dout(new_new_n7109__));
  buf1  g4295(.din(new_new_n7098__), .dout(new_new_n7110__));
  buf1  g4296(.din(new_new_n7110__), .dout(new_new_n7111__));
  buf1  g4297(.din(new_new_n7111__), .dout(new_new_n7112__));
  buf1  g4298(.din(new_new_n7111__), .dout(new_new_n7113__));
  buf1  g4299(.din(new_new_n7110__), .dout(new_new_n7114__));
  buf1  g4300(.din(new_new_n7114__), .dout(new_new_n7115__));
  buf1  g4301(.din(new_new_n7114__), .dout(new_new_n7116__));
  buf1  g4302(.din(new_new_n3279__), .dout(new_new_n7117__));
  buf1  g4303(.din(new_new_n7117__), .dout(new_new_n7118__));
  buf1  g4304(.din(new_new_n7118__), .dout(new_new_n7119__));
  buf1  g4305(.din(new_new_n7119__), .dout(new_new_n7120__));
  buf1  g4306(.din(new_new_n7119__), .dout(new_new_n7121__));
  buf1  g4307(.din(new_new_n7118__), .dout(new_new_n7122__));
  buf1  g4308(.din(new_new_n7117__), .dout(new_new_n7123__));
  buf1  g4309(.din(new_new_n7123__), .dout(new_new_n7124__));
  buf1  g4310(.din(new_new_n7123__), .dout(new_new_n7125__));
  buf1  g4311(.din(new_new_n3278__), .dout(new_new_n7126__));
  buf1  g4312(.din(new_new_n7126__), .dout(new_new_n7127__));
  buf1  g4313(.din(new_new_n7127__), .dout(new_new_n7128__));
  buf1  g4314(.din(new_new_n7128__), .dout(new_new_n7129__));
  buf1  g4315(.din(new_new_n7128__), .dout(new_new_n7130__));
  buf1  g4316(.din(new_new_n7127__), .dout(new_new_n7131__));
  buf1  g4317(.din(new_new_n7126__), .dout(new_new_n7132__));
  buf1  g4318(.din(new_new_n7132__), .dout(new_new_n7133__));
  buf1  g4319(.din(new_new_n7132__), .dout(new_new_n7134__));
  buf1  g4320(.din(new_new_n2506__), .dout(new_new_n7135__));
  buf1  g4321(.din(new_new_n2522__), .dout(new_new_n7136__));
  buf1  g4322(.din(new_new_n4279__), .dout(new_new_n7137__));
  buf1  g4323(.din(new_new_n7137__), .dout(new_new_n7138__));
  buf1  g4324(.din(new_new_n7138__), .dout(new_new_n7139__));
  buf1  g4325(.din(new_new_n7137__), .dout(new_new_n7140__));
  buf1  g4326(.din(new_new_n4252__), .dout(new_new_n7141__));
  buf1  g4327(.din(new_new_n7141__), .dout(new_new_n7142__));
  buf1  g4328(.din(new_new_n7142__), .dout(new_new_n7143__));
  buf1  g4329(.din(new_new_n7141__), .dout(new_new_n7144__));
  buf1  g4330(.din(new_new_n2442__), .dout(new_new_n7145__));
  buf1  g4331(.din(new_new_n2606__), .dout(new_new_n7146__));
  buf1  g4332(.din(new_new_n4284__), .dout(new_new_n7147__));
  buf1  g4333(.din(new_new_n7147__), .dout(new_new_n7148__));
  buf1  g4334(.din(new_new_n7148__), .dout(new_new_n7149__));
  buf1  g4335(.din(new_new_n7147__), .dout(new_new_n7150__));
  buf1  g4336(.din(new_new_n4255__), .dout(new_new_n7151__));
  buf1  g4337(.din(new_new_n7151__), .dout(new_new_n7152__));
  buf1  g4338(.din(new_new_n7152__), .dout(new_new_n7153__));
  buf1  g4339(.din(new_new_n7151__), .dout(new_new_n7154__));
  buf1  g4340(.din(new_new_n2434__), .dout(new_new_n7155__));
  buf1  g4341(.din(new_new_n2598__), .dout(new_new_n7156__));
  buf1  g4342(.din(new_new_n4291__), .dout(new_new_n7157__));
  buf1  g4343(.din(new_new_n7157__), .dout(new_new_n7158__));
  buf1  g4344(.din(new_new_n7158__), .dout(new_new_n7159__));
  buf1  g4345(.din(new_new_n7157__), .dout(new_new_n7160__));
  buf1  g4346(.din(new_new_n4261__), .dout(new_new_n7161__));
  buf1  g4347(.din(new_new_n7161__), .dout(new_new_n7162__));
  buf1  g4348(.din(new_new_n7162__), .dout(new_new_n7163__));
  buf1  g4349(.din(new_new_n7161__), .dout(new_new_n7164__));
  buf1  g4350(.din(new_new_n2591__), .dout(new_new_n7165__));
  buf1  g4351(.din(new_new_n2583__), .dout(new_new_n7166__));
  buf1  g4352(.din(new_new_n4297__), .dout(new_new_n7167__));
  buf1  g4353(.din(new_new_n7167__), .dout(new_new_n7168__));
  buf1  g4354(.din(new_new_n7168__), .dout(new_new_n7169__));
  buf1  g4355(.din(new_new_n7167__), .dout(new_new_n7170__));
  buf1  g4356(.din(new_new_n4234__), .dout(new_new_n7171__));
  buf1  g4357(.din(new_new_n7171__), .dout(new_new_n7172__));
  buf1  g4358(.din(new_new_n7172__), .dout(new_new_n7173__));
  buf1  g4359(.din(new_new_n7171__), .dout(new_new_n7174__));
  buf1  g4360(.din(new_new_n2976__), .dout(new_new_n7175__));
  buf1  g4361(.din(new_new_n3056__), .dout(new_new_n7176__));
  buf1  g4362(.din(new_new_n2945__), .dout(new_new_n7177__));
  buf1  g4363(.din(new_new_n3025__), .dout(new_new_n7178__));
  buf1  g4364(.din(new_new_n2881__), .dout(new_new_n7179__));
  buf1  g4365(.din(new_new_n7179__), .dout(new_new_n7180__));
  buf1  g4366(.din(new_new_n7179__), .dout(new_new_n7181__));
  buf1  g4367(.din(new_new_n2928__), .dout(new_new_n7182__));
  buf1  g4368(.din(new_new_n2936__), .dout(new_new_n7183__));
  buf1  g4369(.din(new_new_n2912__), .dout(new_new_n7184__));
  buf1  g4370(.din(new_new_n2920__), .dout(new_new_n7185__));
  buf1  g4371(.din(new_new_n3347__), .dout(new_new_n7186__));
  buf1  g4372(.din(new_new_n3346__), .dout(new_new_n7187__));
  buf1  g4373(.din(new_new_n2857__), .dout(new_new_n7188__));
  buf1  g4374(.din(new_new_n2856__), .dout(new_new_n7189__));
  buf1  g4375(.din(new_new_n3463__), .dout(new_new_n7190__));
  buf1  g4376(.din(new_new_n4564__), .dout(new_new_n7191__));
  buf1  g4377(.din(new_new_n3083__), .dout(new_new_n7192__));
  buf1  g4378(.din(new_new_n3233__), .dout(new_new_n7193__));
  buf1  g4379(.din(new_new_n4138__), .dout(new_new_n7194__));
  buf1  g4380(.din(new_new_n4143__), .dout(new_new_n7195__));
  buf1  g4381(.din(new_new_n4202__), .dout(new_new_n7196__));
  buf1  g4382(.din(new_new_n4217__), .dout(new_new_n7197__));
  buf1  g4383(.din(new_new_n4318__), .dout(new_new_n7198__));
  buf1  g4384(.din(new_new_n4357__), .dout(new_new_n7199__));
  buf1  g4385(.din(new_new_n2718__), .dout(new_new_n7200__));
  buf1  g4386(.din(new_new_n2726__), .dout(new_new_n7201__));
  buf1  g4387(.din(new_new_n4597__), .dout(new_new_n7202__));
  buf1  g4388(.din(new_new_n7202__), .dout(new_new_n7203__));
  buf1  g4389(.din(new_new_n7203__), .dout(new_new_n7204__));
  buf1  g4390(.din(new_new_n7202__), .dout(new_new_n7205__));
  buf1  g4391(.din(new_new_n4576__), .dout(new_new_n7206__));
  buf1  g4392(.din(new_new_n7206__), .dout(new_new_n7207__));
  buf1  g4393(.din(new_new_n7207__), .dout(new_new_n7208__));
  buf1  g4394(.din(new_new_n7206__), .dout(new_new_n7209__));
  buf1  g4395(.din(new_new_n2538__), .dout(new_new_n7210__));
  buf1  g4396(.din(new_new_n2530__), .dout(new_new_n7211__));
  buf1  g4397(.din(new_new_n4603__), .dout(new_new_n7212__));
  buf1  g4398(.din(new_new_n7212__), .dout(new_new_n7213__));
  buf1  g4399(.din(new_new_n7213__), .dout(new_new_n7214__));
  buf1  g4400(.din(new_new_n7212__), .dout(new_new_n7215__));
  buf1  g4401(.din(new_new_n4580__), .dout(new_new_n7216__));
  buf1  g4402(.din(new_new_n7216__), .dout(new_new_n7217__));
  buf1  g4403(.din(new_new_n7217__), .dout(new_new_n7218__));
  buf1  g4404(.din(new_new_n7216__), .dout(new_new_n7219__));
  buf1  g4405(.din(new_new_n2710__), .dout(new_new_n7220__));
  buf1  g4406(.din(new_new_n2702__), .dout(new_new_n7221__));
  buf1  g4407(.din(new_new_n4609__), .dout(new_new_n7222__));
  buf1  g4408(.din(new_new_n7222__), .dout(new_new_n7223__));
  buf1  g4409(.din(new_new_n7223__), .dout(new_new_n7224__));
  buf1  g4410(.din(new_new_n7222__), .dout(new_new_n7225__));
  buf1  g4411(.din(new_new_n4584__), .dout(new_new_n7226__));
  buf1  g4412(.din(new_new_n7226__), .dout(new_new_n7227__));
  buf1  g4413(.din(new_new_n7227__), .dout(new_new_n7228__));
  buf1  g4414(.din(new_new_n7226__), .dout(new_new_n7229__));
  buf1  g4415(.din(new_new_n2514__), .dout(new_new_n7230__));
  buf1  g4416(.din(new_new_n2678__), .dout(new_new_n7231__));
  buf1  g4417(.din(new_new_n4613__), .dout(new_new_n7232__));
  buf1  g4418(.din(new_new_n7232__), .dout(new_new_n7233__));
  buf1  g4419(.din(new_new_n7233__), .dout(new_new_n7234__));
  buf1  g4420(.din(new_new_n7232__), .dout(new_new_n7235__));
  buf1  g4421(.din(new_new_n4587__), .dout(new_new_n7236__));
  buf1  g4422(.din(new_new_n7236__), .dout(new_new_n7237__));
  buf1  g4423(.din(new_new_n7237__), .dout(new_new_n7238__));
  buf1  g4424(.din(new_new_n7236__), .dout(new_new_n7239__));
  buf1  g4425(.din(new_new_n2984__), .dout(new_new_n7240__));
  buf1  g4426(.din(new_new_n3064__), .dout(new_new_n7241__));
  buf1  g4427(.din(new_new_n2968__), .dout(new_new_n7242__));
  buf1  g4428(.din(new_new_n3048__), .dout(new_new_n7243__));
  buf1  g4429(.din(new_new_n2960__), .dout(new_new_n7244__));
  buf1  g4430(.din(new_new_n3040__), .dout(new_new_n7245__));
  buf1  g4431(.din(new_new_n2952__), .dout(new_new_n7246__));
  buf1  g4432(.din(new_new_n3032__), .dout(new_new_n7247__));
  buf1  g4433(.din(new_new_n4767__), .dout(new_new_n7248__));
  buf1  g4434(.din(new_new_n4766__), .dout(new_new_n7249__));
  buf1  g4435(.din(new_new_n4772__), .dout(new_new_n7250__));
  buf1  g4436(.din(new_new_n2575__), .dout(new_new_n7251__));
  buf1  g4437(.din(new_new_n2427__), .dout(new_new_n7252__));
  buf1  g4438(.din(new_new_n4780__), .dout(new_new_n7253__));
  buf1  g4439(.din(new_new_n7253__), .dout(new_new_n7254__));
  buf1  g4440(.din(new_new_n7253__), .dout(new_new_n7255__));
  buf1  g4441(.din(new_new_n4783__), .dout(new_new_n7256__));
  buf1  g4442(.din(new_new_n7256__), .dout(new_new_n7257__));
  buf1  g4443(.din(new_new_n7256__), .dout(new_new_n7258__));
  buf1  g4444(.din(new_new_n3001__), .dout(new_new_n7259__));
  buf1  g4445(.din(new_new_n2993__), .dout(new_new_n7260__));
  buf1  g4446(.din(new_new_n3619__), .dout(new_new_n7261__));
  buf1  g4447(.din(new_new_n7261__), .dout(new_new_n7262__));
  buf1  g4448(.din(new_new_n7261__), .dout(new_new_n7263__));
  buf1  g4449(.din(new_new_n3965__), .dout(new_new_n7264__));
  buf1  g4450(.din(new_new_n3618__), .dout(new_new_n7265__));
  buf1  g4451(.din(new_new_n7265__), .dout(new_new_n7266__));
  buf1  g4452(.din(new_new_n3964__), .dout(new_new_n7267__));
  buf1  g4453(.din(new_new_n7267__), .dout(new_new_n7268__));
  buf1  g4454(.din(new_new_n4818__), .dout(new_new_n7269__));
  buf1  g4455(.din(new_new_n3555__), .dout(new_new_n7270__));
  buf1  g4456(.din(new_new_n7270__), .dout(new_new_n7271__));
  buf1  g4457(.din(new_new_n7271__), .dout(new_new_n7272__));
  buf1  g4458(.din(new_new_n7270__), .dout(new_new_n7273__));
  buf1  g4459(.din(new_new_n3647__), .dout(new_new_n7274__));
  buf1  g4460(.din(new_new_n2410__), .dout(new_new_n7275__));
  buf1  g4461(.din(new_new_n7275__), .dout(new_new_n7276__));
  buf1  g4462(.din(new_new_n7275__), .dout(new_new_n7277__));
  buf1  g4463(.din(new_new_n3572__), .dout(new_new_n7278__));
  buf1  g4464(.din(new_new_n4825__), .dout(new_new_n7279__));
  buf1  g4465(.din(new_new_n4083__), .dout(new_new_n7280__));
  buf1  g4466(.din(new_new_n4082__), .dout(new_new_n7281__));
  buf1  g4467(.din(new_new_n7281__), .dout(new_new_n7282__));
  buf1  g4468(.din(new_new_n4053__), .dout(new_new_n7283__));
  buf1  g4469(.din(new_new_n4052__), .dout(new_new_n7284__));
  buf1  g4470(.din(new_new_n4078__), .dout(new_new_n7285__));
  buf1  g4471(.din(new_new_n4084__), .dout(new_new_n7286__));
  buf1  g4472(.din(new_new_n7286__), .dout(new_new_n7287__));
  buf1  g4473(.din(new_new_n4088__), .dout(new_new_n7288__));
  buf1  g4474(.din(new_new_n4085__), .dout(new_new_n7289__));
  buf1  g4475(.din(new_new_n3938__), .dout(new_new_n7290__));
  buf1  g4476(.din(new_new_n7290__), .dout(new_new_n7291__));
  buf1  g4477(.din(new_new_n4839__), .dout(new_new_n7292__));
  buf1  g4478(.din(new_new_n7292__), .dout(new_new_n7293__));
  buf1  g4479(.din(new_new_n3939__), .dout(new_new_n7294__));
  buf1  g4480(.din(new_new_n4840__), .dout(new_new_n7295__));
  buf1  g4481(.din(new_new_n3331__), .dout(new_new_n7296__));
  buf1  g4482(.din(new_new_n7296__), .dout(new_new_n7297__));
  buf1  g4483(.din(new_new_n7297__), .dout(new_new_n7298__));
  buf1  g4484(.din(new_new_n7298__), .dout(new_new_n7299__));
  buf1  g4485(.din(new_new_n7298__), .dout(new_new_n7300__));
  buf1  g4486(.din(new_new_n7297__), .dout(new_new_n7301__));
  buf1  g4487(.din(new_new_n7301__), .dout(new_new_n7302__));
  buf1  g4488(.din(new_new_n7301__), .dout(new_new_n7303__));
  buf1  g4489(.din(new_new_n7296__), .dout(new_new_n7304__));
  buf1  g4490(.din(new_new_n7304__), .dout(new_new_n7305__));
  buf1  g4491(.din(new_new_n7304__), .dout(new_new_n7306__));
  buf1  g4492(.din(new_new_n3312__), .dout(new_new_n7307__));
  buf1  g4493(.din(new_new_n7307__), .dout(new_new_n7308__));
  buf1  g4494(.din(new_new_n7308__), .dout(new_new_n7309__));
  buf1  g4495(.din(new_new_n7309__), .dout(new_new_n7310__));
  buf1  g4496(.din(new_new_n7309__), .dout(new_new_n7311__));
  buf1  g4497(.din(new_new_n7308__), .dout(new_new_n7312__));
  buf1  g4498(.din(new_new_n7312__), .dout(new_new_n7313__));
  buf1  g4499(.din(new_new_n7312__), .dout(new_new_n7314__));
  buf1  g4500(.din(new_new_n7307__), .dout(new_new_n7315__));
  buf1  g4501(.din(new_new_n7315__), .dout(new_new_n7316__));
  buf1  g4502(.din(new_new_n7315__), .dout(new_new_n7317__));
  buf1  g4503(.din(new_new_n3644__), .dout(new_new_n7318__));
  buf1  g4504(.din(new_new_n7318__), .dout(new_new_n7319__));
  buf1  g4505(.din(new_new_n4056__), .dout(new_new_n7320__));
  buf1  g4506(.din(new_new_n7320__), .dout(new_new_n7321__));
  buf1  g4507(.din(new_new_n7321__), .dout(new_new_n7322__));
  buf1  g4508(.din(new_new_n7321__), .dout(new_new_n7323__));
  buf1  g4509(.din(new_new_n7320__), .dout(new_new_n7324__));
  buf1  g4510(.din(new_new_n3645__), .dout(new_new_n7325__));
  buf1  g4511(.din(new_new_n4057__), .dout(new_new_n7326__));
  buf1  g4512(.din(new_new_n7326__), .dout(new_new_n7327__));
  buf1  g4513(.din(new_new_n7327__), .dout(new_new_n7328__));
  buf1  g4514(.din(new_new_n7326__), .dout(new_new_n7329__));
  buf1  g4515(.din(new_new_n3948__), .dout(new_new_n7330__));
  buf1  g4516(.din(new_new_n3764__), .dout(new_new_n7331__));
  buf1  g4517(.din(new_new_n4830__), .dout(new_new_n7332__));
  buf1  g4518(.din(new_new_n7332__), .dout(new_new_n7333__));
  buf1  g4519(.din(new_new_n7332__), .dout(new_new_n7334__));
  buf1  g4520(.din(new_new_n4829__), .dout(new_new_n7335__));
  buf1  g4521(.din(new_new_n7335__), .dout(new_new_n7336__));
  buf1  g4522(.din(new_new_n4025__), .dout(new_new_n7337__));
  buf1  g4523(.din(new_new_n4024__), .dout(new_new_n7338__));
  buf1  g4524(.din(new_new_n3988__), .dout(new_new_n7339__));
  buf1  g4525(.din(new_new_n7339__), .dout(new_new_n7340__));
  buf1  g4526(.din(new_new_n7339__), .dout(new_new_n7341__));
  buf1  g4527(.din(new_new_n4029__), .dout(new_new_n7342__));
  buf1  g4528(.din(new_new_n3989__), .dout(new_new_n7343__));
  buf1  g4529(.din(new_new_n7343__), .dout(new_new_n7344__));
  buf1  g4530(.din(new_new_n4028__), .dout(new_new_n7345__));
  buf1  g4531(.din(new_new_n4030__), .dout(new_new_n7346__));
  buf1  g4532(.din(new_new_n7346__), .dout(new_new_n7347__));
  buf1  g4533(.din(new_new_n7347__), .dout(new_new_n7348__));
  buf1  g4534(.din(new_new_n7346__), .dout(new_new_n7349__));
  buf1  g4535(.din(new_new_n4834__), .dout(new_new_n7350__));
  buf1  g4536(.din(new_new_n7350__), .dout(new_new_n7351__));
  buf1  g4537(.din(new_new_n4031__), .dout(new_new_n7352__));
  buf1  g4538(.din(new_new_n7352__), .dout(new_new_n7353__));
  buf1  g4539(.din(new_new_n7352__), .dout(new_new_n7354__));
  buf1  g4540(.din(new_new_n4833__), .dout(new_new_n7355__));
  buf1  g4541(.din(new_new_n4865__), .dout(new_new_n7356__));
  buf1  g4542(.din(new_new_n4864__), .dout(new_new_n7357__));
  buf1  g4543(.din(new_new_n4826__), .dout(new_new_n7358__));
  buf1  g4544(.din(new_new_n3604__), .dout(new_new_n7359__));
  buf1  g4545(.din(new_new_n4876__), .dout(new_new_n7360__));
  buf1  g4546(.din(new_new_n3936__), .dout(new_new_n7361__));
  buf1  g4547(.din(new_new_n7361__), .dout(new_new_n7362__));
  buf1  g4548(.din(new_new_n7361__), .dout(new_new_n7363__));
  buf1  g4549(.din(new_new_n4086__), .dout(new_new_n7364__));
  buf1  g4550(.din(new_new_n7364__), .dout(new_new_n7365__));
  buf1  g4551(.din(new_new_n7364__), .dout(new_new_n7366__));
  buf1  g4552(.din(new_new_n3937__), .dout(new_new_n7367__));
  buf1  g4553(.din(new_new_n4087__), .dout(new_new_n7368__));
  buf1  g4554(.din(new_new_n3590__), .dout(new_new_n7369__));
  buf1  g4555(.din(new_new_n7369__), .dout(new_new_n7370__));
  buf1  g4556(.din(new_new_n3511__), .dout(new_new_n7371__));
  buf1  g4557(.din(new_new_n7371__), .dout(new_new_n7372__));
  buf1  g4558(.din(new_new_n7371__), .dout(new_new_n7373__));
  buf1  g4559(.din(new_new_n3325__), .dout(new_new_n7374__));
  buf1  g4560(.din(new_new_n7374__), .dout(new_new_n7375__));
  buf1  g4561(.din(new_new_n7375__), .dout(new_new_n7376__));
  buf1  g4562(.din(new_new_n7376__), .dout(new_new_n7377__));
  buf1  g4563(.din(new_new_n7376__), .dout(new_new_n7378__));
  buf1  g4564(.din(new_new_n7375__), .dout(new_new_n7379__));
  buf1  g4565(.din(new_new_n7379__), .dout(new_new_n7380__));
  buf1  g4566(.din(new_new_n7374__), .dout(new_new_n7381__));
  buf1  g4567(.din(new_new_n7381__), .dout(new_new_n7382__));
  buf1  g4568(.din(new_new_n7381__), .dout(new_new_n7383__));
  buf1  g4569(.din(new_new_n3510__), .dout(new_new_n7384__));
  buf1  g4570(.din(new_new_n7384__), .dout(new_new_n7385__));
  buf1  g4571(.din(new_new_n7384__), .dout(new_new_n7386__));
  buf1  g4572(.din(new_new_n3318__), .dout(new_new_n7387__));
  buf1  g4573(.din(new_new_n7387__), .dout(new_new_n7388__));
  buf1  g4574(.din(new_new_n7388__), .dout(new_new_n7389__));
  buf1  g4575(.din(new_new_n7389__), .dout(new_new_n7390__));
  buf1  g4576(.din(new_new_n7389__), .dout(new_new_n7391__));
  buf1  g4577(.din(new_new_n7388__), .dout(new_new_n7392__));
  buf1  g4578(.din(new_new_n7392__), .dout(new_new_n7393__));
  buf1  g4579(.din(new_new_n7387__), .dout(new_new_n7394__));
  buf1  g4580(.din(new_new_n7394__), .dout(new_new_n7395__));
  buf1  g4581(.din(new_new_n7394__), .dout(new_new_n7396__));
  buf1  g4582(.din(new_new_n3453__), .dout(new_new_n7397__));
  buf1  g4583(.din(new_new_n7397__), .dout(new_new_n7398__));
  buf1  g4584(.din(new_new_n3452__), .dout(new_new_n7399__));
  buf1  g4585(.din(new_new_n7399__), .dout(new_new_n7400__));
  buf1  g4586(.din(new_new_n3579__), .dout(new_new_n7401__));
  buf1  g4587(.din(new_new_n7401__), .dout(new_new_n7402__));
  buf1  g4588(.din(new_new_n3578__), .dout(new_new_n7403__));
  buf1  g4589(.din(new_new_n7403__), .dout(new_new_n7404__));
  buf1  g4590(.din(new_new_n3178__), .dout(new_new_n7405__));
  buf1  g4591(.din(new_new_n7405__), .dout(new_new_n7406__));
  buf1  g4592(.din(new_new_n7406__), .dout(new_new_n7407__));
  buf1  g4593(.din(new_new_n7405__), .dout(new_new_n7408__));
  buf1  g4594(.din(new_new_n4853__), .dout(new_new_n7409__));
  buf1  g4595(.din(new_new_n7409__), .dout(new_new_n7410__));
  buf1  g4596(.din(new_new_n3179__), .dout(new_new_n7411__));
  buf1  g4597(.din(new_new_n7411__), .dout(new_new_n7412__));
  buf1  g4598(.din(new_new_n7411__), .dout(new_new_n7413__));
  buf1  g4599(.din(new_new_n4852__), .dout(new_new_n7414__));
  buf1  g4600(.din(new_new_n4910__), .dout(new_new_n7415__));
  buf1  g4601(.din(new_new_n4076__), .dout(new_new_n7416__));
  buf1  g4602(.din(new_new_n7416__), .dout(new_new_n7417__));
  buf1  g4603(.din(new_new_n7417__), .dout(new_new_n7418__));
  buf1  g4604(.din(new_new_n7418__), .dout(new_new_n7419__));
  buf1  g4605(.din(new_new_n7418__), .dout(new_new_n7420__));
  buf1  g4606(.din(new_new_n7417__), .dout(new_new_n7421__));
  buf1  g4607(.din(new_new_n7416__), .dout(new_new_n7422__));
  buf1  g4608(.din(new_new_n7422__), .dout(new_new_n7423__));
  buf1  g4609(.din(new_new_n7422__), .dout(new_new_n7424__));
  buf1  g4610(.din(new_new_n4116__), .dout(new_new_n7425__));
  buf1  g4611(.din(new_new_n4077__), .dout(new_new_n7426__));
  buf1  g4612(.din(new_new_n7426__), .dout(new_new_n7427__));
  buf1  g4613(.din(new_new_n7427__), .dout(new_new_n7428__));
  buf1  g4614(.din(new_new_n7428__), .dout(new_new_n7429__));
  buf1  g4615(.din(new_new_n7427__), .dout(new_new_n7430__));
  buf1  g4616(.din(new_new_n7426__), .dout(new_new_n7431__));
  buf1  g4617(.din(new_new_n7431__), .dout(new_new_n7432__));
  buf1  g4618(.din(new_new_n7431__), .dout(new_new_n7433__));
  buf1  g4619(.din(new_new_n4112__), .dout(new_new_n7434__));
  buf1  g4620(.din(new_new_n7434__), .dout(new_new_n7435__));
  buf1  g4621(.din(new_new_n4873__), .dout(new_new_n7436__));
  buf1  g4622(.din(new_new_n7436__), .dout(new_new_n7437__));
  buf1  g4623(.din(new_new_n4114__), .dout(new_new_n7438__));
  buf1  g4624(.din(new_new_n7438__), .dout(new_new_n7439__));
  buf1  g4625(.din(new_new_n4871__), .dout(new_new_n7440__));
  buf1  g4626(.din(new_new_n7440__), .dout(new_new_n7441__));
  buf1  g4627(.din(new_new_n4120__), .dout(new_new_n7442__));
  buf1  g4628(.din(new_new_n4124__), .dout(new_new_n7443__));
  buf1  g4629(.din(new_new_n7443__), .dout(new_new_n7444__));
  buf1  g4630(.din(new_new_n7444__), .dout(new_new_n7445__));
  buf1  g4631(.din(new_new_n7445__), .dout(new_new_n7446__));
  buf1  g4632(.din(new_new_n7445__), .dout(new_new_n7447__));
  buf1  g4633(.din(new_new_n7444__), .dout(new_new_n7448__));
  buf1  g4634(.din(new_new_n7448__), .dout(new_new_n7449__));
  buf1  g4635(.din(new_new_n7448__), .dout(new_new_n7450__));
  buf1  g4636(.din(new_new_n7443__), .dout(new_new_n7451__));
  buf1  g4637(.din(new_new_n7451__), .dout(new_new_n7452__));
  buf1  g4638(.din(new_new_n7451__), .dout(new_new_n7453__));
  buf1  g4639(.din(new_new_n4125__), .dout(new_new_n7454__));
  buf1  g4640(.din(new_new_n7454__), .dout(new_new_n7455__));
  buf1  g4641(.din(new_new_n7455__), .dout(new_new_n7456__));
  buf1  g4642(.din(new_new_n7456__), .dout(new_new_n7457__));
  buf1  g4643(.din(new_new_n7456__), .dout(new_new_n7458__));
  buf1  g4644(.din(new_new_n7455__), .dout(new_new_n7459__));
  buf1  g4645(.din(new_new_n7459__), .dout(new_new_n7460__));
  buf1  g4646(.din(new_new_n7454__), .dout(new_new_n7461__));
  buf1  g4647(.din(new_new_n7461__), .dout(new_new_n7462__));
  buf1  g4648(.din(new_new_n7461__), .dout(new_new_n7463__));
  buf1  g4649(.din(new_new_n4841__), .dout(new_new_n7464__));
  buf1  g4650(.din(new_new_n4868__), .dout(new_new_n7465__));
  buf1  g4651(.din(new_new_n7465__), .dout(new_new_n7466__));
  buf1  g4652(.din(new_new_n4941__), .dout(new_new_n7467__));
  buf1  g4653(.din(new_new_n4869__), .dout(new_new_n7468__));
  buf1  g4654(.din(new_new_n4940__), .dout(new_new_n7469__));
  buf1  g4655(.din(new_new_n4943__), .dout(new_new_n7470__));
  buf1  g4656(.din(new_new_n4942__), .dout(new_new_n7471__));
  buf1  g4657(.din(new_new_n4098__), .dout(new_new_n7472__));
  buf1  g4658(.din(new_new_n4102__), .dout(new_new_n7473__));
  buf1  g4659(.din(new_new_n4831__), .dout(new_new_n7474__));
  buf1  g4660(.din(new_new_n7474__), .dout(new_new_n7475__));
  buf1  g4661(.din(new_new_n4958__), .dout(new_new_n7476__));
  buf1  g4662(.din(new_new_n4832__), .dout(new_new_n7477__));
  buf1  g4663(.din(new_new_n7477__), .dout(new_new_n7478__));
  buf1  g4664(.din(new_new_n7477__), .dout(new_new_n7479__));
  buf1  g4665(.din(new_new_n4959__), .dout(new_new_n7480__));
  buf1  g4666(.din(new_new_n4854__), .dout(new_new_n7481__));
  buf1  g4667(.din(new_new_n7481__), .dout(new_new_n7482__));
  buf1  g4668(.din(new_new_n4966__), .dout(new_new_n7483__));
  buf1  g4669(.din(new_new_n4106__), .dout(new_new_n7484__));
  buf1  g4670(.din(new_new_n4094__), .dout(new_new_n7485__));
  buf1  g4671(.din(new_new_n7485__), .dout(new_new_n7486__));
  buf1  g4672(.din(new_new_n4921__), .dout(new_new_n7487__));
  buf1  g4673(.din(new_new_n7487__), .dout(new_new_n7488__));
  buf1  g4674(.din(new_new_n4110__), .dout(new_new_n7489__));
  buf1  g4675(.din(new_new_n7489__), .dout(new_new_n7490__));
  buf1  g4676(.din(new_new_n4875__), .dout(new_new_n7491__));
  buf1  g4677(.din(new_new_n7491__), .dout(new_new_n7492__));
  buf1  g4678(.din(new_new_n4924__), .dout(new_new_n7493__));
  buf1  g4679(.din(new_new_n7493__), .dout(new_new_n7494__));
  buf1  g4680(.din(new_new_n7493__), .dout(new_new_n7495__));
  buf1  g4681(.din(new_new_n4090__), .dout(new_new_n7496__));
  buf1  g4682(.din(new_new_n4092__), .dout(new_new_n7497__));
  buf1  g4683(.din(new_new_n3174__), .dout(new_new_n7498__));
  buf1  g4684(.din(new_new_n7498__), .dout(new_new_n7499__));
  buf1  g4685(.din(new_new_n4957__), .dout(new_new_n7500__));
  buf1  g4686(.din(new_new_n7500__), .dout(new_new_n7501__));
  buf1  g4687(.din(new_new_n3182__), .dout(new_new_n7502__));
  buf1  g4688(.din(new_new_n7502__), .dout(new_new_n7503__));
  buf1  g4689(.din(new_new_n4951__), .dout(new_new_n7504__));
  buf1  g4690(.din(new_new_n7504__), .dout(new_new_n7505__));
  buf1  g4691(.din(new_new_n3184__), .dout(new_new_n7506__));
  buf1  g4692(.din(new_new_n7506__), .dout(new_new_n7507__));
  buf1  g4693(.din(new_new_n4971__), .dout(new_new_n7508__));
  buf1  g4694(.din(new_new_n7508__), .dout(new_new_n7509__));
  buf1  g4695(.din(new_new_n4096__), .dout(new_new_n7510__));
  buf1  g4696(.din(new_new_n7510__), .dout(new_new_n7511__));
  buf1  g4697(.din(new_new_n4932__), .dout(new_new_n7512__));
  buf1  g4698(.din(new_new_n7512__), .dout(new_new_n7513__));
  buf1  g4699(.din(new_new_n4998__), .dout(new_new_n7514__));
  buf1  g4700(.din(new_new_n4982__), .dout(new_new_n7515__));
  buf1  g4701(.din(new_new_n4984__), .dout(new_new_n7516__));
  buf1  g4702(.din(new_new_n7516__), .dout(new_new_n7517__));
  buf1  g4703(.din(new_new_n3393__), .dout(new_new_n7518__));
  buf1  g4704(.din(new_new_n7518__), .dout(new_new_n7519__));
  buf1  g4705(.din(new_new_n7519__), .dout(new_new_n7520__));
  buf1  g4706(.din(new_new_n7520__), .dout(new_new_n7521__));
  buf1  g4707(.din(new_new_n7520__), .dout(new_new_n7522__));
  buf1  g4708(.din(new_new_n7519__), .dout(new_new_n7523__));
  buf1  g4709(.din(new_new_n7523__), .dout(new_new_n7524__));
  buf1  g4710(.din(new_new_n7518__), .dout(new_new_n7525__));
  buf1  g4711(.din(new_new_n7525__), .dout(new_new_n7526__));
  buf1  g4712(.din(new_new_n7525__), .dout(new_new_n7527__));
  buf1  g4713(.din(new_new_n3392__), .dout(new_new_n7528__));
  buf1  g4714(.din(new_new_n7528__), .dout(new_new_n7529__));
  buf1  g4715(.din(new_new_n7529__), .dout(new_new_n7530__));
  buf1  g4716(.din(new_new_n7530__), .dout(new_new_n7531__));
  buf1  g4717(.din(new_new_n7530__), .dout(new_new_n7532__));
  buf1  g4718(.din(new_new_n7529__), .dout(new_new_n7533__));
  buf1  g4719(.din(new_new_n7533__), .dout(new_new_n7534__));
  buf1  g4720(.din(new_new_n7533__), .dout(new_new_n7535__));
  buf1  g4721(.din(new_new_n7528__), .dout(new_new_n7536__));
  buf1  g4722(.din(new_new_n7536__), .dout(new_new_n7537__));
  buf1  g4723(.din(new_new_n7537__), .dout(new_new_n7538__));
  buf1  g4724(.din(new_new_n7537__), .dout(new_new_n7539__));
  buf1  g4725(.din(new_new_n7536__), .dout(new_new_n7540__));
  buf1  g4726(.din(new_new_n3455__), .dout(new_new_n7541__));
  buf1  g4727(.din(new_new_n7541__), .dout(new_new_n7542__));
  buf1  g4728(.din(new_new_n3454__), .dout(new_new_n7543__));
  buf1  g4729(.din(new_new_n7543__), .dout(new_new_n7544__));
  buf1  g4730(.din(new_new_n3385__), .dout(new_new_n7545__));
  buf1  g4731(.din(new_new_n7545__), .dout(new_new_n7546__));
  buf1  g4732(.din(new_new_n2806__), .dout(new_new_n7547__));
  buf1  g4733(.din(new_new_n3384__), .dout(new_new_n7548__));
  buf1  g4734(.din(new_new_n7548__), .dout(new_new_n7549__));
  buf1  g4735(.din(new_new_n3607__), .dout(new_new_n7550__));
  buf1  g4736(.din(new_new_n3606__), .dout(new_new_n7551__));
  buf1  g4737(.din(new_new_n3608__), .dout(new_new_n7552__));
  buf1  g4738(.din(new_new_n7552__), .dout(new_new_n7553__));
  buf1  g4739(.din(new_new_n3628__), .dout(new_new_n7554__));
  buf1  g4740(.din(new_new_n3980__), .dout(new_new_n7555__));
  buf1  g4741(.din(new_new_n4020__), .dout(new_new_n7556__));
  buf1  g4742(.din(new_new_n3981__), .dout(new_new_n7557__));
  buf1  g4743(.din(new_new_n4021__), .dout(new_new_n7558__));
  buf1  g4744(.din(new_new_n5023__), .dout(new_new_n7559__));
  buf1  g4745(.din(new_new_n5030__), .dout(new_new_n7560__));
  buf1  g4746(.din(new_new_n5024__), .dout(new_new_n7561__));
  buf1  g4747(.din(new_new_n5029__), .dout(new_new_n7562__));
  buf1  g4748(.din(new_new_n3554__), .dout(new_new_n7563__));
  buf1  g4749(.din(new_new_n4821__), .dout(new_new_n7564__));
  buf1  g4750(.din(new_new_n7564__), .dout(new_new_n7565__));
  buf1  g4751(.din(new_new_n5042__), .dout(new_new_n7566__));
  buf1  g4752(.din(new_new_n4822__), .dout(new_new_n7567__));
  buf1  g4753(.din(new_new_n7567__), .dout(new_new_n7568__));
  buf1  g4754(.din(new_new_n5041__), .dout(new_new_n7569__));
  buf1  g4755(.din(new_new_n4909__), .dout(new_new_n7570__));
  buf1  g4756(.din(new_new_n4891__), .dout(new_new_n7571__));
  buf1  g4757(.din(new_new_n4900__), .dout(new_new_n7572__));
  buf1  g4758(.din(new_new_n5059__), .dout(new_new_n7573__));
  buf1  g4759(.din(new_new_n5062__), .dout(new_new_n7574__));
  buf1  g4760(.din(new_new_n5060__), .dout(new_new_n7575__));
  buf1  g4761(.din(new_new_n5061__), .dout(new_new_n7576__));
  buf1  g4762(.din(new_new_n4002__), .dout(new_new_n7577__));
  buf1  g4763(.din(new_new_n3998__), .dout(new_new_n7578__));
  buf1  g4764(.din(new_new_n5069__), .dout(new_new_n7579__));
  buf1  g4765(.din(new_new_n5071__), .dout(new_new_n7580__));
  buf1  g4766(.din(new_new_n5070__), .dout(new_new_n7581__));
  buf1  g4767(.din(new_new_n5072__), .dout(new_new_n7582__));
  buf1  g4768(.din(new_new_n3942__), .dout(new_new_n7583__));
  buf1  g4769(.din(new_new_n7583__), .dout(new_new_n7584__));
  buf1  g4770(.din(new_new_n7583__), .dout(new_new_n7585__));
  buf1  g4771(.din(new_new_n2411__), .dout(new_new_n7586__));
  buf1  g4772(.din(new_new_n3943__), .dout(new_new_n7587__));
  buf1  g4773(.din(new_new_n7587__), .dout(new_new_n7588__));
  buf1  g4774(.din(new_new_n3941__), .dout(new_new_n7589__));
  buf1  g4775(.din(new_new_n7589__), .dout(new_new_n7590__));
  buf1  g4776(.din(new_new_n7589__), .dout(new_new_n7591__));
  buf1  g4777(.din(new_new_n3940__), .dout(new_new_n7592__));
  buf1  g4778(.din(new_new_n7592__), .dout(new_new_n7593__));
  buf1  g4779(.din(new_new_n7593__), .dout(new_new_n7594__));
  buf1  g4780(.din(new_new_n7592__), .dout(new_new_n7595__));
  buf1  g4781(.din(new_new_n5089__), .dout(new_new_n7596__));
  buf1  g4782(.din(new_new_n7596__), .dout(new_new_n7597__));
  buf1  g4783(.din(new_new_n7597__), .dout(new_new_n7598__));
  buf1  g4784(.din(new_new_n7596__), .dout(new_new_n7599__));
  buf1  g4785(.din(new_new_n5088__), .dout(new_new_n7600__));
  buf1  g4786(.din(new_new_n7600__), .dout(new_new_n7601__));
  buf1  g4787(.din(new_new_n7601__), .dout(new_new_n7602__));
  buf1  g4788(.din(new_new_n7600__), .dout(new_new_n7603__));
  buf1  g4789(.din(new_new_n3716__), .dout(new_new_n7604__));
  buf1  g4790(.din(new_new_n3717__), .dout(new_new_n7605__));
  buf1  g4791(.din(new_new_n7605__), .dout(new_new_n7606__));
  buf1  g4792(.din(new_new_n5094__), .dout(new_new_n7607__));
  buf1  g4793(.din(new_new_n4877__), .dout(new_new_n7608__));
  buf1  g4794(.din(new_new_n3148__), .dout(new_new_n7609__));
  buf1  g4795(.din(new_new_n7609__), .dout(new_new_n7610__));
  buf1  g4796(.din(new_new_n5101__), .dout(new_new_n7611__));
  buf1  g4797(.din(new_new_n3616__), .dout(new_new_n7612__));
  buf1  g4798(.din(new_new_n4823__), .dout(new_new_n7613__));
  buf1  g4799(.din(new_new_n5108__), .dout(new_new_n7614__));
  buf1  g4800(.din(new_new_n4882__), .dout(new_new_n7615__));
  buf1  g4801(.din(new_new_n3582__), .dout(new_new_n7616__));
  buf1  g4802(.din(new_new_n5113__), .dout(new_new_n7617__));
  buf1  g4803(.din(new_new_n3126__), .dout(new_new_n7618__));
  buf1  g4804(.din(new_new_n3979__), .dout(new_new_n7619__));
  buf1  g4805(.din(new_new_n7619__), .dout(new_new_n7620__));
  buf1  g4806(.din(new_new_n4847__), .dout(new_new_n7621__));
  buf1  g4807(.din(new_new_n3476__), .dout(new_new_n7622__));
  buf1  g4808(.din(new_new_n7622__), .dout(new_new_n7623__));
  buf1  g4809(.din(new_new_n3477__), .dout(new_new_n7624__));
  buf1  g4810(.din(new_new_n7624__), .dout(new_new_n7625__));
  buf1  g4811(.din(new_new_n3450__), .dout(new_new_n7626__));
  buf1  g4812(.din(new_new_n7626__), .dout(new_new_n7627__));
  buf1  g4813(.din(new_new_n3451__), .dout(new_new_n7628__));
  buf1  g4814(.din(new_new_n7628__), .dout(new_new_n7629__));
  buf1  g4815(.din(new_new_n3478__), .dout(new_new_n7630__));
  buf1  g4816(.din(new_new_n7630__), .dout(new_new_n7631__));
  buf1  g4817(.din(new_new_n3479__), .dout(new_new_n7632__));
  buf1  g4818(.din(new_new_n7632__), .dout(new_new_n7633__));
  buf1  g4819(.din(new_new_n3471__), .dout(new_new_n7634__));
  buf1  g4820(.din(new_new_n7634__), .dout(new_new_n7635__));
  buf1  g4821(.din(new_new_n7634__), .dout(new_new_n7636__));
  buf1  g4822(.din(new_new_n3470__), .dout(new_new_n7637__));
  buf1  g4823(.din(new_new_n7637__), .dout(new_new_n7638__));
  buf1  g4824(.din(new_new_n7637__), .dout(new_new_n7639__));
  buf1  g4825(.din(new_new_n3595__), .dout(new_new_n7640__));
  buf1  g4826(.din(new_new_n7640__), .dout(new_new_n7641__));
  buf1  g4827(.din(new_new_n7640__), .dout(new_new_n7642__));
  buf1  g4828(.din(new_new_n3594__), .dout(new_new_n7643__));
  buf1  g4829(.din(new_new_n7643__), .dout(new_new_n7644__));
  buf1  g4830(.din(new_new_n7643__), .dout(new_new_n7645__));
  buf1  g4831(.din(new_new_n3513__), .dout(new_new_n7646__));
  buf1  g4832(.din(new_new_n7646__), .dout(new_new_n7647__));
  buf1  g4833(.din(new_new_n3512__), .dout(new_new_n7648__));
  buf1  g4834(.din(new_new_n7648__), .dout(new_new_n7649__));
  buf1  g4835(.din(new_new_n3497__), .dout(new_new_n7650__));
  buf1  g4836(.din(new_new_n7650__), .dout(new_new_n7651__));
  buf1  g4837(.din(new_new_n3496__), .dout(new_new_n7652__));
  buf1  g4838(.din(new_new_n7652__), .dout(new_new_n7653__));
  buf1  g4839(.din(new_new_n3969__), .dout(new_new_n7654__));
  buf1  g4840(.din(new_new_n3970__), .dout(new_new_n7655__));
  buf1  g4841(.din(new_new_n3968__), .dout(new_new_n7656__));
  buf1  g4842(.din(new_new_n3971__), .dout(new_new_n7657__));
  buf1  g4843(.din(new_new_n3977__), .dout(new_new_n7658__));
  buf1  g4844(.din(new_new_n3976__), .dout(new_new_n7659__));
  buf1  g4845(.din(new_new_n3978__), .dout(new_new_n7660__));
  buf1  g4846(.din(new_new_n7660__), .dout(new_new_n7661__));
  buf1  g4847(.din(new_new_n5204__), .dout(new_new_n7662__));
  buf1  g4848(.din(new_new_n5209__), .dout(new_new_n7663__));
  buf1  g4849(.din(new_new_n5203__), .dout(new_new_n7664__));
  buf1  g4850(.din(new_new_n5210__), .dout(new_new_n7665__));
  buf1  g4851(.din(new_new_n3967__), .dout(new_new_n7666__));
  buf1  g4852(.din(new_new_n3974__), .dout(new_new_n7667__));
  buf1  g4853(.din(new_new_n3966__), .dout(new_new_n7668__));
  buf1  g4854(.din(new_new_n3975__), .dout(new_new_n7669__));
  buf1  g4855(.din(new_new_n3973__), .dout(new_new_n7670__));
  buf1  g4856(.din(new_new_n4019__), .dout(new_new_n7671__));
  buf1  g4857(.din(new_new_n3972__), .dout(new_new_n7672__));
  buf1  g4858(.din(new_new_n4018__), .dout(new_new_n7673__));
  buf1  g4859(.din(new_new_n5221__), .dout(new_new_n7674__));
  buf1  g4860(.din(new_new_n5228__), .dout(new_new_n7675__));
  buf1  g4861(.din(new_new_n5222__), .dout(new_new_n7676__));
  buf1  g4862(.din(new_new_n5227__), .dout(new_new_n7677__));
  buf1  g4863(.din(new_new_n3098__), .dout(new_new_n7678__));
  buf1  g4864(.din(new_new_n7678__), .dout(new_new_n7679__));
  buf1  g4865(.din(new_new_n3456__), .dout(new_new_n7680__));
  buf1  g4866(.din(new_new_n3099__), .dout(new_new_n7681__));
  buf1  g4867(.din(new_new_n7681__), .dout(new_new_n7682__));
  buf1  g4868(.din(new_new_n3457__), .dout(new_new_n7683__));
  buf1  g4869(.din(new_new_n3614__), .dout(new_new_n7684__));
  buf1  g4870(.din(new_new_n3626__), .dout(new_new_n7685__));
  buf1  g4871(.din(new_new_n3678__), .dout(new_new_n7686__));
  buf1  g4872(.din(new_new_n5279__), .dout(new_new_n7687__));
  buf1  g4873(.din(new_new_n5282__), .dout(new_new_n7688__));
  buf1  g4874(.din(new_new_n3149__), .dout(new_new_n7689__));
  buf1  g4875(.din(new_new_n3540__), .dout(new_new_n7690__));
  buf1  g4876(.din(new_new_n3541__), .dout(new_new_n7691__));
  buf1  g4877(.din(new_new_n5293__), .dout(new_new_n7692__));
  buf1  g4878(.din(new_new_n5296__), .dout(new_new_n7693__));
  buf1  g4879(.din(new_new_n5301__), .dout(new_new_n7694__));
  buf1  g4880(.din(new_new_n5304__), .dout(new_new_n7695__));
  buf1  g4881(.din(new_new_n5322__), .dout(new_new_n7696__));
  buf1  g4882(.din(new_new_n5325__), .dout(new_new_n7697__));
  buf1  g4883(.din(new_new_n5323__), .dout(new_new_n7698__));
  buf1  g4884(.din(new_new_n5324__), .dout(new_new_n7699__));
  buf1  g4885(.din(new_new_n3247__), .dout(new_new_n7700__));
  buf1  g4886(.din(new_new_n7700__), .dout(new_new_n7701__));
  buf1  g4887(.din(new_new_n7700__), .dout(new_new_n7702__));
  buf1  g4888(.din(new_new_n3246__), .dout(new_new_n7703__));
  buf1  g4889(.din(new_new_n7703__), .dout(new_new_n7704__));
  buf1  g4890(.din(new_new_n7703__), .dout(new_new_n7705__));
  buf1  g4891(.din(new_new_n5334__), .dout(new_new_n7706__));
  buf1  g4892(.din(new_new_n5336__), .dout(new_new_n7707__));
  buf1  g4893(.din(new_new_n5335__), .dout(new_new_n7708__));
  buf1  g4894(.din(new_new_n5337__), .dout(new_new_n7709__));
  buf1  g4895(.din(new_new_n5349__), .dout(new_new_n7710__));
  buf1  g4896(.din(new_new_n5348__), .dout(new_new_n7711__));
  buf1  g4897(.din(new_new_n5354__), .dout(new_new_n7712__));
  buf1  g4898(.din(new_new_n5355__), .dout(new_new_n7713__));
  buf1  g4899(.din(new_new_n4976__), .dout(new_new_n7714__));
  buf1  g4900(.din(new_new_n4981__), .dout(new_new_n7715__));
  buf1  g4901(.din(new_new_n7715__), .dout(new_new_n7716__));
  buf1  g4902(.din(new_new_n4922__), .dout(new_new_n7717__));
  buf1  g4903(.din(new_new_n3655__), .dout(new_new_n7718__));
  buf1  g4904(.din(new_new_n4063__), .dout(new_new_n7719__));
  buf1  g4905(.din(new_new_n7719__), .dout(new_new_n7720__));
  buf1  g4906(.din(new_new_n7720__), .dout(new_new_n7721__));
  buf1  g4907(.din(new_new_n7721__), .dout(new_new_n7722__));
  buf1  g4908(.din(new_new_n7721__), .dout(new_new_n7723__));
  buf1  g4909(.din(new_new_n7720__), .dout(new_new_n7724__));
  buf1  g4910(.din(new_new_n7724__), .dout(new_new_n7725__));
  buf1  g4911(.din(new_new_n7724__), .dout(new_new_n7726__));
  buf1  g4912(.din(new_new_n7719__), .dout(new_new_n7727__));
  buf1  g4913(.din(new_new_n7727__), .dout(new_new_n7728__));
  buf1  g4914(.din(new_new_n7728__), .dout(new_new_n7729__));
  buf1  g4915(.din(new_new_n7728__), .dout(new_new_n7730__));
  buf1  g4916(.din(new_new_n7727__), .dout(new_new_n7731__));
  buf1  g4917(.din(new_new_n7731__), .dout(new_new_n7732__));
  buf1  g4918(.din(new_new_n7731__), .dout(new_new_n7733__));
  buf1  g4919(.din(new_new_n3654__), .dout(new_new_n7734__));
  buf1  g4920(.din(new_new_n7734__), .dout(new_new_n7735__));
  buf1  g4921(.din(new_new_n4065__), .dout(new_new_n7736__));
  buf1  g4922(.din(new_new_n7736__), .dout(new_new_n7737__));
  buf1  g4923(.din(new_new_n7737__), .dout(new_new_n7738__));
  buf1  g4924(.din(new_new_n7738__), .dout(new_new_n7739__));
  buf1  g4925(.din(new_new_n7738__), .dout(new_new_n7740__));
  buf1  g4926(.din(new_new_n7737__), .dout(new_new_n7741__));
  buf1  g4927(.din(new_new_n7741__), .dout(new_new_n7742__));
  buf1  g4928(.din(new_new_n7741__), .dout(new_new_n7743__));
  buf1  g4929(.din(new_new_n7736__), .dout(new_new_n7744__));
  buf1  g4930(.din(new_new_n7744__), .dout(new_new_n7745__));
  buf1  g4931(.din(new_new_n7745__), .dout(new_new_n7746__));
  buf1  g4932(.din(new_new_n7745__), .dout(new_new_n7747__));
  buf1  g4933(.din(new_new_n7744__), .dout(new_new_n7748__));
  buf1  g4934(.din(new_new_n7748__), .dout(new_new_n7749__));
  buf1  g4935(.din(new_new_n4066__), .dout(new_new_n7750__));
  buf1  g4936(.din(new_new_n7750__), .dout(new_new_n7751__));
  buf1  g4937(.din(new_new_n7751__), .dout(new_new_n7752__));
  buf1  g4938(.din(new_new_n7752__), .dout(new_new_n7753__));
  buf1  g4939(.din(new_new_n7752__), .dout(new_new_n7754__));
  buf1  g4940(.din(new_new_n7751__), .dout(new_new_n7755__));
  buf1  g4941(.din(new_new_n7755__), .dout(new_new_n7756__));
  buf1  g4942(.din(new_new_n7755__), .dout(new_new_n7757__));
  buf1  g4943(.din(new_new_n7750__), .dout(new_new_n7758__));
  buf1  g4944(.din(new_new_n7758__), .dout(new_new_n7759__));
  buf1  g4945(.din(new_new_n7759__), .dout(new_new_n7760__));
  buf1  g4946(.din(new_new_n7759__), .dout(new_new_n7761__));
  buf1  g4947(.din(new_new_n7758__), .dout(new_new_n7762__));
  buf1  g4948(.din(new_new_n4060__), .dout(new_new_n7763__));
  buf1  g4949(.din(new_new_n7763__), .dout(new_new_n7764__));
  buf1  g4950(.din(new_new_n7764__), .dout(new_new_n7765__));
  buf1  g4951(.din(new_new_n7765__), .dout(new_new_n7766__));
  buf1  g4952(.din(new_new_n7765__), .dout(new_new_n7767__));
  buf1  g4953(.din(new_new_n7764__), .dout(new_new_n7768__));
  buf1  g4954(.din(new_new_n7768__), .dout(new_new_n7769__));
  buf1  g4955(.din(new_new_n7768__), .dout(new_new_n7770__));
  buf1  g4956(.din(new_new_n7763__), .dout(new_new_n7771__));
  buf1  g4957(.din(new_new_n7771__), .dout(new_new_n7772__));
  buf1  g4958(.din(new_new_n7772__), .dout(new_new_n7773__));
  buf1  g4959(.din(new_new_n7772__), .dout(new_new_n7774__));
  buf1  g4960(.din(new_new_n7771__), .dout(new_new_n7775__));
  buf1  g4961(.din(new_new_n7775__), .dout(new_new_n7776__));
  buf1  g4962(.din(new_new_n3665__), .dout(new_new_n7777__));
  buf1  g4963(.din(new_new_n3664__), .dout(new_new_n7778__));
  buf1  g4964(.din(new_new_n7778__), .dout(new_new_n7779__));
  buf1  g4965(.din(new_new_n3752__), .dout(new_new_n7780__));
  buf1  g4966(.din(new_new_n3958__), .dout(new_new_n7781__));
  buf1  g4967(.din(new_new_n3108__), .dout(new_new_n7782__));
  buf1  g4968(.din(new_new_n7782__), .dout(new_new_n7783__));
  buf1  g4969(.din(new_new_n3090__), .dout(new_new_n7784__));
  buf1  g4970(.din(new_new_n3130__), .dout(new_new_n7785__));
  buf1  g4971(.din(new_new_n3132__), .dout(new_new_n7786__));
  buf1  g4972(.din(new_new_n4050__), .dout(new_new_n7787__));
  buf1  g4973(.din(new_new_n7787__), .dout(new_new_n7788__));
  buf1  g4974(.din(new_new_n7787__), .dout(new_new_n7789__));
  buf1  g4975(.din(new_new_n4051__), .dout(new_new_n7790__));
  buf1  g4976(.din(new_new_n7790__), .dout(new_new_n7791__));
  buf1  g4977(.din(new_new_n7790__), .dout(new_new_n7792__));
  buf1  g4978(.din(new_new_n4022__), .dout(new_new_n7793__));
  buf1  g4979(.din(new_new_n4914__), .dout(new_new_n7794__));
  buf1  g4980(.din(new_new_n7794__), .dout(new_new_n7795__));
  buf1  g4981(.din(new_new_n5424__), .dout(new_new_n7796__));
  buf1  g4982(.din(new_new_n7796__), .dout(new_new_n7797__));
  buf1  g4983(.din(new_new_n4049__), .dout(new_new_n7798__));
  buf1  g4984(.din(new_new_n7798__), .dout(new_new_n7799__));
  buf1  g4985(.din(new_new_n7798__), .dout(new_new_n7800__));
  buf1  g4986(.din(new_new_n4879__), .dout(new_new_n7801__));
  buf1  g4987(.din(new_new_n4915__), .dout(new_new_n7802__));
  buf1  g4988(.din(new_new_n7802__), .dout(new_new_n7803__));
  buf1  g4989(.din(new_new_n7802__), .dout(new_new_n7804__));
  buf1  g4990(.din(new_new_n5427__), .dout(new_new_n7805__));
  buf1  g4991(.din(new_new_n3741__), .dout(new_new_n7806__));
  buf1  g4992(.din(new_new_n3740__), .dout(new_new_n7807__));
  buf1  g4993(.din(new_new_n7807__), .dout(new_new_n7808__));
  buf1  g4994(.din(new_new_n3911__), .dout(new_new_n7809__));
  buf1  g4995(.din(new_new_n7809__), .dout(new_new_n7810__));
  buf1  g4996(.din(new_new_n5433__), .dout(new_new_n7811__));
  buf1  g4997(.din(new_new_n3910__), .dout(new_new_n7812__));
  buf1  g4998(.din(new_new_n7812__), .dout(new_new_n7813__));
  buf1  g4999(.din(new_new_n7812__), .dout(new_new_n7814__));
  buf1  g5000(.din(new_new_n5434__), .dout(new_new_n7815__));
  buf1  g5001(.din(new_new_n3742__), .dout(new_new_n7816__));
  buf1  g5002(.din(new_new_n3954__), .dout(new_new_n7817__));
  buf1  g5003(.din(new_new_n4048__), .dout(new_new_n7818__));
  buf1  g5004(.din(new_new_n7818__), .dout(new_new_n7819__));
  buf1  g5005(.din(new_new_n7818__), .dout(new_new_n7820__));
  buf1  g5006(.din(new_new_n5423__), .dout(new_new_n7821__));
  buf1  g5007(.din(new_new_n7821__), .dout(new_new_n7822__));
  buf1  g5008(.din(new_new_n5444__), .dout(new_new_n7823__));
  buf1  g5009(.din(new_new_n7823__), .dout(new_new_n7824__));
  buf1  g5010(.din(new_new_n5443__), .dout(new_new_n7825__));
  buf1  g5011(.din(new_new_n7825__), .dout(new_new_n7826__));
  buf1  g5012(.din(new_new_n5453__), .dout(new_new_n7827__));
  buf1  g5013(.din(new_new_n4838__), .dout(new_new_n7828__));
  buf1  g5014(.din(new_new_n7828__), .dout(new_new_n7829__));
  buf1  g5015(.din(new_new_n5457__), .dout(new_new_n7830__));
  buf1  g5016(.din(new_new_n4837__), .dout(new_new_n7831__));
  buf1  g5017(.din(new_new_n5458__), .dout(new_new_n7832__));
  buf1  g5018(.din(new_new_n3745__), .dout(new_new_n7833__));
  buf1  g5019(.din(new_new_n3744__), .dout(new_new_n7834__));
  buf1  g5020(.din(new_new_n7834__), .dout(new_new_n7835__));
  buf1  g5021(.din(new_new_n7834__), .dout(new_new_n7836__));
  buf1  g5022(.din(new_new_n5464__), .dout(new_new_n7837__));
  buf1  g5023(.din(new_new_n5465__), .dout(new_new_n7838__));
  buf1  g5024(.din(new_new_n4843__), .dout(new_new_n7839__));
  buf1  g5025(.din(new_new_n3746__), .dout(new_new_n7840__));
  buf1  g5026(.din(new_new_n7840__), .dout(new_new_n7841__));
  buf1  g5027(.din(new_new_n5472__), .dout(new_new_n7842__));
  buf1  g5028(.din(new_new_n3747__), .dout(new_new_n7843__));
  buf1  g5029(.din(new_new_n5471__), .dout(new_new_n7844__));
  buf1  g5030(.din(new_new_n5468__), .dout(new_new_n7845__));
  buf1  g5031(.din(new_new_n5478__), .dout(new_new_n7846__));
  buf1  g5032(.din(new_new_n7846__), .dout(new_new_n7847__));
  buf1  g5033(.din(new_new_n5373__), .dout(new_new_n7848__));
  buf1  g5034(.din(new_new_n4995__), .dout(new_new_n7849__));
  buf1  g5035(.din(new_new_n4999__), .dout(new_new_n7850__));
  buf1  g5036(.din(new_new_n3656__), .dout(new_new_n7851__));
  buf1  g5037(.din(new_new_n3114__), .dout(new_new_n7852__));
  buf1  g5038(.din(new_new_n3643__), .dout(new_new_n7853__));
  buf1  g5039(.din(new_new_n3642__), .dout(new_new_n7854__));
  buf1  g5040(.din(new_new_n7854__), .dout(new_new_n7855__));
  buf1  g5041(.din(new_new_n3666__), .dout(new_new_n7856__));
  buf1  g5042(.din(new_new_n3641__), .dout(new_new_n7857__));
  buf1  g5043(.din(new_new_n3640__), .dout(new_new_n7858__));
  buf1  g5044(.din(new_new_n7858__), .dout(new_new_n7859__));
  buf1  g5045(.din(new_new_n3668__), .dout(new_new_n7860__));
  buf1  g5046(.din(new_new_n3639__), .dout(new_new_n7861__));
  buf1  g5047(.din(new_new_n3638__), .dout(new_new_n7862__));
  buf1  g5048(.din(new_new_n7862__), .dout(new_new_n7863__));
  buf1  g5049(.din(new_new_n3670__), .dout(new_new_n7864__));
  buf1  g5050(.din(new_new_n3653__), .dout(new_new_n7865__));
  buf1  g5051(.din(new_new_n3652__), .dout(new_new_n7866__));
  buf1  g5052(.din(new_new_n7866__), .dout(new_new_n7867__));
  buf1  g5053(.din(new_new_n3698__), .dout(new_new_n7868__));
  buf1  g5054(.din(new_new_n3663__), .dout(new_new_n7869__));
  buf1  g5055(.din(new_new_n3662__), .dout(new_new_n7870__));
  buf1  g5056(.din(new_new_n7870__), .dout(new_new_n7871__));
  buf1  g5057(.din(new_new_n3724__), .dout(new_new_n7872__));
  buf1  g5058(.din(new_new_n3661__), .dout(new_new_n7873__));
  buf1  g5059(.din(new_new_n3660__), .dout(new_new_n7874__));
  buf1  g5060(.din(new_new_n7874__), .dout(new_new_n7875__));
  buf1  g5061(.din(new_new_n3726__), .dout(new_new_n7876__));
  buf1  g5062(.din(new_new_n3749__), .dout(new_new_n7877__));
  buf1  g5063(.din(new_new_n3748__), .dout(new_new_n7878__));
  buf1  g5064(.din(new_new_n7878__), .dout(new_new_n7879__));
  buf1  g5065(.din(new_new_n4859__), .dout(new_new_n7880__));
  buf1  g5066(.din(new_new_n7880__), .dout(new_new_n7881__));
  buf1  g5067(.din(new_new_n4858__), .dout(new_new_n7882__));
  buf1  g5068(.din(new_new_n3908__), .dout(new_new_n7883__));
  buf1  g5069(.din(new_new_n5565__), .dout(new_new_n7884__));
  buf1  g5070(.din(new_new_n3909__), .dout(new_new_n7885__));
  buf1  g5071(.din(new_new_n5564__), .dout(new_new_n7886__));
  buf1  g5072(.din(new_new_n5559__), .dout(new_new_n7887__));
  buf1  g5073(.din(new_new_n5574__), .dout(new_new_n7888__));
  buf1  g5074(.din(new_new_n3066__), .dout(new_new_n7889__));
  buf1  g5075(.din(new_new_n4933__), .dout(new_new_n7890__));
  buf1  g5076(.din(new_new_n5584__), .dout(new_new_n7891__));
  buf1  g5077(.din(new_new_n5587__), .dout(new_new_n7892__));
  buf1  g5078(.din(new_new_n4925__), .dout(new_new_n7893__));
  buf1  g5079(.din(new_new_n7893__), .dout(new_new_n7894__));
  buf1  g5080(.din(new_new_n5000__), .dout(new_new_n7895__));
  buf1  g5081(.din(new_new_n5376__), .dout(new_new_n7896__));
  buf1  g5082(.din(new_new_n7896__), .dout(new_new_n7897__));
  buf1  g5083(.din(new_new_n5590__), .dout(new_new_n7898__));
  buf1  g5084(.din(new_new_n5385__), .dout(new_new_n7899__));
  buf1  g5085(.din(new_new_n7899__), .dout(new_new_n7900__));
  buf1  g5086(.din(new_new_n5400__), .dout(new_new_n7901__));
  buf1  g5087(.din(new_new_n7901__), .dout(new_new_n7902__));
  buf1  g5088(.din(new_new_n5394__), .dout(new_new_n7903__));
  buf1  g5089(.din(new_new_n7903__), .dout(new_new_n7904__));
  buf1  g5090(.din(new_new_n5403__), .dout(new_new_n7905__));
  buf1  g5091(.din(new_new_n7905__), .dout(new_new_n7906__));
  buf1  g5092(.din(new_new_n3926__), .dout(new_new_n7907__));
  buf1  g5093(.din(new_new_n7907__), .dout(new_new_n7908__));
  buf1  g5094(.din(new_new_n3927__), .dout(new_new_n7909__));
  buf1  g5095(.din(new_new_n4062__), .dout(new_new_n7910__));
  buf1  g5096(.din(new_new_n7910__), .dout(new_new_n7911__));
  buf1  g5097(.din(new_new_n7911__), .dout(new_new_n7912__));
  buf1  g5098(.din(new_new_n7910__), .dout(new_new_n7913__));
  buf1  g5099(.din(new_new_n4061__), .dout(new_new_n7914__));
  buf1  g5100(.din(new_new_n7914__), .dout(new_new_n7915__));
  buf1  g5101(.din(new_new_n7915__), .dout(new_new_n7916__));
  buf1  g5102(.din(new_new_n7914__), .dout(new_new_n7917__));
  buf1  g5103(.din(new_new_n3961__), .dout(new_new_n7918__));
  buf1  g5104(.din(new_new_n7918__), .dout(new_new_n7919__));
  buf1  g5105(.din(new_new_n7918__), .dout(new_new_n7920__));
  buf1  g5106(.din(new_new_n3960__), .dout(new_new_n7921__));
  buf1  g5107(.din(new_new_n7921__), .dout(new_new_n7922__));
  buf1  g5108(.din(new_new_n7922__), .dout(new_new_n7923__));
  buf1  g5109(.din(new_new_n7921__), .dout(new_new_n7924__));
  buf1  g5110(.din(new_new_n4064__), .dout(new_new_n7925__));
  buf1  g5111(.din(new_new_n7925__), .dout(new_new_n7926__));
  buf1  g5112(.din(new_new_n7925__), .dout(new_new_n7927__));
  buf1  g5113(.din(new_new_n4067__), .dout(new_new_n7928__));
  buf1  g5114(.din(new_new_n7928__), .dout(new_new_n7929__));
  buf1  g5115(.din(new_new_n7928__), .dout(new_new_n7930__));
  buf1  g5116(.din(new_new_n5397__), .dout(new_new_n7931__));
  buf1  g5117(.din(new_new_n7931__), .dout(new_new_n7932__));
  buf1  g5118(.din(new_new_n5622__), .dout(new_new_n7933__));
  buf1  g5119(.din(new_new_n3695__), .dout(new_new_n7934__));
  buf1  g5120(.din(new_new_n3694__), .dout(new_new_n7935__));
  buf1  g5121(.din(new_new_n7935__), .dout(new_new_n7936__));
  buf1  g5122(.din(new_new_n3756__), .dout(new_new_n7937__));
  buf1  g5123(.din(new_new_n3720__), .dout(new_new_n7938__));
  buf1  g5124(.din(new_new_n7938__), .dout(new_new_n7939__));
  buf1  g5125(.din(new_new_n3721__), .dout(new_new_n7940__));
  buf1  g5126(.din(new_new_n3928__), .dout(new_new_n7941__));
  buf1  g5127(.din(new_new_n5633__), .dout(new_new_n7942__));
  buf1  g5128(.din(new_new_n5642__), .dout(new_new_n7943__));
  buf1  g5129(.din(new_new_n3956__), .dout(new_new_n7944__));
  buf1  g5130(.din(new_new_n4945__), .dout(new_new_n7945__));
  buf1  g5131(.din(new_new_n4968__), .dout(new_new_n7946__));
  buf1  g5132(.din(new_new_n4828__), .dout(new_new_n7947__));
  buf1  g5133(.din(new_new_n7947__), .dout(new_new_n7948__));
  buf1  g5134(.din(new_new_n4835__), .dout(new_new_n7949__));
  buf1  g5135(.din(new_new_n4827__), .dout(new_new_n7950__));
  buf1  g5136(.din(new_new_n4836__), .dout(new_new_n7951__));
  buf1  g5137(.din(new_new_n7951__), .dout(new_new_n7952__));
  buf1  g5138(.din(new_new_n3719__), .dout(new_new_n7953__));
  buf1  g5139(.din(new_new_n7953__), .dout(new_new_n7954__));
  buf1  g5140(.din(new_new_n7953__), .dout(new_new_n7955__));
  buf1  g5141(.din(new_new_n3718__), .dout(new_new_n7956__));
  buf1  g5142(.din(new_new_n7956__), .dout(new_new_n7957__));
  buf1  g5143(.din(new_new_n7957__), .dout(new_new_n7958__));
  buf1  g5144(.din(new_new_n7956__), .dout(new_new_n7959__));
  buf1  g5145(.din(new_new_n3924__), .dout(new_new_n7960__));
  buf1  g5146(.din(new_new_n7960__), .dout(new_new_n7961__));
  buf1  g5147(.din(new_new_n3925__), .dout(new_new_n7962__));
  buf1  g5148(.din(new_new_n3283__), .dout(new_new_n7963__));
  buf1  g5149(.din(new_new_n3282__), .dout(new_new_n7964__));
  buf1  g5150(.din(new_new_n4863__), .dout(new_new_n7965__));
  buf1  g5151(.din(new_new_n4974__), .dout(new_new_n7966__));
  buf1  g5152(.din(new_new_n3190__), .dout(new_new_n7967__));
  buf1  g5153(.din(new_new_n5415__), .dout(new_new_n7968__));
  buf1  g5154(.din(new_new_n3192__), .dout(new_new_n7969__));
  buf1  g5155(.din(new_new_n4990__), .dout(new_new_n7970__));
  buf1  g5156(.din(new_new_n5416__), .dout(new_new_n7971__));
  buf1  g5157(.din(new_new_n3118__), .dout(new_new_n7972__));
  buf1  g5158(.din(new_new_n3122__), .dout(new_new_n7973__));
  buf1  g5159(.din(new_new_n5591__), .dout(new_new_n7974__));
  buf1  g5160(.din(new_new_n7974__), .dout(new_new_n7975__));
  buf1  g5161(.din(new_new_n5420__), .dout(new_new_n7976__));
  buf1  g5162(.din(new_new_n7976__), .dout(new_new_n7977__));
  buf1  g5163(.din(new_new_n7976__), .dout(new_new_n7978__));
  buf1  g5164(.din(new_new_n5456__), .dout(new_new_n7979__));
  buf1  g5165(.din(new_new_n7979__), .dout(new_new_n7980__));
  buf1  g5166(.din(new_new_n5481__), .dout(new_new_n7981__));
  buf1  g5167(.din(new_new_n5375__), .dout(new_new_n7982__));
  buf1  g5168(.din(new_new_n5418__), .dout(new_new_n7983__));
  buf1  g5169(.din(new_new_n4991__), .dout(new_new_n7984__));
  buf1  g5170(.din(new_new_n4993__), .dout(new_new_n7985__));
  buf1  g5171(.din(new_new_n5483__), .dout(new_new_n7986__));
  buf1  g5172(.din(new_new_n3180__), .dout(new_new_n7987__));
  buf1  g5173(.din(new_new_n7987__), .dout(new_new_n7988__));
  buf1  g5174(.din(new_new_n5579__), .dout(new_new_n7989__));
  buf1  g5175(.din(new_new_n7989__), .dout(new_new_n7990__));
  buf1  g5176(.din(new_new_n5582__), .dout(new_new_n7991__));
  buf1  g5177(.din(new_new_n5718__), .dout(new_new_n7992__));
  buf1  g5178(.din(new_new_n3188__), .dout(new_new_n7993__));
  buf1  g5179(.din(new_new_n5117__), .dout(new_new_n7994__));
  buf1  g5180(.din(new_new_n5583__), .dout(new_new_n7995__));
  buf1  g5181(.din(new_new_n3172__), .dout(new_new_n7996__));
  buf1  g5182(.din(new_new_n5409__), .dout(new_new_n7997__));
  buf1  g5183(.din(new_new_n5714__), .dout(new_new_n7998__));
  buf1  g5184(.din(new_new_n5715__), .dout(new_new_n7999__));
  buf1  g5185(.din(new_new_n5716__), .dout(new_new_n8000__));
  buf1  g5186(.din(new_new_n2224__), .dout(new_new_n8001__));
  buf1  g5187(.din(new_new_n2288__), .dout(new_new_n8002__));
  buf1  g5188(.din(new_new_n8002__), .dout(new_new_n8003__));
  buf1  g5189(.din(new_new_n8002__), .dout(new_new_n8004__));
  buf1  g5190(.din(new_new_n2289__), .dout(new_new_n8005__));
  buf1  g5191(.din(new_new_n8005__), .dout(new_new_n8006__));
  buf1  g5192(.din(new_new_n2228__), .dout(new_new_n8007__));
  buf1  g5193(.din(new_new_n2254__), .dout(new_new_n8008__));
  buf1  g5194(.din(new_new_n3201__), .dout(new_new_n8009__));
  buf1  g5195(.din(new_new_n8009__), .dout(new_new_n8010__));
  buf1  g5196(.din(new_new_n3208__), .dout(new_new_n8011__));
  buf1  g5197(.din(new_new_n2405__), .dout(new_new_n8012__));
  buf1  g5198(.din(new_new_n8012__), .dout(new_new_n8013__));
  buf1  g5199(.din(new_new_n8012__), .dout(new_new_n8014__));
  buf1  g5200(.din(new_new_n3117__), .dout(new_new_n8015__));
  buf1  g5201(.din(new_new_n4153__), .dout(new_new_n8016__));
  buf1  g5202(.din(new_new_n4191__), .dout(new_new_n8017__));
  buf1  g5203(.din(new_new_n4195__), .dout(new_new_n8018__));
  buf1  g5204(.din(new_new_n4223__), .dout(new_new_n8019__));
  buf1  g5205(.din(new_new_n4224__), .dout(new_new_n8020__));
  always @ (posedge clock) begin
    n2610_lo <= n11762;
    n2613_lo <= n11765;
    n2616_lo <= n11768;
    n2619_lo <= n11771;
    n2622_lo <= n11774;
    n2625_lo <= n11777;
    n2628_lo <= n11780;
    n2634_lo <= n11783;
    n2637_lo <= n11786;
    n2640_lo <= n11789;
    n2643_lo <= n11792;
    n2646_lo <= n11795;
    n2649_lo <= n11798;
    n2652_lo <= n11801;
    n2655_lo <= n11804;
    n2658_lo <= n11807;
    n2661_lo <= n11810;
    n2664_lo <= n11813;
    n2667_lo <= n11816;
    n2670_lo <= n11819;
    n2673_lo <= n11822;
    n2676_lo <= n11825;
    n2679_lo <= n11828;
    n2682_lo <= n11831;
    n2685_lo <= n11834;
    n2688_lo <= n11837;
    n2691_lo <= n11840;
    n2694_lo <= n11843;
    n2697_lo <= n11846;
    n2700_lo <= n11849;
    n2703_lo <= n11852;
    n2706_lo <= n11855;
    n2709_lo <= n11858;
    n2712_lo <= n11861;
    n2715_lo <= n11864;
    n2718_lo <= n11867;
    n2721_lo <= n11870;
    n2724_lo <= n11873;
    n2727_lo <= n11876;
    n2730_lo <= n11879;
    n2733_lo <= n11882;
    n2736_lo <= n11885;
    n2739_lo <= n11888;
    n2742_lo <= n11891;
    n2745_lo <= n11894;
    n2748_lo <= n11897;
    n2751_lo <= n11900;
    n2754_lo <= n11903;
    n2757_lo <= n11906;
    n2760_lo <= n11909;
    n2763_lo <= n11912;
    n2766_lo <= n11915;
    n2769_lo <= n11918;
    n2772_lo <= n11921;
    n2775_lo <= n11924;
    n2778_lo <= n11927;
    n2781_lo <= n11930;
    n2784_lo <= n11933;
    n2787_lo <= n11936;
    n2790_lo <= n11939;
    n2793_lo <= n11942;
    n2796_lo <= n11945;
    n2799_lo <= n11948;
    n2802_lo <= n11951;
    n2805_lo <= n11954;
    n2808_lo <= n11957;
    n2811_lo <= n11960;
    n2814_lo <= n11963;
    n2817_lo <= n11966;
    n2820_lo <= n11969;
    n2823_lo <= n11972;
    n2826_lo <= n11975;
    n2829_lo <= n11978;
    n2832_lo <= n11981;
    n2838_lo <= n11984;
    n2841_lo <= n11987;
    n2844_lo <= n11990;
    n2847_lo <= n11993;
    n2850_lo <= n11996;
    n2853_lo <= n11999;
    n2856_lo <= n12002;
    n2862_lo <= n12005;
    n2865_lo <= n12008;
    n2868_lo <= n12011;
    n2871_lo <= n12014;
    n2874_lo <= n12017;
    n2877_lo <= n12020;
    n2880_lo <= n12023;
    n2883_lo <= n12026;
    n2886_lo <= n12029;
    n2889_lo <= n12032;
    n2892_lo <= n12035;
    n2895_lo <= n12038;
    n2898_lo <= n12041;
    n2901_lo <= n12044;
    n2904_lo <= n12047;
    n2907_lo <= n12050;
    n2910_lo <= n12053;
    n2913_lo <= n12056;
    n2916_lo <= n12059;
    n2919_lo <= n12062;
    n2922_lo <= n12065;
    n2925_lo <= n12068;
    n2928_lo <= n12071;
    n2931_lo <= n12074;
    n2934_lo <= n12077;
    n2937_lo <= n12080;
    n2940_lo <= n12083;
    n2943_lo <= n12086;
    n2946_lo <= n12089;
    n2949_lo <= n12092;
    n2952_lo <= n12095;
    n2955_lo <= n12098;
    n2958_lo <= n12101;
    n2961_lo <= n12104;
    n2964_lo <= n12107;
    n2967_lo <= n12110;
    n2970_lo <= n12113;
    n2973_lo <= n12116;
    n2976_lo <= n12119;
    n2979_lo <= n12122;
    n2982_lo <= n12125;
    n2985_lo <= n12128;
    n2988_lo <= n12131;
    n2991_lo <= n12134;
    n2994_lo <= n12137;
    n2997_lo <= n12140;
    n3000_lo <= n12143;
    n3003_lo <= n12146;
    n3006_lo <= n12149;
    n3009_lo <= n12152;
    n3012_lo <= n12155;
    n3015_lo <= n12158;
    n3018_lo <= n12161;
    n3021_lo <= n12164;
    n3024_lo <= n12167;
    n3027_lo <= n12170;
    n3030_lo <= n12173;
    n3033_lo <= n12176;
    n3036_lo <= n12179;
    n3039_lo <= n12182;
    n3042_lo <= n12185;
    n3045_lo <= n12188;
    n3048_lo <= n12191;
    n3051_lo <= n12194;
    n3054_lo <= n12197;
    n3057_lo <= n12200;
    n3060_lo <= n12203;
    n3063_lo <= n12206;
    n3066_lo <= n12209;
    n3069_lo <= n12212;
    n3072_lo <= n12215;
    n3075_lo <= n12218;
    n3078_lo <= n12221;
    n3081_lo <= n12224;
    n3084_lo <= n12227;
    n3087_lo <= n12230;
    n3090_lo <= n12233;
    n3093_lo <= n12236;
    n3096_lo <= n12239;
    n3099_lo <= n12242;
    n3102_lo <= n12245;
    n3105_lo <= n12248;
    n3108_lo <= n12251;
    n3111_lo <= n12254;
    n3114_lo <= n12257;
    n3117_lo <= n12260;
    n3120_lo <= n12263;
    n3126_lo <= n12266;
    n3129_lo <= n12269;
    n3132_lo <= n12272;
    n3138_lo <= n12275;
    n3141_lo <= n12278;
    n3144_lo <= n12281;
    n3147_lo <= n12284;
    n3150_lo <= n12287;
    n3153_lo <= n12290;
    n3156_lo <= n12293;
    n3162_lo <= n12296;
    n3165_lo <= n12299;
    n3168_lo <= n12302;
    n3174_lo <= n12305;
    n3177_lo <= n12308;
    n3180_lo <= n12311;
    n3186_lo <= n12314;
    n3189_lo <= n12317;
    n3192_lo <= n12320;
    n3195_lo <= n12323;
    n3198_lo <= n12326;
    n3201_lo <= n12329;
    n3204_lo <= n12332;
    n3210_lo <= n12335;
    n3213_lo <= n12338;
    n3216_lo <= n12341;
    n3219_lo <= n12344;
    n3222_lo <= n12347;
    n3225_lo <= n12350;
    n3228_lo <= n12353;
    n3234_lo <= n12356;
    n3237_lo <= n12359;
    n3240_lo <= n12362;
    n3243_lo <= n12365;
    n3246_lo <= n12368;
    n3249_lo <= n12371;
    n3252_lo <= n12374;
    n3255_lo <= n12377;
    n3258_lo <= n12380;
    n3261_lo <= n12383;
    n3264_lo <= n12386;
    n3267_lo <= n12389;
    n3270_lo <= n12392;
    n3273_lo <= n12395;
    n3276_lo <= n12398;
    n3279_lo <= n12401;
    n3282_lo <= n12404;
    n3285_lo <= n12407;
    n3288_lo <= n12410;
    n3294_lo <= n12413;
    n3297_lo <= n12416;
    n3300_lo <= n12419;
    n3306_lo <= n12422;
    n3309_lo <= n12425;
    n3312_lo <= n12428;
    n3318_lo <= n12431;
    n3321_lo <= n12434;
    n3324_lo <= n12437;
    n3330_lo <= n12440;
    n3333_lo <= n12443;
    n3336_lo <= n12446;
    n3339_lo <= n12449;
    n3342_lo <= n12452;
    n3345_lo <= n12455;
    n3348_lo <= n12458;
    n3351_lo <= n12461;
    n3354_lo <= n12464;
    n3357_lo <= n12467;
    n3360_lo <= n12470;
    n3363_lo <= n12473;
    n3366_lo <= n12476;
    n3369_lo <= n12479;
    n3372_lo <= n12482;
    n3375_lo <= n12485;
    n3378_lo <= n12488;
    n3381_lo <= n12491;
    n3384_lo <= n12494;
    n3387_lo <= n12497;
    n3390_lo <= n12500;
    n3393_lo <= n12503;
    n3396_lo <= n12506;
    n3399_lo <= n12509;
    n3402_lo <= n12512;
    n3405_lo <= n12515;
    n3408_lo <= n12518;
    n3411_lo <= n12521;
    n3414_lo <= n12524;
    n3417_lo <= n12527;
    n3420_lo <= n12530;
    n3423_lo <= n12533;
    n3426_lo <= n12536;
    n3429_lo <= n12539;
    n3432_lo <= n12542;
    n3435_lo <= n12545;
    n3438_lo <= n12548;
    n3441_lo <= n12551;
    n3444_lo <= n12554;
    n3447_lo <= n12557;
    n3450_lo <= n12560;
    n3453_lo <= n12563;
    n3456_lo <= n12566;
    n3459_lo <= n12569;
    n3462_lo <= n12572;
    n3465_lo <= n12575;
    n3468_lo <= n12578;
    n3471_lo <= n12581;
    n3474_lo <= n12584;
    n3477_lo <= n12587;
    n3480_lo <= n12590;
    n3483_lo <= n12593;
    n3486_lo <= n12596;
    n3489_lo <= n12599;
    n3492_lo <= n12602;
    n3495_lo <= n12605;
    n3498_lo <= n12608;
    n3501_lo <= n12611;
    n3504_lo <= n12614;
    n3507_lo <= n12617;
    n3510_lo <= n12620;
    n3513_lo <= n12623;
    n3516_lo <= n12626;
    n3519_lo <= n12629;
    n3522_lo <= n12632;
    n3525_lo <= n12635;
    n3528_lo <= n12638;
    n3531_lo <= n12641;
    n3534_lo <= n12644;
    n3537_lo <= n12647;
    n3540_lo <= n12650;
    n3543_lo <= n12653;
    n3546_lo <= n12656;
    n3549_lo <= n12659;
    n3552_lo <= n12662;
    n3555_lo <= n12665;
    n3558_lo <= n12668;
    n3561_lo <= n12671;
    n3564_lo <= n12674;
    n3567_lo <= n12677;
    n3570_lo <= n12680;
    n3573_lo <= n12683;
    n3576_lo <= n12686;
    n3579_lo <= n12689;
    n3582_lo <= n12692;
    n3585_lo <= n12695;
    n3588_lo <= n12698;
    n3591_lo <= n12701;
    n3594_lo <= n12704;
    n3597_lo <= n12707;
    n3600_lo <= n12710;
    n3603_lo <= n12713;
    n3606_lo <= n12716;
    n3609_lo <= n12719;
    n3612_lo <= n12722;
    n3615_lo <= n12725;
    n3618_lo <= n12728;
    n3621_lo <= n12731;
    n3624_lo <= n12734;
    n3627_lo <= n12737;
    n3630_lo <= n12740;
    n3633_lo <= n12743;
    n3636_lo <= n12746;
    n3639_lo <= n12749;
    n3642_lo <= n12752;
    n3645_lo <= n12755;
    n3648_lo <= n12758;
    n3651_lo <= n12761;
    n3654_lo <= n12764;
    n3666_lo <= n12767;
    n3750_lo <= n12770;
    n3762_lo <= n12773;
    n3774_lo <= n12776;
    n3786_lo <= n12779;
    n3789_lo <= n12782;
    n3792_lo <= n12785;
    n3795_lo <= n12788;
    n3798_lo <= n12791;
    n3810_lo <= n12794;
    n3822_lo <= n12797;
    n3834_lo <= n12800;
    n3846_lo <= n12803;
    n3930_lo <= n12806;
    n3933_lo <= n12809;
    n3936_lo <= n12812;
    n3942_lo <= n12815;
    n3945_lo <= n12818;
    n3948_lo <= n12821;
    n3954_lo <= n12824;
    n3957_lo <= n12827;
    n3963_lo <= n12830;
    n3966_lo <= n12833;
    n3969_lo <= n12836;
    n3975_lo <= n12839;
    n3978_lo <= n12842;
    n3990_lo <= n12845;
    n4050_lo <= n12848;
    n4062_lo <= n12851;
    n4098_lo <= n12854;
    n4107_lo <= n12857;
    n4110_lo <= n12860;
    n4122_lo <= n12863;
    n4131_lo <= n12866;
    n4155_lo <= n12869;
    n4158_lo <= n12872;
    n4170_lo <= n12875;
    n4179_lo <= n12878;
    n4182_lo <= n12881;
    n4185_lo <= n12884;
    n4188_lo <= n12887;
    n4194_lo <= n12890;
    n4197_lo <= n12893;
    n4200_lo <= n12896;
    n4206_lo <= n12899;
    n4209_lo <= n12902;
    n4212_lo <= n12905;
    n4215_lo <= n12908;
    n4230_lo <= n12911;
    n4233_lo <= n12914;
    n4236_lo <= n12917;
    n4239_lo <= n12920;
    n4242_lo <= n12923;
    n4254_lo <= n12926;
    n4290_lo <= n12929;
    n4293_lo <= n12932;
    n4302_lo <= n12935;
    n4314_lo <= n12938;
    n4350_lo <= n12941;
    n4362_lo <= n12944;
    n4374_lo <= n12947;
    n4386_lo <= n12950;
    n4398_lo <= n12953;
    n4410_lo <= n12956;
    n4413_lo <= n12959;
    n4416_lo <= n12962;
    n4419_lo <= n12965;
    n4422_lo <= n12968;
    n4425_lo <= n12971;
    n4428_lo <= n12974;
    n4431_lo <= n12977;
    n4434_lo <= n12980;
    n4437_lo <= n12983;
    n4440_lo <= n12986;
    n4443_lo <= n12989;
    n4446_lo <= n12992;
    n4449_lo <= n12995;
    n4452_lo <= n12998;
    n4455_lo <= n13001;
    n4458_lo <= n13004;
    n4461_lo <= n13007;
    n4464_lo <= n13010;
    n4467_lo <= n13013;
    n4470_lo <= n13016;
    n4473_lo <= n13019;
    n4476_lo <= n13022;
    n4479_lo <= n13025;
    n4482_lo <= n13028;
    n4485_lo <= n13031;
    n4488_lo <= n13034;
    n4494_lo <= n13037;
    n4497_lo <= n13040;
    n4500_lo <= n13043;
    n4503_lo <= n13046;
    n4506_lo <= n13049;
    n4509_lo <= n13052;
    n4512_lo <= n13055;
    n4515_lo <= n13058;
    n4518_lo <= n13061;
    n4521_lo <= n13064;
    n4524_lo <= n13067;
    n4527_lo <= n13070;
    n4530_lo <= n13073;
    n4533_lo <= n13076;
    n4536_lo <= n13079;
    n4539_lo <= n13082;
    n4542_lo <= n13085;
    n4545_lo <= n13088;
    n4554_lo <= n13091;
    n4557_lo <= n13094;
    n4560_lo <= n13097;
    n4563_lo <= n13100;
    n4566_lo <= n13103;
    n4569_lo <= n13106;
    n4572_lo <= n13109;
    n4575_lo <= n13112;
    n4578_lo <= n13115;
    n4581_lo <= n13118;
    n4584_lo <= n13121;
    n4587_lo <= n13124;
    n4590_lo <= n13127;
    n4593_lo <= n13130;
    n4596_lo <= n13133;
    n4602_lo <= n13136;
    n4605_lo <= n13139;
    n4608_lo <= n13142;
    n4614_lo <= n13145;
    n4617_lo <= n13148;
    n4620_lo <= n13151;
    n4626_lo <= n13154;
    n4629_lo <= n13157;
    n4632_lo <= n13160;
    n4638_lo <= n13163;
    n4641_lo <= n13166;
    n4644_lo <= n13169;
    n4647_lo <= n13172;
    n4650_lo <= n13175;
    n4653_lo <= n13178;
    n4656_lo <= n13181;
    n4659_lo <= n13184;
    n4662_lo <= n13187;
    n4665_lo <= n13190;
    n4668_lo <= n13193;
    n4671_lo <= n13196;
    n4674_lo <= n13199;
    n4677_lo <= n13202;
    n4680_lo <= n13205;
    n4683_lo <= n13208;
    n4686_lo <= n13211;
    n4689_lo <= n13214;
    n4692_lo <= n13217;
    n4695_lo <= n13220;
    n4698_lo <= n13223;
    n4701_lo <= n13226;
    n4704_lo <= n13229;
    n4707_lo <= n13232;
    n4710_lo <= n13235;
    n4713_lo <= n13238;
    n4716_lo <= n13241;
    n4719_lo <= n13244;
    n4722_lo <= n13247;
    n4725_lo <= n13250;
    n4728_lo <= n13253;
    n4731_lo <= n13256;
    n4734_lo <= n13259;
    n4737_lo <= n13262;
    n4740_lo <= n13265;
    n4743_lo <= n13268;
    n4970_o2 <= n13271;
    n4972_o2 <= n13274;
    n4989_o2 <= n13277;
    n5024_o2 <= n13280;
    n5025_o2 <= n13283;
    n5029_o2 <= n13286;
    n5042_o2 <= n13289;
    n5048_o2 <= n13292;
    n5093_o2 <= n13295;
    n5096_o2 <= n13298;
    n5193_o2 <= n13301;
    n5199_o2 <= n13304;
    n5203_o2 <= n13307;
    n5214_o2 <= n13310;
    n5221_o2 <= n13313;
    n5222_o2 <= n13316;
    n5273_o2 <= n13319;
    n5365_o2 <= n13322;
    n5385_o2 <= n13325;
    n5553_o2 <= n13328;
    n5636_o2 <= n13331;
    n5782_o2 <= n13334;
    n5778_o2 <= n13337;
    n5323_o2 <= n13340;
    n5325_o2 <= n13343;
    n5327_o2 <= n13346;
    n5329_o2 <= n13349;
    n5816_o2 <= n13352;
    n5817_o2 <= n13355;
    n5837_o2 <= n13358;
    n5844_o2 <= n13361;
    n5859_o2 <= n13364;
    n5857_o2 <= n13367;
    n5369_o2 <= n13370;
    n5371_o2 <= n13373;
    n5373_o2 <= n13376;
    n5400_o2 <= n13379;
    n5402_o2 <= n13382;
    n5404_o2 <= n13385;
    n5406_o2 <= n13388;
    n5407_o2 <= n13391;
    n5408_o2 <= n13394;
    n2722_o2 <= n13397;
    n1942_inv <= n13400;
    n5412_o2 <= n13403;
    n1948_inv <= n13406;
    n5557_o2 <= n13409;
    n5558_o2 <= n13412;
    n5559_o2 <= n13415;
    n5564_o2 <= n13418;
    n5565_o2 <= n13421;
    n1966_inv <= n13424;
    n5568_o2 <= n13427;
    n5598_o2 <= n13430;
    n5600_o2 <= n13433;
    n5601_o2 <= n13436;
    n5602_o2 <= n13439;
    n5603_o2 <= n13442;
    n2853_o2 <= n13445;
    n5637_o2 <= n13448;
    n1993_inv <= n13451;
    n1996_inv <= n13454;
    n5635_o2 <= n13457;
    n5640_o2 <= n13460;
    n5641_o2 <= n13463;
    n5642_o2 <= n13466;
    n5650_o2 <= n13469;
    n5652_o2 <= n13472;
    n5653_o2 <= n13475;
    n5654_o2 <= n13478;
    n5655_o2 <= n13481;
    n5657_o2 <= n13484;
    n2029_inv <= n13487;
    n5661_o2 <= n13490;
    n5656_o2 <= n13493;
    n5663_o2 <= n13496;
    n2041_inv <= n13499;
    n5795_o2 <= n13502;
    n5796_o2 <= n13505;
    n5797_o2 <= n13508;
    n5739_o2 <= n13511;
    n5773_o2 <= n13514;
    n2059_inv <= n13517;
    n5799_o2 <= n13520;
    n5802_o2 <= n13523;
    n2068_inv <= n13526;
    n5831_o2 <= n13529;
    n5833_o2 <= n13532;
    n5820_o2 <= n13535;
    n5823_o2 <= n13538;
    n5824_o2 <= n13541;
    n5869_o2 <= n13544;
    n5848_o2 <= n13547;
    n5849_o2 <= n13550;
    n5856_o2 <= n13553;
    n5896_o2 <= n13556;
    n2754_o2 <= n13559;
    n2908_o2 <= n13562;
    n5892_o2 <= n13565;
    n5915_o2 <= n13568;
    n5919_o2 <= n13571;
    n5918_o2 <= n13574;
    n5920_o2 <= n13577;
    n5917_o2 <= n13580;
    lo586_buf_o2 <= n13583;
    n2818_o2 <= n13586;
    n2863_o2 <= n13589;
    n2134_inv <= n13592;
    n2725_o2 <= n13595;
    n3016_o2 <= n13598;
    n3013_o2 <= n13601;
    n2655_o2 <= n13604;
    n2149_inv <= n13607;
    lo562_buf_o2 <= n13610;
    n2155_inv <= n13613;
    n2531_o2 <= n13616;
    n2700_o2 <= n13619;
    n5908_o2 <= n13622;
    n5910_o2 <= n13625;
    n5912_o2 <= n13628;
    n5914_o2 <= n13631;
    n2753_o2 <= n13634;
    n2878_o2 <= n13637;
    n2182_inv <= n13640;
    n5934_o2 <= n13643;
    n5936_o2 <= n13646;
    n5938_o2 <= n13649;
    n2728_o2 <= n13652;
    lo358_buf_o2 <= n13655;
    lo418_buf_o2 <= n13658;
    lo474_buf_o2 <= n13661;
    lo554_buf_o2 <= n13664;
    lo558_buf_o2 <= n13667;
    lo574_buf_o2 <= n13670;
    n2215_inv <= n13673;
    n2218_inv <= n13676;
    n2221_inv <= n13679;
    lo450_buf_o2 <= n13682;
    n2910_o2 <= n13685;
    n2683_o2 <= n13688;
    n2828_o2 <= n13691;
    n2582_o2 <= n13694;
    n2600_o2 <= n13697;
    n2542_o2 <= n13700;
    n2703_o2 <= n13703;
    lo510_buf_o2 <= n13706;
    lo514_buf_o2 <= n13709;
    lo538_buf_o2 <= n13712;
    lo578_buf_o2 <= n13715;
    n2260_inv <= n13718;
    n2666_o2 <= n13721;
    n2667_o2 <= n13724;
    n2660_o2 <= n13727;
    n2272_inv <= n13730;
    lo454_buf_o2 <= n13733;
    n3593_o2 <= n13736;
    n3048_o2 <= n13739;
    lo410_buf_o2 <= n13742;
    lo502_buf_o2 <= n13745;
    lo506_buf_o2 <= n13748;
    lo550_buf_o2 <= n13751;
    lo570_buf_o2 <= n13754;
    lo582_buf_o2 <= n13757;
    n2302_inv <= n13760;
    n2305_inv <= n13763;
    n3499_o2 <= n13766;
    n2311_inv <= n13769;
    n2870_o2 <= n13772;
    n2317_inv <= n13775;
    n2689_o2 <= n13778;
    n2323_inv <= n13781;
    n2662_o2 <= n13784;
    lo350_buf_o2 <= n13787;
    lo498_buf_o2 <= n13790;
    lo518_buf_o2 <= n13793;
    lo522_buf_o2 <= n13796;
    lo598_buf_o2 <= n13799;
    n2344_inv <= n13802;
    n2347_inv <= n13805;
    n2350_inv <= n13808;
    n2353_inv <= n13811;
    n2356_inv <= n13814;
    n2359_inv <= n13817;
    n2872_o2 <= n13820;
    n3313_o2 <= n13823;
    n3273_o2 <= n13826;
    n2848_o2 <= n13829;
    n2893_o2 <= n13832;
    n3267_o2 <= n13835;
    n2925_o2 <= n13838;
    n2839_o2 <= n13841;
    n2831_o2 <= n13844;
    n2558_o2 <= n13847;
    n2562_o2 <= n13850;
    n2825_o2 <= n13853;
    n3263_o2 <= n13856;
    n3517_o2 <= n13859;
    n2873_o2 <= n13862;
    n2926_o2 <= n13865;
    n3261_o2 <= n13868;
    n3268_o2 <= n13871;
    n3274_o2 <= n13874;
    n3314_o2 <= n13877;
    n3571_o2 <= n13880;
    n2950_o2 <= n13883;
    n2951_o2 <= n13886;
    n3022_o2 <= n13889;
    n3023_o2 <= n13892;
    n3057_o2 <= n13895;
    n3058_o2 <= n13898;
    n2931_o2 <= n13901;
    n2911_o2 <= n13904;
    n2959_o2 <= n13907;
    n2960_o2 <= n13910;
    n2922_o2 <= n13913;
    n2888_o2 <= n13916;
    n2889_o2 <= n13919;
    n3051_o2 <= n13922;
    n3052_o2 <= n13925;
    n3063_o2 <= n13928;
    n2845_o2 <= n13931;
    n2476_inv <= n13934;
    n3281_o2 <= n13937;
    n3294_o2 <= n13940;
    n2885_o2 <= n13943;
    n2786_o2 <= n13946;
    n2783_o2 <= n13949;
    n2801_o2 <= n13952;
    n2572_o2 <= n13955;
    n2628_o2 <= n13958;
    n2609_o2 <= n13961;
    n2618_o2 <= n13964;
    n2637_o2 <= n13967;
    n2525_o2 <= n13970;
    n2551_o2 <= n13973;
    n3759_o2 <= n13976;
    n2994_o2 <= n13979;
    n3040_o2 <= n13982;
    n2943_o2 <= n13985;
    n2991_o2 <= n13988;
    n3034_o2 <= n13991;
    n2881_o2 <= n13994;
    n3021_o2 <= n13997;
    n3062_o2 <= n14000;
    n2763_o2 <= n14003;
    n2764_o2 <= n14006;
    n2775_o2 <= n14009;
    n2776_o2 <= n14012;
    n2968_o2 <= n14015;
    n2969_o2 <= n14018;
    n2798_o2 <= n14021;
    n3661_o2 <= n14024;
    n2694_o2 <= n14027;
    n2572_inv <= n14030;
    n2817_o2 <= n14033;
    n2514_o2 <= n14036;
    n2501_o2 <= n14039;
    n2584_inv <= n14042;
    n2505_o2 <= n14045;
    n2492_o2 <= n14048;
    lo546_buf_o2 <= n14051;
    lo590_buf_o2 <= n14054;
    lo594_buf_o2 <= n14057;
    n2602_inv <= n14060;
    n2605_inv <= n14063;
    n2709_o2 <= n14066;
    n2611_inv <= n14069;
    n2614_inv <= n14072;
    n2617_inv <= n14075;
    n2620_inv <= n14078;
    n3590_o2 <= n14081;
    n3591_o2 <= n14084;
    n2629_inv <= n14087;
    n3638_o2 <= n14090;
    n3639_o2 <= n14093;
    n2638_inv <= n14096;
    n2641_inv <= n14099;
    lo458_buf_o2 <= n14102;
    lo482_buf_o2 <= n14105;
    lo566_buf_o2 <= n14108;
    n2718_o2 <= n14111;
    n3707_o2 <= n14114;
    n3671_o2 <= n14117;
    n3680_o2 <= n14120;
    n3749_o2 <= n14123;
    n3716_o2 <= n14126;
    n3692_o2 <= n14129;
    n2591_o2 <= n14132;
    n3478_o2 <= n14135;
    n3610_o2 <= n14138;
    n3611_o2 <= n14141;
    n2686_inv <= n14144;
    n2689_inv <= n14147;
    n2738_o2 <= n14150;
    n3616_o2 <= n14153;
    n3617_o2 <= n14156;
    n3031_o2 <= n14159;
    n2704_inv <= n14162;
    n3562_o2 <= n14165;
    n2502_o2 <= n14168;
    n3560_o2 <= n14171;
    n3554_o2 <= n14174;
    n3555_o2 <= n14177;
    n3536_o2 <= n14180;
    n3537_o2 <= n14183;
    n3508_o2 <= n14186;
    n3650_o2 <= n14189;
    n3740_o2 <= n14192;
    n3484_o2 <= n14195;
    n2740_inv <= n14198;
    n2734_o2 <= n14201;
    n2735_o2 <= n14204;
    n2711_o2 <= n14207;
    lo585_buf_o2 <= n14210;
    n2719_o2 <= n14213;
    n2720_o2 <= n14216;
    n2723_o2 <= n14219;
    n2724_o2 <= n14222;
    n3624_o2 <= n14225;
    n3625_o2 <= n14228;
    n3015_o2 <= n14231;
    n3491_o2 <= n14234;
    n2779_inv <= n14237;
    n2811_o2 <= n14240;
    n3010_o2 <= n14243;
    n3012_o2 <= n14246;
    lo382_buf_o2 <= n14249;
    lo386_buf_o2 <= n14252;
    lo390_buf_o2 <= n14255;
    lo398_buf_o2 <= n14258;
    lo402_buf_o2 <= n14261;
    lo406_buf_o2 <= n14264;
    n3492_o2 <= n14267;
    lo366_buf_o2 <= n14270;
    lo374_buf_o2 <= n14273;
    lo426_buf_o2 <= n14276;
    lo494_buf_o2 <= n14279;
    n2653_o2 <= n14282;
    n2654_o2 <= n14285;
    n2715_o2 <= n14288;
    n2740_o2 <= n14291;
    n2682_o2 <= n14294;
    n2736_o2 <= n14297;
    lo508_buf_o2 <= n14300;
    lo512_buf_o2 <= n14303;
    lo536_buf_o2 <= n14306;
    lo576_buf_o2 <= n14309;
    lo357_buf_o2 <= n14312;
    lo361_buf_o2 <= n14315;
    lo417_buf_o2 <= n14318;
    lo421_buf_o2 <= n14321;
    lo473_buf_o2 <= n14324;
    lo477_buf_o2 <= n14327;
    lo553_buf_o2 <= n14330;
    lo557_buf_o2 <= n14333;
    lo573_buf_o2 <= n14336;
    lo434_buf_o2 <= n14339;
    lo438_buf_o2 <= n14342;
    lo466_buf_o2 <= n14345;
    lo470_buf_o2 <= n14348;
    lo490_buf_o2 <= n14351;
    n2657_o2 <= n14354;
    n2658_o2 <= n14357;
    n2663_o2 <= n14360;
    n2664_o2 <= n14363;
    n2684_o2 <= n14366;
    n2685_o2 <= n14369;
  end
  initial begin
    n2610_lo <= 1'b0;
    n2613_lo <= 1'b0;
    n2616_lo <= 1'b0;
    n2619_lo <= 1'b0;
    n2622_lo <= 1'b0;
    n2625_lo <= 1'b0;
    n2628_lo <= 1'b0;
    n2634_lo <= 1'b0;
    n2637_lo <= 1'b0;
    n2640_lo <= 1'b0;
    n2643_lo <= 1'b0;
    n2646_lo <= 1'b0;
    n2649_lo <= 1'b0;
    n2652_lo <= 1'b0;
    n2655_lo <= 1'b0;
    n2658_lo <= 1'b0;
    n2661_lo <= 1'b0;
    n2664_lo <= 1'b0;
    n2667_lo <= 1'b0;
    n2670_lo <= 1'b0;
    n2673_lo <= 1'b0;
    n2676_lo <= 1'b0;
    n2679_lo <= 1'b0;
    n2682_lo <= 1'b0;
    n2685_lo <= 1'b0;
    n2688_lo <= 1'b0;
    n2691_lo <= 1'b0;
    n2694_lo <= 1'b0;
    n2697_lo <= 1'b0;
    n2700_lo <= 1'b0;
    n2703_lo <= 1'b0;
    n2706_lo <= 1'b0;
    n2709_lo <= 1'b0;
    n2712_lo <= 1'b0;
    n2715_lo <= 1'b0;
    n2718_lo <= 1'b0;
    n2721_lo <= 1'b0;
    n2724_lo <= 1'b0;
    n2727_lo <= 1'b0;
    n2730_lo <= 1'b0;
    n2733_lo <= 1'b0;
    n2736_lo <= 1'b0;
    n2739_lo <= 1'b0;
    n2742_lo <= 1'b0;
    n2745_lo <= 1'b0;
    n2748_lo <= 1'b0;
    n2751_lo <= 1'b0;
    n2754_lo <= 1'b0;
    n2757_lo <= 1'b0;
    n2760_lo <= 1'b0;
    n2763_lo <= 1'b0;
    n2766_lo <= 1'b0;
    n2769_lo <= 1'b0;
    n2772_lo <= 1'b0;
    n2775_lo <= 1'b0;
    n2778_lo <= 1'b0;
    n2781_lo <= 1'b0;
    n2784_lo <= 1'b0;
    n2787_lo <= 1'b0;
    n2790_lo <= 1'b0;
    n2793_lo <= 1'b0;
    n2796_lo <= 1'b0;
    n2799_lo <= 1'b0;
    n2802_lo <= 1'b0;
    n2805_lo <= 1'b0;
    n2808_lo <= 1'b0;
    n2811_lo <= 1'b0;
    n2814_lo <= 1'b0;
    n2817_lo <= 1'b0;
    n2820_lo <= 1'b0;
    n2823_lo <= 1'b0;
    n2826_lo <= 1'b0;
    n2829_lo <= 1'b0;
    n2832_lo <= 1'b0;
    n2838_lo <= 1'b0;
    n2841_lo <= 1'b0;
    n2844_lo <= 1'b0;
    n2847_lo <= 1'b0;
    n2850_lo <= 1'b0;
    n2853_lo <= 1'b0;
    n2856_lo <= 1'b0;
    n2862_lo <= 1'b0;
    n2865_lo <= 1'b0;
    n2868_lo <= 1'b0;
    n2871_lo <= 1'b0;
    n2874_lo <= 1'b0;
    n2877_lo <= 1'b0;
    n2880_lo <= 1'b0;
    n2883_lo <= 1'b0;
    n2886_lo <= 1'b0;
    n2889_lo <= 1'b0;
    n2892_lo <= 1'b0;
    n2895_lo <= 1'b0;
    n2898_lo <= 1'b0;
    n2901_lo <= 1'b0;
    n2904_lo <= 1'b0;
    n2907_lo <= 1'b0;
    n2910_lo <= 1'b0;
    n2913_lo <= 1'b0;
    n2916_lo <= 1'b0;
    n2919_lo <= 1'b0;
    n2922_lo <= 1'b0;
    n2925_lo <= 1'b0;
    n2928_lo <= 1'b0;
    n2931_lo <= 1'b0;
    n2934_lo <= 1'b0;
    n2937_lo <= 1'b0;
    n2940_lo <= 1'b0;
    n2943_lo <= 1'b0;
    n2946_lo <= 1'b0;
    n2949_lo <= 1'b0;
    n2952_lo <= 1'b0;
    n2955_lo <= 1'b0;
    n2958_lo <= 1'b0;
    n2961_lo <= 1'b0;
    n2964_lo <= 1'b0;
    n2967_lo <= 1'b0;
    n2970_lo <= 1'b0;
    n2973_lo <= 1'b0;
    n2976_lo <= 1'b0;
    n2979_lo <= 1'b0;
    n2982_lo <= 1'b0;
    n2985_lo <= 1'b0;
    n2988_lo <= 1'b0;
    n2991_lo <= 1'b0;
    n2994_lo <= 1'b0;
    n2997_lo <= 1'b0;
    n3000_lo <= 1'b0;
    n3003_lo <= 1'b0;
    n3006_lo <= 1'b0;
    n3009_lo <= 1'b0;
    n3012_lo <= 1'b0;
    n3015_lo <= 1'b0;
    n3018_lo <= 1'b0;
    n3021_lo <= 1'b0;
    n3024_lo <= 1'b0;
    n3027_lo <= 1'b0;
    n3030_lo <= 1'b0;
    n3033_lo <= 1'b0;
    n3036_lo <= 1'b0;
    n3039_lo <= 1'b0;
    n3042_lo <= 1'b0;
    n3045_lo <= 1'b0;
    n3048_lo <= 1'b0;
    n3051_lo <= 1'b0;
    n3054_lo <= 1'b0;
    n3057_lo <= 1'b0;
    n3060_lo <= 1'b0;
    n3063_lo <= 1'b0;
    n3066_lo <= 1'b0;
    n3069_lo <= 1'b0;
    n3072_lo <= 1'b0;
    n3075_lo <= 1'b0;
    n3078_lo <= 1'b0;
    n3081_lo <= 1'b0;
    n3084_lo <= 1'b0;
    n3087_lo <= 1'b0;
    n3090_lo <= 1'b0;
    n3093_lo <= 1'b0;
    n3096_lo <= 1'b0;
    n3099_lo <= 1'b0;
    n3102_lo <= 1'b0;
    n3105_lo <= 1'b0;
    n3108_lo <= 1'b0;
    n3111_lo <= 1'b0;
    n3114_lo <= 1'b0;
    n3117_lo <= 1'b0;
    n3120_lo <= 1'b0;
    n3126_lo <= 1'b0;
    n3129_lo <= 1'b0;
    n3132_lo <= 1'b0;
    n3138_lo <= 1'b0;
    n3141_lo <= 1'b0;
    n3144_lo <= 1'b0;
    n3147_lo <= 1'b0;
    n3150_lo <= 1'b0;
    n3153_lo <= 1'b0;
    n3156_lo <= 1'b0;
    n3162_lo <= 1'b0;
    n3165_lo <= 1'b0;
    n3168_lo <= 1'b0;
    n3174_lo <= 1'b0;
    n3177_lo <= 1'b0;
    n3180_lo <= 1'b0;
    n3186_lo <= 1'b0;
    n3189_lo <= 1'b0;
    n3192_lo <= 1'b0;
    n3195_lo <= 1'b0;
    n3198_lo <= 1'b0;
    n3201_lo <= 1'b0;
    n3204_lo <= 1'b0;
    n3210_lo <= 1'b0;
    n3213_lo <= 1'b0;
    n3216_lo <= 1'b0;
    n3219_lo <= 1'b0;
    n3222_lo <= 1'b0;
    n3225_lo <= 1'b0;
    n3228_lo <= 1'b0;
    n3234_lo <= 1'b0;
    n3237_lo <= 1'b0;
    n3240_lo <= 1'b0;
    n3243_lo <= 1'b0;
    n3246_lo <= 1'b0;
    n3249_lo <= 1'b0;
    n3252_lo <= 1'b0;
    n3255_lo <= 1'b0;
    n3258_lo <= 1'b0;
    n3261_lo <= 1'b0;
    n3264_lo <= 1'b0;
    n3267_lo <= 1'b0;
    n3270_lo <= 1'b0;
    n3273_lo <= 1'b0;
    n3276_lo <= 1'b0;
    n3279_lo <= 1'b0;
    n3282_lo <= 1'b0;
    n3285_lo <= 1'b0;
    n3288_lo <= 1'b0;
    n3294_lo <= 1'b0;
    n3297_lo <= 1'b0;
    n3300_lo <= 1'b0;
    n3306_lo <= 1'b0;
    n3309_lo <= 1'b0;
    n3312_lo <= 1'b0;
    n3318_lo <= 1'b0;
    n3321_lo <= 1'b0;
    n3324_lo <= 1'b0;
    n3330_lo <= 1'b0;
    n3333_lo <= 1'b0;
    n3336_lo <= 1'b0;
    n3339_lo <= 1'b0;
    n3342_lo <= 1'b0;
    n3345_lo <= 1'b0;
    n3348_lo <= 1'b0;
    n3351_lo <= 1'b0;
    n3354_lo <= 1'b0;
    n3357_lo <= 1'b0;
    n3360_lo <= 1'b0;
    n3363_lo <= 1'b0;
    n3366_lo <= 1'b0;
    n3369_lo <= 1'b0;
    n3372_lo <= 1'b0;
    n3375_lo <= 1'b0;
    n3378_lo <= 1'b0;
    n3381_lo <= 1'b0;
    n3384_lo <= 1'b0;
    n3387_lo <= 1'b0;
    n3390_lo <= 1'b0;
    n3393_lo <= 1'b0;
    n3396_lo <= 1'b0;
    n3399_lo <= 1'b0;
    n3402_lo <= 1'b0;
    n3405_lo <= 1'b0;
    n3408_lo <= 1'b0;
    n3411_lo <= 1'b0;
    n3414_lo <= 1'b0;
    n3417_lo <= 1'b0;
    n3420_lo <= 1'b0;
    n3423_lo <= 1'b0;
    n3426_lo <= 1'b0;
    n3429_lo <= 1'b0;
    n3432_lo <= 1'b0;
    n3435_lo <= 1'b0;
    n3438_lo <= 1'b0;
    n3441_lo <= 1'b0;
    n3444_lo <= 1'b0;
    n3447_lo <= 1'b0;
    n3450_lo <= 1'b0;
    n3453_lo <= 1'b0;
    n3456_lo <= 1'b0;
    n3459_lo <= 1'b0;
    n3462_lo <= 1'b0;
    n3465_lo <= 1'b0;
    n3468_lo <= 1'b0;
    n3471_lo <= 1'b0;
    n3474_lo <= 1'b0;
    n3477_lo <= 1'b0;
    n3480_lo <= 1'b0;
    n3483_lo <= 1'b0;
    n3486_lo <= 1'b0;
    n3489_lo <= 1'b0;
    n3492_lo <= 1'b0;
    n3495_lo <= 1'b0;
    n3498_lo <= 1'b0;
    n3501_lo <= 1'b0;
    n3504_lo <= 1'b0;
    n3507_lo <= 1'b0;
    n3510_lo <= 1'b0;
    n3513_lo <= 1'b0;
    n3516_lo <= 1'b0;
    n3519_lo <= 1'b0;
    n3522_lo <= 1'b0;
    n3525_lo <= 1'b0;
    n3528_lo <= 1'b0;
    n3531_lo <= 1'b0;
    n3534_lo <= 1'b0;
    n3537_lo <= 1'b0;
    n3540_lo <= 1'b0;
    n3543_lo <= 1'b0;
    n3546_lo <= 1'b0;
    n3549_lo <= 1'b0;
    n3552_lo <= 1'b0;
    n3555_lo <= 1'b0;
    n3558_lo <= 1'b0;
    n3561_lo <= 1'b0;
    n3564_lo <= 1'b0;
    n3567_lo <= 1'b0;
    n3570_lo <= 1'b0;
    n3573_lo <= 1'b0;
    n3576_lo <= 1'b0;
    n3579_lo <= 1'b0;
    n3582_lo <= 1'b0;
    n3585_lo <= 1'b0;
    n3588_lo <= 1'b0;
    n3591_lo <= 1'b0;
    n3594_lo <= 1'b0;
    n3597_lo <= 1'b0;
    n3600_lo <= 1'b0;
    n3603_lo <= 1'b0;
    n3606_lo <= 1'b0;
    n3609_lo <= 1'b0;
    n3612_lo <= 1'b0;
    n3615_lo <= 1'b0;
    n3618_lo <= 1'b0;
    n3621_lo <= 1'b0;
    n3624_lo <= 1'b0;
    n3627_lo <= 1'b0;
    n3630_lo <= 1'b0;
    n3633_lo <= 1'b0;
    n3636_lo <= 1'b0;
    n3639_lo <= 1'b0;
    n3642_lo <= 1'b0;
    n3645_lo <= 1'b0;
    n3648_lo <= 1'b0;
    n3651_lo <= 1'b0;
    n3654_lo <= 1'b0;
    n3666_lo <= 1'b0;
    n3750_lo <= 1'b0;
    n3762_lo <= 1'b0;
    n3774_lo <= 1'b0;
    n3786_lo <= 1'b0;
    n3789_lo <= 1'b0;
    n3792_lo <= 1'b0;
    n3795_lo <= 1'b0;
    n3798_lo <= 1'b0;
    n3810_lo <= 1'b0;
    n3822_lo <= 1'b0;
    n3834_lo <= 1'b0;
    n3846_lo <= 1'b0;
    n3930_lo <= 1'b0;
    n3933_lo <= 1'b0;
    n3936_lo <= 1'b0;
    n3942_lo <= 1'b0;
    n3945_lo <= 1'b0;
    n3948_lo <= 1'b0;
    n3954_lo <= 1'b0;
    n3957_lo <= 1'b0;
    n3963_lo <= 1'b0;
    n3966_lo <= 1'b0;
    n3969_lo <= 1'b0;
    n3975_lo <= 1'b0;
    n3978_lo <= 1'b0;
    n3990_lo <= 1'b0;
    n4050_lo <= 1'b0;
    n4062_lo <= 1'b0;
    n4098_lo <= 1'b0;
    n4107_lo <= 1'b0;
    n4110_lo <= 1'b0;
    n4122_lo <= 1'b0;
    n4131_lo <= 1'b0;
    n4155_lo <= 1'b0;
    n4158_lo <= 1'b0;
    n4170_lo <= 1'b0;
    n4179_lo <= 1'b0;
    n4182_lo <= 1'b0;
    n4185_lo <= 1'b0;
    n4188_lo <= 1'b0;
    n4194_lo <= 1'b0;
    n4197_lo <= 1'b0;
    n4200_lo <= 1'b0;
    n4206_lo <= 1'b0;
    n4209_lo <= 1'b0;
    n4212_lo <= 1'b0;
    n4215_lo <= 1'b0;
    n4230_lo <= 1'b0;
    n4233_lo <= 1'b0;
    n4236_lo <= 1'b0;
    n4239_lo <= 1'b0;
    n4242_lo <= 1'b0;
    n4254_lo <= 1'b0;
    n4290_lo <= 1'b0;
    n4293_lo <= 1'b0;
    n4302_lo <= 1'b0;
    n4314_lo <= 1'b0;
    n4350_lo <= 1'b0;
    n4362_lo <= 1'b0;
    n4374_lo <= 1'b0;
    n4386_lo <= 1'b0;
    n4398_lo <= 1'b0;
    n4410_lo <= 1'b0;
    n4413_lo <= 1'b0;
    n4416_lo <= 1'b0;
    n4419_lo <= 1'b0;
    n4422_lo <= 1'b0;
    n4425_lo <= 1'b0;
    n4428_lo <= 1'b0;
    n4431_lo <= 1'b0;
    n4434_lo <= 1'b0;
    n4437_lo <= 1'b0;
    n4440_lo <= 1'b0;
    n4443_lo <= 1'b0;
    n4446_lo <= 1'b0;
    n4449_lo <= 1'b0;
    n4452_lo <= 1'b0;
    n4455_lo <= 1'b0;
    n4458_lo <= 1'b0;
    n4461_lo <= 1'b0;
    n4464_lo <= 1'b0;
    n4467_lo <= 1'b0;
    n4470_lo <= 1'b0;
    n4473_lo <= 1'b0;
    n4476_lo <= 1'b0;
    n4479_lo <= 1'b0;
    n4482_lo <= 1'b0;
    n4485_lo <= 1'b0;
    n4488_lo <= 1'b0;
    n4494_lo <= 1'b0;
    n4497_lo <= 1'b0;
    n4500_lo <= 1'b0;
    n4503_lo <= 1'b0;
    n4506_lo <= 1'b0;
    n4509_lo <= 1'b0;
    n4512_lo <= 1'b0;
    n4515_lo <= 1'b0;
    n4518_lo <= 1'b0;
    n4521_lo <= 1'b0;
    n4524_lo <= 1'b0;
    n4527_lo <= 1'b0;
    n4530_lo <= 1'b0;
    n4533_lo <= 1'b0;
    n4536_lo <= 1'b0;
    n4539_lo <= 1'b0;
    n4542_lo <= 1'b0;
    n4545_lo <= 1'b0;
    n4554_lo <= 1'b0;
    n4557_lo <= 1'b0;
    n4560_lo <= 1'b0;
    n4563_lo <= 1'b0;
    n4566_lo <= 1'b0;
    n4569_lo <= 1'b0;
    n4572_lo <= 1'b0;
    n4575_lo <= 1'b0;
    n4578_lo <= 1'b0;
    n4581_lo <= 1'b0;
    n4584_lo <= 1'b0;
    n4587_lo <= 1'b0;
    n4590_lo <= 1'b0;
    n4593_lo <= 1'b0;
    n4596_lo <= 1'b0;
    n4602_lo <= 1'b0;
    n4605_lo <= 1'b0;
    n4608_lo <= 1'b0;
    n4614_lo <= 1'b0;
    n4617_lo <= 1'b0;
    n4620_lo <= 1'b0;
    n4626_lo <= 1'b0;
    n4629_lo <= 1'b0;
    n4632_lo <= 1'b0;
    n4638_lo <= 1'b0;
    n4641_lo <= 1'b0;
    n4644_lo <= 1'b0;
    n4647_lo <= 1'b0;
    n4650_lo <= 1'b0;
    n4653_lo <= 1'b0;
    n4656_lo <= 1'b0;
    n4659_lo <= 1'b0;
    n4662_lo <= 1'b0;
    n4665_lo <= 1'b0;
    n4668_lo <= 1'b0;
    n4671_lo <= 1'b0;
    n4674_lo <= 1'b0;
    n4677_lo <= 1'b0;
    n4680_lo <= 1'b0;
    n4683_lo <= 1'b0;
    n4686_lo <= 1'b0;
    n4689_lo <= 1'b0;
    n4692_lo <= 1'b0;
    n4695_lo <= 1'b0;
    n4698_lo <= 1'b0;
    n4701_lo <= 1'b0;
    n4704_lo <= 1'b0;
    n4707_lo <= 1'b0;
    n4710_lo <= 1'b0;
    n4713_lo <= 1'b0;
    n4716_lo <= 1'b0;
    n4719_lo <= 1'b0;
    n4722_lo <= 1'b0;
    n4725_lo <= 1'b0;
    n4728_lo <= 1'b0;
    n4731_lo <= 1'b0;
    n4734_lo <= 1'b0;
    n4737_lo <= 1'b0;
    n4740_lo <= 1'b0;
    n4743_lo <= 1'b0;
    n4970_o2 <= 1'b0;
    n4972_o2 <= 1'b0;
    n4989_o2 <= 1'b0;
    n5024_o2 <= 1'b0;
    n5025_o2 <= 1'b0;
    n5029_o2 <= 1'b0;
    n5042_o2 <= 1'b0;
    n5048_o2 <= 1'b0;
    n5093_o2 <= 1'b0;
    n5096_o2 <= 1'b0;
    n5193_o2 <= 1'b0;
    n5199_o2 <= 1'b0;
    n5203_o2 <= 1'b0;
    n5214_o2 <= 1'b0;
    n5221_o2 <= 1'b0;
    n5222_o2 <= 1'b0;
    n5273_o2 <= 1'b0;
    n5365_o2 <= 1'b0;
    n5385_o2 <= 1'b0;
    n5553_o2 <= 1'b0;
    n5636_o2 <= 1'b0;
    n5782_o2 <= 1'b0;
    n5778_o2 <= 1'b0;
    n5323_o2 <= 1'b0;
    n5325_o2 <= 1'b0;
    n5327_o2 <= 1'b0;
    n5329_o2 <= 1'b0;
    n5816_o2 <= 1'b0;
    n5817_o2 <= 1'b0;
    n5837_o2 <= 1'b0;
    n5844_o2 <= 1'b0;
    n5859_o2 <= 1'b0;
    n5857_o2 <= 1'b0;
    n5369_o2 <= 1'b0;
    n5371_o2 <= 1'b0;
    n5373_o2 <= 1'b0;
    n5400_o2 <= 1'b0;
    n5402_o2 <= 1'b0;
    n5404_o2 <= 1'b0;
    n5406_o2 <= 1'b0;
    n5407_o2 <= 1'b0;
    n5408_o2 <= 1'b0;
    n2722_o2 <= 1'b0;
    n1942_inv <= 1'b0;
    n5412_o2 <= 1'b0;
    n1948_inv <= 1'b0;
    n5557_o2 <= 1'b0;
    n5558_o2 <= 1'b0;
    n5559_o2 <= 1'b0;
    n5564_o2 <= 1'b0;
    n5565_o2 <= 1'b0;
    n1966_inv <= 1'b0;
    n5568_o2 <= 1'b0;
    n5598_o2 <= 1'b0;
    n5600_o2 <= 1'b0;
    n5601_o2 <= 1'b0;
    n5602_o2 <= 1'b0;
    n5603_o2 <= 1'b0;
    n2853_o2 <= 1'b0;
    n5637_o2 <= 1'b0;
    n1993_inv <= 1'b0;
    n1996_inv <= 1'b0;
    n5635_o2 <= 1'b0;
    n5640_o2 <= 1'b0;
    n5641_o2 <= 1'b0;
    n5642_o2 <= 1'b0;
    n5650_o2 <= 1'b0;
    n5652_o2 <= 1'b0;
    n5653_o2 <= 1'b0;
    n5654_o2 <= 1'b0;
    n5655_o2 <= 1'b0;
    n5657_o2 <= 1'b0;
    n2029_inv <= 1'b0;
    n5661_o2 <= 1'b0;
    n5656_o2 <= 1'b0;
    n5663_o2 <= 1'b0;
    n2041_inv <= 1'b0;
    n5795_o2 <= 1'b0;
    n5796_o2 <= 1'b0;
    n5797_o2 <= 1'b0;
    n5739_o2 <= 1'b0;
    n5773_o2 <= 1'b0;
    n2059_inv <= 1'b0;
    n5799_o2 <= 1'b0;
    n5802_o2 <= 1'b0;
    n2068_inv <= 1'b0;
    n5831_o2 <= 1'b0;
    n5833_o2 <= 1'b0;
    n5820_o2 <= 1'b0;
    n5823_o2 <= 1'b0;
    n5824_o2 <= 1'b0;
    n5869_o2 <= 1'b0;
    n5848_o2 <= 1'b0;
    n5849_o2 <= 1'b0;
    n5856_o2 <= 1'b0;
    n5896_o2 <= 1'b0;
    n2754_o2 <= 1'b0;
    n2908_o2 <= 1'b0;
    n5892_o2 <= 1'b0;
    n5915_o2 <= 1'b0;
    n5919_o2 <= 1'b0;
    n5918_o2 <= 1'b0;
    n5920_o2 <= 1'b0;
    n5917_o2 <= 1'b0;
    lo586_buf_o2 <= 1'b0;
    n2818_o2 <= 1'b0;
    n2863_o2 <= 1'b0;
    n2134_inv <= 1'b0;
    n2725_o2 <= 1'b0;
    n3016_o2 <= 1'b0;
    n3013_o2 <= 1'b0;
    n2655_o2 <= 1'b0;
    n2149_inv <= 1'b0;
    lo562_buf_o2 <= 1'b0;
    n2155_inv <= 1'b0;
    n2531_o2 <= 1'b0;
    n2700_o2 <= 1'b0;
    n5908_o2 <= 1'b0;
    n5910_o2 <= 1'b0;
    n5912_o2 <= 1'b0;
    n5914_o2 <= 1'b0;
    n2753_o2 <= 1'b0;
    n2878_o2 <= 1'b0;
    n2182_inv <= 1'b0;
    n5934_o2 <= 1'b0;
    n5936_o2 <= 1'b0;
    n5938_o2 <= 1'b0;
    n2728_o2 <= 1'b0;
    lo358_buf_o2 <= 1'b0;
    lo418_buf_o2 <= 1'b0;
    lo474_buf_o2 <= 1'b0;
    lo554_buf_o2 <= 1'b0;
    lo558_buf_o2 <= 1'b0;
    lo574_buf_o2 <= 1'b0;
    n2215_inv <= 1'b0;
    n2218_inv <= 1'b0;
    n2221_inv <= 1'b0;
    lo450_buf_o2 <= 1'b0;
    n2910_o2 <= 1'b0;
    n2683_o2 <= 1'b0;
    n2828_o2 <= 1'b0;
    n2582_o2 <= 1'b0;
    n2600_o2 <= 1'b0;
    n2542_o2 <= 1'b0;
    n2703_o2 <= 1'b0;
    lo510_buf_o2 <= 1'b0;
    lo514_buf_o2 <= 1'b0;
    lo538_buf_o2 <= 1'b0;
    lo578_buf_o2 <= 1'b0;
    n2260_inv <= 1'b0;
    n2666_o2 <= 1'b0;
    n2667_o2 <= 1'b0;
    n2660_o2 <= 1'b0;
    n2272_inv <= 1'b0;
    lo454_buf_o2 <= 1'b0;
    n3593_o2 <= 1'b0;
    n3048_o2 <= 1'b0;
    lo410_buf_o2 <= 1'b0;
    lo502_buf_o2 <= 1'b0;
    lo506_buf_o2 <= 1'b0;
    lo550_buf_o2 <= 1'b0;
    lo570_buf_o2 <= 1'b0;
    lo582_buf_o2 <= 1'b0;
    n2302_inv <= 1'b0;
    n2305_inv <= 1'b0;
    n3499_o2 <= 1'b0;
    n2311_inv <= 1'b0;
    n2870_o2 <= 1'b0;
    n2317_inv <= 1'b0;
    n2689_o2 <= 1'b0;
    n2323_inv <= 1'b0;
    n2662_o2 <= 1'b0;
    lo350_buf_o2 <= 1'b0;
    lo498_buf_o2 <= 1'b0;
    lo518_buf_o2 <= 1'b0;
    lo522_buf_o2 <= 1'b0;
    lo598_buf_o2 <= 1'b0;
    n2344_inv <= 1'b0;
    n2347_inv <= 1'b0;
    n2350_inv <= 1'b0;
    n2353_inv <= 1'b0;
    n2356_inv <= 1'b0;
    n2359_inv <= 1'b0;
    n2872_o2 <= 1'b0;
    n3313_o2 <= 1'b0;
    n3273_o2 <= 1'b0;
    n2848_o2 <= 1'b0;
    n2893_o2 <= 1'b0;
    n3267_o2 <= 1'b0;
    n2925_o2 <= 1'b0;
    n2839_o2 <= 1'b0;
    n2831_o2 <= 1'b0;
    n2558_o2 <= 1'b0;
    n2562_o2 <= 1'b0;
    n2825_o2 <= 1'b0;
    n3263_o2 <= 1'b0;
    n3517_o2 <= 1'b0;
    n2873_o2 <= 1'b0;
    n2926_o2 <= 1'b0;
    n3261_o2 <= 1'b0;
    n3268_o2 <= 1'b0;
    n3274_o2 <= 1'b0;
    n3314_o2 <= 1'b0;
    n3571_o2 <= 1'b0;
    n2950_o2 <= 1'b0;
    n2951_o2 <= 1'b0;
    n3022_o2 <= 1'b0;
    n3023_o2 <= 1'b0;
    n3057_o2 <= 1'b0;
    n3058_o2 <= 1'b0;
    n2931_o2 <= 1'b0;
    n2911_o2 <= 1'b0;
    n2959_o2 <= 1'b0;
    n2960_o2 <= 1'b0;
    n2922_o2 <= 1'b0;
    n2888_o2 <= 1'b0;
    n2889_o2 <= 1'b0;
    n3051_o2 <= 1'b0;
    n3052_o2 <= 1'b0;
    n3063_o2 <= 1'b0;
    n2845_o2 <= 1'b0;
    n2476_inv <= 1'b0;
    n3281_o2 <= 1'b0;
    n3294_o2 <= 1'b0;
    n2885_o2 <= 1'b0;
    n2786_o2 <= 1'b0;
    n2783_o2 <= 1'b0;
    n2801_o2 <= 1'b0;
    n2572_o2 <= 1'b0;
    n2628_o2 <= 1'b0;
    n2609_o2 <= 1'b0;
    n2618_o2 <= 1'b0;
    n2637_o2 <= 1'b0;
    n2525_o2 <= 1'b0;
    n2551_o2 <= 1'b0;
    n3759_o2 <= 1'b0;
    n2994_o2 <= 1'b0;
    n3040_o2 <= 1'b0;
    n2943_o2 <= 1'b0;
    n2991_o2 <= 1'b0;
    n3034_o2 <= 1'b0;
    n2881_o2 <= 1'b0;
    n3021_o2 <= 1'b0;
    n3062_o2 <= 1'b0;
    n2763_o2 <= 1'b0;
    n2764_o2 <= 1'b0;
    n2775_o2 <= 1'b0;
    n2776_o2 <= 1'b0;
    n2968_o2 <= 1'b0;
    n2969_o2 <= 1'b0;
    n2798_o2 <= 1'b0;
    n3661_o2 <= 1'b0;
    n2694_o2 <= 1'b0;
    n2572_inv <= 1'b0;
    n2817_o2 <= 1'b0;
    n2514_o2 <= 1'b0;
    n2501_o2 <= 1'b0;
    n2584_inv <= 1'b0;
    n2505_o2 <= 1'b0;
    n2492_o2 <= 1'b0;
    lo546_buf_o2 <= 1'b0;
    lo590_buf_o2 <= 1'b0;
    lo594_buf_o2 <= 1'b0;
    n2602_inv <= 1'b0;
    n2605_inv <= 1'b0;
    n2709_o2 <= 1'b0;
    n2611_inv <= 1'b0;
    n2614_inv <= 1'b0;
    n2617_inv <= 1'b0;
    n2620_inv <= 1'b0;
    n3590_o2 <= 1'b0;
    n3591_o2 <= 1'b0;
    n2629_inv <= 1'b0;
    n3638_o2 <= 1'b0;
    n3639_o2 <= 1'b0;
    n2638_inv <= 1'b0;
    n2641_inv <= 1'b0;
    lo458_buf_o2 <= 1'b0;
    lo482_buf_o2 <= 1'b0;
    lo566_buf_o2 <= 1'b0;
    n2718_o2 <= 1'b0;
    n3707_o2 <= 1'b0;
    n3671_o2 <= 1'b0;
    n3680_o2 <= 1'b0;
    n3749_o2 <= 1'b0;
    n3716_o2 <= 1'b0;
    n3692_o2 <= 1'b0;
    n2591_o2 <= 1'b0;
    n3478_o2 <= 1'b0;
    n3610_o2 <= 1'b0;
    n3611_o2 <= 1'b0;
    n2686_inv <= 1'b0;
    n2689_inv <= 1'b0;
    n2738_o2 <= 1'b0;
    n3616_o2 <= 1'b0;
    n3617_o2 <= 1'b0;
    n3031_o2 <= 1'b0;
    n2704_inv <= 1'b0;
    n3562_o2 <= 1'b0;
    n2502_o2 <= 1'b0;
    n3560_o2 <= 1'b0;
    n3554_o2 <= 1'b0;
    n3555_o2 <= 1'b0;
    n3536_o2 <= 1'b0;
    n3537_o2 <= 1'b0;
    n3508_o2 <= 1'b0;
    n3650_o2 <= 1'b0;
    n3740_o2 <= 1'b0;
    n3484_o2 <= 1'b0;
    n2740_inv <= 1'b0;
    n2734_o2 <= 1'b0;
    n2735_o2 <= 1'b0;
    n2711_o2 <= 1'b0;
    lo585_buf_o2 <= 1'b0;
    n2719_o2 <= 1'b0;
    n2720_o2 <= 1'b0;
    n2723_o2 <= 1'b0;
    n2724_o2 <= 1'b0;
    n3624_o2 <= 1'b0;
    n3625_o2 <= 1'b0;
    n3015_o2 <= 1'b0;
    n3491_o2 <= 1'b0;
    n2779_inv <= 1'b0;
    n2811_o2 <= 1'b0;
    n3010_o2 <= 1'b0;
    n3012_o2 <= 1'b0;
    lo382_buf_o2 <= 1'b0;
    lo386_buf_o2 <= 1'b0;
    lo390_buf_o2 <= 1'b0;
    lo398_buf_o2 <= 1'b0;
    lo402_buf_o2 <= 1'b0;
    lo406_buf_o2 <= 1'b0;
    n3492_o2 <= 1'b0;
    lo366_buf_o2 <= 1'b0;
    lo374_buf_o2 <= 1'b0;
    lo426_buf_o2 <= 1'b0;
    lo494_buf_o2 <= 1'b0;
    n2653_o2 <= 1'b0;
    n2654_o2 <= 1'b0;
    n2715_o2 <= 1'b0;
    n2740_o2 <= 1'b0;
    n2682_o2 <= 1'b0;
    n2736_o2 <= 1'b0;
    lo508_buf_o2 <= 1'b0;
    lo512_buf_o2 <= 1'b0;
    lo536_buf_o2 <= 1'b0;
    lo576_buf_o2 <= 1'b0;
    lo357_buf_o2 <= 1'b0;
    lo361_buf_o2 <= 1'b0;
    lo417_buf_o2 <= 1'b0;
    lo421_buf_o2 <= 1'b0;
    lo473_buf_o2 <= 1'b0;
    lo477_buf_o2 <= 1'b0;
    lo553_buf_o2 <= 1'b0;
    lo557_buf_o2 <= 1'b0;
    lo573_buf_o2 <= 1'b0;
    lo434_buf_o2 <= 1'b0;
    lo438_buf_o2 <= 1'b0;
    lo466_buf_o2 <= 1'b0;
    lo470_buf_o2 <= 1'b0;
    lo490_buf_o2 <= 1'b0;
    n2657_o2 <= 1'b0;
    n2658_o2 <= 1'b0;
    n2663_o2 <= 1'b0;
    n2664_o2 <= 1'b0;
    n2684_o2 <= 1'b0;
    n2685_o2 <= 1'b0;
  end
endmodule


