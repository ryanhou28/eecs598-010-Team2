
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  n949_lo,
  n961_lo,
  n973_lo,
  n976_lo,
  n985_lo,
  n997_lo,
  n1009_lo,
  n1021_lo,
  n1024_lo,
  n1033_lo,
  n1036_lo,
  n1045_lo,
  n1057_lo,
  n1069_lo,
  n1081_lo,
  n1093_lo,
  n1105_lo,
  n1117_lo,
  n1129_lo,
  n1132_lo,
  n1141_lo,
  n1144_lo,
  n1156_lo,
  n1159_lo,
  n1165_lo,
  n1168_lo,
  n1180_lo,
  n1189_lo,
  n1192_lo,
  n1201_lo,
  n1204_lo,
  n1216_lo,
  n1228_lo,
  n1231_lo,
  n1237_lo,
  n1240_lo,
  n1243_lo,
  n1249_lo,
  n1252_lo,
  n1255_lo,
  n1261_lo,
  n1264_lo,
  n1267_lo,
  n1273_lo,
  n1276_lo,
  n1279_lo,
  n1282_lo,
  n1285_lo,
  n1288_lo,
  n1291_lo,
  n1294_lo,
  n1297_lo,
  n1300_lo,
  n1303_lo,
  n1309_lo,
  n1312_lo,
  n1315_lo,
  n1318_lo,
  n1321_lo,
  n1324_lo,
  n1333_lo,
  n1874_o2,
  n2180_o2,
  n2372_o2,
  n2190_o2,
  n2191_o2,
  n2212_o2,
  n2213_o2,
  n2214_o2,
  n2215_o2,
  n2275_o2,
  n2276_o2,
  n2290_o2,
  n2291_o2,
  n2681_o2,
  n2680_o2,
  n2683_o2,
  n2684_o2,
  n2686_o2,
  n2319_o2,
  n2320_o2,
  n304_inv,
  G554_o2,
  G557_o2,
  G185_o2,
  G188_o2,
  G191_o2,
  G194_o2,
  G1182_o2,
  G1222_o2,
  G1247_o2,
  G1371_o2,
  G1383_o2,
  G1386_o2,
  n2416_o2,
  n2428_o2,
  n2438_o2,
  n2439_o2,
  n2440_o2,
  n2444_o2,
  n2497_o2,
  n2498_o2,
  n2503_o2,
  n2505_o2,
  n2529_o2,
  n2562_o2,
  n2570_o2,
  n2571_o2,
  n2574_o2,
  n2575_o2,
  G546_o2,
  G550_o2,
  n2633_o2,
  n2639_o2,
  n2642_o2,
  n2645_o2,
  n2679_o2,
  n2662_o2,
  n2724_o2,
  G382_o2,
  G199_o2,
  G202_o2,
  G225_o2,
  G248_o2,
  G260_o2,
  n2716_o2,
  n2737_o2,
  n1174_lo_buf_o2,
  n1198_lo_buf_o2,
  G371_o2,
  G1059_o2,
  n2586_o2,
  n2587_o2,
  n460_inv,
  n2648_o2,
  n2649_o2,
  n2650_o2,
  n2651_o2,
  n2652_o2,
  G365_o2,
  G1496_o2,
  G1502_o2,
  n2700_o2,
  n2701_o2,
  n2733_o2,
  n2734_o2,
  n2744_o2,
  n2747_o2,
  n2754_o2,
  n2755_o2,
  n511_inv,
  G1609_o2,
  G1625_o2,
  G738_o2,
  G755_o2,
  G1511_o2,
  G1522_o2,
  G1538_o2,
  G1549_o2,
  G1563_o2,
  G1584_o2,
  G1576_o2,
  G1598_o2,
  G1395_o2,
  G1410_o2,
  G1420_o2,
  G1434_o2,
  n562_inv,
  n1162_lo_buf_o2,
  n1102_lo_buf_o2,
  G359_o2,
  n982_lo_buf_o2,
  n1030_lo_buf_o2,
  n1042_lo_buf_o2,
  n583_inv,
  G606_o2,
  G1118_o2,
  G1069_o2,
  G1145_o2,
  G1209_o2,
  G1189_o2,
  G1699_o2,
  G1702_o2,
  G1705_o2,
  G1708_o2,
  G1684_o2,
  G1687_o2,
  G1690_o2,
  G1693_o2,
  G1696_o2,
  G1642_o2,
  G1645_o2,
  G1648_o2,
  G1651_o2,
  G1654_o2,
  G1657_o2,
  G1660_o2,
  n1222_lo_buf_o2,
  n1330_lo_buf_o2,
  n658_inv,
  n661_inv,
  n1306_lo_buf_o2,
  n1150_lo_buf_o2,
  G175_o2,
  G241_o2,
  G356_o2,
  G989_o2,
  G984_o2,
  n685_inv,
  n688_inv,
  n958_lo_buf_o2,
  n1114_lo_buf_o2,
  G182_o2,
  G1215_o2,
  G971_o2,
  G938_o2,
  G1198_o2,
  G1203_o2,
  G1218_o2,
  G785_o2,
  G1168_o2,
  G1130_o2,
  G1185_o2,
  G1250_o2,
  G1225_o2,
  G1791_o2,
  G1788_o2,
  G981_o2,
  n745_inv,
  n748_inv,
  G1062_o2,
  n970_lo_buf_o2,
  n1006_lo_buf_o2,
  n1078_lo_buf_o2,
  n1126_lo_buf_o2,
  n766_inv,
  G165_o2,
  n1234_lo_buf_o2,
  n1246_lo_buf_o2,
  n1258_lo_buf_o2,
  n1270_lo_buf_o2,
  G368_o2,
  G428_o2,
  G212_o2,
  G841_o2,
  G788_o2,
  n1186_lo_buf_o2,
  G391_o2,
  G387_o2,
  G645_o2,
  G1140_o2,
  G1178_o2,
  G1370_o2,
  n820_inv,
  G1357_o2,
  G816_o2,
  G1369_o2,
  G901_o2,
  G1056_o2,
  G1107_o2,
  G1087_o2,
  G1135_o2,
  n1018_lo_buf_o2,
  n1090_lo_buf_o2,
  n853_inv,
  G131_o2,
  n859_inv,
  n862_inv,
  G338_o2,
  n1171_lo_buf_o2,
  n1195_lo_buf_o2,
  G419_o2,
  G425_o2,
  G497_o2,
  G416_o2,
  G491_o2,
  G500_o2,
  G353_o2,
  G641_o2,
  G1117_o2,
  G1096_o2,
  G1143_o2,
  G1112_o2,
  n1138_lo_buf_o2,
  n1210_lo_buf_o2,
  G687_o2,
  G541_o2,
  G802_o2,
  G813_o2,
  G810_o2,
  G987_o2,
  G898_o2,
  n946_lo_buf_o2,
  n1054_lo_buf_o2,
  G728_o2,
  G856_o2,
  n949_1_inv,
  G942_o2,
  G1099_o2,
  G1154_o2,
  G1131_o2,
  G1169_o2,
  G134_o2,
  n970_inv,
  G470_o2,
  G344_o2,
  G362_o2,
  G482_o2,
  G660_o2,
  G672_o2,
  n1096_lo_buf_o2,
  G479_o2,
  G669_o2,
  n994_lo_buf_o2,
  n1066_lo_buf_o2,
  n1006_inv,
  G147_o2,
  G473_o2,
  G488_o2,
  G589_o2,
  G663_o2,
  G684_o2,
  G605_o2,
  G774_o2,
  G782_o2,
  G1884,
  G1885,
  G1886,
  G1887,
  G1888,
  G1889,
  G1890,
  G1891,
  G1892,
  G1893,
  G1894,
  G1895,
  G1896,
  G1897,
  G1898,
  G1899,
  G1900,
  G1901,
  G1902,
  G1903,
  G1904,
  G1905,
  G1906,
  G1907,
  G1908,
  n949_li,
  n961_li,
  n973_li,
  n976_li,
  n985_li,
  n997_li,
  n1009_li,
  n1021_li,
  n1024_li,
  n1033_li,
  n1036_li,
  n1045_li,
  n1057_li,
  n1069_li,
  n1081_li,
  n1093_li,
  n1105_li,
  n1117_li,
  n1129_li,
  n1132_li,
  n1141_li,
  n1144_li,
  n1156_li,
  n1159_li,
  n1165_li,
  n1168_li,
  n1180_li,
  n1189_li,
  n1192_li,
  n1201_li,
  n1204_li,
  n1216_li,
  n1228_li,
  n1231_li,
  n1237_li,
  n1240_li,
  n1243_li,
  n1249_li,
  n1252_li,
  n1255_li,
  n1261_li,
  n1264_li,
  n1267_li,
  n1273_li,
  n1276_li,
  n1279_li,
  n1282_li,
  n1285_li,
  n1288_li,
  n1291_li,
  n1294_li,
  n1297_li,
  n1300_li,
  n1303_li,
  n1309_li,
  n1312_li,
  n1315_li,
  n1318_li,
  n1321_li,
  n1324_li,
  n1333_li,
  n1874_i2,
  n2180_i2,
  n2372_i2,
  n2190_i2,
  n2191_i2,
  n2212_i2,
  n2213_i2,
  n2214_i2,
  n2215_i2,
  n2275_i2,
  n2276_i2,
  n2290_i2,
  n2291_i2,
  n2681_i2,
  n2680_i2,
  n2683_i2,
  n2684_i2,
  n2686_i2,
  n2319_i2,
  n2320_i2,
  n2321_i2,
  G554_i2,
  G557_i2,
  G185_i2,
  G188_i2,
  G191_i2,
  G194_i2,
  G1182_i2,
  G1222_i2,
  G1247_i2,
  G1371_i2,
  G1383_i2,
  G1386_i2,
  n2416_i2,
  n2428_i2,
  n2438_i2,
  n2439_i2,
  n2440_i2,
  n2444_i2,
  n2497_i2,
  n2498_i2,
  n2503_i2,
  n2505_i2,
  n2529_i2,
  n2562_i2,
  n2570_i2,
  n2571_i2,
  n2574_i2,
  n2575_i2,
  G546_i2,
  G550_i2,
  n2633_i2,
  n2639_i2,
  n2642_i2,
  n2645_i2,
  n2679_i2,
  n2662_i2,
  n2724_i2,
  G382_i2,
  G199_i2,
  G202_i2,
  G225_i2,
  G248_i2,
  G260_i2,
  n2716_i2,
  n2737_i2,
  n1174_lo_buf_i2,
  n1198_lo_buf_i2,
  G371_i2,
  G1059_i2,
  n2586_i2,
  n2587_i2,
  G1019_i2,
  n2648_i2,
  n2649_i2,
  n2650_i2,
  n2651_i2,
  n2652_i2,
  G365_i2,
  G1496_i2,
  G1502_i2,
  n2700_i2,
  n2701_i2,
  n2733_i2,
  n2734_i2,
  n2744_i2,
  n2747_i2,
  n2754_i2,
  n2755_i2,
  n2756_i2,
  G1609_i2,
  G1625_i2,
  G738_i2,
  G755_i2,
  G1511_i2,
  G1522_i2,
  G1538_i2,
  G1549_i2,
  G1563_i2,
  G1584_i2,
  G1576_i2,
  G1598_i2,
  G1395_i2,
  G1410_i2,
  G1420_i2,
  G1434_i2,
  G1240_i2,
  n1162_lo_buf_i2,
  n1102_lo_buf_i2,
  G359_i2,
  n982_lo_buf_i2,
  n1030_lo_buf_i2,
  n1042_lo_buf_i2,
  G161_i2,
  G606_i2,
  G1118_i2,
  G1069_i2,
  G1145_i2,
  G1209_i2,
  G1189_i2,
  G1699_i2,
  G1702_i2,
  G1705_i2,
  G1708_i2,
  G1684_i2,
  G1687_i2,
  G1690_i2,
  G1693_i2,
  G1696_i2,
  G1642_i2,
  G1645_i2,
  G1648_i2,
  G1651_i2,
  G1654_i2,
  G1657_i2,
  G1660_i2,
  n1222_lo_buf_i2,
  n1330_lo_buf_i2,
  G123_i2,
  G142_i2,
  n1306_lo_buf_i2,
  n1150_lo_buf_i2,
  G175_i2,
  G241_i2,
  G356_i2,
  G989_i2,
  G984_i2,
  G1009_i2,
  G1012_i2,
  n958_lo_buf_i2,
  n1114_lo_buf_i2,
  G182_i2,
  G1215_i2,
  G971_i2,
  G938_i2,
  G1198_i2,
  G1203_i2,
  G1218_i2,
  G785_i2,
  G1168_i2,
  G1130_i2,
  G1185_i2,
  G1250_i2,
  G1225_i2,
  G1791_i2,
  G1788_i2,
  G981_i2,
  G1031_i2,
  G1015_i2,
  G1062_i2,
  n970_lo_buf_i2,
  n1006_lo_buf_i2,
  n1078_lo_buf_i2,
  n1126_lo_buf_i2,
  G116_i2,
  G165_i2,
  n1234_lo_buf_i2,
  n1246_lo_buf_i2,
  n1258_lo_buf_i2,
  n1270_lo_buf_i2,
  G368_i2,
  G428_i2,
  G212_i2,
  G841_i2,
  G788_i2,
  n1186_lo_buf_i2,
  G391_i2,
  G387_i2,
  G645_i2,
  G1140_i2,
  G1178_i2,
  G1370_i2,
  G1205_i2,
  G1357_i2,
  G816_i2,
  G1369_i2,
  G901_i2,
  G1056_i2,
  G1107_i2,
  G1087_i2,
  G1135_i2,
  n1018_lo_buf_i2,
  n1090_lo_buf_i2,
  G119_i2,
  G131_i2,
  G154_i2,
  G169_i2,
  G338_i2,
  n1171_lo_buf_i2,
  n1195_lo_buf_i2,
  G419_i2,
  G425_i2,
  G497_i2,
  G416_i2,
  G491_i2,
  G500_i2,
  G353_i2,
  G641_i2,
  G1117_i2,
  G1096_i2,
  G1143_i2,
  G1112_i2,
  n1138_lo_buf_i2,
  n1210_lo_buf_i2,
  G687_i2,
  G541_i2,
  G802_i2,
  G813_i2,
  G810_i2,
  G987_i2,
  G898_i2,
  n946_lo_buf_i2,
  n1054_lo_buf_i2,
  G728_i2,
  G856_i2,
  G831_i2,
  G942_i2,
  G1099_i2,
  G1154_i2,
  G1131_i2,
  G1169_i2,
  G134_i2,
  G157_i2,
  G470_i2,
  G344_i2,
  G362_i2,
  G482_i2,
  G660_i2,
  G672_i2,
  n1096_lo_buf_i2,
  G479_i2,
  G669_i2,
  n994_lo_buf_i2,
  n1066_lo_buf_i2,
  G112_i2,
  G147_i2,
  G473_i2,
  G488_i2,
  G589_i2,
  G663_i2,
  G684_i2,
  G605_i2,
  G774_i2,
  G782_i2
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input n949_lo;input n961_lo;input n973_lo;input n976_lo;input n985_lo;input n997_lo;input n1009_lo;input n1021_lo;input n1024_lo;input n1033_lo;input n1036_lo;input n1045_lo;input n1057_lo;input n1069_lo;input n1081_lo;input n1093_lo;input n1105_lo;input n1117_lo;input n1129_lo;input n1132_lo;input n1141_lo;input n1144_lo;input n1156_lo;input n1159_lo;input n1165_lo;input n1168_lo;input n1180_lo;input n1189_lo;input n1192_lo;input n1201_lo;input n1204_lo;input n1216_lo;input n1228_lo;input n1231_lo;input n1237_lo;input n1240_lo;input n1243_lo;input n1249_lo;input n1252_lo;input n1255_lo;input n1261_lo;input n1264_lo;input n1267_lo;input n1273_lo;input n1276_lo;input n1279_lo;input n1282_lo;input n1285_lo;input n1288_lo;input n1291_lo;input n1294_lo;input n1297_lo;input n1300_lo;input n1303_lo;input n1309_lo;input n1312_lo;input n1315_lo;input n1318_lo;input n1321_lo;input n1324_lo;input n1333_lo;input n1874_o2;input n2180_o2;input n2372_o2;input n2190_o2;input n2191_o2;input n2212_o2;input n2213_o2;input n2214_o2;input n2215_o2;input n2275_o2;input n2276_o2;input n2290_o2;input n2291_o2;input n2681_o2;input n2680_o2;input n2683_o2;input n2684_o2;input n2686_o2;input n2319_o2;input n2320_o2;input n304_inv;input G554_o2;input G557_o2;input G185_o2;input G188_o2;input G191_o2;input G194_o2;input G1182_o2;input G1222_o2;input G1247_o2;input G1371_o2;input G1383_o2;input G1386_o2;input n2416_o2;input n2428_o2;input n2438_o2;input n2439_o2;input n2440_o2;input n2444_o2;input n2497_o2;input n2498_o2;input n2503_o2;input n2505_o2;input n2529_o2;input n2562_o2;input n2570_o2;input n2571_o2;input n2574_o2;input n2575_o2;input G546_o2;input G550_o2;input n2633_o2;input n2639_o2;input n2642_o2;input n2645_o2;input n2679_o2;input n2662_o2;input n2724_o2;input G382_o2;input G199_o2;input G202_o2;input G225_o2;input G248_o2;input G260_o2;input n2716_o2;input n2737_o2;input n1174_lo_buf_o2;input n1198_lo_buf_o2;input G371_o2;input G1059_o2;input n2586_o2;input n2587_o2;input n460_inv;input n2648_o2;input n2649_o2;input n2650_o2;input n2651_o2;input n2652_o2;input G365_o2;input G1496_o2;input G1502_o2;input n2700_o2;input n2701_o2;input n2733_o2;input n2734_o2;input n2744_o2;input n2747_o2;input n2754_o2;input n2755_o2;input n511_inv;input G1609_o2;input G1625_o2;input G738_o2;input G755_o2;input G1511_o2;input G1522_o2;input G1538_o2;input G1549_o2;input G1563_o2;input G1584_o2;input G1576_o2;input G1598_o2;input G1395_o2;input G1410_o2;input G1420_o2;input G1434_o2;input n562_inv;input n1162_lo_buf_o2;input n1102_lo_buf_o2;input G359_o2;input n982_lo_buf_o2;input n1030_lo_buf_o2;input n1042_lo_buf_o2;input n583_inv;input G606_o2;input G1118_o2;input G1069_o2;input G1145_o2;input G1209_o2;input G1189_o2;input G1699_o2;input G1702_o2;input G1705_o2;input G1708_o2;input G1684_o2;input G1687_o2;input G1690_o2;input G1693_o2;input G1696_o2;input G1642_o2;input G1645_o2;input G1648_o2;input G1651_o2;input G1654_o2;input G1657_o2;input G1660_o2;input n1222_lo_buf_o2;input n1330_lo_buf_o2;input n658_inv;input n661_inv;input n1306_lo_buf_o2;input n1150_lo_buf_o2;input G175_o2;input G241_o2;input G356_o2;input G989_o2;input G984_o2;input n685_inv;input n688_inv;input n958_lo_buf_o2;input n1114_lo_buf_o2;input G182_o2;input G1215_o2;input G971_o2;input G938_o2;input G1198_o2;input G1203_o2;input G1218_o2;input G785_o2;input G1168_o2;input G1130_o2;input G1185_o2;input G1250_o2;input G1225_o2;input G1791_o2;input G1788_o2;input G981_o2;input n745_inv;input n748_inv;input G1062_o2;input n970_lo_buf_o2;input n1006_lo_buf_o2;input n1078_lo_buf_o2;input n1126_lo_buf_o2;input n766_inv;input G165_o2;input n1234_lo_buf_o2;input n1246_lo_buf_o2;input n1258_lo_buf_o2;input n1270_lo_buf_o2;input G368_o2;input G428_o2;input G212_o2;input G841_o2;input G788_o2;input n1186_lo_buf_o2;input G391_o2;input G387_o2;input G645_o2;input G1140_o2;input G1178_o2;input G1370_o2;input n820_inv;input G1357_o2;input G816_o2;input G1369_o2;input G901_o2;input G1056_o2;input G1107_o2;input G1087_o2;input G1135_o2;input n1018_lo_buf_o2;input n1090_lo_buf_o2;input n853_inv;input G131_o2;input n859_inv;input n862_inv;input G338_o2;input n1171_lo_buf_o2;input n1195_lo_buf_o2;input G419_o2;input G425_o2;input G497_o2;input G416_o2;input G491_o2;input G500_o2;input G353_o2;input G641_o2;input G1117_o2;input G1096_o2;input G1143_o2;input G1112_o2;input n1138_lo_buf_o2;input n1210_lo_buf_o2;input G687_o2;input G541_o2;input G802_o2;input G813_o2;input G810_o2;input G987_o2;input G898_o2;input n946_lo_buf_o2;input n1054_lo_buf_o2;input G728_o2;input G856_o2;input n949_1_inv;input G942_o2;input G1099_o2;input G1154_o2;input G1131_o2;input G1169_o2;input G134_o2;input n970_inv;input G470_o2;input G344_o2;input G362_o2;input G482_o2;input G660_o2;input G672_o2;input n1096_lo_buf_o2;input G479_o2;input G669_o2;input n994_lo_buf_o2;input n1066_lo_buf_o2;input n1006_inv;input G147_o2;input G473_o2;input G488_o2;input G589_o2;input G663_o2;input G684_o2;input G605_o2;input G774_o2;input G782_o2;
  output G1884;output G1885;output G1886;output G1887;output G1888;output G1889;output G1890;output G1891;output G1892;output G1893;output G1894;output G1895;output G1896;output G1897;output G1898;output G1899;output G1900;output G1901;output G1902;output G1903;output G1904;output G1905;output G1906;output G1907;output G1908;output n949_li;output n961_li;output n973_li;output n976_li;output n985_li;output n997_li;output n1009_li;output n1021_li;output n1024_li;output n1033_li;output n1036_li;output n1045_li;output n1057_li;output n1069_li;output n1081_li;output n1093_li;output n1105_li;output n1117_li;output n1129_li;output n1132_li;output n1141_li;output n1144_li;output n1156_li;output n1159_li;output n1165_li;output n1168_li;output n1180_li;output n1189_li;output n1192_li;output n1201_li;output n1204_li;output n1216_li;output n1228_li;output n1231_li;output n1237_li;output n1240_li;output n1243_li;output n1249_li;output n1252_li;output n1255_li;output n1261_li;output n1264_li;output n1267_li;output n1273_li;output n1276_li;output n1279_li;output n1282_li;output n1285_li;output n1288_li;output n1291_li;output n1294_li;output n1297_li;output n1300_li;output n1303_li;output n1309_li;output n1312_li;output n1315_li;output n1318_li;output n1321_li;output n1324_li;output n1333_li;output n1874_i2;output n2180_i2;output n2372_i2;output n2190_i2;output n2191_i2;output n2212_i2;output n2213_i2;output n2214_i2;output n2215_i2;output n2275_i2;output n2276_i2;output n2290_i2;output n2291_i2;output n2681_i2;output n2680_i2;output n2683_i2;output n2684_i2;output n2686_i2;output n2319_i2;output n2320_i2;output n2321_i2;output G554_i2;output G557_i2;output G185_i2;output G188_i2;output G191_i2;output G194_i2;output G1182_i2;output G1222_i2;output G1247_i2;output G1371_i2;output G1383_i2;output G1386_i2;output n2416_i2;output n2428_i2;output n2438_i2;output n2439_i2;output n2440_i2;output n2444_i2;output n2497_i2;output n2498_i2;output n2503_i2;output n2505_i2;output n2529_i2;output n2562_i2;output n2570_i2;output n2571_i2;output n2574_i2;output n2575_i2;output G546_i2;output G550_i2;output n2633_i2;output n2639_i2;output n2642_i2;output n2645_i2;output n2679_i2;output n2662_i2;output n2724_i2;output G382_i2;output G199_i2;output G202_i2;output G225_i2;output G248_i2;output G260_i2;output n2716_i2;output n2737_i2;output n1174_lo_buf_i2;output n1198_lo_buf_i2;output G371_i2;output G1059_i2;output n2586_i2;output n2587_i2;output G1019_i2;output n2648_i2;output n2649_i2;output n2650_i2;output n2651_i2;output n2652_i2;output G365_i2;output G1496_i2;output G1502_i2;output n2700_i2;output n2701_i2;output n2733_i2;output n2734_i2;output n2744_i2;output n2747_i2;output n2754_i2;output n2755_i2;output n2756_i2;output G1609_i2;output G1625_i2;output G738_i2;output G755_i2;output G1511_i2;output G1522_i2;output G1538_i2;output G1549_i2;output G1563_i2;output G1584_i2;output G1576_i2;output G1598_i2;output G1395_i2;output G1410_i2;output G1420_i2;output G1434_i2;output G1240_i2;output n1162_lo_buf_i2;output n1102_lo_buf_i2;output G359_i2;output n982_lo_buf_i2;output n1030_lo_buf_i2;output n1042_lo_buf_i2;output G161_i2;output G606_i2;output G1118_i2;output G1069_i2;output G1145_i2;output G1209_i2;output G1189_i2;output G1699_i2;output G1702_i2;output G1705_i2;output G1708_i2;output G1684_i2;output G1687_i2;output G1690_i2;output G1693_i2;output G1696_i2;output G1642_i2;output G1645_i2;output G1648_i2;output G1651_i2;output G1654_i2;output G1657_i2;output G1660_i2;output n1222_lo_buf_i2;output n1330_lo_buf_i2;output G123_i2;output G142_i2;output n1306_lo_buf_i2;output n1150_lo_buf_i2;output G175_i2;output G241_i2;output G356_i2;output G989_i2;output G984_i2;output G1009_i2;output G1012_i2;output n958_lo_buf_i2;output n1114_lo_buf_i2;output G182_i2;output G1215_i2;output G971_i2;output G938_i2;output G1198_i2;output G1203_i2;output G1218_i2;output G785_i2;output G1168_i2;output G1130_i2;output G1185_i2;output G1250_i2;output G1225_i2;output G1791_i2;output G1788_i2;output G981_i2;output G1031_i2;output G1015_i2;output G1062_i2;output n970_lo_buf_i2;output n1006_lo_buf_i2;output n1078_lo_buf_i2;output n1126_lo_buf_i2;output G116_i2;output G165_i2;output n1234_lo_buf_i2;output n1246_lo_buf_i2;output n1258_lo_buf_i2;output n1270_lo_buf_i2;output G368_i2;output G428_i2;output G212_i2;output G841_i2;output G788_i2;output n1186_lo_buf_i2;output G391_i2;output G387_i2;output G645_i2;output G1140_i2;output G1178_i2;output G1370_i2;output G1205_i2;output G1357_i2;output G816_i2;output G1369_i2;output G901_i2;output G1056_i2;output G1107_i2;output G1087_i2;output G1135_i2;output n1018_lo_buf_i2;output n1090_lo_buf_i2;output G119_i2;output G131_i2;output G154_i2;output G169_i2;output G338_i2;output n1171_lo_buf_i2;output n1195_lo_buf_i2;output G419_i2;output G425_i2;output G497_i2;output G416_i2;output G491_i2;output G500_i2;output G353_i2;output G641_i2;output G1117_i2;output G1096_i2;output G1143_i2;output G1112_i2;output n1138_lo_buf_i2;output n1210_lo_buf_i2;output G687_i2;output G541_i2;output G802_i2;output G813_i2;output G810_i2;output G987_i2;output G898_i2;output n946_lo_buf_i2;output n1054_lo_buf_i2;output G728_i2;output G856_i2;output G831_i2;output G942_i2;output G1099_i2;output G1154_i2;output G1131_i2;output G1169_i2;output G134_i2;output G157_i2;output G470_i2;output G344_i2;output G362_i2;output G482_i2;output G660_i2;output G672_i2;output n1096_lo_buf_i2;output G479_i2;output G669_i2;output n994_lo_buf_i2;output n1066_lo_buf_i2;output G112_i2;output G147_i2;output G473_i2;output G488_i2;output G589_i2;output G663_i2;output G684_i2;output G605_i2;output G774_i2;output G782_i2;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire n949_lo_p;
  wire n949_lo_n;
  wire n961_lo_p;
  wire n961_lo_n;
  wire n973_lo_p;
  wire n973_lo_n;
  wire n976_lo_p;
  wire n976_lo_n;
  wire n985_lo_p;
  wire n985_lo_n;
  wire n997_lo_p;
  wire n997_lo_n;
  wire n1009_lo_p;
  wire n1009_lo_n;
  wire n1021_lo_p;
  wire n1021_lo_n;
  wire n1024_lo_p;
  wire n1024_lo_n;
  wire n1033_lo_p;
  wire n1033_lo_n;
  wire n1036_lo_p;
  wire n1036_lo_n;
  wire n1045_lo_p;
  wire n1045_lo_n;
  wire n1057_lo_p;
  wire n1057_lo_n;
  wire n1069_lo_p;
  wire n1069_lo_n;
  wire n1081_lo_p;
  wire n1081_lo_n;
  wire n1093_lo_p;
  wire n1093_lo_n;
  wire n1105_lo_p;
  wire n1105_lo_n;
  wire n1117_lo_p;
  wire n1117_lo_n;
  wire n1129_lo_p;
  wire n1129_lo_n;
  wire n1132_lo_p;
  wire n1132_lo_n;
  wire n1141_lo_p;
  wire n1141_lo_n;
  wire n1144_lo_p;
  wire n1144_lo_n;
  wire n1156_lo_p;
  wire n1156_lo_n;
  wire n1159_lo_p;
  wire n1159_lo_n;
  wire n1165_lo_p;
  wire n1165_lo_n;
  wire n1168_lo_p;
  wire n1168_lo_n;
  wire n1180_lo_p;
  wire n1180_lo_n;
  wire n1189_lo_p;
  wire n1189_lo_n;
  wire n1192_lo_p;
  wire n1192_lo_n;
  wire n1201_lo_p;
  wire n1201_lo_n;
  wire n1204_lo_p;
  wire n1204_lo_n;
  wire n1216_lo_p;
  wire n1216_lo_n;
  wire n1228_lo_p;
  wire n1228_lo_n;
  wire n1231_lo_p;
  wire n1231_lo_n;
  wire n1237_lo_p;
  wire n1237_lo_n;
  wire n1240_lo_p;
  wire n1240_lo_n;
  wire n1243_lo_p;
  wire n1243_lo_n;
  wire n1249_lo_p;
  wire n1249_lo_n;
  wire n1252_lo_p;
  wire n1252_lo_n;
  wire n1255_lo_p;
  wire n1255_lo_n;
  wire n1261_lo_p;
  wire n1261_lo_n;
  wire n1264_lo_p;
  wire n1264_lo_n;
  wire n1267_lo_p;
  wire n1267_lo_n;
  wire n1273_lo_p;
  wire n1273_lo_n;
  wire n1276_lo_p;
  wire n1276_lo_n;
  wire n1279_lo_p;
  wire n1279_lo_n;
  wire n1282_lo_p;
  wire n1282_lo_n;
  wire n1285_lo_p;
  wire n1285_lo_n;
  wire n1288_lo_p;
  wire n1288_lo_n;
  wire n1291_lo_p;
  wire n1291_lo_n;
  wire n1294_lo_p;
  wire n1294_lo_n;
  wire n1297_lo_p;
  wire n1297_lo_n;
  wire n1300_lo_p;
  wire n1300_lo_n;
  wire n1303_lo_p;
  wire n1303_lo_n;
  wire n1309_lo_p;
  wire n1309_lo_n;
  wire n1312_lo_p;
  wire n1312_lo_n;
  wire n1315_lo_p;
  wire n1315_lo_n;
  wire n1318_lo_p;
  wire n1318_lo_n;
  wire n1321_lo_p;
  wire n1321_lo_n;
  wire n1324_lo_p;
  wire n1324_lo_n;
  wire n1333_lo_p;
  wire n1333_lo_n;
  wire n1874_o2_p;
  wire n1874_o2_n;
  wire n2180_o2_p;
  wire n2180_o2_n;
  wire n2372_o2_p;
  wire n2372_o2_n;
  wire n2190_o2_p;
  wire n2190_o2_n;
  wire n2191_o2_p;
  wire n2191_o2_n;
  wire n2212_o2_p;
  wire n2212_o2_n;
  wire n2213_o2_p;
  wire n2213_o2_n;
  wire n2214_o2_p;
  wire n2214_o2_n;
  wire n2215_o2_p;
  wire n2215_o2_n;
  wire n2275_o2_p;
  wire n2275_o2_n;
  wire n2276_o2_p;
  wire n2276_o2_n;
  wire n2290_o2_p;
  wire n2290_o2_n;
  wire n2291_o2_p;
  wire n2291_o2_n;
  wire n2681_o2_p;
  wire n2681_o2_n;
  wire n2680_o2_p;
  wire n2680_o2_n;
  wire n2683_o2_p;
  wire n2683_o2_n;
  wire n2684_o2_p;
  wire n2684_o2_n;
  wire n2686_o2_p;
  wire n2686_o2_n;
  wire n2319_o2_p;
  wire n2319_o2_n;
  wire n2320_o2_p;
  wire n2320_o2_n;
  wire n304_inv_p;
  wire n304_inv_n;
  wire G554_o2_p;
  wire G554_o2_n;
  wire G557_o2_p;
  wire G557_o2_n;
  wire G185_o2_p;
  wire G185_o2_n;
  wire G188_o2_p;
  wire G188_o2_n;
  wire G191_o2_p;
  wire G191_o2_n;
  wire G194_o2_p;
  wire G194_o2_n;
  wire G1182_o2_p;
  wire G1182_o2_n;
  wire G1222_o2_p;
  wire G1222_o2_n;
  wire G1247_o2_p;
  wire G1247_o2_n;
  wire G1371_o2_p;
  wire G1371_o2_n;
  wire G1383_o2_p;
  wire G1383_o2_n;
  wire G1386_o2_p;
  wire G1386_o2_n;
  wire n2416_o2_p;
  wire n2416_o2_n;
  wire n2428_o2_p;
  wire n2428_o2_n;
  wire n2438_o2_p;
  wire n2438_o2_n;
  wire n2439_o2_p;
  wire n2439_o2_n;
  wire n2440_o2_p;
  wire n2440_o2_n;
  wire n2444_o2_p;
  wire n2444_o2_n;
  wire n2497_o2_p;
  wire n2497_o2_n;
  wire n2498_o2_p;
  wire n2498_o2_n;
  wire n2503_o2_p;
  wire n2503_o2_n;
  wire n2505_o2_p;
  wire n2505_o2_n;
  wire n2529_o2_p;
  wire n2529_o2_n;
  wire n2562_o2_p;
  wire n2562_o2_n;
  wire n2570_o2_p;
  wire n2570_o2_n;
  wire n2571_o2_p;
  wire n2571_o2_n;
  wire n2574_o2_p;
  wire n2574_o2_n;
  wire n2575_o2_p;
  wire n2575_o2_n;
  wire G546_o2_p;
  wire G546_o2_n;
  wire G550_o2_p;
  wire G550_o2_n;
  wire n2633_o2_p;
  wire n2633_o2_n;
  wire n2639_o2_p;
  wire n2639_o2_n;
  wire n2642_o2_p;
  wire n2642_o2_n;
  wire n2645_o2_p;
  wire n2645_o2_n;
  wire n2679_o2_p;
  wire n2679_o2_n;
  wire n2662_o2_p;
  wire n2662_o2_n;
  wire n2724_o2_p;
  wire n2724_o2_n;
  wire G382_o2_p;
  wire G382_o2_n;
  wire G199_o2_p;
  wire G199_o2_n;
  wire G202_o2_p;
  wire G202_o2_n;
  wire G225_o2_p;
  wire G225_o2_n;
  wire G248_o2_p;
  wire G248_o2_n;
  wire G260_o2_p;
  wire G260_o2_n;
  wire n2716_o2_p;
  wire n2716_o2_n;
  wire n2737_o2_p;
  wire n2737_o2_n;
  wire n1174_lo_buf_o2_p;
  wire n1174_lo_buf_o2_n;
  wire n1198_lo_buf_o2_p;
  wire n1198_lo_buf_o2_n;
  wire G371_o2_p;
  wire G371_o2_n;
  wire G1059_o2_p;
  wire G1059_o2_n;
  wire n2586_o2_p;
  wire n2586_o2_n;
  wire n2587_o2_p;
  wire n2587_o2_n;
  wire n460_inv_p;
  wire n460_inv_n;
  wire n2648_o2_p;
  wire n2648_o2_n;
  wire n2649_o2_p;
  wire n2649_o2_n;
  wire n2650_o2_p;
  wire n2650_o2_n;
  wire n2651_o2_p;
  wire n2651_o2_n;
  wire n2652_o2_p;
  wire n2652_o2_n;
  wire G365_o2_p;
  wire G365_o2_n;
  wire G1496_o2_p;
  wire G1496_o2_n;
  wire G1502_o2_p;
  wire G1502_o2_n;
  wire n2700_o2_p;
  wire n2700_o2_n;
  wire n2701_o2_p;
  wire n2701_o2_n;
  wire n2733_o2_p;
  wire n2733_o2_n;
  wire n2734_o2_p;
  wire n2734_o2_n;
  wire n2744_o2_p;
  wire n2744_o2_n;
  wire n2747_o2_p;
  wire n2747_o2_n;
  wire n2754_o2_p;
  wire n2754_o2_n;
  wire n2755_o2_p;
  wire n2755_o2_n;
  wire n511_inv_p;
  wire n511_inv_n;
  wire G1609_o2_p;
  wire G1609_o2_n;
  wire G1625_o2_p;
  wire G1625_o2_n;
  wire G738_o2_p;
  wire G738_o2_n;
  wire G755_o2_p;
  wire G755_o2_n;
  wire G1511_o2_p;
  wire G1511_o2_n;
  wire G1522_o2_p;
  wire G1522_o2_n;
  wire G1538_o2_p;
  wire G1538_o2_n;
  wire G1549_o2_p;
  wire G1549_o2_n;
  wire G1563_o2_p;
  wire G1563_o2_n;
  wire G1584_o2_p;
  wire G1584_o2_n;
  wire G1576_o2_p;
  wire G1576_o2_n;
  wire G1598_o2_p;
  wire G1598_o2_n;
  wire G1395_o2_p;
  wire G1395_o2_n;
  wire G1410_o2_p;
  wire G1410_o2_n;
  wire G1420_o2_p;
  wire G1420_o2_n;
  wire G1434_o2_p;
  wire G1434_o2_n;
  wire n562_inv_p;
  wire n562_inv_n;
  wire n1162_lo_buf_o2_p;
  wire n1162_lo_buf_o2_n;
  wire n1102_lo_buf_o2_p;
  wire n1102_lo_buf_o2_n;
  wire G359_o2_p;
  wire G359_o2_n;
  wire n982_lo_buf_o2_p;
  wire n982_lo_buf_o2_n;
  wire n1030_lo_buf_o2_p;
  wire n1030_lo_buf_o2_n;
  wire n1042_lo_buf_o2_p;
  wire n1042_lo_buf_o2_n;
  wire n583_inv_p;
  wire n583_inv_n;
  wire G606_o2_p;
  wire G606_o2_n;
  wire G1118_o2_p;
  wire G1118_o2_n;
  wire G1069_o2_p;
  wire G1069_o2_n;
  wire G1145_o2_p;
  wire G1145_o2_n;
  wire G1209_o2_p;
  wire G1209_o2_n;
  wire G1189_o2_p;
  wire G1189_o2_n;
  wire G1699_o2_p;
  wire G1699_o2_n;
  wire G1702_o2_p;
  wire G1702_o2_n;
  wire G1705_o2_p;
  wire G1705_o2_n;
  wire G1708_o2_p;
  wire G1708_o2_n;
  wire G1684_o2_p;
  wire G1684_o2_n;
  wire G1687_o2_p;
  wire G1687_o2_n;
  wire G1690_o2_p;
  wire G1690_o2_n;
  wire G1693_o2_p;
  wire G1693_o2_n;
  wire G1696_o2_p;
  wire G1696_o2_n;
  wire G1642_o2_p;
  wire G1642_o2_n;
  wire G1645_o2_p;
  wire G1645_o2_n;
  wire G1648_o2_p;
  wire G1648_o2_n;
  wire G1651_o2_p;
  wire G1651_o2_n;
  wire G1654_o2_p;
  wire G1654_o2_n;
  wire G1657_o2_p;
  wire G1657_o2_n;
  wire G1660_o2_p;
  wire G1660_o2_n;
  wire n1222_lo_buf_o2_p;
  wire n1222_lo_buf_o2_n;
  wire n1330_lo_buf_o2_p;
  wire n1330_lo_buf_o2_n;
  wire n658_inv_p;
  wire n658_inv_n;
  wire n661_inv_p;
  wire n661_inv_n;
  wire n1306_lo_buf_o2_p;
  wire n1306_lo_buf_o2_n;
  wire n1150_lo_buf_o2_p;
  wire n1150_lo_buf_o2_n;
  wire G175_o2_p;
  wire G175_o2_n;
  wire G241_o2_p;
  wire G241_o2_n;
  wire G356_o2_p;
  wire G356_o2_n;
  wire G989_o2_p;
  wire G989_o2_n;
  wire G984_o2_p;
  wire G984_o2_n;
  wire n685_inv_p;
  wire n685_inv_n;
  wire n688_inv_p;
  wire n688_inv_n;
  wire n958_lo_buf_o2_p;
  wire n958_lo_buf_o2_n;
  wire n1114_lo_buf_o2_p;
  wire n1114_lo_buf_o2_n;
  wire G182_o2_p;
  wire G182_o2_n;
  wire G1215_o2_p;
  wire G1215_o2_n;
  wire G971_o2_p;
  wire G971_o2_n;
  wire G938_o2_p;
  wire G938_o2_n;
  wire G1198_o2_p;
  wire G1198_o2_n;
  wire G1203_o2_p;
  wire G1203_o2_n;
  wire G1218_o2_p;
  wire G1218_o2_n;
  wire G785_o2_p;
  wire G785_o2_n;
  wire G1168_o2_p;
  wire G1168_o2_n;
  wire G1130_o2_p;
  wire G1130_o2_n;
  wire G1185_o2_p;
  wire G1185_o2_n;
  wire G1250_o2_p;
  wire G1250_o2_n;
  wire G1225_o2_p;
  wire G1225_o2_n;
  wire G1791_o2_p;
  wire G1791_o2_n;
  wire G1788_o2_p;
  wire G1788_o2_n;
  wire G981_o2_p;
  wire G981_o2_n;
  wire n745_inv_p;
  wire n745_inv_n;
  wire n748_inv_p;
  wire n748_inv_n;
  wire G1062_o2_p;
  wire G1062_o2_n;
  wire n970_lo_buf_o2_p;
  wire n970_lo_buf_o2_n;
  wire n1006_lo_buf_o2_p;
  wire n1006_lo_buf_o2_n;
  wire n1078_lo_buf_o2_p;
  wire n1078_lo_buf_o2_n;
  wire n1126_lo_buf_o2_p;
  wire n1126_lo_buf_o2_n;
  wire n766_inv_p;
  wire n766_inv_n;
  wire G165_o2_p;
  wire G165_o2_n;
  wire n1234_lo_buf_o2_p;
  wire n1234_lo_buf_o2_n;
  wire n1246_lo_buf_o2_p;
  wire n1246_lo_buf_o2_n;
  wire n1258_lo_buf_o2_p;
  wire n1258_lo_buf_o2_n;
  wire n1270_lo_buf_o2_p;
  wire n1270_lo_buf_o2_n;
  wire G368_o2_p;
  wire G368_o2_n;
  wire G428_o2_p;
  wire G428_o2_n;
  wire G212_o2_p;
  wire G212_o2_n;
  wire G841_o2_p;
  wire G841_o2_n;
  wire G788_o2_p;
  wire G788_o2_n;
  wire n1186_lo_buf_o2_p;
  wire n1186_lo_buf_o2_n;
  wire G391_o2_p;
  wire G391_o2_n;
  wire G387_o2_p;
  wire G387_o2_n;
  wire G645_o2_p;
  wire G645_o2_n;
  wire G1140_o2_p;
  wire G1140_o2_n;
  wire G1178_o2_p;
  wire G1178_o2_n;
  wire G1370_o2_p;
  wire G1370_o2_n;
  wire n820_inv_p;
  wire n820_inv_n;
  wire G1357_o2_p;
  wire G1357_o2_n;
  wire G816_o2_p;
  wire G816_o2_n;
  wire G1369_o2_p;
  wire G1369_o2_n;
  wire G901_o2_p;
  wire G901_o2_n;
  wire G1056_o2_p;
  wire G1056_o2_n;
  wire G1107_o2_p;
  wire G1107_o2_n;
  wire G1087_o2_p;
  wire G1087_o2_n;
  wire G1135_o2_p;
  wire G1135_o2_n;
  wire n1018_lo_buf_o2_p;
  wire n1018_lo_buf_o2_n;
  wire n1090_lo_buf_o2_p;
  wire n1090_lo_buf_o2_n;
  wire n853_inv_p;
  wire n853_inv_n;
  wire G131_o2_p;
  wire G131_o2_n;
  wire n859_inv_p;
  wire n859_inv_n;
  wire n862_inv_p;
  wire n862_inv_n;
  wire G338_o2_p;
  wire G338_o2_n;
  wire n1171_lo_buf_o2_p;
  wire n1171_lo_buf_o2_n;
  wire n1195_lo_buf_o2_p;
  wire n1195_lo_buf_o2_n;
  wire G419_o2_p;
  wire G419_o2_n;
  wire G425_o2_p;
  wire G425_o2_n;
  wire G497_o2_p;
  wire G497_o2_n;
  wire G416_o2_p;
  wire G416_o2_n;
  wire G491_o2_p;
  wire G491_o2_n;
  wire G500_o2_p;
  wire G500_o2_n;
  wire G353_o2_p;
  wire G353_o2_n;
  wire G641_o2_p;
  wire G641_o2_n;
  wire G1117_o2_p;
  wire G1117_o2_n;
  wire G1096_o2_p;
  wire G1096_o2_n;
  wire G1143_o2_p;
  wire G1143_o2_n;
  wire G1112_o2_p;
  wire G1112_o2_n;
  wire n1138_lo_buf_o2_p;
  wire n1138_lo_buf_o2_n;
  wire n1210_lo_buf_o2_p;
  wire n1210_lo_buf_o2_n;
  wire G687_o2_p;
  wire G687_o2_n;
  wire G541_o2_p;
  wire G541_o2_n;
  wire G802_o2_p;
  wire G802_o2_n;
  wire G813_o2_p;
  wire G813_o2_n;
  wire G810_o2_p;
  wire G810_o2_n;
  wire G987_o2_p;
  wire G987_o2_n;
  wire G898_o2_p;
  wire G898_o2_n;
  wire n946_lo_buf_o2_p;
  wire n946_lo_buf_o2_n;
  wire n1054_lo_buf_o2_p;
  wire n1054_lo_buf_o2_n;
  wire G728_o2_p;
  wire G728_o2_n;
  wire G856_o2_p;
  wire G856_o2_n;
  wire n949_1_inv_p;
  wire n949_1_inv_n;
  wire G942_o2_p;
  wire G942_o2_n;
  wire G1099_o2_p;
  wire G1099_o2_n;
  wire G1154_o2_p;
  wire G1154_o2_n;
  wire G1131_o2_p;
  wire G1131_o2_n;
  wire G1169_o2_p;
  wire G1169_o2_n;
  wire G134_o2_p;
  wire G134_o2_n;
  wire n970_inv_p;
  wire n970_inv_n;
  wire G470_o2_p;
  wire G470_o2_n;
  wire G344_o2_p;
  wire G344_o2_n;
  wire G362_o2_p;
  wire G362_o2_n;
  wire G482_o2_p;
  wire G482_o2_n;
  wire G660_o2_p;
  wire G660_o2_n;
  wire G672_o2_p;
  wire G672_o2_n;
  wire n1096_lo_buf_o2_p;
  wire n1096_lo_buf_o2_n;
  wire G479_o2_p;
  wire G479_o2_n;
  wire G669_o2_p;
  wire G669_o2_n;
  wire n994_lo_buf_o2_p;
  wire n994_lo_buf_o2_n;
  wire n1066_lo_buf_o2_p;
  wire n1066_lo_buf_o2_n;
  wire n1006_inv_p;
  wire n1006_inv_n;
  wire G147_o2_p;
  wire G147_o2_n;
  wire G473_o2_p;
  wire G473_o2_n;
  wire G488_o2_p;
  wire G488_o2_n;
  wire G589_o2_p;
  wire G589_o2_n;
  wire G663_o2_p;
  wire G663_o2_n;
  wire G684_o2_p;
  wire G684_o2_n;
  wire G605_o2_p;
  wire G605_o2_n;
  wire G774_o2_p;
  wire G774_o2_n;
  wire G782_o2_p;
  wire G782_o2_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire g686_p;
  wire g686_n;
  wire g687_p;
  wire g687_n;
  wire g688_p;
  wire g688_n;
  wire g689_p;
  wire g689_n;
  wire g690_p;
  wire g690_n;
  wire g691_p;
  wire g691_n;
  wire g692_p;
  wire g692_n;
  wire g693_p;
  wire g693_n;
  wire g694_p;
  wire g694_n;
  wire g695_p;
  wire g695_n;
  wire g696_p;
  wire g696_n;
  wire g697_p;
  wire g697_n;
  wire g698_p;
  wire g698_n;
  wire g699_p;
  wire g699_n;
  wire g700_p;
  wire g700_n;
  wire g701_p;
  wire g701_n;
  wire g702_p;
  wire g702_n;
  wire g703_p;
  wire g703_n;
  wire g704_p;
  wire g704_n;
  wire g705_p;
  wire g705_n;
  wire g706_p;
  wire g706_n;
  wire g707_p;
  wire g707_n;
  wire g708_p;
  wire g708_n;
  wire g709_p;
  wire g709_n;
  wire g710_p;
  wire g710_n;
  wire g711_p;
  wire g711_n;
  wire g712_p;
  wire g712_n;
  wire g713_p;
  wire g713_n;
  wire g714_p;
  wire g714_n;
  wire g715_p;
  wire g715_n;
  wire g716_p;
  wire g716_n;
  wire g717_p;
  wire g717_n;
  wire g718_p;
  wire g718_n;
  wire g719_p;
  wire g719_n;
  wire g720_p;
  wire g720_n;
  wire g721_p;
  wire g721_n;
  wire g722_p;
  wire g722_n;
  wire g723_p;
  wire g723_n;
  wire g724_p;
  wire g724_n;
  wire g725_p;
  wire g725_n;
  wire g726_p;
  wire g726_n;
  wire g727_p;
  wire g727_n;
  wire g728_p;
  wire g728_n;
  wire g729_p;
  wire g729_n;
  wire g730_p;
  wire g730_n;
  wire g731_p;
  wire g731_n;
  wire g732_p;
  wire g732_n;
  wire g733_p;
  wire g733_n;
  wire g734_p;
  wire g734_n;
  wire g735_p;
  wire g735_n;
  wire g736_p;
  wire g736_n;
  wire g737_p;
  wire g737_n;
  wire g738_p;
  wire g738_n;
  wire g739_p;
  wire g739_n;
  wire g740_p;
  wire g740_n;
  wire g741_p;
  wire g741_n;
  wire g742_p;
  wire g742_n;
  wire g743_p;
  wire g743_n;
  wire g744_p;
  wire g744_n;
  wire g745_p;
  wire g745_n;
  wire g746_p;
  wire g746_n;
  wire g747_p;
  wire g747_n;
  wire g748_p;
  wire g748_n;
  wire g749_p;
  wire g749_n;
  wire g750_p;
  wire g750_n;
  wire g751_p;
  wire g751_n;
  wire g752_p;
  wire g752_n;
  wire g753_p;
  wire g753_n;
  wire g754_p;
  wire g754_n;
  wire g755_p;
  wire g755_n;
  wire g756_p;
  wire g756_n;
  wire g757_p;
  wire g757_n;
  wire g758_p;
  wire g758_n;
  wire g759_p;
  wire g759_n;
  wire g760_p;
  wire g760_n;
  wire g761_p;
  wire g761_n;
  wire g762_p;
  wire g762_n;
  wire g763_p;
  wire g763_n;
  wire g764_p;
  wire g764_n;
  wire g765_p;
  wire g765_n;
  wire g766_p;
  wire g766_n;
  wire g767_p;
  wire g767_n;
  wire g768_p;
  wire g768_n;
  wire g769_p;
  wire g769_n;
  wire g770_p;
  wire g770_n;
  wire g771_p;
  wire g771_n;
  wire g772_p;
  wire g772_n;
  wire g773_p;
  wire g773_n;
  wire g774_p;
  wire g774_n;
  wire g775_p;
  wire g775_n;
  wire g776_p;
  wire g776_n;
  wire g777_p;
  wire g777_n;
  wire g778_p;
  wire g778_n;
  wire g779_p;
  wire g779_n;
  wire g780_p;
  wire g780_n;
  wire g781_p;
  wire g781_n;
  wire g782_p;
  wire g782_n;
  wire g783_p;
  wire g783_n;
  wire g784_p;
  wire g784_n;
  wire g785_p;
  wire g785_n;
  wire g786_p;
  wire g786_n;
  wire g787_p;
  wire g787_n;
  wire g788_p;
  wire g788_n;
  wire g789_p;
  wire g789_n;
  wire g790_p;
  wire g790_n;
  wire g791_p;
  wire g791_n;
  wire g792_p;
  wire g792_n;
  wire g793_p;
  wire g793_n;
  wire g794_p;
  wire g794_n;
  wire g795_p;
  wire g795_n;
  wire g796_p;
  wire g796_n;
  wire g797_p;
  wire g797_n;
  wire g798_p;
  wire g798_n;
  wire g799_p;
  wire g799_n;
  wire g800_p;
  wire g800_n;
  wire g801_p;
  wire g801_n;
  wire g802_p;
  wire g802_n;
  wire g803_p;
  wire g803_n;
  wire g804_p;
  wire g804_n;
  wire g805_p;
  wire g805_n;
  wire g806_p;
  wire g806_n;
  wire g807_p;
  wire g807_n;
  wire g808_p;
  wire g808_n;
  wire g809_p;
  wire g809_n;
  wire g810_p;
  wire g810_n;
  wire g811_p;
  wire g811_n;
  wire g812_p;
  wire g812_n;
  wire g813_p;
  wire g813_n;
  wire g814_p;
  wire g814_n;
  wire g815_p;
  wire g815_n;
  wire g816_p;
  wire g816_n;
  wire g817_p;
  wire g817_n;
  wire g818_p;
  wire g818_n;
  wire g819_p;
  wire g819_n;
  wire g820_p;
  wire g820_n;
  wire g821_p;
  wire g821_n;
  wire g822_p;
  wire g822_n;
  wire g823_p;
  wire g823_n;
  wire g824_p;
  wire g824_n;
  wire g825_p;
  wire g825_n;
  wire g826_p;
  wire g826_n;
  wire g827_p;
  wire g827_n;
  wire g828_p;
  wire g828_n;
  wire g829_p;
  wire g829_n;
  wire g830_p;
  wire g830_n;
  wire g831_p;
  wire g831_n;
  wire g832_p;
  wire g832_n;
  wire g833_p;
  wire g833_n;
  wire g834_p;
  wire g834_n;
  wire g835_p;
  wire g835_n;
  wire g836_p;
  wire g836_n;
  wire g837_p;
  wire g837_n;
  wire g838_p;
  wire g838_n;
  wire g839_p;
  wire g839_n;
  wire g840_p;
  wire g840_n;
  wire g841_p;
  wire g841_n;
  wire g842_p;
  wire g842_n;
  wire g843_p;
  wire g843_n;
  wire g844_p;
  wire g844_n;
  wire g845_p;
  wire g845_n;
  wire g846_p;
  wire g846_n;
  wire g847_p;
  wire g847_n;
  wire g848_p;
  wire g848_n;
  wire g849_p;
  wire g849_n;
  wire g850_p;
  wire g850_n;
  wire g851_p;
  wire g851_n;
  wire g852_p;
  wire g852_n;
  wire g853_p;
  wire g853_n;
  wire g854_p;
  wire g854_n;
  wire g855_p;
  wire g855_n;
  wire g856_p;
  wire g856_n;
  wire g857_p;
  wire g857_n;
  wire g858_p;
  wire g858_n;
  wire g859_p;
  wire g859_n;
  wire g860_p;
  wire g860_n;
  wire g861_p;
  wire g861_n;
  wire g862_p;
  wire g862_n;
  wire g863_p;
  wire g863_n;
  wire g864_p;
  wire g864_n;
  wire g865_p;
  wire g865_n;
  wire g866_p;
  wire g866_n;
  wire g867_p;
  wire g867_n;
  wire g868_p;
  wire g868_n;
  wire g869_p;
  wire g869_n;
  wire g870_p;
  wire g870_n;
  wire g871_p;
  wire g871_n;
  wire g872_p;
  wire g872_n;
  wire g873_p;
  wire g873_n;
  wire g874_p;
  wire g874_n;
  wire g875_p;
  wire g875_n;
  wire g876_p;
  wire g876_n;
  wire g877_p;
  wire g877_n;
  wire g878_p;
  wire g878_n;
  wire g879_p;
  wire g879_n;
  wire g880_p;
  wire g880_n;
  wire g881_p;
  wire g881_n;
  wire g882_p;
  wire g882_n;
  wire g883_p;
  wire g883_n;
  wire g884_p;
  wire g884_n;
  wire g885_p;
  wire g885_n;
  wire g886_p;
  wire g886_n;
  wire g887_p;
  wire g887_n;
  wire g888_p;
  wire g888_n;
  wire G1538_o2_n_spl_;
  wire G1511_o2_n_spl_;
  wire G1538_o2_p_spl_;
  wire G1511_o2_p_spl_;
  wire g359_p_spl_;
  wire g359_p_spl_0;
  wire G1584_o2_p_spl_;
  wire G1584_o2_p_spl_0;
  wire G1584_o2_p_spl_00;
  wire G1584_o2_p_spl_01;
  wire G1584_o2_p_spl_1;
  wire g359_n_spl_;
  wire g359_n_spl_0;
  wire G1584_o2_n_spl_;
  wire G1584_o2_n_spl_0;
  wire G1584_o2_n_spl_00;
  wire G1584_o2_n_spl_1;
  wire G1395_o2_n_spl_;
  wire G1395_o2_n_spl_0;
  wire G1395_o2_n_spl_00;
  wire G1395_o2_n_spl_000;
  wire G1395_o2_n_spl_001;
  wire G1395_o2_n_spl_01;
  wire G1395_o2_n_spl_1;
  wire G1395_o2_n_spl_10;
  wire G1395_o2_n_spl_11;
  wire G1395_o2_p_spl_;
  wire G1395_o2_p_spl_0;
  wire G1395_o2_p_spl_1;
  wire G738_o2_n_spl_;
  wire G738_o2_n_spl_0;
  wire G738_o2_n_spl_00;
  wire G738_o2_n_spl_01;
  wire G738_o2_n_spl_1;
  wire G738_o2_n_spl_10;
  wire G738_o2_n_spl_11;
  wire G738_o2_p_spl_;
  wire G738_o2_p_spl_0;
  wire G738_o2_p_spl_00;
  wire G738_o2_p_spl_01;
  wire G738_o2_p_spl_1;
  wire G738_o2_p_spl_10;
  wire G738_o2_p_spl_11;
  wire G1563_o2_p_spl_;
  wire G1563_o2_p_spl_0;
  wire G1563_o2_p_spl_00;
  wire G1563_o2_p_spl_01;
  wire G1563_o2_p_spl_1;
  wire G1563_o2_n_spl_;
  wire g366_p_spl_;
  wire G1420_o2_n_spl_;
  wire G1420_o2_n_spl_0;
  wire G1420_o2_n_spl_00;
  wire G1420_o2_n_spl_01;
  wire G1420_o2_n_spl_1;
  wire G1420_o2_n_spl_10;
  wire g366_n_spl_;
  wire G1420_o2_p_spl_;
  wire G1420_o2_p_spl_0;
  wire G1420_o2_p_spl_00;
  wire G1420_o2_p_spl_01;
  wire G1420_o2_p_spl_1;
  wire G1410_o2_n_spl_;
  wire G1410_o2_n_spl_0;
  wire G1410_o2_n_spl_00;
  wire G1410_o2_n_spl_1;
  wire G1410_o2_p_spl_;
  wire G1410_o2_p_spl_0;
  wire G1410_o2_p_spl_1;
  wire G1576_o2_p_spl_;
  wire G1576_o2_p_spl_0;
  wire G1576_o2_p_spl_1;
  wire G1576_o2_n_spl_;
  wire G1576_o2_n_spl_0;
  wire G1522_o2_n_spl_;
  wire G1522_o2_n_spl_0;
  wire G1522_o2_p_spl_;
  wire G1522_o2_p_spl_0;
  wire G1598_o2_p_spl_;
  wire G1598_o2_p_spl_0;
  wire G1598_o2_p_spl_1;
  wire G1598_o2_n_spl_;
  wire G1598_o2_n_spl_0;
  wire G1598_o2_n_spl_1;
  wire G755_o2_n_spl_;
  wire G755_o2_n_spl_0;
  wire G755_o2_n_spl_00;
  wire G755_o2_n_spl_01;
  wire G755_o2_n_spl_1;
  wire G755_o2_n_spl_10;
  wire G755_o2_n_spl_11;
  wire G755_o2_p_spl_;
  wire G755_o2_p_spl_0;
  wire G755_o2_p_spl_00;
  wire G755_o2_p_spl_01;
  wire G755_o2_p_spl_1;
  wire G755_o2_p_spl_10;
  wire G755_o2_p_spl_11;
  wire G1549_o2_n_spl_;
  wire G1549_o2_p_spl_;
  wire g390_p_spl_;
  wire g390_n_spl_;
  wire G1434_o2_n_spl_;
  wire G1434_o2_p_spl_;
  wire G1625_o2_p_spl_;
  wire G1625_o2_p_spl_0;
  wire G1625_o2_p_spl_1;
  wire G1625_o2_n_spl_;
  wire g410_p_spl_;
  wire g410_p_spl_0;
  wire g410_p_spl_1;
  wire g410_n_spl_;
  wire g410_n_spl_0;
  wire g410_n_spl_1;
  wire g423_p_spl_;
  wire G1609_o2_p_spl_;
  wire G1609_o2_p_spl_0;
  wire g435_p_spl_;
  wire g435_p_spl_0;
  wire g435_p_spl_1;
  wire g435_n_spl_;
  wire g435_n_spl_0;
  wire g436_p_spl_;
  wire g436_n_spl_;
  wire g484_n_spl_;
  wire n1321_lo_p_spl_;
  wire n1321_lo_p_spl_0;
  wire g488_p_spl_;
  wire g488_p_spl_0;
  wire g488_p_spl_00;
  wire g488_p_spl_01;
  wire g488_p_spl_1;
  wire g488_p_spl_10;
  wire g488_p_spl_11;
  wire g494_p_spl_;
  wire g494_p_spl_0;
  wire g498_p_spl_;
  wire g523_n_spl_;
  wire g523_n_spl_0;
  wire g523_n_spl_00;
  wire g523_n_spl_01;
  wire g523_n_spl_1;
  wire g523_n_spl_10;
  wire g530_n_spl_;
  wire n2372_o2_n_spl_;
  wire g530_p_spl_;
  wire n2372_o2_p_spl_;
  wire n1309_lo_n_spl_;
  wire n1309_lo_n_spl_0;
  wire n1309_lo_n_spl_00;
  wire n1309_lo_n_spl_01;
  wire n1309_lo_n_spl_1;
  wire n1309_lo_p_spl_;
  wire n1309_lo_p_spl_0;
  wire n1309_lo_p_spl_00;
  wire n1309_lo_p_spl_01;
  wire n1309_lo_p_spl_1;
  wire g523_p_spl_;
  wire g523_p_spl_0;
  wire g523_p_spl_00;
  wire g523_p_spl_01;
  wire g523_p_spl_1;
  wire n1333_lo_p_spl_;
  wire n1333_lo_p_spl_0;
  wire n1333_lo_p_spl_00;
  wire n1333_lo_p_spl_1;
  wire g540_n_spl_;
  wire g540_n_spl_0;
  wire g540_n_spl_00;
  wire g540_n_spl_01;
  wire g540_n_spl_1;
  wire g545_p_spl_;
  wire g542_p_spl_;
  wire g545_n_spl_;
  wire g542_n_spl_;
  wire n1333_lo_n_spl_;
  wire n1333_lo_n_spl_0;
  wire n1333_lo_n_spl_1;
  wire G248_o2_n_spl_;
  wire G248_o2_p_spl_;
  wire g584_n_spl_;
  wire g581_p_spl_;
  wire g584_p_spl_;
  wire g581_n_spl_;
  wire g603_n_spl_;
  wire g600_p_spl_;
  wire g603_p_spl_;
  wire g600_n_spl_;
  wire g616_n_spl_;
  wire g614_n_spl_;
  wire g616_p_spl_;
  wire g614_p_spl_;
  wire n2180_o2_p_spl_;
  wire n1874_o2_p_spl_;
  wire n2180_o2_n_spl_;
  wire n1874_o2_n_spl_;
  wire G391_o2_p_spl_;
  wire G391_o2_p_spl_0;
  wire n2724_o2_p_spl_;
  wire G391_o2_n_spl_;
  wire G387_o2_p_spl_;
  wire G387_o2_p_spl_0;
  wire n1162_lo_buf_o2_p_spl_;
  wire G387_o2_n_spl_;
  wire G1140_o2_p_spl_;
  wire G212_o2_n_spl_;
  wire G212_o2_n_spl_0;
  wire G212_o2_n_spl_00;
  wire G212_o2_n_spl_01;
  wire G212_o2_n_spl_1;
  wire G212_o2_p_spl_;
  wire G212_o2_p_spl_0;
  wire G212_o2_p_spl_00;
  wire G212_o2_p_spl_01;
  wire G212_o2_p_spl_1;
  wire G1178_o2_p_spl_;
  wire n820_inv_p_spl_;
  wire n1138_lo_buf_o2_p_spl_;
  wire G241_o2_n_spl_;
  wire G241_o2_n_spl_0;
  wire G241_o2_n_spl_1;
  wire G241_o2_p_spl_;
  wire G241_o2_p_spl_0;
  wire G241_o2_p_spl_1;
  wire n1195_lo_buf_o2_p_spl_;
  wire g633_n_spl_;
  wire g627_p_spl_;
  wire n1234_lo_buf_o2_p_spl_;
  wire n1234_lo_buf_o2_p_spl_0;
  wire g634_p_spl_;
  wire g643_p_spl_;
  wire g643_p_spl_0;
  wire g635_p_spl_;
  wire g646_p_spl_;
  wire g646_p_spl_0;
  wire g636_p_spl_;
  wire n1306_lo_buf_o2_n_spl_;
  wire n2498_o2_n_spl_;
  wire n2498_o2_n_spl_0;
  wire g637_n_spl_;
  wire g637_n_spl_0;
  wire g637_n_spl_1;
  wire g653_p_spl_;
  wire g631_n_spl_;
  wire g628_p_spl_;
  wire g632_n_spl_;
  wire n1246_lo_buf_o2_p_spl_;
  wire n1246_lo_buf_o2_p_spl_0;
  wire n1270_lo_buf_o2_p_spl_;
  wire n1270_lo_buf_o2_p_spl_0;
  wire g629_p_spl_;
  wire n1258_lo_buf_o2_p_spl_;
  wire n1258_lo_buf_o2_p_spl_0;
  wire g630_p_spl_;
  wire g675_n_spl_;
  wire n949_1_inv_n_spl_;
  wire g675_p_spl_;
  wire n949_1_inv_p_spl_;
  wire n949_1_inv_p_spl_0;
  wire g660_n_spl_;
  wire g660_n_spl_0;
  wire g660_n_spl_1;
  wire g647_p_spl_;
  wire g667_p_spl_;
  wire g667_p_spl_0;
  wire g667_p_spl_00;
  wire g667_p_spl_01;
  wire g667_p_spl_1;
  wire g667_p_spl_10;
  wire g674_p_spl_;
  wire g674_p_spl_0;
  wire g674_p_spl_00;
  wire g674_p_spl_01;
  wire g674_p_spl_1;
  wire g674_p_spl_10;
  wire g658_n_spl_;
  wire g658_n_spl_0;
  wire g658_n_spl_1;
  wire g659_n_spl_;
  wire g659_n_spl_0;
  wire g659_n_spl_1;
  wire g648_p_spl_;
  wire g694_p_spl_;
  wire g654_n_spl_;
  wire g654_n_spl_0;
  wire g699_p_spl_;
  wire G669_o2_p_spl_;
  wire G479_o2_p_spl_;
  wire G669_o2_n_spl_;
  wire G479_o2_n_spl_;
  wire G147_o2_p_spl_;
  wire G147_o2_p_spl_0;
  wire G147_o2_p_spl_1;
  wire G147_o2_n_spl_;
  wire G147_o2_n_spl_0;
  wire G147_o2_n_spl_1;
  wire G663_o2_p_spl_;
  wire G473_o2_p_spl_;
  wire G663_o2_n_spl_;
  wire G473_o2_n_spl_;
  wire n994_lo_buf_o2_p_spl_;
  wire n994_lo_buf_o2_p_spl_0;
  wire n994_lo_buf_o2_p_spl_1;
  wire n994_lo_buf_o2_n_spl_;
  wire n1006_inv_p_spl_;
  wire n1006_inv_p_spl_0;
  wire n1006_inv_n_spl_;
  wire g728_n_spl_;
  wire n2737_o2_n_spl_;
  wire g732_n_spl_;
  wire G365_o2_p_spl_;
  wire g736_n_spl_;
  wire n2428_o2_p_spl_;
  wire g736_p_spl_;
  wire n2428_o2_n_spl_;
  wire g745_n_spl_;
  wire g742_n_spl_;
  wire g701_p_spl_;
  wire g701_p_spl_0;
  wire g701_p_spl_00;
  wire g701_p_spl_01;
  wire g701_p_spl_1;
  wire g696_p_spl_;
  wire g691_p_spl_;
  wire g691_p_spl_0;
  wire g691_p_spl_00;
  wire g691_p_spl_01;
  wire g691_p_spl_1;
  wire g691_p_spl_10;
  wire g691_p_spl_11;
  wire g700_p_spl_;
  wire g700_p_spl_0;
  wire g700_p_spl_00;
  wire g700_p_spl_1;
  wire g695_p_spl_;
  wire g695_p_spl_0;
  wire g695_p_spl_00;
  wire g695_p_spl_01;
  wire g695_p_spl_1;
  wire g695_p_spl_10;
  wire g695_p_spl_11;
  wire G338_o2_p_spl_;
  wire n853_inv_p_spl_;
  wire n853_inv_p_spl_0;
  wire G338_o2_n_spl_;
  wire n853_inv_n_spl_;
  wire G684_o2_p_spl_;
  wire G488_o2_p_spl_;
  wire G684_o2_n_spl_;
  wire G488_o2_n_spl_;
  wire n1066_lo_buf_o2_p_spl_;
  wire n1066_lo_buf_o2_p_spl_0;
  wire n1066_lo_buf_o2_p_spl_1;
  wire n2747_o2_p_spl_;
  wire n2744_o2_p_spl_;
  wire n2744_o2_p_spl_0;
  wire n2744_o2_p_spl_1;
  wire n1222_lo_buf_o2_p_spl_;
  wire n1303_lo_p_spl_;
  wire n1303_lo_p_spl_0;
  wire n1303_lo_p_spl_1;
  wire n1210_lo_buf_o2_p_spl_;
  wire n1210_lo_buf_o2_p_spl_0;
  wire n1210_lo_buf_o2_p_spl_1;
  wire G810_o2_p_spl_;
  wire G419_o2_n_spl_;
  wire G810_o2_n_spl_;
  wire G419_o2_p_spl_;
  wire G813_o2_p_spl_;
  wire G425_o2_n_spl_;
  wire G813_o2_n_spl_;
  wire G425_o2_p_spl_;
  wire g780_p_spl_;
  wire g777_n_spl_;
  wire g780_n_spl_;
  wire g777_p_spl_;
  wire n1210_lo_buf_o2_n_spl_;
  wire n1159_lo_p_spl_;
  wire G898_o2_n_spl_;
  wire G641_o2_p_spl_;
  wire G898_o2_p_spl_;
  wire G641_o2_n_spl_;
  wire G802_o2_p_spl_;
  wire G416_o2_n_spl_;
  wire G802_o2_n_spl_;
  wire G416_o2_p_spl_;
  wire g794_p_spl_;
  wire g791_n_spl_;
  wire g794_n_spl_;
  wire g791_p_spl_;
  wire G500_o2_p_spl_;
  wire G497_o2_n_spl_;
  wire G500_o2_n_spl_;
  wire G497_o2_p_spl_;
  wire g800_n_spl_;
  wire n2652_o2_n_spl_;
  wire g800_p_spl_;
  wire n2652_o2_p_spl_;
  wire G687_o2_p_spl_;
  wire G491_o2_p_spl_;
  wire G687_o2_n_spl_;
  wire G491_o2_n_spl_;
  wire g809_n_spl_;
  wire g640_p_spl_;
  wire g640_p_spl_0;
  wire g809_p_spl_;
  wire g640_n_spl_;
  wire g815_n_spl_;
  wire n748_inv_p_spl_;
  wire n748_inv_p_spl_0;
  wire n748_inv_p_spl_1;
  wire g815_p_spl_;
  wire n748_inv_n_spl_;
  wire g827_n_spl_;
  wire g824_p_spl_;
  wire g827_p_spl_;
  wire g824_n_spl_;
  wire n1171_lo_buf_o2_p_spl_;
  wire g832_p_spl_;
  wire n2744_o2_n_spl_;
  wire g832_n_spl_;
  wire g639_p_spl_;
  wire g639_p_spl_0;
  wire n511_inv_p_spl_;
  wire n511_inv_p_spl_0;
  wire g639_n_spl_;
  wire n511_inv_n_spl_;
  wire g844_n_spl_;
  wire G987_o2_n_spl_;
  wire g844_p_spl_;
  wire G987_o2_p_spl_;
  wire G987_o2_p_spl_0;
  wire G134_o2_n_spl_;
  wire G134_o2_n_spl_0;
  wire G134_o2_p_spl_;
  wire G134_o2_p_spl_0;
  wire g854_n_spl_;
  wire G353_o2_p_spl_;
  wire G353_o2_p_spl_0;
  wire g854_p_spl_;
  wire G353_o2_n_spl_;
  wire g678_p_spl_;
  wire n1036_lo_n_spl_;
  wire n1036_lo_n_spl_0;
  wire n1096_lo_buf_o2_p_spl_;
  wire n1096_lo_buf_o2_p_spl_0;
  wire n1096_lo_buf_o2_p_spl_00;
  wire n1096_lo_buf_o2_p_spl_1;
  wire n1036_lo_p_spl_;
  wire n1036_lo_p_spl_0;
  wire n1036_lo_p_spl_1;
  wire n1324_lo_n_spl_;
  wire n1180_lo_p_spl_;
  wire g707_n_spl_;
  wire g707_n_spl_0;
  wire g707_n_spl_00;
  wire g707_n_spl_01;
  wire g707_n_spl_1;
  wire g719_n_spl_;
  wire g719_n_spl_0;
  wire g713_n_spl_;
  wire g713_n_spl_0;
  wire n1144_lo_p_spl_;
  wire n1216_lo_p_spl_;
  wire n1216_lo_p_spl_0;
  wire n1324_lo_p_spl_;
  wire n1324_lo_p_spl_0;
  wire G165_o2_p_spl_;
  wire G165_o2_n_spl_;
  wire n1024_lo_p_spl_;
  wire n1024_lo_p_spl_0;
  wire n1024_lo_p_spl_1;
  wire n1024_lo_n_spl_;
  wire G344_o2_p_spl_;
  wire G344_o2_n_spl_;
  wire n976_lo_p_spl_;
  wire n976_lo_p_spl_0;
  wire n976_lo_p_spl_00;
  wire n976_lo_p_spl_01;
  wire n976_lo_p_spl_1;
  wire n1282_lo_p_spl_;
  wire n1294_lo_p_spl_;
  wire n1318_lo_p_spl_;
  wire n2498_o2_p_spl_;
  wire n2498_o2_p_spl_0;
  wire n2716_o2_p_spl_;
  wire G1059_o2_p_spl_;
  wire n460_inv_p_spl_;
  wire g681_n_spl_;
  wire g684_n_spl_;
  wire g687_n_spl_;
  wire g725_n_spl_;
  wire g725_n_spl_0;
  wire g725_n_spl_1;
  wire G2_p_spl_;
  wire G2_p_spl_0;
  wire G2_p_spl_00;
  wire G2_p_spl_1;
  wire G15_p_spl_;
  wire G15_p_spl_0;
  wire G15_p_spl_00;
  wire G15_p_spl_1;
  wire g764_n_spl_;
  wire g764_n_spl_0;
  wire g770_n_spl_;
  wire g770_n_spl_0;
  wire G3_p_spl_;
  wire G3_p_spl_0;
  wire G3_p_spl_1;
  wire G6_p_spl_;
  wire G6_p_spl_0;
  wire G6_p_spl_1;
  wire G12_p_spl_;
  wire G12_p_spl_0;
  wire G12_p_spl_1;
  wire G16_p_spl_;
  wire G16_p_spl_0;
  wire G16_p_spl_00;
  wire G16_p_spl_1;
  wire n862_inv_p_spl_;
  wire n862_inv_p_spl_0;
  wire g853_n_spl_;
  wire g863_p_spl_;
  wire g863_p_spl_0;
  wire G7_p_spl_;
  wire G7_p_spl_0;
  wire G13_p_spl_;
  wire G13_p_spl_0;
  wire G1_p_spl_;
  wire G10_p_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    n949_lo_p,
    n949_lo
  );


  not

  (
    n949_lo_n,
    n949_lo
  );


  buf

  (
    n961_lo_p,
    n961_lo
  );


  not

  (
    n961_lo_n,
    n961_lo
  );


  buf

  (
    n973_lo_p,
    n973_lo
  );


  not

  (
    n973_lo_n,
    n973_lo
  );


  buf

  (
    n976_lo_p,
    n976_lo
  );


  not

  (
    n976_lo_n,
    n976_lo
  );


  buf

  (
    n985_lo_p,
    n985_lo
  );


  not

  (
    n985_lo_n,
    n985_lo
  );


  buf

  (
    n997_lo_p,
    n997_lo
  );


  not

  (
    n997_lo_n,
    n997_lo
  );


  buf

  (
    n1009_lo_p,
    n1009_lo
  );


  not

  (
    n1009_lo_n,
    n1009_lo
  );


  buf

  (
    n1021_lo_p,
    n1021_lo
  );


  not

  (
    n1021_lo_n,
    n1021_lo
  );


  buf

  (
    n1024_lo_p,
    n1024_lo
  );


  not

  (
    n1024_lo_n,
    n1024_lo
  );


  buf

  (
    n1033_lo_p,
    n1033_lo
  );


  not

  (
    n1033_lo_n,
    n1033_lo
  );


  buf

  (
    n1036_lo_p,
    n1036_lo
  );


  not

  (
    n1036_lo_n,
    n1036_lo
  );


  buf

  (
    n1045_lo_p,
    n1045_lo
  );


  not

  (
    n1045_lo_n,
    n1045_lo
  );


  buf

  (
    n1057_lo_p,
    n1057_lo
  );


  not

  (
    n1057_lo_n,
    n1057_lo
  );


  buf

  (
    n1069_lo_p,
    n1069_lo
  );


  not

  (
    n1069_lo_n,
    n1069_lo
  );


  buf

  (
    n1081_lo_p,
    n1081_lo
  );


  not

  (
    n1081_lo_n,
    n1081_lo
  );


  buf

  (
    n1093_lo_p,
    n1093_lo
  );


  not

  (
    n1093_lo_n,
    n1093_lo
  );


  buf

  (
    n1105_lo_p,
    n1105_lo
  );


  not

  (
    n1105_lo_n,
    n1105_lo
  );


  buf

  (
    n1117_lo_p,
    n1117_lo
  );


  not

  (
    n1117_lo_n,
    n1117_lo
  );


  buf

  (
    n1129_lo_p,
    n1129_lo
  );


  not

  (
    n1129_lo_n,
    n1129_lo
  );


  buf

  (
    n1132_lo_p,
    n1132_lo
  );


  not

  (
    n1132_lo_n,
    n1132_lo
  );


  buf

  (
    n1141_lo_p,
    n1141_lo
  );


  not

  (
    n1141_lo_n,
    n1141_lo
  );


  buf

  (
    n1144_lo_p,
    n1144_lo
  );


  not

  (
    n1144_lo_n,
    n1144_lo
  );


  buf

  (
    n1156_lo_p,
    n1156_lo
  );


  not

  (
    n1156_lo_n,
    n1156_lo
  );


  buf

  (
    n1159_lo_p,
    n1159_lo
  );


  not

  (
    n1159_lo_n,
    n1159_lo
  );


  buf

  (
    n1165_lo_p,
    n1165_lo
  );


  not

  (
    n1165_lo_n,
    n1165_lo
  );


  buf

  (
    n1168_lo_p,
    n1168_lo
  );


  not

  (
    n1168_lo_n,
    n1168_lo
  );


  buf

  (
    n1180_lo_p,
    n1180_lo
  );


  not

  (
    n1180_lo_n,
    n1180_lo
  );


  buf

  (
    n1189_lo_p,
    n1189_lo
  );


  not

  (
    n1189_lo_n,
    n1189_lo
  );


  buf

  (
    n1192_lo_p,
    n1192_lo
  );


  not

  (
    n1192_lo_n,
    n1192_lo
  );


  buf

  (
    n1201_lo_p,
    n1201_lo
  );


  not

  (
    n1201_lo_n,
    n1201_lo
  );


  buf

  (
    n1204_lo_p,
    n1204_lo
  );


  not

  (
    n1204_lo_n,
    n1204_lo
  );


  buf

  (
    n1216_lo_p,
    n1216_lo
  );


  not

  (
    n1216_lo_n,
    n1216_lo
  );


  buf

  (
    n1228_lo_p,
    n1228_lo
  );


  not

  (
    n1228_lo_n,
    n1228_lo
  );


  buf

  (
    n1231_lo_p,
    n1231_lo
  );


  not

  (
    n1231_lo_n,
    n1231_lo
  );


  buf

  (
    n1237_lo_p,
    n1237_lo
  );


  not

  (
    n1237_lo_n,
    n1237_lo
  );


  buf

  (
    n1240_lo_p,
    n1240_lo
  );


  not

  (
    n1240_lo_n,
    n1240_lo
  );


  buf

  (
    n1243_lo_p,
    n1243_lo
  );


  not

  (
    n1243_lo_n,
    n1243_lo
  );


  buf

  (
    n1249_lo_p,
    n1249_lo
  );


  not

  (
    n1249_lo_n,
    n1249_lo
  );


  buf

  (
    n1252_lo_p,
    n1252_lo
  );


  not

  (
    n1252_lo_n,
    n1252_lo
  );


  buf

  (
    n1255_lo_p,
    n1255_lo
  );


  not

  (
    n1255_lo_n,
    n1255_lo
  );


  buf

  (
    n1261_lo_p,
    n1261_lo
  );


  not

  (
    n1261_lo_n,
    n1261_lo
  );


  buf

  (
    n1264_lo_p,
    n1264_lo
  );


  not

  (
    n1264_lo_n,
    n1264_lo
  );


  buf

  (
    n1267_lo_p,
    n1267_lo
  );


  not

  (
    n1267_lo_n,
    n1267_lo
  );


  buf

  (
    n1273_lo_p,
    n1273_lo
  );


  not

  (
    n1273_lo_n,
    n1273_lo
  );


  buf

  (
    n1276_lo_p,
    n1276_lo
  );


  not

  (
    n1276_lo_n,
    n1276_lo
  );


  buf

  (
    n1279_lo_p,
    n1279_lo
  );


  not

  (
    n1279_lo_n,
    n1279_lo
  );


  buf

  (
    n1282_lo_p,
    n1282_lo
  );


  not

  (
    n1282_lo_n,
    n1282_lo
  );


  buf

  (
    n1285_lo_p,
    n1285_lo
  );


  not

  (
    n1285_lo_n,
    n1285_lo
  );


  buf

  (
    n1288_lo_p,
    n1288_lo
  );


  not

  (
    n1288_lo_n,
    n1288_lo
  );


  buf

  (
    n1291_lo_p,
    n1291_lo
  );


  not

  (
    n1291_lo_n,
    n1291_lo
  );


  buf

  (
    n1294_lo_p,
    n1294_lo
  );


  not

  (
    n1294_lo_n,
    n1294_lo
  );


  buf

  (
    n1297_lo_p,
    n1297_lo
  );


  not

  (
    n1297_lo_n,
    n1297_lo
  );


  buf

  (
    n1300_lo_p,
    n1300_lo
  );


  not

  (
    n1300_lo_n,
    n1300_lo
  );


  buf

  (
    n1303_lo_p,
    n1303_lo
  );


  not

  (
    n1303_lo_n,
    n1303_lo
  );


  buf

  (
    n1309_lo_p,
    n1309_lo
  );


  not

  (
    n1309_lo_n,
    n1309_lo
  );


  buf

  (
    n1312_lo_p,
    n1312_lo
  );


  not

  (
    n1312_lo_n,
    n1312_lo
  );


  buf

  (
    n1315_lo_p,
    n1315_lo
  );


  not

  (
    n1315_lo_n,
    n1315_lo
  );


  buf

  (
    n1318_lo_p,
    n1318_lo
  );


  not

  (
    n1318_lo_n,
    n1318_lo
  );


  buf

  (
    n1321_lo_p,
    n1321_lo
  );


  not

  (
    n1321_lo_n,
    n1321_lo
  );


  buf

  (
    n1324_lo_p,
    n1324_lo
  );


  not

  (
    n1324_lo_n,
    n1324_lo
  );


  buf

  (
    n1333_lo_p,
    n1333_lo
  );


  not

  (
    n1333_lo_n,
    n1333_lo
  );


  buf

  (
    n1874_o2_p,
    n1874_o2
  );


  not

  (
    n1874_o2_n,
    n1874_o2
  );


  buf

  (
    n2180_o2_p,
    n2180_o2
  );


  not

  (
    n2180_o2_n,
    n2180_o2
  );


  buf

  (
    n2372_o2_p,
    n2372_o2
  );


  not

  (
    n2372_o2_n,
    n2372_o2
  );


  buf

  (
    n2190_o2_p,
    n2190_o2
  );


  not

  (
    n2190_o2_n,
    n2190_o2
  );


  buf

  (
    n2191_o2_p,
    n2191_o2
  );


  not

  (
    n2191_o2_n,
    n2191_o2
  );


  buf

  (
    n2212_o2_p,
    n2212_o2
  );


  not

  (
    n2212_o2_n,
    n2212_o2
  );


  buf

  (
    n2213_o2_p,
    n2213_o2
  );


  not

  (
    n2213_o2_n,
    n2213_o2
  );


  buf

  (
    n2214_o2_p,
    n2214_o2
  );


  not

  (
    n2214_o2_n,
    n2214_o2
  );


  buf

  (
    n2215_o2_p,
    n2215_o2
  );


  not

  (
    n2215_o2_n,
    n2215_o2
  );


  buf

  (
    n2275_o2_p,
    n2275_o2
  );


  not

  (
    n2275_o2_n,
    n2275_o2
  );


  buf

  (
    n2276_o2_p,
    n2276_o2
  );


  not

  (
    n2276_o2_n,
    n2276_o2
  );


  buf

  (
    n2290_o2_p,
    n2290_o2
  );


  not

  (
    n2290_o2_n,
    n2290_o2
  );


  buf

  (
    n2291_o2_p,
    n2291_o2
  );


  not

  (
    n2291_o2_n,
    n2291_o2
  );


  buf

  (
    n2681_o2_p,
    n2681_o2
  );


  not

  (
    n2681_o2_n,
    n2681_o2
  );


  buf

  (
    n2680_o2_p,
    n2680_o2
  );


  not

  (
    n2680_o2_n,
    n2680_o2
  );


  buf

  (
    n2683_o2_p,
    n2683_o2
  );


  not

  (
    n2683_o2_n,
    n2683_o2
  );


  buf

  (
    n2684_o2_p,
    n2684_o2
  );


  not

  (
    n2684_o2_n,
    n2684_o2
  );


  buf

  (
    n2686_o2_p,
    n2686_o2
  );


  not

  (
    n2686_o2_n,
    n2686_o2
  );


  buf

  (
    n2319_o2_p,
    n2319_o2
  );


  not

  (
    n2319_o2_n,
    n2319_o2
  );


  buf

  (
    n2320_o2_p,
    n2320_o2
  );


  not

  (
    n2320_o2_n,
    n2320_o2
  );


  buf

  (
    n304_inv_p,
    n304_inv
  );


  not

  (
    n304_inv_n,
    n304_inv
  );


  buf

  (
    G554_o2_p,
    G554_o2
  );


  not

  (
    G554_o2_n,
    G554_o2
  );


  buf

  (
    G557_o2_p,
    G557_o2
  );


  not

  (
    G557_o2_n,
    G557_o2
  );


  buf

  (
    G185_o2_p,
    G185_o2
  );


  not

  (
    G185_o2_n,
    G185_o2
  );


  buf

  (
    G188_o2_p,
    G188_o2
  );


  not

  (
    G188_o2_n,
    G188_o2
  );


  buf

  (
    G191_o2_p,
    G191_o2
  );


  not

  (
    G191_o2_n,
    G191_o2
  );


  buf

  (
    G194_o2_p,
    G194_o2
  );


  not

  (
    G194_o2_n,
    G194_o2
  );


  buf

  (
    G1182_o2_p,
    G1182_o2
  );


  not

  (
    G1182_o2_n,
    G1182_o2
  );


  buf

  (
    G1222_o2_p,
    G1222_o2
  );


  not

  (
    G1222_o2_n,
    G1222_o2
  );


  buf

  (
    G1247_o2_p,
    G1247_o2
  );


  not

  (
    G1247_o2_n,
    G1247_o2
  );


  buf

  (
    G1371_o2_p,
    G1371_o2
  );


  not

  (
    G1371_o2_n,
    G1371_o2
  );


  buf

  (
    G1383_o2_p,
    G1383_o2
  );


  not

  (
    G1383_o2_n,
    G1383_o2
  );


  buf

  (
    G1386_o2_p,
    G1386_o2
  );


  not

  (
    G1386_o2_n,
    G1386_o2
  );


  buf

  (
    n2416_o2_p,
    n2416_o2
  );


  not

  (
    n2416_o2_n,
    n2416_o2
  );


  buf

  (
    n2428_o2_p,
    n2428_o2
  );


  not

  (
    n2428_o2_n,
    n2428_o2
  );


  buf

  (
    n2438_o2_p,
    n2438_o2
  );


  not

  (
    n2438_o2_n,
    n2438_o2
  );


  buf

  (
    n2439_o2_p,
    n2439_o2
  );


  not

  (
    n2439_o2_n,
    n2439_o2
  );


  buf

  (
    n2440_o2_p,
    n2440_o2
  );


  not

  (
    n2440_o2_n,
    n2440_o2
  );


  buf

  (
    n2444_o2_p,
    n2444_o2
  );


  not

  (
    n2444_o2_n,
    n2444_o2
  );


  buf

  (
    n2497_o2_p,
    n2497_o2
  );


  not

  (
    n2497_o2_n,
    n2497_o2
  );


  buf

  (
    n2498_o2_p,
    n2498_o2
  );


  not

  (
    n2498_o2_n,
    n2498_o2
  );


  buf

  (
    n2503_o2_p,
    n2503_o2
  );


  not

  (
    n2503_o2_n,
    n2503_o2
  );


  buf

  (
    n2505_o2_p,
    n2505_o2
  );


  not

  (
    n2505_o2_n,
    n2505_o2
  );


  buf

  (
    n2529_o2_p,
    n2529_o2
  );


  not

  (
    n2529_o2_n,
    n2529_o2
  );


  buf

  (
    n2562_o2_p,
    n2562_o2
  );


  not

  (
    n2562_o2_n,
    n2562_o2
  );


  buf

  (
    n2570_o2_p,
    n2570_o2
  );


  not

  (
    n2570_o2_n,
    n2570_o2
  );


  buf

  (
    n2571_o2_p,
    n2571_o2
  );


  not

  (
    n2571_o2_n,
    n2571_o2
  );


  buf

  (
    n2574_o2_p,
    n2574_o2
  );


  not

  (
    n2574_o2_n,
    n2574_o2
  );


  buf

  (
    n2575_o2_p,
    n2575_o2
  );


  not

  (
    n2575_o2_n,
    n2575_o2
  );


  buf

  (
    G546_o2_p,
    G546_o2
  );


  not

  (
    G546_o2_n,
    G546_o2
  );


  buf

  (
    G550_o2_p,
    G550_o2
  );


  not

  (
    G550_o2_n,
    G550_o2
  );


  buf

  (
    n2633_o2_p,
    n2633_o2
  );


  not

  (
    n2633_o2_n,
    n2633_o2
  );


  buf

  (
    n2639_o2_p,
    n2639_o2
  );


  not

  (
    n2639_o2_n,
    n2639_o2
  );


  buf

  (
    n2642_o2_p,
    n2642_o2
  );


  not

  (
    n2642_o2_n,
    n2642_o2
  );


  buf

  (
    n2645_o2_p,
    n2645_o2
  );


  not

  (
    n2645_o2_n,
    n2645_o2
  );


  buf

  (
    n2679_o2_p,
    n2679_o2
  );


  not

  (
    n2679_o2_n,
    n2679_o2
  );


  buf

  (
    n2662_o2_p,
    n2662_o2
  );


  not

  (
    n2662_o2_n,
    n2662_o2
  );


  buf

  (
    n2724_o2_p,
    n2724_o2
  );


  not

  (
    n2724_o2_n,
    n2724_o2
  );


  buf

  (
    G382_o2_p,
    G382_o2
  );


  not

  (
    G382_o2_n,
    G382_o2
  );


  buf

  (
    G199_o2_p,
    G199_o2
  );


  not

  (
    G199_o2_n,
    G199_o2
  );


  buf

  (
    G202_o2_p,
    G202_o2
  );


  not

  (
    G202_o2_n,
    G202_o2
  );


  buf

  (
    G225_o2_p,
    G225_o2
  );


  not

  (
    G225_o2_n,
    G225_o2
  );


  buf

  (
    G248_o2_p,
    G248_o2
  );


  not

  (
    G248_o2_n,
    G248_o2
  );


  buf

  (
    G260_o2_p,
    G260_o2
  );


  not

  (
    G260_o2_n,
    G260_o2
  );


  buf

  (
    n2716_o2_p,
    n2716_o2
  );


  not

  (
    n2716_o2_n,
    n2716_o2
  );


  buf

  (
    n2737_o2_p,
    n2737_o2
  );


  not

  (
    n2737_o2_n,
    n2737_o2
  );


  buf

  (
    n1174_lo_buf_o2_p,
    n1174_lo_buf_o2
  );


  not

  (
    n1174_lo_buf_o2_n,
    n1174_lo_buf_o2
  );


  buf

  (
    n1198_lo_buf_o2_p,
    n1198_lo_buf_o2
  );


  not

  (
    n1198_lo_buf_o2_n,
    n1198_lo_buf_o2
  );


  buf

  (
    G371_o2_p,
    G371_o2
  );


  not

  (
    G371_o2_n,
    G371_o2
  );


  buf

  (
    G1059_o2_p,
    G1059_o2
  );


  not

  (
    G1059_o2_n,
    G1059_o2
  );


  buf

  (
    n2586_o2_p,
    n2586_o2
  );


  not

  (
    n2586_o2_n,
    n2586_o2
  );


  buf

  (
    n2587_o2_p,
    n2587_o2
  );


  not

  (
    n2587_o2_n,
    n2587_o2
  );


  buf

  (
    n460_inv_p,
    n460_inv
  );


  not

  (
    n460_inv_n,
    n460_inv
  );


  buf

  (
    n2648_o2_p,
    n2648_o2
  );


  not

  (
    n2648_o2_n,
    n2648_o2
  );


  buf

  (
    n2649_o2_p,
    n2649_o2
  );


  not

  (
    n2649_o2_n,
    n2649_o2
  );


  buf

  (
    n2650_o2_p,
    n2650_o2
  );


  not

  (
    n2650_o2_n,
    n2650_o2
  );


  buf

  (
    n2651_o2_p,
    n2651_o2
  );


  not

  (
    n2651_o2_n,
    n2651_o2
  );


  buf

  (
    n2652_o2_p,
    n2652_o2
  );


  not

  (
    n2652_o2_n,
    n2652_o2
  );


  buf

  (
    G365_o2_p,
    G365_o2
  );


  not

  (
    G365_o2_n,
    G365_o2
  );


  buf

  (
    G1496_o2_p,
    G1496_o2
  );


  not

  (
    G1496_o2_n,
    G1496_o2
  );


  buf

  (
    G1502_o2_p,
    G1502_o2
  );


  not

  (
    G1502_o2_n,
    G1502_o2
  );


  buf

  (
    n2700_o2_p,
    n2700_o2
  );


  not

  (
    n2700_o2_n,
    n2700_o2
  );


  buf

  (
    n2701_o2_p,
    n2701_o2
  );


  not

  (
    n2701_o2_n,
    n2701_o2
  );


  buf

  (
    n2733_o2_p,
    n2733_o2
  );


  not

  (
    n2733_o2_n,
    n2733_o2
  );


  buf

  (
    n2734_o2_p,
    n2734_o2
  );


  not

  (
    n2734_o2_n,
    n2734_o2
  );


  buf

  (
    n2744_o2_p,
    n2744_o2
  );


  not

  (
    n2744_o2_n,
    n2744_o2
  );


  buf

  (
    n2747_o2_p,
    n2747_o2
  );


  not

  (
    n2747_o2_n,
    n2747_o2
  );


  buf

  (
    n2754_o2_p,
    n2754_o2
  );


  not

  (
    n2754_o2_n,
    n2754_o2
  );


  buf

  (
    n2755_o2_p,
    n2755_o2
  );


  not

  (
    n2755_o2_n,
    n2755_o2
  );


  buf

  (
    n511_inv_p,
    n511_inv
  );


  not

  (
    n511_inv_n,
    n511_inv
  );


  buf

  (
    G1609_o2_p,
    G1609_o2
  );


  not

  (
    G1609_o2_n,
    G1609_o2
  );


  buf

  (
    G1625_o2_p,
    G1625_o2
  );


  not

  (
    G1625_o2_n,
    G1625_o2
  );


  buf

  (
    G738_o2_p,
    G738_o2
  );


  not

  (
    G738_o2_n,
    G738_o2
  );


  buf

  (
    G755_o2_p,
    G755_o2
  );


  not

  (
    G755_o2_n,
    G755_o2
  );


  buf

  (
    G1511_o2_p,
    G1511_o2
  );


  not

  (
    G1511_o2_n,
    G1511_o2
  );


  buf

  (
    G1522_o2_p,
    G1522_o2
  );


  not

  (
    G1522_o2_n,
    G1522_o2
  );


  buf

  (
    G1538_o2_p,
    G1538_o2
  );


  not

  (
    G1538_o2_n,
    G1538_o2
  );


  buf

  (
    G1549_o2_p,
    G1549_o2
  );


  not

  (
    G1549_o2_n,
    G1549_o2
  );


  buf

  (
    G1563_o2_p,
    G1563_o2
  );


  not

  (
    G1563_o2_n,
    G1563_o2
  );


  buf

  (
    G1584_o2_p,
    G1584_o2
  );


  not

  (
    G1584_o2_n,
    G1584_o2
  );


  buf

  (
    G1576_o2_p,
    G1576_o2
  );


  not

  (
    G1576_o2_n,
    G1576_o2
  );


  buf

  (
    G1598_o2_p,
    G1598_o2
  );


  not

  (
    G1598_o2_n,
    G1598_o2
  );


  buf

  (
    G1395_o2_p,
    G1395_o2
  );


  not

  (
    G1395_o2_n,
    G1395_o2
  );


  buf

  (
    G1410_o2_p,
    G1410_o2
  );


  not

  (
    G1410_o2_n,
    G1410_o2
  );


  buf

  (
    G1420_o2_p,
    G1420_o2
  );


  not

  (
    G1420_o2_n,
    G1420_o2
  );


  buf

  (
    G1434_o2_p,
    G1434_o2
  );


  not

  (
    G1434_o2_n,
    G1434_o2
  );


  buf

  (
    n562_inv_p,
    n562_inv
  );


  not

  (
    n562_inv_n,
    n562_inv
  );


  buf

  (
    n1162_lo_buf_o2_p,
    n1162_lo_buf_o2
  );


  not

  (
    n1162_lo_buf_o2_n,
    n1162_lo_buf_o2
  );


  buf

  (
    n1102_lo_buf_o2_p,
    n1102_lo_buf_o2
  );


  not

  (
    n1102_lo_buf_o2_n,
    n1102_lo_buf_o2
  );


  buf

  (
    G359_o2_p,
    G359_o2
  );


  not

  (
    G359_o2_n,
    G359_o2
  );


  buf

  (
    n982_lo_buf_o2_p,
    n982_lo_buf_o2
  );


  not

  (
    n982_lo_buf_o2_n,
    n982_lo_buf_o2
  );


  buf

  (
    n1030_lo_buf_o2_p,
    n1030_lo_buf_o2
  );


  not

  (
    n1030_lo_buf_o2_n,
    n1030_lo_buf_o2
  );


  buf

  (
    n1042_lo_buf_o2_p,
    n1042_lo_buf_o2
  );


  not

  (
    n1042_lo_buf_o2_n,
    n1042_lo_buf_o2
  );


  buf

  (
    n583_inv_p,
    n583_inv
  );


  not

  (
    n583_inv_n,
    n583_inv
  );


  buf

  (
    G606_o2_p,
    G606_o2
  );


  not

  (
    G606_o2_n,
    G606_o2
  );


  buf

  (
    G1118_o2_p,
    G1118_o2
  );


  not

  (
    G1118_o2_n,
    G1118_o2
  );


  buf

  (
    G1069_o2_p,
    G1069_o2
  );


  not

  (
    G1069_o2_n,
    G1069_o2
  );


  buf

  (
    G1145_o2_p,
    G1145_o2
  );


  not

  (
    G1145_o2_n,
    G1145_o2
  );


  buf

  (
    G1209_o2_p,
    G1209_o2
  );


  not

  (
    G1209_o2_n,
    G1209_o2
  );


  buf

  (
    G1189_o2_p,
    G1189_o2
  );


  not

  (
    G1189_o2_n,
    G1189_o2
  );


  buf

  (
    G1699_o2_p,
    G1699_o2
  );


  not

  (
    G1699_o2_n,
    G1699_o2
  );


  buf

  (
    G1702_o2_p,
    G1702_o2
  );


  not

  (
    G1702_o2_n,
    G1702_o2
  );


  buf

  (
    G1705_o2_p,
    G1705_o2
  );


  not

  (
    G1705_o2_n,
    G1705_o2
  );


  buf

  (
    G1708_o2_p,
    G1708_o2
  );


  not

  (
    G1708_o2_n,
    G1708_o2
  );


  buf

  (
    G1684_o2_p,
    G1684_o2
  );


  not

  (
    G1684_o2_n,
    G1684_o2
  );


  buf

  (
    G1687_o2_p,
    G1687_o2
  );


  not

  (
    G1687_o2_n,
    G1687_o2
  );


  buf

  (
    G1690_o2_p,
    G1690_o2
  );


  not

  (
    G1690_o2_n,
    G1690_o2
  );


  buf

  (
    G1693_o2_p,
    G1693_o2
  );


  not

  (
    G1693_o2_n,
    G1693_o2
  );


  buf

  (
    G1696_o2_p,
    G1696_o2
  );


  not

  (
    G1696_o2_n,
    G1696_o2
  );


  buf

  (
    G1642_o2_p,
    G1642_o2
  );


  not

  (
    G1642_o2_n,
    G1642_o2
  );


  buf

  (
    G1645_o2_p,
    G1645_o2
  );


  not

  (
    G1645_o2_n,
    G1645_o2
  );


  buf

  (
    G1648_o2_p,
    G1648_o2
  );


  not

  (
    G1648_o2_n,
    G1648_o2
  );


  buf

  (
    G1651_o2_p,
    G1651_o2
  );


  not

  (
    G1651_o2_n,
    G1651_o2
  );


  buf

  (
    G1654_o2_p,
    G1654_o2
  );


  not

  (
    G1654_o2_n,
    G1654_o2
  );


  buf

  (
    G1657_o2_p,
    G1657_o2
  );


  not

  (
    G1657_o2_n,
    G1657_o2
  );


  buf

  (
    G1660_o2_p,
    G1660_o2
  );


  not

  (
    G1660_o2_n,
    G1660_o2
  );


  buf

  (
    n1222_lo_buf_o2_p,
    n1222_lo_buf_o2
  );


  not

  (
    n1222_lo_buf_o2_n,
    n1222_lo_buf_o2
  );


  buf

  (
    n1330_lo_buf_o2_p,
    n1330_lo_buf_o2
  );


  not

  (
    n1330_lo_buf_o2_n,
    n1330_lo_buf_o2
  );


  buf

  (
    n658_inv_p,
    n658_inv
  );


  not

  (
    n658_inv_n,
    n658_inv
  );


  buf

  (
    n661_inv_p,
    n661_inv
  );


  not

  (
    n661_inv_n,
    n661_inv
  );


  buf

  (
    n1306_lo_buf_o2_p,
    n1306_lo_buf_o2
  );


  not

  (
    n1306_lo_buf_o2_n,
    n1306_lo_buf_o2
  );


  buf

  (
    n1150_lo_buf_o2_p,
    n1150_lo_buf_o2
  );


  not

  (
    n1150_lo_buf_o2_n,
    n1150_lo_buf_o2
  );


  buf

  (
    G175_o2_p,
    G175_o2
  );


  not

  (
    G175_o2_n,
    G175_o2
  );


  buf

  (
    G241_o2_p,
    G241_o2
  );


  not

  (
    G241_o2_n,
    G241_o2
  );


  buf

  (
    G356_o2_p,
    G356_o2
  );


  not

  (
    G356_o2_n,
    G356_o2
  );


  buf

  (
    G989_o2_p,
    G989_o2
  );


  not

  (
    G989_o2_n,
    G989_o2
  );


  buf

  (
    G984_o2_p,
    G984_o2
  );


  not

  (
    G984_o2_n,
    G984_o2
  );


  buf

  (
    n685_inv_p,
    n685_inv
  );


  not

  (
    n685_inv_n,
    n685_inv
  );


  buf

  (
    n688_inv_p,
    n688_inv
  );


  not

  (
    n688_inv_n,
    n688_inv
  );


  buf

  (
    n958_lo_buf_o2_p,
    n958_lo_buf_o2
  );


  not

  (
    n958_lo_buf_o2_n,
    n958_lo_buf_o2
  );


  buf

  (
    n1114_lo_buf_o2_p,
    n1114_lo_buf_o2
  );


  not

  (
    n1114_lo_buf_o2_n,
    n1114_lo_buf_o2
  );


  buf

  (
    G182_o2_p,
    G182_o2
  );


  not

  (
    G182_o2_n,
    G182_o2
  );


  buf

  (
    G1215_o2_p,
    G1215_o2
  );


  not

  (
    G1215_o2_n,
    G1215_o2
  );


  buf

  (
    G971_o2_p,
    G971_o2
  );


  not

  (
    G971_o2_n,
    G971_o2
  );


  buf

  (
    G938_o2_p,
    G938_o2
  );


  not

  (
    G938_o2_n,
    G938_o2
  );


  buf

  (
    G1198_o2_p,
    G1198_o2
  );


  not

  (
    G1198_o2_n,
    G1198_o2
  );


  buf

  (
    G1203_o2_p,
    G1203_o2
  );


  not

  (
    G1203_o2_n,
    G1203_o2
  );


  buf

  (
    G1218_o2_p,
    G1218_o2
  );


  not

  (
    G1218_o2_n,
    G1218_o2
  );


  buf

  (
    G785_o2_p,
    G785_o2
  );


  not

  (
    G785_o2_n,
    G785_o2
  );


  buf

  (
    G1168_o2_p,
    G1168_o2
  );


  not

  (
    G1168_o2_n,
    G1168_o2
  );


  buf

  (
    G1130_o2_p,
    G1130_o2
  );


  not

  (
    G1130_o2_n,
    G1130_o2
  );


  buf

  (
    G1185_o2_p,
    G1185_o2
  );


  not

  (
    G1185_o2_n,
    G1185_o2
  );


  buf

  (
    G1250_o2_p,
    G1250_o2
  );


  not

  (
    G1250_o2_n,
    G1250_o2
  );


  buf

  (
    G1225_o2_p,
    G1225_o2
  );


  not

  (
    G1225_o2_n,
    G1225_o2
  );


  buf

  (
    G1791_o2_p,
    G1791_o2
  );


  not

  (
    G1791_o2_n,
    G1791_o2
  );


  buf

  (
    G1788_o2_p,
    G1788_o2
  );


  not

  (
    G1788_o2_n,
    G1788_o2
  );


  buf

  (
    G981_o2_p,
    G981_o2
  );


  not

  (
    G981_o2_n,
    G981_o2
  );


  buf

  (
    n745_inv_p,
    n745_inv
  );


  not

  (
    n745_inv_n,
    n745_inv
  );


  buf

  (
    n748_inv_p,
    n748_inv
  );


  not

  (
    n748_inv_n,
    n748_inv
  );


  buf

  (
    G1062_o2_p,
    G1062_o2
  );


  not

  (
    G1062_o2_n,
    G1062_o2
  );


  buf

  (
    n970_lo_buf_o2_p,
    n970_lo_buf_o2
  );


  not

  (
    n970_lo_buf_o2_n,
    n970_lo_buf_o2
  );


  buf

  (
    n1006_lo_buf_o2_p,
    n1006_lo_buf_o2
  );


  not

  (
    n1006_lo_buf_o2_n,
    n1006_lo_buf_o2
  );


  buf

  (
    n1078_lo_buf_o2_p,
    n1078_lo_buf_o2
  );


  not

  (
    n1078_lo_buf_o2_n,
    n1078_lo_buf_o2
  );


  buf

  (
    n1126_lo_buf_o2_p,
    n1126_lo_buf_o2
  );


  not

  (
    n1126_lo_buf_o2_n,
    n1126_lo_buf_o2
  );


  buf

  (
    n766_inv_p,
    n766_inv
  );


  not

  (
    n766_inv_n,
    n766_inv
  );


  buf

  (
    G165_o2_p,
    G165_o2
  );


  not

  (
    G165_o2_n,
    G165_o2
  );


  buf

  (
    n1234_lo_buf_o2_p,
    n1234_lo_buf_o2
  );


  not

  (
    n1234_lo_buf_o2_n,
    n1234_lo_buf_o2
  );


  buf

  (
    n1246_lo_buf_o2_p,
    n1246_lo_buf_o2
  );


  not

  (
    n1246_lo_buf_o2_n,
    n1246_lo_buf_o2
  );


  buf

  (
    n1258_lo_buf_o2_p,
    n1258_lo_buf_o2
  );


  not

  (
    n1258_lo_buf_o2_n,
    n1258_lo_buf_o2
  );


  buf

  (
    n1270_lo_buf_o2_p,
    n1270_lo_buf_o2
  );


  not

  (
    n1270_lo_buf_o2_n,
    n1270_lo_buf_o2
  );


  buf

  (
    G368_o2_p,
    G368_o2
  );


  not

  (
    G368_o2_n,
    G368_o2
  );


  buf

  (
    G428_o2_p,
    G428_o2
  );


  not

  (
    G428_o2_n,
    G428_o2
  );


  buf

  (
    G212_o2_p,
    G212_o2
  );


  not

  (
    G212_o2_n,
    G212_o2
  );


  buf

  (
    G841_o2_p,
    G841_o2
  );


  not

  (
    G841_o2_n,
    G841_o2
  );


  buf

  (
    G788_o2_p,
    G788_o2
  );


  not

  (
    G788_o2_n,
    G788_o2
  );


  buf

  (
    n1186_lo_buf_o2_p,
    n1186_lo_buf_o2
  );


  not

  (
    n1186_lo_buf_o2_n,
    n1186_lo_buf_o2
  );


  buf

  (
    G391_o2_p,
    G391_o2
  );


  not

  (
    G391_o2_n,
    G391_o2
  );


  buf

  (
    G387_o2_p,
    G387_o2
  );


  not

  (
    G387_o2_n,
    G387_o2
  );


  buf

  (
    G645_o2_p,
    G645_o2
  );


  not

  (
    G645_o2_n,
    G645_o2
  );


  buf

  (
    G1140_o2_p,
    G1140_o2
  );


  not

  (
    G1140_o2_n,
    G1140_o2
  );


  buf

  (
    G1178_o2_p,
    G1178_o2
  );


  not

  (
    G1178_o2_n,
    G1178_o2
  );


  buf

  (
    G1370_o2_p,
    G1370_o2
  );


  not

  (
    G1370_o2_n,
    G1370_o2
  );


  buf

  (
    n820_inv_p,
    n820_inv
  );


  not

  (
    n820_inv_n,
    n820_inv
  );


  buf

  (
    G1357_o2_p,
    G1357_o2
  );


  not

  (
    G1357_o2_n,
    G1357_o2
  );


  buf

  (
    G816_o2_p,
    G816_o2
  );


  not

  (
    G816_o2_n,
    G816_o2
  );


  buf

  (
    G1369_o2_p,
    G1369_o2
  );


  not

  (
    G1369_o2_n,
    G1369_o2
  );


  buf

  (
    G901_o2_p,
    G901_o2
  );


  not

  (
    G901_o2_n,
    G901_o2
  );


  buf

  (
    G1056_o2_p,
    G1056_o2
  );


  not

  (
    G1056_o2_n,
    G1056_o2
  );


  buf

  (
    G1107_o2_p,
    G1107_o2
  );


  not

  (
    G1107_o2_n,
    G1107_o2
  );


  buf

  (
    G1087_o2_p,
    G1087_o2
  );


  not

  (
    G1087_o2_n,
    G1087_o2
  );


  buf

  (
    G1135_o2_p,
    G1135_o2
  );


  not

  (
    G1135_o2_n,
    G1135_o2
  );


  buf

  (
    n1018_lo_buf_o2_p,
    n1018_lo_buf_o2
  );


  not

  (
    n1018_lo_buf_o2_n,
    n1018_lo_buf_o2
  );


  buf

  (
    n1090_lo_buf_o2_p,
    n1090_lo_buf_o2
  );


  not

  (
    n1090_lo_buf_o2_n,
    n1090_lo_buf_o2
  );


  buf

  (
    n853_inv_p,
    n853_inv
  );


  not

  (
    n853_inv_n,
    n853_inv
  );


  buf

  (
    G131_o2_p,
    G131_o2
  );


  not

  (
    G131_o2_n,
    G131_o2
  );


  buf

  (
    n859_inv_p,
    n859_inv
  );


  not

  (
    n859_inv_n,
    n859_inv
  );


  buf

  (
    n862_inv_p,
    n862_inv
  );


  not

  (
    n862_inv_n,
    n862_inv
  );


  buf

  (
    G338_o2_p,
    G338_o2
  );


  not

  (
    G338_o2_n,
    G338_o2
  );


  buf

  (
    n1171_lo_buf_o2_p,
    n1171_lo_buf_o2
  );


  not

  (
    n1171_lo_buf_o2_n,
    n1171_lo_buf_o2
  );


  buf

  (
    n1195_lo_buf_o2_p,
    n1195_lo_buf_o2
  );


  not

  (
    n1195_lo_buf_o2_n,
    n1195_lo_buf_o2
  );


  buf

  (
    G419_o2_p,
    G419_o2
  );


  not

  (
    G419_o2_n,
    G419_o2
  );


  buf

  (
    G425_o2_p,
    G425_o2
  );


  not

  (
    G425_o2_n,
    G425_o2
  );


  buf

  (
    G497_o2_p,
    G497_o2
  );


  not

  (
    G497_o2_n,
    G497_o2
  );


  buf

  (
    G416_o2_p,
    G416_o2
  );


  not

  (
    G416_o2_n,
    G416_o2
  );


  buf

  (
    G491_o2_p,
    G491_o2
  );


  not

  (
    G491_o2_n,
    G491_o2
  );


  buf

  (
    G500_o2_p,
    G500_o2
  );


  not

  (
    G500_o2_n,
    G500_o2
  );


  buf

  (
    G353_o2_p,
    G353_o2
  );


  not

  (
    G353_o2_n,
    G353_o2
  );


  buf

  (
    G641_o2_p,
    G641_o2
  );


  not

  (
    G641_o2_n,
    G641_o2
  );


  buf

  (
    G1117_o2_p,
    G1117_o2
  );


  not

  (
    G1117_o2_n,
    G1117_o2
  );


  buf

  (
    G1096_o2_p,
    G1096_o2
  );


  not

  (
    G1096_o2_n,
    G1096_o2
  );


  buf

  (
    G1143_o2_p,
    G1143_o2
  );


  not

  (
    G1143_o2_n,
    G1143_o2
  );


  buf

  (
    G1112_o2_p,
    G1112_o2
  );


  not

  (
    G1112_o2_n,
    G1112_o2
  );


  buf

  (
    n1138_lo_buf_o2_p,
    n1138_lo_buf_o2
  );


  not

  (
    n1138_lo_buf_o2_n,
    n1138_lo_buf_o2
  );


  buf

  (
    n1210_lo_buf_o2_p,
    n1210_lo_buf_o2
  );


  not

  (
    n1210_lo_buf_o2_n,
    n1210_lo_buf_o2
  );


  buf

  (
    G687_o2_p,
    G687_o2
  );


  not

  (
    G687_o2_n,
    G687_o2
  );


  buf

  (
    G541_o2_p,
    G541_o2
  );


  not

  (
    G541_o2_n,
    G541_o2
  );


  buf

  (
    G802_o2_p,
    G802_o2
  );


  not

  (
    G802_o2_n,
    G802_o2
  );


  buf

  (
    G813_o2_p,
    G813_o2
  );


  not

  (
    G813_o2_n,
    G813_o2
  );


  buf

  (
    G810_o2_p,
    G810_o2
  );


  not

  (
    G810_o2_n,
    G810_o2
  );


  buf

  (
    G987_o2_p,
    G987_o2
  );


  not

  (
    G987_o2_n,
    G987_o2
  );


  buf

  (
    G898_o2_p,
    G898_o2
  );


  not

  (
    G898_o2_n,
    G898_o2
  );


  buf

  (
    n946_lo_buf_o2_p,
    n946_lo_buf_o2
  );


  not

  (
    n946_lo_buf_o2_n,
    n946_lo_buf_o2
  );


  buf

  (
    n1054_lo_buf_o2_p,
    n1054_lo_buf_o2
  );


  not

  (
    n1054_lo_buf_o2_n,
    n1054_lo_buf_o2
  );


  buf

  (
    G728_o2_p,
    G728_o2
  );


  not

  (
    G728_o2_n,
    G728_o2
  );


  buf

  (
    G856_o2_p,
    G856_o2
  );


  not

  (
    G856_o2_n,
    G856_o2
  );


  buf

  (
    n949_1_inv_p,
    n949_1_inv
  );


  not

  (
    n949_1_inv_n,
    n949_1_inv
  );


  buf

  (
    G942_o2_p,
    G942_o2
  );


  not

  (
    G942_o2_n,
    G942_o2
  );


  buf

  (
    G1099_o2_p,
    G1099_o2
  );


  not

  (
    G1099_o2_n,
    G1099_o2
  );


  buf

  (
    G1154_o2_p,
    G1154_o2
  );


  not

  (
    G1154_o2_n,
    G1154_o2
  );


  buf

  (
    G1131_o2_p,
    G1131_o2
  );


  not

  (
    G1131_o2_n,
    G1131_o2
  );


  buf

  (
    G1169_o2_p,
    G1169_o2
  );


  not

  (
    G1169_o2_n,
    G1169_o2
  );


  buf

  (
    G134_o2_p,
    G134_o2
  );


  not

  (
    G134_o2_n,
    G134_o2
  );


  buf

  (
    n970_inv_p,
    n970_inv
  );


  not

  (
    n970_inv_n,
    n970_inv
  );


  buf

  (
    G470_o2_p,
    G470_o2
  );


  not

  (
    G470_o2_n,
    G470_o2
  );


  buf

  (
    G344_o2_p,
    G344_o2
  );


  not

  (
    G344_o2_n,
    G344_o2
  );


  buf

  (
    G362_o2_p,
    G362_o2
  );


  not

  (
    G362_o2_n,
    G362_o2
  );


  buf

  (
    G482_o2_p,
    G482_o2
  );


  not

  (
    G482_o2_n,
    G482_o2
  );


  buf

  (
    G660_o2_p,
    G660_o2
  );


  not

  (
    G660_o2_n,
    G660_o2
  );


  buf

  (
    G672_o2_p,
    G672_o2
  );


  not

  (
    G672_o2_n,
    G672_o2
  );


  buf

  (
    n1096_lo_buf_o2_p,
    n1096_lo_buf_o2
  );


  not

  (
    n1096_lo_buf_o2_n,
    n1096_lo_buf_o2
  );


  buf

  (
    G479_o2_p,
    G479_o2
  );


  not

  (
    G479_o2_n,
    G479_o2
  );


  buf

  (
    G669_o2_p,
    G669_o2
  );


  not

  (
    G669_o2_n,
    G669_o2
  );


  buf

  (
    n994_lo_buf_o2_p,
    n994_lo_buf_o2
  );


  not

  (
    n994_lo_buf_o2_n,
    n994_lo_buf_o2
  );


  buf

  (
    n1066_lo_buf_o2_p,
    n1066_lo_buf_o2
  );


  not

  (
    n1066_lo_buf_o2_n,
    n1066_lo_buf_o2
  );


  buf

  (
    n1006_inv_p,
    n1006_inv
  );


  not

  (
    n1006_inv_n,
    n1006_inv
  );


  buf

  (
    G147_o2_p,
    G147_o2
  );


  not

  (
    G147_o2_n,
    G147_o2
  );


  buf

  (
    G473_o2_p,
    G473_o2
  );


  not

  (
    G473_o2_n,
    G473_o2
  );


  buf

  (
    G488_o2_p,
    G488_o2
  );


  not

  (
    G488_o2_n,
    G488_o2
  );


  buf

  (
    G589_o2_p,
    G589_o2
  );


  not

  (
    G589_o2_n,
    G589_o2
  );


  buf

  (
    G663_o2_p,
    G663_o2
  );


  not

  (
    G663_o2_n,
    G663_o2
  );


  buf

  (
    G684_o2_p,
    G684_o2
  );


  not

  (
    G684_o2_n,
    G684_o2
  );


  buf

  (
    G605_o2_p,
    G605_o2
  );


  not

  (
    G605_o2_n,
    G605_o2
  );


  buf

  (
    G774_o2_p,
    G774_o2
  );


  not

  (
    G774_o2_n,
    G774_o2
  );


  buf

  (
    G782_o2_p,
    G782_o2
  );


  not

  (
    G782_o2_n,
    G782_o2
  );


  and

  (
    g359_p,
    G1538_o2_n_spl_,
    G1511_o2_n_spl_
  );


  or

  (
    g359_n,
    G1538_o2_p_spl_,
    G1511_o2_p_spl_
  );


  and

  (
    g360_p,
    g359_p_spl_0,
    G1584_o2_p_spl_00
  );


  or

  (
    g360_n,
    g359_n_spl_0,
    G1584_o2_n_spl_00
  );


  and

  (
    g361_p,
    g360_p,
    G1395_o2_n_spl_000
  );


  or

  (
    g361_n,
    g360_n,
    G1395_o2_p_spl_0
  );


  and

  (
    g362_p,
    g361_p,
    G738_o2_n_spl_00
  );


  or

  (
    g362_n,
    g361_n,
    G738_o2_p_spl_00
  );


  and

  (
    g363_p,
    g362_p,
    n949_lo_p
  );


  and

  (
    g364_p,
    g362_n,
    n949_lo_n
  );


  or

  (
    g365_n,
    g364_p,
    g363_p
  );


  and

  (
    g366_p,
    g359_p_spl_0,
    G1563_o2_p_spl_00
  );


  or

  (
    g366_n,
    g359_n_spl_0,
    G1563_o2_n_spl_
  );


  and

  (
    g367_p,
    g366_p_spl_,
    G1420_o2_n_spl_00
  );


  or

  (
    g367_n,
    g366_n_spl_,
    G1420_o2_p_spl_00
  );


  and

  (
    g368_p,
    g367_p,
    G738_o2_n_spl_00
  );


  or

  (
    g368_n,
    g367_n,
    G738_o2_p_spl_00
  );


  and

  (
    g369_p,
    g368_p,
    n961_lo_p
  );


  and

  (
    g370_p,
    g368_n,
    n961_lo_n
  );


  or

  (
    g371_n,
    g370_p,
    g369_p
  );


  and

  (
    g372_p,
    g366_p_spl_,
    G1410_o2_n_spl_00
  );


  or

  (
    g372_n,
    g366_n_spl_,
    G1410_o2_p_spl_0
  );


  and

  (
    g373_p,
    g372_p,
    G738_o2_n_spl_01
  );


  or

  (
    g373_n,
    g372_n,
    G738_o2_p_spl_01
  );


  and

  (
    g374_p,
    g373_p,
    n973_lo_p
  );


  and

  (
    g375_p,
    g373_n,
    n973_lo_n
  );


  or

  (
    g376_n,
    g375_p,
    g374_p
  );


  and

  (
    g377_p,
    g359_p_spl_,
    G1576_o2_p_spl_0
  );


  or

  (
    g377_n,
    g359_n_spl_,
    G1576_o2_n_spl_0
  );


  and

  (
    g378_p,
    g377_p,
    G1395_o2_n_spl_000
  );


  or

  (
    g378_n,
    g377_n,
    G1395_o2_p_spl_0
  );


  and

  (
    g379_p,
    g378_p,
    G738_o2_n_spl_01
  );


  or

  (
    g379_n,
    g378_n,
    G738_o2_p_spl_01
  );


  and

  (
    g380_p,
    g379_p,
    n985_lo_p
  );


  and

  (
    g381_p,
    g379_n,
    n985_lo_n
  );


  or

  (
    g382_n,
    g381_p,
    g380_p
  );


  and

  (
    g383_p,
    G1538_o2_n_spl_,
    G1522_o2_n_spl_0
  );


  or

  (
    g383_n,
    G1538_o2_p_spl_,
    G1522_o2_p_spl_0
  );


  and

  (
    g384_p,
    g383_p,
    G1598_o2_p_spl_0
  );


  or

  (
    g384_n,
    g383_n,
    G1598_o2_n_spl_0
  );


  and

  (
    g385_p,
    g384_p,
    G1410_o2_n_spl_00
  );


  or

  (
    g385_n,
    g384_n,
    G1410_o2_p_spl_0
  );


  and

  (
    g386_p,
    g385_p,
    G755_o2_n_spl_00
  );


  or

  (
    g386_n,
    g385_n,
    G755_o2_p_spl_00
  );


  and

  (
    g387_p,
    g386_p,
    n1057_lo_p
  );


  and

  (
    g388_p,
    g386_n,
    n1057_lo_n
  );


  or

  (
    g389_n,
    g388_p,
    g387_p
  );


  and

  (
    g390_p,
    G1549_o2_n_spl_,
    G1522_o2_n_spl_0
  );


  or

  (
    g390_n,
    G1549_o2_p_spl_,
    G1522_o2_p_spl_0
  );


  and

  (
    g391_p,
    g390_p_spl_,
    G1584_o2_p_spl_00
  );


  or

  (
    g391_n,
    g390_n_spl_,
    G1584_o2_n_spl_00
  );


  and

  (
    g392_p,
    g391_p,
    G1434_o2_n_spl_
  );


  or

  (
    g392_n,
    g391_n,
    G1434_o2_p_spl_
  );


  and

  (
    g393_p,
    g392_p,
    G755_o2_n_spl_00
  );


  or

  (
    g393_n,
    g392_n,
    G755_o2_p_spl_00
  );


  and

  (
    g394_p,
    g393_p,
    n1117_lo_p
  );


  and

  (
    g395_p,
    g393_n,
    n1117_lo_n
  );


  or

  (
    g396_n,
    g395_p,
    g394_p
  );


  and

  (
    g397_p,
    g390_p_spl_,
    G1598_o2_p_spl_0
  );


  or

  (
    g397_n,
    g390_n_spl_,
    G1598_o2_n_spl_0
  );


  and

  (
    g398_p,
    g397_p,
    G1420_o2_n_spl_00
  );


  or

  (
    g398_n,
    g397_n,
    G1420_o2_p_spl_00
  );


  and

  (
    g399_p,
    g398_p,
    G755_o2_n_spl_01
  );


  or

  (
    g399_n,
    g398_n,
    G755_o2_p_spl_01
  );


  and

  (
    g400_p,
    g399_p,
    n1129_lo_p
  );


  and

  (
    g401_p,
    g399_n,
    n1129_lo_n
  );


  or

  (
    g402_n,
    g401_p,
    g400_p
  );


  and

  (
    g403_p,
    G1511_o2_n_spl_,
    G1625_o2_p_spl_0
  );


  or

  (
    g403_n,
    G1511_o2_p_spl_,
    G1625_o2_n_spl_
  );


  and

  (
    g404_p,
    g403_p,
    G1584_o2_p_spl_01
  );


  or

  (
    g404_n,
    g403_n,
    G1584_o2_n_spl_0
  );


  and

  (
    g405_p,
    g404_p,
    G1420_o2_n_spl_01
  );


  or

  (
    g405_n,
    g404_n,
    G1420_o2_p_spl_01
  );


  and

  (
    g406_p,
    g405_p,
    G738_o2_n_spl_10
  );


  or

  (
    g406_n,
    g405_n,
    G738_o2_p_spl_10
  );


  and

  (
    g407_p,
    g406_p,
    n997_lo_p
  );


  and

  (
    g408_p,
    g406_n,
    n997_lo_n
  );


  or

  (
    g409_n,
    g408_p,
    g407_p
  );


  and

  (
    g410_p,
    G1522_o2_n_spl_,
    G1625_o2_p_spl_0
  );


  or

  (
    g410_n,
    G1522_o2_p_spl_,
    G1625_o2_n_spl_
  );


  and

  (
    g411_p,
    g410_p_spl_0,
    G1584_o2_p_spl_01
  );


  or

  (
    g411_n,
    g410_n_spl_0,
    G1584_o2_n_spl_1
  );


  and

  (
    g412_p,
    g411_p,
    G1410_o2_n_spl_0
  );


  or

  (
    g412_n,
    g411_n,
    G1410_o2_p_spl_1
  );


  and

  (
    g413_p,
    g412_p,
    G738_o2_n_spl_10
  );


  or

  (
    g413_n,
    g412_n,
    G738_o2_p_spl_10
  );


  and

  (
    g414_p,
    g413_p,
    n1009_lo_p
  );


  and

  (
    g415_p,
    g413_n,
    n1009_lo_n
  );


  or

  (
    g416_n,
    g415_p,
    g414_p
  );


  and

  (
    g417_p,
    g410_p_spl_0,
    G1598_o2_p_spl_1
  );


  or

  (
    g417_n,
    g410_n_spl_0,
    G1598_o2_n_spl_1
  );


  and

  (
    g418_p,
    g417_p,
    G1395_o2_n_spl_001
  );


  or

  (
    g418_n,
    g417_n,
    G1395_o2_p_spl_1
  );


  and

  (
    g419_p,
    g418_p,
    G738_o2_n_spl_11
  );


  or

  (
    g419_n,
    g418_n,
    G738_o2_p_spl_11
  );


  and

  (
    g420_p,
    g419_p,
    n1021_lo_p
  );


  and

  (
    g421_p,
    g419_n,
    n1021_lo_n
  );


  or

  (
    g422_n,
    g421_p,
    g420_p
  );


  and

  (
    g423_p,
    g410_p_spl_1,
    G1563_o2_p_spl_00
  );


  or

  (
    g423_n,
    g410_n_spl_1,
    G1563_o2_n_spl_
  );


  and

  (
    g424_p,
    g423_p_spl_,
    G1434_o2_n_spl_
  );


  or

  (
    g424_n,
    g423_n,
    G1434_o2_p_spl_
  );


  and

  (
    g425_p,
    g424_p,
    G738_o2_n_spl_11
  );


  or

  (
    g425_n,
    g424_n,
    G738_o2_p_spl_11
  );


  and

  (
    g426_p,
    g425_p,
    n1033_lo_p
  );


  and

  (
    g427_p,
    g425_n,
    n1033_lo_n
  );


  or

  (
    g428_n,
    g427_p,
    g426_p
  );


  and

  (
    g429_p,
    g410_p_spl_1,
    G1576_o2_p_spl_0
  );


  or

  (
    g429_n,
    g410_n_spl_1,
    G1576_o2_n_spl_0
  );


  and

  (
    g430_p,
    g429_p,
    G1420_o2_n_spl_01
  );


  or

  (
    g430_n,
    g429_n,
    G1420_o2_p_spl_01
  );


  and

  (
    g431_p,
    g430_p,
    G755_o2_n_spl_01
  );


  or

  (
    g431_n,
    g430_n,
    G755_o2_p_spl_01
  );


  and

  (
    g432_p,
    g431_p,
    n1045_lo_p
  );


  and

  (
    g433_p,
    g431_n,
    n1045_lo_n
  );


  or

  (
    g434_n,
    g433_p,
    g432_p
  );


  and

  (
    g435_p,
    G1549_o2_n_spl_,
    G1609_o2_p_spl_0
  );


  or

  (
    g435_n,
    G1549_o2_p_spl_,
    G1609_o2_n
  );


  and

  (
    g436_p,
    g435_p_spl_0,
    G1584_o2_p_spl_1
  );


  or

  (
    g436_n,
    g435_n_spl_0,
    G1584_o2_n_spl_1
  );


  and

  (
    g437_p,
    g436_p_spl_,
    G1420_o2_n_spl_10
  );


  or

  (
    g437_n,
    g436_n_spl_,
    G1420_o2_p_spl_1
  );


  and

  (
    g438_p,
    g437_p,
    G755_o2_n_spl_10
  );


  or

  (
    g438_n,
    g437_n,
    G755_o2_p_spl_10
  );


  and

  (
    g439_p,
    g438_p,
    n1069_lo_p
  );


  and

  (
    g440_p,
    g438_n,
    n1069_lo_n
  );


  or

  (
    g441_n,
    g440_p,
    g439_p
  );


  and

  (
    g442_p,
    g436_p_spl_,
    G1410_o2_n_spl_1
  );


  or

  (
    g442_n,
    g436_n_spl_,
    G1410_o2_p_spl_1
  );


  and

  (
    g443_p,
    g442_p,
    G755_o2_n_spl_10
  );


  or

  (
    g443_n,
    g442_n,
    G755_o2_p_spl_10
  );


  and

  (
    g444_p,
    g443_p,
    n1081_lo_p
  );


  and

  (
    g445_p,
    g443_n,
    n1081_lo_n
  );


  or

  (
    g446_n,
    g445_p,
    g444_p
  );


  and

  (
    g447_p,
    g435_p_spl_0,
    G1598_o2_p_spl_1
  );


  or

  (
    g447_n,
    g435_n_spl_0,
    G1598_o2_n_spl_1
  );


  and

  (
    g448_p,
    g447_p,
    G1395_o2_n_spl_001
  );


  or

  (
    g448_n,
    g447_n,
    G1395_o2_p_spl_1
  );


  and

  (
    g449_p,
    g448_p,
    G755_o2_n_spl_11
  );


  or

  (
    g449_n,
    g448_n,
    G755_o2_p_spl_11
  );


  and

  (
    g450_p,
    g449_p,
    n1093_lo_p
  );


  and

  (
    g451_p,
    g449_n,
    n1093_lo_n
  );


  or

  (
    g452_n,
    g451_p,
    g450_p
  );


  and

  (
    g453_p,
    g435_p_spl_1,
    G1576_o2_p_spl_1
  );


  or

  (
    g453_n,
    g435_n_spl_,
    G1576_o2_n_spl_
  );


  and

  (
    g454_p,
    g453_p,
    G1420_o2_n_spl_10
  );


  or

  (
    g454_n,
    g453_n,
    G1420_o2_p_spl_1
  );


  and

  (
    g455_p,
    g454_p,
    G755_o2_n_spl_11
  );


  or

  (
    g455_n,
    g454_n,
    G755_o2_p_spl_11
  );


  and

  (
    g456_p,
    g455_p,
    n1105_lo_p
  );


  and

  (
    g457_p,
    g455_n,
    n1105_lo_n
  );


  or

  (
    g458_n,
    g457_p,
    g456_p
  );


  or

  (
    g459_n,
    G1247_o2_p,
    G557_o2_p
  );


  or

  (
    g460_n,
    G1247_o2_n,
    G557_o2_n
  );


  and

  (
    g461_p,
    g460_n,
    g459_n
  );


  or

  (
    g462_n,
    G1182_o2_n,
    G194_o2_p
  );


  or

  (
    g463_n,
    G1182_o2_p,
    G194_o2_n
  );


  and

  (
    g464_p,
    g463_n,
    g462_n
  );


  or

  (
    g465_n,
    G1222_o2_n,
    G191_o2_p
  );


  or

  (
    g466_n,
    G1222_o2_p,
    G191_o2_n
  );


  and

  (
    g467_p,
    g466_n,
    g465_n
  );


  or

  (
    g468_n,
    G1371_o2_p,
    G188_o2_p
  );


  or

  (
    g469_n,
    G1371_o2_n,
    G188_o2_n
  );


  and

  (
    g470_p,
    g469_n,
    g468_n
  );


  or

  (
    g471_n,
    G1386_o2_n,
    G185_o2_p
  );


  or

  (
    g472_n,
    G1386_o2_p,
    G185_o2_n
  );


  and

  (
    g473_p,
    g472_n,
    g471_n
  );


  or

  (
    g474_n,
    G1383_o2_p,
    G554_o2_p
  );


  or

  (
    g475_n,
    G1383_o2_n,
    G554_o2_n
  );


  and

  (
    g476_p,
    g475_n,
    g474_n
  );


  and

  (
    g477_p,
    g464_p,
    g461_p
  );


  and

  (
    g478_p,
    g477_p,
    g467_p
  );


  and

  (
    g479_p,
    g478_p,
    g470_p
  );


  and

  (
    g480_p,
    g479_p,
    G546_o2_n
  );


  and

  (
    g481_p,
    g480_p,
    g473_p
  );


  and

  (
    g482_p,
    g481_p,
    g476_p
  );


  and

  (
    g483_p,
    g482_p,
    G550_o2_n
  );


  or

  (
    g484_n,
    g483_p,
    G260_o2_p
  );


  or

  (
    g485_n,
    g484_n_spl_,
    n1321_lo_p_spl_0
  );


  or

  (
    g486_n,
    g485_n,
    n1321_lo_p_spl_0
  );


  and

  (
    g487_p,
    G260_o2_n,
    G225_o2_n
  );


  and

  (
    g488_p,
    g487_p,
    G382_o2_n
  );


  and

  (
    g489_p,
    g423_p_spl_,
    G1395_o2_n_spl_01
  );


  and

  (
    g490_p,
    g489_p,
    g488_p_spl_00
  );


  and

  (
    g491_p,
    g435_p_spl_1,
    G1563_o2_p_spl_01
  );


  and

  (
    g492_p,
    g491_p,
    G1395_o2_n_spl_01
  );


  and

  (
    g493_p,
    g492_p,
    g488_p_spl_00
  );


  and

  (
    g494_p,
    G1625_o2_p_spl_1,
    G1609_o2_p_spl_0
  );


  and

  (
    g495_p,
    g494_p_spl_0,
    G1584_o2_p_spl_1
  );


  and

  (
    g496_p,
    g495_p,
    G1395_o2_n_spl_10
  );


  and

  (
    g497_p,
    g496_p,
    g488_p_spl_01
  );


  and

  (
    g498_p,
    g494_p_spl_0,
    G1563_o2_p_spl_01
  );


  and

  (
    g499_p,
    g498_p_spl_,
    G1420_o2_n_spl_1
  );


  and

  (
    g500_p,
    g499_p,
    g488_p_spl_01
  );


  and

  (
    g501_p,
    g498_p_spl_,
    G1410_o2_n_spl_1
  );


  and

  (
    g502_p,
    g501_p,
    g488_p_spl_10
  );


  and

  (
    g503_p,
    g494_p_spl_,
    G1576_o2_p_spl_1
  );


  and

  (
    g504_p,
    g503_p,
    G1395_o2_n_spl_10
  );


  and

  (
    g505_p,
    g504_p,
    g488_p_spl_10
  );


  and

  (
    g506_p,
    G1502_o2_n,
    G550_o2_p
  );


  and

  (
    g507_p,
    g506_p,
    G1609_o2_p_spl_
  );


  and

  (
    g508_p,
    g507_p,
    G1563_o2_p_spl_1
  );


  and

  (
    g509_p,
    g508_p,
    G1395_o2_n_spl_11
  );


  and

  (
    g510_p,
    g509_p,
    g488_p_spl_11
  );


  and

  (
    g511_p,
    G1496_o2_p,
    G546_o2_p
  );


  and

  (
    g512_p,
    g511_p,
    G1625_o2_p_spl_1
  );


  and

  (
    g513_p,
    g512_p,
    G1563_o2_p_spl_1
  );


  and

  (
    g514_p,
    g513_p,
    G1395_o2_n_spl_11
  );


  and

  (
    g515_p,
    g514_p,
    g488_p_spl_11
  );


  or

  (
    g516_n,
    g493_p,
    g490_p
  );


  or

  (
    g517_n,
    g516_n,
    g497_p
  );


  or

  (
    g518_n,
    g517_n,
    g500_p
  );


  or

  (
    g519_n,
    g518_n,
    g502_p
  );


  or

  (
    g520_n,
    g519_n,
    g505_p
  );


  or

  (
    g521_n,
    g520_n,
    g510_p
  );


  or

  (
    g522_n,
    g521_n,
    g515_p
  );


  and

  (
    g523_p,
    G1788_o2_n,
    G1791_o2_n
  );


  or

  (
    g523_n,
    G1788_o2_p,
    G1791_o2_p
  );


  or

  (
    g524_n,
    g523_n_spl_00,
    g522_n
  );


  or

  (
    g525_n,
    g484_n_spl_,
    n1321_lo_n
  );


  or

  (
    g526_n,
    g525_n,
    g524_n
  );


  and

  (
    g527_p,
    g526_n,
    g486_n
  );


  and

  (
    g528_p,
    G785_o2_p,
    G1145_o2_p
  );


  or

  (
    g528_n,
    G785_o2_n,
    G1145_o2_n
  );


  and

  (
    g529_p,
    G1185_o2_n,
    G606_o2_n
  );


  or

  (
    g529_n,
    G1185_o2_p,
    G606_o2_p
  );


  and

  (
    g530_p,
    g529_n,
    g528_n
  );


  or

  (
    g530_n,
    g529_p,
    g528_p
  );


  and

  (
    g531_p,
    g530_n_spl_,
    n2372_o2_n_spl_
  );


  or

  (
    g531_n,
    g530_p_spl_,
    n2372_o2_p_spl_
  );


  and

  (
    g532_p,
    g530_p_spl_,
    n2372_o2_p_spl_
  );


  or

  (
    g532_n,
    g530_n_spl_,
    n2372_o2_n_spl_
  );


  and

  (
    g533_p,
    g532_n,
    g531_n
  );


  or

  (
    g533_n,
    g532_p,
    g531_p
  );


  and

  (
    g534_p,
    n2680_o2_p,
    n1141_lo_p
  );


  or

  (
    g534_n,
    n2680_o2_n,
    n1141_lo_n
  );


  and

  (
    g535_p,
    g534_p,
    n1309_lo_n_spl_00
  );


  or

  (
    g535_n,
    g534_n,
    n1309_lo_p_spl_00
  );


  and

  (
    g536_p,
    g535_p,
    g523_n_spl_00
  );


  or

  (
    g536_n,
    g535_n,
    g523_p_spl_00
  );


  and

  (
    g537_p,
    g536_n,
    g533_n
  );


  and

  (
    g538_p,
    g536_p,
    g533_p
  );


  or

  (
    g539_n,
    g538_p,
    g537_p
  );


  or

  (
    g540_n,
    n1333_lo_p_spl_00,
    n1321_lo_p_spl_
  );


  and

  (
    g541_p,
    g540_n_spl_00,
    g539_n
  );


  and

  (
    g542_p,
    G938_o2_n,
    G971_o2_n
  );


  or

  (
    g542_n,
    G938_o2_p,
    G971_o2_p
  );


  and

  (
    g543_p,
    G1168_o2_p,
    G1209_o2_p
  );


  or

  (
    g543_n,
    G1168_o2_n,
    G1209_o2_n
  );


  and

  (
    g544_p,
    G1250_o2_n,
    G1118_o2_n
  );


  or

  (
    g544_n,
    G1250_o2_p,
    G1118_o2_p
  );


  and

  (
    g545_p,
    g544_n,
    g543_n
  );


  or

  (
    g545_n,
    g544_p,
    g543_p
  );


  and

  (
    g546_p,
    g545_p_spl_,
    g542_p_spl_
  );


  or

  (
    g546_n,
    g545_n_spl_,
    g542_n_spl_
  );


  and

  (
    g547_p,
    g545_n_spl_,
    g542_n_spl_
  );


  or

  (
    g547_n,
    g545_p_spl_,
    g542_p_spl_
  );


  and

  (
    g548_p,
    g547_n,
    g546_n
  );


  or

  (
    g548_n,
    g547_p,
    g546_p
  );


  and

  (
    g549_p,
    n1309_lo_n_spl_00,
    n1237_lo_p
  );


  or

  (
    g549_n,
    n1309_lo_p_spl_00,
    n1237_lo_n
  );


  and

  (
    g550_p,
    g549_p,
    g523_n_spl_01
  );


  or

  (
    g550_n,
    g549_n,
    g523_p_spl_00
  );


  and

  (
    g551_p,
    g550_n,
    g548_n
  );


  and

  (
    g552_p,
    g550_p,
    g548_p
  );


  or

  (
    g553_n,
    g552_p,
    g551_p
  );


  and

  (
    g554_p,
    g553_n,
    g540_n_spl_00
  );


  and

  (
    g555_p,
    n1309_lo_n_spl_01,
    n1261_lo_p
  );


  or

  (
    g555_n,
    n1309_lo_p_spl_01,
    n1261_lo_n
  );


  and

  (
    g556_p,
    g555_p,
    g523_n_spl_01
  );


  or

  (
    g556_n,
    g555_n,
    g523_p_spl_01
  );


  and

  (
    g557_p,
    g556_n,
    n2684_o2_n
  );


  and

  (
    g558_p,
    g556_p,
    n2684_o2_p
  );


  or

  (
    g559_n,
    g558_p,
    g557_p
  );


  and

  (
    g560_p,
    g559_n,
    g540_n_spl_01
  );


  and

  (
    g561_p,
    n1309_lo_n_spl_01,
    n1273_lo_p
  );


  or

  (
    g561_n,
    n1309_lo_p_spl_01,
    n1273_lo_n
  );


  and

  (
    g562_p,
    g561_p,
    g523_n_spl_10
  );


  or

  (
    g562_n,
    g561_n,
    g523_p_spl_01
  );


  and

  (
    g563_p,
    g562_n,
    n2683_o2_n
  );


  and

  (
    g564_p,
    g562_p,
    n2683_o2_p
  );


  or

  (
    g565_n,
    g564_p,
    g563_p
  );


  and

  (
    g566_p,
    g565_n,
    g540_n_spl_01
  );


  and

  (
    g567_p,
    n2681_o2_p,
    n1165_lo_p
  );


  or

  (
    g567_n,
    n2681_o2_n,
    n1165_lo_n
  );


  and

  (
    g568_p,
    g567_p,
    n1309_lo_n_spl_1
  );


  or

  (
    g568_n,
    g567_n,
    n1309_lo_p_spl_1
  );


  and

  (
    g569_p,
    g568_p,
    g523_n_spl_10
  );


  or

  (
    g569_n,
    g568_n,
    g523_p_spl_1
  );


  and

  (
    g570_p,
    g569_n,
    n2686_o2_p
  );


  and

  (
    g571_p,
    g569_p,
    n2686_o2_n
  );


  or

  (
    g572_n,
    g571_p,
    g570_p
  );


  and

  (
    g573_p,
    g572_n,
    g540_n_spl_1
  );


  and

  (
    g574_p,
    G1645_o2_n,
    G1642_o2_n
  );


  or

  (
    g574_n,
    G1645_o2_p,
    G1642_o2_p
  );


  and

  (
    g575_p,
    g574_p,
    G1648_o2_n
  );


  or

  (
    g575_n,
    g574_n,
    G1648_o2_p
  );


  and

  (
    g576_p,
    g575_p,
    G1651_o2_n
  );


  or

  (
    g576_n,
    g575_n,
    G1651_o2_p
  );


  and

  (
    g577_p,
    g576_p,
    G1684_o2_n
  );


  or

  (
    g577_n,
    g576_n,
    G1684_o2_p
  );


  and

  (
    g578_p,
    g577_p,
    G1687_o2_n
  );


  or

  (
    g578_n,
    g577_n,
    G1687_o2_p
  );


  and

  (
    g579_p,
    g578_p,
    G1690_o2_n
  );


  or

  (
    g579_n,
    g578_n,
    G1690_o2_p
  );


  and

  (
    g580_p,
    g579_p,
    G1693_o2_n
  );


  or

  (
    g580_n,
    g579_n,
    G1693_o2_p
  );


  and

  (
    g581_p,
    g580_n,
    n1333_lo_n_spl_0
  );


  or

  (
    g581_n,
    g580_p,
    n1333_lo_p_spl_00
  );


  and

  (
    g582_p,
    G1198_o2_p,
    G1215_o2_n
  );


  or

  (
    g582_n,
    G1198_o2_n,
    G1215_o2_p
  );


  and

  (
    g583_p,
    G248_o2_n_spl_,
    G199_o2_n
  );


  or

  (
    g583_n,
    G248_o2_p_spl_,
    G199_o2_p
  );


  and

  (
    g584_p,
    g583_n,
    g582_p
  );


  or

  (
    g584_n,
    g583_p,
    g582_n
  );


  and

  (
    g585_p,
    g584_n_spl_,
    g581_p_spl_
  );


  or

  (
    g585_n,
    g584_p_spl_,
    g581_n_spl_
  );


  and

  (
    g586_p,
    g584_p_spl_,
    g581_n_spl_
  );


  or

  (
    g586_n,
    g584_n_spl_,
    g581_p_spl_
  );


  and

  (
    g587_p,
    g586_n,
    g585_n
  );


  or

  (
    g587_n,
    g586_p,
    g585_p
  );


  and

  (
    g588_p,
    n1285_lo_p,
    n1189_lo_p
  );


  or

  (
    g588_n,
    n1285_lo_n,
    n1189_lo_n
  );


  and

  (
    g589_p,
    g588_n,
    n1333_lo_n_spl_0
  );


  or

  (
    g589_n,
    g588_p,
    n1333_lo_p_spl_0
  );


  and

  (
    g590_p,
    g589_n,
    g587_n
  );


  and

  (
    g591_p,
    g589_p,
    g587_p
  );


  or

  (
    g592_n,
    g591_p,
    g590_p
  );


  and

  (
    g593_p,
    G1654_o2_n,
    G1696_o2_n
  );


  or

  (
    g593_n,
    G1654_o2_p,
    G1696_o2_p
  );


  and

  (
    g594_p,
    g593_p,
    G1699_o2_n
  );


  or

  (
    g594_n,
    g593_n,
    G1699_o2_p
  );


  and

  (
    g595_p,
    g594_p,
    G1702_o2_n
  );


  or

  (
    g595_n,
    g594_n,
    G1702_o2_p
  );


  and

  (
    g596_p,
    g595_p,
    G1705_o2_n
  );


  or

  (
    g596_n,
    g595_n,
    G1705_o2_p
  );


  and

  (
    g597_p,
    g596_p,
    G1708_o2_n
  );


  or

  (
    g597_n,
    g596_n,
    G1708_o2_p
  );


  and

  (
    g598_p,
    g597_p,
    G1657_o2_n
  );


  or

  (
    g598_n,
    g597_n,
    G1657_o2_p
  );


  and

  (
    g599_p,
    g598_p,
    G1660_o2_n
  );


  or

  (
    g599_n,
    g598_n,
    G1660_o2_p
  );


  and

  (
    g600_p,
    g599_n,
    n1333_lo_n_spl_1
  );


  or

  (
    g600_n,
    g599_p,
    n1333_lo_p_spl_1
  );


  and

  (
    g601_p,
    G248_o2_n_spl_,
    G202_o2_n
  );


  or

  (
    g601_n,
    G248_o2_p_spl_,
    G202_o2_p
  );


  and

  (
    g602_p,
    G1218_o2_p,
    G1203_o2_n
  );


  or

  (
    g602_n,
    G1218_o2_n,
    G1203_o2_p
  );


  and

  (
    g603_p,
    g602_p,
    g601_n
  );


  or

  (
    g603_n,
    g602_n,
    g601_p
  );


  and

  (
    g604_p,
    g603_n_spl_,
    g600_p_spl_
  );


  or

  (
    g604_n,
    g603_p_spl_,
    g600_n_spl_
  );


  and

  (
    g605_p,
    g603_p_spl_,
    g600_n_spl_
  );


  or

  (
    g605_n,
    g603_n_spl_,
    g600_p_spl_
  );


  and

  (
    g606_p,
    g605_n,
    g604_n
  );


  or

  (
    g606_n,
    g605_p,
    g604_p
  );


  and

  (
    g607_p,
    n1297_lo_p,
    n1201_lo_p
  );


  or

  (
    g607_n,
    n1297_lo_n,
    n1201_lo_n
  );


  and

  (
    g608_p,
    g607_n,
    n1333_lo_n_spl_1
  );


  or

  (
    g608_n,
    g607_p,
    n1333_lo_p_spl_1
  );


  and

  (
    g609_p,
    g608_n,
    g606_n
  );


  and

  (
    g610_p,
    g608_p,
    g606_p
  );


  or

  (
    g611_n,
    g610_p,
    g609_p
  );


  and

  (
    g612_p,
    G1130_o2_n,
    G1189_o2_p
  );


  or

  (
    g612_n,
    G1130_o2_p,
    G1189_o2_n
  );


  and

  (
    g613_p,
    G1225_o2_n,
    G1069_o2_p
  );


  or

  (
    g613_n,
    G1225_o2_p,
    G1069_o2_n
  );


  and

  (
    g614_p,
    g613_n,
    g612_n
  );


  or

  (
    g614_n,
    g613_p,
    g612_p
  );


  and

  (
    g615_p,
    n1309_lo_n_spl_1,
    n1249_lo_p
  );


  or

  (
    g615_n,
    n1309_lo_p_spl_1,
    n1249_lo_n
  );


  and

  (
    g616_p,
    g615_p,
    g523_n_spl_1
  );


  or

  (
    g616_n,
    g615_n,
    g523_p_spl_1
  );


  and

  (
    g617_p,
    g616_n_spl_,
    g614_n_spl_
  );


  or

  (
    g617_n,
    g616_p_spl_,
    g614_p_spl_
  );


  and

  (
    g618_p,
    g616_p_spl_,
    g614_p_spl_
  );


  or

  (
    g618_n,
    g616_n_spl_,
    g614_n_spl_
  );


  and

  (
    g619_p,
    g618_n,
    g617_n
  );


  or

  (
    g619_n,
    g618_p,
    g617_p
  );


  and

  (
    g620_p,
    n2180_o2_p_spl_,
    n1874_o2_p_spl_
  );


  or

  (
    g620_n,
    n2180_o2_n_spl_,
    n1874_o2_n_spl_
  );


  and

  (
    g621_p,
    n2180_o2_n_spl_,
    n1874_o2_n_spl_
  );


  or

  (
    g621_n,
    n2180_o2_p_spl_,
    n1874_o2_p_spl_
  );


  and

  (
    g622_p,
    g621_n,
    g620_n
  );


  or

  (
    g622_n,
    g621_p,
    g620_p
  );


  and

  (
    g623_p,
    g622_p,
    g619_n
  );


  and

  (
    g624_p,
    g622_n,
    g619_p
  );


  or

  (
    g625_n,
    g624_p,
    g623_p
  );


  and

  (
    g626_p,
    g625_n,
    g540_n_spl_1
  );


  and

  (
    g627_p,
    G391_o2_p_spl_0,
    n2724_o2_p_spl_
  );


  or

  (
    g627_n,
    G391_o2_n_spl_,
    n2724_o2_n
  );


  and

  (
    g628_p,
    G387_o2_p_spl_0,
    n1162_lo_buf_o2_p_spl_
  );


  or

  (
    g628_n,
    G387_o2_n_spl_,
    n1162_lo_buf_o2_n
  );


  and

  (
    g629_p,
    G1140_o2_p_spl_,
    G212_o2_n_spl_00
  );


  or

  (
    g629_n,
    G1140_o2_n,
    G212_o2_p_spl_00
  );


  and

  (
    g630_p,
    G1178_o2_p_spl_,
    G212_o2_n_spl_00
  );


  or

  (
    g630_n,
    G1178_o2_n,
    G212_o2_p_spl_00
  );


  and

  (
    g631_p,
    n820_inv_n,
    G212_o2_n_spl_01
  );


  or

  (
    g631_n,
    n820_inv_p_spl_,
    G212_o2_p_spl_01
  );


  and

  (
    g632_p,
    G1357_o2_n,
    G212_o2_n_spl_01
  );


  or

  (
    g632_n,
    G1357_o2_p,
    G212_o2_p_spl_01
  );


  and

  (
    g633_p,
    G1369_o2_n,
    G212_o2_n_spl_1
  );


  or

  (
    g633_n,
    G1369_o2_p,
    G212_o2_p_spl_1
  );


  and

  (
    g634_p,
    G1370_o2_p,
    G212_o2_n_spl_1
  );


  or

  (
    g634_n,
    G1370_o2_n,
    G212_o2_p_spl_1
  );


  and

  (
    g635_p,
    G391_o2_p_spl_0,
    n2529_o2_p
  );


  or

  (
    g635_n,
    G391_o2_n_spl_,
    n2529_o2_n
  );


  and

  (
    g636_p,
    G387_o2_p_spl_0,
    n1174_lo_buf_o2_p
  );


  or

  (
    g636_n,
    G387_o2_n_spl_,
    n1174_lo_buf_o2_n
  );


  or

  (
    g637_n,
    G182_o2_p,
    n2497_o2_n
  );


  and

  (
    g638_p,
    n1138_lo_buf_o2_p_spl_,
    G175_o2_n
  );


  or

  (
    g638_n,
    n1138_lo_buf_o2_n,
    G175_o2_p
  );


  and

  (
    g639_p,
    g638_p,
    G241_o2_n_spl_0
  );


  or

  (
    g639_n,
    g638_n,
    G241_o2_p_spl_0
  );


  and

  (
    g640_p,
    n1195_lo_buf_o2_p_spl_,
    G241_o2_n_spl_0
  );


  or

  (
    g640_n,
    n1195_lo_buf_o2_n,
    G241_o2_p_spl_0
  );


  or

  (
    g641_n,
    g633_n_spl_,
    g627_p_spl_
  );


  or

  (
    g642_n,
    g633_p,
    g627_n
  );


  and

  (
    g643_p,
    g642_n,
    g641_n
  );


  or

  (
    g644_n,
    g634_n,
    n1234_lo_buf_o2_p_spl_0
  );


  or

  (
    g645_n,
    g634_p_spl_,
    n1234_lo_buf_o2_n
  );


  and

  (
    g646_p,
    g645_n,
    g644_n
  );


  and

  (
    g647_p,
    g643_p_spl_0,
    g635_p_spl_
  );


  and

  (
    g648_p,
    g646_p_spl_0,
    g636_p_spl_
  );


  and

  (
    g649_p,
    n1306_lo_buf_o2_n_spl_,
    n1282_lo_n
  );


  and

  (
    g650_p,
    g649_p,
    n2498_o2_n_spl_0
  );


  and

  (
    g651_p,
    g650_p,
    g637_n_spl_0
  );


  and

  (
    g652_p,
    n2498_o2_n_spl_0,
    n1318_lo_n
  );


  and

  (
    g653_p,
    g652_p,
    g637_n_spl_0
  );


  or

  (
    g654_n,
    g653_p_spl_,
    g651_p
  );


  and

  (
    g655_p,
    n1306_lo_buf_o2_n_spl_,
    n1294_lo_n
  );


  and

  (
    g656_p,
    g655_p,
    n2498_o2_n_spl_
  );


  and

  (
    g657_p,
    g656_p,
    g637_n_spl_1
  );


  or

  (
    g658_n,
    g657_p,
    g653_p_spl_
  );


  or

  (
    g659_n,
    g643_p_spl_0,
    g635_n
  );


  or

  (
    g660_n,
    g646_p_spl_0,
    g636_n
  );


  or

  (
    g661_n,
    g631_n_spl_,
    g628_p_spl_
  );


  or

  (
    g662_n,
    g631_p,
    g628_n
  );


  and

  (
    g663_p,
    g662_n,
    g661_n
  );


  or

  (
    g664_n,
    g632_n_spl_,
    n1246_lo_buf_o2_p_spl_0
  );


  or

  (
    g665_n,
    g632_p,
    n1246_lo_buf_o2_n
  );


  and

  (
    g666_p,
    g665_n,
    g664_n
  );


  and

  (
    g667_p,
    g666_p,
    g663_p
  );


  or

  (
    g668_n,
    g629_n,
    n1270_lo_buf_o2_p_spl_0
  );


  or

  (
    g669_n,
    g629_p_spl_,
    n1270_lo_buf_o2_n
  );


  and

  (
    g670_p,
    g669_n,
    g668_n
  );


  or

  (
    g671_n,
    g630_n,
    n1258_lo_buf_o2_p_spl_0
  );


  or

  (
    g672_n,
    g630_p_spl_,
    n1258_lo_buf_o2_n
  );


  and

  (
    g673_p,
    g672_n,
    g671_n
  );


  and

  (
    g674_p,
    g673_p,
    g670_p
  );


  and

  (
    g675_p,
    G1112_o2_n,
    G1143_o2_p
  );


  or

  (
    g675_n,
    G1112_o2_p,
    G1143_o2_n
  );


  and

  (
    g676_p,
    g675_n_spl_,
    n949_1_inv_n_spl_
  );


  or

  (
    g676_n,
    g675_p_spl_,
    n949_1_inv_p_spl_0
  );


  and

  (
    g677_p,
    g675_p_spl_,
    n949_1_inv_p_spl_0
  );


  or

  (
    g677_n,
    g675_n_spl_,
    n949_1_inv_n_spl_
  );


  and

  (
    g678_p,
    g677_n,
    g676_n
  );


  or

  (
    g678_n,
    g677_p,
    g676_p
  );


  and

  (
    g679_p,
    n2570_o2_n,
    n2562_o2_p
  );


  and

  (
    g680_p,
    n2570_o2_p,
    n2562_o2_n
  );


  or

  (
    g681_n,
    g680_p,
    g679_p
  );


  and

  (
    g682_p,
    n2645_o2_p,
    n2633_o2_n
  );


  and

  (
    g683_p,
    n2645_o2_n,
    n2633_o2_p
  );


  or

  (
    g684_n,
    g683_p,
    g682_p
  );


  and

  (
    g685_p,
    n2642_o2_p,
    n2639_o2_n
  );


  and

  (
    g686_p,
    n2642_o2_n,
    n2639_o2_p
  );


  or

  (
    g687_n,
    g686_p,
    g685_p
  );


  and

  (
    g688_p,
    g660_n_spl_0,
    g647_p_spl_
  );


  and

  (
    g689_p,
    g688_p,
    g667_p_spl_00
  );


  and

  (
    g690_p,
    g689_p,
    g674_p_spl_00
  );


  and

  (
    g691_p,
    g690_p,
    g658_n_spl_0
  );


  and

  (
    g692_p,
    g659_n_spl_0,
    g648_p_spl_
  );


  and

  (
    g693_p,
    g692_p,
    g667_p_spl_00
  );


  and

  (
    g694_p,
    g693_p,
    g674_p_spl_00
  );


  and

  (
    g695_p,
    g694_p_spl_,
    g654_n_spl_0
  );


  and

  (
    g696_p,
    g694_p_spl_,
    g658_n_spl_0
  );


  and

  (
    g697_p,
    g660_n_spl_0,
    g659_n_spl_0
  );


  and

  (
    g698_p,
    g697_p,
    g667_p_spl_01
  );


  and

  (
    g699_p,
    g698_p,
    g674_p_spl_01
  );


  and

  (
    g700_p,
    g699_p_spl_,
    g654_n_spl_0
  );


  and

  (
    g701_p,
    g699_p_spl_,
    g658_n_spl_1
  );


  and

  (
    g702_p,
    G669_o2_p_spl_,
    G479_o2_p_spl_
  );


  or

  (
    g702_n,
    G669_o2_n_spl_,
    G479_o2_n_spl_
  );


  and

  (
    g703_p,
    G669_o2_n_spl_,
    G479_o2_n_spl_
  );


  or

  (
    g703_n,
    G669_o2_p_spl_,
    G479_o2_p_spl_
  );


  and

  (
    g704_p,
    g703_n,
    g702_n
  );


  or

  (
    g704_n,
    g703_p,
    g702_p
  );


  and

  (
    g705_p,
    g704_n,
    G147_o2_p_spl_0
  );


  and

  (
    g706_p,
    g704_p,
    G147_o2_n_spl_0
  );


  or

  (
    g707_n,
    g706_p,
    g705_p
  );


  and

  (
    g708_p,
    G663_o2_p_spl_,
    G473_o2_p_spl_
  );


  or

  (
    g708_n,
    G663_o2_n_spl_,
    G473_o2_n_spl_
  );


  and

  (
    g709_p,
    G663_o2_n_spl_,
    G473_o2_n_spl_
  );


  or

  (
    g709_n,
    G663_o2_p_spl_,
    G473_o2_p_spl_
  );


  and

  (
    g710_p,
    g709_n,
    g708_n
  );


  or

  (
    g710_n,
    g709_p,
    g708_p
  );


  and

  (
    g711_p,
    g710_n,
    n994_lo_buf_o2_p_spl_0
  );


  and

  (
    g712_p,
    g710_p,
    n994_lo_buf_o2_n_spl_
  );


  or

  (
    g713_n,
    g712_p,
    g711_p
  );


  and

  (
    g714_p,
    G774_o2_p,
    G470_o2_p
  );


  or

  (
    g714_n,
    G774_o2_n,
    G470_o2_n
  );


  and

  (
    g715_p,
    G589_o2_n,
    G660_o2_n
  );


  or

  (
    g715_n,
    G589_o2_p,
    G660_o2_p
  );


  and

  (
    g716_p,
    g715_n,
    g714_n
  );


  or

  (
    g716_n,
    g715_p,
    g714_p
  );


  and

  (
    g717_p,
    g716_n,
    n1006_inv_p_spl_0
  );


  and

  (
    g718_p,
    g716_p,
    n1006_inv_n_spl_
  );


  or

  (
    g719_n,
    g718_p,
    g717_p
  );


  and

  (
    g720_p,
    G782_o2_p,
    G482_o2_p
  );


  or

  (
    g720_n,
    G782_o2_n,
    G482_o2_n
  );


  and

  (
    g721_p,
    G605_o2_n,
    G672_o2_n
  );


  or

  (
    g721_n,
    G605_o2_p,
    G672_o2_p
  );


  and

  (
    g722_p,
    g721_n,
    g720_n
  );


  or

  (
    g722_n,
    g721_p,
    g720_p
  );


  and

  (
    g723_p,
    g722_n,
    G147_o2_p_spl_0
  );


  and

  (
    g724_p,
    g722_p,
    G147_o2_n_spl_0
  );


  or

  (
    g725_n,
    g724_p,
    g723_p
  );


  and

  (
    g726_p,
    n2574_o2_p,
    n2571_o2_p
  );


  and

  (
    g727_p,
    n2574_o2_n,
    n2571_o2_n
  );


  or

  (
    g728_n,
    g727_p,
    g726_p
  );


  or

  (
    g729_n,
    g728_n_spl_,
    n2737_o2_n_spl_
  );


  and

  (
    g730_p,
    n2662_o2_p,
    n2503_o2_p
  );


  and

  (
    g731_p,
    n2662_o2_n,
    n2503_o2_n
  );


  or

  (
    g732_n,
    g731_p,
    g730_p
  );


  or

  (
    g733_n,
    g732_n_spl_,
    G365_o2_p_spl_
  );


  and

  (
    g734_p,
    g732_n_spl_,
    G365_o2_p_spl_
  );


  and

  (
    g735_p,
    g728_n_spl_,
    n2737_o2_n_spl_
  );


  and

  (
    g736_p,
    G788_o2_p,
    G841_o2_n
  );


  or

  (
    g736_n,
    G788_o2_n,
    G841_o2_p
  );


  and

  (
    g737_p,
    g736_n_spl_,
    n2428_o2_p_spl_
  );


  or

  (
    g737_n,
    g736_p_spl_,
    n2428_o2_n_spl_
  );


  and

  (
    g738_p,
    g736_p_spl_,
    n2428_o2_n_spl_
  );


  or

  (
    g738_n,
    g736_n_spl_,
    n2428_o2_p_spl_
  );


  and

  (
    g739_p,
    g738_n,
    g737_n
  );


  or

  (
    g739_n,
    g738_p,
    g737_p
  );


  and

  (
    g740_p,
    g739_p,
    n2575_o2_p
  );


  and

  (
    g741_p,
    g739_n,
    n2575_o2_n
  );


  or

  (
    g742_n,
    g741_p,
    g740_p
  );


  and

  (
    g743_p,
    n2505_o2_n,
    n2444_o2_p
  );


  and

  (
    g744_p,
    n2505_o2_p,
    n2444_o2_n
  );


  or

  (
    g745_n,
    g744_p,
    g743_p
  );


  and

  (
    g746_p,
    g745_n_spl_,
    g742_n_spl_
  );


  or

  (
    g747_n,
    g745_n_spl_,
    g742_n_spl_
  );


  or

  (
    g748_n,
    g701_p_spl_00,
    g696_p_spl_
  );


  or

  (
    g749_n,
    g748_n,
    g691_p_spl_00
  );


  or

  (
    g750_n,
    g749_n,
    g691_p_spl_00
  );


  or

  (
    g751_n,
    g750_n,
    g691_p_spl_01
  );


  or

  (
    g752_n,
    g751_n,
    g691_p_spl_01
  );


  or

  (
    g753_n,
    g752_n,
    g701_p_spl_00
  );


  or

  (
    g754_n,
    g753_n,
    g701_p_spl_01
  );


  or

  (
    g755_n,
    g700_p_spl_00,
    g695_p_spl_00
  );


  or

  (
    g756_n,
    g755_n,
    g695_p_spl_00
  );


  or

  (
    g757_n,
    g756_n,
    g695_p_spl_01
  );


  or

  (
    g758_n,
    g757_n,
    g695_p_spl_01
  );


  and

  (
    g759_p,
    G338_o2_p_spl_,
    n853_inv_p_spl_0
  );


  or

  (
    g759_n,
    G338_o2_n_spl_,
    n853_inv_n_spl_
  );


  and

  (
    g760_p,
    G338_o2_n_spl_,
    n853_inv_n_spl_
  );


  or

  (
    g760_n,
    G338_o2_p_spl_,
    n853_inv_p_spl_0
  );


  and

  (
    g761_p,
    g760_n,
    g759_n
  );


  or

  (
    g761_n,
    g760_p,
    g759_p
  );


  and

  (
    g762_p,
    g761_n,
    n1006_inv_p_spl_0
  );


  and

  (
    g763_p,
    g761_p,
    n1006_inv_n_spl_
  );


  or

  (
    g764_n,
    g763_p,
    g762_p
  );


  and

  (
    g765_p,
    G684_o2_p_spl_,
    G488_o2_p_spl_
  );


  or

  (
    g765_n,
    G684_o2_n_spl_,
    G488_o2_n_spl_
  );


  and

  (
    g766_p,
    G684_o2_n_spl_,
    G488_o2_n_spl_
  );


  or

  (
    g766_n,
    G684_o2_p_spl_,
    G488_o2_p_spl_
  );


  and

  (
    g767_p,
    g766_n,
    g765_n
  );


  or

  (
    g767_n,
    g766_p,
    g765_p
  );


  and

  (
    g768_p,
    g767_n,
    n1066_lo_buf_o2_p_spl_0
  );


  and

  (
    g769_p,
    g767_p,
    n1066_lo_buf_o2_n
  );


  or

  (
    g770_n,
    g769_p,
    g768_p
  );


  and

  (
    g771_p,
    n2747_o2_p_spl_,
    n2744_o2_p_spl_0
  );


  or

  (
    g772_n,
    n2747_o2_p_spl_,
    n2744_o2_p_spl_0
  );


  or

  (
    g773_n,
    n1222_lo_buf_o2_p_spl_,
    n1303_lo_p_spl_0
  );


  or

  (
    g774_n,
    n1210_lo_buf_o2_p_spl_0,
    n1303_lo_p_spl_0
  );


  and

  (
    g775_p,
    G810_o2_p_spl_,
    G419_o2_n_spl_
  );


  or

  (
    g775_n,
    G810_o2_n_spl_,
    G419_o2_p_spl_
  );


  and

  (
    g776_p,
    G810_o2_n_spl_,
    G419_o2_p_spl_
  );


  or

  (
    g776_n,
    G810_o2_p_spl_,
    G419_o2_n_spl_
  );


  and

  (
    g777_p,
    g776_n,
    g775_n
  );


  or

  (
    g777_n,
    g776_p,
    g775_p
  );


  and

  (
    g778_p,
    G813_o2_p_spl_,
    G425_o2_n_spl_
  );


  or

  (
    g778_n,
    G813_o2_n_spl_,
    G425_o2_p_spl_
  );


  and

  (
    g779_p,
    G813_o2_n_spl_,
    G425_o2_p_spl_
  );


  or

  (
    g779_n,
    G813_o2_p_spl_,
    G425_o2_n_spl_
  );


  and

  (
    g780_p,
    g779_n,
    g778_n
  );


  or

  (
    g780_n,
    g779_p,
    g778_p
  );


  and

  (
    g781_p,
    g780_p_spl_,
    g777_n_spl_
  );


  or

  (
    g781_n,
    g780_n_spl_,
    g777_p_spl_
  );


  and

  (
    g782_p,
    g780_n_spl_,
    g777_p_spl_
  );


  or

  (
    g782_n,
    g780_p_spl_,
    g777_n_spl_
  );


  and

  (
    g783_p,
    g782_n,
    g781_n
  );


  or

  (
    g783_n,
    g782_p,
    g781_p
  );


  and

  (
    g784_p,
    n1210_lo_buf_o2_n_spl_,
    n1159_lo_p_spl_
  );


  or

  (
    g784_n,
    n1210_lo_buf_o2_p_spl_0,
    n1159_lo_n
  );


  and

  (
    g785_p,
    g784_p,
    G241_o2_n_spl_1
  );


  or

  (
    g785_n,
    g784_n,
    G241_o2_p_spl_1
  );


  and

  (
    g786_p,
    g785_n,
    g783_n
  );


  and

  (
    g787_p,
    g785_p,
    g783_p
  );


  or

  (
    g788_n,
    g787_p,
    g786_p
  );


  and

  (
    g789_p,
    G898_o2_n_spl_,
    G641_o2_p_spl_
  );


  or

  (
    g789_n,
    G898_o2_p_spl_,
    G641_o2_n_spl_
  );


  and

  (
    g790_p,
    G898_o2_p_spl_,
    G641_o2_n_spl_
  );


  or

  (
    g790_n,
    G898_o2_n_spl_,
    G641_o2_p_spl_
  );


  and

  (
    g791_p,
    g790_n,
    g789_n
  );


  or

  (
    g791_n,
    g790_p,
    g789_p
  );


  and

  (
    g792_p,
    G802_o2_p_spl_,
    G416_o2_n_spl_
  );


  or

  (
    g792_n,
    G802_o2_n_spl_,
    G416_o2_p_spl_
  );


  and

  (
    g793_p,
    G802_o2_n_spl_,
    G416_o2_p_spl_
  );


  or

  (
    g793_n,
    G802_o2_p_spl_,
    G416_o2_n_spl_
  );


  and

  (
    g794_p,
    g793_n,
    g792_n
  );


  or

  (
    g794_n,
    g793_p,
    g792_p
  );


  and

  (
    g795_p,
    g794_p_spl_,
    g791_n_spl_
  );


  or

  (
    g795_n,
    g794_n_spl_,
    g791_p_spl_
  );


  and

  (
    g796_p,
    g794_n_spl_,
    g791_p_spl_
  );


  or

  (
    g796_n,
    g794_p_spl_,
    g791_n_spl_
  );


  and

  (
    g797_p,
    g796_n,
    g795_n
  );


  or

  (
    g797_n,
    g796_p,
    g795_p
  );


  and

  (
    g798_p,
    G500_o2_p_spl_,
    G497_o2_n_spl_
  );


  or

  (
    g798_n,
    G500_o2_n_spl_,
    G497_o2_p_spl_
  );


  and

  (
    g799_p,
    G500_o2_n_spl_,
    G497_o2_p_spl_
  );


  or

  (
    g799_n,
    G500_o2_p_spl_,
    G497_o2_n_spl_
  );


  and

  (
    g800_p,
    g799_n,
    g798_n
  );


  or

  (
    g800_n,
    g799_p,
    g798_p
  );


  and

  (
    g801_p,
    g800_n_spl_,
    n2652_o2_n_spl_
  );


  or

  (
    g801_n,
    g800_p_spl_,
    n2652_o2_p_spl_
  );


  and

  (
    g802_p,
    g800_p_spl_,
    n2652_o2_p_spl_
  );


  or

  (
    g802_n,
    g800_n_spl_,
    n2652_o2_n_spl_
  );


  and

  (
    g803_p,
    g802_n,
    g801_n
  );


  or

  (
    g803_n,
    g802_p,
    g801_p
  );


  and

  (
    g804_p,
    g803_p,
    g797_n
  );


  and

  (
    g805_p,
    g803_n,
    g797_p
  );


  or

  (
    g806_n,
    g805_p,
    g804_p
  );


  and

  (
    g807_p,
    G687_o2_p_spl_,
    G491_o2_p_spl_
  );


  or

  (
    g807_n,
    G687_o2_n_spl_,
    G491_o2_n_spl_
  );


  and

  (
    g808_p,
    G687_o2_n_spl_,
    G491_o2_n_spl_
  );


  or

  (
    g808_n,
    G687_o2_p_spl_,
    G491_o2_p_spl_
  );


  and

  (
    g809_p,
    g808_n,
    g807_n
  );


  or

  (
    g809_n,
    g808_p,
    g807_p
  );


  and

  (
    g810_p,
    g809_n_spl_,
    g640_p_spl_0
  );


  or

  (
    g810_n,
    g809_p_spl_,
    g640_n_spl_
  );


  and

  (
    g811_p,
    g809_p_spl_,
    g640_n_spl_
  );


  or

  (
    g811_n,
    g809_n_spl_,
    g640_p_spl_0
  );


  and

  (
    g812_p,
    g811_n,
    g810_n
  );


  or

  (
    g812_n,
    g811_p,
    g810_p
  );


  and

  (
    g813_p,
    G1169_o2_p,
    G1056_o2_n
  );


  or

  (
    g813_n,
    G1169_o2_n,
    G1056_o2_p
  );


  and

  (
    g814_p,
    G1099_o2_p,
    G1135_o2_n
  );


  or

  (
    g814_n,
    G1099_o2_n,
    G1135_o2_p
  );


  and

  (
    g815_p,
    g814_n,
    g813_n
  );


  or

  (
    g815_n,
    g814_p,
    g813_p
  );


  and

  (
    g816_p,
    g815_n_spl_,
    n748_inv_p_spl_0
  );


  or

  (
    g816_n,
    g815_p_spl_,
    n748_inv_n_spl_
  );


  and

  (
    g817_p,
    g815_p_spl_,
    n748_inv_n_spl_
  );


  or

  (
    g817_n,
    g815_n_spl_,
    n748_inv_p_spl_0
  );


  and

  (
    g818_p,
    g817_n,
    g816_n
  );


  or

  (
    g818_n,
    g817_p,
    g816_p
  );


  and

  (
    g819_p,
    g818_n,
    g812_n
  );


  and

  (
    g820_p,
    g818_p,
    g812_p
  );


  or

  (
    g821_n,
    g820_p,
    g819_p
  );


  and

  (
    g822_p,
    G728_o2_p,
    G901_o2_n
  );


  or

  (
    g822_n,
    G728_o2_n,
    G901_o2_p
  );


  and

  (
    g823_p,
    G942_o2_p,
    G645_o2_n
  );


  or

  (
    g823_n,
    G942_o2_n,
    G645_o2_p
  );


  and

  (
    g824_p,
    g823_n,
    g822_n
  );


  or

  (
    g824_n,
    g823_p,
    g822_p
  );


  and

  (
    g825_p,
    G541_o2_n,
    G816_o2_p
  );


  or

  (
    g825_n,
    G541_o2_p,
    G816_o2_n
  );


  and

  (
    g826_p,
    G856_o2_n,
    G428_o2_p
  );


  or

  (
    g826_n,
    G856_o2_p,
    G428_o2_n
  );


  and

  (
    g827_p,
    g826_n,
    g825_n
  );


  or

  (
    g827_n,
    g826_p,
    g825_p
  );


  and

  (
    g828_p,
    g827_n_spl_,
    g824_p_spl_
  );


  or

  (
    g828_n,
    g827_p_spl_,
    g824_n_spl_
  );


  and

  (
    g829_p,
    g827_p_spl_,
    g824_n_spl_
  );


  or

  (
    g829_n,
    g827_n_spl_,
    g824_p_spl_
  );


  and

  (
    g830_p,
    g829_n,
    g828_n
  );


  or

  (
    g830_n,
    g829_p,
    g828_p
  );


  and

  (
    g831_p,
    n1210_lo_buf_o2_n_spl_,
    n1171_lo_buf_o2_p_spl_
  );


  or

  (
    g831_n,
    n1210_lo_buf_o2_p_spl_1,
    n1171_lo_buf_o2_n
  );


  and

  (
    g832_p,
    g831_p,
    G241_o2_n_spl_1
  );


  or

  (
    g832_n,
    g831_n,
    G241_o2_p_spl_1
  );


  and

  (
    g833_p,
    g832_p_spl_,
    n2744_o2_n_spl_
  );


  or

  (
    g833_n,
    g832_n_spl_,
    n2744_o2_p_spl_1
  );


  and

  (
    g834_p,
    g832_n_spl_,
    n2744_o2_p_spl_1
  );


  or

  (
    g834_n,
    g832_p_spl_,
    n2744_o2_n_spl_
  );


  and

  (
    g835_p,
    g834_n,
    g833_n
  );


  or

  (
    g835_n,
    g834_p,
    g833_p
  );


  or

  (
    g836_n,
    g835_p,
    g830_p
  );


  or

  (
    g837_n,
    g835_n,
    g830_n
  );


  and

  (
    g838_p,
    g837_n,
    g836_n
  );


  and

  (
    g839_p,
    g639_p_spl_0,
    n511_inv_p_spl_0
  );


  or

  (
    g839_n,
    g639_n_spl_,
    n511_inv_n_spl_
  );


  and

  (
    g840_p,
    g639_n_spl_,
    n511_inv_n_spl_
  );


  or

  (
    g840_n,
    g639_p_spl_0,
    n511_inv_p_spl_0
  );


  and

  (
    g841_p,
    g840_n,
    g839_n
  );


  or

  (
    g841_n,
    g840_p,
    g839_p
  );


  and

  (
    g842_p,
    G1154_o2_n,
    G1087_o2_p
  );


  or

  (
    g842_n,
    G1154_o2_p,
    G1087_o2_n
  );


  and

  (
    g843_p,
    G1131_o2_n,
    G1107_o2_p
  );


  or

  (
    g843_n,
    G1131_o2_p,
    G1107_o2_n
  );


  and

  (
    g844_p,
    g843_n,
    g842_n
  );


  or

  (
    g844_n,
    g843_p,
    g842_p
  );


  and

  (
    g845_p,
    g844_n_spl_,
    G987_o2_n_spl_
  );


  or

  (
    g845_n,
    g844_p_spl_,
    G987_o2_p_spl_0
  );


  and

  (
    g846_p,
    g844_p_spl_,
    G987_o2_p_spl_0
  );


  or

  (
    g846_n,
    g844_n_spl_,
    G987_o2_n_spl_
  );


  and

  (
    g847_p,
    g846_n,
    g845_n
  );


  or

  (
    g847_n,
    g846_p,
    g845_p
  );


  or

  (
    g848_n,
    g847_p,
    g841_n
  );


  or

  (
    g849_n,
    g847_n,
    g841_p
  );


  and

  (
    g850_p,
    g849_n,
    g848_n
  );


  and

  (
    g851_p,
    G147_o2_p_spl_1,
    G134_o2_n_spl_0
  );


  and

  (
    g852_p,
    G147_o2_n_spl_1,
    G134_o2_p_spl_0
  );


  or

  (
    g853_n,
    g852_p,
    g851_p
  );


  and

  (
    g854_p,
    G1096_o2_n,
    G1117_o2_n
  );


  or

  (
    g854_n,
    G1096_o2_p,
    G1117_o2_p
  );


  and

  (
    g855_p,
    g854_n_spl_,
    G353_o2_p_spl_0
  );


  or

  (
    g855_n,
    g854_p_spl_,
    G353_o2_n_spl_
  );


  and

  (
    g856_p,
    g854_p_spl_,
    G353_o2_n_spl_
  );


  or

  (
    g856_n,
    g854_n_spl_,
    G353_o2_p_spl_0
  );


  and

  (
    g857_p,
    g856_n,
    g855_n
  );


  or

  (
    g857_n,
    g856_p,
    g855_p
  );


  and

  (
    g858_p,
    g857_p,
    g678_n
  );


  and

  (
    g859_p,
    g857_n,
    g678_p_spl_
  );


  or

  (
    g860_n,
    g859_p,
    g858_p
  );


  or

  (
    g861_n,
    n1096_lo_buf_o2_n,
    n1036_lo_n_spl_0
  );


  or

  (
    g862_n,
    n1096_lo_buf_o2_p_spl_00,
    n1036_lo_p_spl_0
  );


  and

  (
    g863_p,
    g862_n,
    g861_n
  );


  and

  (
    g864_p,
    n1324_lo_n_spl_,
    n1180_lo_p_spl_
  );


  and

  (
    g865_p,
    g707_n_spl_00,
    n1036_lo_n_spl_0
  );


  or

  (
    g866_n,
    g707_n_spl_00,
    n1036_lo_n_spl_
  );


  or

  (
    g867_n,
    g719_n_spl_0,
    g713_n_spl_0
  );


  and

  (
    g868_p,
    g719_n_spl_0,
    g713_n_spl_0
  );


  and

  (
    g869_p,
    n1216_lo_n,
    n1144_lo_p_spl_
  );


  or

  (
    g869_n,
    n1216_lo_p_spl_0,
    n1144_lo_n
  );


  and

  (
    g870_p,
    g869_p,
    n1324_lo_n_spl_
  );


  or

  (
    g870_n,
    g869_n,
    n1324_lo_p_spl_0
  );


  and

  (
    g871_p,
    g870_n,
    G165_o2_p_spl_
  );


  and

  (
    g872_p,
    g870_p,
    G165_o2_n_spl_
  );


  or

  (
    g873_n,
    g872_p,
    g871_p
  );


  and

  (
    g874_p,
    G147_o2_n_spl_1,
    G165_o2_p_spl_
  );


  and

  (
    g875_p,
    G147_o2_p_spl_1,
    G165_o2_n_spl_
  );


  or

  (
    g876_n,
    g875_p,
    g874_p
  );


  and

  (
    g877_p,
    G131_o2_n,
    n1024_lo_p_spl_0
  );


  and

  (
    g878_p,
    G131_o2_p,
    n1024_lo_n_spl_
  );


  or

  (
    g879_n,
    g878_p,
    g877_p
  );


  and

  (
    g880_p,
    G344_o2_p_spl_,
    G134_o2_p_spl_0
  );


  or

  (
    g880_n,
    G344_o2_n_spl_,
    G134_o2_n_spl_0
  );


  and

  (
    g881_p,
    G344_o2_n_spl_,
    G134_o2_n_spl_
  );


  or

  (
    g881_n,
    G344_o2_p_spl_,
    G134_o2_p_spl_
  );


  and

  (
    g882_p,
    g881_n,
    g880_n
  );


  or

  (
    g882_n,
    g881_p,
    g880_p
  );


  and

  (
    g883_p,
    g882_n,
    n994_lo_buf_o2_p_spl_0
  );


  and

  (
    g884_p,
    g882_p,
    n994_lo_buf_o2_n_spl_
  );


  or

  (
    g885_n,
    g884_p,
    g883_p
  );


  and

  (
    g886_p,
    n1024_lo_p_spl_0,
    n976_lo_n
  );


  and

  (
    g887_p,
    n1024_lo_n_spl_,
    n976_lo_p_spl_00
  );


  or

  (
    g888_n,
    g887_p,
    g886_p
  );


  buf

  (
    G1884,
    g365_n
  );


  buf

  (
    G1885,
    g371_n
  );


  buf

  (
    G1886,
    g376_n
  );


  buf

  (
    G1887,
    g382_n
  );


  buf

  (
    G1888,
    g389_n
  );


  buf

  (
    G1889,
    g396_n
  );


  buf

  (
    G1890,
    g402_n
  );


  buf

  (
    G1891,
    g409_n
  );


  buf

  (
    G1892,
    g416_n
  );


  buf

  (
    G1893,
    g422_n
  );


  buf

  (
    G1894,
    g428_n
  );


  buf

  (
    G1895,
    g434_n
  );


  buf

  (
    G1896,
    g441_n
  );


  buf

  (
    G1897,
    g446_n
  );


  buf

  (
    G1898,
    g452_n
  );


  buf

  (
    G1899,
    g458_n
  );


  buf

  (
    G1900,
    g527_p
  );


  buf

  (
    G1901,
    g541_p
  );


  buf

  (
    G1902,
    g554_p
  );


  buf

  (
    G1903,
    g560_p
  );


  buf

  (
    G1904,
    g566_p
  );


  buf

  (
    G1905,
    g573_p
  );


  buf

  (
    G1906,
    g592_n
  );


  buf

  (
    G1907,
    g611_n
  );


  buf

  (
    G1908,
    g626_p
  );


  buf

  (
    n949_li,
    n2290_o2_p
  );


  buf

  (
    n961_li,
    n2190_o2_p
  );


  buf

  (
    n973_li,
    n2212_o2_p
  );


  buf

  (
    n976_li,
    G4_p
  );


  buf

  (
    n985_li,
    n2438_o2_p
  );


  buf

  (
    n997_li,
    n2319_o2_p
  );


  buf

  (
    n1009_li,
    n2213_o2_p
  );


  buf

  (
    n1021_li,
    n2275_o2_p
  );


  buf

  (
    n1024_li,
    G8_p
  );


  buf

  (
    n1033_li,
    n2439_o2_p
  );


  buf

  (
    n1036_li,
    G9_p
  );


  buf

  (
    n1045_li,
    n2440_o2_p
  );


  buf

  (
    n1057_li,
    n2291_o2_p
  );


  buf

  (
    n1069_li,
    n2320_o2_p
  );


  buf

  (
    n1081_li,
    n2214_o2_p
  );


  buf

  (
    n1093_li,
    n2276_o2_p
  );


  buf

  (
    n1105_li,
    n2416_o2_p
  );


  buf

  (
    n1117_li,
    n2191_o2_p
  );


  buf

  (
    n1129_li,
    n2215_o2_p
  );


  buf

  (
    n1132_li,
    G17_p
  );


  buf

  (
    n1141_li,
    n2724_o2_p_spl_
  );


  buf

  (
    n1144_li,
    G18_p
  );


  buf

  (
    n1156_li,
    G19_p
  );


  buf

  (
    n1159_li,
    n1156_lo_p
  );


  buf

  (
    n1165_li,
    n1162_lo_buf_o2_p_spl_
  );


  buf

  (
    n1168_li,
    G20_p
  );


  buf

  (
    n1180_li,
    G21_p
  );


  buf

  (
    n1189_li,
    n2679_o2_p
  );


  buf

  (
    n1192_li,
    G22_p
  );


  buf

  (
    n1201_li,
    n1198_lo_buf_o2_p
  );


  buf

  (
    n1204_li,
    G23_p
  );


  buf

  (
    n1216_li,
    G24_p
  );


  buf

  (
    n1228_li,
    G25_p
  );


  buf

  (
    n1231_li,
    n1228_lo_p
  );


  buf

  (
    n1237_li,
    n1234_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1240_li,
    G26_p
  );


  buf

  (
    n1243_li,
    n1240_lo_p
  );


  buf

  (
    n1249_li,
    n1246_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1252_li,
    G27_p
  );


  buf

  (
    n1255_li,
    n1252_lo_p
  );


  buf

  (
    n1261_li,
    n1258_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1264_li,
    G28_p
  );


  buf

  (
    n1267_li,
    n1264_lo_p
  );


  buf

  (
    n1273_li,
    n1270_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1276_li,
    G29_p
  );


  buf

  (
    n1279_li,
    n1276_lo_p
  );


  buf

  (
    n1282_li,
    n1279_lo_p
  );


  buf

  (
    n1285_li,
    n1282_lo_p_spl_
  );


  buf

  (
    n1288_li,
    G30_p
  );


  buf

  (
    n1291_li,
    n1288_lo_p
  );


  buf

  (
    n1294_li,
    n1291_lo_p
  );


  buf

  (
    n1297_li,
    n1294_lo_p_spl_
  );


  buf

  (
    n1300_li,
    G31_p
  );


  buf

  (
    n1303_li,
    n1300_lo_p
  );


  buf

  (
    n1309_li,
    n1306_lo_buf_o2_p
  );


  buf

  (
    n1312_li,
    G32_p
  );


  buf

  (
    n1315_li,
    n1312_lo_p
  );


  buf

  (
    n1318_li,
    n1315_lo_p
  );


  buf

  (
    n1321_li,
    n1318_lo_p_spl_
  );


  buf

  (
    n1324_li,
    G33_p
  );


  buf

  (
    n1333_li,
    n2498_o2_p_spl_0
  );


  buf

  (
    n1874_i2,
    n304_inv_p
  );


  buf

  (
    n2180_i2,
    G371_o2_p
  );


  buf

  (
    n2372_i2,
    n562_inv_p
  );


  buf

  (
    n2190_i2,
    n2586_o2_p
  );


  buf

  (
    n2191_i2,
    n2587_o2_p
  );


  buf

  (
    n2212_i2,
    n2648_o2_p
  );


  buf

  (
    n2213_i2,
    n2649_o2_p
  );


  buf

  (
    n2214_i2,
    n2650_o2_p
  );


  buf

  (
    n2215_i2,
    n2651_o2_p
  );


  buf

  (
    n2275_i2,
    n2700_o2_p
  );


  buf

  (
    n2276_i2,
    n2701_o2_p
  );


  buf

  (
    n2290_i2,
    n2733_o2_p
  );


  buf

  (
    n2291_i2,
    n2734_o2_p
  );


  buf

  (
    n2681_i2,
    G387_o2_p_spl_
  );


  buf

  (
    n2680_i2,
    G391_o2_p_spl_
  );


  buf

  (
    n2683_i2,
    G1140_o2_p_spl_
  );


  buf

  (
    n2684_i2,
    G1178_o2_p_spl_
  );


  buf

  (
    n2686_i2,
    n820_inv_p_spl_
  );


  buf

  (
    n2319_i2,
    n2754_o2_p
  );


  buf

  (
    n2320_i2,
    n2755_o2_p
  );


  buf

  (
    n2321_i2,
    n511_inv_p_spl_
  );


  buf

  (
    G554_i2,
    g627_p_spl_
  );


  buf

  (
    G557_i2,
    g628_p_spl_
  );


  buf

  (
    G185_i2,
    n1234_lo_buf_o2_p_spl_
  );


  buf

  (
    G188_i2,
    n1246_lo_buf_o2_p_spl_
  );


  buf

  (
    G191_i2,
    n1258_lo_buf_o2_p_spl_
  );


  buf

  (
    G194_i2,
    n1270_lo_buf_o2_p_spl_
  );


  buf

  (
    G1182_i2,
    g629_p_spl_
  );


  buf

  (
    G1222_i2,
    g630_p_spl_
  );


  buf

  (
    G1247_i2,
    g631_n_spl_
  );


  buf

  (
    G1371_i2,
    g632_n_spl_
  );


  buf

  (
    G1383_i2,
    g633_n_spl_
  );


  buf

  (
    G1386_i2,
    g634_p_spl_
  );


  buf

  (
    n2416_i2,
    n1102_lo_buf_o2_p
  );


  buf

  (
    n2428_i2,
    G359_o2_p
  );


  buf

  (
    n2438_i2,
    n982_lo_buf_o2_p
  );


  buf

  (
    n2439_i2,
    n1030_lo_buf_o2_p
  );


  buf

  (
    n2440_i2,
    n1042_lo_buf_o2_p
  );


  buf

  (
    n2444_i2,
    n583_inv_p
  );


  buf

  (
    n2497_i2,
    n1222_lo_buf_o2_p_spl_
  );


  buf

  (
    n2498_i2,
    n1330_lo_buf_o2_p
  );


  buf

  (
    n2503_i2,
    n658_inv_p
  );


  buf

  (
    n2505_i2,
    n661_inv_p
  );


  buf

  (
    n2529_i2,
    n1150_lo_buf_o2_p
  );


  buf

  (
    n2562_i2,
    G356_o2_p
  );


  buf

  (
    n2570_i2,
    G989_o2_p
  );


  buf

  (
    n2571_i2,
    G984_o2_p
  );


  buf

  (
    n2574_i2,
    n685_inv_p
  );


  buf

  (
    n2575_i2,
    n688_inv_p
  );


  buf

  (
    G546_i2,
    g635_p_spl_
  );


  buf

  (
    G550_i2,
    g636_p_spl_
  );


  buf

  (
    n2633_i2,
    G981_o2_p
  );


  buf

  (
    n2639_i2,
    n745_inv_p
  );


  buf

  (
    n2642_i2,
    n748_inv_p_spl_1
  );


  buf

  (
    n2645_i2,
    G1062_o2_p
  );


  buf

  (
    n2679_i2,
    n1186_lo_buf_o2_p
  );


  buf

  (
    n2662_i2,
    G368_o2_p
  );


  buf

  (
    n2724_i2,
    n1138_lo_buf_o2_p_spl_
  );


  not

  (
    G382_i2,
    g637_n_spl_1
  );


  buf

  (
    G199_i2,
    n1282_lo_p_spl_
  );


  buf

  (
    G202_i2,
    n1294_lo_p_spl_
  );


  buf

  (
    G225_i2,
    n1318_lo_p_spl_
  );


  buf

  (
    G248_i2,
    n2498_o2_p_spl_0
  );


  buf

  (
    G260_i2,
    n2498_o2_p_spl_
  );


  buf

  (
    n2716_i2,
    G353_o2_p_spl_
  );


  buf

  (
    n2737_i2,
    n949_1_inv_p_spl_
  );


  buf

  (
    n1174_lo_buf_i2,
    n1171_lo_buf_o2_p_spl_
  );


  buf

  (
    n1198_lo_buf_i2,
    n1195_lo_buf_o2_p_spl_
  );


  buf

  (
    G371_i2,
    g639_p_spl_
  );


  buf

  (
    G1059_i2,
    n748_inv_p_spl_1
  );


  buf

  (
    n2586_i2,
    n958_lo_buf_o2_p
  );


  buf

  (
    n2587_i2,
    n1114_lo_buf_o2_p
  );


  buf

  (
    G1019_i2,
    G987_o2_p_spl_
  );


  buf

  (
    n2648_i2,
    n970_lo_buf_o2_p
  );


  buf

  (
    n2649_i2,
    n1006_lo_buf_o2_p
  );


  buf

  (
    n2650_i2,
    n1078_lo_buf_o2_p
  );


  buf

  (
    n2651_i2,
    n1126_lo_buf_o2_p
  );


  buf

  (
    n2652_i2,
    n766_inv_p
  );


  buf

  (
    G365_i2,
    g640_p_spl_
  );


  buf

  (
    G1496_i2,
    g643_p_spl_
  );


  not

  (
    G1502_i2,
    g646_p_spl_
  );


  buf

  (
    n2700_i2,
    n1018_lo_buf_o2_p
  );


  buf

  (
    n2701_i2,
    n1090_lo_buf_o2_p
  );


  buf

  (
    n2733_i2,
    n946_lo_buf_o2_p
  );


  buf

  (
    n2734_i2,
    n1054_lo_buf_o2_p
  );


  buf

  (
    n2744_i2,
    n970_inv_p
  );


  buf

  (
    n2747_i2,
    G362_o2_p
  );


  buf

  (
    n2754_i2,
    n994_lo_buf_o2_p_spl_1
  );


  buf

  (
    n2755_i2,
    n1066_lo_buf_o2_p_spl_0
  );


  buf

  (
    n2756_i2,
    n1006_inv_p_spl_
  );


  buf

  (
    G1609_i2,
    g647_p_spl_
  );


  buf

  (
    G1625_i2,
    g648_p_spl_
  );


  not

  (
    G738_i2,
    g654_n_spl_
  );


  not

  (
    G755_i2,
    g658_n_spl_1
  );


  not

  (
    G1511_i2,
    g659_n_spl_1
  );


  not

  (
    G1522_i2,
    g659_n_spl_1
  );


  not

  (
    G1538_i2,
    g660_n_spl_1
  );


  not

  (
    G1549_i2,
    g660_n_spl_1
  );


  buf

  (
    G1563_i2,
    g667_p_spl_01
  );


  buf

  (
    G1584_i2,
    g667_p_spl_10
  );


  buf

  (
    G1576_i2,
    g667_p_spl_10
  );


  buf

  (
    G1598_i2,
    g667_p_spl_1
  );


  not

  (
    G1395_i2,
    g674_p_spl_01
  );


  not

  (
    G1410_i2,
    g674_p_spl_10
  );


  not

  (
    G1420_i2,
    g674_p_spl_10
  );


  not

  (
    G1434_i2,
    g674_p_spl_1
  );


  buf

  (
    G1240_i2,
    g678_p_spl_
  );


  buf

  (
    n1162_lo_buf_i2,
    n1159_lo_p_spl_
  );


  buf

  (
    n1102_lo_buf_i2,
    n1096_lo_buf_o2_p_spl_00
  );


  buf

  (
    G359_i2,
    n1066_lo_buf_o2_p_spl_1
  );


  buf

  (
    n982_lo_buf_i2,
    n976_lo_p_spl_00
  );


  buf

  (
    n1030_lo_buf_i2,
    n1024_lo_p_spl_1
  );


  buf

  (
    n1042_lo_buf_i2,
    n1036_lo_p_spl_0
  );


  buf

  (
    G161_i2,
    n1096_lo_buf_o2_p_spl_0
  );


  buf

  (
    G606_i2,
    n2716_o2_p_spl_
  );


  buf

  (
    G1118_i2,
    G1059_o2_p_spl_
  );


  buf

  (
    G1069_i2,
    n460_inv_p_spl_
  );


  buf

  (
    G1145_i2,
    g681_n_spl_
  );


  buf

  (
    G1209_i2,
    g684_n_spl_
  );


  buf

  (
    G1189_i2,
    g687_n_spl_
  );


  buf

  (
    G1699_i2,
    g691_p_spl_10
  );


  buf

  (
    G1702_i2,
    g691_p_spl_10
  );


  buf

  (
    G1705_i2,
    g691_p_spl_11
  );


  buf

  (
    G1708_i2,
    g691_p_spl_11
  );


  buf

  (
    G1684_i2,
    g695_p_spl_10
  );


  buf

  (
    G1687_i2,
    g695_p_spl_10
  );


  buf

  (
    G1690_i2,
    g695_p_spl_11
  );


  buf

  (
    G1693_i2,
    g695_p_spl_11
  );


  buf

  (
    G1696_i2,
    g696_p_spl_
  );


  buf

  (
    G1642_i2,
    g700_p_spl_00
  );


  buf

  (
    G1645_i2,
    g700_p_spl_0
  );


  buf

  (
    G1648_i2,
    g700_p_spl_1
  );


  buf

  (
    G1651_i2,
    g700_p_spl_1
  );


  buf

  (
    G1654_i2,
    g701_p_spl_01
  );


  buf

  (
    G1657_i2,
    g701_p_spl_1
  );


  buf

  (
    G1660_i2,
    g701_p_spl_1
  );


  buf

  (
    n1222_lo_buf_i2,
    n1216_lo_p_spl_0
  );


  buf

  (
    n1330_lo_buf_i2,
    n1324_lo_p_spl_0
  );


  buf

  (
    G123_i2,
    n976_lo_p_spl_01
  );


  buf

  (
    G142_i2,
    n1036_lo_p_spl_1
  );


  buf

  (
    n1306_lo_buf_i2,
    n1303_lo_p_spl_1
  );


  buf

  (
    n1150_lo_buf_i2,
    n1144_lo_p_spl_
  );


  buf

  (
    G175_i2,
    n1216_lo_p_spl_
  );


  buf

  (
    G241_i2,
    n1324_lo_p_spl_
  );


  buf

  (
    G356_i2,
    n1036_lo_p_spl_1
  );


  buf

  (
    G989_i2,
    g707_n_spl_01
  );


  buf

  (
    G984_i2,
    g713_n_spl_
  );


  buf

  (
    G1009_i2,
    g719_n_spl_
  );


  buf

  (
    G1012_i2,
    g725_n_spl_0
  );


  buf

  (
    n958_lo_buf_i2,
    G2_p_spl_00
  );


  buf

  (
    n1114_lo_buf_i2,
    G15_p_spl_00
  );


  buf

  (
    G182_i2,
    n1210_lo_buf_o2_p_spl_1
  );


  not

  (
    G1215_i2,
    g729_n
  );


  not

  (
    G971_i2,
    g733_n
  );


  buf

  (
    G938_i2,
    g734_p
  );


  not

  (
    G1198_i2,
    g735_p
  );


  buf

  (
    G1203_i2,
    g746_p
  );


  buf

  (
    G1218_i2,
    g747_n
  );


  buf

  (
    G785_i2,
    n2716_o2_p_spl_
  );


  buf

  (
    G1168_i2,
    G1059_o2_p_spl_
  );


  buf

  (
    G1130_i2,
    n460_inv_p_spl_
  );


  buf

  (
    G1185_i2,
    g681_n_spl_
  );


  buf

  (
    G1250_i2,
    g684_n_spl_
  );


  buf

  (
    G1225_i2,
    g687_n_spl_
  );


  buf

  (
    G1791_i2,
    g754_n
  );


  buf

  (
    G1788_i2,
    g758_n
  );


  buf

  (
    G981_i2,
    g764_n_spl_0
  );


  buf

  (
    G1031_i2,
    g707_n_spl_01
  );


  buf

  (
    G1015_i2,
    g770_n_spl_0
  );


  buf

  (
    G1062_i2,
    g725_n_spl_0
  );


  buf

  (
    n970_lo_buf_i2,
    G3_p_spl_0
  );


  buf

  (
    n1006_lo_buf_i2,
    G6_p_spl_0
  );


  buf

  (
    n1078_lo_buf_i2,
    G12_p_spl_0
  );


  buf

  (
    n1126_lo_buf_i2,
    G16_p_spl_00
  );


  buf

  (
    G116_i2,
    G2_p_spl_00
  );


  buf

  (
    G165_i2,
    G15_p_spl_00
  );


  buf

  (
    n1234_lo_buf_i2,
    n1231_lo_p
  );


  buf

  (
    n1246_lo_buf_i2,
    n1243_lo_p
  );


  buf

  (
    n1258_lo_buf_i2,
    n1255_lo_p
  );


  buf

  (
    n1270_lo_buf_i2,
    n1267_lo_p
  );


  buf

  (
    G368_i2,
    n1096_lo_buf_o2_p_spl_1
  );


  buf

  (
    G428_i2,
    n976_lo_p_spl_01
  );


  buf

  (
    G212_i2,
    n1303_lo_p_spl_1
  );


  buf

  (
    G841_i2,
    g771_p
  );


  buf

  (
    G788_i2,
    g772_n
  );


  buf

  (
    n1186_lo_buf_i2,
    n1180_lo_p_spl_
  );


  buf

  (
    G391_i2,
    g773_n
  );


  buf

  (
    G387_i2,
    g774_n
  );


  buf

  (
    G645_i2,
    n862_inv_p_spl_0
  );


  buf

  (
    G1140_i2,
    g788_n
  );


  buf

  (
    G1178_i2,
    g806_n
  );


  buf

  (
    G1370_i2,
    g821_n
  );


  buf

  (
    G1205_i2,
    g838_p
  );


  buf

  (
    G1357_i2,
    g850_p
  );


  buf

  (
    G816_i2,
    g853_n_spl_
  );


  buf

  (
    G1369_i2,
    g860_n
  );


  buf

  (
    G901_i2,
    g863_p_spl_0
  );


  buf

  (
    G1056_i2,
    g764_n_spl_0
  );


  buf

  (
    G1107_i2,
    g707_n_spl_1
  );


  buf

  (
    G1087_i2,
    g770_n_spl_0
  );


  buf

  (
    G1135_i2,
    g725_n_spl_1
  );


  buf

  (
    n1018_lo_buf_i2,
    G7_p_spl_0
  );


  buf

  (
    n1090_lo_buf_i2,
    G13_p_spl_0
  );


  buf

  (
    G119_i2,
    G3_p_spl_0
  );


  buf

  (
    G131_i2,
    G6_p_spl_0
  );


  buf

  (
    G154_i2,
    G12_p_spl_0
  );


  buf

  (
    G169_i2,
    G16_p_spl_00
  );


  buf

  (
    G338_i2,
    G2_p_spl_0
  );


  buf

  (
    n1171_lo_buf_i2,
    n1168_lo_p
  );


  buf

  (
    n1195_lo_buf_i2,
    n1192_lo_p
  );


  buf

  (
    G419_i2,
    n853_inv_p_spl_
  );


  buf

  (
    G425_i2,
    n859_inv_p
  );


  buf

  (
    G497_i2,
    n994_lo_buf_o2_p_spl_1
  );


  buf

  (
    G416_i2,
    n1066_lo_buf_o2_p_spl_1
  );


  buf

  (
    G491_i2,
    n976_lo_p_spl_1
  );


  buf

  (
    G500_i2,
    n1024_lo_p_spl_1
  );


  buf

  (
    G353_i2,
    g864_p
  );


  buf

  (
    G641_i2,
    n862_inv_p_spl_0
  );


  buf

  (
    G1117_i2,
    g865_p
  );


  not

  (
    G1096_i2,
    g866_n
  );


  buf

  (
    G1143_i2,
    g867_n
  );


  buf

  (
    G1112_i2,
    g868_p
  );


  buf

  (
    n1138_lo_buf_i2,
    n1132_lo_p
  );


  buf

  (
    n1210_lo_buf_i2,
    n1204_lo_p
  );


  buf

  (
    G687_i2,
    n1096_lo_buf_o2_p_spl_1
  );


  buf

  (
    G541_i2,
    n976_lo_p_spl_1
  );


  buf

  (
    G802_i2,
    g873_n
  );


  buf

  (
    G813_i2,
    g876_n
  );


  buf

  (
    G810_i2,
    g879_n
  );


  buf

  (
    G987_i2,
    g885_n
  );


  buf

  (
    G898_i2,
    g863_p_spl_0
  );


  buf

  (
    n946_lo_buf_i2,
    G1_p_spl_
  );


  buf

  (
    n1054_lo_buf_i2,
    G10_p_spl_
  );


  buf

  (
    G728_i2,
    n862_inv_p_spl_
  );


  buf

  (
    G856_i2,
    g853_n_spl_
  );


  buf

  (
    G831_i2,
    g888_n
  );


  buf

  (
    G942_i2,
    g863_p_spl_
  );


  buf

  (
    G1099_i2,
    g764_n_spl_
  );


  buf

  (
    G1154_i2,
    g707_n_spl_1
  );


  buf

  (
    G1131_i2,
    g770_n_spl_
  );


  buf

  (
    G1169_i2,
    g725_n_spl_1
  );


  buf

  (
    G134_i2,
    G7_p_spl_0
  );


  buf

  (
    G157_i2,
    G13_p_spl_0
  );


  buf

  (
    G470_i2,
    G3_p_spl_1
  );


  buf

  (
    G344_i2,
    G6_p_spl_1
  );


  buf

  (
    G362_i2,
    G12_p_spl_1
  );


  buf

  (
    G482_i2,
    G16_p_spl_0
  );


  buf

  (
    G660_i2,
    G2_p_spl_1
  );


  buf

  (
    G672_i2,
    G15_p_spl_0
  );


  buf

  (
    n1096_lo_buf_i2,
    G14_p
  );


  buf

  (
    G479_i2,
    G16_p_spl_1
  );


  buf

  (
    G669_i2,
    G15_p_spl_1
  );


  buf

  (
    n994_lo_buf_i2,
    G5_p
  );


  buf

  (
    n1066_lo_buf_i2,
    G11_p
  );


  buf

  (
    G112_i2,
    G1_p_spl_
  );


  buf

  (
    G147_i2,
    G10_p_spl_
  );


  buf

  (
    G473_i2,
    G7_p_spl_
  );


  buf

  (
    G488_i2,
    G13_p_spl_
  );


  buf

  (
    G589_i2,
    G3_p_spl_1
  );


  buf

  (
    G663_i2,
    G6_p_spl_1
  );


  buf

  (
    G684_i2,
    G12_p_spl_1
  );


  buf

  (
    G605_i2,
    G16_p_spl_1
  );


  buf

  (
    G774_i2,
    G2_p_spl_1
  );


  buf

  (
    G782_i2,
    G15_p_spl_1
  );


  buf

  (
    G1538_o2_n_spl_,
    G1538_o2_n
  );


  buf

  (
    G1511_o2_n_spl_,
    G1511_o2_n
  );


  buf

  (
    G1538_o2_p_spl_,
    G1538_o2_p
  );


  buf

  (
    G1511_o2_p_spl_,
    G1511_o2_p
  );


  buf

  (
    g359_p_spl_,
    g359_p
  );


  buf

  (
    g359_p_spl_0,
    g359_p_spl_
  );


  buf

  (
    G1584_o2_p_spl_,
    G1584_o2_p
  );


  buf

  (
    G1584_o2_p_spl_0,
    G1584_o2_p_spl_
  );


  buf

  (
    G1584_o2_p_spl_00,
    G1584_o2_p_spl_0
  );


  buf

  (
    G1584_o2_p_spl_01,
    G1584_o2_p_spl_0
  );


  buf

  (
    G1584_o2_p_spl_1,
    G1584_o2_p_spl_
  );


  buf

  (
    g359_n_spl_,
    g359_n
  );


  buf

  (
    g359_n_spl_0,
    g359_n_spl_
  );


  buf

  (
    G1584_o2_n_spl_,
    G1584_o2_n
  );


  buf

  (
    G1584_o2_n_spl_0,
    G1584_o2_n_spl_
  );


  buf

  (
    G1584_o2_n_spl_00,
    G1584_o2_n_spl_0
  );


  buf

  (
    G1584_o2_n_spl_1,
    G1584_o2_n_spl_
  );


  buf

  (
    G1395_o2_n_spl_,
    G1395_o2_n
  );


  buf

  (
    G1395_o2_n_spl_0,
    G1395_o2_n_spl_
  );


  buf

  (
    G1395_o2_n_spl_00,
    G1395_o2_n_spl_0
  );


  buf

  (
    G1395_o2_n_spl_000,
    G1395_o2_n_spl_00
  );


  buf

  (
    G1395_o2_n_spl_001,
    G1395_o2_n_spl_00
  );


  buf

  (
    G1395_o2_n_spl_01,
    G1395_o2_n_spl_0
  );


  buf

  (
    G1395_o2_n_spl_1,
    G1395_o2_n_spl_
  );


  buf

  (
    G1395_o2_n_spl_10,
    G1395_o2_n_spl_1
  );


  buf

  (
    G1395_o2_n_spl_11,
    G1395_o2_n_spl_1
  );


  buf

  (
    G1395_o2_p_spl_,
    G1395_o2_p
  );


  buf

  (
    G1395_o2_p_spl_0,
    G1395_o2_p_spl_
  );


  buf

  (
    G1395_o2_p_spl_1,
    G1395_o2_p_spl_
  );


  buf

  (
    G738_o2_n_spl_,
    G738_o2_n
  );


  buf

  (
    G738_o2_n_spl_0,
    G738_o2_n_spl_
  );


  buf

  (
    G738_o2_n_spl_00,
    G738_o2_n_spl_0
  );


  buf

  (
    G738_o2_n_spl_01,
    G738_o2_n_spl_0
  );


  buf

  (
    G738_o2_n_spl_1,
    G738_o2_n_spl_
  );


  buf

  (
    G738_o2_n_spl_10,
    G738_o2_n_spl_1
  );


  buf

  (
    G738_o2_n_spl_11,
    G738_o2_n_spl_1
  );


  buf

  (
    G738_o2_p_spl_,
    G738_o2_p
  );


  buf

  (
    G738_o2_p_spl_0,
    G738_o2_p_spl_
  );


  buf

  (
    G738_o2_p_spl_00,
    G738_o2_p_spl_0
  );


  buf

  (
    G738_o2_p_spl_01,
    G738_o2_p_spl_0
  );


  buf

  (
    G738_o2_p_spl_1,
    G738_o2_p_spl_
  );


  buf

  (
    G738_o2_p_spl_10,
    G738_o2_p_spl_1
  );


  buf

  (
    G738_o2_p_spl_11,
    G738_o2_p_spl_1
  );


  buf

  (
    G1563_o2_p_spl_,
    G1563_o2_p
  );


  buf

  (
    G1563_o2_p_spl_0,
    G1563_o2_p_spl_
  );


  buf

  (
    G1563_o2_p_spl_00,
    G1563_o2_p_spl_0
  );


  buf

  (
    G1563_o2_p_spl_01,
    G1563_o2_p_spl_0
  );


  buf

  (
    G1563_o2_p_spl_1,
    G1563_o2_p_spl_
  );


  buf

  (
    G1563_o2_n_spl_,
    G1563_o2_n
  );


  buf

  (
    g366_p_spl_,
    g366_p
  );


  buf

  (
    G1420_o2_n_spl_,
    G1420_o2_n
  );


  buf

  (
    G1420_o2_n_spl_0,
    G1420_o2_n_spl_
  );


  buf

  (
    G1420_o2_n_spl_00,
    G1420_o2_n_spl_0
  );


  buf

  (
    G1420_o2_n_spl_01,
    G1420_o2_n_spl_0
  );


  buf

  (
    G1420_o2_n_spl_1,
    G1420_o2_n_spl_
  );


  buf

  (
    G1420_o2_n_spl_10,
    G1420_o2_n_spl_1
  );


  buf

  (
    g366_n_spl_,
    g366_n
  );


  buf

  (
    G1420_o2_p_spl_,
    G1420_o2_p
  );


  buf

  (
    G1420_o2_p_spl_0,
    G1420_o2_p_spl_
  );


  buf

  (
    G1420_o2_p_spl_00,
    G1420_o2_p_spl_0
  );


  buf

  (
    G1420_o2_p_spl_01,
    G1420_o2_p_spl_0
  );


  buf

  (
    G1420_o2_p_spl_1,
    G1420_o2_p_spl_
  );


  buf

  (
    G1410_o2_n_spl_,
    G1410_o2_n
  );


  buf

  (
    G1410_o2_n_spl_0,
    G1410_o2_n_spl_
  );


  buf

  (
    G1410_o2_n_spl_00,
    G1410_o2_n_spl_0
  );


  buf

  (
    G1410_o2_n_spl_1,
    G1410_o2_n_spl_
  );


  buf

  (
    G1410_o2_p_spl_,
    G1410_o2_p
  );


  buf

  (
    G1410_o2_p_spl_0,
    G1410_o2_p_spl_
  );


  buf

  (
    G1410_o2_p_spl_1,
    G1410_o2_p_spl_
  );


  buf

  (
    G1576_o2_p_spl_,
    G1576_o2_p
  );


  buf

  (
    G1576_o2_p_spl_0,
    G1576_o2_p_spl_
  );


  buf

  (
    G1576_o2_p_spl_1,
    G1576_o2_p_spl_
  );


  buf

  (
    G1576_o2_n_spl_,
    G1576_o2_n
  );


  buf

  (
    G1576_o2_n_spl_0,
    G1576_o2_n_spl_
  );


  buf

  (
    G1522_o2_n_spl_,
    G1522_o2_n
  );


  buf

  (
    G1522_o2_n_spl_0,
    G1522_o2_n_spl_
  );


  buf

  (
    G1522_o2_p_spl_,
    G1522_o2_p
  );


  buf

  (
    G1522_o2_p_spl_0,
    G1522_o2_p_spl_
  );


  buf

  (
    G1598_o2_p_spl_,
    G1598_o2_p
  );


  buf

  (
    G1598_o2_p_spl_0,
    G1598_o2_p_spl_
  );


  buf

  (
    G1598_o2_p_spl_1,
    G1598_o2_p_spl_
  );


  buf

  (
    G1598_o2_n_spl_,
    G1598_o2_n
  );


  buf

  (
    G1598_o2_n_spl_0,
    G1598_o2_n_spl_
  );


  buf

  (
    G1598_o2_n_spl_1,
    G1598_o2_n_spl_
  );


  buf

  (
    G755_o2_n_spl_,
    G755_o2_n
  );


  buf

  (
    G755_o2_n_spl_0,
    G755_o2_n_spl_
  );


  buf

  (
    G755_o2_n_spl_00,
    G755_o2_n_spl_0
  );


  buf

  (
    G755_o2_n_spl_01,
    G755_o2_n_spl_0
  );


  buf

  (
    G755_o2_n_spl_1,
    G755_o2_n_spl_
  );


  buf

  (
    G755_o2_n_spl_10,
    G755_o2_n_spl_1
  );


  buf

  (
    G755_o2_n_spl_11,
    G755_o2_n_spl_1
  );


  buf

  (
    G755_o2_p_spl_,
    G755_o2_p
  );


  buf

  (
    G755_o2_p_spl_0,
    G755_o2_p_spl_
  );


  buf

  (
    G755_o2_p_spl_00,
    G755_o2_p_spl_0
  );


  buf

  (
    G755_o2_p_spl_01,
    G755_o2_p_spl_0
  );


  buf

  (
    G755_o2_p_spl_1,
    G755_o2_p_spl_
  );


  buf

  (
    G755_o2_p_spl_10,
    G755_o2_p_spl_1
  );


  buf

  (
    G755_o2_p_spl_11,
    G755_o2_p_spl_1
  );


  buf

  (
    G1549_o2_n_spl_,
    G1549_o2_n
  );


  buf

  (
    G1549_o2_p_spl_,
    G1549_o2_p
  );


  buf

  (
    g390_p_spl_,
    g390_p
  );


  buf

  (
    g390_n_spl_,
    g390_n
  );


  buf

  (
    G1434_o2_n_spl_,
    G1434_o2_n
  );


  buf

  (
    G1434_o2_p_spl_,
    G1434_o2_p
  );


  buf

  (
    G1625_o2_p_spl_,
    G1625_o2_p
  );


  buf

  (
    G1625_o2_p_spl_0,
    G1625_o2_p_spl_
  );


  buf

  (
    G1625_o2_p_spl_1,
    G1625_o2_p_spl_
  );


  buf

  (
    G1625_o2_n_spl_,
    G1625_o2_n
  );


  buf

  (
    g410_p_spl_,
    g410_p
  );


  buf

  (
    g410_p_spl_0,
    g410_p_spl_
  );


  buf

  (
    g410_p_spl_1,
    g410_p_spl_
  );


  buf

  (
    g410_n_spl_,
    g410_n
  );


  buf

  (
    g410_n_spl_0,
    g410_n_spl_
  );


  buf

  (
    g410_n_spl_1,
    g410_n_spl_
  );


  buf

  (
    g423_p_spl_,
    g423_p
  );


  buf

  (
    G1609_o2_p_spl_,
    G1609_o2_p
  );


  buf

  (
    G1609_o2_p_spl_0,
    G1609_o2_p_spl_
  );


  buf

  (
    g435_p_spl_,
    g435_p
  );


  buf

  (
    g435_p_spl_0,
    g435_p_spl_
  );


  buf

  (
    g435_p_spl_1,
    g435_p_spl_
  );


  buf

  (
    g435_n_spl_,
    g435_n
  );


  buf

  (
    g435_n_spl_0,
    g435_n_spl_
  );


  buf

  (
    g436_p_spl_,
    g436_p
  );


  buf

  (
    g436_n_spl_,
    g436_n
  );


  buf

  (
    g484_n_spl_,
    g484_n
  );


  buf

  (
    n1321_lo_p_spl_,
    n1321_lo_p
  );


  buf

  (
    n1321_lo_p_spl_0,
    n1321_lo_p_spl_
  );


  buf

  (
    g488_p_spl_,
    g488_p
  );


  buf

  (
    g488_p_spl_0,
    g488_p_spl_
  );


  buf

  (
    g488_p_spl_00,
    g488_p_spl_0
  );


  buf

  (
    g488_p_spl_01,
    g488_p_spl_0
  );


  buf

  (
    g488_p_spl_1,
    g488_p_spl_
  );


  buf

  (
    g488_p_spl_10,
    g488_p_spl_1
  );


  buf

  (
    g488_p_spl_11,
    g488_p_spl_1
  );


  buf

  (
    g494_p_spl_,
    g494_p
  );


  buf

  (
    g494_p_spl_0,
    g494_p_spl_
  );


  buf

  (
    g498_p_spl_,
    g498_p
  );


  buf

  (
    g523_n_spl_,
    g523_n
  );


  buf

  (
    g523_n_spl_0,
    g523_n_spl_
  );


  buf

  (
    g523_n_spl_00,
    g523_n_spl_0
  );


  buf

  (
    g523_n_spl_01,
    g523_n_spl_0
  );


  buf

  (
    g523_n_spl_1,
    g523_n_spl_
  );


  buf

  (
    g523_n_spl_10,
    g523_n_spl_1
  );


  buf

  (
    g530_n_spl_,
    g530_n
  );


  buf

  (
    n2372_o2_n_spl_,
    n2372_o2_n
  );


  buf

  (
    g530_p_spl_,
    g530_p
  );


  buf

  (
    n2372_o2_p_spl_,
    n2372_o2_p
  );


  buf

  (
    n1309_lo_n_spl_,
    n1309_lo_n
  );


  buf

  (
    n1309_lo_n_spl_0,
    n1309_lo_n_spl_
  );


  buf

  (
    n1309_lo_n_spl_00,
    n1309_lo_n_spl_0
  );


  buf

  (
    n1309_lo_n_spl_01,
    n1309_lo_n_spl_0
  );


  buf

  (
    n1309_lo_n_spl_1,
    n1309_lo_n_spl_
  );


  buf

  (
    n1309_lo_p_spl_,
    n1309_lo_p
  );


  buf

  (
    n1309_lo_p_spl_0,
    n1309_lo_p_spl_
  );


  buf

  (
    n1309_lo_p_spl_00,
    n1309_lo_p_spl_0
  );


  buf

  (
    n1309_lo_p_spl_01,
    n1309_lo_p_spl_0
  );


  buf

  (
    n1309_lo_p_spl_1,
    n1309_lo_p_spl_
  );


  buf

  (
    g523_p_spl_,
    g523_p
  );


  buf

  (
    g523_p_spl_0,
    g523_p_spl_
  );


  buf

  (
    g523_p_spl_00,
    g523_p_spl_0
  );


  buf

  (
    g523_p_spl_01,
    g523_p_spl_0
  );


  buf

  (
    g523_p_spl_1,
    g523_p_spl_
  );


  buf

  (
    n1333_lo_p_spl_,
    n1333_lo_p
  );


  buf

  (
    n1333_lo_p_spl_0,
    n1333_lo_p_spl_
  );


  buf

  (
    n1333_lo_p_spl_00,
    n1333_lo_p_spl_0
  );


  buf

  (
    n1333_lo_p_spl_1,
    n1333_lo_p_spl_
  );


  buf

  (
    g540_n_spl_,
    g540_n
  );


  buf

  (
    g540_n_spl_0,
    g540_n_spl_
  );


  buf

  (
    g540_n_spl_00,
    g540_n_spl_0
  );


  buf

  (
    g540_n_spl_01,
    g540_n_spl_0
  );


  buf

  (
    g540_n_spl_1,
    g540_n_spl_
  );


  buf

  (
    g545_p_spl_,
    g545_p
  );


  buf

  (
    g542_p_spl_,
    g542_p
  );


  buf

  (
    g545_n_spl_,
    g545_n
  );


  buf

  (
    g542_n_spl_,
    g542_n
  );


  buf

  (
    n1333_lo_n_spl_,
    n1333_lo_n
  );


  buf

  (
    n1333_lo_n_spl_0,
    n1333_lo_n_spl_
  );


  buf

  (
    n1333_lo_n_spl_1,
    n1333_lo_n_spl_
  );


  buf

  (
    G248_o2_n_spl_,
    G248_o2_n
  );


  buf

  (
    G248_o2_p_spl_,
    G248_o2_p
  );


  buf

  (
    g584_n_spl_,
    g584_n
  );


  buf

  (
    g581_p_spl_,
    g581_p
  );


  buf

  (
    g584_p_spl_,
    g584_p
  );


  buf

  (
    g581_n_spl_,
    g581_n
  );


  buf

  (
    g603_n_spl_,
    g603_n
  );


  buf

  (
    g600_p_spl_,
    g600_p
  );


  buf

  (
    g603_p_spl_,
    g603_p
  );


  buf

  (
    g600_n_spl_,
    g600_n
  );


  buf

  (
    g616_n_spl_,
    g616_n
  );


  buf

  (
    g614_n_spl_,
    g614_n
  );


  buf

  (
    g616_p_spl_,
    g616_p
  );


  buf

  (
    g614_p_spl_,
    g614_p
  );


  buf

  (
    n2180_o2_p_spl_,
    n2180_o2_p
  );


  buf

  (
    n1874_o2_p_spl_,
    n1874_o2_p
  );


  buf

  (
    n2180_o2_n_spl_,
    n2180_o2_n
  );


  buf

  (
    n1874_o2_n_spl_,
    n1874_o2_n
  );


  buf

  (
    G391_o2_p_spl_,
    G391_o2_p
  );


  buf

  (
    G391_o2_p_spl_0,
    G391_o2_p_spl_
  );


  buf

  (
    n2724_o2_p_spl_,
    n2724_o2_p
  );


  buf

  (
    G391_o2_n_spl_,
    G391_o2_n
  );


  buf

  (
    G387_o2_p_spl_,
    G387_o2_p
  );


  buf

  (
    G387_o2_p_spl_0,
    G387_o2_p_spl_
  );


  buf

  (
    n1162_lo_buf_o2_p_spl_,
    n1162_lo_buf_o2_p
  );


  buf

  (
    G387_o2_n_spl_,
    G387_o2_n
  );


  buf

  (
    G1140_o2_p_spl_,
    G1140_o2_p
  );


  buf

  (
    G212_o2_n_spl_,
    G212_o2_n
  );


  buf

  (
    G212_o2_n_spl_0,
    G212_o2_n_spl_
  );


  buf

  (
    G212_o2_n_spl_00,
    G212_o2_n_spl_0
  );


  buf

  (
    G212_o2_n_spl_01,
    G212_o2_n_spl_0
  );


  buf

  (
    G212_o2_n_spl_1,
    G212_o2_n_spl_
  );


  buf

  (
    G212_o2_p_spl_,
    G212_o2_p
  );


  buf

  (
    G212_o2_p_spl_0,
    G212_o2_p_spl_
  );


  buf

  (
    G212_o2_p_spl_00,
    G212_o2_p_spl_0
  );


  buf

  (
    G212_o2_p_spl_01,
    G212_o2_p_spl_0
  );


  buf

  (
    G212_o2_p_spl_1,
    G212_o2_p_spl_
  );


  buf

  (
    G1178_o2_p_spl_,
    G1178_o2_p
  );


  buf

  (
    n820_inv_p_spl_,
    n820_inv_p
  );


  buf

  (
    n1138_lo_buf_o2_p_spl_,
    n1138_lo_buf_o2_p
  );


  buf

  (
    G241_o2_n_spl_,
    G241_o2_n
  );


  buf

  (
    G241_o2_n_spl_0,
    G241_o2_n_spl_
  );


  buf

  (
    G241_o2_n_spl_1,
    G241_o2_n_spl_
  );


  buf

  (
    G241_o2_p_spl_,
    G241_o2_p
  );


  buf

  (
    G241_o2_p_spl_0,
    G241_o2_p_spl_
  );


  buf

  (
    G241_o2_p_spl_1,
    G241_o2_p_spl_
  );


  buf

  (
    n1195_lo_buf_o2_p_spl_,
    n1195_lo_buf_o2_p
  );


  buf

  (
    g633_n_spl_,
    g633_n
  );


  buf

  (
    g627_p_spl_,
    g627_p
  );


  buf

  (
    n1234_lo_buf_o2_p_spl_,
    n1234_lo_buf_o2_p
  );


  buf

  (
    n1234_lo_buf_o2_p_spl_0,
    n1234_lo_buf_o2_p_spl_
  );


  buf

  (
    g634_p_spl_,
    g634_p
  );


  buf

  (
    g643_p_spl_,
    g643_p
  );


  buf

  (
    g643_p_spl_0,
    g643_p_spl_
  );


  buf

  (
    g635_p_spl_,
    g635_p
  );


  buf

  (
    g646_p_spl_,
    g646_p
  );


  buf

  (
    g646_p_spl_0,
    g646_p_spl_
  );


  buf

  (
    g636_p_spl_,
    g636_p
  );


  buf

  (
    n1306_lo_buf_o2_n_spl_,
    n1306_lo_buf_o2_n
  );


  buf

  (
    n2498_o2_n_spl_,
    n2498_o2_n
  );


  buf

  (
    n2498_o2_n_spl_0,
    n2498_o2_n_spl_
  );


  buf

  (
    g637_n_spl_,
    g637_n
  );


  buf

  (
    g637_n_spl_0,
    g637_n_spl_
  );


  buf

  (
    g637_n_spl_1,
    g637_n_spl_
  );


  buf

  (
    g653_p_spl_,
    g653_p
  );


  buf

  (
    g631_n_spl_,
    g631_n
  );


  buf

  (
    g628_p_spl_,
    g628_p
  );


  buf

  (
    g632_n_spl_,
    g632_n
  );


  buf

  (
    n1246_lo_buf_o2_p_spl_,
    n1246_lo_buf_o2_p
  );


  buf

  (
    n1246_lo_buf_o2_p_spl_0,
    n1246_lo_buf_o2_p_spl_
  );


  buf

  (
    n1270_lo_buf_o2_p_spl_,
    n1270_lo_buf_o2_p
  );


  buf

  (
    n1270_lo_buf_o2_p_spl_0,
    n1270_lo_buf_o2_p_spl_
  );


  buf

  (
    g629_p_spl_,
    g629_p
  );


  buf

  (
    n1258_lo_buf_o2_p_spl_,
    n1258_lo_buf_o2_p
  );


  buf

  (
    n1258_lo_buf_o2_p_spl_0,
    n1258_lo_buf_o2_p_spl_
  );


  buf

  (
    g630_p_spl_,
    g630_p
  );


  buf

  (
    g675_n_spl_,
    g675_n
  );


  buf

  (
    n949_1_inv_n_spl_,
    n949_1_inv_n
  );


  buf

  (
    g675_p_spl_,
    g675_p
  );


  buf

  (
    n949_1_inv_p_spl_,
    n949_1_inv_p
  );


  buf

  (
    n949_1_inv_p_spl_0,
    n949_1_inv_p_spl_
  );


  buf

  (
    g660_n_spl_,
    g660_n
  );


  buf

  (
    g660_n_spl_0,
    g660_n_spl_
  );


  buf

  (
    g660_n_spl_1,
    g660_n_spl_
  );


  buf

  (
    g647_p_spl_,
    g647_p
  );


  buf

  (
    g667_p_spl_,
    g667_p
  );


  buf

  (
    g667_p_spl_0,
    g667_p_spl_
  );


  buf

  (
    g667_p_spl_00,
    g667_p_spl_0
  );


  buf

  (
    g667_p_spl_01,
    g667_p_spl_0
  );


  buf

  (
    g667_p_spl_1,
    g667_p_spl_
  );


  buf

  (
    g667_p_spl_10,
    g667_p_spl_1
  );


  buf

  (
    g674_p_spl_,
    g674_p
  );


  buf

  (
    g674_p_spl_0,
    g674_p_spl_
  );


  buf

  (
    g674_p_spl_00,
    g674_p_spl_0
  );


  buf

  (
    g674_p_spl_01,
    g674_p_spl_0
  );


  buf

  (
    g674_p_spl_1,
    g674_p_spl_
  );


  buf

  (
    g674_p_spl_10,
    g674_p_spl_1
  );


  buf

  (
    g658_n_spl_,
    g658_n
  );


  buf

  (
    g658_n_spl_0,
    g658_n_spl_
  );


  buf

  (
    g658_n_spl_1,
    g658_n_spl_
  );


  buf

  (
    g659_n_spl_,
    g659_n
  );


  buf

  (
    g659_n_spl_0,
    g659_n_spl_
  );


  buf

  (
    g659_n_spl_1,
    g659_n_spl_
  );


  buf

  (
    g648_p_spl_,
    g648_p
  );


  buf

  (
    g694_p_spl_,
    g694_p
  );


  buf

  (
    g654_n_spl_,
    g654_n
  );


  buf

  (
    g654_n_spl_0,
    g654_n_spl_
  );


  buf

  (
    g699_p_spl_,
    g699_p
  );


  buf

  (
    G669_o2_p_spl_,
    G669_o2_p
  );


  buf

  (
    G479_o2_p_spl_,
    G479_o2_p
  );


  buf

  (
    G669_o2_n_spl_,
    G669_o2_n
  );


  buf

  (
    G479_o2_n_spl_,
    G479_o2_n
  );


  buf

  (
    G147_o2_p_spl_,
    G147_o2_p
  );


  buf

  (
    G147_o2_p_spl_0,
    G147_o2_p_spl_
  );


  buf

  (
    G147_o2_p_spl_1,
    G147_o2_p_spl_
  );


  buf

  (
    G147_o2_n_spl_,
    G147_o2_n
  );


  buf

  (
    G147_o2_n_spl_0,
    G147_o2_n_spl_
  );


  buf

  (
    G147_o2_n_spl_1,
    G147_o2_n_spl_
  );


  buf

  (
    G663_o2_p_spl_,
    G663_o2_p
  );


  buf

  (
    G473_o2_p_spl_,
    G473_o2_p
  );


  buf

  (
    G663_o2_n_spl_,
    G663_o2_n
  );


  buf

  (
    G473_o2_n_spl_,
    G473_o2_n
  );


  buf

  (
    n994_lo_buf_o2_p_spl_,
    n994_lo_buf_o2_p
  );


  buf

  (
    n994_lo_buf_o2_p_spl_0,
    n994_lo_buf_o2_p_spl_
  );


  buf

  (
    n994_lo_buf_o2_p_spl_1,
    n994_lo_buf_o2_p_spl_
  );


  buf

  (
    n994_lo_buf_o2_n_spl_,
    n994_lo_buf_o2_n
  );


  buf

  (
    n1006_inv_p_spl_,
    n1006_inv_p
  );


  buf

  (
    n1006_inv_p_spl_0,
    n1006_inv_p_spl_
  );


  buf

  (
    n1006_inv_n_spl_,
    n1006_inv_n
  );


  buf

  (
    g728_n_spl_,
    g728_n
  );


  buf

  (
    n2737_o2_n_spl_,
    n2737_o2_n
  );


  buf

  (
    g732_n_spl_,
    g732_n
  );


  buf

  (
    G365_o2_p_spl_,
    G365_o2_p
  );


  buf

  (
    g736_n_spl_,
    g736_n
  );


  buf

  (
    n2428_o2_p_spl_,
    n2428_o2_p
  );


  buf

  (
    g736_p_spl_,
    g736_p
  );


  buf

  (
    n2428_o2_n_spl_,
    n2428_o2_n
  );


  buf

  (
    g745_n_spl_,
    g745_n
  );


  buf

  (
    g742_n_spl_,
    g742_n
  );


  buf

  (
    g701_p_spl_,
    g701_p
  );


  buf

  (
    g701_p_spl_0,
    g701_p_spl_
  );


  buf

  (
    g701_p_spl_00,
    g701_p_spl_0
  );


  buf

  (
    g701_p_spl_01,
    g701_p_spl_0
  );


  buf

  (
    g701_p_spl_1,
    g701_p_spl_
  );


  buf

  (
    g696_p_spl_,
    g696_p
  );


  buf

  (
    g691_p_spl_,
    g691_p
  );


  buf

  (
    g691_p_spl_0,
    g691_p_spl_
  );


  buf

  (
    g691_p_spl_00,
    g691_p_spl_0
  );


  buf

  (
    g691_p_spl_01,
    g691_p_spl_0
  );


  buf

  (
    g691_p_spl_1,
    g691_p_spl_
  );


  buf

  (
    g691_p_spl_10,
    g691_p_spl_1
  );


  buf

  (
    g691_p_spl_11,
    g691_p_spl_1
  );


  buf

  (
    g700_p_spl_,
    g700_p
  );


  buf

  (
    g700_p_spl_0,
    g700_p_spl_
  );


  buf

  (
    g700_p_spl_00,
    g700_p_spl_0
  );


  buf

  (
    g700_p_spl_1,
    g700_p_spl_
  );


  buf

  (
    g695_p_spl_,
    g695_p
  );


  buf

  (
    g695_p_spl_0,
    g695_p_spl_
  );


  buf

  (
    g695_p_spl_00,
    g695_p_spl_0
  );


  buf

  (
    g695_p_spl_01,
    g695_p_spl_0
  );


  buf

  (
    g695_p_spl_1,
    g695_p_spl_
  );


  buf

  (
    g695_p_spl_10,
    g695_p_spl_1
  );


  buf

  (
    g695_p_spl_11,
    g695_p_spl_1
  );


  buf

  (
    G338_o2_p_spl_,
    G338_o2_p
  );


  buf

  (
    n853_inv_p_spl_,
    n853_inv_p
  );


  buf

  (
    n853_inv_p_spl_0,
    n853_inv_p_spl_
  );


  buf

  (
    G338_o2_n_spl_,
    G338_o2_n
  );


  buf

  (
    n853_inv_n_spl_,
    n853_inv_n
  );


  buf

  (
    G684_o2_p_spl_,
    G684_o2_p
  );


  buf

  (
    G488_o2_p_spl_,
    G488_o2_p
  );


  buf

  (
    G684_o2_n_spl_,
    G684_o2_n
  );


  buf

  (
    G488_o2_n_spl_,
    G488_o2_n
  );


  buf

  (
    n1066_lo_buf_o2_p_spl_,
    n1066_lo_buf_o2_p
  );


  buf

  (
    n1066_lo_buf_o2_p_spl_0,
    n1066_lo_buf_o2_p_spl_
  );


  buf

  (
    n1066_lo_buf_o2_p_spl_1,
    n1066_lo_buf_o2_p_spl_
  );


  buf

  (
    n2747_o2_p_spl_,
    n2747_o2_p
  );


  buf

  (
    n2744_o2_p_spl_,
    n2744_o2_p
  );


  buf

  (
    n2744_o2_p_spl_0,
    n2744_o2_p_spl_
  );


  buf

  (
    n2744_o2_p_spl_1,
    n2744_o2_p_spl_
  );


  buf

  (
    n1222_lo_buf_o2_p_spl_,
    n1222_lo_buf_o2_p
  );


  buf

  (
    n1303_lo_p_spl_,
    n1303_lo_p
  );


  buf

  (
    n1303_lo_p_spl_0,
    n1303_lo_p_spl_
  );


  buf

  (
    n1303_lo_p_spl_1,
    n1303_lo_p_spl_
  );


  buf

  (
    n1210_lo_buf_o2_p_spl_,
    n1210_lo_buf_o2_p
  );


  buf

  (
    n1210_lo_buf_o2_p_spl_0,
    n1210_lo_buf_o2_p_spl_
  );


  buf

  (
    n1210_lo_buf_o2_p_spl_1,
    n1210_lo_buf_o2_p_spl_
  );


  buf

  (
    G810_o2_p_spl_,
    G810_o2_p
  );


  buf

  (
    G419_o2_n_spl_,
    G419_o2_n
  );


  buf

  (
    G810_o2_n_spl_,
    G810_o2_n
  );


  buf

  (
    G419_o2_p_spl_,
    G419_o2_p
  );


  buf

  (
    G813_o2_p_spl_,
    G813_o2_p
  );


  buf

  (
    G425_o2_n_spl_,
    G425_o2_n
  );


  buf

  (
    G813_o2_n_spl_,
    G813_o2_n
  );


  buf

  (
    G425_o2_p_spl_,
    G425_o2_p
  );


  buf

  (
    g780_p_spl_,
    g780_p
  );


  buf

  (
    g777_n_spl_,
    g777_n
  );


  buf

  (
    g780_n_spl_,
    g780_n
  );


  buf

  (
    g777_p_spl_,
    g777_p
  );


  buf

  (
    n1210_lo_buf_o2_n_spl_,
    n1210_lo_buf_o2_n
  );


  buf

  (
    n1159_lo_p_spl_,
    n1159_lo_p
  );


  buf

  (
    G898_o2_n_spl_,
    G898_o2_n
  );


  buf

  (
    G641_o2_p_spl_,
    G641_o2_p
  );


  buf

  (
    G898_o2_p_spl_,
    G898_o2_p
  );


  buf

  (
    G641_o2_n_spl_,
    G641_o2_n
  );


  buf

  (
    G802_o2_p_spl_,
    G802_o2_p
  );


  buf

  (
    G416_o2_n_spl_,
    G416_o2_n
  );


  buf

  (
    G802_o2_n_spl_,
    G802_o2_n
  );


  buf

  (
    G416_o2_p_spl_,
    G416_o2_p
  );


  buf

  (
    g794_p_spl_,
    g794_p
  );


  buf

  (
    g791_n_spl_,
    g791_n
  );


  buf

  (
    g794_n_spl_,
    g794_n
  );


  buf

  (
    g791_p_spl_,
    g791_p
  );


  buf

  (
    G500_o2_p_spl_,
    G500_o2_p
  );


  buf

  (
    G497_o2_n_spl_,
    G497_o2_n
  );


  buf

  (
    G500_o2_n_spl_,
    G500_o2_n
  );


  buf

  (
    G497_o2_p_spl_,
    G497_o2_p
  );


  buf

  (
    g800_n_spl_,
    g800_n
  );


  buf

  (
    n2652_o2_n_spl_,
    n2652_o2_n
  );


  buf

  (
    g800_p_spl_,
    g800_p
  );


  buf

  (
    n2652_o2_p_spl_,
    n2652_o2_p
  );


  buf

  (
    G687_o2_p_spl_,
    G687_o2_p
  );


  buf

  (
    G491_o2_p_spl_,
    G491_o2_p
  );


  buf

  (
    G687_o2_n_spl_,
    G687_o2_n
  );


  buf

  (
    G491_o2_n_spl_,
    G491_o2_n
  );


  buf

  (
    g809_n_spl_,
    g809_n
  );


  buf

  (
    g640_p_spl_,
    g640_p
  );


  buf

  (
    g640_p_spl_0,
    g640_p_spl_
  );


  buf

  (
    g809_p_spl_,
    g809_p
  );


  buf

  (
    g640_n_spl_,
    g640_n
  );


  buf

  (
    g815_n_spl_,
    g815_n
  );


  buf

  (
    n748_inv_p_spl_,
    n748_inv_p
  );


  buf

  (
    n748_inv_p_spl_0,
    n748_inv_p_spl_
  );


  buf

  (
    n748_inv_p_spl_1,
    n748_inv_p_spl_
  );


  buf

  (
    g815_p_spl_,
    g815_p
  );


  buf

  (
    n748_inv_n_spl_,
    n748_inv_n
  );


  buf

  (
    g827_n_spl_,
    g827_n
  );


  buf

  (
    g824_p_spl_,
    g824_p
  );


  buf

  (
    g827_p_spl_,
    g827_p
  );


  buf

  (
    g824_n_spl_,
    g824_n
  );


  buf

  (
    n1171_lo_buf_o2_p_spl_,
    n1171_lo_buf_o2_p
  );


  buf

  (
    g832_p_spl_,
    g832_p
  );


  buf

  (
    n2744_o2_n_spl_,
    n2744_o2_n
  );


  buf

  (
    g832_n_spl_,
    g832_n
  );


  buf

  (
    g639_p_spl_,
    g639_p
  );


  buf

  (
    g639_p_spl_0,
    g639_p_spl_
  );


  buf

  (
    n511_inv_p_spl_,
    n511_inv_p
  );


  buf

  (
    n511_inv_p_spl_0,
    n511_inv_p_spl_
  );


  buf

  (
    g639_n_spl_,
    g639_n
  );


  buf

  (
    n511_inv_n_spl_,
    n511_inv_n
  );


  buf

  (
    g844_n_spl_,
    g844_n
  );


  buf

  (
    G987_o2_n_spl_,
    G987_o2_n
  );


  buf

  (
    g844_p_spl_,
    g844_p
  );


  buf

  (
    G987_o2_p_spl_,
    G987_o2_p
  );


  buf

  (
    G987_o2_p_spl_0,
    G987_o2_p_spl_
  );


  buf

  (
    G134_o2_n_spl_,
    G134_o2_n
  );


  buf

  (
    G134_o2_n_spl_0,
    G134_o2_n_spl_
  );


  buf

  (
    G134_o2_p_spl_,
    G134_o2_p
  );


  buf

  (
    G134_o2_p_spl_0,
    G134_o2_p_spl_
  );


  buf

  (
    g854_n_spl_,
    g854_n
  );


  buf

  (
    G353_o2_p_spl_,
    G353_o2_p
  );


  buf

  (
    G353_o2_p_spl_0,
    G353_o2_p_spl_
  );


  buf

  (
    g854_p_spl_,
    g854_p
  );


  buf

  (
    G353_o2_n_spl_,
    G353_o2_n
  );


  buf

  (
    g678_p_spl_,
    g678_p
  );


  buf

  (
    n1036_lo_n_spl_,
    n1036_lo_n
  );


  buf

  (
    n1036_lo_n_spl_0,
    n1036_lo_n_spl_
  );


  buf

  (
    n1096_lo_buf_o2_p_spl_,
    n1096_lo_buf_o2_p
  );


  buf

  (
    n1096_lo_buf_o2_p_spl_0,
    n1096_lo_buf_o2_p_spl_
  );


  buf

  (
    n1096_lo_buf_o2_p_spl_00,
    n1096_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1096_lo_buf_o2_p_spl_1,
    n1096_lo_buf_o2_p_spl_
  );


  buf

  (
    n1036_lo_p_spl_,
    n1036_lo_p
  );


  buf

  (
    n1036_lo_p_spl_0,
    n1036_lo_p_spl_
  );


  buf

  (
    n1036_lo_p_spl_1,
    n1036_lo_p_spl_
  );


  buf

  (
    n1324_lo_n_spl_,
    n1324_lo_n
  );


  buf

  (
    n1180_lo_p_spl_,
    n1180_lo_p
  );


  buf

  (
    g707_n_spl_,
    g707_n
  );


  buf

  (
    g707_n_spl_0,
    g707_n_spl_
  );


  buf

  (
    g707_n_spl_00,
    g707_n_spl_0
  );


  buf

  (
    g707_n_spl_01,
    g707_n_spl_0
  );


  buf

  (
    g707_n_spl_1,
    g707_n_spl_
  );


  buf

  (
    g719_n_spl_,
    g719_n
  );


  buf

  (
    g719_n_spl_0,
    g719_n_spl_
  );


  buf

  (
    g713_n_spl_,
    g713_n
  );


  buf

  (
    g713_n_spl_0,
    g713_n_spl_
  );


  buf

  (
    n1144_lo_p_spl_,
    n1144_lo_p
  );


  buf

  (
    n1216_lo_p_spl_,
    n1216_lo_p
  );


  buf

  (
    n1216_lo_p_spl_0,
    n1216_lo_p_spl_
  );


  buf

  (
    n1324_lo_p_spl_,
    n1324_lo_p
  );


  buf

  (
    n1324_lo_p_spl_0,
    n1324_lo_p_spl_
  );


  buf

  (
    G165_o2_p_spl_,
    G165_o2_p
  );


  buf

  (
    G165_o2_n_spl_,
    G165_o2_n
  );


  buf

  (
    n1024_lo_p_spl_,
    n1024_lo_p
  );


  buf

  (
    n1024_lo_p_spl_0,
    n1024_lo_p_spl_
  );


  buf

  (
    n1024_lo_p_spl_1,
    n1024_lo_p_spl_
  );


  buf

  (
    n1024_lo_n_spl_,
    n1024_lo_n
  );


  buf

  (
    G344_o2_p_spl_,
    G344_o2_p
  );


  buf

  (
    G344_o2_n_spl_,
    G344_o2_n
  );


  buf

  (
    n976_lo_p_spl_,
    n976_lo_p
  );


  buf

  (
    n976_lo_p_spl_0,
    n976_lo_p_spl_
  );


  buf

  (
    n976_lo_p_spl_00,
    n976_lo_p_spl_0
  );


  buf

  (
    n976_lo_p_spl_01,
    n976_lo_p_spl_0
  );


  buf

  (
    n976_lo_p_spl_1,
    n976_lo_p_spl_
  );


  buf

  (
    n1282_lo_p_spl_,
    n1282_lo_p
  );


  buf

  (
    n1294_lo_p_spl_,
    n1294_lo_p
  );


  buf

  (
    n1318_lo_p_spl_,
    n1318_lo_p
  );


  buf

  (
    n2498_o2_p_spl_,
    n2498_o2_p
  );


  buf

  (
    n2498_o2_p_spl_0,
    n2498_o2_p_spl_
  );


  buf

  (
    n2716_o2_p_spl_,
    n2716_o2_p
  );


  buf

  (
    G1059_o2_p_spl_,
    G1059_o2_p
  );


  buf

  (
    n460_inv_p_spl_,
    n460_inv_p
  );


  buf

  (
    g681_n_spl_,
    g681_n
  );


  buf

  (
    g684_n_spl_,
    g684_n
  );


  buf

  (
    g687_n_spl_,
    g687_n
  );


  buf

  (
    g725_n_spl_,
    g725_n
  );


  buf

  (
    g725_n_spl_0,
    g725_n_spl_
  );


  buf

  (
    g725_n_spl_1,
    g725_n_spl_
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G2_p_spl_0,
    G2_p_spl_
  );


  buf

  (
    G2_p_spl_00,
    G2_p_spl_0
  );


  buf

  (
    G2_p_spl_1,
    G2_p_spl_
  );


  buf

  (
    G15_p_spl_,
    G15_p
  );


  buf

  (
    G15_p_spl_0,
    G15_p_spl_
  );


  buf

  (
    G15_p_spl_00,
    G15_p_spl_0
  );


  buf

  (
    G15_p_spl_1,
    G15_p_spl_
  );


  buf

  (
    g764_n_spl_,
    g764_n
  );


  buf

  (
    g764_n_spl_0,
    g764_n_spl_
  );


  buf

  (
    g770_n_spl_,
    g770_n
  );


  buf

  (
    g770_n_spl_0,
    g770_n_spl_
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G3_p_spl_0,
    G3_p_spl_
  );


  buf

  (
    G3_p_spl_1,
    G3_p_spl_
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G6_p_spl_0,
    G6_p_spl_
  );


  buf

  (
    G6_p_spl_1,
    G6_p_spl_
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G12_p_spl_0,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_1,
    G12_p_spl_
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    G16_p_spl_0,
    G16_p_spl_
  );


  buf

  (
    G16_p_spl_00,
    G16_p_spl_0
  );


  buf

  (
    G16_p_spl_1,
    G16_p_spl_
  );


  buf

  (
    n862_inv_p_spl_,
    n862_inv_p
  );


  buf

  (
    n862_inv_p_spl_0,
    n862_inv_p_spl_
  );


  buf

  (
    g853_n_spl_,
    g853_n
  );


  buf

  (
    g863_p_spl_,
    g863_p
  );


  buf

  (
    g863_p_spl_0,
    g863_p_spl_
  );


  buf

  (
    G7_p_spl_,
    G7_p
  );


  buf

  (
    G7_p_spl_0,
    G7_p_spl_
  );


  buf

  (
    G13_p_spl_,
    G13_p
  );


  buf

  (
    G13_p_spl_0,
    G13_p_spl_
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G10_p_spl_,
    G10_p
  );


endmodule
