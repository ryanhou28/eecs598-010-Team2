



module pe_comb(input_f, input_w, psum_reg, enable, reset, psum_next, output_f);input enable;
  input reset;
  
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  
  
  wire enable;
  
  input [7:0] input_f;
  wire [7:0] input_f;
  
  
  wire [7:0] input_psum;
  
  input [7:0] input_w;
  wire [7:0] input_w;
  
  
  
  wire [7:0] mac1.adder1.A ;
  
  
  
  wire [7:0] mac1.adder1.B ;
  
  
  
  wire [1:0] mac1.adder1.C ;
  
  
  
  wire [7:0] mac1.adder1.SUM ;
  
  
  
  wire [3:0] mac1.adder1.cla1.A ;
  
  
  
  wire [3:0] mac1.adder1.cla1.B ;
  
  
  wire mac1.adder1.cla1.CIN ;
  
  
  
  wire mac1.adder1.cla1.COUT ;
  
  
  
  wire mac1.adder1.cla1.fa0.a ;
  
  
  
  wire mac1.adder1.cla1.fa0.b ;
  
  
  wire mac1.adder1.cla1.fa0.cin ;
  
  
  
  wire mac1.adder1.cla1.fa1.a ;
  
  
  
  wire mac1.adder1.cla1.fa1.b ;
  
  
  
  wire mac1.adder1.cla1.fa2.a ;
  
  
  
  wire mac1.adder1.cla1.fa2.b ;
  
  
  
  wire mac1.adder1.cla1.fa3.a ;
  
  
  
  wire mac1.adder1.cla1.fa3.b ;
  
  
  
  wire [3:0] mac1.adder1.cla2.A ;
  
  
  
  wire [3:0] mac1.adder1.cla2.B ;
  
  
  
  wire mac1.adder1.cla2.CIN ;
  
  
  
  wire mac1.adder1.cla2.COUT ;
  
  
  
  wire mac1.adder1.cla2.fa0.a ;
  
  
  
  wire mac1.adder1.cla2.fa0.b ;
  
  
  
  wire mac1.adder1.cla2.fa0.cin ;
  
  
  
  wire mac1.adder1.cla2.fa1.a ;
  
  
  
  wire mac1.adder1.cla2.fa1.b ;
  
  
  
  wire mac1.adder1.cla2.fa2.a ;
  
  
  
  wire mac1.adder1.cla2.fa2.b ;
  
  
  
  wire mac1.adder1.cla2.fa3.a ;
  
  
  
  wire mac1.adder1.cla2.fa3.b ;
  
  
  
  wire [7:0] mac1.adder1.sat_sum ;
  
  
  
  wire [7:0] mac1.adder_out ;
  
  
  wire [7:0] mac1.input_f ;
  
  
  
  wire [7:0] mac1.input_psum ;
  
  
  wire [7:0] mac1.input_w ;
  
  
  wire [7:0] mac1.mult1.a ;
  
  
  wire [7:0] mac1.mult1.b ;
  
  
  
  wire [7:0] mac1.mult1.product ;
  
  
  
  wire [7:0] mac1.mult_out ;
  
  
  
  wire [7:0] mac1.output_f ;
  
  
  wire [7:0] mac_out;
  
  output [7:0] output_f;
  wire [7:0] output_f;
  
  output [7:0] psum_next;
  wire [7:0] psum_next;
  
  input [7:0] psum_reg;
  wire [7:0] psum_reg;
  
  
  wire [7:0] relu1.input_f ;
  
  
  wire [7:0] relu1.output_f ;
  
  
  wire reset;
  
  
  nand (_0383_, input_f[0], input_f[0]);
  
  
  nand (_0394_, input_f[1], input_f[1]);
  
  
  nand (_0405_, input_f[2], input_f[2]);
  
  
  nand (_0416_, input_f[3], input_f[3]);
  
  
  nand (_0427_, input_f[4], input_f[4]);
  
  
  nand (_0438_, input_f[5], input_f[5]);
  
  
  nand (_0449_, input_f[6], input_f[6]);
  
  
  nand (_0460_, input_f[7], input_f[7]);
  
  
  nand (_0471_, input_w[7], input_w[7]);
  
  
  nand (_0482_, reset, reset);
  
  
  nand (_0493_, enable, enable);
  nand (_0504_, _0482_, psum_reg[7]);
  
  
  nand (_0515_, _0504_, _0504_);
  nand (_0526_, _0493_, _0515_);
  nand (_0537_, input_f[7], input_w[1]);
  nand (_0548_, input_f[7], input_w[0]);
  
  
  nand (_0559_, _0548_, _0548_);
  nand (_0570_, input_w[1], _0559_);
  
  
  nand (_0581_, _0570_, _0570_);
  nand (_0592_, input_f[7], input_w[2]);
  
  
  nand (_0603_, _0592_, _0592_);
  nand (_0614_, _0537_, _0548_);
  
  
  nand (_0625_, _0614_, _0614_);
  nand (_0636_, _0570_, _0614_);
  
  
  nand (_0647_, _0636_, _0636_);
  nand (_0658_, _0592_, _0636_);
  nand (_0669_, _0603_, _0647_);
  nand (_0680_, _0658_, _0669_);
  nand (_0691_, input_w[2], _0581_);
  
  
  nand (_0702_, _0691_, _0691_);
  nand (_0713_, _0592_, _0625_);
  
  
  nand (_0724_, _0713_, _0713_);
  nand (_0735_, _0691_, _0713_);
  
  
  nand (_0746_, _0735_, _0735_);
  nand (_0757_, input_f[5], input_w[5]);
  
  
  nand (_0768_, _0757_, _0757_);
  nand (_0779_, input_f[7], input_w[3]);
  
  
  nand (_0790_, _0779_, _0779_);
  nand (_0801_, input_f[6], input_w[4]);
  
  
  nand (_0812_, _0801_, _0801_);
  nand (_0823_, input_f[7], input_w[4]);
  nand (_0834_, input_f[6], input_w[3]);
  nand (_0845_, _0790_, _0812_);
  nand (_0856_, _0779_, _0801_);
  nand (_0867_, _0845_, _0856_);
  
  
  nand (_0878_, _0867_, _0867_);
  nand (_0889_, _0768_, _0878_);
  nand (_0900_, _0757_, _0867_);
  nand (_0911_, _0889_, _0900_);
  
  
  nand (_0922_, _0911_, _0911_);
  nand (_0933_, _0746_, _0922_);
  nand (_0944_, _0691_, _0933_);
  
  
  nand (_0954_, _0944_, _0944_);
  nand (_0964_, input_w[4], _0790_);
  nand (_0974_, _0779_, _0823_);
  nand (_0984_, _0964_, _0974_);
  
  
  nand (_0009_, _0984_, _0984_);
  nand (_0015_, input_f[6], input_w[5]);
  
  
  nand (_0025_, _0015_, _0015_);
  nand (_0034_, _0009_, _0025_);
  nand (_0037_, _0984_, _0015_);
  nand (_0038_, _0034_, _0037_);
  
  
  nand (_0039_, _0038_, _0038_);
  nand (_0040_, _0746_, _0039_);
  nand (_0041_, _0735_, _0038_);
  nand (_0042_, _0040_, _0041_);
  
  
  nand (_0043_, _0042_, _0042_);
  nand (_0044_, _0944_, _0043_);
  nand (_0045_, input_f[4], input_w[6]);
  
  
  nand (_0046_, _0045_, _0045_);
  nand (_0047_, _0416_, input_w[7]);
  
  
  nand (_0048_, _0047_, _0047_);
  nand (_0049_, _0046_, _0048_);
  
  
  nand (_0050_, _0049_, _0049_);
  nand (_0051_, _0845_, _0889_);
  
  
  nand (_0052_, _0051_, _0051_);
  nand (_0053_, input_f[5], input_w[6]);
  
  
  nand (_0054_, _0053_, _0053_);
  nand (_0055_, _0427_, input_w[7]);
  
  
  nand (_0056_, _0055_, _0055_);
  nand (_0057_, _0054_, _0056_);
  
  
  nand (_0058_, _0057_, _0057_);
  nand (_0059_, _0053_, _0055_);
  nand (_0060_, _0057_, _0059_);
  
  
  nand (_0061_, _0060_, _0060_);
  nand (_0062_, _0051_, _0061_);
  nand (_0063_, _0052_, _0060_);
  nand (_0064_, _0062_, _0063_);
  
  
  nand (_0065_, _0064_, _0064_);
  nand (_0066_, _0050_, _0065_);
  nand (_0067_, _0049_, _0064_);
  nand (_0068_, _0066_, _0067_);
  
  
  nand (_0069_, _0068_, _0068_);
  nand (_0070_, _0954_, _0042_);
  nand (_0071_, _0044_, _0070_);
  
  
  nand (_0072_, _0071_, _0071_);
  nand (_0073_, _0069_, _0072_);
  nand (_0074_, _0044_, _0073_);
  
  
  nand (_0075_, _0074_, _0074_);
  nand (_0076_, _0964_, _0034_);
  
  
  nand (_0077_, _0076_, _0076_);
  nand (_0078_, input_f[6], input_w[6]);
  
  
  nand (_0079_, _0078_, _0078_);
  nand (_0080_, _0438_, input_w[7]);
  
  
  nand (_0081_, _0080_, _0080_);
  nand (_0082_, _0079_, _0081_);
  
  
  nand (_0083_, _0082_, _0082_);
  nand (_0084_, _0078_, _0080_);
  nand (_0085_, _0082_, _0084_);
  
  
  nand (_0086_, _0085_, _0085_);
  nand (_0087_, _0076_, _0086_);
  nand (_0088_, _0077_, _0085_);
  nand (_0089_, _0087_, _0088_);
  
  
  nand (_0090_, _0089_, _0089_);
  nand (_0091_, _0058_, _0090_);
  nand (_0092_, _0057_, _0089_);
  nand (_0093_, _0091_, _0092_);
  
  
  nand (_0094_, _0093_, _0093_);
  nand (_0095_, input_f[7], input_w[5]);
  
  
  nand (_0096_, _0095_, _0095_);
  nand (_0097_, _0009_, _0096_);
  nand (_0098_, _0984_, _0095_);
  nand (_0099_, _0097_, _0098_);
  
  
  nand (_0100_, _0099_, _0099_);
  nand (_0101_, _0735_, _0099_);
  nand (_0102_, _0746_, _0100_);
  nand (_0103_, _0101_, _0102_);
  
  
  nand (_0104_, _0103_, _0103_);
  nand (_0105_, _0691_, _0040_);
  
  
  nand (_0106_, _0105_, _0105_);
  nand (_0107_, _0104_, _0105_);
  nand (_0108_, _0103_, _0106_);
  nand (_0109_, _0107_, _0108_);
  
  
  nand (_0110_, _0109_, _0109_);
  nand (_0111_, _0094_, _0110_);
  nand (_0112_, _0093_, _0109_);
  nand (_0113_, _0111_, _0112_);
  
  
  nand (_0114_, _0113_, _0113_);
  nand (_0115_, _0074_, _0114_);
  nand (_0116_, _0062_, _0066_);
  
  
  nand (_0117_, _0116_, _0116_);
  nand (_0118_, _0075_, _0113_);
  nand (_0119_, _0115_, _0118_);
  
  
  nand (_0120_, _0119_, _0119_);
  nand (_0121_, _0116_, _0120_);
  nand (_0122_, _0115_, _0121_);
  
  
  nand (_0123_, _0122_, _0122_);
  nand (_0124_, _0087_, _0091_);
  
  
  nand (_0125_, _0124_, _0124_);
  nand (_0126_, _0107_, _0111_);
  
  
  nand (_0127_, _0126_, _0126_);
  nand (_0128_, _0702_, _0100_);
  nand (_0129_, _0724_, _0099_);
  nand (_0130_, _0128_, _0129_);
  
  
  nand (_0131_, _0130_, _0130_);
  nand (_0132_, _0964_, _0097_);
  
  
  nand (_0133_, _0132_, _0132_);
  nand (_0134_, input_f[7], input_w[6]);
  
  
  nand (_0135_, _0134_, _0134_);
  nand (_0136_, _0449_, input_w[7]);
  
  
  nand (_0137_, _0136_, _0136_);
  nand (_0138_, _0135_, _0137_);
  nand (_0139_, _0134_, _0136_);
  nand (_0140_, _0138_, _0139_);
  
  
  nand (_0141_, _0140_, _0140_);
  nand (_0142_, _0132_, _0141_);
  nand (_0143_, _0133_, _0140_);
  nand (_0144_, _0142_, _0143_);
  
  
  nand (_0145_, _0144_, _0144_);
  nand (_0146_, _0083_, _0145_);
  nand (_0147_, _0082_, _0144_);
  nand (_0148_, _0146_, _0147_);
  
  
  nand (_0149_, _0148_, _0148_);
  nand (_0150_, _0131_, _0149_);
  nand (_0151_, _0130_, _0148_);
  nand (_0152_, _0150_, _0151_);
  
  
  nand (_0153_, _0152_, _0152_);
  nand (_0154_, _0126_, _0153_);
  nand (_0155_, _0127_, _0152_);
  nand (_0156_, _0154_, _0155_);
  
  
  nand (_0157_, _0156_, _0156_);
  nand (_0158_, _0124_, _0157_);
  nand (_0159_, _0125_, _0156_);
  nand (_0160_, _0158_, _0159_);
  
  
  nand (_0161_, _0160_, _0160_);
  nand (_0162_, _0122_, _0161_);
  nand (_0163_, input_f[4], input_w[5]);
  
  
  nand (_0164_, _0163_, _0163_);
  nand (_0165_, input_f[5], input_w[4]);
  nand (_0166_, input_f[5], input_w[3]);
  
  
  nand (_0167_, _0166_, _0166_);
  nand (_0168_, _0812_, _0167_);
  nand (_0169_, _0834_, _0165_);
  nand (_0170_, _0168_, _0169_);
  
  
  nand (_0171_, _0170_, _0170_);
  nand (_0172_, _0164_, _0171_);
  nand (_0173_, _0163_, _0170_);
  nand (_0174_, _0172_, _0173_);
  
  
  nand (_0175_, _0174_, _0174_);
  nand (_0176_, input_f[6], input_w[2]);
  
  
  nand (_0177_, _0176_, _0176_);
  nand (_0178_, _0647_, _0177_);
  nand (_0179_, _0570_, _0178_);
  
  
  nand (_0180_, _0179_, _0179_);
  nand (_0181_, _0680_, _0180_);
  nand (_0182_, _0691_, _0181_);
  
  
  nand (_0183_, _0182_, _0182_);
  nand (_0184_, _0175_, _0183_);
  nand (_0185_, _0691_, _0184_);
  
  
  nand (_0186_, _0185_, _0185_);
  nand (_0187_, _0735_, _0911_);
  nand (_0188_, _0933_, _0187_);
  
  
  nand (_0189_, _0188_, _0188_);
  nand (_0190_, _0185_, _0189_);
  nand (_0191_, input_f[3], input_w[6]);
  
  
  nand (_0192_, _0191_, _0191_);
  nand (_0193_, _0405_, input_w[7]);
  
  
  nand (_0194_, _0193_, _0193_);
  nand (_0195_, _0192_, _0194_);
  
  
  nand (_0196_, _0195_, _0195_);
  nand (_0197_, _0168_, _0172_);
  
  
  nand (_0198_, _0197_, _0197_);
  nand (_0199_, _0045_, _0047_);
  nand (_0200_, _0049_, _0199_);
  
  
  nand (_0201_, _0200_, _0200_);
  nand (_0202_, _0197_, _0201_);
  nand (_0203_, _0198_, _0200_);
  nand (_0204_, _0202_, _0203_);
  
  
  nand (_0205_, _0204_, _0204_);
  nand (_0206_, _0196_, _0205_);
  nand (_0207_, _0195_, _0204_);
  nand (_0208_, _0206_, _0207_);
  
  
  nand (_0209_, _0208_, _0208_);
  nand (_0210_, _0186_, _0188_);
  nand (_0211_, _0190_, _0210_);
  
  
  nand (_0212_, _0211_, _0211_);
  nand (_0213_, _0209_, _0212_);
  nand (_0214_, _0190_, _0213_);
  
  
  nand (_0215_, _0214_, _0214_);
  nand (_0216_, _0068_, _0071_);
  nand (_0217_, _0073_, _0216_);
  
  
  nand (_0218_, _0217_, _0217_);
  nand (_0219_, _0214_, _0218_);
  nand (_0220_, _0202_, _0206_);
  
  
  nand (_0221_, _0220_, _0220_);
  nand (_0222_, _0215_, _0217_);
  nand (_0223_, _0219_, _0222_);
  
  
  nand (_0224_, _0223_, _0223_);
  nand (_0225_, _0220_, _0224_);
  nand (_0226_, _0219_, _0225_);
  
  
  nand (_0227_, _0226_, _0226_);
  nand (_0228_, _0117_, _0119_);
  nand (_0229_, _0121_, _0228_);
  
  
  nand (_0230_, _0229_, _0229_);
  nand (_0231_, _0226_, _0230_);
  nand (_0232_, input_w[7], _0559_);
  nand (_0233_, input_f[6], input_w[1]);
  
  
  nand (_0234_, _0233_, _0233_);
  nand (_0235_, _0471_, _0548_);
  nand (_0236_, _0232_, _0235_);
  
  
  nand (_0237_, _0236_, _0236_);
  nand (_0238_, _0234_, _0237_);
  nand (_0239_, _0232_, _0238_);
  
  
  nand (_0240_, _0239_, _0239_);
  nand (_0241_, _0636_, _0176_);
  nand (_0242_, _0178_, _0241_);
  
  
  nand (_0243_, _0242_, _0242_);
  nand (_0244_, _0239_, _0243_);
  nand (_0245_, input_f[3], input_w[5]);
  
  
  nand (_0246_, _0245_, _0245_);
  nand (_0247_, input_f[4], input_w[4]);
  
  
  nand (_0248_, _0247_, _0247_);
  nand (_0249_, input_f[4], input_w[3]);
  nand (_0250_, _0167_, _0248_);
  nand (_0251_, _0166_, _0247_);
  nand (_0252_, _0250_, _0251_);
  
  
  nand (_0253_, _0252_, _0252_);
  nand (_0254_, _0246_, _0253_);
  nand (_0255_, _0245_, _0252_);
  nand (_0256_, _0254_, _0255_);
  
  
  nand (_0257_, _0256_, _0256_);
  nand (_0258_, _0240_, _0242_);
  nand (_0259_, _0244_, _0258_);
  
  
  nand (_0260_, _0259_, _0259_);
  nand (_0261_, _0257_, _0260_);
  nand (_0262_, _0244_, _0261_);
  
  
  nand (_0263_, _0262_, _0262_);
  nand (_0264_, _0174_, _0182_);
  nand (_0265_, _0184_, _0264_);
  
  
  nand (_0266_, _0265_, _0265_);
  nand (_0267_, _0262_, _0266_);
  nand (_0268_, input_f[2], input_w[6]);
  
  
  nand (_0269_, _0268_, _0268_);
  nand (_0270_, _0394_, input_w[7]);
  
  
  nand (_0271_, _0270_, _0270_);
  nand (_0272_, _0269_, _0271_);
  
  
  nand (_0273_, _0272_, _0272_);
  nand (_0274_, _0250_, _0254_);
  
  
  nand (_0275_, _0274_, _0274_);
  nand (_0276_, _0191_, _0193_);
  nand (_0277_, _0195_, _0276_);
  
  
  nand (_0278_, _0277_, _0277_);
  nand (_0279_, _0274_, _0278_);
  nand (_0280_, _0275_, _0277_);
  nand (_0281_, _0279_, _0280_);
  
  
  nand (_0282_, _0281_, _0281_);
  nand (_0283_, _0273_, _0282_);
  nand (_0284_, _0272_, _0281_);
  nand (_0285_, _0283_, _0284_);
  
  
  nand (_0286_, _0285_, _0285_);
  nand (_0287_, _0263_, _0265_);
  nand (_0288_, _0267_, _0287_);
  
  
  nand (_0289_, _0288_, _0288_);
  nand (_0290_, _0286_, _0289_);
  nand (_0291_, _0267_, _0290_);
  
  
  nand (_0292_, _0291_, _0291_);
  nand (_0293_, _0208_, _0211_);
  nand (_0294_, _0213_, _0293_);
  
  
  nand (_0295_, _0294_, _0294_);
  nand (_0296_, _0291_, _0295_);
  nand (_0297_, _0279_, _0283_);
  
  
  nand (_0298_, _0297_, _0297_);
  nand (_0299_, _0292_, _0294_);
  nand (_0300_, _0296_, _0299_);
  
  
  nand (_0301_, _0300_, _0300_);
  nand (_0302_, _0297_, _0301_);
  nand (_0303_, _0296_, _0302_);
  
  
  nand (_0304_, _0303_, _0303_);
  nand (_0305_, _0221_, _0223_);
  nand (_0306_, _0225_, _0305_);
  
  
  nand (_0307_, _0306_, _0306_);
  nand (_0308_, _0303_, _0307_);
  nand (_0309_, _0304_, _0306_);
  nand (_0310_, _0308_, _0309_);
  
  
  nand (_0311_, _0310_, _0310_);
  nand (_0312_, input_f[6], input_w[0]);
  nand (_0313_, input_f[5], input_w[1]);
  nand (_0314_, input_f[5], input_w[0]);
  
  
  nand (_0315_, _0314_, _0314_);
  nand (_0316_, _0234_, _0315_);
  nand (_0317_, input_f[4], input_w[2]);
  
  
  nand (_0318_, _0317_, _0317_);
  nand (_0319_, _0312_, _0313_);
  nand (_0320_, _0316_, _0319_);
  
  
  nand (_0321_, _0320_, _0320_);
  nand (_0322_, _0318_, _0321_);
  nand (_0323_, _0316_, _0322_);
  
  
  nand (_0324_, _0323_, _0323_);
  nand (_0325_, _0233_, _0236_);
  nand (_0326_, _0238_, _0325_);
  
  
  nand (_0327_, _0326_, _0326_);
  nand (_0328_, _0323_, _0327_);
  nand (_0329_, _0324_, _0326_);
  nand (_0330_, _0328_, _0329_);
  
  
  nand (_0331_, _0330_, _0330_);
  nand (_0332_, input_f[3], input_w[4]);
  
  
  nand (_0333_, _0332_, _0332_);
  nand (_0334_, input_f[5], input_w[2]);
  nand (_0335_, _0167_, _0318_);
  nand (_0336_, _0249_, _0334_);
  nand (_0337_, _0335_, _0336_);
  
  
  nand (_0338_, _0337_, _0337_);
  nand (_0339_, _0333_, _0338_);
  nand (_0340_, _0332_, _0337_);
  nand (_0341_, _0339_, _0340_);
  
  
  nand (_0342_, _0341_, _0341_);
  nand (_0343_, _0331_, _0342_);
  nand (_0344_, _0328_, _0343_);
  
  
  nand (_0345_, _0344_, _0344_);
  nand (_0346_, _0256_, _0259_);
  nand (_0347_, _0261_, _0346_);
  
  
  nand (_0348_, _0347_, _0347_);
  nand (_0349_, _0344_, _0348_);
  nand (_0350_, input_f[2], input_w[5]);
  nand (_0351_, input_f[1], input_w[6]);
  nand (_0352_, input_f[1], input_w[5]);
  
  
  nand (_0353_, _0352_, _0352_);
  nand (_0354_, _0269_, _0353_);
  nand (_0355_, _0383_, input_w[7]);
  
  
  nand (_0356_, _0355_, _0355_);
  nand (_0357_, _0350_, _0351_);
  nand (_0358_, _0354_, _0357_);
  
  
  nand (_0359_, _0358_, _0358_);
  nand (_0360_, _0356_, _0359_);
  nand (_0361_, _0354_, _0360_);
  
  
  nand (_0362_, _0361_, _0361_);
  nand (_0363_, _0335_, _0339_);
  
  
  nand (_0364_, _0363_, _0363_);
  nand (_0365_, _0268_, _0270_);
  nand (_0366_, _0272_, _0365_);
  
  
  nand (_0367_, _0366_, _0366_);
  nand (_0368_, _0363_, _0367_);
  nand (_0369_, _0364_, _0366_);
  nand (_0370_, _0368_, _0369_);
  
  
  nand (_0371_, _0370_, _0370_);
  nand (_0372_, _0361_, _0371_);
  nand (_0373_, _0362_, _0370_);
  nand (_0374_, _0372_, _0373_);
  
  
  nand (_0375_, _0374_, _0374_);
  nand (_0376_, _0345_, _0347_);
  nand (_0377_, _0349_, _0376_);
  
  
  nand (_0378_, _0377_, _0377_);
  nand (_0379_, _0375_, _0378_);
  nand (_0380_, _0349_, _0379_);
  
  
  nand (_0381_, _0380_, _0380_);
  nand (_0382_, _0285_, _0288_);
  nand (_0384_, _0290_, _0382_);
  
  
  nand (_0385_, _0384_, _0384_);
  nand (_0386_, _0380_, _0385_);
  nand (_0387_, _0368_, _0372_);
  
  
  nand (_0388_, _0387_, _0387_);
  nand (_0389_, _0381_, _0384_);
  nand (_0390_, _0386_, _0389_);
  
  
  nand (_0391_, _0390_, _0390_);
  nand (_0392_, _0387_, _0391_);
  nand (_0393_, _0386_, _0392_);
  
  
  nand (_0395_, _0393_, _0393_);
  nand (_0396_, _0298_, _0300_);
  nand (_0397_, _0302_, _0396_);
  
  
  nand (_0398_, _0397_, _0397_);
  nand (_0399_, _0393_, _0398_);
  nand (_0400_, _0395_, _0397_);
  nand (_0401_, _0399_, _0400_);
  
  
  nand (_0402_, _0401_, _0401_);
  nand (_0403_, input_f[4], input_w[1]);
  
  
  nand (_0404_, _0403_, _0403_);
  nand (_0406_, input_f[4], input_w[0]);
  
  
  nand (_0407_, _0406_, _0406_);
  nand (_0408_, _0315_, _0404_);
  nand (_0409_, input_f[3], input_w[2]);
  
  
  nand (_0410_, _0409_, _0409_);
  nand (_0411_, _0314_, _0403_);
  nand (_0412_, _0408_, _0411_);
  
  
  nand (_0413_, _0412_, _0412_);
  nand (_0414_, _0410_, _0413_);
  nand (_0415_, _0408_, _0414_);
  
  
  nand (_0417_, _0415_, _0415_);
  nand (_0418_, _0317_, _0320_);
  nand (_0419_, _0322_, _0418_);
  
  
  nand (_0420_, _0419_, _0419_);
  nand (_0421_, _0415_, _0420_);
  nand (_0422_, input_f[3], input_w[3]);
  nand (_0423_, input_f[2], input_w[4]);
  nand (_0424_, input_f[2], input_w[3]);
  
  
  nand (_0425_, _0424_, _0424_);
  nand (_0426_, _0333_, _0425_);
  nand (_0428_, _0422_, _0423_);
  nand (_0429_, _0426_, _0428_);
  
  
  nand (_0430_, _0429_, _0429_);
  nand (_0431_, _0353_, _0430_);
  nand (_0432_, _0352_, _0429_);
  nand (_0433_, _0431_, _0432_);
  
  
  nand (_0434_, _0433_, _0433_);
  nand (_0435_, _0417_, _0419_);
  nand (_0436_, _0421_, _0435_);
  
  
  nand (_0437_, _0436_, _0436_);
  nand (_0439_, _0434_, _0437_);
  nand (_0440_, _0421_, _0439_);
  
  
  nand (_0441_, _0440_, _0440_);
  nand (_0442_, _0330_, _0341_);
  nand (_0443_, _0343_, _0442_);
  
  
  nand (_0444_, _0443_, _0443_);
  nand (_0445_, _0440_, _0444_);
  nand (_0446_, _0441_, _0443_);
  nand (_0447_, _0445_, _0446_);
  
  
  nand (_0448_, _0447_, _0447_);
  nand (_0450_, _0426_, _0431_);
  
  
  nand (_0451_, _0450_, _0450_);
  nand (_0452_, _0355_, _0358_);
  nand (_0453_, _0360_, _0452_);
  
  
  nand (_0454_, _0453_, _0453_);
  nand (_0455_, _0450_, _0454_);
  
  
  nand (_0456_, _0455_, _0455_);
  nand (_0457_, _0451_, _0453_);
  nand (_0458_, _0455_, _0457_);
  
  
  nand (_0459_, _0458_, _0458_);
  nand (_0461_, _0448_, _0459_);
  nand (_0462_, _0445_, _0461_);
  
  
  nand (_0463_, _0462_, _0462_);
  nand (_0464_, _0374_, _0377_);
  nand (_0465_, _0379_, _0464_);
  
  
  nand (_0466_, _0465_, _0465_);
  nand (_0467_, _0462_, _0466_);
  nand (_0468_, _0463_, _0465_);
  nand (_0469_, _0467_, _0468_);
  
  
  nand (_0470_, _0469_, _0469_);
  nand (_0472_, _0456_, _0470_);
  nand (_0473_, _0467_, _0472_);
  
  
  nand (_0474_, _0473_, _0473_);
  nand (_0475_, _0388_, _0390_);
  nand (_0476_, _0392_, _0475_);
  
  
  nand (_0477_, _0476_, _0476_);
  nand (_0478_, _0473_, _0477_);
  nand (_0479_, input_f[3], input_w[1]);
  
  
  nand (_0480_, _0479_, _0479_);
  nand (_0481_, input_f[3], input_w[0]);
  nand (_0483_, _0407_, _0480_);
  nand (_0484_, input_f[2], input_w[2]);
  
  
  nand (_0485_, _0484_, _0484_);
  nand (_0486_, _0406_, _0479_);
  nand (_0487_, _0483_, _0486_);
  
  
  nand (_0488_, _0487_, _0487_);
  nand (_0489_, _0485_, _0488_);
  nand (_0490_, _0483_, _0489_);
  
  
  nand (_0491_, _0490_, _0490_);
  nand (_0492_, _0409_, _0412_);
  nand (_0494_, _0414_, _0492_);
  
  
  nand (_0495_, _0494_, _0494_);
  nand (_0496_, _0490_, _0495_);
  nand (_0497_, input_f[0], input_w[5]);
  
  
  nand (_0498_, _0497_, _0497_);
  nand (_0499_, input_f[1], input_w[4]);
  
  
  nand (_0500_, _0499_, _0499_);
  nand (_0501_, input_f[1], input_w[3]);
  nand (_0502_, _0425_, _0500_);
  nand (_0503_, _0424_, _0499_);
  nand (_0505_, _0502_, _0503_);
  
  
  nand (_0506_, _0505_, _0505_);
  nand (_0507_, _0498_, _0506_);
  nand (_0508_, _0497_, _0505_);
  nand (_0509_, _0507_, _0508_);
  
  
  nand (_0510_, _0509_, _0509_);
  nand (_0511_, _0491_, _0494_);
  nand (_0512_, _0496_, _0511_);
  
  
  nand (_0513_, _0512_, _0512_);
  nand (_0514_, _0510_, _0513_);
  nand (_0516_, _0496_, _0514_);
  
  
  nand (_0517_, _0516_, _0516_);
  nand (_0518_, _0433_, _0436_);
  nand (_0519_, _0439_, _0518_);
  
  
  nand (_0520_, _0519_, _0519_);
  nand (_0521_, _0516_, _0520_);
  nand (_0522_, _0502_, _0507_);
  
  
  nand (_0523_, _0522_, _0522_);
  nand (_0524_, input_f[0], input_w[6]);
  
  
  nand (_0525_, _0524_, _0524_);
  nand (_0527_, _0522_, _0525_);
  
  
  nand (_0528_, _0527_, _0527_);
  nand (_0529_, _0523_, _0524_);
  nand (_0530_, _0527_, _0529_);
  
  
  nand (_0531_, _0530_, _0530_);
  nand (_0532_, _0517_, _0519_);
  nand (_0533_, _0521_, _0532_);
  
  
  nand (_0534_, _0533_, _0533_);
  nand (_0535_, _0531_, _0534_);
  nand (_0536_, _0521_, _0535_);
  
  
  nand (_0538_, _0536_, _0536_);
  nand (_0539_, _0447_, _0458_);
  nand (_0540_, _0461_, _0539_);
  
  
  nand (_0541_, _0540_, _0540_);
  nand (_0542_, _0536_, _0541_);
  nand (_0543_, _0538_, _0540_);
  nand (_0544_, _0542_, _0543_);
  
  
  nand (_0545_, _0544_, _0544_);
  nand (_0546_, _0528_, _0545_);
  nand (_0547_, _0542_, _0546_);
  
  
  nand (_0549_, _0547_, _0547_);
  nand (_0550_, _0455_, _0469_);
  nand (_0551_, _0472_, _0550_);
  
  
  nand (_0552_, _0551_, _0551_);
  nand (_0553_, _0547_, _0552_);
  nand (_0554_, input_f[2], input_w[1]);
  nand (_0555_, input_f[2], input_w[0]);
  
  
  nand (_0556_, _0555_, _0555_);
  nand (_0557_, _0480_, _0556_);
  nand (_0558_, input_f[1], input_w[2]);
  
  
  nand (_0560_, _0558_, _0558_);
  nand (_0561_, _0481_, _0554_);
  nand (_0562_, _0557_, _0561_);
  
  
  nand (_0563_, _0562_, _0562_);
  nand (_0564_, _0560_, _0563_);
  nand (_0565_, _0557_, _0564_);
  
  
  nand (_0566_, _0565_, _0565_);
  nand (_0567_, _0484_, _0487_);
  nand (_0568_, _0489_, _0567_);
  
  
  nand (_0569_, _0568_, _0568_);
  nand (_0571_, _0565_, _0569_);
  nand (_0572_, input_f[0], input_w[4]);
  nand (_0573_, input_f[0], input_w[3]);
  
  
  nand (_0574_, _0573_, _0573_);
  nand (_0575_, _0500_, _0574_);
  
  
  nand (_0576_, _0575_, _0575_);
  nand (_0577_, _0501_, _0572_);
  nand (_0578_, _0575_, _0577_);
  
  
  nand (_0579_, _0578_, _0578_);
  nand (_0580_, _0566_, _0568_);
  nand (_0582_, _0571_, _0580_);
  
  
  nand (_0583_, _0582_, _0582_);
  nand (_0584_, _0579_, _0583_);
  nand (_0585_, _0571_, _0584_);
  
  
  nand (_0586_, _0585_, _0585_);
  nand (_0587_, _0509_, _0512_);
  nand (_0588_, _0514_, _0587_);
  
  
  nand (_0589_, _0588_, _0588_);
  nand (_0590_, _0585_, _0589_);
  nand (_0591_, _0586_, _0588_);
  nand (_0593_, _0590_, _0591_);
  
  
  nand (_0594_, _0593_, _0593_);
  nand (_0595_, _0576_, _0594_);
  nand (_0596_, _0590_, _0595_);
  
  
  nand (_0597_, _0596_, _0596_);
  nand (_0598_, _0530_, _0533_);
  nand (_0599_, _0535_, _0598_);
  
  
  nand (_0600_, _0599_, _0599_);
  nand (_0601_, _0596_, _0600_);
  
  
  nand (_0602_, _0601_, _0601_);
  nand (_0604_, _0527_, _0544_);
  nand (_0605_, _0546_, _0604_);
  
  
  nand (_0606_, _0605_, _0605_);
  nand (_0607_, _0602_, _0606_);
  nand (_0608_, input_f[1], input_w[1]);
  
  
  nand (_0609_, _0608_, _0608_);
  nand (_0610_, input_f[1], input_w[0]);
  nand (_0611_, _0556_, _0609_);
  nand (_0612_, input_f[0], input_w[2]);
  
  
  nand (_0613_, _0612_, _0612_);
  nand (_0615_, _0555_, _0608_);
  nand (_0616_, _0611_, _0615_);
  
  
  nand (_0617_, _0616_, _0616_);
  nand (_0618_, _0613_, _0617_);
  nand (_0619_, _0611_, _0618_);
  
  
  nand (_0620_, _0619_, _0619_);
  nand (_0621_, _0558_, _0562_);
  nand (_0622_, _0564_, _0621_);
  
  
  nand (_0623_, _0622_, _0622_);
  nand (_0624_, _0619_, _0623_);
  nand (_0626_, _0620_, _0622_);
  nand (_0627_, _0624_, _0626_);
  
  
  nand (_0628_, _0627_, _0627_);
  nand (_0629_, _0574_, _0628_);
  nand (_0630_, _0624_, _0629_);
  
  
  nand (_0631_, _0630_, _0630_);
  nand (_0632_, _0578_, _0582_);
  nand (_0633_, _0584_, _0632_);
  
  
  nand (_0634_, _0633_, _0633_);
  nand (_0635_, _0630_, _0634_);
  
  
  nand (_0637_, _0635_, _0635_);
  nand (_0638_, _0575_, _0593_);
  nand (_0639_, _0595_, _0638_);
  
  
  nand (_0640_, _0639_, _0639_);
  nand (_0641_, _0637_, _0640_);
  
  
  nand (_0642_, _0641_, _0641_);
  nand (_0643_, _0597_, _0599_);
  nand (_0644_, _0601_, _0643_);
  
  
  nand (_0645_, _0644_, _0644_);
  nand (_0646_, _0642_, _0645_);
  nand (_0648_, input_f[0], input_w[1]);
  nand (_0649_, input_f[0], input_w[0]);
  
  
  nand (_0650_, _0649_, _0649_);
  nand (_0651_, _0609_, _0650_);
  
  
  nand (_0652_, _0651_, _0651_);
  nand (_0653_, _0612_, _0616_);
  nand (_0654_, _0618_, _0653_);
  
  
  nand (_0655_, _0654_, _0654_);
  nand (_0656_, _0652_, _0655_);
  
  
  nand (_0657_, _0656_, _0656_);
  nand (_0659_, _0573_, _0627_);
  nand (_0660_, _0629_, _0659_);
  
  
  nand (_0661_, _0660_, _0660_);
  nand (_0662_, _0657_, _0661_);
  
  
  nand (_0663_, _0662_, _0662_);
  nand (_0664_, _0631_, _0633_);
  nand (_0665_, _0635_, _0664_);
  
  
  nand (_0666_, _0665_, _0665_);
  nand (_0667_, _0663_, _0666_);
  
  
  nand (_0668_, _0667_, _0667_);
  nand (_0670_, _0635_, _0639_);
  nand (_0671_, _0641_, _0670_);
  
  
  nand (_0672_, _0671_, _0671_);
  nand (_0673_, _0668_, _0672_);
  
  
  nand (_0674_, _0673_, _0673_);
  nand (_0675_, _0641_, _0644_);
  nand (_0676_, _0646_, _0675_);
  
  
  nand (_0677_, _0676_, _0676_);
  nand (_0678_, _0674_, _0677_);
  nand (_0679_, _0646_, _0678_);
  
  
  nand (_0681_, _0679_, _0679_);
  nand (_0682_, _0601_, _0605_);
  nand (_0683_, _0607_, _0682_);
  
  
  nand (_0684_, _0683_, _0683_);
  nand (_0685_, _0679_, _0684_);
  nand (_0686_, _0607_, _0685_);
  
  
  nand (_0687_, _0686_, _0686_);
  nand (_0688_, _0549_, _0551_);
  nand (_0689_, _0553_, _0688_);
  
  
  nand (_0690_, _0689_, _0689_);
  nand (_0692_, _0686_, _0690_);
  nand (_0693_, _0553_, _0692_);
  
  
  nand (_0694_, _0693_, _0693_);
  nand (_0695_, _0474_, _0476_);
  nand (_0696_, _0478_, _0695_);
  
  
  nand (_0697_, _0696_, _0696_);
  nand (_0698_, _0693_, _0697_);
  nand (_0699_, _0478_, _0698_);
  
  
  nand (_0700_, _0699_, _0699_);
  nand (_0701_, _0402_, _0699_);
  nand (_0703_, _0399_, _0701_);
  
  
  nand (_0704_, _0703_, _0703_);
  nand (_0705_, _0311_, _0703_);
  nand (_0706_, _0308_, _0705_);
  
  
  nand (_0707_, _0706_, _0706_);
  nand (_0708_, _0227_, _0229_);
  nand (_0709_, _0231_, _0708_);
  
  
  nand (_0710_, _0709_, _0709_);
  nand (_0711_, _0706_, _0710_);
  nand (_0712_, _0231_, _0711_);
  
  
  nand (_0714_, _0712_, _0712_);
  nand (_0715_, _0123_, _0160_);
  nand (_0716_, _0162_, _0715_);
  
  
  nand (_0717_, _0716_, _0716_);
  nand (_0718_, _0712_, _0717_);
  nand (_0719_, _0162_, _0718_);
  
  
  nand (_0720_, _0719_, _0719_);
  nand (_0721_, _0154_, _0158_);
  
  
  nand (_0722_, _0721_, _0721_);
  nand (_0723_, _0142_, _0146_);
  
  
  nand (_0725_, _0723_, _0723_);
  nand (_0726_, _0460_, input_w[7]);
  nand (_0727_, _0134_, _0726_);
  nand (_0728_, _0138_, _0727_);
  
  
  nand (_0729_, _0728_, _0728_);
  nand (_0730_, _0133_, _0728_);
  
  
  nand (_0731_, _0730_, _0730_);
  nand (_0732_, _0132_, _0729_);
  nand (_0733_, _0730_, _0732_);
  
  
  nand (_0734_, _0733_, _0733_);
  nand (_0736_, _0131_, _0733_);
  nand (_0737_, _0130_, _0734_);
  nand (_0738_, _0736_, _0737_);
  
  
  nand (_0739_, _0738_, _0738_);
  nand (_0740_, _0128_, _0150_);
  
  
  nand (_0741_, _0740_, _0740_);
  nand (_0742_, _0738_, _0740_);
  nand (_0743_, _0739_, _0741_);
  nand (_0744_, _0742_, _0743_);
  
  
  nand (_0745_, _0744_, _0744_);
  nand (_0747_, _0723_, _0745_);
  nand (_0748_, _0725_, _0744_);
  nand (_0749_, _0747_, _0748_);
  
  
  nand (_0750_, _0749_, _0749_);
  nand (_0751_, _0721_, _0750_);
  nand (_0752_, _0722_, _0749_);
  nand (_0753_, _0751_, _0752_);
  
  
  nand (_0754_, _0753_, _0753_);
  nand (_0755_, _0719_, _0754_);
  nand (_0756_, _0742_, _0747_);
  
  
  nand (_0758_, _0756_, _0756_);
  nand (_0759_, _0128_, _0736_);
  
  
  nand (_0760_, _0759_, _0759_);
  nand (_0761_, _0731_, _0759_);
  nand (_0762_, _0730_, _0760_);
  nand (_0763_, _0761_, _0762_);
  nand (_0764_, _0758_, _0763_);
  nand (_0765_, _0730_, _0759_);
  nand (_0766_, _0764_, _0765_);
  nand (_0767_, _0751_, _0766_);
  
  
  nand (_0769_, _0767_, _0767_);
  nand (_0770_, _0755_, _0769_);
  
  
  nand (_0771_, _0770_, _0770_);
  nand (_0772_, _0720_, _0753_);
  nand (_0773_, _0755_, _0772_);
  nand (_0774_, _0714_, _0716_);
  nand (_0775_, _0718_, _0774_);
  
  
  nand (_0776_, _0775_, _0775_);
  nand (_0777_, _0707_, _0709_);
  nand (_0778_, _0711_, _0777_);
  
  
  nand (_0780_, _0778_, _0778_);
  nand (_0781_, _0310_, _0704_);
  nand (_0782_, _0705_, _0781_);
  
  
  nand (_0783_, _0782_, _0782_);
  nand (_0784_, _0401_, _0700_);
  nand (_0785_, _0701_, _0784_);
  
  
  nand (_0786_, _0785_, _0785_);
  nand (_0787_, _0681_, _0683_);
  nand (_0788_, _0685_, _0787_);
  
  
  nand (_0789_, _0788_, _0788_);
  nand (_0791_, _0687_, _0689_);
  nand (_0792_, _0692_, _0791_);
  
  
  nand (_0793_, _0792_, _0792_);
  nand (_0794_, _0788_, _0792_);
  
  
  nand (_0795_, _0794_, _0794_);
  nand (_0796_, _0694_, _0696_);
  nand (_0797_, _0698_, _0796_);
  
  
  nand (_0798_, _0797_, _0797_);
  nand (_0799_, _0795_, _0797_);
  
  
  nand (_0800_, _0799_, _0799_);
  nand (_0802_, _0785_, _0800_);
  
  
  nand (_0803_, _0802_, _0802_);
  nand (_0804_, _0782_, _0803_);
  
  
  nand (_0805_, _0804_, _0804_);
  nand (_0806_, _0778_, _0805_);
  
  
  nand (_0807_, _0806_, _0806_);
  nand (_0808_, _0775_, _0807_);
  
  
  nand (_0809_, _0808_, _0808_);
  nand (_0810_, _0773_, _0809_);
  nand (_0811_, _0770_, _0810_);
  nand (_0813_, _0789_, _0793_);
  
  
  nand (_0814_, _0813_, _0813_);
  nand (_0815_, _0798_, _0814_);
  
  
  nand (_0816_, _0815_, _0815_);
  nand (_0817_, _0786_, _0816_);
  
  
  nand (_0818_, _0817_, _0817_);
  nand (_0819_, _0783_, _0818_);
  
  
  nand (_0820_, _0819_, _0819_);
  nand (_0821_, _0780_, _0820_);
  
  
  nand (_0822_, _0821_, _0821_);
  nand (_0824_, _0776_, _0822_);
  nand (_0825_, _0771_, _0824_);
  nand (_0826_, _0673_, _0676_);
  nand (_0827_, _0678_, _0826_);
  
  
  nand (_0828_, _0827_, _0827_);
  nand (_0829_, _0825_, _0828_);
  nand (_0830_, _0811_, _0829_);
  
  
  nand (_0831_, _0830_, _0830_);
  nand (_0832_, _0482_, psum_reg[6]);
  
  
  nand (_0833_, _0832_, _0832_);
  nand (_0835_, _0830_, _0833_);
  nand (_0836_, _0667_, _0671_);
  nand (_0837_, _0673_, _0836_);
  
  
  nand (_0838_, _0837_, _0837_);
  nand (_0839_, _0825_, _0838_);
  nand (_0840_, _0811_, _0839_);
  
  
  nand (_0841_, _0840_, _0840_);
  nand (_0842_, _0482_, psum_reg[5]);
  
  
  nand (_0843_, _0842_, _0842_);
  nand (_0844_, _0840_, _0843_);
  nand (_0846_, _0662_, _0665_);
  nand (_0847_, _0667_, _0846_);
  
  
  nand (_0848_, _0847_, _0847_);
  nand (_0849_, _0825_, _0848_);
  nand (_0850_, _0811_, _0849_);
  
  
  nand (_0851_, _0850_, _0850_);
  nand (_0852_, _0482_, psum_reg[4]);
  
  
  nand (_0853_, _0852_, _0852_);
  nand (_0854_, _0850_, _0853_);
  nand (_0855_, _0851_, _0852_);
  nand (_0857_, _0854_, _0855_);
  
  
  nand (_0858_, _0857_, _0857_);
  nand (_0859_, _0656_, _0660_);
  nand (_0860_, _0662_, _0859_);
  
  
  nand (_0861_, _0860_, _0860_);
  nand (_0862_, _0825_, _0861_);
  nand (_0863_, _0811_, _0862_);
  
  
  nand (_0864_, _0863_, _0863_);
  nand (_0865_, _0482_, psum_reg[3]);
  
  
  nand (_0866_, _0865_, _0865_);
  nand (_0868_, _0863_, _0866_);
  nand (_0869_, _0864_, _0865_);
  nand (_0870_, _0651_, _0654_);
  nand (_0871_, _0656_, _0870_);
  
  
  nand (_0872_, _0871_, _0871_);
  nand (_0873_, _0825_, _0872_);
  nand (_0874_, _0811_, _0873_);
  
  
  nand (_0875_, _0874_, _0874_);
  nand (_0876_, _0482_, psum_reg[2]);
  
  
  nand (_0877_, _0876_, _0876_);
  nand (_0879_, _0874_, _0877_);
  nand (_0880_, _0875_, _0876_);
  nand (_0881_, _0482_, psum_reg[1]);
  
  
  nand (_0882_, _0881_, _0881_);
  nand (_0883_, _0610_, _0648_);
  nand (_0884_, _0651_, _0883_);
  
  
  nand (_0885_, _0884_, _0884_);
  nand (_0886_, _0811_, _0884_);
  nand (_0887_, _0825_, _0885_);
  nand (_0888_, _0811_, _0887_);
  nand (_0890_, _0825_, _0886_);
  nand (_0891_, _0882_, _0888_);
  nand (_0892_, _0881_, _0890_);
  nand (_0893_, psum_reg[0], _0482_);
  
  
  nand (_0894_, _0893_, _0893_);
  nand (_0895_, _0649_, _0811_);
  nand (_0896_, _0650_, _0825_);
  nand (_0897_, _0811_, _0896_);
  nand (_0898_, _0825_, _0895_);
  nand (_0899_, _0894_, _0897_);
  
  
  nand (_0901_, _0899_, _0899_);
  nand (_0902_, _0892_, _0901_);
  nand (_0903_, _0891_, _0899_);
  nand (_0904_, _0892_, _0903_);
  nand (_0905_, _0891_, _0902_);
  nand (_0906_, _0880_, _0905_);
  nand (_0907_, _0879_, _0904_);
  nand (_0908_, _0880_, _0907_);
  nand (_0909_, _0879_, _0906_);
  nand (_0910_, _0869_, _0909_);
  nand (_0912_, _0868_, _0908_);
  nand (_0913_, _0869_, _0912_);
  nand (_0914_, _0868_, _0910_);
  nand (_0915_, _0858_, _0914_);
  nand (_0916_, _0854_, _0915_);
  
  
  nand (_0917_, _0916_, _0916_);
  nand (_0918_, _0841_, _0842_);
  nand (_0919_, _0844_, _0918_);
  
  
  nand (_0920_, _0919_, _0919_);
  nand (_0921_, _0916_, _0920_);
  nand (_0923_, _0844_, _0921_);
  
  
  nand (_0924_, _0923_, _0923_);
  nand (_0925_, _0831_, _0832_);
  nand (_0926_, _0835_, _0925_);
  
  
  nand (_0927_, _0926_, _0926_);
  nand (_0928_, _0923_, _0927_);
  nand (_0929_, _0835_, _0928_);
  
  
  nand (_0930_, _0929_, _0929_);
  nand (_0931_, _0504_, _0770_);
  
  
  nand (_0932_, _0931_, _0931_);
  nand (_0934_, _0929_, _0932_);
  nand (_0935_, enable, _0934_);
  
  
  nand (_0936_, _0935_, _0935_);
  nand (_0937_, _0515_, _0771_);
  nand (_0938_, _0931_, _0937_);
  
  
  nand (_0939_, _0938_, _0938_);
  nand (_0940_, _0929_, _0938_);
  nand (_0941_, _0930_, _0939_);
  nand (_0942_, _0930_, _0938_);
  nand (_0943_, _0929_, _0939_);
  nand (_0945_, _0942_, _0943_);
  nand (_0946_, _0940_, _0941_);
  nand (_0947_, _0937_, _0945_);
  nand (_0948_, _0936_, _0947_);
  nand (psum_next[7], _0526_, _0948_);
  
  
  nand (_0949_, psum_next[7], psum_next[7]);
  nand (_0950_, _0493_, _0842_);
  nand (_0951_, _0931_, _0946_);
  nand (_0952_, _0947_, _0951_);
  nand (_0953_, _0917_, _0919_);
  nand (_0955_, _0921_, _0953_);
  
  
  nand (_0956_, _0955_, _0955_);
  nand (_0957_, _0952_, _0956_);
  nand (_0958_, _0936_, _0957_);
  nand (_0959_, _0950_, _0958_);
  
  
  nand (psum_next[5], _0959_, _0959_);
  nand (_0960_, _0868_, _0869_);
  
  
  nand (_0961_, _0960_, _0960_);
  nand (_0962_, _0908_, _0961_);
  nand (_0963_, _0909_, _0960_);
  nand (_0965_, _0962_, _0963_);
  nand (_0966_, _0952_, _0965_);
  nand (_0967_, _0936_, _0966_);
  nand (_0968_, _0493_, _0865_);
  nand (_0969_, _0967_, _0968_);
  
  
  nand (psum_next[3], _0969_, _0969_);
  nand (_0970_, _0493_, _0832_);
  nand (_0971_, _0924_, _0926_);
  nand (_0972_, _0928_, _0971_);
  
  
  nand (_0973_, _0972_, _0972_);
  nand (_0975_, _0952_, _0973_);
  nand (_0976_, _0936_, _0975_);
  nand (_0977_, _0970_, _0976_);
  
  
  nand (psum_next[6], _0977_, _0977_);
  nand (_0978_, _0857_, _0913_);
  nand (_0979_, _0915_, _0978_);
  
  
  nand (_0980_, _0979_, _0979_);
  nand (_0981_, _0952_, _0980_);
  nand (_0982_, _0936_, _0981_);
  nand (_0983_, _0493_, _0852_);
  nand (_0000_, _0982_, _0983_);
  
  
  nand (psum_next[4], _0000_, _0000_);
  nand (_0001_, _0879_, _0880_);
  
  
  nand (_0002_, _0001_, _0001_);
  nand (_0003_, _0904_, _0002_);
  nand (_0004_, _0905_, _0001_);
  nand (_0005_, _0003_, _0004_);
  nand (_0006_, _0952_, _0005_);
  nand (_0007_, _0936_, _0006_);
  nand (_0008_, _0493_, _0876_);
  nand (_0010_, _0007_, _0008_);
  
  
  nand (psum_next[2], _0010_, _0010_);
  nand (_0011_, _0949_, psum_next[6]);
  
  
  nand (output_f[6], _0011_, _0011_);
  nand (_0012_, _0949_, psum_next[5]);
  
  
  nand (output_f[5], _0012_, _0012_);
  nand (_0013_, _0949_, psum_next[4]);
  
  
  nand (output_f[4], _0013_, _0013_);
  nand (_0014_, _0949_, psum_next[3]);
  
  
  nand (output_f[3], _0014_, _0014_);
  nand (_0016_, _0949_, psum_next[2]);
  
  
  nand (output_f[2], _0016_, _0016_);
  nand (_0017_, _0891_, _0892_);
  
  
  nand (_0018_, _0017_, _0017_);
  nand (_0019_, _0899_, _0018_);
  nand (_0020_, _0901_, _0017_);
  nand (_0021_, _0019_, _0020_);
  nand (_0022_, _0952_, _0021_);
  nand (_0023_, _0936_, _0022_);
  nand (_0024_, _0493_, _0881_);
  nand (_0026_, _0023_, _0024_);
  
  
  nand (psum_next[1], _0026_, _0026_);
  nand (_0027_, _0949_, psum_next[1]);
  
  
  nand (output_f[1], _0027_, _0027_);
  nand (_0028_, _0893_, _0898_);
  nand (_0029_, _0899_, _0028_);
  
  
  nand (_0030_, _0029_, _0029_);
  nand (_0031_, _0952_, _0030_);
  nand (_0032_, _0936_, _0031_);
  nand (_0033_, _0493_, _0893_);
  nand (_0035_, _0032_, _0033_);
  
  
  nand (psum_next[0], _0035_, _0035_);
  nand (_0036_, _0949_, psum_next[0]);
  
  
  nand (output_f[0], _0036_, _0036_);
  assign mac1.output_f[0] = mac1.adder1.SUM[0];
  assign mac1.output_f[1] = mac1.adder1.SUM[1];
  assign mac1.output_f[2] = mac1.adder1.SUM[2];
  assign mac1.output_f[3] = mac1.adder1.SUM[3];
  assign mac1.output_f[4] = mac1.adder1.SUM[4];
  assign mac1.output_f[5] = mac1.adder1.SUM[5];
  assign mac1.output_f[6] = mac1.adder1.SUM[6];
  assign mac1.output_f[7] = mac1.adder1.SUM[7];
  assign mac1.mult_out[0] = mac1.adder1.A[0];
  assign mac1.mult_out[1] = mac1.adder1.A[1];
  assign mac1.mult_out[2] = mac1.adder1.A[2];
  assign mac1.mult_out[3] = mac1.adder1.A[3];
  assign mac1.mult_out[4] = mac1.adder1.A[4];
  assign mac1.mult_out[5] = mac1.adder1.A[5];
  assign mac1.mult_out[6] = mac1.adder1.A[6];
  assign mac1.mult_out[7] = mac1.adder1.A[7];
  assign mac1.input_w[0] = input_w[0];
  assign mac1.input_w[1] = input_w[1];
  assign mac1.input_w[2] = input_w[2];
  assign mac1.input_w[3] = input_w[3];
  assign mac1.input_w[4] = input_w[4];
  assign mac1.input_w[5] = input_w[5];
  assign mac1.input_w[6] = input_w[6];
  assign mac1.input_w[7] = input_w[7];
  assign mac1.input_psum[0] = mac1.adder1.B[0];
  assign mac1.input_psum[1] = mac1.adder1.B[1];
  assign mac1.input_psum[2] = mac1.adder1.B[2];
  assign mac1.input_psum[3] = mac1.adder1.B[3];
  assign mac1.input_psum[4] = mac1.adder1.B[4];
  assign mac1.input_psum[5] = mac1.adder1.B[5];
  assign mac1.input_psum[6] = mac1.adder1.B[6];
  assign mac1.input_psum[7] = mac1.adder1.B[7];
  assign mac1.input_f[0] = input_f[0];
  assign mac1.input_f[1] = input_f[1];
  assign mac1.input_f[2] = input_f[2];
  assign mac1.input_f[3] = input_f[3];
  assign mac1.input_f[4] = input_f[4];
  assign mac1.input_f[5] = input_f[5];
  assign mac1.input_f[6] = input_f[6];
  assign mac1.input_f[7] = input_f[7];
  assign mac1.adder_out[0] = mac1.adder1.SUM[0];
  assign mac1.adder_out[1] = mac1.adder1.SUM[1];
  assign mac1.adder_out[2] = mac1.adder1.SUM[2];
  assign mac1.adder_out[3] = mac1.adder1.SUM[3];
  assign mac1.adder_out[4] = mac1.adder1.SUM[4];
  assign mac1.adder_out[5] = mac1.adder1.SUM[5];
  assign mac1.adder_out[6] = mac1.adder1.SUM[6];
  assign mac1.adder_out[7] = mac1.adder1.SUM[7];
  assign mac1.mult1.a[0] = input_f[0];
  assign mac1.mult1.a[1] = input_f[1];
  assign mac1.mult1.a[2] = input_f[2];
  assign mac1.mult1.a[3] = input_f[3];
  assign mac1.mult1.a[4] = input_f[4];
  assign mac1.mult1.a[5] = input_f[5];
  assign mac1.mult1.a[6] = input_f[6];
  assign mac1.mult1.a[7] = input_f[7];
  assign mac1.mult1.b[0]  = input_w[0];
  assign mac1.mult1.b[1]  = input_w[1];
  assign mac1.mult1.b[2]  = input_w[2];
  assign mac1.mult1.b[3]  = input_w[3];
  assign mac1.mult1.b[4]  = input_w[4];
  assign mac1.mult1.b[5]  = input_w[5];
  assign mac1.mult1.b[6]  = input_w[6];
  assign mac1.mult1.b[7]  = input_w[7];
  assign mac1.mult1.product[0] = mac1.adder1.A[0];
  assign mac1.mult1.product[1] = mac1.adder1.A[1];
  assign mac1.mult1.product[2] = mac1.adder1.A[2];
  assign mac1.mult1.product[3] = mac1.adder1.A[3];
  assign mac1.mult1.product[4] = mac1.adder1.A[4];
  assign mac1.mult1.product[5] = mac1.adder1.A[5];
  assign mac1.mult1.product[6] = mac1.adder1.A[6];
  assign mac1.mult1.product[7] = mac1.adder1.A[7];
  assign mac1.adder1.cla1.COUT  = mac1.adder1.C[0];
  assign mac1.adder1.cla1.CIN  = 1'h0;
  assign mac1.adder1.cla1.B[0] = mac1.adder1.B[0];
  assign mac1.adder1.cla1.B[1] = mac1.adder1.B[1];
  assign mac1.adder1.cla1.B[2] = mac1.adder1.B[2];
  assign mac1.adder1.cla1.B[3] = mac1.adder1.B[3];
  assign mac1.adder1.cla1.A[0] = mac1.adder1.A[0];
  assign mac1.adder1.cla1.A[1] = mac1.adder1.A[1];
  assign mac1.adder1.cla1.A[2] = mac1.adder1.A[2];
  assign mac1.adder1.cla1.A[3] = mac1.adder1.A[3];
  assign mac1.adder1.cla1.fa3.a  = mac1.adder1.A[3];
  assign mac1.adder1.cla1.fa3.b  = mac1.adder1.B[3];
  assign mac1.adder1.cla1.fa2.a  = mac1.adder1.A[2];
  assign mac1.adder1.cla1.fa2.b  = mac1.adder1.B[2];
  assign mac1.adder1.cla1.fa1.a  = mac1.adder1.A[1];
  assign mac1.adder1.cla1.fa1.b  = mac1.adder1.B[1];
  assign mac1.adder1.cla1.fa0.a  = mac1.adder1.A[0];
  assign mac1.adder1.cla1.fa0.b  = mac1.adder1.B[0];
  assign mac1.adder1.cla1.fa0.cin  = 1'h0;
  assign mac1.adder1.cla2.COUT  = mac1.adder1.C[1];
  assign mac1.adder1.cla2.CIN  = mac1.adder1.C[0];
  assign mac1.adder1.cla2.B[0] = mac1.adder1.B[4];
  assign mac1.adder1.cla2.B[1] = mac1.adder1.B[5];
  assign mac1.adder1.cla2.B[2] = mac1.adder1.B[6];
  assign mac1.adder1.cla2.B[3] = mac1.adder1.B[7];
  assign mac1.adder1.cla2.A[0] = mac1.adder1.A[4];
  assign mac1.adder1.cla2.A[1] = mac1.adder1.A[5];
  assign mac1.adder1.cla2.A[2] = mac1.adder1.A[6];
  assign mac1.adder1.cla2.A[3] = mac1.adder1.A[7];
  assign mac1.adder1.cla2.fa3.a  = mac1.adder1.A[7];
  assign mac1.adder1.cla2.fa3.b  = mac1.adder1.B[7];
  assign mac1.adder1.cla2.fa2.a  = mac1.adder1.A[6];
  assign mac1.adder1.cla2.fa2.b  = mac1.adder1.B[6];
  assign mac1.adder1.cla2.fa1.a  = mac1.adder1.A[5];
  assign mac1.adder1.cla2.fa1.b  = mac1.adder1.B[5];
  assign mac1.adder1.cla2.fa0.a  = mac1.adder1.A[4];
  assign mac1.adder1.cla2.fa0.b  = mac1.adder1.B[4];
  assign mac1.adder1.cla2.fa0.cin  = mac1.adder1.C[0];
  assign mac1.adder1.sat_sum[7] = mac1.adder1.A[7];
  assign mac1.adder1.sat_sum[5] = mac1.adder1.sat_sum[6];
  assign mac1.adder1.sat_sum[4] = mac1.adder1.sat_sum[6];
  assign mac1.adder1.sat_sum[3] = mac1.adder1.sat_sum[6];
  assign mac1.adder1.sat_sum[2] = mac1.adder1.sat_sum[6];
  assign mac1.adder1.sat_sum[1] = mac1.adder1.sat_sum[6];
  assign mac1.adder1.sat_sum[0] = mac1.adder1.sat_sum[6];
  assign relu1.output_f[7]  = 1'h0;
  assign relu1.output_f[6] = output_f[6];
  assign relu1.output_f[5] = output_f[5];
  assign relu1.output_f[4] = output_f[4];
  assign relu1.output_f[3] = output_f[3];
  assign relu1.output_f[2] = output_f[2];
  assign relu1.output_f[1] = output_f[1];
  assign relu1.output_f[0] = output_f[0];
  assign relu1.input_f[0] = psum_next[0];
  assign relu1.input_f[1] = psum_next[1];
  assign relu1.input_f[2] = psum_next[2];
  assign relu1.input_f[3] = psum_next[3];
  assign relu1.input_f[4] = psum_next[4];
  assign relu1.input_f[5] = psum_next[5];
  assign relu1.input_f[6] = psum_next[6];
  assign relu1.input_f[7] = psum_next[7];
  assign input_psum[0] = mac1.adder1.B[0];
  assign input_psum[1] = mac1.adder1.B[1];
  assign input_psum[2] = mac1.adder1.B[2];
  assign input_psum[3] = mac1.adder1.B[3];
  assign input_psum[4] = mac1.adder1.B[4];
  assign input_psum[5] = mac1.adder1.B[5];
  assign input_psum[6] = mac1.adder1.B[6];
  assign input_psum[7] = mac1.adder1.B[7];
  assign mac_out[0] = mac1.adder1.SUM[0];
  assign mac_out[1] = mac1.adder1.SUM[1];
  assign mac_out[2] = mac1.adder1.SUM[2];
  assign mac_out[3] = mac1.adder1.SUM[3];
  assign mac_out[4] = mac1.adder1.SUM[4];
  assign mac_out[5] = mac1.adder1.SUM[5];
  assign mac_out[6] = mac1.adder1.SUM[6];
  assign mac_out[7] = mac1.adder1.SUM[7];
  assign output_f[7] = 1'h0;
endmodule
