module c6288(G1,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,
  G24,G25,G26,G27,G28,G29,G3,G30,G31,G32,G4,G5,G6,G6257,G6258,G6259,G6260,
  G6261,G6262,G6263,G6264,G6265,G6266,G6267,G6268,G6269,G6270,G6271,G6272,
  G6273,G6274,G6275,G6276,G6277,G6278,G6279,G6280,G6281,G6282,G6283,G6284,
  G6285,G6286,G6287,G6288,G7,G8,G9);
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
  G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32;
output G6257,G6258,G6259,G6260,G6261,G6262,G6263,G6264,G6265,G6266,G6267,G6268,
  G6269,G6270,G6271,G6272,G6273,G6274,G6275,G6276,G6277,G6278,G6279,G6280,
  G6281,G6282,G6283,G6284,G6285,G6286,G6287,G6288;

  wire G545,G548,G551,G554,G557,G560,G563,G566,G569,G572,G575,G578,G581,G584,
    G587,G590,G593,G596,G599,G602,G605,G608,G611,G614,G617,G620,G623,G626,G629,
    G632,G635,G638,G641,G644,G647,G650,G653,G656,G659,G662,G665,G668,G671,G674,
    G677,G680,G683,G686,G689,G692,G695,G698,G701,G704,G707,G710,G713,G716,G719,
    G722,G725,G728,G731,G734,G737,G740,G743,G746,G749,G752,G755,G758,G761,G764,
    G767,G770,G773,G776,G779,G782,G785,G788,G791,G794,G797,G800,G803,G806,G809,
    G812,G815,G818,G821,G824,G827,G830,G833,G836,G839,G842,G845,G848,G851,G854,
    G857,G860,G863,G866,G869,G872,G875,G878,G881,G884,G887,G890,G893,G896,G899,
    G902,G905,G908,G911,G914,G917,G920,G923,G926,G929,G932,G935,G938,G941,G944,
    G947,G950,G953,G956,G959,G962,G965,G968,G971,G974,G977,G980,G983,G986,G989,
    G992,G995,G998,G1001,G1004,G1007,G1010,G1013,G1016,G1019,G1022,G1025,G1028,
    G1031,G1034,G1037,G1040,G1043,G1046,G1049,G1052,G1055,G1058,G1061,G1064,
    G1067,G1070,G1073,G1076,G1079,G1082,G1085,G1088,G1091,G1094,G1097,G1100,
    G1103,G1106,G1109,G1112,G1115,G1118,G1121,G1124,G1127,G1130,G1133,G1136,
    G1139,G1142,G1145,G1148,G1151,G1154,G1157,G1160,G1163,G1166,G1169,G1172,
    G1175,G1178,G1181,G1184,G1187,G1190,G1193,G1196,G1199,G1202,G1205,G1208,
    G1211,G1214,G1217,G1220,G1223,G1226,G1229,G1232,G1235,G1238,G1241,G1244,
    G1247,G1250,G1253,G1256,G1259,G1262,G1265,G1268,G1271,G1274,G1277,G1280,
    G1283,G1286,G1289,G1292,G1295,G1298,G1301,G1304,G1307,G1310,G1314,G1318,
    G1322,G1326,G1330,G1334,G1338,G1342,G1346,G1350,G1354,G1358,G1362,G1366,
    G1370,G1371,G1372,G1373,G1374,G1375,G1376,G1377,G1378,G1379,G1380,G1381,
    G1382,G1383,G1384,G1385,G1386,G1387,G1388,G1389,G1390,G1391,G1392,G1393,
    G1394,G1395,G1396,G1397,G1398,G1399,G1400,G1403,G1406,G1409,G1412,G1415,
    G1418,G1421,G1424,G1427,G1430,G1433,G1436,G1439,G1442,G1445,G1449,G1453,
    G1457,G1461,G1465,G1469,G1473,G1477,G1481,G1485,G1489,G1493,G1497,G1501,
    G1505,G1506,G1507,G1510,G1511,G1512,G1515,G1516,G1517,G1520,G1521,G1522,
    G1525,G1526,G1527,G1530,G1531,G1532,G1535,G1536,G1537,G1540,G1541,G1542,
    G1545,G1546,G1547,G1550,G1551,G1552,G1555,G1556,G1557,G1560,G1561,G1562,
    G1565,G1566,G1567,G1570,G1571,G1572,G1575,G1576,G1577,G1580,G1583,G1586,
    G1589,G1592,G1595,G1598,G1601,G1604,G1607,G1610,G1613,G1616,G1619,G1622,
    G1626,G1630,G1634,G1638,G1642,G1646,G1650,G1654,G1658,G1662,G1666,G1670,
    G1674,G1678,G1682,G1683,G1684,G1685,G1686,G1687,G1688,G1689,G1690,G1691,
    G1692,G1693,G1694,G1695,G1696,G1697,G1698,G1699,G1700,G1701,G1702,G1703,
    G1704,G1705,G1706,G1707,G1708,G1709,G1710,G1711,G1712,G1715,G1718,G1721,
    G1724,G1727,G1730,G1733,G1736,G1739,G1742,G1745,G1748,G1751,G1754,G1757,
    G1761,G1765,G1769,G1773,G1777,G1781,G1785,G1789,G1793,G1797,G1801,G1805,
    G1809,G1813,G1817,G1818,G1819,G1822,G1823,G1824,G1827,G1828,G1829,G1832,
    G1833,G1834,G1837,G1838,G1839,G1842,G1843,G1844,G1847,G1848,G1849,G1852,
    G1853,G1854,G1857,G1858,G1859,G1862,G1863,G1864,G1867,G1868,G1869,G1872,
    G1873,G1874,G1877,G1878,G1879,G1882,G1883,G1884,G1887,G1888,G1889,G1892,
    G1895,G1899,G1902,G1905,G1908,G1911,G1914,G1917,G1920,G1923,G1926,G1929,
    G1932,G1935,G1938,G1942,G1943,G1944,G1948,G1952,G1956,G1960,G1964,G1968,
    G1972,G1976,G1980,G1984,G1988,G1992,G1996,G1997,G1998,G2001,G2002,G2003,
    G2004,G2005,G2006,G2007,G2008,G2009,G2010,G2011,G2012,G2013,G2014,G2015,
    G2016,G2017,G2018,G2019,G2020,G2021,G2022,G2023,G2024,G2025,G2026,G2027,
    G2030,G2034,G2037,G2040,G2043,G2046,G2049,G2052,G2055,G2058,G2061,G2064,
    G2067,G2070,G2073,G2077,G2078,G2079,G2082,G2086,G2090,G2094,G2098,G2102,
    G2106,G2110,G2114,G2118,G2122,G2126,G2130,G2134,G2135,G2136,G2139,G2142,
    G2146,G2147,G2148,G2151,G2152,G2153,G2156,G2157,G2158,G2161,G2162,G2163,
    G2166,G2167,G2168,G2171,G2172,G2173,G2176,G2177,G2178,G2181,G2182,G2183,
    G2186,G2187,G2188,G2191,G2192,G2193,G2196,G2197,G2198,G2201,G2202,G2203,
    G2206,G2207,G2208,G2211,G2214,G2218,G2219,G2220,G2223,G2226,G2229,G2232,
    G2235,G2238,G2241,G2244,G2247,G2250,G2253,G2256,G2260,G2261,G2262,G2265,
    G2269,G2273,G2277,G2281,G2285,G2289,G2293,G2297,G2301,G2305,G2309,G2313,
    G2314,G2315,G2318,G2322,G2323,G2324,G2325,G2326,G2327,G2328,G2329,G2330,
    G2331,G2332,G2333,G2334,G2335,G2336,G2337,G2338,G2339,G2340,G2341,G2342,
    G2343,G2344,G2345,G2346,G2349,G2353,G2354,G2355,G2358,G2361,G2364,G2367,
    G2370,G2373,G2376,G2379,G2382,G2385,G2388,G2391,G2394,G2398,G2399,G2400,
    G2403,G2406,G2410,G2414,G2418,G2422,G2426,G2430,G2434,G2438,G2442,G2446,
    G2450,G2454,G2458,G2459,G2460,G2463,G2466,G2470,G2471,G2472,G2473,G2474,
    G2477,G2478,G2479,G2482,G2483,G2484,G2487,G2488,G2489,G2492,G2493,G2494,
    G2497,G2498,G2499,G2502,G2503,G2504,G2507,G2508,G2509,G2512,G2513,G2514,
    G2517,G2518,G2519,G2522,G2523,G2524,G2527,G2528,G2529,G2532,G2535,G2539,
    G2540,G2541,G2544,G2547,G2550,G2553,G2556,G2559,G2562,G2565,G2568,G2571,
    G2574,G2577,G2581,G2582,G2583,G2586,G2590,G2594,G2598,G2602,G2606,G2610,
    G2614,G2618,G2622,G2626,G2630,G2634,G2635,G2636,G2639,G2643,G2644,G2645,
    G2648,G2649,G2650,G2651,G2652,G2653,G2654,G2655,G2656,G2657,G2658,G2659,
    G2660,G2661,G2662,G2663,G2664,G2665,G2666,G2667,G2668,G2669,G2670,G2673,
    G2677,G2678,G2679,G2682,G2685,G2689,G2692,G2695,G2698,G2701,G2704,G2707,
    G2710,G2713,G2716,G2719,G2722,G2726,G2727,G2728,G2731,G2734,G2738,G2739,
    G2740,G2744,G2748,G2752,G2756,G2760,G2764,G2768,G2772,G2776,G2780,G2784,
    G2785,G2786,G2789,G2792,G2796,G2797,G2798,G2801,G2802,G2803,G2806,G2807,
    G2808,G2811,G2812,G2813,G2816,G2817,G2818,G2821,G2822,G2823,G2826,G2827,
    G2828,G2831,G2832,G2833,G2836,G2837,G2838,G2841,G2842,G2843,G2846,G2847,
    G2848,G2851,G2852,G2853,G2856,G2859,G2863,G2864,G2865,G2868,G2872,G2875,
    G2878,G2881,G2884,G2887,G2890,G2893,G2896,G2899,G2902,G2906,G2907,G2908,
    G2911,G2915,G2916,G2917,G2920,G2924,G2928,G2932,G2936,G2940,G2944,G2948,
    G2952,G2956,G2960,G2961,G2962,G2965,G2969,G2970,G2971,G2974,G2977,G2981,
    G2982,G2983,G2984,G2985,G2986,G2987,G2988,G2989,G2990,G2991,G2992,G2993,
    G2994,G2995,G2996,G2997,G2998,G2999,G3000,G3001,G3004,G3008,G3009,G3010,
    G3013,G3016,G3020,G3021,G3022,G3025,G3028,G3031,G3034,G3037,G3040,G3043,
    G3046,G3049,G3052,G3056,G3057,G3058,G3061,G3064,G3068,G3069,G3070,G3073,
    G3077,G3081,G3085,G3089,G3093,G3097,G3101,G3105,G3109,G3113,G3114,G3115,
    G3118,G3121,G3125,G3126,G3127,G3130,G3134,G3135,G3136,G3139,G3140,G3141,
    G3144,G3145,G3146,G3149,G3150,G3151,G3154,G3155,G3156,G3159,G3160,G3161,
    G3164,G3165,G3166,G3169,G3170,G3171,G3174,G3175,G3176,G3179,G3180,G3181,
    G3184,G3187,G3191,G3192,G3193,G3196,G3200,G3201,G3202,G3205,G3208,G3211,
    G3214,G3217,G3220,G3223,G3226,G3229,G3232,G3236,G3237,G3238,G3241,G3245,
    G3246,G3247,G3250,G3253,G3257,G3261,G3265,G3269,G3273,G3277,G3281,G3285,
    G3289,G3293,G3294,G3295,G3298,G3302,G3303,G3304,G3307,G3310,G3314,G3315,
    G3316,G3317,G3318,G3319,G3320,G3321,G3322,G3323,G3324,G3325,G3326,G3327,
    G3328,G3329,G3330,G3331,G3332,G3333,G3334,G3337,G3341,G3342,G3343,G3346,
    G3349,G3353,G3354,G3355,G3358,G3361,G3364,G3367,G3370,G3373,G3376,G3379,
    G3382,G3385,G3389,G3390,G3391,G3394,G3397,G3401,G3402,G3403,G3406,G3410,
    G3414,G3418,G3422,G3426,G3430,G3434,G3438,G3442,G3446,G3447,G3448,G3451,
    G3454,G3458,G3459,G3460,G3463,G3467,G3468,G3469,G3472,G3473,G3474,G3477,
    G3478,G3479,G3482,G3483,G3484,G3487,G3488,G3489,G3492,G3493,G3494,G3497,
    G3498,G3499,G3502,G3503,G3504,G3507,G3508,G3509,G3512,G3513,G3514,G3517,
    G3520,G3524,G3525,G3526,G3529,G3533,G3534,G3535,G3538,G3541,G3545,G3548,
    G3551,G3554,G3557,G3560,G3563,G3566,G3569,G3573,G3574,G3575,G3578,G3582,
    G3583,G3584,G3587,G3590,G3594,G3595,G3596,G3600,G3604,G3608,G3612,G3616,
    G3620,G3624,G3628,G3629,G3630,G3633,G3637,G3638,G3639,G3642,G3645,G3649,
    G3650,G3651,G3654,G3655,G3656,G3657,G3658,G3659,G3660,G3661,G3662,G3663,
    G3664,G3665,G3666,G3667,G3668,G3669,G3670,G3673,G3677,G3678,G3679,G3682,
    G3685,G3689,G3690,G3691,G3694,G3698,G3701,G3704,G3707,G3710,G3713,G3716,
    G3719,G3722,G3726,G3727,G3728,G3731,G3734,G3738,G3739,G3740,G3743,G3747,
    G3748,G3749,G3752,G3756,G3760,G3764,G3768,G3772,G3776,G3780,G3784,G3785,
    G3786,G3789,G3792,G3796,G3797,G3798,G3801,G3805,G3806,G3807,G3810,G3813,
    G3817,G3818,G3819,G3822,G3823,G3824,G3827,G3828,G3829,G3832,G3833,G3834,
    G3837,G3838,G3839,G3842,G3843,G3844,G3847,G3848,G3849,G3852,G3853,G3854,
    G3857,G3860,G3864,G3865,G3866,G3869,G3873,G3874,G3875,G3878,G3881,G3885,
    G3886,G3887,G3890,G3893,G3896,G3899,G3902,G3905,G3908,G3912,G3913,G3914,
    G3917,G3921,G3922,G3923,G3926,G3929,G3933,G3934,G3935,G3938,G3942,G3946,
    G3950,G3954,G3958,G3962,G3966,G3967,G3968,G3971,G3975,G3976,G3977,G3980,
    G3983,G3987,G3988,G3989,G3992,G3996,G3997,G3998,G3999,G4000,G4001,G4002,
    G4003,G4004,G4005,G4006,G4007,G4008,G4009,G4010,G4013,G4017,G4018,G4019,
    G4022,G4025,G4029,G4030,G4031,G4034,G4038,G4039,G4040,G4043,G4046,G4049,
    G4052,G4055,G4058,G4061,G4064,G4068,G4069,G4070,G4073,G4076,G4080,G4081,
    G4082,G4085,G4089,G4090,G4091,G4094,G4097,G4101,G4105,G4109,G4113,G4117,
    G4121,G4125,G4129,G4130,G4131,G4134,G4137,G4141,G4142,G4143,G4146,G4150,
    G4151,G4152,G4155,G4158,G4162,G4163,G4164,G4165,G4166,G4169,G4170,G4171,
    G4174,G4175,G4176,G4179,G4180,G4181,G4184,G4185,G4186,G4189,G4190,G4191,
    G4194,G4195,G4196,G4199,G4202,G4206,G4207,G4208,G4211,G4215,G4216,G4217,
    G4220,G4223,G4227,G4228,G4229,G4232,G4235,G4238,G4241,G4244,G4247,G4250,
    G4254,G4255,G4256,G4259,G4263,G4264,G4265,G4268,G4271,G4275,G4276,G4277,
    G4280,G4284,G4288,G4292,G4296,G4300,G4304,G4308,G4309,G4310,G4313,G4317,
    G4318,G4319,G4322,G4325,G4329,G4330,G4331,G4334,G4338,G4339,G4340,G4343,
    G4344,G4345,G4346,G4347,G4348,G4349,G4350,G4351,G4352,G4353,G4354,G4355,
    G4358,G4362,G4363,G4364,G4367,G4370,G4374,G4375,G4376,G4379,G4383,G4384,
    G4385,G4388,G4391,G4395,G4398,G4401,G4404,G4407,G4410,G4413,G4417,G4418,
    G4419,G4422,G4425,G4429,G4430,G4431,G4434,G4438,G4439,G4440,G4443,G4446,
    G4450,G4451,G4452,G4456,G4460,G4464,G4468,G4472,G4476,G4477,G4478,G4481,
    G4484,G4488,G4489,G4490,G4493,G4497,G4498,G4499,G4502,G4505,G4509,G4510,
    G4511,G4514,G4515,G4516,G4519,G4520,G4521,G4524,G4525,G4526,G4529,G4530,
    G4531,G4534,G4535,G4536,G4539,G4540,G4541,G4544,G4547,G4551,G4552,G4553,
    G4556,G4560,G4561,G4562,G4565,G4568,G4572,G4573,G4574,G4577,G4581,G4584,
    G4587,G4590,G4593,G4596,G4600,G4601,G4602,G4605,G4609,G4610,G4611,G4614,
    G4617,G4621,G4622,G4623,G4626,G4630,G4631,G4632,G4635,G4639,G4643,G4647,
    G4651,G4655,G4656,G4657,G4660,G4664,G4665,G4666,G4669,G4672,G4676,G4677,
    G4678,G4681,G4685,G4686,G4687,G4690,G4693,G4697,G4698,G4699,G4700,G4701,
    G4702,G4703,G4704,G4705,G4706,G4707,G4710,G4714,G4715,G4716,G4719,G4722,
    G4726,G4727,G4728,G4731,G4735,G4736,G4737,G4740,G4743,G4747,G4748,G4749,
    G4752,G4755,G4758,G4761,G4764,G4768,G4769,G4770,G4773,G4776,G4780,G4781,
    G4782,G4785,G4789,G4790,G4791,G4794,G4797,G4801,G4802,G4803,G4806,G4810,
    G4814,G4818,G4822,G4826,G4827,G4828,G4831,G4834,G4838,G4839,G4840,G4843,
    G4847,G4848,G4849,G4852,G4855,G4859,G4860,G4861,G4864,G4868,G4869,G4870,
    G4873,G4874,G4875,G4878,G4879,G4880,G4883,G4884,G4885,G4888,G4889,G4890,
    G4893,G4896,G4900,G4901,G4902,G4905,G4909,G4910,G4911,G4914,G4917,G4921,
    G4922,G4923,G4926,G4930,G4931,G4932,G4935,G4938,G4941,G4944,G4947,G4951,
    G4952,G4953,G4956,G4960,G4961,G4962,G4965,G4968,G4972,G4973,G4974,G4977,
    G4981,G4982,G4983,G4986,G4989,G4993,G4997,G5001,G5005,G5009,G5010,G5011,
    G5014,G5018,G5019,G5020,G5023,G5026,G5030,G5031,G5032,G5035,G5039,G5040,
    G5041,G5044,G5047,G5051,G5052,G5053,G5054,G5055,G5056,G5057,G5058,G5059,
    G5060,G5061,G5064,G5068,G5069,G5070,G5073,G5076,G5080,G5081,G5082,G5085,
    G5089,G5090,G5091,G5094,G5097,G5101,G5102,G5103,G5106,G5109,G5112,G5115,
    G5118,G5122,G5123,G5124,G5127,G5130,G5134,G5135,G5136,G5139,G5143,G5144,
    G5145,G5148,G5151,G5155,G5156,G5157,G5160,G5164,G5168,G5172,G5176,G5180,
    G5181,G5182,G5185,G5188,G5192,G5193,G5194,G5197,G5201,G5202,G5203,G5206,
    G5209,G5213,G5214,G5215,G5218,G5222,G5223,G5224,G5227,G5228,G5229,G5232,
    G5233,G5234,G5237,G5238,G5239,G5242,G5243,G5244,G5247,G5250,G5254,G5255,
    G5256,G5259,G5263,G5264,G5265,G5268,G5271,G5275,G5276,G5277,G5280,G5284,
    G5285,G5286,G5289,G5292,G5296,G5299,G5302,G5305,G5309,G5310,G5311,G5314,
    G5318,G5319,G5320,G5323,G5326,G5330,G5331,G5332,G5335,G5339,G5340,G5341,
    G5344,G5347,G5351,G5352,G5353,G5357,G5361,G5365,G5366,G5367,G5370,G5374,
    G5375,G5376,G5379,G5382,G5386,G5387,G5388,G5391,G5395,G5396,G5397,G5400,
    G5403,G5407,G5408,G5409,G5412,G5413,G5414,G5415,G5416,G5417,G5418,G5421,
    G5425,G5426,G5427,G5430,G5433,G5437,G5438,G5439,G5442,G5446,G5447,G5448,
    G5451,G5454,G5458,G5459,G5460,G5463,G5467,G5470,G5473,G5476,G5480,G5481,
    G5482,G5485,G5488,G5492,G5493,G5494,G5497,G5501,G5502,G5503,G5506,G5509,
    G5513,G5514,G5515,G5518,G5522,G5523,G5524,G5527,G5531,G5535,G5539,G5540,
    G5541,G5544,G5547,G5551,G5552,G5553,G5556,G5560,G5561,G5562,G5565,G5568,
    G5572,G5573,G5574,G5577,G5581,G5582,G5583,G5586,G5589,G5593,G5594,G5595,
    G5598,G5599,G5600,G5603,G5604,G5605,G5608,G5611,G5615,G5616,G5617,G5620,
    G5624,G5625,G5626,G5629,G5632,G5636,G5637,G5638,G5641,G5645,G5646,G5647,
    G5650,G5653,G5657,G5658,G5659,G5662,G5665,G5669,G5670,G5671,G5674,G5678,
    G5679,G5680,G5683,G5686,G5690,G5691,G5692,G5695,G5699,G5700,G5701,G5704,
    G5707,G5711,G5712,G5713,G5716,G5720,G5724,G5725,G5726,G5729,G5733,G5734,
    G5735,G5738,G5741,G5745,G5746,G5747,G5750,G5754,G5755,G5756,G5759,G5762,
    G5766,G5767,G5768,G5771,G5772,G5773,G5774,G5775,G5778,G5782,G5783,G5784,
    G5787,G5790,G5794,G5795,G5796,G5799,G5803,G5804,G5805,G5808,G5811,G5815,
    G5816,G5817,G5820,G5823,G5826,G5830,G5831,G5832,G5835,G5838,G5842,G5843,
    G5844,G5847,G5851,G5852,G5853,G5856,G5859,G5863,G5864,G5865,G5868,G5872,
    G5876,G5877,G5878,G5881,G5884,G5888,G5889,G5890,G5893,G5897,G5898,G5899,
    G5902,G5905,G5909,G5910,G5911,G5914,G5915,G5916,G5919,G5920,G5921,G5924,
    G5927,G5931,G5932,G5933,G5936,G5940,G5941,G5942,G5945,G5948,G5952,G5953,
    G5954,G5957,G5960,G5964,G5965,G5966,G5969,G5973,G5974,G5975,G5978,G5981,
    G5985,G5986,G5987,G5990,G5994,G5995,G5996,G5999,G6003,G6004,G6005,G6008,
    G6011,G6015,G6016,G6017,G6020,G6021,G6022,G6025,G6029,G6030,G6031,G6034,
    G6037,G6041,G6042,G6043,G6046,G6049,G6053,G6054,G6055,G6058,G6061,G6065,
    G6066,G6067,G6070,G6074,G6075,G6076,G6079,G6082,G6086,G6087,G6088,G6091,
    G6092,G6093,G6096,G6099,G6103,G6104,G6105,G6108,G6112,G6113,G6114,G6117,
    G6118,G6119,G6122,G6125,G6129,G6130,G6131,G6134,G6138,G6139,G6140,G6143,
    G6147,G6148,G6149,G6152,G6156,G6157,G6158,G6161,G6165,G6166,G6167,G6170,
    G6174,G6175,G6176,G6179,G6183,G6184,G6185,G6188,G6192,G6193,G6194,G6197,
    G6201,G6202,G6203,G6206,G6210,G6211,G6212,G6215,G6219,G6220,G6221,G6224,
    G6228,G6229,G6230,G6233,G6237,G6238,G6239,G6242,G6246,G6247,G6248,G6251,
    G6255,G6256;

  and (G545,G1,G18);
  and (G548,G1,G19);
  and (G551,G1,G20);
  and (G554,G1,G21);
  and (G557,G1,G22);
  and (G560,G1,G23);
  and (G563,G1,G24);
  and (G566,G1,G25);
  and (G569,G1,G26);
  and (G572,G1,G27);
  and (G575,G1,G28);
  and (G578,G1,G29);
  and (G581,G1,G30);
  and (G584,G1,G31);
  and (G587,G1,G32);
  and (G590,G2,G17);
  and (G593,G2,G18);
  and (G596,G2,G19);
  and (G599,G2,G20);
  and (G602,G2,G21);
  and (G605,G2,G22);
  and (G608,G2,G23);
  and (G611,G2,G24);
  and (G614,G2,G25);
  and (G617,G2,G26);
  and (G620,G2,G27);
  and (G623,G2,G28);
  and (G626,G2,G29);
  and (G629,G2,G30);
  and (G632,G2,G31);
  and (G635,G2,G32);
  and (G638,G3,G17);
  and (G641,G3,G18);
  and (G644,G3,G19);
  and (G647,G3,G20);
  and (G650,G3,G21);
  and (G653,G3,G22);
  and (G656,G3,G23);
  and (G659,G3,G24);
  and (G662,G3,G25);
  and (G665,G3,G26);
  and (G668,G3,G27);
  and (G671,G3,G28);
  and (G674,G3,G29);
  and (G677,G3,G30);
  and (G680,G3,G31);
  and (G683,G3,G32);
  and (G686,G4,G17);
  and (G689,G4,G18);
  and (G692,G4,G19);
  and (G695,G4,G20);
  and (G698,G4,G21);
  and (G701,G4,G22);
  and (G704,G4,G23);
  and (G707,G4,G24);
  and (G710,G4,G25);
  and (G713,G4,G26);
  and (G716,G4,G27);
  and (G719,G4,G28);
  and (G722,G4,G29);
  and (G725,G4,G30);
  and (G728,G4,G31);
  and (G731,G4,G32);
  and (G734,G5,G17);
  and (G737,G5,G18);
  and (G740,G5,G19);
  and (G743,G5,G20);
  and (G746,G5,G21);
  and (G749,G5,G22);
  and (G752,G5,G23);
  and (G755,G5,G24);
  and (G758,G5,G25);
  and (G761,G5,G26);
  and (G764,G5,G27);
  and (G767,G5,G28);
  and (G770,G5,G29);
  and (G773,G5,G30);
  and (G776,G5,G31);
  and (G779,G5,G32);
  and (G782,G6,G17);
  and (G785,G6,G18);
  and (G788,G6,G19);
  and (G791,G6,G20);
  and (G794,G6,G21);
  and (G797,G6,G22);
  and (G800,G6,G23);
  and (G803,G6,G24);
  and (G806,G6,G25);
  and (G809,G6,G26);
  and (G812,G6,G27);
  and (G815,G6,G28);
  and (G818,G6,G29);
  and (G821,G6,G30);
  and (G824,G6,G31);
  and (G827,G6,G32);
  and (G830,G7,G17);
  and (G833,G7,G18);
  and (G836,G7,G19);
  and (G839,G7,G20);
  and (G842,G7,G21);
  and (G845,G7,G22);
  and (G848,G7,G23);
  and (G851,G7,G24);
  and (G854,G7,G25);
  and (G857,G7,G26);
  and (G860,G7,G27);
  and (G863,G7,G28);
  and (G866,G7,G29);
  and (G869,G7,G30);
  and (G872,G7,G31);
  and (G875,G7,G32);
  and (G878,G8,G17);
  and (G881,G8,G18);
  and (G884,G8,G19);
  and (G887,G8,G20);
  and (G890,G8,G21);
  and (G893,G8,G22);
  and (G896,G8,G23);
  and (G899,G8,G24);
  and (G902,G8,G25);
  and (G905,G8,G26);
  and (G908,G8,G27);
  and (G911,G8,G28);
  and (G914,G8,G29);
  and (G917,G8,G30);
  and (G920,G8,G31);
  and (G923,G8,G32);
  and (G926,G9,G17);
  and (G929,G9,G18);
  and (G932,G9,G19);
  and (G935,G9,G20);
  and (G938,G9,G21);
  and (G941,G9,G22);
  and (G944,G9,G23);
  and (G947,G9,G24);
  and (G950,G9,G25);
  and (G953,G9,G26);
  and (G956,G9,G27);
  and (G959,G9,G28);
  and (G962,G9,G29);
  and (G965,G9,G30);
  and (G968,G9,G31);
  and (G971,G9,G32);
  and (G974,G10,G17);
  and (G977,G10,G18);
  and (G980,G10,G19);
  and (G983,G10,G20);
  and (G986,G10,G21);
  and (G989,G10,G22);
  and (G992,G10,G23);
  and (G995,G10,G24);
  and (G998,G10,G25);
  and (G1001,G10,G26);
  and (G1004,G10,G27);
  and (G1007,G10,G28);
  and (G1010,G10,G29);
  and (G1013,G10,G30);
  and (G1016,G10,G31);
  and (G1019,G10,G32);
  and (G1022,G11,G17);
  and (G1025,G11,G18);
  and (G1028,G11,G19);
  and (G1031,G11,G20);
  and (G1034,G11,G21);
  and (G1037,G11,G22);
  and (G1040,G11,G23);
  and (G1043,G11,G24);
  and (G1046,G11,G25);
  and (G1049,G11,G26);
  and (G1052,G11,G27);
  and (G1055,G11,G28);
  and (G1058,G11,G29);
  and (G1061,G11,G30);
  and (G1064,G11,G31);
  and (G1067,G11,G32);
  and (G1070,G12,G17);
  and (G1073,G12,G18);
  and (G1076,G12,G19);
  and (G1079,G12,G20);
  and (G1082,G12,G21);
  and (G1085,G12,G22);
  and (G1088,G12,G23);
  and (G1091,G12,G24);
  and (G1094,G12,G25);
  and (G1097,G12,G26);
  and (G1100,G12,G27);
  and (G1103,G12,G28);
  and (G1106,G12,G29);
  and (G1109,G12,G30);
  and (G1112,G12,G31);
  and (G1115,G12,G32);
  and (G1118,G13,G17);
  and (G1121,G13,G18);
  and (G1124,G13,G19);
  and (G1127,G13,G20);
  and (G1130,G13,G21);
  and (G1133,G13,G22);
  and (G1136,G13,G23);
  and (G1139,G13,G24);
  and (G1142,G13,G25);
  and (G1145,G13,G26);
  and (G1148,G13,G27);
  and (G1151,G13,G28);
  and (G1154,G13,G29);
  and (G1157,G13,G30);
  and (G1160,G13,G31);
  and (G1163,G13,G32);
  and (G1166,G14,G17);
  and (G1169,G14,G18);
  and (G1172,G14,G19);
  and (G1175,G14,G20);
  and (G1178,G14,G21);
  and (G1181,G14,G22);
  and (G1184,G14,G23);
  and (G1187,G14,G24);
  and (G1190,G14,G25);
  and (G1193,G14,G26);
  and (G1196,G14,G27);
  and (G1199,G14,G28);
  and (G1202,G14,G29);
  and (G1205,G14,G30);
  and (G1208,G14,G31);
  and (G1211,G14,G32);
  and (G1214,G15,G17);
  and (G1217,G15,G18);
  and (G1220,G15,G19);
  and (G1223,G15,G20);
  and (G1226,G15,G21);
  and (G1229,G15,G22);
  and (G1232,G15,G23);
  and (G1235,G15,G24);
  and (G1238,G15,G25);
  and (G1241,G15,G26);
  and (G1244,G15,G27);
  and (G1247,G15,G28);
  and (G1250,G15,G29);
  and (G1253,G15,G30);
  and (G1256,G15,G31);
  and (G1259,G15,G32);
  and (G1262,G16,G17);
  and (G1265,G16,G18);
  and (G1268,G16,G19);
  and (G1271,G16,G20);
  and (G1274,G16,G21);
  and (G1277,G16,G22);
  and (G1280,G16,G23);
  and (G1283,G16,G24);
  and (G1286,G16,G25);
  and (G1289,G16,G26);
  and (G1292,G16,G27);
  and (G1295,G16,G28);
  and (G1298,G16,G29);
  and (G1301,G16,G30);
  and (G1304,G16,G31);
  and (G1307,G16,G32);
  not (G1310,G590);
  not (G1314,G638);
  not (G1318,G686);
  not (G1322,G734);
  not (G1326,G782);
  not (G1330,G830);
  not (G1334,G878);
  not (G1338,G926);
  not (G1342,G974);
  not (G1346,G1022);
  not (G1350,G1070);
  not (G1354,G1118);
  not (G1358,G1166);
  not (G1362,G1214);
  not (G1366,G1262);
  nor (G1370,G590,G1310);
  not (G1371,G1310);
  nor (G1372,G638,G1314);
  not (G1373,G1314);
  nor (G1374,G686,G1318);
  not (G1375,G1318);
  nor (G1376,G734,G1322);
  not (G1377,G1322);
  nor (G1378,G782,G1326);
  not (G1379,G1326);
  nor (G1380,G830,G1330);
  not (G1381,G1330);
  nor (G1382,G878,G1334);
  not (G1383,G1334);
  nor (G1384,G926,G1338);
  not (G1385,G1338);
  nor (G1386,G974,G1342);
  not (G1387,G1342);
  nor (G1388,G1022,G1346);
  not (G1389,G1346);
  nor (G1390,G1070,G1350);
  not (G1391,G1350);
  nor (G1392,G1118,G1354);
  not (G1393,G1354);
  nor (G1394,G1166,G1358);
  not (G1395,G1358);
  nor (G1396,G1214,G1362);
  not (G1397,G1362);
  nor (G1398,G1262,G1366);
  not (G1399,G1366);
  nor (G1400,G1370,G1371);
  nor (G1403,G1372,G1373);
  nor (G1406,G1374,G1375);
  nor (G1409,G1376,G1377);
  nor (G1412,G1378,G1379);
  nor (G1415,G1380,G1381);
  nor (G1418,G1382,G1383);
  nor (G1421,G1384,G1385);
  nor (G1424,G1386,G1387);
  nor (G1427,G1388,G1389);
  nor (G1430,G1390,G1391);
  nor (G1433,G1392,G1393);
  nor (G1436,G1394,G1395);
  nor (G1439,G1396,G1397);
  nor (G1442,G1398,G1399);
  nor (G1445,G1400,G545);
  nor (G1449,G1403,G593);
  nor (G1453,G1406,G641);
  nor (G1457,G1409,G689);
  nor (G1461,G1412,G737);
  nor (G1465,G1415,G785);
  nor (G1469,G1418,G833);
  nor (G1473,G1421,G881);
  nor (G1477,G1424,G929);
  nor (G1481,G1427,G977);
  nor (G1485,G1430,G1025);
  nor (G1489,G1433,G1073);
  nor (G1493,G1436,G1121);
  nor (G1497,G1439,G1169);
  nor (G1501,G1442,G1217);
  nor (G1505,G1400,G1445);
  nor (G1506,G1445,G545);
  nor (G1507,G1310,G1445);
  nor (G1510,G1403,G1449);
  nor (G1511,G1449,G593);
  nor (G1512,G1314,G1449);
  nor (G1515,G1406,G1453);
  nor (G1516,G1453,G641);
  nor (G1517,G1318,G1453);
  nor (G1520,G1409,G1457);
  nor (G1521,G1457,G689);
  nor (G1522,G1322,G1457);
  nor (G1525,G1412,G1461);
  nor (G1526,G1461,G737);
  nor (G1527,G1326,G1461);
  nor (G1530,G1415,G1465);
  nor (G1531,G1465,G785);
  nor (G1532,G1330,G1465);
  nor (G1535,G1418,G1469);
  nor (G1536,G1469,G833);
  nor (G1537,G1334,G1469);
  nor (G1540,G1421,G1473);
  nor (G1541,G1473,G881);
  nor (G1542,G1338,G1473);
  nor (G1545,G1424,G1477);
  nor (G1546,G1477,G929);
  nor (G1547,G1342,G1477);
  nor (G1550,G1427,G1481);
  nor (G1551,G1481,G977);
  nor (G1552,G1346,G1481);
  nor (G1555,G1430,G1485);
  nor (G1556,G1485,G1025);
  nor (G1557,G1350,G1485);
  nor (G1560,G1433,G1489);
  nor (G1561,G1489,G1073);
  nor (G1562,G1354,G1489);
  nor (G1565,G1436,G1493);
  nor (G1566,G1493,G1121);
  nor (G1567,G1358,G1493);
  nor (G1570,G1439,G1497);
  nor (G1571,G1497,G1169);
  nor (G1572,G1362,G1497);
  nor (G1575,G1442,G1501);
  nor (G1576,G1501,G1217);
  nor (G1577,G1366,G1501);
  nor (G1580,G1510,G1511);
  nor (G1583,G1515,G1516);
  nor (G1586,G1520,G1521);
  nor (G1589,G1525,G1526);
  nor (G1592,G1530,G1531);
  nor (G1595,G1535,G1536);
  nor (G1598,G1540,G1541);
  nor (G1601,G1545,G1546);
  nor (G1604,G1550,G1551);
  nor (G1607,G1555,G1556);
  nor (G1610,G1560,G1561);
  nor (G1613,G1565,G1566);
  nor (G1616,G1570,G1571);
  nor (G1619,G1575,G1576);
  nor (G1622,G1265,G1577);
  nor (G1626,G1580,G1507);
  nor (G1630,G1583,G1512);
  nor (G1634,G1586,G1517);
  nor (G1638,G1589,G1522);
  nor (G1642,G1592,G1527);
  nor (G1646,G1595,G1532);
  nor (G1650,G1598,G1537);
  nor (G1654,G1601,G1542);
  nor (G1658,G1604,G1547);
  nor (G1662,G1607,G1552);
  nor (G1666,G1610,G1557);
  nor (G1670,G1613,G1562);
  nor (G1674,G1616,G1567);
  nor (G1678,G1619,G1572);
  nor (G1682,G1265,G1622);
  nor (G1683,G1622,G1577);
  nor (G1684,G1580,G1626);
  nor (G1685,G1626,G1507);
  nor (G1686,G1583,G1630);
  nor (G1687,G1630,G1512);
  nor (G1688,G1586,G1634);
  nor (G1689,G1634,G1517);
  nor (G1690,G1589,G1638);
  nor (G1691,G1638,G1522);
  nor (G1692,G1592,G1642);
  nor (G1693,G1642,G1527);
  nor (G1694,G1595,G1646);
  nor (G1695,G1646,G1532);
  nor (G1696,G1598,G1650);
  nor (G1697,G1650,G1537);
  nor (G1698,G1601,G1654);
  nor (G1699,G1654,G1542);
  nor (G1700,G1604,G1658);
  nor (G1701,G1658,G1547);
  nor (G1702,G1607,G1662);
  nor (G1703,G1662,G1552);
  nor (G1704,G1610,G1666);
  nor (G1705,G1666,G1557);
  nor (G1706,G1613,G1670);
  nor (G1707,G1670,G1562);
  nor (G1708,G1616,G1674);
  nor (G1709,G1674,G1567);
  nor (G1710,G1619,G1678);
  nor (G1711,G1678,G1572);
  nor (G1712,G1682,G1683);
  nor (G1715,G1684,G1685);
  nor (G1718,G1686,G1687);
  nor (G1721,G1688,G1689);
  nor (G1724,G1690,G1691);
  nor (G1727,G1692,G1693);
  nor (G1730,G1694,G1695);
  nor (G1733,G1696,G1697);
  nor (G1736,G1698,G1699);
  nor (G1739,G1700,G1701);
  nor (G1742,G1702,G1703);
  nor (G1745,G1704,G1705);
  nor (G1748,G1706,G1707);
  nor (G1751,G1708,G1709);
  nor (G1754,G1710,G1711);
  nor (G1757,G1712,G1220);
  nor (G1761,G1715,G548);
  nor (G1765,G1718,G596);
  nor (G1769,G1721,G644);
  nor (G1773,G1724,G692);
  nor (G1777,G1727,G740);
  nor (G1781,G1730,G788);
  nor (G1785,G1733,G836);
  nor (G1789,G1736,G884);
  nor (G1793,G1739,G932);
  nor (G1797,G1742,G980);
  nor (G1801,G1745,G1028);
  nor (G1805,G1748,G1076);
  nor (G1809,G1751,G1124);
  nor (G1813,G1754,G1172);
  nor (G1817,G1712,G1757);
  nor (G1818,G1757,G1220);
  nor (G1819,G1622,G1757);
  nor (G1822,G1715,G1761);
  nor (G1823,G1761,G548);
  nor (G1824,G1626,G1761);
  nor (G1827,G1718,G1765);
  nor (G1828,G1765,G596);
  nor (G1829,G1630,G1765);
  nor (G1832,G1721,G1769);
  nor (G1833,G1769,G644);
  nor (G1834,G1634,G1769);
  nor (G1837,G1724,G1773);
  nor (G1838,G1773,G692);
  nor (G1839,G1638,G1773);
  nor (G1842,G1727,G1777);
  nor (G1843,G1777,G740);
  nor (G1844,G1642,G1777);
  nor (G1847,G1730,G1781);
  nor (G1848,G1781,G788);
  nor (G1849,G1646,G1781);
  nor (G1852,G1733,G1785);
  nor (G1853,G1785,G836);
  nor (G1854,G1650,G1785);
  nor (G1857,G1736,G1789);
  nor (G1858,G1789,G884);
  nor (G1859,G1654,G1789);
  nor (G1862,G1739,G1793);
  nor (G1863,G1793,G932);
  nor (G1864,G1658,G1793);
  nor (G1867,G1742,G1797);
  nor (G1868,G1797,G980);
  nor (G1869,G1662,G1797);
  nor (G1872,G1745,G1801);
  nor (G1873,G1801,G1028);
  nor (G1874,G1666,G1801);
  nor (G1877,G1748,G1805);
  nor (G1878,G1805,G1076);
  nor (G1879,G1670,G1805);
  nor (G1882,G1751,G1809);
  nor (G1883,G1809,G1124);
  nor (G1884,G1674,G1809);
  nor (G1887,G1754,G1813);
  nor (G1888,G1813,G1172);
  nor (G1889,G1678,G1813);
  nor (G1892,G1817,G1818);
  nor (G1895,G1268,G1819);
  nor (G1899,G1827,G1828);
  nor (G1902,G1832,G1833);
  nor (G1905,G1837,G1838);
  nor (G1908,G1842,G1843);
  nor (G1911,G1847,G1848);
  nor (G1914,G1852,G1853);
  nor (G1917,G1857,G1858);
  nor (G1920,G1862,G1863);
  nor (G1923,G1867,G1868);
  nor (G1926,G1872,G1873);
  nor (G1929,G1877,G1878);
  nor (G1932,G1882,G1883);
  nor (G1935,G1887,G1888);
  nor (G1938,G1892,G1889);
  nor (G1942,G1268,G1895);
  nor (G1943,G1895,G1819);
  nor (G1944,G1899,G1824);
  nor (G1948,G1902,G1829);
  nor (G1952,G1905,G1834);
  nor (G1956,G1908,G1839);
  nor (G1960,G1911,G1844);
  nor (G1964,G1914,G1849);
  nor (G1968,G1917,G1854);
  nor (G1972,G1920,G1859);
  nor (G1976,G1923,G1864);
  nor (G1980,G1926,G1869);
  nor (G1984,G1929,G1874);
  nor (G1988,G1932,G1879);
  nor (G1992,G1935,G1884);
  nor (G1996,G1892,G1938);
  nor (G1997,G1938,G1889);
  nor (G1998,G1942,G1943);
  nor (G2001,G1899,G1944);
  nor (G2002,G1944,G1824);
  nor (G2003,G1902,G1948);
  nor (G2004,G1948,G1829);
  nor (G2005,G1905,G1952);
  nor (G2006,G1952,G1834);
  nor (G2007,G1908,G1956);
  nor (G2008,G1956,G1839);
  nor (G2009,G1911,G1960);
  nor (G2010,G1960,G1844);
  nor (G2011,G1914,G1964);
  nor (G2012,G1964,G1849);
  nor (G2013,G1917,G1968);
  nor (G2014,G1968,G1854);
  nor (G2015,G1920,G1972);
  nor (G2016,G1972,G1859);
  nor (G2017,G1923,G1976);
  nor (G2018,G1976,G1864);
  nor (G2019,G1926,G1980);
  nor (G2020,G1980,G1869);
  nor (G2021,G1929,G1984);
  nor (G2022,G1984,G1874);
  nor (G2023,G1932,G1988);
  nor (G2024,G1988,G1879);
  nor (G2025,G1935,G1992);
  nor (G2026,G1992,G1884);
  nor (G2027,G1996,G1997);
  nor (G2030,G1998,G1223);
  nor (G2034,G2001,G2002);
  nor (G2037,G2003,G2004);
  nor (G2040,G2005,G2006);
  nor (G2043,G2007,G2008);
  nor (G2046,G2009,G2010);
  nor (G2049,G2011,G2012);
  nor (G2052,G2013,G2014);
  nor (G2055,G2015,G2016);
  nor (G2058,G2017,G2018);
  nor (G2061,G2019,G2020);
  nor (G2064,G2021,G2022);
  nor (G2067,G2023,G2024);
  nor (G2070,G2025,G2026);
  nor (G2073,G2027,G1175);
  nor (G2077,G1998,G2030);
  nor (G2078,G2030,G1223);
  nor (G2079,G1895,G2030);
  nor (G2082,G2034,G551);
  nor (G2086,G2037,G599);
  nor (G2090,G2040,G647);
  nor (G2094,G2043,G695);
  nor (G2098,G2046,G743);
  nor (G2102,G2049,G791);
  nor (G2106,G2052,G839);
  nor (G2110,G2055,G887);
  nor (G2114,G2058,G935);
  nor (G2118,G2061,G983);
  nor (G2122,G2064,G1031);
  nor (G2126,G2067,G1079);
  nor (G2130,G2070,G1127);
  nor (G2134,G2027,G2073);
  nor (G2135,G2073,G1175);
  nor (G2136,G1938,G2073);
  nor (G2139,G2077,G2078);
  nor (G2142,G1271,G2079);
  nor (G2146,G2034,G2082);
  nor (G2147,G2082,G551);
  nor (G2148,G1944,G2082);
  nor (G2151,G2037,G2086);
  nor (G2152,G2086,G599);
  nor (G2153,G1948,G2086);
  nor (G2156,G2040,G2090);
  nor (G2157,G2090,G647);
  nor (G2158,G1952,G2090);
  nor (G2161,G2043,G2094);
  nor (G2162,G2094,G695);
  nor (G2163,G1956,G2094);
  nor (G2166,G2046,G2098);
  nor (G2167,G2098,G743);
  nor (G2168,G1960,G2098);
  nor (G2171,G2049,G2102);
  nor (G2172,G2102,G791);
  nor (G2173,G1964,G2102);
  nor (G2176,G2052,G2106);
  nor (G2177,G2106,G839);
  nor (G2178,G1968,G2106);
  nor (G2181,G2055,G2110);
  nor (G2182,G2110,G887);
  nor (G2183,G1972,G2110);
  nor (G2186,G2058,G2114);
  nor (G2187,G2114,G935);
  nor (G2188,G1976,G2114);
  nor (G2191,G2061,G2118);
  nor (G2192,G2118,G983);
  nor (G2193,G1980,G2118);
  nor (G2196,G2064,G2122);
  nor (G2197,G2122,G1031);
  nor (G2198,G1984,G2122);
  nor (G2201,G2067,G2126);
  nor (G2202,G2126,G1079);
  nor (G2203,G1988,G2126);
  nor (G2206,G2070,G2130);
  nor (G2207,G2130,G1127);
  nor (G2208,G1992,G2130);
  nor (G2211,G2134,G2135);
  nor (G2214,G2139,G2136);
  nor (G2218,G1271,G2142);
  nor (G2219,G2142,G2079);
  nor (G2220,G2151,G2152);
  nor (G2223,G2156,G2157);
  nor (G2226,G2161,G2162);
  nor (G2229,G2166,G2167);
  nor (G2232,G2171,G2172);
  nor (G2235,G2176,G2177);
  nor (G2238,G2181,G2182);
  nor (G2241,G2186,G2187);
  nor (G2244,G2191,G2192);
  nor (G2247,G2196,G2197);
  nor (G2250,G2201,G2202);
  nor (G2253,G2206,G2207);
  nor (G2256,G2211,G2208);
  nor (G2260,G2139,G2214);
  nor (G2261,G2214,G2136);
  nor (G2262,G2218,G2219);
  nor (G2265,G2220,G2148);
  nor (G2269,G2223,G2153);
  nor (G2273,G2226,G2158);
  nor (G2277,G2229,G2163);
  nor (G2281,G2232,G2168);
  nor (G2285,G2235,G2173);
  nor (G2289,G2238,G2178);
  nor (G2293,G2241,G2183);
  nor (G2297,G2244,G2188);
  nor (G2301,G2247,G2193);
  nor (G2305,G2250,G2198);
  nor (G2309,G2253,G2203);
  nor (G2313,G2211,G2256);
  nor (G2314,G2256,G2208);
  nor (G2315,G2260,G2261);
  nor (G2318,G2262,G1226);
  nor (G2322,G2220,G2265);
  nor (G2323,G2265,G2148);
  nor (G2324,G2223,G2269);
  nor (G2325,G2269,G2153);
  nor (G2326,G2226,G2273);
  nor (G2327,G2273,G2158);
  nor (G2328,G2229,G2277);
  nor (G2329,G2277,G2163);
  nor (G2330,G2232,G2281);
  nor (G2331,G2281,G2168);
  nor (G2332,G2235,G2285);
  nor (G2333,G2285,G2173);
  nor (G2334,G2238,G2289);
  nor (G2335,G2289,G2178);
  nor (G2336,G2241,G2293);
  nor (G2337,G2293,G2183);
  nor (G2338,G2244,G2297);
  nor (G2339,G2297,G2188);
  nor (G2340,G2247,G2301);
  nor (G2341,G2301,G2193);
  nor (G2342,G2250,G2305);
  nor (G2343,G2305,G2198);
  nor (G2344,G2253,G2309);
  nor (G2345,G2309,G2203);
  nor (G2346,G2313,G2314);
  nor (G2349,G2315,G1178);
  nor (G2353,G2262,G2318);
  nor (G2354,G2318,G1226);
  nor (G2355,G2142,G2318);
  nor (G2358,G2322,G2323);
  nor (G2361,G2324,G2325);
  nor (G2364,G2326,G2327);
  nor (G2367,G2328,G2329);
  nor (G2370,G2330,G2331);
  nor (G2373,G2332,G2333);
  nor (G2376,G2334,G2335);
  nor (G2379,G2336,G2337);
  nor (G2382,G2338,G2339);
  nor (G2385,G2340,G2341);
  nor (G2388,G2342,G2343);
  nor (G2391,G2344,G2345);
  nor (G2394,G2346,G1130);
  nor (G2398,G2315,G2349);
  nor (G2399,G2349,G1178);
  nor (G2400,G2214,G2349);
  nor (G2403,G2353,G2354);
  nor (G2406,G1274,G2355);
  nor (G2410,G2358,G554);
  nor (G2414,G2361,G602);
  nor (G2418,G2364,G650);
  nor (G2422,G2367,G698);
  nor (G2426,G2370,G746);
  nor (G2430,G2373,G794);
  nor (G2434,G2376,G842);
  nor (G2438,G2379,G890);
  nor (G2442,G2382,G938);
  nor (G2446,G2385,G986);
  nor (G2450,G2388,G1034);
  nor (G2454,G2391,G1082);
  nor (G2458,G2346,G2394);
  nor (G2459,G2394,G1130);
  nor (G2460,G2256,G2394);
  nor (G2463,G2398,G2399);
  nor (G2466,G2403,G2400);
  nor (G2470,G1274,G2406);
  nor (G2471,G2406,G2355);
  nor (G2472,G2358,G2410);
  nor (G2473,G2410,G554);
  nor (G2474,G2265,G2410);
  nor (G2477,G2361,G2414);
  nor (G2478,G2414,G602);
  nor (G2479,G2269,G2414);
  nor (G2482,G2364,G2418);
  nor (G2483,G2418,G650);
  nor (G2484,G2273,G2418);
  nor (G2487,G2367,G2422);
  nor (G2488,G2422,G698);
  nor (G2489,G2277,G2422);
  nor (G2492,G2370,G2426);
  nor (G2493,G2426,G746);
  nor (G2494,G2281,G2426);
  nor (G2497,G2373,G2430);
  nor (G2498,G2430,G794);
  nor (G2499,G2285,G2430);
  nor (G2502,G2376,G2434);
  nor (G2503,G2434,G842);
  nor (G2504,G2289,G2434);
  nor (G2507,G2379,G2438);
  nor (G2508,G2438,G890);
  nor (G2509,G2293,G2438);
  nor (G2512,G2382,G2442);
  nor (G2513,G2442,G938);
  nor (G2514,G2297,G2442);
  nor (G2517,G2385,G2446);
  nor (G2518,G2446,G986);
  nor (G2519,G2301,G2446);
  nor (G2522,G2388,G2450);
  nor (G2523,G2450,G1034);
  nor (G2524,G2305,G2450);
  nor (G2527,G2391,G2454);
  nor (G2528,G2454,G1082);
  nor (G2529,G2309,G2454);
  nor (G2532,G2458,G2459);
  nor (G2535,G2463,G2460);
  nor (G2539,G2403,G2466);
  nor (G2540,G2466,G2400);
  nor (G2541,G2470,G2471);
  nor (G2544,G2477,G2478);
  nor (G2547,G2482,G2483);
  nor (G2550,G2487,G2488);
  nor (G2553,G2492,G2493);
  nor (G2556,G2497,G2498);
  nor (G2559,G2502,G2503);
  nor (G2562,G2507,G2508);
  nor (G2565,G2512,G2513);
  nor (G2568,G2517,G2518);
  nor (G2571,G2522,G2523);
  nor (G2574,G2527,G2528);
  nor (G2577,G2532,G2529);
  nor (G2581,G2463,G2535);
  nor (G2582,G2535,G2460);
  nor (G2583,G2539,G2540);
  nor (G2586,G2541,G1229);
  nor (G2590,G2544,G2474);
  nor (G2594,G2547,G2479);
  nor (G2598,G2550,G2484);
  nor (G2602,G2553,G2489);
  nor (G2606,G2556,G2494);
  nor (G2610,G2559,G2499);
  nor (G2614,G2562,G2504);
  nor (G2618,G2565,G2509);
  nor (G2622,G2568,G2514);
  nor (G2626,G2571,G2519);
  nor (G2630,G2574,G2524);
  nor (G2634,G2532,G2577);
  nor (G2635,G2577,G2529);
  nor (G2636,G2581,G2582);
  nor (G2639,G2583,G1181);
  nor (G2643,G2541,G2586);
  nor (G2644,G2586,G1229);
  nor (G2645,G2406,G2586);
  nor (G2648,G2544,G2590);
  nor (G2649,G2590,G2474);
  nor (G2650,G2547,G2594);
  nor (G2651,G2594,G2479);
  nor (G2652,G2550,G2598);
  nor (G2653,G2598,G2484);
  nor (G2654,G2553,G2602);
  nor (G2655,G2602,G2489);
  nor (G2656,G2556,G2606);
  nor (G2657,G2606,G2494);
  nor (G2658,G2559,G2610);
  nor (G2659,G2610,G2499);
  nor (G2660,G2562,G2614);
  nor (G2661,G2614,G2504);
  nor (G2662,G2565,G2618);
  nor (G2663,G2618,G2509);
  nor (G2664,G2568,G2622);
  nor (G2665,G2622,G2514);
  nor (G2666,G2571,G2626);
  nor (G2667,G2626,G2519);
  nor (G2668,G2574,G2630);
  nor (G2669,G2630,G2524);
  nor (G2670,G2634,G2635);
  nor (G2673,G2636,G1133);
  nor (G2677,G2583,G2639);
  nor (G2678,G2639,G1181);
  nor (G2679,G2466,G2639);
  nor (G2682,G2643,G2644);
  nor (G2685,G1277,G2645);
  nor (G2689,G2648,G2649);
  nor (G2692,G2650,G2651);
  nor (G2695,G2652,G2653);
  nor (G2698,G2654,G2655);
  nor (G2701,G2656,G2657);
  nor (G2704,G2658,G2659);
  nor (G2707,G2660,G2661);
  nor (G2710,G2662,G2663);
  nor (G2713,G2664,G2665);
  nor (G2716,G2666,G2667);
  nor (G2719,G2668,G2669);
  nor (G2722,G2670,G1085);
  nor (G2726,G2636,G2673);
  nor (G2727,G2673,G1133);
  nor (G2728,G2535,G2673);
  nor (G2731,G2677,G2678);
  nor (G2734,G2682,G2679);
  nor (G2738,G1277,G2685);
  nor (G2739,G2685,G2645);
  nor (G2740,G2689,G557);
  nor (G2744,G2692,G605);
  nor (G2748,G2695,G653);
  nor (G2752,G2698,G701);
  nor (G2756,G2701,G749);
  nor (G2760,G2704,G797);
  nor (G2764,G2707,G845);
  nor (G2768,G2710,G893);
  nor (G2772,G2713,G941);
  nor (G2776,G2716,G989);
  nor (G2780,G2719,G1037);
  nor (G2784,G2670,G2722);
  nor (G2785,G2722,G1085);
  nor (G2786,G2577,G2722);
  nor (G2789,G2726,G2727);
  nor (G2792,G2731,G2728);
  nor (G2796,G2682,G2734);
  nor (G2797,G2734,G2679);
  nor (G2798,G2738,G2739);
  nor (G2801,G2689,G2740);
  nor (G2802,G2740,G557);
  nor (G2803,G2590,G2740);
  nor (G2806,G2692,G2744);
  nor (G2807,G2744,G605);
  nor (G2808,G2594,G2744);
  nor (G2811,G2695,G2748);
  nor (G2812,G2748,G653);
  nor (G2813,G2598,G2748);
  nor (G2816,G2698,G2752);
  nor (G2817,G2752,G701);
  nor (G2818,G2602,G2752);
  nor (G2821,G2701,G2756);
  nor (G2822,G2756,G749);
  nor (G2823,G2606,G2756);
  nor (G2826,G2704,G2760);
  nor (G2827,G2760,G797);
  nor (G2828,G2610,G2760);
  nor (G2831,G2707,G2764);
  nor (G2832,G2764,G845);
  nor (G2833,G2614,G2764);
  nor (G2836,G2710,G2768);
  nor (G2837,G2768,G893);
  nor (G2838,G2618,G2768);
  nor (G2841,G2713,G2772);
  nor (G2842,G2772,G941);
  nor (G2843,G2622,G2772);
  nor (G2846,G2716,G2776);
  nor (G2847,G2776,G989);
  nor (G2848,G2626,G2776);
  nor (G2851,G2719,G2780);
  nor (G2852,G2780,G1037);
  nor (G2853,G2630,G2780);
  nor (G2856,G2784,G2785);
  nor (G2859,G2789,G2786);
  nor (G2863,G2731,G2792);
  nor (G2864,G2792,G2728);
  nor (G2865,G2796,G2797);
  nor (G2868,G2798,G1232);
  nor (G2872,G2806,G2807);
  nor (G2875,G2811,G2812);
  nor (G2878,G2816,G2817);
  nor (G2881,G2821,G2822);
  nor (G2884,G2826,G2827);
  nor (G2887,G2831,G2832);
  nor (G2890,G2836,G2837);
  nor (G2893,G2841,G2842);
  nor (G2896,G2846,G2847);
  nor (G2899,G2851,G2852);
  nor (G2902,G2856,G2853);
  nor (G2906,G2789,G2859);
  nor (G2907,G2859,G2786);
  nor (G2908,G2863,G2864);
  nor (G2911,G2865,G1184);
  nor (G2915,G2798,G2868);
  nor (G2916,G2868,G1232);
  nor (G2917,G2685,G2868);
  nor (G2920,G2872,G2803);
  nor (G2924,G2875,G2808);
  nor (G2928,G2878,G2813);
  nor (G2932,G2881,G2818);
  nor (G2936,G2884,G2823);
  nor (G2940,G2887,G2828);
  nor (G2944,G2890,G2833);
  nor (G2948,G2893,G2838);
  nor (G2952,G2896,G2843);
  nor (G2956,G2899,G2848);
  nor (G2960,G2856,G2902);
  nor (G2961,G2902,G2853);
  nor (G2962,G2906,G2907);
  nor (G2965,G2908,G1136);
  nor (G2969,G2865,G2911);
  nor (G2970,G2911,G1184);
  nor (G2971,G2734,G2911);
  nor (G2974,G2915,G2916);
  nor (G2977,G1280,G2917);
  nor (G2981,G2872,G2920);
  nor (G2982,G2920,G2803);
  nor (G2983,G2875,G2924);
  nor (G2984,G2924,G2808);
  nor (G2985,G2878,G2928);
  nor (G2986,G2928,G2813);
  nor (G2987,G2881,G2932);
  nor (G2988,G2932,G2818);
  nor (G2989,G2884,G2936);
  nor (G2990,G2936,G2823);
  nor (G2991,G2887,G2940);
  nor (G2992,G2940,G2828);
  nor (G2993,G2890,G2944);
  nor (G2994,G2944,G2833);
  nor (G2995,G2893,G2948);
  nor (G2996,G2948,G2838);
  nor (G2997,G2896,G2952);
  nor (G2998,G2952,G2843);
  nor (G2999,G2899,G2956);
  nor (G3000,G2956,G2848);
  nor (G3001,G2960,G2961);
  nor (G3004,G2962,G1088);
  nor (G3008,G2908,G2965);
  nor (G3009,G2965,G1136);
  nor (G3010,G2792,G2965);
  nor (G3013,G2969,G2970);
  nor (G3016,G2974,G2971);
  nor (G3020,G1280,G2977);
  nor (G3021,G2977,G2917);
  nor (G3022,G2981,G2982);
  nor (G3025,G2983,G2984);
  nor (G3028,G2985,G2986);
  nor (G3031,G2987,G2988);
  nor (G3034,G2989,G2990);
  nor (G3037,G2991,G2992);
  nor (G3040,G2993,G2994);
  nor (G3043,G2995,G2996);
  nor (G3046,G2997,G2998);
  nor (G3049,G2999,G3000);
  nor (G3052,G3001,G1040);
  nor (G3056,G2962,G3004);
  nor (G3057,G3004,G1088);
  nor (G3058,G2859,G3004);
  nor (G3061,G3008,G3009);
  nor (G3064,G3013,G3010);
  nor (G3068,G2974,G3016);
  nor (G3069,G3016,G2971);
  nor (G3070,G3020,G3021);
  nor (G3073,G3022,G560);
  nor (G3077,G3025,G608);
  nor (G3081,G3028,G656);
  nor (G3085,G3031,G704);
  nor (G3089,G3034,G752);
  nor (G3093,G3037,G800);
  nor (G3097,G3040,G848);
  nor (G3101,G3043,G896);
  nor (G3105,G3046,G944);
  nor (G3109,G3049,G992);
  nor (G3113,G3001,G3052);
  nor (G3114,G3052,G1040);
  nor (G3115,G2902,G3052);
  nor (G3118,G3056,G3057);
  nor (G3121,G3061,G3058);
  nor (G3125,G3013,G3064);
  nor (G3126,G3064,G3010);
  nor (G3127,G3068,G3069);
  nor (G3130,G3070,G1235);
  nor (G3134,G3022,G3073);
  nor (G3135,G3073,G560);
  nor (G3136,G2920,G3073);
  nor (G3139,G3025,G3077);
  nor (G3140,G3077,G608);
  nor (G3141,G2924,G3077);
  nor (G3144,G3028,G3081);
  nor (G3145,G3081,G656);
  nor (G3146,G2928,G3081);
  nor (G3149,G3031,G3085);
  nor (G3150,G3085,G704);
  nor (G3151,G2932,G3085);
  nor (G3154,G3034,G3089);
  nor (G3155,G3089,G752);
  nor (G3156,G2936,G3089);
  nor (G3159,G3037,G3093);
  nor (G3160,G3093,G800);
  nor (G3161,G2940,G3093);
  nor (G3164,G3040,G3097);
  nor (G3165,G3097,G848);
  nor (G3166,G2944,G3097);
  nor (G3169,G3043,G3101);
  nor (G3170,G3101,G896);
  nor (G3171,G2948,G3101);
  nor (G3174,G3046,G3105);
  nor (G3175,G3105,G944);
  nor (G3176,G2952,G3105);
  nor (G3179,G3049,G3109);
  nor (G3180,G3109,G992);
  nor (G3181,G2956,G3109);
  nor (G3184,G3113,G3114);
  nor (G3187,G3118,G3115);
  nor (G3191,G3061,G3121);
  nor (G3192,G3121,G3058);
  nor (G3193,G3125,G3126);
  nor (G3196,G3127,G1187);
  nor (G3200,G3070,G3130);
  nor (G3201,G3130,G1235);
  nor (G3202,G2977,G3130);
  nor (G3205,G3139,G3140);
  nor (G3208,G3144,G3145);
  nor (G3211,G3149,G3150);
  nor (G3214,G3154,G3155);
  nor (G3217,G3159,G3160);
  nor (G3220,G3164,G3165);
  nor (G3223,G3169,G3170);
  nor (G3226,G3174,G3175);
  nor (G3229,G3179,G3180);
  nor (G3232,G3184,G3181);
  nor (G3236,G3118,G3187);
  nor (G3237,G3187,G3115);
  nor (G3238,G3191,G3192);
  nor (G3241,G3193,G1139);
  nor (G3245,G3127,G3196);
  nor (G3246,G3196,G1187);
  nor (G3247,G3016,G3196);
  nor (G3250,G3200,G3201);
  nor (G3253,G1283,G3202);
  nor (G3257,G3205,G3136);
  nor (G3261,G3208,G3141);
  nor (G3265,G3211,G3146);
  nor (G3269,G3214,G3151);
  nor (G3273,G3217,G3156);
  nor (G3277,G3220,G3161);
  nor (G3281,G3223,G3166);
  nor (G3285,G3226,G3171);
  nor (G3289,G3229,G3176);
  nor (G3293,G3184,G3232);
  nor (G3294,G3232,G3181);
  nor (G3295,G3236,G3237);
  nor (G3298,G3238,G1091);
  nor (G3302,G3193,G3241);
  nor (G3303,G3241,G1139);
  nor (G3304,G3064,G3241);
  nor (G3307,G3245,G3246);
  nor (G3310,G3250,G3247);
  nor (G3314,G1283,G3253);
  nor (G3315,G3253,G3202);
  nor (G3316,G3205,G3257);
  nor (G3317,G3257,G3136);
  nor (G3318,G3208,G3261);
  nor (G3319,G3261,G3141);
  nor (G3320,G3211,G3265);
  nor (G3321,G3265,G3146);
  nor (G3322,G3214,G3269);
  nor (G3323,G3269,G3151);
  nor (G3324,G3217,G3273);
  nor (G3325,G3273,G3156);
  nor (G3326,G3220,G3277);
  nor (G3327,G3277,G3161);
  nor (G3328,G3223,G3281);
  nor (G3329,G3281,G3166);
  nor (G3330,G3226,G3285);
  nor (G3331,G3285,G3171);
  nor (G3332,G3229,G3289);
  nor (G3333,G3289,G3176);
  nor (G3334,G3293,G3294);
  nor (G3337,G3295,G1043);
  nor (G3341,G3238,G3298);
  nor (G3342,G3298,G1091);
  nor (G3343,G3121,G3298);
  nor (G3346,G3302,G3303);
  nor (G3349,G3307,G3304);
  nor (G3353,G3250,G3310);
  nor (G3354,G3310,G3247);
  nor (G3355,G3314,G3315);
  nor (G3358,G3316,G3317);
  nor (G3361,G3318,G3319);
  nor (G3364,G3320,G3321);
  nor (G3367,G3322,G3323);
  nor (G3370,G3324,G3325);
  nor (G3373,G3326,G3327);
  nor (G3376,G3328,G3329);
  nor (G3379,G3330,G3331);
  nor (G3382,G3332,G3333);
  nor (G3385,G3334,G995);
  nor (G3389,G3295,G3337);
  nor (G3390,G3337,G1043);
  nor (G3391,G3187,G3337);
  nor (G3394,G3341,G3342);
  nor (G3397,G3346,G3343);
  nor (G3401,G3307,G3349);
  nor (G3402,G3349,G3304);
  nor (G3403,G3353,G3354);
  nor (G3406,G3355,G1238);
  nor (G3410,G3358,G563);
  nor (G3414,G3361,G611);
  nor (G3418,G3364,G659);
  nor (G3422,G3367,G707);
  nor (G3426,G3370,G755);
  nor (G3430,G3373,G803);
  nor (G3434,G3376,G851);
  nor (G3438,G3379,G899);
  nor (G3442,G3382,G947);
  nor (G3446,G3334,G3385);
  nor (G3447,G3385,G995);
  nor (G3448,G3232,G3385);
  nor (G3451,G3389,G3390);
  nor (G3454,G3394,G3391);
  nor (G3458,G3346,G3397);
  nor (G3459,G3397,G3343);
  nor (G3460,G3401,G3402);
  nor (G3463,G3403,G1190);
  nor (G3467,G3355,G3406);
  nor (G3468,G3406,G1238);
  nor (G3469,G3253,G3406);
  nor (G3472,G3358,G3410);
  nor (G3473,G3410,G563);
  nor (G3474,G3257,G3410);
  nor (G3477,G3361,G3414);
  nor (G3478,G3414,G611);
  nor (G3479,G3261,G3414);
  nor (G3482,G3364,G3418);
  nor (G3483,G3418,G659);
  nor (G3484,G3265,G3418);
  nor (G3487,G3367,G3422);
  nor (G3488,G3422,G707);
  nor (G3489,G3269,G3422);
  nor (G3492,G3370,G3426);
  nor (G3493,G3426,G755);
  nor (G3494,G3273,G3426);
  nor (G3497,G3373,G3430);
  nor (G3498,G3430,G803);
  nor (G3499,G3277,G3430);
  nor (G3502,G3376,G3434);
  nor (G3503,G3434,G851);
  nor (G3504,G3281,G3434);
  nor (G3507,G3379,G3438);
  nor (G3508,G3438,G899);
  nor (G3509,G3285,G3438);
  nor (G3512,G3382,G3442);
  nor (G3513,G3442,G947);
  nor (G3514,G3289,G3442);
  nor (G3517,G3446,G3447);
  nor (G3520,G3451,G3448);
  nor (G3524,G3394,G3454);
  nor (G3525,G3454,G3391);
  nor (G3526,G3458,G3459);
  nor (G3529,G3460,G1142);
  nor (G3533,G3403,G3463);
  nor (G3534,G3463,G1190);
  nor (G3535,G3310,G3463);
  nor (G3538,G3467,G3468);
  nor (G3541,G1286,G3469);
  nor (G3545,G3477,G3478);
  nor (G3548,G3482,G3483);
  nor (G3551,G3487,G3488);
  nor (G3554,G3492,G3493);
  nor (G3557,G3497,G3498);
  nor (G3560,G3502,G3503);
  nor (G3563,G3507,G3508);
  nor (G3566,G3512,G3513);
  nor (G3569,G3517,G3514);
  nor (G3573,G3451,G3520);
  nor (G3574,G3520,G3448);
  nor (G3575,G3524,G3525);
  nor (G3578,G3526,G1094);
  nor (G3582,G3460,G3529);
  nor (G3583,G3529,G1142);
  nor (G3584,G3349,G3529);
  nor (G3587,G3533,G3534);
  nor (G3590,G3538,G3535);
  nor (G3594,G1286,G3541);
  nor (G3595,G3541,G3469);
  nor (G3596,G3545,G3474);
  nor (G3600,G3548,G3479);
  nor (G3604,G3551,G3484);
  nor (G3608,G3554,G3489);
  nor (G3612,G3557,G3494);
  nor (G3616,G3560,G3499);
  nor (G3620,G3563,G3504);
  nor (G3624,G3566,G3509);
  nor (G3628,G3517,G3569);
  nor (G3629,G3569,G3514);
  nor (G3630,G3573,G3574);
  nor (G3633,G3575,G1046);
  nor (G3637,G3526,G3578);
  nor (G3638,G3578,G1094);
  nor (G3639,G3397,G3578);
  nor (G3642,G3582,G3583);
  nor (G3645,G3587,G3584);
  nor (G3649,G3538,G3590);
  nor (G3650,G3590,G3535);
  nor (G3651,G3594,G3595);
  nor (G3654,G3545,G3596);
  nor (G3655,G3596,G3474);
  nor (G3656,G3548,G3600);
  nor (G3657,G3600,G3479);
  nor (G3658,G3551,G3604);
  nor (G3659,G3604,G3484);
  nor (G3660,G3554,G3608);
  nor (G3661,G3608,G3489);
  nor (G3662,G3557,G3612);
  nor (G3663,G3612,G3494);
  nor (G3664,G3560,G3616);
  nor (G3665,G3616,G3499);
  nor (G3666,G3563,G3620);
  nor (G3667,G3620,G3504);
  nor (G3668,G3566,G3624);
  nor (G3669,G3624,G3509);
  nor (G3670,G3628,G3629);
  nor (G3673,G3630,G998);
  nor (G3677,G3575,G3633);
  nor (G3678,G3633,G1046);
  nor (G3679,G3454,G3633);
  nor (G3682,G3637,G3638);
  nor (G3685,G3642,G3639);
  nor (G3689,G3587,G3645);
  nor (G3690,G3645,G3584);
  nor (G3691,G3649,G3650);
  nor (G3694,G3651,G1241);
  nor (G3698,G3654,G3655);
  nor (G3701,G3656,G3657);
  nor (G3704,G3658,G3659);
  nor (G3707,G3660,G3661);
  nor (G3710,G3662,G3663);
  nor (G3713,G3664,G3665);
  nor (G3716,G3666,G3667);
  nor (G3719,G3668,G3669);
  nor (G3722,G3670,G950);
  nor (G3726,G3630,G3673);
  nor (G3727,G3673,G998);
  nor (G3728,G3520,G3673);
  nor (G3731,G3677,G3678);
  nor (G3734,G3682,G3679);
  nor (G3738,G3642,G3685);
  nor (G3739,G3685,G3639);
  nor (G3740,G3689,G3690);
  nor (G3743,G3691,G1193);
  nor (G3747,G3651,G3694);
  nor (G3748,G3694,G1241);
  nor (G3749,G3541,G3694);
  nor (G3752,G3698,G566);
  nor (G3756,G3701,G614);
  nor (G3760,G3704,G662);
  nor (G3764,G3707,G710);
  nor (G3768,G3710,G758);
  nor (G3772,G3713,G806);
  nor (G3776,G3716,G854);
  nor (G3780,G3719,G902);
  nor (G3784,G3670,G3722);
  nor (G3785,G3722,G950);
  nor (G3786,G3569,G3722);
  nor (G3789,G3726,G3727);
  nor (G3792,G3731,G3728);
  nor (G3796,G3682,G3734);
  nor (G3797,G3734,G3679);
  nor (G3798,G3738,G3739);
  nor (G3801,G3740,G1145);
  nor (G3805,G3691,G3743);
  nor (G3806,G3743,G1193);
  nor (G3807,G3590,G3743);
  nor (G3810,G3747,G3748);
  nor (G3813,G1289,G3749);
  nor (G3817,G3698,G3752);
  nor (G3818,G3752,G566);
  nor (G3819,G3596,G3752);
  nor (G3822,G3701,G3756);
  nor (G3823,G3756,G614);
  nor (G3824,G3600,G3756);
  nor (G3827,G3704,G3760);
  nor (G3828,G3760,G662);
  nor (G3829,G3604,G3760);
  nor (G3832,G3707,G3764);
  nor (G3833,G3764,G710);
  nor (G3834,G3608,G3764);
  nor (G3837,G3710,G3768);
  nor (G3838,G3768,G758);
  nor (G3839,G3612,G3768);
  nor (G3842,G3713,G3772);
  nor (G3843,G3772,G806);
  nor (G3844,G3616,G3772);
  nor (G3847,G3716,G3776);
  nor (G3848,G3776,G854);
  nor (G3849,G3620,G3776);
  nor (G3852,G3719,G3780);
  nor (G3853,G3780,G902);
  nor (G3854,G3624,G3780);
  nor (G3857,G3784,G3785);
  nor (G3860,G3789,G3786);
  nor (G3864,G3731,G3792);
  nor (G3865,G3792,G3728);
  nor (G3866,G3796,G3797);
  nor (G3869,G3798,G1097);
  nor (G3873,G3740,G3801);
  nor (G3874,G3801,G1145);
  nor (G3875,G3645,G3801);
  nor (G3878,G3805,G3806);
  nor (G3881,G3810,G3807);
  nor (G3885,G1289,G3813);
  nor (G3886,G3813,G3749);
  nor (G3887,G3822,G3823);
  nor (G3890,G3827,G3828);
  nor (G3893,G3832,G3833);
  nor (G3896,G3837,G3838);
  nor (G3899,G3842,G3843);
  nor (G3902,G3847,G3848);
  nor (G3905,G3852,G3853);
  nor (G3908,G3857,G3854);
  nor (G3912,G3789,G3860);
  nor (G3913,G3860,G3786);
  nor (G3914,G3864,G3865);
  nor (G3917,G3866,G1049);
  nor (G3921,G3798,G3869);
  nor (G3922,G3869,G1097);
  nor (G3923,G3685,G3869);
  nor (G3926,G3873,G3874);
  nor (G3929,G3878,G3875);
  nor (G3933,G3810,G3881);
  nor (G3934,G3881,G3807);
  nor (G3935,G3885,G3886);
  nor (G3938,G3887,G3819);
  nor (G3942,G3890,G3824);
  nor (G3946,G3893,G3829);
  nor (G3950,G3896,G3834);
  nor (G3954,G3899,G3839);
  nor (G3958,G3902,G3844);
  nor (G3962,G3905,G3849);
  nor (G3966,G3857,G3908);
  nor (G3967,G3908,G3854);
  nor (G3968,G3912,G3913);
  nor (G3971,G3914,G1001);
  nor (G3975,G3866,G3917);
  nor (G3976,G3917,G1049);
  nor (G3977,G3734,G3917);
  nor (G3980,G3921,G3922);
  nor (G3983,G3926,G3923);
  nor (G3987,G3878,G3929);
  nor (G3988,G3929,G3875);
  nor (G3989,G3933,G3934);
  nor (G3992,G3935,G1244);
  nor (G3996,G3887,G3938);
  nor (G3997,G3938,G3819);
  nor (G3998,G3890,G3942);
  nor (G3999,G3942,G3824);
  nor (G4000,G3893,G3946);
  nor (G4001,G3946,G3829);
  nor (G4002,G3896,G3950);
  nor (G4003,G3950,G3834);
  nor (G4004,G3899,G3954);
  nor (G4005,G3954,G3839);
  nor (G4006,G3902,G3958);
  nor (G4007,G3958,G3844);
  nor (G4008,G3905,G3962);
  nor (G4009,G3962,G3849);
  nor (G4010,G3966,G3967);
  nor (G4013,G3968,G953);
  nor (G4017,G3914,G3971);
  nor (G4018,G3971,G1001);
  nor (G4019,G3792,G3971);
  nor (G4022,G3975,G3976);
  nor (G4025,G3980,G3977);
  nor (G4029,G3926,G3983);
  nor (G4030,G3983,G3923);
  nor (G4031,G3987,G3988);
  nor (G4034,G3989,G1196);
  nor (G4038,G3935,G3992);
  nor (G4039,G3992,G1244);
  nor (G4040,G3813,G3992);
  nor (G4043,G3996,G3997);
  nor (G4046,G3998,G3999);
  nor (G4049,G4000,G4001);
  nor (G4052,G4002,G4003);
  nor (G4055,G4004,G4005);
  nor (G4058,G4006,G4007);
  nor (G4061,G4008,G4009);
  nor (G4064,G4010,G905);
  nor (G4068,G3968,G4013);
  nor (G4069,G4013,G953);
  nor (G4070,G3860,G4013);
  nor (G4073,G4017,G4018);
  nor (G4076,G4022,G4019);
  nor (G4080,G3980,G4025);
  nor (G4081,G4025,G3977);
  nor (G4082,G4029,G4030);
  nor (G4085,G4031,G1148);
  nor (G4089,G3989,G4034);
  nor (G4090,G4034,G1196);
  nor (G4091,G3881,G4034);
  nor (G4094,G4038,G4039);
  nor (G4097,G1292,G4040);
  nor (G4101,G4043,G569);
  nor (G4105,G4046,G617);
  nor (G4109,G4049,G665);
  nor (G4113,G4052,G713);
  nor (G4117,G4055,G761);
  nor (G4121,G4058,G809);
  nor (G4125,G4061,G857);
  nor (G4129,G4010,G4064);
  nor (G4130,G4064,G905);
  nor (G4131,G3908,G4064);
  nor (G4134,G4068,G4069);
  nor (G4137,G4073,G4070);
  nor (G4141,G4022,G4076);
  nor (G4142,G4076,G4019);
  nor (G4143,G4080,G4081);
  nor (G4146,G4082,G1100);
  nor (G4150,G4031,G4085);
  nor (G4151,G4085,G1148);
  nor (G4152,G3929,G4085);
  nor (G4155,G4089,G4090);
  nor (G4158,G4094,G4091);
  nor (G4162,G1292,G4097);
  nor (G4163,G4097,G4040);
  nor (G4164,G4043,G4101);
  nor (G4165,G4101,G569);
  nor (G4166,G3938,G4101);
  nor (G4169,G4046,G4105);
  nor (G4170,G4105,G617);
  nor (G4171,G3942,G4105);
  nor (G4174,G4049,G4109);
  nor (G4175,G4109,G665);
  nor (G4176,G3946,G4109);
  nor (G4179,G4052,G4113);
  nor (G4180,G4113,G713);
  nor (G4181,G3950,G4113);
  nor (G4184,G4055,G4117);
  nor (G4185,G4117,G761);
  nor (G4186,G3954,G4117);
  nor (G4189,G4058,G4121);
  nor (G4190,G4121,G809);
  nor (G4191,G3958,G4121);
  nor (G4194,G4061,G4125);
  nor (G4195,G4125,G857);
  nor (G4196,G3962,G4125);
  nor (G4199,G4129,G4130);
  nor (G4202,G4134,G4131);
  nor (G4206,G4073,G4137);
  nor (G4207,G4137,G4070);
  nor (G4208,G4141,G4142);
  nor (G4211,G4143,G1052);
  nor (G4215,G4082,G4146);
  nor (G4216,G4146,G1100);
  nor (G4217,G3983,G4146);
  nor (G4220,G4150,G4151);
  nor (G4223,G4155,G4152);
  nor (G4227,G4094,G4158);
  nor (G4228,G4158,G4091);
  nor (G4229,G4162,G4163);
  nor (G4232,G4169,G4170);
  nor (G4235,G4174,G4175);
  nor (G4238,G4179,G4180);
  nor (G4241,G4184,G4185);
  nor (G4244,G4189,G4190);
  nor (G4247,G4194,G4195);
  nor (G4250,G4199,G4196);
  nor (G4254,G4134,G4202);
  nor (G4255,G4202,G4131);
  nor (G4256,G4206,G4207);
  nor (G4259,G4208,G1004);
  nor (G4263,G4143,G4211);
  nor (G4264,G4211,G1052);
  nor (G4265,G4025,G4211);
  nor (G4268,G4215,G4216);
  nor (G4271,G4220,G4217);
  nor (G4275,G4155,G4223);
  nor (G4276,G4223,G4152);
  nor (G4277,G4227,G4228);
  nor (G4280,G4229,G1247);
  nor (G4284,G4232,G4166);
  nor (G4288,G4235,G4171);
  nor (G4292,G4238,G4176);
  nor (G4296,G4241,G4181);
  nor (G4300,G4244,G4186);
  nor (G4304,G4247,G4191);
  nor (G4308,G4199,G4250);
  nor (G4309,G4250,G4196);
  nor (G4310,G4254,G4255);
  nor (G4313,G4256,G956);
  nor (G4317,G4208,G4259);
  nor (G4318,G4259,G1004);
  nor (G4319,G4076,G4259);
  nor (G4322,G4263,G4264);
  nor (G4325,G4268,G4265);
  nor (G4329,G4220,G4271);
  nor (G4330,G4271,G4217);
  nor (G4331,G4275,G4276);
  nor (G4334,G4277,G1199);
  nor (G4338,G4229,G4280);
  nor (G4339,G4280,G1247);
  nor (G4340,G4097,G4280);
  nor (G4343,G4232,G4284);
  nor (G4344,G4284,G4166);
  nor (G4345,G4235,G4288);
  nor (G4346,G4288,G4171);
  nor (G4347,G4238,G4292);
  nor (G4348,G4292,G4176);
  nor (G4349,G4241,G4296);
  nor (G4350,G4296,G4181);
  nor (G4351,G4244,G4300);
  nor (G4352,G4300,G4186);
  nor (G4353,G4247,G4304);
  nor (G4354,G4304,G4191);
  nor (G4355,G4308,G4309);
  nor (G4358,G4310,G908);
  nor (G4362,G4256,G4313);
  nor (G4363,G4313,G956);
  nor (G4364,G4137,G4313);
  nor (G4367,G4317,G4318);
  nor (G4370,G4322,G4319);
  nor (G4374,G4268,G4325);
  nor (G4375,G4325,G4265);
  nor (G4376,G4329,G4330);
  nor (G4379,G4331,G1151);
  nor (G4383,G4277,G4334);
  nor (G4384,G4334,G1199);
  nor (G4385,G4158,G4334);
  nor (G4388,G4338,G4339);
  nor (G4391,G1295,G4340);
  nor (G4395,G4343,G4344);
  nor (G4398,G4345,G4346);
  nor (G4401,G4347,G4348);
  nor (G4404,G4349,G4350);
  nor (G4407,G4351,G4352);
  nor (G4410,G4353,G4354);
  nor (G4413,G4355,G860);
  nor (G4417,G4310,G4358);
  nor (G4418,G4358,G908);
  nor (G4419,G4202,G4358);
  nor (G4422,G4362,G4363);
  nor (G4425,G4367,G4364);
  nor (G4429,G4322,G4370);
  nor (G4430,G4370,G4319);
  nor (G4431,G4374,G4375);
  nor (G4434,G4376,G1103);
  nor (G4438,G4331,G4379);
  nor (G4439,G4379,G1151);
  nor (G4440,G4223,G4379);
  nor (G4443,G4383,G4384);
  nor (G4446,G4388,G4385);
  nor (G4450,G1295,G4391);
  nor (G4451,G4391,G4340);
  nor (G4452,G4395,G572);
  nor (G4456,G4398,G620);
  nor (G4460,G4401,G668);
  nor (G4464,G4404,G716);
  nor (G4468,G4407,G764);
  nor (G4472,G4410,G812);
  nor (G4476,G4355,G4413);
  nor (G4477,G4413,G860);
  nor (G4478,G4250,G4413);
  nor (G4481,G4417,G4418);
  nor (G4484,G4422,G4419);
  nor (G4488,G4367,G4425);
  nor (G4489,G4425,G4364);
  nor (G4490,G4429,G4430);
  nor (G4493,G4431,G1055);
  nor (G4497,G4376,G4434);
  nor (G4498,G4434,G1103);
  nor (G4499,G4271,G4434);
  nor (G4502,G4438,G4439);
  nor (G4505,G4443,G4440);
  nor (G4509,G4388,G4446);
  nor (G4510,G4446,G4385);
  nor (G4511,G4450,G4451);
  nor (G4514,G4395,G4452);
  nor (G4515,G4452,G572);
  nor (G4516,G4284,G4452);
  nor (G4519,G4398,G4456);
  nor (G4520,G4456,G620);
  nor (G4521,G4288,G4456);
  nor (G4524,G4401,G4460);
  nor (G4525,G4460,G668);
  nor (G4526,G4292,G4460);
  nor (G4529,G4404,G4464);
  nor (G4530,G4464,G716);
  nor (G4531,G4296,G4464);
  nor (G4534,G4407,G4468);
  nor (G4535,G4468,G764);
  nor (G4536,G4300,G4468);
  nor (G4539,G4410,G4472);
  nor (G4540,G4472,G812);
  nor (G4541,G4304,G4472);
  nor (G4544,G4476,G4477);
  nor (G4547,G4481,G4478);
  nor (G4551,G4422,G4484);
  nor (G4552,G4484,G4419);
  nor (G4553,G4488,G4489);
  nor (G4556,G4490,G1007);
  nor (G4560,G4431,G4493);
  nor (G4561,G4493,G1055);
  nor (G4562,G4325,G4493);
  nor (G4565,G4497,G4498);
  nor (G4568,G4502,G4499);
  nor (G4572,G4443,G4505);
  nor (G4573,G4505,G4440);
  nor (G4574,G4509,G4510);
  nor (G4577,G4511,G1250);
  nor (G4581,G4519,G4520);
  nor (G4584,G4524,G4525);
  nor (G4587,G4529,G4530);
  nor (G4590,G4534,G4535);
  nor (G4593,G4539,G4540);
  nor (G4596,G4544,G4541);
  nor (G4600,G4481,G4547);
  nor (G4601,G4547,G4478);
  nor (G4602,G4551,G4552);
  nor (G4605,G4553,G959);
  nor (G4609,G4490,G4556);
  nor (G4610,G4556,G1007);
  nor (G4611,G4370,G4556);
  nor (G4614,G4560,G4561);
  nor (G4617,G4565,G4562);
  nor (G4621,G4502,G4568);
  nor (G4622,G4568,G4499);
  nor (G4623,G4572,G4573);
  nor (G4626,G4574,G1202);
  nor (G4630,G4511,G4577);
  nor (G4631,G4577,G1250);
  nor (G4632,G4391,G4577);
  nor (G4635,G4581,G4516);
  nor (G4639,G4584,G4521);
  nor (G4643,G4587,G4526);
  nor (G4647,G4590,G4531);
  nor (G4651,G4593,G4536);
  nor (G4655,G4544,G4596);
  nor (G4656,G4596,G4541);
  nor (G4657,G4600,G4601);
  nor (G4660,G4602,G911);
  nor (G4664,G4553,G4605);
  nor (G4665,G4605,G959);
  nor (G4666,G4425,G4605);
  nor (G4669,G4609,G4610);
  nor (G4672,G4614,G4611);
  nor (G4676,G4565,G4617);
  nor (G4677,G4617,G4562);
  nor (G4678,G4621,G4622);
  nor (G4681,G4623,G1154);
  nor (G4685,G4574,G4626);
  nor (G4686,G4626,G1202);
  nor (G4687,G4446,G4626);
  nor (G4690,G4630,G4631);
  nor (G4693,G1298,G4632);
  nor (G4697,G4581,G4635);
  nor (G4698,G4635,G4516);
  nor (G4699,G4584,G4639);
  nor (G4700,G4639,G4521);
  nor (G4701,G4587,G4643);
  nor (G4702,G4643,G4526);
  nor (G4703,G4590,G4647);
  nor (G4704,G4647,G4531);
  nor (G4705,G4593,G4651);
  nor (G4706,G4651,G4536);
  nor (G4707,G4655,G4656);
  nor (G4710,G4657,G863);
  nor (G4714,G4602,G4660);
  nor (G4715,G4660,G911);
  nor (G4716,G4484,G4660);
  nor (G4719,G4664,G4665);
  nor (G4722,G4669,G4666);
  nor (G4726,G4614,G4672);
  nor (G4727,G4672,G4611);
  nor (G4728,G4676,G4677);
  nor (G4731,G4678,G1106);
  nor (G4735,G4623,G4681);
  nor (G4736,G4681,G1154);
  nor (G4737,G4505,G4681);
  nor (G4740,G4685,G4686);
  nor (G4743,G4690,G4687);
  nor (G4747,G1298,G4693);
  nor (G4748,G4693,G4632);
  nor (G4749,G4697,G4698);
  nor (G4752,G4699,G4700);
  nor (G4755,G4701,G4702);
  nor (G4758,G4703,G4704);
  nor (G4761,G4705,G4706);
  nor (G4764,G4707,G815);
  nor (G4768,G4657,G4710);
  nor (G4769,G4710,G863);
  nor (G4770,G4547,G4710);
  nor (G4773,G4714,G4715);
  nor (G4776,G4719,G4716);
  nor (G4780,G4669,G4722);
  nor (G4781,G4722,G4666);
  nor (G4782,G4726,G4727);
  nor (G4785,G4728,G1058);
  nor (G4789,G4678,G4731);
  nor (G4790,G4731,G1106);
  nor (G4791,G4568,G4731);
  nor (G4794,G4735,G4736);
  nor (G4797,G4740,G4737);
  nor (G4801,G4690,G4743);
  nor (G4802,G4743,G4687);
  nor (G4803,G4747,G4748);
  nor (G4806,G4749,G575);
  nor (G4810,G4752,G623);
  nor (G4814,G4755,G671);
  nor (G4818,G4758,G719);
  nor (G4822,G4761,G767);
  nor (G4826,G4707,G4764);
  nor (G4827,G4764,G815);
  nor (G4828,G4596,G4764);
  nor (G4831,G4768,G4769);
  nor (G4834,G4773,G4770);
  nor (G4838,G4719,G4776);
  nor (G4839,G4776,G4716);
  nor (G4840,G4780,G4781);
  nor (G4843,G4782,G1010);
  nor (G4847,G4728,G4785);
  nor (G4848,G4785,G1058);
  nor (G4849,G4617,G4785);
  nor (G4852,G4789,G4790);
  nor (G4855,G4794,G4791);
  nor (G4859,G4740,G4797);
  nor (G4860,G4797,G4737);
  nor (G4861,G4801,G4802);
  nor (G4864,G4803,G1253);
  nor (G4868,G4749,G4806);
  nor (G4869,G4806,G575);
  nor (G4870,G4635,G4806);
  nor (G4873,G4752,G4810);
  nor (G4874,G4810,G623);
  nor (G4875,G4639,G4810);
  nor (G4878,G4755,G4814);
  nor (G4879,G4814,G671);
  nor (G4880,G4643,G4814);
  nor (G4883,G4758,G4818);
  nor (G4884,G4818,G719);
  nor (G4885,G4647,G4818);
  nor (G4888,G4761,G4822);
  nor (G4889,G4822,G767);
  nor (G4890,G4651,G4822);
  nor (G4893,G4826,G4827);
  nor (G4896,G4831,G4828);
  nor (G4900,G4773,G4834);
  nor (G4901,G4834,G4770);
  nor (G4902,G4838,G4839);
  nor (G4905,G4840,G962);
  nor (G4909,G4782,G4843);
  nor (G4910,G4843,G1010);
  nor (G4911,G4672,G4843);
  nor (G4914,G4847,G4848);
  nor (G4917,G4852,G4849);
  nor (G4921,G4794,G4855);
  nor (G4922,G4855,G4791);
  nor (G4923,G4859,G4860);
  nor (G4926,G4861,G1205);
  nor (G4930,G4803,G4864);
  nor (G4931,G4864,G1253);
  nor (G4932,G4693,G4864);
  nor (G4935,G4873,G4874);
  nor (G4938,G4878,G4879);
  nor (G4941,G4883,G4884);
  nor (G4944,G4888,G4889);
  nor (G4947,G4893,G4890);
  nor (G4951,G4831,G4896);
  nor (G4952,G4896,G4828);
  nor (G4953,G4900,G4901);
  nor (G4956,G4902,G914);
  nor (G4960,G4840,G4905);
  nor (G4961,G4905,G962);
  nor (G4962,G4722,G4905);
  nor (G4965,G4909,G4910);
  nor (G4968,G4914,G4911);
  nor (G4972,G4852,G4917);
  nor (G4973,G4917,G4849);
  nor (G4974,G4921,G4922);
  nor (G4977,G4923,G1157);
  nor (G4981,G4861,G4926);
  nor (G4982,G4926,G1205);
  nor (G4983,G4743,G4926);
  nor (G4986,G4930,G4931);
  nor (G4989,G1301,G4932);
  nor (G4993,G4935,G4870);
  nor (G4997,G4938,G4875);
  nor (G5001,G4941,G4880);
  nor (G5005,G4944,G4885);
  nor (G5009,G4893,G4947);
  nor (G5010,G4947,G4890);
  nor (G5011,G4951,G4952);
  nor (G5014,G4953,G866);
  nor (G5018,G4902,G4956);
  nor (G5019,G4956,G914);
  nor (G5020,G4776,G4956);
  nor (G5023,G4960,G4961);
  nor (G5026,G4965,G4962);
  nor (G5030,G4914,G4968);
  nor (G5031,G4968,G4911);
  nor (G5032,G4972,G4973);
  nor (G5035,G4974,G1109);
  nor (G5039,G4923,G4977);
  nor (G5040,G4977,G1157);
  nor (G5041,G4797,G4977);
  nor (G5044,G4981,G4982);
  nor (G5047,G4986,G4983);
  nor (G5051,G1301,G4989);
  nor (G5052,G4989,G4932);
  nor (G5053,G4935,G4993);
  nor (G5054,G4993,G4870);
  nor (G5055,G4938,G4997);
  nor (G5056,G4997,G4875);
  nor (G5057,G4941,G5001);
  nor (G5058,G5001,G4880);
  nor (G5059,G4944,G5005);
  nor (G5060,G5005,G4885);
  nor (G5061,G5009,G5010);
  nor (G5064,G5011,G818);
  nor (G5068,G4953,G5014);
  nor (G5069,G5014,G866);
  nor (G5070,G4834,G5014);
  nor (G5073,G5018,G5019);
  nor (G5076,G5023,G5020);
  nor (G5080,G4965,G5026);
  nor (G5081,G5026,G4962);
  nor (G5082,G5030,G5031);
  nor (G5085,G5032,G1061);
  nor (G5089,G4974,G5035);
  nor (G5090,G5035,G1109);
  nor (G5091,G4855,G5035);
  nor (G5094,G5039,G5040);
  nor (G5097,G5044,G5041);
  nor (G5101,G4986,G5047);
  nor (G5102,G5047,G4983);
  nor (G5103,G5051,G5052);
  nor (G5106,G5053,G5054);
  nor (G5109,G5055,G5056);
  nor (G5112,G5057,G5058);
  nor (G5115,G5059,G5060);
  nor (G5118,G5061,G770);
  nor (G5122,G5011,G5064);
  nor (G5123,G5064,G818);
  nor (G5124,G4896,G5064);
  nor (G5127,G5068,G5069);
  nor (G5130,G5073,G5070);
  nor (G5134,G5023,G5076);
  nor (G5135,G5076,G5020);
  nor (G5136,G5080,G5081);
  nor (G5139,G5082,G1013);
  nor (G5143,G5032,G5085);
  nor (G5144,G5085,G1061);
  nor (G5145,G4917,G5085);
  nor (G5148,G5089,G5090);
  nor (G5151,G5094,G5091);
  nor (G5155,G5044,G5097);
  nor (G5156,G5097,G5041);
  nor (G5157,G5101,G5102);
  nor (G5160,G5103,G1256);
  nor (G5164,G5106,G578);
  nor (G5168,G5109,G626);
  nor (G5172,G5112,G674);
  nor (G5176,G5115,G722);
  nor (G5180,G5061,G5118);
  nor (G5181,G5118,G770);
  nor (G5182,G4947,G5118);
  nor (G5185,G5122,G5123);
  nor (G5188,G5127,G5124);
  nor (G5192,G5073,G5130);
  nor (G5193,G5130,G5070);
  nor (G5194,G5134,G5135);
  nor (G5197,G5136,G965);
  nor (G5201,G5082,G5139);
  nor (G5202,G5139,G1013);
  nor (G5203,G4968,G5139);
  nor (G5206,G5143,G5144);
  nor (G5209,G5148,G5145);
  nor (G5213,G5094,G5151);
  nor (G5214,G5151,G5091);
  nor (G5215,G5155,G5156);
  nor (G5218,G5157,G1208);
  nor (G5222,G5103,G5160);
  nor (G5223,G5160,G1256);
  nor (G5224,G4989,G5160);
  nor (G5227,G5106,G5164);
  nor (G5228,G5164,G578);
  nor (G5229,G4993,G5164);
  nor (G5232,G5109,G5168);
  nor (G5233,G5168,G626);
  nor (G5234,G4997,G5168);
  nor (G5237,G5112,G5172);
  nor (G5238,G5172,G674);
  nor (G5239,G5001,G5172);
  nor (G5242,G5115,G5176);
  nor (G5243,G5176,G722);
  nor (G5244,G5005,G5176);
  nor (G5247,G5180,G5181);
  nor (G5250,G5185,G5182);
  nor (G5254,G5127,G5188);
  nor (G5255,G5188,G5124);
  nor (G5256,G5192,G5193);
  nor (G5259,G5194,G917);
  nor (G5263,G5136,G5197);
  nor (G5264,G5197,G965);
  nor (G5265,G5026,G5197);
  nor (G5268,G5201,G5202);
  nor (G5271,G5206,G5203);
  nor (G5275,G5148,G5209);
  nor (G5276,G5209,G5145);
  nor (G5277,G5213,G5214);
  nor (G5280,G5215,G1160);
  nor (G5284,G5157,G5218);
  nor (G5285,G5218,G1208);
  nor (G5286,G5047,G5218);
  nor (G5289,G5222,G5223);
  nor (G5292,G1304,G5224);
  nor (G5296,G5232,G5233);
  nor (G5299,G5237,G5238);
  nor (G5302,G5242,G5243);
  nor (G5305,G5247,G5244);
  nor (G5309,G5185,G5250);
  nor (G5310,G5250,G5182);
  nor (G5311,G5254,G5255);
  nor (G5314,G5256,G869);
  nor (G5318,G5194,G5259);
  nor (G5319,G5259,G917);
  nor (G5320,G5076,G5259);
  nor (G5323,G5263,G5264);
  nor (G5326,G5268,G5265);
  nor (G5330,G5206,G5271);
  nor (G5331,G5271,G5203);
  nor (G5332,G5275,G5276);
  nor (G5335,G5277,G1112);
  nor (G5339,G5215,G5280);
  nor (G5340,G5280,G1160);
  nor (G5341,G5097,G5280);
  nor (G5344,G5284,G5285);
  nor (G5347,G5289,G5286);
  nor (G5351,G1304,G5292);
  nor (G5352,G5292,G5224);
  nor (G5353,G5296,G5229);
  nor (G5357,G5299,G5234);
  nor (G5361,G5302,G5239);
  nor (G5365,G5247,G5305);
  nor (G5366,G5305,G5244);
  nor (G5367,G5309,G5310);
  nor (G5370,G5311,G821);
  nor (G5374,G5256,G5314);
  nor (G5375,G5314,G869);
  nor (G5376,G5130,G5314);
  nor (G5379,G5318,G5319);
  nor (G5382,G5323,G5320);
  nor (G5386,G5268,G5326);
  nor (G5387,G5326,G5265);
  nor (G5388,G5330,G5331);
  nor (G5391,G5332,G1064);
  nor (G5395,G5277,G5335);
  nor (G5396,G5335,G1112);
  nor (G5397,G5151,G5335);
  nor (G5400,G5339,G5340);
  nor (G5403,G5344,G5341);
  nor (G5407,G5289,G5347);
  nor (G5408,G5347,G5286);
  nor (G5409,G5351,G5352);
  nor (G5412,G5296,G5353);
  nor (G5413,G5353,G5229);
  nor (G5414,G5299,G5357);
  nor (G5415,G5357,G5234);
  nor (G5416,G5302,G5361);
  nor (G5417,G5361,G5239);
  nor (G5418,G5365,G5366);
  nor (G5421,G5367,G773);
  nor (G5425,G5311,G5370);
  nor (G5426,G5370,G821);
  nor (G5427,G5188,G5370);
  nor (G5430,G5374,G5375);
  nor (G5433,G5379,G5376);
  nor (G5437,G5323,G5382);
  nor (G5438,G5382,G5320);
  nor (G5439,G5386,G5387);
  nor (G5442,G5388,G1016);
  nor (G5446,G5332,G5391);
  nor (G5447,G5391,G1064);
  nor (G5448,G5209,G5391);
  nor (G5451,G5395,G5396);
  nor (G5454,G5400,G5397);
  nor (G5458,G5344,G5403);
  nor (G5459,G5403,G5341);
  nor (G5460,G5407,G5408);
  nor (G5463,G5409,G1259);
  nor (G5467,G5412,G5413);
  nor (G5470,G5414,G5415);
  nor (G5473,G5416,G5417);
  nor (G5476,G5418,G725);
  nor (G5480,G5367,G5421);
  nor (G5481,G5421,G773);
  nor (G5482,G5250,G5421);
  nor (G5485,G5425,G5426);
  nor (G5488,G5430,G5427);
  nor (G5492,G5379,G5433);
  nor (G5493,G5433,G5376);
  nor (G5494,G5437,G5438);
  nor (G5497,G5439,G968);
  nor (G5501,G5388,G5442);
  nor (G5502,G5442,G1016);
  nor (G5503,G5271,G5442);
  nor (G5506,G5446,G5447);
  nor (G5509,G5451,G5448);
  nor (G5513,G5400,G5454);
  nor (G5514,G5454,G5397);
  nor (G5515,G5458,G5459);
  nor (G5518,G5460,G1211);
  nor (G5522,G5409,G5463);
  nor (G5523,G5463,G1259);
  nor (G5524,G5292,G5463);
  nor (G5527,G5467,G581);
  nor (G5531,G5470,G629);
  nor (G5535,G5473,G677);
  nor (G5539,G5418,G5476);
  nor (G5540,G5476,G725);
  nor (G5541,G5305,G5476);
  nor (G5544,G5480,G5481);
  nor (G5547,G5485,G5482);
  nor (G5551,G5430,G5488);
  nor (G5552,G5488,G5427);
  nor (G5553,G5492,G5493);
  nor (G5556,G5494,G920);
  nor (G5560,G5439,G5497);
  nor (G5561,G5497,G968);
  nor (G5562,G5326,G5497);
  nor (G5565,G5501,G5502);
  nor (G5568,G5506,G5503);
  nor (G5572,G5451,G5509);
  nor (G5573,G5509,G5448);
  nor (G5574,G5513,G5514);
  nor (G5577,G5515,G1163);
  nor (G5581,G5460,G5518);
  nor (G5582,G5518,G1211);
  nor (G5583,G5347,G5518);
  nor (G5586,G5522,G5523);
  nor (G5589,G1307,G5524);
  nor (G5593,G5467,G5527);
  nor (G5594,G5527,G581);
  nor (G5595,G5353,G5527);
  nor (G5598,G5470,G5531);
  nor (G5599,G5531,G629);
  nor (G5600,G5357,G5531);
  nor (G5603,G5473,G5535);
  nor (G5604,G5535,G677);
  nor (G5605,G5361,G5535);
  nor (G5608,G5539,G5540);
  nor (G5611,G5544,G5541);
  nor (G5615,G5485,G5547);
  nor (G5616,G5547,G5482);
  nor (G5617,G5551,G5552);
  nor (G5620,G5553,G872);
  nor (G5624,G5494,G5556);
  nor (G5625,G5556,G920);
  nor (G5626,G5382,G5556);
  nor (G5629,G5560,G5561);
  nor (G5632,G5565,G5562);
  nor (G5636,G5506,G5568);
  nor (G5637,G5568,G5503);
  nor (G5638,G5572,G5573);
  nor (G5641,G5574,G1115);
  nor (G5645,G5515,G5577);
  nor (G5646,G5577,G1163);
  nor (G5647,G5403,G5577);
  nor (G5650,G5581,G5582);
  nor (G5653,G5586,G5583);
  nor (G5657,G1307,G5589);
  nor (G5658,G5589,G5524);
  nor (G5659,G5598,G5599);
  nor (G5662,G5603,G5604);
  nor (G5665,G5608,G5605);
  nor (G5669,G5544,G5611);
  nor (G5670,G5611,G5541);
  nor (G5671,G5615,G5616);
  nor (G5674,G5617,G824);
  nor (G5678,G5553,G5620);
  nor (G5679,G5620,G872);
  nor (G5680,G5433,G5620);
  nor (G5683,G5624,G5625);
  nor (G5686,G5629,G5626);
  nor (G5690,G5565,G5632);
  nor (G5691,G5632,G5562);
  nor (G5692,G5636,G5637);
  nor (G5695,G5638,G1067);
  nor (G5699,G5574,G5641);
  nor (G5700,G5641,G1115);
  nor (G5701,G5454,G5641);
  nor (G5704,G5645,G5646);
  nor (G5707,G5650,G5647);
  nor (G5711,G5586,G5653);
  nor (G5712,G5653,G5583);
  nor (G5713,G5657,G5658);
  nor (G5716,G5659,G5595);
  nor (G5720,G5662,G5600);
  nor (G5724,G5608,G5665);
  nor (G5725,G5665,G5605);
  nor (G5726,G5669,G5670);
  nor (G5729,G5671,G776);
  nor (G5733,G5617,G5674);
  nor (G5734,G5674,G824);
  nor (G5735,G5488,G5674);
  nor (G5738,G5678,G5679);
  nor (G5741,G5683,G5680);
  nor (G5745,G5629,G5686);
  nor (G5746,G5686,G5626);
  nor (G5747,G5690,G5691);
  nor (G5750,G5692,G1019);
  nor (G5754,G5638,G5695);
  nor (G5755,G5695,G1067);
  nor (G5756,G5509,G5695);
  nor (G5759,G5699,G5700);
  nor (G5762,G5704,G5701);
  nor (G5766,G5650,G5707);
  nor (G5767,G5707,G5647);
  nor (G5768,G5711,G5712);
  nor (G5771,G5659,G5716);
  nor (G5772,G5716,G5595);
  nor (G5773,G5662,G5720);
  nor (G5774,G5720,G5600);
  nor (G5775,G5724,G5725);
  nor (G5778,G5726,G728);
  nor (G5782,G5671,G5729);
  nor (G5783,G5729,G776);
  nor (G5784,G5547,G5729);
  nor (G5787,G5733,G5734);
  nor (G5790,G5738,G5735);
  nor (G5794,G5683,G5741);
  nor (G5795,G5741,G5680);
  nor (G5796,G5745,G5746);
  nor (G5799,G5747,G971);
  nor (G5803,G5692,G5750);
  nor (G5804,G5750,G1019);
  nor (G5805,G5568,G5750);
  nor (G5808,G5754,G5755);
  nor (G5811,G5759,G5756);
  nor (G5815,G5704,G5762);
  nor (G5816,G5762,G5701);
  nor (G5817,G5766,G5767);
  nor (G5820,G5771,G5772);
  nor (G5823,G5773,G5774);
  nor (G5826,G5775,G680);
  nor (G5830,G5726,G5778);
  nor (G5831,G5778,G728);
  nor (G5832,G5611,G5778);
  nor (G5835,G5782,G5783);
  nor (G5838,G5787,G5784);
  nor (G5842,G5738,G5790);
  nor (G5843,G5790,G5735);
  nor (G5844,G5794,G5795);
  nor (G5847,G5796,G923);
  nor (G5851,G5747,G5799);
  nor (G5852,G5799,G971);
  nor (G5853,G5632,G5799);
  nor (G5856,G5803,G5804);
  nor (G5859,G5808,G5805);
  nor (G5863,G5759,G5811);
  nor (G5864,G5811,G5756);
  nor (G5865,G5815,G5816);
  nor (G5868,G5820,G584);
  nor (G5872,G5823,G632);
  nor (G5876,G5775,G5826);
  nor (G5877,G5826,G680);
  nor (G5878,G5665,G5826);
  nor (G5881,G5830,G5831);
  nor (G5884,G5835,G5832);
  nor (G5888,G5787,G5838);
  nor (G5889,G5838,G5784);
  nor (G5890,G5842,G5843);
  nor (G5893,G5844,G875);
  nor (G5897,G5796,G5847);
  nor (G5898,G5847,G923);
  nor (G5899,G5686,G5847);
  nor (G5902,G5851,G5852);
  nor (G5905,G5856,G5853);
  nor (G5909,G5808,G5859);
  nor (G5910,G5859,G5805);
  nor (G5911,G5863,G5864);
  nor (G5914,G5820,G5868);
  nor (G5915,G5868,G584);
  nor (G5916,G5716,G5868);
  nor (G5919,G5823,G5872);
  nor (G5920,G5872,G632);
  nor (G5921,G5720,G5872);
  nor (G5924,G5876,G5877);
  nor (G5927,G5881,G5878);
  nor (G5931,G5835,G5884);
  nor (G5932,G5884,G5832);
  nor (G5933,G5888,G5889);
  nor (G5936,G5890,G827);
  nor (G5940,G5844,G5893);
  nor (G5941,G5893,G875);
  nor (G5942,G5741,G5893);
  nor (G5945,G5897,G5898);
  nor (G5948,G5902,G5899);
  nor (G5952,G5856,G5905);
  nor (G5953,G5905,G5853);
  nor (G5954,G5909,G5910);
  nor (G5957,G5919,G5920);
  nor (G5960,G5924,G5921);
  nor (G5964,G5881,G5927);
  nor (G5965,G5927,G5878);
  nor (G5966,G5931,G5932);
  nor (G5969,G5933,G779);
  nor (G5973,G5890,G5936);
  nor (G5974,G5936,G827);
  nor (G5975,G5790,G5936);
  nor (G5978,G5940,G5941);
  nor (G5981,G5945,G5942);
  nor (G5985,G5902,G5948);
  nor (G5986,G5948,G5899);
  nor (G5987,G5952,G5953);
  nor (G5990,G5957,G5916);
  nor (G5994,G5924,G5960);
  nor (G5995,G5960,G5921);
  nor (G5996,G5964,G5965);
  nor (G5999,G5966,G731);
  nor (G6003,G5933,G5969);
  nor (G6004,G5969,G779);
  nor (G6005,G5838,G5969);
  nor (G6008,G5973,G5974);
  nor (G6011,G5978,G5975);
  nor (G6015,G5945,G5981);
  nor (G6016,G5981,G5942);
  nor (G6017,G5985,G5986);
  nor (G6020,G5957,G5990);
  nor (G6021,G5990,G5916);
  nor (G6022,G5994,G5995);
  nor (G6025,G5996,G683);
  nor (G6029,G5966,G5999);
  nor (G6030,G5999,G731);
  nor (G6031,G5884,G5999);
  nor (G6034,G6003,G6004);
  nor (G6037,G6008,G6005);
  nor (G6041,G5978,G6011);
  nor (G6042,G6011,G5975);
  nor (G6043,G6015,G6016);
  nor (G6046,G6020,G6021);
  nor (G6049,G6022,G635);
  nor (G6053,G5996,G6025);
  nor (G6054,G6025,G683);
  nor (G6055,G5927,G6025);
  nor (G6058,G6029,G6030);
  nor (G6061,G6034,G6031);
  nor (G6065,G6008,G6037);
  nor (G6066,G6037,G6005);
  nor (G6067,G6041,G6042);
  nor (G6070,G6046,G587);
  nor (G6074,G6022,G6049);
  nor (G6075,G6049,G635);
  nor (G6076,G5960,G6049);
  nor (G6079,G6053,G6054);
  nor (G6082,G6058,G6055);
  nor (G6086,G6034,G6061);
  nor (G6087,G6061,G6031);
  nor (G6088,G6065,G6066);
  nor (G6091,G6046,G6070);
  nor (G6092,G6070,G587);
  nor (G6093,G5990,G6070);
  nor (G6096,G6074,G6075);
  nor (G6099,G6079,G6076);
  nor (G6103,G6058,G6082);
  nor (G6104,G6082,G6055);
  nor (G6105,G6086,G6087);
  nor (G6108,G6096,G6093);
  nor (G6112,G6079,G6099);
  nor (G6113,G6099,G6076);
  nor (G6114,G6103,G6104);
  nor (G6117,G6096,G6108);
  nor (G6118,G6108,G6093);
  nor (G6119,G6112,G6113);
  nor (G6122,G6117,G6118);
  not (G6125,G6122);
  nor (G6129,G6122,G6125);
  not (G6130,G6125);
  nor (G6131,G6108,G6125);
  nor (G6134,G6119,G6131);
  nor (G6138,G6119,G6134);
  nor (G6139,G6134,G6131);
  nor (G6140,G6099,G6134);
  nor (G6143,G6114,G6140);
  nor (G6147,G6114,G6143);
  nor (G6148,G6143,G6140);
  nor (G6149,G6082,G6143);
  nor (G6152,G6105,G6149);
  nor (G6156,G6105,G6152);
  nor (G6157,G6152,G6149);
  nor (G6158,G6061,G6152);
  nor (G6161,G6088,G6158);
  nor (G6165,G6088,G6161);
  nor (G6166,G6161,G6158);
  nor (G6167,G6037,G6161);
  nor (G6170,G6067,G6167);
  nor (G6174,G6067,G6170);
  nor (G6175,G6170,G6167);
  nor (G6176,G6011,G6170);
  nor (G6179,G6043,G6176);
  nor (G6183,G6043,G6179);
  nor (G6184,G6179,G6176);
  nor (G6185,G5981,G6179);
  nor (G6188,G6017,G6185);
  nor (G6192,G6017,G6188);
  nor (G6193,G6188,G6185);
  nor (G6194,G5948,G6188);
  nor (G6197,G5987,G6194);
  nor (G6201,G5987,G6197);
  nor (G6202,G6197,G6194);
  nor (G6203,G5905,G6197);
  nor (G6206,G5954,G6203);
  nor (G6210,G5954,G6206);
  nor (G6211,G6206,G6203);
  nor (G6212,G5859,G6206);
  nor (G6215,G5911,G6212);
  nor (G6219,G5911,G6215);
  nor (G6220,G6215,G6212);
  nor (G6221,G5811,G6215);
  nor (G6224,G5865,G6221);
  nor (G6228,G5865,G6224);
  nor (G6229,G6224,G6221);
  nor (G6230,G5762,G6224);
  nor (G6233,G5817,G6230);
  nor (G6237,G5817,G6233);
  nor (G6238,G6233,G6230);
  nor (G6239,G5707,G6233);
  nor (G6242,G5768,G6239);
  nor (G6246,G5768,G6242);
  nor (G6247,G6242,G6239);
  nor (G6248,G5653,G6242);
  nor (G6251,G5713,G6248);
  nor (G6255,G5713,G6251);
  nor (G6256,G6251,G6248);
  and (G6257,G1,G17);
  nor (G6258,G1505,G1506);
  nor (G6259,G1822,G1823);
  nor (G6260,G2146,G2147);
  nor (G6261,G2472,G2473);
  nor (G6262,G2801,G2802);
  nor (G6263,G3134,G3135);
  nor (G6264,G3472,G3473);
  nor (G6265,G3817,G3818);
  nor (G6266,G4164,G4165);
  nor (G6267,G4514,G4515);
  nor (G6268,G4868,G4869);
  nor (G6269,G5227,G5228);
  nor (G6270,G5593,G5594);
  nor (G6271,G5914,G5915);
  nor (G6272,G6091,G6092);
  nor (G6273,G6129,G6130);
  nor (G6274,G6138,G6139);
  nor (G6275,G6147,G6148);
  nor (G6276,G6156,G6157);
  nor (G6277,G6165,G6166);
  nor (G6278,G6174,G6175);
  nor (G6279,G6183,G6184);
  nor (G6280,G6192,G6193);
  nor (G6281,G6201,G6202);
  nor (G6282,G6210,G6211);
  nor (G6283,G6219,G6220);
  nor (G6284,G6228,G6229);
  nor (G6285,G6237,G6238);
  nor (G6286,G6246,G6247);
  nor (G6287,G5589,G6251);
  nor (G6288,G6255,G6256);

endmodule
