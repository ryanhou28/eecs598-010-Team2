module c1355(G1,G10,G11,G12,G13,G1324,G1325,G1326,G1327,G1328,G1329,G1330,
  G1331,G1332,G1333,G1334,G1335,G1336,G1337,G1338,G1339,G1340,G1341,G1342,
  G1343,G1344,G1345,G1346,G1347,G1348,G1349,G1350,G1351,G1352,G1353,G1354,
  G1355,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G3,
  G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G4,G40,G41,G5,G6,G7,G8,G9);
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
  G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,
  G40,G41;
output G1324,G1325,G1326,G1327,G1328,G1329,G1330,G1331,G1332,G1333,G1334,G1335,
  G1336,G1337,G1338,G1339,G1340,G1341,G1342,G1343,G1344,G1345,G1346,G1347,
  G1348,G1349,G1350,G1351,G1352,G1353,G1354,G1355;

  wire G242,G245,G248,G251,G254,G257,G260,G263,G266,G269,G272,G275,G278,G281,
    G284,G287,G290,G293,G296,G299,G302,G305,G308,G311,G314,G317,G320,G323,G326,
    G329,G332,G335,G338,G341,G344,G347,G350,G353,G356,G359,G362,G363,G364,G365,
    G366,G367,G368,G369,G370,G371,G372,G373,G374,G375,G376,G377,G378,G379,G380,
    G381,G382,G383,G384,G385,G386,G387,G388,G389,G390,G391,G392,G393,G394,G395,
    G396,G397,G398,G399,G400,G401,G402,G403,G404,G405,G406,G407,G408,G409,G410,
    G411,G412,G413,G414,G415,G416,G417,G418,G419,G420,G421,G422,G423,G424,G425,
    G426,G429,G432,G435,G438,G441,G444,G447,G450,G453,G456,G459,G462,G465,G468,
    G471,G474,G477,G480,G483,G486,G489,G492,G495,G498,G501,G504,G507,G510,G513,
    G516,G519,G522,G525,G528,G531,G534,G537,G540,G543,G546,G549,G552,G555,G558,
    G561,G564,G567,G570,G571,G572,G573,G574,G575,G576,G577,G578,G579,G580,G581,
    G582,G583,G584,G585,G586,G587,G588,G589,G590,G591,G592,G593,G594,G595,G596,
    G597,G598,G599,G600,G601,G602,G607,G612,G617,G622,G627,G632,G637,G642,G645,
    G648,G651,G654,G657,G660,G663,G666,G669,G672,G675,G678,G681,G684,G687,G690,
    G691,G692,G693,G694,G695,G696,G697,G698,G699,G700,G701,G702,G703,G704,G705,
    G706,G709,G712,G715,G718,G721,G724,G727,G730,G733,G736,G739,G742,G745,G748,
    G751,G754,G755,G756,G757,G758,G759,G760,G761,G762,G763,G764,G765,G766,G767,
    G768,G769,G770,G773,G776,G779,G782,G785,G788,G791,G794,G797,G800,G803,G806,
    G809,G812,G815,G818,G819,G820,G821,G822,G823,G824,G825,G826,G827,G828,G829,
    G830,G831,G832,G833,G834,G847,G860,G873,G886,G899,G912,G925,G938,G939,G940,
    G941,G942,G943,G944,G945,G946,G947,G948,G949,G950,G951,G952,G953,G954,G955,
    G956,G957,G958,G959,G960,G961,G962,G963,G964,G965,G966,G967,G968,G969,G970,
    G971,G972,G973,G974,G975,G976,G977,G978,G979,G980,G981,G982,G983,G984,G985,
    G986,G991,G996,G1001,G1006,G1011,G1016,G1021,G1026,G1031,G1036,G1039,G1042,
    G1045,G1048,G1051,G1054,G1057,G1060,G1063,G1066,G1069,G1072,G1075,G1078,
    G1081,G1084,G1087,G1090,G1093,G1096,G1099,G1102,G1105,G1108,G1111,G1114,
    G1117,G1120,G1123,G1126,G1129,G1132,G1135,G1138,G1141,G1144,G1147,G1150,
    G1153,G1156,G1159,G1162,G1165,G1168,G1171,G1174,G1177,G1180,G1183,G1186,
    G1189,G1192,G1195,G1198,G1201,G1204,G1207,G1210,G1213,G1216,G1219,G1222,
    G1225,G1228,G1229,G1230,G1231,G1232,G1233,G1234,G1235,G1236,G1237,G1238,
    G1239,G1240,G1241,G1242,G1243,G1244,G1245,G1246,G1247,G1248,G1249,G1250,
    G1251,G1252,G1253,G1254,G1255,G1256,G1257,G1258,G1259,G1260,G1261,G1262,
    G1263,G1264,G1265,G1266,G1267,G1268,G1269,G1270,G1271,G1272,G1273,G1274,
    G1275,G1276,G1277,G1278,G1279,G1280,G1281,G1282,G1283,G1284,G1285,G1286,
    G1287,G1288,G1289,G1290,G1291,G1292,G1293,G1294,G1295,G1296,G1297,G1298,
    G1299,G1300,G1301,G1302,G1303,G1304,G1305,G1306,G1307,G1308,G1309,G1310,
    G1311,G1312,G1313,G1314,G1315,G1316,G1317,G1318,G1319,G1320,G1321,G1322,
    G1323;

  and (G242,G33,G41);
  and (G245,G34,G41);
  and (G248,G35,G41);
  and (G251,G36,G41);
  and (G254,G37,G41);
  and (G257,G38,G41);
  and (G260,G39,G41);
  and (G263,G40,G41);
  nand (G266,G1,G2);
  nand (G269,G3,G4);
  nand (G272,G5,G6);
  nand (G275,G7,G8);
  nand (G278,G9,G10);
  nand (G281,G11,G12);
  nand (G284,G13,G14);
  nand (G287,G15,G16);
  nand (G290,G17,G18);
  nand (G293,G19,G20);
  nand (G296,G21,G22);
  nand (G299,G23,G24);
  nand (G302,G25,G26);
  nand (G305,G27,G28);
  nand (G308,G29,G30);
  nand (G311,G31,G32);
  nand (G314,G1,G5);
  nand (G317,G9,G13);
  nand (G320,G2,G6);
  nand (G323,G10,G14);
  nand (G326,G3,G7);
  nand (G329,G11,G15);
  nand (G332,G4,G8);
  nand (G335,G12,G16);
  nand (G338,G17,G21);
  nand (G341,G25,G29);
  nand (G344,G18,G22);
  nand (G347,G26,G30);
  nand (G350,G19,G23);
  nand (G353,G27,G31);
  nand (G356,G20,G24);
  nand (G359,G28,G32);
  nand (G362,G1,G266);
  nand (G363,G2,G266);
  nand (G364,G3,G269);
  nand (G365,G4,G269);
  nand (G366,G5,G272);
  nand (G367,G6,G272);
  nand (G368,G7,G275);
  nand (G369,G8,G275);
  nand (G370,G9,G278);
  nand (G371,G10,G278);
  nand (G372,G11,G281);
  nand (G373,G12,G281);
  nand (G374,G13,G284);
  nand (G375,G14,G284);
  nand (G376,G15,G287);
  nand (G377,G16,G287);
  nand (G378,G17,G290);
  nand (G379,G18,G290);
  nand (G380,G19,G293);
  nand (G381,G20,G293);
  nand (G382,G21,G296);
  nand (G383,G22,G296);
  nand (G384,G23,G299);
  nand (G385,G24,G299);
  nand (G386,G25,G302);
  nand (G387,G26,G302);
  nand (G388,G27,G305);
  nand (G389,G28,G305);
  nand (G390,G29,G308);
  nand (G391,G30,G308);
  nand (G392,G31,G311);
  nand (G393,G32,G311);
  nand (G394,G1,G314);
  nand (G395,G5,G314);
  nand (G396,G9,G317);
  nand (G397,G13,G317);
  nand (G398,G2,G320);
  nand (G399,G6,G320);
  nand (G400,G10,G323);
  nand (G401,G14,G323);
  nand (G402,G3,G326);
  nand (G403,G7,G326);
  nand (G404,G11,G329);
  nand (G405,G15,G329);
  nand (G406,G4,G332);
  nand (G407,G8,G332);
  nand (G408,G12,G335);
  nand (G409,G16,G335);
  nand (G410,G17,G338);
  nand (G411,G21,G338);
  nand (G412,G25,G341);
  nand (G413,G29,G341);
  nand (G414,G18,G344);
  nand (G415,G22,G344);
  nand (G416,G26,G347);
  nand (G417,G30,G347);
  nand (G418,G19,G350);
  nand (G419,G23,G350);
  nand (G420,G27,G353);
  nand (G421,G31,G353);
  nand (G422,G20,G356);
  nand (G423,G24,G356);
  nand (G424,G28,G359);
  nand (G425,G32,G359);
  nand (G426,G362,G363);
  nand (G429,G364,G365);
  nand (G432,G366,G367);
  nand (G435,G368,G369);
  nand (G438,G370,G371);
  nand (G441,G372,G373);
  nand (G444,G374,G375);
  nand (G447,G376,G377);
  nand (G450,G378,G379);
  nand (G453,G380,G381);
  nand (G456,G382,G383);
  nand (G459,G384,G385);
  nand (G462,G386,G387);
  nand (G465,G388,G389);
  nand (G468,G390,G391);
  nand (G471,G392,G393);
  nand (G474,G394,G395);
  nand (G477,G396,G397);
  nand (G480,G398,G399);
  nand (G483,G400,G401);
  nand (G486,G402,G403);
  nand (G489,G404,G405);
  nand (G492,G406,G407);
  nand (G495,G408,G409);
  nand (G498,G410,G411);
  nand (G501,G412,G413);
  nand (G504,G414,G415);
  nand (G507,G416,G417);
  nand (G510,G418,G419);
  nand (G513,G420,G421);
  nand (G516,G422,G423);
  nand (G519,G424,G425);
  nand (G522,G426,G429);
  nand (G525,G432,G435);
  nand (G528,G438,G441);
  nand (G531,G444,G447);
  nand (G534,G450,G453);
  nand (G537,G456,G459);
  nand (G540,G462,G465);
  nand (G543,G468,G471);
  nand (G546,G474,G477);
  nand (G549,G480,G483);
  nand (G552,G486,G489);
  nand (G555,G492,G495);
  nand (G558,G498,G501);
  nand (G561,G504,G507);
  nand (G564,G510,G513);
  nand (G567,G516,G519);
  nand (G570,G426,G522);
  nand (G571,G429,G522);
  nand (G572,G432,G525);
  nand (G573,G435,G525);
  nand (G574,G438,G528);
  nand (G575,G441,G528);
  nand (G576,G444,G531);
  nand (G577,G447,G531);
  nand (G578,G450,G534);
  nand (G579,G453,G534);
  nand (G580,G456,G537);
  nand (G581,G459,G537);
  nand (G582,G462,G540);
  nand (G583,G465,G540);
  nand (G584,G468,G543);
  nand (G585,G471,G543);
  nand (G586,G474,G546);
  nand (G587,G477,G546);
  nand (G588,G480,G549);
  nand (G589,G483,G549);
  nand (G590,G486,G552);
  nand (G591,G489,G552);
  nand (G592,G492,G555);
  nand (G593,G495,G555);
  nand (G594,G498,G558);
  nand (G595,G501,G558);
  nand (G596,G504,G561);
  nand (G597,G507,G561);
  nand (G598,G510,G564);
  nand (G599,G513,G564);
  nand (G600,G516,G567);
  nand (G601,G519,G567);
  nand (G602,G570,G571);
  nand (G607,G572,G573);
  nand (G612,G574,G575);
  nand (G617,G576,G577);
  nand (G622,G578,G579);
  nand (G627,G580,G581);
  nand (G632,G582,G583);
  nand (G637,G584,G585);
  nand (G642,G586,G587);
  nand (G645,G588,G589);
  nand (G648,G590,G591);
  nand (G651,G592,G593);
  nand (G654,G594,G595);
  nand (G657,G596,G597);
  nand (G660,G598,G599);
  nand (G663,G600,G601);
  nand (G666,G602,G607);
  nand (G669,G612,G617);
  nand (G672,G602,G612);
  nand (G675,G607,G617);
  nand (G678,G622,G627);
  nand (G681,G632,G637);
  nand (G684,G622,G632);
  nand (G687,G627,G637);
  nand (G690,G602,G666);
  nand (G691,G607,G666);
  nand (G692,G612,G669);
  nand (G693,G617,G669);
  nand (G694,G602,G672);
  nand (G695,G612,G672);
  nand (G696,G607,G675);
  nand (G697,G617,G675);
  nand (G698,G622,G678);
  nand (G699,G627,G678);
  nand (G700,G632,G681);
  nand (G701,G637,G681);
  nand (G702,G622,G684);
  nand (G703,G632,G684);
  nand (G704,G627,G687);
  nand (G705,G637,G687);
  nand (G706,G690,G691);
  nand (G709,G692,G693);
  nand (G712,G694,G695);
  nand (G715,G696,G697);
  nand (G718,G698,G699);
  nand (G721,G700,G701);
  nand (G724,G702,G703);
  nand (G727,G704,G705);
  nand (G730,G242,G718);
  nand (G733,G245,G721);
  nand (G736,G248,G724);
  nand (G739,G251,G727);
  nand (G742,G254,G706);
  nand (G745,G257,G709);
  nand (G748,G260,G712);
  nand (G751,G263,G715);
  nand (G754,G242,G730);
  nand (G755,G718,G730);
  nand (G756,G245,G733);
  nand (G757,G721,G733);
  nand (G758,G248,G736);
  nand (G759,G724,G736);
  nand (G760,G251,G739);
  nand (G761,G727,G739);
  nand (G762,G254,G742);
  nand (G763,G706,G742);
  nand (G764,G257,G745);
  nand (G765,G709,G745);
  nand (G766,G260,G748);
  nand (G767,G712,G748);
  nand (G768,G263,G751);
  nand (G769,G715,G751);
  nand (G770,G754,G755);
  nand (G773,G756,G757);
  nand (G776,G758,G759);
  nand (G779,G760,G761);
  nand (G782,G762,G763);
  nand (G785,G764,G765);
  nand (G788,G766,G767);
  nand (G791,G768,G769);
  nand (G794,G642,G770);
  nand (G797,G645,G773);
  nand (G800,G648,G776);
  nand (G803,G651,G779);
  nand (G806,G654,G782);
  nand (G809,G657,G785);
  nand (G812,G660,G788);
  nand (G815,G663,G791);
  nand (G818,G642,G794);
  nand (G819,G770,G794);
  nand (G820,G645,G797);
  nand (G821,G773,G797);
  nand (G822,G648,G800);
  nand (G823,G776,G800);
  nand (G824,G651,G803);
  nand (G825,G779,G803);
  nand (G826,G654,G806);
  nand (G827,G782,G806);
  nand (G828,G657,G809);
  nand (G829,G785,G809);
  nand (G830,G660,G812);
  nand (G831,G788,G812);
  nand (G832,G663,G815);
  nand (G833,G791,G815);
  nand (G834,G818,G819);
  nand (G847,G820,G821);
  nand (G860,G822,G823);
  nand (G873,G824,G825);
  nand (G886,G828,G829);
  nand (G899,G832,G833);
  nand (G912,G830,G831);
  nand (G925,G826,G827);
  not (G938,G834);
  not (G939,G847);
  not (G940,G860);
  not (G941,G834);
  not (G942,G847);
  not (G943,G873);
  not (G944,G834);
  not (G945,G860);
  not (G946,G873);
  not (G947,G847);
  not (G948,G860);
  not (G949,G873);
  not (G950,G886);
  not (G951,G899);
  not (G952,G886);
  not (G953,G912);
  not (G954,G925);
  not (G955,G899);
  not (G956,G925);
  not (G957,G912);
  not (G958,G925);
  not (G959,G886);
  not (G960,G912);
  not (G961,G925);
  not (G962,G886);
  not (G963,G899);
  not (G964,G925);
  not (G965,G912);
  not (G966,G899);
  not (G967,G886);
  not (G968,G912);
  not (G969,G899);
  not (G970,G847);
  not (G971,G873);
  not (G972,G847);
  not (G973,G860);
  not (G974,G834);
  not (G975,G873);
  not (G976,G834);
  not (G977,G860);
  and (G978,G938,G939,G940,G873);
  and (G979,G941,G942,G860,G943);
  and (G980,G944,G847,G945,G946);
  and (G981,G834,G947,G948,G949);
  and (G982,G958,G959,G960,G899);
  and (G983,G961,G962,G912,G963);
  and (G984,G964,G886,G965,G966);
  and (G985,G925,G967,G968,G969);
  or (G986,G978,G979,G980,G981);
  or (G991,G982,G983,G984,G985);
  and (G996,G925,G950,G912,G951,G986);
  and (G1001,G925,G952,G953,G899,G986);
  and (G1006,G954,G886,G912,G955,G986);
  and (G1011,G956,G886,G957,G899,G986);
  and (G1016,G834,G970,G860,G971,G991);
  and (G1021,G834,G972,G973,G873,G991);
  and (G1026,G974,G847,G860,G975,G991);
  and (G1031,G976,G847,G977,G873,G991);
  and (G1036,G834,G996);
  and (G1039,G847,G996);
  and (G1042,G860,G996);
  and (G1045,G873,G996);
  and (G1048,G834,G1001);
  and (G1051,G847,G1001);
  and (G1054,G860,G1001);
  and (G1057,G873,G1001);
  and (G1060,G834,G1006);
  and (G1063,G847,G1006);
  and (G1066,G860,G1006);
  and (G1069,G873,G1006);
  and (G1072,G834,G1011);
  and (G1075,G847,G1011);
  and (G1078,G860,G1011);
  and (G1081,G873,G1011);
  and (G1084,G925,G1016);
  and (G1087,G886,G1016);
  and (G1090,G912,G1016);
  and (G1093,G899,G1016);
  and (G1096,G925,G1021);
  and (G1099,G886,G1021);
  and (G1102,G912,G1021);
  and (G1105,G899,G1021);
  and (G1108,G925,G1026);
  and (G1111,G886,G1026);
  and (G1114,G912,G1026);
  and (G1117,G899,G1026);
  and (G1120,G925,G1031);
  and (G1123,G886,G1031);
  and (G1126,G912,G1031);
  and (G1129,G899,G1031);
  nand (G1132,G1,G1036);
  nand (G1135,G2,G1039);
  nand (G1138,G3,G1042);
  nand (G1141,G4,G1045);
  nand (G1144,G5,G1048);
  nand (G1147,G6,G1051);
  nand (G1150,G7,G1054);
  nand (G1153,G8,G1057);
  nand (G1156,G9,G1060);
  nand (G1159,G10,G1063);
  nand (G1162,G11,G1066);
  nand (G1165,G12,G1069);
  nand (G1168,G13,G1072);
  nand (G1171,G14,G1075);
  nand (G1174,G15,G1078);
  nand (G1177,G16,G1081);
  nand (G1180,G17,G1084);
  nand (G1183,G18,G1087);
  nand (G1186,G19,G1090);
  nand (G1189,G20,G1093);
  nand (G1192,G21,G1096);
  nand (G1195,G22,G1099);
  nand (G1198,G23,G1102);
  nand (G1201,G24,G1105);
  nand (G1204,G25,G1108);
  nand (G1207,G26,G1111);
  nand (G1210,G27,G1114);
  nand (G1213,G28,G1117);
  nand (G1216,G29,G1120);
  nand (G1219,G30,G1123);
  nand (G1222,G31,G1126);
  nand (G1225,G32,G1129);
  nand (G1228,G1,G1132);
  nand (G1229,G1036,G1132);
  nand (G1230,G2,G1135);
  nand (G1231,G1039,G1135);
  nand (G1232,G3,G1138);
  nand (G1233,G1042,G1138);
  nand (G1234,G4,G1141);
  nand (G1235,G1045,G1141);
  nand (G1236,G5,G1144);
  nand (G1237,G1048,G1144);
  nand (G1238,G6,G1147);
  nand (G1239,G1051,G1147);
  nand (G1240,G7,G1150);
  nand (G1241,G1054,G1150);
  nand (G1242,G8,G1153);
  nand (G1243,G1057,G1153);
  nand (G1244,G9,G1156);
  nand (G1245,G1060,G1156);
  nand (G1246,G10,G1159);
  nand (G1247,G1063,G1159);
  nand (G1248,G11,G1162);
  nand (G1249,G1066,G1162);
  nand (G1250,G12,G1165);
  nand (G1251,G1069,G1165);
  nand (G1252,G13,G1168);
  nand (G1253,G1072,G1168);
  nand (G1254,G14,G1171);
  nand (G1255,G1075,G1171);
  nand (G1256,G15,G1174);
  nand (G1257,G1078,G1174);
  nand (G1258,G16,G1177);
  nand (G1259,G1081,G1177);
  nand (G1260,G17,G1180);
  nand (G1261,G1084,G1180);
  nand (G1262,G18,G1183);
  nand (G1263,G1087,G1183);
  nand (G1264,G19,G1186);
  nand (G1265,G1090,G1186);
  nand (G1266,G20,G1189);
  nand (G1267,G1093,G1189);
  nand (G1268,G21,G1192);
  nand (G1269,G1096,G1192);
  nand (G1270,G22,G1195);
  nand (G1271,G1099,G1195);
  nand (G1272,G23,G1198);
  nand (G1273,G1102,G1198);
  nand (G1274,G24,G1201);
  nand (G1275,G1105,G1201);
  nand (G1276,G25,G1204);
  nand (G1277,G1108,G1204);
  nand (G1278,G26,G1207);
  nand (G1279,G1111,G1207);
  nand (G1280,G27,G1210);
  nand (G1281,G1114,G1210);
  nand (G1282,G28,G1213);
  nand (G1283,G1117,G1213);
  nand (G1284,G29,G1216);
  nand (G1285,G1120,G1216);
  nand (G1286,G30,G1219);
  nand (G1287,G1123,G1219);
  nand (G1288,G31,G1222);
  nand (G1289,G1126,G1222);
  nand (G1290,G32,G1225);
  nand (G1291,G1129,G1225);
  nand (G1292,G1228,G1229);
  nand (G1293,G1230,G1231);
  nand (G1294,G1232,G1233);
  nand (G1295,G1234,G1235);
  nand (G1296,G1236,G1237);
  nand (G1297,G1238,G1239);
  nand (G1298,G1240,G1241);
  nand (G1299,G1242,G1243);
  nand (G1300,G1244,G1245);
  nand (G1301,G1246,G1247);
  nand (G1302,G1248,G1249);
  nand (G1303,G1250,G1251);
  nand (G1304,G1252,G1253);
  nand (G1305,G1254,G1255);
  nand (G1306,G1256,G1257);
  nand (G1307,G1258,G1259);
  nand (G1308,G1260,G1261);
  nand (G1309,G1262,G1263);
  nand (G1310,G1264,G1265);
  nand (G1311,G1266,G1267);
  nand (G1312,G1268,G1269);
  nand (G1313,G1270,G1271);
  nand (G1314,G1272,G1273);
  nand (G1315,G1274,G1275);
  nand (G1316,G1276,G1277);
  nand (G1317,G1278,G1279);
  nand (G1318,G1280,G1281);
  nand (G1319,G1282,G1283);
  nand (G1320,G1284,G1285);
  nand (G1321,G1286,G1287);
  nand (G1322,G1288,G1289);
  nand (G1323,G1290,G1291);
  not (G1324,G1292);
  not (G1325,G1293);
  not (G1326,G1294);
  not (G1327,G1295);
  not (G1328,G1296);
  not (G1329,G1297);
  not (G1330,G1298);
  not (G1331,G1299);
  not (G1332,G1300);
  not (G1333,G1301);
  not (G1334,G1302);
  not (G1335,G1303);
  not (G1336,G1304);
  not (G1337,G1305);
  not (G1338,G1306);
  not (G1339,G1307);
  not (G1340,G1308);
  not (G1341,G1309);
  not (G1342,G1310);
  not (G1343,G1311);
  not (G1344,G1312);
  not (G1345,G1313);
  not (G1346,G1314);
  not (G1347,G1315);
  not (G1348,G1316);
  not (G1349,G1317);
  not (G1350,G1318);
  not (G1351,G1319);
  not (G1352,G1320);
  not (G1353,G1321);
  not (G1354,G1322);
  not (G1355,G1323);

endmodule
