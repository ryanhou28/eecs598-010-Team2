// Benchmark "mymod" written by ABC on Wed Nov  1 23:37:45 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41,
    G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
    G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
    G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
    G1354, G1355  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
    G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
    G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
    G1354, G1355;
  reg n621_lo, n630_lo, n633_lo, n642_lo, n645_lo, n654_lo, n657_lo,
    n666_lo, n669_lo, n678_lo, n681_lo, n690_lo, n693_lo, n702_lo, n705_lo,
    n714_lo, n717_lo, n726_lo, n729_lo, n738_lo, n741_lo, n750_lo, n753_lo,
    n762_lo, n765_lo, n774_lo, n777_lo, n786_lo, n789_lo, n798_lo, n801_lo,
    n810_lo, n813_lo, n822_lo, n825_lo, n834_lo, n837_lo, n846_lo, n849_lo,
    n858_lo, n861_lo, n870_lo, n873_lo, n882_lo, n885_lo, n894_lo, n897_lo,
    n906_lo, n909_lo, n918_lo, n921_lo, n930_lo, n933_lo, n942_lo, n945_lo,
    n954_lo, n957_lo, n966_lo, n969_lo, n978_lo, n981_lo, n990_lo, n993_lo,
    n1002_lo, n1005_lo, n1017_lo, n1029_lo, n1041_lo, n1053_lo, n1065_lo,
    n1077_lo, n1089_lo, n1101_lo, n602_o2, n639_o2, n678_o2, n658_o2,
    n783_o2, n802_o2, n726_o2, n763_o2, n1644_o2, n1645_o2, n1646_o2,
    n1647_o2, n1648_o2, n1649_o2, n1650_o2, n1651_o2, n1652_o2, n1653_o2,
    n1654_o2, n1655_o2, n1656_o2, n1657_o2, n1658_o2, n1659_o2, n1660_o2,
    n1661_o2, n1662_o2, n1663_o2, n1664_o2, n1665_o2, n1666_o2, n1667_o2,
    n1668_o2, n1669_o2, n1670_o2, n1671_o2, n1672_o2, n1673_o2, n1674_o2,
    n1675_o2, n685_o2, n680_o2, n822_o2, n843_o2, n842_o2, n681_o2,
    n684_o2, n686_o2, n823_o2, n683_o2, n688_o2, n803_o2, n862_o2, n764_o2,
    n863_o2, n886_o2, lo002_buf_o2, lo006_buf_o2, lo010_buf_o2,
    lo014_buf_o2, lo018_buf_o2, lo022_buf_o2, lo026_buf_o2, lo030_buf_o2,
    lo034_buf_o2, lo038_buf_o2, lo042_buf_o2, lo046_buf_o2, lo050_buf_o2,
    lo054_buf_o2, lo058_buf_o2, lo062_buf_o2, lo066_buf_o2, lo070_buf_o2,
    lo074_buf_o2, lo078_buf_o2, lo082_buf_o2, lo086_buf_o2, lo090_buf_o2,
    lo094_buf_o2, lo098_buf_o2, lo102_buf_o2, lo106_buf_o2, lo110_buf_o2,
    lo114_buf_o2, lo118_buf_o2, lo122_buf_o2, lo126_buf_o2, n600_o2,
    n601_o2, n637_o2, n638_o2, n676_o2, n677_o2, n656_o2, n657_o2, n781_o2,
    n782_o2, n800_o2, n801_o2, n724_o2, n725_o2, n761_o2, n762_o2,
    lo129_buf_o2, lo133_buf_o2, lo137_buf_o2, lo141_buf_o2, lo145_buf_o2,
    lo149_buf_o2, lo153_buf_o2, lo157_buf_o2, lo161_buf_o2, n571_o2,
    n708_o2, n608_o2, n665_o2, n705_o2, n645_o2, n745_o2, n742_o2, n568_o2,
    n717_o2, n605_o2, n662_o2, n714_o2, n642_o2, n754_o2, n751_o2, n584_o2,
    n770_o2, n789_o2, n581_o2, n695_o2, n732_o2, n593_o2, n590_o2, n630_o2,
    n767_o2, n786_o2, n627_o2, n692_o2, n729_o2, n621_o2, n618_o2;
  wire new_n510_, new_n512_, new_n514_, new_n516_, new_n518_, new_n520_,
    new_n522_, new_n524_, new_n526_, new_n528_, new_n530_, new_n532_,
    new_n534_, new_n536_, new_n538_, new_n540_, new_n542_, new_n544_,
    new_n546_, new_n548_, new_n550_, new_n552_, new_n554_, new_n556_,
    new_n558_, new_n560_, new_n562_, new_n564_, new_n566_, new_n568_,
    new_n570_, new_n572_, new_n574_, new_n576_, new_n578_, new_n580_,
    new_n582_, new_n584_, new_n586_, new_n588_, new_n590_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n724_, new_n726_, new_n728_,
    new_n730_, new_n732_, new_n734_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n758_, new_n760_,
    new_n762_, new_n764_, new_n766_, new_n768_, new_n770_, new_n772_,
    new_n774_, new_n776_, new_n778_, new_n780_, new_n782_, new_n784_,
    new_n786_, new_n788_, new_n790_, new_n792_, new_n794_, new_n796_,
    new_n798_, new_n800_, new_n802_, new_n804_, new_n806_, new_n808_,
    new_n810_, new_n812_, new_n814_, new_n816_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n854_, new_n856_, new_n858_, new_n860_,
    new_n862_, new_n864_, new_n866_, new_n868_, new_n870_, new_n872_,
    new_n874_, new_n876_, new_n878_, new_n880_, new_n882_, new_n884_,
    new_n886_, new_n888_, new_n890_, new_n892_, new_n894_, new_n896_,
    new_n898_, new_n900_, new_n902_, new_n904_, new_n906_, new_n908_,
    new_n910_, new_n912_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_,
    new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_,
    new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_,
    new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_,
    new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_,
    new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_,
    new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_,
    new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_,
    new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_,
    new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_,
    new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_,
    new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_,
    new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_,
    new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_,
    new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_,
    new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_,
    new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_,
    new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_,
    new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_,
    new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_,
    new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_,
    new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_,
    new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_,
    new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_,
    new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_,
    new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_,
    new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_,
    new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_,
    new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_,
    new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_,
    new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_,
    new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_,
    new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_,
    new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_,
    new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_,
    new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_,
    new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_,
    new_n1834_, new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_,
    new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_,
    new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_,
    new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_,
    new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_,
    new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_,
    new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_,
    new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_,
    new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_,
    new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_,
    new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_,
    new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_,
    new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_,
    new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_,
    new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_,
    new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_,
    new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_,
    new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_,
    new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_,
    new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_,
    new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_,
    new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_,
    new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_,
    new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_,
    new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_,
    new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_,
    new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_,
    new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_,
    new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_,
    new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_,
    new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_,
    new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_,
    new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_,
    new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_,
    new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_,
    new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_,
    new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_,
    new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_,
    new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_,
    new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_,
    new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_,
    new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_,
    new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_,
    new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_,
    new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_,
    new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_,
    new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_,
    new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_,
    new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_,
    new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_,
    new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_,
    n1699_li000_li000, n1708_li003_li003, n1711_li004_li004,
    n1720_li007_li007, n1723_li008_li008, n1732_li011_li011,
    n1735_li012_li012, n1744_li015_li015, n1747_li016_li016,
    n1756_li019_li019, n1759_li020_li020, n1768_li023_li023,
    n1771_li024_li024, n1780_li027_li027, n1783_li028_li028,
    n1792_li031_li031, n1795_li032_li032, n1804_li035_li035,
    n1807_li036_li036, n1816_li039_li039, n1819_li040_li040,
    n1828_li043_li043, n1831_li044_li044, n1840_li047_li047,
    n1843_li048_li048, n1852_li051_li051, n1855_li052_li052,
    n1864_li055_li055, n1867_li056_li056, n1876_li059_li059,
    n1879_li060_li060, n1888_li063_li063, n1891_li064_li064,
    n1900_li067_li067, n1903_li068_li068, n1912_li071_li071,
    n1915_li072_li072, n1924_li075_li075, n1927_li076_li076,
    n1936_li079_li079, n1939_li080_li080, n1948_li083_li083,
    n1951_li084_li084, n1960_li087_li087, n1963_li088_li088,
    n1972_li091_li091, n1975_li092_li092, n1984_li095_li095,
    n1987_li096_li096, n1996_li099_li099, n1999_li100_li100,
    n2008_li103_li103, n2011_li104_li104, n2020_li107_li107,
    n2023_li108_li108, n2032_li111_li111, n2035_li112_li112,
    n2044_li115_li115, n2047_li116_li116, n2056_li119_li119,
    n2059_li120_li120, n2068_li123_li123, n2071_li124_li124,
    n2080_li127_li127, n2083_li128_li128, n2095_li132_li132,
    n2107_li136_li136, n2119_li140_li140, n2131_li144_li144,
    n2143_li148_li148, n2155_li152_li152, n2167_li156_li156,
    n2179_li160_li160, n602_i2, n639_i2, n678_i2, n658_i2, n783_i2,
    n802_i2, n726_i2, n763_i2, n1644_i2, n1645_i2, n1646_i2, n1647_i2,
    n1648_i2, n1649_i2, n1650_i2, n1651_i2, n1652_i2, n1653_i2, n1654_i2,
    n1655_i2, n1656_i2, n1657_i2, n1658_i2, n1659_i2, n1660_i2, n1661_i2,
    n1662_i2, n1663_i2, n1664_i2, n1665_i2, n1666_i2, n1667_i2, n1668_i2,
    n1669_i2, n1670_i2, n1671_i2, n1672_i2, n1673_i2, n1674_i2, n1675_i2,
    n685_i2, n680_i2, n822_i2, n843_i2, n842_i2, n681_i2, n684_i2, n686_i2,
    n823_i2, n683_i2, n688_i2, n803_i2, n862_i2, n764_i2, n863_i2, n886_i2,
    lo002_buf_i2, lo006_buf_i2, lo010_buf_i2, lo014_buf_i2, lo018_buf_i2,
    lo022_buf_i2, lo026_buf_i2, lo030_buf_i2, lo034_buf_i2, lo038_buf_i2,
    lo042_buf_i2, lo046_buf_i2, lo050_buf_i2, lo054_buf_i2, lo058_buf_i2,
    lo062_buf_i2, lo066_buf_i2, lo070_buf_i2, lo074_buf_i2, lo078_buf_i2,
    lo082_buf_i2, lo086_buf_i2, lo090_buf_i2, lo094_buf_i2, lo098_buf_i2,
    lo102_buf_i2, lo106_buf_i2, lo110_buf_i2, lo114_buf_i2, lo118_buf_i2,
    lo122_buf_i2, lo126_buf_i2, n600_i2, n601_i2, n637_i2, n638_i2,
    n676_i2, n677_i2, n656_i2, n657_i2, n781_i2, n782_i2, n800_i2, n801_i2,
    n724_i2, n725_i2, n761_i2, n762_i2, lo129_buf_i2, lo133_buf_i2,
    lo137_buf_i2, lo141_buf_i2, lo145_buf_i2, lo149_buf_i2, lo153_buf_i2,
    lo157_buf_i2, lo161_buf_i2, n571_i2, n708_i2, n608_i2, n665_i2,
    n705_i2, n645_i2, n745_i2, n742_i2, n568_i2, n717_i2, n605_i2, n662_i2,
    n714_i2, n642_i2, n754_i2, n751_i2, n584_i2, n770_i2, n789_i2, n581_i2,
    n695_i2, n732_i2, n593_i2, n590_i2, n630_i2, n767_i2, n786_i2, n627_i2,
    n692_i2, n729_i2, n621_i2, n618_i2;
  assign new_n510_ = G1;
  assign new_n512_ = G2;
  assign new_n514_ = G3;
  assign new_n516_ = G4;
  assign new_n518_ = G5;
  assign new_n520_ = G6;
  assign new_n522_ = G7;
  assign new_n524_ = G8;
  assign new_n526_ = G9;
  assign new_n528_ = G10;
  assign new_n530_ = G11;
  assign new_n532_ = G12;
  assign new_n534_ = G13;
  assign new_n536_ = G14;
  assign new_n538_ = G15;
  assign new_n540_ = G16;
  assign new_n542_ = G17;
  assign new_n544_ = G18;
  assign new_n546_ = G19;
  assign new_n548_ = G20;
  assign new_n550_ = G21;
  assign new_n552_ = G22;
  assign new_n554_ = G23;
  assign new_n556_ = G24;
  assign new_n558_ = G25;
  assign new_n560_ = G26;
  assign new_n562_ = G27;
  assign new_n564_ = G28;
  assign new_n566_ = G29;
  assign new_n568_ = G30;
  assign new_n570_ = G31;
  assign new_n572_ = G32;
  assign new_n574_ = G33;
  assign new_n576_ = G34;
  assign new_n578_ = G35;
  assign new_n580_ = G36;
  assign new_n582_ = G37;
  assign new_n584_ = G38;
  assign new_n586_ = G39;
  assign new_n588_ = G40;
  assign new_n590_ = G41;
  assign new_n592_ = n621_lo;
  assign new_n593_ = ~n621_lo;
  assign new_n594_ = n630_lo;
  assign new_n595_ = ~n630_lo;
  assign new_n596_ = n633_lo;
  assign new_n597_ = ~n633_lo;
  assign new_n598_ = n642_lo;
  assign new_n599_ = ~n642_lo;
  assign new_n600_ = n645_lo;
  assign new_n601_ = ~n645_lo;
  assign new_n602_ = n654_lo;
  assign new_n603_ = ~n654_lo;
  assign new_n604_ = n657_lo;
  assign new_n605_ = ~n657_lo;
  assign new_n606_ = n666_lo;
  assign new_n607_ = ~n666_lo;
  assign new_n608_ = n669_lo;
  assign new_n609_ = ~n669_lo;
  assign new_n610_ = n678_lo;
  assign new_n611_ = ~n678_lo;
  assign new_n612_ = n681_lo;
  assign new_n613_ = ~n681_lo;
  assign new_n614_ = n690_lo;
  assign new_n615_ = ~n690_lo;
  assign new_n616_ = n693_lo;
  assign new_n617_ = ~n693_lo;
  assign new_n618_ = n702_lo;
  assign new_n619_ = ~n702_lo;
  assign new_n620_ = n705_lo;
  assign new_n621_ = ~n705_lo;
  assign new_n622_ = n714_lo;
  assign new_n623_ = ~n714_lo;
  assign new_n624_ = n717_lo;
  assign new_n625_ = ~n717_lo;
  assign new_n626_ = n726_lo;
  assign new_n627_ = ~n726_lo;
  assign new_n628_ = n729_lo;
  assign new_n629_ = ~n729_lo;
  assign new_n630_ = n738_lo;
  assign new_n631_ = ~n738_lo;
  assign new_n632_ = n741_lo;
  assign new_n633_ = ~n741_lo;
  assign new_n634_ = n750_lo;
  assign new_n635_ = ~n750_lo;
  assign new_n636_ = n753_lo;
  assign new_n637_ = ~n753_lo;
  assign new_n638_ = n762_lo;
  assign new_n639_ = ~n762_lo;
  assign new_n640_ = n765_lo;
  assign new_n641_ = ~n765_lo;
  assign new_n642_ = n774_lo;
  assign new_n643_ = ~n774_lo;
  assign new_n644_ = n777_lo;
  assign new_n645_ = ~n777_lo;
  assign new_n646_ = n786_lo;
  assign new_n647_ = ~n786_lo;
  assign new_n648_ = n789_lo;
  assign new_n649_ = ~n789_lo;
  assign new_n650_ = n798_lo;
  assign new_n651_ = ~n798_lo;
  assign new_n652_ = n801_lo;
  assign new_n653_ = ~n801_lo;
  assign new_n654_ = n810_lo;
  assign new_n655_ = ~n810_lo;
  assign new_n656_ = n813_lo;
  assign new_n657_ = ~n813_lo;
  assign new_n658_ = n822_lo;
  assign new_n659_ = ~n822_lo;
  assign new_n660_ = n825_lo;
  assign new_n661_ = ~n825_lo;
  assign new_n662_ = n834_lo;
  assign new_n663_ = ~n834_lo;
  assign new_n664_ = n837_lo;
  assign new_n665_ = ~n837_lo;
  assign new_n666_ = n846_lo;
  assign new_n667_ = ~n846_lo;
  assign new_n668_ = n849_lo;
  assign new_n669_ = ~n849_lo;
  assign new_n670_ = n858_lo;
  assign new_n671_ = ~n858_lo;
  assign new_n672_ = n861_lo;
  assign new_n673_ = ~n861_lo;
  assign new_n674_ = n870_lo;
  assign new_n675_ = ~n870_lo;
  assign new_n676_ = n873_lo;
  assign new_n677_ = ~n873_lo;
  assign new_n678_ = n882_lo;
  assign new_n679_ = ~n882_lo;
  assign new_n680_ = n885_lo;
  assign new_n681_ = ~n885_lo;
  assign new_n682_ = n894_lo;
  assign new_n683_ = ~n894_lo;
  assign new_n684_ = n897_lo;
  assign new_n685_ = ~n897_lo;
  assign new_n686_ = n906_lo;
  assign new_n687_ = ~n906_lo;
  assign new_n688_ = n909_lo;
  assign new_n689_ = ~n909_lo;
  assign new_n690_ = n918_lo;
  assign new_n691_ = ~n918_lo;
  assign new_n692_ = n921_lo;
  assign new_n693_ = ~n921_lo;
  assign new_n694_ = n930_lo;
  assign new_n695_ = ~n930_lo;
  assign new_n696_ = n933_lo;
  assign new_n697_ = ~n933_lo;
  assign new_n698_ = n942_lo;
  assign new_n699_ = ~n942_lo;
  assign new_n700_ = n945_lo;
  assign new_n701_ = ~n945_lo;
  assign new_n702_ = n954_lo;
  assign new_n703_ = ~n954_lo;
  assign new_n704_ = n957_lo;
  assign new_n705_ = ~n957_lo;
  assign new_n706_ = n966_lo;
  assign new_n707_ = ~n966_lo;
  assign new_n708_ = n969_lo;
  assign new_n709_ = ~n969_lo;
  assign new_n710_ = n978_lo;
  assign new_n711_ = ~n978_lo;
  assign new_n712_ = n981_lo;
  assign new_n713_ = ~n981_lo;
  assign new_n714_ = n990_lo;
  assign new_n715_ = ~n990_lo;
  assign new_n716_ = n993_lo;
  assign new_n717_ = ~n993_lo;
  assign new_n718_ = n1002_lo;
  assign new_n719_ = ~n1002_lo;
  assign new_n720_ = n1005_lo;
  assign new_n722_ = n1017_lo;
  assign new_n724_ = n1029_lo;
  assign new_n726_ = n1041_lo;
  assign new_n728_ = n1053_lo;
  assign new_n730_ = n1065_lo;
  assign new_n732_ = n1077_lo;
  assign new_n734_ = n1089_lo;
  assign new_n736_ = n1101_lo;
  assign new_n738_ = n602_o2;
  assign new_n739_ = ~n602_o2;
  assign new_n740_ = n639_o2;
  assign new_n741_ = ~n639_o2;
  assign new_n742_ = n678_o2;
  assign new_n743_ = ~n678_o2;
  assign new_n744_ = n658_o2;
  assign new_n745_ = ~n658_o2;
  assign new_n746_ = n783_o2;
  assign new_n747_ = ~n783_o2;
  assign new_n748_ = n802_o2;
  assign new_n749_ = ~n802_o2;
  assign new_n750_ = n726_o2;
  assign new_n751_ = ~n726_o2;
  assign new_n752_ = n763_o2;
  assign new_n753_ = ~n763_o2;
  assign new_n754_ = n1644_o2;
  assign new_n756_ = n1645_o2;
  assign new_n758_ = n1646_o2;
  assign new_n760_ = n1647_o2;
  assign new_n762_ = n1648_o2;
  assign new_n764_ = n1649_o2;
  assign new_n766_ = n1650_o2;
  assign new_n768_ = n1651_o2;
  assign new_n770_ = n1652_o2;
  assign new_n772_ = n1653_o2;
  assign new_n774_ = n1654_o2;
  assign new_n776_ = n1655_o2;
  assign new_n778_ = n1656_o2;
  assign new_n780_ = n1657_o2;
  assign new_n782_ = n1658_o2;
  assign new_n784_ = n1659_o2;
  assign new_n786_ = n1660_o2;
  assign new_n788_ = n1661_o2;
  assign new_n790_ = n1662_o2;
  assign new_n792_ = n1663_o2;
  assign new_n794_ = n1664_o2;
  assign new_n796_ = n1665_o2;
  assign new_n798_ = n1666_o2;
  assign new_n800_ = n1667_o2;
  assign new_n802_ = n1668_o2;
  assign new_n804_ = n1669_o2;
  assign new_n806_ = n1670_o2;
  assign new_n808_ = n1671_o2;
  assign new_n810_ = n1672_o2;
  assign new_n812_ = n1673_o2;
  assign new_n814_ = n1674_o2;
  assign new_n816_ = n1675_o2;
  assign new_n818_ = n685_o2;
  assign new_n819_ = ~n685_o2;
  assign new_n820_ = n680_o2;
  assign new_n821_ = ~n680_o2;
  assign new_n822_ = n822_o2;
  assign new_n823_ = ~n822_o2;
  assign new_n824_ = n843_o2;
  assign new_n825_ = ~n843_o2;
  assign new_n826_ = n842_o2;
  assign new_n827_ = ~n842_o2;
  assign new_n828_ = n681_o2;
  assign new_n829_ = ~n681_o2;
  assign new_n830_ = n684_o2;
  assign new_n831_ = ~n684_o2;
  assign new_n832_ = n686_o2;
  assign new_n833_ = ~n686_o2;
  assign new_n834_ = n823_o2;
  assign new_n835_ = ~n823_o2;
  assign new_n836_ = n683_o2;
  assign new_n837_ = ~n683_o2;
  assign new_n838_ = n688_o2;
  assign new_n839_ = ~n688_o2;
  assign new_n840_ = n803_o2;
  assign new_n841_ = ~n803_o2;
  assign new_n842_ = n862_o2;
  assign new_n843_ = ~n862_o2;
  assign new_n844_ = n764_o2;
  assign new_n845_ = ~n764_o2;
  assign new_n846_ = n863_o2;
  assign new_n847_ = ~n863_o2;
  assign new_n848_ = n886_o2;
  assign new_n849_ = ~n886_o2;
  assign new_n850_ = lo002_buf_o2;
  assign new_n852_ = lo006_buf_o2;
  assign new_n854_ = lo010_buf_o2;
  assign new_n856_ = lo014_buf_o2;
  assign new_n858_ = lo018_buf_o2;
  assign new_n860_ = lo022_buf_o2;
  assign new_n862_ = lo026_buf_o2;
  assign new_n864_ = lo030_buf_o2;
  assign new_n866_ = lo034_buf_o2;
  assign new_n868_ = lo038_buf_o2;
  assign new_n870_ = lo042_buf_o2;
  assign new_n872_ = lo046_buf_o2;
  assign new_n874_ = lo050_buf_o2;
  assign new_n876_ = lo054_buf_o2;
  assign new_n878_ = lo058_buf_o2;
  assign new_n880_ = lo062_buf_o2;
  assign new_n882_ = lo066_buf_o2;
  assign new_n884_ = lo070_buf_o2;
  assign new_n886_ = lo074_buf_o2;
  assign new_n888_ = lo078_buf_o2;
  assign new_n890_ = lo082_buf_o2;
  assign new_n892_ = lo086_buf_o2;
  assign new_n894_ = lo090_buf_o2;
  assign new_n896_ = lo094_buf_o2;
  assign new_n898_ = lo098_buf_o2;
  assign new_n900_ = lo102_buf_o2;
  assign new_n902_ = lo106_buf_o2;
  assign new_n904_ = lo110_buf_o2;
  assign new_n906_ = lo114_buf_o2;
  assign new_n908_ = lo118_buf_o2;
  assign new_n910_ = lo122_buf_o2;
  assign new_n912_ = lo126_buf_o2;
  assign new_n914_ = n600_o2;
  assign new_n915_ = ~n600_o2;
  assign new_n916_ = n601_o2;
  assign new_n917_ = ~n601_o2;
  assign new_n918_ = n637_o2;
  assign new_n919_ = ~n637_o2;
  assign new_n920_ = n638_o2;
  assign new_n921_ = ~n638_o2;
  assign new_n922_ = n676_o2;
  assign new_n923_ = ~n676_o2;
  assign new_n924_ = n677_o2;
  assign new_n925_ = ~n677_o2;
  assign new_n926_ = n656_o2;
  assign new_n927_ = ~n656_o2;
  assign new_n928_ = n657_o2;
  assign new_n929_ = ~n657_o2;
  assign new_n930_ = n781_o2;
  assign new_n931_ = ~n781_o2;
  assign new_n932_ = n782_o2;
  assign new_n933_ = ~n782_o2;
  assign new_n934_ = n800_o2;
  assign new_n935_ = ~n800_o2;
  assign new_n936_ = n801_o2;
  assign new_n937_ = ~n801_o2;
  assign new_n938_ = n724_o2;
  assign new_n939_ = ~n724_o2;
  assign new_n940_ = n725_o2;
  assign new_n941_ = ~n725_o2;
  assign new_n942_ = n761_o2;
  assign new_n943_ = ~n761_o2;
  assign new_n944_ = n762_o2;
  assign new_n945_ = ~n762_o2;
  assign new_n946_ = lo129_buf_o2;
  assign new_n947_ = ~lo129_buf_o2;
  assign new_n948_ = lo133_buf_o2;
  assign new_n949_ = ~lo133_buf_o2;
  assign new_n950_ = lo137_buf_o2;
  assign new_n951_ = ~lo137_buf_o2;
  assign new_n952_ = lo141_buf_o2;
  assign new_n953_ = ~lo141_buf_o2;
  assign new_n954_ = lo145_buf_o2;
  assign new_n955_ = ~lo145_buf_o2;
  assign new_n956_ = lo149_buf_o2;
  assign new_n957_ = ~lo149_buf_o2;
  assign new_n958_ = lo153_buf_o2;
  assign new_n959_ = ~lo153_buf_o2;
  assign new_n960_ = lo157_buf_o2;
  assign new_n961_ = ~lo157_buf_o2;
  assign new_n962_ = lo161_buf_o2;
  assign new_n963_ = ~lo161_buf_o2;
  assign new_n964_ = n571_o2;
  assign new_n965_ = ~n571_o2;
  assign new_n966_ = n708_o2;
  assign new_n967_ = ~n708_o2;
  assign new_n968_ = n608_o2;
  assign new_n969_ = ~n608_o2;
  assign new_n970_ = n665_o2;
  assign new_n971_ = ~n665_o2;
  assign new_n972_ = n705_o2;
  assign new_n973_ = ~n705_o2;
  assign new_n974_ = n645_o2;
  assign new_n975_ = ~n645_o2;
  assign new_n976_ = n745_o2;
  assign new_n977_ = ~n745_o2;
  assign new_n978_ = n742_o2;
  assign new_n979_ = ~n742_o2;
  assign new_n980_ = n568_o2;
  assign new_n981_ = ~n568_o2;
  assign new_n982_ = n717_o2;
  assign new_n983_ = ~n717_o2;
  assign new_n984_ = n605_o2;
  assign new_n985_ = ~n605_o2;
  assign new_n986_ = n662_o2;
  assign new_n987_ = ~n662_o2;
  assign new_n988_ = n714_o2;
  assign new_n989_ = ~n714_o2;
  assign new_n990_ = n642_o2;
  assign new_n991_ = ~n642_o2;
  assign new_n992_ = n754_o2;
  assign new_n993_ = ~n754_o2;
  assign new_n994_ = n751_o2;
  assign new_n995_ = ~n751_o2;
  assign new_n996_ = n584_o2;
  assign new_n997_ = ~n584_o2;
  assign new_n998_ = n770_o2;
  assign new_n999_ = ~n770_o2;
  assign new_n1000_ = n789_o2;
  assign new_n1001_ = ~n789_o2;
  assign new_n1002_ = n581_o2;
  assign new_n1003_ = ~n581_o2;
  assign new_n1004_ = n695_o2;
  assign new_n1005_ = ~n695_o2;
  assign new_n1006_ = n732_o2;
  assign new_n1007_ = ~n732_o2;
  assign new_n1008_ = n593_o2;
  assign new_n1009_ = ~n593_o2;
  assign new_n1010_ = n590_o2;
  assign new_n1011_ = ~n590_o2;
  assign new_n1012_ = n630_o2;
  assign new_n1013_ = ~n630_o2;
  assign new_n1014_ = n767_o2;
  assign new_n1015_ = ~n767_o2;
  assign new_n1016_ = n786_o2;
  assign new_n1017_ = ~n786_o2;
  assign new_n1018_ = n627_o2;
  assign new_n1019_ = ~n627_o2;
  assign new_n1020_ = n692_o2;
  assign new_n1021_ = ~n692_o2;
  assign new_n1022_ = n729_o2;
  assign new_n1023_ = ~n729_o2;
  assign new_n1024_ = n621_o2;
  assign new_n1025_ = ~n621_o2;
  assign new_n1026_ = n618_o2;
  assign new_n1027_ = ~n618_o2;
  assign new_n1028_ = new_n837_ & new_n839_;
  assign new_n1029_ = new_n836_ | new_n838_;
  assign new_n1030_ = new_n840_ & new_n844_;
  assign new_n1031_ = new_n841_ | new_n845_;
  assign new_n1032_ = new_n1787_ & new_n1030_;
  assign new_n1033_ = new_n1790_ | new_n1031_;
  assign new_n1034_ = new_n1793_ & new_n1796_;
  assign new_n1035_ = new_n1799_ | new_n1802_;
  assign new_n1036_ = new_n595_ | new_n1034_;
  assign new_n1037_ = new_n594_ | new_n1035_;
  assign new_n1038_ = new_n1036_ & new_n1037_;
  assign new_n1039_ = new_n1806_ & new_n1796_;
  assign new_n1040_ = new_n1810_ | new_n1802_;
  assign new_n1041_ = new_n599_ | new_n1039_;
  assign new_n1042_ = new_n598_ | new_n1040_;
  assign new_n1043_ = new_n1041_ & new_n1042_;
  assign new_n1044_ = new_n1814_ & new_n1797_;
  assign new_n1045_ = new_n1819_ | new_n1803_;
  assign new_n1046_ = new_n603_ | new_n1044_;
  assign new_n1047_ = new_n602_ | new_n1045_;
  assign new_n1048_ = new_n1046_ & new_n1047_;
  assign new_n1049_ = new_n1823_ & new_n1797_;
  assign new_n1050_ = new_n1826_ | new_n1803_;
  assign new_n1051_ = new_n607_ | new_n1049_;
  assign new_n1052_ = new_n606_ | new_n1050_;
  assign new_n1053_ = new_n1051_ & new_n1052_;
  assign new_n1054_ = new_n822_ & new_n835_;
  assign new_n1055_ = new_n823_ | new_n834_;
  assign new_n1056_ = new_n1787_ & new_n1054_;
  assign new_n1057_ = new_n1790_ | new_n1055_;
  assign new_n1058_ = new_n1793_ & new_n1829_;
  assign new_n1059_ = new_n1799_ | new_n1832_;
  assign new_n1060_ = new_n611_ | new_n1058_;
  assign new_n1061_ = new_n610_ | new_n1059_;
  assign new_n1062_ = new_n1060_ & new_n1061_;
  assign new_n1063_ = new_n1806_ & new_n1829_;
  assign new_n1064_ = new_n1810_ | new_n1832_;
  assign new_n1065_ = new_n615_ | new_n1063_;
  assign new_n1066_ = new_n614_ | new_n1064_;
  assign new_n1067_ = new_n1065_ & new_n1066_;
  assign new_n1068_ = new_n1814_ & new_n1830_;
  assign new_n1069_ = new_n1819_ | new_n1833_;
  assign new_n1070_ = new_n619_ | new_n1068_;
  assign new_n1071_ = new_n618_ | new_n1069_;
  assign new_n1072_ = new_n1070_ & new_n1071_;
  assign new_n1073_ = new_n1823_ & new_n1830_;
  assign new_n1074_ = new_n1826_ | new_n1833_;
  assign new_n1075_ = new_n623_ | new_n1073_;
  assign new_n1076_ = new_n622_ | new_n1074_;
  assign new_n1077_ = new_n1075_ & new_n1076_;
  assign new_n1078_ = new_n825_ & new_n826_;
  assign new_n1079_ = new_n824_ | new_n827_;
  assign new_n1080_ = new_n1788_ & new_n1078_;
  assign new_n1081_ = new_n1791_ | new_n1079_;
  assign new_n1082_ = new_n1794_ & new_n1835_;
  assign new_n1083_ = new_n1800_ | new_n1838_;
  assign new_n1084_ = new_n627_ | new_n1082_;
  assign new_n1085_ = new_n626_ | new_n1083_;
  assign new_n1086_ = new_n1084_ & new_n1085_;
  assign new_n1087_ = new_n1805_ & new_n1835_;
  assign new_n1088_ = new_n1809_ | new_n1838_;
  assign new_n1089_ = new_n631_ | new_n1087_;
  assign new_n1090_ = new_n630_ | new_n1088_;
  assign new_n1091_ = new_n1089_ & new_n1090_;
  assign new_n1092_ = new_n1815_ & new_n1836_;
  assign new_n1093_ = new_n1820_ | new_n1839_;
  assign new_n1094_ = new_n635_ | new_n1092_;
  assign new_n1095_ = new_n634_ | new_n1093_;
  assign new_n1096_ = new_n1094_ & new_n1095_;
  assign new_n1097_ = new_n1824_ & new_n1836_;
  assign new_n1098_ = new_n1827_ | new_n1839_;
  assign new_n1099_ = new_n639_ | new_n1097_;
  assign new_n1100_ = new_n638_ | new_n1098_;
  assign new_n1101_ = new_n1099_ & new_n1100_;
  assign new_n1102_ = new_n842_ & new_n846_;
  assign new_n1103_ = new_n843_ | new_n847_;
  assign new_n1104_ = new_n1788_ & new_n1102_;
  assign new_n1105_ = new_n1791_ | new_n1103_;
  assign new_n1106_ = new_n1794_ & new_n1841_;
  assign new_n1107_ = new_n1800_ | new_n1844_;
  assign new_n1108_ = new_n643_ | new_n1106_;
  assign new_n1109_ = new_n642_ | new_n1107_;
  assign new_n1110_ = new_n1108_ & new_n1109_;
  assign new_n1111_ = new_n1807_ & new_n1841_;
  assign new_n1112_ = new_n1811_ | new_n1844_;
  assign new_n1113_ = new_n647_ | new_n1111_;
  assign new_n1114_ = new_n646_ | new_n1112_;
  assign new_n1115_ = new_n1113_ & new_n1114_;
  assign new_n1116_ = new_n1815_ & new_n1842_;
  assign new_n1117_ = new_n1820_ | new_n1845_;
  assign new_n1118_ = new_n651_ | new_n1116_;
  assign new_n1119_ = new_n650_ | new_n1117_;
  assign new_n1120_ = new_n1118_ & new_n1119_;
  assign new_n1121_ = new_n1824_ & new_n1842_;
  assign new_n1122_ = new_n1827_ | new_n1845_;
  assign new_n1123_ = new_n655_ | new_n1121_;
  assign new_n1124_ = new_n654_ | new_n1122_;
  assign new_n1125_ = new_n1123_ & new_n1124_;
  assign new_n1126_ = new_n832_ & new_n1847_;
  assign new_n1127_ = new_n833_ | new_n1850_;
  assign new_n1128_ = new_n1816_ & new_n1126_;
  assign new_n1129_ = new_n1821_ | new_n1127_;
  assign new_n1130_ = new_n1853_ & new_n1856_;
  assign new_n1131_ = new_n1859_ | new_n1862_;
  assign new_n1132_ = new_n659_ | new_n1130_;
  assign new_n1133_ = new_n658_ | new_n1131_;
  assign new_n1134_ = new_n1132_ & new_n1133_;
  assign new_n1135_ = new_n1865_ & new_n1856_;
  assign new_n1136_ = new_n1868_ | new_n1862_;
  assign new_n1137_ = new_n663_ | new_n1135_;
  assign new_n1138_ = new_n662_ | new_n1136_;
  assign new_n1139_ = new_n1137_ & new_n1138_;
  assign new_n1140_ = new_n1871_ & new_n1857_;
  assign new_n1141_ = new_n1874_ | new_n1863_;
  assign new_n1142_ = new_n667_ | new_n1140_;
  assign new_n1143_ = new_n666_ | new_n1141_;
  assign new_n1144_ = new_n1142_ & new_n1143_;
  assign new_n1145_ = new_n1877_ & new_n1857_;
  assign new_n1146_ = new_n1880_ | new_n1863_;
  assign new_n1147_ = new_n671_ | new_n1145_;
  assign new_n1148_ = new_n670_ | new_n1146_;
  assign new_n1149_ = new_n1147_ & new_n1148_;
  assign new_n1150_ = new_n818_ & new_n820_;
  assign new_n1151_ = new_n819_ | new_n821_;
  assign new_n1152_ = new_n1847_ & new_n1150_;
  assign new_n1153_ = new_n1850_ | new_n1151_;
  assign new_n1154_ = new_n1853_ & new_n1883_;
  assign new_n1155_ = new_n1859_ | new_n1886_;
  assign new_n1156_ = new_n675_ | new_n1154_;
  assign new_n1157_ = new_n674_ | new_n1155_;
  assign new_n1158_ = new_n1156_ & new_n1157_;
  assign new_n1159_ = new_n1865_ & new_n1883_;
  assign new_n1160_ = new_n1868_ | new_n1886_;
  assign new_n1161_ = new_n679_ | new_n1159_;
  assign new_n1162_ = new_n678_ | new_n1160_;
  assign new_n1163_ = new_n1161_ & new_n1162_;
  assign new_n1164_ = new_n1871_ & new_n1884_;
  assign new_n1165_ = new_n1874_ | new_n1887_;
  assign new_n1166_ = new_n683_ | new_n1164_;
  assign new_n1167_ = new_n682_ | new_n1165_;
  assign new_n1168_ = new_n1166_ & new_n1167_;
  assign new_n1169_ = new_n1877_ & new_n1884_;
  assign new_n1170_ = new_n1880_ | new_n1887_;
  assign new_n1171_ = new_n687_ | new_n1169_;
  assign new_n1172_ = new_n686_ | new_n1170_;
  assign new_n1173_ = new_n1171_ & new_n1172_;
  assign new_n1174_ = new_n1816_ & new_n830_;
  assign new_n1175_ = new_n1821_ | new_n831_;
  assign new_n1176_ = new_n1848_ & new_n1174_;
  assign new_n1177_ = new_n1851_ | new_n1175_;
  assign new_n1178_ = new_n1854_ & new_n1889_;
  assign new_n1179_ = new_n1860_ | new_n1892_;
  assign new_n1180_ = new_n691_ | new_n1178_;
  assign new_n1181_ = new_n690_ | new_n1179_;
  assign new_n1182_ = new_n1180_ & new_n1181_;
  assign new_n1183_ = new_n1866_ & new_n1889_;
  assign new_n1184_ = new_n1869_ | new_n1892_;
  assign new_n1185_ = new_n695_ | new_n1183_;
  assign new_n1186_ = new_n694_ | new_n1184_;
  assign new_n1187_ = new_n1185_ & new_n1186_;
  assign new_n1188_ = new_n1872_ & new_n1890_;
  assign new_n1189_ = new_n1875_ | new_n1893_;
  assign new_n1190_ = new_n699_ | new_n1188_;
  assign new_n1191_ = new_n698_ | new_n1189_;
  assign new_n1192_ = new_n1190_ & new_n1191_;
  assign new_n1193_ = new_n1878_ & new_n1890_;
  assign new_n1194_ = new_n1881_ | new_n1893_;
  assign new_n1195_ = new_n703_ | new_n1193_;
  assign new_n1196_ = new_n702_ | new_n1194_;
  assign new_n1197_ = new_n1195_ & new_n1196_;
  assign new_n1198_ = new_n1807_ & new_n828_;
  assign new_n1199_ = new_n1811_ | new_n829_;
  assign new_n1200_ = new_n1848_ & new_n1198_;
  assign new_n1201_ = new_n1851_ | new_n1199_;
  assign new_n1202_ = new_n1854_ & new_n1895_;
  assign new_n1203_ = new_n1860_ | new_n1898_;
  assign new_n1204_ = new_n707_ | new_n1202_;
  assign new_n1205_ = new_n706_ | new_n1203_;
  assign new_n1206_ = new_n1204_ & new_n1205_;
  assign new_n1207_ = new_n1866_ & new_n1895_;
  assign new_n1208_ = new_n1869_ | new_n1898_;
  assign new_n1209_ = new_n711_ | new_n1207_;
  assign new_n1210_ = new_n710_ | new_n1208_;
  assign new_n1211_ = new_n1209_ & new_n1210_;
  assign new_n1212_ = new_n1872_ & new_n1896_;
  assign new_n1213_ = new_n1875_ | new_n1899_;
  assign new_n1214_ = new_n715_ | new_n1212_;
  assign new_n1215_ = new_n714_ | new_n1213_;
  assign new_n1216_ = new_n1214_ & new_n1215_;
  assign new_n1217_ = new_n1878_ & new_n1896_;
  assign new_n1218_ = new_n1881_ | new_n1899_;
  assign new_n1219_ = new_n719_ | new_n1217_;
  assign new_n1220_ = new_n718_ | new_n1218_;
  assign new_n1221_ = new_n1219_ & new_n1220_;
  assign new_n1222_ = new_n915_ & new_n917_;
  assign new_n1223_ = new_n914_ | new_n916_;
  assign new_n1224_ = new_n919_ & new_n921_;
  assign new_n1225_ = new_n918_ | new_n920_;
  assign new_n1226_ = new_n923_ & new_n925_;
  assign new_n1227_ = new_n922_ | new_n924_;
  assign new_n1228_ = new_n927_ & new_n929_;
  assign new_n1229_ = new_n926_ | new_n928_;
  assign new_n1230_ = new_n931_ & new_n933_;
  assign new_n1231_ = new_n930_ | new_n932_;
  assign new_n1232_ = new_n935_ & new_n937_;
  assign new_n1233_ = new_n934_ | new_n936_;
  assign new_n1234_ = new_n939_ & new_n941_;
  assign new_n1235_ = new_n938_ | new_n940_;
  assign new_n1236_ = new_n943_ & new_n945_;
  assign new_n1237_ = new_n942_ | new_n944_;
  assign new_n1238_ = new_n1222_ | new_n1901_;
  assign new_n1239_ = new_n1903_ | new_n1228_;
  assign new_n1240_ = new_n1905_ | new_n1907_;
  assign new_n1241_ = new_n1905_ & new_n1907_;
  assign new_n1242_ = new_n1909_ | new_n1911_;
  assign new_n1243_ = new_n1913_ | new_n1915_;
  assign new_n1244_ = new_n1917_ | new_n1918_;
  assign new_n1245_ = new_n1917_ | new_n1920_;
  assign new_n1246_ = new_n1224_ | new_n1921_;
  assign new_n1247_ = new_n1920_ | new_n1922_;
  assign new_n1248_ = new_n1913_ & new_n1915_;
  assign new_n1249_ = new_n1924_ | new_n1926_;
  assign new_n1250_ = new_n1226_ | new_n1921_;
  assign new_n1251_ = new_n1927_ & new_n1250_;
  assign new_n1252_ = new_n1901_ | new_n1251_;
  assign new_n1253_ = new_n1928_ & new_n1929_;
  assign new_n1254_ = new_n1903_ | new_n1253_;
  assign new_n1255_ = new_n1909_ & new_n1912_;
  assign new_n1256_ = new_n1904_ & new_n1924_;
  assign new_n1257_ = new_n1926_ & new_n1906_;
  assign new_n1258_ = new_n1914_ & new_n1911_;
  assign new_n1259_ = new_n1930_ & new_n1931_;
  assign new_n1260_ = new_n1932_ | new_n1259_;
  assign new_n1261_ = new_n1241_ & new_n1933_;
  assign new_n1262_ = new_n1248_ | new_n1261_;
  assign new_n1263_ = new_n1260_ & new_n1262_;
  assign new_n1264_ = new_n1934_ & new_n1935_;
  assign new_n1265_ = new_n1936_ | new_n1937_;
  assign new_n1266_ = new_n1936_ & new_n1937_;
  assign new_n1267_ = new_n1934_ | new_n1935_;
  assign new_n1268_ = new_n1265_ & new_n1267_;
  assign new_n1269_ = new_n1264_ | new_n1266_;
  assign new_n1270_ = new_n946_ & new_n1940_;
  assign new_n1271_ = new_n947_ | new_n1947_;
  assign new_n1272_ = new_n1269_ & new_n1270_;
  assign new_n1273_ = new_n1268_ & new_n1271_;
  assign new_n1274_ = new_n1272_ | new_n1273_;
  assign new_n1275_ = new_n1952_ & new_n1953_;
  assign new_n1276_ = new_n1954_ | new_n1955_;
  assign new_n1277_ = new_n1954_ & new_n1955_;
  assign new_n1278_ = new_n1952_ | new_n1953_;
  assign new_n1279_ = new_n1276_ & new_n1278_;
  assign new_n1280_ = new_n1275_ | new_n1277_;
  assign new_n1281_ = new_n1956_ & new_n1957_;
  assign new_n1282_ = new_n1958_ | new_n1959_;
  assign new_n1283_ = new_n1958_ & new_n1959_;
  assign new_n1284_ = new_n1956_ | new_n1957_;
  assign new_n1285_ = new_n1282_ & new_n1284_;
  assign new_n1286_ = new_n1281_ | new_n1283_;
  assign new_n1287_ = new_n1960_ & new_n1961_;
  assign new_n1288_ = new_n1962_ & new_n1963_;
  assign new_n1289_ = new_n1287_ | new_n1288_;
  assign new_n1290_ = new_n1964_ & new_n1965_;
  assign new_n1291_ = new_n1964_ | new_n1965_;
  assign new_n1292_ = new_n1966_ & new_n1967_;
  assign new_n1293_ = new_n1968_ | new_n1969_;
  assign new_n1294_ = new_n1968_ & new_n1969_;
  assign new_n1295_ = new_n1966_ | new_n1967_;
  assign new_n1296_ = new_n1293_ & new_n1295_;
  assign new_n1297_ = new_n1292_ | new_n1294_;
  assign new_n1298_ = new_n948_ & new_n1940_;
  assign new_n1299_ = new_n949_ | new_n1947_;
  assign new_n1300_ = new_n1297_ & new_n1298_;
  assign new_n1301_ = new_n1296_ & new_n1299_;
  assign new_n1302_ = new_n1300_ | new_n1301_;
  assign new_n1303_ = new_n1970_ & new_n1971_;
  assign new_n1304_ = new_n1972_ | new_n1973_;
  assign new_n1305_ = new_n1972_ & new_n1973_;
  assign new_n1306_ = new_n1970_ | new_n1971_;
  assign new_n1307_ = new_n1304_ & new_n1306_;
  assign new_n1308_ = new_n1303_ | new_n1305_;
  assign new_n1309_ = new_n1974_ & new_n1975_;
  assign new_n1310_ = new_n1976_ | new_n1977_;
  assign new_n1311_ = new_n1976_ & new_n1977_;
  assign new_n1312_ = new_n1974_ | new_n1975_;
  assign new_n1313_ = new_n1310_ & new_n1312_;
  assign new_n1314_ = new_n1309_ | new_n1311_;
  assign new_n1315_ = new_n1978_ & new_n1979_;
  assign new_n1316_ = new_n1980_ & new_n1981_;
  assign new_n1317_ = new_n1315_ | new_n1316_;
  assign new_n1318_ = new_n1982_ & new_n1983_;
  assign new_n1319_ = new_n1982_ | new_n1983_;
  assign new_n1320_ = new_n1984_ & new_n1985_;
  assign new_n1321_ = new_n1986_ | new_n1987_;
  assign new_n1322_ = new_n1986_ & new_n1987_;
  assign new_n1323_ = new_n1984_ | new_n1985_;
  assign new_n1324_ = new_n1321_ & new_n1323_;
  assign new_n1325_ = new_n1320_ | new_n1322_;
  assign new_n1326_ = new_n950_ & new_n1941_;
  assign new_n1327_ = new_n951_ | new_n1948_;
  assign new_n1328_ = new_n1325_ & new_n1326_;
  assign new_n1329_ = new_n1324_ & new_n1327_;
  assign new_n1330_ = new_n1328_ | new_n1329_;
  assign new_n1331_ = new_n1960_ & new_n1979_;
  assign new_n1332_ = new_n1962_ & new_n1981_;
  assign new_n1333_ = new_n1331_ | new_n1332_;
  assign new_n1334_ = new_n1988_ & new_n1989_;
  assign new_n1335_ = new_n1988_ | new_n1989_;
  assign new_n1336_ = new_n1990_ & new_n1991_;
  assign new_n1337_ = new_n1992_ | new_n1993_;
  assign new_n1338_ = new_n1992_ & new_n1993_;
  assign new_n1339_ = new_n1990_ | new_n1991_;
  assign new_n1340_ = new_n1337_ & new_n1339_;
  assign new_n1341_ = new_n1336_ | new_n1338_;
  assign new_n1342_ = new_n952_ & new_n1941_;
  assign new_n1343_ = new_n953_ | new_n1948_;
  assign new_n1344_ = new_n1341_ & new_n1342_;
  assign new_n1345_ = new_n1340_ & new_n1343_;
  assign new_n1346_ = new_n1344_ | new_n1345_;
  assign new_n1347_ = new_n1963_ & new_n1980_;
  assign new_n1348_ = new_n1961_ & new_n1978_;
  assign new_n1349_ = new_n1347_ | new_n1348_;
  assign new_n1350_ = new_n1994_ & new_n1995_;
  assign new_n1351_ = new_n1994_ | new_n1995_;
  assign new_n1352_ = new_n1996_ & new_n1997_;
  assign new_n1353_ = new_n1998_ | new_n1999_;
  assign new_n1354_ = new_n1998_ & new_n1999_;
  assign new_n1355_ = new_n1996_ | new_n1997_;
  assign new_n1356_ = new_n1353_ & new_n1355_;
  assign new_n1357_ = new_n1352_ | new_n1354_;
  assign new_n1358_ = new_n954_ & new_n1943_;
  assign new_n1359_ = new_n955_ | new_n1950_;
  assign new_n1360_ = new_n1357_ & new_n1358_;
  assign new_n1361_ = new_n1356_ & new_n1359_;
  assign new_n1362_ = new_n1360_ | new_n1361_;
  assign new_n1363_ = new_n2000_ & new_n2001_;
  assign new_n1364_ = new_n2002_ | new_n2003_;
  assign new_n1365_ = new_n2002_ & new_n2003_;
  assign new_n1366_ = new_n2000_ | new_n2001_;
  assign new_n1367_ = new_n1364_ & new_n1366_;
  assign new_n1368_ = new_n1363_ | new_n1365_;
  assign new_n1369_ = new_n2004_ & new_n2005_;
  assign new_n1370_ = new_n2006_ | new_n2007_;
  assign new_n1371_ = new_n2006_ & new_n2007_;
  assign new_n1372_ = new_n2004_ | new_n2005_;
  assign new_n1373_ = new_n1370_ & new_n1372_;
  assign new_n1374_ = new_n1369_ | new_n1371_;
  assign new_n1375_ = new_n2008_ & new_n2009_;
  assign new_n1376_ = new_n2010_ & new_n2011_;
  assign new_n1377_ = new_n1375_ | new_n1376_;
  assign new_n1378_ = new_n2012_ & new_n2013_;
  assign new_n1379_ = new_n2012_ | new_n2013_;
  assign new_n1380_ = new_n2014_ & new_n2015_;
  assign new_n1381_ = new_n2016_ | new_n2017_;
  assign new_n1382_ = new_n2016_ & new_n2017_;
  assign new_n1383_ = new_n2014_ | new_n2015_;
  assign new_n1384_ = new_n1381_ & new_n1383_;
  assign new_n1385_ = new_n1380_ | new_n1382_;
  assign new_n1386_ = new_n956_ & new_n1943_;
  assign new_n1387_ = new_n957_ | new_n1950_;
  assign new_n1388_ = new_n1385_ & new_n1386_;
  assign new_n1389_ = new_n1384_ & new_n1387_;
  assign new_n1390_ = new_n1388_ | new_n1389_;
  assign new_n1391_ = new_n2018_ & new_n2019_;
  assign new_n1392_ = new_n2020_ | new_n2021_;
  assign new_n1393_ = new_n2020_ & new_n2021_;
  assign new_n1394_ = new_n2018_ | new_n2019_;
  assign new_n1395_ = new_n1392_ & new_n1394_;
  assign new_n1396_ = new_n1391_ | new_n1393_;
  assign new_n1397_ = new_n2022_ & new_n2023_;
  assign new_n1398_ = new_n2024_ | new_n2025_;
  assign new_n1399_ = new_n2024_ & new_n2025_;
  assign new_n1400_ = new_n2022_ | new_n2023_;
  assign new_n1401_ = new_n1398_ & new_n1400_;
  assign new_n1402_ = new_n1397_ | new_n1399_;
  assign new_n1403_ = new_n2026_ & new_n2027_;
  assign new_n1404_ = new_n2028_ & new_n2029_;
  assign new_n1405_ = new_n1403_ | new_n1404_;
  assign new_n1406_ = new_n2030_ & new_n2031_;
  assign new_n1407_ = new_n2030_ | new_n2031_;
  assign new_n1408_ = new_n2032_ & new_n2033_;
  assign new_n1409_ = new_n2034_ | new_n2035_;
  assign new_n1410_ = new_n2034_ & new_n2035_;
  assign new_n1411_ = new_n2032_ | new_n2033_;
  assign new_n1412_ = new_n1409_ & new_n1411_;
  assign new_n1413_ = new_n1408_ | new_n1410_;
  assign new_n1414_ = new_n958_ & new_n1944_;
  assign new_n1415_ = new_n959_ | new_n1951_;
  assign new_n1416_ = new_n1413_ & new_n1414_;
  assign new_n1417_ = new_n1412_ & new_n1415_;
  assign new_n1418_ = new_n1416_ | new_n1417_;
  assign new_n1419_ = new_n2008_ & new_n2028_;
  assign new_n1420_ = new_n2010_ & new_n2026_;
  assign new_n1421_ = new_n1419_ | new_n1420_;
  assign new_n1422_ = new_n2036_ & new_n2037_;
  assign new_n1423_ = new_n2036_ | new_n2037_;
  assign new_n1424_ = new_n2038_ & new_n2039_;
  assign new_n1425_ = new_n2040_ | new_n2041_;
  assign new_n1426_ = new_n2040_ & new_n2041_;
  assign new_n1427_ = new_n2038_ | new_n2039_;
  assign new_n1428_ = new_n1425_ & new_n1427_;
  assign new_n1429_ = new_n1424_ | new_n1426_;
  assign new_n1430_ = new_n960_ & new_n1944_;
  assign new_n1431_ = new_n961_ | new_n1951_;
  assign new_n1432_ = new_n1429_ & new_n1430_;
  assign new_n1433_ = new_n1428_ & new_n1431_;
  assign new_n1434_ = new_n1432_ | new_n1433_;
  assign new_n1435_ = new_n2011_ & new_n2027_;
  assign new_n1436_ = new_n2009_ & new_n2029_;
  assign new_n1437_ = new_n1435_ | new_n1436_;
  assign new_n1438_ = new_n2042_ & new_n2043_;
  assign new_n1439_ = new_n2042_ | new_n2043_;
  assign new_n1440_ = new_n2045_ | new_n2047_;
  assign new_n1441_ = new_n2048_ | new_n2049_;
  assign new_n1442_ = new_n1440_ & new_n1441_;
  assign new_n1443_ = new_n2045_ | new_n2051_;
  assign new_n1444_ = new_n2048_ | new_n2052_;
  assign new_n1445_ = new_n1443_ & new_n1444_;
  assign new_n1446_ = new_n2051_ | new_n2054_;
  assign new_n1447_ = new_n2052_ | new_n2055_;
  assign new_n1448_ = new_n1446_ & new_n1447_;
  assign new_n1449_ = new_n2057_ | new_n2059_;
  assign new_n1450_ = new_n2060_ | new_n2061_;
  assign new_n1451_ = new_n1449_ & new_n1450_;
  assign new_n1452_ = new_n2057_ & new_n2062_;
  assign new_n1453_ = new_n2060_ & new_n2064_;
  assign new_n1454_ = new_n1452_ | new_n1453_;
  assign new_n1455_ = new_n2064_ | new_n2066_;
  assign new_n1456_ = new_n2062_ | new_n2067_;
  assign new_n1457_ = new_n1455_ & new_n1456_;
  assign new_n1458_ = new_n2047_ | new_n2054_;
  assign new_n1459_ = new_n2049_ | new_n2055_;
  assign new_n1460_ = new_n1458_ & new_n1459_;
  assign new_n1461_ = new_n2059_ & new_n2067_;
  assign new_n1462_ = new_n2061_ & new_n2066_;
  assign new_n1463_ = new_n1461_ | new_n1462_;
  assign new_n1464_ = new_n2069_ & new_n2070_;
  assign new_n1465_ = new_n2071_ & new_n2073_;
  assign new_n1466_ = new_n1464_ | new_n1465_;
  assign new_n1467_ = new_n2069_ | new_n2075_;
  assign new_n1468_ = new_n2071_ | new_n2076_;
  assign new_n1469_ = new_n1467_ & new_n1468_;
  assign new_n1470_ = new_n2075_ & new_n2077_;
  assign new_n1471_ = new_n2076_ & new_n2079_;
  assign new_n1472_ = new_n1470_ | new_n1471_;
  assign new_n1473_ = new_n2081_ & new_n2082_;
  assign new_n1474_ = new_n2083_ & new_n2085_;
  assign new_n1475_ = new_n1473_ | new_n1474_;
  assign new_n1476_ = new_n2081_ & new_n2086_;
  assign new_n1477_ = new_n2083_ & new_n2088_;
  assign new_n1478_ = new_n1476_ | new_n1477_;
  assign new_n1479_ = new_n2088_ & new_n2089_;
  assign new_n1480_ = new_n2086_ & new_n2091_;
  assign new_n1481_ = new_n1479_ | new_n1480_;
  assign new_n1482_ = new_n2073_ | new_n2079_;
  assign new_n1483_ = new_n2070_ | new_n2077_;
  assign new_n1484_ = new_n1482_ & new_n1483_;
  assign new_n1485_ = new_n2085_ & new_n2089_;
  assign new_n1486_ = new_n2082_ & new_n2091_;
  assign new_n1487_ = new_n1485_ | new_n1486_;
  assign new_n1488_ = new_n2093_ | new_n2095_;
  assign new_n1489_ = new_n2096_ | new_n2097_;
  assign new_n1490_ = new_n1488_ & new_n1489_;
  assign new_n1491_ = new_n2093_ | new_n2099_;
  assign new_n1492_ = new_n2096_ | new_n2100_;
  assign new_n1493_ = new_n1491_ & new_n1492_;
  assign new_n1494_ = new_n2095_ | new_n2102_;
  assign new_n1495_ = new_n2097_ | new_n2103_;
  assign new_n1496_ = new_n1494_ & new_n1495_;
  assign new_n1497_ = new_n2105_ & new_n2106_;
  assign new_n1498_ = new_n2107_ & new_n2109_;
  assign new_n1499_ = new_n1497_ | new_n1498_;
  assign new_n1500_ = new_n2105_ | new_n2111_;
  assign new_n1501_ = new_n2107_ | new_n2112_;
  assign new_n1502_ = new_n1500_ & new_n1501_;
  assign new_n1503_ = new_n2109_ | new_n2114_;
  assign new_n1504_ = new_n2106_ | new_n2115_;
  assign new_n1505_ = new_n1503_ & new_n1504_;
  assign new_n1506_ = new_n2099_ | new_n2102_;
  assign new_n1507_ = new_n2100_ | new_n2103_;
  assign new_n1508_ = new_n1506_ & new_n1507_;
  assign new_n1509_ = new_n2111_ & new_n2115_;
  assign new_n1510_ = new_n2112_ & new_n2114_;
  assign new_n1511_ = new_n1509_ | new_n1510_;
  assign new_n1512_ = new_n2117_ | new_n2119_;
  assign new_n1513_ = new_n2120_ | new_n2121_;
  assign new_n1514_ = new_n1512_ & new_n1513_;
  assign new_n1515_ = new_n2117_ & new_n2122_;
  assign new_n1516_ = new_n2120_ & new_n2124_;
  assign new_n1517_ = new_n1515_ | new_n1516_;
  assign new_n1518_ = new_n2119_ & new_n2125_;
  assign new_n1519_ = new_n2121_ & new_n2127_;
  assign new_n1520_ = new_n1518_ | new_n1519_;
  assign new_n1521_ = new_n2129_ & new_n2130_;
  assign new_n1522_ = new_n2131_ & new_n2133_;
  assign new_n1523_ = new_n1521_ | new_n1522_;
  assign new_n1524_ = new_n2129_ & new_n2134_;
  assign new_n1525_ = new_n2131_ & new_n2136_;
  assign new_n1526_ = new_n1524_ | new_n1525_;
  assign new_n1527_ = new_n2133_ & new_n2137_;
  assign new_n1528_ = new_n2130_ & new_n2139_;
  assign new_n1529_ = new_n1527_ | new_n1528_;
  assign new_n1530_ = new_n2124_ | new_n2127_;
  assign new_n1531_ = new_n2122_ | new_n2125_;
  assign new_n1532_ = new_n1530_ & new_n1531_;
  assign new_n1533_ = new_n2136_ & new_n2137_;
  assign new_n1534_ = new_n2134_ & new_n2139_;
  assign new_n1535_ = new_n1533_ | new_n1534_;
  assign G1324 = new_n1038_;
  assign G1325 = new_n1043_;
  assign G1326 = new_n1048_;
  assign G1327 = new_n1053_;
  assign G1328 = new_n1062_;
  assign G1329 = new_n1067_;
  assign G1330 = new_n1072_;
  assign G1331 = new_n1077_;
  assign G1332 = new_n1086_;
  assign G1333 = new_n1091_;
  assign G1334 = new_n1096_;
  assign G1335 = new_n1101_;
  assign G1336 = new_n1110_;
  assign G1337 = new_n1115_;
  assign G1338 = new_n1120_;
  assign G1339 = new_n1125_;
  assign G1340 = new_n1134_;
  assign G1341 = new_n1139_;
  assign G1342 = new_n1144_;
  assign G1343 = new_n1149_;
  assign G1344 = new_n1158_;
  assign G1345 = new_n1163_;
  assign G1346 = new_n1168_;
  assign G1347 = new_n1173_;
  assign G1348 = new_n1182_;
  assign G1349 = new_n1187_;
  assign G1350 = new_n1192_;
  assign G1351 = new_n1197_;
  assign G1352 = new_n1206_;
  assign G1353 = new_n1211_;
  assign G1354 = new_n1216_;
  assign G1355 = new_n1221_;
  assign n1699_li000_li000 = new_n510_;
  assign n1708_li003_li003 = new_n754_;
  assign n1711_li004_li004 = new_n512_;
  assign n1720_li007_li007 = new_n756_;
  assign n1723_li008_li008 = new_n514_;
  assign n1732_li011_li011 = new_n758_;
  assign n1735_li012_li012 = new_n516_;
  assign n1744_li015_li015 = new_n760_;
  assign n1747_li016_li016 = new_n518_;
  assign n1756_li019_li019 = new_n762_;
  assign n1759_li020_li020 = new_n520_;
  assign n1768_li023_li023 = new_n764_;
  assign n1771_li024_li024 = new_n522_;
  assign n1780_li027_li027 = new_n766_;
  assign n1783_li028_li028 = new_n524_;
  assign n1792_li031_li031 = new_n768_;
  assign n1795_li032_li032 = new_n526_;
  assign n1804_li035_li035 = new_n770_;
  assign n1807_li036_li036 = new_n528_;
  assign n1816_li039_li039 = new_n772_;
  assign n1819_li040_li040 = new_n530_;
  assign n1828_li043_li043 = new_n774_;
  assign n1831_li044_li044 = new_n532_;
  assign n1840_li047_li047 = new_n776_;
  assign n1843_li048_li048 = new_n534_;
  assign n1852_li051_li051 = new_n778_;
  assign n1855_li052_li052 = new_n536_;
  assign n1864_li055_li055 = new_n780_;
  assign n1867_li056_li056 = new_n538_;
  assign n1876_li059_li059 = new_n782_;
  assign n1879_li060_li060 = new_n540_;
  assign n1888_li063_li063 = new_n784_;
  assign n1891_li064_li064 = new_n542_;
  assign n1900_li067_li067 = new_n786_;
  assign n1903_li068_li068 = new_n544_;
  assign n1912_li071_li071 = new_n788_;
  assign n1915_li072_li072 = new_n546_;
  assign n1924_li075_li075 = new_n790_;
  assign n1927_li076_li076 = new_n548_;
  assign n1936_li079_li079 = new_n792_;
  assign n1939_li080_li080 = new_n550_;
  assign n1948_li083_li083 = new_n794_;
  assign n1951_li084_li084 = new_n552_;
  assign n1960_li087_li087 = new_n796_;
  assign n1963_li088_li088 = new_n554_;
  assign n1972_li091_li091 = new_n798_;
  assign n1975_li092_li092 = new_n556_;
  assign n1984_li095_li095 = new_n800_;
  assign n1987_li096_li096 = new_n558_;
  assign n1996_li099_li099 = new_n802_;
  assign n1999_li100_li100 = new_n560_;
  assign n2008_li103_li103 = new_n804_;
  assign n2011_li104_li104 = new_n562_;
  assign n2020_li107_li107 = new_n806_;
  assign n2023_li108_li108 = new_n564_;
  assign n2032_li111_li111 = new_n808_;
  assign n2035_li112_li112 = new_n566_;
  assign n2044_li115_li115 = new_n810_;
  assign n2047_li116_li116 = new_n568_;
  assign n2056_li119_li119 = new_n812_;
  assign n2059_li120_li120 = new_n570_;
  assign n2068_li123_li123 = new_n814_;
  assign n2071_li124_li124 = new_n572_;
  assign n2080_li127_li127 = new_n816_;
  assign n2083_li128_li128 = new_n574_;
  assign n2095_li132_li132 = new_n576_;
  assign n2107_li136_li136 = new_n578_;
  assign n2119_li140_li140 = new_n580_;
  assign n2131_li144_li144 = new_n582_;
  assign n2143_li148_li148 = new_n584_;
  assign n2155_li152_li152 = new_n586_;
  assign n2167_li156_li156 = new_n588_;
  assign n2179_li160_li160 = new_n590_;
  assign n602_i2 = new_n1916_;
  assign n639_i2 = new_n1900_;
  assign n678_i2 = new_n1902_;
  assign n658_i2 = new_n1919_;
  assign n783_i2 = new_n1908_;
  assign n802_i2 = new_n1923_;
  assign n726_i2 = new_n1925_;
  assign n763_i2 = new_n1910_;
  assign n1644_i2 = new_n850_;
  assign n1645_i2 = new_n852_;
  assign n1646_i2 = new_n854_;
  assign n1647_i2 = new_n856_;
  assign n1648_i2 = new_n858_;
  assign n1649_i2 = new_n860_;
  assign n1650_i2 = new_n862_;
  assign n1651_i2 = new_n864_;
  assign n1652_i2 = new_n866_;
  assign n1653_i2 = new_n868_;
  assign n1654_i2 = new_n870_;
  assign n1655_i2 = new_n872_;
  assign n1656_i2 = new_n874_;
  assign n1657_i2 = new_n876_;
  assign n1658_i2 = new_n878_;
  assign n1659_i2 = new_n880_;
  assign n1660_i2 = new_n882_;
  assign n1661_i2 = new_n884_;
  assign n1662_i2 = new_n886_;
  assign n1663_i2 = new_n888_;
  assign n1664_i2 = new_n890_;
  assign n1665_i2 = new_n892_;
  assign n1666_i2 = new_n894_;
  assign n1667_i2 = new_n896_;
  assign n1668_i2 = new_n898_;
  assign n1669_i2 = new_n900_;
  assign n1670_i2 = new_n902_;
  assign n1671_i2 = new_n904_;
  assign n1672_i2 = new_n906_;
  assign n1673_i2 = new_n908_;
  assign n1674_i2 = new_n910_;
  assign n1675_i2 = new_n912_;
  assign n685_i2 = ~new_n1922_;
  assign n680_i2 = ~new_n1918_;
  assign n822_i2 = ~new_n1930_;
  assign n843_i2 = new_n1931_;
  assign n842_i2 = ~new_n1933_;
  assign n681_i2 = ~new_n1927_;
  assign n684_i2 = ~new_n1928_;
  assign n686_i2 = ~new_n1929_;
  assign n823_i2 = new_n1932_;
  assign n683_i2 = ~new_n1252_;
  assign n688_i2 = ~new_n1254_;
  assign n803_i2 = new_n1255_;
  assign n862_i2 = new_n1256_;
  assign n764_i2 = new_n1257_;
  assign n863_i2 = new_n1258_;
  assign n886_i2 = new_n1263_;
  assign lo002_buf_i2 = new_n2044_;
  assign lo006_buf_i2 = new_n2050_;
  assign lo010_buf_i2 = new_n2056_;
  assign lo014_buf_i2 = new_n2063_;
  assign lo018_buf_i2 = new_n2046_;
  assign lo022_buf_i2 = new_n2053_;
  assign lo026_buf_i2 = new_n2058_;
  assign lo030_buf_i2 = new_n2065_;
  assign lo034_buf_i2 = new_n2068_;
  assign lo038_buf_i2 = new_n2074_;
  assign lo042_buf_i2 = new_n2080_;
  assign lo046_buf_i2 = new_n2087_;
  assign lo050_buf_i2 = new_n2072_;
  assign lo054_buf_i2 = new_n2078_;
  assign lo058_buf_i2 = new_n2084_;
  assign lo062_buf_i2 = new_n2090_;
  assign lo066_buf_i2 = new_n2092_;
  assign lo070_buf_i2 = new_n2094_;
  assign lo074_buf_i2 = new_n2104_;
  assign lo078_buf_i2 = new_n2108_;
  assign lo082_buf_i2 = new_n2098_;
  assign lo086_buf_i2 = new_n2101_;
  assign lo090_buf_i2 = new_n2110_;
  assign lo094_buf_i2 = new_n2113_;
  assign lo098_buf_i2 = new_n2116_;
  assign lo102_buf_i2 = new_n2118_;
  assign lo106_buf_i2 = new_n2128_;
  assign lo110_buf_i2 = new_n2132_;
  assign lo114_buf_i2 = new_n2123_;
  assign lo118_buf_i2 = new_n2126_;
  assign lo122_buf_i2 = new_n2135_;
  assign lo126_buf_i2 = new_n2138_;
  assign n600_i2 = new_n1290_;
  assign n601_i2 = ~new_n1291_;
  assign n637_i2 = new_n1318_;
  assign n638_i2 = ~new_n1319_;
  assign n676_i2 = new_n1334_;
  assign n677_i2 = ~new_n1335_;
  assign n656_i2 = new_n1350_;
  assign n657_i2 = ~new_n1351_;
  assign n781_i2 = new_n1378_;
  assign n782_i2 = ~new_n1379_;
  assign n800_i2 = new_n1406_;
  assign n801_i2 = ~new_n1407_;
  assign n724_i2 = new_n1422_;
  assign n725_i2 = ~new_n1423_;
  assign n761_i2 = new_n1438_;
  assign n762_i2 = ~new_n1439_;
  assign lo129_buf_i2 = new_n720_;
  assign lo133_buf_i2 = new_n722_;
  assign lo137_buf_i2 = new_n724_;
  assign lo141_buf_i2 = new_n726_;
  assign lo145_buf_i2 = new_n728_;
  assign lo149_buf_i2 = new_n730_;
  assign lo153_buf_i2 = new_n732_;
  assign lo157_buf_i2 = new_n734_;
  assign lo161_buf_i2 = new_n736_;
  assign n571_i2 = new_n1442_;
  assign n708_i2 = new_n1445_;
  assign n608_i2 = new_n1448_;
  assign n665_i2 = new_n1451_;
  assign n705_i2 = new_n1454_;
  assign n645_i2 = new_n1457_;
  assign n745_i2 = new_n1460_;
  assign n742_i2 = new_n1463_;
  assign n568_i2 = new_n1466_;
  assign n717_i2 = new_n1469_;
  assign n605_i2 = new_n1472_;
  assign n662_i2 = new_n1475_;
  assign n714_i2 = new_n1478_;
  assign n642_i2 = new_n1481_;
  assign n754_i2 = new_n1484_;
  assign n751_i2 = new_n1487_;
  assign n584_i2 = new_n1490_;
  assign n770_i2 = new_n1493_;
  assign n789_i2 = new_n1496_;
  assign n581_i2 = new_n1499_;
  assign n695_i2 = new_n1502_;
  assign n732_i2 = new_n1505_;
  assign n593_i2 = new_n1508_;
  assign n590_i2 = new_n1511_;
  assign n630_i2 = new_n1514_;
  assign n767_i2 = new_n1517_;
  assign n786_i2 = new_n1520_;
  assign n627_i2 = new_n1523_;
  assign n692_i2 = new_n1526_;
  assign n729_i2 = new_n1529_;
  assign n621_i2 = new_n1532_;
  assign n618_i2 = new_n1535_;
  assign new_n1786_ = new_n1029_;
  assign new_n1787_ = new_n1786_;
  assign new_n1788_ = new_n1786_;
  assign new_n1789_ = new_n1028_;
  assign new_n1790_ = new_n1789_;
  assign new_n1791_ = new_n1789_;
  assign new_n1792_ = new_n738_;
  assign new_n1793_ = new_n1792_;
  assign new_n1794_ = new_n1792_;
  assign new_n1795_ = new_n1032_;
  assign new_n1796_ = new_n1795_;
  assign new_n1797_ = new_n1795_;
  assign new_n1798_ = new_n739_;
  assign new_n1799_ = new_n1798_;
  assign new_n1800_ = new_n1798_;
  assign new_n1801_ = new_n1033_;
  assign new_n1802_ = new_n1801_;
  assign new_n1803_ = new_n1801_;
  assign new_n1804_ = new_n740_;
  assign new_n1805_ = new_n1804_;
  assign new_n1806_ = new_n1805_;
  assign new_n1807_ = new_n1804_;
  assign new_n1808_ = new_n741_;
  assign new_n1809_ = new_n1808_;
  assign new_n1810_ = new_n1809_;
  assign new_n1811_ = new_n1808_;
  assign new_n1812_ = new_n742_;
  assign new_n1813_ = new_n1812_;
  assign new_n1814_ = new_n1813_;
  assign new_n1815_ = new_n1813_;
  assign new_n1816_ = new_n1812_;
  assign new_n1817_ = new_n743_;
  assign new_n1818_ = new_n1817_;
  assign new_n1819_ = new_n1818_;
  assign new_n1820_ = new_n1818_;
  assign new_n1821_ = new_n1817_;
  assign new_n1822_ = new_n744_;
  assign new_n1823_ = new_n1822_;
  assign new_n1824_ = new_n1822_;
  assign new_n1825_ = new_n745_;
  assign new_n1826_ = new_n1825_;
  assign new_n1827_ = new_n1825_;
  assign new_n1828_ = new_n1056_;
  assign new_n1829_ = new_n1828_;
  assign new_n1830_ = new_n1828_;
  assign new_n1831_ = new_n1057_;
  assign new_n1832_ = new_n1831_;
  assign new_n1833_ = new_n1831_;
  assign new_n1834_ = new_n1080_;
  assign new_n1835_ = new_n1834_;
  assign new_n1836_ = new_n1834_;
  assign new_n1837_ = new_n1081_;
  assign new_n1838_ = new_n1837_;
  assign new_n1839_ = new_n1837_;
  assign new_n1840_ = new_n1104_;
  assign new_n1841_ = new_n1840_;
  assign new_n1842_ = new_n1840_;
  assign new_n1843_ = new_n1105_;
  assign new_n1844_ = new_n1843_;
  assign new_n1845_ = new_n1843_;
  assign new_n1846_ = new_n848_;
  assign new_n1847_ = new_n1846_;
  assign new_n1848_ = new_n1846_;
  assign new_n1849_ = new_n849_;
  assign new_n1850_ = new_n1849_;
  assign new_n1851_ = new_n1849_;
  assign new_n1852_ = new_n746_;
  assign new_n1853_ = new_n1852_;
  assign new_n1854_ = new_n1852_;
  assign new_n1855_ = new_n1128_;
  assign new_n1856_ = new_n1855_;
  assign new_n1857_ = new_n1855_;
  assign new_n1858_ = new_n747_;
  assign new_n1859_ = new_n1858_;
  assign new_n1860_ = new_n1858_;
  assign new_n1861_ = new_n1129_;
  assign new_n1862_ = new_n1861_;
  assign new_n1863_ = new_n1861_;
  assign new_n1864_ = new_n748_;
  assign new_n1865_ = new_n1864_;
  assign new_n1866_ = new_n1864_;
  assign new_n1867_ = new_n749_;
  assign new_n1868_ = new_n1867_;
  assign new_n1869_ = new_n1867_;
  assign new_n1870_ = new_n750_;
  assign new_n1871_ = new_n1870_;
  assign new_n1872_ = new_n1870_;
  assign new_n1873_ = new_n751_;
  assign new_n1874_ = new_n1873_;
  assign new_n1875_ = new_n1873_;
  assign new_n1876_ = new_n752_;
  assign new_n1877_ = new_n1876_;
  assign new_n1878_ = new_n1876_;
  assign new_n1879_ = new_n753_;
  assign new_n1880_ = new_n1879_;
  assign new_n1881_ = new_n1879_;
  assign new_n1882_ = new_n1152_;
  assign new_n1883_ = new_n1882_;
  assign new_n1884_ = new_n1882_;
  assign new_n1885_ = new_n1153_;
  assign new_n1886_ = new_n1885_;
  assign new_n1887_ = new_n1885_;
  assign new_n1888_ = new_n1176_;
  assign new_n1889_ = new_n1888_;
  assign new_n1890_ = new_n1888_;
  assign new_n1891_ = new_n1177_;
  assign new_n1892_ = new_n1891_;
  assign new_n1893_ = new_n1891_;
  assign new_n1894_ = new_n1200_;
  assign new_n1895_ = new_n1894_;
  assign new_n1896_ = new_n1894_;
  assign new_n1897_ = new_n1201_;
  assign new_n1898_ = new_n1897_;
  assign new_n1899_ = new_n1897_;
  assign new_n1900_ = new_n1225_;
  assign new_n1901_ = new_n1900_;
  assign new_n1902_ = new_n1227_;
  assign new_n1903_ = new_n1902_;
  assign new_n1904_ = new_n1230_;
  assign new_n1905_ = new_n1904_;
  assign new_n1906_ = new_n1236_;
  assign new_n1907_ = new_n1906_;
  assign new_n1908_ = new_n1231_;
  assign new_n1909_ = new_n1908_;
  assign new_n1910_ = new_n1237_;
  assign new_n1911_ = new_n1910_;
  assign new_n1912_ = new_n1232_;
  assign new_n1913_ = new_n1912_;
  assign new_n1914_ = new_n1234_;
  assign new_n1915_ = new_n1914_;
  assign new_n1916_ = new_n1223_;
  assign new_n1917_ = new_n1916_;
  assign new_n1918_ = new_n1239_;
  assign new_n1919_ = new_n1229_;
  assign new_n1920_ = new_n1919_;
  assign new_n1921_ = new_n1245_;
  assign new_n1922_ = new_n1238_;
  assign new_n1923_ = new_n1233_;
  assign new_n1924_ = new_n1923_;
  assign new_n1925_ = new_n1235_;
  assign new_n1926_ = new_n1925_;
  assign new_n1927_ = new_n1244_;
  assign new_n1928_ = new_n1246_;
  assign new_n1929_ = new_n1247_;
  assign new_n1930_ = new_n1240_;
  assign new_n1931_ = new_n1242_;
  assign new_n1932_ = new_n1249_;
  assign new_n1933_ = new_n1243_;
  assign new_n1934_ = new_n964_;
  assign new_n1935_ = new_n981_;
  assign new_n1936_ = new_n965_;
  assign new_n1937_ = new_n980_;
  assign new_n1938_ = new_n962_;
  assign new_n1939_ = new_n1938_;
  assign new_n1940_ = new_n1939_;
  assign new_n1941_ = new_n1939_;
  assign new_n1942_ = new_n1938_;
  assign new_n1943_ = new_n1942_;
  assign new_n1944_ = new_n1942_;
  assign new_n1945_ = new_n963_;
  assign new_n1946_ = new_n1945_;
  assign new_n1947_ = new_n1946_;
  assign new_n1948_ = new_n1946_;
  assign new_n1949_ = new_n1945_;
  assign new_n1950_ = new_n1949_;
  assign new_n1951_ = new_n1949_;
  assign new_n1952_ = new_n996_;
  assign new_n1953_ = new_n1003_;
  assign new_n1954_ = new_n997_;
  assign new_n1955_ = new_n1002_;
  assign new_n1956_ = new_n1008_;
  assign new_n1957_ = new_n1011_;
  assign new_n1958_ = new_n1009_;
  assign new_n1959_ = new_n1010_;
  assign new_n1960_ = new_n1279_;
  assign new_n1961_ = new_n1286_;
  assign new_n1962_ = new_n1280_;
  assign new_n1963_ = new_n1285_;
  assign new_n1964_ = new_n1274_;
  assign new_n1965_ = new_n1289_;
  assign new_n1966_ = new_n968_;
  assign new_n1967_ = new_n985_;
  assign new_n1968_ = new_n969_;
  assign new_n1969_ = new_n984_;
  assign new_n1970_ = new_n1024_;
  assign new_n1971_ = new_n1027_;
  assign new_n1972_ = new_n1025_;
  assign new_n1973_ = new_n1026_;
  assign new_n1974_ = new_n1012_;
  assign new_n1975_ = new_n1019_;
  assign new_n1976_ = new_n1013_;
  assign new_n1977_ = new_n1018_;
  assign new_n1978_ = new_n1307_;
  assign new_n1979_ = new_n1314_;
  assign new_n1980_ = new_n1308_;
  assign new_n1981_ = new_n1313_;
  assign new_n1982_ = new_n1302_;
  assign new_n1983_ = new_n1317_;
  assign new_n1984_ = new_n970_;
  assign new_n1985_ = new_n987_;
  assign new_n1986_ = new_n971_;
  assign new_n1987_ = new_n986_;
  assign new_n1988_ = new_n1330_;
  assign new_n1989_ = new_n1333_;
  assign new_n1990_ = new_n974_;
  assign new_n1991_ = new_n991_;
  assign new_n1992_ = new_n975_;
  assign new_n1993_ = new_n990_;
  assign new_n1994_ = new_n1346_;
  assign new_n1995_ = new_n1349_;
  assign new_n1996_ = new_n998_;
  assign new_n1997_ = new_n1015_;
  assign new_n1998_ = new_n999_;
  assign new_n1999_ = new_n1014_;
  assign new_n2000_ = new_n966_;
  assign new_n2001_ = new_n973_;
  assign new_n2002_ = new_n967_;
  assign new_n2003_ = new_n972_;
  assign new_n2004_ = new_n976_;
  assign new_n2005_ = new_n979_;
  assign new_n2006_ = new_n977_;
  assign new_n2007_ = new_n978_;
  assign new_n2008_ = new_n1367_;
  assign new_n2009_ = new_n1374_;
  assign new_n2010_ = new_n1368_;
  assign new_n2011_ = new_n1373_;
  assign new_n2012_ = new_n1362_;
  assign new_n2013_ = new_n1377_;
  assign new_n2014_ = new_n1000_;
  assign new_n2015_ = new_n1017_;
  assign new_n2016_ = new_n1001_;
  assign new_n2017_ = new_n1016_;
  assign new_n2018_ = new_n982_;
  assign new_n2019_ = new_n989_;
  assign new_n2020_ = new_n983_;
  assign new_n2021_ = new_n988_;
  assign new_n2022_ = new_n992_;
  assign new_n2023_ = new_n995_;
  assign new_n2024_ = new_n993_;
  assign new_n2025_ = new_n994_;
  assign new_n2026_ = new_n1395_;
  assign new_n2027_ = new_n1402_;
  assign new_n2028_ = new_n1396_;
  assign new_n2029_ = new_n1401_;
  assign new_n2030_ = new_n1390_;
  assign new_n2031_ = new_n1405_;
  assign new_n2032_ = new_n1004_;
  assign new_n2033_ = new_n1021_;
  assign new_n2034_ = new_n1005_;
  assign new_n2035_ = new_n1020_;
  assign new_n2036_ = new_n1418_;
  assign new_n2037_ = new_n1421_;
  assign new_n2038_ = new_n1006_;
  assign new_n2039_ = new_n1023_;
  assign new_n2040_ = new_n1007_;
  assign new_n2041_ = new_n1022_;
  assign new_n2042_ = new_n1434_;
  assign new_n2043_ = new_n1437_;
  assign new_n2044_ = new_n592_;
  assign new_n2045_ = new_n2044_;
  assign new_n2046_ = new_n608_;
  assign new_n2047_ = new_n2046_;
  assign new_n2048_ = new_n593_;
  assign new_n2049_ = new_n609_;
  assign new_n2050_ = new_n596_;
  assign new_n2051_ = new_n2050_;
  assign new_n2052_ = new_n597_;
  assign new_n2053_ = new_n612_;
  assign new_n2054_ = new_n2053_;
  assign new_n2055_ = new_n613_;
  assign new_n2056_ = new_n600_;
  assign new_n2057_ = new_n2056_;
  assign new_n2058_ = new_n616_;
  assign new_n2059_ = new_n2058_;
  assign new_n2060_ = new_n601_;
  assign new_n2061_ = new_n617_;
  assign new_n2062_ = new_n605_;
  assign new_n2063_ = new_n604_;
  assign new_n2064_ = new_n2063_;
  assign new_n2065_ = new_n620_;
  assign new_n2066_ = new_n2065_;
  assign new_n2067_ = new_n621_;
  assign new_n2068_ = new_n624_;
  assign new_n2069_ = new_n2068_;
  assign new_n2070_ = new_n641_;
  assign new_n2071_ = new_n625_;
  assign new_n2072_ = new_n640_;
  assign new_n2073_ = new_n2072_;
  assign new_n2074_ = new_n628_;
  assign new_n2075_ = new_n2074_;
  assign new_n2076_ = new_n629_;
  assign new_n2077_ = new_n645_;
  assign new_n2078_ = new_n644_;
  assign new_n2079_ = new_n2078_;
  assign new_n2080_ = new_n632_;
  assign new_n2081_ = new_n2080_;
  assign new_n2082_ = new_n649_;
  assign new_n2083_ = new_n633_;
  assign new_n2084_ = new_n648_;
  assign new_n2085_ = new_n2084_;
  assign new_n2086_ = new_n637_;
  assign new_n2087_ = new_n636_;
  assign new_n2088_ = new_n2087_;
  assign new_n2089_ = new_n653_;
  assign new_n2090_ = new_n652_;
  assign new_n2091_ = new_n2090_;
  assign new_n2092_ = new_n656_;
  assign new_n2093_ = new_n2092_;
  assign new_n2094_ = new_n660_;
  assign new_n2095_ = new_n2094_;
  assign new_n2096_ = new_n657_;
  assign new_n2097_ = new_n661_;
  assign new_n2098_ = new_n672_;
  assign new_n2099_ = new_n2098_;
  assign new_n2100_ = new_n673_;
  assign new_n2101_ = new_n676_;
  assign new_n2102_ = new_n2101_;
  assign new_n2103_ = new_n677_;
  assign new_n2104_ = new_n664_;
  assign new_n2105_ = new_n2104_;
  assign new_n2106_ = new_n669_;
  assign new_n2107_ = new_n665_;
  assign new_n2108_ = new_n668_;
  assign new_n2109_ = new_n2108_;
  assign new_n2110_ = new_n680_;
  assign new_n2111_ = new_n2110_;
  assign new_n2112_ = new_n681_;
  assign new_n2113_ = new_n684_;
  assign new_n2114_ = new_n2113_;
  assign new_n2115_ = new_n685_;
  assign new_n2116_ = new_n688_;
  assign new_n2117_ = new_n2116_;
  assign new_n2118_ = new_n692_;
  assign new_n2119_ = new_n2118_;
  assign new_n2120_ = new_n689_;
  assign new_n2121_ = new_n693_;
  assign new_n2122_ = new_n705_;
  assign new_n2123_ = new_n704_;
  assign new_n2124_ = new_n2123_;
  assign new_n2125_ = new_n709_;
  assign new_n2126_ = new_n708_;
  assign new_n2127_ = new_n2126_;
  assign new_n2128_ = new_n696_;
  assign new_n2129_ = new_n2128_;
  assign new_n2130_ = new_n701_;
  assign new_n2131_ = new_n697_;
  assign new_n2132_ = new_n700_;
  assign new_n2133_ = new_n2132_;
  assign new_n2134_ = new_n713_;
  assign new_n2135_ = new_n712_;
  assign new_n2136_ = new_n2135_;
  assign new_n2137_ = new_n717_;
  assign new_n2138_ = new_n716_;
  assign new_n2139_ = new_n2138_;
  always @ (posedge clock) begin
    n621_lo <= n1699_li000_li000;
    n630_lo <= n1708_li003_li003;
    n633_lo <= n1711_li004_li004;
    n642_lo <= n1720_li007_li007;
    n645_lo <= n1723_li008_li008;
    n654_lo <= n1732_li011_li011;
    n657_lo <= n1735_li012_li012;
    n666_lo <= n1744_li015_li015;
    n669_lo <= n1747_li016_li016;
    n678_lo <= n1756_li019_li019;
    n681_lo <= n1759_li020_li020;
    n690_lo <= n1768_li023_li023;
    n693_lo <= n1771_li024_li024;
    n702_lo <= n1780_li027_li027;
    n705_lo <= n1783_li028_li028;
    n714_lo <= n1792_li031_li031;
    n717_lo <= n1795_li032_li032;
    n726_lo <= n1804_li035_li035;
    n729_lo <= n1807_li036_li036;
    n738_lo <= n1816_li039_li039;
    n741_lo <= n1819_li040_li040;
    n750_lo <= n1828_li043_li043;
    n753_lo <= n1831_li044_li044;
    n762_lo <= n1840_li047_li047;
    n765_lo <= n1843_li048_li048;
    n774_lo <= n1852_li051_li051;
    n777_lo <= n1855_li052_li052;
    n786_lo <= n1864_li055_li055;
    n789_lo <= n1867_li056_li056;
    n798_lo <= n1876_li059_li059;
    n801_lo <= n1879_li060_li060;
    n810_lo <= n1888_li063_li063;
    n813_lo <= n1891_li064_li064;
    n822_lo <= n1900_li067_li067;
    n825_lo <= n1903_li068_li068;
    n834_lo <= n1912_li071_li071;
    n837_lo <= n1915_li072_li072;
    n846_lo <= n1924_li075_li075;
    n849_lo <= n1927_li076_li076;
    n858_lo <= n1936_li079_li079;
    n861_lo <= n1939_li080_li080;
    n870_lo <= n1948_li083_li083;
    n873_lo <= n1951_li084_li084;
    n882_lo <= n1960_li087_li087;
    n885_lo <= n1963_li088_li088;
    n894_lo <= n1972_li091_li091;
    n897_lo <= n1975_li092_li092;
    n906_lo <= n1984_li095_li095;
    n909_lo <= n1987_li096_li096;
    n918_lo <= n1996_li099_li099;
    n921_lo <= n1999_li100_li100;
    n930_lo <= n2008_li103_li103;
    n933_lo <= n2011_li104_li104;
    n942_lo <= n2020_li107_li107;
    n945_lo <= n2023_li108_li108;
    n954_lo <= n2032_li111_li111;
    n957_lo <= n2035_li112_li112;
    n966_lo <= n2044_li115_li115;
    n969_lo <= n2047_li116_li116;
    n978_lo <= n2056_li119_li119;
    n981_lo <= n2059_li120_li120;
    n990_lo <= n2068_li123_li123;
    n993_lo <= n2071_li124_li124;
    n1002_lo <= n2080_li127_li127;
    n1005_lo <= n2083_li128_li128;
    n1017_lo <= n2095_li132_li132;
    n1029_lo <= n2107_li136_li136;
    n1041_lo <= n2119_li140_li140;
    n1053_lo <= n2131_li144_li144;
    n1065_lo <= n2143_li148_li148;
    n1077_lo <= n2155_li152_li152;
    n1089_lo <= n2167_li156_li156;
    n1101_lo <= n2179_li160_li160;
    n602_o2 <= n602_i2;
    n639_o2 <= n639_i2;
    n678_o2 <= n678_i2;
    n658_o2 <= n658_i2;
    n783_o2 <= n783_i2;
    n802_o2 <= n802_i2;
    n726_o2 <= n726_i2;
    n763_o2 <= n763_i2;
    n1644_o2 <= n1644_i2;
    n1645_o2 <= n1645_i2;
    n1646_o2 <= n1646_i2;
    n1647_o2 <= n1647_i2;
    n1648_o2 <= n1648_i2;
    n1649_o2 <= n1649_i2;
    n1650_o2 <= n1650_i2;
    n1651_o2 <= n1651_i2;
    n1652_o2 <= n1652_i2;
    n1653_o2 <= n1653_i2;
    n1654_o2 <= n1654_i2;
    n1655_o2 <= n1655_i2;
    n1656_o2 <= n1656_i2;
    n1657_o2 <= n1657_i2;
    n1658_o2 <= n1658_i2;
    n1659_o2 <= n1659_i2;
    n1660_o2 <= n1660_i2;
    n1661_o2 <= n1661_i2;
    n1662_o2 <= n1662_i2;
    n1663_o2 <= n1663_i2;
    n1664_o2 <= n1664_i2;
    n1665_o2 <= n1665_i2;
    n1666_o2 <= n1666_i2;
    n1667_o2 <= n1667_i2;
    n1668_o2 <= n1668_i2;
    n1669_o2 <= n1669_i2;
    n1670_o2 <= n1670_i2;
    n1671_o2 <= n1671_i2;
    n1672_o2 <= n1672_i2;
    n1673_o2 <= n1673_i2;
    n1674_o2 <= n1674_i2;
    n1675_o2 <= n1675_i2;
    n685_o2 <= n685_i2;
    n680_o2 <= n680_i2;
    n822_o2 <= n822_i2;
    n843_o2 <= n843_i2;
    n842_o2 <= n842_i2;
    n681_o2 <= n681_i2;
    n684_o2 <= n684_i2;
    n686_o2 <= n686_i2;
    n823_o2 <= n823_i2;
    n683_o2 <= n683_i2;
    n688_o2 <= n688_i2;
    n803_o2 <= n803_i2;
    n862_o2 <= n862_i2;
    n764_o2 <= n764_i2;
    n863_o2 <= n863_i2;
    n886_o2 <= n886_i2;
    lo002_buf_o2 <= lo002_buf_i2;
    lo006_buf_o2 <= lo006_buf_i2;
    lo010_buf_o2 <= lo010_buf_i2;
    lo014_buf_o2 <= lo014_buf_i2;
    lo018_buf_o2 <= lo018_buf_i2;
    lo022_buf_o2 <= lo022_buf_i2;
    lo026_buf_o2 <= lo026_buf_i2;
    lo030_buf_o2 <= lo030_buf_i2;
    lo034_buf_o2 <= lo034_buf_i2;
    lo038_buf_o2 <= lo038_buf_i2;
    lo042_buf_o2 <= lo042_buf_i2;
    lo046_buf_o2 <= lo046_buf_i2;
    lo050_buf_o2 <= lo050_buf_i2;
    lo054_buf_o2 <= lo054_buf_i2;
    lo058_buf_o2 <= lo058_buf_i2;
    lo062_buf_o2 <= lo062_buf_i2;
    lo066_buf_o2 <= lo066_buf_i2;
    lo070_buf_o2 <= lo070_buf_i2;
    lo074_buf_o2 <= lo074_buf_i2;
    lo078_buf_o2 <= lo078_buf_i2;
    lo082_buf_o2 <= lo082_buf_i2;
    lo086_buf_o2 <= lo086_buf_i2;
    lo090_buf_o2 <= lo090_buf_i2;
    lo094_buf_o2 <= lo094_buf_i2;
    lo098_buf_o2 <= lo098_buf_i2;
    lo102_buf_o2 <= lo102_buf_i2;
    lo106_buf_o2 <= lo106_buf_i2;
    lo110_buf_o2 <= lo110_buf_i2;
    lo114_buf_o2 <= lo114_buf_i2;
    lo118_buf_o2 <= lo118_buf_i2;
    lo122_buf_o2 <= lo122_buf_i2;
    lo126_buf_o2 <= lo126_buf_i2;
    n600_o2 <= n600_i2;
    n601_o2 <= n601_i2;
    n637_o2 <= n637_i2;
    n638_o2 <= n638_i2;
    n676_o2 <= n676_i2;
    n677_o2 <= n677_i2;
    n656_o2 <= n656_i2;
    n657_o2 <= n657_i2;
    n781_o2 <= n781_i2;
    n782_o2 <= n782_i2;
    n800_o2 <= n800_i2;
    n801_o2 <= n801_i2;
    n724_o2 <= n724_i2;
    n725_o2 <= n725_i2;
    n761_o2 <= n761_i2;
    n762_o2 <= n762_i2;
    lo129_buf_o2 <= lo129_buf_i2;
    lo133_buf_o2 <= lo133_buf_i2;
    lo137_buf_o2 <= lo137_buf_i2;
    lo141_buf_o2 <= lo141_buf_i2;
    lo145_buf_o2 <= lo145_buf_i2;
    lo149_buf_o2 <= lo149_buf_i2;
    lo153_buf_o2 <= lo153_buf_i2;
    lo157_buf_o2 <= lo157_buf_i2;
    lo161_buf_o2 <= lo161_buf_i2;
    n571_o2 <= n571_i2;
    n708_o2 <= n708_i2;
    n608_o2 <= n608_i2;
    n665_o2 <= n665_i2;
    n705_o2 <= n705_i2;
    n645_o2 <= n645_i2;
    n745_o2 <= n745_i2;
    n742_o2 <= n742_i2;
    n568_o2 <= n568_i2;
    n717_o2 <= n717_i2;
    n605_o2 <= n605_i2;
    n662_o2 <= n662_i2;
    n714_o2 <= n714_i2;
    n642_o2 <= n642_i2;
    n754_o2 <= n754_i2;
    n751_o2 <= n751_i2;
    n584_o2 <= n584_i2;
    n770_o2 <= n770_i2;
    n789_o2 <= n789_i2;
    n581_o2 <= n581_i2;
    n695_o2 <= n695_i2;
    n732_o2 <= n732_i2;
    n593_o2 <= n593_i2;
    n590_o2 <= n590_i2;
    n630_o2 <= n630_i2;
    n767_o2 <= n767_i2;
    n786_o2 <= n786_i2;
    n627_o2 <= n627_i2;
    n692_o2 <= n692_i2;
    n729_o2 <= n729_i2;
    n621_o2 <= n621_i2;
    n618_o2 <= n618_i2;
  end
  initial begin
    n621_lo <= 1'b0;
    n630_lo <= 1'b0;
    n633_lo <= 1'b0;
    n642_lo <= 1'b0;
    n645_lo <= 1'b0;
    n654_lo <= 1'b0;
    n657_lo <= 1'b0;
    n666_lo <= 1'b0;
    n669_lo <= 1'b0;
    n678_lo <= 1'b0;
    n681_lo <= 1'b0;
    n690_lo <= 1'b0;
    n693_lo <= 1'b0;
    n702_lo <= 1'b0;
    n705_lo <= 1'b0;
    n714_lo <= 1'b0;
    n717_lo <= 1'b0;
    n726_lo <= 1'b0;
    n729_lo <= 1'b0;
    n738_lo <= 1'b0;
    n741_lo <= 1'b0;
    n750_lo <= 1'b0;
    n753_lo <= 1'b0;
    n762_lo <= 1'b0;
    n765_lo <= 1'b0;
    n774_lo <= 1'b0;
    n777_lo <= 1'b0;
    n786_lo <= 1'b0;
    n789_lo <= 1'b0;
    n798_lo <= 1'b0;
    n801_lo <= 1'b0;
    n810_lo <= 1'b0;
    n813_lo <= 1'b0;
    n822_lo <= 1'b0;
    n825_lo <= 1'b0;
    n834_lo <= 1'b0;
    n837_lo <= 1'b0;
    n846_lo <= 1'b0;
    n849_lo <= 1'b0;
    n858_lo <= 1'b0;
    n861_lo <= 1'b0;
    n870_lo <= 1'b0;
    n873_lo <= 1'b0;
    n882_lo <= 1'b0;
    n885_lo <= 1'b0;
    n894_lo <= 1'b0;
    n897_lo <= 1'b0;
    n906_lo <= 1'b0;
    n909_lo <= 1'b0;
    n918_lo <= 1'b0;
    n921_lo <= 1'b0;
    n930_lo <= 1'b0;
    n933_lo <= 1'b0;
    n942_lo <= 1'b0;
    n945_lo <= 1'b0;
    n954_lo <= 1'b0;
    n957_lo <= 1'b0;
    n966_lo <= 1'b0;
    n969_lo <= 1'b0;
    n978_lo <= 1'b0;
    n981_lo <= 1'b0;
    n990_lo <= 1'b0;
    n993_lo <= 1'b0;
    n1002_lo <= 1'b0;
    n1005_lo <= 1'b0;
    n1017_lo <= 1'b0;
    n1029_lo <= 1'b0;
    n1041_lo <= 1'b0;
    n1053_lo <= 1'b0;
    n1065_lo <= 1'b0;
    n1077_lo <= 1'b0;
    n1089_lo <= 1'b0;
    n1101_lo <= 1'b0;
    n602_o2 <= 1'b0;
    n639_o2 <= 1'b0;
    n678_o2 <= 1'b0;
    n658_o2 <= 1'b0;
    n783_o2 <= 1'b0;
    n802_o2 <= 1'b0;
    n726_o2 <= 1'b0;
    n763_o2 <= 1'b0;
    n1644_o2 <= 1'b0;
    n1645_o2 <= 1'b0;
    n1646_o2 <= 1'b0;
    n1647_o2 <= 1'b0;
    n1648_o2 <= 1'b0;
    n1649_o2 <= 1'b0;
    n1650_o2 <= 1'b0;
    n1651_o2 <= 1'b0;
    n1652_o2 <= 1'b0;
    n1653_o2 <= 1'b0;
    n1654_o2 <= 1'b0;
    n1655_o2 <= 1'b0;
    n1656_o2 <= 1'b0;
    n1657_o2 <= 1'b0;
    n1658_o2 <= 1'b0;
    n1659_o2 <= 1'b0;
    n1660_o2 <= 1'b0;
    n1661_o2 <= 1'b0;
    n1662_o2 <= 1'b0;
    n1663_o2 <= 1'b0;
    n1664_o2 <= 1'b0;
    n1665_o2 <= 1'b0;
    n1666_o2 <= 1'b0;
    n1667_o2 <= 1'b0;
    n1668_o2 <= 1'b0;
    n1669_o2 <= 1'b0;
    n1670_o2 <= 1'b0;
    n1671_o2 <= 1'b0;
    n1672_o2 <= 1'b0;
    n1673_o2 <= 1'b0;
    n1674_o2 <= 1'b0;
    n1675_o2 <= 1'b0;
    n685_o2 <= 1'b0;
    n680_o2 <= 1'b0;
    n822_o2 <= 1'b0;
    n843_o2 <= 1'b0;
    n842_o2 <= 1'b0;
    n681_o2 <= 1'b0;
    n684_o2 <= 1'b0;
    n686_o2 <= 1'b0;
    n823_o2 <= 1'b0;
    n683_o2 <= 1'b0;
    n688_o2 <= 1'b0;
    n803_o2 <= 1'b0;
    n862_o2 <= 1'b0;
    n764_o2 <= 1'b0;
    n863_o2 <= 1'b0;
    n886_o2 <= 1'b0;
    lo002_buf_o2 <= 1'b0;
    lo006_buf_o2 <= 1'b0;
    lo010_buf_o2 <= 1'b0;
    lo014_buf_o2 <= 1'b0;
    lo018_buf_o2 <= 1'b0;
    lo022_buf_o2 <= 1'b0;
    lo026_buf_o2 <= 1'b0;
    lo030_buf_o2 <= 1'b0;
    lo034_buf_o2 <= 1'b0;
    lo038_buf_o2 <= 1'b0;
    lo042_buf_o2 <= 1'b0;
    lo046_buf_o2 <= 1'b0;
    lo050_buf_o2 <= 1'b0;
    lo054_buf_o2 <= 1'b0;
    lo058_buf_o2 <= 1'b0;
    lo062_buf_o2 <= 1'b0;
    lo066_buf_o2 <= 1'b0;
    lo070_buf_o2 <= 1'b0;
    lo074_buf_o2 <= 1'b0;
    lo078_buf_o2 <= 1'b0;
    lo082_buf_o2 <= 1'b0;
    lo086_buf_o2 <= 1'b0;
    lo090_buf_o2 <= 1'b0;
    lo094_buf_o2 <= 1'b0;
    lo098_buf_o2 <= 1'b0;
    lo102_buf_o2 <= 1'b0;
    lo106_buf_o2 <= 1'b0;
    lo110_buf_o2 <= 1'b0;
    lo114_buf_o2 <= 1'b0;
    lo118_buf_o2 <= 1'b0;
    lo122_buf_o2 <= 1'b0;
    lo126_buf_o2 <= 1'b0;
    n600_o2 <= 1'b0;
    n601_o2 <= 1'b0;
    n637_o2 <= 1'b0;
    n638_o2 <= 1'b0;
    n676_o2 <= 1'b0;
    n677_o2 <= 1'b0;
    n656_o2 <= 1'b0;
    n657_o2 <= 1'b0;
    n781_o2 <= 1'b0;
    n782_o2 <= 1'b0;
    n800_o2 <= 1'b0;
    n801_o2 <= 1'b0;
    n724_o2 <= 1'b0;
    n725_o2 <= 1'b0;
    n761_o2 <= 1'b0;
    n762_o2 <= 1'b0;
    lo129_buf_o2 <= 1'b0;
    lo133_buf_o2 <= 1'b0;
    lo137_buf_o2 <= 1'b0;
    lo141_buf_o2 <= 1'b0;
    lo145_buf_o2 <= 1'b0;
    lo149_buf_o2 <= 1'b0;
    lo153_buf_o2 <= 1'b0;
    lo157_buf_o2 <= 1'b0;
    lo161_buf_o2 <= 1'b0;
    n571_o2 <= 1'b0;
    n708_o2 <= 1'b0;
    n608_o2 <= 1'b0;
    n665_o2 <= 1'b0;
    n705_o2 <= 1'b0;
    n645_o2 <= 1'b0;
    n745_o2 <= 1'b0;
    n742_o2 <= 1'b0;
    n568_o2 <= 1'b0;
    n717_o2 <= 1'b0;
    n605_o2 <= 1'b0;
    n662_o2 <= 1'b0;
    n714_o2 <= 1'b0;
    n642_o2 <= 1'b0;
    n754_o2 <= 1'b0;
    n751_o2 <= 1'b0;
    n584_o2 <= 1'b0;
    n770_o2 <= 1'b0;
    n789_o2 <= 1'b0;
    n581_o2 <= 1'b0;
    n695_o2 <= 1'b0;
    n732_o2 <= 1'b0;
    n593_o2 <= 1'b0;
    n590_o2 <= 1'b0;
    n630_o2 <= 1'b0;
    n767_o2 <= 1'b0;
    n786_o2 <= 1'b0;
    n627_o2 <= 1'b0;
    n692_o2 <= 1'b0;
    n729_o2 <= 1'b0;
    n621_o2 <= 1'b0;
    n618_o2 <= 1'b0;
  end
endmodule


