
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  n205_lo,
  n214_lo,
  n217_lo,
  n226_lo,
  n229_lo,
  n232_lo,
  n238_lo,
  n241_lo,
  n250_lo,
  n253_lo,
  n256_lo,
  n262_lo,
  n265_lo,
  n274_lo,
  n277_lo,
  n280_lo,
  n286_lo,
  n289_lo,
  n298_lo,
  n301_lo,
  n304_lo,
  n310_lo,
  n313_lo,
  n322_lo,
  n325_lo,
  n328_lo,
  n334_lo,
  n337_lo,
  n346_lo,
  n349_lo,
  n352_lo,
  n358_lo,
  n361_lo,
  n370_lo,
  n373_lo,
  n376_lo,
  n382_lo,
  n385_lo,
  n394_lo,
  n397_lo,
  n400_lo,
  n406_lo,
  n409_lo,
  n418_lo,
  n421_lo,
  n424_lo,
  n430_lo,
  n433_lo,
  n442_lo,
  n445_lo,
  n448_lo,
  n454_lo,
  n457_lo,
  n466_lo,
  n469_lo,
  n472_lo,
  n478_lo,
  n481_lo,
  n490_lo,
  n493_lo,
  n496_lo,
  n502_lo,
  n505_lo,
  n514_lo,
  n517_lo,
  n520_lo,
  n526_lo,
  n529_lo,
  n538_lo,
  n541_lo,
  n544_lo,
  n550_lo,
  n553_lo,
  n562_lo,
  n565_lo,
  n568_lo,
  n574_lo,
  n577_lo,
  n586_lo,
  n589_lo,
  n592_lo,
  n598_lo,
  n601_lo,
  n610_lo,
  n613_lo,
  n616_lo,
  n622_lo,
  n625_lo,
  n628_lo,
  n634_lo,
  n316_inv,
  n319_inv,
  n997_o2,
  n998_o2,
  n999_o2,
  n1000_o2,
  n1001_o2,
  n1002_o2,
  n1003_o2,
  n1004_o2,
  n1005_o2,
  n1015_o2,
  n1016_o2,
  n1017_o2,
  n1018_o2,
  n1019_o2,
  n1020_o2,
  n1021_o2,
  n1022_o2,
  n1023_o2,
  n376_1_inv,
  n235_lo_buf_o2,
  n283_lo_buf_o2,
  n331_lo_buf_o2,
  n379_lo_buf_o2,
  n427_lo_buf_o2,
  n475_lo_buf_o2,
  n523_lo_buf_o2,
  n571_lo_buf_o2,
  n619_lo_buf_o2,
  n406_1_inv,
  G223_o2,
  G226_o2,
  G229_o2,
  G232_o2,
  G235_o2,
  G238_o2,
  G242_o2,
  G246_o2,
  G250_o2,
  n259_lo_buf_o2,
  n307_lo_buf_o2,
  n355_lo_buf_o2,
  n403_lo_buf_o2,
  n451_lo_buf_o2,
  n499_lo_buf_o2,
  n547_lo_buf_o2,
  n595_lo_buf_o2,
  n631_lo_buf_o2,
  G213_o2,
  G318_o2,
  G358_o2,
  G259_o2,
  G263_o2,
  G266_o2,
  G269_o2,
  G272_o2,
  G275_o2,
  G278_o2,
  G281_o2,
  G284_o2,
  n211_lo_buf_o2,
  n247_lo_buf_o2,
  n295_lo_buf_o2,
  n343_lo_buf_o2,
  n391_lo_buf_o2,
  n439_lo_buf_o2,
  n487_lo_buf_o2,
  n535_lo_buf_o2,
  n583_lo_buf_o2,
  G158_o2,
  G184_o2,
  G186_o2,
  G188_o2,
  G190_o2,
  G192_o2,
  G194_o2,
  G196_o2,
  G198_o2,
  n223_lo_buf_o2,
  n271_lo_buf_o2,
  n319_lo_buf_o2,
  n367_lo_buf_o2,
  n415_lo_buf_o2,
  n463_lo_buf_o2,
  n511_lo_buf_o2,
  n559_lo_buf_o2,
  n607_lo_buf_o2,
  n580_inv,
  G154_o2,
  G159_o2,
  G162_o2,
  G165_o2,
  G168_o2,
  G171_o2,
  G174_o2,
  G177_o2,
  G180_o2,
  G426,
  G427,
  G428,
  G429,
  G430,
  G431,
  G432,
  n205_li,
  n214_li,
  n217_li,
  n226_li,
  n229_li,
  n232_li,
  n238_li,
  n241_li,
  n250_li,
  n253_li,
  n256_li,
  n262_li,
  n265_li,
  n274_li,
  n277_li,
  n280_li,
  n286_li,
  n289_li,
  n298_li,
  n301_li,
  n304_li,
  n310_li,
  n313_li,
  n322_li,
  n325_li,
  n328_li,
  n334_li,
  n337_li,
  n346_li,
  n349_li,
  n352_li,
  n358_li,
  n361_li,
  n370_li,
  n373_li,
  n376_li,
  n382_li,
  n385_li,
  n394_li,
  n397_li,
  n400_li,
  n406_li,
  n409_li,
  n418_li,
  n421_li,
  n424_li,
  n430_li,
  n433_li,
  n442_li,
  n445_li,
  n448_li,
  n454_li,
  n457_li,
  n466_li,
  n469_li,
  n472_li,
  n478_li,
  n481_li,
  n490_li,
  n493_li,
  n496_li,
  n502_li,
  n505_li,
  n514_li,
  n517_li,
  n520_li,
  n526_li,
  n529_li,
  n538_li,
  n541_li,
  n544_li,
  n550_li,
  n553_li,
  n562_li,
  n565_li,
  n568_li,
  n574_li,
  n577_li,
  n586_li,
  n589_li,
  n592_li,
  n598_li,
  n601_li,
  n610_li,
  n613_li,
  n616_li,
  n622_li,
  n625_li,
  n628_li,
  n634_li,
  n919_i2,
  n1024_i2,
  n997_i2,
  n998_i2,
  n999_i2,
  n1000_i2,
  n1001_i2,
  n1002_i2,
  n1003_i2,
  n1004_i2,
  n1005_i2,
  n1015_i2,
  n1016_i2,
  n1017_i2,
  n1018_i2,
  n1019_i2,
  n1020_i2,
  n1021_i2,
  n1022_i2,
  n1023_i2,
  G199_i2,
  n235_lo_buf_i2,
  n283_lo_buf_i2,
  n331_lo_buf_i2,
  n379_lo_buf_i2,
  n427_lo_buf_i2,
  n475_lo_buf_i2,
  n523_lo_buf_i2,
  n571_lo_buf_i2,
  n619_lo_buf_i2,
  G355_i2,
  G223_i2,
  G226_i2,
  G229_i2,
  G232_i2,
  G235_i2,
  G238_i2,
  G242_i2,
  G246_i2,
  G250_i2,
  n259_lo_buf_i2,
  n307_lo_buf_i2,
  n355_lo_buf_i2,
  n403_lo_buf_i2,
  n451_lo_buf_i2,
  n499_lo_buf_i2,
  n547_lo_buf_i2,
  n595_lo_buf_i2,
  n631_lo_buf_i2,
  G213_i2,
  G318_i2,
  G358_i2,
  G259_i2,
  G263_i2,
  G266_i2,
  G269_i2,
  G272_i2,
  G275_i2,
  G278_i2,
  G281_i2,
  G284_i2,
  n211_lo_buf_i2,
  n247_lo_buf_i2,
  n295_lo_buf_i2,
  n343_lo_buf_i2,
  n391_lo_buf_i2,
  n439_lo_buf_i2,
  n487_lo_buf_i2,
  n535_lo_buf_i2,
  n583_lo_buf_i2,
  G158_i2,
  G184_i2,
  G186_i2,
  G188_i2,
  G190_i2,
  G192_i2,
  G194_i2,
  G196_i2,
  G198_i2,
  n223_lo_buf_i2,
  n271_lo_buf_i2,
  n319_lo_buf_i2,
  n367_lo_buf_i2,
  n415_lo_buf_i2,
  n463_lo_buf_i2,
  n511_lo_buf_i2,
  n559_lo_buf_i2,
  n607_lo_buf_i2,
  G295_i2,
  G154_i2,
  G159_i2,
  G162_i2,
  G165_i2,
  G168_i2,
  G171_i2,
  G174_i2,
  G177_i2,
  G180_i2
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input n205_lo;input n214_lo;input n217_lo;input n226_lo;input n229_lo;input n232_lo;input n238_lo;input n241_lo;input n250_lo;input n253_lo;input n256_lo;input n262_lo;input n265_lo;input n274_lo;input n277_lo;input n280_lo;input n286_lo;input n289_lo;input n298_lo;input n301_lo;input n304_lo;input n310_lo;input n313_lo;input n322_lo;input n325_lo;input n328_lo;input n334_lo;input n337_lo;input n346_lo;input n349_lo;input n352_lo;input n358_lo;input n361_lo;input n370_lo;input n373_lo;input n376_lo;input n382_lo;input n385_lo;input n394_lo;input n397_lo;input n400_lo;input n406_lo;input n409_lo;input n418_lo;input n421_lo;input n424_lo;input n430_lo;input n433_lo;input n442_lo;input n445_lo;input n448_lo;input n454_lo;input n457_lo;input n466_lo;input n469_lo;input n472_lo;input n478_lo;input n481_lo;input n490_lo;input n493_lo;input n496_lo;input n502_lo;input n505_lo;input n514_lo;input n517_lo;input n520_lo;input n526_lo;input n529_lo;input n538_lo;input n541_lo;input n544_lo;input n550_lo;input n553_lo;input n562_lo;input n565_lo;input n568_lo;input n574_lo;input n577_lo;input n586_lo;input n589_lo;input n592_lo;input n598_lo;input n601_lo;input n610_lo;input n613_lo;input n616_lo;input n622_lo;input n625_lo;input n628_lo;input n634_lo;input n316_inv;input n319_inv;input n997_o2;input n998_o2;input n999_o2;input n1000_o2;input n1001_o2;input n1002_o2;input n1003_o2;input n1004_o2;input n1005_o2;input n1015_o2;input n1016_o2;input n1017_o2;input n1018_o2;input n1019_o2;input n1020_o2;input n1021_o2;input n1022_o2;input n1023_o2;input n376_1_inv;input n235_lo_buf_o2;input n283_lo_buf_o2;input n331_lo_buf_o2;input n379_lo_buf_o2;input n427_lo_buf_o2;input n475_lo_buf_o2;input n523_lo_buf_o2;input n571_lo_buf_o2;input n619_lo_buf_o2;input n406_1_inv;input G223_o2;input G226_o2;input G229_o2;input G232_o2;input G235_o2;input G238_o2;input G242_o2;input G246_o2;input G250_o2;input n259_lo_buf_o2;input n307_lo_buf_o2;input n355_lo_buf_o2;input n403_lo_buf_o2;input n451_lo_buf_o2;input n499_lo_buf_o2;input n547_lo_buf_o2;input n595_lo_buf_o2;input n631_lo_buf_o2;input G213_o2;input G318_o2;input G358_o2;input G259_o2;input G263_o2;input G266_o2;input G269_o2;input G272_o2;input G275_o2;input G278_o2;input G281_o2;input G284_o2;input n211_lo_buf_o2;input n247_lo_buf_o2;input n295_lo_buf_o2;input n343_lo_buf_o2;input n391_lo_buf_o2;input n439_lo_buf_o2;input n487_lo_buf_o2;input n535_lo_buf_o2;input n583_lo_buf_o2;input G158_o2;input G184_o2;input G186_o2;input G188_o2;input G190_o2;input G192_o2;input G194_o2;input G196_o2;input G198_o2;input n223_lo_buf_o2;input n271_lo_buf_o2;input n319_lo_buf_o2;input n367_lo_buf_o2;input n415_lo_buf_o2;input n463_lo_buf_o2;input n511_lo_buf_o2;input n559_lo_buf_o2;input n607_lo_buf_o2;input n580_inv;input G154_o2;input G159_o2;input G162_o2;input G165_o2;input G168_o2;input G171_o2;input G174_o2;input G177_o2;input G180_o2;
  output G426;output G427;output G428;output G429;output G430;output G431;output G432;output n205_li;output n214_li;output n217_li;output n226_li;output n229_li;output n232_li;output n238_li;output n241_li;output n250_li;output n253_li;output n256_li;output n262_li;output n265_li;output n274_li;output n277_li;output n280_li;output n286_li;output n289_li;output n298_li;output n301_li;output n304_li;output n310_li;output n313_li;output n322_li;output n325_li;output n328_li;output n334_li;output n337_li;output n346_li;output n349_li;output n352_li;output n358_li;output n361_li;output n370_li;output n373_li;output n376_li;output n382_li;output n385_li;output n394_li;output n397_li;output n400_li;output n406_li;output n409_li;output n418_li;output n421_li;output n424_li;output n430_li;output n433_li;output n442_li;output n445_li;output n448_li;output n454_li;output n457_li;output n466_li;output n469_li;output n472_li;output n478_li;output n481_li;output n490_li;output n493_li;output n496_li;output n502_li;output n505_li;output n514_li;output n517_li;output n520_li;output n526_li;output n529_li;output n538_li;output n541_li;output n544_li;output n550_li;output n553_li;output n562_li;output n565_li;output n568_li;output n574_li;output n577_li;output n586_li;output n589_li;output n592_li;output n598_li;output n601_li;output n610_li;output n613_li;output n616_li;output n622_li;output n625_li;output n628_li;output n634_li;output n919_i2;output n1024_i2;output n997_i2;output n998_i2;output n999_i2;output n1000_i2;output n1001_i2;output n1002_i2;output n1003_i2;output n1004_i2;output n1005_i2;output n1015_i2;output n1016_i2;output n1017_i2;output n1018_i2;output n1019_i2;output n1020_i2;output n1021_i2;output n1022_i2;output n1023_i2;output G199_i2;output n235_lo_buf_i2;output n283_lo_buf_i2;output n331_lo_buf_i2;output n379_lo_buf_i2;output n427_lo_buf_i2;output n475_lo_buf_i2;output n523_lo_buf_i2;output n571_lo_buf_i2;output n619_lo_buf_i2;output G355_i2;output G223_i2;output G226_i2;output G229_i2;output G232_i2;output G235_i2;output G238_i2;output G242_i2;output G246_i2;output G250_i2;output n259_lo_buf_i2;output n307_lo_buf_i2;output n355_lo_buf_i2;output n403_lo_buf_i2;output n451_lo_buf_i2;output n499_lo_buf_i2;output n547_lo_buf_i2;output n595_lo_buf_i2;output n631_lo_buf_i2;output G213_i2;output G318_i2;output G358_i2;output G259_i2;output G263_i2;output G266_i2;output G269_i2;output G272_i2;output G275_i2;output G278_i2;output G281_i2;output G284_i2;output n211_lo_buf_i2;output n247_lo_buf_i2;output n295_lo_buf_i2;output n343_lo_buf_i2;output n391_lo_buf_i2;output n439_lo_buf_i2;output n487_lo_buf_i2;output n535_lo_buf_i2;output n583_lo_buf_i2;output G158_i2;output G184_i2;output G186_i2;output G188_i2;output G190_i2;output G192_i2;output G194_i2;output G196_i2;output G198_i2;output n223_lo_buf_i2;output n271_lo_buf_i2;output n319_lo_buf_i2;output n367_lo_buf_i2;output n415_lo_buf_i2;output n463_lo_buf_i2;output n511_lo_buf_i2;output n559_lo_buf_i2;output n607_lo_buf_i2;output G295_i2;output G154_i2;output G159_i2;output G162_i2;output G165_i2;output G168_i2;output G171_i2;output G174_i2;output G177_i2;output G180_i2;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire n205_lo_p;
  wire n205_lo_n;
  wire n214_lo_p;
  wire n214_lo_n;
  wire n217_lo_p;
  wire n217_lo_n;
  wire n226_lo_p;
  wire n226_lo_n;
  wire n229_lo_p;
  wire n229_lo_n;
  wire n232_lo_p;
  wire n232_lo_n;
  wire n238_lo_p;
  wire n238_lo_n;
  wire n241_lo_p;
  wire n241_lo_n;
  wire n250_lo_p;
  wire n250_lo_n;
  wire n253_lo_p;
  wire n253_lo_n;
  wire n256_lo_p;
  wire n256_lo_n;
  wire n262_lo_p;
  wire n262_lo_n;
  wire n265_lo_p;
  wire n265_lo_n;
  wire n274_lo_p;
  wire n274_lo_n;
  wire n277_lo_p;
  wire n277_lo_n;
  wire n280_lo_p;
  wire n280_lo_n;
  wire n286_lo_p;
  wire n286_lo_n;
  wire n289_lo_p;
  wire n289_lo_n;
  wire n298_lo_p;
  wire n298_lo_n;
  wire n301_lo_p;
  wire n301_lo_n;
  wire n304_lo_p;
  wire n304_lo_n;
  wire n310_lo_p;
  wire n310_lo_n;
  wire n313_lo_p;
  wire n313_lo_n;
  wire n322_lo_p;
  wire n322_lo_n;
  wire n325_lo_p;
  wire n325_lo_n;
  wire n328_lo_p;
  wire n328_lo_n;
  wire n334_lo_p;
  wire n334_lo_n;
  wire n337_lo_p;
  wire n337_lo_n;
  wire n346_lo_p;
  wire n346_lo_n;
  wire n349_lo_p;
  wire n349_lo_n;
  wire n352_lo_p;
  wire n352_lo_n;
  wire n358_lo_p;
  wire n358_lo_n;
  wire n361_lo_p;
  wire n361_lo_n;
  wire n370_lo_p;
  wire n370_lo_n;
  wire n373_lo_p;
  wire n373_lo_n;
  wire n376_lo_p;
  wire n376_lo_n;
  wire n382_lo_p;
  wire n382_lo_n;
  wire n385_lo_p;
  wire n385_lo_n;
  wire n394_lo_p;
  wire n394_lo_n;
  wire n397_lo_p;
  wire n397_lo_n;
  wire n400_lo_p;
  wire n400_lo_n;
  wire n406_lo_p;
  wire n406_lo_n;
  wire n409_lo_p;
  wire n409_lo_n;
  wire n418_lo_p;
  wire n418_lo_n;
  wire n421_lo_p;
  wire n421_lo_n;
  wire n424_lo_p;
  wire n424_lo_n;
  wire n430_lo_p;
  wire n430_lo_n;
  wire n433_lo_p;
  wire n433_lo_n;
  wire n442_lo_p;
  wire n442_lo_n;
  wire n445_lo_p;
  wire n445_lo_n;
  wire n448_lo_p;
  wire n448_lo_n;
  wire n454_lo_p;
  wire n454_lo_n;
  wire n457_lo_p;
  wire n457_lo_n;
  wire n466_lo_p;
  wire n466_lo_n;
  wire n469_lo_p;
  wire n469_lo_n;
  wire n472_lo_p;
  wire n472_lo_n;
  wire n478_lo_p;
  wire n478_lo_n;
  wire n481_lo_p;
  wire n481_lo_n;
  wire n490_lo_p;
  wire n490_lo_n;
  wire n493_lo_p;
  wire n493_lo_n;
  wire n496_lo_p;
  wire n496_lo_n;
  wire n502_lo_p;
  wire n502_lo_n;
  wire n505_lo_p;
  wire n505_lo_n;
  wire n514_lo_p;
  wire n514_lo_n;
  wire n517_lo_p;
  wire n517_lo_n;
  wire n520_lo_p;
  wire n520_lo_n;
  wire n526_lo_p;
  wire n526_lo_n;
  wire n529_lo_p;
  wire n529_lo_n;
  wire n538_lo_p;
  wire n538_lo_n;
  wire n541_lo_p;
  wire n541_lo_n;
  wire n544_lo_p;
  wire n544_lo_n;
  wire n550_lo_p;
  wire n550_lo_n;
  wire n553_lo_p;
  wire n553_lo_n;
  wire n562_lo_p;
  wire n562_lo_n;
  wire n565_lo_p;
  wire n565_lo_n;
  wire n568_lo_p;
  wire n568_lo_n;
  wire n574_lo_p;
  wire n574_lo_n;
  wire n577_lo_p;
  wire n577_lo_n;
  wire n586_lo_p;
  wire n586_lo_n;
  wire n589_lo_p;
  wire n589_lo_n;
  wire n592_lo_p;
  wire n592_lo_n;
  wire n598_lo_p;
  wire n598_lo_n;
  wire n601_lo_p;
  wire n601_lo_n;
  wire n610_lo_p;
  wire n610_lo_n;
  wire n613_lo_p;
  wire n613_lo_n;
  wire n616_lo_p;
  wire n616_lo_n;
  wire n622_lo_p;
  wire n622_lo_n;
  wire n625_lo_p;
  wire n625_lo_n;
  wire n628_lo_p;
  wire n628_lo_n;
  wire n634_lo_p;
  wire n634_lo_n;
  wire n316_inv_p;
  wire n316_inv_n;
  wire n319_inv_p;
  wire n319_inv_n;
  wire n997_o2_p;
  wire n997_o2_n;
  wire n998_o2_p;
  wire n998_o2_n;
  wire n999_o2_p;
  wire n999_o2_n;
  wire n1000_o2_p;
  wire n1000_o2_n;
  wire n1001_o2_p;
  wire n1001_o2_n;
  wire n1002_o2_p;
  wire n1002_o2_n;
  wire n1003_o2_p;
  wire n1003_o2_n;
  wire n1004_o2_p;
  wire n1004_o2_n;
  wire n1005_o2_p;
  wire n1005_o2_n;
  wire n1015_o2_p;
  wire n1015_o2_n;
  wire n1016_o2_p;
  wire n1016_o2_n;
  wire n1017_o2_p;
  wire n1017_o2_n;
  wire n1018_o2_p;
  wire n1018_o2_n;
  wire n1019_o2_p;
  wire n1019_o2_n;
  wire n1020_o2_p;
  wire n1020_o2_n;
  wire n1021_o2_p;
  wire n1021_o2_n;
  wire n1022_o2_p;
  wire n1022_o2_n;
  wire n1023_o2_p;
  wire n1023_o2_n;
  wire n376_1_inv_p;
  wire n376_1_inv_n;
  wire n235_lo_buf_o2_p;
  wire n235_lo_buf_o2_n;
  wire n283_lo_buf_o2_p;
  wire n283_lo_buf_o2_n;
  wire n331_lo_buf_o2_p;
  wire n331_lo_buf_o2_n;
  wire n379_lo_buf_o2_p;
  wire n379_lo_buf_o2_n;
  wire n427_lo_buf_o2_p;
  wire n427_lo_buf_o2_n;
  wire n475_lo_buf_o2_p;
  wire n475_lo_buf_o2_n;
  wire n523_lo_buf_o2_p;
  wire n523_lo_buf_o2_n;
  wire n571_lo_buf_o2_p;
  wire n571_lo_buf_o2_n;
  wire n619_lo_buf_o2_p;
  wire n619_lo_buf_o2_n;
  wire n406_1_inv_p;
  wire n406_1_inv_n;
  wire G223_o2_p;
  wire G223_o2_n;
  wire G226_o2_p;
  wire G226_o2_n;
  wire G229_o2_p;
  wire G229_o2_n;
  wire G232_o2_p;
  wire G232_o2_n;
  wire G235_o2_p;
  wire G235_o2_n;
  wire G238_o2_p;
  wire G238_o2_n;
  wire G242_o2_p;
  wire G242_o2_n;
  wire G246_o2_p;
  wire G246_o2_n;
  wire G250_o2_p;
  wire G250_o2_n;
  wire n259_lo_buf_o2_p;
  wire n259_lo_buf_o2_n;
  wire n307_lo_buf_o2_p;
  wire n307_lo_buf_o2_n;
  wire n355_lo_buf_o2_p;
  wire n355_lo_buf_o2_n;
  wire n403_lo_buf_o2_p;
  wire n403_lo_buf_o2_n;
  wire n451_lo_buf_o2_p;
  wire n451_lo_buf_o2_n;
  wire n499_lo_buf_o2_p;
  wire n499_lo_buf_o2_n;
  wire n547_lo_buf_o2_p;
  wire n547_lo_buf_o2_n;
  wire n595_lo_buf_o2_p;
  wire n595_lo_buf_o2_n;
  wire n631_lo_buf_o2_p;
  wire n631_lo_buf_o2_n;
  wire G213_o2_p;
  wire G213_o2_n;
  wire G318_o2_p;
  wire G318_o2_n;
  wire G358_o2_p;
  wire G358_o2_n;
  wire G259_o2_p;
  wire G259_o2_n;
  wire G263_o2_p;
  wire G263_o2_n;
  wire G266_o2_p;
  wire G266_o2_n;
  wire G269_o2_p;
  wire G269_o2_n;
  wire G272_o2_p;
  wire G272_o2_n;
  wire G275_o2_p;
  wire G275_o2_n;
  wire G278_o2_p;
  wire G278_o2_n;
  wire G281_o2_p;
  wire G281_o2_n;
  wire G284_o2_p;
  wire G284_o2_n;
  wire n211_lo_buf_o2_p;
  wire n211_lo_buf_o2_n;
  wire n247_lo_buf_o2_p;
  wire n247_lo_buf_o2_n;
  wire n295_lo_buf_o2_p;
  wire n295_lo_buf_o2_n;
  wire n343_lo_buf_o2_p;
  wire n343_lo_buf_o2_n;
  wire n391_lo_buf_o2_p;
  wire n391_lo_buf_o2_n;
  wire n439_lo_buf_o2_p;
  wire n439_lo_buf_o2_n;
  wire n487_lo_buf_o2_p;
  wire n487_lo_buf_o2_n;
  wire n535_lo_buf_o2_p;
  wire n535_lo_buf_o2_n;
  wire n583_lo_buf_o2_p;
  wire n583_lo_buf_o2_n;
  wire G158_o2_p;
  wire G158_o2_n;
  wire G184_o2_p;
  wire G184_o2_n;
  wire G186_o2_p;
  wire G186_o2_n;
  wire G188_o2_p;
  wire G188_o2_n;
  wire G190_o2_p;
  wire G190_o2_n;
  wire G192_o2_p;
  wire G192_o2_n;
  wire G194_o2_p;
  wire G194_o2_n;
  wire G196_o2_p;
  wire G196_o2_n;
  wire G198_o2_p;
  wire G198_o2_n;
  wire n223_lo_buf_o2_p;
  wire n223_lo_buf_o2_n;
  wire n271_lo_buf_o2_p;
  wire n271_lo_buf_o2_n;
  wire n319_lo_buf_o2_p;
  wire n319_lo_buf_o2_n;
  wire n367_lo_buf_o2_p;
  wire n367_lo_buf_o2_n;
  wire n415_lo_buf_o2_p;
  wire n415_lo_buf_o2_n;
  wire n463_lo_buf_o2_p;
  wire n463_lo_buf_o2_n;
  wire n511_lo_buf_o2_p;
  wire n511_lo_buf_o2_n;
  wire n559_lo_buf_o2_p;
  wire n559_lo_buf_o2_n;
  wire n607_lo_buf_o2_p;
  wire n607_lo_buf_o2_n;
  wire n580_inv_p;
  wire n580_inv_n;
  wire G154_o2_p;
  wire G154_o2_n;
  wire G159_o2_p;
  wire G159_o2_n;
  wire G162_o2_p;
  wire G162_o2_n;
  wire G165_o2_p;
  wire G165_o2_n;
  wire G168_o2_p;
  wire G168_o2_n;
  wire G171_o2_p;
  wire G171_o2_n;
  wire G174_o2_p;
  wire G174_o2_n;
  wire G177_o2_p;
  wire G177_o2_n;
  wire G180_o2_p;
  wire G180_o2_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire G213_o2_n_spl_;
  wire G213_o2_n_spl_0;
  wire G213_o2_n_spl_00;
  wire G213_o2_n_spl_1;
  wire G318_o2_n_spl_;
  wire G318_o2_n_spl_0;
  wire G318_o2_n_spl_00;
  wire G318_o2_n_spl_1;
  wire G358_o2_n_spl_;
  wire G358_o2_n_spl_0;
  wire G358_o2_n_spl_00;
  wire G358_o2_n_spl_1;
  wire G213_o2_p_spl_;
  wire G213_o2_p_spl_0;
  wire G213_o2_p_spl_00;
  wire G213_o2_p_spl_01;
  wire G213_o2_p_spl_1;
  wire G213_o2_p_spl_10;
  wire G213_o2_p_spl_11;
  wire G318_o2_p_spl_;
  wire G318_o2_p_spl_0;
  wire G318_o2_p_spl_00;
  wire G318_o2_p_spl_01;
  wire G318_o2_p_spl_1;
  wire G318_o2_p_spl_10;
  wire G318_o2_p_spl_11;
  wire G358_o2_p_spl_;
  wire G358_o2_p_spl_0;
  wire G358_o2_p_spl_00;
  wire G358_o2_p_spl_01;
  wire G358_o2_p_spl_1;
  wire G358_o2_p_spl_10;
  wire G358_o2_p_spl_11;
  wire g236_n_spl_;
  wire g279_p_spl_;
  wire g279_p_spl_0;
  wire g248_n_spl_;
  wire g254_n_spl_;
  wire g260_n_spl_;
  wire g266_n_spl_;
  wire g272_n_spl_;
  wire g242_p_spl_;
  wire g287_n_spl_;
  wire g248_p_spl_;
  wire g290_n_spl_;
  wire g254_p_spl_;
  wire g292_n_spl_;
  wire G159_o2_n_spl_;
  wire G154_o2_n_spl_;
  wire G159_o2_p_spl_;
  wire G154_o2_p_spl_;
  wire G162_o2_n_spl_;
  wire G162_o2_p_spl_;
  wire G165_o2_n_spl_;
  wire G165_o2_p_spl_;
  wire G168_o2_n_spl_;
  wire G168_o2_p_spl_;
  wire G171_o2_n_spl_;
  wire G171_o2_p_spl_;
  wire G174_o2_n_spl_;
  wire G174_o2_p_spl_;
  wire G177_o2_n_spl_;
  wire G177_o2_p_spl_;
  wire G180_o2_n_spl_;
  wire G180_o2_p_spl_;
  wire n580_inv_n_spl_;
  wire n580_inv_n_spl_0;
  wire n580_inv_n_spl_00;
  wire n580_inv_n_spl_000;
  wire n580_inv_n_spl_01;
  wire n580_inv_n_spl_1;
  wire n580_inv_n_spl_10;
  wire n580_inv_n_spl_11;
  wire n580_inv_p_spl_;
  wire n580_inv_p_spl_0;
  wire n580_inv_p_spl_00;
  wire n580_inv_p_spl_000;
  wire n580_inv_p_spl_001;
  wire n580_inv_p_spl_01;
  wire n580_inv_p_spl_010;
  wire n580_inv_p_spl_1;
  wire n580_inv_p_spl_10;
  wire n580_inv_p_spl_11;
  wire g309_p_spl_;
  wire g309_p_spl_0;
  wire g309_p_spl_00;
  wire g309_p_spl_000;
  wire g309_p_spl_01;
  wire g309_p_spl_1;
  wire g309_p_spl_10;
  wire g309_p_spl_11;
  wire g309_n_spl_;
  wire g309_n_spl_0;
  wire g309_n_spl_00;
  wire g309_n_spl_000;
  wire g309_n_spl_001;
  wire g309_n_spl_01;
  wire g309_n_spl_1;
  wire g309_n_spl_10;
  wire g309_n_spl_11;
  wire n223_lo_buf_o2_p_spl_;
  wire n223_lo_buf_o2_p_spl_0;
  wire g365_n_spl_;
  wire n271_lo_buf_o2_p_spl_;
  wire n271_lo_buf_o2_p_spl_0;
  wire g368_n_spl_;
  wire n319_lo_buf_o2_p_spl_;
  wire n319_lo_buf_o2_p_spl_0;
  wire g371_n_spl_;
  wire n367_lo_buf_o2_p_spl_;
  wire n367_lo_buf_o2_p_spl_0;
  wire g374_n_spl_;
  wire n415_lo_buf_o2_p_spl_;
  wire n415_lo_buf_o2_p_spl_0;
  wire g377_n_spl_;
  wire n463_lo_buf_o2_p_spl_;
  wire n463_lo_buf_o2_p_spl_0;
  wire g380_n_spl_;
  wire n511_lo_buf_o2_p_spl_;
  wire n511_lo_buf_o2_p_spl_0;
  wire g383_n_spl_;
  wire n559_lo_buf_o2_p_spl_;
  wire n559_lo_buf_o2_p_spl_0;
  wire g386_n_spl_;
  wire n607_lo_buf_o2_p_spl_;
  wire n607_lo_buf_o2_p_spl_0;
  wire g389_n_spl_;
  wire g393_p_spl_;
  wire g391_p_spl_;
  wire g395_p_spl_;
  wire g397_p_spl_;
  wire g399_p_spl_;
  wire g401_p_spl_;
  wire g403_p_spl_;
  wire g405_p_spl_;
  wire g407_p_spl_;
  wire n217_lo_p_spl_;
  wire n265_lo_p_spl_;
  wire n313_lo_p_spl_;
  wire n361_lo_p_spl_;
  wire n409_lo_p_spl_;
  wire n457_lo_p_spl_;
  wire n505_lo_p_spl_;
  wire n553_lo_p_spl_;
  wire n601_lo_p_spl_;
  wire n376_1_inv_p_spl_;
  wire g362_n_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    n205_lo_p,
    n205_lo
  );


  not

  (
    n205_lo_n,
    n205_lo
  );


  buf

  (
    n214_lo_p,
    n214_lo
  );


  not

  (
    n214_lo_n,
    n214_lo
  );


  buf

  (
    n217_lo_p,
    n217_lo
  );


  not

  (
    n217_lo_n,
    n217_lo
  );


  buf

  (
    n226_lo_p,
    n226_lo
  );


  not

  (
    n226_lo_n,
    n226_lo
  );


  buf

  (
    n229_lo_p,
    n229_lo
  );


  not

  (
    n229_lo_n,
    n229_lo
  );


  buf

  (
    n232_lo_p,
    n232_lo
  );


  not

  (
    n232_lo_n,
    n232_lo
  );


  buf

  (
    n238_lo_p,
    n238_lo
  );


  not

  (
    n238_lo_n,
    n238_lo
  );


  buf

  (
    n241_lo_p,
    n241_lo
  );


  not

  (
    n241_lo_n,
    n241_lo
  );


  buf

  (
    n250_lo_p,
    n250_lo
  );


  not

  (
    n250_lo_n,
    n250_lo
  );


  buf

  (
    n253_lo_p,
    n253_lo
  );


  not

  (
    n253_lo_n,
    n253_lo
  );


  buf

  (
    n256_lo_p,
    n256_lo
  );


  not

  (
    n256_lo_n,
    n256_lo
  );


  buf

  (
    n262_lo_p,
    n262_lo
  );


  not

  (
    n262_lo_n,
    n262_lo
  );


  buf

  (
    n265_lo_p,
    n265_lo
  );


  not

  (
    n265_lo_n,
    n265_lo
  );


  buf

  (
    n274_lo_p,
    n274_lo
  );


  not

  (
    n274_lo_n,
    n274_lo
  );


  buf

  (
    n277_lo_p,
    n277_lo
  );


  not

  (
    n277_lo_n,
    n277_lo
  );


  buf

  (
    n280_lo_p,
    n280_lo
  );


  not

  (
    n280_lo_n,
    n280_lo
  );


  buf

  (
    n286_lo_p,
    n286_lo
  );


  not

  (
    n286_lo_n,
    n286_lo
  );


  buf

  (
    n289_lo_p,
    n289_lo
  );


  not

  (
    n289_lo_n,
    n289_lo
  );


  buf

  (
    n298_lo_p,
    n298_lo
  );


  not

  (
    n298_lo_n,
    n298_lo
  );


  buf

  (
    n301_lo_p,
    n301_lo
  );


  not

  (
    n301_lo_n,
    n301_lo
  );


  buf

  (
    n304_lo_p,
    n304_lo
  );


  not

  (
    n304_lo_n,
    n304_lo
  );


  buf

  (
    n310_lo_p,
    n310_lo
  );


  not

  (
    n310_lo_n,
    n310_lo
  );


  buf

  (
    n313_lo_p,
    n313_lo
  );


  not

  (
    n313_lo_n,
    n313_lo
  );


  buf

  (
    n322_lo_p,
    n322_lo
  );


  not

  (
    n322_lo_n,
    n322_lo
  );


  buf

  (
    n325_lo_p,
    n325_lo
  );


  not

  (
    n325_lo_n,
    n325_lo
  );


  buf

  (
    n328_lo_p,
    n328_lo
  );


  not

  (
    n328_lo_n,
    n328_lo
  );


  buf

  (
    n334_lo_p,
    n334_lo
  );


  not

  (
    n334_lo_n,
    n334_lo
  );


  buf

  (
    n337_lo_p,
    n337_lo
  );


  not

  (
    n337_lo_n,
    n337_lo
  );


  buf

  (
    n346_lo_p,
    n346_lo
  );


  not

  (
    n346_lo_n,
    n346_lo
  );


  buf

  (
    n349_lo_p,
    n349_lo
  );


  not

  (
    n349_lo_n,
    n349_lo
  );


  buf

  (
    n352_lo_p,
    n352_lo
  );


  not

  (
    n352_lo_n,
    n352_lo
  );


  buf

  (
    n358_lo_p,
    n358_lo
  );


  not

  (
    n358_lo_n,
    n358_lo
  );


  buf

  (
    n361_lo_p,
    n361_lo
  );


  not

  (
    n361_lo_n,
    n361_lo
  );


  buf

  (
    n370_lo_p,
    n370_lo
  );


  not

  (
    n370_lo_n,
    n370_lo
  );


  buf

  (
    n373_lo_p,
    n373_lo
  );


  not

  (
    n373_lo_n,
    n373_lo
  );


  buf

  (
    n376_lo_p,
    n376_lo
  );


  not

  (
    n376_lo_n,
    n376_lo
  );


  buf

  (
    n382_lo_p,
    n382_lo
  );


  not

  (
    n382_lo_n,
    n382_lo
  );


  buf

  (
    n385_lo_p,
    n385_lo
  );


  not

  (
    n385_lo_n,
    n385_lo
  );


  buf

  (
    n394_lo_p,
    n394_lo
  );


  not

  (
    n394_lo_n,
    n394_lo
  );


  buf

  (
    n397_lo_p,
    n397_lo
  );


  not

  (
    n397_lo_n,
    n397_lo
  );


  buf

  (
    n400_lo_p,
    n400_lo
  );


  not

  (
    n400_lo_n,
    n400_lo
  );


  buf

  (
    n406_lo_p,
    n406_lo
  );


  not

  (
    n406_lo_n,
    n406_lo
  );


  buf

  (
    n409_lo_p,
    n409_lo
  );


  not

  (
    n409_lo_n,
    n409_lo
  );


  buf

  (
    n418_lo_p,
    n418_lo
  );


  not

  (
    n418_lo_n,
    n418_lo
  );


  buf

  (
    n421_lo_p,
    n421_lo
  );


  not

  (
    n421_lo_n,
    n421_lo
  );


  buf

  (
    n424_lo_p,
    n424_lo
  );


  not

  (
    n424_lo_n,
    n424_lo
  );


  buf

  (
    n430_lo_p,
    n430_lo
  );


  not

  (
    n430_lo_n,
    n430_lo
  );


  buf

  (
    n433_lo_p,
    n433_lo
  );


  not

  (
    n433_lo_n,
    n433_lo
  );


  buf

  (
    n442_lo_p,
    n442_lo
  );


  not

  (
    n442_lo_n,
    n442_lo
  );


  buf

  (
    n445_lo_p,
    n445_lo
  );


  not

  (
    n445_lo_n,
    n445_lo
  );


  buf

  (
    n448_lo_p,
    n448_lo
  );


  not

  (
    n448_lo_n,
    n448_lo
  );


  buf

  (
    n454_lo_p,
    n454_lo
  );


  not

  (
    n454_lo_n,
    n454_lo
  );


  buf

  (
    n457_lo_p,
    n457_lo
  );


  not

  (
    n457_lo_n,
    n457_lo
  );


  buf

  (
    n466_lo_p,
    n466_lo
  );


  not

  (
    n466_lo_n,
    n466_lo
  );


  buf

  (
    n469_lo_p,
    n469_lo
  );


  not

  (
    n469_lo_n,
    n469_lo
  );


  buf

  (
    n472_lo_p,
    n472_lo
  );


  not

  (
    n472_lo_n,
    n472_lo
  );


  buf

  (
    n478_lo_p,
    n478_lo
  );


  not

  (
    n478_lo_n,
    n478_lo
  );


  buf

  (
    n481_lo_p,
    n481_lo
  );


  not

  (
    n481_lo_n,
    n481_lo
  );


  buf

  (
    n490_lo_p,
    n490_lo
  );


  not

  (
    n490_lo_n,
    n490_lo
  );


  buf

  (
    n493_lo_p,
    n493_lo
  );


  not

  (
    n493_lo_n,
    n493_lo
  );


  buf

  (
    n496_lo_p,
    n496_lo
  );


  not

  (
    n496_lo_n,
    n496_lo
  );


  buf

  (
    n502_lo_p,
    n502_lo
  );


  not

  (
    n502_lo_n,
    n502_lo
  );


  buf

  (
    n505_lo_p,
    n505_lo
  );


  not

  (
    n505_lo_n,
    n505_lo
  );


  buf

  (
    n514_lo_p,
    n514_lo
  );


  not

  (
    n514_lo_n,
    n514_lo
  );


  buf

  (
    n517_lo_p,
    n517_lo
  );


  not

  (
    n517_lo_n,
    n517_lo
  );


  buf

  (
    n520_lo_p,
    n520_lo
  );


  not

  (
    n520_lo_n,
    n520_lo
  );


  buf

  (
    n526_lo_p,
    n526_lo
  );


  not

  (
    n526_lo_n,
    n526_lo
  );


  buf

  (
    n529_lo_p,
    n529_lo
  );


  not

  (
    n529_lo_n,
    n529_lo
  );


  buf

  (
    n538_lo_p,
    n538_lo
  );


  not

  (
    n538_lo_n,
    n538_lo
  );


  buf

  (
    n541_lo_p,
    n541_lo
  );


  not

  (
    n541_lo_n,
    n541_lo
  );


  buf

  (
    n544_lo_p,
    n544_lo
  );


  not

  (
    n544_lo_n,
    n544_lo
  );


  buf

  (
    n550_lo_p,
    n550_lo
  );


  not

  (
    n550_lo_n,
    n550_lo
  );


  buf

  (
    n553_lo_p,
    n553_lo
  );


  not

  (
    n553_lo_n,
    n553_lo
  );


  buf

  (
    n562_lo_p,
    n562_lo
  );


  not

  (
    n562_lo_n,
    n562_lo
  );


  buf

  (
    n565_lo_p,
    n565_lo
  );


  not

  (
    n565_lo_n,
    n565_lo
  );


  buf

  (
    n568_lo_p,
    n568_lo
  );


  not

  (
    n568_lo_n,
    n568_lo
  );


  buf

  (
    n574_lo_p,
    n574_lo
  );


  not

  (
    n574_lo_n,
    n574_lo
  );


  buf

  (
    n577_lo_p,
    n577_lo
  );


  not

  (
    n577_lo_n,
    n577_lo
  );


  buf

  (
    n586_lo_p,
    n586_lo
  );


  not

  (
    n586_lo_n,
    n586_lo
  );


  buf

  (
    n589_lo_p,
    n589_lo
  );


  not

  (
    n589_lo_n,
    n589_lo
  );


  buf

  (
    n592_lo_p,
    n592_lo
  );


  not

  (
    n592_lo_n,
    n592_lo
  );


  buf

  (
    n598_lo_p,
    n598_lo
  );


  not

  (
    n598_lo_n,
    n598_lo
  );


  buf

  (
    n601_lo_p,
    n601_lo
  );


  not

  (
    n601_lo_n,
    n601_lo
  );


  buf

  (
    n610_lo_p,
    n610_lo
  );


  not

  (
    n610_lo_n,
    n610_lo
  );


  buf

  (
    n613_lo_p,
    n613_lo
  );


  not

  (
    n613_lo_n,
    n613_lo
  );


  buf

  (
    n616_lo_p,
    n616_lo
  );


  not

  (
    n616_lo_n,
    n616_lo
  );


  buf

  (
    n622_lo_p,
    n622_lo
  );


  not

  (
    n622_lo_n,
    n622_lo
  );


  buf

  (
    n625_lo_p,
    n625_lo
  );


  not

  (
    n625_lo_n,
    n625_lo
  );


  buf

  (
    n628_lo_p,
    n628_lo
  );


  not

  (
    n628_lo_n,
    n628_lo
  );


  buf

  (
    n634_lo_p,
    n634_lo
  );


  not

  (
    n634_lo_n,
    n634_lo
  );


  buf

  (
    n316_inv_p,
    n316_inv
  );


  not

  (
    n316_inv_n,
    n316_inv
  );


  buf

  (
    n319_inv_p,
    n319_inv
  );


  not

  (
    n319_inv_n,
    n319_inv
  );


  buf

  (
    n997_o2_p,
    n997_o2
  );


  not

  (
    n997_o2_n,
    n997_o2
  );


  buf

  (
    n998_o2_p,
    n998_o2
  );


  not

  (
    n998_o2_n,
    n998_o2
  );


  buf

  (
    n999_o2_p,
    n999_o2
  );


  not

  (
    n999_o2_n,
    n999_o2
  );


  buf

  (
    n1000_o2_p,
    n1000_o2
  );


  not

  (
    n1000_o2_n,
    n1000_o2
  );


  buf

  (
    n1001_o2_p,
    n1001_o2
  );


  not

  (
    n1001_o2_n,
    n1001_o2
  );


  buf

  (
    n1002_o2_p,
    n1002_o2
  );


  not

  (
    n1002_o2_n,
    n1002_o2
  );


  buf

  (
    n1003_o2_p,
    n1003_o2
  );


  not

  (
    n1003_o2_n,
    n1003_o2
  );


  buf

  (
    n1004_o2_p,
    n1004_o2
  );


  not

  (
    n1004_o2_n,
    n1004_o2
  );


  buf

  (
    n1005_o2_p,
    n1005_o2
  );


  not

  (
    n1005_o2_n,
    n1005_o2
  );


  buf

  (
    n1015_o2_p,
    n1015_o2
  );


  not

  (
    n1015_o2_n,
    n1015_o2
  );


  buf

  (
    n1016_o2_p,
    n1016_o2
  );


  not

  (
    n1016_o2_n,
    n1016_o2
  );


  buf

  (
    n1017_o2_p,
    n1017_o2
  );


  not

  (
    n1017_o2_n,
    n1017_o2
  );


  buf

  (
    n1018_o2_p,
    n1018_o2
  );


  not

  (
    n1018_o2_n,
    n1018_o2
  );


  buf

  (
    n1019_o2_p,
    n1019_o2
  );


  not

  (
    n1019_o2_n,
    n1019_o2
  );


  buf

  (
    n1020_o2_p,
    n1020_o2
  );


  not

  (
    n1020_o2_n,
    n1020_o2
  );


  buf

  (
    n1021_o2_p,
    n1021_o2
  );


  not

  (
    n1021_o2_n,
    n1021_o2
  );


  buf

  (
    n1022_o2_p,
    n1022_o2
  );


  not

  (
    n1022_o2_n,
    n1022_o2
  );


  buf

  (
    n1023_o2_p,
    n1023_o2
  );


  not

  (
    n1023_o2_n,
    n1023_o2
  );


  buf

  (
    n376_1_inv_p,
    n376_1_inv
  );


  not

  (
    n376_1_inv_n,
    n376_1_inv
  );


  buf

  (
    n235_lo_buf_o2_p,
    n235_lo_buf_o2
  );


  not

  (
    n235_lo_buf_o2_n,
    n235_lo_buf_o2
  );


  buf

  (
    n283_lo_buf_o2_p,
    n283_lo_buf_o2
  );


  not

  (
    n283_lo_buf_o2_n,
    n283_lo_buf_o2
  );


  buf

  (
    n331_lo_buf_o2_p,
    n331_lo_buf_o2
  );


  not

  (
    n331_lo_buf_o2_n,
    n331_lo_buf_o2
  );


  buf

  (
    n379_lo_buf_o2_p,
    n379_lo_buf_o2
  );


  not

  (
    n379_lo_buf_o2_n,
    n379_lo_buf_o2
  );


  buf

  (
    n427_lo_buf_o2_p,
    n427_lo_buf_o2
  );


  not

  (
    n427_lo_buf_o2_n,
    n427_lo_buf_o2
  );


  buf

  (
    n475_lo_buf_o2_p,
    n475_lo_buf_o2
  );


  not

  (
    n475_lo_buf_o2_n,
    n475_lo_buf_o2
  );


  buf

  (
    n523_lo_buf_o2_p,
    n523_lo_buf_o2
  );


  not

  (
    n523_lo_buf_o2_n,
    n523_lo_buf_o2
  );


  buf

  (
    n571_lo_buf_o2_p,
    n571_lo_buf_o2
  );


  not

  (
    n571_lo_buf_o2_n,
    n571_lo_buf_o2
  );


  buf

  (
    n619_lo_buf_o2_p,
    n619_lo_buf_o2
  );


  not

  (
    n619_lo_buf_o2_n,
    n619_lo_buf_o2
  );


  buf

  (
    n406_1_inv_p,
    n406_1_inv
  );


  not

  (
    n406_1_inv_n,
    n406_1_inv
  );


  buf

  (
    G223_o2_p,
    G223_o2
  );


  not

  (
    G223_o2_n,
    G223_o2
  );


  buf

  (
    G226_o2_p,
    G226_o2
  );


  not

  (
    G226_o2_n,
    G226_o2
  );


  buf

  (
    G229_o2_p,
    G229_o2
  );


  not

  (
    G229_o2_n,
    G229_o2
  );


  buf

  (
    G232_o2_p,
    G232_o2
  );


  not

  (
    G232_o2_n,
    G232_o2
  );


  buf

  (
    G235_o2_p,
    G235_o2
  );


  not

  (
    G235_o2_n,
    G235_o2
  );


  buf

  (
    G238_o2_p,
    G238_o2
  );


  not

  (
    G238_o2_n,
    G238_o2
  );


  buf

  (
    G242_o2_p,
    G242_o2
  );


  not

  (
    G242_o2_n,
    G242_o2
  );


  buf

  (
    G246_o2_p,
    G246_o2
  );


  not

  (
    G246_o2_n,
    G246_o2
  );


  buf

  (
    G250_o2_p,
    G250_o2
  );


  not

  (
    G250_o2_n,
    G250_o2
  );


  buf

  (
    n259_lo_buf_o2_p,
    n259_lo_buf_o2
  );


  not

  (
    n259_lo_buf_o2_n,
    n259_lo_buf_o2
  );


  buf

  (
    n307_lo_buf_o2_p,
    n307_lo_buf_o2
  );


  not

  (
    n307_lo_buf_o2_n,
    n307_lo_buf_o2
  );


  buf

  (
    n355_lo_buf_o2_p,
    n355_lo_buf_o2
  );


  not

  (
    n355_lo_buf_o2_n,
    n355_lo_buf_o2
  );


  buf

  (
    n403_lo_buf_o2_p,
    n403_lo_buf_o2
  );


  not

  (
    n403_lo_buf_o2_n,
    n403_lo_buf_o2
  );


  buf

  (
    n451_lo_buf_o2_p,
    n451_lo_buf_o2
  );


  not

  (
    n451_lo_buf_o2_n,
    n451_lo_buf_o2
  );


  buf

  (
    n499_lo_buf_o2_p,
    n499_lo_buf_o2
  );


  not

  (
    n499_lo_buf_o2_n,
    n499_lo_buf_o2
  );


  buf

  (
    n547_lo_buf_o2_p,
    n547_lo_buf_o2
  );


  not

  (
    n547_lo_buf_o2_n,
    n547_lo_buf_o2
  );


  buf

  (
    n595_lo_buf_o2_p,
    n595_lo_buf_o2
  );


  not

  (
    n595_lo_buf_o2_n,
    n595_lo_buf_o2
  );


  buf

  (
    n631_lo_buf_o2_p,
    n631_lo_buf_o2
  );


  not

  (
    n631_lo_buf_o2_n,
    n631_lo_buf_o2
  );


  buf

  (
    G213_o2_p,
    G213_o2
  );


  not

  (
    G213_o2_n,
    G213_o2
  );


  buf

  (
    G318_o2_p,
    G318_o2
  );


  not

  (
    G318_o2_n,
    G318_o2
  );


  buf

  (
    G358_o2_p,
    G358_o2
  );


  not

  (
    G358_o2_n,
    G358_o2
  );


  buf

  (
    G259_o2_p,
    G259_o2
  );


  not

  (
    G259_o2_n,
    G259_o2
  );


  buf

  (
    G263_o2_p,
    G263_o2
  );


  not

  (
    G263_o2_n,
    G263_o2
  );


  buf

  (
    G266_o2_p,
    G266_o2
  );


  not

  (
    G266_o2_n,
    G266_o2
  );


  buf

  (
    G269_o2_p,
    G269_o2
  );


  not

  (
    G269_o2_n,
    G269_o2
  );


  buf

  (
    G272_o2_p,
    G272_o2
  );


  not

  (
    G272_o2_n,
    G272_o2
  );


  buf

  (
    G275_o2_p,
    G275_o2
  );


  not

  (
    G275_o2_n,
    G275_o2
  );


  buf

  (
    G278_o2_p,
    G278_o2
  );


  not

  (
    G278_o2_n,
    G278_o2
  );


  buf

  (
    G281_o2_p,
    G281_o2
  );


  not

  (
    G281_o2_n,
    G281_o2
  );


  buf

  (
    G284_o2_p,
    G284_o2
  );


  not

  (
    G284_o2_n,
    G284_o2
  );


  buf

  (
    n211_lo_buf_o2_p,
    n211_lo_buf_o2
  );


  not

  (
    n211_lo_buf_o2_n,
    n211_lo_buf_o2
  );


  buf

  (
    n247_lo_buf_o2_p,
    n247_lo_buf_o2
  );


  not

  (
    n247_lo_buf_o2_n,
    n247_lo_buf_o2
  );


  buf

  (
    n295_lo_buf_o2_p,
    n295_lo_buf_o2
  );


  not

  (
    n295_lo_buf_o2_n,
    n295_lo_buf_o2
  );


  buf

  (
    n343_lo_buf_o2_p,
    n343_lo_buf_o2
  );


  not

  (
    n343_lo_buf_o2_n,
    n343_lo_buf_o2
  );


  buf

  (
    n391_lo_buf_o2_p,
    n391_lo_buf_o2
  );


  not

  (
    n391_lo_buf_o2_n,
    n391_lo_buf_o2
  );


  buf

  (
    n439_lo_buf_o2_p,
    n439_lo_buf_o2
  );


  not

  (
    n439_lo_buf_o2_n,
    n439_lo_buf_o2
  );


  buf

  (
    n487_lo_buf_o2_p,
    n487_lo_buf_o2
  );


  not

  (
    n487_lo_buf_o2_n,
    n487_lo_buf_o2
  );


  buf

  (
    n535_lo_buf_o2_p,
    n535_lo_buf_o2
  );


  not

  (
    n535_lo_buf_o2_n,
    n535_lo_buf_o2
  );


  buf

  (
    n583_lo_buf_o2_p,
    n583_lo_buf_o2
  );


  not

  (
    n583_lo_buf_o2_n,
    n583_lo_buf_o2
  );


  buf

  (
    G158_o2_p,
    G158_o2
  );


  not

  (
    G158_o2_n,
    G158_o2
  );


  buf

  (
    G184_o2_p,
    G184_o2
  );


  not

  (
    G184_o2_n,
    G184_o2
  );


  buf

  (
    G186_o2_p,
    G186_o2
  );


  not

  (
    G186_o2_n,
    G186_o2
  );


  buf

  (
    G188_o2_p,
    G188_o2
  );


  not

  (
    G188_o2_n,
    G188_o2
  );


  buf

  (
    G190_o2_p,
    G190_o2
  );


  not

  (
    G190_o2_n,
    G190_o2
  );


  buf

  (
    G192_o2_p,
    G192_o2
  );


  not

  (
    G192_o2_n,
    G192_o2
  );


  buf

  (
    G194_o2_p,
    G194_o2
  );


  not

  (
    G194_o2_n,
    G194_o2
  );


  buf

  (
    G196_o2_p,
    G196_o2
  );


  not

  (
    G196_o2_n,
    G196_o2
  );


  buf

  (
    G198_o2_p,
    G198_o2
  );


  not

  (
    G198_o2_n,
    G198_o2
  );


  buf

  (
    n223_lo_buf_o2_p,
    n223_lo_buf_o2
  );


  not

  (
    n223_lo_buf_o2_n,
    n223_lo_buf_o2
  );


  buf

  (
    n271_lo_buf_o2_p,
    n271_lo_buf_o2
  );


  not

  (
    n271_lo_buf_o2_n,
    n271_lo_buf_o2
  );


  buf

  (
    n319_lo_buf_o2_p,
    n319_lo_buf_o2
  );


  not

  (
    n319_lo_buf_o2_n,
    n319_lo_buf_o2
  );


  buf

  (
    n367_lo_buf_o2_p,
    n367_lo_buf_o2
  );


  not

  (
    n367_lo_buf_o2_n,
    n367_lo_buf_o2
  );


  buf

  (
    n415_lo_buf_o2_p,
    n415_lo_buf_o2
  );


  not

  (
    n415_lo_buf_o2_n,
    n415_lo_buf_o2
  );


  buf

  (
    n463_lo_buf_o2_p,
    n463_lo_buf_o2
  );


  not

  (
    n463_lo_buf_o2_n,
    n463_lo_buf_o2
  );


  buf

  (
    n511_lo_buf_o2_p,
    n511_lo_buf_o2
  );


  not

  (
    n511_lo_buf_o2_n,
    n511_lo_buf_o2
  );


  buf

  (
    n559_lo_buf_o2_p,
    n559_lo_buf_o2
  );


  not

  (
    n559_lo_buf_o2_n,
    n559_lo_buf_o2
  );


  buf

  (
    n607_lo_buf_o2_p,
    n607_lo_buf_o2
  );


  not

  (
    n607_lo_buf_o2_n,
    n607_lo_buf_o2
  );


  buf

  (
    n580_inv_p,
    n580_inv
  );


  not

  (
    n580_inv_n,
    n580_inv
  );


  buf

  (
    G154_o2_p,
    G154_o2
  );


  not

  (
    G154_o2_n,
    G154_o2
  );


  buf

  (
    G159_o2_p,
    G159_o2
  );


  not

  (
    G159_o2_n,
    G159_o2
  );


  buf

  (
    G162_o2_p,
    G162_o2
  );


  not

  (
    G162_o2_n,
    G162_o2
  );


  buf

  (
    G165_o2_p,
    G165_o2
  );


  not

  (
    G165_o2_n,
    G165_o2
  );


  buf

  (
    G168_o2_p,
    G168_o2
  );


  not

  (
    G168_o2_n,
    G168_o2
  );


  buf

  (
    G171_o2_p,
    G171_o2
  );


  not

  (
    G171_o2_n,
    G171_o2
  );


  buf

  (
    G174_o2_p,
    G174_o2
  );


  not

  (
    G174_o2_n,
    G174_o2
  );


  buf

  (
    G177_o2_p,
    G177_o2
  );


  not

  (
    G177_o2_n,
    G177_o2
  );


  buf

  (
    G180_o2_p,
    G180_o2
  );


  not

  (
    G180_o2_n,
    G180_o2
  );


  or

  (
    g225_n,
    G213_o2_n_spl_00,
    n214_lo_n
  );


  or

  (
    g226_n,
    G318_o2_n_spl_00,
    n238_lo_n
  );


  or

  (
    g227_n,
    G358_o2_n_spl_00,
    n262_lo_n
  );


  and

  (
    g228_p,
    g225_n,
    n226_lo_p
  );


  and

  (
    g229_p,
    g228_p,
    g226_n
  );


  and

  (
    g230_p,
    g229_p,
    g227_n
  );


  and

  (
    g231_p,
    G213_o2_p_spl_00,
    n250_lo_p
  );


  and

  (
    g232_p,
    G318_o2_p_spl_00,
    n286_lo_p
  );


  and

  (
    g233_p,
    G358_o2_p_spl_00,
    n310_lo_p
  );


  or

  (
    g234_n,
    g232_p,
    g231_p
  );


  or

  (
    g235_n,
    g234_n,
    g233_p
  );


  or

  (
    g236_n,
    g235_n,
    n274_lo_n
  );


  and

  (
    g237_p,
    G213_o2_p_spl_00,
    n298_lo_p
  );


  or

  (
    g237_n,
    G213_o2_n_spl_00,
    n298_lo_n
  );


  and

  (
    g238_p,
    G318_o2_p_spl_00,
    n334_lo_p
  );


  or

  (
    g238_n,
    G318_o2_n_spl_00,
    n334_lo_n
  );


  and

  (
    g239_p,
    G358_o2_p_spl_00,
    n358_lo_p
  );


  or

  (
    g239_n,
    G358_o2_n_spl_00,
    n358_lo_n
  );


  and

  (
    g240_p,
    g238_n,
    g237_n
  );


  or

  (
    g240_n,
    g238_p,
    g237_p
  );


  and

  (
    g241_p,
    g240_p,
    g239_n
  );


  or

  (
    g241_n,
    g240_n,
    g239_p
  );


  and

  (
    g242_p,
    g241_p,
    n322_lo_p
  );


  or

  (
    g242_n,
    g241_n,
    n322_lo_n
  );


  and

  (
    g243_p,
    G213_o2_p_spl_01,
    n346_lo_p
  );


  or

  (
    g243_n,
    G213_o2_n_spl_0,
    n346_lo_n
  );


  and

  (
    g244_p,
    G318_o2_p_spl_01,
    n382_lo_p
  );


  or

  (
    g244_n,
    G318_o2_n_spl_0,
    n382_lo_n
  );


  and

  (
    g245_p,
    G358_o2_p_spl_01,
    n406_lo_p
  );


  or

  (
    g245_n,
    G358_o2_n_spl_0,
    n406_lo_n
  );


  and

  (
    g246_p,
    g244_n,
    g243_n
  );


  or

  (
    g246_n,
    g244_p,
    g243_p
  );


  and

  (
    g247_p,
    g246_p,
    g245_n
  );


  or

  (
    g247_n,
    g246_n,
    g245_p
  );


  and

  (
    g248_p,
    g247_p,
    n370_lo_p
  );


  or

  (
    g248_n,
    g247_n,
    n370_lo_n
  );


  and

  (
    g249_p,
    G213_o2_p_spl_01,
    n394_lo_p
  );


  or

  (
    g249_n,
    G213_o2_n_spl_1,
    n394_lo_n
  );


  and

  (
    g250_p,
    G318_o2_p_spl_01,
    n430_lo_p
  );


  or

  (
    g250_n,
    G318_o2_n_spl_1,
    n430_lo_n
  );


  and

  (
    g251_p,
    G358_o2_p_spl_01,
    n454_lo_p
  );


  or

  (
    g251_n,
    G358_o2_n_spl_1,
    n454_lo_n
  );


  and

  (
    g252_p,
    g250_n,
    g249_n
  );


  or

  (
    g252_n,
    g250_p,
    g249_p
  );


  and

  (
    g253_p,
    g252_p,
    g251_n
  );


  or

  (
    g253_n,
    g252_n,
    g251_p
  );


  and

  (
    g254_p,
    g253_p,
    n418_lo_p
  );


  or

  (
    g254_n,
    g253_n,
    n418_lo_n
  );


  and

  (
    g255_p,
    G213_o2_p_spl_10,
    n442_lo_p
  );


  and

  (
    g256_p,
    G318_o2_p_spl_10,
    n478_lo_p
  );


  and

  (
    g257_p,
    G358_o2_p_spl_10,
    n502_lo_p
  );


  or

  (
    g258_n,
    g256_p,
    g255_p
  );


  or

  (
    g259_n,
    g258_n,
    g257_p
  );


  or

  (
    g260_n,
    g259_n,
    n466_lo_n
  );


  and

  (
    g261_p,
    G213_o2_p_spl_10,
    n490_lo_p
  );


  or

  (
    g261_n,
    G213_o2_n_spl_1,
    n490_lo_n
  );


  and

  (
    g262_p,
    G318_o2_p_spl_10,
    n526_lo_p
  );


  or

  (
    g262_n,
    G318_o2_n_spl_1,
    n526_lo_n
  );


  and

  (
    g263_p,
    G358_o2_p_spl_10,
    n550_lo_p
  );


  or

  (
    g263_n,
    G358_o2_n_spl_1,
    n550_lo_n
  );


  and

  (
    g264_p,
    g262_n,
    g261_n
  );


  or

  (
    g264_n,
    g262_p,
    g261_p
  );


  and

  (
    g265_p,
    g264_p,
    g263_n
  );


  or

  (
    g265_n,
    g264_n,
    g263_p
  );


  and

  (
    g266_p,
    g265_p,
    n514_lo_p
  );


  or

  (
    g266_n,
    g265_n,
    n514_lo_n
  );


  and

  (
    g267_p,
    G213_o2_p_spl_11,
    n538_lo_p
  );


  and

  (
    g268_p,
    G318_o2_p_spl_11,
    n574_lo_p
  );


  and

  (
    g269_p,
    G358_o2_p_spl_11,
    n598_lo_p
  );


  or

  (
    g270_n,
    g268_p,
    g267_p
  );


  or

  (
    g271_n,
    g270_n,
    g269_p
  );


  or

  (
    g272_n,
    g271_n,
    n562_lo_n
  );


  and

  (
    g273_p,
    G213_o2_p_spl_11,
    n586_lo_p
  );


  and

  (
    g274_p,
    G318_o2_p_spl_11,
    n622_lo_p
  );


  and

  (
    g275_p,
    G358_o2_p_spl_11,
    n634_lo_p
  );


  or

  (
    g276_n,
    g274_p,
    g273_p
  );


  or

  (
    g277_n,
    g276_n,
    g275_p
  );


  or

  (
    g278_n,
    g277_n,
    n610_lo_n
  );


  and

  (
    g279_p,
    g242_n,
    g236_n_spl_
  );


  and

  (
    g280_p,
    g279_p_spl_0,
    g248_n_spl_
  );


  and

  (
    g281_p,
    g280_p,
    g254_n_spl_
  );


  and

  (
    g282_p,
    g281_p,
    g260_n_spl_
  );


  and

  (
    g283_p,
    g282_p,
    g266_n_spl_
  );


  and

  (
    g284_p,
    g283_p,
    g272_n_spl_
  );


  and

  (
    g285_p,
    g284_p,
    g278_n
  );


  or

  (
    g286_n,
    g285_p,
    g230_p
  );


  or

  (
    g287_n,
    g248_n_spl_,
    g242_p_spl_
  );


  and

  (
    g288_p,
    g287_n_spl_,
    g279_p_spl_0
  );


  and

  (
    g289_p,
    g288_p,
    g254_n_spl_
  );


  or

  (
    g290_n,
    g248_p_spl_,
    g242_p_spl_
  );


  or

  (
    g291_n,
    g290_n_spl_,
    g260_n_spl_
  );


  or

  (
    g292_n,
    g291_n,
    g254_p_spl_
  );


  or

  (
    g293_n,
    g254_p_spl_,
    g248_p_spl_
  );


  or

  (
    g294_n,
    g293_n,
    g266_n_spl_
  );


  and

  (
    g295_p,
    g292_n_spl_,
    g279_p_spl_
  );


  and

  (
    g296_p,
    g295_p,
    g294_n
  );


  or

  (
    g297_n,
    g290_n_spl_,
    g266_p
  );


  or

  (
    g298_n,
    g297_n,
    g272_n_spl_
  );


  and

  (
    g299_p,
    g287_n_spl_,
    g236_n_spl_
  );


  and

  (
    g300_p,
    g299_p,
    g292_n_spl_
  );


  and

  (
    g301_p,
    g300_p,
    g298_n
  );


  and

  (
    g302_p,
    G159_o2_n_spl_,
    G154_o2_n_spl_
  );


  or

  (
    g302_n,
    G159_o2_p_spl_,
    G154_o2_p_spl_
  );


  and

  (
    g303_p,
    g302_p,
    G162_o2_n_spl_
  );


  or

  (
    g303_n,
    g302_n,
    G162_o2_p_spl_
  );


  and

  (
    g304_p,
    g303_p,
    G165_o2_n_spl_
  );


  or

  (
    g304_n,
    g303_n,
    G165_o2_p_spl_
  );


  and

  (
    g305_p,
    g304_p,
    G168_o2_n_spl_
  );


  or

  (
    g305_n,
    g304_n,
    G168_o2_p_spl_
  );


  and

  (
    g306_p,
    g305_p,
    G171_o2_n_spl_
  );


  or

  (
    g306_n,
    g305_n,
    G171_o2_p_spl_
  );


  and

  (
    g307_p,
    g306_p,
    G174_o2_n_spl_
  );


  or

  (
    g307_n,
    g306_n,
    G174_o2_p_spl_
  );


  and

  (
    g308_p,
    g307_p,
    G177_o2_n_spl_
  );


  or

  (
    g308_n,
    g307_n,
    G177_o2_p_spl_
  );


  and

  (
    g309_p,
    g308_p,
    G180_o2_n_spl_
  );


  or

  (
    g309_n,
    g308_n,
    G180_o2_p_spl_
  );


  and

  (
    g310_p,
    n580_inv_n_spl_000,
    G259_o2_n
  );


  and

  (
    g311_p,
    n580_inv_p_spl_000,
    G259_o2_p
  );


  or

  (
    g312_n,
    g311_p,
    g310_p
  );


  and

  (
    g313_p,
    G158_o2_p,
    G223_o2_n
  );


  and

  (
    g314_p,
    g313_p,
    g312_n
  );


  and

  (
    g315_p,
    n580_inv_n_spl_000,
    G263_o2_n
  );


  and

  (
    g316_p,
    n580_inv_p_spl_000,
    G263_o2_p
  );


  or

  (
    g317_n,
    g316_p,
    g315_p
  );


  and

  (
    g318_p,
    G184_o2_p,
    G226_o2_n
  );


  and

  (
    g319_p,
    g318_p,
    g317_n
  );


  and

  (
    g320_p,
    n580_inv_n_spl_00,
    G266_o2_n
  );


  and

  (
    g321_p,
    n580_inv_p_spl_001,
    G266_o2_p
  );


  or

  (
    g322_n,
    g321_p,
    g320_p
  );


  and

  (
    g323_p,
    G186_o2_p,
    G229_o2_n
  );


  and

  (
    g324_p,
    g323_p,
    g322_n
  );


  and

  (
    g325_p,
    n580_inv_n_spl_01,
    G269_o2_n
  );


  and

  (
    g326_p,
    n580_inv_p_spl_001,
    G269_o2_p
  );


  or

  (
    g327_n,
    g326_p,
    g325_p
  );


  and

  (
    g328_p,
    G188_o2_p,
    G232_o2_n
  );


  and

  (
    g329_p,
    g328_p,
    g327_n
  );


  and

  (
    g330_p,
    n580_inv_n_spl_01,
    G272_o2_n
  );


  and

  (
    g331_p,
    n580_inv_p_spl_010,
    G272_o2_p
  );


  or

  (
    g332_n,
    g331_p,
    g330_p
  );


  and

  (
    g333_p,
    G190_o2_p,
    G235_o2_n
  );


  and

  (
    g334_p,
    g333_p,
    g332_n
  );


  and

  (
    g335_p,
    n580_inv_n_spl_10,
    G275_o2_n
  );


  and

  (
    g336_p,
    n580_inv_p_spl_010,
    G275_o2_p
  );


  or

  (
    g337_n,
    g336_p,
    g335_p
  );


  and

  (
    g338_p,
    G192_o2_p,
    G238_o2_n
  );


  and

  (
    g339_p,
    g338_p,
    g337_n
  );


  and

  (
    g340_p,
    n580_inv_n_spl_10,
    G278_o2_n
  );


  and

  (
    g341_p,
    n580_inv_p_spl_01,
    G278_o2_p
  );


  or

  (
    g342_n,
    g341_p,
    g340_p
  );


  and

  (
    g343_p,
    G194_o2_p,
    G242_o2_n
  );


  and

  (
    g344_p,
    g343_p,
    g342_n
  );


  and

  (
    g345_p,
    n580_inv_n_spl_11,
    G281_o2_n
  );


  and

  (
    g346_p,
    n580_inv_p_spl_10,
    G281_o2_p
  );


  or

  (
    g347_n,
    g346_p,
    g345_p
  );


  and

  (
    g348_p,
    G196_o2_p,
    G246_o2_n
  );


  and

  (
    g349_p,
    g348_p,
    g347_n
  );


  and

  (
    g350_p,
    n580_inv_n_spl_11,
    G284_o2_n
  );


  and

  (
    g351_p,
    n580_inv_p_spl_10,
    G284_o2_p
  );


  or

  (
    g352_n,
    g351_p,
    g350_p
  );


  and

  (
    g353_p,
    G198_o2_p,
    G250_o2_n
  );


  and

  (
    g354_p,
    g353_p,
    g352_n
  );


  or

  (
    g355_n,
    g319_p,
    g314_p
  );


  or

  (
    g356_n,
    g355_n,
    g324_p
  );


  or

  (
    g357_n,
    g356_n,
    g329_p
  );


  or

  (
    g358_n,
    g357_n,
    g334_p
  );


  or

  (
    g359_n,
    g358_n,
    g339_p
  );


  or

  (
    g360_n,
    g359_n,
    g344_p
  );


  or

  (
    g361_n,
    g360_n,
    g349_p
  );


  or

  (
    g362_n,
    g361_n,
    g354_p
  );


  and

  (
    g363_p,
    g309_p_spl_000,
    G154_o2_n_spl_
  );


  and

  (
    g364_p,
    g309_n_spl_000,
    G154_o2_p_spl_
  );


  or

  (
    g365_n,
    g364_p,
    g363_p
  );


  and

  (
    g366_p,
    g309_p_spl_000,
    G159_o2_n_spl_
  );


  and

  (
    g367_p,
    g309_n_spl_000,
    G159_o2_p_spl_
  );


  or

  (
    g368_n,
    g367_p,
    g366_p
  );


  and

  (
    g369_p,
    g309_p_spl_00,
    G162_o2_n_spl_
  );


  and

  (
    g370_p,
    g309_n_spl_001,
    G162_o2_p_spl_
  );


  or

  (
    g371_n,
    g370_p,
    g369_p
  );


  and

  (
    g372_p,
    g309_p_spl_01,
    G165_o2_n_spl_
  );


  and

  (
    g373_p,
    g309_n_spl_001,
    G165_o2_p_spl_
  );


  or

  (
    g374_n,
    g373_p,
    g372_p
  );


  and

  (
    g375_p,
    g309_p_spl_01,
    G168_o2_n_spl_
  );


  and

  (
    g376_p,
    g309_n_spl_01,
    G168_o2_p_spl_
  );


  or

  (
    g377_n,
    g376_p,
    g375_p
  );


  and

  (
    g378_p,
    g309_p_spl_10,
    G171_o2_n_spl_
  );


  and

  (
    g379_p,
    g309_n_spl_01,
    G171_o2_p_spl_
  );


  or

  (
    g380_n,
    g379_p,
    g378_p
  );


  and

  (
    g381_p,
    g309_p_spl_10,
    G174_o2_n_spl_
  );


  and

  (
    g382_p,
    g309_n_spl_10,
    G174_o2_p_spl_
  );


  or

  (
    g383_n,
    g382_p,
    g381_p
  );


  and

  (
    g384_p,
    g309_p_spl_11,
    G177_o2_n_spl_
  );


  and

  (
    g385_p,
    g309_n_spl_10,
    G177_o2_p_spl_
  );


  or

  (
    g386_n,
    g385_p,
    g384_p
  );


  and

  (
    g387_p,
    g309_p_spl_11,
    G180_o2_n_spl_
  );


  and

  (
    g388_p,
    g309_n_spl_11,
    G180_o2_p_spl_
  );


  or

  (
    g389_n,
    g388_p,
    g387_p
  );


  and

  (
    g390_p,
    n223_lo_buf_o2_p_spl_0,
    n232_lo_n
  );


  and

  (
    g391_p,
    g390_p,
    g365_n_spl_
  );


  and

  (
    g392_p,
    n271_lo_buf_o2_p_spl_0,
    n280_lo_n
  );


  and

  (
    g393_p,
    g392_p,
    g368_n_spl_
  );


  and

  (
    g394_p,
    n319_lo_buf_o2_p_spl_0,
    n328_lo_n
  );


  and

  (
    g395_p,
    g394_p,
    g371_n_spl_
  );


  and

  (
    g396_p,
    n367_lo_buf_o2_p_spl_0,
    n376_lo_n
  );


  and

  (
    g397_p,
    g396_p,
    g374_n_spl_
  );


  and

  (
    g398_p,
    n415_lo_buf_o2_p_spl_0,
    n424_lo_n
  );


  and

  (
    g399_p,
    g398_p,
    g377_n_spl_
  );


  and

  (
    g400_p,
    n463_lo_buf_o2_p_spl_0,
    n472_lo_n
  );


  and

  (
    g401_p,
    g400_p,
    g380_n_spl_
  );


  and

  (
    g402_p,
    n511_lo_buf_o2_p_spl_0,
    n520_lo_n
  );


  and

  (
    g403_p,
    g402_p,
    g383_n_spl_
  );


  and

  (
    g404_p,
    n559_lo_buf_o2_p_spl_0,
    n568_lo_n
  );


  and

  (
    g405_p,
    g404_p,
    g386_n_spl_
  );


  and

  (
    g406_p,
    n607_lo_buf_o2_p_spl_0,
    n616_lo_n
  );


  and

  (
    g407_p,
    g406_p,
    g389_n_spl_
  );


  and

  (
    g408_p,
    n223_lo_buf_o2_p_spl_0,
    n256_lo_n
  );


  and

  (
    g409_p,
    n271_lo_buf_o2_p_spl_0,
    n304_lo_n
  );


  and

  (
    g410_p,
    n319_lo_buf_o2_p_spl_0,
    n352_lo_n
  );


  and

  (
    g411_p,
    n367_lo_buf_o2_p_spl_0,
    n400_lo_n
  );


  and

  (
    g412_p,
    n415_lo_buf_o2_p_spl_0,
    n448_lo_n
  );


  and

  (
    g413_p,
    n463_lo_buf_o2_p_spl_0,
    n496_lo_n
  );


  and

  (
    g414_p,
    n511_lo_buf_o2_p_spl_0,
    n544_lo_n
  );


  and

  (
    g415_p,
    n559_lo_buf_o2_p_spl_0,
    n592_lo_n
  );


  and

  (
    g416_p,
    n607_lo_buf_o2_p_spl_0,
    n628_lo_n
  );


  or

  (
    g417_n,
    g393_p_spl_,
    g391_p_spl_
  );


  or

  (
    g418_n,
    g417_n,
    g395_p_spl_
  );


  or

  (
    g419_n,
    g418_n,
    g397_p_spl_
  );


  or

  (
    g420_n,
    g419_n,
    g399_p_spl_
  );


  or

  (
    g421_n,
    g420_n,
    g401_p_spl_
  );


  or

  (
    g422_n,
    g421_n,
    g403_p_spl_
  );


  or

  (
    g423_n,
    g422_n,
    g405_p_spl_
  );


  or

  (
    g424_n,
    g423_n,
    g407_p_spl_
  );


  and

  (
    g425_p,
    n217_lo_p_spl_,
    n205_lo_n
  );


  and

  (
    g426_p,
    n265_lo_p_spl_,
    n241_lo_n
  );


  and

  (
    g427_p,
    n313_lo_p_spl_,
    n289_lo_n
  );


  and

  (
    g428_p,
    n361_lo_p_spl_,
    n337_lo_n
  );


  and

  (
    g429_p,
    n409_lo_p_spl_,
    n385_lo_n
  );


  and

  (
    g430_p,
    n457_lo_p_spl_,
    n433_lo_n
  );


  and

  (
    g431_p,
    n505_lo_p_spl_,
    n481_lo_n
  );


  and

  (
    g432_p,
    n553_lo_p_spl_,
    n529_lo_n
  );


  and

  (
    g433_p,
    n601_lo_p_spl_,
    n577_lo_n
  );


  buf

  (
    G426,
    n316_inv_p
  );


  buf

  (
    G427,
    n319_inv_p
  );


  buf

  (
    G428,
    n406_1_inv_p
  );


  not

  (
    G429,
    g286_n
  );


  not

  (
    G430,
    g289_p
  );


  not

  (
    G431,
    g296_p
  );


  not

  (
    G432,
    g301_p
  );


  buf

  (
    n205_li,
    G1_p
  );


  buf

  (
    n214_li,
    n997_o2_p
  );


  buf

  (
    n217_li,
    G2_p
  );


  buf

  (
    n226_li,
    n1015_o2_p
  );


  buf

  (
    n229_li,
    G3_p
  );


  buf

  (
    n232_li,
    n229_lo_p
  );


  buf

  (
    n238_li,
    n235_lo_buf_o2_p
  );


  buf

  (
    n241_li,
    G4_p
  );


  buf

  (
    n250_li,
    n998_o2_p
  );


  buf

  (
    n253_li,
    G5_p
  );


  buf

  (
    n256_li,
    n253_lo_p
  );


  buf

  (
    n262_li,
    n259_lo_buf_o2_p
  );


  buf

  (
    n265_li,
    G6_p
  );


  buf

  (
    n274_li,
    n1016_o2_p
  );


  buf

  (
    n277_li,
    G7_p
  );


  buf

  (
    n280_li,
    n277_lo_p
  );


  buf

  (
    n286_li,
    n283_lo_buf_o2_p
  );


  buf

  (
    n289_li,
    G8_p
  );


  buf

  (
    n298_li,
    n999_o2_p
  );


  buf

  (
    n301_li,
    G9_p
  );


  buf

  (
    n304_li,
    n301_lo_p
  );


  buf

  (
    n310_li,
    n307_lo_buf_o2_p
  );


  buf

  (
    n313_li,
    G10_p
  );


  buf

  (
    n322_li,
    n1017_o2_p
  );


  buf

  (
    n325_li,
    G11_p
  );


  buf

  (
    n328_li,
    n325_lo_p
  );


  buf

  (
    n334_li,
    n331_lo_buf_o2_p
  );


  buf

  (
    n337_li,
    G12_p
  );


  buf

  (
    n346_li,
    n1000_o2_p
  );


  buf

  (
    n349_li,
    G13_p
  );


  buf

  (
    n352_li,
    n349_lo_p
  );


  buf

  (
    n358_li,
    n355_lo_buf_o2_p
  );


  buf

  (
    n361_li,
    G14_p
  );


  buf

  (
    n370_li,
    n1018_o2_p
  );


  buf

  (
    n373_li,
    G15_p
  );


  buf

  (
    n376_li,
    n373_lo_p
  );


  buf

  (
    n382_li,
    n379_lo_buf_o2_p
  );


  buf

  (
    n385_li,
    G16_p
  );


  buf

  (
    n394_li,
    n1001_o2_p
  );


  buf

  (
    n397_li,
    G17_p
  );


  buf

  (
    n400_li,
    n397_lo_p
  );


  buf

  (
    n406_li,
    n403_lo_buf_o2_p
  );


  buf

  (
    n409_li,
    G18_p
  );


  buf

  (
    n418_li,
    n1019_o2_p
  );


  buf

  (
    n421_li,
    G19_p
  );


  buf

  (
    n424_li,
    n421_lo_p
  );


  buf

  (
    n430_li,
    n427_lo_buf_o2_p
  );


  buf

  (
    n433_li,
    G20_p
  );


  buf

  (
    n442_li,
    n1002_o2_p
  );


  buf

  (
    n445_li,
    G21_p
  );


  buf

  (
    n448_li,
    n445_lo_p
  );


  buf

  (
    n454_li,
    n451_lo_buf_o2_p
  );


  buf

  (
    n457_li,
    G22_p
  );


  buf

  (
    n466_li,
    n1020_o2_p
  );


  buf

  (
    n469_li,
    G23_p
  );


  buf

  (
    n472_li,
    n469_lo_p
  );


  buf

  (
    n478_li,
    n475_lo_buf_o2_p
  );


  buf

  (
    n481_li,
    G24_p
  );


  buf

  (
    n490_li,
    n1003_o2_p
  );


  buf

  (
    n493_li,
    G25_p
  );


  buf

  (
    n496_li,
    n493_lo_p
  );


  buf

  (
    n502_li,
    n499_lo_buf_o2_p
  );


  buf

  (
    n505_li,
    G26_p
  );


  buf

  (
    n514_li,
    n1021_o2_p
  );


  buf

  (
    n517_li,
    G27_p
  );


  buf

  (
    n520_li,
    n517_lo_p
  );


  buf

  (
    n526_li,
    n523_lo_buf_o2_p
  );


  buf

  (
    n529_li,
    G28_p
  );


  buf

  (
    n538_li,
    n1004_o2_p
  );


  buf

  (
    n541_li,
    G29_p
  );


  buf

  (
    n544_li,
    n541_lo_p
  );


  buf

  (
    n550_li,
    n547_lo_buf_o2_p
  );


  buf

  (
    n553_li,
    G30_p
  );


  buf

  (
    n562_li,
    n1022_o2_p
  );


  buf

  (
    n565_li,
    G31_p
  );


  buf

  (
    n568_li,
    n565_lo_p
  );


  buf

  (
    n574_li,
    n571_lo_buf_o2_p
  );


  buf

  (
    n577_li,
    G32_p
  );


  buf

  (
    n586_li,
    n1005_o2_p
  );


  buf

  (
    n589_li,
    G33_p
  );


  buf

  (
    n592_li,
    n589_lo_p
  );


  buf

  (
    n598_li,
    n595_lo_buf_o2_p
  );


  buf

  (
    n601_li,
    G34_p
  );


  buf

  (
    n610_li,
    n1023_o2_p
  );


  buf

  (
    n613_li,
    G35_p
  );


  buf

  (
    n616_li,
    n613_lo_p
  );


  buf

  (
    n622_li,
    n619_lo_buf_o2_p
  );


  buf

  (
    n625_li,
    G36_p
  );


  buf

  (
    n628_li,
    n625_lo_p
  );


  buf

  (
    n634_li,
    n631_lo_buf_o2_p
  );


  buf

  (
    n919_i2,
    n376_1_inv_p_spl_
  );


  buf

  (
    n1024_i2,
    n580_inv_p_spl_11
  );


  buf

  (
    n997_i2,
    n211_lo_buf_o2_p
  );


  buf

  (
    n998_i2,
    n247_lo_buf_o2_p
  );


  buf

  (
    n999_i2,
    n295_lo_buf_o2_p
  );


  buf

  (
    n1000_i2,
    n343_lo_buf_o2_p
  );


  buf

  (
    n1001_i2,
    n391_lo_buf_o2_p
  );


  buf

  (
    n1002_i2,
    n439_lo_buf_o2_p
  );


  buf

  (
    n1003_i2,
    n487_lo_buf_o2_p
  );


  buf

  (
    n1004_i2,
    n535_lo_buf_o2_p
  );


  buf

  (
    n1005_i2,
    n583_lo_buf_o2_p
  );


  buf

  (
    n1015_i2,
    n223_lo_buf_o2_p_spl_
  );


  buf

  (
    n1016_i2,
    n271_lo_buf_o2_p_spl_
  );


  buf

  (
    n1017_i2,
    n319_lo_buf_o2_p_spl_
  );


  buf

  (
    n1018_i2,
    n367_lo_buf_o2_p_spl_
  );


  buf

  (
    n1019_i2,
    n415_lo_buf_o2_p_spl_
  );


  buf

  (
    n1020_i2,
    n463_lo_buf_o2_p_spl_
  );


  buf

  (
    n1021_i2,
    n511_lo_buf_o2_p_spl_
  );


  buf

  (
    n1022_i2,
    n559_lo_buf_o2_p_spl_
  );


  buf

  (
    n1023_i2,
    n607_lo_buf_o2_p_spl_
  );


  buf

  (
    G199_i2,
    g309_n_spl_11
  );


  buf

  (
    n235_lo_buf_i2,
    n232_lo_p
  );


  buf

  (
    n283_lo_buf_i2,
    n280_lo_p
  );


  buf

  (
    n331_lo_buf_i2,
    n328_lo_p
  );


  buf

  (
    n379_lo_buf_i2,
    n376_lo_p
  );


  buf

  (
    n427_lo_buf_i2,
    n424_lo_p
  );


  buf

  (
    n475_lo_buf_i2,
    n472_lo_p
  );


  buf

  (
    n523_lo_buf_i2,
    n520_lo_p
  );


  buf

  (
    n571_lo_buf_i2,
    n568_lo_p
  );


  buf

  (
    n619_lo_buf_i2,
    n616_lo_p
  );


  buf

  (
    G355_i2,
    g362_n_spl_
  );


  not

  (
    G223_i2,
    g365_n_spl_
  );


  not

  (
    G226_i2,
    g368_n_spl_
  );


  not

  (
    G229_i2,
    g371_n_spl_
  );


  not

  (
    G232_i2,
    g374_n_spl_
  );


  not

  (
    G235_i2,
    g377_n_spl_
  );


  not

  (
    G238_i2,
    g380_n_spl_
  );


  not

  (
    G242_i2,
    g383_n_spl_
  );


  not

  (
    G246_i2,
    g386_n_spl_
  );


  not

  (
    G250_i2,
    g389_n_spl_
  );


  buf

  (
    n259_lo_buf_i2,
    n256_lo_p
  );


  buf

  (
    n307_lo_buf_i2,
    n304_lo_p
  );


  buf

  (
    n355_lo_buf_i2,
    n352_lo_p
  );


  buf

  (
    n403_lo_buf_i2,
    n400_lo_p
  );


  buf

  (
    n451_lo_buf_i2,
    n448_lo_p
  );


  buf

  (
    n499_lo_buf_i2,
    n496_lo_p
  );


  buf

  (
    n547_lo_buf_i2,
    n544_lo_p
  );


  buf

  (
    n595_lo_buf_i2,
    n592_lo_p
  );


  buf

  (
    n631_lo_buf_i2,
    n628_lo_p
  );


  buf

  (
    G213_i2,
    n376_1_inv_p_spl_
  );


  buf

  (
    G318_i2,
    n580_inv_p_spl_11
  );


  buf

  (
    G358_i2,
    g362_n_spl_
  );


  buf

  (
    G259_i2,
    g391_p_spl_
  );


  buf

  (
    G263_i2,
    g393_p_spl_
  );


  buf

  (
    G266_i2,
    g395_p_spl_
  );


  buf

  (
    G269_i2,
    g397_p_spl_
  );


  buf

  (
    G272_i2,
    g399_p_spl_
  );


  buf

  (
    G275_i2,
    g401_p_spl_
  );


  buf

  (
    G278_i2,
    g403_p_spl_
  );


  buf

  (
    G281_i2,
    g405_p_spl_
  );


  buf

  (
    G284_i2,
    g407_p_spl_
  );


  buf

  (
    n211_lo_buf_i2,
    n205_lo_p
  );


  buf

  (
    n247_lo_buf_i2,
    n241_lo_p
  );


  buf

  (
    n295_lo_buf_i2,
    n289_lo_p
  );


  buf

  (
    n343_lo_buf_i2,
    n337_lo_p
  );


  buf

  (
    n391_lo_buf_i2,
    n385_lo_p
  );


  buf

  (
    n439_lo_buf_i2,
    n433_lo_p
  );


  buf

  (
    n487_lo_buf_i2,
    n481_lo_p
  );


  buf

  (
    n535_lo_buf_i2,
    n529_lo_p
  );


  buf

  (
    n583_lo_buf_i2,
    n577_lo_p
  );


  buf

  (
    G158_i2,
    g408_p
  );


  buf

  (
    G184_i2,
    g409_p
  );


  buf

  (
    G186_i2,
    g410_p
  );


  buf

  (
    G188_i2,
    g411_p
  );


  buf

  (
    G190_i2,
    g412_p
  );


  buf

  (
    G192_i2,
    g413_p
  );


  buf

  (
    G194_i2,
    g414_p
  );


  buf

  (
    G196_i2,
    g415_p
  );


  buf

  (
    G198_i2,
    g416_p
  );


  buf

  (
    n223_lo_buf_i2,
    n217_lo_p_spl_
  );


  buf

  (
    n271_lo_buf_i2,
    n265_lo_p_spl_
  );


  buf

  (
    n319_lo_buf_i2,
    n313_lo_p_spl_
  );


  buf

  (
    n367_lo_buf_i2,
    n361_lo_p_spl_
  );


  buf

  (
    n415_lo_buf_i2,
    n409_lo_p_spl_
  );


  buf

  (
    n463_lo_buf_i2,
    n457_lo_p_spl_
  );


  buf

  (
    n511_lo_buf_i2,
    n505_lo_p_spl_
  );


  buf

  (
    n559_lo_buf_i2,
    n553_lo_p_spl_
  );


  buf

  (
    n607_lo_buf_i2,
    n601_lo_p_spl_
  );


  buf

  (
    G295_i2,
    g424_n
  );


  buf

  (
    G154_i2,
    g425_p
  );


  buf

  (
    G159_i2,
    g426_p
  );


  buf

  (
    G162_i2,
    g427_p
  );


  buf

  (
    G165_i2,
    g428_p
  );


  buf

  (
    G168_i2,
    g429_p
  );


  buf

  (
    G171_i2,
    g430_p
  );


  buf

  (
    G174_i2,
    g431_p
  );


  buf

  (
    G177_i2,
    g432_p
  );


  buf

  (
    G180_i2,
    g433_p
  );


  buf

  (
    G213_o2_n_spl_,
    G213_o2_n
  );


  buf

  (
    G213_o2_n_spl_0,
    G213_o2_n_spl_
  );


  buf

  (
    G213_o2_n_spl_00,
    G213_o2_n_spl_0
  );


  buf

  (
    G213_o2_n_spl_1,
    G213_o2_n_spl_
  );


  buf

  (
    G318_o2_n_spl_,
    G318_o2_n
  );


  buf

  (
    G318_o2_n_spl_0,
    G318_o2_n_spl_
  );


  buf

  (
    G318_o2_n_spl_00,
    G318_o2_n_spl_0
  );


  buf

  (
    G318_o2_n_spl_1,
    G318_o2_n_spl_
  );


  buf

  (
    G358_o2_n_spl_,
    G358_o2_n
  );


  buf

  (
    G358_o2_n_spl_0,
    G358_o2_n_spl_
  );


  buf

  (
    G358_o2_n_spl_00,
    G358_o2_n_spl_0
  );


  buf

  (
    G358_o2_n_spl_1,
    G358_o2_n_spl_
  );


  buf

  (
    G213_o2_p_spl_,
    G213_o2_p
  );


  buf

  (
    G213_o2_p_spl_0,
    G213_o2_p_spl_
  );


  buf

  (
    G213_o2_p_spl_00,
    G213_o2_p_spl_0
  );


  buf

  (
    G213_o2_p_spl_01,
    G213_o2_p_spl_0
  );


  buf

  (
    G213_o2_p_spl_1,
    G213_o2_p_spl_
  );


  buf

  (
    G213_o2_p_spl_10,
    G213_o2_p_spl_1
  );


  buf

  (
    G213_o2_p_spl_11,
    G213_o2_p_spl_1
  );


  buf

  (
    G318_o2_p_spl_,
    G318_o2_p
  );


  buf

  (
    G318_o2_p_spl_0,
    G318_o2_p_spl_
  );


  buf

  (
    G318_o2_p_spl_00,
    G318_o2_p_spl_0
  );


  buf

  (
    G318_o2_p_spl_01,
    G318_o2_p_spl_0
  );


  buf

  (
    G318_o2_p_spl_1,
    G318_o2_p_spl_
  );


  buf

  (
    G318_o2_p_spl_10,
    G318_o2_p_spl_1
  );


  buf

  (
    G318_o2_p_spl_11,
    G318_o2_p_spl_1
  );


  buf

  (
    G358_o2_p_spl_,
    G358_o2_p
  );


  buf

  (
    G358_o2_p_spl_0,
    G358_o2_p_spl_
  );


  buf

  (
    G358_o2_p_spl_00,
    G358_o2_p_spl_0
  );


  buf

  (
    G358_o2_p_spl_01,
    G358_o2_p_spl_0
  );


  buf

  (
    G358_o2_p_spl_1,
    G358_o2_p_spl_
  );


  buf

  (
    G358_o2_p_spl_10,
    G358_o2_p_spl_1
  );


  buf

  (
    G358_o2_p_spl_11,
    G358_o2_p_spl_1
  );


  buf

  (
    g236_n_spl_,
    g236_n
  );


  buf

  (
    g279_p_spl_,
    g279_p
  );


  buf

  (
    g279_p_spl_0,
    g279_p_spl_
  );


  buf

  (
    g248_n_spl_,
    g248_n
  );


  buf

  (
    g254_n_spl_,
    g254_n
  );


  buf

  (
    g260_n_spl_,
    g260_n
  );


  buf

  (
    g266_n_spl_,
    g266_n
  );


  buf

  (
    g272_n_spl_,
    g272_n
  );


  buf

  (
    g242_p_spl_,
    g242_p
  );


  buf

  (
    g287_n_spl_,
    g287_n
  );


  buf

  (
    g248_p_spl_,
    g248_p
  );


  buf

  (
    g290_n_spl_,
    g290_n
  );


  buf

  (
    g254_p_spl_,
    g254_p
  );


  buf

  (
    g292_n_spl_,
    g292_n
  );


  buf

  (
    G159_o2_n_spl_,
    G159_o2_n
  );


  buf

  (
    G154_o2_n_spl_,
    G154_o2_n
  );


  buf

  (
    G159_o2_p_spl_,
    G159_o2_p
  );


  buf

  (
    G154_o2_p_spl_,
    G154_o2_p
  );


  buf

  (
    G162_o2_n_spl_,
    G162_o2_n
  );


  buf

  (
    G162_o2_p_spl_,
    G162_o2_p
  );


  buf

  (
    G165_o2_n_spl_,
    G165_o2_n
  );


  buf

  (
    G165_o2_p_spl_,
    G165_o2_p
  );


  buf

  (
    G168_o2_n_spl_,
    G168_o2_n
  );


  buf

  (
    G168_o2_p_spl_,
    G168_o2_p
  );


  buf

  (
    G171_o2_n_spl_,
    G171_o2_n
  );


  buf

  (
    G171_o2_p_spl_,
    G171_o2_p
  );


  buf

  (
    G174_o2_n_spl_,
    G174_o2_n
  );


  buf

  (
    G174_o2_p_spl_,
    G174_o2_p
  );


  buf

  (
    G177_o2_n_spl_,
    G177_o2_n
  );


  buf

  (
    G177_o2_p_spl_,
    G177_o2_p
  );


  buf

  (
    G180_o2_n_spl_,
    G180_o2_n
  );


  buf

  (
    G180_o2_p_spl_,
    G180_o2_p
  );


  buf

  (
    n580_inv_n_spl_,
    n580_inv_n
  );


  buf

  (
    n580_inv_n_spl_0,
    n580_inv_n_spl_
  );


  buf

  (
    n580_inv_n_spl_00,
    n580_inv_n_spl_0
  );


  buf

  (
    n580_inv_n_spl_000,
    n580_inv_n_spl_00
  );


  buf

  (
    n580_inv_n_spl_01,
    n580_inv_n_spl_0
  );


  buf

  (
    n580_inv_n_spl_1,
    n580_inv_n_spl_
  );


  buf

  (
    n580_inv_n_spl_10,
    n580_inv_n_spl_1
  );


  buf

  (
    n580_inv_n_spl_11,
    n580_inv_n_spl_1
  );


  buf

  (
    n580_inv_p_spl_,
    n580_inv_p
  );


  buf

  (
    n580_inv_p_spl_0,
    n580_inv_p_spl_
  );


  buf

  (
    n580_inv_p_spl_00,
    n580_inv_p_spl_0
  );


  buf

  (
    n580_inv_p_spl_000,
    n580_inv_p_spl_00
  );


  buf

  (
    n580_inv_p_spl_001,
    n580_inv_p_spl_00
  );


  buf

  (
    n580_inv_p_spl_01,
    n580_inv_p_spl_0
  );


  buf

  (
    n580_inv_p_spl_010,
    n580_inv_p_spl_01
  );


  buf

  (
    n580_inv_p_spl_1,
    n580_inv_p_spl_
  );


  buf

  (
    n580_inv_p_spl_10,
    n580_inv_p_spl_1
  );


  buf

  (
    n580_inv_p_spl_11,
    n580_inv_p_spl_1
  );


  buf

  (
    g309_p_spl_,
    g309_p
  );


  buf

  (
    g309_p_spl_0,
    g309_p_spl_
  );


  buf

  (
    g309_p_spl_00,
    g309_p_spl_0
  );


  buf

  (
    g309_p_spl_000,
    g309_p_spl_00
  );


  buf

  (
    g309_p_spl_01,
    g309_p_spl_0
  );


  buf

  (
    g309_p_spl_1,
    g309_p_spl_
  );


  buf

  (
    g309_p_spl_10,
    g309_p_spl_1
  );


  buf

  (
    g309_p_spl_11,
    g309_p_spl_1
  );


  buf

  (
    g309_n_spl_,
    g309_n
  );


  buf

  (
    g309_n_spl_0,
    g309_n_spl_
  );


  buf

  (
    g309_n_spl_00,
    g309_n_spl_0
  );


  buf

  (
    g309_n_spl_000,
    g309_n_spl_00
  );


  buf

  (
    g309_n_spl_001,
    g309_n_spl_00
  );


  buf

  (
    g309_n_spl_01,
    g309_n_spl_0
  );


  buf

  (
    g309_n_spl_1,
    g309_n_spl_
  );


  buf

  (
    g309_n_spl_10,
    g309_n_spl_1
  );


  buf

  (
    g309_n_spl_11,
    g309_n_spl_1
  );


  buf

  (
    n223_lo_buf_o2_p_spl_,
    n223_lo_buf_o2_p
  );


  buf

  (
    n223_lo_buf_o2_p_spl_0,
    n223_lo_buf_o2_p_spl_
  );


  buf

  (
    g365_n_spl_,
    g365_n
  );


  buf

  (
    n271_lo_buf_o2_p_spl_,
    n271_lo_buf_o2_p
  );


  buf

  (
    n271_lo_buf_o2_p_spl_0,
    n271_lo_buf_o2_p_spl_
  );


  buf

  (
    g368_n_spl_,
    g368_n
  );


  buf

  (
    n319_lo_buf_o2_p_spl_,
    n319_lo_buf_o2_p
  );


  buf

  (
    n319_lo_buf_o2_p_spl_0,
    n319_lo_buf_o2_p_spl_
  );


  buf

  (
    g371_n_spl_,
    g371_n
  );


  buf

  (
    n367_lo_buf_o2_p_spl_,
    n367_lo_buf_o2_p
  );


  buf

  (
    n367_lo_buf_o2_p_spl_0,
    n367_lo_buf_o2_p_spl_
  );


  buf

  (
    g374_n_spl_,
    g374_n
  );


  buf

  (
    n415_lo_buf_o2_p_spl_,
    n415_lo_buf_o2_p
  );


  buf

  (
    n415_lo_buf_o2_p_spl_0,
    n415_lo_buf_o2_p_spl_
  );


  buf

  (
    g377_n_spl_,
    g377_n
  );


  buf

  (
    n463_lo_buf_o2_p_spl_,
    n463_lo_buf_o2_p
  );


  buf

  (
    n463_lo_buf_o2_p_spl_0,
    n463_lo_buf_o2_p_spl_
  );


  buf

  (
    g380_n_spl_,
    g380_n
  );


  buf

  (
    n511_lo_buf_o2_p_spl_,
    n511_lo_buf_o2_p
  );


  buf

  (
    n511_lo_buf_o2_p_spl_0,
    n511_lo_buf_o2_p_spl_
  );


  buf

  (
    g383_n_spl_,
    g383_n
  );


  buf

  (
    n559_lo_buf_o2_p_spl_,
    n559_lo_buf_o2_p
  );


  buf

  (
    n559_lo_buf_o2_p_spl_0,
    n559_lo_buf_o2_p_spl_
  );


  buf

  (
    g386_n_spl_,
    g386_n
  );


  buf

  (
    n607_lo_buf_o2_p_spl_,
    n607_lo_buf_o2_p
  );


  buf

  (
    n607_lo_buf_o2_p_spl_0,
    n607_lo_buf_o2_p_spl_
  );


  buf

  (
    g389_n_spl_,
    g389_n
  );


  buf

  (
    g393_p_spl_,
    g393_p
  );


  buf

  (
    g391_p_spl_,
    g391_p
  );


  buf

  (
    g395_p_spl_,
    g395_p
  );


  buf

  (
    g397_p_spl_,
    g397_p
  );


  buf

  (
    g399_p_spl_,
    g399_p
  );


  buf

  (
    g401_p_spl_,
    g401_p
  );


  buf

  (
    g403_p_spl_,
    g403_p
  );


  buf

  (
    g405_p_spl_,
    g405_p
  );


  buf

  (
    g407_p_spl_,
    g407_p
  );


  buf

  (
    n217_lo_p_spl_,
    n217_lo_p
  );


  buf

  (
    n265_lo_p_spl_,
    n265_lo_p
  );


  buf

  (
    n313_lo_p_spl_,
    n313_lo_p
  );


  buf

  (
    n361_lo_p_spl_,
    n361_lo_p
  );


  buf

  (
    n409_lo_p_spl_,
    n409_lo_p
  );


  buf

  (
    n457_lo_p_spl_,
    n457_lo_p
  );


  buf

  (
    n505_lo_p_spl_,
    n505_lo_p
  );


  buf

  (
    n553_lo_p_spl_,
    n553_lo_p
  );


  buf

  (
    n601_lo_p_spl_,
    n601_lo_p
  );


  buf

  (
    n376_1_inv_p_spl_,
    n376_1_inv_p
  );


  buf

  (
    g362_n_spl_,
    g362_n
  );


endmodule
