// Benchmark "mymod" written by ABC on Sun Oct 29 19:31:59 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58,
    G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70, G71, G72,
    G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86,
    G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G109, G110, G111, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G124,
    G125, G126, G127, G128, G129, G130, G131, G132, G133, G134, G135, G136,
    G137, G138, G139, G140, G141, G142, G143, G144, G145, G146, G147, G148,
    G149, G150, G151, G152, G153, G154, G155, G156, G157, G158, G159, G160,
    G161, G162, G163, G164, G165, G166, G167, G168, G169, G170, G171, G172,
    G173, G174, G175, G176, G177, G178,
    G5193, G5194, G5195, G5196, G5197, G5198, G5199, G5200, G5201, G5202,
    G5203, G5204, G5205, G5206, G5207, G5208, G5209, G5210, G5211, G5212,
    G5213, G5214, G5215, G5216, G5217, G5218, G5219, G5220, G5221, G5222,
    G5223, G5224, G5225, G5226, G5227, G5228, G5229, G5230, G5231, G5232,
    G5233, G5234, G5235, G5236, G5237, G5238, G5239, G5240, G5241, G5242,
    G5243, G5244, G5245, G5246, G5247, G5248, G5249, G5250, G5251, G5252,
    G5253, G5254, G5255, G5256, G5257, G5258, G5259, G5260, G5261, G5262,
    G5263, G5264, G5265, G5266, G5267, G5268, G5269, G5270, G5271, G5272,
    G5273, G5274, G5275, G5276, G5277, G5278, G5279, G5280, G5281, G5282,
    G5283, G5284, G5285, G5286, G5287, G5288, G5289, G5290, G5291, G5292,
    G5293, G5294, G5295, G5296, G5297, G5298, G5299, G5300, G5301, G5302,
    G5303, G5304, G5305, G5306, G5307, G5308, G5309, G5310, G5311, G5312,
    G5313, G5314, G5315  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70,
    G71, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98,
    G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G110,
    G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G133, G134,
    G135, G136, G137, G138, G139, G140, G141, G142, G143, G144, G145, G146,
    G147, G148, G149, G150, G151, G152, G153, G154, G155, G156, G157, G158,
    G159, G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G170,
    G171, G172, G173, G174, G175, G176, G177, G178;
  output G5193, G5194, G5195, G5196, G5197, G5198, G5199, G5200, G5201, G5202,
    G5203, G5204, G5205, G5206, G5207, G5208, G5209, G5210, G5211, G5212,
    G5213, G5214, G5215, G5216, G5217, G5218, G5219, G5220, G5221, G5222,
    G5223, G5224, G5225, G5226, G5227, G5228, G5229, G5230, G5231, G5232,
    G5233, G5234, G5235, G5236, G5237, G5238, G5239, G5240, G5241, G5242,
    G5243, G5244, G5245, G5246, G5247, G5248, G5249, G5250, G5251, G5252,
    G5253, G5254, G5255, G5256, G5257, G5258, G5259, G5260, G5261, G5262,
    G5263, G5264, G5265, G5266, G5267, G5268, G5269, G5270, G5271, G5272,
    G5273, G5274, G5275, G5276, G5277, G5278, G5279, G5280, G5281, G5282,
    G5283, G5284, G5285, G5286, G5287, G5288, G5289, G5290, G5291, G5292,
    G5293, G5294, G5295, G5296, G5297, G5298, G5299, G5300, G5301, G5302,
    G5303, G5304, G5305, G5306, G5307, G5308, G5309, G5310, G5311, G5312,
    G5313, G5314, G5315;
  reg n2610_lo, n2613_lo, n2616_lo, n2619_lo, n2622_lo, n2625_lo, n2628_lo,
    n2631_lo, n2634_lo, n2637_lo, n2640_lo, n2643_lo, n2646_lo, n2649_lo,
    n2652_lo, n2655_lo, n2658_lo, n2661_lo, n2664_lo, n2667_lo, n2670_lo,
    n2673_lo, n2676_lo, n2679_lo, n2682_lo, n2685_lo, n2688_lo, n2691_lo,
    n2694_lo, n2697_lo, n2700_lo, n2703_lo, n2706_lo, n2709_lo, n2712_lo,
    n2715_lo, n2718_lo, n2721_lo, n2724_lo, n2727_lo, n2730_lo, n2733_lo,
    n2736_lo, n2739_lo, n2742_lo, n2745_lo, n2748_lo, n2751_lo, n2754_lo,
    n2757_lo, n2760_lo, n2763_lo, n2766_lo, n2769_lo, n2772_lo, n2775_lo,
    n2778_lo, n2781_lo, n2784_lo, n2787_lo, n2790_lo, n2793_lo, n2796_lo,
    n2799_lo, n2802_lo, n2805_lo, n2808_lo, n2811_lo, n2814_lo, n2817_lo,
    n2820_lo, n2823_lo, n2826_lo, n2829_lo, n2832_lo, n2835_lo, n2838_lo,
    n2841_lo, n2844_lo, n2847_lo, n2850_lo, n2853_lo, n2856_lo, n2859_lo,
    n2862_lo, n2865_lo, n2868_lo, n2871_lo, n2874_lo, n2877_lo, n2880_lo,
    n2883_lo, n2886_lo, n2889_lo, n2892_lo, n2895_lo, n2898_lo, n2901_lo,
    n2904_lo, n2907_lo, n2910_lo, n2913_lo, n2916_lo, n2919_lo, n2922_lo,
    n2925_lo, n2928_lo, n2931_lo, n2934_lo, n2937_lo, n2940_lo, n2943_lo,
    n2946_lo, n2949_lo, n2952_lo, n2955_lo, n2958_lo, n2961_lo, n2964_lo,
    n2967_lo, n2970_lo, n2973_lo, n2976_lo, n2979_lo, n2982_lo, n2985_lo,
    n2988_lo, n2991_lo, n2994_lo, n2997_lo, n3000_lo, n3003_lo, n3006_lo,
    n3009_lo, n3012_lo, n3015_lo, n3018_lo, n3021_lo, n3024_lo, n3027_lo,
    n3030_lo, n3033_lo, n3036_lo, n3039_lo, n3042_lo, n3045_lo, n3048_lo,
    n3051_lo, n3054_lo, n3057_lo, n3060_lo, n3063_lo, n3066_lo, n3069_lo,
    n3072_lo, n3075_lo, n3078_lo, n3081_lo, n3084_lo, n3087_lo, n3090_lo,
    n3093_lo, n3096_lo, n3099_lo, n3102_lo, n3105_lo, n3108_lo, n3111_lo,
    n3114_lo, n3117_lo, n3120_lo, n3123_lo, n3126_lo, n3129_lo, n3132_lo,
    n3135_lo, n3138_lo, n3141_lo, n3144_lo, n3147_lo, n3150_lo, n3153_lo,
    n3156_lo, n3159_lo, n3162_lo, n3165_lo, n3168_lo, n3171_lo, n3174_lo,
    n3177_lo, n3180_lo, n3183_lo, n3186_lo, n3189_lo, n3192_lo, n3195_lo,
    n3198_lo, n3201_lo, n3204_lo, n3207_lo, n3210_lo, n3213_lo, n3216_lo,
    n3219_lo, n3222_lo, n3225_lo, n3228_lo, n3231_lo, n3234_lo, n3237_lo,
    n3240_lo, n3243_lo, n3246_lo, n3249_lo, n3252_lo, n3255_lo, n3258_lo,
    n3261_lo, n3264_lo, n3267_lo, n3270_lo, n3273_lo, n3276_lo, n3279_lo,
    n3282_lo, n3285_lo, n3288_lo, n3291_lo, n3294_lo, n3297_lo, n3300_lo,
    n3303_lo, n3306_lo, n3309_lo, n3312_lo, n3315_lo, n3318_lo, n3321_lo,
    n3324_lo, n3327_lo, n3330_lo, n3333_lo, n3336_lo, n3339_lo, n3342_lo,
    n3345_lo, n3348_lo, n3351_lo, n3354_lo, n3357_lo, n3360_lo, n3363_lo,
    n3366_lo, n3369_lo, n3372_lo, n3375_lo, n3378_lo, n3381_lo, n3384_lo,
    n3387_lo, n3390_lo, n3393_lo, n3396_lo, n3399_lo, n3402_lo, n3405_lo,
    n3408_lo, n3411_lo, n3414_lo, n3417_lo, n3420_lo, n3423_lo, n3426_lo,
    n3429_lo, n3432_lo, n3435_lo, n3438_lo, n3441_lo, n3444_lo, n3447_lo,
    n3450_lo, n3453_lo, n3456_lo, n3459_lo, n3462_lo, n3465_lo, n3468_lo,
    n3471_lo, n3474_lo, n3477_lo, n3480_lo, n3483_lo, n3486_lo, n3489_lo,
    n3492_lo, n3495_lo, n3498_lo, n3501_lo, n3504_lo, n3507_lo, n3510_lo,
    n3513_lo, n3516_lo, n3519_lo, n3522_lo, n3525_lo, n3528_lo, n3531_lo,
    n3534_lo, n3537_lo, n3540_lo, n3543_lo, n3546_lo, n3549_lo, n3552_lo,
    n3555_lo, n3558_lo, n3561_lo, n3564_lo, n3567_lo, n3570_lo, n3573_lo,
    n3576_lo, n3579_lo, n3582_lo, n3585_lo, n3588_lo, n3591_lo, n3594_lo,
    n3597_lo, n3600_lo, n3603_lo, n3606_lo, n3609_lo, n3612_lo, n3615_lo,
    n3618_lo, n3621_lo, n3624_lo, n3627_lo, n3630_lo, n3633_lo, n3636_lo,
    n3639_lo, n3642_lo, n3645_lo, n3648_lo, n3651_lo, n3654_lo, n3657_lo,
    n3666_lo, n3669_lo, n3678_lo, n3687_lo, n3690_lo, n3702_lo, n3711_lo,
    n3714_lo, n3726_lo, n3735_lo, n3738_lo, n3750_lo, n3753_lo, n3759_lo,
    n3762_lo, n3765_lo, n3774_lo, n3777_lo, n3786_lo, n3789_lo, n3792_lo,
    n3795_lo, n3798_lo, n3801_lo, n3810_lo, n3813_lo, n3822_lo, n3825_lo,
    n3834_lo, n3843_lo, n3846_lo, n3867_lo, n3891_lo, n3915_lo, n3930_lo,
    n3933_lo, n3936_lo, n3942_lo, n3945_lo, n3948_lo, n3954_lo, n3957_lo,
    n3963_lo, n3966_lo, n3969_lo, n3975_lo, n3978_lo, n3987_lo, n3990_lo,
    n4002_lo, n4011_lo, n4014_lo, n4026_lo, n4035_lo, n4038_lo, n4050_lo,
    n4053_lo, n4059_lo, n4062_lo, n4065_lo, n4098_lo, n4107_lo, n4119_lo,
    n4131_lo, n4143_lo, n4155_lo, n4167_lo, n4179_lo, n4182_lo, n4185_lo,
    n4188_lo, n4194_lo, n4197_lo, n4200_lo, n4206_lo, n4209_lo, n4212_lo,
    n4215_lo, n4227_lo, n4230_lo, n4233_lo, n4236_lo, n4239_lo, n4242_lo,
    n4251_lo, n4263_lo, n4275_lo, n4278_lo, n4287_lo, n4290_lo, n4293_lo,
    n4299_lo, n4302_lo, n4305_lo, n4311_lo, n4314_lo, n4323_lo, n4326_lo,
    n4335_lo, n4338_lo, n4347_lo, n4350_lo, n4359_lo, n4362_lo, n4365_lo,
    n4371_lo, n4374_lo, n4383_lo, n4395_lo, n4407_lo, n4410_lo, n4413_lo,
    n4416_lo, n4419_lo, n4422_lo, n4425_lo, n4428_lo, n4431_lo, n4434_lo,
    n4437_lo, n4440_lo, n4443_lo, n4446_lo, n4449_lo, n4452_lo, n4455_lo,
    n4458_lo, n4461_lo, n4464_lo, n4467_lo, n4470_lo, n4473_lo, n4476_lo,
    n4479_lo, n4482_lo, n4485_lo, n4488_lo, n4494_lo, n4497_lo, n4500_lo,
    n4503_lo, n4506_lo, n4509_lo, n4512_lo, n4515_lo, n4518_lo, n4521_lo,
    n4524_lo, n4527_lo, n4530_lo, n4533_lo, n4536_lo, n4539_lo, n4542_lo,
    n4545_lo, n4548_lo, n4554_lo, n4557_lo, n4560_lo, n4563_lo, n4566_lo,
    n4569_lo, n4572_lo, n4575_lo, n4578_lo, n4581_lo, n4584_lo, n4587_lo,
    n4590_lo, n4593_lo, n4596_lo, n4599_lo, n4602_lo, n4605_lo, n4608_lo,
    n4611_lo, n4614_lo, n4617_lo, n4620_lo, n4623_lo, n4626_lo, n4629_lo,
    n4632_lo, n4635_lo, n4638_lo, n4641_lo, n4644_lo, n4647_lo, n4650_lo,
    n4653_lo, n4656_lo, n4659_lo, n4662_lo, n4665_lo, n4668_lo, n4671_lo,
    n4674_lo, n4677_lo, n4680_lo, n4683_lo, n4686_lo, n4689_lo, n4692_lo,
    n4695_lo, n4698_lo, n4701_lo, n4704_lo, n4707_lo, n4710_lo, n4713_lo,
    n4716_lo, n4719_lo, n4722_lo, n4725_lo, n4728_lo, n4731_lo, n4734_lo,
    n4737_lo, n4740_lo, n4743_lo, n6382_o2, n6383_o2, n6419_o2, n6420_o2,
    n6435_o2, n6436_o2, n6448_o2, n6449_o2, n6613_o2, n6614_o2, n6641_o2,
    n6658_o2, n6757_o2, n6756_o2, n7116_o2, n7156_o2, n6549_o2, n6550_o2,
    n7357_o2, n7358_o2, n7359_o2, n7360_o2, n6621_o2, n6623_o2, n6625_o2,
    n6626_o2, n6627_o2, n6628_o2, n6629_o2, n6630_o2, n6669_o2, n7449_o2,
    n7450_o2, n7451_o2, n7452_o2, n6682_o2, n6683_o2, n6684_o2, n6685_o2,
    n7463_o2, n6686_o2, n6687_o2, n6688_o2, n6689_o2, n6772_o2, n6773_o2,
    n6774_o2, n6775_o2, G3467_o2, G2810_o2, n6833_o2, n6945_o2, n6947_o2,
    n6949_o2, n6951_o2, n6888_o2, n6889_o2, n6936_o2, n6954_o2, n6955_o2,
    n6956_o2, n6957_o2, n6958_o2, n6982_o2, n6984_o2, n6974_o2, n6975_o2,
    n6999_o2, n7015_o2, n7016_o2, n7017_o2, n7018_o2, n7005_o2, n7019_o2,
    n7022_o2, n7023_o2, n7132_o2, n7133_o2, n7135_o2, n7136_o2, n7175_o2,
    n7155_o2, G3060_o2, n7383_o2, G3802_o2, G3859_o2, n7355_o2, n7356_o2,
    G4054_o2, G4068_o2, n7384_o2, n7387_o2, n7388_o2, n7389_o2, n7386_o2,
    n7453_o2, n7431_o2, n7432_o2, n7433_o2, n7430_o2, n7485_o2, n7486_o2,
    G2508_o2, G2486_o2, n2326_inv, n2329_inv, n3756_lo_buf_o2,
    n4056_lo_buf_o2, G3474_o2, n2341_inv, n7396_o2, n7398_o2, n7400_o2,
    n7401_o2, n7402_o2, n7403_o2, n7404_o2, n7405_o2, G2711_o2, n2371_inv,
    n7490_o2, n7527_o2, n7528_o2, n7529_o2, n7530_o2, n7523_o2, n7524_o2,
    n7525_o2, n7526_o2, n4296_lo_buf_o2, n4368_lo_buf_o2, G2466_o2,
    G2404_o2, n7534_o2, n7535_o2, n7536_o2, n7533_o2, G1060_o2, G963_o2,
    G2448_o2, G2685_o2, G2679_o2, G2774_o2, G2780_o2, G2759_o2, G2737_o2,
    G2850_o2, G3393_o2, G3404_o2, G3559_o2, G2744_o2, n3708_lo_buf_o2,
    n3840_lo_buf_o2, n4008_lo_buf_o2, n4104_lo_buf_o2, G1821_o2, G1734_o2,
    G3517_o2, G3533_o2, G3629_o2, G3645_o2, n2497_inv, G2731_o2, G2844_o2,
    n3732_lo_buf_o2, n4032_lo_buf_o2, G3552_o2, G2271_o2, n4248_lo_buf_o2,
    n4332_lo_buf_o2, n4344_lo_buf_o2, n4380_lo_buf_o2, G2398_o2, G2480_o2,
    G2418_o2, G1455_o2, G1449_o2, G1452_o2, G1425_o2, G1428_o2, G1419_o2,
    G1422_o2, n4308_lo_buf_o2, G2675_o2, G3035_o2, G3026_o2, G3029_o2,
    G3032_o2, G2999_o2, G3002_o2, G2770_o2, G3008_o2, G2073_o2, G2752_o2,
    G3005_o2, G5108_o2, G5135_o2, G5111_o2, G5138_o2, G3415_o2, G3386_o2,
    G3570_o2, G2430_o2, G3495_o2, G3621_o2, n4284_lo_buf_o2,
    n4356_lo_buf_o2, G2472_o2, G2410_o2, n3960_lo_buf_o2, n3972_lo_buf_o2,
    n2647_inv, n2650_inv, n3684_lo_buf_o2, n4080_lo_buf_o2,
    n4092_lo_buf_o2, n2662_inv, n2665_inv, G1147_o2, G2705_o2, G2693_o2,
    G2696_o2, G2700_o2, G2915_o2, G2966_o2, G2540_o2, G2788_o2, G2792_o2,
    G2797_o2, G2804_o2, G1038_o2, G1044_o2, G1090_o2, G1096_o2, G1029_o2,
    G3942_o2, G3954_o2, G4011_o2, G4017_o2, G1141_o2, G1081_o2, G2146_o2,
    G2145_o2, G2144_o2, G2143_o2, G2142_o2, G2141_o2, G2140_o2, G2139_o2,
    G3769_o2, G3773_o2, G3768_o2, G4101_o2, G3161_o2, G4143_o2, G3828_o2,
    G3831_o2, G3334_o2, G3335_o2, G3180_o2, G3340_o2, G3339_o2, G3341_o2,
    G3234_o2, G3829_o2, G3338_o2, G3336_o2, G3770_o2, G3918_o2, G3774_o2,
    G3921_o2, G3832_o2, G3993_o2, G2076_o2, G2071_o2, G2072_o2, G2069_o2,
    G2070_o2, G2067_o2, G2068_o2, G4095_o2, G3272_o2, G3269_o2, G3270_o2,
    G3271_o2, G3265_o2, G3266_o2, G4137_o2, G3268_o2, G2361_o2, G3228_o2,
    G3267_o2, G2336_o2, G3459_o2, G3428_o2, G3438_o2, G3449_o2, G3421_o2,
    G3576_o2, G3303_o2, G3583_o2, G3594_o2, G3674_o2, G3685_o2, G4504_o2,
    G4180_o2, G5123_o2, G5142_o2, G5126_o2, G5144_o2, G3912_o2, G4417_o2,
    G4420_o2, G3969_o2, G4023_o2, G2720_o2, G2837_o2, n2965_inv, n2968_inv,
    n2971_inv, n2974_inv, G1876_o2, G4996_o2, G4984_o2, G4920_o2, G4923_o2,
    G4930_o2, G4933_o2, n4320_lo_buf_o2, G2424_o2, G3317_o2, G3503_o2,
    G3485_o2, G3611_o2, n3864_lo_buf_o2, n3888_lo_buf_o2, n4116_lo_buf_o2,
    n4128_lo_buf_o2, n4140_lo_buf_o2, n4152_lo_buf_o2, G1815_o2, G1728_o2,
    G1035_o2, G1041_o2, G1087_o2, G1093_o2, G1132_o2, G1108_o2, G1138_o2,
    G1114_o2, G1807_o2, G2108_o2, G1126_o2, G1899_o2, G2134_o2, G1852_o2,
    G2116_o2, G2543_o2, G2727_o2, G2715_o2, G2832_o2, G1873_o2, G3291_o2,
    G5025_o2, G5036_o2, G3132_o2, G5038_o2, G5039_o2, n3118_inv, n3121_inv,
    n3124_inv, n3127_inv, n3984_lo_buf_o2, G1802_o2, G1804_o2, G1849_o2,
    G1851_o2, G2492_o2, G1799_o2, G4231_o2, G4234_o2, G4245_o2, G4247_o2,
    G1894_o2, G1846_o2, G4238_o2, G4249_o2, G2293_o2, G5022_o2, G5006_o2,
    G4944_o2, G4946_o2, G4954_o2, G4956_o2, G3546_o2, G3658_o2, G1344_o2,
    G2921_o2, n3912_lo_buf_o2, G1835_o2, G3810_o2, G3866_o2, G3811_o2,
    G2269_o2, G3812_o2, G3867_o2, G3868_o2, G3809_o2, G3716_o2, G4529_o2,
    G4670_o2, G4493_o2, G4580_o2, G3822_o2, G3877_o2, G4131_o2, G4170_o2,
    G4051_o2, G4065_o2, G4697_o2, G4706_o2, G2460_o2, G2454_o2, G2392_o2,
    G2386_o2, n4260_lo_buf_o2, n4272_lo_buf_o2, n4392_lo_buf_o2,
    n4404_lo_buf_o2, G1512_o2, G3135_o2, G2379_o2, n4164_lo_buf_o2,
    n4176_lo_buf_o2, n4224_lo_buf_o2, G2975_o2, G2978_o2, G2933_o2,
    G2936_o2, G1356_o2, G1359_o2, G1398_o2, G1401_o2;
  wire new_new_n2328__, new_new_n2330__, new_new_n2332__, new_new_n2334__,
    new_new_n2336__, new_new_n2338__, new_new_n2340__, new_new_n2342__,
    new_new_n2344__, new_new_n2346__, new_new_n2348__, new_new_n2350__,
    new_new_n2352__, new_new_n2354__, new_new_n2356__, new_new_n2358__,
    new_new_n2360__, new_new_n2362__, new_new_n2364__, new_new_n2366__,
    new_new_n2368__, new_new_n2370__, new_new_n2372__, new_new_n2374__,
    new_new_n2376__, new_new_n2378__, new_new_n2380__, new_new_n2382__,
    new_new_n2384__, new_new_n2386__, new_new_n2388__, new_new_n2390__,
    new_new_n2392__, new_new_n2394__, new_new_n2396__, new_new_n2398__,
    new_new_n2400__, new_new_n2402__, new_new_n2404__, new_new_n2406__,
    new_new_n2408__, new_new_n2410__, new_new_n2412__, new_new_n2414__,
    new_new_n2416__, new_new_n2418__, new_new_n2420__, new_new_n2422__,
    new_new_n2424__, new_new_n2426__, new_new_n2428__, new_new_n2430__,
    new_new_n2432__, new_new_n2434__, new_new_n2436__, new_new_n2438__,
    new_new_n2440__, new_new_n2442__, new_new_n2444__, new_new_n2446__,
    new_new_n2448__, new_new_n2450__, new_new_n2452__, new_new_n2454__,
    new_new_n2456__, new_new_n2458__, new_new_n2460__, new_new_n2462__,
    new_new_n2464__, new_new_n2466__, new_new_n2468__, new_new_n2470__,
    new_new_n2472__, new_new_n2474__, new_new_n2476__, new_new_n2478__,
    new_new_n2480__, new_new_n2482__, new_new_n2484__, new_new_n2486__,
    new_new_n2488__, new_new_n2490__, new_new_n2492__, new_new_n2494__,
    new_new_n2496__, new_new_n2498__, new_new_n2500__, new_new_n2502__,
    new_new_n2504__, new_new_n2506__, new_new_n2508__, new_new_n2510__,
    new_new_n2512__, new_new_n2514__, new_new_n2516__, new_new_n2518__,
    new_new_n2520__, new_new_n2522__, new_new_n2524__, new_new_n2526__,
    new_new_n2528__, new_new_n2530__, new_new_n2532__, new_new_n2534__,
    new_new_n2536__, new_new_n2538__, new_new_n2540__, new_new_n2542__,
    new_new_n2544__, new_new_n2546__, new_new_n2548__, new_new_n2550__,
    new_new_n2552__, new_new_n2554__, new_new_n2556__, new_new_n2558__,
    new_new_n2560__, new_new_n2562__, new_new_n2564__, new_new_n2566__,
    new_new_n2568__, new_new_n2570__, new_new_n2572__, new_new_n2573__,
    new_new_n2574__, new_new_n2575__, new_new_n2576__, new_new_n2578__,
    new_new_n2580__, new_new_n2582__, new_new_n2584__, new_new_n2586__,
    new_new_n2588__, new_new_n2590__, new_new_n2592__, new_new_n2594__,
    new_new_n2596__, new_new_n2598__, new_new_n2600__, new_new_n2602__,
    new_new_n2604__, new_new_n2606__, new_new_n2608__, new_new_n2610__,
    new_new_n2612__, new_new_n2614__, new_new_n2616__, new_new_n2618__,
    new_new_n2620__, new_new_n2622__, new_new_n2624__, new_new_n2626__,
    new_new_n2628__, new_new_n2630__, new_new_n2632__, new_new_n2634__,
    new_new_n2636__, new_new_n2638__, new_new_n2640__, new_new_n2642__,
    new_new_n2644__, new_new_n2646__, new_new_n2648__, new_new_n2650__,
    new_new_n2652__, new_new_n2654__, new_new_n2656__, new_new_n2658__,
    new_new_n2660__, new_new_n2662__, new_new_n2664__, new_new_n2666__,
    new_new_n2668__, new_new_n2670__, new_new_n2672__, new_new_n2674__,
    new_new_n2676__, new_new_n2678__, new_new_n2680__, new_new_n2682__,
    new_new_n2684__, new_new_n2686__, new_new_n2688__, new_new_n2690__,
    new_new_n2691__, new_new_n2692__, new_new_n2694__, new_new_n2696__,
    new_new_n2698__, new_new_n2699__, new_new_n2700__, new_new_n2702__,
    new_new_n2704__, new_new_n2706__, new_new_n2708__, new_new_n2710__,
    new_new_n2712__, new_new_n2714__, new_new_n2716__, new_new_n2718__,
    new_new_n2720__, new_new_n2722__, new_new_n2724__, new_new_n2726__,
    new_new_n2728__, new_new_n2730__, new_new_n2732__, new_new_n2734__,
    new_new_n2736__, new_new_n2739__, new_new_n2740__, new_new_n2742__,
    new_new_n2744__, new_new_n2747__, new_new_n2748__, new_new_n2750__,
    new_new_n2752__, new_new_n2755__, new_new_n2756__, new_new_n2758__,
    new_new_n2760__, new_new_n2763__, new_new_n2764__, new_new_n2766__,
    new_new_n2768__, new_new_n2770__, new_new_n2771__, new_new_n2772__,
    new_new_n2774__, new_new_n2776__, new_new_n2778__, new_new_n2779__,
    new_new_n2780__, new_new_n2782__, new_new_n2784__, new_new_n2787__,
    new_new_n2788__, new_new_n2790__, new_new_n2792__, new_new_n2794__,
    new_new_n2796__, new_new_n2798__, new_new_n2800__, new_new_n2802__,
    new_new_n2804__, new_new_n2806__, new_new_n2808__, new_new_n2810__,
    new_new_n2812__, new_new_n2814__, new_new_n2816__, new_new_n2818__,
    new_new_n2820__, new_new_n2822__, new_new_n2824__, new_new_n2826__,
    new_new_n2828__, new_new_n2830__, new_new_n2832__, new_new_n2834__,
    new_new_n2836__, new_new_n2838__, new_new_n2840__, new_new_n2842__,
    new_new_n2844__, new_new_n2846__, new_new_n2848__, new_new_n2850__,
    new_new_n2851__, new_new_n2852__, new_new_n2854__, new_new_n2856__,
    new_new_n2858__, new_new_n2860__, new_new_n2862__, new_new_n2864__,
    new_new_n2866__, new_new_n2868__, new_new_n2870__, new_new_n2872__,
    new_new_n2874__, new_new_n2876__, new_new_n2878__, new_new_n2880__,
    new_new_n2882__, new_new_n2884__, new_new_n2886__, new_new_n2888__,
    new_new_n2890__, new_new_n2892__, new_new_n2894__, new_new_n2896__,
    new_new_n2898__, new_new_n2900__, new_new_n2902__, new_new_n2904__,
    new_new_n2907__, new_new_n2908__, new_new_n2910__, new_new_n2912__,
    new_new_n2915__, new_new_n2916__, new_new_n2918__, new_new_n2920__,
    new_new_n2923__, new_new_n2924__, new_new_n2926__, new_new_n2928__,
    new_new_n2931__, new_new_n2932__, new_new_n2934__, new_new_n2936__,
    new_new_n2939__, new_new_n2940__, new_new_n2942__, new_new_n2944__,
    new_new_n2947__, new_new_n2948__, new_new_n2950__, new_new_n2952__,
    new_new_n2955__, new_new_n2956__, new_new_n2958__, new_new_n2960__,
    new_new_n2963__, new_new_n2964__, new_new_n2966__, new_new_n2968__,
    new_new_n2970__, new_new_n2972__, new_new_n2974__, new_new_n2976__,
    new_new_n2978__, new_new_n2980__, new_new_n2982__, new_new_n2984__,
    new_new_n2986__, new_new_n2988__, new_new_n2990__, new_new_n2992__,
    new_new_n2994__, new_new_n2996__, new_new_n2998__, new_new_n3000__,
    new_new_n3002__, new_new_n3004__, new_new_n3006__, new_new_n3008__,
    new_new_n3010__, new_new_n3012__, new_new_n3014__, new_new_n3016__,
    new_new_n3018__, new_new_n3020__, new_new_n3022__, new_new_n3024__,
    new_new_n3026__, new_new_n3028__, new_new_n3030__, new_new_n3032__,
    new_new_n3034__, new_new_n3036__, new_new_n3038__, new_new_n3040__,
    new_new_n3042__, new_new_n3044__, new_new_n3046__, new_new_n3048__,
    new_new_n3050__, new_new_n3052__, new_new_n3054__, new_new_n3056__,
    new_new_n3058__, new_new_n3060__, new_new_n3062__, new_new_n3064__,
    new_new_n3066__, new_new_n3068__, new_new_n3070__, new_new_n3072__,
    new_new_n3075__, new_new_n3076__, new_new_n3078__, new_new_n3080__,
    new_new_n3082__, new_new_n3084__, new_new_n3086__, new_new_n3088__,
    new_new_n3091__, new_new_n3092__, new_new_n3094__, new_new_n3096__,
    new_new_n3098__, new_new_n3100__, new_new_n3102__, new_new_n3104__,
    new_new_n3106__, new_new_n3108__, new_new_n3110__, new_new_n3112__,
    new_new_n3114__, new_new_n3116__, new_new_n3118__, new_new_n3120__,
    new_new_n3122__, new_new_n3124__, new_new_n3126__, new_new_n3128__,
    new_new_n3130__, new_new_n3132__, new_new_n3134__, new_new_n3136__,
    new_new_n3138__, new_new_n3140__, new_new_n3142__, new_new_n3144__,
    new_new_n3146__, new_new_n3148__, new_new_n3150__, new_new_n3152__,
    new_new_n3154__, new_new_n3156__, new_new_n3158__, new_new_n3160__,
    new_new_n3162__, new_new_n3164__, new_new_n3166__, new_new_n3168__,
    new_new_n3170__, new_new_n3171__, new_new_n3172__, new_new_n3174__,
    new_new_n3176__, new_new_n3179__, new_new_n3180__, new_new_n3182__,
    new_new_n3184__, new_new_n3186__, new_new_n3188__, new_new_n3190__,
    new_new_n3192__, new_new_n3194__, new_new_n3196__, new_new_n3198__,
    new_new_n3200__, new_new_n3203__, new_new_n3204__, new_new_n3206__,
    new_new_n3208__, new_new_n3210__, new_new_n3211__, new_new_n3212__,
    new_new_n3214__, new_new_n3216__, new_new_n3218__, new_new_n3220__,
    new_new_n3222__, new_new_n3224__, new_new_n3226__, new_new_n3228__,
    new_new_n3230__, new_new_n3232__, new_new_n3234__, new_new_n3236__,
    new_new_n3238__, new_new_n3240__, new_new_n3242__, new_new_n3244__,
    new_new_n3246__, new_new_n3248__, new_new_n3250__, new_new_n3252__,
    new_new_n3254__, new_new_n3256__, new_new_n3258__, new_new_n3260__,
    new_new_n3262__, new_new_n3264__, new_new_n3266__, new_new_n3268__,
    new_new_n3270__, new_new_n3272__, new_new_n3274__, new_new_n3276__,
    new_new_n3278__, new_new_n3280__, new_new_n3282__, new_new_n3284__,
    new_new_n3286__, new_new_n3288__, new_new_n3290__, new_new_n3292__,
    new_new_n3294__, new_new_n3296__, new_new_n3298__, new_new_n3300__,
    new_new_n3302__, new_new_n3304__, new_new_n3306__, new_new_n3308__,
    new_new_n3310__, new_new_n3312__, new_new_n3314__, new_new_n3316__,
    new_new_n3318__, new_new_n3320__, new_new_n3322__, new_new_n3324__,
    new_new_n3326__, new_new_n3328__, new_new_n3330__, new_new_n3332__,
    new_new_n3334__, new_new_n3336__, new_new_n3338__, new_new_n3340__,
    new_new_n3342__, new_new_n3344__, new_new_n3346__, new_new_n3348__,
    new_new_n3350__, new_new_n3352__, new_new_n3354__, new_new_n3356__,
    new_new_n3358__, new_new_n3360__, new_new_n3362__, new_new_n3364__,
    new_new_n3366__, new_new_n3368__, new_new_n3370__, new_new_n3372__,
    new_new_n3374__, new_new_n3376__, new_new_n3378__, new_new_n3380__,
    new_new_n3382__, new_new_n3384__, new_new_n3386__, new_new_n3388__,
    new_new_n3390__, new_new_n3391__, new_new_n3392__, new_new_n3394__,
    new_new_n3395__, new_new_n3396__, new_new_n3397__, new_new_n3398__,
    new_new_n3399__, new_new_n3400__, new_new_n3401__, new_new_n3402__,
    new_new_n3403__, new_new_n3404__, new_new_n3405__, new_new_n3406__,
    new_new_n3408__, new_new_n3409__, new_new_n3410__, new_new_n3411__,
    new_new_n3412__, new_new_n3414__, new_new_n3415__, new_new_n3416__,
    new_new_n3418__, new_new_n3420__, new_new_n3422__, new_new_n3424__,
    new_new_n3427__, new_new_n3428__, new_new_n3430__, new_new_n3431__,
    new_new_n3432__, new_new_n3434__, new_new_n3435__, new_new_n3436__,
    new_new_n3438__, new_new_n3440__, new_new_n3441__, new_new_n3442__,
    new_new_n3443__, new_new_n3444__, new_new_n3445__, new_new_n3446__,
    new_new_n3447__, new_new_n3448__, new_new_n3449__, new_new_n3450__,
    new_new_n3451__, new_new_n3452__, new_new_n3454__, new_new_n3456__,
    new_new_n3457__, new_new_n3458__, new_new_n3460__, new_new_n3462__,
    new_new_n3463__, new_new_n3464__, new_new_n3466__, new_new_n3468__,
    new_new_n3469__, new_new_n3470__, new_new_n3472__, new_new_n3474__,
    new_new_n3475__, new_new_n3476__, new_new_n3478__, new_new_n3479__,
    new_new_n3480__, new_new_n3482__, new_new_n3483__, new_new_n3484__,
    new_new_n3485__, new_new_n3486__, new_new_n3487__, new_new_n3488__,
    new_new_n3489__, new_new_n3490__, new_new_n3491__, new_new_n3492__,
    new_new_n3493__, new_new_n3494__, new_new_n3496__, new_new_n3497__,
    new_new_n3498__, new_new_n3499__, new_new_n3500__, new_new_n3502__,
    new_new_n3503__, new_new_n3504__, new_new_n3505__, new_new_n3507__,
    new_new_n3508__, new_new_n3509__, new_new_n3511__, new_new_n3512__,
    new_new_n3513__, new_new_n3515__, new_new_n3516__, new_new_n3517__,
    new_new_n3519__, new_new_n3520__, new_new_n3522__, new_new_n3524__,
    new_new_n3525__, new_new_n3526__, new_new_n3528__, new_new_n3530__,
    new_new_n3532__, new_new_n3534__, new_new_n3536__, new_new_n3538__,
    new_new_n3540__, new_new_n3541__, new_new_n3542__, new_new_n3544__,
    new_new_n3546__, new_new_n3549__, new_new_n3550__, new_new_n3551__,
    new_new_n3552__, new_new_n3553__, new_new_n3554__, new_new_n3555__,
    new_new_n3556__, new_new_n3557__, new_new_n3558__, new_new_n3559__,
    new_new_n3560__, new_new_n3561__, new_new_n3562__, new_new_n3564__,
    new_new_n3565__, new_new_n3566__, new_new_n3567__, new_new_n3568__,
    new_new_n3570__, new_new_n3571__, new_new_n3572__, new_new_n3573__,
    new_new_n3574__, new_new_n3576__, new_new_n3577__, new_new_n3578__,
    new_new_n3579__, new_new_n3580__, new_new_n3581__, new_new_n3582__,
    new_new_n3583__, new_new_n3584__, new_new_n3585__, new_new_n3586__,
    new_new_n3587__, new_new_n3588__, new_new_n3589__, new_new_n3590__,
    new_new_n3592__, new_new_n3593__, new_new_n3594__, new_new_n3595__,
    new_new_n3596__, new_new_n3597__, new_new_n3598__, new_new_n3599__,
    new_new_n3600__, new_new_n3601__, new_new_n3602__, new_new_n3603__,
    new_new_n3604__, new_new_n3606__, new_new_n3608__, new_new_n3611__,
    new_new_n3612__, new_new_n3614__, new_new_n3616__, new_new_n3618__,
    new_new_n3619__, new_new_n3620__, new_new_n3622__, new_new_n3624__,
    new_new_n3626__, new_new_n3627__, new_new_n3628__, new_new_n3630__,
    new_new_n3632__, new_new_n3635__, new_new_n3636__, new_new_n3638__,
    new_new_n3640__, new_new_n3643__, new_new_n3644__, new_new_n3646__,
    new_new_n3648__, new_new_n3650__, new_new_n3651__, new_new_n3652__,
    new_new_n3654__, new_new_n3656__, new_new_n3657__, new_new_n3658__,
    new_new_n3660__, new_new_n3662__, new_new_n3664__, new_new_n3665__,
    new_new_n3666__, new_new_n3668__, new_new_n3670__, new_new_n3672__,
    new_new_n3673__, new_new_n3674__, new_new_n3676__, new_new_n3678__,
    new_new_n3680__, new_new_n3681__, new_new_n3682__, new_new_n3684__,
    new_new_n3686__, new_new_n3688__, new_new_n3689__, new_new_n3690__,
    new_new_n3692__, new_new_n3694__, new_new_n3695__, new_new_n3696__,
    new_new_n3698__, new_new_n3700__, new_new_n3702__, new_new_n3703__,
    new_new_n3704__, new_new_n3706__, new_new_n3708__, new_new_n3710__,
    new_new_n3712__, new_new_n3714__, new_new_n3716__, new_new_n3719__,
    new_new_n3720__, new_new_n3722__, new_new_n3724__, new_new_n3727__,
    new_new_n3728__, new_new_n3730__, new_new_n3732__, new_new_n3735__,
    new_new_n3736__, new_new_n3738__, new_new_n3740__, new_new_n3742__,
    new_new_n3744__, new_new_n3746__, new_new_n3748__, new_new_n3750__,
    new_new_n3752__, new_new_n3754__, new_new_n3756__, new_new_n3758__,
    new_new_n3759__, new_new_n3760__, new_new_n3762__, new_new_n3764__,
    new_new_n3766__, new_new_n3767__, new_new_n3768__, new_new_n3770__,
    new_new_n3772__, new_new_n3774__, new_new_n3775__, new_new_n3776__,
    new_new_n3778__, new_new_n3780__, new_new_n3782__, new_new_n3783__,
    new_new_n3784__, new_new_n3786__, new_new_n3788__, new_new_n3790__,
    new_new_n3791__, new_new_n3792__, new_new_n3794__, new_new_n3796__,
    new_new_n3798__, new_new_n3799__, new_new_n3800__, new_new_n3802__,
    new_new_n3804__, new_new_n3806__, new_new_n3807__, new_new_n3808__,
    new_new_n3810__, new_new_n3812__, new_new_n3814__, new_new_n3815__,
    new_new_n3816__, new_new_n3818__, new_new_n3820__, new_new_n3823__,
    new_new_n3825__, new_new_n3827__, new_new_n3829__, new_new_n3831__,
    new_new_n3833__, new_new_n3835__, new_new_n3837__, new_new_n3839__,
    new_new_n3841__, new_new_n3842__, new_new_n3845__, new_new_n3846__,
    new_new_n3848__, new_new_n3849__, new_new_n3850__, new_new_n3851__,
    new_new_n3853__, new_new_n3854__, new_new_n3855__, new_new_n3857__,
    new_new_n3858__, new_new_n3859__, new_new_n3860__, new_new_n3862__,
    new_new_n3864__, new_new_n3866__, new_new_n3868__, new_new_n3869__,
    new_new_n3870__, new_new_n3871__, new_new_n3872__, new_new_n3873__,
    new_new_n3874__, new_new_n3876__, new_new_n3877__, new_new_n3878__,
    new_new_n3880__, new_new_n3882__, new_new_n3883__, new_new_n3884__,
    new_new_n3885__, new_new_n3886__, new_new_n3887__, new_new_n3889__,
    new_new_n3891__, new_new_n3892__, new_new_n3893__, new_new_n3894__,
    new_new_n3895__, new_new_n3896__, new_new_n3897__, new_new_n3898__,
    new_new_n3899__, new_new_n3900__, new_new_n3901__, new_new_n3902__,
    new_new_n3903__, new_new_n3904__, new_new_n3905__, new_new_n3906__,
    new_new_n3907__, new_new_n3908__, new_new_n3909__, new_new_n3910__,
    new_new_n3911__, new_new_n3912__, new_new_n3913__, new_new_n3914__,
    new_new_n3916__, new_new_n3917__, new_new_n3918__, new_new_n3919__,
    new_new_n3921__, new_new_n3922__, new_new_n3924__, new_new_n3926__,
    new_new_n3927__, new_new_n3928__, new_new_n3929__, new_new_n3930__,
    new_new_n3931__, new_new_n3932__, new_new_n3934__, new_new_n3935__,
    new_new_n3936__, new_new_n3937__, new_new_n3938__, new_new_n3939__,
    new_new_n3940__, new_new_n3941__, new_new_n3942__, new_new_n3943__,
    new_new_n3944__, new_new_n3945__, new_new_n3946__, new_new_n3947__,
    new_new_n3948__, new_new_n3949__, new_new_n3950__, new_new_n3951__,
    new_new_n3952__, new_new_n3953__, new_new_n3954__, new_new_n3955__,
    new_new_n3956__, new_new_n3957__, new_new_n3958__, new_new_n3959__,
    new_new_n3960__, new_new_n3961__, new_new_n3962__, new_new_n3963__,
    new_new_n3964__, new_new_n3965__, new_new_n3966__, new_new_n3967__,
    new_new_n3968__, new_new_n3969__, new_new_n3970__, new_new_n3971__,
    new_new_n3972__, new_new_n3973__, new_new_n3974__, new_new_n3975__,
    new_new_n3976__, new_new_n3977__, new_new_n3978__, new_new_n3979__,
    new_new_n3980__, new_new_n3981__, new_new_n3982__, new_new_n3983__,
    new_new_n3984__, new_new_n3985__, new_new_n3986__, new_new_n3987__,
    new_new_n3989__, new_new_n3990__, new_new_n3991__, new_new_n3993__,
    new_new_n3995__, new_new_n3996__, new_new_n3998__, new_new_n4001__,
    new_new_n4003__, new_new_n4004__, new_new_n4005__, new_new_n4006__,
    new_new_n4007__, new_new_n4008__, new_new_n4010__, new_new_n4012__,
    new_new_n4013__, new_new_n4014__, new_new_n4015__, new_new_n4016__,
    new_new_n4017__, new_new_n4018__, new_new_n4020__, new_new_n4022__,
    new_new_n4023__, new_new_n4024__, new_new_n4026__, new_new_n4028__,
    new_new_n4030__, new_new_n4031__, new_new_n4032__, new_new_n4034__,
    new_new_n4036__, new_new_n4037__, new_new_n4038__, new_new_n4040__,
    new_new_n4041__, new_new_n4042__, new_new_n4043__, new_new_n4044__,
    new_new_n4046__, new_new_n4048__, new_new_n4050__, new_new_n4052__,
    new_new_n4054__, new_new_n4056__, new_new_n4058__, new_new_n4060__,
    new_new_n4062__, new_new_n4064__, new_new_n4066__, new_new_n4068__,
    new_new_n4070__, new_new_n4072__, new_new_n4074__, new_new_n4076__,
    new_new_n4078__, new_new_n4080__, new_new_n4082__, new_new_n4083__,
    new_new_n4084__, new_new_n4085__, new_new_n4086__, new_new_n4087__,
    new_new_n4088__, new_new_n4089__, new_new_n4090__, new_new_n4092__,
    new_new_n4094__, new_new_n4096__, new_new_n4098__, new_new_n4099__,
    new_new_n4100__, new_new_n4101__, new_new_n4102__, new_new_n4104__,
    new_new_n4105__, new_new_n4106__, new_new_n4107__, new_new_n4108__,
    new_new_n4109__, new_new_n4110__, new_new_n4111__, new_new_n4112__,
    new_new_n4113__, new_new_n4114__, new_new_n4116__, new_new_n4118__,
    new_new_n4119__, new_new_n4120__, new_new_n4121__, new_new_n4122__,
    new_new_n4123__, new_new_n4124__, new_new_n4126__, new_new_n4128__,
    new_new_n4129__, new_new_n4130__, new_new_n4132__, new_new_n4134__,
    new_new_n4135__, new_new_n4136__, new_new_n4137__, new_new_n4138__,
    new_new_n4140__, new_new_n4141__, new_new_n4142__, new_new_n4144__,
    new_new_n4145__, new_new_n4146__, new_new_n4148__, new_new_n4150__,
    new_new_n4152__, new_new_n4154__, new_new_n4156__, new_new_n4157__,
    new_new_n4158__, new_new_n4160__, new_new_n4162__, new_new_n4164__,
    new_new_n4166__, new_new_n4168__, new_new_n4170__, new_new_n4172__,
    new_new_n4174__, new_new_n4175__, new_new_n4176__, new_new_n4177__,
    new_new_n4178__, new_new_n4179__, new_new_n4180__, new_new_n4181__,
    new_new_n4182__, new_new_n4183__, new_new_n4184__, new_new_n4185__,
    new_new_n4186__, new_new_n4187__, new_new_n4188__, new_new_n4189__,
    new_new_n4190__, new_new_n4191__, new_new_n4192__, new_new_n4193__,
    new_new_n4194__, new_new_n4195__, new_new_n4196__, new_new_n4197__,
    new_new_n4198__, new_new_n4199__, new_new_n4200__, new_new_n4201__,
    new_new_n4202__, new_new_n4203__, new_new_n4204__, new_new_n4205__,
    new_new_n4206__, new_new_n4207__, new_new_n4208__, new_new_n4209__,
    new_new_n4210__, new_new_n4211__, new_new_n4212__, new_new_n4213__,
    new_new_n4214__, new_new_n4217__, new_new_n4219__, new_new_n4221__,
    new_new_n4222__, new_new_n4223__, new_new_n4224__, new_new_n4225__,
    new_new_n4226__, new_new_n4227__, new_new_n4228__, new_new_n4229__,
    new_new_n4230__, new_new_n4231__, new_new_n4232__, new_new_n4233__,
    new_new_n4234__, new_new_n4235__, new_new_n4236__, new_new_n4237__,
    new_new_n4238__, new_new_n4239__, new_new_n4240__, new_new_n4241__,
    new_new_n4242__, new_new_n4243__, new_new_n4244__, new_new_n4246__,
    new_new_n4247__, new_new_n4248__, new_new_n4250__, new_new_n4252__,
    new_new_n4253__, new_new_n4254__, new_new_n4255__, new_new_n4256__,
    new_new_n4257__, new_new_n4258__, new_new_n4259__, new_new_n4260__,
    new_new_n4261__, new_new_n4262__, new_new_n4263__, new_new_n4264__,
    new_new_n4265__, new_new_n4266__, new_new_n4267__, new_new_n4268__,
    new_new_n4269__, new_new_n4270__, new_new_n4271__, new_new_n4272__,
    new_new_n4273__, new_new_n4274__, new_new_n4275__, new_new_n4276__,
    new_new_n4277__, new_new_n4278__, new_new_n4279__, new_new_n4280__,
    new_new_n4281__, new_new_n4282__, new_new_n4283__, new_new_n4284__,
    new_new_n4285__, new_new_n4286__, new_new_n4287__, new_new_n4288__,
    new_new_n4289__, new_new_n4290__, new_new_n4291__, new_new_n4292__,
    new_new_n4293__, new_new_n4294__, new_new_n4295__, new_new_n4296__,
    new_new_n4297__, new_new_n4298__, new_new_n4299__, new_new_n4300__,
    new_new_n4301__, new_new_n4302__, new_new_n4303__, new_new_n4304__,
    new_new_n4305__, new_new_n4306__, new_new_n4307__, new_new_n4308__,
    new_new_n4309__, new_new_n4310__, new_new_n4311__, new_new_n4312__,
    new_new_n4313__, new_new_n4314__, new_new_n4315__, new_new_n4316__,
    new_new_n4317__, new_new_n4318__, new_new_n4319__, new_new_n4320__,
    new_new_n4321__, new_new_n4322__, new_new_n4323__, new_new_n4324__,
    new_new_n4325__, new_new_n4326__, new_new_n4327__, new_new_n4328__,
    new_new_n4329__, new_new_n4330__, new_new_n4331__, new_new_n4332__,
    new_new_n4333__, new_new_n4334__, new_new_n4335__, new_new_n4336__,
    new_new_n4337__, new_new_n4338__, new_new_n4339__, new_new_n4340__,
    new_new_n4341__, new_new_n4342__, new_new_n4343__, new_new_n4344__,
    new_new_n4345__, new_new_n4346__, new_new_n4347__, new_new_n4348__,
    new_new_n4349__, new_new_n4350__, new_new_n4351__, new_new_n4352__,
    new_new_n4353__, new_new_n4354__, new_new_n4355__, new_new_n4356__,
    new_new_n4357__, new_new_n4358__, new_new_n4359__, new_new_n4360__,
    new_new_n4361__, new_new_n4362__, new_new_n4363__, new_new_n4364__,
    new_new_n4365__, new_new_n4366__, new_new_n4367__, new_new_n4368__,
    new_new_n4369__, new_new_n4370__, new_new_n4371__, new_new_n4372__,
    new_new_n4373__, new_new_n4374__, new_new_n4375__, new_new_n4376__,
    new_new_n4377__, new_new_n4378__, new_new_n4379__, new_new_n4380__,
    new_new_n4381__, new_new_n4382__, new_new_n4383__, new_new_n4384__,
    new_new_n4385__, new_new_n4386__, new_new_n4387__, new_new_n4388__,
    new_new_n4389__, new_new_n4390__, new_new_n4391__, new_new_n4392__,
    new_new_n4393__, new_new_n4394__, new_new_n4395__, new_new_n4396__,
    new_new_n4397__, new_new_n4398__, new_new_n4399__, new_new_n4400__,
    new_new_n4401__, new_new_n4402__, new_new_n4403__, new_new_n4404__,
    new_new_n4405__, new_new_n4406__, new_new_n4407__, new_new_n4408__,
    new_new_n4409__, new_new_n4410__, new_new_n4411__, new_new_n4412__,
    new_new_n4413__, new_new_n4414__, new_new_n4415__, new_new_n4416__,
    new_new_n4417__, new_new_n4418__, new_new_n4419__, new_new_n4420__,
    new_new_n4421__, new_new_n4422__, new_new_n4423__, new_new_n4424__,
    new_new_n4425__, new_new_n4426__, new_new_n4427__, new_new_n4428__,
    new_new_n4429__, new_new_n4430__, new_new_n4431__, new_new_n4432__,
    new_new_n4433__, new_new_n4434__, new_new_n4435__, new_new_n4437__,
    new_new_n4438__, new_new_n4440__, new_new_n4442__, new_new_n4444__,
    new_new_n4445__, new_new_n4446__, new_new_n4447__, new_new_n4448__,
    new_new_n4449__, new_new_n4450__, new_new_n4451__, new_new_n4452__,
    new_new_n4453__, new_new_n4454__, new_new_n4455__, new_new_n4456__,
    new_new_n4457__, new_new_n4458__, new_new_n4459__, new_new_n4460__,
    new_new_n4461__, new_new_n4462__, new_new_n4463__, new_new_n4464__,
    new_new_n4465__, new_new_n4466__, new_new_n4467__, new_new_n4468__,
    new_new_n4469__, new_new_n4470__, new_new_n4471__, new_new_n4472__,
    new_new_n4473__, new_new_n4474__, new_new_n4475__, new_new_n4476__,
    new_new_n4477__, new_new_n4478__, new_new_n4479__, new_new_n4480__,
    new_new_n4481__, new_new_n4482__, new_new_n4483__, new_new_n4484__,
    new_new_n4486__, new_new_n4488__, new_new_n4489__, new_new_n4490__,
    new_new_n4491__, new_new_n4492__, new_new_n4494__, new_new_n4496__,
    new_new_n4498__, new_new_n4500__, new_new_n4502__, new_new_n4504__,
    new_new_n4505__, new_new_n4506__, new_new_n4507__, new_new_n4508__,
    new_new_n4509__, new_new_n4510__, new_new_n4511__, new_new_n4512__,
    new_new_n4513__, new_new_n4514__, new_new_n4515__, new_new_n4516__,
    new_new_n4517__, new_new_n4518__, new_new_n4519__, new_new_n4520__,
    new_new_n4521__, new_new_n4522__, new_new_n4523__, new_new_n4524__,
    new_new_n4525__, new_new_n4526__, new_new_n4527__, new_new_n4528__,
    new_new_n4529__, new_new_n4530__, new_new_n4531__, new_new_n4532__,
    new_new_n4533__, new_new_n4534__, new_new_n4535__, new_new_n4536__,
    new_new_n4537__, new_new_n4538__, new_new_n4539__, new_new_n4540__,
    new_new_n4541__, new_new_n4542__, new_new_n4543__, new_new_n4544__,
    new_new_n4545__, new_new_n4546__, new_new_n4547__, new_new_n4548__,
    new_new_n4549__, new_new_n4550__, new_new_n4551__, new_new_n4552__,
    new_new_n4553__, new_new_n4554__, new_new_n4555__, new_new_n4556__,
    new_new_n4557__, new_new_n4558__, new_new_n4559__, new_new_n4560__,
    new_new_n4561__, new_new_n4562__, new_new_n4563__, new_new_n4564__,
    new_new_n4565__, new_new_n4566__, new_new_n4567__, new_new_n4568__,
    new_new_n4570__, new_new_n4571__, new_new_n4572__, new_new_n4573__,
    new_new_n4574__, new_new_n4575__, new_new_n4576__, new_new_n4577__,
    new_new_n4578__, new_new_n4579__, new_new_n4580__, new_new_n4581__,
    new_new_n4582__, new_new_n4583__, new_new_n4584__, new_new_n4585__,
    new_new_n4586__, new_new_n4587__, new_new_n4588__, new_new_n4589__,
    new_new_n4590__, new_new_n4591__, new_new_n4592__, new_new_n4593__,
    new_new_n4594__, new_new_n4595__, new_new_n4596__, new_new_n4597__,
    new_new_n4598__, new_new_n4599__, new_new_n4600__, new_new_n4601__,
    new_new_n4602__, new_new_n4603__, new_new_n4604__, new_new_n4605__,
    new_new_n4606__, new_new_n4607__, new_new_n4608__, new_new_n4609__,
    new_new_n4610__, new_new_n4611__, new_new_n4612__, new_new_n4613__,
    new_new_n4614__, new_new_n4615__, new_new_n4616__, new_new_n4617__,
    new_new_n4618__, new_new_n4619__, new_new_n4620__, new_new_n4622__,
    new_new_n4623__, new_new_n4624__, new_new_n4625__, new_new_n4626__,
    new_new_n4627__, new_new_n4628__, new_new_n4629__, new_new_n4630__,
    new_new_n4631__, new_new_n4632__, new_new_n4633__, new_new_n4634__,
    new_new_n4635__, new_new_n4636__, new_new_n4637__, new_new_n4638__,
    new_new_n4639__, new_new_n4640__, new_new_n4641__, new_new_n4642__,
    new_new_n4643__, new_new_n4644__, new_new_n4645__, new_new_n4646__,
    new_new_n4647__, new_new_n4648__, new_new_n4649__, new_new_n4650__,
    new_new_n4651__, new_new_n4652__, new_new_n4653__, new_new_n4654__,
    new_new_n4655__, new_new_n4656__, new_new_n4657__, new_new_n4658__,
    new_new_n4659__, new_new_n4660__, new_new_n4661__, new_new_n4662__,
    new_new_n4663__, new_new_n4664__, new_new_n4665__, new_new_n4666__,
    new_new_n4667__, new_new_n4668__, new_new_n4669__, new_new_n4670__,
    new_new_n4671__, new_new_n4672__, new_new_n4673__, new_new_n4674__,
    new_new_n4675__, new_new_n4676__, new_new_n4677__, new_new_n4678__,
    new_new_n4679__, new_new_n4680__, new_new_n4681__, new_new_n4682__,
    new_new_n4683__, new_new_n4684__, new_new_n4685__, new_new_n4686__,
    new_new_n4687__, new_new_n4688__, new_new_n4689__, new_new_n4690__,
    new_new_n4691__, new_new_n4692__, new_new_n4693__, new_new_n4694__,
    new_new_n4695__, new_new_n4696__, new_new_n4697__, new_new_n4698__,
    new_new_n4699__, new_new_n4700__, new_new_n4701__, new_new_n4702__,
    new_new_n4703__, new_new_n4704__, new_new_n4705__, new_new_n4706__,
    new_new_n4707__, new_new_n4708__, new_new_n4709__, new_new_n4710__,
    new_new_n4711__, new_new_n4712__, new_new_n4713__, new_new_n4714__,
    new_new_n4715__, new_new_n4716__, new_new_n4717__, new_new_n4718__,
    new_new_n4719__, new_new_n4720__, new_new_n4721__, new_new_n4722__,
    new_new_n4723__, new_new_n4724__, new_new_n4725__, new_new_n4726__,
    new_new_n4727__, new_new_n4728__, new_new_n4729__, new_new_n4730__,
    new_new_n4731__, new_new_n4732__, new_new_n4733__, new_new_n4734__,
    new_new_n4735__, new_new_n4736__, new_new_n4737__, new_new_n4738__,
    new_new_n4739__, new_new_n4740__, new_new_n4741__, new_new_n4742__,
    new_new_n4743__, new_new_n4744__, new_new_n4745__, new_new_n4746__,
    new_new_n4747__, new_new_n4748__, new_new_n4749__, new_new_n4750__,
    new_new_n4751__, new_new_n4752__, new_new_n4753__, new_new_n4754__,
    new_new_n4755__, new_new_n4756__, new_new_n4757__, new_new_n4758__,
    new_new_n4759__, new_new_n4760__, new_new_n4761__, new_new_n4762__,
    new_new_n4763__, new_new_n4764__, new_new_n4765__, new_new_n4766__,
    new_new_n4767__, new_new_n4768__, new_new_n4769__, new_new_n4770__,
    new_new_n4771__, new_new_n4772__, new_new_n4773__, new_new_n4774__,
    new_new_n4775__, new_new_n4776__, new_new_n4777__, new_new_n4778__,
    new_new_n4779__, new_new_n4780__, new_new_n4781__, new_new_n4782__,
    new_new_n4783__, new_new_n4784__, new_new_n4785__, new_new_n4786__,
    new_new_n4787__, new_new_n4788__, new_new_n4789__, new_new_n4790__,
    new_new_n4791__, new_new_n4792__, new_new_n4793__, new_new_n4794__,
    new_new_n4795__, new_new_n4796__, new_new_n4797__, new_new_n4798__,
    new_new_n4799__, new_new_n4800__, new_new_n4801__, new_new_n4802__,
    new_new_n4803__, new_new_n4804__, new_new_n4805__, new_new_n4806__,
    new_new_n4807__, new_new_n4808__, new_new_n4809__, new_new_n4810__,
    new_new_n4811__, new_new_n4812__, new_new_n4813__, new_new_n4814__,
    new_new_n4815__, new_new_n4816__, new_new_n4817__, new_new_n4818__,
    new_new_n4819__, new_new_n4820__, new_new_n4821__, new_new_n4822__,
    new_new_n4823__, new_new_n4824__, new_new_n4825__, new_new_n4826__,
    new_new_n4827__, new_new_n4828__, new_new_n4829__, new_new_n4830__,
    new_new_n4831__, new_new_n4832__, new_new_n4833__, new_new_n4834__,
    new_new_n4835__, new_new_n4836__, new_new_n4837__, new_new_n4838__,
    new_new_n4839__, new_new_n4840__, new_new_n4841__, new_new_n4842__,
    new_new_n4843__, new_new_n4844__, new_new_n4845__, new_new_n4846__,
    new_new_n4847__, new_new_n4848__, new_new_n4849__, new_new_n4850__,
    new_new_n4851__, new_new_n4852__, new_new_n4853__, new_new_n4854__,
    new_new_n4855__, new_new_n4856__, new_new_n4857__, new_new_n4858__,
    new_new_n4859__, new_new_n4860__, new_new_n4861__, new_new_n4862__,
    new_new_n4863__, new_new_n4864__, new_new_n4865__, new_new_n4866__,
    new_new_n4867__, new_new_n4868__, new_new_n4869__, new_new_n4870__,
    new_new_n4871__, new_new_n4872__, new_new_n4873__, new_new_n4874__,
    new_new_n4875__, new_new_n4876__, new_new_n4877__, new_new_n4878__,
    new_new_n4879__, new_new_n4880__, new_new_n4881__, new_new_n4882__,
    new_new_n4883__, new_new_n4884__, new_new_n4885__, new_new_n4886__,
    new_new_n4887__, new_new_n4888__, new_new_n4889__, new_new_n4890__,
    new_new_n4891__, new_new_n4892__, new_new_n4893__, new_new_n4894__,
    new_new_n4895__, new_new_n4896__, new_new_n4897__, new_new_n4898__,
    new_new_n4899__, new_new_n4900__, new_new_n4901__, new_new_n4902__,
    new_new_n4903__, new_new_n4904__, new_new_n4905__, new_new_n4906__,
    new_new_n4907__, new_new_n4908__, new_new_n4909__, new_new_n4910__,
    new_new_n4911__, new_new_n4912__, new_new_n4913__, new_new_n4914__,
    new_new_n4915__, new_new_n4916__, new_new_n4917__, new_new_n4918__,
    new_new_n4919__, new_new_n4920__, new_new_n4921__, new_new_n4922__,
    new_new_n4923__, new_new_n4924__, new_new_n4925__, new_new_n4926__,
    new_new_n4927__, new_new_n4928__, new_new_n4929__, new_new_n4930__,
    new_new_n4931__, new_new_n4932__, new_new_n4933__, new_new_n4934__,
    new_new_n4935__, new_new_n4936__, new_new_n4937__, new_new_n4938__,
    new_new_n4939__, new_new_n4940__, new_new_n4941__, new_new_n4942__,
    new_new_n4943__, new_new_n4944__, new_new_n4945__, new_new_n4946__,
    new_new_n4947__, new_new_n4948__, new_new_n4949__, new_new_n4950__,
    new_new_n4951__, new_new_n4952__, new_new_n4953__, new_new_n4954__,
    new_new_n4955__, new_new_n4956__, new_new_n4957__, new_new_n4958__,
    new_new_n4959__, new_new_n4960__, new_new_n4961__, new_new_n4962__,
    new_new_n4963__, new_new_n4964__, new_new_n4965__, new_new_n4966__,
    new_new_n4967__, new_new_n4968__, new_new_n4969__, new_new_n4970__,
    new_new_n4971__, new_new_n4972__, new_new_n4973__, new_new_n4974__,
    new_new_n4975__, new_new_n4976__, new_new_n4977__, new_new_n4978__,
    new_new_n4979__, new_new_n4980__, new_new_n4981__, new_new_n4982__,
    new_new_n4983__, new_new_n4984__, new_new_n4985__, new_new_n4986__,
    new_new_n4987__, new_new_n4988__, new_new_n4989__, new_new_n4990__,
    new_new_n4991__, new_new_n4992__, new_new_n4993__, new_new_n4994__,
    new_new_n4995__, new_new_n4996__, new_new_n4997__, new_new_n4998__,
    new_new_n4999__, new_new_n5000__, new_new_n5001__, new_new_n5002__,
    new_new_n5003__, new_new_n5004__, new_new_n5005__, new_new_n5006__,
    new_new_n5007__, new_new_n5008__, new_new_n5009__, new_new_n5010__,
    new_new_n5011__, new_new_n5012__, new_new_n5013__, new_new_n5014__,
    new_new_n5015__, new_new_n5016__, new_new_n5017__, new_new_n5018__,
    new_new_n5019__, new_new_n5020__, new_new_n5021__, new_new_n5022__,
    new_new_n5023__, new_new_n5024__, new_new_n5025__, new_new_n5026__,
    new_new_n5027__, new_new_n5028__, new_new_n5029__, new_new_n5030__,
    new_new_n5031__, new_new_n5032__, new_new_n5033__, new_new_n5034__,
    new_new_n5035__, new_new_n5036__, new_new_n5037__, new_new_n5038__,
    new_new_n5039__, new_new_n5040__, new_new_n5041__, new_new_n5042__,
    new_new_n5043__, new_new_n5044__, new_new_n5045__, new_new_n5046__,
    new_new_n5047__, new_new_n5048__, new_new_n5049__, new_new_n5050__,
    new_new_n5051__, new_new_n5052__, new_new_n5053__, new_new_n5054__,
    new_new_n5055__, new_new_n5056__, new_new_n5057__, new_new_n5058__,
    new_new_n5059__, new_new_n5060__, new_new_n5061__, new_new_n5062__,
    new_new_n5063__, new_new_n5064__, new_new_n5065__, new_new_n5066__,
    new_new_n5067__, new_new_n5068__, new_new_n5069__, new_new_n5070__,
    new_new_n5071__, new_new_n5072__, new_new_n5073__, new_new_n5074__,
    new_new_n5075__, new_new_n5076__, new_new_n5077__, new_new_n5078__,
    new_new_n5079__, new_new_n5080__, new_new_n5081__, new_new_n5082__,
    new_new_n5083__, new_new_n5084__, new_new_n5085__, new_new_n5086__,
    new_new_n5087__, new_new_n5088__, new_new_n5089__, new_new_n5090__,
    new_new_n5091__, new_new_n5092__, new_new_n5093__, new_new_n5094__,
    new_new_n5095__, new_new_n5096__, new_new_n5097__, new_new_n5098__,
    new_new_n5099__, new_new_n5100__, new_new_n5101__, new_new_n5102__,
    new_new_n5103__, new_new_n5104__, new_new_n5105__, new_new_n5106__,
    new_new_n5107__, new_new_n5108__, new_new_n5109__, new_new_n5110__,
    new_new_n5111__, new_new_n5112__, new_new_n5113__, new_new_n5114__,
    new_new_n5115__, new_new_n5116__, new_new_n5117__, new_new_n5118__,
    new_new_n5119__, new_new_n5120__, new_new_n5121__, new_new_n5122__,
    new_new_n5123__, new_new_n5124__, new_new_n5125__, new_new_n5126__,
    new_new_n5127__, new_new_n5128__, new_new_n5129__, new_new_n5130__,
    new_new_n5131__, new_new_n5132__, new_new_n5133__, new_new_n5134__,
    new_new_n5135__, new_new_n5136__, new_new_n5137__, new_new_n5138__,
    new_new_n5139__, new_new_n5140__, new_new_n5141__, new_new_n5142__,
    new_new_n5143__, new_new_n5144__, new_new_n5145__, new_new_n5146__,
    new_new_n5147__, new_new_n5148__, new_new_n5149__, new_new_n5150__,
    new_new_n5151__, new_new_n5152__, new_new_n5153__, new_new_n5154__,
    new_new_n5155__, new_new_n5156__, new_new_n5157__, new_new_n5158__,
    new_new_n5159__, new_new_n5160__, new_new_n5161__, new_new_n5162__,
    new_new_n5163__, new_new_n5164__, new_new_n5165__, new_new_n5166__,
    new_new_n5167__, new_new_n5168__, new_new_n5169__, new_new_n5170__,
    new_new_n5171__, new_new_n5172__, new_new_n5173__, new_new_n5174__,
    new_new_n5175__, new_new_n5176__, new_new_n5177__, new_new_n5178__,
    new_new_n5179__, new_new_n5180__, new_new_n5181__, new_new_n5182__,
    new_new_n5183__, new_new_n5184__, new_new_n5185__, new_new_n5186__,
    new_new_n5187__, new_new_n5188__, new_new_n5189__, new_new_n5190__,
    new_new_n5191__, new_new_n5192__, new_new_n5193__, new_new_n5194__,
    new_new_n5195__, new_new_n5196__, new_new_n5197__, new_new_n5198__,
    new_new_n5199__, new_new_n5200__, new_new_n5201__, new_new_n5202__,
    new_new_n5203__, new_new_n5204__, new_new_n5205__, new_new_n5206__,
    new_new_n5207__, new_new_n5208__, new_new_n5209__, new_new_n5210__,
    new_new_n5211__, new_new_n5212__, new_new_n5213__, new_new_n5214__,
    new_new_n5215__, new_new_n5216__, new_new_n5217__, new_new_n5218__,
    new_new_n5219__, new_new_n5220__, new_new_n5221__, new_new_n5222__,
    new_new_n5223__, new_new_n5224__, new_new_n5225__, new_new_n5226__,
    new_new_n5227__, new_new_n5228__, new_new_n5229__, new_new_n5230__,
    new_new_n5231__, new_new_n5232__, new_new_n5233__, new_new_n5234__,
    new_new_n5235__, new_new_n5236__, new_new_n5237__, new_new_n5238__,
    new_new_n5239__, new_new_n5240__, new_new_n5241__, new_new_n5242__,
    new_new_n5243__, new_new_n5244__, new_new_n5245__, new_new_n5246__,
    new_new_n5247__, new_new_n5248__, new_new_n5249__, new_new_n5250__,
    new_new_n5251__, new_new_n5252__, new_new_n5253__, new_new_n5254__,
    new_new_n5255__, new_new_n5256__, new_new_n5257__, new_new_n5258__,
    new_new_n5259__, new_new_n5260__, new_new_n5261__, new_new_n5262__,
    new_new_n5263__, new_new_n5264__, new_new_n5265__, new_new_n5266__,
    new_new_n5267__, new_new_n5268__, new_new_n5269__, new_new_n5270__,
    new_new_n5271__, new_new_n5272__, new_new_n5273__, new_new_n5274__,
    new_new_n5275__, new_new_n5276__, new_new_n5277__, new_new_n5278__,
    new_new_n5279__, new_new_n5280__, new_new_n5281__, new_new_n5282__,
    new_new_n5283__, new_new_n5284__, new_new_n5285__, new_new_n5286__,
    new_new_n5287__, new_new_n5288__, new_new_n5289__, new_new_n5290__,
    new_new_n5291__, new_new_n5292__, new_new_n5293__, new_new_n5294__,
    new_new_n5295__, new_new_n5296__, new_new_n5297__, new_new_n5298__,
    new_new_n5299__, new_new_n5300__, new_new_n5301__, new_new_n5302__,
    new_new_n5303__, new_new_n5304__, new_new_n5305__, new_new_n5306__,
    new_new_n5307__, new_new_n5308__, new_new_n5309__, new_new_n5310__,
    new_new_n5311__, new_new_n5312__, new_new_n5313__, new_new_n5314__,
    new_new_n5315__, new_new_n5316__, new_new_n5317__, new_new_n5318__,
    new_new_n5319__, new_new_n5320__, new_new_n5321__, new_new_n5322__,
    new_new_n5323__, new_new_n5324__, new_new_n5325__, new_new_n5326__,
    new_new_n5327__, new_new_n5328__, new_new_n5329__, new_new_n5330__,
    new_new_n5331__, new_new_n5332__, new_new_n5333__, new_new_n5334__,
    new_new_n5335__, new_new_n5336__, new_new_n5337__, new_new_n5338__,
    new_new_n5339__, new_new_n5340__, new_new_n5341__, new_new_n5342__,
    new_new_n5343__, new_new_n5344__, new_new_n5345__, new_new_n5346__,
    new_new_n5347__, new_new_n5348__, new_new_n5349__, new_new_n5350__,
    new_new_n5351__, new_new_n5352__, new_new_n5353__, new_new_n5354__,
    new_new_n5355__, new_new_n5356__, new_new_n5357__, new_new_n5358__,
    new_new_n5359__, new_new_n5360__, new_new_n5361__, new_new_n5362__,
    new_new_n5363__, new_new_n5364__, new_new_n5365__, new_new_n5366__,
    new_new_n5367__, new_new_n5368__, new_new_n5369__, new_new_n5370__,
    new_new_n5371__, new_new_n5372__, new_new_n5373__, new_new_n5374__,
    new_new_n5375__, new_new_n5376__, new_new_n5377__, new_new_n5378__,
    new_new_n5379__, new_new_n5380__, new_new_n5381__, new_new_n5382__,
    new_new_n5383__, new_new_n5384__, new_new_n5385__, new_new_n5386__,
    new_new_n5387__, new_new_n5388__, new_new_n5389__, new_new_n5390__,
    new_new_n5391__, new_new_n5392__, new_new_n5393__, new_new_n5394__,
    new_new_n5395__, new_new_n5396__, new_new_n5397__, new_new_n5398__,
    new_new_n5399__, new_new_n5400__, new_new_n5401__, new_new_n5402__,
    new_new_n5403__, new_new_n5404__, new_new_n5405__, new_new_n5406__,
    new_new_n5407__, new_new_n5408__, new_new_n5409__, new_new_n5410__,
    new_new_n5411__, new_new_n5412__, new_new_n5413__, new_new_n5414__,
    new_new_n5415__, new_new_n5416__, new_new_n5417__, new_new_n5418__,
    new_new_n5419__, new_new_n5420__, new_new_n5421__, new_new_n5422__,
    new_new_n5423__, new_new_n5424__, new_new_n5425__, new_new_n5426__,
    new_new_n5427__, new_new_n5428__, new_new_n5429__, new_new_n5430__,
    new_new_n5431__, new_new_n5432__, new_new_n5433__, new_new_n5434__,
    new_new_n5435__, new_new_n5436__, new_new_n5437__, new_new_n5438__,
    new_new_n5439__, new_new_n5440__, new_new_n5441__, new_new_n5442__,
    new_new_n5443__, new_new_n5444__, new_new_n5445__, new_new_n5446__,
    new_new_n5447__, new_new_n5448__, new_new_n5449__, new_new_n5450__,
    new_new_n5451__, new_new_n5452__, new_new_n5453__, new_new_n5454__,
    new_new_n5455__, new_new_n5456__, new_new_n5457__, new_new_n5458__,
    new_new_n5459__, new_new_n5460__, new_new_n5461__, new_new_n5462__,
    new_new_n5463__, new_new_n5464__, new_new_n5465__, new_new_n5466__,
    new_new_n5467__, new_new_n5468__, new_new_n5469__, new_new_n5470__,
    new_new_n5471__, new_new_n5472__, new_new_n5473__, new_new_n5474__,
    new_new_n5475__, new_new_n5476__, new_new_n5477__, new_new_n5478__,
    new_new_n5479__, new_new_n5480__, new_new_n5481__, new_new_n5482__,
    new_new_n5483__, new_new_n5484__, new_new_n5485__, new_new_n5486__,
    new_new_n5487__, new_new_n5488__, new_new_n5489__, new_new_n5490__,
    new_new_n5491__, new_new_n5492__, new_new_n5493__, new_new_n5494__,
    new_new_n5495__, new_new_n5496__, new_new_n5497__, new_new_n5498__,
    new_new_n5499__, new_new_n5500__, new_new_n5501__, new_new_n5502__,
    new_new_n5503__, new_new_n5504__, new_new_n5505__, new_new_n5506__,
    new_new_n5507__, new_new_n5508__, new_new_n5509__, new_new_n5510__,
    new_new_n5511__, new_new_n5512__, new_new_n5513__, new_new_n5514__,
    new_new_n5515__, new_new_n5516__, new_new_n5517__, new_new_n5518__,
    new_new_n5519__, new_new_n5520__, new_new_n5521__, new_new_n5522__,
    new_new_n5523__, new_new_n5524__, new_new_n5525__, new_new_n5526__,
    new_new_n5527__, new_new_n5528__, new_new_n5529__, new_new_n5530__,
    new_new_n5531__, new_new_n5532__, new_new_n5533__, new_new_n5534__,
    new_new_n5535__, new_new_n5536__, new_new_n5537__, new_new_n5538__,
    new_new_n5539__, new_new_n5540__, new_new_n5541__, new_new_n5542__,
    new_new_n5543__, new_new_n5544__, new_new_n5545__, new_new_n5546__,
    new_new_n5547__, new_new_n5548__, new_new_n5549__, new_new_n5550__,
    new_new_n5551__, new_new_n5552__, new_new_n5553__, new_new_n5554__,
    new_new_n5555__, new_new_n5556__, new_new_n5557__, new_new_n5558__,
    new_new_n5559__, new_new_n5560__, new_new_n5561__, new_new_n5562__,
    new_new_n5563__, new_new_n5564__, new_new_n5565__, new_new_n5566__,
    new_new_n5567__, new_new_n5568__, new_new_n5569__, new_new_n5570__,
    new_new_n5571__, new_new_n5572__, new_new_n5573__, new_new_n5574__,
    new_new_n5575__, new_new_n5576__, new_new_n5577__, new_new_n5578__,
    new_new_n5579__, new_new_n5580__, new_new_n5581__, new_new_n5582__,
    new_new_n5583__, new_new_n5584__, new_new_n5585__, new_new_n5586__,
    new_new_n5587__, new_new_n5588__, new_new_n5589__, new_new_n5590__,
    new_new_n5591__, new_new_n5592__, new_new_n5593__, new_new_n5594__,
    new_new_n5595__, new_new_n5596__, new_new_n5597__, new_new_n5598__,
    new_new_n5599__, new_new_n5600__, new_new_n5601__, new_new_n5602__,
    new_new_n5603__, new_new_n5604__, new_new_n5605__, new_new_n5606__,
    new_new_n5607__, new_new_n5608__, new_new_n5609__, new_new_n5610__,
    new_new_n5611__, new_new_n5612__, new_new_n5613__, new_new_n5614__,
    new_new_n5615__, new_new_n5616__, new_new_n5617__, new_new_n5618__,
    new_new_n5619__, new_new_n5620__, new_new_n5621__, new_new_n5622__,
    new_new_n5623__, new_new_n5624__, new_new_n5625__, new_new_n5626__,
    new_new_n5627__, new_new_n5628__, new_new_n5629__, new_new_n5630__,
    new_new_n5631__, new_new_n5632__, new_new_n5633__, new_new_n5634__,
    new_new_n5635__, new_new_n5636__, new_new_n5637__, new_new_n5638__,
    new_new_n5639__, new_new_n5640__, new_new_n5641__, new_new_n5642__,
    new_new_n5643__, new_new_n5644__, new_new_n5645__, new_new_n5646__,
    new_new_n5647__, new_new_n5648__, new_new_n5649__, new_new_n5650__,
    new_new_n5651__, new_new_n5652__, new_new_n5653__, new_new_n5654__,
    new_new_n5655__, new_new_n5656__, new_new_n5657__, new_new_n5658__,
    new_new_n5659__, new_new_n5660__, new_new_n5661__, new_new_n5662__,
    new_new_n5663__, new_new_n5664__, new_new_n5665__, new_new_n5666__,
    new_new_n5667__, new_new_n5668__, new_new_n5669__, new_new_n5670__,
    new_new_n5671__, new_new_n5672__, new_new_n5673__, new_new_n5674__,
    new_new_n5675__, new_new_n5676__, new_new_n5677__, new_new_n5678__,
    new_new_n5679__, new_new_n5680__, new_new_n5681__, new_new_n5682__,
    new_new_n5683__, new_new_n5684__, new_new_n5685__, new_new_n5686__,
    new_new_n5687__, new_new_n5688__, new_new_n5689__, new_new_n5690__,
    new_new_n5691__, new_new_n5692__, new_new_n5693__, new_new_n5694__,
    new_new_n5695__, new_new_n5696__, new_new_n5697__, new_new_n5698__,
    new_new_n5699__, new_new_n5700__, new_new_n5701__, new_new_n5702__,
    new_new_n5703__, new_new_n5704__, new_new_n5705__, new_new_n5706__,
    new_new_n5707__, new_new_n5708__, new_new_n5709__, new_new_n5710__,
    new_new_n5711__, new_new_n5712__, new_new_n5713__, new_new_n5714__,
    new_new_n5715__, new_new_n5716__, new_new_n5717__, new_new_n5718__,
    new_new_n5719__, new_new_n5720__, new_new_n5721__, new_new_n5722__,
    new_new_n5723__, new_new_n5724__, new_new_n5725__, new_new_n5726__,
    new_new_n5727__, new_new_n5728__, new_new_n5729__, new_new_n5730__,
    new_new_n5731__, new_new_n5732__, new_new_n5733__, new_new_n5734__,
    new_new_n5735__, new_new_n5736__, new_new_n5737__, new_new_n5738__,
    new_new_n5739__, new_new_n5740__, new_new_n5741__, new_new_n5742__,
    new_new_n5743__, new_new_n5744__, new_new_n5745__, new_new_n5746__,
    new_new_n5747__, new_new_n5748__, new_new_n5749__, new_new_n5750__,
    new_new_n5751__, new_new_n5752__, new_new_n5753__, new_new_n5754__,
    new_new_n5755__, new_new_n5756__, new_new_n5757__, new_new_n5758__,
    new_new_n5759__, new_new_n5760__, new_new_n5761__, new_new_n5762__,
    new_new_n5763__, new_new_n5764__, new_new_n5765__, new_new_n5766__,
    new_new_n5767__, new_new_n5768__, new_new_n5769__, new_new_n5770__,
    new_new_n5771__, new_new_n5772__, new_new_n5773__, new_new_n5774__,
    new_new_n5775__, new_new_n5776__, new_new_n5777__, new_new_n5778__,
    new_new_n5779__, new_new_n5780__, new_new_n5781__, new_new_n5782__,
    new_new_n5783__, new_new_n5784__, new_new_n5785__, new_new_n5786__,
    new_new_n5787__, new_new_n5788__, new_new_n5789__, new_new_n5790__,
    new_new_n5791__, new_new_n5792__, new_new_n5793__, new_new_n5794__,
    new_new_n5795__, new_new_n5796__, new_new_n5797__, new_new_n5798__,
    new_new_n5799__, new_new_n5800__, new_new_n5801__, new_new_n5802__,
    new_new_n5803__, new_new_n5804__, new_new_n5805__, new_new_n5806__,
    new_new_n5807__, new_new_n5808__, new_new_n5809__, new_new_n5810__,
    new_new_n5811__, new_new_n5812__, new_new_n5813__, new_new_n5814__,
    new_new_n5815__, new_new_n5816__, new_new_n5817__, new_new_n5818__,
    new_new_n5819__, new_new_n5820__, new_new_n5821__, new_new_n5822__,
    new_new_n5823__, new_new_n5824__, new_new_n5825__, new_new_n5826__,
    new_new_n5827__, new_new_n5828__, new_new_n5829__, new_new_n5830__,
    new_new_n5831__, new_new_n5832__, new_new_n5833__, new_new_n5834__,
    new_new_n5835__, new_new_n5836__, new_new_n5837__, new_new_n5838__,
    new_new_n5839__, new_new_n5840__, new_new_n5841__, new_new_n5842__,
    new_new_n5843__, new_new_n5844__, new_new_n5845__, new_new_n5846__,
    new_new_n5847__, new_new_n5848__, new_new_n5849__, new_new_n5850__,
    new_new_n5851__, new_new_n5852__, new_new_n5853__, new_new_n5854__,
    new_new_n5855__, new_new_n5856__, new_new_n5857__, new_new_n5858__,
    new_new_n5859__, new_new_n5860__, new_new_n5861__, new_new_n5862__,
    new_new_n5863__, new_new_n5864__, new_new_n5865__, new_new_n5866__,
    new_new_n5867__, new_new_n5868__, new_new_n5869__, new_new_n5870__,
    new_new_n5871__, new_new_n5872__, new_new_n5873__, new_new_n5874__,
    new_new_n5875__, new_new_n5876__, new_new_n5877__, new_new_n5878__,
    new_new_n5879__, new_new_n5880__, new_new_n5881__, new_new_n5882__,
    new_new_n5883__, new_new_n5884__, new_new_n5885__, new_new_n5886__,
    new_new_n5887__, new_new_n5888__, new_new_n5889__, new_new_n5890__,
    new_new_n5891__, new_new_n5892__, new_new_n5893__, new_new_n5894__,
    new_new_n5895__, new_new_n5896__, new_new_n5897__, new_new_n5898__,
    new_new_n5899__, new_new_n5900__, new_new_n5901__, new_new_n5902__,
    new_new_n5903__, new_new_n5904__, new_new_n5905__, new_new_n5906__,
    new_new_n5907__, new_new_n5908__, new_new_n5909__, new_new_n5910__,
    new_new_n5911__, new_new_n5912__, new_new_n5913__, new_new_n5914__,
    new_new_n5915__, new_new_n5916__, new_new_n5917__, new_new_n5918__,
    new_new_n5919__, new_new_n5920__, new_new_n5921__, new_new_n5922__,
    new_new_n5923__, new_new_n5924__, new_new_n5925__, new_new_n5926__,
    new_new_n5927__, new_new_n5928__, new_new_n5929__, new_new_n5930__,
    new_new_n5931__, new_new_n5932__, new_new_n5933__, new_new_n5934__,
    new_new_n5935__, new_new_n5936__, new_new_n5937__, new_new_n5938__,
    new_new_n5939__, new_new_n5940__, new_new_n5941__, new_new_n5942__,
    new_new_n5943__, new_new_n5944__, new_new_n5945__, new_new_n5946__,
    new_new_n5947__, new_new_n5948__, new_new_n5949__, new_new_n5950__,
    new_new_n5951__, new_new_n5952__, new_new_n5953__, new_new_n5954__,
    new_new_n5955__, new_new_n5956__, new_new_n5957__, new_new_n5958__,
    new_new_n5959__, new_new_n5960__, new_new_n5961__, new_new_n5962__,
    new_new_n5963__, new_new_n5964__, new_new_n5965__, new_new_n5966__,
    new_new_n5967__, new_new_n5968__, new_new_n5969__, new_new_n5970__,
    new_new_n5971__, new_new_n5972__, new_new_n5973__, new_new_n5974__,
    new_new_n5975__, new_new_n5976__, new_new_n5977__, new_new_n5978__,
    new_new_n5979__, new_new_n5980__, new_new_n5981__, new_new_n5982__,
    new_new_n5983__, new_new_n5984__, new_new_n5985__, new_new_n5986__,
    new_new_n5987__, new_new_n5988__, new_new_n5989__, new_new_n5990__,
    new_new_n5991__, new_new_n5992__, new_new_n5993__, new_new_n5994__,
    new_new_n5995__, new_new_n5996__, new_new_n5997__, new_new_n5998__,
    new_new_n5999__, new_new_n6000__, new_new_n6001__, new_new_n6002__,
    new_new_n6003__, new_new_n6004__, new_new_n6005__, new_new_n6006__,
    new_new_n6007__, new_new_n6008__, new_new_n6009__, new_new_n6010__,
    new_new_n6011__, new_new_n6012__, new_new_n6013__, new_new_n6014__,
    new_new_n6015__, new_new_n6016__, new_new_n6017__, new_new_n6018__,
    new_new_n6019__, new_new_n6020__, new_new_n6021__, new_new_n6022__,
    new_new_n6023__, new_new_n6024__, new_new_n6025__, new_new_n6026__,
    new_new_n6027__, new_new_n6028__, new_new_n6029__, new_new_n6030__,
    new_new_n6031__, new_new_n6032__, new_new_n6033__, new_new_n6034__,
    new_new_n6035__, new_new_n6036__, new_new_n6037__, new_new_n6038__,
    new_new_n6039__, new_new_n6040__, new_new_n6041__, new_new_n6042__,
    new_new_n6043__, new_new_n6044__, new_new_n6045__, new_new_n6046__,
    new_new_n6047__, new_new_n6048__, new_new_n6049__, new_new_n6050__,
    new_new_n6051__, new_new_n6052__, new_new_n6053__, new_new_n6054__,
    new_new_n6055__, new_new_n6056__, new_new_n6057__, new_new_n6058__,
    new_new_n6059__, new_new_n6060__, new_new_n6061__, new_new_n6062__,
    new_new_n6063__, new_new_n6064__, new_new_n6065__, new_new_n6066__,
    new_new_n6067__, new_new_n6068__, new_new_n6069__, new_new_n6070__,
    new_new_n6071__, new_new_n6072__, new_new_n6073__, new_new_n6074__,
    new_new_n6075__, new_new_n6076__, new_new_n6077__, new_new_n6078__,
    new_new_n6079__, new_new_n6080__, new_new_n6081__, new_new_n6082__,
    new_new_n6083__, new_new_n6084__, new_new_n6085__, new_new_n6086__,
    new_new_n6087__, new_new_n6088__, new_new_n6089__, new_new_n6090__,
    new_new_n6091__, new_new_n6092__, new_new_n6093__, new_new_n6094__,
    new_new_n6095__, new_new_n6096__, new_new_n6097__, new_new_n6098__,
    new_new_n6099__, new_new_n6100__, new_new_n6101__, new_new_n6102__,
    new_new_n6103__, new_new_n6104__, new_new_n6105__, new_new_n6106__,
    new_new_n6107__, new_new_n6108__, new_new_n6109__, new_new_n6110__,
    new_new_n6111__, new_new_n6112__, new_new_n6113__, new_new_n6114__,
    new_new_n6115__, new_new_n6116__, new_new_n6117__, new_new_n6118__,
    new_new_n6119__, new_new_n6120__, new_new_n6121__, new_new_n6122__,
    new_new_n6123__, new_new_n6124__, new_new_n6125__, new_new_n6126__,
    new_new_n6127__, new_new_n6128__, new_new_n6129__, new_new_n6130__,
    new_new_n6131__, new_new_n6132__, new_new_n6133__, new_new_n6134__,
    new_new_n6135__, new_new_n6136__, new_new_n6137__, new_new_n6138__,
    new_new_n6139__, new_new_n6140__, new_new_n6141__, new_new_n6142__,
    new_new_n6143__, new_new_n6144__, new_new_n6145__, new_new_n6146__,
    new_new_n6147__, new_new_n6148__, new_new_n6149__, new_new_n6150__,
    new_new_n6151__, new_new_n6152__, new_new_n6153__, new_new_n6154__,
    new_new_n6155__, new_new_n6156__, new_new_n6157__, new_new_n6158__,
    new_new_n6159__, new_new_n6160__, new_new_n6161__, new_new_n6162__,
    new_new_n6163__, new_new_n6164__, new_new_n6165__, new_new_n6166__,
    new_new_n6167__, new_new_n6168__, new_new_n6169__, new_new_n6170__,
    new_new_n6171__, new_new_n6172__, new_new_n6173__, new_new_n6174__,
    new_new_n6175__, new_new_n6176__, new_new_n6177__, new_new_n6178__,
    new_new_n6179__, new_new_n6180__, new_new_n6181__, new_new_n6182__,
    new_new_n6183__, new_new_n6184__, new_new_n6185__, new_new_n6186__,
    new_new_n6187__, new_new_n6188__, new_new_n6189__, new_new_n6190__,
    new_new_n6191__, new_new_n6192__, new_new_n6193__, new_new_n6194__,
    new_new_n6195__, new_new_n6196__, new_new_n6197__, new_new_n6198__,
    new_new_n6199__, new_new_n6200__, new_new_n6201__, new_new_n6202__,
    new_new_n6203__, new_new_n6204__, new_new_n6205__, new_new_n6206__,
    new_new_n6207__, new_new_n6208__, new_new_n6209__, new_new_n6210__,
    new_new_n6211__, new_new_n6212__, new_new_n6213__, new_new_n6214__,
    new_new_n6215__, new_new_n6216__, new_new_n6217__, new_new_n6218__,
    new_new_n6219__, new_new_n6220__, new_new_n6221__, new_new_n6222__,
    new_new_n6223__, new_new_n6224__, new_new_n6225__, new_new_n6226__,
    new_new_n6227__, new_new_n6228__, new_new_n6229__, new_new_n6230__,
    new_new_n6231__, new_new_n6232__, new_new_n6233__, new_new_n6234__,
    new_new_n6235__, new_new_n6236__, new_new_n6237__, new_new_n6238__,
    new_new_n6239__, new_new_n6240__, new_new_n6241__, new_new_n6242__,
    new_new_n6243__, new_new_n6244__, new_new_n6245__, new_new_n6246__,
    new_new_n6247__, new_new_n6248__, new_new_n6249__, new_new_n6250__,
    new_new_n6251__, new_new_n6252__, new_new_n6253__, new_new_n6254__,
    new_new_n6255__, new_new_n6256__, new_new_n6257__, new_new_n6258__,
    new_new_n6259__, new_new_n6260__, new_new_n6261__, new_new_n6262__,
    new_new_n6263__, new_new_n6264__, new_new_n6265__, new_new_n6266__,
    new_new_n6267__, new_new_n6268__, new_new_n6269__, new_new_n6270__,
    new_new_n6271__, new_new_n6272__, new_new_n6273__, new_new_n6274__,
    new_new_n6275__, new_new_n6276__, new_new_n6277__, new_new_n6278__,
    new_new_n6279__, new_new_n6280__, new_new_n6281__, new_new_n6282__,
    new_new_n6283__, new_new_n6284__, new_new_n6285__, new_new_n6286__,
    new_new_n6287__, new_new_n6288__, new_new_n6289__, new_new_n6290__,
    new_new_n6291__, new_new_n6292__, new_new_n6293__, new_new_n6294__,
    new_new_n6295__, new_new_n6296__, new_new_n6297__, new_new_n6298__,
    new_new_n6299__, new_new_n6300__, new_new_n6301__, new_new_n6302__,
    new_new_n6303__, new_new_n6304__, new_new_n6305__, new_new_n6306__,
    new_new_n6307__, new_new_n6308__, new_new_n6309__, new_new_n6310__,
    new_new_n6311__, new_new_n6312__, new_new_n6313__, new_new_n6314__,
    new_new_n6315__, new_new_n6316__, new_new_n6317__, new_new_n6318__,
    new_new_n6319__, new_new_n6320__, new_new_n6321__, new_new_n6322__,
    new_new_n6323__, new_new_n6324__, new_new_n6325__, new_new_n6326__,
    new_new_n6327__, new_new_n6328__, new_new_n6329__, new_new_n6330__,
    new_new_n6331__, new_new_n6332__, new_new_n6333__, new_new_n6334__,
    new_new_n6335__, new_new_n6336__, new_new_n6337__, new_new_n6338__,
    new_new_n6339__, new_new_n6340__, new_new_n6341__, new_new_n6342__,
    new_new_n6343__, new_new_n6344__, new_new_n6345__, new_new_n6346__,
    new_new_n6347__, new_new_n6348__, new_new_n6349__, new_new_n6350__,
    new_new_n6351__, new_new_n6352__, new_new_n6353__, new_new_n6354__,
    new_new_n6355__, new_new_n6356__, new_new_n6357__, new_new_n6358__,
    new_new_n6359__, new_new_n6360__, new_new_n6361__, new_new_n6362__,
    new_new_n6363__, new_new_n6364__, new_new_n6365__, new_new_n6366__,
    new_new_n6367__, new_new_n6368__, new_new_n6369__, new_new_n6370__,
    new_new_n6371__, new_new_n6372__, new_new_n6373__, new_new_n6374__,
    new_new_n6375__, new_new_n6376__, new_new_n6377__, new_new_n6378__,
    new_new_n6379__, new_new_n6380__, new_new_n6381__, new_new_n6382__,
    new_new_n6383__, new_new_n6384__, new_new_n6385__, new_new_n6386__,
    new_new_n6387__, new_new_n6388__, new_new_n6389__, new_new_n6390__,
    new_new_n6391__, new_new_n6392__, new_new_n6393__, new_new_n6394__,
    new_new_n6395__, new_new_n6396__, new_new_n6397__, new_new_n6398__,
    new_new_n6399__, new_new_n6400__, new_new_n6401__, new_new_n6402__,
    new_new_n6403__, new_new_n6404__, new_new_n6405__, new_new_n6406__,
    new_new_n6407__, new_new_n6408__, new_new_n6409__, new_new_n6410__,
    new_new_n6411__, new_new_n6412__, new_new_n6413__, new_new_n6414__,
    new_new_n6415__, new_new_n6416__, new_new_n6417__, new_new_n6418__,
    new_new_n6419__, new_new_n6420__, new_new_n6421__, new_new_n6422__,
    new_new_n6423__, new_new_n6424__, new_new_n6425__, new_new_n6426__,
    new_new_n6427__, new_new_n6428__, new_new_n6429__, new_new_n6430__,
    new_new_n6431__, new_new_n6432__, new_new_n6433__, new_new_n6434__,
    new_new_n6435__, new_new_n6436__, new_new_n6437__, new_new_n6438__,
    new_new_n6439__, new_new_n6440__, new_new_n6441__, new_new_n6442__,
    new_new_n6443__, new_new_n6444__, new_new_n6445__, new_new_n6446__,
    new_new_n6447__, new_new_n6448__, new_new_n6449__, new_new_n6450__,
    new_new_n6451__, new_new_n6452__, new_new_n6453__, new_new_n6454__,
    new_new_n6455__, new_new_n6456__, new_new_n6457__, new_new_n6458__,
    new_new_n6459__, new_new_n6460__, new_new_n6461__, new_new_n6462__,
    new_new_n6463__, new_new_n6464__, new_new_n6465__, new_new_n6466__,
    new_new_n6467__, new_new_n6468__, new_new_n6469__, new_new_n6470__,
    new_new_n6471__, new_new_n6472__, new_new_n6473__, new_new_n6474__,
    new_new_n6475__, new_new_n6476__, new_new_n6477__, new_new_n6478__,
    new_new_n6479__, new_new_n6480__, new_new_n6481__, new_new_n6482__,
    new_new_n6483__, new_new_n6484__, new_new_n6485__, new_new_n6486__,
    new_new_n6487__, new_new_n6488__, new_new_n6489__, new_new_n6490__,
    new_new_n6491__, new_new_n6492__, new_new_n6493__, new_new_n6494__,
    new_new_n6495__, new_new_n6496__, new_new_n6497__, new_new_n6498__,
    new_new_n6499__, new_new_n6500__, new_new_n6501__, new_new_n6502__,
    new_new_n6503__, new_new_n6504__, new_new_n6505__, new_new_n6506__,
    new_new_n6507__, new_new_n6508__, new_new_n6509__, new_new_n6510__,
    new_new_n6511__, new_new_n6512__, new_new_n6513__, new_new_n6514__,
    new_new_n6515__, new_new_n6516__, new_new_n6517__, new_new_n6518__,
    new_new_n6519__, new_new_n6520__, new_new_n6521__, new_new_n6522__,
    new_new_n6523__, new_new_n6524__, new_new_n6525__, new_new_n6526__,
    new_new_n6527__, new_new_n6528__, new_new_n6529__, new_new_n6530__,
    new_new_n6531__, new_new_n6532__, new_new_n6533__, new_new_n6534__,
    new_new_n6535__, new_new_n6536__, new_new_n6537__, new_new_n6538__,
    new_new_n6539__, new_new_n6540__, new_new_n6541__, new_new_n6542__,
    new_new_n6543__, new_new_n6544__, new_new_n6545__, new_new_n6546__,
    new_new_n6547__, new_new_n6548__, new_new_n6549__, new_new_n6550__,
    new_new_n6551__, new_new_n6552__, new_new_n6553__, new_new_n6554__,
    new_new_n6555__, new_new_n6556__, new_new_n6557__, new_new_n6558__,
    new_new_n6559__, new_new_n6560__, new_new_n6561__, new_new_n6562__,
    new_new_n6563__, new_new_n6564__, new_new_n6565__, new_new_n6566__,
    new_new_n6567__, new_new_n6568__, new_new_n6569__, new_new_n6570__,
    new_new_n6571__, new_new_n6572__, new_new_n6573__, new_new_n6574__,
    new_new_n6575__, new_new_n6576__, new_new_n6577__, new_new_n6578__,
    new_new_n6579__, new_new_n6580__, new_new_n6581__, new_new_n6582__,
    new_new_n6583__, new_new_n6584__, new_new_n6585__, new_new_n6586__,
    new_new_n6587__, new_new_n6588__, new_new_n6589__, new_new_n6590__,
    new_new_n6591__, new_new_n6592__, new_new_n6593__, new_new_n6594__,
    new_new_n6595__, new_new_n6596__, new_new_n6597__, new_new_n6598__,
    new_new_n6599__, new_new_n6600__, new_new_n6601__, new_new_n6602__,
    new_new_n6603__, new_new_n6604__, new_new_n6605__, new_new_n6606__,
    new_new_n6607__, new_new_n6608__, new_new_n6609__, new_new_n6610__,
    new_new_n6611__, new_new_n6612__, new_new_n6613__, new_new_n6614__,
    new_new_n6615__, new_new_n6616__, new_new_n6617__, new_new_n6618__,
    new_new_n6619__, new_new_n6620__, new_new_n6621__, new_new_n6622__,
    new_new_n6623__, new_new_n6624__, new_new_n6625__, new_new_n6626__,
    new_new_n6627__, new_new_n6628__, new_new_n6629__, new_new_n6630__,
    new_new_n6631__, new_new_n6632__, new_new_n6633__, new_new_n6634__,
    new_new_n6635__, new_new_n6636__, new_new_n6637__, new_new_n6638__,
    new_new_n6639__, new_new_n6640__, new_new_n6641__, new_new_n6642__,
    new_new_n6643__, new_new_n6644__, new_new_n6645__, new_new_n6646__,
    new_new_n6647__, new_new_n6648__, new_new_n6649__, new_new_n6650__,
    new_new_n6651__, new_new_n6652__, new_new_n6653__, new_new_n6654__,
    new_new_n6655__, new_new_n6656__, new_new_n6657__, new_new_n6658__,
    new_new_n6659__, new_new_n6660__, new_new_n6661__, new_new_n6662__,
    new_new_n6663__, new_new_n6664__, new_new_n6665__, new_new_n6666__,
    new_new_n6667__, new_new_n6668__, new_new_n6669__, new_new_n6670__,
    new_new_n6671__, new_new_n6672__, new_new_n6673__, new_new_n6674__,
    new_new_n6675__, new_new_n6676__, new_new_n6677__, new_new_n6678__,
    new_new_n6679__, new_new_n6680__, new_new_n6681__, new_new_n6682__,
    new_new_n6683__, new_new_n6684__, new_new_n6685__, new_new_n6686__,
    new_new_n6687__, new_new_n6688__, new_new_n6689__, new_new_n6690__,
    new_new_n6691__, new_new_n6692__, new_new_n6693__, new_new_n6694__,
    new_new_n6695__, new_new_n6696__, new_new_n6697__, new_new_n6698__,
    new_new_n6699__, new_new_n6700__, new_new_n6701__, new_new_n6702__,
    new_new_n6703__, new_new_n6704__, new_new_n6705__, new_new_n6706__,
    new_new_n6707__, new_new_n6708__, new_new_n6709__, new_new_n6710__,
    new_new_n6711__, new_new_n6712__, new_new_n6713__, new_new_n6714__,
    new_new_n6715__, new_new_n6716__, new_new_n6717__, new_new_n6718__,
    new_new_n6719__, new_new_n6720__, new_new_n6721__, new_new_n6722__,
    new_new_n6723__, new_new_n6724__, new_new_n6725__, new_new_n6726__,
    new_new_n6727__, new_new_n6728__, new_new_n6729__, new_new_n6730__,
    new_new_n6731__, new_new_n6732__, new_new_n6733__, new_new_n6734__,
    new_new_n6735__, new_new_n6736__, new_new_n6737__, new_new_n6738__,
    new_new_n6739__, new_new_n6740__, new_new_n6741__, new_new_n6742__,
    new_new_n6743__, new_new_n6744__, new_new_n6745__, new_new_n6746__,
    new_new_n6747__, new_new_n6748__, new_new_n6749__, new_new_n6750__,
    new_new_n6751__, new_new_n6752__, new_new_n6753__, new_new_n6754__,
    new_new_n6755__, new_new_n6756__, new_new_n6757__, new_new_n6758__,
    new_new_n6759__, new_new_n6760__, new_new_n6761__, new_new_n6762__,
    new_new_n6763__, new_new_n6764__, new_new_n6765__, new_new_n6766__,
    new_new_n6767__, new_new_n6768__, new_new_n6769__, new_new_n6770__,
    new_new_n6771__, new_new_n6772__, new_new_n6773__, new_new_n6774__,
    new_new_n6775__, new_new_n6776__, new_new_n6777__, new_new_n6778__,
    new_new_n6779__, new_new_n6780__, new_new_n6781__, new_new_n6782__,
    new_new_n6783__, new_new_n6784__, new_new_n6785__, new_new_n6786__,
    new_new_n6787__, new_new_n6788__, new_new_n6789__, new_new_n6790__,
    new_new_n6791__, new_new_n6792__, new_new_n6793__, new_new_n6794__,
    new_new_n6795__, new_new_n6796__, new_new_n6797__, new_new_n6798__,
    new_new_n6799__, new_new_n6800__, new_new_n6801__, new_new_n6802__,
    new_new_n6803__, new_new_n6804__, new_new_n6805__, new_new_n6806__,
    new_new_n6807__, new_new_n6808__, new_new_n6809__, new_new_n6810__,
    new_new_n6811__, new_new_n6812__, new_new_n6813__, new_new_n6814__,
    new_new_n6815__, new_new_n6816__, new_new_n6817__, new_new_n6818__,
    new_new_n6819__, new_new_n6820__, new_new_n6821__, new_new_n6822__,
    new_new_n6823__, new_new_n6824__, new_new_n6825__, new_new_n6826__,
    new_new_n6827__, new_new_n6828__, new_new_n6829__, new_new_n6830__,
    new_new_n6831__, new_new_n6832__, new_new_n6833__, new_new_n6834__,
    new_new_n6835__, new_new_n6836__, new_new_n6837__, new_new_n6838__,
    new_new_n6839__, new_new_n6840__, new_new_n6841__, new_new_n6842__,
    new_new_n6843__, new_new_n6844__, new_new_n6845__, new_new_n6846__,
    new_new_n6847__, new_new_n6848__, new_new_n6849__, new_new_n6850__,
    new_new_n6851__, new_new_n6852__, new_new_n6853__, new_new_n6854__,
    new_new_n6855__, new_new_n6856__, new_new_n6857__, new_new_n6858__,
    new_new_n6859__, new_new_n6860__, new_new_n6861__, new_new_n6862__,
    new_new_n6863__, new_new_n6864__, new_new_n6865__, new_new_n6866__,
    new_new_n6867__, new_new_n6868__, new_new_n6869__, new_new_n6870__,
    new_new_n6871__, new_new_n6872__, new_new_n6873__, new_new_n6874__,
    new_new_n6875__, new_new_n6876__, new_new_n6877__, new_new_n6878__,
    new_new_n6879__, new_new_n6880__, new_new_n6881__, new_new_n6882__,
    new_new_n6883__, new_new_n6884__, new_new_n6885__, new_new_n6886__,
    new_new_n6887__, new_new_n6888__, new_new_n6889__, new_new_n6890__,
    new_new_n6891__, new_new_n6892__, new_new_n6893__, new_new_n6894__,
    new_new_n6895__, new_new_n6896__, new_new_n6897__, new_new_n6898__,
    new_new_n6899__, new_new_n6900__, new_new_n6901__, new_new_n6902__,
    new_new_n6903__, new_new_n6904__, new_new_n6905__, new_new_n6906__,
    new_new_n6907__, new_new_n6908__, new_new_n6909__, new_new_n6910__,
    new_new_n6911__, new_new_n6912__, new_new_n6913__, new_new_n6914__,
    new_new_n6915__, new_new_n6916__, new_new_n6917__, new_new_n6918__,
    new_new_n6919__, new_new_n6920__, new_new_n6921__, new_new_n6922__,
    new_new_n6923__, new_new_n6924__, new_new_n6925__, new_new_n6926__,
    new_new_n6927__, new_new_n6928__, new_new_n6929__, new_new_n6930__,
    new_new_n6931__, new_new_n6932__, new_new_n6933__, new_new_n6934__,
    new_new_n6935__, new_new_n6936__, new_new_n6937__, new_new_n6938__,
    new_new_n6939__, new_new_n6940__, new_new_n6941__, new_new_n6942__,
    new_new_n6943__, new_new_n6944__, new_new_n6945__, new_new_n6946__,
    new_new_n6947__, new_new_n6948__, new_new_n6949__, new_new_n6950__,
    new_new_n6951__, new_new_n6952__, new_new_n6953__, new_new_n6954__,
    new_new_n6955__, new_new_n6956__, new_new_n6957__, new_new_n6958__,
    new_new_n6959__, new_new_n6960__, new_new_n6961__, new_new_n6962__,
    new_new_n6963__, new_new_n6964__, new_new_n6965__, new_new_n6966__,
    new_new_n6967__, new_new_n6968__, new_new_n6969__, new_new_n6970__,
    new_new_n6971__, new_new_n6972__, new_new_n6973__, new_new_n6974__,
    new_new_n6975__, new_new_n6976__, new_new_n6977__, new_new_n6978__,
    new_new_n6979__, new_new_n6980__, new_new_n6981__, new_new_n6982__,
    new_new_n6983__, new_new_n6984__, new_new_n6985__, new_new_n6986__,
    new_new_n6987__, new_new_n6988__, new_new_n6989__, new_new_n6990__,
    new_new_n6991__, new_new_n6992__, new_new_n6993__, new_new_n6994__,
    new_new_n6995__, new_new_n6996__, new_new_n6997__, new_new_n6998__,
    new_new_n6999__, new_new_n7000__, new_new_n7001__, new_new_n7002__,
    new_new_n7003__, new_new_n7004__, new_new_n7005__, new_new_n7006__,
    new_new_n7007__, new_new_n7008__, new_new_n7009__, new_new_n7010__,
    new_new_n7011__, new_new_n7012__, new_new_n7013__, new_new_n7014__,
    new_new_n7015__, new_new_n7016__, new_new_n7017__, new_new_n7018__,
    new_new_n7019__, new_new_n7020__, new_new_n7021__, new_new_n7022__,
    new_new_n7023__, new_new_n7024__, new_new_n7025__, new_new_n7026__,
    new_new_n7027__, new_new_n7028__, new_new_n7029__, new_new_n7030__,
    new_new_n7031__, new_new_n7032__, new_new_n7033__, new_new_n7034__,
    new_new_n7035__, new_new_n7036__, new_new_n7037__, new_new_n7038__,
    new_new_n7039__, new_new_n7040__, new_new_n7041__, new_new_n7042__,
    new_new_n7043__, new_new_n7044__, new_new_n7045__, new_new_n7046__,
    new_new_n7047__, new_new_n7048__, new_new_n7049__, new_new_n7050__,
    new_new_n7051__, new_new_n7052__, new_new_n7053__, new_new_n7054__,
    new_new_n7055__, new_new_n7056__, new_new_n7057__, new_new_n7058__,
    new_new_n7059__, new_new_n7060__, new_new_n7061__, new_new_n7062__,
    new_new_n7063__, new_new_n7064__, new_new_n7065__, new_new_n7066__,
    new_new_n7067__, new_new_n7068__, new_new_n7069__, new_new_n7070__,
    new_new_n7071__, new_new_n7072__, new_new_n7073__, new_new_n7074__,
    new_new_n7075__, new_new_n7076__, new_new_n7077__, new_new_n7078__,
    new_new_n7079__, new_new_n7080__, new_new_n7081__, new_new_n7082__,
    new_new_n7083__, new_new_n7084__, new_new_n7085__, new_new_n7086__,
    new_new_n7087__, new_new_n7088__, new_new_n7089__, new_new_n7090__,
    new_new_n7091__, new_new_n7092__, new_new_n7093__, new_new_n7094__,
    new_new_n7095__, new_new_n7096__, new_new_n7097__, new_new_n7098__,
    new_new_n7099__, new_new_n7100__, new_new_n7101__, new_new_n7102__,
    new_new_n7103__, new_new_n7104__, new_new_n7105__, new_new_n7106__,
    new_new_n7107__, new_new_n7108__, new_new_n7109__, new_new_n7110__,
    new_new_n7111__, new_new_n7112__, new_new_n7113__, new_new_n7114__,
    new_new_n7115__, new_new_n7116__, new_new_n7117__, new_new_n7118__,
    new_new_n7119__, new_new_n7120__, new_new_n7121__, new_new_n7122__,
    new_new_n7123__, new_new_n7124__, new_new_n7125__, new_new_n7126__,
    new_new_n7127__, new_new_n7128__, new_new_n7129__, new_new_n7130__,
    new_new_n7131__, new_new_n7132__, new_new_n7133__, new_new_n7134__,
    new_new_n7135__, new_new_n7136__, new_new_n7137__, new_new_n7138__,
    new_new_n7139__, new_new_n7140__, new_new_n7141__, new_new_n7142__,
    new_new_n7143__, new_new_n7144__, new_new_n7145__, new_new_n7146__,
    new_new_n7147__, new_new_n7148__, new_new_n7149__, new_new_n7150__,
    new_new_n7151__, new_new_n7152__, new_new_n7153__, new_new_n7154__,
    new_new_n7155__, new_new_n7156__, new_new_n7157__, new_new_n7158__,
    new_new_n7159__, new_new_n7160__, new_new_n7161__, new_new_n7162__,
    new_new_n7163__, new_new_n7164__, new_new_n7165__, new_new_n7166__,
    new_new_n7167__, new_new_n7168__, new_new_n7169__, new_new_n7170__,
    new_new_n7171__, new_new_n7172__, new_new_n7173__, new_new_n7174__,
    new_new_n7175__, new_new_n7176__, new_new_n7177__, new_new_n7178__,
    new_new_n7179__, new_new_n7180__, new_new_n7181__, new_new_n7182__,
    new_new_n7183__, new_new_n7184__, new_new_n7185__, new_new_n7186__,
    new_new_n7187__, new_new_n7188__, new_new_n7189__, new_new_n7190__,
    new_new_n7191__, new_new_n7192__, new_new_n7193__, new_new_n7194__,
    new_new_n7195__, new_new_n7196__, new_new_n7197__, new_new_n7198__,
    new_new_n7199__, new_new_n7200__, new_new_n7201__, new_new_n7202__,
    new_new_n7203__, new_new_n7204__, new_new_n7205__, new_new_n7206__,
    new_new_n7207__, new_new_n7208__, new_new_n7209__, new_new_n7210__,
    new_new_n7211__, new_new_n7212__, new_new_n7213__, new_new_n7214__,
    new_new_n7215__, new_new_n7216__, new_new_n7217__, new_new_n7218__,
    new_new_n7219__, new_new_n7220__, new_new_n7221__, new_new_n7222__,
    new_new_n7223__, new_new_n7224__, new_new_n7225__, new_new_n7226__,
    new_new_n7227__, new_new_n7228__, new_new_n7229__, new_new_n7230__,
    new_new_n7231__, new_new_n7232__, new_new_n7233__, new_new_n7234__,
    new_new_n7235__, new_new_n7236__, new_new_n7237__, new_new_n7238__,
    new_new_n7239__, new_new_n7240__, new_new_n7241__, new_new_n7242__,
    new_new_n7243__, new_new_n7244__, new_new_n7245__, new_new_n7246__,
    new_new_n7247__, new_new_n7248__, new_new_n7249__, new_new_n7250__,
    new_new_n7251__, new_new_n7252__, new_new_n7253__, new_new_n7254__,
    new_new_n7255__, new_new_n7256__, new_new_n7257__, new_new_n7258__,
    new_new_n7259__, new_new_n7260__, new_new_n7261__, new_new_n7262__,
    new_new_n7263__, new_new_n7264__, new_new_n7265__, new_new_n7266__,
    new_new_n7267__, new_new_n7268__, new_new_n7269__, new_new_n7270__,
    new_new_n7271__, new_new_n7272__, new_new_n7273__, new_new_n7274__,
    new_new_n7275__, new_new_n7276__, new_new_n7277__, new_new_n7278__,
    new_new_n7279__, new_new_n7280__, new_new_n7281__, new_new_n7282__,
    new_new_n7283__, new_new_n7284__, new_new_n7285__, new_new_n7286__,
    new_new_n7287__, new_new_n7288__, new_new_n7289__, new_new_n7290__,
    new_new_n7291__, new_new_n7292__, new_new_n7293__, new_new_n7294__,
    new_new_n7295__, new_new_n7296__, new_new_n7297__, new_new_n7298__,
    new_new_n7299__, new_new_n7300__, new_new_n7301__, new_new_n7302__,
    new_new_n7303__, new_new_n7304__, new_new_n7305__, new_new_n7306__,
    new_new_n8443__, new_new_n8444__, new_new_n8445__, new_new_n8446__,
    new_new_n8447__, new_new_n8448__, new_new_n8449__, new_new_n8450__,
    new_new_n8451__, new_new_n8452__, new_new_n8453__, new_new_n8454__,
    new_new_n8455__, new_new_n8456__, new_new_n8457__, new_new_n8458__,
    new_new_n8459__, new_new_n8460__, new_new_n8461__, new_new_n8462__,
    new_new_n8463__, new_new_n8464__, new_new_n8465__, new_new_n8466__,
    new_new_n8467__, new_new_n8468__, new_new_n8469__, new_new_n8470__,
    new_new_n8471__, new_new_n8472__, new_new_n8473__, new_new_n8474__,
    new_new_n8475__, new_new_n8476__, new_new_n8477__, new_new_n8478__,
    new_new_n8479__, new_new_n8480__, new_new_n8481__, new_new_n8482__,
    new_new_n8483__, new_new_n8484__, new_new_n8485__, new_new_n8486__,
    new_new_n8487__, new_new_n8488__, new_new_n8489__, new_new_n8490__,
    new_new_n8491__, new_new_n8492__, new_new_n8493__, new_new_n8494__,
    new_new_n8495__, new_new_n8496__, new_new_n8497__, new_new_n8498__,
    new_new_n8499__, new_new_n8500__, new_new_n8501__, new_new_n8502__,
    new_new_n8503__, new_new_n8504__, new_new_n8505__, new_new_n8506__,
    new_new_n8507__, new_new_n8508__, new_new_n8509__, new_new_n8510__,
    new_new_n8511__, new_new_n8512__, new_new_n8513__, new_new_n8514__,
    new_new_n8515__, new_new_n8516__, new_new_n8517__, new_new_n8518__,
    new_new_n8519__, new_new_n8520__, new_new_n8521__, new_new_n8522__,
    new_new_n8523__, new_new_n8524__, new_new_n8525__, new_new_n8526__,
    new_new_n8527__, new_new_n8528__, new_new_n8529__, new_new_n8530__,
    new_new_n8531__, new_new_n8532__, new_new_n8533__, new_new_n8534__,
    new_new_n8535__, new_new_n8536__, new_new_n8537__, new_new_n8538__,
    new_new_n8539__, new_new_n8540__, new_new_n8541__, new_new_n8542__,
    new_new_n8543__, new_new_n8544__, new_new_n8545__, new_new_n8546__,
    new_new_n8547__, new_new_n8548__, new_new_n8549__, new_new_n8550__,
    new_new_n8551__, new_new_n8552__, new_new_n8553__, new_new_n8554__,
    new_new_n8555__, new_new_n8556__, new_new_n8557__, new_new_n8558__,
    new_new_n8559__, new_new_n8560__, new_new_n8561__, new_new_n8562__,
    new_new_n8563__, new_new_n8564__, new_new_n8565__, new_new_n8566__,
    new_new_n8567__, new_new_n8568__, new_new_n8569__, new_new_n8570__,
    new_new_n8571__, new_new_n8572__, new_new_n8573__, new_new_n8574__,
    new_new_n8575__, new_new_n8576__, new_new_n8577__, new_new_n8578__,
    new_new_n8579__, new_new_n8580__, new_new_n8581__, new_new_n8582__,
    new_new_n8583__, new_new_n8584__, new_new_n8585__, new_new_n8586__,
    new_new_n8587__, new_new_n8588__, new_new_n8589__, new_new_n8590__,
    new_new_n8591__, new_new_n8592__, new_new_n8593__, new_new_n8594__,
    new_new_n8595__, new_new_n8596__, new_new_n8597__, new_new_n8598__,
    new_new_n8599__, new_new_n8600__, new_new_n8601__, new_new_n8602__,
    new_new_n8603__, new_new_n8604__, new_new_n8605__, new_new_n8606__,
    new_new_n8607__, new_new_n8608__, new_new_n8609__, new_new_n8610__,
    new_new_n8611__, new_new_n8612__, new_new_n8613__, new_new_n8614__,
    new_new_n8615__, new_new_n8616__, new_new_n8617__, new_new_n8618__,
    new_new_n8619__, new_new_n8620__, new_new_n8621__, new_new_n8622__,
    new_new_n8623__, new_new_n8624__, new_new_n8625__, new_new_n8626__,
    new_new_n8627__, new_new_n8628__, new_new_n8629__, new_new_n8630__,
    new_new_n8631__, new_new_n8632__, new_new_n8633__, new_new_n8634__,
    new_new_n8635__, new_new_n8636__, new_new_n8637__, new_new_n8638__,
    new_new_n8639__, new_new_n8640__, new_new_n8641__, new_new_n8642__,
    new_new_n8643__, new_new_n8644__, new_new_n8645__, new_new_n8646__,
    new_new_n8647__, new_new_n8648__, new_new_n8649__, new_new_n8650__,
    new_new_n8651__, new_new_n8652__, new_new_n8653__, new_new_n8654__,
    new_new_n8655__, new_new_n8656__, new_new_n8657__, new_new_n8658__,
    new_new_n8659__, new_new_n8660__, new_new_n8661__, new_new_n8662__,
    new_new_n8663__, new_new_n8664__, new_new_n8665__, new_new_n8666__,
    new_new_n8667__, new_new_n8668__, new_new_n8669__, new_new_n8670__,
    new_new_n8671__, new_new_n8672__, new_new_n8673__, new_new_n8674__,
    new_new_n8675__, new_new_n8676__, new_new_n8677__, new_new_n8678__,
    new_new_n8679__, new_new_n8680__, new_new_n8681__, new_new_n8682__,
    new_new_n8683__, new_new_n8684__, new_new_n8685__, new_new_n8686__,
    new_new_n8687__, new_new_n8688__, new_new_n8689__, new_new_n8690__,
    new_new_n8691__, new_new_n8692__, new_new_n8693__, new_new_n8694__,
    new_new_n8695__, new_new_n8696__, new_new_n8697__, new_new_n8698__,
    new_new_n8699__, new_new_n8700__, new_new_n8701__, new_new_n8702__,
    new_new_n8703__, new_new_n8704__, new_new_n8705__, new_new_n8706__,
    new_new_n8707__, new_new_n8708__, new_new_n8709__, new_new_n8710__,
    new_new_n8711__, new_new_n8712__, new_new_n8713__, new_new_n8714__,
    new_new_n8715__, new_new_n8716__, new_new_n8717__, new_new_n8718__,
    new_new_n8719__, new_new_n8720__, new_new_n8721__, new_new_n8722__,
    new_new_n8723__, new_new_n8724__, new_new_n8725__, new_new_n8726__,
    new_new_n8727__, new_new_n8728__, new_new_n8729__, new_new_n8730__,
    new_new_n8731__, new_new_n8732__, new_new_n8733__, new_new_n8734__,
    new_new_n8735__, new_new_n8736__, new_new_n8737__, new_new_n8738__,
    new_new_n8739__, new_new_n8740__, new_new_n8741__, new_new_n8742__,
    new_new_n8743__, new_new_n8744__, new_new_n8745__, new_new_n8746__,
    new_new_n8747__, new_new_n8748__, new_new_n8749__, new_new_n8750__,
    new_new_n8751__, new_new_n8752__, new_new_n8753__, new_new_n8754__,
    new_new_n8755__, new_new_n8756__, new_new_n8757__, new_new_n8758__,
    new_new_n8759__, new_new_n8760__, new_new_n8761__, new_new_n8762__,
    new_new_n8763__, new_new_n8764__, new_new_n8765__, new_new_n8766__,
    new_new_n8767__, new_new_n8768__, new_new_n8769__, new_new_n8770__,
    new_new_n8771__, new_new_n8772__, new_new_n8773__, new_new_n8774__,
    new_new_n8775__, new_new_n8776__, new_new_n8777__, new_new_n8778__,
    new_new_n8779__, new_new_n8780__, new_new_n8781__, new_new_n8782__,
    new_new_n8783__, new_new_n8784__, new_new_n8785__, new_new_n8786__,
    new_new_n8787__, new_new_n8788__, new_new_n8789__, new_new_n8790__,
    new_new_n8791__, new_new_n8792__, new_new_n8793__, new_new_n8794__,
    new_new_n8795__, new_new_n8796__, new_new_n8797__, new_new_n8798__,
    new_new_n8799__, new_new_n8800__, new_new_n8801__, new_new_n8802__,
    new_new_n8803__, new_new_n8804__, new_new_n8805__, new_new_n8806__,
    new_new_n8807__, new_new_n8808__, new_new_n8809__, new_new_n8810__,
    new_new_n8811__, new_new_n8812__, new_new_n8813__, new_new_n8814__,
    new_new_n8815__, new_new_n8816__, new_new_n8817__, new_new_n8818__,
    new_new_n8819__, new_new_n8820__, new_new_n8821__, new_new_n8822__,
    new_new_n8823__, new_new_n8824__, new_new_n8825__, new_new_n8826__,
    new_new_n8827__, new_new_n8828__, new_new_n8829__, new_new_n8830__,
    new_new_n8831__, new_new_n8832__, new_new_n8833__, new_new_n8834__,
    new_new_n8835__, new_new_n8836__, new_new_n8837__, new_new_n8838__,
    new_new_n8839__, new_new_n8840__, new_new_n8841__, new_new_n8842__,
    new_new_n8843__, new_new_n8844__, new_new_n8845__, new_new_n8846__,
    new_new_n8847__, new_new_n8848__, new_new_n8849__, new_new_n8850__,
    new_new_n8851__, new_new_n8852__, new_new_n8853__, new_new_n8854__,
    new_new_n8855__, new_new_n8856__, new_new_n8857__, new_new_n8858__,
    new_new_n8859__, new_new_n8860__, new_new_n8861__, new_new_n8862__,
    new_new_n8863__, new_new_n8864__, new_new_n8865__, new_new_n8866__,
    new_new_n8867__, new_new_n8868__, new_new_n8869__, new_new_n8870__,
    new_new_n8871__, new_new_n8872__, new_new_n8873__, new_new_n8874__,
    new_new_n8875__, new_new_n8876__, new_new_n8877__, new_new_n8878__,
    new_new_n8879__, new_new_n8880__, new_new_n8881__, new_new_n8882__,
    new_new_n8883__, new_new_n8884__, new_new_n8885__, new_new_n8886__,
    new_new_n8887__, new_new_n8888__, new_new_n8889__, new_new_n8890__,
    new_new_n8891__, new_new_n8892__, new_new_n8893__, new_new_n8894__,
    new_new_n8895__, new_new_n8896__, new_new_n8897__, new_new_n8898__,
    new_new_n8899__, new_new_n8900__, new_new_n8901__, new_new_n8902__,
    new_new_n8903__, new_new_n8904__, new_new_n8905__, new_new_n8906__,
    new_new_n8907__, new_new_n8908__, new_new_n8909__, new_new_n8910__,
    new_new_n8911__, new_new_n8912__, new_new_n8913__, new_new_n8914__,
    new_new_n8915__, new_new_n8916__, new_new_n8917__, new_new_n8918__,
    new_new_n8919__, new_new_n8920__, new_new_n8921__, new_new_n8922__,
    new_new_n8923__, new_new_n8924__, new_new_n8925__, new_new_n8926__,
    new_new_n8927__, new_new_n8928__, new_new_n8929__, new_new_n8930__,
    new_new_n8931__, new_new_n8932__, new_new_n8933__, new_new_n8934__,
    new_new_n8935__, new_new_n8936__, new_new_n8937__, new_new_n8938__,
    new_new_n8939__, new_new_n8940__, new_new_n8941__, new_new_n8942__,
    new_new_n8943__, new_new_n8944__, new_new_n8945__, new_new_n8946__,
    new_new_n8947__, new_new_n8948__, new_new_n8949__, new_new_n8950__,
    new_new_n8951__, new_new_n8952__, new_new_n8953__, new_new_n8954__,
    new_new_n8955__, new_new_n8956__, new_new_n8957__, new_new_n8958__,
    new_new_n8959__, new_new_n8960__, new_new_n8961__, new_new_n8962__,
    new_new_n8963__, new_new_n8964__, new_new_n8965__, new_new_n8966__,
    new_new_n8967__, new_new_n8968__, new_new_n8969__, new_new_n8970__,
    new_new_n8971__, new_new_n8972__, new_new_n8973__, new_new_n8974__,
    new_new_n8975__, new_new_n8976__, new_new_n8977__, new_new_n8978__,
    new_new_n8979__, new_new_n8980__, new_new_n8981__, new_new_n8982__,
    new_new_n8983__, new_new_n8984__, new_new_n8985__, new_new_n8986__,
    new_new_n8987__, new_new_n8988__, new_new_n8989__, new_new_n8990__,
    new_new_n8991__, new_new_n8992__, new_new_n8993__, new_new_n8994__,
    new_new_n8995__, new_new_n8996__, new_new_n8997__, new_new_n8998__,
    new_new_n8999__, new_new_n9000__, new_new_n9001__, new_new_n9002__,
    new_new_n9003__, new_new_n9004__, new_new_n9005__, new_new_n9006__,
    new_new_n9007__, new_new_n9008__, new_new_n9009__, new_new_n9010__,
    new_new_n9011__, new_new_n9012__, new_new_n9013__, new_new_n9014__,
    new_new_n9015__, new_new_n9016__, new_new_n9017__, new_new_n9018__,
    new_new_n9019__, new_new_n9020__, new_new_n9021__, new_new_n9022__,
    new_new_n9023__, new_new_n9024__, new_new_n9025__, new_new_n9026__,
    new_new_n9027__, new_new_n9028__, new_new_n9029__, new_new_n9030__,
    new_new_n9031__, new_new_n9032__, new_new_n9033__, new_new_n9034__,
    new_new_n9035__, new_new_n9036__, new_new_n9037__, new_new_n9038__,
    new_new_n9039__, new_new_n9040__, new_new_n9041__, new_new_n9042__,
    new_new_n9043__, new_new_n9044__, new_new_n9045__, new_new_n9046__,
    new_new_n9047__, new_new_n9048__, new_new_n9049__, new_new_n9050__,
    new_new_n9051__, new_new_n9052__, new_new_n9053__, new_new_n9054__,
    new_new_n9055__, new_new_n9056__, new_new_n9057__, new_new_n9058__,
    new_new_n9059__, new_new_n9060__, new_new_n9061__, new_new_n9062__,
    new_new_n9063__, new_new_n9064__, new_new_n9065__, new_new_n9066__,
    new_new_n9067__, new_new_n9068__, new_new_n9069__, new_new_n9070__,
    new_new_n9071__, new_new_n9072__, new_new_n9073__, new_new_n9074__,
    new_new_n9075__, new_new_n9076__, new_new_n9077__, new_new_n9078__,
    new_new_n9079__, new_new_n9080__, new_new_n9081__, new_new_n9082__,
    new_new_n9083__, new_new_n9084__, new_new_n9085__, new_new_n9086__,
    new_new_n9087__, new_new_n9088__, new_new_n9089__, new_new_n9090__,
    new_new_n9091__, new_new_n9092__, new_new_n9093__, new_new_n9094__,
    new_new_n9095__, new_new_n9096__, new_new_n9097__, new_new_n9098__,
    new_new_n9099__, new_new_n9100__, new_new_n9101__, new_new_n9102__,
    new_new_n9103__, new_new_n9104__, new_new_n9105__, new_new_n9106__,
    new_new_n9107__, new_new_n9108__, new_new_n9109__, new_new_n9110__,
    new_new_n9111__, new_new_n9112__, new_new_n9113__, new_new_n9114__,
    new_new_n9115__, new_new_n9116__, new_new_n9117__, new_new_n9118__,
    new_new_n9119__, new_new_n9120__, new_new_n9121__, new_new_n9122__,
    new_new_n9123__, new_new_n9124__, new_new_n9125__, new_new_n9126__,
    new_new_n9127__, new_new_n9128__, new_new_n9129__, new_new_n9130__,
    new_new_n9131__, new_new_n9132__, new_new_n9133__, new_new_n9134__,
    new_new_n9135__, new_new_n9136__, new_new_n9137__, new_new_n9138__,
    new_new_n9139__, new_new_n9140__, new_new_n9141__, new_new_n9142__,
    new_new_n9143__, new_new_n9144__, new_new_n9145__, new_new_n9146__,
    new_new_n9147__, new_new_n9148__, new_new_n9149__, new_new_n9150__,
    new_new_n9151__, new_new_n9152__, new_new_n9153__, new_new_n9154__,
    new_new_n9155__, new_new_n9156__, new_new_n9157__, new_new_n9158__,
    new_new_n9159__, new_new_n9160__, new_new_n9161__, new_new_n9162__,
    new_new_n9163__, new_new_n9164__, new_new_n9165__, new_new_n9166__,
    new_new_n9167__, new_new_n9168__, new_new_n9169__, new_new_n9170__,
    new_new_n9171__, new_new_n9172__, new_new_n9173__, new_new_n9174__,
    new_new_n9175__, new_new_n9176__, new_new_n9177__, new_new_n9178__,
    new_new_n9179__, new_new_n9180__, new_new_n9181__, new_new_n9182__,
    new_new_n9183__, new_new_n9184__, new_new_n9185__, new_new_n9186__,
    new_new_n9187__, new_new_n9188__, new_new_n9189__, new_new_n9190__,
    new_new_n9191__, new_new_n9192__, new_new_n9193__, new_new_n9194__,
    new_new_n9195__, new_new_n9196__, new_new_n9197__, new_new_n9198__,
    new_new_n9199__, new_new_n9200__, new_new_n9201__, new_new_n9202__,
    new_new_n9203__, new_new_n9204__, new_new_n9205__, new_new_n9206__,
    new_new_n9207__, new_new_n9208__, new_new_n9209__, new_new_n9210__,
    new_new_n9211__, new_new_n9212__, new_new_n9213__, new_new_n9214__,
    new_new_n9215__, new_new_n9216__, new_new_n9217__, new_new_n9218__,
    new_new_n9219__, new_new_n9220__, new_new_n9221__, new_new_n9222__,
    new_new_n9223__, new_new_n9224__, new_new_n9225__, new_new_n9226__,
    new_new_n9227__, new_new_n9228__, new_new_n9229__, new_new_n9230__,
    new_new_n9231__, new_new_n9232__, new_new_n9233__, new_new_n9234__,
    new_new_n9235__, new_new_n9236__, new_new_n9237__, new_new_n9238__,
    new_new_n9239__, new_new_n9240__, new_new_n9241__, new_new_n9242__,
    new_new_n9243__, new_new_n9244__, new_new_n9245__, new_new_n9246__,
    new_new_n9247__, new_new_n9248__, new_new_n9249__, new_new_n9250__,
    new_new_n9251__, new_new_n9252__, new_new_n9253__, new_new_n9254__,
    new_new_n9255__, new_new_n9256__, new_new_n9257__, new_new_n9258__,
    new_new_n9259__, new_new_n9260__, new_new_n9261__, new_new_n9262__,
    new_new_n9263__, new_new_n9264__, new_new_n9265__, new_new_n9266__,
    new_new_n9267__, new_new_n9268__, new_new_n9269__, new_new_n9270__,
    new_new_n9271__, new_new_n9272__, new_new_n9273__, new_new_n9274__,
    new_new_n9275__, new_new_n9276__, new_new_n9277__, new_new_n9278__,
    new_new_n9279__, new_new_n9280__, new_new_n9281__, new_new_n9282__,
    new_new_n9283__, new_new_n9284__, new_new_n9285__, new_new_n9286__,
    new_new_n9287__, new_new_n9288__, new_new_n9289__, new_new_n9290__,
    new_new_n9291__, new_new_n9292__, new_new_n9293__, new_new_n9294__,
    new_new_n9295__, new_new_n9296__, new_new_n9297__, new_new_n9298__,
    new_new_n9299__, new_new_n9300__, new_new_n9301__, new_new_n9302__,
    new_new_n9303__, new_new_n9304__, new_new_n9305__, new_new_n9306__,
    new_new_n9307__, new_new_n9308__, new_new_n9309__, new_new_n9310__,
    new_new_n9311__, new_new_n9312__, new_new_n9313__, new_new_n9314__,
    new_new_n9315__, new_new_n9316__, new_new_n9317__, new_new_n9318__,
    new_new_n9319__, new_new_n9320__, new_new_n9321__, new_new_n9322__,
    new_new_n9323__, new_new_n9324__, new_new_n9325__, new_new_n9326__,
    new_new_n9327__, new_new_n9328__, new_new_n9329__, new_new_n9330__,
    new_new_n9331__, new_new_n9332__, new_new_n9333__, new_new_n9334__,
    new_new_n9335__, new_new_n9336__, new_new_n9337__, new_new_n9338__,
    new_new_n9339__, new_new_n9340__, new_new_n9341__, new_new_n9342__,
    new_new_n9343__, new_new_n9344__, new_new_n9345__, new_new_n9346__,
    new_new_n9347__, new_new_n9348__, new_new_n9349__, new_new_n9350__,
    new_new_n9351__, new_new_n9352__, new_new_n9353__, new_new_n9354__,
    new_new_n9355__, new_new_n9356__, new_new_n9357__, new_new_n9358__,
    new_new_n9359__, new_new_n9360__, new_new_n9361__, new_new_n9362__,
    new_new_n9363__, new_new_n9364__, new_new_n9365__, new_new_n9366__,
    new_new_n9367__, new_new_n9368__, new_new_n9369__, new_new_n9370__,
    new_new_n9371__, new_new_n9372__, new_new_n9373__, new_new_n9374__,
    new_new_n9375__, new_new_n9376__, new_new_n9377__, new_new_n9378__,
    new_new_n9379__, new_new_n9380__, new_new_n9381__, new_new_n9382__,
    new_new_n9383__, new_new_n9384__, new_new_n9385__, new_new_n9386__,
    new_new_n9387__, new_new_n9388__, new_new_n9389__, new_new_n9390__,
    new_new_n9391__, new_new_n9392__, new_new_n9393__, new_new_n9394__,
    new_new_n9395__, new_new_n9396__, new_new_n9397__, new_new_n9398__,
    new_new_n9399__, new_new_n9400__, new_new_n9401__, new_new_n9402__,
    new_new_n9403__, new_new_n9404__, new_new_n9405__, new_new_n9406__,
    new_new_n9407__, new_new_n9408__, new_new_n9409__, new_new_n9410__,
    new_new_n9411__, new_new_n9412__, new_new_n9413__, new_new_n9414__,
    new_new_n9415__, new_new_n9416__, new_new_n9417__, new_new_n9418__,
    new_new_n9419__, new_new_n9420__, new_new_n9421__, new_new_n9422__,
    new_new_n9423__, new_new_n9424__, new_new_n9425__, new_new_n9426__,
    new_new_n9427__, new_new_n9428__, new_new_n9429__, new_new_n9430__,
    new_new_n9431__, new_new_n9432__, new_new_n9433__, new_new_n9434__,
    new_new_n9435__, new_new_n9436__, new_new_n9437__, new_new_n9438__,
    new_new_n9439__, new_new_n9440__, new_new_n9441__, new_new_n9442__,
    new_new_n9443__, new_new_n9444__, new_new_n9445__, new_new_n9446__,
    new_new_n9447__, new_new_n9448__, new_new_n9449__, new_new_n9450__,
    new_new_n9451__, new_new_n9452__, new_new_n9453__, new_new_n9454__,
    new_new_n9455__, new_new_n9456__, new_new_n9457__, new_new_n9458__,
    new_new_n9459__, new_new_n9460__, new_new_n9461__, new_new_n9462__,
    new_new_n9463__, new_new_n9464__, new_new_n9465__, new_new_n9466__,
    new_new_n9467__, new_new_n9468__, new_new_n9469__, new_new_n9470__,
    new_new_n9471__, new_new_n9472__, new_new_n9473__, new_new_n9474__,
    new_new_n9475__, new_new_n9476__, new_new_n9477__, new_new_n9478__,
    new_new_n9479__, new_new_n9480__, new_new_n9481__, new_new_n9482__,
    new_new_n9483__, new_new_n9484__, new_new_n9485__, new_new_n9486__,
    new_new_n9487__, new_new_n9488__, new_new_n9489__, new_new_n9490__,
    new_new_n9491__, new_new_n9492__, new_new_n9493__, new_new_n9494__,
    new_new_n9495__, new_new_n9496__, new_new_n9497__, new_new_n9498__,
    new_new_n9499__, new_new_n9500__, new_new_n9501__, new_new_n9502__,
    new_new_n9503__, new_new_n9504__, new_new_n9505__, new_new_n9506__,
    new_new_n9507__, new_new_n9508__, new_new_n9509__, new_new_n9510__,
    new_new_n9511__, new_new_n9512__, new_new_n9513__, new_new_n9514__,
    new_new_n9515__, new_new_n9516__, new_new_n9517__, new_new_n9518__,
    new_new_n9519__, new_new_n9520__, new_new_n9521__, new_new_n9522__,
    new_new_n9523__, new_new_n9524__, new_new_n9525__, new_new_n9526__,
    new_new_n9527__, new_new_n9528__, new_new_n9529__, new_new_n9530__,
    new_new_n9531__, new_new_n9532__, new_new_n9533__, new_new_n9534__,
    new_new_n9535__, new_new_n9536__, new_new_n9537__, new_new_n9538__,
    new_new_n9539__, new_new_n9540__, new_new_n9541__, new_new_n9542__,
    new_new_n9543__, new_new_n9544__, new_new_n9545__, new_new_n9546__,
    new_new_n9547__, new_new_n9548__, new_new_n9549__, new_new_n9550__,
    new_new_n9551__, new_new_n9552__, new_new_n9553__, new_new_n9554__,
    new_new_n9555__, new_new_n9556__, new_new_n9557__, new_new_n9558__,
    new_new_n9559__, new_new_n9560__, new_new_n9561__, new_new_n9562__,
    new_new_n9563__, new_new_n9564__, new_new_n9565__, new_new_n9566__,
    new_new_n9567__, new_new_n9568__, new_new_n9569__, new_new_n9570__,
    new_new_n9571__, new_new_n9572__, new_new_n9573__, new_new_n9574__,
    new_new_n9575__, new_new_n9576__, new_new_n9577__, new_new_n9578__,
    new_new_n9579__, new_new_n9580__, new_new_n9581__, new_new_n9582__,
    new_new_n9583__, new_new_n9584__, new_new_n9585__, new_new_n9586__,
    new_new_n9587__, new_new_n9588__, new_new_n9589__, new_new_n9590__,
    new_new_n9591__, new_new_n9592__, new_new_n9593__, new_new_n9594__,
    new_new_n9595__, new_new_n9596__, new_new_n9597__, new_new_n9598__,
    new_new_n9599__, new_new_n9600__, new_new_n9601__, new_new_n9602__,
    new_new_n9603__, new_new_n9604__, new_new_n9605__, new_new_n9606__,
    new_new_n9607__, new_new_n9608__, new_new_n9609__, new_new_n9610__,
    new_new_n9611__, new_new_n9612__, new_new_n9613__, new_new_n9614__,
    new_new_n9615__, new_new_n9616__, new_new_n9617__, new_new_n9618__,
    new_new_n9619__, new_new_n9620__, new_new_n9621__, new_new_n9622__,
    new_new_n9623__, new_new_n9624__, new_new_n9625__, new_new_n9626__,
    new_new_n9627__, new_new_n9628__, new_new_n9629__, new_new_n9630__,
    new_new_n9631__, new_new_n9632__, new_new_n9633__, new_new_n9634__,
    new_new_n9635__, new_new_n9636__, new_new_n9637__, new_new_n9638__,
    new_new_n9639__, new_new_n9640__, new_new_n9641__, new_new_n9642__,
    new_new_n9643__, new_new_n9644__, new_new_n9645__, new_new_n9646__,
    new_new_n9647__, new_new_n9648__, new_new_n9649__, new_new_n9650__,
    new_new_n9651__, new_new_n9652__, new_new_n9653__, new_new_n9654__,
    new_new_n9655__, new_new_n9656__, new_new_n9657__, new_new_n9658__,
    new_new_n9659__, new_new_n9660__, new_new_n9661__, new_new_n9662__,
    new_new_n9663__, new_new_n9664__, new_new_n9665__, new_new_n9666__,
    new_new_n9667__, new_new_n9668__, new_new_n9669__, new_new_n9670__,
    new_new_n9671__, new_new_n9672__, new_new_n9673__, new_new_n9674__,
    new_new_n9675__, new_new_n9676__, new_new_n9677__, new_new_n9678__,
    new_new_n9679__, new_new_n9680__, new_new_n9681__, new_new_n9682__,
    new_new_n9683__, new_new_n9684__, new_new_n9685__, new_new_n9686__,
    new_new_n9687__, new_new_n9688__, new_new_n9689__, new_new_n9690__,
    new_new_n9691__, new_new_n9692__, new_new_n9693__, new_new_n9694__,
    new_new_n9695__, new_new_n9696__, new_new_n9697__, new_new_n9698__,
    new_new_n9699__, new_new_n9700__, new_new_n9701__, new_new_n9702__,
    new_new_n9703__, new_new_n9704__, new_new_n9705__, new_new_n9706__,
    new_new_n9707__, new_new_n9708__, new_new_n9709__, new_new_n9710__,
    new_new_n9711__, new_new_n9712__, new_new_n9713__, new_new_n9714__,
    new_new_n9715__, new_new_n9716__, new_new_n9717__, new_new_n9718__,
    new_new_n9719__, new_new_n9720__, new_new_n9721__, new_new_n9722__,
    new_new_n9723__, new_new_n9724__, new_new_n9725__, new_new_n9726__,
    new_new_n9727__, new_new_n9728__, new_new_n9729__, new_new_n9730__,
    new_new_n9731__, new_new_n9732__, new_new_n9733__, new_new_n9734__,
    new_new_n9735__, new_new_n9736__, new_new_n9737__, new_new_n9738__,
    new_new_n9739__, new_new_n9740__, new_new_n9741__, new_new_n9742__,
    new_new_n9743__, new_new_n9744__, new_new_n9745__, new_new_n9746__,
    new_new_n9747__, new_new_n9748__, new_new_n9749__, new_new_n9750__,
    new_new_n9751__, new_new_n9752__, new_new_n9753__, new_new_n9754__,
    new_new_n9755__, new_new_n9756__, new_new_n9757__, new_new_n9758__,
    new_new_n9759__, new_new_n9760__, new_new_n9761__, new_new_n9762__,
    new_new_n9763__, new_new_n9764__, new_new_n9765__, new_new_n9766__,
    new_new_n9767__, new_new_n9768__, new_new_n9769__, new_new_n9770__,
    new_new_n9771__, new_new_n9772__, new_new_n9773__, new_new_n9774__,
    new_new_n9775__, new_new_n9776__, new_new_n9777__, new_new_n9778__,
    new_new_n9779__, new_new_n9780__, new_new_n9781__, new_new_n9782__,
    new_new_n9783__, new_new_n9784__, new_new_n9785__, new_new_n9786__,
    new_new_n9787__, new_new_n9788__, new_new_n9789__, new_new_n9790__,
    new_new_n9791__, new_new_n9792__, new_new_n9793__, new_new_n9794__,
    new_new_n9795__, new_new_n9796__, new_new_n9797__, new_new_n9798__,
    new_new_n9799__, new_new_n9800__, new_new_n9801__, new_new_n9802__,
    new_new_n9803__, new_new_n9804__, new_new_n9805__, new_new_n9806__,
    new_new_n9807__, new_new_n9808__, new_new_n9809__, new_new_n9810__,
    new_new_n9811__, new_new_n9812__, new_new_n9813__, new_new_n9814__,
    new_new_n9815__, new_new_n9816__, new_new_n9817__, new_new_n9818__,
    new_new_n9819__, new_new_n9820__, new_new_n9821__, new_new_n9822__,
    new_new_n9823__, new_new_n9824__, new_new_n9825__, new_new_n9826__,
    new_new_n9827__, new_new_n9828__, new_new_n9829__, new_new_n9830__,
    new_new_n9831__, new_new_n9832__, new_new_n9833__, new_new_n9834__,
    new_new_n9835__, new_new_n9836__, new_new_n9837__, new_new_n9838__,
    new_new_n9839__, new_new_n9840__, new_new_n9841__, new_new_n9842__,
    new_new_n9843__, new_new_n9844__, new_new_n9845__, new_new_n9846__,
    new_new_n9847__, new_new_n9848__, new_new_n9849__, new_new_n9850__,
    new_new_n9851__, new_new_n9852__, new_new_n9853__, new_new_n9854__,
    new_new_n9855__, new_new_n9856__, new_new_n9857__, new_new_n9858__,
    new_new_n9859__, new_new_n9860__, new_new_n9861__, new_new_n9862__,
    new_new_n9863__, new_new_n9864__, new_new_n9865__, new_new_n9866__,
    new_new_n9867__, new_new_n9868__, new_new_n9869__, new_new_n9870__,
    new_new_n9871__, new_new_n9872__, new_new_n9873__, new_new_n9874__,
    new_new_n9875__, new_new_n9876__, new_new_n9877__, new_new_n9878__,
    new_new_n9879__, new_new_n9880__, new_new_n9881__, new_new_n9882__,
    new_new_n9883__, new_new_n9884__, new_new_n9885__, new_new_n9886__,
    new_new_n9887__, new_new_n9888__, new_new_n9889__, new_new_n9890__,
    new_new_n9891__, new_new_n9892__, new_new_n9893__, new_new_n9894__,
    new_new_n9895__, new_new_n9896__, new_new_n9897__, new_new_n9898__,
    new_new_n9899__, new_new_n9900__, new_new_n9901__, new_new_n9902__,
    new_new_n9903__, new_new_n9904__, new_new_n9905__, new_new_n9906__,
    new_new_n9907__, new_new_n9908__, new_new_n9909__, new_new_n9910__,
    new_new_n9911__, new_new_n9912__, new_new_n9913__, new_new_n9914__,
    new_new_n9915__, new_new_n9916__, new_new_n9917__, new_new_n9918__,
    new_new_n9919__, new_new_n9920__, new_new_n9921__, new_new_n9922__,
    new_new_n9923__, new_new_n9924__, new_new_n9925__, new_new_n9926__,
    new_new_n9927__, new_new_n9928__, new_new_n9929__, new_new_n9930__,
    new_new_n9931__, new_new_n9932__, new_new_n9933__, new_new_n9934__,
    new_new_n9935__, new_new_n9936__, new_new_n9937__, new_new_n9938__,
    new_new_n9939__, new_new_n9940__, new_new_n9941__, new_new_n9942__,
    new_new_n9943__, new_new_n9944__, new_new_n9945__, new_new_n9946__,
    new_new_n9947__, new_new_n9948__, new_new_n9949__, new_new_n9950__,
    new_new_n9951__, new_new_n9952__, new_new_n9953__, new_new_n9954__,
    new_new_n9955__, new_new_n9956__, new_new_n9957__, new_new_n9958__,
    new_new_n9959__, new_new_n9960__, new_new_n9961__, new_new_n9962__,
    new_new_n9963__, new_new_n9964__, new_new_n9965__, new_new_n9966__,
    new_new_n9967__, new_new_n9968__, new_new_n9969__, new_new_n9970__,
    new_new_n9971__, new_new_n9972__, new_new_n9973__, new_new_n9974__,
    new_new_n9975__, new_new_n9976__, new_new_n9977__, new_new_n9978__,
    new_new_n9979__, new_new_n9980__, new_new_n9981__, new_new_n9982__,
    new_new_n9983__, new_new_n9984__, new_new_n9985__, new_new_n9986__,
    new_new_n9987__, new_new_n9988__, new_new_n9989__, new_new_n9990__,
    new_new_n9991__, new_new_n9992__, new_new_n9993__, new_new_n9994__,
    new_new_n9995__, new_new_n9996__, new_new_n9997__, new_new_n9998__,
    new_new_n9999__, new_new_n10000__, new_new_n10001__, new_new_n10002__,
    new_new_n10003__, new_new_n10004__, new_new_n10005__, new_new_n10006__,
    new_new_n10007__, new_new_n10008__, new_new_n10009__, new_new_n10010__,
    new_new_n10011__, new_new_n10012__, new_new_n10013__, new_new_n10014__,
    new_new_n10015__, new_new_n10016__, new_new_n10017__, new_new_n10018__,
    new_new_n10019__, new_new_n10020__, new_new_n10021__, new_new_n10022__,
    new_new_n10023__, new_new_n10024__, new_new_n10025__, new_new_n10026__,
    new_new_n10027__, new_new_n10028__, new_new_n10029__, new_new_n10030__,
    new_new_n10031__, new_new_n10032__, new_new_n10033__, new_new_n10034__,
    new_new_n10035__, new_new_n10036__, new_new_n10037__, new_new_n10038__,
    new_new_n10039__, new_new_n10040__, new_new_n10041__, new_new_n10042__,
    new_new_n10043__, new_new_n10044__, new_new_n10045__, new_new_n10046__,
    new_new_n10047__, new_new_n10048__, new_new_n10049__, new_new_n10050__,
    new_new_n10051__, new_new_n10052__, new_new_n10053__, new_new_n10054__,
    new_new_n10055__, new_new_n10056__, new_new_n10057__, new_new_n10058__,
    new_new_n10059__, new_new_n10060__, new_new_n10061__, new_new_n10062__,
    new_new_n10063__, new_new_n10064__, new_new_n10065__, new_new_n10066__,
    new_new_n10067__, new_new_n10068__, new_new_n10069__, new_new_n10070__,
    new_new_n10071__, new_new_n10072__, new_new_n10073__, new_new_n10074__,
    new_new_n10075__, new_new_n10076__, new_new_n10077__, new_new_n10078__,
    new_new_n10079__, new_new_n10080__, new_new_n10081__, new_new_n10082__,
    new_new_n10083__, new_new_n10084__, new_new_n10085__, new_new_n10086__,
    new_new_n10087__, new_new_n10088__, new_new_n10089__, new_new_n10090__,
    new_new_n10091__, new_new_n10092__, new_new_n10093__, new_new_n10094__,
    new_new_n10095__, new_new_n10096__, new_new_n10097__, new_new_n10098__,
    new_new_n10099__, new_new_n10100__, new_new_n10101__, new_new_n10102__,
    new_new_n10103__, new_new_n10104__, new_new_n10105__, new_new_n10106__,
    new_new_n10107__, new_new_n10108__, new_new_n10109__, new_new_n10110__,
    new_new_n10111__, new_new_n10112__, new_new_n10113__, new_new_n10114__,
    new_new_n10115__, new_new_n10116__, new_new_n10117__, new_new_n10118__,
    new_new_n10119__, new_new_n10120__, new_new_n10121__, new_new_n10122__,
    new_new_n10123__, new_new_n10124__, new_new_n10125__, new_new_n10126__,
    new_new_n10127__, new_new_n10128__, new_new_n10129__, new_new_n10130__,
    new_new_n10131__, new_new_n10132__, new_new_n10133__, new_new_n10134__,
    new_new_n10135__, new_new_n10136__, new_new_n10137__, new_new_n10138__,
    new_new_n10139__, new_new_n10140__, new_new_n10141__, new_new_n10142__,
    new_new_n10143__, new_new_n10144__, new_new_n10145__, new_new_n10146__,
    new_new_n10147__, new_new_n10148__, new_new_n10149__, new_new_n10150__,
    new_new_n10151__, new_new_n10152__, new_new_n10153__, new_new_n10154__,
    new_new_n10155__, new_new_n10156__, new_new_n10157__, new_new_n10158__,
    new_new_n10159__, new_new_n10160__, new_new_n10161__, new_new_n10162__,
    new_new_n10163__, new_new_n10164__, new_new_n10165__, new_new_n10166__,
    new_new_n10167__, new_new_n10168__, new_new_n10169__, new_new_n10170__,
    new_new_n10171__, new_new_n10172__, new_new_n10173__, new_new_n10174__,
    new_new_n10175__, new_new_n10176__, new_new_n10177__, new_new_n10178__,
    new_new_n10179__, new_new_n10180__, new_new_n10181__, new_new_n10182__,
    new_new_n10183__, new_new_n10184__, new_new_n10185__, new_new_n10186__,
    new_new_n10187__, new_new_n10188__, new_new_n10189__, new_new_n10190__,
    new_new_n10191__, new_new_n10192__, new_new_n10193__, new_new_n10194__,
    new_new_n10195__, new_new_n10196__, new_new_n10197__, new_new_n10198__,
    new_new_n10199__, new_new_n10200__, new_new_n10201__, new_new_n10202__,
    new_new_n10203__, new_new_n10204__, new_new_n10205__, new_new_n10206__,
    new_new_n10207__, new_new_n10208__, new_new_n10209__, new_new_n10210__,
    new_new_n10211__, new_new_n10212__, new_new_n10213__, new_new_n10214__,
    new_new_n10215__, new_new_n10216__, new_new_n10217__, new_new_n10218__,
    new_new_n10219__, new_new_n10220__, new_new_n10221__, new_new_n10222__,
    new_new_n10223__, new_new_n10224__, new_new_n10225__, new_new_n10226__,
    new_new_n10227__, new_new_n10228__, new_new_n10229__, new_new_n10230__,
    new_new_n10231__, new_new_n10232__, new_new_n10233__, new_new_n10234__,
    new_new_n10235__, new_new_n10236__, new_new_n10237__, new_new_n10238__,
    new_new_n10239__, new_new_n10240__, new_new_n10241__, new_new_n10242__,
    new_new_n10243__, new_new_n10244__, new_new_n10245__, new_new_n10246__,
    new_new_n10247__, new_new_n10248__, new_new_n10249__, new_new_n10250__,
    new_new_n10251__, new_new_n10252__, new_new_n10253__, new_new_n10254__,
    new_new_n10255__, new_new_n10256__, new_new_n10257__, new_new_n10258__,
    new_new_n10259__, new_new_n10260__, new_new_n10261__, new_new_n10262__,
    new_new_n10263__, new_new_n10264__, new_new_n10265__, new_new_n10266__,
    new_new_n10267__, new_new_n10268__, new_new_n10269__, new_new_n10270__,
    new_new_n10271__, new_new_n10272__, new_new_n10273__, new_new_n10274__,
    new_new_n10275__, new_new_n10276__, new_new_n10277__, new_new_n10278__,
    new_new_n10279__, new_new_n10280__, new_new_n10281__, new_new_n10282__,
    new_new_n10283__, new_new_n10284__, new_new_n10285__, new_new_n10286__,
    new_new_n10287__, new_new_n10288__, new_new_n10289__, new_new_n10290__,
    new_new_n10291__, new_new_n10292__, new_new_n10293__, new_new_n10294__,
    new_new_n10295__, new_new_n10296__, new_new_n10297__, new_new_n10298__,
    new_new_n10299__, new_new_n10300__, new_new_n10301__, new_new_n10302__,
    new_new_n10303__, new_new_n10304__, new_new_n10305__, new_new_n10306__,
    new_new_n10307__, new_new_n10308__, new_new_n10309__, new_new_n10310__,
    new_new_n10311__, new_new_n10312__, new_new_n10313__, new_new_n10314__,
    new_new_n10315__, new_new_n10316__, new_new_n10317__, new_new_n10318__,
    new_new_n10319__, new_new_n10320__, new_new_n10321__, new_new_n10322__,
    new_new_n10323__, new_new_n10324__, new_new_n10325__, new_new_n10326__,
    new_new_n10327__, new_new_n10328__, new_new_n10329__, new_new_n10330__,
    new_new_n10331__, new_new_n10332__, new_new_n10333__, new_new_n10334__,
    new_new_n10335__, new_new_n10336__, new_new_n10337__, new_new_n10338__,
    new_new_n10339__, new_new_n10340__, new_new_n10341__, new_new_n10342__,
    new_new_n10343__, new_new_n10344__, new_new_n10345__, new_new_n10346__,
    new_new_n10347__, new_new_n10348__, new_new_n10349__, new_new_n10350__,
    new_new_n10351__, new_new_n10352__, new_new_n10353__, new_new_n10354__,
    new_new_n10355__, new_new_n10356__, new_new_n10357__, new_new_n10358__,
    new_new_n10359__, new_new_n10360__, new_new_n10361__, new_new_n10362__,
    new_new_n10363__, new_new_n10364__, new_new_n10365__, new_new_n10366__,
    new_new_n10367__, new_new_n10368__, new_new_n10369__, new_new_n10370__,
    new_new_n10371__, new_new_n10372__, new_new_n10373__, new_new_n10374__,
    new_new_n10375__, new_new_n10376__, new_new_n10377__, new_new_n10378__,
    new_new_n10379__, new_new_n10380__, new_new_n10381__, new_new_n10382__,
    new_new_n10383__, new_new_n10384__, new_new_n10385__, new_new_n10386__,
    new_new_n10387__, new_new_n10388__, new_new_n10389__, new_new_n10390__,
    new_new_n10391__, new_new_n10392__, new_new_n10393__, new_new_n10394__,
    new_new_n10395__, new_new_n10396__, new_new_n10397__, new_new_n10398__,
    new_new_n10399__, new_new_n10400__, new_new_n10401__, new_new_n10402__,
    new_new_n10403__, new_new_n10404__, new_new_n10405__, new_new_n10406__,
    new_new_n10407__, new_new_n10408__, new_new_n10409__, new_new_n10410__,
    new_new_n10411__, new_new_n10412__, new_new_n10413__, new_new_n10414__,
    new_new_n10415__, new_new_n10416__, new_new_n10417__, new_new_n10418__,
    new_new_n10419__, new_new_n10420__, new_new_n10421__, new_new_n10422__,
    new_new_n10423__, new_new_n10424__, new_new_n10425__, new_new_n10426__,
    new_new_n10427__, new_new_n10428__, new_new_n10429__, new_new_n10430__,
    new_new_n10431__, new_new_n10432__, new_new_n10433__, new_new_n10434__,
    new_new_n10435__, new_new_n10436__, new_new_n10437__, new_new_n10438__,
    new_new_n10439__, new_new_n10440__, new_new_n10441__, new_new_n10442__,
    new_new_n10443__, new_new_n10444__, new_new_n10445__, new_new_n10446__,
    new_new_n10447__, new_new_n10448__, new_new_n10449__, new_new_n10450__,
    new_new_n10451__, new_new_n10452__, new_new_n10453__, new_new_n10454__,
    new_new_n10455__, new_new_n10456__, new_new_n10457__, new_new_n10458__,
    new_new_n10459__, new_new_n10460__, new_new_n10461__, new_new_n10462__,
    new_new_n10463__, new_new_n10464__, new_new_n10465__, new_new_n10466__,
    new_new_n10467__, new_new_n10468__, new_new_n10469__, new_new_n10470__,
    new_new_n10471__, new_new_n10472__, new_new_n10473__, new_new_n10474__,
    new_new_n10475__, new_new_n10476__, new_new_n10477__, new_new_n10478__,
    new_new_n10479__, new_new_n10480__, new_new_n10481__, new_new_n10482__,
    new_new_n10483__, new_new_n10484__, new_new_n10485__, new_new_n10486__,
    new_new_n10487__, new_new_n10488__, new_new_n10489__, new_new_n10490__,
    new_new_n10491__, new_new_n10492__, new_new_n10493__, new_new_n10494__,
    new_new_n10495__, new_new_n10496__, new_new_n10497__, new_new_n10498__,
    new_new_n10499__, new_new_n10500__, new_new_n10501__, new_new_n10502__,
    new_new_n10503__, new_new_n10504__, new_new_n10505__, new_new_n10506__,
    new_new_n10507__, new_new_n10508__, new_new_n10509__, new_new_n10510__,
    new_new_n10511__, new_new_n10512__, new_new_n10513__, new_new_n10514__,
    new_new_n10515__, new_new_n10516__, new_new_n10517__, new_new_n10518__,
    new_new_n10519__, new_new_n10520__, new_new_n10521__, new_new_n10522__,
    new_new_n10523__, new_new_n10524__, new_new_n10525__, new_new_n10526__,
    new_new_n10527__, new_new_n10528__, new_new_n10529__, new_new_n10530__,
    new_new_n10531__, new_new_n10532__, new_new_n10533__, new_new_n10534__,
    new_new_n10535__, new_new_n10536__, new_new_n10537__, new_new_n10538__,
    new_new_n10539__, new_new_n10540__, new_new_n10541__, new_new_n10542__,
    new_new_n10543__, new_new_n10544__, new_new_n10545__, new_new_n10546__,
    new_new_n10547__, new_new_n10548__, new_new_n10549__, new_new_n10550__,
    new_new_n10551__, new_new_n10552__, new_new_n10553__, new_new_n10554__,
    new_new_n10555__, new_new_n10556__, new_new_n10557__, new_new_n10558__,
    new_new_n10559__, new_new_n10560__, new_new_n10561__, new_new_n10562__,
    new_new_n10563__, new_new_n10564__, n16425, n16428, n16431, n16434,
    n16437, n16440, n16443, n16446, n16449, n16452, n16455, n16458, n16461,
    n16464, n16467, n16470, n16473, n16476, n16479, n16482, n16485, n16488,
    n16491, n16494, n16497, n16500, n16503, n16506, n16509, n16512, n16515,
    n16518, n16521, n16524, n16527, n16530, n16533, n16536, n16539, n16542,
    n16545, n16548, n16551, n16554, n16557, n16560, n16563, n16566, n16569,
    n16572, n16575, n16578, n16581, n16584, n16587, n16590, n16593, n16596,
    n16599, n16602, n16605, n16608, n16611, n16614, n16617, n16620, n16623,
    n16626, n16629, n16632, n16635, n16638, n16641, n16644, n16647, n16650,
    n16653, n16656, n16659, n16662, n16665, n16668, n16671, n16674, n16677,
    n16680, n16683, n16686, n16689, n16692, n16695, n16698, n16701, n16704,
    n16707, n16710, n16713, n16716, n16719, n16722, n16725, n16728, n16731,
    n16734, n16737, n16740, n16743, n16746, n16749, n16752, n16755, n16758,
    n16761, n16764, n16767, n16770, n16773, n16776, n16779, n16782, n16785,
    n16788, n16791, n16794, n16797, n16800, n16803, n16806, n16809, n16812,
    n16815, n16818, n16821, n16824, n16827, n16830, n16833, n16836, n16839,
    n16842, n16845, n16848, n16851, n16854, n16857, n16860, n16863, n16866,
    n16869, n16872, n16875, n16878, n16881, n16884, n16887, n16890, n16893,
    n16896, n16899, n16902, n16905, n16908, n16911, n16914, n16917, n16920,
    n16923, n16926, n16929, n16932, n16935, n16938, n16941, n16944, n16947,
    n16950, n16953, n16956, n16959, n16962, n16965, n16968, n16971, n16974,
    n16977, n16980, n16983, n16986, n16989, n16992, n16995, n16998, n17001,
    n17004, n17007, n17010, n17013, n17016, n17019, n17022, n17025, n17028,
    n17031, n17034, n17037, n17040, n17043, n17046, n17049, n17052, n17055,
    n17058, n17061, n17064, n17067, n17070, n17073, n17076, n17079, n17082,
    n17085, n17088, n17091, n17094, n17097, n17100, n17103, n17106, n17109,
    n17112, n17115, n17118, n17121, n17124, n17127, n17130, n17133, n17136,
    n17139, n17142, n17145, n17148, n17151, n17154, n17157, n17160, n17163,
    n17166, n17169, n17172, n17175, n17178, n17181, n17184, n17187, n17190,
    n17193, n17196, n17199, n17202, n17205, n17208, n17211, n17214, n17217,
    n17220, n17223, n17226, n17229, n17232, n17235, n17238, n17241, n17244,
    n17247, n17250, n17253, n17256, n17259, n17262, n17265, n17268, n17271,
    n17274, n17277, n17280, n17283, n17286, n17289, n17292, n17295, n17298,
    n17301, n17304, n17307, n17310, n17313, n17316, n17319, n17322, n17325,
    n17328, n17331, n17334, n17337, n17340, n17343, n17346, n17349, n17352,
    n17355, n17358, n17361, n17364, n17367, n17370, n17373, n17376, n17379,
    n17382, n17385, n17388, n17391, n17394, n17397, n17400, n17403, n17406,
    n17409, n17412, n17415, n17418, n17421, n17424, n17427, n17430, n17433,
    n17436, n17439, n17442, n17445, n17448, n17451, n17454, n17457, n17460,
    n17463, n17466, n17469, n17472, n17475, n17478, n17481, n17484, n17487,
    n17490, n17493, n17496, n17499, n17502, n17505, n17508, n17511, n17514,
    n17517, n17520, n17523, n17526, n17529, n17532, n17535, n17538, n17541,
    n17544, n17547, n17550, n17553, n17556, n17559, n17562, n17565, n17568,
    n17571, n17574, n17577, n17580, n17583, n17586, n17589, n17592, n17595,
    n17598, n17601, n17604, n17607, n17610, n17613, n17616, n17619, n17622,
    n17625, n17628, n17631, n17634, n17637, n17640, n17643, n17646, n17649,
    n17652, n17655, n17658, n17661, n17664, n17667, n17670, n17673, n17676,
    n17679, n17682, n17685, n17688, n17691, n17694, n17697, n17700, n17703,
    n17706, n17709, n17712, n17715, n17718, n17721, n17724, n17727, n17730,
    n17733, n17736, n17739, n17742, n17745, n17748, n17751, n17754, n17757,
    n17760, n17763, n17766, n17769, n17772, n17775, n17778, n17781, n17784,
    n17787, n17790, n17793, n17796, n17799, n17802, n17805, n17808, n17811,
    n17814, n17817, n17820, n17823, n17826, n17829, n17832, n17835, n17838,
    n17841, n17844, n17847, n17850, n17853, n17856, n17859, n17862, n17865,
    n17868, n17871, n17874, n17877, n17880, n17883, n17886, n17889, n17892,
    n17895, n17898, n17901, n17904, n17907, n17910, n17913, n17916, n17919,
    n17922, n17925, n17928, n17931, n17934, n17937, n17940, n17943, n17946,
    n17949, n17952, n17955, n17958, n17961, n17964, n17967, n17970, n17973,
    n17976, n17979, n17982, n17985, n17988, n17991, n17994, n17997, n18000,
    n18003, n18006, n18009, n18012, n18015, n18018, n18021, n18024, n18027,
    n18030, n18033, n18036, n18039, n18042, n18045, n18048, n18051, n18054,
    n18057, n18060, n18063, n18066, n18069, n18072, n18075, n18078, n18081,
    n18084, n18087, n18090, n18093, n18096, n18099, n18102, n18105, n18108,
    n18111, n18114, n18117, n18120, n18123, n18126, n18129, n18132, n18135,
    n18138, n18141, n18144, n18147, n18150, n18153, n18156, n18159, n18162,
    n18165, n18168, n18171, n18174, n18177, n18180, n18183, n18186, n18189,
    n18192, n18195, n18198, n18201, n18204, n18207, n18210, n18213, n18216,
    n18219, n18222, n18225, n18228, n18231, n18234, n18237, n18240, n18243,
    n18246, n18249, n18252, n18255, n18258, n18261, n18264, n18267, n18270,
    n18273, n18276, n18279, n18282, n18285, n18288, n18291, n18294, n18297,
    n18300, n18303, n18306, n18309, n18312, n18315, n18318, n18321, n18324,
    n18327, n18330, n18333, n18336, n18339, n18342, n18345, n18348, n18351,
    n18354, n18357, n18360, n18363, n18366, n18369, n18372, n18375, n18378,
    n18381, n18384, n18387, n18390, n18393, n18396, n18399, n18402, n18405,
    n18408, n18411, n18414, n18417, n18420, n18423, n18426, n18429, n18432,
    n18435, n18438, n18441, n18444, n18447, n18450, n18453, n18456, n18459,
    n18462, n18465, n18468, n18471, n18474, n18477, n18480, n18483, n18486,
    n18489, n18492, n18495, n18498, n18501, n18504, n18507, n18510, n18513,
    n18516, n18519, n18522, n18525, n18528, n18531, n18534, n18537, n18540,
    n18543, n18546, n18549, n18552, n18555, n18558, n18561, n18564, n18567,
    n18570, n18573, n18576, n18579, n18582, n18585, n18588, n18591, n18594,
    n18597, n18600, n18603, n18606, n18609, n18612, n18615, n18618, n18621,
    n18624, n18627, n18630, n18633, n18636, n18639, n18642, n18645, n18648,
    n18651, n18654, n18657, n18660, n18663, n18666, n18669, n18672, n18675,
    n18678, n18681, n18684, n18687, n18690, n18693, n18696, n18699, n18702,
    n18705, n18708, n18711, n18714, n18717, n18720, n18723, n18726, n18729,
    n18732, n18735, n18738, n18741, n18744, n18747, n18750, n18753, n18756,
    n18759, n18762, n18765, n18768, n18771, n18774, n18777, n18780, n18783,
    n18786, n18789, n18792, n18795, n18798, n18801, n18804, n18807, n18810,
    n18813, n18816, n18819, n18822, n18825, n18828, n18831, n18834, n18837,
    n18840, n18843, n18846, n18849, n18852, n18855, n18858, n18861, n18864,
    n18867, n18870, n18873, n18876, n18879, n18882, n18885, n18888, n18891,
    n18894, n18897, n18900, n18903, n18906, n18909, n18912, n18915, n18918,
    n18921, n18924, n18927, n18930, n18933, n18936, n18939, n18942, n18945,
    n18948, n18951, n18954, n18957, n18960, n18963, n18966, n18969, n18972,
    n18975, n18978, n18981, n18984, n18987, n18990, n18993, n18996, n18999,
    n19002, n19005, n19008, n19011, n19014, n19017, n19020, n19023, n19026,
    n19029, n19032, n19035, n19038, n19041, n19044, n19047, n19050, n19053,
    n19056, n19059, n19062, n19065, n19068, n19071, n19074, n19077, n19080,
    n19083, n19086, n19089, n19092, n19095, n19098, n19101, n19104, n19107,
    n19110, n19113, n19116, n19119, n19122, n19125, n19128, n19131, n19134,
    n19137, n19140, n19143, n19146, n19149, n19152, n19155, n19158, n19161,
    n19164, n19167, n19170, n19173, n19176, n19179, n19182, n19185, n19188,
    n19191, n19194, n19197, n19200, n19203, n19206, n19209, n19212, n19215,
    n19218, n19221, n19224, n19227, n19230, n19233, n19236, n19239, n19242,
    n19245, n19248, n19251, n19254, n19257, n19260, n19263, n19266, n19269,
    n19272, n19275, n19278, n19281, n19284, n19287, n19290, n19293, n19296,
    n19299, n19302, n19305, n19308, n19311, n19314, n19317, n19320, n19323,
    n19326, n19329, n19332, n19335, n19338, n19341, n19344, n19347, n19350,
    n19353, n19356, n19359, n19362, n19365, n19368, n19371, n19374, n19377,
    n19380, n19383, n19386, n19389, n19392, n19395, n19398, n19401, n19404,
    n19407, n19410, n19413, n19416, n19419, n19422, n19425, n19428, n19431,
    n19434, n19437, n19440, n19443, n19446, n19449, n19452, n19455, n19458,
    n19461;
  buf1  g0000(.din(G1), .dout(new_new_n2328__));
  buf1  g0001(.din(G2), .dout(new_new_n2330__));
  buf1  g0002(.din(G3), .dout(new_new_n2332__));
  buf1  g0003(.din(G4), .dout(new_new_n2334__));
  buf1  g0004(.din(G5), .dout(new_new_n2336__));
  buf1  g0005(.din(G6), .dout(new_new_n2338__));
  buf1  g0006(.din(G7), .dout(new_new_n2340__));
  buf1  g0007(.din(G8), .dout(new_new_n2342__));
  buf1  g0008(.din(G9), .dout(new_new_n2344__));
  buf1  g0009(.din(G10), .dout(new_new_n2346__));
  buf1  g0010(.din(G11), .dout(new_new_n2348__));
  buf1  g0011(.din(G12), .dout(new_new_n2350__));
  buf1  g0012(.din(G13), .dout(new_new_n2352__));
  buf1  g0013(.din(G14), .dout(new_new_n2354__));
  buf1  g0014(.din(G15), .dout(new_new_n2356__));
  buf1  g0015(.din(G16), .dout(new_new_n2358__));
  buf1  g0016(.din(G17), .dout(new_new_n2360__));
  buf1  g0017(.din(G18), .dout(new_new_n2362__));
  buf1  g0018(.din(G19), .dout(new_new_n2364__));
  buf1  g0019(.din(G20), .dout(new_new_n2366__));
  buf1  g0020(.din(G21), .dout(new_new_n2368__));
  buf1  g0021(.din(G22), .dout(new_new_n2370__));
  buf1  g0022(.din(G23), .dout(new_new_n2372__));
  buf1  g0023(.din(G24), .dout(new_new_n2374__));
  buf1  g0024(.din(G25), .dout(new_new_n2376__));
  buf1  g0025(.din(G26), .dout(new_new_n2378__));
  buf1  g0026(.din(G27), .dout(new_new_n2380__));
  buf1  g0027(.din(G28), .dout(new_new_n2382__));
  buf1  g0028(.din(G29), .dout(new_new_n2384__));
  buf1  g0029(.din(G30), .dout(new_new_n2386__));
  buf1  g0030(.din(G31), .dout(new_new_n2388__));
  buf1  g0031(.din(G32), .dout(new_new_n2390__));
  buf1  g0032(.din(G33), .dout(new_new_n2392__));
  buf1  g0033(.din(G34), .dout(new_new_n2394__));
  buf1  g0034(.din(G35), .dout(new_new_n2396__));
  buf1  g0035(.din(G36), .dout(new_new_n2398__));
  buf1  g0036(.din(G37), .dout(new_new_n2400__));
  buf1  g0037(.din(G38), .dout(new_new_n2402__));
  buf1  g0038(.din(G39), .dout(new_new_n2404__));
  buf1  g0039(.din(G40), .dout(new_new_n2406__));
  buf1  g0040(.din(G41), .dout(new_new_n2408__));
  buf1  g0041(.din(G42), .dout(new_new_n2410__));
  buf1  g0042(.din(G43), .dout(new_new_n2412__));
  buf1  g0043(.din(G44), .dout(new_new_n2414__));
  buf1  g0044(.din(G45), .dout(new_new_n2416__));
  buf1  g0045(.din(G46), .dout(new_new_n2418__));
  buf1  g0046(.din(G47), .dout(new_new_n2420__));
  buf1  g0047(.din(G48), .dout(new_new_n2422__));
  buf1  g0048(.din(G49), .dout(new_new_n2424__));
  buf1  g0049(.din(G50), .dout(new_new_n2426__));
  buf1  g0050(.din(G51), .dout(new_new_n2428__));
  buf1  g0051(.din(G52), .dout(new_new_n2430__));
  buf1  g0052(.din(G53), .dout(new_new_n2432__));
  buf1  g0053(.din(G54), .dout(new_new_n2434__));
  buf1  g0054(.din(G55), .dout(new_new_n2436__));
  buf1  g0055(.din(G56), .dout(new_new_n2438__));
  buf1  g0056(.din(G57), .dout(new_new_n2440__));
  buf1  g0057(.din(G58), .dout(new_new_n2442__));
  buf1  g0058(.din(G59), .dout(new_new_n2444__));
  buf1  g0059(.din(G60), .dout(new_new_n2446__));
  buf1  g0060(.din(G61), .dout(new_new_n2448__));
  buf1  g0061(.din(G62), .dout(new_new_n2450__));
  buf1  g0062(.din(G63), .dout(new_new_n2452__));
  buf1  g0063(.din(G64), .dout(new_new_n2454__));
  buf1  g0064(.din(G65), .dout(new_new_n2456__));
  buf1  g0065(.din(G66), .dout(new_new_n2458__));
  buf1  g0066(.din(G67), .dout(new_new_n2460__));
  buf1  g0067(.din(G68), .dout(new_new_n2462__));
  buf1  g0068(.din(G69), .dout(new_new_n2464__));
  buf1  g0069(.din(G70), .dout(new_new_n2466__));
  buf1  g0070(.din(G71), .dout(new_new_n2468__));
  buf1  g0071(.din(G72), .dout(new_new_n2470__));
  buf1  g0072(.din(G73), .dout(new_new_n2472__));
  buf1  g0073(.din(G74), .dout(new_new_n2474__));
  buf1  g0074(.din(G75), .dout(new_new_n2476__));
  buf1  g0075(.din(G76), .dout(new_new_n2478__));
  buf1  g0076(.din(G77), .dout(new_new_n2480__));
  buf1  g0077(.din(G78), .dout(new_new_n2482__));
  buf1  g0078(.din(G79), .dout(new_new_n2484__));
  buf1  g0079(.din(G80), .dout(new_new_n2486__));
  buf1  g0080(.din(G81), .dout(new_new_n2488__));
  buf1  g0081(.din(G82), .dout(new_new_n2490__));
  buf1  g0082(.din(G83), .dout(new_new_n2492__));
  buf1  g0083(.din(G84), .dout(new_new_n2494__));
  buf1  g0084(.din(G85), .dout(new_new_n2496__));
  buf1  g0085(.din(G86), .dout(new_new_n2498__));
  buf1  g0086(.din(G87), .dout(new_new_n2500__));
  buf1  g0087(.din(G88), .dout(new_new_n2502__));
  buf1  g0088(.din(G89), .dout(new_new_n2504__));
  buf1  g0089(.din(G90), .dout(new_new_n2506__));
  buf1  g0090(.din(G91), .dout(new_new_n2508__));
  buf1  g0091(.din(G92), .dout(new_new_n2510__));
  buf1  g0092(.din(G93), .dout(new_new_n2512__));
  buf1  g0093(.din(G94), .dout(new_new_n2514__));
  buf1  g0094(.din(G95), .dout(new_new_n2516__));
  buf1  g0095(.din(G96), .dout(new_new_n2518__));
  buf1  g0096(.din(G97), .dout(new_new_n2520__));
  buf1  g0097(.din(G98), .dout(new_new_n2522__));
  buf1  g0098(.din(G99), .dout(new_new_n2524__));
  buf1  g0099(.din(G100), .dout(new_new_n2526__));
  buf1  g0100(.din(G101), .dout(new_new_n2528__));
  buf1  g0101(.din(G102), .dout(new_new_n2530__));
  buf1  g0102(.din(G103), .dout(new_new_n2532__));
  buf1  g0103(.din(G104), .dout(new_new_n2534__));
  buf1  g0104(.din(G105), .dout(new_new_n2536__));
  buf1  g0105(.din(G106), .dout(new_new_n2538__));
  buf1  g0106(.din(G107), .dout(new_new_n2540__));
  buf1  g0107(.din(G108), .dout(new_new_n2542__));
  buf1  g0108(.din(G109), .dout(new_new_n2544__));
  buf1  g0109(.din(G110), .dout(new_new_n2546__));
  buf1  g0110(.din(G111), .dout(new_new_n2548__));
  buf1  g0111(.din(G112), .dout(new_new_n2550__));
  buf1  g0112(.din(G113), .dout(new_new_n2552__));
  buf1  g0113(.din(G114), .dout(new_new_n2554__));
  buf1  g0114(.din(G115), .dout(new_new_n2556__));
  buf1  g0115(.din(G116), .dout(new_new_n2558__));
  buf1  g0116(.din(G117), .dout(new_new_n2560__));
  buf1  g0117(.din(G118), .dout(new_new_n2562__));
  buf1  g0118(.din(G119), .dout(new_new_n2564__));
  buf1  g0119(.din(G120), .dout(new_new_n2566__));
  buf1  g0120(.din(G121), .dout(new_new_n2568__));
  buf1  g0121(.din(G122), .dout(new_new_n2570__));
  buf1  g0122(.din(G123), .dout(new_new_n2572__));
  not1  g0123(.din(G123), .dout(new_new_n2573__));
  buf1  g0124(.din(G124), .dout(new_new_n2574__));
  not1  g0125(.din(G124), .dout(new_new_n2575__));
  buf1  g0126(.din(G125), .dout(new_new_n2576__));
  buf1  g0127(.din(G126), .dout(new_new_n2578__));
  buf1  g0128(.din(G127), .dout(new_new_n2580__));
  buf1  g0129(.din(G128), .dout(new_new_n2582__));
  buf1  g0130(.din(G129), .dout(new_new_n2584__));
  buf1  g0131(.din(G130), .dout(new_new_n2586__));
  buf1  g0132(.din(G131), .dout(new_new_n2588__));
  buf1  g0133(.din(G132), .dout(new_new_n2590__));
  buf1  g0134(.din(G133), .dout(new_new_n2592__));
  buf1  g0135(.din(G134), .dout(new_new_n2594__));
  buf1  g0136(.din(G135), .dout(new_new_n2596__));
  buf1  g0137(.din(G136), .dout(new_new_n2598__));
  buf1  g0138(.din(G137), .dout(new_new_n2600__));
  buf1  g0139(.din(G138), .dout(new_new_n2602__));
  buf1  g0140(.din(G139), .dout(new_new_n2604__));
  buf1  g0141(.din(G140), .dout(new_new_n2606__));
  buf1  g0142(.din(G141), .dout(new_new_n2608__));
  buf1  g0143(.din(G142), .dout(new_new_n2610__));
  buf1  g0144(.din(G143), .dout(new_new_n2612__));
  buf1  g0145(.din(G144), .dout(new_new_n2614__));
  buf1  g0146(.din(G145), .dout(new_new_n2616__));
  buf1  g0147(.din(G146), .dout(new_new_n2618__));
  buf1  g0148(.din(G147), .dout(new_new_n2620__));
  buf1  g0149(.din(G148), .dout(new_new_n2622__));
  buf1  g0150(.din(G149), .dout(new_new_n2624__));
  buf1  g0151(.din(G150), .dout(new_new_n2626__));
  buf1  g0152(.din(G151), .dout(new_new_n2628__));
  buf1  g0153(.din(G152), .dout(new_new_n2630__));
  buf1  g0154(.din(G153), .dout(new_new_n2632__));
  buf1  g0155(.din(G154), .dout(new_new_n2634__));
  buf1  g0156(.din(G155), .dout(new_new_n2636__));
  buf1  g0157(.din(G156), .dout(new_new_n2638__));
  buf1  g0158(.din(G157), .dout(new_new_n2640__));
  buf1  g0159(.din(G158), .dout(new_new_n2642__));
  buf1  g0160(.din(G159), .dout(new_new_n2644__));
  buf1  g0161(.din(G160), .dout(new_new_n2646__));
  buf1  g0162(.din(G161), .dout(new_new_n2648__));
  buf1  g0163(.din(G162), .dout(new_new_n2650__));
  buf1  g0164(.din(G163), .dout(new_new_n2652__));
  buf1  g0165(.din(G164), .dout(new_new_n2654__));
  buf1  g0166(.din(G165), .dout(new_new_n2656__));
  buf1  g0167(.din(G166), .dout(new_new_n2658__));
  buf1  g0168(.din(G167), .dout(new_new_n2660__));
  buf1  g0169(.din(G168), .dout(new_new_n2662__));
  buf1  g0170(.din(G169), .dout(new_new_n2664__));
  buf1  g0171(.din(G170), .dout(new_new_n2666__));
  buf1  g0172(.din(G171), .dout(new_new_n2668__));
  buf1  g0173(.din(G172), .dout(new_new_n2670__));
  buf1  g0174(.din(G173), .dout(new_new_n2672__));
  buf1  g0175(.din(G174), .dout(new_new_n2674__));
  buf1  g0176(.din(G175), .dout(new_new_n2676__));
  buf1  g0177(.din(G176), .dout(new_new_n2678__));
  buf1  g0178(.din(G177), .dout(new_new_n2680__));
  buf1  g0179(.din(G178), .dout(new_new_n2682__));
  buf1  g0180(.din(n2610_lo), .dout(new_new_n2684__));
  buf1  g0181(.din(n2613_lo), .dout(new_new_n2686__));
  buf1  g0182(.din(n2616_lo), .dout(new_new_n2688__));
  buf1  g0183(.din(n2619_lo), .dout(new_new_n2690__));
  not1  g0184(.din(n2619_lo), .dout(new_new_n2691__));
  buf1  g0185(.din(n2622_lo), .dout(new_new_n2692__));
  buf1  g0186(.din(n2625_lo), .dout(new_new_n2694__));
  buf1  g0187(.din(n2628_lo), .dout(new_new_n2696__));
  buf1  g0188(.din(n2631_lo), .dout(new_new_n2698__));
  not1  g0189(.din(n2631_lo), .dout(new_new_n2699__));
  buf1  g0190(.din(n2634_lo), .dout(new_new_n2700__));
  buf1  g0191(.din(n2637_lo), .dout(new_new_n2702__));
  buf1  g0192(.din(n2640_lo), .dout(new_new_n2704__));
  buf1  g0193(.din(n2643_lo), .dout(new_new_n2706__));
  buf1  g0194(.din(n2646_lo), .dout(new_new_n2708__));
  buf1  g0195(.din(n2649_lo), .dout(new_new_n2710__));
  buf1  g0196(.din(n2652_lo), .dout(new_new_n2712__));
  buf1  g0197(.din(n2655_lo), .dout(new_new_n2714__));
  buf1  g0198(.din(n2658_lo), .dout(new_new_n2716__));
  buf1  g0199(.din(n2661_lo), .dout(new_new_n2718__));
  buf1  g0200(.din(n2664_lo), .dout(new_new_n2720__));
  buf1  g0201(.din(n2667_lo), .dout(new_new_n2722__));
  buf1  g0202(.din(n2670_lo), .dout(new_new_n2724__));
  buf1  g0203(.din(n2673_lo), .dout(new_new_n2726__));
  buf1  g0204(.din(n2676_lo), .dout(new_new_n2728__));
  buf1  g0205(.din(n2679_lo), .dout(new_new_n2730__));
  buf1  g0206(.din(n2682_lo), .dout(new_new_n2732__));
  buf1  g0207(.din(n2685_lo), .dout(new_new_n2734__));
  buf1  g0208(.din(n2688_lo), .dout(new_new_n2736__));
  not1  g0209(.din(n2691_lo), .dout(new_new_n2739__));
  buf1  g0210(.din(n2694_lo), .dout(new_new_n2740__));
  buf1  g0211(.din(n2697_lo), .dout(new_new_n2742__));
  buf1  g0212(.din(n2700_lo), .dout(new_new_n2744__));
  not1  g0213(.din(n2703_lo), .dout(new_new_n2747__));
  buf1  g0214(.din(n2706_lo), .dout(new_new_n2748__));
  buf1  g0215(.din(n2709_lo), .dout(new_new_n2750__));
  buf1  g0216(.din(n2712_lo), .dout(new_new_n2752__));
  not1  g0217(.din(n2715_lo), .dout(new_new_n2755__));
  buf1  g0218(.din(n2718_lo), .dout(new_new_n2756__));
  buf1  g0219(.din(n2721_lo), .dout(new_new_n2758__));
  buf1  g0220(.din(n2724_lo), .dout(new_new_n2760__));
  not1  g0221(.din(n2727_lo), .dout(new_new_n2763__));
  buf1  g0222(.din(n2730_lo), .dout(new_new_n2764__));
  buf1  g0223(.din(n2733_lo), .dout(new_new_n2766__));
  buf1  g0224(.din(n2736_lo), .dout(new_new_n2768__));
  buf1  g0225(.din(n2739_lo), .dout(new_new_n2770__));
  not1  g0226(.din(n2739_lo), .dout(new_new_n2771__));
  buf1  g0227(.din(n2742_lo), .dout(new_new_n2772__));
  buf1  g0228(.din(n2745_lo), .dout(new_new_n2774__));
  buf1  g0229(.din(n2748_lo), .dout(new_new_n2776__));
  buf1  g0230(.din(n2751_lo), .dout(new_new_n2778__));
  not1  g0231(.din(n2751_lo), .dout(new_new_n2779__));
  buf1  g0232(.din(n2754_lo), .dout(new_new_n2780__));
  buf1  g0233(.din(n2757_lo), .dout(new_new_n2782__));
  buf1  g0234(.din(n2760_lo), .dout(new_new_n2784__));
  not1  g0235(.din(n2763_lo), .dout(new_new_n2787__));
  buf1  g0236(.din(n2766_lo), .dout(new_new_n2788__));
  buf1  g0237(.din(n2769_lo), .dout(new_new_n2790__));
  buf1  g0238(.din(n2772_lo), .dout(new_new_n2792__));
  buf1  g0239(.din(n2775_lo), .dout(new_new_n2794__));
  buf1  g0240(.din(n2778_lo), .dout(new_new_n2796__));
  buf1  g0241(.din(n2781_lo), .dout(new_new_n2798__));
  buf1  g0242(.din(n2784_lo), .dout(new_new_n2800__));
  buf1  g0243(.din(n2787_lo), .dout(new_new_n2802__));
  buf1  g0244(.din(n2790_lo), .dout(new_new_n2804__));
  buf1  g0245(.din(n2793_lo), .dout(new_new_n2806__));
  buf1  g0246(.din(n2796_lo), .dout(new_new_n2808__));
  buf1  g0247(.din(n2799_lo), .dout(new_new_n2810__));
  buf1  g0248(.din(n2802_lo), .dout(new_new_n2812__));
  buf1  g0249(.din(n2805_lo), .dout(new_new_n2814__));
  buf1  g0250(.din(n2808_lo), .dout(new_new_n2816__));
  buf1  g0251(.din(n2811_lo), .dout(new_new_n2818__));
  buf1  g0252(.din(n2814_lo), .dout(new_new_n2820__));
  buf1  g0253(.din(n2817_lo), .dout(new_new_n2822__));
  buf1  g0254(.din(n2820_lo), .dout(new_new_n2824__));
  buf1  g0255(.din(n2823_lo), .dout(new_new_n2826__));
  buf1  g0256(.din(n2826_lo), .dout(new_new_n2828__));
  buf1  g0257(.din(n2829_lo), .dout(new_new_n2830__));
  buf1  g0258(.din(n2832_lo), .dout(new_new_n2832__));
  buf1  g0259(.din(n2835_lo), .dout(new_new_n2834__));
  buf1  g0260(.din(n2838_lo), .dout(new_new_n2836__));
  buf1  g0261(.din(n2841_lo), .dout(new_new_n2838__));
  buf1  g0262(.din(n2844_lo), .dout(new_new_n2840__));
  buf1  g0263(.din(n2847_lo), .dout(new_new_n2842__));
  buf1  g0264(.din(n2850_lo), .dout(new_new_n2844__));
  buf1  g0265(.din(n2853_lo), .dout(new_new_n2846__));
  buf1  g0266(.din(n2856_lo), .dout(new_new_n2848__));
  buf1  g0267(.din(n2859_lo), .dout(new_new_n2850__));
  not1  g0268(.din(n2859_lo), .dout(new_new_n2851__));
  buf1  g0269(.din(n2862_lo), .dout(new_new_n2852__));
  buf1  g0270(.din(n2865_lo), .dout(new_new_n2854__));
  buf1  g0271(.din(n2868_lo), .dout(new_new_n2856__));
  buf1  g0272(.din(n2871_lo), .dout(new_new_n2858__));
  buf1  g0273(.din(n2874_lo), .dout(new_new_n2860__));
  buf1  g0274(.din(n2877_lo), .dout(new_new_n2862__));
  buf1  g0275(.din(n2880_lo), .dout(new_new_n2864__));
  buf1  g0276(.din(n2883_lo), .dout(new_new_n2866__));
  buf1  g0277(.din(n2886_lo), .dout(new_new_n2868__));
  buf1  g0278(.din(n2889_lo), .dout(new_new_n2870__));
  buf1  g0279(.din(n2892_lo), .dout(new_new_n2872__));
  buf1  g0280(.din(n2895_lo), .dout(new_new_n2874__));
  buf1  g0281(.din(n2898_lo), .dout(new_new_n2876__));
  buf1  g0282(.din(n2901_lo), .dout(new_new_n2878__));
  buf1  g0283(.din(n2904_lo), .dout(new_new_n2880__));
  buf1  g0284(.din(n2907_lo), .dout(new_new_n2882__));
  buf1  g0285(.din(n2910_lo), .dout(new_new_n2884__));
  buf1  g0286(.din(n2913_lo), .dout(new_new_n2886__));
  buf1  g0287(.din(n2916_lo), .dout(new_new_n2888__));
  buf1  g0288(.din(n2919_lo), .dout(new_new_n2890__));
  buf1  g0289(.din(n2922_lo), .dout(new_new_n2892__));
  buf1  g0290(.din(n2925_lo), .dout(new_new_n2894__));
  buf1  g0291(.din(n2928_lo), .dout(new_new_n2896__));
  buf1  g0292(.din(n2931_lo), .dout(new_new_n2898__));
  buf1  g0293(.din(n2934_lo), .dout(new_new_n2900__));
  buf1  g0294(.din(n2937_lo), .dout(new_new_n2902__));
  buf1  g0295(.din(n2940_lo), .dout(new_new_n2904__));
  not1  g0296(.din(n2943_lo), .dout(new_new_n2907__));
  buf1  g0297(.din(n2946_lo), .dout(new_new_n2908__));
  buf1  g0298(.din(n2949_lo), .dout(new_new_n2910__));
  buf1  g0299(.din(n2952_lo), .dout(new_new_n2912__));
  not1  g0300(.din(n2955_lo), .dout(new_new_n2915__));
  buf1  g0301(.din(n2958_lo), .dout(new_new_n2916__));
  buf1  g0302(.din(n2961_lo), .dout(new_new_n2918__));
  buf1  g0303(.din(n2964_lo), .dout(new_new_n2920__));
  not1  g0304(.din(n2967_lo), .dout(new_new_n2923__));
  buf1  g0305(.din(n2970_lo), .dout(new_new_n2924__));
  buf1  g0306(.din(n2973_lo), .dout(new_new_n2926__));
  buf1  g0307(.din(n2976_lo), .dout(new_new_n2928__));
  not1  g0308(.din(n2979_lo), .dout(new_new_n2931__));
  buf1  g0309(.din(n2982_lo), .dout(new_new_n2932__));
  buf1  g0310(.din(n2985_lo), .dout(new_new_n2934__));
  buf1  g0311(.din(n2988_lo), .dout(new_new_n2936__));
  not1  g0312(.din(n2991_lo), .dout(new_new_n2939__));
  buf1  g0313(.din(n2994_lo), .dout(new_new_n2940__));
  buf1  g0314(.din(n2997_lo), .dout(new_new_n2942__));
  buf1  g0315(.din(n3000_lo), .dout(new_new_n2944__));
  not1  g0316(.din(n3003_lo), .dout(new_new_n2947__));
  buf1  g0317(.din(n3006_lo), .dout(new_new_n2948__));
  buf1  g0318(.din(n3009_lo), .dout(new_new_n2950__));
  buf1  g0319(.din(n3012_lo), .dout(new_new_n2952__));
  not1  g0320(.din(n3015_lo), .dout(new_new_n2955__));
  buf1  g0321(.din(n3018_lo), .dout(new_new_n2956__));
  buf1  g0322(.din(n3021_lo), .dout(new_new_n2958__));
  buf1  g0323(.din(n3024_lo), .dout(new_new_n2960__));
  not1  g0324(.din(n3027_lo), .dout(new_new_n2963__));
  buf1  g0325(.din(n3030_lo), .dout(new_new_n2964__));
  buf1  g0326(.din(n3033_lo), .dout(new_new_n2966__));
  buf1  g0327(.din(n3036_lo), .dout(new_new_n2968__));
  buf1  g0328(.din(n3039_lo), .dout(new_new_n2970__));
  buf1  g0329(.din(n3042_lo), .dout(new_new_n2972__));
  buf1  g0330(.din(n3045_lo), .dout(new_new_n2974__));
  buf1  g0331(.din(n3048_lo), .dout(new_new_n2976__));
  buf1  g0332(.din(n3051_lo), .dout(new_new_n2978__));
  buf1  g0333(.din(n3054_lo), .dout(new_new_n2980__));
  buf1  g0334(.din(n3057_lo), .dout(new_new_n2982__));
  buf1  g0335(.din(n3060_lo), .dout(new_new_n2984__));
  buf1  g0336(.din(n3063_lo), .dout(new_new_n2986__));
  buf1  g0337(.din(n3066_lo), .dout(new_new_n2988__));
  buf1  g0338(.din(n3069_lo), .dout(new_new_n2990__));
  buf1  g0339(.din(n3072_lo), .dout(new_new_n2992__));
  buf1  g0340(.din(n3075_lo), .dout(new_new_n2994__));
  buf1  g0341(.din(n3078_lo), .dout(new_new_n2996__));
  buf1  g0342(.din(n3081_lo), .dout(new_new_n2998__));
  buf1  g0343(.din(n3084_lo), .dout(new_new_n3000__));
  buf1  g0344(.din(n3087_lo), .dout(new_new_n3002__));
  buf1  g0345(.din(n3090_lo), .dout(new_new_n3004__));
  buf1  g0346(.din(n3093_lo), .dout(new_new_n3006__));
  buf1  g0347(.din(n3096_lo), .dout(new_new_n3008__));
  buf1  g0348(.din(n3099_lo), .dout(new_new_n3010__));
  buf1  g0349(.din(n3102_lo), .dout(new_new_n3012__));
  buf1  g0350(.din(n3105_lo), .dout(new_new_n3014__));
  buf1  g0351(.din(n3108_lo), .dout(new_new_n3016__));
  buf1  g0352(.din(n3111_lo), .dout(new_new_n3018__));
  buf1  g0353(.din(n3114_lo), .dout(new_new_n3020__));
  buf1  g0354(.din(n3117_lo), .dout(new_new_n3022__));
  buf1  g0355(.din(n3120_lo), .dout(new_new_n3024__));
  buf1  g0356(.din(n3123_lo), .dout(new_new_n3026__));
  buf1  g0357(.din(n3126_lo), .dout(new_new_n3028__));
  buf1  g0358(.din(n3129_lo), .dout(new_new_n3030__));
  buf1  g0359(.din(n3132_lo), .dout(new_new_n3032__));
  buf1  g0360(.din(n3135_lo), .dout(new_new_n3034__));
  buf1  g0361(.din(n3138_lo), .dout(new_new_n3036__));
  buf1  g0362(.din(n3141_lo), .dout(new_new_n3038__));
  buf1  g0363(.din(n3144_lo), .dout(new_new_n3040__));
  buf1  g0364(.din(n3147_lo), .dout(new_new_n3042__));
  buf1  g0365(.din(n3150_lo), .dout(new_new_n3044__));
  buf1  g0366(.din(n3153_lo), .dout(new_new_n3046__));
  buf1  g0367(.din(n3156_lo), .dout(new_new_n3048__));
  buf1  g0368(.din(n3159_lo), .dout(new_new_n3050__));
  buf1  g0369(.din(n3162_lo), .dout(new_new_n3052__));
  buf1  g0370(.din(n3165_lo), .dout(new_new_n3054__));
  buf1  g0371(.din(n3168_lo), .dout(new_new_n3056__));
  buf1  g0372(.din(n3171_lo), .dout(new_new_n3058__));
  buf1  g0373(.din(n3174_lo), .dout(new_new_n3060__));
  buf1  g0374(.din(n3177_lo), .dout(new_new_n3062__));
  buf1  g0375(.din(n3180_lo), .dout(new_new_n3064__));
  buf1  g0376(.din(n3183_lo), .dout(new_new_n3066__));
  buf1  g0377(.din(n3186_lo), .dout(new_new_n3068__));
  buf1  g0378(.din(n3189_lo), .dout(new_new_n3070__));
  buf1  g0379(.din(n3192_lo), .dout(new_new_n3072__));
  not1  g0380(.din(n3195_lo), .dout(new_new_n3075__));
  buf1  g0381(.din(n3198_lo), .dout(new_new_n3076__));
  buf1  g0382(.din(n3201_lo), .dout(new_new_n3078__));
  buf1  g0383(.din(n3204_lo), .dout(new_new_n3080__));
  buf1  g0384(.din(n3207_lo), .dout(new_new_n3082__));
  buf1  g0385(.din(n3210_lo), .dout(new_new_n3084__));
  buf1  g0386(.din(n3213_lo), .dout(new_new_n3086__));
  buf1  g0387(.din(n3216_lo), .dout(new_new_n3088__));
  not1  g0388(.din(n3219_lo), .dout(new_new_n3091__));
  buf1  g0389(.din(n3222_lo), .dout(new_new_n3092__));
  buf1  g0390(.din(n3225_lo), .dout(new_new_n3094__));
  buf1  g0391(.din(n3228_lo), .dout(new_new_n3096__));
  buf1  g0392(.din(n3231_lo), .dout(new_new_n3098__));
  buf1  g0393(.din(n3234_lo), .dout(new_new_n3100__));
  buf1  g0394(.din(n3237_lo), .dout(new_new_n3102__));
  buf1  g0395(.din(n3240_lo), .dout(new_new_n3104__));
  buf1  g0396(.din(n3243_lo), .dout(new_new_n3106__));
  buf1  g0397(.din(n3246_lo), .dout(new_new_n3108__));
  buf1  g0398(.din(n3249_lo), .dout(new_new_n3110__));
  buf1  g0399(.din(n3252_lo), .dout(new_new_n3112__));
  buf1  g0400(.din(n3255_lo), .dout(new_new_n3114__));
  buf1  g0401(.din(n3258_lo), .dout(new_new_n3116__));
  buf1  g0402(.din(n3261_lo), .dout(new_new_n3118__));
  buf1  g0403(.din(n3264_lo), .dout(new_new_n3120__));
  buf1  g0404(.din(n3267_lo), .dout(new_new_n3122__));
  buf1  g0405(.din(n3270_lo), .dout(new_new_n3124__));
  buf1  g0406(.din(n3273_lo), .dout(new_new_n3126__));
  buf1  g0407(.din(n3276_lo), .dout(new_new_n3128__));
  buf1  g0408(.din(n3279_lo), .dout(new_new_n3130__));
  buf1  g0409(.din(n3282_lo), .dout(new_new_n3132__));
  buf1  g0410(.din(n3285_lo), .dout(new_new_n3134__));
  buf1  g0411(.din(n3288_lo), .dout(new_new_n3136__));
  buf1  g0412(.din(n3291_lo), .dout(new_new_n3138__));
  buf1  g0413(.din(n3294_lo), .dout(new_new_n3140__));
  buf1  g0414(.din(n3297_lo), .dout(new_new_n3142__));
  buf1  g0415(.din(n3300_lo), .dout(new_new_n3144__));
  buf1  g0416(.din(n3303_lo), .dout(new_new_n3146__));
  buf1  g0417(.din(n3306_lo), .dout(new_new_n3148__));
  buf1  g0418(.din(n3309_lo), .dout(new_new_n3150__));
  buf1  g0419(.din(n3312_lo), .dout(new_new_n3152__));
  buf1  g0420(.din(n3315_lo), .dout(new_new_n3154__));
  buf1  g0421(.din(n3318_lo), .dout(new_new_n3156__));
  buf1  g0422(.din(n3321_lo), .dout(new_new_n3158__));
  buf1  g0423(.din(n3324_lo), .dout(new_new_n3160__));
  buf1  g0424(.din(n3327_lo), .dout(new_new_n3162__));
  buf1  g0425(.din(n3330_lo), .dout(new_new_n3164__));
  buf1  g0426(.din(n3333_lo), .dout(new_new_n3166__));
  buf1  g0427(.din(n3336_lo), .dout(new_new_n3168__));
  buf1  g0428(.din(n3339_lo), .dout(new_new_n3170__));
  not1  g0429(.din(n3339_lo), .dout(new_new_n3171__));
  buf1  g0430(.din(n3342_lo), .dout(new_new_n3172__));
  buf1  g0431(.din(n3345_lo), .dout(new_new_n3174__));
  buf1  g0432(.din(n3348_lo), .dout(new_new_n3176__));
  not1  g0433(.din(n3351_lo), .dout(new_new_n3179__));
  buf1  g0434(.din(n3354_lo), .dout(new_new_n3180__));
  buf1  g0435(.din(n3357_lo), .dout(new_new_n3182__));
  buf1  g0436(.din(n3360_lo), .dout(new_new_n3184__));
  buf1  g0437(.din(n3363_lo), .dout(new_new_n3186__));
  buf1  g0438(.din(n3366_lo), .dout(new_new_n3188__));
  buf1  g0439(.din(n3369_lo), .dout(new_new_n3190__));
  buf1  g0440(.din(n3372_lo), .dout(new_new_n3192__));
  buf1  g0441(.din(n3375_lo), .dout(new_new_n3194__));
  buf1  g0442(.din(n3378_lo), .dout(new_new_n3196__));
  buf1  g0443(.din(n3381_lo), .dout(new_new_n3198__));
  buf1  g0444(.din(n3384_lo), .dout(new_new_n3200__));
  not1  g0445(.din(n3387_lo), .dout(new_new_n3203__));
  buf1  g0446(.din(n3390_lo), .dout(new_new_n3204__));
  buf1  g0447(.din(n3393_lo), .dout(new_new_n3206__));
  buf1  g0448(.din(n3396_lo), .dout(new_new_n3208__));
  buf1  g0449(.din(n3399_lo), .dout(new_new_n3210__));
  not1  g0450(.din(n3399_lo), .dout(new_new_n3211__));
  buf1  g0451(.din(n3402_lo), .dout(new_new_n3212__));
  buf1  g0452(.din(n3405_lo), .dout(new_new_n3214__));
  buf1  g0453(.din(n3408_lo), .dout(new_new_n3216__));
  buf1  g0454(.din(n3411_lo), .dout(new_new_n3218__));
  buf1  g0455(.din(n3414_lo), .dout(new_new_n3220__));
  buf1  g0456(.din(n3417_lo), .dout(new_new_n3222__));
  buf1  g0457(.din(n3420_lo), .dout(new_new_n3224__));
  buf1  g0458(.din(n3423_lo), .dout(new_new_n3226__));
  buf1  g0459(.din(n3426_lo), .dout(new_new_n3228__));
  buf1  g0460(.din(n3429_lo), .dout(new_new_n3230__));
  buf1  g0461(.din(n3432_lo), .dout(new_new_n3232__));
  buf1  g0462(.din(n3435_lo), .dout(new_new_n3234__));
  buf1  g0463(.din(n3438_lo), .dout(new_new_n3236__));
  buf1  g0464(.din(n3441_lo), .dout(new_new_n3238__));
  buf1  g0465(.din(n3444_lo), .dout(new_new_n3240__));
  buf1  g0466(.din(n3447_lo), .dout(new_new_n3242__));
  buf1  g0467(.din(n3450_lo), .dout(new_new_n3244__));
  buf1  g0468(.din(n3453_lo), .dout(new_new_n3246__));
  buf1  g0469(.din(n3456_lo), .dout(new_new_n3248__));
  buf1  g0470(.din(n3459_lo), .dout(new_new_n3250__));
  buf1  g0471(.din(n3462_lo), .dout(new_new_n3252__));
  buf1  g0472(.din(n3465_lo), .dout(new_new_n3254__));
  buf1  g0473(.din(n3468_lo), .dout(new_new_n3256__));
  buf1  g0474(.din(n3471_lo), .dout(new_new_n3258__));
  buf1  g0475(.din(n3474_lo), .dout(new_new_n3260__));
  buf1  g0476(.din(n3477_lo), .dout(new_new_n3262__));
  buf1  g0477(.din(n3480_lo), .dout(new_new_n3264__));
  buf1  g0478(.din(n3483_lo), .dout(new_new_n3266__));
  buf1  g0479(.din(n3486_lo), .dout(new_new_n3268__));
  buf1  g0480(.din(n3489_lo), .dout(new_new_n3270__));
  buf1  g0481(.din(n3492_lo), .dout(new_new_n3272__));
  buf1  g0482(.din(n3495_lo), .dout(new_new_n3274__));
  buf1  g0483(.din(n3498_lo), .dout(new_new_n3276__));
  buf1  g0484(.din(n3501_lo), .dout(new_new_n3278__));
  buf1  g0485(.din(n3504_lo), .dout(new_new_n3280__));
  buf1  g0486(.din(n3507_lo), .dout(new_new_n3282__));
  buf1  g0487(.din(n3510_lo), .dout(new_new_n3284__));
  buf1  g0488(.din(n3513_lo), .dout(new_new_n3286__));
  buf1  g0489(.din(n3516_lo), .dout(new_new_n3288__));
  buf1  g0490(.din(n3519_lo), .dout(new_new_n3290__));
  buf1  g0491(.din(n3522_lo), .dout(new_new_n3292__));
  buf1  g0492(.din(n3525_lo), .dout(new_new_n3294__));
  buf1  g0493(.din(n3528_lo), .dout(new_new_n3296__));
  buf1  g0494(.din(n3531_lo), .dout(new_new_n3298__));
  buf1  g0495(.din(n3534_lo), .dout(new_new_n3300__));
  buf1  g0496(.din(n3537_lo), .dout(new_new_n3302__));
  buf1  g0497(.din(n3540_lo), .dout(new_new_n3304__));
  buf1  g0498(.din(n3543_lo), .dout(new_new_n3306__));
  buf1  g0499(.din(n3546_lo), .dout(new_new_n3308__));
  buf1  g0500(.din(n3549_lo), .dout(new_new_n3310__));
  buf1  g0501(.din(n3552_lo), .dout(new_new_n3312__));
  buf1  g0502(.din(n3555_lo), .dout(new_new_n3314__));
  buf1  g0503(.din(n3558_lo), .dout(new_new_n3316__));
  buf1  g0504(.din(n3561_lo), .dout(new_new_n3318__));
  buf1  g0505(.din(n3564_lo), .dout(new_new_n3320__));
  buf1  g0506(.din(n3567_lo), .dout(new_new_n3322__));
  buf1  g0507(.din(n3570_lo), .dout(new_new_n3324__));
  buf1  g0508(.din(n3573_lo), .dout(new_new_n3326__));
  buf1  g0509(.din(n3576_lo), .dout(new_new_n3328__));
  buf1  g0510(.din(n3579_lo), .dout(new_new_n3330__));
  buf1  g0511(.din(n3582_lo), .dout(new_new_n3332__));
  buf1  g0512(.din(n3585_lo), .dout(new_new_n3334__));
  buf1  g0513(.din(n3588_lo), .dout(new_new_n3336__));
  buf1  g0514(.din(n3591_lo), .dout(new_new_n3338__));
  buf1  g0515(.din(n3594_lo), .dout(new_new_n3340__));
  buf1  g0516(.din(n3597_lo), .dout(new_new_n3342__));
  buf1  g0517(.din(n3600_lo), .dout(new_new_n3344__));
  buf1  g0518(.din(n3603_lo), .dout(new_new_n3346__));
  buf1  g0519(.din(n3606_lo), .dout(new_new_n3348__));
  buf1  g0520(.din(n3609_lo), .dout(new_new_n3350__));
  buf1  g0521(.din(n3612_lo), .dout(new_new_n3352__));
  buf1  g0522(.din(n3615_lo), .dout(new_new_n3354__));
  buf1  g0523(.din(n3618_lo), .dout(new_new_n3356__));
  buf1  g0524(.din(n3621_lo), .dout(new_new_n3358__));
  buf1  g0525(.din(n3624_lo), .dout(new_new_n3360__));
  buf1  g0526(.din(n3627_lo), .dout(new_new_n3362__));
  buf1  g0527(.din(n3630_lo), .dout(new_new_n3364__));
  buf1  g0528(.din(n3633_lo), .dout(new_new_n3366__));
  buf1  g0529(.din(n3636_lo), .dout(new_new_n3368__));
  buf1  g0530(.din(n3639_lo), .dout(new_new_n3370__));
  buf1  g0531(.din(n3642_lo), .dout(new_new_n3372__));
  buf1  g0532(.din(n3645_lo), .dout(new_new_n3374__));
  buf1  g0533(.din(n3648_lo), .dout(new_new_n3376__));
  buf1  g0534(.din(n3651_lo), .dout(new_new_n3378__));
  buf1  g0535(.din(n3654_lo), .dout(new_new_n3380__));
  buf1  g0536(.din(n3657_lo), .dout(new_new_n3382__));
  buf1  g0537(.din(n3666_lo), .dout(new_new_n3384__));
  buf1  g0538(.din(n3669_lo), .dout(new_new_n3386__));
  buf1  g0539(.din(n3678_lo), .dout(new_new_n3388__));
  buf1  g0540(.din(n3687_lo), .dout(new_new_n3390__));
  not1  g0541(.din(n3687_lo), .dout(new_new_n3391__));
  buf1  g0542(.din(n3690_lo), .dout(new_new_n3392__));
  buf1  g0543(.din(n3702_lo), .dout(new_new_n3394__));
  not1  g0544(.din(n3702_lo), .dout(new_new_n3395__));
  buf1  g0545(.din(n3711_lo), .dout(new_new_n3396__));
  not1  g0546(.din(n3711_lo), .dout(new_new_n3397__));
  buf1  g0547(.din(n3714_lo), .dout(new_new_n3398__));
  not1  g0548(.din(n3714_lo), .dout(new_new_n3399__));
  buf1  g0549(.din(n3726_lo), .dout(new_new_n3400__));
  not1  g0550(.din(n3726_lo), .dout(new_new_n3401__));
  buf1  g0551(.din(n3735_lo), .dout(new_new_n3402__));
  not1  g0552(.din(n3735_lo), .dout(new_new_n3403__));
  buf1  g0553(.din(n3738_lo), .dout(new_new_n3404__));
  not1  g0554(.din(n3738_lo), .dout(new_new_n3405__));
  buf1  g0555(.din(n3750_lo), .dout(new_new_n3406__));
  buf1  g0556(.din(n3753_lo), .dout(new_new_n3408__));
  not1  g0557(.din(n3753_lo), .dout(new_new_n3409__));
  buf1  g0558(.din(n3759_lo), .dout(new_new_n3410__));
  not1  g0559(.din(n3759_lo), .dout(new_new_n3411__));
  buf1  g0560(.din(n3762_lo), .dout(new_new_n3412__));
  buf1  g0561(.din(n3765_lo), .dout(new_new_n3414__));
  not1  g0562(.din(n3765_lo), .dout(new_new_n3415__));
  buf1  g0563(.din(n3774_lo), .dout(new_new_n3416__));
  buf1  g0564(.din(n3777_lo), .dout(new_new_n3418__));
  buf1  g0565(.din(n3786_lo), .dout(new_new_n3420__));
  buf1  g0566(.din(n3789_lo), .dout(new_new_n3422__));
  buf1  g0567(.din(n3792_lo), .dout(new_new_n3424__));
  not1  g0568(.din(n3795_lo), .dout(new_new_n3427__));
  buf1  g0569(.din(n3798_lo), .dout(new_new_n3428__));
  buf1  g0570(.din(n3801_lo), .dout(new_new_n3430__));
  not1  g0571(.din(n3801_lo), .dout(new_new_n3431__));
  buf1  g0572(.din(n3810_lo), .dout(new_new_n3432__));
  buf1  g0573(.din(n3813_lo), .dout(new_new_n3434__));
  not1  g0574(.din(n3813_lo), .dout(new_new_n3435__));
  buf1  g0575(.din(n3822_lo), .dout(new_new_n3436__));
  buf1  g0576(.din(n3825_lo), .dout(new_new_n3438__));
  buf1  g0577(.din(n3834_lo), .dout(new_new_n3440__));
  not1  g0578(.din(n3834_lo), .dout(new_new_n3441__));
  buf1  g0579(.din(n3843_lo), .dout(new_new_n3442__));
  not1  g0580(.din(n3843_lo), .dout(new_new_n3443__));
  buf1  g0581(.din(n3846_lo), .dout(new_new_n3444__));
  not1  g0582(.din(n3846_lo), .dout(new_new_n3445__));
  buf1  g0583(.din(n3867_lo), .dout(new_new_n3446__));
  not1  g0584(.din(n3867_lo), .dout(new_new_n3447__));
  buf1  g0585(.din(n3891_lo), .dout(new_new_n3448__));
  not1  g0586(.din(n3891_lo), .dout(new_new_n3449__));
  buf1  g0587(.din(n3915_lo), .dout(new_new_n3450__));
  not1  g0588(.din(n3915_lo), .dout(new_new_n3451__));
  buf1  g0589(.din(n3930_lo), .dout(new_new_n3452__));
  buf1  g0590(.din(n3933_lo), .dout(new_new_n3454__));
  buf1  g0591(.din(n3936_lo), .dout(new_new_n3456__));
  not1  g0592(.din(n3936_lo), .dout(new_new_n3457__));
  buf1  g0593(.din(n3942_lo), .dout(new_new_n3458__));
  buf1  g0594(.din(n3945_lo), .dout(new_new_n3460__));
  buf1  g0595(.din(n3948_lo), .dout(new_new_n3462__));
  not1  g0596(.din(n3948_lo), .dout(new_new_n3463__));
  buf1  g0597(.din(n3954_lo), .dout(new_new_n3464__));
  buf1  g0598(.din(n3957_lo), .dout(new_new_n3466__));
  buf1  g0599(.din(n3963_lo), .dout(new_new_n3468__));
  not1  g0600(.din(n3963_lo), .dout(new_new_n3469__));
  buf1  g0601(.din(n3966_lo), .dout(new_new_n3470__));
  buf1  g0602(.din(n3969_lo), .dout(new_new_n3472__));
  buf1  g0603(.din(n3975_lo), .dout(new_new_n3474__));
  not1  g0604(.din(n3975_lo), .dout(new_new_n3475__));
  buf1  g0605(.din(n3978_lo), .dout(new_new_n3476__));
  buf1  g0606(.din(n3987_lo), .dout(new_new_n3478__));
  not1  g0607(.din(n3987_lo), .dout(new_new_n3479__));
  buf1  g0608(.din(n3990_lo), .dout(new_new_n3480__));
  buf1  g0609(.din(n4002_lo), .dout(new_new_n3482__));
  not1  g0610(.din(n4002_lo), .dout(new_new_n3483__));
  buf1  g0611(.din(n4011_lo), .dout(new_new_n3484__));
  not1  g0612(.din(n4011_lo), .dout(new_new_n3485__));
  buf1  g0613(.din(n4014_lo), .dout(new_new_n3486__));
  not1  g0614(.din(n4014_lo), .dout(new_new_n3487__));
  buf1  g0615(.din(n4026_lo), .dout(new_new_n3488__));
  not1  g0616(.din(n4026_lo), .dout(new_new_n3489__));
  buf1  g0617(.din(n4035_lo), .dout(new_new_n3490__));
  not1  g0618(.din(n4035_lo), .dout(new_new_n3491__));
  buf1  g0619(.din(n4038_lo), .dout(new_new_n3492__));
  not1  g0620(.din(n4038_lo), .dout(new_new_n3493__));
  buf1  g0621(.din(n4050_lo), .dout(new_new_n3494__));
  buf1  g0622(.din(n4053_lo), .dout(new_new_n3496__));
  not1  g0623(.din(n4053_lo), .dout(new_new_n3497__));
  buf1  g0624(.din(n4059_lo), .dout(new_new_n3498__));
  not1  g0625(.din(n4059_lo), .dout(new_new_n3499__));
  buf1  g0626(.din(n4062_lo), .dout(new_new_n3500__));
  buf1  g0627(.din(n4065_lo), .dout(new_new_n3502__));
  not1  g0628(.din(n4065_lo), .dout(new_new_n3503__));
  buf1  g0629(.din(n4098_lo), .dout(new_new_n3504__));
  not1  g0630(.din(n4098_lo), .dout(new_new_n3505__));
  not1  g0631(.din(n4107_lo), .dout(new_new_n3507__));
  buf1  g0632(.din(n4119_lo), .dout(new_new_n3508__));
  not1  g0633(.din(n4119_lo), .dout(new_new_n3509__));
  not1  g0634(.din(n4131_lo), .dout(new_new_n3511__));
  buf1  g0635(.din(n4143_lo), .dout(new_new_n3512__));
  not1  g0636(.din(n4143_lo), .dout(new_new_n3513__));
  not1  g0637(.din(n4155_lo), .dout(new_new_n3515__));
  buf1  g0638(.din(n4167_lo), .dout(new_new_n3516__));
  not1  g0639(.din(n4167_lo), .dout(new_new_n3517__));
  not1  g0640(.din(n4179_lo), .dout(new_new_n3519__));
  buf1  g0641(.din(n4182_lo), .dout(new_new_n3520__));
  buf1  g0642(.din(n4185_lo), .dout(new_new_n3522__));
  buf1  g0643(.din(n4188_lo), .dout(new_new_n3524__));
  not1  g0644(.din(n4188_lo), .dout(new_new_n3525__));
  buf1  g0645(.din(n4194_lo), .dout(new_new_n3526__));
  buf1  g0646(.din(n4197_lo), .dout(new_new_n3528__));
  buf1  g0647(.din(n4200_lo), .dout(new_new_n3530__));
  buf1  g0648(.din(n4206_lo), .dout(new_new_n3532__));
  buf1  g0649(.din(n4209_lo), .dout(new_new_n3534__));
  buf1  g0650(.din(n4212_lo), .dout(new_new_n3536__));
  buf1  g0651(.din(n4215_lo), .dout(new_new_n3538__));
  buf1  g0652(.din(n4227_lo), .dout(new_new_n3540__));
  not1  g0653(.din(n4227_lo), .dout(new_new_n3541__));
  buf1  g0654(.din(n4230_lo), .dout(new_new_n3542__));
  buf1  g0655(.din(n4233_lo), .dout(new_new_n3544__));
  buf1  g0656(.din(n4236_lo), .dout(new_new_n3546__));
  not1  g0657(.din(n4239_lo), .dout(new_new_n3549__));
  buf1  g0658(.din(n4242_lo), .dout(new_new_n3550__));
  not1  g0659(.din(n4242_lo), .dout(new_new_n3551__));
  buf1  g0660(.din(n4251_lo), .dout(new_new_n3552__));
  not1  g0661(.din(n4251_lo), .dout(new_new_n3553__));
  buf1  g0662(.din(n4263_lo), .dout(new_new_n3554__));
  not1  g0663(.din(n4263_lo), .dout(new_new_n3555__));
  buf1  g0664(.din(n4275_lo), .dout(new_new_n3556__));
  not1  g0665(.din(n4275_lo), .dout(new_new_n3557__));
  buf1  g0666(.din(n4278_lo), .dout(new_new_n3558__));
  not1  g0667(.din(n4278_lo), .dout(new_new_n3559__));
  buf1  g0668(.din(n4287_lo), .dout(new_new_n3560__));
  not1  g0669(.din(n4287_lo), .dout(new_new_n3561__));
  buf1  g0670(.din(n4290_lo), .dout(new_new_n3562__));
  buf1  g0671(.din(n4293_lo), .dout(new_new_n3564__));
  not1  g0672(.din(n4293_lo), .dout(new_new_n3565__));
  buf1  g0673(.din(n4299_lo), .dout(new_new_n3566__));
  not1  g0674(.din(n4299_lo), .dout(new_new_n3567__));
  buf1  g0675(.din(n4302_lo), .dout(new_new_n3568__));
  buf1  g0676(.din(n4305_lo), .dout(new_new_n3570__));
  not1  g0677(.din(n4305_lo), .dout(new_new_n3571__));
  buf1  g0678(.din(n4311_lo), .dout(new_new_n3572__));
  not1  g0679(.din(n4311_lo), .dout(new_new_n3573__));
  buf1  g0680(.din(n4314_lo), .dout(new_new_n3574__));
  buf1  g0681(.din(n4323_lo), .dout(new_new_n3576__));
  not1  g0682(.din(n4323_lo), .dout(new_new_n3577__));
  buf1  g0683(.din(n4326_lo), .dout(new_new_n3578__));
  not1  g0684(.din(n4326_lo), .dout(new_new_n3579__));
  buf1  g0685(.din(n4335_lo), .dout(new_new_n3580__));
  not1  g0686(.din(n4335_lo), .dout(new_new_n3581__));
  buf1  g0687(.din(n4338_lo), .dout(new_new_n3582__));
  not1  g0688(.din(n4338_lo), .dout(new_new_n3583__));
  buf1  g0689(.din(n4347_lo), .dout(new_new_n3584__));
  not1  g0690(.din(n4347_lo), .dout(new_new_n3585__));
  buf1  g0691(.din(n4350_lo), .dout(new_new_n3586__));
  not1  g0692(.din(n4350_lo), .dout(new_new_n3587__));
  buf1  g0693(.din(n4359_lo), .dout(new_new_n3588__));
  not1  g0694(.din(n4359_lo), .dout(new_new_n3589__));
  buf1  g0695(.din(n4362_lo), .dout(new_new_n3590__));
  buf1  g0696(.din(n4365_lo), .dout(new_new_n3592__));
  not1  g0697(.din(n4365_lo), .dout(new_new_n3593__));
  buf1  g0698(.din(n4371_lo), .dout(new_new_n3594__));
  not1  g0699(.din(n4371_lo), .dout(new_new_n3595__));
  buf1  g0700(.din(n4374_lo), .dout(new_new_n3596__));
  not1  g0701(.din(n4374_lo), .dout(new_new_n3597__));
  buf1  g0702(.din(n4383_lo), .dout(new_new_n3598__));
  not1  g0703(.din(n4383_lo), .dout(new_new_n3599__));
  buf1  g0704(.din(n4395_lo), .dout(new_new_n3600__));
  not1  g0705(.din(n4395_lo), .dout(new_new_n3601__));
  buf1  g0706(.din(n4407_lo), .dout(new_new_n3602__));
  not1  g0707(.din(n4407_lo), .dout(new_new_n3603__));
  buf1  g0708(.din(n4410_lo), .dout(new_new_n3604__));
  buf1  g0709(.din(n4413_lo), .dout(new_new_n3606__));
  buf1  g0710(.din(n4416_lo), .dout(new_new_n3608__));
  not1  g0711(.din(n4419_lo), .dout(new_new_n3611__));
  buf1  g0712(.din(n4422_lo), .dout(new_new_n3612__));
  buf1  g0713(.din(n4425_lo), .dout(new_new_n3614__));
  buf1  g0714(.din(n4428_lo), .dout(new_new_n3616__));
  buf1  g0715(.din(n4431_lo), .dout(new_new_n3618__));
  not1  g0716(.din(n4431_lo), .dout(new_new_n3619__));
  buf1  g0717(.din(n4434_lo), .dout(new_new_n3620__));
  buf1  g0718(.din(n4437_lo), .dout(new_new_n3622__));
  buf1  g0719(.din(n4440_lo), .dout(new_new_n3624__));
  buf1  g0720(.din(n4443_lo), .dout(new_new_n3626__));
  not1  g0721(.din(n4443_lo), .dout(new_new_n3627__));
  buf1  g0722(.din(n4446_lo), .dout(new_new_n3628__));
  buf1  g0723(.din(n4449_lo), .dout(new_new_n3630__));
  buf1  g0724(.din(n4452_lo), .dout(new_new_n3632__));
  not1  g0725(.din(n4455_lo), .dout(new_new_n3635__));
  buf1  g0726(.din(n4458_lo), .dout(new_new_n3636__));
  buf1  g0727(.din(n4461_lo), .dout(new_new_n3638__));
  buf1  g0728(.din(n4464_lo), .dout(new_new_n3640__));
  not1  g0729(.din(n4467_lo), .dout(new_new_n3643__));
  buf1  g0730(.din(n4470_lo), .dout(new_new_n3644__));
  buf1  g0731(.din(n4473_lo), .dout(new_new_n3646__));
  buf1  g0732(.din(n4476_lo), .dout(new_new_n3648__));
  buf1  g0733(.din(n4479_lo), .dout(new_new_n3650__));
  not1  g0734(.din(n4479_lo), .dout(new_new_n3651__));
  buf1  g0735(.din(n4482_lo), .dout(new_new_n3652__));
  buf1  g0736(.din(n4485_lo), .dout(new_new_n3654__));
  buf1  g0737(.din(n4488_lo), .dout(new_new_n3656__));
  not1  g0738(.din(n4488_lo), .dout(new_new_n3657__));
  buf1  g0739(.din(n4494_lo), .dout(new_new_n3658__));
  buf1  g0740(.din(n4497_lo), .dout(new_new_n3660__));
  buf1  g0741(.din(n4500_lo), .dout(new_new_n3662__));
  buf1  g0742(.din(n4503_lo), .dout(new_new_n3664__));
  not1  g0743(.din(n4503_lo), .dout(new_new_n3665__));
  buf1  g0744(.din(n4506_lo), .dout(new_new_n3666__));
  buf1  g0745(.din(n4509_lo), .dout(new_new_n3668__));
  buf1  g0746(.din(n4512_lo), .dout(new_new_n3670__));
  buf1  g0747(.din(n4515_lo), .dout(new_new_n3672__));
  not1  g0748(.din(n4515_lo), .dout(new_new_n3673__));
  buf1  g0749(.din(n4518_lo), .dout(new_new_n3674__));
  buf1  g0750(.din(n4521_lo), .dout(new_new_n3676__));
  buf1  g0751(.din(n4524_lo), .dout(new_new_n3678__));
  buf1  g0752(.din(n4527_lo), .dout(new_new_n3680__));
  not1  g0753(.din(n4527_lo), .dout(new_new_n3681__));
  buf1  g0754(.din(n4530_lo), .dout(new_new_n3682__));
  buf1  g0755(.din(n4533_lo), .dout(new_new_n3684__));
  buf1  g0756(.din(n4536_lo), .dout(new_new_n3686__));
  buf1  g0757(.din(n4539_lo), .dout(new_new_n3688__));
  not1  g0758(.din(n4539_lo), .dout(new_new_n3689__));
  buf1  g0759(.din(n4542_lo), .dout(new_new_n3690__));
  buf1  g0760(.din(n4545_lo), .dout(new_new_n3692__));
  buf1  g0761(.din(n4548_lo), .dout(new_new_n3694__));
  not1  g0762(.din(n4548_lo), .dout(new_new_n3695__));
  buf1  g0763(.din(n4554_lo), .dout(new_new_n3696__));
  buf1  g0764(.din(n4557_lo), .dout(new_new_n3698__));
  buf1  g0765(.din(n4560_lo), .dout(new_new_n3700__));
  buf1  g0766(.din(n4563_lo), .dout(new_new_n3702__));
  not1  g0767(.din(n4563_lo), .dout(new_new_n3703__));
  buf1  g0768(.din(n4566_lo), .dout(new_new_n3704__));
  buf1  g0769(.din(n4569_lo), .dout(new_new_n3706__));
  buf1  g0770(.din(n4572_lo), .dout(new_new_n3708__));
  buf1  g0771(.din(n4575_lo), .dout(new_new_n3710__));
  buf1  g0772(.din(n4578_lo), .dout(new_new_n3712__));
  buf1  g0773(.din(n4581_lo), .dout(new_new_n3714__));
  buf1  g0774(.din(n4584_lo), .dout(new_new_n3716__));
  not1  g0775(.din(n4587_lo), .dout(new_new_n3719__));
  buf1  g0776(.din(n4590_lo), .dout(new_new_n3720__));
  buf1  g0777(.din(n4593_lo), .dout(new_new_n3722__));
  buf1  g0778(.din(n4596_lo), .dout(new_new_n3724__));
  not1  g0779(.din(n4599_lo), .dout(new_new_n3727__));
  buf1  g0780(.din(n4602_lo), .dout(new_new_n3728__));
  buf1  g0781(.din(n4605_lo), .dout(new_new_n3730__));
  buf1  g0782(.din(n4608_lo), .dout(new_new_n3732__));
  not1  g0783(.din(n4611_lo), .dout(new_new_n3735__));
  buf1  g0784(.din(n4614_lo), .dout(new_new_n3736__));
  buf1  g0785(.din(n4617_lo), .dout(new_new_n3738__));
  buf1  g0786(.din(n4620_lo), .dout(new_new_n3740__));
  buf1  g0787(.din(n4623_lo), .dout(new_new_n3742__));
  buf1  g0788(.din(n4626_lo), .dout(new_new_n3744__));
  buf1  g0789(.din(n4629_lo), .dout(new_new_n3746__));
  buf1  g0790(.din(n4632_lo), .dout(new_new_n3748__));
  buf1  g0791(.din(n4635_lo), .dout(new_new_n3750__));
  buf1  g0792(.din(n4638_lo), .dout(new_new_n3752__));
  buf1  g0793(.din(n4641_lo), .dout(new_new_n3754__));
  buf1  g0794(.din(n4644_lo), .dout(new_new_n3756__));
  buf1  g0795(.din(n4647_lo), .dout(new_new_n3758__));
  not1  g0796(.din(n4647_lo), .dout(new_new_n3759__));
  buf1  g0797(.din(n4650_lo), .dout(new_new_n3760__));
  buf1  g0798(.din(n4653_lo), .dout(new_new_n3762__));
  buf1  g0799(.din(n4656_lo), .dout(new_new_n3764__));
  buf1  g0800(.din(n4659_lo), .dout(new_new_n3766__));
  not1  g0801(.din(n4659_lo), .dout(new_new_n3767__));
  buf1  g0802(.din(n4662_lo), .dout(new_new_n3768__));
  buf1  g0803(.din(n4665_lo), .dout(new_new_n3770__));
  buf1  g0804(.din(n4668_lo), .dout(new_new_n3772__));
  buf1  g0805(.din(n4671_lo), .dout(new_new_n3774__));
  not1  g0806(.din(n4671_lo), .dout(new_new_n3775__));
  buf1  g0807(.din(n4674_lo), .dout(new_new_n3776__));
  buf1  g0808(.din(n4677_lo), .dout(new_new_n3778__));
  buf1  g0809(.din(n4680_lo), .dout(new_new_n3780__));
  buf1  g0810(.din(n4683_lo), .dout(new_new_n3782__));
  not1  g0811(.din(n4683_lo), .dout(new_new_n3783__));
  buf1  g0812(.din(n4686_lo), .dout(new_new_n3784__));
  buf1  g0813(.din(n4689_lo), .dout(new_new_n3786__));
  buf1  g0814(.din(n4692_lo), .dout(new_new_n3788__));
  buf1  g0815(.din(n4695_lo), .dout(new_new_n3790__));
  not1  g0816(.din(n4695_lo), .dout(new_new_n3791__));
  buf1  g0817(.din(n4698_lo), .dout(new_new_n3792__));
  buf1  g0818(.din(n4701_lo), .dout(new_new_n3794__));
  buf1  g0819(.din(n4704_lo), .dout(new_new_n3796__));
  buf1  g0820(.din(n4707_lo), .dout(new_new_n3798__));
  not1  g0821(.din(n4707_lo), .dout(new_new_n3799__));
  buf1  g0822(.din(n4710_lo), .dout(new_new_n3800__));
  buf1  g0823(.din(n4713_lo), .dout(new_new_n3802__));
  buf1  g0824(.din(n4716_lo), .dout(new_new_n3804__));
  buf1  g0825(.din(n4719_lo), .dout(new_new_n3806__));
  not1  g0826(.din(n4719_lo), .dout(new_new_n3807__));
  buf1  g0827(.din(n4722_lo), .dout(new_new_n3808__));
  buf1  g0828(.din(n4725_lo), .dout(new_new_n3810__));
  buf1  g0829(.din(n4728_lo), .dout(new_new_n3812__));
  buf1  g0830(.din(n4731_lo), .dout(new_new_n3814__));
  not1  g0831(.din(n4731_lo), .dout(new_new_n3815__));
  buf1  g0832(.din(n4734_lo), .dout(new_new_n3816__));
  buf1  g0833(.din(n4737_lo), .dout(new_new_n3818__));
  buf1  g0834(.din(n4740_lo), .dout(new_new_n3820__));
  not1  g0835(.din(n4743_lo), .dout(new_new_n3823__));
  not1  g0836(.din(n6382_o2), .dout(new_new_n3825__));
  not1  g0837(.din(n6383_o2), .dout(new_new_n3827__));
  not1  g0838(.din(n6419_o2), .dout(new_new_n3829__));
  not1  g0839(.din(n6420_o2), .dout(new_new_n3831__));
  not1  g0840(.din(n6435_o2), .dout(new_new_n3833__));
  not1  g0841(.din(n6436_o2), .dout(new_new_n3835__));
  not1  g0842(.din(n6448_o2), .dout(new_new_n3837__));
  not1  g0843(.din(n6449_o2), .dout(new_new_n3839__));
  not1  g0844(.din(n6613_o2), .dout(new_new_n3841__));
  buf1  g0845(.din(n6614_o2), .dout(new_new_n3842__));
  not1  g0846(.din(n6641_o2), .dout(new_new_n3845__));
  buf1  g0847(.din(n6658_o2), .dout(new_new_n3846__));
  buf1  g0848(.din(n6757_o2), .dout(new_new_n3848__));
  not1  g0849(.din(n6757_o2), .dout(new_new_n3849__));
  buf1  g0850(.din(n6756_o2), .dout(new_new_n3850__));
  not1  g0851(.din(n6756_o2), .dout(new_new_n3851__));
  not1  g0852(.din(n7116_o2), .dout(new_new_n3853__));
  buf1  g0853(.din(n7156_o2), .dout(new_new_n3854__));
  not1  g0854(.din(n7156_o2), .dout(new_new_n3855__));
  not1  g0855(.din(n6549_o2), .dout(new_new_n3857__));
  buf1  g0856(.din(n6550_o2), .dout(new_new_n3858__));
  not1  g0857(.din(n6550_o2), .dout(new_new_n3859__));
  buf1  g0858(.din(n7357_o2), .dout(new_new_n3860__));
  buf1  g0859(.din(n7358_o2), .dout(new_new_n3862__));
  buf1  g0860(.din(n7359_o2), .dout(new_new_n3864__));
  buf1  g0861(.din(n7360_o2), .dout(new_new_n3866__));
  buf1  g0862(.din(n6621_o2), .dout(new_new_n3868__));
  not1  g0863(.din(n6621_o2), .dout(new_new_n3869__));
  buf1  g0864(.din(n6623_o2), .dout(new_new_n3870__));
  not1  g0865(.din(n6623_o2), .dout(new_new_n3871__));
  buf1  g0866(.din(n6625_o2), .dout(new_new_n3872__));
  not1  g0867(.din(n6625_o2), .dout(new_new_n3873__));
  buf1  g0868(.din(n6626_o2), .dout(new_new_n3874__));
  buf1  g0869(.din(n6627_o2), .dout(new_new_n3876__));
  not1  g0870(.din(n6627_o2), .dout(new_new_n3877__));
  buf1  g0871(.din(n6628_o2), .dout(new_new_n3878__));
  buf1  g0872(.din(n6629_o2), .dout(new_new_n3880__));
  buf1  g0873(.din(n6630_o2), .dout(new_new_n3882__));
  not1  g0874(.din(n6630_o2), .dout(new_new_n3883__));
  buf1  g0875(.din(n6669_o2), .dout(new_new_n3884__));
  not1  g0876(.din(n6669_o2), .dout(new_new_n3885__));
  buf1  g0877(.din(n7449_o2), .dout(new_new_n3886__));
  not1  g0878(.din(n7449_o2), .dout(new_new_n3887__));
  not1  g0879(.din(n7450_o2), .dout(new_new_n3889__));
  not1  g0880(.din(n7451_o2), .dout(new_new_n3891__));
  buf1  g0881(.din(n7452_o2), .dout(new_new_n3892__));
  not1  g0882(.din(n7452_o2), .dout(new_new_n3893__));
  buf1  g0883(.din(n6682_o2), .dout(new_new_n3894__));
  not1  g0884(.din(n6682_o2), .dout(new_new_n3895__));
  buf1  g0885(.din(n6683_o2), .dout(new_new_n3896__));
  not1  g0886(.din(n6683_o2), .dout(new_new_n3897__));
  buf1  g0887(.din(n6684_o2), .dout(new_new_n3898__));
  not1  g0888(.din(n6684_o2), .dout(new_new_n3899__));
  buf1  g0889(.din(n6685_o2), .dout(new_new_n3900__));
  not1  g0890(.din(n6685_o2), .dout(new_new_n3901__));
  buf1  g0891(.din(n7463_o2), .dout(new_new_n3902__));
  not1  g0892(.din(n7463_o2), .dout(new_new_n3903__));
  buf1  g0893(.din(n6686_o2), .dout(new_new_n3904__));
  not1  g0894(.din(n6686_o2), .dout(new_new_n3905__));
  buf1  g0895(.din(n6687_o2), .dout(new_new_n3906__));
  not1  g0896(.din(n6687_o2), .dout(new_new_n3907__));
  buf1  g0897(.din(n6688_o2), .dout(new_new_n3908__));
  not1  g0898(.din(n6688_o2), .dout(new_new_n3909__));
  buf1  g0899(.din(n6689_o2), .dout(new_new_n3910__));
  not1  g0900(.din(n6689_o2), .dout(new_new_n3911__));
  buf1  g0901(.din(n6772_o2), .dout(new_new_n3912__));
  not1  g0902(.din(n6772_o2), .dout(new_new_n3913__));
  buf1  g0903(.din(n6773_o2), .dout(new_new_n3914__));
  buf1  g0904(.din(n6774_o2), .dout(new_new_n3916__));
  not1  g0905(.din(n6774_o2), .dout(new_new_n3917__));
  buf1  g0906(.din(n6775_o2), .dout(new_new_n3918__));
  not1  g0907(.din(n6775_o2), .dout(new_new_n3919__));
  not1  g0908(.din(G3467_o2), .dout(new_new_n3921__));
  buf1  g0909(.din(G2810_o2), .dout(new_new_n3922__));
  buf1  g0910(.din(n6833_o2), .dout(new_new_n3924__));
  buf1  g0911(.din(n6945_o2), .dout(new_new_n3926__));
  not1  g0912(.din(n6945_o2), .dout(new_new_n3927__));
  buf1  g0913(.din(n6947_o2), .dout(new_new_n3928__));
  not1  g0914(.din(n6947_o2), .dout(new_new_n3929__));
  buf1  g0915(.din(n6949_o2), .dout(new_new_n3930__));
  not1  g0916(.din(n6949_o2), .dout(new_new_n3931__));
  buf1  g0917(.din(n6951_o2), .dout(new_new_n3932__));
  buf1  g0918(.din(n6888_o2), .dout(new_new_n3934__));
  not1  g0919(.din(n6888_o2), .dout(new_new_n3935__));
  buf1  g0920(.din(n6889_o2), .dout(new_new_n3936__));
  not1  g0921(.din(n6889_o2), .dout(new_new_n3937__));
  buf1  g0922(.din(n6936_o2), .dout(new_new_n3938__));
  not1  g0923(.din(n6936_o2), .dout(new_new_n3939__));
  buf1  g0924(.din(n6954_o2), .dout(new_new_n3940__));
  not1  g0925(.din(n6954_o2), .dout(new_new_n3941__));
  buf1  g0926(.din(n6955_o2), .dout(new_new_n3942__));
  not1  g0927(.din(n6955_o2), .dout(new_new_n3943__));
  buf1  g0928(.din(n6956_o2), .dout(new_new_n3944__));
  not1  g0929(.din(n6956_o2), .dout(new_new_n3945__));
  buf1  g0930(.din(n6957_o2), .dout(new_new_n3946__));
  not1  g0931(.din(n6957_o2), .dout(new_new_n3947__));
  buf1  g0932(.din(n6958_o2), .dout(new_new_n3948__));
  not1  g0933(.din(n6958_o2), .dout(new_new_n3949__));
  buf1  g0934(.din(n6982_o2), .dout(new_new_n3950__));
  not1  g0935(.din(n6982_o2), .dout(new_new_n3951__));
  buf1  g0936(.din(n6984_o2), .dout(new_new_n3952__));
  not1  g0937(.din(n6984_o2), .dout(new_new_n3953__));
  buf1  g0938(.din(n6974_o2), .dout(new_new_n3954__));
  not1  g0939(.din(n6974_o2), .dout(new_new_n3955__));
  buf1  g0940(.din(n6975_o2), .dout(new_new_n3956__));
  not1  g0941(.din(n6975_o2), .dout(new_new_n3957__));
  buf1  g0942(.din(n6999_o2), .dout(new_new_n3958__));
  not1  g0943(.din(n6999_o2), .dout(new_new_n3959__));
  buf1  g0944(.din(n7015_o2), .dout(new_new_n3960__));
  not1  g0945(.din(n7015_o2), .dout(new_new_n3961__));
  buf1  g0946(.din(n7016_o2), .dout(new_new_n3962__));
  not1  g0947(.din(n7016_o2), .dout(new_new_n3963__));
  buf1  g0948(.din(n7017_o2), .dout(new_new_n3964__));
  not1  g0949(.din(n7017_o2), .dout(new_new_n3965__));
  buf1  g0950(.din(n7018_o2), .dout(new_new_n3966__));
  not1  g0951(.din(n7018_o2), .dout(new_new_n3967__));
  buf1  g0952(.din(n7005_o2), .dout(new_new_n3968__));
  not1  g0953(.din(n7005_o2), .dout(new_new_n3969__));
  buf1  g0954(.din(n7019_o2), .dout(new_new_n3970__));
  not1  g0955(.din(n7019_o2), .dout(new_new_n3971__));
  buf1  g0956(.din(n7022_o2), .dout(new_new_n3972__));
  not1  g0957(.din(n7022_o2), .dout(new_new_n3973__));
  buf1  g0958(.din(n7023_o2), .dout(new_new_n3974__));
  not1  g0959(.din(n7023_o2), .dout(new_new_n3975__));
  buf1  g0960(.din(n7132_o2), .dout(new_new_n3976__));
  not1  g0961(.din(n7132_o2), .dout(new_new_n3977__));
  buf1  g0962(.din(n7133_o2), .dout(new_new_n3978__));
  not1  g0963(.din(n7133_o2), .dout(new_new_n3979__));
  buf1  g0964(.din(n7135_o2), .dout(new_new_n3980__));
  not1  g0965(.din(n7135_o2), .dout(new_new_n3981__));
  buf1  g0966(.din(n7136_o2), .dout(new_new_n3982__));
  not1  g0967(.din(n7136_o2), .dout(new_new_n3983__));
  buf1  g0968(.din(n7175_o2), .dout(new_new_n3984__));
  not1  g0969(.din(n7175_o2), .dout(new_new_n3985__));
  buf1  g0970(.din(n7155_o2), .dout(new_new_n3986__));
  not1  g0971(.din(n7155_o2), .dout(new_new_n3987__));
  not1  g0972(.din(G3060_o2), .dout(new_new_n3989__));
  buf1  g0973(.din(n7383_o2), .dout(new_new_n3990__));
  not1  g0974(.din(n7383_o2), .dout(new_new_n3991__));
  not1  g0975(.din(G3802_o2), .dout(new_new_n3993__));
  not1  g0976(.din(G3859_o2), .dout(new_new_n3995__));
  buf1  g0977(.din(n7355_o2), .dout(new_new_n3996__));
  buf1  g0978(.din(n7356_o2), .dout(new_new_n3998__));
  not1  g0979(.din(G4054_o2), .dout(new_new_n4001__));
  not1  g0980(.din(G4068_o2), .dout(new_new_n4003__));
  buf1  g0981(.din(n7384_o2), .dout(new_new_n4004__));
  not1  g0982(.din(n7384_o2), .dout(new_new_n4005__));
  buf1  g0983(.din(n7387_o2), .dout(new_new_n4006__));
  not1  g0984(.din(n7387_o2), .dout(new_new_n4007__));
  buf1  g0985(.din(n7388_o2), .dout(new_new_n4008__));
  buf1  g0986(.din(n7389_o2), .dout(new_new_n4010__));
  buf1  g0987(.din(n7386_o2), .dout(new_new_n4012__));
  not1  g0988(.din(n7386_o2), .dout(new_new_n4013__));
  buf1  g0989(.din(n7453_o2), .dout(new_new_n4014__));
  not1  g0990(.din(n7453_o2), .dout(new_new_n4015__));
  buf1  g0991(.din(n7431_o2), .dout(new_new_n4016__));
  not1  g0992(.din(n7431_o2), .dout(new_new_n4017__));
  buf1  g0993(.din(n7432_o2), .dout(new_new_n4018__));
  buf1  g0994(.din(n7433_o2), .dout(new_new_n4020__));
  buf1  g0995(.din(n7430_o2), .dout(new_new_n4022__));
  not1  g0996(.din(n7430_o2), .dout(new_new_n4023__));
  buf1  g0997(.din(n7485_o2), .dout(new_new_n4024__));
  buf1  g0998(.din(n7486_o2), .dout(new_new_n4026__));
  buf1  g0999(.din(G2508_o2), .dout(new_new_n4028__));
  buf1  g1000(.din(G2486_o2), .dout(new_new_n4030__));
  not1  g1001(.din(G2486_o2), .dout(new_new_n4031__));
  buf1  g1002(.din(n2326_inv), .dout(new_new_n4032__));
  buf1  g1003(.din(n2329_inv), .dout(new_new_n4034__));
  buf1  g1004(.din(n3756_lo_buf_o2), .dout(new_new_n4036__));
  not1  g1005(.din(n3756_lo_buf_o2), .dout(new_new_n4037__));
  buf1  g1006(.din(n4056_lo_buf_o2), .dout(new_new_n4038__));
  buf1  g1007(.din(G3474_o2), .dout(new_new_n4040__));
  not1  g1008(.din(G3474_o2), .dout(new_new_n4041__));
  buf1  g1009(.din(n2341_inv), .dout(new_new_n4042__));
  not1  g1010(.din(n2341_inv), .dout(new_new_n4043__));
  buf1  g1011(.din(n7396_o2), .dout(new_new_n4044__));
  buf1  g1012(.din(n7398_o2), .dout(new_new_n4046__));
  buf1  g1013(.din(n7400_o2), .dout(new_new_n4048__));
  buf1  g1014(.din(n7401_o2), .dout(new_new_n4050__));
  buf1  g1015(.din(n7402_o2), .dout(new_new_n4052__));
  buf1  g1016(.din(n7403_o2), .dout(new_new_n4054__));
  buf1  g1017(.din(n7404_o2), .dout(new_new_n4056__));
  buf1  g1018(.din(n7405_o2), .dout(new_new_n4058__));
  buf1  g1019(.din(G2711_o2), .dout(new_new_n4060__));
  buf1  g1020(.din(n2371_inv), .dout(new_new_n4062__));
  buf1  g1021(.din(n7490_o2), .dout(new_new_n4064__));
  buf1  g1022(.din(n7527_o2), .dout(new_new_n4066__));
  buf1  g1023(.din(n7528_o2), .dout(new_new_n4068__));
  buf1  g1024(.din(n7529_o2), .dout(new_new_n4070__));
  buf1  g1025(.din(n7530_o2), .dout(new_new_n4072__));
  buf1  g1026(.din(n7523_o2), .dout(new_new_n4074__));
  buf1  g1027(.din(n7524_o2), .dout(new_new_n4076__));
  buf1  g1028(.din(n7525_o2), .dout(new_new_n4078__));
  buf1  g1029(.din(n7526_o2), .dout(new_new_n4080__));
  buf1  g1030(.din(n4296_lo_buf_o2), .dout(new_new_n4082__));
  not1  g1031(.din(n4296_lo_buf_o2), .dout(new_new_n4083__));
  buf1  g1032(.din(n4368_lo_buf_o2), .dout(new_new_n4084__));
  not1  g1033(.din(n4368_lo_buf_o2), .dout(new_new_n4085__));
  buf1  g1034(.din(G2466_o2), .dout(new_new_n4086__));
  not1  g1035(.din(G2466_o2), .dout(new_new_n4087__));
  buf1  g1036(.din(G2404_o2), .dout(new_new_n4088__));
  not1  g1037(.din(G2404_o2), .dout(new_new_n4089__));
  buf1  g1038(.din(n7534_o2), .dout(new_new_n4090__));
  buf1  g1039(.din(n7535_o2), .dout(new_new_n4092__));
  buf1  g1040(.din(n7536_o2), .dout(new_new_n4094__));
  buf1  g1041(.din(n7533_o2), .dout(new_new_n4096__));
  buf1  g1042(.din(G1060_o2), .dout(new_new_n4098__));
  not1  g1043(.din(G1060_o2), .dout(new_new_n4099__));
  buf1  g1044(.din(G963_o2), .dout(new_new_n4100__));
  not1  g1045(.din(G963_o2), .dout(new_new_n4101__));
  buf1  g1046(.din(G2448_o2), .dout(new_new_n4102__));
  buf1  g1047(.din(G2685_o2), .dout(new_new_n4104__));
  not1  g1048(.din(G2685_o2), .dout(new_new_n4105__));
  buf1  g1049(.din(G2679_o2), .dout(new_new_n4106__));
  not1  g1050(.din(G2679_o2), .dout(new_new_n4107__));
  buf1  g1051(.din(G2774_o2), .dout(new_new_n4108__));
  not1  g1052(.din(G2774_o2), .dout(new_new_n4109__));
  buf1  g1053(.din(G2780_o2), .dout(new_new_n4110__));
  not1  g1054(.din(G2780_o2), .dout(new_new_n4111__));
  buf1  g1055(.din(G2759_o2), .dout(new_new_n4112__));
  not1  g1056(.din(G2759_o2), .dout(new_new_n4113__));
  buf1  g1057(.din(G2737_o2), .dout(new_new_n4114__));
  buf1  g1058(.din(G2850_o2), .dout(new_new_n4116__));
  buf1  g1059(.din(G3393_o2), .dout(new_new_n4118__));
  not1  g1060(.din(G3393_o2), .dout(new_new_n4119__));
  buf1  g1061(.din(G3404_o2), .dout(new_new_n4120__));
  not1  g1062(.din(G3404_o2), .dout(new_new_n4121__));
  buf1  g1063(.din(G3559_o2), .dout(new_new_n4122__));
  not1  g1064(.din(G3559_o2), .dout(new_new_n4123__));
  buf1  g1065(.din(G2744_o2), .dout(new_new_n4124__));
  buf1  g1066(.din(n3708_lo_buf_o2), .dout(new_new_n4126__));
  buf1  g1067(.din(n3840_lo_buf_o2), .dout(new_new_n4128__));
  not1  g1068(.din(n3840_lo_buf_o2), .dout(new_new_n4129__));
  buf1  g1069(.din(n4008_lo_buf_o2), .dout(new_new_n4130__));
  buf1  g1070(.din(n4104_lo_buf_o2), .dout(new_new_n4132__));
  buf1  g1071(.din(G1821_o2), .dout(new_new_n4134__));
  not1  g1072(.din(G1821_o2), .dout(new_new_n4135__));
  buf1  g1073(.din(G1734_o2), .dout(new_new_n4136__));
  not1  g1074(.din(G1734_o2), .dout(new_new_n4137__));
  buf1  g1075(.din(G3517_o2), .dout(new_new_n4138__));
  buf1  g1076(.din(G3533_o2), .dout(new_new_n4140__));
  not1  g1077(.din(G3533_o2), .dout(new_new_n4141__));
  buf1  g1078(.din(G3629_o2), .dout(new_new_n4142__));
  buf1  g1079(.din(G3645_o2), .dout(new_new_n4144__));
  not1  g1080(.din(G3645_o2), .dout(new_new_n4145__));
  buf1  g1081(.din(n2497_inv), .dout(new_new_n4146__));
  buf1  g1082(.din(G2731_o2), .dout(new_new_n4148__));
  buf1  g1083(.din(G2844_o2), .dout(new_new_n4150__));
  buf1  g1084(.din(n3732_lo_buf_o2), .dout(new_new_n4152__));
  buf1  g1085(.din(n4032_lo_buf_o2), .dout(new_new_n4154__));
  buf1  g1086(.din(G3552_o2), .dout(new_new_n4156__));
  not1  g1087(.din(G3552_o2), .dout(new_new_n4157__));
  buf1  g1088(.din(G2271_o2), .dout(new_new_n4158__));
  buf1  g1089(.din(n4248_lo_buf_o2), .dout(new_new_n4160__));
  buf1  g1090(.din(n4332_lo_buf_o2), .dout(new_new_n4162__));
  buf1  g1091(.din(n4344_lo_buf_o2), .dout(new_new_n4164__));
  buf1  g1092(.din(n4380_lo_buf_o2), .dout(new_new_n4166__));
  buf1  g1093(.din(G2398_o2), .dout(new_new_n4168__));
  buf1  g1094(.din(G2480_o2), .dout(new_new_n4170__));
  buf1  g1095(.din(G2418_o2), .dout(new_new_n4172__));
  buf1  g1096(.din(G1455_o2), .dout(new_new_n4174__));
  not1  g1097(.din(G1455_o2), .dout(new_new_n4175__));
  buf1  g1098(.din(G1449_o2), .dout(new_new_n4176__));
  not1  g1099(.din(G1449_o2), .dout(new_new_n4177__));
  buf1  g1100(.din(G1452_o2), .dout(new_new_n4178__));
  not1  g1101(.din(G1452_o2), .dout(new_new_n4179__));
  buf1  g1102(.din(G1425_o2), .dout(new_new_n4180__));
  not1  g1103(.din(G1425_o2), .dout(new_new_n4181__));
  buf1  g1104(.din(G1428_o2), .dout(new_new_n4182__));
  not1  g1105(.din(G1428_o2), .dout(new_new_n4183__));
  buf1  g1106(.din(G1419_o2), .dout(new_new_n4184__));
  not1  g1107(.din(G1419_o2), .dout(new_new_n4185__));
  buf1  g1108(.din(G1422_o2), .dout(new_new_n4186__));
  not1  g1109(.din(G1422_o2), .dout(new_new_n4187__));
  buf1  g1110(.din(n4308_lo_buf_o2), .dout(new_new_n4188__));
  not1  g1111(.din(n4308_lo_buf_o2), .dout(new_new_n4189__));
  buf1  g1112(.din(G2675_o2), .dout(new_new_n4190__));
  not1  g1113(.din(G2675_o2), .dout(new_new_n4191__));
  buf1  g1114(.din(G3035_o2), .dout(new_new_n4192__));
  not1  g1115(.din(G3035_o2), .dout(new_new_n4193__));
  buf1  g1116(.din(G3026_o2), .dout(new_new_n4194__));
  not1  g1117(.din(G3026_o2), .dout(new_new_n4195__));
  buf1  g1118(.din(G3029_o2), .dout(new_new_n4196__));
  not1  g1119(.din(G3029_o2), .dout(new_new_n4197__));
  buf1  g1120(.din(G3032_o2), .dout(new_new_n4198__));
  not1  g1121(.din(G3032_o2), .dout(new_new_n4199__));
  buf1  g1122(.din(G2999_o2), .dout(new_new_n4200__));
  not1  g1123(.din(G2999_o2), .dout(new_new_n4201__));
  buf1  g1124(.din(G3002_o2), .dout(new_new_n4202__));
  not1  g1125(.din(G3002_o2), .dout(new_new_n4203__));
  buf1  g1126(.din(G2770_o2), .dout(new_new_n4204__));
  not1  g1127(.din(G2770_o2), .dout(new_new_n4205__));
  buf1  g1128(.din(G3008_o2), .dout(new_new_n4206__));
  not1  g1129(.din(G3008_o2), .dout(new_new_n4207__));
  buf1  g1130(.din(G2073_o2), .dout(new_new_n4208__));
  not1  g1131(.din(G2073_o2), .dout(new_new_n4209__));
  buf1  g1132(.din(G2752_o2), .dout(new_new_n4210__));
  not1  g1133(.din(G2752_o2), .dout(new_new_n4211__));
  buf1  g1134(.din(G3005_o2), .dout(new_new_n4212__));
  not1  g1135(.din(G3005_o2), .dout(new_new_n4213__));
  buf1  g1136(.din(G5108_o2), .dout(new_new_n4214__));
  not1  g1137(.din(G5135_o2), .dout(new_new_n4217__));
  not1  g1138(.din(G5111_o2), .dout(new_new_n4219__));
  not1  g1139(.din(G5138_o2), .dout(new_new_n4221__));
  buf1  g1140(.din(G3415_o2), .dout(new_new_n4222__));
  not1  g1141(.din(G3415_o2), .dout(new_new_n4223__));
  buf1  g1142(.din(G3386_o2), .dout(new_new_n4224__));
  not1  g1143(.din(G3386_o2), .dout(new_new_n4225__));
  buf1  g1144(.din(G3570_o2), .dout(new_new_n4226__));
  not1  g1145(.din(G3570_o2), .dout(new_new_n4227__));
  buf1  g1146(.din(G2430_o2), .dout(new_new_n4228__));
  not1  g1147(.din(G2430_o2), .dout(new_new_n4229__));
  buf1  g1148(.din(G3495_o2), .dout(new_new_n4230__));
  not1  g1149(.din(G3495_o2), .dout(new_new_n4231__));
  buf1  g1150(.din(G3621_o2), .dout(new_new_n4232__));
  not1  g1151(.din(G3621_o2), .dout(new_new_n4233__));
  buf1  g1152(.din(n4284_lo_buf_o2), .dout(new_new_n4234__));
  not1  g1153(.din(n4284_lo_buf_o2), .dout(new_new_n4235__));
  buf1  g1154(.din(n4356_lo_buf_o2), .dout(new_new_n4236__));
  not1  g1155(.din(n4356_lo_buf_o2), .dout(new_new_n4237__));
  buf1  g1156(.din(G2472_o2), .dout(new_new_n4238__));
  not1  g1157(.din(G2472_o2), .dout(new_new_n4239__));
  buf1  g1158(.din(G2410_o2), .dout(new_new_n4240__));
  not1  g1159(.din(G2410_o2), .dout(new_new_n4241__));
  buf1  g1160(.din(n3960_lo_buf_o2), .dout(new_new_n4242__));
  not1  g1161(.din(n3960_lo_buf_o2), .dout(new_new_n4243__));
  buf1  g1162(.din(n3972_lo_buf_o2), .dout(new_new_n4244__));
  buf1  g1163(.din(n2647_inv), .dout(new_new_n4246__));
  not1  g1164(.din(n2647_inv), .dout(new_new_n4247__));
  buf1  g1165(.din(n2650_inv), .dout(new_new_n4248__));
  buf1  g1166(.din(n3684_lo_buf_o2), .dout(new_new_n4250__));
  buf1  g1167(.din(n4080_lo_buf_o2), .dout(new_new_n4252__));
  not1  g1168(.din(n4080_lo_buf_o2), .dout(new_new_n4253__));
  buf1  g1169(.din(n4092_lo_buf_o2), .dout(new_new_n4254__));
  not1  g1170(.din(n4092_lo_buf_o2), .dout(new_new_n4255__));
  buf1  g1171(.din(n2662_inv), .dout(new_new_n4256__));
  not1  g1172(.din(n2662_inv), .dout(new_new_n4257__));
  buf1  g1173(.din(n2665_inv), .dout(new_new_n4258__));
  not1  g1174(.din(n2665_inv), .dout(new_new_n4259__));
  buf1  g1175(.din(G1147_o2), .dout(new_new_n4260__));
  not1  g1176(.din(G1147_o2), .dout(new_new_n4261__));
  buf1  g1177(.din(G2705_o2), .dout(new_new_n4262__));
  not1  g1178(.din(G2705_o2), .dout(new_new_n4263__));
  buf1  g1179(.din(G2693_o2), .dout(new_new_n4264__));
  not1  g1180(.din(G2693_o2), .dout(new_new_n4265__));
  buf1  g1181(.din(G2696_o2), .dout(new_new_n4266__));
  not1  g1182(.din(G2696_o2), .dout(new_new_n4267__));
  buf1  g1183(.din(G2700_o2), .dout(new_new_n4268__));
  not1  g1184(.din(G2700_o2), .dout(new_new_n4269__));
  buf1  g1185(.din(G2915_o2), .dout(new_new_n4270__));
  not1  g1186(.din(G2915_o2), .dout(new_new_n4271__));
  buf1  g1187(.din(G2966_o2), .dout(new_new_n4272__));
  not1  g1188(.din(G2966_o2), .dout(new_new_n4273__));
  buf1  g1189(.din(G2540_o2), .dout(new_new_n4274__));
  not1  g1190(.din(G2540_o2), .dout(new_new_n4275__));
  buf1  g1191(.din(G2788_o2), .dout(new_new_n4276__));
  not1  g1192(.din(G2788_o2), .dout(new_new_n4277__));
  buf1  g1193(.din(G2792_o2), .dout(new_new_n4278__));
  not1  g1194(.din(G2792_o2), .dout(new_new_n4279__));
  buf1  g1195(.din(G2797_o2), .dout(new_new_n4280__));
  not1  g1196(.din(G2797_o2), .dout(new_new_n4281__));
  buf1  g1197(.din(G2804_o2), .dout(new_new_n4282__));
  not1  g1198(.din(G2804_o2), .dout(new_new_n4283__));
  buf1  g1199(.din(G1038_o2), .dout(new_new_n4284__));
  not1  g1200(.din(G1038_o2), .dout(new_new_n4285__));
  buf1  g1201(.din(G1044_o2), .dout(new_new_n4286__));
  not1  g1202(.din(G1044_o2), .dout(new_new_n4287__));
  buf1  g1203(.din(G1090_o2), .dout(new_new_n4288__));
  not1  g1204(.din(G1090_o2), .dout(new_new_n4289__));
  buf1  g1205(.din(G1096_o2), .dout(new_new_n4290__));
  not1  g1206(.din(G1096_o2), .dout(new_new_n4291__));
  buf1  g1207(.din(G1029_o2), .dout(new_new_n4292__));
  not1  g1208(.din(G1029_o2), .dout(new_new_n4293__));
  buf1  g1209(.din(G3942_o2), .dout(new_new_n4294__));
  not1  g1210(.din(G3942_o2), .dout(new_new_n4295__));
  buf1  g1211(.din(G3954_o2), .dout(new_new_n4296__));
  not1  g1212(.din(G3954_o2), .dout(new_new_n4297__));
  buf1  g1213(.din(G4011_o2), .dout(new_new_n4298__));
  not1  g1214(.din(G4011_o2), .dout(new_new_n4299__));
  buf1  g1215(.din(G4017_o2), .dout(new_new_n4300__));
  not1  g1216(.din(G4017_o2), .dout(new_new_n4301__));
  buf1  g1217(.din(G1141_o2), .dout(new_new_n4302__));
  not1  g1218(.din(G1141_o2), .dout(new_new_n4303__));
  buf1  g1219(.din(G1081_o2), .dout(new_new_n4304__));
  not1  g1220(.din(G1081_o2), .dout(new_new_n4305__));
  buf1  g1221(.din(G2146_o2), .dout(new_new_n4306__));
  not1  g1222(.din(G2146_o2), .dout(new_new_n4307__));
  buf1  g1223(.din(G2145_o2), .dout(new_new_n4308__));
  not1  g1224(.din(G2145_o2), .dout(new_new_n4309__));
  buf1  g1225(.din(G2144_o2), .dout(new_new_n4310__));
  not1  g1226(.din(G2144_o2), .dout(new_new_n4311__));
  buf1  g1227(.din(G2143_o2), .dout(new_new_n4312__));
  not1  g1228(.din(G2143_o2), .dout(new_new_n4313__));
  buf1  g1229(.din(G2142_o2), .dout(new_new_n4314__));
  not1  g1230(.din(G2142_o2), .dout(new_new_n4315__));
  buf1  g1231(.din(G2141_o2), .dout(new_new_n4316__));
  not1  g1232(.din(G2141_o2), .dout(new_new_n4317__));
  buf1  g1233(.din(G2140_o2), .dout(new_new_n4318__));
  not1  g1234(.din(G2140_o2), .dout(new_new_n4319__));
  buf1  g1235(.din(G2139_o2), .dout(new_new_n4320__));
  not1  g1236(.din(G2139_o2), .dout(new_new_n4321__));
  buf1  g1237(.din(G3769_o2), .dout(new_new_n4322__));
  not1  g1238(.din(G3769_o2), .dout(new_new_n4323__));
  buf1  g1239(.din(G3773_o2), .dout(new_new_n4324__));
  not1  g1240(.din(G3773_o2), .dout(new_new_n4325__));
  buf1  g1241(.din(G3768_o2), .dout(new_new_n4326__));
  not1  g1242(.din(G3768_o2), .dout(new_new_n4327__));
  buf1  g1243(.din(G4101_o2), .dout(new_new_n4328__));
  not1  g1244(.din(G4101_o2), .dout(new_new_n4329__));
  buf1  g1245(.din(G3161_o2), .dout(new_new_n4330__));
  not1  g1246(.din(G3161_o2), .dout(new_new_n4331__));
  buf1  g1247(.din(G4143_o2), .dout(new_new_n4332__));
  not1  g1248(.din(G4143_o2), .dout(new_new_n4333__));
  buf1  g1249(.din(G3828_o2), .dout(new_new_n4334__));
  not1  g1250(.din(G3828_o2), .dout(new_new_n4335__));
  buf1  g1251(.din(G3831_o2), .dout(new_new_n4336__));
  not1  g1252(.din(G3831_o2), .dout(new_new_n4337__));
  buf1  g1253(.din(G3334_o2), .dout(new_new_n4338__));
  not1  g1254(.din(G3334_o2), .dout(new_new_n4339__));
  buf1  g1255(.din(G3335_o2), .dout(new_new_n4340__));
  not1  g1256(.din(G3335_o2), .dout(new_new_n4341__));
  buf1  g1257(.din(G3180_o2), .dout(new_new_n4342__));
  not1  g1258(.din(G3180_o2), .dout(new_new_n4343__));
  buf1  g1259(.din(G3340_o2), .dout(new_new_n4344__));
  not1  g1260(.din(G3340_o2), .dout(new_new_n4345__));
  buf1  g1261(.din(G3339_o2), .dout(new_new_n4346__));
  not1  g1262(.din(G3339_o2), .dout(new_new_n4347__));
  buf1  g1263(.din(G3341_o2), .dout(new_new_n4348__));
  not1  g1264(.din(G3341_o2), .dout(new_new_n4349__));
  buf1  g1265(.din(G3234_o2), .dout(new_new_n4350__));
  not1  g1266(.din(G3234_o2), .dout(new_new_n4351__));
  buf1  g1267(.din(G3829_o2), .dout(new_new_n4352__));
  not1  g1268(.din(G3829_o2), .dout(new_new_n4353__));
  buf1  g1269(.din(G3338_o2), .dout(new_new_n4354__));
  not1  g1270(.din(G3338_o2), .dout(new_new_n4355__));
  buf1  g1271(.din(G3336_o2), .dout(new_new_n4356__));
  not1  g1272(.din(G3336_o2), .dout(new_new_n4357__));
  buf1  g1273(.din(G3770_o2), .dout(new_new_n4358__));
  not1  g1274(.din(G3770_o2), .dout(new_new_n4359__));
  buf1  g1275(.din(G3918_o2), .dout(new_new_n4360__));
  not1  g1276(.din(G3918_o2), .dout(new_new_n4361__));
  buf1  g1277(.din(G3774_o2), .dout(new_new_n4362__));
  not1  g1278(.din(G3774_o2), .dout(new_new_n4363__));
  buf1  g1279(.din(G3921_o2), .dout(new_new_n4364__));
  not1  g1280(.din(G3921_o2), .dout(new_new_n4365__));
  buf1  g1281(.din(G3832_o2), .dout(new_new_n4366__));
  not1  g1282(.din(G3832_o2), .dout(new_new_n4367__));
  buf1  g1283(.din(G3993_o2), .dout(new_new_n4368__));
  not1  g1284(.din(G3993_o2), .dout(new_new_n4369__));
  buf1  g1285(.din(G2076_o2), .dout(new_new_n4370__));
  not1  g1286(.din(G2076_o2), .dout(new_new_n4371__));
  buf1  g1287(.din(G2071_o2), .dout(new_new_n4372__));
  not1  g1288(.din(G2071_o2), .dout(new_new_n4373__));
  buf1  g1289(.din(G2072_o2), .dout(new_new_n4374__));
  not1  g1290(.din(G2072_o2), .dout(new_new_n4375__));
  buf1  g1291(.din(G2069_o2), .dout(new_new_n4376__));
  not1  g1292(.din(G2069_o2), .dout(new_new_n4377__));
  buf1  g1293(.din(G2070_o2), .dout(new_new_n4378__));
  not1  g1294(.din(G2070_o2), .dout(new_new_n4379__));
  buf1  g1295(.din(G2067_o2), .dout(new_new_n4380__));
  not1  g1296(.din(G2067_o2), .dout(new_new_n4381__));
  buf1  g1297(.din(G2068_o2), .dout(new_new_n4382__));
  not1  g1298(.din(G2068_o2), .dout(new_new_n4383__));
  buf1  g1299(.din(G4095_o2), .dout(new_new_n4384__));
  not1  g1300(.din(G4095_o2), .dout(new_new_n4385__));
  buf1  g1301(.din(G3272_o2), .dout(new_new_n4386__));
  not1  g1302(.din(G3272_o2), .dout(new_new_n4387__));
  buf1  g1303(.din(G3269_o2), .dout(new_new_n4388__));
  not1  g1304(.din(G3269_o2), .dout(new_new_n4389__));
  buf1  g1305(.din(G3270_o2), .dout(new_new_n4390__));
  not1  g1306(.din(G3270_o2), .dout(new_new_n4391__));
  buf1  g1307(.din(G3271_o2), .dout(new_new_n4392__));
  not1  g1308(.din(G3271_o2), .dout(new_new_n4393__));
  buf1  g1309(.din(G3265_o2), .dout(new_new_n4394__));
  not1  g1310(.din(G3265_o2), .dout(new_new_n4395__));
  buf1  g1311(.din(G3266_o2), .dout(new_new_n4396__));
  not1  g1312(.din(G3266_o2), .dout(new_new_n4397__));
  buf1  g1313(.din(G4137_o2), .dout(new_new_n4398__));
  not1  g1314(.din(G4137_o2), .dout(new_new_n4399__));
  buf1  g1315(.din(G3268_o2), .dout(new_new_n4400__));
  not1  g1316(.din(G3268_o2), .dout(new_new_n4401__));
  buf1  g1317(.din(G2361_o2), .dout(new_new_n4402__));
  not1  g1318(.din(G2361_o2), .dout(new_new_n4403__));
  buf1  g1319(.din(G3228_o2), .dout(new_new_n4404__));
  not1  g1320(.din(G3228_o2), .dout(new_new_n4405__));
  buf1  g1321(.din(G3267_o2), .dout(new_new_n4406__));
  not1  g1322(.din(G3267_o2), .dout(new_new_n4407__));
  buf1  g1323(.din(G2336_o2), .dout(new_new_n4408__));
  not1  g1324(.din(G2336_o2), .dout(new_new_n4409__));
  buf1  g1325(.din(G3459_o2), .dout(new_new_n4410__));
  not1  g1326(.din(G3459_o2), .dout(new_new_n4411__));
  buf1  g1327(.din(G3428_o2), .dout(new_new_n4412__));
  not1  g1328(.din(G3428_o2), .dout(new_new_n4413__));
  buf1  g1329(.din(G3438_o2), .dout(new_new_n4414__));
  not1  g1330(.din(G3438_o2), .dout(new_new_n4415__));
  buf1  g1331(.din(G3449_o2), .dout(new_new_n4416__));
  not1  g1332(.din(G3449_o2), .dout(new_new_n4417__));
  buf1  g1333(.din(G3421_o2), .dout(new_new_n4418__));
  not1  g1334(.din(G3421_o2), .dout(new_new_n4419__));
  buf1  g1335(.din(G3576_o2), .dout(new_new_n4420__));
  not1  g1336(.din(G3576_o2), .dout(new_new_n4421__));
  buf1  g1337(.din(G3303_o2), .dout(new_new_n4422__));
  not1  g1338(.din(G3303_o2), .dout(new_new_n4423__));
  buf1  g1339(.din(G3583_o2), .dout(new_new_n4424__));
  not1  g1340(.din(G3583_o2), .dout(new_new_n4425__));
  buf1  g1341(.din(G3594_o2), .dout(new_new_n4426__));
  not1  g1342(.din(G3594_o2), .dout(new_new_n4427__));
  buf1  g1343(.din(G3674_o2), .dout(new_new_n4428__));
  not1  g1344(.din(G3674_o2), .dout(new_new_n4429__));
  buf1  g1345(.din(G3685_o2), .dout(new_new_n4430__));
  not1  g1346(.din(G3685_o2), .dout(new_new_n4431__));
  buf1  g1347(.din(G4504_o2), .dout(new_new_n4432__));
  not1  g1348(.din(G4504_o2), .dout(new_new_n4433__));
  buf1  g1349(.din(G4180_o2), .dout(new_new_n4434__));
  not1  g1350(.din(G4180_o2), .dout(new_new_n4435__));
  not1  g1351(.din(G5123_o2), .dout(new_new_n4437__));
  buf1  g1352(.din(G5142_o2), .dout(new_new_n4438__));
  buf1  g1353(.din(G5126_o2), .dout(new_new_n4440__));
  buf1  g1354(.din(G5144_o2), .dout(new_new_n4442__));
  buf1  g1355(.din(G3912_o2), .dout(new_new_n4444__));
  not1  g1356(.din(G3912_o2), .dout(new_new_n4445__));
  buf1  g1357(.din(G4417_o2), .dout(new_new_n4446__));
  not1  g1358(.din(G4417_o2), .dout(new_new_n4447__));
  buf1  g1359(.din(G4420_o2), .dout(new_new_n4448__));
  not1  g1360(.din(G4420_o2), .dout(new_new_n4449__));
  buf1  g1361(.din(G3969_o2), .dout(new_new_n4450__));
  not1  g1362(.din(G3969_o2), .dout(new_new_n4451__));
  buf1  g1363(.din(G4023_o2), .dout(new_new_n4452__));
  not1  g1364(.din(G4023_o2), .dout(new_new_n4453__));
  buf1  g1365(.din(G2720_o2), .dout(new_new_n4454__));
  not1  g1366(.din(G2720_o2), .dout(new_new_n4455__));
  buf1  g1367(.din(G2837_o2), .dout(new_new_n4456__));
  not1  g1368(.din(G2837_o2), .dout(new_new_n4457__));
  buf1  g1369(.din(n2965_inv), .dout(new_new_n4458__));
  not1  g1370(.din(n2965_inv), .dout(new_new_n4459__));
  buf1  g1371(.din(n2968_inv), .dout(new_new_n4460__));
  not1  g1372(.din(n2968_inv), .dout(new_new_n4461__));
  buf1  g1373(.din(n2971_inv), .dout(new_new_n4462__));
  not1  g1374(.din(n2971_inv), .dout(new_new_n4463__));
  buf1  g1375(.din(n2974_inv), .dout(new_new_n4464__));
  not1  g1376(.din(n2974_inv), .dout(new_new_n4465__));
  buf1  g1377(.din(G1876_o2), .dout(new_new_n4466__));
  not1  g1378(.din(G1876_o2), .dout(new_new_n4467__));
  buf1  g1379(.din(G4996_o2), .dout(new_new_n4468__));
  not1  g1380(.din(G4996_o2), .dout(new_new_n4469__));
  buf1  g1381(.din(G4984_o2), .dout(new_new_n4470__));
  not1  g1382(.din(G4984_o2), .dout(new_new_n4471__));
  buf1  g1383(.din(G4920_o2), .dout(new_new_n4472__));
  not1  g1384(.din(G4920_o2), .dout(new_new_n4473__));
  buf1  g1385(.din(G4923_o2), .dout(new_new_n4474__));
  not1  g1386(.din(G4923_o2), .dout(new_new_n4475__));
  buf1  g1387(.din(G4930_o2), .dout(new_new_n4476__));
  not1  g1388(.din(G4930_o2), .dout(new_new_n4477__));
  buf1  g1389(.din(G4933_o2), .dout(new_new_n4478__));
  not1  g1390(.din(G4933_o2), .dout(new_new_n4479__));
  buf1  g1391(.din(n4320_lo_buf_o2), .dout(new_new_n4480__));
  not1  g1392(.din(n4320_lo_buf_o2), .dout(new_new_n4481__));
  buf1  g1393(.din(G2424_o2), .dout(new_new_n4482__));
  not1  g1394(.din(G2424_o2), .dout(new_new_n4483__));
  buf1  g1395(.din(G3317_o2), .dout(new_new_n4484__));
  buf1  g1396(.din(G3503_o2), .dout(new_new_n4486__));
  buf1  g1397(.din(G3485_o2), .dout(new_new_n4488__));
  not1  g1398(.din(G3485_o2), .dout(new_new_n4489__));
  buf1  g1399(.din(G3611_o2), .dout(new_new_n4490__));
  not1  g1400(.din(G3611_o2), .dout(new_new_n4491__));
  buf1  g1401(.din(n3864_lo_buf_o2), .dout(new_new_n4492__));
  buf1  g1402(.din(n3888_lo_buf_o2), .dout(new_new_n4494__));
  buf1  g1403(.din(n4116_lo_buf_o2), .dout(new_new_n4496__));
  buf1  g1404(.din(n4128_lo_buf_o2), .dout(new_new_n4498__));
  buf1  g1405(.din(n4140_lo_buf_o2), .dout(new_new_n4500__));
  buf1  g1406(.din(n4152_lo_buf_o2), .dout(new_new_n4502__));
  buf1  g1407(.din(G1815_o2), .dout(new_new_n4504__));
  not1  g1408(.din(G1815_o2), .dout(new_new_n4505__));
  buf1  g1409(.din(G1728_o2), .dout(new_new_n4506__));
  not1  g1410(.din(G1728_o2), .dout(new_new_n4507__));
  buf1  g1411(.din(G1035_o2), .dout(new_new_n4508__));
  not1  g1412(.din(G1035_o2), .dout(new_new_n4509__));
  buf1  g1413(.din(G1041_o2), .dout(new_new_n4510__));
  not1  g1414(.din(G1041_o2), .dout(new_new_n4511__));
  buf1  g1415(.din(G1087_o2), .dout(new_new_n4512__));
  not1  g1416(.din(G1087_o2), .dout(new_new_n4513__));
  buf1  g1417(.din(G1093_o2), .dout(new_new_n4514__));
  not1  g1418(.din(G1093_o2), .dout(new_new_n4515__));
  buf1  g1419(.din(G1132_o2), .dout(new_new_n4516__));
  not1  g1420(.din(G1132_o2), .dout(new_new_n4517__));
  buf1  g1421(.din(G1108_o2), .dout(new_new_n4518__));
  not1  g1422(.din(G1108_o2), .dout(new_new_n4519__));
  buf1  g1423(.din(G1138_o2), .dout(new_new_n4520__));
  not1  g1424(.din(G1138_o2), .dout(new_new_n4521__));
  buf1  g1425(.din(G1114_o2), .dout(new_new_n4522__));
  not1  g1426(.din(G1114_o2), .dout(new_new_n4523__));
  buf1  g1427(.din(G1807_o2), .dout(new_new_n4524__));
  not1  g1428(.din(G1807_o2), .dout(new_new_n4525__));
  buf1  g1429(.din(G2108_o2), .dout(new_new_n4526__));
  not1  g1430(.din(G2108_o2), .dout(new_new_n4527__));
  buf1  g1431(.din(G1126_o2), .dout(new_new_n4528__));
  not1  g1432(.din(G1126_o2), .dout(new_new_n4529__));
  buf1  g1433(.din(G1899_o2), .dout(new_new_n4530__));
  not1  g1434(.din(G1899_o2), .dout(new_new_n4531__));
  buf1  g1435(.din(G2134_o2), .dout(new_new_n4532__));
  not1  g1436(.din(G2134_o2), .dout(new_new_n4533__));
  buf1  g1437(.din(G1852_o2), .dout(new_new_n4534__));
  not1  g1438(.din(G1852_o2), .dout(new_new_n4535__));
  buf1  g1439(.din(G2116_o2), .dout(new_new_n4536__));
  not1  g1440(.din(G2116_o2), .dout(new_new_n4537__));
  buf1  g1441(.din(G2543_o2), .dout(new_new_n4538__));
  not1  g1442(.din(G2543_o2), .dout(new_new_n4539__));
  buf1  g1443(.din(G2727_o2), .dout(new_new_n4540__));
  not1  g1444(.din(G2727_o2), .dout(new_new_n4541__));
  buf1  g1445(.din(G2715_o2), .dout(new_new_n4542__));
  not1  g1446(.din(G2715_o2), .dout(new_new_n4543__));
  buf1  g1447(.din(G2832_o2), .dout(new_new_n4544__));
  not1  g1448(.din(G2832_o2), .dout(new_new_n4545__));
  buf1  g1449(.din(G1873_o2), .dout(new_new_n4546__));
  not1  g1450(.din(G1873_o2), .dout(new_new_n4547__));
  buf1  g1451(.din(G3291_o2), .dout(new_new_n4548__));
  not1  g1452(.din(G3291_o2), .dout(new_new_n4549__));
  buf1  g1453(.din(G5025_o2), .dout(new_new_n4550__));
  not1  g1454(.din(G5025_o2), .dout(new_new_n4551__));
  buf1  g1455(.din(G5036_o2), .dout(new_new_n4552__));
  not1  g1456(.din(G5036_o2), .dout(new_new_n4553__));
  buf1  g1457(.din(G3132_o2), .dout(new_new_n4554__));
  not1  g1458(.din(G3132_o2), .dout(new_new_n4555__));
  buf1  g1459(.din(G5038_o2), .dout(new_new_n4556__));
  not1  g1460(.din(G5038_o2), .dout(new_new_n4557__));
  buf1  g1461(.din(G5039_o2), .dout(new_new_n4558__));
  not1  g1462(.din(G5039_o2), .dout(new_new_n4559__));
  buf1  g1463(.din(n3118_inv), .dout(new_new_n4560__));
  not1  g1464(.din(n3118_inv), .dout(new_new_n4561__));
  buf1  g1465(.din(n3121_inv), .dout(new_new_n4562__));
  not1  g1466(.din(n3121_inv), .dout(new_new_n4563__));
  buf1  g1467(.din(n3124_inv), .dout(new_new_n4564__));
  not1  g1468(.din(n3124_inv), .dout(new_new_n4565__));
  buf1  g1469(.din(n3127_inv), .dout(new_new_n4566__));
  not1  g1470(.din(n3127_inv), .dout(new_new_n4567__));
  buf1  g1471(.din(n3984_lo_buf_o2), .dout(new_new_n4568__));
  buf1  g1472(.din(G1802_o2), .dout(new_new_n4570__));
  not1  g1473(.din(G1802_o2), .dout(new_new_n4571__));
  buf1  g1474(.din(G1804_o2), .dout(new_new_n4572__));
  not1  g1475(.din(G1804_o2), .dout(new_new_n4573__));
  buf1  g1476(.din(G1849_o2), .dout(new_new_n4574__));
  not1  g1477(.din(G1849_o2), .dout(new_new_n4575__));
  buf1  g1478(.din(G1851_o2), .dout(new_new_n4576__));
  not1  g1479(.din(G1851_o2), .dout(new_new_n4577__));
  buf1  g1480(.din(G2492_o2), .dout(new_new_n4578__));
  not1  g1481(.din(G2492_o2), .dout(new_new_n4579__));
  buf1  g1482(.din(G1799_o2), .dout(new_new_n4580__));
  not1  g1483(.din(G1799_o2), .dout(new_new_n4581__));
  buf1  g1484(.din(G4231_o2), .dout(new_new_n4582__));
  not1  g1485(.din(G4231_o2), .dout(new_new_n4583__));
  buf1  g1486(.din(G4234_o2), .dout(new_new_n4584__));
  not1  g1487(.din(G4234_o2), .dout(new_new_n4585__));
  buf1  g1488(.din(G4245_o2), .dout(new_new_n4586__));
  not1  g1489(.din(G4245_o2), .dout(new_new_n4587__));
  buf1  g1490(.din(G4247_o2), .dout(new_new_n4588__));
  not1  g1491(.din(G4247_o2), .dout(new_new_n4589__));
  buf1  g1492(.din(G1894_o2), .dout(new_new_n4590__));
  not1  g1493(.din(G1894_o2), .dout(new_new_n4591__));
  buf1  g1494(.din(G1846_o2), .dout(new_new_n4592__));
  not1  g1495(.din(G1846_o2), .dout(new_new_n4593__));
  buf1  g1496(.din(G4238_o2), .dout(new_new_n4594__));
  not1  g1497(.din(G4238_o2), .dout(new_new_n4595__));
  buf1  g1498(.din(G4249_o2), .dout(new_new_n4596__));
  not1  g1499(.din(G4249_o2), .dout(new_new_n4597__));
  buf1  g1500(.din(G2293_o2), .dout(new_new_n4598__));
  not1  g1501(.din(G2293_o2), .dout(new_new_n4599__));
  buf1  g1502(.din(G5022_o2), .dout(new_new_n4600__));
  not1  g1503(.din(G5022_o2), .dout(new_new_n4601__));
  buf1  g1504(.din(G5006_o2), .dout(new_new_n4602__));
  not1  g1505(.din(G5006_o2), .dout(new_new_n4603__));
  buf1  g1506(.din(G4944_o2), .dout(new_new_n4604__));
  not1  g1507(.din(G4944_o2), .dout(new_new_n4605__));
  buf1  g1508(.din(G4946_o2), .dout(new_new_n4606__));
  not1  g1509(.din(G4946_o2), .dout(new_new_n4607__));
  buf1  g1510(.din(G4954_o2), .dout(new_new_n4608__));
  not1  g1511(.din(G4954_o2), .dout(new_new_n4609__));
  buf1  g1512(.din(G4956_o2), .dout(new_new_n4610__));
  not1  g1513(.din(G4956_o2), .dout(new_new_n4611__));
  buf1  g1514(.din(G3546_o2), .dout(new_new_n4612__));
  not1  g1515(.din(G3546_o2), .dout(new_new_n4613__));
  buf1  g1516(.din(G3658_o2), .dout(new_new_n4614__));
  not1  g1517(.din(G3658_o2), .dout(new_new_n4615__));
  buf1  g1518(.din(G1344_o2), .dout(new_new_n4616__));
  not1  g1519(.din(G1344_o2), .dout(new_new_n4617__));
  buf1  g1520(.din(G2921_o2), .dout(new_new_n4618__));
  not1  g1521(.din(G2921_o2), .dout(new_new_n4619__));
  buf1  g1522(.din(n3912_lo_buf_o2), .dout(new_new_n4620__));
  buf1  g1523(.din(G1835_o2), .dout(new_new_n4622__));
  not1  g1524(.din(G1835_o2), .dout(new_new_n4623__));
  buf1  g1525(.din(G3810_o2), .dout(new_new_n4624__));
  not1  g1526(.din(G3810_o2), .dout(new_new_n4625__));
  buf1  g1527(.din(G3866_o2), .dout(new_new_n4626__));
  not1  g1528(.din(G3866_o2), .dout(new_new_n4627__));
  buf1  g1529(.din(G3811_o2), .dout(new_new_n4628__));
  not1  g1530(.din(G3811_o2), .dout(new_new_n4629__));
  buf1  g1531(.din(G2269_o2), .dout(new_new_n4630__));
  not1  g1532(.din(G2269_o2), .dout(new_new_n4631__));
  buf1  g1533(.din(G3812_o2), .dout(new_new_n4632__));
  not1  g1534(.din(G3812_o2), .dout(new_new_n4633__));
  buf1  g1535(.din(G3867_o2), .dout(new_new_n4634__));
  not1  g1536(.din(G3867_o2), .dout(new_new_n4635__));
  buf1  g1537(.din(G3868_o2), .dout(new_new_n4636__));
  not1  g1538(.din(G3868_o2), .dout(new_new_n4637__));
  buf1  g1539(.din(G3809_o2), .dout(new_new_n4638__));
  not1  g1540(.din(G3809_o2), .dout(new_new_n4639__));
  buf1  g1541(.din(G3716_o2), .dout(new_new_n4640__));
  not1  g1542(.din(G3716_o2), .dout(new_new_n4641__));
  buf1  g1543(.din(G4529_o2), .dout(new_new_n4642__));
  not1  g1544(.din(G4529_o2), .dout(new_new_n4643__));
  buf1  g1545(.din(G4670_o2), .dout(new_new_n4644__));
  not1  g1546(.din(G4670_o2), .dout(new_new_n4645__));
  buf1  g1547(.din(G4493_o2), .dout(new_new_n4646__));
  not1  g1548(.din(G4493_o2), .dout(new_new_n4647__));
  buf1  g1549(.din(G4580_o2), .dout(new_new_n4648__));
  not1  g1550(.din(G4580_o2), .dout(new_new_n4649__));
  buf1  g1551(.din(G3822_o2), .dout(new_new_n4650__));
  not1  g1552(.din(G3822_o2), .dout(new_new_n4651__));
  buf1  g1553(.din(G3877_o2), .dout(new_new_n4652__));
  not1  g1554(.din(G3877_o2), .dout(new_new_n4653__));
  buf1  g1555(.din(G4131_o2), .dout(new_new_n4654__));
  not1  g1556(.din(G4131_o2), .dout(new_new_n4655__));
  buf1  g1557(.din(G4170_o2), .dout(new_new_n4656__));
  not1  g1558(.din(G4170_o2), .dout(new_new_n4657__));
  buf1  g1559(.din(G4051_o2), .dout(new_new_n4658__));
  not1  g1560(.din(G4051_o2), .dout(new_new_n4659__));
  buf1  g1561(.din(G4065_o2), .dout(new_new_n4660__));
  not1  g1562(.din(G4065_o2), .dout(new_new_n4661__));
  buf1  g1563(.din(G4697_o2), .dout(new_new_n4662__));
  not1  g1564(.din(G4697_o2), .dout(new_new_n4663__));
  buf1  g1565(.din(G4706_o2), .dout(new_new_n4664__));
  not1  g1566(.din(G4706_o2), .dout(new_new_n4665__));
  buf1  g1567(.din(G2460_o2), .dout(new_new_n4666__));
  not1  g1568(.din(G2460_o2), .dout(new_new_n4667__));
  buf1  g1569(.din(G2454_o2), .dout(new_new_n4668__));
  not1  g1570(.din(G2454_o2), .dout(new_new_n4669__));
  buf1  g1571(.din(G2392_o2), .dout(new_new_n4670__));
  not1  g1572(.din(G2392_o2), .dout(new_new_n4671__));
  buf1  g1573(.din(G2386_o2), .dout(new_new_n4672__));
  not1  g1574(.din(G2386_o2), .dout(new_new_n4673__));
  buf1  g1575(.din(n4260_lo_buf_o2), .dout(new_new_n4674__));
  not1  g1576(.din(n4260_lo_buf_o2), .dout(new_new_n4675__));
  buf1  g1577(.din(n4272_lo_buf_o2), .dout(new_new_n4676__));
  not1  g1578(.din(n4272_lo_buf_o2), .dout(new_new_n4677__));
  buf1  g1579(.din(n4392_lo_buf_o2), .dout(new_new_n4678__));
  not1  g1580(.din(n4392_lo_buf_o2), .dout(new_new_n4679__));
  buf1  g1581(.din(n4404_lo_buf_o2), .dout(new_new_n4680__));
  not1  g1582(.din(n4404_lo_buf_o2), .dout(new_new_n4681__));
  buf1  g1583(.din(G1512_o2), .dout(new_new_n4682__));
  not1  g1584(.din(G1512_o2), .dout(new_new_n4683__));
  buf1  g1585(.din(G3135_o2), .dout(new_new_n4684__));
  not1  g1586(.din(G3135_o2), .dout(new_new_n4685__));
  buf1  g1587(.din(G2379_o2), .dout(new_new_n4686__));
  not1  g1588(.din(G2379_o2), .dout(new_new_n4687__));
  buf1  g1589(.din(n4164_lo_buf_o2), .dout(new_new_n4688__));
  not1  g1590(.din(n4164_lo_buf_o2), .dout(new_new_n4689__));
  buf1  g1591(.din(n4176_lo_buf_o2), .dout(new_new_n4690__));
  not1  g1592(.din(n4176_lo_buf_o2), .dout(new_new_n4691__));
  buf1  g1593(.din(n4224_lo_buf_o2), .dout(new_new_n4692__));
  not1  g1594(.din(n4224_lo_buf_o2), .dout(new_new_n4693__));
  buf1  g1595(.din(G2975_o2), .dout(new_new_n4694__));
  not1  g1596(.din(G2975_o2), .dout(new_new_n4695__));
  buf1  g1597(.din(G2978_o2), .dout(new_new_n4696__));
  not1  g1598(.din(G2978_o2), .dout(new_new_n4697__));
  buf1  g1599(.din(G2933_o2), .dout(new_new_n4698__));
  not1  g1600(.din(G2933_o2), .dout(new_new_n4699__));
  buf1  g1601(.din(G2936_o2), .dout(new_new_n4700__));
  not1  g1602(.din(G2936_o2), .dout(new_new_n4701__));
  buf1  g1603(.din(G1356_o2), .dout(new_new_n4702__));
  not1  g1604(.din(G1356_o2), .dout(new_new_n4703__));
  buf1  g1605(.din(G1359_o2), .dout(new_new_n4704__));
  not1  g1606(.din(G1359_o2), .dout(new_new_n4705__));
  buf1  g1607(.din(G1398_o2), .dout(new_new_n4706__));
  not1  g1608(.din(G1398_o2), .dout(new_new_n4707__));
  buf1  g1609(.din(G1401_o2), .dout(new_new_n4708__));
  not1  g1610(.din(G1401_o2), .dout(new_new_n4709__));
  and1  g1611(.dina(new_new_n3650__), .dinb(new_new_n3626__), .dout(new_new_n4710__));
  and1  g1612(.dina(new_new_n3218__), .dinb(new_new_n8443__), .dout(new_new_n4711__));
  and1  g1613(.dina(new_new_n3538__), .dinb(new_new_n8444__), .dout(new_new_n4712__));
  and1  g1614(.dina(new_new_n8445__), .dinb(new_new_n3186__), .dout(new_new_n4713__));
  or1   g1615(.dina(new_new_n3710__), .dinb(new_new_n8446__), .dout(new_new_n4714__));
  or1   g1616(.dina(new_new_n8447__), .dinb(new_new_n8448__), .dout(new_new_n4715__));
  and1  g1617(.dina(new_new_n2778__), .dinb(new_new_n2770__), .dout(new_new_n4716__));
  or1   g1618(.dina(new_new_n2779__), .dinb(new_new_n8446__), .dout(new_new_n4717__));
  or1   g1619(.dina(new_new_n8452__), .dinb(new_new_n3203__), .dout(new_new_n4718__));
  or1   g1620(.dina(new_new_n8463__), .dinb(new_new_n2955__), .dout(new_new_n4719__));
  or1   g1621(.dina(new_new_n8470__), .dinb(new_new_n2947__), .dout(new_new_n4720__));
  and1  g1622(.dina(new_new_n4720__), .dinb(new_new_n4719__), .dout(new_new_n4721__));
  or1   g1623(.dina(new_new_n4721__), .dinb(new_new_n8452__), .dout(new_new_n4722__));
  or1   g1624(.dina(new_new_n8463__), .dinb(new_new_n2787__), .dout(new_new_n4723__));
  or1   g1625(.dina(new_new_n8470__), .dinb(new_new_n2963__), .dout(new_new_n4724__));
  and1  g1626(.dina(new_new_n4724__), .dinb(new_new_n4723__), .dout(new_new_n4725__));
  or1   g1627(.dina(new_new_n4725__), .dinb(new_new_n8453__), .dout(new_new_n4726__));
  or1   g1628(.dina(new_new_n8464__), .dinb(new_new_n8475__), .dout(new_new_n4727__));
  or1   g1629(.dina(new_new_n8471__), .dinb(new_new_n8475__), .dout(new_new_n4728__));
  and1  g1630(.dina(new_new_n4728__), .dinb(new_new_n4727__), .dout(new_new_n4729__));
  or1   g1631(.dina(new_new_n4729__), .dinb(new_new_n8453__), .dout(new_new_n4730__));
  or1   g1632(.dina(new_new_n8464__), .dinb(new_new_n2747__), .dout(new_new_n4731__));
  or1   g1633(.dina(new_new_n4731__), .dinb(new_new_n8455__), .dout(new_new_n4732__));
  or1   g1634(.dina(new_new_n8471__), .dinb(new_new_n2755__), .dout(new_new_n4733__));
  or1   g1635(.dina(new_new_n4733__), .dinb(new_new_n8455__), .dout(new_new_n4734__));
  or1   g1636(.dina(new_new_n8476__), .dinb(new_new_n8466__), .dout(new_new_n4735__));
  or1   g1637(.dina(new_new_n8476__), .dinb(new_new_n8473__), .dout(new_new_n4736__));
  and1  g1638(.dina(new_new_n4734__), .dinb(new_new_n4732__), .dout(new_new_n4737__));
  and1  g1639(.dina(new_new_n4737__), .dinb(new_new_n8478__), .dout(new_new_n4738__));
  and1  g1640(.dina(new_new_n4738__), .dinb(new_new_n8481__), .dout(new_new_n4739__));
  or1   g1641(.dina(new_new_n4739__), .dinb(new_new_n8485__), .dout(new_new_n4740__));
  or1   g1642(.dina(new_new_n8466__), .dinb(new_new_n2763__), .dout(new_new_n4741__));
  or1   g1643(.dina(new_new_n4741__), .dinb(new_new_n8456__), .dout(new_new_n4742__));
  or1   g1644(.dina(new_new_n8473__), .dinb(new_new_n2923__), .dout(new_new_n4743__));
  or1   g1645(.dina(new_new_n4743__), .dinb(new_new_n8456__), .dout(new_new_n4744__));
  and1  g1646(.dina(new_new_n4744__), .dinb(new_new_n4742__), .dout(new_new_n4745__));
  and1  g1647(.dina(new_new_n4745__), .dinb(new_new_n8478__), .dout(new_new_n4746__));
  and1  g1648(.dina(new_new_n4746__), .dinb(new_new_n8481__), .dout(new_new_n4747__));
  or1   g1649(.dina(new_new_n4747__), .dinb(new_new_n8485__), .dout(new_new_n4748__));
  or1   g1650(.dina(new_new_n8467__), .dinb(new_new_n2907__), .dout(new_new_n4749__));
  or1   g1651(.dina(new_new_n4749__), .dinb(new_new_n8459__), .dout(new_new_n4750__));
  or1   g1652(.dina(new_new_n8474__), .dinb(new_new_n2739__), .dout(new_new_n4751__));
  or1   g1653(.dina(new_new_n4751__), .dinb(new_new_n8459__), .dout(new_new_n4752__));
  and1  g1654(.dina(new_new_n4752__), .dinb(new_new_n4750__), .dout(new_new_n4753__));
  and1  g1655(.dina(new_new_n4753__), .dinb(new_new_n8479__), .dout(new_new_n4754__));
  and1  g1656(.dina(new_new_n4754__), .dinb(new_new_n8482__), .dout(new_new_n4755__));
  or1   g1657(.dina(new_new_n4755__), .dinb(new_new_n8484__), .dout(new_new_n4756__));
  or1   g1658(.dina(new_new_n8467__), .dinb(new_new_n2931__), .dout(new_new_n4757__));
  or1   g1659(.dina(new_new_n4757__), .dinb(new_new_n8458__), .dout(new_new_n4758__));
  or1   g1660(.dina(new_new_n8474__), .dinb(new_new_n2915__), .dout(new_new_n4759__));
  or1   g1661(.dina(new_new_n4759__), .dinb(new_new_n8460__), .dout(new_new_n4760__));
  and1  g1662(.dina(new_new_n4760__), .dinb(new_new_n4758__), .dout(new_new_n4761__));
  and1  g1663(.dina(new_new_n4761__), .dinb(new_new_n8479__), .dout(new_new_n4762__));
  and1  g1664(.dina(new_new_n4762__), .dinb(new_new_n8482__), .dout(new_new_n4763__));
  or1   g1665(.dina(new_new_n4763__), .dinb(new_new_n8486__), .dout(new_new_n4764__));
  or1   g1666(.dina(new_new_n8488__), .dinb(new_new_n8489__), .dout(new_new_n4765__));
  or1   g1667(.dina(new_new_n4765__), .dinb(new_new_n8490__), .dout(new_new_n4766__));
  or1   g1668(.dina(new_new_n8492__), .dinb(new_new_n8489__), .dout(new_new_n4767__));
  or1   g1669(.dina(new_new_n4767__), .dinb(new_new_n8493__), .dout(new_new_n4768__));
  and1  g1670(.dina(new_new_n4768__), .dinb(new_new_n4766__), .dout(new_new_n4769__));
  and1  g1671(.dina(new_new_n8495__), .dinb(new_new_n8493__), .dout(new_new_n4770__));
  and1  g1672(.dina(new_new_n8497__), .dinb(new_new_n8490__), .dout(new_new_n4771__));
  or1   g1673(.dina(new_new_n4771__), .dinb(new_new_n4770__), .dout(new_new_n4772__));
  or1   g1674(.dina(new_new_n4772__), .dinb(new_new_n3588__), .dout(new_new_n4773__));
  and1  g1675(.dina(new_new_n4773__), .dinb(new_new_n4769__), .dout(new_new_n4774__));
  or1   g1676(.dina(new_new_n8488__), .dinb(new_new_n8498__), .dout(new_new_n4775__));
  or1   g1677(.dina(new_new_n4775__), .dinb(new_new_n8499__), .dout(new_new_n4776__));
  or1   g1678(.dina(new_new_n8492__), .dinb(new_new_n8498__), .dout(new_new_n4777__));
  or1   g1679(.dina(new_new_n4777__), .dinb(new_new_n8500__), .dout(new_new_n4778__));
  and1  g1680(.dina(new_new_n4778__), .dinb(new_new_n4776__), .dout(new_new_n4779__));
  and1  g1681(.dina(new_new_n8495__), .dinb(new_new_n8500__), .dout(new_new_n4780__));
  and1  g1682(.dina(new_new_n8497__), .dinb(new_new_n8499__), .dout(new_new_n4781__));
  or1   g1683(.dina(new_new_n4781__), .dinb(new_new_n4780__), .dout(new_new_n4782__));
  or1   g1684(.dina(new_new_n4782__), .dinb(new_new_n3584__), .dout(new_new_n4783__));
  and1  g1685(.dina(new_new_n4783__), .dinb(new_new_n4779__), .dout(new_new_n4784__));
  or1   g1686(.dina(new_new_n8487__), .dinb(new_new_n3478__), .dout(new_new_n4785__));
  or1   g1687(.dina(new_new_n8491__), .dinb(new_new_n3479__), .dout(new_new_n4786__));
  and1  g1688(.dina(new_new_n4786__), .dinb(new_new_n4785__), .dout(new_new_n4787__));
  and1  g1689(.dina(new_new_n8494__), .dinb(new_new_n8502__), .dout(new_new_n4788__));
  or1   g1690(.dina(new_new_n3886__), .dinb(new_new_n8503__), .dout(new_new_n4789__));
  and1  g1691(.dina(new_new_n8496__), .dinb(new_new_n8503__), .dout(new_new_n4790__));
  or1   g1692(.dina(new_new_n3892__), .dinb(new_new_n8502__), .dout(new_new_n4791__));
  and1  g1693(.dina(new_new_n4791__), .dinb(new_new_n4789__), .dout(new_new_n4792__));
  or1   g1694(.dina(new_new_n4790__), .dinb(new_new_n4788__), .dout(new_new_n4793__));
  or1   g1695(.dina(new_new_n8504__), .dinb(new_new_n8505__), .dout(new_new_n4794__));
  or1   g1696(.dina(new_new_n4794__), .dinb(new_new_n8506__), .dout(new_new_n4795__));
  or1   g1697(.dina(new_new_n4795__), .dinb(new_new_n4793__), .dout(new_new_n4796__));
  or1   g1698(.dina(new_new_n8510__), .dinb(new_new_n8518__), .dout(new_new_n4797__));
  or1   g1699(.dina(new_new_n4797__), .dinb(new_new_n8519__), .dout(new_new_n4798__));
  or1   g1700(.dina(new_new_n8523__), .dinb(new_new_n8518__), .dout(new_new_n4799__));
  or1   g1701(.dina(new_new_n4799__), .dinb(new_new_n8530__), .dout(new_new_n4800__));
  and1  g1702(.dina(new_new_n4800__), .dinb(new_new_n4798__), .dout(new_new_n4801__));
  and1  g1703(.dina(new_new_n8534__), .dinb(new_new_n8530__), .dout(new_new_n4802__));
  and1  g1704(.dina(new_new_n8545__), .dinb(new_new_n8519__), .dout(new_new_n4803__));
  or1   g1705(.dina(new_new_n4803__), .dinb(new_new_n4802__), .dout(new_new_n4804__));
  or1   g1706(.dina(new_new_n4804__), .dinb(new_new_n3602__), .dout(new_new_n4805__));
  and1  g1707(.dina(new_new_n4805__), .dinb(new_new_n4801__), .dout(new_new_n4806__));
  or1   g1708(.dina(new_new_n8510__), .dinb(new_new_n8552__), .dout(new_new_n4807__));
  or1   g1709(.dina(new_new_n4807__), .dinb(new_new_n8553__), .dout(new_new_n4808__));
  or1   g1710(.dina(new_new_n8523__), .dinb(new_new_n8552__), .dout(new_new_n4809__));
  or1   g1711(.dina(new_new_n4809__), .dinb(new_new_n8554__), .dout(new_new_n4810__));
  and1  g1712(.dina(new_new_n4810__), .dinb(new_new_n4808__), .dout(new_new_n4811__));
  and1  g1713(.dina(new_new_n8534__), .dinb(new_new_n8554__), .dout(new_new_n4812__));
  and1  g1714(.dina(new_new_n8545__), .dinb(new_new_n8553__), .dout(new_new_n4813__));
  or1   g1715(.dina(new_new_n4813__), .dinb(new_new_n4812__), .dout(new_new_n4814__));
  or1   g1716(.dina(new_new_n4814__), .dinb(new_new_n3600__), .dout(new_new_n4815__));
  and1  g1717(.dina(new_new_n4815__), .dinb(new_new_n4811__), .dout(new_new_n4816__));
  or1   g1718(.dina(new_new_n8511__), .dinb(new_new_n3599__), .dout(new_new_n4817__));
  or1   g1719(.dina(new_new_n8535__), .dinb(new_new_n3598__), .dout(new_new_n4818__));
  and1  g1720(.dina(new_new_n4818__), .dinb(new_new_n4817__), .dout(new_new_n4819__));
  or1   g1721(.dina(new_new_n8511__), .dinb(new_new_n8556__), .dout(new_new_n4820__));
  or1   g1722(.dina(new_new_n4820__), .dinb(new_new_n8557__), .dout(new_new_n4821__));
  or1   g1723(.dina(new_new_n8524__), .dinb(new_new_n8556__), .dout(new_new_n4822__));
  or1   g1724(.dina(new_new_n4822__), .dinb(new_new_n8558__), .dout(new_new_n4823__));
  and1  g1725(.dina(new_new_n4823__), .dinb(new_new_n4821__), .dout(new_new_n4824__));
  and1  g1726(.dina(new_new_n8535__), .dinb(new_new_n8558__), .dout(new_new_n4825__));
  and1  g1727(.dina(new_new_n8546__), .dinb(new_new_n8557__), .dout(new_new_n4826__));
  or1   g1728(.dina(new_new_n4826__), .dinb(new_new_n4825__), .dout(new_new_n4827__));
  or1   g1729(.dina(new_new_n4827__), .dinb(new_new_n8559__), .dout(new_new_n4828__));
  and1  g1730(.dina(new_new_n4828__), .dinb(new_new_n4824__), .dout(new_new_n4829__));
  or1   g1731(.dina(new_new_n8560__), .dinb(new_new_n8561__), .dout(new_new_n4830__));
  or1   g1732(.dina(new_new_n4830__), .dinb(new_new_n8562__), .dout(new_new_n4831__));
  or1   g1733(.dina(new_new_n4831__), .dinb(new_new_n8563__), .dout(new_new_n4832__));
  or1   g1734(.dina(new_new_n4832__), .dinb(new_new_n4796__), .dout(new_new_n4833__));
  or1   g1735(.dina(new_new_n4833__), .dinb(new_new_n4028__), .dout(new_new_n4834__));
  or1   g1736(.dina(new_new_n8513__), .dinb(new_new_n8565__), .dout(new_new_n4835__));
  or1   g1737(.dina(new_new_n4835__), .dinb(new_new_n8566__), .dout(new_new_n4836__));
  or1   g1738(.dina(new_new_n8524__), .dinb(new_new_n8565__), .dout(new_new_n4837__));
  or1   g1739(.dina(new_new_n4837__), .dinb(new_new_n8567__), .dout(new_new_n4838__));
  and1  g1740(.dina(new_new_n4838__), .dinb(new_new_n4836__), .dout(new_new_n4839__));
  and1  g1741(.dina(new_new_n8537__), .dinb(new_new_n8567__), .dout(new_new_n4840__));
  and1  g1742(.dina(new_new_n8546__), .dinb(new_new_n8566__), .dout(new_new_n4841__));
  or1   g1743(.dina(new_new_n4841__), .dinb(new_new_n4840__), .dout(new_new_n4842__));
  or1   g1744(.dina(new_new_n4842__), .dinb(new_new_n8568__), .dout(new_new_n4843__));
  and1  g1745(.dina(new_new_n4843__), .dinb(new_new_n4839__), .dout(new_new_n4844__));
  or1   g1746(.dina(new_new_n8513__), .dinb(new_new_n8569__), .dout(new_new_n4845__));
  or1   g1747(.dina(new_new_n4845__), .dinb(new_new_n8570__), .dout(new_new_n4846__));
  or1   g1748(.dina(new_new_n8526__), .dinb(new_new_n8569__), .dout(new_new_n4847__));
  or1   g1749(.dina(new_new_n4847__), .dinb(new_new_n8571__), .dout(new_new_n4848__));
  and1  g1750(.dina(new_new_n4848__), .dinb(new_new_n4846__), .dout(new_new_n4849__));
  and1  g1751(.dina(new_new_n8537__), .dinb(new_new_n8571__), .dout(new_new_n4850__));
  and1  g1752(.dina(new_new_n8548__), .dinb(new_new_n8570__), .dout(new_new_n4851__));
  or1   g1753(.dina(new_new_n4851__), .dinb(new_new_n4850__), .dout(new_new_n4852__));
  or1   g1754(.dina(new_new_n4852__), .dinb(new_new_n3560__), .dout(new_new_n4853__));
  and1  g1755(.dina(new_new_n4853__), .dinb(new_new_n4849__), .dout(new_new_n4854__));
  or1   g1756(.dina(new_new_n8514__), .dinb(new_new_n8572__), .dout(new_new_n4855__));
  or1   g1757(.dina(new_new_n4855__), .dinb(new_new_n8573__), .dout(new_new_n4856__));
  or1   g1758(.dina(new_new_n8526__), .dinb(new_new_n8572__), .dout(new_new_n4857__));
  or1   g1759(.dina(new_new_n4857__), .dinb(new_new_n8574__), .dout(new_new_n4858__));
  and1  g1760(.dina(new_new_n4858__), .dinb(new_new_n4856__), .dout(new_new_n4859__));
  and1  g1761(.dina(new_new_n8538__), .dinb(new_new_n8574__), .dout(new_new_n4860__));
  and1  g1762(.dina(new_new_n8548__), .dinb(new_new_n8573__), .dout(new_new_n4861__));
  or1   g1763(.dina(new_new_n4861__), .dinb(new_new_n4860__), .dout(new_new_n4862__));
  or1   g1764(.dina(new_new_n4862__), .dinb(new_new_n3580__), .dout(new_new_n4863__));
  and1  g1765(.dina(new_new_n4863__), .dinb(new_new_n4859__), .dout(new_new_n4864__));
  or1   g1766(.dina(new_new_n8514__), .dinb(new_new_n8575__), .dout(new_new_n4865__));
  or1   g1767(.dina(new_new_n4865__), .dinb(new_new_n8576__), .dout(new_new_n4866__));
  or1   g1768(.dina(new_new_n8525__), .dinb(new_new_n8575__), .dout(new_new_n4867__));
  or1   g1769(.dina(new_new_n4867__), .dinb(new_new_n8577__), .dout(new_new_n4868__));
  and1  g1770(.dina(new_new_n4868__), .dinb(new_new_n4866__), .dout(new_new_n4869__));
  and1  g1771(.dina(new_new_n8538__), .dinb(new_new_n8577__), .dout(new_new_n4870__));
  and1  g1772(.dina(new_new_n8547__), .dinb(new_new_n8576__), .dout(new_new_n4871__));
  or1   g1773(.dina(new_new_n4871__), .dinb(new_new_n4870__), .dout(new_new_n4872__));
  or1   g1774(.dina(new_new_n4872__), .dinb(new_new_n3576__), .dout(new_new_n4873__));
  and1  g1775(.dina(new_new_n4873__), .dinb(new_new_n4869__), .dout(new_new_n4874__));
  or1   g1776(.dina(new_new_n8578__), .dinb(new_new_n8579__), .dout(new_new_n4875__));
  or1   g1777(.dina(new_new_n4875__), .dinb(new_new_n8580__), .dout(new_new_n4876__));
  or1   g1778(.dina(new_new_n4876__), .dinb(new_new_n8581__), .dout(new_new_n4877__));
  or1   g1779(.dina(new_new_n8516__), .dinb(new_new_n8582__), .dout(new_new_n4878__));
  or1   g1780(.dina(new_new_n4878__), .dinb(new_new_n8583__), .dout(new_new_n4879__));
  or1   g1781(.dina(new_new_n8528__), .dinb(new_new_n8582__), .dout(new_new_n4880__));
  or1   g1782(.dina(new_new_n4880__), .dinb(new_new_n8584__), .dout(new_new_n4881__));
  and1  g1783(.dina(new_new_n4881__), .dinb(new_new_n4879__), .dout(new_new_n4882__));
  and1  g1784(.dina(new_new_n8540__), .dinb(new_new_n8584__), .dout(new_new_n4883__));
  and1  g1785(.dina(new_new_n8550__), .dinb(new_new_n8583__), .dout(new_new_n4884__));
  or1   g1786(.dina(new_new_n4884__), .dinb(new_new_n4883__), .dout(new_new_n4885__));
  or1   g1787(.dina(new_new_n4885__), .dinb(new_new_n3540__), .dout(new_new_n4886__));
  and1  g1788(.dina(new_new_n4886__), .dinb(new_new_n4882__), .dout(new_new_n4887__));
  or1   g1789(.dina(new_new_n8516__), .dinb(new_new_n8585__), .dout(new_new_n4888__));
  or1   g1790(.dina(new_new_n4888__), .dinb(new_new_n8586__), .dout(new_new_n4889__));
  or1   g1791(.dina(new_new_n8528__), .dinb(new_new_n8585__), .dout(new_new_n4890__));
  or1   g1792(.dina(new_new_n4890__), .dinb(new_new_n8587__), .dout(new_new_n4891__));
  and1  g1793(.dina(new_new_n4891__), .dinb(new_new_n4889__), .dout(new_new_n4892__));
  and1  g1794(.dina(new_new_n8540__), .dinb(new_new_n8587__), .dout(new_new_n4893__));
  and1  g1795(.dina(new_new_n8550__), .dinb(new_new_n8586__), .dout(new_new_n4894__));
  or1   g1796(.dina(new_new_n4894__), .dinb(new_new_n4893__), .dout(new_new_n4895__));
  or1   g1797(.dina(new_new_n4895__), .dinb(new_new_n3556__), .dout(new_new_n4896__));
  and1  g1798(.dina(new_new_n4896__), .dinb(new_new_n4892__), .dout(new_new_n4897__));
  or1   g1799(.dina(new_new_n8517__), .dinb(new_new_n8588__), .dout(new_new_n4898__));
  or1   g1800(.dina(new_new_n4898__), .dinb(new_new_n8589__), .dout(new_new_n4899__));
  or1   g1801(.dina(new_new_n8529__), .dinb(new_new_n8588__), .dout(new_new_n4900__));
  or1   g1802(.dina(new_new_n4900__), .dinb(new_new_n8590__), .dout(new_new_n4901__));
  and1  g1803(.dina(new_new_n4901__), .dinb(new_new_n4899__), .dout(new_new_n4902__));
  and1  g1804(.dina(new_new_n8541__), .dinb(new_new_n8590__), .dout(new_new_n4903__));
  and1  g1805(.dina(new_new_n8551__), .dinb(new_new_n8589__), .dout(new_new_n4904__));
  or1   g1806(.dina(new_new_n4904__), .dinb(new_new_n4903__), .dout(new_new_n4905__));
  or1   g1807(.dina(new_new_n4905__), .dinb(new_new_n3554__), .dout(new_new_n4906__));
  and1  g1808(.dina(new_new_n4906__), .dinb(new_new_n4902__), .dout(new_new_n4907__));
  or1   g1809(.dina(new_new_n8517__), .dinb(new_new_n8591__), .dout(new_new_n4908__));
  or1   g1810(.dina(new_new_n4908__), .dinb(new_new_n8592__), .dout(new_new_n4909__));
  or1   g1811(.dina(new_new_n8529__), .dinb(new_new_n8591__), .dout(new_new_n4910__));
  or1   g1812(.dina(new_new_n4910__), .dinb(new_new_n8593__), .dout(new_new_n4911__));
  and1  g1813(.dina(new_new_n4911__), .dinb(new_new_n4909__), .dout(new_new_n4912__));
  and1  g1814(.dina(new_new_n8541__), .dinb(new_new_n8593__), .dout(new_new_n4913__));
  and1  g1815(.dina(new_new_n8551__), .dinb(new_new_n8592__), .dout(new_new_n4914__));
  or1   g1816(.dina(new_new_n4914__), .dinb(new_new_n4913__), .dout(new_new_n4915__));
  or1   g1817(.dina(new_new_n4915__), .dinb(new_new_n3552__), .dout(new_new_n4916__));
  and1  g1818(.dina(new_new_n4916__), .dinb(new_new_n4912__), .dout(new_new_n4917__));
  or1   g1819(.dina(new_new_n8594__), .dinb(new_new_n8595__), .dout(new_new_n4918__));
  or1   g1820(.dina(new_new_n4918__), .dinb(new_new_n8596__), .dout(new_new_n4919__));
  or1   g1821(.dina(new_new_n4919__), .dinb(new_new_n8597__), .dout(new_new_n4920__));
  or1   g1822(.dina(new_new_n4920__), .dinb(new_new_n4877__), .dout(new_new_n4921__));
  or1   g1823(.dina(new_new_n4921__), .dinb(new_new_n3989__), .dout(new_new_n4922__));
  or1   g1824(.dina(new_new_n3837__), .dinb(new_new_n8598__), .dout(new_new_n4923__));
  or1   g1825(.dina(new_new_n4923__), .dinb(new_new_n8600__), .dout(new_new_n4924__));
  or1   g1826(.dina(new_new_n4924__), .dinb(new_new_n8602__), .dout(new_new_n4925__));
  or1   g1827(.dina(new_new_n8604__), .dinb(new_new_n3993__), .dout(new_new_n4926__));
  or1   g1828(.dina(new_new_n8605__), .dinb(new_new_n8607__), .dout(new_new_n4927__));
  or1   g1829(.dina(new_new_n4927__), .dinb(new_new_n8610__), .dout(new_new_n4928__));
  or1   g1830(.dina(new_new_n4928__), .dinb(new_new_n8613__), .dout(new_new_n4929__));
  and1  g1831(.dina(new_new_n8619__), .dinb(new_new_n8625__), .dout(new_new_n4930__));
  or1   g1832(.dina(new_new_n8629__), .dinb(new_new_n8635__), .dout(new_new_n4931__));
  and1  g1833(.dina(new_new_n4930__), .dinb(new_new_n8638__), .dout(new_new_n4932__));
  or1   g1834(.dina(new_new_n4931__), .dinb(new_new_n8643__), .dout(new_new_n4933__));
  and1  g1835(.dina(new_new_n4932__), .dinb(new_new_n8648__), .dout(new_new_n4934__));
  or1   g1836(.dina(new_new_n4933__), .dinb(new_new_n8653__), .dout(new_new_n4935__));
  and1  g1837(.dina(new_new_n4934__), .dinb(new_new_n8658__), .dout(new_new_n4936__));
  or1   g1838(.dina(new_new_n4935__), .dinb(new_new_n8663__), .dout(new_new_n4937__));
  or1   g1839(.dina(new_new_n8666__), .dinb(new_new_n8667__), .dout(new_new_n4938__));
  or1   g1840(.dina(new_new_n3839__), .dinb(new_new_n8668__), .dout(new_new_n4939__));
  or1   g1841(.dina(new_new_n4939__), .dinb(new_new_n8670__), .dout(new_new_n4940__));
  or1   g1842(.dina(new_new_n4940__), .dinb(new_new_n8672__), .dout(new_new_n4941__));
  or1   g1843(.dina(new_new_n8674__), .dinb(new_new_n3995__), .dout(new_new_n4942__));
  or1   g1844(.dina(new_new_n8675__), .dinb(new_new_n8677__), .dout(new_new_n4943__));
  or1   g1845(.dina(new_new_n4943__), .dinb(new_new_n8680__), .dout(new_new_n4944__));
  or1   g1846(.dina(new_new_n4944__), .dinb(new_new_n8683__), .dout(new_new_n4945__));
  and1  g1847(.dina(new_new_n8688__), .dinb(new_new_n8694__), .dout(new_new_n4946__));
  or1   g1848(.dina(new_new_n8698__), .dinb(new_new_n8704__), .dout(new_new_n4947__));
  and1  g1849(.dina(new_new_n4946__), .dinb(new_new_n8707__), .dout(new_new_n4948__));
  or1   g1850(.dina(new_new_n4947__), .dinb(new_new_n8712__), .dout(new_new_n4949__));
  and1  g1851(.dina(new_new_n4948__), .dinb(new_new_n8717__), .dout(new_new_n4950__));
  or1   g1852(.dina(new_new_n4949__), .dinb(new_new_n8722__), .dout(new_new_n4951__));
  and1  g1853(.dina(new_new_n4950__), .dinb(new_new_n8727__), .dout(new_new_n4952__));
  or1   g1854(.dina(new_new_n4951__), .dinb(new_new_n8732__), .dout(new_new_n4953__));
  or1   g1855(.dina(new_new_n8735__), .dinb(new_new_n8736__), .dout(new_new_n4954__));
  and1  g1856(.dina(new_new_n4380__), .dinb(new_new_n4187__), .dout(new_new_n4955__));
  or1   g1857(.dina(new_new_n4381__), .dinb(new_new_n4186__), .dout(new_new_n4956__));
  and1  g1858(.dina(new_new_n4382__), .dinb(new_new_n4185__), .dout(new_new_n4957__));
  or1   g1859(.dina(new_new_n4383__), .dinb(new_new_n4184__), .dout(new_new_n4958__));
  and1  g1860(.dina(new_new_n4958__), .dinb(new_new_n4956__), .dout(new_new_n4959__));
  or1   g1861(.dina(new_new_n4957__), .dinb(new_new_n4955__), .dout(new_new_n4960__));
  and1  g1862(.dina(new_new_n4376__), .dinb(new_new_n4183__), .dout(new_new_n4961__));
  or1   g1863(.dina(new_new_n4377__), .dinb(new_new_n4182__), .dout(new_new_n4962__));
  and1  g1864(.dina(new_new_n4378__), .dinb(new_new_n4181__), .dout(new_new_n4963__));
  or1   g1865(.dina(new_new_n4379__), .dinb(new_new_n4180__), .dout(new_new_n4964__));
  and1  g1866(.dina(new_new_n4964__), .dinb(new_new_n4962__), .dout(new_new_n4965__));
  or1   g1867(.dina(new_new_n4963__), .dinb(new_new_n4961__), .dout(new_new_n4966__));
  and1  g1868(.dina(new_new_n8737__), .dinb(new_new_n8738__), .dout(new_new_n4967__));
  or1   g1869(.dina(new_new_n8739__), .dinb(new_new_n8740__), .dout(new_new_n4968__));
  and1  g1870(.dina(new_new_n8739__), .dinb(new_new_n8740__), .dout(new_new_n4969__));
  or1   g1871(.dina(new_new_n8737__), .dinb(new_new_n8738__), .dout(new_new_n4970__));
  and1  g1872(.dina(new_new_n4970__), .dinb(new_new_n4968__), .dout(new_new_n4971__));
  or1   g1873(.dina(new_new_n4969__), .dinb(new_new_n4967__), .dout(new_new_n4972__));
  and1  g1874(.dina(new_new_n4321__), .dinb(new_new_n4319__), .dout(new_new_n4973__));
  or1   g1875(.dina(new_new_n4320__), .dinb(new_new_n4318__), .dout(new_new_n4974__));
  and1  g1876(.dina(new_new_n4317__), .dinb(new_new_n4315__), .dout(new_new_n4975__));
  or1   g1877(.dina(new_new_n4316__), .dinb(new_new_n4314__), .dout(new_new_n4976__));
  and1  g1878(.dina(new_new_n8742__), .dinb(new_new_n8745__), .dout(new_new_n4977__));
  or1   g1879(.dina(new_new_n8748__), .dinb(new_new_n8751__), .dout(new_new_n4978__));
  and1  g1880(.dina(new_new_n4977__), .dinb(new_new_n8754__), .dout(new_new_n4979__));
  or1   g1881(.dina(new_new_n4978__), .dinb(new_new_n8757__), .dout(new_new_n4980__));
  and1  g1882(.dina(new_new_n8742__), .dinb(new_new_n8751__), .dout(new_new_n4981__));
  or1   g1883(.dina(new_new_n8748__), .dinb(new_new_n8745__), .dout(new_new_n4982__));
  and1  g1884(.dina(new_new_n4981__), .dinb(new_new_n8757__), .dout(new_new_n4983__));
  or1   g1885(.dina(new_new_n4982__), .dinb(new_new_n8754__), .dout(new_new_n4984__));
  and1  g1886(.dina(new_new_n4984__), .dinb(new_new_n4980__), .dout(new_new_n4985__));
  or1   g1887(.dina(new_new_n4983__), .dinb(new_new_n4979__), .dout(new_new_n4986__));
  and1  g1888(.dina(new_new_n8749__), .dinb(new_new_n8752__), .dout(new_new_n4987__));
  or1   g1889(.dina(new_new_n8743__), .dinb(new_new_n8746__), .dout(new_new_n4988__));
  and1  g1890(.dina(new_new_n4987__), .dinb(new_new_n8755__), .dout(new_new_n4989__));
  or1   g1891(.dina(new_new_n4988__), .dinb(new_new_n8758__), .dout(new_new_n4990__));
  and1  g1892(.dina(new_new_n8749__), .dinb(new_new_n8746__), .dout(new_new_n4991__));
  or1   g1893(.dina(new_new_n8743__), .dinb(new_new_n8752__), .dout(new_new_n4992__));
  and1  g1894(.dina(new_new_n4991__), .dinb(new_new_n8758__), .dout(new_new_n4993__));
  or1   g1895(.dina(new_new_n4992__), .dinb(new_new_n8755__), .dout(new_new_n4994__));
  and1  g1896(.dina(new_new_n4994__), .dinb(new_new_n4990__), .dout(new_new_n4995__));
  or1   g1897(.dina(new_new_n4993__), .dinb(new_new_n4989__), .dout(new_new_n4996__));
  and1  g1898(.dina(new_new_n4995__), .dinb(new_new_n4985__), .dout(new_new_n4997__));
  or1   g1899(.dina(new_new_n4996__), .dinb(new_new_n4986__), .dout(new_new_n4998__));
  and1  g1900(.dina(new_new_n4997__), .dinb(new_new_n4972__), .dout(new_new_n4999__));
  and1  g1901(.dina(new_new_n4998__), .dinb(new_new_n4971__), .dout(new_new_n5000__));
  or1   g1902(.dina(new_new_n5000__), .dinb(new_new_n4999__), .dout(new_new_n5001__));
  and1  g1903(.dina(new_new_n4372__), .dinb(new_new_n4179__), .dout(new_new_n5002__));
  or1   g1904(.dina(new_new_n4373__), .dinb(new_new_n4178__), .dout(new_new_n5003__));
  and1  g1905(.dina(new_new_n4374__), .dinb(new_new_n4177__), .dout(new_new_n5004__));
  or1   g1906(.dina(new_new_n4375__), .dinb(new_new_n4176__), .dout(new_new_n5005__));
  and1  g1907(.dina(new_new_n5005__), .dinb(new_new_n5003__), .dout(new_new_n5006__));
  or1   g1908(.dina(new_new_n5004__), .dinb(new_new_n5002__), .dout(new_new_n5007__));
  and1  g1909(.dina(new_new_n4403__), .dinb(new_new_n4175__), .dout(new_new_n5008__));
  or1   g1910(.dina(new_new_n4402__), .dinb(new_new_n4174__), .dout(new_new_n5009__));
  and1  g1911(.dina(new_new_n4370__), .dinb(new_new_n4208__), .dout(new_new_n5010__));
  or1   g1912(.dina(new_new_n4371__), .dinb(new_new_n4209__), .dout(new_new_n5011__));
  and1  g1913(.dina(new_new_n5011__), .dinb(new_new_n5009__), .dout(new_new_n5012__));
  or1   g1914(.dina(new_new_n5010__), .dinb(new_new_n5008__), .dout(new_new_n5013__));
  and1  g1915(.dina(new_new_n8759__), .dinb(new_new_n8760__), .dout(new_new_n5014__));
  or1   g1916(.dina(new_new_n8761__), .dinb(new_new_n8762__), .dout(new_new_n5015__));
  and1  g1917(.dina(new_new_n8761__), .dinb(new_new_n8762__), .dout(new_new_n5016__));
  or1   g1918(.dina(new_new_n8759__), .dinb(new_new_n8760__), .dout(new_new_n5017__));
  and1  g1919(.dina(new_new_n5017__), .dinb(new_new_n5015__), .dout(new_new_n5018__));
  or1   g1920(.dina(new_new_n5016__), .dinb(new_new_n5014__), .dout(new_new_n5019__));
  and1  g1921(.dina(new_new_n4313__), .dinb(new_new_n4311__), .dout(new_new_n5020__));
  or1   g1922(.dina(new_new_n4312__), .dinb(new_new_n4310__), .dout(new_new_n5021__));
  and1  g1923(.dina(new_new_n4309__), .dinb(new_new_n4307__), .dout(new_new_n5022__));
  or1   g1924(.dina(new_new_n4308__), .dinb(new_new_n4306__), .dout(new_new_n5023__));
  and1  g1925(.dina(new_new_n8764__), .dinb(new_new_n8767__), .dout(new_new_n5024__));
  or1   g1926(.dina(new_new_n8770__), .dinb(new_new_n8773__), .dout(new_new_n5025__));
  and1  g1927(.dina(new_new_n5024__), .dinb(new_new_n8776__), .dout(new_new_n5026__));
  or1   g1928(.dina(new_new_n5025__), .dinb(new_new_n8779__), .dout(new_new_n5027__));
  and1  g1929(.dina(new_new_n8764__), .dinb(new_new_n8773__), .dout(new_new_n5028__));
  or1   g1930(.dina(new_new_n8770__), .dinb(new_new_n8767__), .dout(new_new_n5029__));
  and1  g1931(.dina(new_new_n5028__), .dinb(new_new_n8779__), .dout(new_new_n5030__));
  or1   g1932(.dina(new_new_n5029__), .dinb(new_new_n8776__), .dout(new_new_n5031__));
  and1  g1933(.dina(new_new_n5031__), .dinb(new_new_n5027__), .dout(new_new_n5032__));
  or1   g1934(.dina(new_new_n5030__), .dinb(new_new_n5026__), .dout(new_new_n5033__));
  and1  g1935(.dina(new_new_n8771__), .dinb(new_new_n8774__), .dout(new_new_n5034__));
  or1   g1936(.dina(new_new_n8765__), .dinb(new_new_n8768__), .dout(new_new_n5035__));
  and1  g1937(.dina(new_new_n5034__), .dinb(new_new_n8777__), .dout(new_new_n5036__));
  or1   g1938(.dina(new_new_n5035__), .dinb(new_new_n8780__), .dout(new_new_n5037__));
  and1  g1939(.dina(new_new_n8771__), .dinb(new_new_n8768__), .dout(new_new_n5038__));
  or1   g1940(.dina(new_new_n8765__), .dinb(new_new_n8774__), .dout(new_new_n5039__));
  and1  g1941(.dina(new_new_n5038__), .dinb(new_new_n8780__), .dout(new_new_n5040__));
  or1   g1942(.dina(new_new_n5039__), .dinb(new_new_n8777__), .dout(new_new_n5041__));
  and1  g1943(.dina(new_new_n5041__), .dinb(new_new_n5037__), .dout(new_new_n5042__));
  or1   g1944(.dina(new_new_n5040__), .dinb(new_new_n5036__), .dout(new_new_n5043__));
  and1  g1945(.dina(new_new_n5042__), .dinb(new_new_n5032__), .dout(new_new_n5044__));
  or1   g1946(.dina(new_new_n5043__), .dinb(new_new_n5033__), .dout(new_new_n5045__));
  and1  g1947(.dina(new_new_n5044__), .dinb(new_new_n5019__), .dout(new_new_n5046__));
  and1  g1948(.dina(new_new_n5045__), .dinb(new_new_n5018__), .dout(new_new_n5047__));
  or1   g1949(.dina(new_new_n5047__), .dinb(new_new_n5046__), .dout(new_new_n5048__));
  or1   g1950(.dina(new_new_n3853__), .dinb(new_new_n8782__), .dout(new_new_n5049__));
  or1   g1951(.dina(new_new_n8602__), .dinb(new_new_n3845__), .dout(new_new_n5050__));
  or1   g1952(.dina(new_new_n8603__), .dinb(new_new_n8600__), .dout(new_new_n5051__));
  or1   g1953(.dina(new_new_n5051__), .dinb(new_new_n3833__), .dout(new_new_n5052__));
  or1   g1954(.dina(new_new_n8603__), .dinb(new_new_n8598__), .dout(new_new_n5053__));
  or1   g1955(.dina(new_new_n5053__), .dinb(new_new_n3825__), .dout(new_new_n5054__));
  or1   g1956(.dina(new_new_n5054__), .dinb(new_new_n8599__), .dout(new_new_n5055__));
  and1  g1957(.dina(new_new_n5050__), .dinb(new_new_n8783__), .dout(new_new_n5056__));
  and1  g1958(.dina(new_new_n5056__), .dinb(new_new_n5052__), .dout(new_new_n5057__));
  and1  g1959(.dina(new_new_n5057__), .dinb(new_new_n5055__), .dout(new_new_n5058__));
  or1   g1960(.dina(new_new_n8604__), .dinb(new_new_n4001__), .dout(new_new_n5059__));
  and1  g1961(.dina(new_new_n5059__), .dinb(new_new_n5058__), .dout(new_new_n5060__));
  or1   g1962(.dina(new_new_n8613__), .dinb(new_new_n8784__), .dout(new_new_n5061__));
  or1   g1963(.dina(new_new_n8614__), .dinb(new_new_n8607__), .dout(new_new_n5062__));
  or1   g1964(.dina(new_new_n5062__), .dinb(new_new_n8785__), .dout(new_new_n5063__));
  or1   g1965(.dina(new_new_n8614__), .dinb(new_new_n8610__), .dout(new_new_n5064__));
  or1   g1966(.dina(new_new_n5064__), .dinb(new_new_n8786__), .dout(new_new_n5065__));
  or1   g1967(.dina(new_new_n5065__), .dinb(new_new_n8608__), .dout(new_new_n5066__));
  and1  g1968(.dina(new_new_n5061__), .dinb(new_new_n8788__), .dout(new_new_n5067__));
  and1  g1969(.dina(new_new_n5067__), .dinb(new_new_n5063__), .dout(new_new_n5068__));
  and1  g1970(.dina(new_new_n5068__), .dinb(new_new_n5066__), .dout(new_new_n5069__));
  and1  g1971(.dina(new_new_n3850__), .dinb(new_new_n8559__), .dout(new_new_n5070__));
  or1   g1972(.dina(new_new_n3851__), .dinb(new_new_n8555__), .dout(new_new_n5071__));
  and1  g1973(.dina(new_new_n8648__), .dinb(new_new_n8790__), .dout(new_new_n5072__));
  or1   g1974(.dina(new_new_n8653__), .dinb(new_new_n8791__), .dout(new_new_n5073__));
  and1  g1975(.dina(new_new_n8619__), .dinb(new_new_n8649__), .dout(new_new_n5074__));
  or1   g1976(.dina(new_new_n8629__), .dinb(new_new_n8654__), .dout(new_new_n5075__));
  and1  g1977(.dina(new_new_n5074__), .dinb(new_new_n8793__), .dout(new_new_n5076__));
  or1   g1978(.dina(new_new_n5075__), .dinb(new_new_n8795__), .dout(new_new_n5077__));
  and1  g1979(.dina(new_new_n8638__), .dinb(new_new_n8649__), .dout(new_new_n5078__));
  or1   g1980(.dina(new_new_n8643__), .dinb(new_new_n8654__), .dout(new_new_n5079__));
  and1  g1981(.dina(new_new_n5078__), .dinb(new_new_n8797__), .dout(new_new_n5080__));
  or1   g1982(.dina(new_new_n5079__), .dinb(new_new_n8799__), .dout(new_new_n5081__));
  and1  g1983(.dina(new_new_n5080__), .dinb(new_new_n8618__), .dout(new_new_n5082__));
  or1   g1984(.dina(new_new_n5081__), .dinb(new_new_n8628__), .dout(new_new_n5083__));
  and1  g1985(.dina(new_new_n8658__), .dinb(new_new_n8639__), .dout(new_new_n5084__));
  or1   g1986(.dina(new_new_n8663__), .dinb(new_new_n8644__), .dout(new_new_n5085__));
  and1  g1987(.dina(new_new_n8800__), .dinb(new_new_n8650__), .dout(new_new_n5086__));
  or1   g1988(.dina(new_new_n8801__), .dinb(new_new_n8655__), .dout(new_new_n5087__));
  and1  g1989(.dina(new_new_n5086__), .dinb(new_new_n8803__), .dout(new_new_n5088__));
  or1   g1990(.dina(new_new_n5087__), .dinb(new_new_n8806__), .dout(new_new_n5089__));
  and1  g1991(.dina(new_new_n5088__), .dinb(new_new_n8620__), .dout(new_new_n5090__));
  or1   g1992(.dina(new_new_n5089__), .dinb(new_new_n8630__), .dout(new_new_n5091__));
  and1  g1993(.dina(new_new_n5073__), .dinb(new_new_n5071__), .dout(new_new_n5092__));
  or1   g1994(.dina(new_new_n5072__), .dinb(new_new_n5070__), .dout(new_new_n5093__));
  and1  g1995(.dina(new_new_n5092__), .dinb(new_new_n5077__), .dout(new_new_n5094__));
  or1   g1996(.dina(new_new_n5093__), .dinb(new_new_n5076__), .dout(new_new_n5095__));
  and1  g1997(.dina(new_new_n5094__), .dinb(new_new_n5083__), .dout(new_new_n5096__));
  or1   g1998(.dina(new_new_n5095__), .dinb(new_new_n5082__), .dout(new_new_n5097__));
  and1  g1999(.dina(new_new_n5096__), .dinb(new_new_n5091__), .dout(new_new_n5098__));
  or1   g2000(.dina(new_new_n5097__), .dinb(new_new_n5090__), .dout(new_new_n5099__));
  or1   g2001(.dina(new_new_n8808__), .dinb(new_new_n8667__), .dout(new_new_n5100__));
  and1  g2002(.dina(new_new_n5100__), .dinb(new_new_n5069__), .dout(new_new_n5101__));
  or1   g2003(.dina(new_new_n8683__), .dinb(new_new_n8809__), .dout(new_new_n5102__));
  or1   g2004(.dina(new_new_n8682__), .dinb(new_new_n8677__), .dout(new_new_n5103__));
  or1   g2005(.dina(new_new_n5103__), .dinb(new_new_n8810__), .dout(new_new_n5104__));
  or1   g2006(.dina(new_new_n8684__), .dinb(new_new_n8680__), .dout(new_new_n5105__));
  or1   g2007(.dina(new_new_n5105__), .dinb(new_new_n8811__), .dout(new_new_n5106__));
  or1   g2008(.dina(new_new_n5106__), .dinb(new_new_n8678__), .dout(new_new_n5107__));
  and1  g2009(.dina(new_new_n5102__), .dinb(new_new_n8783__), .dout(new_new_n5108__));
  and1  g2010(.dina(new_new_n5108__), .dinb(new_new_n5104__), .dout(new_new_n5109__));
  and1  g2011(.dina(new_new_n5109__), .dinb(new_new_n5107__), .dout(new_new_n5110__));
  and1  g2012(.dina(new_new_n3848__), .dinb(new_new_n8568__), .dout(new_new_n5111__));
  or1   g2013(.dina(new_new_n3849__), .dinb(new_new_n8564__), .dout(new_new_n5112__));
  and1  g2014(.dina(new_new_n8717__), .dinb(new_new_n8812__), .dout(new_new_n5113__));
  or1   g2015(.dina(new_new_n8722__), .dinb(new_new_n8813__), .dout(new_new_n5114__));
  and1  g2016(.dina(new_new_n8718__), .dinb(new_new_n8688__), .dout(new_new_n5115__));
  or1   g2017(.dina(new_new_n8723__), .dinb(new_new_n8698__), .dout(new_new_n5116__));
  and1  g2018(.dina(new_new_n5115__), .dinb(new_new_n8815__), .dout(new_new_n5117__));
  or1   g2019(.dina(new_new_n5116__), .dinb(new_new_n8817__), .dout(new_new_n5118__));
  and1  g2020(.dina(new_new_n8718__), .dinb(new_new_n8707__), .dout(new_new_n5119__));
  or1   g2021(.dina(new_new_n8723__), .dinb(new_new_n8712__), .dout(new_new_n5120__));
  and1  g2022(.dina(new_new_n5119__), .dinb(new_new_n8819__), .dout(new_new_n5121__));
  or1   g2023(.dina(new_new_n5120__), .dinb(new_new_n8821__), .dout(new_new_n5122__));
  and1  g2024(.dina(new_new_n5121__), .dinb(new_new_n8687__), .dout(new_new_n5123__));
  or1   g2025(.dina(new_new_n5122__), .dinb(new_new_n8697__), .dout(new_new_n5124__));
  and1  g2026(.dina(new_new_n8727__), .dinb(new_new_n8708__), .dout(new_new_n5125__));
  or1   g2027(.dina(new_new_n8732__), .dinb(new_new_n8713__), .dout(new_new_n5126__));
  and1  g2028(.dina(new_new_n8822__), .dinb(new_new_n8719__), .dout(new_new_n5127__));
  or1   g2029(.dina(new_new_n8823__), .dinb(new_new_n8724__), .dout(new_new_n5128__));
  and1  g2030(.dina(new_new_n5127__), .dinb(new_new_n8825__), .dout(new_new_n5129__));
  or1   g2031(.dina(new_new_n5128__), .dinb(new_new_n8828__), .dout(new_new_n5130__));
  and1  g2032(.dina(new_new_n5129__), .dinb(new_new_n8689__), .dout(new_new_n5131__));
  or1   g2033(.dina(new_new_n5130__), .dinb(new_new_n8699__), .dout(new_new_n5132__));
  and1  g2034(.dina(new_new_n5114__), .dinb(new_new_n5112__), .dout(new_new_n5133__));
  or1   g2035(.dina(new_new_n5113__), .dinb(new_new_n5111__), .dout(new_new_n5134__));
  and1  g2036(.dina(new_new_n5133__), .dinb(new_new_n5118__), .dout(new_new_n5135__));
  or1   g2037(.dina(new_new_n5134__), .dinb(new_new_n5117__), .dout(new_new_n5136__));
  and1  g2038(.dina(new_new_n5135__), .dinb(new_new_n5124__), .dout(new_new_n5137__));
  or1   g2039(.dina(new_new_n5136__), .dinb(new_new_n5123__), .dout(new_new_n5138__));
  and1  g2040(.dina(new_new_n5137__), .dinb(new_new_n5132__), .dout(new_new_n5139__));
  or1   g2041(.dina(new_new_n5138__), .dinb(new_new_n5131__), .dout(new_new_n5140__));
  or1   g2042(.dina(new_new_n8830__), .dinb(new_new_n8736__), .dout(new_new_n5141__));
  and1  g2043(.dina(new_new_n5141__), .dinb(new_new_n5110__), .dout(new_new_n5142__));
  or1   g2044(.dina(new_new_n8672__), .dinb(new_new_n3846__), .dout(new_new_n5143__));
  or1   g2045(.dina(new_new_n8673__), .dinb(new_new_n8670__), .dout(new_new_n5144__));
  or1   g2046(.dina(new_new_n5144__), .dinb(new_new_n3835__), .dout(new_new_n5145__));
  or1   g2047(.dina(new_new_n8673__), .dinb(new_new_n8668__), .dout(new_new_n5146__));
  or1   g2048(.dina(new_new_n5146__), .dinb(new_new_n3827__), .dout(new_new_n5147__));
  or1   g2049(.dina(new_new_n5147__), .dinb(new_new_n8669__), .dout(new_new_n5148__));
  and1  g2050(.dina(new_new_n5143__), .dinb(new_new_n8788__), .dout(new_new_n5149__));
  and1  g2051(.dina(new_new_n5149__), .dinb(new_new_n5145__), .dout(new_new_n5150__));
  and1  g2052(.dina(new_new_n5150__), .dinb(new_new_n5148__), .dout(new_new_n5151__));
  or1   g2053(.dina(new_new_n8674__), .dinb(new_new_n4003__), .dout(new_new_n5152__));
  and1  g2054(.dina(new_new_n5152__), .dinb(new_new_n5151__), .dout(new_new_n5153__));
  or1   g2055(.dina(new_new_n8831__), .dinb(new_new_n3516__), .dout(new_new_n5154__));
  or1   g2056(.dina(new_new_n8832__), .dinb(new_new_n3517__), .dout(new_new_n5155__));
  and1  g2057(.dina(new_new_n5155__), .dinb(new_new_n5154__), .dout(new_new_n5156__));
  and1  g2058(.dina(new_new_n5156__), .dinb(new_new_n8838__), .dout(new_new_n5157__));
  and1  g2059(.dina(new_new_n5157__), .dinb(new_new_n8878__), .dout(new_new_n5158__));
  and1  g2060(.dina(new_new_n8635__), .dinb(new_new_n8914__), .dout(new_new_n5159__));
  and1  g2061(.dina(new_new_n8625__), .dinb(new_new_n8916__), .dout(new_new_n5160__));
  or1   g2062(.dina(new_new_n5160__), .dinb(new_new_n5159__), .dout(new_new_n5161__));
  and1  g2063(.dina(new_new_n8917__), .dinb(new_new_n8922__), .dout(new_new_n5162__));
  and1  g2064(.dina(new_new_n5162__), .dinb(new_new_n8878__), .dout(new_new_n5163__));
  and1  g2065(.dina(new_new_n8838__), .dinb(new_new_n3162__), .dout(new_new_n5164__));
  and1  g2066(.dina(new_new_n5164__), .dinb(new_new_n8945__), .dout(new_new_n5165__));
  or1   g2067(.dina(new_new_n5163__), .dinb(new_new_n5158__), .dout(new_new_n5166__));
  or1   g2068(.dina(new_new_n5166__), .dinb(new_new_n5165__), .dout(new_new_n5167__));
  and1  g2069(.dina(new_new_n8561__), .dinb(new_new_n8839__), .dout(new_new_n5168__));
  and1  g2070(.dina(new_new_n5168__), .dinb(new_new_n8879__), .dout(new_new_n5169__));
  and1  g2071(.dina(new_new_n8624__), .dinb(new_new_n8914__), .dout(new_new_n5170__));
  or1   g2072(.dina(new_new_n8634__), .dinb(new_new_n8916__), .dout(new_new_n5171__));
  and1  g2073(.dina(new_new_n8965__), .dinb(new_new_n8806__), .dout(new_new_n5172__));
  or1   g2074(.dina(new_new_n8967__), .dinb(new_new_n8803__), .dout(new_new_n5173__));
  and1  g2075(.dina(new_new_n5172__), .dinb(new_new_n8664__), .dout(new_new_n5174__));
  and1  g2076(.dina(new_new_n5173__), .dinb(new_new_n8659__), .dout(new_new_n5175__));
  or1   g2077(.dina(new_new_n5175__), .dinb(new_new_n5174__), .dout(new_new_n5176__));
  and1  g2078(.dina(new_new_n8968__), .dinb(new_new_n8922__), .dout(new_new_n5177__));
  and1  g2079(.dina(new_new_n5177__), .dinb(new_new_n8879__), .dout(new_new_n5178__));
  and1  g2080(.dina(new_new_n8839__), .dinb(new_new_n3146__), .dout(new_new_n5179__));
  and1  g2081(.dina(new_new_n5179__), .dinb(new_new_n8945__), .dout(new_new_n5180__));
  or1   g2082(.dina(new_new_n5178__), .dinb(new_new_n5169__), .dout(new_new_n5181__));
  or1   g2083(.dina(new_new_n5181__), .dinb(new_new_n5180__), .dout(new_new_n5182__));
  and1  g2084(.dina(new_new_n8595__), .dinb(new_new_n8841__), .dout(new_new_n5183__));
  and1  g2085(.dina(new_new_n5183__), .dinb(new_new_n8881__), .dout(new_new_n5184__));
  and1  g2086(.dina(new_new_n8704__), .dinb(new_new_n8970__), .dout(new_new_n5185__));
  and1  g2087(.dina(new_new_n8694__), .dinb(new_new_n8972__), .dout(new_new_n5186__));
  or1   g2088(.dina(new_new_n5186__), .dinb(new_new_n5185__), .dout(new_new_n5187__));
  and1  g2089(.dina(new_new_n8973__), .dinb(new_new_n8923__), .dout(new_new_n5188__));
  and1  g2090(.dina(new_new_n5188__), .dinb(new_new_n8881__), .dout(new_new_n5189__));
  and1  g2091(.dina(new_new_n8841__), .dinb(new_new_n3066__), .dout(new_new_n5190__));
  and1  g2092(.dina(new_new_n5190__), .dinb(new_new_n8946__), .dout(new_new_n5191__));
  or1   g2093(.dina(new_new_n5189__), .dinb(new_new_n5184__), .dout(new_new_n5192__));
  or1   g2094(.dina(new_new_n5192__), .dinb(new_new_n5191__), .dout(new_new_n5193__));
  and1  g2095(.dina(new_new_n8974__), .dinb(new_new_n8975__), .dout(new_new_n5194__));
  or1   g2096(.dina(new_new_n8976__), .dinb(new_new_n8977__), .dout(new_new_n5195__));
  and1  g2097(.dina(new_new_n8976__), .dinb(new_new_n8977__), .dout(new_new_n5196__));
  or1   g2098(.dina(new_new_n8974__), .dinb(new_new_n8975__), .dout(new_new_n5197__));
  and1  g2099(.dina(new_new_n5197__), .dinb(new_new_n5195__), .dout(new_new_n5198__));
  or1   g2100(.dina(new_new_n5196__), .dinb(new_new_n5194__), .dout(new_new_n5199__));
  and1  g2101(.dina(new_new_n4936__), .dinb(new_new_n8913__), .dout(new_new_n5200__));
  or1   g2102(.dina(new_new_n8666__), .dinb(new_new_n8915__), .dout(new_new_n5201__));
  and1  g2103(.dina(new_new_n5201__), .dinb(new_new_n8808__), .dout(new_new_n5202__));
  or1   g2104(.dina(new_new_n5200__), .dinb(new_new_n5099__), .dout(new_new_n5203__));
  and1  g2105(.dina(new_new_n8980__), .dinb(new_new_n5198__), .dout(new_new_n5204__));
  or1   g2106(.dina(new_new_n8984__), .dinb(new_new_n5199__), .dout(new_new_n5205__));
  and1  g2107(.dina(new_new_n4331__), .dinb(new_new_n8784__), .dout(new_new_n5206__));
  or1   g2108(.dina(new_new_n4330__), .dinb(new_new_n4205__), .dout(new_new_n5207__));
  and1  g2109(.dina(new_new_n5206__), .dinb(new_new_n4335__), .dout(new_new_n5208__));
  or1   g2110(.dina(new_new_n5207__), .dinb(new_new_n4334__), .dout(new_new_n5209__));
  and1  g2111(.dina(new_new_n5208__), .dinb(new_new_n4353__), .dout(new_new_n5210__));
  or1   g2112(.dina(new_new_n5209__), .dinb(new_new_n4352__), .dout(new_new_n5211__));
  and1  g2113(.dina(new_new_n8986__), .dinb(new_new_n8615__), .dout(new_new_n5212__));
  or1   g2114(.dina(new_new_n8987__), .dinb(new_new_n8988__), .dout(new_new_n5213__));
  and1  g2115(.dina(new_new_n8987__), .dinb(new_new_n8988__), .dout(new_new_n5214__));
  or1   g2116(.dina(new_new_n8986__), .dinb(new_new_n8615__), .dout(new_new_n5215__));
  and1  g2117(.dina(new_new_n5215__), .dinb(new_new_n5213__), .dout(new_new_n5216__));
  or1   g2118(.dina(new_new_n5214__), .dinb(new_new_n5212__), .dout(new_new_n5217__));
  and1  g2119(.dina(new_new_n5217__), .dinb(new_new_n8984__), .dout(new_new_n5218__));
  or1   g2120(.dina(new_new_n5216__), .dinb(new_new_n8980__), .dout(new_new_n5219__));
  and1  g2121(.dina(new_new_n5219__), .dinb(new_new_n5205__), .dout(new_new_n5220__));
  or1   g2122(.dina(new_new_n5218__), .dinb(new_new_n5204__), .dout(new_new_n5221__));
  and1  g2123(.dina(new_new_n8991__), .dinb(new_new_n8997__), .dout(new_new_n5222__));
  and1  g2124(.dina(new_new_n5222__), .dinb(new_new_n9016__), .dout(new_new_n5223__));
  and1  g2125(.dina(new_new_n9033__), .dinb(new_new_n9039__), .dout(new_new_n5224__));
  and1  g2126(.dina(new_new_n5224__), .dinb(new_new_n9016__), .dout(new_new_n5225__));
  and1  g2127(.dina(new_new_n8997__), .dinb(new_new_n9054__), .dout(new_new_n5226__));
  and1  g2128(.dina(new_new_n5226__), .dinb(new_new_n9059__), .dout(new_new_n5227__));
  and1  g2129(.dina(new_new_n9039__), .dinb(new_new_n9074__), .dout(new_new_n5228__));
  and1  g2130(.dina(new_new_n5228__), .dinb(new_new_n9059__), .dout(new_new_n5229__));
  or1   g2131(.dina(new_new_n5225__), .dinb(new_new_n5223__), .dout(new_new_n5230__));
  or1   g2132(.dina(new_new_n5230__), .dinb(new_new_n5227__), .dout(new_new_n5231__));
  or1   g2133(.dina(new_new_n5231__), .dinb(new_new_n5229__), .dout(new_new_n5232__));
  and1  g2134(.dina(new_new_n8563__), .dinb(new_new_n8842__), .dout(new_new_n5233__));
  and1  g2135(.dina(new_new_n5233__), .dinb(new_new_n8882__), .dout(new_new_n5234__));
  and1  g2136(.dina(new_new_n8620__), .dinb(new_new_n8793__), .dout(new_new_n5235__));
  or1   g2137(.dina(new_new_n8630__), .dinb(new_new_n8795__), .dout(new_new_n5236__));
  and1  g2138(.dina(new_new_n8639__), .dinb(new_new_n8797__), .dout(new_new_n5237__));
  or1   g2139(.dina(new_new_n8644__), .dinb(new_new_n8799__), .dout(new_new_n5238__));
  and1  g2140(.dina(new_new_n9075__), .dinb(new_new_n8622__), .dout(new_new_n5239__));
  or1   g2141(.dina(new_new_n9076__), .dinb(new_new_n8632__), .dout(new_new_n5240__));
  and1  g2142(.dina(new_new_n8800__), .dinb(new_new_n8804__), .dout(new_new_n5241__));
  or1   g2143(.dina(new_new_n8801__), .dinb(new_new_n8807__), .dout(new_new_n5242__));
  and1  g2144(.dina(new_new_n9077__), .dinb(new_new_n8622__), .dout(new_new_n5243__));
  or1   g2145(.dina(new_new_n9078__), .dinb(new_new_n8632__), .dout(new_new_n5244__));
  and1  g2146(.dina(new_new_n8967__), .dinb(new_new_n8640__), .dout(new_new_n5245__));
  or1   g2147(.dina(new_new_n8965__), .dinb(new_new_n8645__), .dout(new_new_n5246__));
  and1  g2148(.dina(new_new_n5245__), .dinb(new_new_n8659__), .dout(new_new_n5247__));
  or1   g2149(.dina(new_new_n5246__), .dinb(new_new_n8664__), .dout(new_new_n5248__));
  and1  g2150(.dina(new_new_n9079__), .dinb(new_new_n8623__), .dout(new_new_n5249__));
  or1   g2151(.dina(new_new_n9080__), .dinb(new_new_n8633__), .dout(new_new_n5250__));
  and1  g2152(.dina(new_new_n5236__), .dinb(new_new_n8791__), .dout(new_new_n5251__));
  or1   g2153(.dina(new_new_n5235__), .dinb(new_new_n8790__), .dout(new_new_n5252__));
  and1  g2154(.dina(new_new_n5251__), .dinb(new_new_n5240__), .dout(new_new_n5253__));
  or1   g2155(.dina(new_new_n5252__), .dinb(new_new_n5239__), .dout(new_new_n5254__));
  and1  g2156(.dina(new_new_n5253__), .dinb(new_new_n5244__), .dout(new_new_n5255__));
  or1   g2157(.dina(new_new_n5254__), .dinb(new_new_n5243__), .dout(new_new_n5256__));
  and1  g2158(.dina(new_new_n5255__), .dinb(new_new_n5250__), .dout(new_new_n5257__));
  or1   g2159(.dina(new_new_n5256__), .dinb(new_new_n5249__), .dout(new_new_n5258__));
  and1  g2160(.dina(new_new_n5257__), .dinb(new_new_n8655__), .dout(new_new_n5259__));
  and1  g2161(.dina(new_new_n5258__), .dinb(new_new_n8650__), .dout(new_new_n5260__));
  or1   g2162(.dina(new_new_n5260__), .dinb(new_new_n5259__), .dout(new_new_n5261__));
  and1  g2163(.dina(new_new_n9081__), .dinb(new_new_n8923__), .dout(new_new_n5262__));
  and1  g2164(.dina(new_new_n5262__), .dinb(new_new_n8882__), .dout(new_new_n5263__));
  and1  g2165(.dina(new_new_n8842__), .dinb(new_new_n2834__), .dout(new_new_n5264__));
  and1  g2166(.dina(new_new_n5264__), .dinb(new_new_n8946__), .dout(new_new_n5265__));
  or1   g2167(.dina(new_new_n5263__), .dinb(new_new_n5234__), .dout(new_new_n5266__));
  or1   g2168(.dina(new_new_n5266__), .dinb(new_new_n5265__), .dout(new_new_n5267__));
  and1  g2169(.dina(new_new_n8562__), .dinb(new_new_n8845__), .dout(new_new_n5268__));
  and1  g2170(.dina(new_new_n5268__), .dinb(new_new_n8885__), .dout(new_new_n5269__));
  and1  g2171(.dina(new_new_n9076__), .dinb(new_new_n8794__), .dout(new_new_n5270__));
  or1   g2172(.dina(new_new_n9075__), .dinb(new_new_n8792__), .dout(new_new_n5271__));
  and1  g2173(.dina(new_new_n5270__), .dinb(new_new_n9078__), .dout(new_new_n5272__));
  or1   g2174(.dina(new_new_n5271__), .dinb(new_new_n9077__), .dout(new_new_n5273__));
  and1  g2175(.dina(new_new_n5272__), .dinb(new_new_n9080__), .dout(new_new_n5274__));
  or1   g2176(.dina(new_new_n5273__), .dinb(new_new_n9079__), .dout(new_new_n5275__));
  and1  g2177(.dina(new_new_n5274__), .dinb(new_new_n8633__), .dout(new_new_n5276__));
  and1  g2178(.dina(new_new_n5275__), .dinb(new_new_n8623__), .dout(new_new_n5277__));
  or1   g2179(.dina(new_new_n5277__), .dinb(new_new_n5276__), .dout(new_new_n5278__));
  and1  g2180(.dina(new_new_n9082__), .dinb(new_new_n8925__), .dout(new_new_n5279__));
  and1  g2181(.dina(new_new_n5279__), .dinb(new_new_n8885__), .dout(new_new_n5280__));
  and1  g2182(.dina(new_new_n8845__), .dinb(new_new_n3154__), .dout(new_new_n5281__));
  and1  g2183(.dina(new_new_n5281__), .dinb(new_new_n8948__), .dout(new_new_n5282__));
  or1   g2184(.dina(new_new_n5280__), .dinb(new_new_n5269__), .dout(new_new_n5283__));
  or1   g2185(.dina(new_new_n5283__), .dinb(new_new_n5282__), .dout(new_new_n5284__));
  and1  g2186(.dina(new_new_n8560__), .dinb(new_new_n8846__), .dout(new_new_n5285__));
  and1  g2187(.dina(new_new_n5285__), .dinb(new_new_n8886__), .dout(new_new_n5286__));
  and1  g2188(.dina(new_new_n8660__), .dinb(new_new_n8804__), .dout(new_new_n5287__));
  or1   g2189(.dina(new_new_n8665__), .dinb(new_new_n8807__), .dout(new_new_n5288__));
  and1  g2190(.dina(new_new_n8966__), .dinb(new_new_n8660__), .dout(new_new_n5289__));
  or1   g2191(.dina(new_new_n8964__), .dinb(new_new_n8665__), .dout(new_new_n5290__));
  and1  g2192(.dina(new_new_n5288__), .dinb(new_new_n8798__), .dout(new_new_n5291__));
  or1   g2193(.dina(new_new_n5287__), .dinb(new_new_n8796__), .dout(new_new_n5292__));
  and1  g2194(.dina(new_new_n5291__), .dinb(new_new_n5290__), .dout(new_new_n5293__));
  or1   g2195(.dina(new_new_n5292__), .dinb(new_new_n5289__), .dout(new_new_n5294__));
  and1  g2196(.dina(new_new_n5293__), .dinb(new_new_n8645__), .dout(new_new_n5295__));
  and1  g2197(.dina(new_new_n5294__), .dinb(new_new_n8640__), .dout(new_new_n5296__));
  or1   g2198(.dina(new_new_n5296__), .dinb(new_new_n5295__), .dout(new_new_n5297__));
  and1  g2199(.dina(new_new_n9083__), .dinb(new_new_n8925__), .dout(new_new_n5298__));
  and1  g2200(.dina(new_new_n5298__), .dinb(new_new_n8886__), .dout(new_new_n5299__));
  and1  g2201(.dina(new_new_n8846__), .dinb(new_new_n3082__), .dout(new_new_n5300__));
  and1  g2202(.dina(new_new_n5300__), .dinb(new_new_n8948__), .dout(new_new_n5301__));
  or1   g2203(.dina(new_new_n5299__), .dinb(new_new_n5286__), .dout(new_new_n5302__));
  or1   g2204(.dina(new_new_n5302__), .dinb(new_new_n5301__), .dout(new_new_n5303__));
  and1  g2205(.dina(new_new_n8991__), .dinb(new_new_n9088__), .dout(new_new_n5304__));
  and1  g2206(.dina(new_new_n5304__), .dinb(new_new_n9107__), .dout(new_new_n5305__));
  and1  g2207(.dina(new_new_n9033__), .dinb(new_new_n9126__), .dout(new_new_n5306__));
  and1  g2208(.dina(new_new_n5306__), .dinb(new_new_n9107__), .dout(new_new_n5307__));
  and1  g2209(.dina(new_new_n9088__), .dinb(new_new_n9054__), .dout(new_new_n5308__));
  and1  g2210(.dina(new_new_n5308__), .dinb(new_new_n9145__), .dout(new_new_n5309__));
  and1  g2211(.dina(new_new_n9126__), .dinb(new_new_n9074__), .dout(new_new_n5310__));
  and1  g2212(.dina(new_new_n5310__), .dinb(new_new_n9145__), .dout(new_new_n5311__));
  or1   g2213(.dina(new_new_n5307__), .dinb(new_new_n5305__), .dout(new_new_n5312__));
  or1   g2214(.dina(new_new_n5312__), .dinb(new_new_n5309__), .dout(new_new_n5313__));
  or1   g2215(.dina(new_new_n5313__), .dinb(new_new_n5311__), .dout(new_new_n5314__));
  and1  g2216(.dina(new_new_n8579__), .dinb(new_new_n8848__), .dout(new_new_n5315__));
  and1  g2217(.dina(new_new_n5315__), .dinb(new_new_n8888__), .dout(new_new_n5316__));
  and1  g2218(.dina(new_new_n8689__), .dinb(new_new_n8815__), .dout(new_new_n5317__));
  or1   g2219(.dina(new_new_n8699__), .dinb(new_new_n8817__), .dout(new_new_n5318__));
  and1  g2220(.dina(new_new_n8708__), .dinb(new_new_n8819__), .dout(new_new_n5319__));
  or1   g2221(.dina(new_new_n8713__), .dinb(new_new_n8821__), .dout(new_new_n5320__));
  and1  g2222(.dina(new_new_n9160__), .dinb(new_new_n8691__), .dout(new_new_n5321__));
  or1   g2223(.dina(new_new_n9161__), .dinb(new_new_n8701__), .dout(new_new_n5322__));
  and1  g2224(.dina(new_new_n8822__), .dinb(new_new_n8825__), .dout(new_new_n5323__));
  or1   g2225(.dina(new_new_n8823__), .dinb(new_new_n8828__), .dout(new_new_n5324__));
  and1  g2226(.dina(new_new_n9162__), .dinb(new_new_n8691__), .dout(new_new_n5325__));
  or1   g2227(.dina(new_new_n9163__), .dinb(new_new_n8701__), .dout(new_new_n5326__));
  and1  g2228(.dina(new_new_n8693__), .dinb(new_new_n8970__), .dout(new_new_n5327__));
  or1   g2229(.dina(new_new_n8703__), .dinb(new_new_n8972__), .dout(new_new_n5328__));
  and1  g2230(.dina(new_new_n9165__), .dinb(new_new_n8709__), .dout(new_new_n5329__));
  or1   g2231(.dina(new_new_n9167__), .dinb(new_new_n8714__), .dout(new_new_n5330__));
  and1  g2232(.dina(new_new_n5329__), .dinb(new_new_n8728__), .dout(new_new_n5331__));
  or1   g2233(.dina(new_new_n5330__), .dinb(new_new_n8733__), .dout(new_new_n5332__));
  and1  g2234(.dina(new_new_n9168__), .dinb(new_new_n8692__), .dout(new_new_n5333__));
  or1   g2235(.dina(new_new_n9169__), .dinb(new_new_n8702__), .dout(new_new_n5334__));
  and1  g2236(.dina(new_new_n5318__), .dinb(new_new_n8813__), .dout(new_new_n5335__));
  or1   g2237(.dina(new_new_n5317__), .dinb(new_new_n8812__), .dout(new_new_n5336__));
  and1  g2238(.dina(new_new_n5335__), .dinb(new_new_n5322__), .dout(new_new_n5337__));
  or1   g2239(.dina(new_new_n5336__), .dinb(new_new_n5321__), .dout(new_new_n5338__));
  and1  g2240(.dina(new_new_n5337__), .dinb(new_new_n5326__), .dout(new_new_n5339__));
  or1   g2241(.dina(new_new_n5338__), .dinb(new_new_n5325__), .dout(new_new_n5340__));
  and1  g2242(.dina(new_new_n5339__), .dinb(new_new_n5334__), .dout(new_new_n5341__));
  or1   g2243(.dina(new_new_n5340__), .dinb(new_new_n5333__), .dout(new_new_n5342__));
  and1  g2244(.dina(new_new_n5341__), .dinb(new_new_n8724__), .dout(new_new_n5343__));
  and1  g2245(.dina(new_new_n5342__), .dinb(new_new_n8719__), .dout(new_new_n5344__));
  or1   g2246(.dina(new_new_n5344__), .dinb(new_new_n5343__), .dout(new_new_n5345__));
  and1  g2247(.dina(new_new_n9170__), .dinb(new_new_n8926__), .dout(new_new_n5346__));
  and1  g2248(.dina(new_new_n5346__), .dinb(new_new_n8888__), .dout(new_new_n5347__));
  and1  g2249(.dina(new_new_n8848__), .dinb(new_new_n3106__), .dout(new_new_n5348__));
  and1  g2250(.dina(new_new_n5348__), .dinb(new_new_n8949__), .dout(new_new_n5349__));
  or1   g2251(.dina(new_new_n5347__), .dinb(new_new_n5316__), .dout(new_new_n5350__));
  or1   g2252(.dina(new_new_n5350__), .dinb(new_new_n5349__), .dout(new_new_n5351__));
  and1  g2253(.dina(new_new_n8597__), .dinb(new_new_n8849__), .dout(new_new_n5352__));
  and1  g2254(.dina(new_new_n5352__), .dinb(new_new_n8889__), .dout(new_new_n5353__));
  and1  g2255(.dina(new_new_n9161__), .dinb(new_new_n8816__), .dout(new_new_n5354__));
  or1   g2256(.dina(new_new_n9160__), .dinb(new_new_n8814__), .dout(new_new_n5355__));
  and1  g2257(.dina(new_new_n5354__), .dinb(new_new_n9163__), .dout(new_new_n5356__));
  or1   g2258(.dina(new_new_n5355__), .dinb(new_new_n9162__), .dout(new_new_n5357__));
  and1  g2259(.dina(new_new_n5356__), .dinb(new_new_n9169__), .dout(new_new_n5358__));
  or1   g2260(.dina(new_new_n5357__), .dinb(new_new_n9168__), .dout(new_new_n5359__));
  and1  g2261(.dina(new_new_n5358__), .dinb(new_new_n8702__), .dout(new_new_n5360__));
  and1  g2262(.dina(new_new_n5359__), .dinb(new_new_n8692__), .dout(new_new_n5361__));
  or1   g2263(.dina(new_new_n5361__), .dinb(new_new_n5360__), .dout(new_new_n5362__));
  and1  g2264(.dina(new_new_n9171__), .dinb(new_new_n8926__), .dout(new_new_n5363__));
  and1  g2265(.dina(new_new_n5363__), .dinb(new_new_n8889__), .dout(new_new_n5364__));
  and1  g2266(.dina(new_new_n8849__), .dinb(new_new_n3138__), .dout(new_new_n5365__));
  and1  g2267(.dina(new_new_n5365__), .dinb(new_new_n8949__), .dout(new_new_n5366__));
  or1   g2268(.dina(new_new_n5364__), .dinb(new_new_n5353__), .dout(new_new_n5367__));
  or1   g2269(.dina(new_new_n5367__), .dinb(new_new_n5366__), .dout(new_new_n5368__));
  and1  g2270(.dina(new_new_n8596__), .dinb(new_new_n8853__), .dout(new_new_n5369__));
  and1  g2271(.dina(new_new_n5369__), .dinb(new_new_n8893__), .dout(new_new_n5370__));
  and1  g2272(.dina(new_new_n8728__), .dinb(new_new_n8826__), .dout(new_new_n5371__));
  or1   g2273(.dina(new_new_n8733__), .dinb(new_new_n8829__), .dout(new_new_n5372__));
  and1  g2274(.dina(new_new_n9165__), .dinb(new_new_n8729__), .dout(new_new_n5373__));
  or1   g2275(.dina(new_new_n9167__), .dinb(new_new_n8734__), .dout(new_new_n5374__));
  and1  g2276(.dina(new_new_n5372__), .dinb(new_new_n8820__), .dout(new_new_n5375__));
  or1   g2277(.dina(new_new_n5371__), .dinb(new_new_n8818__), .dout(new_new_n5376__));
  and1  g2278(.dina(new_new_n5375__), .dinb(new_new_n5374__), .dout(new_new_n5377__));
  or1   g2279(.dina(new_new_n5376__), .dinb(new_new_n5373__), .dout(new_new_n5378__));
  and1  g2280(.dina(new_new_n5377__), .dinb(new_new_n8714__), .dout(new_new_n5379__));
  and1  g2281(.dina(new_new_n5378__), .dinb(new_new_n8709__), .dout(new_new_n5380__));
  or1   g2282(.dina(new_new_n5380__), .dinb(new_new_n5379__), .dout(new_new_n5381__));
  and1  g2283(.dina(new_new_n9172__), .dinb(new_new_n8929__), .dout(new_new_n5382__));
  and1  g2284(.dina(new_new_n5382__), .dinb(new_new_n8893__), .dout(new_new_n5383__));
  and1  g2285(.dina(new_new_n8853__), .dinb(new_new_n3130__), .dout(new_new_n5384__));
  and1  g2286(.dina(new_new_n5384__), .dinb(new_new_n8952__), .dout(new_new_n5385__));
  or1   g2287(.dina(new_new_n5383__), .dinb(new_new_n5370__), .dout(new_new_n5386__));
  or1   g2288(.dina(new_new_n5386__), .dinb(new_new_n5385__), .dout(new_new_n5387__));
  and1  g2289(.dina(new_new_n8594__), .dinb(new_new_n8852__), .dout(new_new_n5388__));
  and1  g2290(.dina(new_new_n5388__), .dinb(new_new_n8892__), .dout(new_new_n5389__));
  and1  g2291(.dina(new_new_n9166__), .dinb(new_new_n8829__), .dout(new_new_n5390__));
  or1   g2292(.dina(new_new_n9164__), .dinb(new_new_n8826__), .dout(new_new_n5391__));
  and1  g2293(.dina(new_new_n5390__), .dinb(new_new_n8734__), .dout(new_new_n5392__));
  and1  g2294(.dina(new_new_n5391__), .dinb(new_new_n8729__), .dout(new_new_n5393__));
  or1   g2295(.dina(new_new_n5393__), .dinb(new_new_n5392__), .dout(new_new_n5394__));
  and1  g2296(.dina(new_new_n9173__), .dinb(new_new_n8929__), .dout(new_new_n5395__));
  and1  g2297(.dina(new_new_n5395__), .dinb(new_new_n8894__), .dout(new_new_n5396__));
  and1  g2298(.dina(new_new_n8854__), .dinb(new_new_n3122__), .dout(new_new_n5397__));
  and1  g2299(.dina(new_new_n5397__), .dinb(new_new_n8952__), .dout(new_new_n5398__));
  or1   g2300(.dina(new_new_n5396__), .dinb(new_new_n5389__), .dout(new_new_n5399__));
  or1   g2301(.dina(new_new_n5399__), .dinb(new_new_n5398__), .dout(new_new_n5400__));
  and1  g2302(.dina(new_new_n4394__), .dinb(new_new_n4203__), .dout(new_new_n5401__));
  or1   g2303(.dina(new_new_n4395__), .dinb(new_new_n4202__), .dout(new_new_n5402__));
  and1  g2304(.dina(new_new_n4396__), .dinb(new_new_n4201__), .dout(new_new_n5403__));
  or1   g2305(.dina(new_new_n4397__), .dinb(new_new_n4200__), .dout(new_new_n5404__));
  and1  g2306(.dina(new_new_n5404__), .dinb(new_new_n5402__), .dout(new_new_n5405__));
  or1   g2307(.dina(new_new_n5403__), .dinb(new_new_n5401__), .dout(new_new_n5406__));
  and1  g2308(.dina(new_new_n4406__), .dinb(new_new_n4207__), .dout(new_new_n5407__));
  or1   g2309(.dina(new_new_n4407__), .dinb(new_new_n4206__), .dout(new_new_n5408__));
  and1  g2310(.dina(new_new_n4400__), .dinb(new_new_n4213__), .dout(new_new_n5409__));
  or1   g2311(.dina(new_new_n4401__), .dinb(new_new_n4212__), .dout(new_new_n5410__));
  and1  g2312(.dina(new_new_n5410__), .dinb(new_new_n5408__), .dout(new_new_n5411__));
  or1   g2313(.dina(new_new_n5409__), .dinb(new_new_n5407__), .dout(new_new_n5412__));
  and1  g2314(.dina(new_new_n9174__), .dinb(new_new_n9175__), .dout(new_new_n5413__));
  or1   g2315(.dina(new_new_n9176__), .dinb(new_new_n9177__), .dout(new_new_n5414__));
  and1  g2316(.dina(new_new_n9176__), .dinb(new_new_n9177__), .dout(new_new_n5415__));
  or1   g2317(.dina(new_new_n9174__), .dinb(new_new_n9175__), .dout(new_new_n5416__));
  and1  g2318(.dina(new_new_n5416__), .dinb(new_new_n5414__), .dout(new_new_n5417__));
  or1   g2319(.dina(new_new_n5415__), .dinb(new_new_n5413__), .dout(new_new_n5418__));
  and1  g2320(.dina(new_new_n4341__), .dinb(new_new_n4339__), .dout(new_new_n5419__));
  or1   g2321(.dina(new_new_n4340__), .dinb(new_new_n4338__), .dout(new_new_n5420__));
  and1  g2322(.dina(new_new_n4357__), .dinb(new_new_n4342__), .dout(new_new_n5421__));
  or1   g2323(.dina(new_new_n4356__), .dinb(new_new_n4343__), .dout(new_new_n5422__));
  and1  g2324(.dina(new_new_n9179__), .dinb(new_new_n9182__), .dout(new_new_n5423__));
  or1   g2325(.dina(new_new_n9185__), .dinb(new_new_n9188__), .dout(new_new_n5424__));
  and1  g2326(.dina(new_new_n5423__), .dinb(new_new_n9191__), .dout(new_new_n5425__));
  or1   g2327(.dina(new_new_n5424__), .dinb(new_new_n9194__), .dout(new_new_n5426__));
  and1  g2328(.dina(new_new_n9179__), .dinb(new_new_n9188__), .dout(new_new_n5427__));
  or1   g2329(.dina(new_new_n9185__), .dinb(new_new_n9182__), .dout(new_new_n5428__));
  and1  g2330(.dina(new_new_n5427__), .dinb(new_new_n9194__), .dout(new_new_n5429__));
  or1   g2331(.dina(new_new_n5428__), .dinb(new_new_n9191__), .dout(new_new_n5430__));
  and1  g2332(.dina(new_new_n5430__), .dinb(new_new_n5426__), .dout(new_new_n5431__));
  or1   g2333(.dina(new_new_n5429__), .dinb(new_new_n5425__), .dout(new_new_n5432__));
  and1  g2334(.dina(new_new_n9186__), .dinb(new_new_n9189__), .dout(new_new_n5433__));
  or1   g2335(.dina(new_new_n9180__), .dinb(new_new_n9183__), .dout(new_new_n5434__));
  and1  g2336(.dina(new_new_n5433__), .dinb(new_new_n9192__), .dout(new_new_n5435__));
  or1   g2337(.dina(new_new_n5434__), .dinb(new_new_n9195__), .dout(new_new_n5436__));
  and1  g2338(.dina(new_new_n9186__), .dinb(new_new_n9183__), .dout(new_new_n5437__));
  or1   g2339(.dina(new_new_n9180__), .dinb(new_new_n9189__), .dout(new_new_n5438__));
  and1  g2340(.dina(new_new_n5437__), .dinb(new_new_n9195__), .dout(new_new_n5439__));
  or1   g2341(.dina(new_new_n5438__), .dinb(new_new_n9192__), .dout(new_new_n5440__));
  and1  g2342(.dina(new_new_n5440__), .dinb(new_new_n5436__), .dout(new_new_n5441__));
  or1   g2343(.dina(new_new_n5439__), .dinb(new_new_n5435__), .dout(new_new_n5442__));
  and1  g2344(.dina(new_new_n5441__), .dinb(new_new_n5431__), .dout(new_new_n5443__));
  or1   g2345(.dina(new_new_n5442__), .dinb(new_new_n5432__), .dout(new_new_n5444__));
  and1  g2346(.dina(new_new_n5443__), .dinb(new_new_n5418__), .dout(new_new_n5445__));
  and1  g2347(.dina(new_new_n5444__), .dinb(new_new_n5417__), .dout(new_new_n5446__));
  or1   g2348(.dina(new_new_n5446__), .dinb(new_new_n5445__), .dout(new_new_n5447__));
  and1  g2349(.dina(new_new_n4388__), .dinb(new_new_n4197__), .dout(new_new_n5448__));
  or1   g2350(.dina(new_new_n4389__), .dinb(new_new_n4196__), .dout(new_new_n5449__));
  and1  g2351(.dina(new_new_n4390__), .dinb(new_new_n4195__), .dout(new_new_n5450__));
  or1   g2352(.dina(new_new_n4391__), .dinb(new_new_n4194__), .dout(new_new_n5451__));
  and1  g2353(.dina(new_new_n5451__), .dinb(new_new_n5449__), .dout(new_new_n5452__));
  or1   g2354(.dina(new_new_n5450__), .dinb(new_new_n5448__), .dout(new_new_n5453__));
  and1  g2355(.dina(new_new_n4392__), .dinb(new_new_n4193__), .dout(new_new_n5454__));
  or1   g2356(.dina(new_new_n4393__), .dinb(new_new_n4192__), .dout(new_new_n5455__));
  and1  g2357(.dina(new_new_n4386__), .dinb(new_new_n4199__), .dout(new_new_n5456__));
  or1   g2358(.dina(new_new_n4387__), .dinb(new_new_n4198__), .dout(new_new_n5457__));
  and1  g2359(.dina(new_new_n5457__), .dinb(new_new_n5455__), .dout(new_new_n5458__));
  or1   g2360(.dina(new_new_n5456__), .dinb(new_new_n5454__), .dout(new_new_n5459__));
  and1  g2361(.dina(new_new_n9196__), .dinb(new_new_n9197__), .dout(new_new_n5460__));
  or1   g2362(.dina(new_new_n9198__), .dinb(new_new_n9199__), .dout(new_new_n5461__));
  and1  g2363(.dina(new_new_n9198__), .dinb(new_new_n9199__), .dout(new_new_n5462__));
  or1   g2364(.dina(new_new_n9196__), .dinb(new_new_n9197__), .dout(new_new_n5463__));
  and1  g2365(.dina(new_new_n5463__), .dinb(new_new_n5461__), .dout(new_new_n5464__));
  or1   g2366(.dina(new_new_n5462__), .dinb(new_new_n5460__), .dout(new_new_n5465__));
  and1  g2367(.dina(new_new_n4355__), .dinb(new_new_n4347__), .dout(new_new_n5466__));
  or1   g2368(.dina(new_new_n4354__), .dinb(new_new_n4346__), .dout(new_new_n5467__));
  and1  g2369(.dina(new_new_n4349__), .dinb(new_new_n4345__), .dout(new_new_n5468__));
  or1   g2370(.dina(new_new_n4348__), .dinb(new_new_n4344__), .dout(new_new_n5469__));
  and1  g2371(.dina(new_new_n9201__), .dinb(new_new_n9204__), .dout(new_new_n5470__));
  or1   g2372(.dina(new_new_n9207__), .dinb(new_new_n9210__), .dout(new_new_n5471__));
  and1  g2373(.dina(new_new_n5470__), .dinb(new_new_n9213__), .dout(new_new_n5472__));
  or1   g2374(.dina(new_new_n5471__), .dinb(new_new_n9216__), .dout(new_new_n5473__));
  and1  g2375(.dina(new_new_n9201__), .dinb(new_new_n9210__), .dout(new_new_n5474__));
  or1   g2376(.dina(new_new_n9207__), .dinb(new_new_n9204__), .dout(new_new_n5475__));
  and1  g2377(.dina(new_new_n5474__), .dinb(new_new_n9216__), .dout(new_new_n5476__));
  or1   g2378(.dina(new_new_n5475__), .dinb(new_new_n9213__), .dout(new_new_n5477__));
  and1  g2379(.dina(new_new_n5477__), .dinb(new_new_n5473__), .dout(new_new_n5478__));
  or1   g2380(.dina(new_new_n5476__), .dinb(new_new_n5472__), .dout(new_new_n5479__));
  and1  g2381(.dina(new_new_n9208__), .dinb(new_new_n9211__), .dout(new_new_n5480__));
  or1   g2382(.dina(new_new_n9202__), .dinb(new_new_n9205__), .dout(new_new_n5481__));
  and1  g2383(.dina(new_new_n5480__), .dinb(new_new_n9214__), .dout(new_new_n5482__));
  or1   g2384(.dina(new_new_n5481__), .dinb(new_new_n9217__), .dout(new_new_n5483__));
  and1  g2385(.dina(new_new_n9208__), .dinb(new_new_n9205__), .dout(new_new_n5484__));
  or1   g2386(.dina(new_new_n9202__), .dinb(new_new_n9211__), .dout(new_new_n5485__));
  and1  g2387(.dina(new_new_n5484__), .dinb(new_new_n9217__), .dout(new_new_n5486__));
  or1   g2388(.dina(new_new_n5485__), .dinb(new_new_n9214__), .dout(new_new_n5487__));
  and1  g2389(.dina(new_new_n5487__), .dinb(new_new_n5483__), .dout(new_new_n5488__));
  or1   g2390(.dina(new_new_n5486__), .dinb(new_new_n5482__), .dout(new_new_n5489__));
  and1  g2391(.dina(new_new_n5488__), .dinb(new_new_n5478__), .dout(new_new_n5490__));
  or1   g2392(.dina(new_new_n5489__), .dinb(new_new_n5479__), .dout(new_new_n5491__));
  and1  g2393(.dina(new_new_n5490__), .dinb(new_new_n5465__), .dout(new_new_n5492__));
  and1  g2394(.dina(new_new_n5491__), .dinb(new_new_n5464__), .dout(new_new_n5493__));
  or1   g2395(.dina(new_new_n5493__), .dinb(new_new_n5492__), .dout(new_new_n5494__));
  and1  g2396(.dina(new_new_n4952__), .dinb(new_new_n8969__), .dout(new_new_n5495__));
  or1   g2397(.dina(new_new_n8735__), .dinb(new_new_n8971__), .dout(new_new_n5496__));
  and1  g2398(.dina(new_new_n5496__), .dinb(new_new_n8830__), .dout(new_new_n5497__));
  or1   g2399(.dina(new_new_n5495__), .dinb(new_new_n5140__), .dout(new_new_n5498__));
  and1  g2400(.dina(new_new_n9219__), .dinb(new_new_n4222__), .dout(new_new_n5499__));
  and1  g2401(.dina(new_new_n9222__), .dinb(new_new_n8675__), .dout(new_new_n5500__));
  or1   g2402(.dina(new_new_n5500__), .dinb(new_new_n5499__), .dout(new_new_n5501__));
  and1  g2403(.dina(new_new_n8679__), .dinb(new_new_n4104__), .dout(new_new_n5502__));
  and1  g2404(.dina(new_new_n4120__), .dinb(new_new_n8811__), .dout(new_new_n5503__));
  or1   g2405(.dina(new_new_n5503__), .dinb(new_new_n5502__), .dout(new_new_n5504__));
  and1  g2406(.dina(new_new_n5504__), .dinb(new_new_n9219__), .dout(new_new_n5505__));
  or1   g2407(.dina(new_new_n4364__), .dinb(new_new_n4271__), .dout(new_new_n5506__));
  or1   g2408(.dina(new_new_n4365__), .dinb(new_new_n4270__), .dout(new_new_n5507__));
  and1  g2409(.dina(new_new_n5507__), .dinb(new_new_n5506__), .dout(new_new_n5508__));
  and1  g2410(.dina(new_new_n5508__), .dinb(new_new_n9222__), .dout(new_new_n5509__));
  or1   g2411(.dina(new_new_n5509__), .dinb(new_new_n5505__), .dout(new_new_n5510__));
  or1   g2412(.dina(new_new_n4360__), .dinb(new_new_n4329__), .dout(new_new_n5511__));
  or1   g2413(.dina(new_new_n4361__), .dinb(new_new_n4328__), .dout(new_new_n5512__));
  and1  g2414(.dina(new_new_n5512__), .dinb(new_new_n5511__), .dout(new_new_n5513__));
  and1  g2415(.dina(new_new_n5513__), .dinb(new_new_n9220__), .dout(new_new_n5514__));
  and1  g2416(.dina(new_new_n4325__), .dinb(new_new_n8810__), .dout(new_new_n5515__));
  or1   g2417(.dina(new_new_n4324__), .dinb(new_new_n4106__), .dout(new_new_n5516__));
  and1  g2418(.dina(new_new_n5515__), .dinb(new_new_n4363__), .dout(new_new_n5517__));
  or1   g2419(.dina(new_new_n5516__), .dinb(new_new_n4362__), .dout(new_new_n5518__));
  and1  g2420(.dina(new_new_n5517__), .dinb(new_new_n8678__), .dout(new_new_n5519__));
  and1  g2421(.dina(new_new_n5518__), .dinb(new_new_n4118__), .dout(new_new_n5520__));
  or1   g2422(.dina(new_new_n5520__), .dinb(new_new_n5519__), .dout(new_new_n5521__));
  and1  g2423(.dina(new_new_n5521__), .dinb(new_new_n9223__), .dout(new_new_n5522__));
  or1   g2424(.dina(new_new_n5522__), .dinb(new_new_n5514__), .dout(new_new_n5523__));
  or1   g2425(.dina(new_new_n4444__), .dinb(new_new_n4385__), .dout(new_new_n5524__));
  or1   g2426(.dina(new_new_n4445__), .dinb(new_new_n4384__), .dout(new_new_n5525__));
  and1  g2427(.dina(new_new_n5525__), .dinb(new_new_n5524__), .dout(new_new_n5526__));
  and1  g2428(.dina(new_new_n5526__), .dinb(new_new_n9220__), .dout(new_new_n5527__));
  and1  g2429(.dina(new_new_n4327__), .dinb(new_new_n8809__), .dout(new_new_n5528__));
  or1   g2430(.dina(new_new_n4326__), .dinb(new_new_n4190__), .dout(new_new_n5529__));
  and1  g2431(.dina(new_new_n5528__), .dinb(new_new_n4323__), .dout(new_new_n5530__));
  or1   g2432(.dina(new_new_n5529__), .dinb(new_new_n4322__), .dout(new_new_n5531__));
  and1  g2433(.dina(new_new_n5530__), .dinb(new_new_n4359__), .dout(new_new_n5532__));
  or1   g2434(.dina(new_new_n5531__), .dinb(new_new_n4358__), .dout(new_new_n5533__));
  and1  g2435(.dina(new_new_n5532__), .dinb(new_new_n8684__), .dout(new_new_n5534__));
  and1  g2436(.dina(new_new_n5533__), .dinb(new_new_n4224__), .dout(new_new_n5535__));
  or1   g2437(.dina(new_new_n5535__), .dinb(new_new_n5534__), .dout(new_new_n5536__));
  and1  g2438(.dina(new_new_n5536__), .dinb(new_new_n9223__), .dout(new_new_n5537__));
  or1   g2439(.dina(new_new_n5537__), .dinb(new_new_n5527__), .dout(new_new_n5538__));
  or1   g2440(.dina(new_new_n9173__), .dinb(new_new_n8973__), .dout(new_new_n5539__));
  or1   g2441(.dina(new_new_n5539__), .dinb(new_new_n9172__), .dout(new_new_n5540__));
  or1   g2442(.dina(new_new_n5540__), .dinb(new_new_n9171__), .dout(new_new_n5541__));
  or1   g2443(.dina(new_new_n5541__), .dinb(new_new_n9170__), .dout(new_new_n5542__));
  or1   g2444(.dina(new_new_n5542__), .dinb(new_new_n9224__), .dout(new_new_n5543__));
  or1   g2445(.dina(new_new_n5543__), .dinb(new_new_n9225__), .dout(new_new_n5544__));
  or1   g2446(.dina(new_new_n5544__), .dinb(new_new_n9226__), .dout(new_new_n5545__));
  or1   g2447(.dina(new_new_n5545__), .dinb(new_new_n9227__), .dout(new_new_n5546__));
  and1  g2448(.dina(new_new_n8979__), .dinb(new_new_n4226__), .dout(new_new_n5547__));
  and1  g2449(.dina(new_new_n8983__), .dinb(new_new_n8605__), .dout(new_new_n5548__));
  or1   g2450(.dina(new_new_n5548__), .dinb(new_new_n5547__), .dout(new_new_n5549__));
  and1  g2451(.dina(new_new_n8609__), .dinb(new_new_n4110__), .dout(new_new_n5550__));
  and1  g2452(.dina(new_new_n4122__), .dinb(new_new_n8786__), .dout(new_new_n5551__));
  or1   g2453(.dina(new_new_n5551__), .dinb(new_new_n5550__), .dout(new_new_n5552__));
  and1  g2454(.dina(new_new_n5552__), .dinb(new_new_n8981__), .dout(new_new_n5553__));
  or1   g2455(.dina(new_new_n4368__), .dinb(new_new_n4273__), .dout(new_new_n5554__));
  or1   g2456(.dina(new_new_n4369__), .dinb(new_new_n4272__), .dout(new_new_n5555__));
  and1  g2457(.dina(new_new_n5555__), .dinb(new_new_n5554__), .dout(new_new_n5556__));
  and1  g2458(.dina(new_new_n5556__), .dinb(new_new_n8985__), .dout(new_new_n5557__));
  or1   g2459(.dina(new_new_n5557__), .dinb(new_new_n5553__), .dout(new_new_n5558__));
  or1   g2460(.dina(new_new_n4351__), .dinb(new_new_n4333__), .dout(new_new_n5559__));
  or1   g2461(.dina(new_new_n4350__), .dinb(new_new_n4332__), .dout(new_new_n5560__));
  and1  g2462(.dina(new_new_n5560__), .dinb(new_new_n5559__), .dout(new_new_n5561__));
  and1  g2463(.dina(new_new_n5561__), .dinb(new_new_n8981__), .dout(new_new_n5562__));
  and1  g2464(.dina(new_new_n4337__), .dinb(new_new_n8785__), .dout(new_new_n5563__));
  or1   g2465(.dina(new_new_n4336__), .dinb(new_new_n4108__), .dout(new_new_n5564__));
  and1  g2466(.dina(new_new_n5563__), .dinb(new_new_n4367__), .dout(new_new_n5565__));
  or1   g2467(.dina(new_new_n5564__), .dinb(new_new_n4366__), .dout(new_new_n5566__));
  and1  g2468(.dina(new_new_n5565__), .dinb(new_new_n8608__), .dout(new_new_n5567__));
  and1  g2469(.dina(new_new_n5566__), .dinb(new_new_n4113__), .dout(new_new_n5568__));
  or1   g2470(.dina(new_new_n5568__), .dinb(new_new_n5567__), .dout(new_new_n5569__));
  and1  g2471(.dina(new_new_n5569__), .dinb(new_new_n8985__), .dout(new_new_n5570__));
  or1   g2472(.dina(new_new_n5570__), .dinb(new_new_n5562__), .dout(new_new_n5571__));
  or1   g2473(.dina(new_new_n8968__), .dinb(new_new_n8917__), .dout(new_new_n5572__));
  or1   g2474(.dina(new_new_n5572__), .dinb(new_new_n9083__), .dout(new_new_n5573__));
  or1   g2475(.dina(new_new_n5573__), .dinb(new_new_n9082__), .dout(new_new_n5574__));
  or1   g2476(.dina(new_new_n5574__), .dinb(new_new_n9081__), .dout(new_new_n5575__));
  or1   g2477(.dina(new_new_n5575__), .dinb(new_new_n9228__), .dout(new_new_n5576__));
  or1   g2478(.dina(new_new_n5576__), .dinb(new_new_n9229__), .dout(new_new_n5577__));
  or1   g2479(.dina(new_new_n5577__), .dinb(new_new_n9230__), .dout(new_new_n5578__));
  or1   g2480(.dina(new_new_n5578__), .dinb(new_new_n9232__), .dout(new_new_n5579__));
  and1  g2481(.dina(new_new_n8990__), .dinb(new_new_n9238__), .dout(new_new_n5580__));
  and1  g2482(.dina(new_new_n5580__), .dinb(new_new_n9257__), .dout(new_new_n5581__));
  and1  g2483(.dina(new_new_n9032__), .dinb(new_new_n9276__), .dout(new_new_n5582__));
  and1  g2484(.dina(new_new_n5582__), .dinb(new_new_n9257__), .dout(new_new_n5583__));
  and1  g2485(.dina(new_new_n9238__), .dinb(new_new_n9291__), .dout(new_new_n5584__));
  and1  g2486(.dina(new_new_n5584__), .dinb(new_new_n9296__), .dout(new_new_n5585__));
  and1  g2487(.dina(new_new_n9276__), .dinb(new_new_n9311__), .dout(new_new_n5586__));
  and1  g2488(.dina(new_new_n5586__), .dinb(new_new_n9296__), .dout(new_new_n5587__));
  or1   g2489(.dina(new_new_n5583__), .dinb(new_new_n5581__), .dout(new_new_n5588__));
  or1   g2490(.dina(new_new_n5588__), .dinb(new_new_n5585__), .dout(new_new_n5589__));
  or1   g2491(.dina(new_new_n5589__), .dinb(new_new_n5587__), .dout(new_new_n5590__));
  and1  g2492(.dina(new_new_n5590__), .dinb(new_new_n9316__), .dout(new_new_n5591__));
  and1  g2493(.dina(new_new_n8992__), .dinb(new_new_n9336__), .dout(new_new_n5592__));
  and1  g2494(.dina(new_new_n5592__), .dinb(new_new_n9355__), .dout(new_new_n5593__));
  and1  g2495(.dina(new_new_n9034__), .dinb(new_new_n9374__), .dout(new_new_n5594__));
  and1  g2496(.dina(new_new_n5594__), .dinb(new_new_n9355__), .dout(new_new_n5595__));
  and1  g2497(.dina(new_new_n9336__), .dinb(new_new_n9291__), .dout(new_new_n5596__));
  and1  g2498(.dina(new_new_n5596__), .dinb(new_new_n9393__), .dout(new_new_n5597__));
  and1  g2499(.dina(new_new_n9374__), .dinb(new_new_n9311__), .dout(new_new_n5598__));
  and1  g2500(.dina(new_new_n5598__), .dinb(new_new_n9393__), .dout(new_new_n5599__));
  or1   g2501(.dina(new_new_n5595__), .dinb(new_new_n5593__), .dout(new_new_n5600__));
  or1   g2502(.dina(new_new_n5600__), .dinb(new_new_n5597__), .dout(new_new_n5601__));
  or1   g2503(.dina(new_new_n5601__), .dinb(new_new_n5599__), .dout(new_new_n5602__));
  and1  g2504(.dina(new_new_n5602__), .dinb(new_new_n9316__), .dout(new_new_n5603__));
  and1  g2505(.dina(new_new_n9410__), .dinb(new_new_n8998__), .dout(new_new_n5604__));
  and1  g2506(.dina(new_new_n5604__), .dinb(new_new_n9017__), .dout(new_new_n5605__));
  and1  g2507(.dina(new_new_n9414__), .dinb(new_new_n9040__), .dout(new_new_n5606__));
  and1  g2508(.dina(new_new_n5606__), .dinb(new_new_n9017__), .dout(new_new_n5607__));
  and1  g2509(.dina(new_new_n8998__), .dinb(new_new_n9416__), .dout(new_new_n5608__));
  and1  g2510(.dina(new_new_n5608__), .dinb(new_new_n9060__), .dout(new_new_n5609__));
  and1  g2511(.dina(new_new_n9040__), .dinb(new_new_n9417__), .dout(new_new_n5610__));
  and1  g2512(.dina(new_new_n5610__), .dinb(new_new_n9060__), .dout(new_new_n5611__));
  or1   g2513(.dina(new_new_n5607__), .dinb(new_new_n5605__), .dout(new_new_n5612__));
  or1   g2514(.dina(new_new_n5612__), .dinb(new_new_n5609__), .dout(new_new_n5613__));
  or1   g2515(.dina(new_new_n5613__), .dinb(new_new_n5611__), .dout(new_new_n5614__));
  and1  g2516(.dina(new_new_n9420__), .dinb(new_new_n9000__), .dout(new_new_n5615__));
  and1  g2517(.dina(new_new_n5615__), .dinb(new_new_n9019__), .dout(new_new_n5616__));
  and1  g2518(.dina(new_new_n9424__), .dinb(new_new_n9042__), .dout(new_new_n5617__));
  and1  g2519(.dina(new_new_n5617__), .dinb(new_new_n9019__), .dout(new_new_n5618__));
  and1  g2520(.dina(new_new_n9000__), .dinb(new_new_n9426__), .dout(new_new_n5619__));
  and1  g2521(.dina(new_new_n5619__), .dinb(new_new_n9062__), .dout(new_new_n5620__));
  and1  g2522(.dina(new_new_n9042__), .dinb(new_new_n9427__), .dout(new_new_n5621__));
  and1  g2523(.dina(new_new_n5621__), .dinb(new_new_n9062__), .dout(new_new_n5622__));
  or1   g2524(.dina(new_new_n5618__), .dinb(new_new_n5616__), .dout(new_new_n5623__));
  or1   g2525(.dina(new_new_n5623__), .dinb(new_new_n5620__), .dout(new_new_n5624__));
  or1   g2526(.dina(new_new_n5624__), .dinb(new_new_n5622__), .dout(new_new_n5625__));
  and1  g2527(.dina(new_new_n9430__), .dinb(new_new_n9001__), .dout(new_new_n5626__));
  and1  g2528(.dina(new_new_n5626__), .dinb(new_new_n9020__), .dout(new_new_n5627__));
  and1  g2529(.dina(new_new_n9434__), .dinb(new_new_n9043__), .dout(new_new_n5628__));
  and1  g2530(.dina(new_new_n5628__), .dinb(new_new_n9020__), .dout(new_new_n5629__));
  and1  g2531(.dina(new_new_n9001__), .dinb(new_new_n9436__), .dout(new_new_n5630__));
  and1  g2532(.dina(new_new_n5630__), .dinb(new_new_n9063__), .dout(new_new_n5631__));
  and1  g2533(.dina(new_new_n9043__), .dinb(new_new_n9437__), .dout(new_new_n5632__));
  and1  g2534(.dina(new_new_n5632__), .dinb(new_new_n9063__), .dout(new_new_n5633__));
  or1   g2535(.dina(new_new_n5629__), .dinb(new_new_n5627__), .dout(new_new_n5634__));
  or1   g2536(.dina(new_new_n5634__), .dinb(new_new_n5631__), .dout(new_new_n5635__));
  or1   g2537(.dina(new_new_n5635__), .dinb(new_new_n5633__), .dout(new_new_n5636__));
  and1  g2538(.dina(new_new_n9440__), .dinb(new_new_n9003__), .dout(new_new_n5637__));
  and1  g2539(.dina(new_new_n5637__), .dinb(new_new_n9022__), .dout(new_new_n5638__));
  and1  g2540(.dina(new_new_n9444__), .dinb(new_new_n9045__), .dout(new_new_n5639__));
  and1  g2541(.dina(new_new_n5639__), .dinb(new_new_n9022__), .dout(new_new_n5640__));
  and1  g2542(.dina(new_new_n9003__), .dinb(new_new_n9446__), .dout(new_new_n5641__));
  and1  g2543(.dina(new_new_n5641__), .dinb(new_new_n9065__), .dout(new_new_n5642__));
  and1  g2544(.dina(new_new_n9045__), .dinb(new_new_n9447__), .dout(new_new_n5643__));
  and1  g2545(.dina(new_new_n5643__), .dinb(new_new_n9065__), .dout(new_new_n5644__));
  or1   g2546(.dina(new_new_n5640__), .dinb(new_new_n5638__), .dout(new_new_n5645__));
  or1   g2547(.dina(new_new_n5645__), .dinb(new_new_n5642__), .dout(new_new_n5646__));
  or1   g2548(.dina(new_new_n5646__), .dinb(new_new_n5644__), .dout(new_new_n5647__));
  and1  g2549(.dina(new_new_n9410__), .dinb(new_new_n9089__), .dout(new_new_n5648__));
  and1  g2550(.dina(new_new_n5648__), .dinb(new_new_n9108__), .dout(new_new_n5649__));
  and1  g2551(.dina(new_new_n9414__), .dinb(new_new_n9127__), .dout(new_new_n5650__));
  and1  g2552(.dina(new_new_n5650__), .dinb(new_new_n9108__), .dout(new_new_n5651__));
  and1  g2553(.dina(new_new_n9089__), .dinb(new_new_n9416__), .dout(new_new_n5652__));
  and1  g2554(.dina(new_new_n5652__), .dinb(new_new_n9146__), .dout(new_new_n5653__));
  and1  g2555(.dina(new_new_n9127__), .dinb(new_new_n9417__), .dout(new_new_n5654__));
  and1  g2556(.dina(new_new_n5654__), .dinb(new_new_n9146__), .dout(new_new_n5655__));
  or1   g2557(.dina(new_new_n5651__), .dinb(new_new_n5649__), .dout(new_new_n5656__));
  or1   g2558(.dina(new_new_n5656__), .dinb(new_new_n5653__), .dout(new_new_n5657__));
  or1   g2559(.dina(new_new_n5657__), .dinb(new_new_n5655__), .dout(new_new_n5658__));
  and1  g2560(.dina(new_new_n9420__), .dinb(new_new_n9091__), .dout(new_new_n5659__));
  and1  g2561(.dina(new_new_n5659__), .dinb(new_new_n9110__), .dout(new_new_n5660__));
  and1  g2562(.dina(new_new_n9424__), .dinb(new_new_n9129__), .dout(new_new_n5661__));
  and1  g2563(.dina(new_new_n5661__), .dinb(new_new_n9110__), .dout(new_new_n5662__));
  and1  g2564(.dina(new_new_n9091__), .dinb(new_new_n9426__), .dout(new_new_n5663__));
  and1  g2565(.dina(new_new_n5663__), .dinb(new_new_n9148__), .dout(new_new_n5664__));
  and1  g2566(.dina(new_new_n9129__), .dinb(new_new_n9427__), .dout(new_new_n5665__));
  and1  g2567(.dina(new_new_n5665__), .dinb(new_new_n9148__), .dout(new_new_n5666__));
  or1   g2568(.dina(new_new_n5662__), .dinb(new_new_n5660__), .dout(new_new_n5667__));
  or1   g2569(.dina(new_new_n5667__), .dinb(new_new_n5664__), .dout(new_new_n5668__));
  or1   g2570(.dina(new_new_n5668__), .dinb(new_new_n5666__), .dout(new_new_n5669__));
  and1  g2571(.dina(new_new_n9430__), .dinb(new_new_n9092__), .dout(new_new_n5670__));
  and1  g2572(.dina(new_new_n5670__), .dinb(new_new_n9111__), .dout(new_new_n5671__));
  and1  g2573(.dina(new_new_n9434__), .dinb(new_new_n9130__), .dout(new_new_n5672__));
  and1  g2574(.dina(new_new_n5672__), .dinb(new_new_n9111__), .dout(new_new_n5673__));
  and1  g2575(.dina(new_new_n9092__), .dinb(new_new_n9436__), .dout(new_new_n5674__));
  and1  g2576(.dina(new_new_n5674__), .dinb(new_new_n9149__), .dout(new_new_n5675__));
  and1  g2577(.dina(new_new_n9130__), .dinb(new_new_n9437__), .dout(new_new_n5676__));
  and1  g2578(.dina(new_new_n5676__), .dinb(new_new_n9149__), .dout(new_new_n5677__));
  or1   g2579(.dina(new_new_n5673__), .dinb(new_new_n5671__), .dout(new_new_n5678__));
  or1   g2580(.dina(new_new_n5678__), .dinb(new_new_n5675__), .dout(new_new_n5679__));
  or1   g2581(.dina(new_new_n5679__), .dinb(new_new_n5677__), .dout(new_new_n5680__));
  and1  g2582(.dina(new_new_n9440__), .dinb(new_new_n9094__), .dout(new_new_n5681__));
  and1  g2583(.dina(new_new_n5681__), .dinb(new_new_n9113__), .dout(new_new_n5682__));
  and1  g2584(.dina(new_new_n9444__), .dinb(new_new_n9132__), .dout(new_new_n5683__));
  and1  g2585(.dina(new_new_n5683__), .dinb(new_new_n9113__), .dout(new_new_n5684__));
  and1  g2586(.dina(new_new_n9094__), .dinb(new_new_n9446__), .dout(new_new_n5685__));
  and1  g2587(.dina(new_new_n5685__), .dinb(new_new_n9151__), .dout(new_new_n5686__));
  and1  g2588(.dina(new_new_n9132__), .dinb(new_new_n9447__), .dout(new_new_n5687__));
  and1  g2589(.dina(new_new_n5687__), .dinb(new_new_n9151__), .dout(new_new_n5688__));
  or1   g2590(.dina(new_new_n5684__), .dinb(new_new_n5682__), .dout(new_new_n5689__));
  or1   g2591(.dina(new_new_n5689__), .dinb(new_new_n5686__), .dout(new_new_n5690__));
  or1   g2592(.dina(new_new_n5690__), .dinb(new_new_n5688__), .dout(new_new_n5691__));
  and1  g2593(.dina(new_new_n9409__), .dinb(new_new_n9239__), .dout(new_new_n5692__));
  and1  g2594(.dina(new_new_n5692__), .dinb(new_new_n9258__), .dout(new_new_n5693__));
  and1  g2595(.dina(new_new_n9413__), .dinb(new_new_n9277__), .dout(new_new_n5694__));
  and1  g2596(.dina(new_new_n5694__), .dinb(new_new_n9258__), .dout(new_new_n5695__));
  and1  g2597(.dina(new_new_n9239__), .dinb(new_new_n9448__), .dout(new_new_n5696__));
  and1  g2598(.dina(new_new_n5696__), .dinb(new_new_n9297__), .dout(new_new_n5697__));
  and1  g2599(.dina(new_new_n9277__), .dinb(new_new_n9449__), .dout(new_new_n5698__));
  and1  g2600(.dina(new_new_n5698__), .dinb(new_new_n9297__), .dout(new_new_n5699__));
  or1   g2601(.dina(new_new_n5695__), .dinb(new_new_n5693__), .dout(new_new_n5700__));
  or1   g2602(.dina(new_new_n5700__), .dinb(new_new_n5697__), .dout(new_new_n5701__));
  or1   g2603(.dina(new_new_n5701__), .dinb(new_new_n5699__), .dout(new_new_n5702__));
  and1  g2604(.dina(new_new_n5702__), .dinb(new_new_n9317__), .dout(new_new_n5703__));
  and1  g2605(.dina(new_new_n9439__), .dinb(new_new_n9241__), .dout(new_new_n5704__));
  and1  g2606(.dina(new_new_n5704__), .dinb(new_new_n9260__), .dout(new_new_n5705__));
  and1  g2607(.dina(new_new_n9443__), .dinb(new_new_n9279__), .dout(new_new_n5706__));
  and1  g2608(.dina(new_new_n5706__), .dinb(new_new_n9260__), .dout(new_new_n5707__));
  and1  g2609(.dina(new_new_n9241__), .dinb(new_new_n9450__), .dout(new_new_n5708__));
  and1  g2610(.dina(new_new_n5708__), .dinb(new_new_n9299__), .dout(new_new_n5709__));
  and1  g2611(.dina(new_new_n9279__), .dinb(new_new_n9451__), .dout(new_new_n5710__));
  and1  g2612(.dina(new_new_n5710__), .dinb(new_new_n9299__), .dout(new_new_n5711__));
  or1   g2613(.dina(new_new_n5707__), .dinb(new_new_n5705__), .dout(new_new_n5712__));
  or1   g2614(.dina(new_new_n5712__), .dinb(new_new_n5709__), .dout(new_new_n5713__));
  or1   g2615(.dina(new_new_n5713__), .dinb(new_new_n5711__), .dout(new_new_n5714__));
  and1  g2616(.dina(new_new_n5714__), .dinb(new_new_n9317__), .dout(new_new_n5715__));
  and1  g2617(.dina(new_new_n9429__), .dinb(new_new_n9242__), .dout(new_new_n5716__));
  and1  g2618(.dina(new_new_n5716__), .dinb(new_new_n9261__), .dout(new_new_n5717__));
  and1  g2619(.dina(new_new_n9433__), .dinb(new_new_n9280__), .dout(new_new_n5718__));
  and1  g2620(.dina(new_new_n5718__), .dinb(new_new_n9261__), .dout(new_new_n5719__));
  and1  g2621(.dina(new_new_n9242__), .dinb(new_new_n9452__), .dout(new_new_n5720__));
  and1  g2622(.dina(new_new_n5720__), .dinb(new_new_n9300__), .dout(new_new_n5721__));
  and1  g2623(.dina(new_new_n9280__), .dinb(new_new_n9453__), .dout(new_new_n5722__));
  and1  g2624(.dina(new_new_n5722__), .dinb(new_new_n9300__), .dout(new_new_n5723__));
  or1   g2625(.dina(new_new_n5719__), .dinb(new_new_n5717__), .dout(new_new_n5724__));
  or1   g2626(.dina(new_new_n5724__), .dinb(new_new_n5721__), .dout(new_new_n5725__));
  or1   g2627(.dina(new_new_n5725__), .dinb(new_new_n5723__), .dout(new_new_n5726__));
  and1  g2628(.dina(new_new_n5726__), .dinb(new_new_n9319__), .dout(new_new_n5727__));
  and1  g2629(.dina(new_new_n9419__), .dinb(new_new_n9244__), .dout(new_new_n5728__));
  and1  g2630(.dina(new_new_n5728__), .dinb(new_new_n9263__), .dout(new_new_n5729__));
  and1  g2631(.dina(new_new_n9423__), .dinb(new_new_n9282__), .dout(new_new_n5730__));
  and1  g2632(.dina(new_new_n5730__), .dinb(new_new_n9263__), .dout(new_new_n5731__));
  and1  g2633(.dina(new_new_n9244__), .dinb(new_new_n9454__), .dout(new_new_n5732__));
  and1  g2634(.dina(new_new_n5732__), .dinb(new_new_n9302__), .dout(new_new_n5733__));
  and1  g2635(.dina(new_new_n9282__), .dinb(new_new_n9455__), .dout(new_new_n5734__));
  and1  g2636(.dina(new_new_n5734__), .dinb(new_new_n9302__), .dout(new_new_n5735__));
  or1   g2637(.dina(new_new_n5731__), .dinb(new_new_n5729__), .dout(new_new_n5736__));
  or1   g2638(.dina(new_new_n5736__), .dinb(new_new_n5733__), .dout(new_new_n5737__));
  or1   g2639(.dina(new_new_n5737__), .dinb(new_new_n5735__), .dout(new_new_n5738__));
  and1  g2640(.dina(new_new_n5738__), .dinb(new_new_n9319__), .dout(new_new_n5739__));
  and1  g2641(.dina(new_new_n9411__), .dinb(new_new_n9337__), .dout(new_new_n5740__));
  and1  g2642(.dina(new_new_n5740__), .dinb(new_new_n9356__), .dout(new_new_n5741__));
  and1  g2643(.dina(new_new_n9415__), .dinb(new_new_n9375__), .dout(new_new_n5742__));
  and1  g2644(.dina(new_new_n5742__), .dinb(new_new_n9356__), .dout(new_new_n5743__));
  and1  g2645(.dina(new_new_n9337__), .dinb(new_new_n9448__), .dout(new_new_n5744__));
  and1  g2646(.dina(new_new_n5744__), .dinb(new_new_n9394__), .dout(new_new_n5745__));
  and1  g2647(.dina(new_new_n9375__), .dinb(new_new_n9449__), .dout(new_new_n5746__));
  and1  g2648(.dina(new_new_n5746__), .dinb(new_new_n9394__), .dout(new_new_n5747__));
  or1   g2649(.dina(new_new_n5743__), .dinb(new_new_n5741__), .dout(new_new_n5748__));
  or1   g2650(.dina(new_new_n5748__), .dinb(new_new_n5745__), .dout(new_new_n5749__));
  or1   g2651(.dina(new_new_n5749__), .dinb(new_new_n5747__), .dout(new_new_n5750__));
  and1  g2652(.dina(new_new_n5750__), .dinb(new_new_n9320__), .dout(new_new_n5751__));
  and1  g2653(.dina(new_new_n9441__), .dinb(new_new_n9339__), .dout(new_new_n5752__));
  and1  g2654(.dina(new_new_n5752__), .dinb(new_new_n9358__), .dout(new_new_n5753__));
  and1  g2655(.dina(new_new_n9445__), .dinb(new_new_n9377__), .dout(new_new_n5754__));
  and1  g2656(.dina(new_new_n5754__), .dinb(new_new_n9358__), .dout(new_new_n5755__));
  and1  g2657(.dina(new_new_n9339__), .dinb(new_new_n9450__), .dout(new_new_n5756__));
  and1  g2658(.dina(new_new_n5756__), .dinb(new_new_n9396__), .dout(new_new_n5757__));
  and1  g2659(.dina(new_new_n9377__), .dinb(new_new_n9451__), .dout(new_new_n5758__));
  and1  g2660(.dina(new_new_n5758__), .dinb(new_new_n9396__), .dout(new_new_n5759__));
  or1   g2661(.dina(new_new_n5755__), .dinb(new_new_n5753__), .dout(new_new_n5760__));
  or1   g2662(.dina(new_new_n5760__), .dinb(new_new_n5757__), .dout(new_new_n5761__));
  or1   g2663(.dina(new_new_n5761__), .dinb(new_new_n5759__), .dout(new_new_n5762__));
  and1  g2664(.dina(new_new_n5762__), .dinb(new_new_n9320__), .dout(new_new_n5763__));
  and1  g2665(.dina(new_new_n9431__), .dinb(new_new_n9340__), .dout(new_new_n5764__));
  and1  g2666(.dina(new_new_n5764__), .dinb(new_new_n9359__), .dout(new_new_n5765__));
  and1  g2667(.dina(new_new_n9435__), .dinb(new_new_n9378__), .dout(new_new_n5766__));
  and1  g2668(.dina(new_new_n5766__), .dinb(new_new_n9359__), .dout(new_new_n5767__));
  and1  g2669(.dina(new_new_n9340__), .dinb(new_new_n9452__), .dout(new_new_n5768__));
  and1  g2670(.dina(new_new_n5768__), .dinb(new_new_n9397__), .dout(new_new_n5769__));
  and1  g2671(.dina(new_new_n9378__), .dinb(new_new_n9453__), .dout(new_new_n5770__));
  and1  g2672(.dina(new_new_n5770__), .dinb(new_new_n9397__), .dout(new_new_n5771__));
  or1   g2673(.dina(new_new_n5767__), .dinb(new_new_n5765__), .dout(new_new_n5772__));
  or1   g2674(.dina(new_new_n5772__), .dinb(new_new_n5769__), .dout(new_new_n5773__));
  or1   g2675(.dina(new_new_n5773__), .dinb(new_new_n5771__), .dout(new_new_n5774__));
  and1  g2676(.dina(new_new_n5774__), .dinb(new_new_n9323__), .dout(new_new_n5775__));
  and1  g2677(.dina(new_new_n9421__), .dinb(new_new_n9342__), .dout(new_new_n5776__));
  and1  g2678(.dina(new_new_n5776__), .dinb(new_new_n9361__), .dout(new_new_n5777__));
  and1  g2679(.dina(new_new_n9425__), .dinb(new_new_n9380__), .dout(new_new_n5778__));
  and1  g2680(.dina(new_new_n5778__), .dinb(new_new_n9361__), .dout(new_new_n5779__));
  and1  g2681(.dina(new_new_n9342__), .dinb(new_new_n9454__), .dout(new_new_n5780__));
  and1  g2682(.dina(new_new_n5780__), .dinb(new_new_n9399__), .dout(new_new_n5781__));
  and1  g2683(.dina(new_new_n9380__), .dinb(new_new_n9455__), .dout(new_new_n5782__));
  and1  g2684(.dina(new_new_n5782__), .dinb(new_new_n9399__), .dout(new_new_n5783__));
  or1   g2685(.dina(new_new_n5779__), .dinb(new_new_n5777__), .dout(new_new_n5784__));
  or1   g2686(.dina(new_new_n5784__), .dinb(new_new_n5781__), .dout(new_new_n5785__));
  or1   g2687(.dina(new_new_n5785__), .dinb(new_new_n5783__), .dout(new_new_n5786__));
  and1  g2688(.dina(new_new_n5786__), .dinb(new_new_n9323__), .dout(new_new_n5787__));
  or1   g2689(.dina(new_new_n3823__), .dinb(new_new_n3179__), .dout(new_new_n5788__));
  and1  g2690(.dina(new_new_n9456__), .dinb(new_new_n9457__), .dout(new_new_n5789__));
  and1  g2691(.dina(new_new_n5789__), .dinb(new_new_n9458__), .dout(new_new_n5790__));
  and1  g2692(.dina(new_new_n9459__), .dinb(new_new_n9460__), .dout(new_new_n5791__));
  or1   g2693(.dina(new_new_n8789__), .dinb(new_new_n9461__), .dout(new_new_n5792__));
  and1  g2694(.dina(new_new_n9462__), .dinb(new_new_n9459__), .dout(new_new_n5793__));
  or1   g2695(.dina(new_new_n9463__), .dinb(new_new_n8789__), .dout(new_new_n5794__));
  and1  g2696(.dina(new_new_n9462__), .dinb(new_new_n9460__), .dout(new_new_n5795__));
  or1   g2697(.dina(new_new_n9463__), .dinb(new_new_n9461__), .dout(new_new_n5796__));
  and1  g2698(.dina(new_new_n5796__), .dinb(new_new_n5794__), .dout(new_new_n5797__));
  or1   g2699(.dina(new_new_n5795__), .dinb(new_new_n5793__), .dout(new_new_n5798__));
  and1  g2700(.dina(new_new_n9464__), .dinb(new_new_n9465__), .dout(new_new_n5799__));
  and1  g2701(.dina(new_new_n5799__), .dinb(new_new_n9458__), .dout(new_new_n5800__));
  and1  g2702(.dina(new_new_n9457__), .dinb(new_new_n9466__), .dout(new_new_n5801__));
  and1  g2703(.dina(new_new_n5801__), .dinb(new_new_n9467__), .dout(new_new_n5802__));
  and1  g2704(.dina(new_new_n9232__), .dinb(new_new_n9465__), .dout(new_new_n5803__));
  and1  g2705(.dina(new_new_n5803__), .dinb(new_new_n9467__), .dout(new_new_n5804__));
  or1   g2706(.dina(new_new_n5800__), .dinb(new_new_n5790__), .dout(new_new_n5805__));
  or1   g2707(.dina(new_new_n5805__), .dinb(new_new_n5802__), .dout(new_new_n5806__));
  or1   g2708(.dina(new_new_n5806__), .dinb(new_new_n5804__), .dout(new_new_n5807__));
  and1  g2709(.dina(new_new_n5807__), .dinb(new_new_n5788__), .dout(new_new_n5808__));
  or1   g2710(.dina(new_new_n5797__), .dinb(new_new_n9468__), .dout(new_new_n5809__));
  and1  g2711(.dina(new_new_n9469__), .dinb(new_new_n9464__), .dout(new_new_n5810__));
  and1  g2712(.dina(new_new_n9469__), .dinb(new_new_n9233__), .dout(new_new_n5811__));
  or1   g2713(.dina(new_new_n5811__), .dinb(new_new_n5810__), .dout(new_new_n5812__));
  and1  g2714(.dina(new_new_n9456__), .dinb(new_new_n8854__), .dout(new_new_n5813__));
  and1  g2715(.dina(new_new_n5813__), .dinb(new_new_n8894__), .dout(new_new_n5814__));
  and1  g2716(.dina(new_new_n9233__), .dinb(new_new_n8930__), .dout(new_new_n5815__));
  and1  g2717(.dina(new_new_n5815__), .dinb(new_new_n8896__), .dout(new_new_n5816__));
  and1  g2718(.dina(new_new_n8856__), .dinb(new_new_n9466__), .dout(new_new_n5817__));
  and1  g2719(.dina(new_new_n5817__), .dinb(new_new_n8953__), .dout(new_new_n5818__));
  or1   g2720(.dina(new_new_n5816__), .dinb(new_new_n5814__), .dout(new_new_n5819__));
  or1   g2721(.dina(new_new_n5819__), .dinb(new_new_n5818__), .dout(new_new_n5820__));
  and1  g2722(.dina(new_new_n8506__), .dinb(new_new_n8856__), .dout(new_new_n5821__));
  and1  g2723(.dina(new_new_n5821__), .dinb(new_new_n8896__), .dout(new_new_n5822__));
  and1  g2724(.dina(new_new_n9230__), .dinb(new_new_n8930__), .dout(new_new_n5823__));
  and1  g2725(.dina(new_new_n5823__), .dinb(new_new_n8897__), .dout(new_new_n5824__));
  and1  g2726(.dina(new_new_n8857__), .dinb(new_new_n3098__), .dout(new_new_n5825__));
  and1  g2727(.dina(new_new_n5825__), .dinb(new_new_n8953__), .dout(new_new_n5826__));
  or1   g2728(.dina(new_new_n5824__), .dinb(new_new_n5822__), .dout(new_new_n5827__));
  or1   g2729(.dina(new_new_n5827__), .dinb(new_new_n5826__), .dout(new_new_n5828__));
  and1  g2730(.dina(new_new_n8504__), .dinb(new_new_n8857__), .dout(new_new_n5829__));
  and1  g2731(.dina(new_new_n5829__), .dinb(new_new_n8897__), .dout(new_new_n5830__));
  and1  g2732(.dina(new_new_n9229__), .dinb(new_new_n8932__), .dout(new_new_n5831__));
  and1  g2733(.dina(new_new_n5831__), .dinb(new_new_n8901__), .dout(new_new_n5832__));
  and1  g2734(.dina(new_new_n8861__), .dinb(new_new_n3058__), .dout(new_new_n5833__));
  and1  g2735(.dina(new_new_n5833__), .dinb(new_new_n8955__), .dout(new_new_n5834__));
  or1   g2736(.dina(new_new_n5832__), .dinb(new_new_n5830__), .dout(new_new_n5835__));
  or1   g2737(.dina(new_new_n5835__), .dinb(new_new_n5834__), .dout(new_new_n5836__));
  and1  g2738(.dina(new_new_n8505__), .dinb(new_new_n8861__), .dout(new_new_n5837__));
  and1  g2739(.dina(new_new_n5837__), .dinb(new_new_n8901__), .dout(new_new_n5838__));
  and1  g2740(.dina(new_new_n9228__), .dinb(new_new_n8932__), .dout(new_new_n5839__));
  and1  g2741(.dina(new_new_n5839__), .dinb(new_new_n8902__), .dout(new_new_n5840__));
  and1  g2742(.dina(new_new_n8862__), .dinb(new_new_n3026__), .dout(new_new_n5841__));
  and1  g2743(.dina(new_new_n5841__), .dinb(new_new_n8955__), .dout(new_new_n5842__));
  or1   g2744(.dina(new_new_n5840__), .dinb(new_new_n5838__), .dout(new_new_n5843__));
  or1   g2745(.dina(new_new_n5843__), .dinb(new_new_n5842__), .dout(new_new_n5844__));
  or1   g2746(.dina(new_new_n9470__), .dinb(new_new_n8448__), .dout(new_new_n5845__));
  or1   g2747(.dina(new_new_n5845__), .dinb(new_new_n8447__), .dout(new_new_n5846__));
  or1   g2748(.dina(new_new_n5846__), .dinb(new_new_n9471__), .dout(new_new_n5847__));
  or1   g2749(.dina(new_new_n9472__), .dinb(new_new_n9473__), .dout(new_new_n5848__));
  or1   g2750(.dina(new_new_n5848__), .dinb(new_new_n9474__), .dout(new_new_n5849__));
  or1   g2751(.dina(new_new_n5849__), .dinb(new_new_n9475__), .dout(new_new_n5850__));
  or1   g2752(.dina(new_new_n5850__), .dinb(new_new_n9476__), .dout(new_new_n5851__));
  or1   g2753(.dina(new_new_n5851__), .dinb(new_new_n5847__), .dout(new_new_n5852__));
  or1   g2754(.dina(new_new_n5852__), .dinb(new_new_n9477__), .dout(new_new_n5853__));
  or1   g2755(.dina(new_new_n8831__), .dinb(new_new_n8782__), .dout(new_new_n5854__));
  or1   g2756(.dina(new_new_n5854__), .dinb(new_new_n9478__), .dout(new_new_n5855__));
  or1   g2757(.dina(new_new_n8832__), .dinb(new_new_n8781__), .dout(new_new_n5856__));
  or1   g2758(.dina(new_new_n5856__), .dinb(new_new_n9479__), .dout(new_new_n5857__));
  and1  g2759(.dina(new_new_n5857__), .dinb(new_new_n5855__), .dout(new_new_n5858__));
  and1  g2760(.dina(new_new_n3889__), .dinb(new_new_n9479__), .dout(new_new_n5859__));
  and1  g2761(.dina(new_new_n3891__), .dinb(new_new_n9478__), .dout(new_new_n5860__));
  or1   g2762(.dina(new_new_n5860__), .dinb(new_new_n5859__), .dout(new_new_n5861__));
  or1   g2763(.dina(new_new_n5861__), .dinb(new_new_n3572__), .dout(new_new_n5862__));
  and1  g2764(.dina(new_new_n5862__), .dinb(new_new_n5858__), .dout(new_new_n5863__));
  and1  g2765(.dina(new_new_n5863__), .dinb(new_new_n8862__), .dout(new_new_n5864__));
  and1  g2766(.dina(new_new_n5864__), .dinb(new_new_n8902__), .dout(new_new_n5865__));
  and1  g2767(.dina(new_new_n9227__), .dinb(new_new_n8933__), .dout(new_new_n5866__));
  and1  g2768(.dina(new_new_n5866__), .dinb(new_new_n8904__), .dout(new_new_n5867__));
  and1  g2769(.dina(new_new_n8864__), .dinb(new_new_n3050__), .dout(new_new_n5868__));
  and1  g2770(.dina(new_new_n5868__), .dinb(new_new_n8956__), .dout(new_new_n5869__));
  or1   g2771(.dina(new_new_n5867__), .dinb(new_new_n5865__), .dout(new_new_n5870__));
  or1   g2772(.dina(new_new_n5870__), .dinb(new_new_n5869__), .dout(new_new_n5871__));
  and1  g2773(.dina(new_new_n8581__), .dinb(new_new_n8864__), .dout(new_new_n5872__));
  and1  g2774(.dina(new_new_n5872__), .dinb(new_new_n8904__), .dout(new_new_n5873__));
  and1  g2775(.dina(new_new_n9226__), .dinb(new_new_n8933__), .dout(new_new_n5874__));
  and1  g2776(.dina(new_new_n5874__), .dinb(new_new_n8905__), .dout(new_new_n5875__));
  and1  g2777(.dina(new_new_n8865__), .dinb(new_new_n3042__), .dout(new_new_n5876__));
  and1  g2778(.dina(new_new_n5876__), .dinb(new_new_n8956__), .dout(new_new_n5877__));
  or1   g2779(.dina(new_new_n5875__), .dinb(new_new_n5873__), .dout(new_new_n5878__));
  or1   g2780(.dina(new_new_n5878__), .dinb(new_new_n5877__), .dout(new_new_n5879__));
  and1  g2781(.dina(new_new_n8580__), .dinb(new_new_n8865__), .dout(new_new_n5880__));
  and1  g2782(.dina(new_new_n5880__), .dinb(new_new_n8905__), .dout(new_new_n5881__));
  and1  g2783(.dina(new_new_n9225__), .dinb(new_new_n8936__), .dout(new_new_n5882__));
  and1  g2784(.dina(new_new_n5882__), .dinb(new_new_n8908__), .dout(new_new_n5883__));
  and1  g2785(.dina(new_new_n8868__), .dinb(new_new_n2842__), .dout(new_new_n5884__));
  and1  g2786(.dina(new_new_n5884__), .dinb(new_new_n8959__), .dout(new_new_n5885__));
  or1   g2787(.dina(new_new_n5883__), .dinb(new_new_n5881__), .dout(new_new_n5886__));
  or1   g2788(.dina(new_new_n5886__), .dinb(new_new_n5885__), .dout(new_new_n5887__));
  and1  g2789(.dina(new_new_n8578__), .dinb(new_new_n8868__), .dout(new_new_n5888__));
  and1  g2790(.dina(new_new_n5888__), .dinb(new_new_n8908__), .dout(new_new_n5889__));
  and1  g2791(.dina(new_new_n9224__), .dinb(new_new_n8936__), .dout(new_new_n5890__));
  and1  g2792(.dina(new_new_n5890__), .dinb(new_new_n8909__), .dout(new_new_n5891__));
  and1  g2793(.dina(new_new_n8869__), .dinb(new_new_n3034__), .dout(new_new_n5892__));
  and1  g2794(.dina(new_new_n5892__), .dinb(new_new_n8959__), .dout(new_new_n5893__));
  or1   g2795(.dina(new_new_n5891__), .dinb(new_new_n5889__), .dout(new_new_n5894__));
  or1   g2796(.dina(new_new_n5894__), .dinb(new_new_n5893__), .dout(new_new_n5895__));
  and1  g2797(.dina(new_new_n9482__), .dinb(new_new_n9095__), .dout(new_new_n5896__));
  and1  g2798(.dina(new_new_n5896__), .dinb(new_new_n9114__), .dout(new_new_n5897__));
  and1  g2799(.dina(new_new_n9486__), .dinb(new_new_n9133__), .dout(new_new_n5898__));
  and1  g2800(.dina(new_new_n5898__), .dinb(new_new_n9114__), .dout(new_new_n5899__));
  and1  g2801(.dina(new_new_n9095__), .dinb(new_new_n9488__), .dout(new_new_n5900__));
  and1  g2802(.dina(new_new_n5900__), .dinb(new_new_n9152__), .dout(new_new_n5901__));
  and1  g2803(.dina(new_new_n9133__), .dinb(new_new_n9489__), .dout(new_new_n5902__));
  and1  g2804(.dina(new_new_n5902__), .dinb(new_new_n9152__), .dout(new_new_n5903__));
  or1   g2805(.dina(new_new_n5899__), .dinb(new_new_n5897__), .dout(new_new_n5904__));
  or1   g2806(.dina(new_new_n5904__), .dinb(new_new_n5901__), .dout(new_new_n5905__));
  or1   g2807(.dina(new_new_n5905__), .dinb(new_new_n5903__), .dout(new_new_n5906__));
  and1  g2808(.dina(new_new_n9482__), .dinb(new_new_n9004__), .dout(new_new_n5907__));
  and1  g2809(.dina(new_new_n5907__), .dinb(new_new_n9023__), .dout(new_new_n5908__));
  and1  g2810(.dina(new_new_n9486__), .dinb(new_new_n9046__), .dout(new_new_n5909__));
  and1  g2811(.dina(new_new_n5909__), .dinb(new_new_n9023__), .dout(new_new_n5910__));
  and1  g2812(.dina(new_new_n9004__), .dinb(new_new_n9488__), .dout(new_new_n5911__));
  and1  g2813(.dina(new_new_n5911__), .dinb(new_new_n9066__), .dout(new_new_n5912__));
  and1  g2814(.dina(new_new_n9046__), .dinb(new_new_n9489__), .dout(new_new_n5913__));
  and1  g2815(.dina(new_new_n5913__), .dinb(new_new_n9066__), .dout(new_new_n5914__));
  or1   g2816(.dina(new_new_n5910__), .dinb(new_new_n5908__), .dout(new_new_n5915__));
  or1   g2817(.dina(new_new_n5915__), .dinb(new_new_n5912__), .dout(new_new_n5916__));
  or1   g2818(.dina(new_new_n5916__), .dinb(new_new_n5914__), .dout(new_new_n5917__));
  and1  g2819(.dina(new_new_n9492__), .dinb(new_new_n9007__), .dout(new_new_n5918__));
  and1  g2820(.dina(new_new_n5918__), .dinb(new_new_n9026__), .dout(new_new_n5919__));
  and1  g2821(.dina(new_new_n9496__), .dinb(new_new_n9049__), .dout(new_new_n5920__));
  and1  g2822(.dina(new_new_n5920__), .dinb(new_new_n9026__), .dout(new_new_n5921__));
  and1  g2823(.dina(new_new_n9007__), .dinb(new_new_n9498__), .dout(new_new_n5922__));
  and1  g2824(.dina(new_new_n5922__), .dinb(new_new_n9069__), .dout(new_new_n5923__));
  and1  g2825(.dina(new_new_n9049__), .dinb(new_new_n9499__), .dout(new_new_n5924__));
  and1  g2826(.dina(new_new_n5924__), .dinb(new_new_n9069__), .dout(new_new_n5925__));
  or1   g2827(.dina(new_new_n5921__), .dinb(new_new_n5919__), .dout(new_new_n5926__));
  or1   g2828(.dina(new_new_n5926__), .dinb(new_new_n5923__), .dout(new_new_n5927__));
  or1   g2829(.dina(new_new_n5927__), .dinb(new_new_n5925__), .dout(new_new_n5928__));
  and1  g2830(.dina(new_new_n9502__), .dinb(new_new_n9008__), .dout(new_new_n5929__));
  and1  g2831(.dina(new_new_n5929__), .dinb(new_new_n9027__), .dout(new_new_n5930__));
  and1  g2832(.dina(new_new_n9506__), .dinb(new_new_n9050__), .dout(new_new_n5931__));
  and1  g2833(.dina(new_new_n5931__), .dinb(new_new_n9027__), .dout(new_new_n5932__));
  and1  g2834(.dina(new_new_n9008__), .dinb(new_new_n9508__), .dout(new_new_n5933__));
  and1  g2835(.dina(new_new_n5933__), .dinb(new_new_n9070__), .dout(new_new_n5934__));
  and1  g2836(.dina(new_new_n9050__), .dinb(new_new_n9509__), .dout(new_new_n5935__));
  and1  g2837(.dina(new_new_n5935__), .dinb(new_new_n9070__), .dout(new_new_n5936__));
  or1   g2838(.dina(new_new_n5932__), .dinb(new_new_n5930__), .dout(new_new_n5937__));
  or1   g2839(.dina(new_new_n5937__), .dinb(new_new_n5934__), .dout(new_new_n5938__));
  or1   g2840(.dina(new_new_n5938__), .dinb(new_new_n5936__), .dout(new_new_n5939__));
  and1  g2841(.dina(new_new_n9512__), .dinb(new_new_n9010__), .dout(new_new_n5940__));
  and1  g2842(.dina(new_new_n5940__), .dinb(new_new_n9029__), .dout(new_new_n5941__));
  and1  g2843(.dina(new_new_n9516__), .dinb(new_new_n9052__), .dout(new_new_n5942__));
  and1  g2844(.dina(new_new_n5942__), .dinb(new_new_n9029__), .dout(new_new_n5943__));
  and1  g2845(.dina(new_new_n9010__), .dinb(new_new_n9518__), .dout(new_new_n5944__));
  and1  g2846(.dina(new_new_n5944__), .dinb(new_new_n9072__), .dout(new_new_n5945__));
  and1  g2847(.dina(new_new_n9052__), .dinb(new_new_n9519__), .dout(new_new_n5946__));
  and1  g2848(.dina(new_new_n5946__), .dinb(new_new_n9072__), .dout(new_new_n5947__));
  or1   g2849(.dina(new_new_n5943__), .dinb(new_new_n5941__), .dout(new_new_n5948__));
  or1   g2850(.dina(new_new_n5948__), .dinb(new_new_n5945__), .dout(new_new_n5949__));
  or1   g2851(.dina(new_new_n5949__), .dinb(new_new_n5947__), .dout(new_new_n5950__));
  and1  g2852(.dina(new_new_n9492__), .dinb(new_new_n9098__), .dout(new_new_n5951__));
  and1  g2853(.dina(new_new_n5951__), .dinb(new_new_n9117__), .dout(new_new_n5952__));
  and1  g2854(.dina(new_new_n9496__), .dinb(new_new_n9136__), .dout(new_new_n5953__));
  and1  g2855(.dina(new_new_n5953__), .dinb(new_new_n9117__), .dout(new_new_n5954__));
  and1  g2856(.dina(new_new_n9098__), .dinb(new_new_n9498__), .dout(new_new_n5955__));
  and1  g2857(.dina(new_new_n5955__), .dinb(new_new_n9155__), .dout(new_new_n5956__));
  and1  g2858(.dina(new_new_n9136__), .dinb(new_new_n9499__), .dout(new_new_n5957__));
  and1  g2859(.dina(new_new_n5957__), .dinb(new_new_n9155__), .dout(new_new_n5958__));
  or1   g2860(.dina(new_new_n5954__), .dinb(new_new_n5952__), .dout(new_new_n5959__));
  or1   g2861(.dina(new_new_n5959__), .dinb(new_new_n5956__), .dout(new_new_n5960__));
  or1   g2862(.dina(new_new_n5960__), .dinb(new_new_n5958__), .dout(new_new_n5961__));
  and1  g2863(.dina(new_new_n9502__), .dinb(new_new_n9099__), .dout(new_new_n5962__));
  and1  g2864(.dina(new_new_n5962__), .dinb(new_new_n9118__), .dout(new_new_n5963__));
  and1  g2865(.dina(new_new_n9506__), .dinb(new_new_n9137__), .dout(new_new_n5964__));
  and1  g2866(.dina(new_new_n5964__), .dinb(new_new_n9118__), .dout(new_new_n5965__));
  and1  g2867(.dina(new_new_n9099__), .dinb(new_new_n9508__), .dout(new_new_n5966__));
  and1  g2868(.dina(new_new_n5966__), .dinb(new_new_n9156__), .dout(new_new_n5967__));
  and1  g2869(.dina(new_new_n9137__), .dinb(new_new_n9509__), .dout(new_new_n5968__));
  and1  g2870(.dina(new_new_n5968__), .dinb(new_new_n9156__), .dout(new_new_n5969__));
  or1   g2871(.dina(new_new_n5965__), .dinb(new_new_n5963__), .dout(new_new_n5970__));
  or1   g2872(.dina(new_new_n5970__), .dinb(new_new_n5967__), .dout(new_new_n5971__));
  or1   g2873(.dina(new_new_n5971__), .dinb(new_new_n5969__), .dout(new_new_n5972__));
  and1  g2874(.dina(new_new_n9512__), .dinb(new_new_n9101__), .dout(new_new_n5973__));
  and1  g2875(.dina(new_new_n5973__), .dinb(new_new_n9120__), .dout(new_new_n5974__));
  and1  g2876(.dina(new_new_n9516__), .dinb(new_new_n9139__), .dout(new_new_n5975__));
  and1  g2877(.dina(new_new_n5975__), .dinb(new_new_n9120__), .dout(new_new_n5976__));
  and1  g2878(.dina(new_new_n9101__), .dinb(new_new_n9518__), .dout(new_new_n5977__));
  and1  g2879(.dina(new_new_n5977__), .dinb(new_new_n9158__), .dout(new_new_n5978__));
  and1  g2880(.dina(new_new_n9139__), .dinb(new_new_n9519__), .dout(new_new_n5979__));
  and1  g2881(.dina(new_new_n5979__), .dinb(new_new_n9158__), .dout(new_new_n5980__));
  or1   g2882(.dina(new_new_n5976__), .dinb(new_new_n5974__), .dout(new_new_n5981__));
  or1   g2883(.dina(new_new_n5981__), .dinb(new_new_n5978__), .dout(new_new_n5982__));
  or1   g2884(.dina(new_new_n5982__), .dinb(new_new_n5980__), .dout(new_new_n5983__));
  and1  g2885(.dina(new_new_n9511__), .dinb(new_new_n9245__), .dout(new_new_n5984__));
  and1  g2886(.dina(new_new_n5984__), .dinb(new_new_n9264__), .dout(new_new_n5985__));
  and1  g2887(.dina(new_new_n9515__), .dinb(new_new_n9283__), .dout(new_new_n5986__));
  and1  g2888(.dina(new_new_n5986__), .dinb(new_new_n9264__), .dout(new_new_n5987__));
  and1  g2889(.dina(new_new_n9245__), .dinb(new_new_n9520__), .dout(new_new_n5988__));
  and1  g2890(.dina(new_new_n5988__), .dinb(new_new_n9303__), .dout(new_new_n5989__));
  and1  g2891(.dina(new_new_n9283__), .dinb(new_new_n9521__), .dout(new_new_n5990__));
  and1  g2892(.dina(new_new_n5990__), .dinb(new_new_n9303__), .dout(new_new_n5991__));
  or1   g2893(.dina(new_new_n5987__), .dinb(new_new_n5985__), .dout(new_new_n5992__));
  or1   g2894(.dina(new_new_n5992__), .dinb(new_new_n5989__), .dout(new_new_n5993__));
  or1   g2895(.dina(new_new_n5993__), .dinb(new_new_n5991__), .dout(new_new_n5994__));
  and1  g2896(.dina(new_new_n5994__), .dinb(new_new_n9322__), .dout(new_new_n5995__));
  and1  g2897(.dina(new_new_n9501__), .dinb(new_new_n9248__), .dout(new_new_n5996__));
  and1  g2898(.dina(new_new_n5996__), .dinb(new_new_n9267__), .dout(new_new_n5997__));
  and1  g2899(.dina(new_new_n9505__), .dinb(new_new_n9286__), .dout(new_new_n5998__));
  and1  g2900(.dina(new_new_n5998__), .dinb(new_new_n9267__), .dout(new_new_n5999__));
  and1  g2901(.dina(new_new_n9248__), .dinb(new_new_n9522__), .dout(new_new_n6000__));
  and1  g2902(.dina(new_new_n6000__), .dinb(new_new_n9306__), .dout(new_new_n6001__));
  and1  g2903(.dina(new_new_n9286__), .dinb(new_new_n9523__), .dout(new_new_n6002__));
  and1  g2904(.dina(new_new_n6002__), .dinb(new_new_n9306__), .dout(new_new_n6003__));
  or1   g2905(.dina(new_new_n5999__), .dinb(new_new_n5997__), .dout(new_new_n6004__));
  or1   g2906(.dina(new_new_n6004__), .dinb(new_new_n6001__), .dout(new_new_n6005__));
  or1   g2907(.dina(new_new_n6005__), .dinb(new_new_n6003__), .dout(new_new_n6006__));
  and1  g2908(.dina(new_new_n6006__), .dinb(new_new_n9324__), .dout(new_new_n6007__));
  and1  g2909(.dina(new_new_n9491__), .dinb(new_new_n9249__), .dout(new_new_n6008__));
  and1  g2910(.dina(new_new_n6008__), .dinb(new_new_n9268__), .dout(new_new_n6009__));
  and1  g2911(.dina(new_new_n9495__), .dinb(new_new_n9287__), .dout(new_new_n6010__));
  and1  g2912(.dina(new_new_n6010__), .dinb(new_new_n9268__), .dout(new_new_n6011__));
  and1  g2913(.dina(new_new_n9249__), .dinb(new_new_n9524__), .dout(new_new_n6012__));
  and1  g2914(.dina(new_new_n6012__), .dinb(new_new_n9307__), .dout(new_new_n6013__));
  and1  g2915(.dina(new_new_n9287__), .dinb(new_new_n9525__), .dout(new_new_n6014__));
  and1  g2916(.dina(new_new_n6014__), .dinb(new_new_n9307__), .dout(new_new_n6015__));
  or1   g2917(.dina(new_new_n6011__), .dinb(new_new_n6009__), .dout(new_new_n6016__));
  or1   g2918(.dina(new_new_n6016__), .dinb(new_new_n6013__), .dout(new_new_n6017__));
  or1   g2919(.dina(new_new_n6017__), .dinb(new_new_n6015__), .dout(new_new_n6018__));
  and1  g2920(.dina(new_new_n6018__), .dinb(new_new_n9324__), .dout(new_new_n6019__));
  and1  g2921(.dina(new_new_n9481__), .dinb(new_new_n9251__), .dout(new_new_n6020__));
  and1  g2922(.dina(new_new_n6020__), .dinb(new_new_n9270__), .dout(new_new_n6021__));
  and1  g2923(.dina(new_new_n9485__), .dinb(new_new_n9289__), .dout(new_new_n6022__));
  and1  g2924(.dina(new_new_n6022__), .dinb(new_new_n9270__), .dout(new_new_n6023__));
  and1  g2925(.dina(new_new_n9251__), .dinb(new_new_n9526__), .dout(new_new_n6024__));
  and1  g2926(.dina(new_new_n6024__), .dinb(new_new_n9309__), .dout(new_new_n6025__));
  and1  g2927(.dina(new_new_n9289__), .dinb(new_new_n9527__), .dout(new_new_n6026__));
  and1  g2928(.dina(new_new_n6026__), .dinb(new_new_n9309__), .dout(new_new_n6027__));
  or1   g2929(.dina(new_new_n6023__), .dinb(new_new_n6021__), .dout(new_new_n6028__));
  or1   g2930(.dina(new_new_n6028__), .dinb(new_new_n6025__), .dout(new_new_n6029__));
  or1   g2931(.dina(new_new_n6029__), .dinb(new_new_n6027__), .dout(new_new_n6030__));
  and1  g2932(.dina(new_new_n6030__), .dinb(new_new_n9327__), .dout(new_new_n6031__));
  and1  g2933(.dina(new_new_n9513__), .dinb(new_new_n9343__), .dout(new_new_n6032__));
  and1  g2934(.dina(new_new_n6032__), .dinb(new_new_n9362__), .dout(new_new_n6033__));
  and1  g2935(.dina(new_new_n9517__), .dinb(new_new_n9381__), .dout(new_new_n6034__));
  and1  g2936(.dina(new_new_n6034__), .dinb(new_new_n9362__), .dout(new_new_n6035__));
  and1  g2937(.dina(new_new_n9343__), .dinb(new_new_n9520__), .dout(new_new_n6036__));
  and1  g2938(.dina(new_new_n6036__), .dinb(new_new_n9400__), .dout(new_new_n6037__));
  and1  g2939(.dina(new_new_n9381__), .dinb(new_new_n9521__), .dout(new_new_n6038__));
  and1  g2940(.dina(new_new_n6038__), .dinb(new_new_n9400__), .dout(new_new_n6039__));
  or1   g2941(.dina(new_new_n6035__), .dinb(new_new_n6033__), .dout(new_new_n6040__));
  or1   g2942(.dina(new_new_n6040__), .dinb(new_new_n6037__), .dout(new_new_n6041__));
  or1   g2943(.dina(new_new_n6041__), .dinb(new_new_n6039__), .dout(new_new_n6042__));
  and1  g2944(.dina(new_new_n6042__), .dinb(new_new_n9327__), .dout(new_new_n6043__));
  and1  g2945(.dina(new_new_n9503__), .dinb(new_new_n9346__), .dout(new_new_n6044__));
  and1  g2946(.dina(new_new_n6044__), .dinb(new_new_n9365__), .dout(new_new_n6045__));
  and1  g2947(.dina(new_new_n9507__), .dinb(new_new_n9384__), .dout(new_new_n6046__));
  and1  g2948(.dina(new_new_n6046__), .dinb(new_new_n9365__), .dout(new_new_n6047__));
  and1  g2949(.dina(new_new_n9346__), .dinb(new_new_n9522__), .dout(new_new_n6048__));
  and1  g2950(.dina(new_new_n6048__), .dinb(new_new_n9403__), .dout(new_new_n6049__));
  and1  g2951(.dina(new_new_n9384__), .dinb(new_new_n9523__), .dout(new_new_n6050__));
  and1  g2952(.dina(new_new_n6050__), .dinb(new_new_n9403__), .dout(new_new_n6051__));
  or1   g2953(.dina(new_new_n6047__), .dinb(new_new_n6045__), .dout(new_new_n6052__));
  or1   g2954(.dina(new_new_n6052__), .dinb(new_new_n6049__), .dout(new_new_n6053__));
  or1   g2955(.dina(new_new_n6053__), .dinb(new_new_n6051__), .dout(new_new_n6054__));
  and1  g2956(.dina(new_new_n6054__), .dinb(new_new_n9328__), .dout(new_new_n6055__));
  and1  g2957(.dina(new_new_n9493__), .dinb(new_new_n9347__), .dout(new_new_n6056__));
  and1  g2958(.dina(new_new_n6056__), .dinb(new_new_n9366__), .dout(new_new_n6057__));
  and1  g2959(.dina(new_new_n9497__), .dinb(new_new_n9385__), .dout(new_new_n6058__));
  and1  g2960(.dina(new_new_n6058__), .dinb(new_new_n9366__), .dout(new_new_n6059__));
  and1  g2961(.dina(new_new_n9347__), .dinb(new_new_n9524__), .dout(new_new_n6060__));
  and1  g2962(.dina(new_new_n6060__), .dinb(new_new_n9404__), .dout(new_new_n6061__));
  and1  g2963(.dina(new_new_n9385__), .dinb(new_new_n9525__), .dout(new_new_n6062__));
  and1  g2964(.dina(new_new_n6062__), .dinb(new_new_n9404__), .dout(new_new_n6063__));
  or1   g2965(.dina(new_new_n6059__), .dinb(new_new_n6057__), .dout(new_new_n6064__));
  or1   g2966(.dina(new_new_n6064__), .dinb(new_new_n6061__), .dout(new_new_n6065__));
  or1   g2967(.dina(new_new_n6065__), .dinb(new_new_n6063__), .dout(new_new_n6066__));
  and1  g2968(.dina(new_new_n6066__), .dinb(new_new_n9328__), .dout(new_new_n6067__));
  and1  g2969(.dina(new_new_n9483__), .dinb(new_new_n9349__), .dout(new_new_n6068__));
  and1  g2970(.dina(new_new_n6068__), .dinb(new_new_n9368__), .dout(new_new_n6069__));
  and1  g2971(.dina(new_new_n9487__), .dinb(new_new_n9387__), .dout(new_new_n6070__));
  and1  g2972(.dina(new_new_n6070__), .dinb(new_new_n9368__), .dout(new_new_n6071__));
  and1  g2973(.dina(new_new_n9349__), .dinb(new_new_n9526__), .dout(new_new_n6072__));
  and1  g2974(.dina(new_new_n6072__), .dinb(new_new_n9406__), .dout(new_new_n6073__));
  and1  g2975(.dina(new_new_n9387__), .dinb(new_new_n9527__), .dout(new_new_n6074__));
  and1  g2976(.dina(new_new_n6074__), .dinb(new_new_n9406__), .dout(new_new_n6075__));
  or1   g2977(.dina(new_new_n6071__), .dinb(new_new_n6069__), .dout(new_new_n6076__));
  or1   g2978(.dina(new_new_n6076__), .dinb(new_new_n6073__), .dout(new_new_n6077__));
  or1   g2979(.dina(new_new_n6077__), .dinb(new_new_n6075__), .dout(new_new_n6078__));
  and1  g2980(.dina(new_new_n6078__), .dinb(new_new_n9330__), .dout(new_new_n6079__));
  and1  g2981(.dina(new_new_n4449__), .dinb(new_new_n4435__), .dout(new_new_n6080__));
  and1  g2982(.dina(new_new_n4448__), .dinb(new_new_n4434__), .dout(new_new_n6081__));
  or1   g2983(.dina(new_new_n6081__), .dinb(new_new_n6080__), .dout(new_new_n6082__));
  or1   g2984(.dina(new_new_n9528__), .dinb(new_new_n8937__), .dout(new_new_n6083__));
  or1   g2985(.dina(new_new_n6083__), .dinb(new_new_n8960__), .dout(new_new_n6084__));
  or1   g2986(.dina(new_new_n4440__), .dinb(new_new_n4221__), .dout(new_new_n6085__));
  or1   g2987(.dina(new_new_n4442__), .dinb(new_new_n4219__), .dout(new_new_n6086__));
  and1  g2988(.dina(new_new_n6086__), .dinb(new_new_n6085__), .dout(new_new_n6087__));
  or1   g2989(.dina(new_new_n9529__), .dinb(new_new_n8869__), .dout(new_new_n6088__));
  or1   g2990(.dina(new_new_n6088__), .dinb(new_new_n8960__), .dout(new_new_n6089__));
  or1   g2991(.dina(new_new_n8937__), .dinb(new_new_n3091__), .dout(new_new_n6090__));
  or1   g2992(.dina(new_new_n6090__), .dinb(new_new_n8909__), .dout(new_new_n6091__));
  or1   g2993(.dina(new_new_n8911__), .dinb(new_new_n8871__), .dout(new_new_n6092__));
  and1  g2994(.dina(new_new_n6089__), .dinb(new_new_n6084__), .dout(new_new_n6093__));
  and1  g2995(.dina(new_new_n6093__), .dinb(new_new_n6091__), .dout(new_new_n6094__));
  and1  g2996(.dina(new_new_n6094__), .dinb(new_new_n9530__), .dout(new_new_n6095__));
  and1  g2997(.dina(new_new_n4446__), .dinb(new_new_n4433__), .dout(new_new_n6096__));
  and1  g2998(.dina(new_new_n4447__), .dinb(new_new_n4432__), .dout(new_new_n6097__));
  or1   g2999(.dina(new_new_n6097__), .dinb(new_new_n6096__), .dout(new_new_n6098__));
  or1   g3000(.dina(new_new_n9531__), .dinb(new_new_n8939__), .dout(new_new_n6099__));
  or1   g3001(.dina(new_new_n6099__), .dinb(new_new_n8962__), .dout(new_new_n6100__));
  or1   g3002(.dina(new_new_n4437__), .dinb(new_new_n4217__), .dout(new_new_n6101__));
  or1   g3003(.dina(new_new_n4438__), .dinb(new_new_n4214__), .dout(new_new_n6102__));
  and1  g3004(.dina(new_new_n6102__), .dinb(new_new_n6101__), .dout(new_new_n6103__));
  or1   g3005(.dina(new_new_n9532__), .dinb(new_new_n8871__), .dout(new_new_n6104__));
  or1   g3006(.dina(new_new_n6104__), .dinb(new_new_n8962__), .dout(new_new_n6105__));
  or1   g3007(.dina(new_new_n8939__), .dinb(new_new_n3075__), .dout(new_new_n6106__));
  or1   g3008(.dina(new_new_n6106__), .dinb(new_new_n8911__), .dout(new_new_n6107__));
  and1  g3009(.dina(new_new_n6105__), .dinb(new_new_n6100__), .dout(new_new_n6108__));
  and1  g3010(.dina(new_new_n6108__), .dinb(new_new_n6107__), .dout(new_new_n6109__));
  and1  g3011(.dina(new_new_n6109__), .dinb(new_new_n9530__), .dout(new_new_n6110__));
  and1  g3012(.dina(new_new_n9528__), .dinb(new_new_n8872__), .dout(new_new_n6111__));
  and1  g3013(.dina(new_new_n9529__), .dinb(new_new_n8940__), .dout(new_new_n6112__));
  or1   g3014(.dina(new_new_n6112__), .dinb(new_new_n6111__), .dout(new_new_n6113__));
  and1  g3015(.dina(new_new_n6113__), .dinb(new_new_n8912__), .dout(new_new_n6114__));
  and1  g3016(.dina(new_new_n8963__), .dinb(new_new_n2978__), .dout(new_new_n6115__));
  or1   g3017(.dina(new_new_n6115__), .dinb(new_new_n6114__), .dout(new_new_n6116__));
  and1  g3018(.dina(new_new_n9534__), .dinb(new_new_n9011__), .dout(new_new_n6117__));
  and1  g3019(.dina(new_new_n6117__), .dinb(new_new_n9030__), .dout(new_new_n6118__));
  and1  g3020(.dina(new_new_n9531__), .dinb(new_new_n8872__), .dout(new_new_n6119__));
  and1  g3021(.dina(new_new_n9532__), .dinb(new_new_n8940__), .dout(new_new_n6120__));
  or1   g3022(.dina(new_new_n6120__), .dinb(new_new_n6119__), .dout(new_new_n6121__));
  and1  g3023(.dina(new_new_n6121__), .dinb(new_new_n8912__), .dout(new_new_n6122__));
  and1  g3024(.dina(new_new_n8963__), .dinb(new_new_n2986__), .dout(new_new_n6123__));
  or1   g3025(.dina(new_new_n6123__), .dinb(new_new_n6122__), .dout(new_new_n6124__));
  and1  g3026(.dina(new_new_n9537__), .dinb(new_new_n9053__), .dout(new_new_n6125__));
  and1  g3027(.dina(new_new_n6125__), .dinb(new_new_n9030__), .dout(new_new_n6126__));
  and1  g3028(.dina(new_new_n9011__), .dinb(new_new_n9539__), .dout(new_new_n6127__));
  and1  g3029(.dina(new_new_n6127__), .dinb(new_new_n9073__), .dout(new_new_n6128__));
  and1  g3030(.dina(new_new_n9053__), .dinb(new_new_n9540__), .dout(new_new_n6129__));
  and1  g3031(.dina(new_new_n6129__), .dinb(new_new_n9073__), .dout(new_new_n6130__));
  or1   g3032(.dina(new_new_n6126__), .dinb(new_new_n6118__), .dout(new_new_n6131__));
  or1   g3033(.dina(new_new_n6131__), .dinb(new_new_n6128__), .dout(new_new_n6132__));
  or1   g3034(.dina(new_new_n6132__), .dinb(new_new_n6130__), .dout(new_new_n6133__));
  and1  g3035(.dina(new_new_n9534__), .dinb(new_new_n9102__), .dout(new_new_n6134__));
  and1  g3036(.dina(new_new_n6134__), .dinb(new_new_n9121__), .dout(new_new_n6135__));
  and1  g3037(.dina(new_new_n9537__), .dinb(new_new_n9140__), .dout(new_new_n6136__));
  and1  g3038(.dina(new_new_n6136__), .dinb(new_new_n9121__), .dout(new_new_n6137__));
  and1  g3039(.dina(new_new_n9102__), .dinb(new_new_n9539__), .dout(new_new_n6138__));
  and1  g3040(.dina(new_new_n6138__), .dinb(new_new_n9159__), .dout(new_new_n6139__));
  and1  g3041(.dina(new_new_n9140__), .dinb(new_new_n9540__), .dout(new_new_n6140__));
  and1  g3042(.dina(new_new_n6140__), .dinb(new_new_n9159__), .dout(new_new_n6141__));
  or1   g3043(.dina(new_new_n6137__), .dinb(new_new_n6135__), .dout(new_new_n6142__));
  or1   g3044(.dina(new_new_n6142__), .dinb(new_new_n6139__), .dout(new_new_n6143__));
  or1   g3045(.dina(new_new_n6143__), .dinb(new_new_n6141__), .dout(new_new_n6144__));
  and1  g3046(.dina(new_new_n9535__), .dinb(new_new_n9252__), .dout(new_new_n6145__));
  and1  g3047(.dina(new_new_n6145__), .dinb(new_new_n9271__), .dout(new_new_n6146__));
  and1  g3048(.dina(new_new_n9538__), .dinb(new_new_n9290__), .dout(new_new_n6147__));
  and1  g3049(.dina(new_new_n6147__), .dinb(new_new_n9271__), .dout(new_new_n6148__));
  and1  g3050(.dina(new_new_n9252__), .dinb(new_new_n9541__), .dout(new_new_n6149__));
  and1  g3051(.dina(new_new_n6149__), .dinb(new_new_n9310__), .dout(new_new_n6150__));
  and1  g3052(.dina(new_new_n9290__), .dinb(new_new_n9542__), .dout(new_new_n6151__));
  and1  g3053(.dina(new_new_n6151__), .dinb(new_new_n9310__), .dout(new_new_n6152__));
  or1   g3054(.dina(new_new_n6148__), .dinb(new_new_n6146__), .dout(new_new_n6153__));
  or1   g3055(.dina(new_new_n6153__), .dinb(new_new_n6150__), .dout(new_new_n6154__));
  or1   g3056(.dina(new_new_n6154__), .dinb(new_new_n6152__), .dout(new_new_n6155__));
  and1  g3057(.dina(new_new_n6155__), .dinb(new_new_n9330__), .dout(new_new_n6156__));
  and1  g3058(.dina(new_new_n9535__), .dinb(new_new_n9350__), .dout(new_new_n6157__));
  and1  g3059(.dina(new_new_n6157__), .dinb(new_new_n9369__), .dout(new_new_n6158__));
  and1  g3060(.dina(new_new_n9538__), .dinb(new_new_n9388__), .dout(new_new_n6159__));
  and1  g3061(.dina(new_new_n6159__), .dinb(new_new_n9369__), .dout(new_new_n6160__));
  and1  g3062(.dina(new_new_n9350__), .dinb(new_new_n9541__), .dout(new_new_n6161__));
  and1  g3063(.dina(new_new_n6161__), .dinb(new_new_n9407__), .dout(new_new_n6162__));
  and1  g3064(.dina(new_new_n9388__), .dinb(new_new_n9542__), .dout(new_new_n6163__));
  and1  g3065(.dina(new_new_n6163__), .dinb(new_new_n9407__), .dout(new_new_n6164__));
  or1   g3066(.dina(new_new_n6160__), .dinb(new_new_n6158__), .dout(new_new_n6165__));
  or1   g3067(.dina(new_new_n6165__), .dinb(new_new_n6162__), .dout(new_new_n6166__));
  or1   g3068(.dina(new_new_n6166__), .dinb(new_new_n6164__), .dout(new_new_n6167__));
  and1  g3069(.dina(new_new_n6167__), .dinb(new_new_n9331__), .dout(new_new_n6168__));
  and1  g3070(.dina(new_new_n4555__), .dinb(new_new_n4549__), .dout(new_new_n6169__));
  or1   g3071(.dina(new_new_n4554__), .dinb(new_new_n4548__), .dout(new_new_n6170__));
  and1  g3072(.dina(new_new_n9545__), .dinb(new_new_n9552__), .dout(new_new_n6171__));
  or1   g3073(.dina(new_new_n9557__), .dinb(new_new_n9563__), .dout(new_new_n6172__));
  and1  g3074(.dina(new_new_n6171__), .dinb(new_new_n4466__), .dout(new_new_n6173__));
  or1   g3075(.dina(new_new_n6172__), .dinb(new_new_n4467__), .dout(new_new_n6174__));
  and1  g3076(.dina(new_new_n9567__), .dinb(new_new_n9552__), .dout(new_new_n6175__));
  or1   g3077(.dina(new_new_n9573__), .dinb(new_new_n9563__), .dout(new_new_n6176__));
  and1  g3078(.dina(new_new_n6175__), .dinb(new_new_n4599__), .dout(new_new_n6177__));
  or1   g3079(.dina(new_new_n6176__), .dinb(new_new_n4598__), .dout(new_new_n6178__));
  and1  g3080(.dina(new_new_n6178__), .dinb(new_new_n6174__), .dout(new_new_n6179__));
  or1   g3081(.dina(new_new_n6177__), .dinb(new_new_n6173__), .dout(new_new_n6180__));
  and1  g3082(.dina(new_new_n9580__), .dinb(new_new_n9585__), .dout(new_new_n6181__));
  or1   g3083(.dina(new_new_n9589__), .dinb(new_new_n9594__), .dout(new_new_n6182__));
  and1  g3084(.dina(new_new_n9597__), .dinb(new_new_n9594__), .dout(new_new_n6183__));
  or1   g3085(.dina(new_new_n9603__), .dinb(new_new_n9585__), .dout(new_new_n6184__));
  and1  g3086(.dina(new_new_n6184__), .dinb(new_new_n6182__), .dout(new_new_n6185__));
  or1   g3087(.dina(new_new_n6183__), .dinb(new_new_n6181__), .dout(new_new_n6186__));
  and1  g3088(.dina(new_new_n6185__), .dinb(new_new_n9564__), .dout(new_new_n6187__));
  or1   g3089(.dina(new_new_n6186__), .dinb(new_new_n9551__), .dout(new_new_n6188__));
  and1  g3090(.dina(new_new_n6188__), .dinb(new_new_n6179__), .dout(new_new_n6189__));
  or1   g3091(.dina(new_new_n6187__), .dinb(new_new_n6180__), .dout(new_new_n6190__));
  and1  g3092(.dina(new_new_n3958__), .dinb(new_new_n9608__), .dout(new_new_n6191__));
  or1   g3093(.dina(new_new_n3959__), .dinb(new_new_n9609__), .dout(new_new_n6192__));
  and1  g3094(.dina(new_new_n6191__), .dinb(new_new_n9612__), .dout(new_new_n6193__));
  or1   g3095(.dina(new_new_n6192__), .dinb(new_new_n9618__), .dout(new_new_n6194__));
  and1  g3096(.dina(new_new_n6193__), .dinb(new_new_n9624__), .dout(new_new_n6195__));
  or1   g3097(.dina(new_new_n6194__), .dinb(new_new_n9629__), .dout(new_new_n6196__));
  and1  g3098(.dina(new_new_n6195__), .dinb(new_new_n9634__), .dout(new_new_n6197__));
  or1   g3099(.dina(new_new_n6196__), .dinb(new_new_n9638__), .dout(new_new_n6198__));
  and1  g3100(.dina(new_new_n3987__), .dinb(new_new_n9640__), .dout(new_new_n6199__));
  or1   g3101(.dina(new_new_n3986__), .dinb(new_new_n9641__), .dout(new_new_n6200__));
  and1  g3102(.dina(new_new_n6199__), .dinb(new_new_n9644__), .dout(new_new_n6201__));
  or1   g3103(.dina(new_new_n6200__), .dinb(new_new_n9650__), .dout(new_new_n6202__));
  and1  g3104(.dina(new_new_n6201__), .dinb(new_new_n9656__), .dout(new_new_n6203__));
  or1   g3105(.dina(new_new_n6202__), .dinb(new_new_n9661__), .dout(new_new_n6204__));
  and1  g3106(.dina(new_new_n6203__), .dinb(new_new_n9666__), .dout(new_new_n6205__));
  or1   g3107(.dina(new_new_n6204__), .dinb(new_new_n9670__), .dout(new_new_n6206__));
  and1  g3108(.dina(new_new_n9673__), .dinb(new_new_n9676__), .dout(new_new_n6207__));
  or1   g3109(.dina(new_new_n9679__), .dinb(new_new_n9681__), .dout(new_new_n6208__));
  and1  g3110(.dina(new_new_n9634__), .dinb(new_new_n4016__), .dout(new_new_n6209__));
  or1   g3111(.dina(new_new_n9638__), .dinb(new_new_n4017__), .dout(new_new_n6210__));
  and1  g3112(.dina(new_new_n9633__), .dinb(new_new_n9624__), .dout(new_new_n6211__));
  or1   g3113(.dina(new_new_n9637__), .dinb(new_new_n9629__), .dout(new_new_n6212__));
  and1  g3114(.dina(new_new_n6211__), .dinb(new_new_n3954__), .dout(new_new_n6213__));
  or1   g3115(.dina(new_new_n6212__), .dinb(new_new_n3955__), .dout(new_new_n6214__));
  and1  g3116(.dina(new_new_n9635__), .dinb(new_new_n9612__), .dout(new_new_n6215__));
  or1   g3117(.dina(new_new_n9639__), .dinb(new_new_n9618__), .dout(new_new_n6216__));
  and1  g3118(.dina(new_new_n6215__), .dinb(new_new_n3934__), .dout(new_new_n6217__));
  or1   g3119(.dina(new_new_n6216__), .dinb(new_new_n3935__), .dout(new_new_n6218__));
  and1  g3120(.dina(new_new_n6217__), .dinb(new_new_n9625__), .dout(new_new_n6219__));
  or1   g3121(.dina(new_new_n6218__), .dinb(new_new_n9630__), .dout(new_new_n6220__));
  and1  g3122(.dina(new_new_n9608__), .dinb(new_new_n9613__), .dout(new_new_n6221__));
  or1   g3123(.dina(new_new_n9609__), .dinb(new_new_n9619__), .dout(new_new_n6222__));
  and1  g3124(.dina(new_new_n6221__), .dinb(new_new_n9635__), .dout(new_new_n6223__));
  or1   g3125(.dina(new_new_n6222__), .dinb(new_new_n9639__), .dout(new_new_n6224__));
  and1  g3126(.dina(new_new_n6223__), .dinb(new_new_n3938__), .dout(new_new_n6225__));
  or1   g3127(.dina(new_new_n6224__), .dinb(new_new_n3939__), .dout(new_new_n6226__));
  and1  g3128(.dina(new_new_n6225__), .dinb(new_new_n9625__), .dout(new_new_n6227__));
  or1   g3129(.dina(new_new_n6226__), .dinb(new_new_n9630__), .dout(new_new_n6228__));
  and1  g3130(.dina(new_new_n6210__), .dinb(new_new_n6208__), .dout(new_new_n6229__));
  or1   g3131(.dina(new_new_n6209__), .dinb(new_new_n6207__), .dout(new_new_n6230__));
  and1  g3132(.dina(new_new_n6229__), .dinb(new_new_n6214__), .dout(new_new_n6231__));
  or1   g3133(.dina(new_new_n6230__), .dinb(new_new_n6213__), .dout(new_new_n6232__));
  and1  g3134(.dina(new_new_n6231__), .dinb(new_new_n6220__), .dout(new_new_n6233__));
  or1   g3135(.dina(new_new_n6232__), .dinb(new_new_n6219__), .dout(new_new_n6234__));
  and1  g3136(.dina(new_new_n6233__), .dinb(new_new_n6228__), .dout(new_new_n6235__));
  or1   g3137(.dina(new_new_n6234__), .dinb(new_new_n6227__), .dout(new_new_n6236__));
  and1  g3138(.dina(new_new_n9683__), .dinb(new_new_n9686__), .dout(new_new_n6237__));
  or1   g3139(.dina(new_new_n9689__), .dinb(new_new_n9691__), .dout(new_new_n6238__));
  and1  g3140(.dina(new_new_n9666__), .dinb(new_new_n4022__), .dout(new_new_n6239__));
  or1   g3141(.dina(new_new_n9670__), .dinb(new_new_n4023__), .dout(new_new_n6240__));
  and1  g3142(.dina(new_new_n9665__), .dinb(new_new_n9656__), .dout(new_new_n6241__));
  or1   g3143(.dina(new_new_n9669__), .dinb(new_new_n9661__), .dout(new_new_n6242__));
  and1  g3144(.dina(new_new_n6241__), .dinb(new_new_n3956__), .dout(new_new_n6243__));
  or1   g3145(.dina(new_new_n6242__), .dinb(new_new_n3957__), .dout(new_new_n6244__));
  and1  g3146(.dina(new_new_n9667__), .dinb(new_new_n9644__), .dout(new_new_n6245__));
  or1   g3147(.dina(new_new_n9671__), .dinb(new_new_n9650__), .dout(new_new_n6246__));
  and1  g3148(.dina(new_new_n6245__), .dinb(new_new_n3936__), .dout(new_new_n6247__));
  or1   g3149(.dina(new_new_n6246__), .dinb(new_new_n3937__), .dout(new_new_n6248__));
  and1  g3150(.dina(new_new_n6247__), .dinb(new_new_n9657__), .dout(new_new_n6249__));
  or1   g3151(.dina(new_new_n6248__), .dinb(new_new_n9662__), .dout(new_new_n6250__));
  and1  g3152(.dina(new_new_n9640__), .dinb(new_new_n9645__), .dout(new_new_n6251__));
  or1   g3153(.dina(new_new_n9641__), .dinb(new_new_n9651__), .dout(new_new_n6252__));
  and1  g3154(.dina(new_new_n6251__), .dinb(new_new_n9667__), .dout(new_new_n6253__));
  or1   g3155(.dina(new_new_n6252__), .dinb(new_new_n9671__), .dout(new_new_n6254__));
  and1  g3156(.dina(new_new_n6253__), .dinb(new_new_n3949__), .dout(new_new_n6255__));
  or1   g3157(.dina(new_new_n6254__), .dinb(new_new_n3948__), .dout(new_new_n6256__));
  and1  g3158(.dina(new_new_n6255__), .dinb(new_new_n9657__), .dout(new_new_n6257__));
  or1   g3159(.dina(new_new_n6256__), .dinb(new_new_n9662__), .dout(new_new_n6258__));
  and1  g3160(.dina(new_new_n6240__), .dinb(new_new_n6238__), .dout(new_new_n6259__));
  or1   g3161(.dina(new_new_n6239__), .dinb(new_new_n6237__), .dout(new_new_n6260__));
  and1  g3162(.dina(new_new_n6259__), .dinb(new_new_n6244__), .dout(new_new_n6261__));
  or1   g3163(.dina(new_new_n6260__), .dinb(new_new_n6243__), .dout(new_new_n6262__));
  and1  g3164(.dina(new_new_n6261__), .dinb(new_new_n6250__), .dout(new_new_n6263__));
  or1   g3165(.dina(new_new_n6262__), .dinb(new_new_n6249__), .dout(new_new_n6264__));
  and1  g3166(.dina(new_new_n6263__), .dinb(new_new_n6258__), .dout(new_new_n6265__));
  or1   g3167(.dina(new_new_n6264__), .dinb(new_new_n6257__), .dout(new_new_n6266__));
  and1  g3168(.dina(new_new_n9545__), .dinb(new_new_n9693__), .dout(new_new_n6267__));
  or1   g3169(.dina(new_new_n9557__), .dinb(new_new_n9695__), .dout(new_new_n6268__));
  and1  g3170(.dina(new_new_n9567__), .dinb(new_new_n9695__), .dout(new_new_n6269__));
  or1   g3171(.dina(new_new_n9573__), .dinb(new_new_n9693__), .dout(new_new_n6270__));
  and1  g3172(.dina(new_new_n6270__), .dinb(new_new_n6268__), .dout(new_new_n6271__));
  or1   g3173(.dina(new_new_n6269__), .dinb(new_new_n6267__), .dout(new_new_n6272__));
  and1  g3174(.dina(new_new_n4631__), .dinb(new_new_n4623__), .dout(new_new_n6273__));
  or1   g3175(.dina(new_new_n4630__), .dinb(new_new_n4622__), .dout(new_new_n6274__));
  and1  g3176(.dina(new_new_n4682__), .dinb(new_new_n4619__), .dout(new_new_n6275__));
  or1   g3177(.dina(new_new_n4683__), .dinb(new_new_n4618__), .dout(new_new_n6276__));
  and1  g3178(.dina(new_new_n4684__), .dinb(new_new_n4617__), .dout(new_new_n6277__));
  or1   g3179(.dina(new_new_n4685__), .dinb(new_new_n4616__), .dout(new_new_n6278__));
  and1  g3180(.dina(new_new_n6278__), .dinb(new_new_n6276__), .dout(new_new_n6279__));
  or1   g3181(.dina(new_new_n6277__), .dinb(new_new_n6275__), .dout(new_new_n6280__));
  and1  g3182(.dina(new_new_n9697__), .dinb(new_new_n9698__), .dout(new_new_n6281__));
  or1   g3183(.dina(new_new_n4483__), .dinb(new_new_n4481__), .dout(new_new_n6282__));
  and1  g3184(.dina(new_new_n9699__), .dinb(new_new_n9702__), .dout(new_new_n6283__));
  or1   g3185(.dina(new_new_n4135__), .dinb(new_new_n9704__), .dout(new_new_n6284__));
  and1  g3186(.dina(new_new_n9705__), .dinb(new_new_n3502__), .dout(new_new_n6285__));
  or1   g3187(.dina(new_new_n4098__), .dinb(new_new_n3503__), .dout(new_new_n6286__));
  and1  g3188(.dina(new_new_n6286__), .dinb(new_new_n6284__), .dout(new_new_n6287__));
  or1   g3189(.dina(new_new_n6285__), .dinb(new_new_n6283__), .dout(new_new_n6288__));
  and1  g3190(.dina(new_new_n9706__), .dinb(new_new_n9709__), .dout(new_new_n6289__));
  or1   g3191(.dina(new_new_n4137__), .dinb(new_new_n9711__), .dout(new_new_n6290__));
  and1  g3192(.dina(new_new_n9712__), .dinb(new_new_n3414__), .dout(new_new_n6291__));
  or1   g3193(.dina(new_new_n4100__), .dinb(new_new_n3415__), .dout(new_new_n6292__));
  and1  g3194(.dina(new_new_n6292__), .dinb(new_new_n6290__), .dout(new_new_n6293__));
  or1   g3195(.dina(new_new_n6291__), .dinb(new_new_n6289__), .dout(new_new_n6294__));
  and1  g3196(.dina(new_new_n9713__), .dinb(new_new_n9715__), .dout(new_new_n6295__));
  or1   g3197(.dina(new_new_n4689__), .dinb(new_new_n9716__), .dout(new_new_n6296__));
  and1  g3198(.dina(new_new_n9717__), .dinb(new_new_n9718__), .dout(new_new_n6297__));
  or1   g3199(.dina(new_new_n4691__), .dinb(new_new_n9720__), .dout(new_new_n6298__));
  and1  g3200(.dina(new_new_n6298__), .dinb(new_new_n6296__), .dout(new_new_n6299__));
  or1   g3201(.dina(new_new_n6297__), .dinb(new_new_n6295__), .dout(new_new_n6300__));
  and1  g3202(.dina(new_new_n9722__), .dinb(new_new_n9726__), .dout(new_new_n6301__));
  and1  g3203(.dina(new_new_n9731__), .dinb(new_new_n9734__), .dout(new_new_n6302__));
  or1   g3204(.dina(new_new_n9738__), .dinb(new_new_n9741__), .dout(new_new_n6303__));
  or1   g3205(.dina(new_new_n9744__), .dinb(new_new_n9747__), .dout(new_new_n6304__));
  and1  g3206(.dina(new_new_n9749__), .dinb(new_new_n9750__), .dout(new_new_n6305__));
  or1   g3207(.dina(new_new_n4677__), .dinb(new_new_n4673__), .dout(new_new_n6306__));
  and1  g3208(.dina(new_new_n9751__), .dinb(new_new_n9752__), .dout(new_new_n6307__));
  or1   g3209(.dina(new_new_n4681__), .dinb(new_new_n4669__), .dout(new_new_n6308__));
  and1  g3210(.dina(new_new_n9754__), .dinb(new_new_n9756__), .dout(new_new_n6309__));
  and1  g3211(.dina(new_new_n9758__), .dinb(new_new_n9761__), .dout(new_new_n6310__));
  or1   g3212(.dina(new_new_n6310__), .dinb(new_new_n6309__), .dout(new_new_n6311__));
  and1  g3213(.dina(new_new_n9731__), .dinb(new_new_n9765__), .dout(new_new_n6312__));
  and1  g3214(.dina(new_new_n9767__), .dinb(new_new_n9734__), .dout(new_new_n6313__));
  or1   g3215(.dina(new_new_n6313__), .dinb(new_new_n6312__), .dout(new_new_n6314__));
  and1  g3216(.dina(new_new_n9769__), .dinb(new_new_n9741__), .dout(new_new_n6315__));
  or1   g3217(.dina(new_new_n9738__), .dinb(new_new_n9773__), .dout(new_new_n6316__));
  and1  g3218(.dina(new_new_n9737__), .dinb(new_new_n9773__), .dout(new_new_n6317__));
  or1   g3219(.dina(new_new_n9769__), .dinb(new_new_n9742__), .dout(new_new_n6318__));
  and1  g3220(.dina(new_new_n6318__), .dinb(new_new_n6316__), .dout(new_new_n6319__));
  or1   g3221(.dina(new_new_n6317__), .dinb(new_new_n6315__), .dout(new_new_n6320__));
  and1  g3222(.dina(new_new_n9778__), .dinb(new_new_n9782__), .dout(new_new_n6321__));
  or1   g3223(.dina(new_new_n9785__), .dinb(new_new_n9788__), .dout(new_new_n6322__));
  and1  g3224(.dina(new_new_n9790__), .dinb(new_new_n9791__), .dout(new_new_n6323__));
  or1   g3225(.dina(new_new_n9792__), .dinb(new_new_n9793__), .dout(new_new_n6324__));
  and1  g3226(.dina(new_new_n9792__), .dinb(new_new_n9793__), .dout(new_new_n6325__));
  or1   g3227(.dina(new_new_n9790__), .dinb(new_new_n9791__), .dout(new_new_n6326__));
  and1  g3228(.dina(new_new_n6326__), .dinb(new_new_n6324__), .dout(new_new_n6327__));
  or1   g3229(.dina(new_new_n6325__), .dinb(new_new_n6323__), .dout(new_new_n6328__));
  and1  g3230(.dina(new_new_n9794__), .dinb(new_new_n9795__), .dout(new_new_n6329__));
  or1   g3231(.dina(new_new_n9796__), .dinb(new_new_n9797__), .dout(new_new_n6330__));
  and1  g3232(.dina(new_new_n9796__), .dinb(new_new_n9797__), .dout(new_new_n6331__));
  or1   g3233(.dina(new_new_n9794__), .dinb(new_new_n9795__), .dout(new_new_n6332__));
  and1  g3234(.dina(new_new_n6332__), .dinb(new_new_n6330__), .dout(new_new_n6333__));
  or1   g3235(.dina(new_new_n6331__), .dinb(new_new_n6329__), .dout(new_new_n6334__));
  and1  g3236(.dina(new_new_n9798__), .dinb(new_new_n9799__), .dout(new_new_n6335__));
  or1   g3237(.dina(new_new_n9800__), .dinb(new_new_n9801__), .dout(new_new_n6336__));
  and1  g3238(.dina(new_new_n9800__), .dinb(new_new_n9801__), .dout(new_new_n6337__));
  or1   g3239(.dina(new_new_n9798__), .dinb(new_new_n9799__), .dout(new_new_n6338__));
  and1  g3240(.dina(new_new_n6338__), .dinb(new_new_n6336__), .dout(new_new_n6339__));
  or1   g3241(.dina(new_new_n6337__), .dinb(new_new_n6335__), .dout(new_new_n6340__));
  and1  g3242(.dina(new_new_n9802__), .dinb(new_new_n9803__), .dout(new_new_n6341__));
  or1   g3243(.dina(new_new_n9804__), .dinb(new_new_n9805__), .dout(new_new_n6342__));
  and1  g3244(.dina(new_new_n9804__), .dinb(new_new_n9805__), .dout(new_new_n6343__));
  or1   g3245(.dina(new_new_n9802__), .dinb(new_new_n9803__), .dout(new_new_n6344__));
  and1  g3246(.dina(new_new_n6344__), .dinb(new_new_n6342__), .dout(new_new_n6345__));
  or1   g3247(.dina(new_new_n6343__), .dinb(new_new_n6341__), .dout(new_new_n6346__));
  and1  g3248(.dina(new_new_n9806__), .dinb(new_new_n9807__), .dout(new_new_n6347__));
  or1   g3249(.dina(new_new_n4675__), .dinb(new_new_n4671__), .dout(new_new_n6348__));
  and1  g3250(.dina(new_new_n9808__), .dinb(new_new_n9809__), .dout(new_new_n6349__));
  or1   g3251(.dina(new_new_n4679__), .dinb(new_new_n4667__), .dout(new_new_n6350__));
  and1  g3252(.dina(new_new_n9778__), .dinb(new_new_n9788__), .dout(new_new_n6351__));
  or1   g3253(.dina(new_new_n9785__), .dinb(new_new_n9782__), .dout(new_new_n6352__));
  and1  g3254(.dina(new_new_n9786__), .dinb(new_new_n9781__), .dout(new_new_n6353__));
  or1   g3255(.dina(new_new_n9777__), .dinb(new_new_n9789__), .dout(new_new_n6354__));
  and1  g3256(.dina(new_new_n6354__), .dinb(new_new_n6352__), .dout(new_new_n6355__));
  or1   g3257(.dina(new_new_n6353__), .dinb(new_new_n6351__), .dout(new_new_n6356__));
  and1  g3258(.dina(new_new_n9718__), .dinb(new_new_n9810__), .dout(new_new_n6357__));
  or1   g3259(.dina(new_new_n9720__), .dinb(new_new_n3505__), .dout(new_new_n6358__));
  and1  g3260(.dina(new_new_n6358__), .dinb(new_new_n9716__), .dout(new_new_n6359__));
  or1   g3261(.dina(new_new_n6357__), .dinb(new_new_n9715__), .dout(new_new_n6360__));
  and1  g3262(.dina(new_new_n9811__), .dinb(new_new_n9812__), .dout(new_new_n6361__));
  or1   g3263(.dina(new_new_n4507__), .dinb(new_new_n3441__), .dout(new_new_n6362__));
  and1  g3264(.dina(new_new_n4259__), .dinb(new_new_n3444__), .dout(new_new_n6363__));
  or1   g3265(.dina(new_new_n9813__), .dinb(new_new_n3445__), .dout(new_new_n6364__));
  and1  g3266(.dina(new_new_n6364__), .dinb(new_new_n6362__), .dout(new_new_n6365__));
  or1   g3267(.dina(new_new_n6363__), .dinb(new_new_n6361__), .dout(new_new_n6366__));
  and1  g3268(.dina(new_new_n9816__), .dinb(new_new_n9820__), .dout(new_new_n6367__));
  or1   g3269(.dina(new_new_n9823__), .dinb(new_new_n3483__), .dout(new_new_n6368__));
  and1  g3270(.dina(new_new_n9823__), .dinb(new_new_n3486__), .dout(new_new_n6369__));
  or1   g3271(.dina(new_new_n9816__), .dinb(new_new_n3487__), .dout(new_new_n6370__));
  and1  g3272(.dina(new_new_n6370__), .dinb(new_new_n6368__), .dout(new_new_n6371__));
  or1   g3273(.dina(new_new_n6369__), .dinb(new_new_n6367__), .dout(new_new_n6372__));
  and1  g3274(.dina(new_new_n9827__), .dinb(new_new_n9831__), .dout(new_new_n6373__));
  or1   g3275(.dina(new_new_n9834__), .dinb(new_new_n3395__), .dout(new_new_n6374__));
  and1  g3276(.dina(new_new_n9834__), .dinb(new_new_n3398__), .dout(new_new_n6375__));
  or1   g3277(.dina(new_new_n9827__), .dinb(new_new_n3399__), .dout(new_new_n6376__));
  and1  g3278(.dina(new_new_n6376__), .dinb(new_new_n6374__), .dout(new_new_n6377__));
  or1   g3279(.dina(new_new_n6375__), .dinb(new_new_n6373__), .dout(new_new_n6378__));
  and1  g3280(.dina(new_new_n9754__), .dinb(new_new_n9761__), .dout(new_new_n6379__));
  and1  g3281(.dina(new_new_n4607__), .dinb(new_new_n4297__), .dout(new_new_n6380__));
  or1   g3282(.dina(new_new_n4606__), .dinb(new_new_n4296__), .dout(new_new_n6381__));
  and1  g3283(.dina(new_new_n4584__), .dinb(new_new_n4474__), .dout(new_new_n6382__));
  or1   g3284(.dina(new_new_n4585__), .dinb(new_new_n4475__), .dout(new_new_n6383__));
  and1  g3285(.dina(new_new_n6383__), .dinb(new_new_n6381__), .dout(new_new_n6384__));
  or1   g3286(.dina(new_new_n6382__), .dinb(new_new_n6380__), .dout(new_new_n6385__));
  and1  g3287(.dina(new_new_n9836__), .dinb(new_new_n9838__), .dout(new_new_n6386__));
  or1   g3288(.dina(new_new_n9840__), .dinb(new_new_n9843__), .dout(new_new_n6387__));
  and1  g3289(.dina(new_new_n9840__), .dinb(new_new_n9843__), .dout(new_new_n6388__));
  or1   g3290(.dina(new_new_n9836__), .dinb(new_new_n9838__), .dout(new_new_n6389__));
  and1  g3291(.dina(new_new_n6389__), .dinb(new_new_n6387__), .dout(new_new_n6390__));
  or1   g3292(.dina(new_new_n6388__), .dinb(new_new_n6386__), .dout(new_new_n6391__));
  or1   g3293(.dina(new_new_n6391__), .dinb(new_new_n9846__), .dout(new_new_n6392__));
  or1   g3294(.dina(new_new_n6390__), .dinb(new_new_n9847__), .dout(new_new_n6393__));
  and1  g3295(.dina(new_new_n6393__), .dinb(new_new_n6392__), .dout(new_new_n6394__));
  or1   g3296(.dina(new_new_n9848__), .dinb(new_new_n9850__), .dout(new_new_n6395__));
  or1   g3297(.dina(new_new_n6395__), .dinb(new_new_n9852__), .dout(new_new_n6396__));
  and1  g3298(.dina(new_new_n4605__), .dinb(new_new_n4295__), .dout(new_new_n6397__));
  or1   g3299(.dina(new_new_n4604__), .dinb(new_new_n4294__), .dout(new_new_n6398__));
  and1  g3300(.dina(new_new_n4582__), .dinb(new_new_n4472__), .dout(new_new_n6399__));
  or1   g3301(.dina(new_new_n4583__), .dinb(new_new_n4473__), .dout(new_new_n6400__));
  and1  g3302(.dina(new_new_n6400__), .dinb(new_new_n6398__), .dout(new_new_n6401__));
  or1   g3303(.dina(new_new_n6399__), .dinb(new_new_n6397__), .dout(new_new_n6402__));
  and1  g3304(.dina(new_new_n9853__), .dinb(new_new_n9839__), .dout(new_new_n6403__));
  or1   g3305(.dina(new_new_n9854__), .dinb(new_new_n9842__), .dout(new_new_n6404__));
  and1  g3306(.dina(new_new_n9854__), .dinb(new_new_n9844__), .dout(new_new_n6405__));
  or1   g3307(.dina(new_new_n9853__), .dinb(new_new_n9839__), .dout(new_new_n6406__));
  and1  g3308(.dina(new_new_n6406__), .dinb(new_new_n6404__), .dout(new_new_n6407__));
  or1   g3309(.dina(new_new_n6405__), .dinb(new_new_n6403__), .dout(new_new_n6408__));
  or1   g3310(.dina(new_new_n6408__), .dinb(new_new_n9846__), .dout(new_new_n6409__));
  or1   g3311(.dina(new_new_n6407__), .dinb(new_new_n9847__), .dout(new_new_n6410__));
  and1  g3312(.dina(new_new_n6410__), .dinb(new_new_n6409__), .dout(new_new_n6411__));
  or1   g3313(.dina(new_new_n9855__), .dinb(new_new_n9856__), .dout(new_new_n6412__));
  or1   g3314(.dina(new_new_n6412__), .dinb(new_new_n9852__), .dout(new_new_n6413__));
  and1  g3315(.dina(new_new_n9856__), .dinb(new_new_n6198__), .dout(new_new_n6414__));
  or1   g3316(.dina(new_new_n9850__), .dinb(new_new_n9857__), .dout(new_new_n6415__));
  or1   g3317(.dina(new_new_n6415__), .dinb(new_new_n9848__), .dout(new_new_n6416__));
  or1   g3318(.dina(new_new_n6416__), .dinb(new_new_n9859__), .dout(new_new_n6417__));
  or1   g3319(.dina(new_new_n6414__), .dinb(new_new_n9855__), .dout(new_new_n6418__));
  or1   g3320(.dina(new_new_n6418__), .dinb(new_new_n9859__), .dout(new_new_n6419__));
  and1  g3321(.dina(new_new_n6413__), .dinb(new_new_n6396__), .dout(new_new_n6420__));
  and1  g3322(.dina(new_new_n6420__), .dinb(new_new_n6417__), .dout(new_new_n6421__));
  and1  g3323(.dina(new_new_n6421__), .dinb(new_new_n6419__), .dout(new_new_n6422__));
  and1  g3324(.dina(new_new_n4556__), .dinb(new_new_n4551__), .dout(new_new_n6423__));
  or1   g3325(.dina(new_new_n4557__), .dinb(new_new_n4550__), .dout(new_new_n6424__));
  and1  g3326(.dina(new_new_n9860__), .dinb(new_new_n9619__), .dout(new_new_n6425__));
  or1   g3327(.dina(new_new_n9861__), .dinb(new_new_n9613__), .dout(new_new_n6426__));
  and1  g3328(.dina(new_new_n9861__), .dinb(new_new_n9615__), .dout(new_new_n6427__));
  or1   g3329(.dina(new_new_n9860__), .dinb(new_new_n9621__), .dout(new_new_n6428__));
  and1  g3330(.dina(new_new_n6428__), .dinb(new_new_n6426__), .dout(new_new_n6429__));
  or1   g3331(.dina(new_new_n6427__), .dinb(new_new_n6425__), .dout(new_new_n6430__));
  or1   g3332(.dina(new_new_n6430__), .dinb(new_new_n9626__), .dout(new_new_n6431__));
  or1   g3333(.dina(new_new_n6429__), .dinb(new_new_n9631__), .dout(new_new_n6432__));
  and1  g3334(.dina(new_new_n6432__), .dinb(new_new_n6431__), .dout(new_new_n6433__));
  and1  g3335(.dina(new_new_n6433__), .dinb(new_new_n9858__), .dout(new_new_n6434__));
  and1  g3336(.dina(new_new_n4600__), .dinb(new_new_n4451__), .dout(new_new_n6435__));
  or1   g3337(.dina(new_new_n4601__), .dinb(new_new_n4450__), .dout(new_new_n6436__));
  and1  g3338(.dina(new_new_n4594__), .dinb(new_new_n4469__), .dout(new_new_n6437__));
  or1   g3339(.dina(new_new_n4595__), .dinb(new_new_n4468__), .dout(new_new_n6438__));
  and1  g3340(.dina(new_new_n6438__), .dinb(new_new_n6436__), .dout(new_new_n6439__));
  or1   g3341(.dina(new_new_n6437__), .dinb(new_new_n6435__), .dout(new_new_n6440__));
  and1  g3342(.dina(new_new_n9862__), .dinb(new_new_n9621__), .dout(new_new_n6441__));
  or1   g3343(.dina(new_new_n9863__), .dinb(new_new_n9615__), .dout(new_new_n6442__));
  and1  g3344(.dina(new_new_n9863__), .dinb(new_new_n9614__), .dout(new_new_n6443__));
  or1   g3345(.dina(new_new_n9862__), .dinb(new_new_n9620__), .dout(new_new_n6444__));
  and1  g3346(.dina(new_new_n6444__), .dinb(new_new_n6442__), .dout(new_new_n6445__));
  or1   g3347(.dina(new_new_n6443__), .dinb(new_new_n6441__), .dout(new_new_n6446__));
  and1  g3348(.dina(new_new_n6445__), .dinb(new_new_n9631__), .dout(new_new_n6447__));
  and1  g3349(.dina(new_new_n6446__), .dinb(new_new_n9626__), .dout(new_new_n6448__));
  or1   g3350(.dina(new_new_n6448__), .dinb(new_new_n6447__), .dout(new_new_n6449__));
  and1  g3351(.dina(new_new_n6449__), .dinb(new_new_n9851__), .dout(new_new_n6450__));
  or1   g3352(.dina(new_new_n6450__), .dinb(new_new_n6434__), .dout(new_new_n6451__));
  and1  g3353(.dina(new_new_n4610__), .dinb(new_new_n4301__), .dout(new_new_n6452__));
  or1   g3354(.dina(new_new_n4611__), .dinb(new_new_n4300__), .dout(new_new_n6453__));
  and1  g3355(.dina(new_new_n4588__), .dinb(new_new_n4479__), .dout(new_new_n6454__));
  or1   g3356(.dina(new_new_n4589__), .dinb(new_new_n4478__), .dout(new_new_n6455__));
  and1  g3357(.dina(new_new_n6455__), .dinb(new_new_n6453__), .dout(new_new_n6456__));
  or1   g3358(.dina(new_new_n6454__), .dinb(new_new_n6452__), .dout(new_new_n6457__));
  and1  g3359(.dina(new_new_n9864__), .dinb(new_new_n9868__), .dout(new_new_n6458__));
  or1   g3360(.dina(new_new_n9874__), .dinb(new_new_n9876__), .dout(new_new_n6459__));
  and1  g3361(.dina(new_new_n9874__), .dinb(new_new_n9876__), .dout(new_new_n6460__));
  or1   g3362(.dina(new_new_n9864__), .dinb(new_new_n9868__), .dout(new_new_n6461__));
  and1  g3363(.dina(new_new_n6461__), .dinb(new_new_n6459__), .dout(new_new_n6462__));
  or1   g3364(.dina(new_new_n6460__), .dinb(new_new_n6458__), .dout(new_new_n6463__));
  and1  g3365(.dina(new_new_n6462__), .dinb(new_new_n9879__), .dout(new_new_n6464__));
  and1  g3366(.dina(new_new_n6463__), .dinb(new_new_n9880__), .dout(new_new_n6465__));
  or1   g3367(.dina(new_new_n6465__), .dinb(new_new_n6464__), .dout(new_new_n6466__));
  and1  g3368(.dina(new_new_n9881__), .dinb(new_new_n9882__), .dout(new_new_n6467__));
  and1  g3369(.dina(new_new_n6467__), .dinb(new_new_n9884__), .dout(new_new_n6468__));
  and1  g3370(.dina(new_new_n4608__), .dinb(new_new_n4299__), .dout(new_new_n6469__));
  or1   g3371(.dina(new_new_n4609__), .dinb(new_new_n4298__), .dout(new_new_n6470__));
  and1  g3372(.dina(new_new_n4586__), .dinb(new_new_n4477__), .dout(new_new_n6471__));
  or1   g3373(.dina(new_new_n4587__), .dinb(new_new_n4476__), .dout(new_new_n6472__));
  and1  g3374(.dina(new_new_n6472__), .dinb(new_new_n6470__), .dout(new_new_n6473__));
  or1   g3375(.dina(new_new_n6471__), .dinb(new_new_n6469__), .dout(new_new_n6474__));
  and1  g3376(.dina(new_new_n9885__), .dinb(new_new_n9869__), .dout(new_new_n6475__));
  or1   g3377(.dina(new_new_n9886__), .dinb(new_new_n9877__), .dout(new_new_n6476__));
  and1  g3378(.dina(new_new_n9886__), .dinb(new_new_n9877__), .dout(new_new_n6477__));
  or1   g3379(.dina(new_new_n9885__), .dinb(new_new_n9869__), .dout(new_new_n6478__));
  and1  g3380(.dina(new_new_n6478__), .dinb(new_new_n6476__), .dout(new_new_n6479__));
  or1   g3381(.dina(new_new_n6477__), .dinb(new_new_n6475__), .dout(new_new_n6480__));
  and1  g3382(.dina(new_new_n6479__), .dinb(new_new_n9879__), .dout(new_new_n6481__));
  and1  g3383(.dina(new_new_n6480__), .dinb(new_new_n9880__), .dout(new_new_n6482__));
  or1   g3384(.dina(new_new_n6482__), .dinb(new_new_n6481__), .dout(new_new_n6483__));
  and1  g3385(.dina(new_new_n9887__), .dinb(new_new_n9889__), .dout(new_new_n6484__));
  and1  g3386(.dina(new_new_n6484__), .dinb(new_new_n9884__), .dout(new_new_n6485__));
  and1  g3387(.dina(new_new_n9882__), .dinb(new_new_n6206__), .dout(new_new_n6486__));
  or1   g3388(.dina(new_new_n9889__), .dinb(new_new_n9890__), .dout(new_new_n6487__));
  and1  g3389(.dina(new_new_n6486__), .dinb(new_new_n9881__), .dout(new_new_n6488__));
  and1  g3390(.dina(new_new_n6488__), .dinb(new_new_n9892__), .dout(new_new_n6489__));
  and1  g3391(.dina(new_new_n6487__), .dinb(new_new_n9887__), .dout(new_new_n6490__));
  and1  g3392(.dina(new_new_n6490__), .dinb(new_new_n9892__), .dout(new_new_n6491__));
  or1   g3393(.dina(new_new_n6485__), .dinb(new_new_n6468__), .dout(new_new_n6492__));
  or1   g3394(.dina(new_new_n6492__), .dinb(new_new_n6489__), .dout(new_new_n6493__));
  or1   g3395(.dina(new_new_n6493__), .dinb(new_new_n6491__), .dout(new_new_n6494__));
  and1  g3396(.dina(new_new_n4558__), .dinb(new_new_n4553__), .dout(new_new_n6495__));
  or1   g3397(.dina(new_new_n4559__), .dinb(new_new_n4552__), .dout(new_new_n6496__));
  and1  g3398(.dina(new_new_n9893__), .dinb(new_new_n9651__), .dout(new_new_n6497__));
  or1   g3399(.dina(new_new_n9894__), .dinb(new_new_n9645__), .dout(new_new_n6498__));
  and1  g3400(.dina(new_new_n9894__), .dinb(new_new_n9647__), .dout(new_new_n6499__));
  or1   g3401(.dina(new_new_n9893__), .dinb(new_new_n9653__), .dout(new_new_n6500__));
  and1  g3402(.dina(new_new_n6500__), .dinb(new_new_n6498__), .dout(new_new_n6501__));
  or1   g3403(.dina(new_new_n6499__), .dinb(new_new_n6497__), .dout(new_new_n6502__));
  or1   g3404(.dina(new_new_n6502__), .dinb(new_new_n9658__), .dout(new_new_n6503__));
  or1   g3405(.dina(new_new_n6501__), .dinb(new_new_n9663__), .dout(new_new_n6504__));
  and1  g3406(.dina(new_new_n6504__), .dinb(new_new_n6503__), .dout(new_new_n6505__));
  and1  g3407(.dina(new_new_n6505__), .dinb(new_new_n9883__), .dout(new_new_n6506__));
  and1  g3408(.dina(new_new_n4602__), .dinb(new_new_n4453__), .dout(new_new_n6507__));
  or1   g3409(.dina(new_new_n4603__), .dinb(new_new_n4452__), .dout(new_new_n6508__));
  and1  g3410(.dina(new_new_n4596__), .dinb(new_new_n4471__), .dout(new_new_n6509__));
  or1   g3411(.dina(new_new_n4597__), .dinb(new_new_n4470__), .dout(new_new_n6510__));
  and1  g3412(.dina(new_new_n6510__), .dinb(new_new_n6508__), .dout(new_new_n6511__));
  or1   g3413(.dina(new_new_n6509__), .dinb(new_new_n6507__), .dout(new_new_n6512__));
  and1  g3414(.dina(new_new_n9895__), .dinb(new_new_n9653__), .dout(new_new_n6513__));
  or1   g3415(.dina(new_new_n9896__), .dinb(new_new_n9647__), .dout(new_new_n6514__));
  and1  g3416(.dina(new_new_n9896__), .dinb(new_new_n9646__), .dout(new_new_n6515__));
  or1   g3417(.dina(new_new_n9895__), .dinb(new_new_n9652__), .dout(new_new_n6516__));
  and1  g3418(.dina(new_new_n6516__), .dinb(new_new_n6514__), .dout(new_new_n6517__));
  or1   g3419(.dina(new_new_n6515__), .dinb(new_new_n6513__), .dout(new_new_n6518__));
  and1  g3420(.dina(new_new_n6517__), .dinb(new_new_n9663__), .dout(new_new_n6519__));
  and1  g3421(.dina(new_new_n6518__), .dinb(new_new_n9658__), .dout(new_new_n6520__));
  or1   g3422(.dina(new_new_n6520__), .dinb(new_new_n6519__), .dout(new_new_n6521__));
  and1  g3423(.dina(new_new_n6521__), .dinb(new_new_n9891__), .dout(new_new_n6522__));
  or1   g3424(.dina(new_new_n6522__), .dinb(new_new_n6506__), .dout(new_new_n6523__));
  and1  g3425(.dina(new_new_n9722__), .dinb(new_new_n9898__), .dout(new_new_n6524__));
  and1  g3426(.dina(new_new_n9900__), .dinb(new_new_n9726__), .dout(new_new_n6525__));
  or1   g3427(.dina(new_new_n6525__), .dinb(new_new_n6524__), .dout(new_new_n6526__));
  and1  g3428(.dina(new_new_n9902__), .dinb(new_new_n9564__), .dout(new_new_n6527__));
  and1  g3429(.dina(new_new_n9903__), .dinb(new_new_n9553__), .dout(new_new_n6528__));
  or1   g3430(.dina(new_new_n6528__), .dinb(new_new_n6527__), .dout(new_new_n6529__));
  and1  g3431(.dina(new_new_n9905__), .dinb(new_new_n9747__), .dout(new_new_n6530__));
  and1  g3432(.dina(new_new_n9744__), .dinb(new_new_n9909__), .dout(new_new_n6531__));
  or1   g3433(.dina(new_new_n6531__), .dinb(new_new_n6530__), .dout(new_new_n6532__));
  and1  g3434(.dina(new_new_n9706__), .dinb(new_new_n9914__), .dout(new_new_n6533__));
  and1  g3435(.dina(new_new_n9712__), .dinb(new_new_n3386__), .dout(new_new_n6534__));
  or1   g3436(.dina(new_new_n6534__), .dinb(new_new_n6533__), .dout(new_new_n6535__));
  and1  g3437(.dina(new_new_n6293__), .dinb(new_new_n9917__), .dout(new_new_n6536__));
  and1  g3438(.dina(new_new_n9919__), .dinb(new_new_n3565__), .dout(new_new_n6537__));
  or1   g3439(.dina(new_new_n6537__), .dinb(new_new_n6536__), .dout(new_new_n6538__));
  and1  g3440(.dina(new_new_n6287__), .dinb(new_new_n9921__), .dout(new_new_n6539__));
  and1  g3441(.dina(new_new_n9923__), .dinb(new_new_n3593__), .dout(new_new_n6540__));
  or1   g3442(.dina(new_new_n6540__), .dinb(new_new_n6539__), .dout(new_new_n6541__));
  and1  g3443(.dina(new_new_n9817__), .dinb(new_new_n9924__), .dout(new_new_n6542__));
  or1   g3444(.dina(new_new_n9822__), .dinb(new_new_n3489__), .dout(new_new_n6543__));
  and1  g3445(.dina(new_new_n9824__), .dinb(new_new_n3492__), .dout(new_new_n6544__));
  or1   g3446(.dina(new_new_n9817__), .dinb(new_new_n3493__), .dout(new_new_n6545__));
  and1  g3447(.dina(new_new_n6545__), .dinb(new_new_n6543__), .dout(new_new_n6546__));
  or1   g3448(.dina(new_new_n6544__), .dinb(new_new_n6542__), .dout(new_new_n6547__));
  and1  g3449(.dina(new_new_n9828__), .dinb(new_new_n9925__), .dout(new_new_n6548__));
  or1   g3450(.dina(new_new_n9833__), .dinb(new_new_n3401__), .dout(new_new_n6549__));
  and1  g3451(.dina(new_new_n9835__), .dinb(new_new_n3404__), .dout(new_new_n6550__));
  or1   g3452(.dina(new_new_n9828__), .dinb(new_new_n3405__), .dout(new_new_n6551__));
  and1  g3453(.dina(new_new_n6551__), .dinb(new_new_n6549__), .dout(new_new_n6552__));
  or1   g3454(.dina(new_new_n6550__), .dinb(new_new_n6548__), .dout(new_new_n6553__));
  and1  g3455(.dina(new_new_n9927__), .dinb(new_new_n9931__), .dout(new_new_n6554__));
  and1  g3456(.dina(new_new_n9935__), .dinb(new_new_n9938__), .dout(new_new_n6555__));
  and1  g3457(.dina(new_new_n9941__), .dinb(new_new_n9945__), .dout(new_new_n6556__));
  and1  g3458(.dina(new_new_n9949__), .dinb(new_new_n9953__), .dout(new_new_n6557__));
  or1   g3459(.dina(new_new_n9723__), .dinb(new_new_n9727__), .dout(new_new_n6558__));
  or1   g3460(.dina(new_new_n9905__), .dinb(new_new_n9909__), .dout(new_new_n6559__));
  and1  g3461(.dina(new_new_n9957__), .dinb(new_new_n9960__), .dout(new_new_n6560__));
  and1  g3462(.dina(new_new_n9963__), .dinb(new_new_n9966__), .dout(new_new_n6561__));
  and1  g3463(.dina(new_new_n9970__), .dinb(new_new_n9973__), .dout(new_new_n6562__));
  and1  g3464(.dina(new_new_n9976__), .dinb(new_new_n3869__), .dout(new_new_n6563__));
  and1  g3465(.dina(new_new_n3871__), .dinb(new_new_n9977__), .dout(new_new_n6564__));
  and1  g3466(.dina(new_new_n9980__), .dinb(new_new_n9982__), .dout(new_new_n6565__));
  and1  g3467(.dina(new_new_n9985__), .dinb(new_new_n9988__), .dout(new_new_n6566__));
  and1  g3468(.dina(new_new_n9989__), .dinb(new_new_n3873__), .dout(new_new_n6567__));
  and1  g3469(.dina(new_new_n3877__), .dinb(new_new_n9990__), .dout(new_new_n6568__));
  and1  g3470(.dina(new_new_n9692__), .dinb(new_new_n9991__), .dout(new_new_n6569__));
  and1  g3471(.dina(new_new_n9696__), .dinb(new_new_n3525__), .dout(new_new_n6570__));
  and1  g3472(.dina(new_new_n9993__), .dinb(new_new_n9995__), .dout(new_new_n6571__));
  and1  g3473(.dina(new_new_n9997__), .dinb(new_new_n10000__), .dout(new_new_n6572__));
  and1  g3474(.dina(new_new_n10000__), .dinb(new_new_n10003__), .dout(new_new_n6573__));
  or1   g3475(.dina(new_new_n9997__), .dinb(new_new_n10003__), .dout(new_new_n6574__));
  or1   g3476(.dina(new_new_n10005__), .dinb(new_new_n10008__), .dout(new_new_n6575__));
  or1   g3477(.dina(new_new_n6319__), .dinb(new_new_n10013__), .dout(new_new_n6576__));
  and1  g3478(.dina(new_new_n10015__), .dinb(new_new_n10005__), .dout(new_new_n6577__));
  or1   g3479(.dina(new_new_n10015__), .dinb(new_new_n10008__), .dout(new_new_n6578__));
  and1  g3480(.dina(new_new_n9970__), .dinb(new_new_n10016__), .dout(new_new_n6579__));
  and1  g3481(.dina(new_new_n10017__), .dinb(new_new_n9963__), .dout(new_new_n6580__));
  and1  g3482(.dina(new_new_n3880__), .dinb(new_new_n9991__), .dout(new_new_n6581__));
  and1  g3483(.dina(new_new_n3857__), .dinb(new_new_n3530__), .dout(new_new_n6582__));
  or1   g3484(.dina(new_new_n6582__), .dinb(new_new_n6581__), .dout(new_new_n6583__));
  or1   g3485(.dina(new_new_n10018__), .dinb(new_new_n10020__), .dout(new_new_n6584__));
  and1  g3486(.dina(new_new_n9753__), .dinb(new_new_n9767__), .dout(new_new_n6585__));
  and1  g3487(.dina(new_new_n9673__), .dinb(new_new_n9900__), .dout(new_new_n6586__));
  and1  g3488(.dina(new_new_n9758__), .dinb(new_new_n9730__), .dout(new_new_n6587__));
  and1  g3489(.dina(new_new_n10022__), .dinb(new_new_n10024__), .dout(new_new_n6588__));
  and1  g3490(.dina(new_new_n10025__), .dinb(new_new_n4031__), .dout(new_new_n6589__));
  and1  g3491(.dina(new_new_n9679__), .dinb(new_new_n9723__), .dout(new_new_n6590__));
  and1  g3492(.dina(new_new_n10018__), .dinb(new_new_n10020__), .dout(new_new_n6591__));
  and1  g3493(.dina(new_new_n10026__), .dinb(new_new_n9993__), .dout(new_new_n6592__));
  and1  g3494(.dina(new_new_n10027__), .dinb(new_new_n9999__), .dout(new_new_n6593__));
  or1   g3495(.dina(new_new_n10028__), .dinb(new_new_n10029__), .dout(new_new_n6594__));
  or1   g3496(.dina(new_new_n6594__), .dinb(new_new_n10030__), .dout(new_new_n6595__));
  and1  g3497(.dina(new_new_n10031__), .dinb(new_new_n10009__), .dout(new_new_n6596__));
  and1  g3498(.dina(new_new_n6596__), .dinb(new_new_n10032__), .dout(new_new_n6597__));
  and1  g3499(.dina(new_new_n10033__), .dinb(new_new_n3929__), .dout(new_new_n6598__));
  and1  g3500(.dina(new_new_n4037__), .dinb(new_new_n10034__), .dout(new_new_n6599__));
  or1   g3501(.dina(new_new_n6599__), .dinb(new_new_n6598__), .dout(new_new_n6600__));
  and1  g3502(.dina(new_new_n9927__), .dinb(new_new_n10036__), .dout(new_new_n6601__));
  and1  g3503(.dina(new_new_n3919__), .dinb(new_new_n9931__), .dout(new_new_n6602__));
  or1   g3504(.dina(new_new_n6602__), .dinb(new_new_n6601__), .dout(new_new_n6603__));
  and1  g3505(.dina(new_new_n9935__), .dinb(new_new_n10038__), .dout(new_new_n6604__));
  and1  g3506(.dina(new_new_n3971__), .dinb(new_new_n9938__), .dout(new_new_n6605__));
  or1   g3507(.dina(new_new_n6605__), .dinb(new_new_n6604__), .dout(new_new_n6606__));
  and1  g3508(.dina(new_new_n9941__), .dinb(new_new_n10040__), .dout(new_new_n6607__));
  and1  g3509(.dina(new_new_n3909__), .dinb(new_new_n9945__), .dout(new_new_n6608__));
  or1   g3510(.dina(new_new_n6608__), .dinb(new_new_n6607__), .dout(new_new_n6609__));
  and1  g3511(.dina(new_new_n9949__), .dinb(new_new_n10043__), .dout(new_new_n6610__));
  and1  g3512(.dina(new_new_n3911__), .dinb(new_new_n9953__), .dout(new_new_n6611__));
  or1   g3513(.dina(new_new_n6611__), .dinb(new_new_n6610__), .dout(new_new_n6612__));
  and1  g3514(.dina(new_new_n9674__), .dinb(new_new_n9681__), .dout(new_new_n6613__));
  and1  g3515(.dina(new_new_n9678__), .dinb(new_new_n9676__), .dout(new_new_n6614__));
  or1   g3516(.dina(new_new_n6614__), .dinb(new_new_n6613__), .dout(new_new_n6615__));
  and1  g3517(.dina(new_new_n9683__), .dinb(new_new_n9691__), .dout(new_new_n6616__));
  and1  g3518(.dina(new_new_n9689__), .dinb(new_new_n9686__), .dout(new_new_n6617__));
  or1   g3519(.dina(new_new_n6617__), .dinb(new_new_n6616__), .dout(new_new_n6618__));
  and1  g3520(.dina(new_new_n9957__), .dinb(new_new_n10046__), .dout(new_new_n6619__));
  and1  g3521(.dina(new_new_n10047__), .dinb(new_new_n9960__), .dout(new_new_n6620__));
  or1   g3522(.dina(new_new_n6620__), .dinb(new_new_n6619__), .dout(new_new_n6621__));
  and1  g3523(.dina(new_new_n9962__), .dinb(new_new_n10049__), .dout(new_new_n6622__));
  and1  g3524(.dina(new_new_n10016__), .dinb(new_new_n9966__), .dout(new_new_n6623__));
  or1   g3525(.dina(new_new_n6623__), .dinb(new_new_n6622__), .dout(new_new_n6624__));
  and1  g3526(.dina(new_new_n9969__), .dinb(new_new_n10052__), .dout(new_new_n6625__));
  and1  g3527(.dina(new_new_n10017__), .dinb(new_new_n9973__), .dout(new_new_n6626__));
  or1   g3528(.dina(new_new_n6626__), .dinb(new_new_n6625__), .dout(new_new_n6627__));
  and1  g3529(.dina(new_new_n9684__), .dinb(new_new_n10047__), .dout(new_new_n6628__));
  and1  g3530(.dina(new_new_n9688__), .dinb(new_new_n9956__), .dout(new_new_n6629__));
  or1   g3531(.dina(new_new_n6629__), .dinb(new_new_n6628__), .dout(new_new_n6630__));
  and1  g3532(.dina(new_new_n3882__), .dinb(new_new_n9982__), .dout(new_new_n6631__));
  or1   g3533(.dina(new_new_n3883__), .dinb(new_new_n9988__), .dout(new_new_n6632__));
  and1  g3534(.dina(new_new_n3859__), .dinb(new_new_n3462__), .dout(new_new_n6633__));
  or1   g3535(.dina(new_new_n3858__), .dinb(new_new_n3463__), .dout(new_new_n6634__));
  and1  g3536(.dina(new_new_n6634__), .dinb(new_new_n6632__), .dout(new_new_n6635__));
  or1   g3537(.dina(new_new_n6633__), .dinb(new_new_n6631__), .dout(new_new_n6636__));
  or1   g3538(.dina(new_new_n6636__), .dinb(new_new_n9902__), .dout(new_new_n6637__));
  or1   g3539(.dina(new_new_n6635__), .dinb(new_new_n9903__), .dout(new_new_n6638__));
  and1  g3540(.dina(new_new_n6638__), .dinb(new_new_n6637__), .dout(new_new_n6639__));
  and1  g3541(.dina(new_new_n10056__), .dinb(new_new_n9727__), .dout(new_new_n6640__));
  or1   g3542(.dina(new_new_n10061__), .dinb(new_new_n9898__), .dout(new_new_n6641__));
  and1  g3543(.dina(new_new_n6640__), .dinb(new_new_n10065__), .dout(new_new_n6642__));
  or1   g3544(.dina(new_new_n6641__), .dinb(new_new_n10066__), .dout(new_new_n6643__));
  and1  g3545(.dina(new_new_n10069__), .dinb(new_new_n9729__), .dout(new_new_n6644__));
  or1   g3546(.dina(new_new_n10074__), .dinb(new_new_n9899__), .dout(new_new_n6645__));
  and1  g3547(.dina(new_new_n6644__), .dinb(new_new_n10066__), .dout(new_new_n6646__));
  or1   g3548(.dina(new_new_n6645__), .dinb(new_new_n10065__), .dout(new_new_n6647__));
  and1  g3549(.dina(new_new_n6647__), .dinb(new_new_n6643__), .dout(new_new_n6648__));
  or1   g3550(.dina(new_new_n6646__), .dinb(new_new_n6642__), .dout(new_new_n6649__));
  and1  g3551(.dina(new_new_n10080__), .dinb(new_new_n10085__), .dout(new_new_n6650__));
  or1   g3552(.dina(new_new_n10089__), .dinb(new_new_n10096__), .dout(new_new_n6651__));
  and1  g3553(.dina(new_new_n10100__), .dinb(new_new_n10096__), .dout(new_new_n6652__));
  or1   g3554(.dina(new_new_n10108__), .dinb(new_new_n10085__), .dout(new_new_n6653__));
  and1  g3555(.dina(new_new_n6653__), .dinb(new_new_n6651__), .dout(new_new_n6654__));
  or1   g3556(.dina(new_new_n6652__), .dinb(new_new_n6650__), .dout(new_new_n6655__));
  and1  g3557(.dina(new_new_n6654__), .dinb(new_new_n9899__), .dout(new_new_n6656__));
  or1   g3558(.dina(new_new_n6655__), .dinb(new_new_n9729__), .dout(new_new_n6657__));
  and1  g3559(.dina(new_new_n6657__), .dinb(new_new_n6648__), .dout(new_new_n6658__));
  or1   g3560(.dina(new_new_n6656__), .dinb(new_new_n6649__), .dout(new_new_n6659__));
  and1  g3561(.dina(new_new_n10056__), .dinb(new_new_n9735__), .dout(new_new_n6660__));
  or1   g3562(.dina(new_new_n10061__), .dinb(new_new_n9765__), .dout(new_new_n6661__));
  and1  g3563(.dina(new_new_n6660__), .dinb(new_new_n10113__), .dout(new_new_n6662__));
  or1   g3564(.dina(new_new_n6661__), .dinb(new_new_n10114__), .dout(new_new_n6663__));
  and1  g3565(.dina(new_new_n10069__), .dinb(new_new_n9735__), .dout(new_new_n6664__));
  or1   g3566(.dina(new_new_n10074__), .dinb(new_new_n9766__), .dout(new_new_n6665__));
  and1  g3567(.dina(new_new_n6664__), .dinb(new_new_n10114__), .dout(new_new_n6666__));
  or1   g3568(.dina(new_new_n6665__), .dinb(new_new_n10113__), .dout(new_new_n6667__));
  and1  g3569(.dina(new_new_n6667__), .dinb(new_new_n6663__), .dout(new_new_n6668__));
  or1   g3570(.dina(new_new_n6666__), .dinb(new_new_n6662__), .dout(new_new_n6669__));
  and1  g3571(.dina(new_new_n10080__), .dinb(new_new_n10115__), .dout(new_new_n6670__));
  or1   g3572(.dina(new_new_n10089__), .dinb(new_new_n10118__), .dout(new_new_n6671__));
  and1  g3573(.dina(new_new_n10100__), .dinb(new_new_n10118__), .dout(new_new_n6672__));
  or1   g3574(.dina(new_new_n10108__), .dinb(new_new_n10115__), .dout(new_new_n6673__));
  and1  g3575(.dina(new_new_n6673__), .dinb(new_new_n6671__), .dout(new_new_n6674__));
  or1   g3576(.dina(new_new_n6672__), .dinb(new_new_n6670__), .dout(new_new_n6675__));
  and1  g3577(.dina(new_new_n6674__), .dinb(new_new_n9766__), .dout(new_new_n6676__));
  or1   g3578(.dina(new_new_n6675__), .dinb(new_new_n9736__), .dout(new_new_n6677__));
  and1  g3579(.dina(new_new_n6677__), .dinb(new_new_n6668__), .dout(new_new_n6678__));
  or1   g3580(.dina(new_new_n6676__), .dinb(new_new_n6669__), .dout(new_new_n6679__));
  and1  g3581(.dina(new_new_n10120__), .dinb(new_new_n10121__), .dout(new_new_n6680__));
  or1   g3582(.dina(new_new_n10122__), .dinb(new_new_n10123__), .dout(new_new_n6681__));
  and1  g3583(.dina(new_new_n10122__), .dinb(new_new_n10123__), .dout(new_new_n6682__));
  or1   g3584(.dina(new_new_n10120__), .dinb(new_new_n10121__), .dout(new_new_n6683__));
  and1  g3585(.dina(new_new_n6683__), .dinb(new_new_n6681__), .dout(new_new_n6684__));
  or1   g3586(.dina(new_new_n6682__), .dinb(new_new_n6680__), .dout(new_new_n6685__));
  and1  g3587(.dina(new_new_n10057__), .dinb(new_new_n9762__), .dout(new_new_n6686__));
  or1   g3588(.dina(new_new_n10062__), .dinb(new_new_n9756__), .dout(new_new_n6687__));
  and1  g3589(.dina(new_new_n6686__), .dinb(new_new_n10124__), .dout(new_new_n6688__));
  or1   g3590(.dina(new_new_n6687__), .dinb(new_new_n10125__), .dout(new_new_n6689__));
  and1  g3591(.dina(new_new_n10070__), .dinb(new_new_n9762__), .dout(new_new_n6690__));
  or1   g3592(.dina(new_new_n10075__), .dinb(new_new_n9757__), .dout(new_new_n6691__));
  and1  g3593(.dina(new_new_n6690__), .dinb(new_new_n10125__), .dout(new_new_n6692__));
  or1   g3594(.dina(new_new_n6691__), .dinb(new_new_n10124__), .dout(new_new_n6693__));
  and1  g3595(.dina(new_new_n6693__), .dinb(new_new_n6689__), .dout(new_new_n6694__));
  or1   g3596(.dina(new_new_n6692__), .dinb(new_new_n6688__), .dout(new_new_n6695__));
  and1  g3597(.dina(new_new_n10081__), .dinb(new_new_n10126__), .dout(new_new_n6696__));
  or1   g3598(.dina(new_new_n10088__), .dinb(new_new_n10129__), .dout(new_new_n6697__));
  and1  g3599(.dina(new_new_n10101__), .dinb(new_new_n10129__), .dout(new_new_n6698__));
  or1   g3600(.dina(new_new_n10107__), .dinb(new_new_n10126__), .dout(new_new_n6699__));
  and1  g3601(.dina(new_new_n6699__), .dinb(new_new_n6697__), .dout(new_new_n6700__));
  or1   g3602(.dina(new_new_n6698__), .dinb(new_new_n6696__), .dout(new_new_n6701__));
  and1  g3603(.dina(new_new_n6700__), .dinb(new_new_n9757__), .dout(new_new_n6702__));
  or1   g3604(.dina(new_new_n6701__), .dinb(new_new_n9763__), .dout(new_new_n6703__));
  and1  g3605(.dina(new_new_n6703__), .dinb(new_new_n6694__), .dout(new_new_n6704__));
  or1   g3606(.dina(new_new_n6702__), .dinb(new_new_n6695__), .dout(new_new_n6705__));
  and1  g3607(.dina(new_new_n10131__), .dinb(new_new_n10132__), .dout(new_new_n6706__));
  or1   g3608(.dina(new_new_n10133__), .dinb(new_new_n10135__), .dout(new_new_n6707__));
  and1  g3609(.dina(new_new_n10133__), .dinb(new_new_n10135__), .dout(new_new_n6708__));
  or1   g3610(.dina(new_new_n10131__), .dinb(new_new_n10132__), .dout(new_new_n6709__));
  and1  g3611(.dina(new_new_n6709__), .dinb(new_new_n6707__), .dout(new_new_n6710__));
  or1   g3612(.dina(new_new_n6708__), .dinb(new_new_n6706__), .dout(new_new_n6711__));
  or1   g3613(.dina(new_new_n6711__), .dinb(new_new_n6684__), .dout(new_new_n6712__));
  or1   g3614(.dina(new_new_n6710__), .dinb(new_new_n6685__), .dout(new_new_n6713__));
  and1  g3615(.dina(new_new_n6713__), .dinb(new_new_n6712__), .dout(new_new_n6714__));
  and1  g3616(.dina(new_new_n9546__), .dinb(new_new_n9910__), .dout(new_new_n6715__));
  or1   g3617(.dina(new_new_n9556__), .dinb(new_new_n9746__), .dout(new_new_n6716__));
  and1  g3618(.dina(new_new_n6715__), .dinb(new_new_n10136__), .dout(new_new_n6717__));
  or1   g3619(.dina(new_new_n6716__), .dinb(new_new_n10137__), .dout(new_new_n6718__));
  and1  g3620(.dina(new_new_n9568__), .dinb(new_new_n9910__), .dout(new_new_n6719__));
  or1   g3621(.dina(new_new_n9574__), .dinb(new_new_n9748__), .dout(new_new_n6720__));
  and1  g3622(.dina(new_new_n6719__), .dinb(new_new_n10137__), .dout(new_new_n6721__));
  or1   g3623(.dina(new_new_n6720__), .dinb(new_new_n10136__), .dout(new_new_n6722__));
  and1  g3624(.dina(new_new_n6722__), .dinb(new_new_n6718__), .dout(new_new_n6723__));
  or1   g3625(.dina(new_new_n6721__), .dinb(new_new_n6717__), .dout(new_new_n6724__));
  and1  g3626(.dina(new_new_n9580__), .dinb(new_new_n10138__), .dout(new_new_n6725__));
  or1   g3627(.dina(new_new_n9589__), .dinb(new_new_n10141__), .dout(new_new_n6726__));
  and1  g3628(.dina(new_new_n9597__), .dinb(new_new_n10141__), .dout(new_new_n6727__));
  or1   g3629(.dina(new_new_n9603__), .dinb(new_new_n10138__), .dout(new_new_n6728__));
  and1  g3630(.dina(new_new_n6728__), .dinb(new_new_n6726__), .dout(new_new_n6729__));
  or1   g3631(.dina(new_new_n6727__), .dinb(new_new_n6725__), .dout(new_new_n6730__));
  and1  g3632(.dina(new_new_n6729__), .dinb(new_new_n9748__), .dout(new_new_n6731__));
  or1   g3633(.dina(new_new_n6730__), .dinb(new_new_n9911__), .dout(new_new_n6732__));
  and1  g3634(.dina(new_new_n6732__), .dinb(new_new_n6723__), .dout(new_new_n6733__));
  or1   g3635(.dina(new_new_n6731__), .dinb(new_new_n6724__), .dout(new_new_n6734__));
  and1  g3636(.dina(new_new_n9546__), .dinb(new_new_n9774__), .dout(new_new_n6735__));
  or1   g3637(.dina(new_new_n9558__), .dinb(new_new_n9742__), .dout(new_new_n6736__));
  and1  g3638(.dina(new_new_n6735__), .dinb(new_new_n10143__), .dout(new_new_n6737__));
  or1   g3639(.dina(new_new_n6736__), .dinb(new_new_n10144__), .dout(new_new_n6738__));
  and1  g3640(.dina(new_new_n9568__), .dinb(new_new_n9774__), .dout(new_new_n6739__));
  or1   g3641(.dina(new_new_n9574__), .dinb(new_new_n9743__), .dout(new_new_n6740__));
  and1  g3642(.dina(new_new_n6739__), .dinb(new_new_n10144__), .dout(new_new_n6741__));
  or1   g3643(.dina(new_new_n6740__), .dinb(new_new_n10143__), .dout(new_new_n6742__));
  and1  g3644(.dina(new_new_n6742__), .dinb(new_new_n6738__), .dout(new_new_n6743__));
  or1   g3645(.dina(new_new_n6741__), .dinb(new_new_n6737__), .dout(new_new_n6744__));
  and1  g3646(.dina(new_new_n9581__), .dinb(new_new_n10145__), .dout(new_new_n6745__));
  or1   g3647(.dina(new_new_n9588__), .dinb(new_new_n10148__), .dout(new_new_n6746__));
  and1  g3648(.dina(new_new_n9598__), .dinb(new_new_n10148__), .dout(new_new_n6747__));
  or1   g3649(.dina(new_new_n9604__), .dinb(new_new_n10145__), .dout(new_new_n6748__));
  and1  g3650(.dina(new_new_n6748__), .dinb(new_new_n6746__), .dout(new_new_n6749__));
  or1   g3651(.dina(new_new_n6747__), .dinb(new_new_n6745__), .dout(new_new_n6750__));
  and1  g3652(.dina(new_new_n6749__), .dinb(new_new_n9743__), .dout(new_new_n6751__));
  or1   g3653(.dina(new_new_n6750__), .dinb(new_new_n9775__), .dout(new_new_n6752__));
  and1  g3654(.dina(new_new_n6752__), .dinb(new_new_n6743__), .dout(new_new_n6753__));
  or1   g3655(.dina(new_new_n6751__), .dinb(new_new_n6744__), .dout(new_new_n6754__));
  and1  g3656(.dina(new_new_n10150__), .dinb(new_new_n10151__), .dout(new_new_n6755__));
  or1   g3657(.dina(new_new_n10152__), .dinb(new_new_n10153__), .dout(new_new_n6756__));
  and1  g3658(.dina(new_new_n10152__), .dinb(new_new_n10153__), .dout(new_new_n6757__));
  or1   g3659(.dina(new_new_n10150__), .dinb(new_new_n10151__), .dout(new_new_n6758__));
  and1  g3660(.dina(new_new_n6758__), .dinb(new_new_n6756__), .dout(new_new_n6759__));
  or1   g3661(.dina(new_new_n6757__), .dinb(new_new_n6755__), .dout(new_new_n6760__));
  and1  g3662(.dina(new_new_n9548__), .dinb(new_new_n10154__), .dout(new_new_n6761__));
  or1   g3663(.dina(new_new_n9558__), .dinb(new_new_n10157__), .dout(new_new_n6762__));
  and1  g3664(.dina(new_new_n9570__), .dinb(new_new_n10157__), .dout(new_new_n6763__));
  or1   g3665(.dina(new_new_n9576__), .dinb(new_new_n10154__), .dout(new_new_n6764__));
  and1  g3666(.dina(new_new_n6764__), .dinb(new_new_n6762__), .dout(new_new_n6765__));
  or1   g3667(.dina(new_new_n6763__), .dinb(new_new_n6761__), .dout(new_new_n6766__));
  and1  g3668(.dina(new_new_n9581__), .dinb(new_new_n10159__), .dout(new_new_n6767__));
  or1   g3669(.dina(new_new_n9590__), .dinb(new_new_n10162__), .dout(new_new_n6768__));
  and1  g3670(.dina(new_new_n9598__), .dinb(new_new_n10162__), .dout(new_new_n6769__));
  or1   g3671(.dina(new_new_n9604__), .dinb(new_new_n10159__), .dout(new_new_n6770__));
  and1  g3672(.dina(new_new_n6770__), .dinb(new_new_n6768__), .dout(new_new_n6771__));
  or1   g3673(.dina(new_new_n6769__), .dinb(new_new_n6767__), .dout(new_new_n6772__));
  and1  g3674(.dina(new_new_n10164__), .dinb(new_new_n10165__), .dout(new_new_n6773__));
  or1   g3675(.dina(new_new_n10166__), .dinb(new_new_n10167__), .dout(new_new_n6774__));
  and1  g3676(.dina(new_new_n10166__), .dinb(new_new_n10167__), .dout(new_new_n6775__));
  or1   g3677(.dina(new_new_n10164__), .dinb(new_new_n10165__), .dout(new_new_n6776__));
  and1  g3678(.dina(new_new_n6776__), .dinb(new_new_n6774__), .dout(new_new_n6777__));
  or1   g3679(.dina(new_new_n6775__), .dinb(new_new_n6773__), .dout(new_new_n6778__));
  or1   g3680(.dina(new_new_n6778__), .dinb(new_new_n6759__), .dout(new_new_n6779__));
  or1   g3681(.dina(new_new_n6777__), .dinb(new_new_n6760__), .dout(new_new_n6780__));
  and1  g3682(.dina(new_new_n6780__), .dinb(new_new_n6779__), .dout(new_new_n6781__));
  and1  g3683(.dina(new_new_n10057__), .dinb(new_new_n9932__), .dout(new_new_n6782__));
  or1   g3684(.dina(new_new_n10062__), .dinb(new_new_n10036__), .dout(new_new_n6783__));
  and1  g3685(.dina(new_new_n6782__), .dinb(new_new_n9980__), .dout(new_new_n6784__));
  or1   g3686(.dina(new_new_n6783__), .dinb(new_new_n9985__), .dout(new_new_n6785__));
  and1  g3687(.dina(new_new_n10070__), .dinb(new_new_n9932__), .dout(new_new_n6786__));
  or1   g3688(.dina(new_new_n10075__), .dinb(new_new_n10037__), .dout(new_new_n6787__));
  and1  g3689(.dina(new_new_n6786__), .dinb(new_new_n9986__), .dout(new_new_n6788__));
  or1   g3690(.dina(new_new_n6787__), .dinb(new_new_n9979__), .dout(new_new_n6789__));
  and1  g3691(.dina(new_new_n6789__), .dinb(new_new_n6785__), .dout(new_new_n6790__));
  or1   g3692(.dina(new_new_n6788__), .dinb(new_new_n6784__), .dout(new_new_n6791__));
  and1  g3693(.dina(new_new_n10081__), .dinb(new_new_n9981__), .dout(new_new_n6792__));
  or1   g3694(.dina(new_new_n10090__), .dinb(new_new_n9986__), .dout(new_new_n6793__));
  and1  g3695(.dina(new_new_n10101__), .dinb(new_new_n9987__), .dout(new_new_n6794__));
  or1   g3696(.dina(new_new_n10109__), .dinb(new_new_n9981__), .dout(new_new_n6795__));
  and1  g3697(.dina(new_new_n6795__), .dinb(new_new_n6793__), .dout(new_new_n6796__));
  or1   g3698(.dina(new_new_n6794__), .dinb(new_new_n6792__), .dout(new_new_n6797__));
  and1  g3699(.dina(new_new_n6796__), .dinb(new_new_n10037__), .dout(new_new_n6798__));
  or1   g3700(.dina(new_new_n6797__), .dinb(new_new_n9933__), .dout(new_new_n6799__));
  and1  g3701(.dina(new_new_n6799__), .dinb(new_new_n6790__), .dout(new_new_n6800__));
  or1   g3702(.dina(new_new_n6798__), .dinb(new_new_n6791__), .dout(new_new_n6801__));
  and1  g3703(.dina(new_new_n10058__), .dinb(new_new_n9954__), .dout(new_new_n6802__));
  or1   g3704(.dina(new_new_n10064__), .dinb(new_new_n10043__), .dout(new_new_n6803__));
  and1  g3705(.dina(new_new_n6802__), .dinb(new_new_n4287__), .dout(new_new_n6804__));
  or1   g3706(.dina(new_new_n6803__), .dinb(new_new_n4286__), .dout(new_new_n6805__));
  and1  g3707(.dina(new_new_n10071__), .dinb(new_new_n9954__), .dout(new_new_n6806__));
  or1   g3708(.dina(new_new_n10077__), .dinb(new_new_n10044__), .dout(new_new_n6807__));
  and1  g3709(.dina(new_new_n6806__), .dinb(new_new_n4572__), .dout(new_new_n6808__));
  or1   g3710(.dina(new_new_n6807__), .dinb(new_new_n4573__), .dout(new_new_n6809__));
  and1  g3711(.dina(new_new_n6809__), .dinb(new_new_n6805__), .dout(new_new_n6810__));
  or1   g3712(.dina(new_new_n6808__), .dinb(new_new_n6804__), .dout(new_new_n6811__));
  and1  g3713(.dina(new_new_n10083__), .dinb(new_new_n10168__), .dout(new_new_n6812__));
  or1   g3714(.dina(new_new_n10090__), .dinb(new_new_n10169__), .dout(new_new_n6813__));
  and1  g3715(.dina(new_new_n10103__), .dinb(new_new_n10169__), .dout(new_new_n6814__));
  or1   g3716(.dina(new_new_n10109__), .dinb(new_new_n10168__), .dout(new_new_n6815__));
  and1  g3717(.dina(new_new_n6815__), .dinb(new_new_n6813__), .dout(new_new_n6816__));
  or1   g3718(.dina(new_new_n6814__), .dinb(new_new_n6812__), .dout(new_new_n6817__));
  and1  g3719(.dina(new_new_n6816__), .dinb(new_new_n10044__), .dout(new_new_n6818__));
  or1   g3720(.dina(new_new_n6817__), .dinb(new_new_n9955__), .dout(new_new_n6819__));
  and1  g3721(.dina(new_new_n6819__), .dinb(new_new_n6810__), .dout(new_new_n6820__));
  or1   g3722(.dina(new_new_n6818__), .dinb(new_new_n6811__), .dout(new_new_n6821__));
  and1  g3723(.dina(new_new_n10058__), .dinb(new_new_n9946__), .dout(new_new_n6822__));
  or1   g3724(.dina(new_new_n10064__), .dinb(new_new_n10040__), .dout(new_new_n6823__));
  and1  g3725(.dina(new_new_n6822__), .dinb(new_new_n4285__), .dout(new_new_n6824__));
  or1   g3726(.dina(new_new_n6823__), .dinb(new_new_n4284__), .dout(new_new_n6825__));
  and1  g3727(.dina(new_new_n10071__), .dinb(new_new_n9946__), .dout(new_new_n6826__));
  or1   g3728(.dina(new_new_n10077__), .dinb(new_new_n10041__), .dout(new_new_n6827__));
  and1  g3729(.dina(new_new_n6826__), .dinb(new_new_n4570__), .dout(new_new_n6828__));
  or1   g3730(.dina(new_new_n6827__), .dinb(new_new_n4571__), .dout(new_new_n6829__));
  and1  g3731(.dina(new_new_n6829__), .dinb(new_new_n6825__), .dout(new_new_n6830__));
  or1   g3732(.dina(new_new_n6828__), .dinb(new_new_n6824__), .dout(new_new_n6831__));
  and1  g3733(.dina(new_new_n10083__), .dinb(new_new_n10170__), .dout(new_new_n6832__));
  or1   g3734(.dina(new_new_n10092__), .dinb(new_new_n10171__), .dout(new_new_n6833__));
  and1  g3735(.dina(new_new_n10103__), .dinb(new_new_n10171__), .dout(new_new_n6834__));
  or1   g3736(.dina(new_new_n10111__), .dinb(new_new_n10170__), .dout(new_new_n6835__));
  and1  g3737(.dina(new_new_n6835__), .dinb(new_new_n6833__), .dout(new_new_n6836__));
  or1   g3738(.dina(new_new_n6834__), .dinb(new_new_n6832__), .dout(new_new_n6837__));
  and1  g3739(.dina(new_new_n6836__), .dinb(new_new_n10041__), .dout(new_new_n6838__));
  or1   g3740(.dina(new_new_n6837__), .dinb(new_new_n9947__), .dout(new_new_n6839__));
  and1  g3741(.dina(new_new_n6839__), .dinb(new_new_n6830__), .dout(new_new_n6840__));
  or1   g3742(.dina(new_new_n6838__), .dinb(new_new_n6831__), .dout(new_new_n6841__));
  and1  g3743(.dina(new_new_n10172__), .dinb(new_new_n10173__), .dout(new_new_n6842__));
  or1   g3744(.dina(new_new_n10174__), .dinb(new_new_n10175__), .dout(new_new_n6843__));
  and1  g3745(.dina(new_new_n10174__), .dinb(new_new_n10175__), .dout(new_new_n6844__));
  or1   g3746(.dina(new_new_n10172__), .dinb(new_new_n10173__), .dout(new_new_n6845__));
  and1  g3747(.dina(new_new_n6845__), .dinb(new_new_n6843__), .dout(new_new_n6846__));
  or1   g3748(.dina(new_new_n6844__), .dinb(new_new_n6842__), .dout(new_new_n6847__));
  and1  g3749(.dina(new_new_n4527__), .dinb(new_new_n4525__), .dout(new_new_n6848__));
  or1   g3750(.dina(new_new_n4526__), .dinb(new_new_n4524__), .dout(new_new_n6849__));
  and1  g3751(.dina(new_new_n10084__), .dinb(new_new_n4293__), .dout(new_new_n6850__));
  or1   g3752(.dina(new_new_n10092__), .dinb(new_new_n4292__), .dout(new_new_n6851__));
  and1  g3753(.dina(new_new_n4580__), .dinb(new_new_n10104__), .dout(new_new_n6852__));
  or1   g3754(.dina(new_new_n4581__), .dinb(new_new_n10111__), .dout(new_new_n6853__));
  and1  g3755(.dina(new_new_n6853__), .dinb(new_new_n6851__), .dout(new_new_n6854__));
  or1   g3756(.dina(new_new_n6852__), .dinb(new_new_n6850__), .dout(new_new_n6855__));
  and1  g3757(.dina(new_new_n6854__), .dinb(new_new_n10038__), .dout(new_new_n6856__));
  or1   g3758(.dina(new_new_n6855__), .dinb(new_new_n9939__), .dout(new_new_n6857__));
  and1  g3759(.dina(new_new_n6857__), .dinb(new_new_n6848__), .dout(new_new_n6858__));
  or1   g3760(.dina(new_new_n6856__), .dinb(new_new_n6849__), .dout(new_new_n6859__));
  and1  g3761(.dina(new_new_n4533__), .dinb(new_new_n4531__), .dout(new_new_n6860__));
  or1   g3762(.dina(new_new_n4532__), .dinb(new_new_n4530__), .dout(new_new_n6861__));
  and1  g3763(.dina(new_new_n10084__), .dinb(new_new_n4303__), .dout(new_new_n6862__));
  or1   g3764(.dina(new_new_n10093__), .dinb(new_new_n4302__), .dout(new_new_n6863__));
  and1  g3765(.dina(new_new_n4590__), .dinb(new_new_n10104__), .dout(new_new_n6864__));
  or1   g3766(.dina(new_new_n4591__), .dinb(new_new_n10112__), .dout(new_new_n6865__));
  and1  g3767(.dina(new_new_n6865__), .dinb(new_new_n6863__), .dout(new_new_n6866__));
  or1   g3768(.dina(new_new_n6864__), .dinb(new_new_n6862__), .dout(new_new_n6867__));
  and1  g3769(.dina(new_new_n6866__), .dinb(new_new_n9680__), .dout(new_new_n6868__));
  or1   g3770(.dina(new_new_n6867__), .dinb(new_new_n9677__), .dout(new_new_n6869__));
  and1  g3771(.dina(new_new_n6869__), .dinb(new_new_n6860__), .dout(new_new_n6870__));
  or1   g3772(.dina(new_new_n6868__), .dinb(new_new_n6861__), .dout(new_new_n6871__));
  and1  g3773(.dina(new_new_n10176__), .dinb(new_new_n10177__), .dout(new_new_n6872__));
  or1   g3774(.dina(new_new_n10178__), .dinb(new_new_n10179__), .dout(new_new_n6873__));
  and1  g3775(.dina(new_new_n10178__), .dinb(new_new_n10179__), .dout(new_new_n6874__));
  or1   g3776(.dina(new_new_n10176__), .dinb(new_new_n10177__), .dout(new_new_n6875__));
  and1  g3777(.dina(new_new_n6875__), .dinb(new_new_n6873__), .dout(new_new_n6876__));
  or1   g3778(.dina(new_new_n6874__), .dinb(new_new_n6872__), .dout(new_new_n6877__));
  or1   g3779(.dina(new_new_n10180__), .dinb(new_new_n10181__), .dout(new_new_n6878__));
  or1   g3780(.dina(new_new_n6878__), .dinb(new_new_n10182__), .dout(new_new_n6879__));
  or1   g3781(.dina(new_new_n10180__), .dinb(new_new_n10183__), .dout(new_new_n6880__));
  or1   g3782(.dina(new_new_n6880__), .dinb(new_new_n10184__), .dout(new_new_n6881__));
  and1  g3783(.dina(new_new_n6881__), .dinb(new_new_n6879__), .dout(new_new_n6882__));
  or1   g3784(.dina(new_new_n10185__), .dinb(new_new_n10183__), .dout(new_new_n6883__));
  or1   g3785(.dina(new_new_n6883__), .dinb(new_new_n10182__), .dout(new_new_n6884__));
  or1   g3786(.dina(new_new_n10185__), .dinb(new_new_n10181__), .dout(new_new_n6885__));
  or1   g3787(.dina(new_new_n6885__), .dinb(new_new_n10184__), .dout(new_new_n6886__));
  and1  g3788(.dina(new_new_n6886__), .dinb(new_new_n6884__), .dout(new_new_n6887__));
  and1  g3789(.dina(new_new_n6887__), .dinb(new_new_n6882__), .dout(new_new_n6888__));
  and1  g3790(.dina(new_new_n9548__), .dinb(new_new_n9974__), .dout(new_new_n6889__));
  or1   g3791(.dina(new_new_n9560__), .dinb(new_new_n10052__), .dout(new_new_n6890__));
  and1  g3792(.dina(new_new_n6889__), .dinb(new_new_n4291__), .dout(new_new_n6891__));
  or1   g3793(.dina(new_new_n6890__), .dinb(new_new_n4290__), .dout(new_new_n6892__));
  and1  g3794(.dina(new_new_n9570__), .dinb(new_new_n9974__), .dout(new_new_n6893__));
  or1   g3795(.dina(new_new_n9576__), .dinb(new_new_n10053__), .dout(new_new_n6894__));
  and1  g3796(.dina(new_new_n6893__), .dinb(new_new_n4576__), .dout(new_new_n6895__));
  or1   g3797(.dina(new_new_n6894__), .dinb(new_new_n4577__), .dout(new_new_n6896__));
  and1  g3798(.dina(new_new_n6896__), .dinb(new_new_n6892__), .dout(new_new_n6897__));
  or1   g3799(.dina(new_new_n6895__), .dinb(new_new_n6891__), .dout(new_new_n6898__));
  and1  g3800(.dina(new_new_n9583__), .dinb(new_new_n10186__), .dout(new_new_n6899__));
  or1   g3801(.dina(new_new_n9590__), .dinb(new_new_n10187__), .dout(new_new_n6900__));
  and1  g3802(.dina(new_new_n9600__), .dinb(new_new_n10187__), .dout(new_new_n6901__));
  or1   g3803(.dina(new_new_n9606__), .dinb(new_new_n10186__), .dout(new_new_n6902__));
  and1  g3804(.dina(new_new_n6902__), .dinb(new_new_n6900__), .dout(new_new_n6903__));
  or1   g3805(.dina(new_new_n6901__), .dinb(new_new_n6899__), .dout(new_new_n6904__));
  and1  g3806(.dina(new_new_n6903__), .dinb(new_new_n10053__), .dout(new_new_n6905__));
  or1   g3807(.dina(new_new_n6904__), .dinb(new_new_n9975__), .dout(new_new_n6906__));
  and1  g3808(.dina(new_new_n6906__), .dinb(new_new_n6897__), .dout(new_new_n6907__));
  or1   g3809(.dina(new_new_n6905__), .dinb(new_new_n6898__), .dout(new_new_n6908__));
  and1  g3810(.dina(new_new_n9549__), .dinb(new_new_n9967__), .dout(new_new_n6909__));
  or1   g3811(.dina(new_new_n9560__), .dinb(new_new_n10049__), .dout(new_new_n6910__));
  and1  g3812(.dina(new_new_n6909__), .dinb(new_new_n4289__), .dout(new_new_n6911__));
  or1   g3813(.dina(new_new_n6910__), .dinb(new_new_n4288__), .dout(new_new_n6912__));
  and1  g3814(.dina(new_new_n9569__), .dinb(new_new_n9967__), .dout(new_new_n6913__));
  or1   g3815(.dina(new_new_n9577__), .dinb(new_new_n10050__), .dout(new_new_n6914__));
  and1  g3816(.dina(new_new_n6913__), .dinb(new_new_n4574__), .dout(new_new_n6915__));
  or1   g3817(.dina(new_new_n6914__), .dinb(new_new_n4575__), .dout(new_new_n6916__));
  and1  g3818(.dina(new_new_n6916__), .dinb(new_new_n6912__), .dout(new_new_n6917__));
  or1   g3819(.dina(new_new_n6915__), .dinb(new_new_n6911__), .dout(new_new_n6918__));
  and1  g3820(.dina(new_new_n9583__), .dinb(new_new_n10188__), .dout(new_new_n6919__));
  or1   g3821(.dina(new_new_n9592__), .dinb(new_new_n10189__), .dout(new_new_n6920__));
  and1  g3822(.dina(new_new_n9600__), .dinb(new_new_n10189__), .dout(new_new_n6921__));
  or1   g3823(.dina(new_new_n9606__), .dinb(new_new_n10188__), .dout(new_new_n6922__));
  and1  g3824(.dina(new_new_n6922__), .dinb(new_new_n6920__), .dout(new_new_n6923__));
  or1   g3825(.dina(new_new_n6921__), .dinb(new_new_n6919__), .dout(new_new_n6924__));
  and1  g3826(.dina(new_new_n6923__), .dinb(new_new_n10050__), .dout(new_new_n6925__));
  or1   g3827(.dina(new_new_n6924__), .dinb(new_new_n9968__), .dout(new_new_n6926__));
  and1  g3828(.dina(new_new_n6926__), .dinb(new_new_n6917__), .dout(new_new_n6927__));
  or1   g3829(.dina(new_new_n6925__), .dinb(new_new_n6918__), .dout(new_new_n6928__));
  and1  g3830(.dina(new_new_n10190__), .dinb(new_new_n10191__), .dout(new_new_n6929__));
  or1   g3831(.dina(new_new_n10192__), .dinb(new_new_n10193__), .dout(new_new_n6930__));
  and1  g3832(.dina(new_new_n10192__), .dinb(new_new_n10193__), .dout(new_new_n6931__));
  or1   g3833(.dina(new_new_n10190__), .dinb(new_new_n10191__), .dout(new_new_n6932__));
  and1  g3834(.dina(new_new_n6932__), .dinb(new_new_n6930__), .dout(new_new_n6933__));
  or1   g3835(.dina(new_new_n6931__), .dinb(new_new_n6929__), .dout(new_new_n6934__));
  and1  g3836(.dina(new_new_n9549__), .dinb(new_new_n9959__), .dout(new_new_n6935__));
  or1   g3837(.dina(new_new_n9561__), .dinb(new_new_n10046__), .dout(new_new_n6936__));
  and1  g3838(.dina(new_new_n9592__), .dinb(new_new_n10045__), .dout(new_new_n6937__));
  or1   g3839(.dina(new_new_n9584__), .dinb(new_new_n9961__), .dout(new_new_n6938__));
  and1  g3840(.dina(new_new_n6938__), .dinb(new_new_n6936__), .dout(new_new_n6939__));
  or1   g3841(.dina(new_new_n6937__), .dinb(new_new_n6935__), .dout(new_new_n6940__));
  and1  g3842(.dina(new_new_n4537__), .dinb(new_new_n4535__), .dout(new_new_n6941__));
  or1   g3843(.dina(new_new_n4536__), .dinb(new_new_n4534__), .dout(new_new_n6942__));
  and1  g3844(.dina(new_new_n9584__), .dinb(new_new_n4305__), .dout(new_new_n6943__));
  or1   g3845(.dina(new_new_n9593__), .dinb(new_new_n4304__), .dout(new_new_n6944__));
  and1  g3846(.dina(new_new_n4592__), .dinb(new_new_n9599__), .dout(new_new_n6945__));
  or1   g3847(.dina(new_new_n4593__), .dinb(new_new_n9607__), .dout(new_new_n6946__));
  and1  g3848(.dina(new_new_n6946__), .dinb(new_new_n6944__), .dout(new_new_n6947__));
  or1   g3849(.dina(new_new_n6945__), .dinb(new_new_n6943__), .dout(new_new_n6948__));
  and1  g3850(.dina(new_new_n6947__), .dinb(new_new_n9690__), .dout(new_new_n6949__));
  or1   g3851(.dina(new_new_n6948__), .dinb(new_new_n9687__), .dout(new_new_n6950__));
  and1  g3852(.dina(new_new_n6950__), .dinb(new_new_n6941__), .dout(new_new_n6951__));
  or1   g3853(.dina(new_new_n6949__), .dinb(new_new_n6942__), .dout(new_new_n6952__));
  and1  g3854(.dina(new_new_n10194__), .dinb(new_new_n10195__), .dout(new_new_n6953__));
  or1   g3855(.dina(new_new_n10196__), .dinb(new_new_n10197__), .dout(new_new_n6954__));
  and1  g3856(.dina(new_new_n10196__), .dinb(new_new_n10197__), .dout(new_new_n6955__));
  or1   g3857(.dina(new_new_n10194__), .dinb(new_new_n10195__), .dout(new_new_n6956__));
  and1  g3858(.dina(new_new_n6956__), .dinb(new_new_n6954__), .dout(new_new_n6957__));
  or1   g3859(.dina(new_new_n6955__), .dinb(new_new_n6953__), .dout(new_new_n6958__));
  and1  g3860(.dina(new_new_n10198__), .dinb(new_new_n10199__), .dout(new_new_n6959__));
  and1  g3861(.dina(new_new_n6959__), .dinb(new_new_n10200__), .dout(new_new_n6960__));
  and1  g3862(.dina(new_new_n10198__), .dinb(new_new_n10202__), .dout(new_new_n6961__));
  and1  g3863(.dina(new_new_n6961__), .dinb(new_new_n10203__), .dout(new_new_n6962__));
  or1   g3864(.dina(new_new_n6962__), .dinb(new_new_n6960__), .dout(new_new_n6963__));
  and1  g3865(.dina(new_new_n10204__), .dinb(new_new_n10202__), .dout(new_new_n6964__));
  and1  g3866(.dina(new_new_n6964__), .dinb(new_new_n10200__), .dout(new_new_n6965__));
  and1  g3867(.dina(new_new_n10204__), .dinb(new_new_n10199__), .dout(new_new_n6966__));
  and1  g3868(.dina(new_new_n6966__), .dinb(new_new_n10203__), .dout(new_new_n6967__));
  or1   g3869(.dina(new_new_n6967__), .dinb(new_new_n6965__), .dout(new_new_n6968__));
  or1   g3870(.dina(new_new_n6968__), .dinb(new_new_n6963__), .dout(new_new_n6969__));
  and1  g3871(.dina(new_new_n10206__), .dinb(new_new_n10208__), .dout(new_new_n6970__));
  and1  g3872(.dina(new_new_n10210__), .dinb(new_new_n10212__), .dout(new_new_n6971__));
  and1  g3873(.dina(new_new_n4639__), .dinb(new_new_n4541__), .dout(new_new_n6972__));
  or1   g3874(.dina(new_new_n4638__), .dinb(new_new_n10213__), .dout(new_new_n6973__));
  and1  g3875(.dina(new_new_n6972__), .dinb(new_new_n4625__), .dout(new_new_n6974__));
  or1   g3876(.dina(new_new_n6973__), .dinb(new_new_n4624__), .dout(new_new_n6975__));
  and1  g3877(.dina(new_new_n6974__), .dinb(new_new_n4629__), .dout(new_new_n6976__));
  or1   g3878(.dina(new_new_n6975__), .dinb(new_new_n4628__), .dout(new_new_n6977__));
  and1  g3879(.dina(new_new_n6976__), .dinb(new_new_n4633__), .dout(new_new_n6978__));
  or1   g3880(.dina(new_new_n6977__), .dinb(new_new_n4632__), .dout(new_new_n6979__));
  and1  g3881(.dina(new_new_n4648__), .dinb(new_new_n4645__), .dout(new_new_n6980__));
  or1   g3882(.dina(new_new_n4649__), .dinb(new_new_n4644__), .dout(new_new_n6981__));
  and1  g3883(.dina(new_new_n10214__), .dinb(new_new_n10215__), .dout(new_new_n6982__));
  or1   g3884(.dina(new_new_n10216__), .dinb(new_new_n10217__), .dout(new_new_n6983__));
  and1  g3885(.dina(new_new_n10216__), .dinb(new_new_n10217__), .dout(new_new_n6984__));
  or1   g3886(.dina(new_new_n10214__), .dinb(new_new_n10215__), .dout(new_new_n6985__));
  and1  g3887(.dina(new_new_n6985__), .dinb(new_new_n6983__), .dout(new_new_n6986__));
  or1   g3888(.dina(new_new_n6984__), .dinb(new_new_n6982__), .dout(new_new_n6987__));
  and1  g3889(.dina(new_new_n10218__), .dinb(new_new_n10220__), .dout(new_new_n6988__));
  or1   g3890(.dina(new_new_n10222__), .dinb(new_new_n10225__), .dout(new_new_n6989__));
  and1  g3891(.dina(new_new_n10222__), .dinb(new_new_n10225__), .dout(new_new_n6990__));
  or1   g3892(.dina(new_new_n10218__), .dinb(new_new_n10220__), .dout(new_new_n6991__));
  and1  g3893(.dina(new_new_n6991__), .dinb(new_new_n6989__), .dout(new_new_n6992__));
  or1   g3894(.dina(new_new_n6990__), .dinb(new_new_n6988__), .dout(new_new_n6993__));
  or1   g3895(.dina(new_new_n6993__), .dinb(new_new_n10228__), .dout(new_new_n6994__));
  or1   g3896(.dina(new_new_n6992__), .dinb(new_new_n10229__), .dout(new_new_n6995__));
  and1  g3897(.dina(new_new_n6995__), .dinb(new_new_n6994__), .dout(new_new_n6996__));
  and1  g3898(.dina(new_new_n4641__), .dinb(new_new_n4539__), .dout(new_new_n6997__));
  or1   g3899(.dina(new_new_n4640__), .dinb(new_new_n10230__), .dout(new_new_n6998__));
  and1  g3900(.dina(new_new_n6997__), .dinb(new_new_n4627__), .dout(new_new_n6999__));
  or1   g3901(.dina(new_new_n6998__), .dinb(new_new_n4626__), .dout(new_new_n7000__));
  and1  g3902(.dina(new_new_n6999__), .dinb(new_new_n4635__), .dout(new_new_n7001__));
  or1   g3903(.dina(new_new_n7000__), .dinb(new_new_n4634__), .dout(new_new_n7002__));
  and1  g3904(.dina(new_new_n7001__), .dinb(new_new_n4637__), .dout(new_new_n7003__));
  or1   g3905(.dina(new_new_n7002__), .dinb(new_new_n4636__), .dout(new_new_n7004__));
  and1  g3906(.dina(new_new_n4647__), .dinb(new_new_n4643__), .dout(new_new_n7005__));
  or1   g3907(.dina(new_new_n4646__), .dinb(new_new_n4642__), .dout(new_new_n7006__));
  and1  g3908(.dina(new_new_n10231__), .dinb(new_new_n10232__), .dout(new_new_n7007__));
  or1   g3909(.dina(new_new_n10233__), .dinb(new_new_n10234__), .dout(new_new_n7008__));
  and1  g3910(.dina(new_new_n10233__), .dinb(new_new_n10234__), .dout(new_new_n7009__));
  or1   g3911(.dina(new_new_n10231__), .dinb(new_new_n10232__), .dout(new_new_n7010__));
  and1  g3912(.dina(new_new_n7010__), .dinb(new_new_n7008__), .dout(new_new_n7011__));
  or1   g3913(.dina(new_new_n7009__), .dinb(new_new_n7007__), .dout(new_new_n7012__));
  and1  g3914(.dina(new_new_n10235__), .dinb(new_new_n10238__), .dout(new_new_n7013__));
  or1   g3915(.dina(new_new_n10240__), .dinb(new_new_n10242__), .dout(new_new_n7014__));
  and1  g3916(.dina(new_new_n10240__), .dinb(new_new_n10242__), .dout(new_new_n7015__));
  or1   g3917(.dina(new_new_n10235__), .dinb(new_new_n10238__), .dout(new_new_n7016__));
  and1  g3918(.dina(new_new_n7016__), .dinb(new_new_n7014__), .dout(new_new_n7017__));
  or1   g3919(.dina(new_new_n7015__), .dinb(new_new_n7013__), .dout(new_new_n7018__));
  or1   g3920(.dina(new_new_n7018__), .dinb(new_new_n10245__), .dout(new_new_n7019__));
  or1   g3921(.dina(new_new_n7017__), .dinb(new_new_n10246__), .dout(new_new_n7020__));
  and1  g3922(.dina(new_new_n7020__), .dinb(new_new_n7019__), .dout(new_new_n7021__));
  and1  g3923(.dina(new_new_n10248__), .dinb(new_new_n10250__), .dout(new_new_n7022__));
  or1   g3924(.dina(new_new_n10252__), .dinb(new_new_n4543__), .dout(new_new_n7023__));
  and1  g3925(.dina(new_new_n10255__), .dinb(new_new_n10260__), .dout(new_new_n7024__));
  or1   g3926(.dina(new_new_n10262__), .dinb(new_new_n10264__), .dout(new_new_n7025__));
  and1  g3927(.dina(new_new_n7024__), .dinb(new_new_n10248__), .dout(new_new_n7026__));
  or1   g3928(.dina(new_new_n7025__), .dinb(new_new_n10252__), .dout(new_new_n7027__));
  and1  g3929(.dina(new_new_n10266__), .dinb(new_new_n10255__), .dout(new_new_n7028__));
  or1   g3930(.dina(new_new_n10269__), .dinb(new_new_n10262__), .dout(new_new_n7029__));
  and1  g3931(.dina(new_new_n7028__), .dinb(new_new_n10249__), .dout(new_new_n7030__));
  or1   g3932(.dina(new_new_n7029__), .dinb(new_new_n10251__), .dout(new_new_n7031__));
  and1  g3933(.dina(new_new_n7023__), .dinb(new_new_n6282__), .dout(new_new_n7032__));
  or1   g3934(.dina(new_new_n7022__), .dinb(new_new_n10270__), .dout(new_new_n7033__));
  and1  g3935(.dina(new_new_n7032__), .dinb(new_new_n7027__), .dout(new_new_n7034__));
  or1   g3936(.dina(new_new_n7033__), .dinb(new_new_n7026__), .dout(new_new_n7035__));
  and1  g3937(.dina(new_new_n10272__), .dinb(new_new_n7031__), .dout(new_new_n7036__));
  or1   g3938(.dina(new_new_n10274__), .dinb(new_new_n7030__), .dout(new_new_n7037__));
  and1  g3939(.dina(new_new_n10276__), .dinb(new_new_n4651__), .dout(new_new_n7038__));
  or1   g3940(.dina(new_new_n10278__), .dinb(new_new_n4650__), .dout(new_new_n7039__));
  and1  g3941(.dina(new_new_n4241__), .dinb(new_new_n4235__), .dout(new_new_n7040__));
  or1   g3942(.dina(new_new_n10279__), .dinb(new_new_n10280__), .dout(new_new_n7041__));
  and1  g3943(.dina(new_new_n10281__), .dinb(new_new_n10282__), .dout(new_new_n7042__));
  or1   g3944(.dina(new_new_n10283__), .dinb(new_new_n10284__), .dout(new_new_n7043__));
  and1  g3945(.dina(new_new_n10283__), .dinb(new_new_n10284__), .dout(new_new_n7044__));
  or1   g3946(.dina(new_new_n10281__), .dinb(new_new_n10282__), .dout(new_new_n7045__));
  and1  g3947(.dina(new_new_n7045__), .dinb(new_new_n7043__), .dout(new_new_n7046__));
  or1   g3948(.dina(new_new_n7044__), .dinb(new_new_n7042__), .dout(new_new_n7047__));
  and1  g3949(.dina(new_new_n10285__), .dinb(new_new_n10286__), .dout(new_new_n7048__));
  or1   g3950(.dina(new_new_n10287__), .dinb(new_new_n10288__), .dout(new_new_n7049__));
  and1  g3951(.dina(new_new_n10287__), .dinb(new_new_n10288__), .dout(new_new_n7050__));
  or1   g3952(.dina(new_new_n10285__), .dinb(new_new_n10286__), .dout(new_new_n7051__));
  and1  g3953(.dina(new_new_n7051__), .dinb(new_new_n7049__), .dout(new_new_n7052__));
  or1   g3954(.dina(new_new_n7050__), .dinb(new_new_n7048__), .dout(new_new_n7053__));
  and1  g3955(.dina(new_new_n7052__), .dinb(new_new_n10269__), .dout(new_new_n7054__));
  and1  g3956(.dina(new_new_n7053__), .dinb(new_new_n10266__), .dout(new_new_n7055__));
  or1   g3957(.dina(new_new_n7055__), .dinb(new_new_n7054__), .dout(new_new_n7056__));
  and1  g3958(.dina(new_new_n10276__), .dinb(new_new_n10260__), .dout(new_new_n7057__));
  or1   g3959(.dina(new_new_n10278__), .dinb(new_new_n10264__), .dout(new_new_n7058__));
  and1  g3960(.dina(new_new_n10277__), .dinb(new_new_n10263__), .dout(new_new_n7059__));
  or1   g3961(.dina(new_new_n10275__), .dinb(new_new_n10261__), .dout(new_new_n7060__));
  and1  g3962(.dina(new_new_n7060__), .dinb(new_new_n7058__), .dout(new_new_n7061__));
  or1   g3963(.dina(new_new_n7059__), .dinb(new_new_n7057__), .dout(new_new_n7062__));
  and1  g3964(.dina(new_new_n10289__), .dinb(new_new_n10272__), .dout(new_new_n7063__));
  or1   g3965(.dina(new_new_n10290__), .dinb(new_new_n10274__), .dout(new_new_n7064__));
  and1  g3966(.dina(new_new_n10290__), .dinb(new_new_n10273__), .dout(new_new_n7065__));
  or1   g3967(.dina(new_new_n10289__), .dinb(new_new_n10271__), .dout(new_new_n7066__));
  and1  g3968(.dina(new_new_n7066__), .dinb(new_new_n7064__), .dout(new_new_n7067__));
  or1   g3969(.dina(new_new_n7065__), .dinb(new_new_n7063__), .dout(new_new_n7068__));
  and1  g3970(.dina(new_new_n7067__), .dinb(new_new_n10268__), .dout(new_new_n7069__));
  and1  g3971(.dina(new_new_n7068__), .dinb(new_new_n10267__), .dout(new_new_n7070__));
  or1   g3972(.dina(new_new_n7070__), .dinb(new_new_n7069__), .dout(new_new_n7071__));
  and1  g3973(.dina(new_new_n10292__), .dinb(new_new_n10294__), .dout(new_new_n7072__));
  or1   g3974(.dina(new_new_n10297__), .dinb(new_new_n4545__), .dout(new_new_n7073__));
  and1  g3975(.dina(new_new_n10303__), .dinb(new_new_n10308__), .dout(new_new_n7074__));
  or1   g3976(.dina(new_new_n10310__), .dinb(new_new_n10312__), .dout(new_new_n7075__));
  and1  g3977(.dina(new_new_n7074__), .dinb(new_new_n10292__), .dout(new_new_n7076__));
  or1   g3978(.dina(new_new_n7075__), .dinb(new_new_n10297__), .dout(new_new_n7077__));
  and1  g3979(.dina(new_new_n10314__), .dinb(new_new_n10303__), .dout(new_new_n7078__));
  or1   g3980(.dina(new_new_n10317__), .dinb(new_new_n10310__), .dout(new_new_n7079__));
  and1  g3981(.dina(new_new_n7078__), .dinb(new_new_n10293__), .dout(new_new_n7080__));
  or1   g3982(.dina(new_new_n7079__), .dinb(new_new_n10298__), .dout(new_new_n7081__));
  and1  g3983(.dina(new_new_n7073__), .dinb(new_new_n10298__), .dout(new_new_n7082__));
  or1   g3984(.dina(new_new_n7072__), .dinb(new_new_n10293__), .dout(new_new_n7083__));
  and1  g3985(.dina(new_new_n7082__), .dinb(new_new_n7077__), .dout(new_new_n7084__));
  or1   g3986(.dina(new_new_n7083__), .dinb(new_new_n7076__), .dout(new_new_n7085__));
  and1  g3987(.dina(new_new_n10319__), .dinb(new_new_n7081__), .dout(new_new_n7086__));
  or1   g3988(.dina(new_new_n10321__), .dinb(new_new_n7080__), .dout(new_new_n7087__));
  and1  g3989(.dina(new_new_n10323__), .dinb(new_new_n4653__), .dout(new_new_n7088__));
  or1   g3990(.dina(new_new_n10325__), .dinb(new_new_n4652__), .dout(new_new_n7089__));
  and1  g3991(.dina(new_new_n4239__), .dinb(new_new_n4237__), .dout(new_new_n7090__));
  or1   g3992(.dina(new_new_n10326__), .dinb(new_new_n10327__), .dout(new_new_n7091__));
  and1  g3993(.dina(new_new_n10328__), .dinb(new_new_n10329__), .dout(new_new_n7092__));
  or1   g3994(.dina(new_new_n10330__), .dinb(new_new_n10331__), .dout(new_new_n7093__));
  and1  g3995(.dina(new_new_n10330__), .dinb(new_new_n10331__), .dout(new_new_n7094__));
  or1   g3996(.dina(new_new_n10328__), .dinb(new_new_n10329__), .dout(new_new_n7095__));
  and1  g3997(.dina(new_new_n7095__), .dinb(new_new_n7093__), .dout(new_new_n7096__));
  or1   g3998(.dina(new_new_n7094__), .dinb(new_new_n7092__), .dout(new_new_n7097__));
  and1  g3999(.dina(new_new_n10332__), .dinb(new_new_n10333__), .dout(new_new_n7098__));
  or1   g4000(.dina(new_new_n10334__), .dinb(new_new_n10335__), .dout(new_new_n7099__));
  and1  g4001(.dina(new_new_n10334__), .dinb(new_new_n10335__), .dout(new_new_n7100__));
  or1   g4002(.dina(new_new_n10332__), .dinb(new_new_n10333__), .dout(new_new_n7101__));
  and1  g4003(.dina(new_new_n7101__), .dinb(new_new_n7099__), .dout(new_new_n7102__));
  or1   g4004(.dina(new_new_n7100__), .dinb(new_new_n7098__), .dout(new_new_n7103__));
  or1   g4005(.dina(new_new_n7103__), .dinb(new_new_n10314__), .dout(new_new_n7104__));
  or1   g4006(.dina(new_new_n7102__), .dinb(new_new_n10317__), .dout(new_new_n7105__));
  and1  g4007(.dina(new_new_n7105__), .dinb(new_new_n7104__), .dout(new_new_n7106__));
  and1  g4008(.dina(new_new_n10323__), .dinb(new_new_n10308__), .dout(new_new_n7107__));
  or1   g4009(.dina(new_new_n10325__), .dinb(new_new_n10312__), .dout(new_new_n7108__));
  and1  g4010(.dina(new_new_n10324__), .dinb(new_new_n10311__), .dout(new_new_n7109__));
  or1   g4011(.dina(new_new_n10322__), .dinb(new_new_n10309__), .dout(new_new_n7110__));
  and1  g4012(.dina(new_new_n7110__), .dinb(new_new_n7108__), .dout(new_new_n7111__));
  or1   g4013(.dina(new_new_n7109__), .dinb(new_new_n7107__), .dout(new_new_n7112__));
  and1  g4014(.dina(new_new_n10336__), .dinb(new_new_n10319__), .dout(new_new_n7113__));
  or1   g4015(.dina(new_new_n10337__), .dinb(new_new_n10321__), .dout(new_new_n7114__));
  and1  g4016(.dina(new_new_n10337__), .dinb(new_new_n10320__), .dout(new_new_n7115__));
  or1   g4017(.dina(new_new_n10336__), .dinb(new_new_n10318__), .dout(new_new_n7116__));
  and1  g4018(.dina(new_new_n7116__), .dinb(new_new_n7114__), .dout(new_new_n7117__));
  or1   g4019(.dina(new_new_n7115__), .dinb(new_new_n7113__), .dout(new_new_n7118__));
  or1   g4020(.dina(new_new_n7118__), .dinb(new_new_n10315__), .dout(new_new_n7119__));
  or1   g4021(.dina(new_new_n7117__), .dinb(new_new_n10316__), .dout(new_new_n7120__));
  and1  g4022(.dina(new_new_n7120__), .dinb(new_new_n7119__), .dout(new_new_n7121__));
  and1  g4023(.dina(new_new_n9830__), .dinb(new_new_n10338__), .dout(new_new_n7122__));
  and1  g4024(.dina(new_new_n9835__), .dinb(new_new_n3392__), .dout(new_new_n7123__));
  or1   g4025(.dina(new_new_n7123__), .dinb(new_new_n7122__), .dout(new_new_n7124__));
  and1  g4026(.dina(new_new_n10340__), .dinb(new_new_n10342__), .dout(new_new_n7125__));
  or1   g4027(.dina(new_new_n10344__), .dinb(new_new_n10346__), .dout(new_new_n7126__));
  and1  g4028(.dina(new_new_n10344__), .dinb(new_new_n10346__), .dout(new_new_n7127__));
  or1   g4029(.dina(new_new_n10340__), .dinb(new_new_n10342__), .dout(new_new_n7128__));
  and1  g4030(.dina(new_new_n7128__), .dinb(new_new_n7126__), .dout(new_new_n7129__));
  or1   g4031(.dina(new_new_n7127__), .dinb(new_new_n7125__), .dout(new_new_n7130__));
  and1  g4032(.dina(new_new_n6365__), .dinb(new_new_n10348__), .dout(new_new_n7131__));
  and1  g4033(.dina(new_new_n10350__), .dinb(new_new_n3551__), .dout(new_new_n7132__));
  or1   g4034(.dina(new_new_n7132__), .dinb(new_new_n7131__), .dout(new_new_n7133__));
  and1  g4035(.dina(new_new_n6377__), .dinb(new_new_n10352__), .dout(new_new_n7134__));
  and1  g4036(.dina(new_new_n10354__), .dinb(new_new_n3579__), .dout(new_new_n7135__));
  or1   g4037(.dina(new_new_n7135__), .dinb(new_new_n7134__), .dout(new_new_n7136__));
  and1  g4038(.dina(new_new_n6371__), .dinb(new_new_n10356__), .dout(new_new_n7137__));
  and1  g4039(.dina(new_new_n10358__), .dinb(new_new_n3583__), .dout(new_new_n7138__));
  or1   g4040(.dina(new_new_n7138__), .dinb(new_new_n7137__), .dout(new_new_n7139__));
  and1  g4041(.dina(new_new_n10360__), .dinb(new_new_n10362__), .dout(new_new_n7140__));
  and1  g4042(.dina(new_new_n7140__), .dinb(new_new_n4129__), .dout(new_new_n7141__));
  and1  g4043(.dina(new_new_n10360__), .dinb(new_new_n10364__), .dout(new_new_n7142__));
  and1  g4044(.dina(new_new_n7142__), .dinb(new_new_n10366__), .dout(new_new_n7143__));
  and1  g4045(.dina(new_new_n9917__), .dinb(new_new_n10362__), .dout(new_new_n7144__));
  and1  g4046(.dina(new_new_n7144__), .dinb(new_new_n9711__), .dout(new_new_n7145__));
  and1  g4047(.dina(new_new_n9918__), .dinb(new_new_n10364__), .dout(new_new_n7146__));
  and1  g4048(.dina(new_new_n7146__), .dinb(new_new_n9709__), .dout(new_new_n7147__));
  and1  g4049(.dina(new_new_n9921__), .dinb(new_new_n10361__), .dout(new_new_n7148__));
  and1  g4050(.dina(new_new_n7148__), .dinb(new_new_n9704__), .dout(new_new_n7149__));
  and1  g4051(.dina(new_new_n9922__), .dinb(new_new_n10363__), .dout(new_new_n7150__));
  and1  g4052(.dina(new_new_n7150__), .dinb(new_new_n9702__), .dout(new_new_n7151__));
  or1   g4053(.dina(new_new_n10339__), .dinb(new_new_n10345__), .dout(new_new_n7152__));
  and1  g4054(.dina(new_new_n10350__), .dinb(new_new_n10348__), .dout(new_new_n7153__));
  and1  g4055(.dina(new_new_n10354__), .dinb(new_new_n10352__), .dout(new_new_n7154__));
  and1  g4056(.dina(new_new_n10358__), .dinb(new_new_n10356__), .dout(new_new_n7155__));
  and1  g4057(.dina(new_new_n10369__), .dinb(new_new_n10370__), .dout(new_new_n7156__));
  and1  g4058(.dina(new_new_n10371__), .dinb(new_new_n10372__), .dout(new_new_n7157__));
  or1   g4059(.dina(new_new_n10373__), .dinb(new_new_n10374__), .dout(new_new_n7158__));
  and1  g4060(.dina(new_new_n10373__), .dinb(new_new_n10374__), .dout(new_new_n7159__));
  or1   g4061(.dina(new_new_n10371__), .dinb(new_new_n10372__), .dout(new_new_n7160__));
  and1  g4062(.dina(new_new_n7160__), .dinb(new_new_n7158__), .dout(new_new_n7161__));
  or1   g4063(.dina(new_new_n7159__), .dinb(new_new_n7157__), .dout(new_new_n7162__));
  and1  g4064(.dina(new_new_n10375__), .dinb(new_new_n10221__), .dout(new_new_n7163__));
  or1   g4065(.dina(new_new_n10376__), .dinb(new_new_n10224__), .dout(new_new_n7164__));
  and1  g4066(.dina(new_new_n10376__), .dinb(new_new_n10226__), .dout(new_new_n7165__));
  or1   g4067(.dina(new_new_n10375__), .dinb(new_new_n10221__), .dout(new_new_n7166__));
  and1  g4068(.dina(new_new_n7166__), .dinb(new_new_n7164__), .dout(new_new_n7167__));
  or1   g4069(.dina(new_new_n7165__), .dinb(new_new_n7163__), .dout(new_new_n7168__));
  and1  g4070(.dina(new_new_n7167__), .dinb(new_new_n10229__), .dout(new_new_n7169__));
  and1  g4071(.dina(new_new_n7168__), .dinb(new_new_n10228__), .dout(new_new_n7170__));
  or1   g4072(.dina(new_new_n7170__), .dinb(new_new_n7169__), .dout(new_new_n7171__));
  and1  g4073(.dina(new_new_n10377__), .dinb(new_new_n10380__), .dout(new_new_n7172__));
  and1  g4074(.dina(new_new_n10382__), .dinb(new_new_n10383__), .dout(new_new_n7173__));
  or1   g4075(.dina(new_new_n10384__), .dinb(new_new_n10385__), .dout(new_new_n7174__));
  and1  g4076(.dina(new_new_n10384__), .dinb(new_new_n10385__), .dout(new_new_n7175__));
  or1   g4077(.dina(new_new_n10382__), .dinb(new_new_n10383__), .dout(new_new_n7176__));
  and1  g4078(.dina(new_new_n7176__), .dinb(new_new_n7174__), .dout(new_new_n7177__));
  or1   g4079(.dina(new_new_n7175__), .dinb(new_new_n7173__), .dout(new_new_n7178__));
  and1  g4080(.dina(new_new_n10386__), .dinb(new_new_n10237__), .dout(new_new_n7179__));
  or1   g4081(.dina(new_new_n10387__), .dinb(new_new_n10243__), .dout(new_new_n7180__));
  and1  g4082(.dina(new_new_n10387__), .dinb(new_new_n10243__), .dout(new_new_n7181__));
  or1   g4083(.dina(new_new_n10386__), .dinb(new_new_n10239__), .dout(new_new_n7182__));
  and1  g4084(.dina(new_new_n7182__), .dinb(new_new_n7180__), .dout(new_new_n7183__));
  or1   g4085(.dina(new_new_n7181__), .dinb(new_new_n7179__), .dout(new_new_n7184__));
  and1  g4086(.dina(new_new_n7183__), .dinb(new_new_n10246__), .dout(new_new_n7185__));
  and1  g4087(.dina(new_new_n7184__), .dinb(new_new_n10245__), .dout(new_new_n7186__));
  or1   g4088(.dina(new_new_n7186__), .dinb(new_new_n7185__), .dout(new_new_n7187__));
  and1  g4089(.dina(new_new_n10388__), .dinb(new_new_n10391__), .dout(new_new_n7188__));
  or1   g4090(.dina(new_new_n10369__), .dinb(new_new_n10370__), .dout(new_new_n7189__));
  or1   g4091(.dina(new_new_n10377__), .dinb(new_new_n10380__), .dout(new_new_n7190__));
  or1   g4092(.dina(new_new_n10388__), .dinb(new_new_n10391__), .dout(new_new_n7191__));
  and1  g4093(.dina(new_new_n9699__), .dinb(new_new_n10393__), .dout(new_new_n7192__));
  and1  g4094(.dina(new_new_n9705__), .dinb(new_new_n10394__), .dout(new_new_n7193__));
  or1   g4095(.dina(new_new_n7193__), .dinb(new_new_n7192__), .dout(new_new_n7194__));
  and1  g4096(.dina(new_new_n6552__), .dinb(new_new_n10208__), .dout(new_new_n7195__));
  and1  g4097(.dina(new_new_n10206__), .dinb(new_new_n3559__), .dout(new_new_n7196__));
  or1   g4098(.dina(new_new_n7196__), .dinb(new_new_n7195__), .dout(new_new_n7197__));
  and1  g4099(.dina(new_new_n6546__), .dinb(new_new_n10212__), .dout(new_new_n7198__));
  and1  g4100(.dina(new_new_n10210__), .dinb(new_new_n3587__), .dout(new_new_n7199__));
  or1   g4101(.dina(new_new_n7199__), .dinb(new_new_n7198__), .dout(new_new_n7200__));
  and1  g4102(.dina(new_new_n9824__), .dinb(new_new_n3480__), .dout(new_new_n7201__));
  and1  g4103(.dina(new_new_n10396__), .dinb(new_new_n10399__), .dout(new_new_n7202__));
  or1   g4104(.dina(new_new_n10401__), .dinb(new_new_n10402__), .dout(new_new_n7203__));
  and1  g4105(.dina(new_new_n10403__), .dinb(new_new_n10406__), .dout(new_new_n7204__));
  and1  g4106(.dina(new_new_n10409__), .dinb(new_new_n10411__), .dout(new_new_n7205__));
  or1   g4107(.dina(new_new_n10413__), .dinb(new_new_n10414__), .dout(new_new_n7206__));
  or1   g4108(.dina(new_new_n10415__), .dinb(new_new_n10417__), .dout(new_new_n7207__));
  and1  g4109(.dina(new_new_n10421__), .dinb(new_new_n10396__), .dout(new_new_n7208__));
  or1   g4110(.dina(new_new_n10425__), .dinb(new_new_n10401__), .dout(new_new_n7209__));
  and1  g4111(.dina(new_new_n7208__), .dinb(new_new_n10428__), .dout(new_new_n7210__));
  or1   g4112(.dina(new_new_n7209__), .dinb(new_new_n10431__), .dout(new_new_n7211__));
  and1  g4113(.dina(new_new_n10433__), .dinb(new_new_n10406__), .dout(new_new_n7212__));
  and1  g4114(.dina(new_new_n9819__), .dinb(new_new_n10434__), .dout(new_new_n7213__));
  and1  g4115(.dina(new_new_n10436__), .dinb(new_new_n10397__), .dout(new_new_n7214__));
  or1   g4116(.dina(new_new_n6355__), .dinb(new_new_n10400__), .dout(new_new_n7215__));
  and1  g4117(.dina(new_new_n10437__), .dinb(new_new_n10405__), .dout(new_new_n7216__));
  and1  g4118(.dina(new_new_n7216__), .dinb(new_new_n10421__), .dout(new_new_n7217__));
  and1  g4119(.dina(new_new_n10439__), .dinb(new_new_n10409__), .dout(new_new_n7218__));
  or1   g4120(.dina(new_new_n10441__), .dinb(new_new_n10413__), .dout(new_new_n7219__));
  and1  g4121(.dina(new_new_n7218__), .dinb(new_new_n10444__), .dout(new_new_n7220__));
  or1   g4122(.dina(new_new_n7219__), .dinb(new_new_n10448__), .dout(new_new_n7221__));
  or1   g4123(.dina(new_new_n10453__), .dinb(new_new_n10417__), .dout(new_new_n7222__));
  or1   g4124(.dina(new_new_n10412__), .dinb(new_new_n10448__), .dout(new_new_n7223__));
  or1   g4125(.dina(new_new_n10454__), .dinb(new_new_n10418__), .dout(new_new_n7224__));
  or1   g4126(.dina(new_new_n7224__), .dinb(new_new_n10441__), .dout(new_new_n7225__));
  and1  g4127(.dina(new_new_n10407__), .dinb(new_new_n10456__), .dout(new_new_n7226__));
  or1   g4128(.dina(new_new_n10418__), .dinb(new_new_n10457__), .dout(new_new_n7227__));
  or1   g4129(.dina(new_new_n10454__), .dinb(new_new_n10442__), .dout(new_new_n7228__));
  and1  g4130(.dina(new_new_n10415__), .dinb(new_new_n10457__), .dout(new_new_n7229__));
  or1   g4131(.dina(new_new_n7205__), .dinb(new_new_n10458__), .dout(new_new_n7230__));
  and1  g4132(.dina(new_new_n7229__), .dinb(new_new_n10453__), .dout(new_new_n7231__));
  or1   g4133(.dina(new_new_n7230__), .dinb(new_new_n7220__), .dout(new_new_n7232__));
  and1  g4134(.dina(new_new_n10460__), .dinb(new_new_n7228__), .dout(new_new_n7233__));
  and1  g4135(.dina(new_new_n10439__), .dinb(new_new_n10444__), .dout(new_new_n7234__));
  or1   g4136(.dina(new_new_n10442__), .dinb(new_new_n10449__), .dout(new_new_n7235__));
  and1  g4137(.dina(new_new_n7235__), .dinb(new_new_n10414__), .dout(new_new_n7236__));
  or1   g4138(.dina(new_new_n10461__), .dinb(new_new_n10411__), .dout(new_new_n7237__));
  or1   g4139(.dina(new_new_n10462__), .dinb(new_new_n10461__), .dout(new_new_n7238__));
  or1   g4140(.dina(new_new_n10463__), .dinb(new_new_n10464__), .dout(new_new_n7239__));
  and1  g4141(.dina(new_new_n10422__), .dinb(new_new_n10428__), .dout(new_new_n7240__));
  or1   g4142(.dina(new_new_n10425__), .dinb(new_new_n10431__), .dout(new_new_n7241__));
  and1  g4143(.dina(new_new_n7241__), .dinb(new_new_n10402__), .dout(new_new_n7242__));
  or1   g4144(.dina(new_new_n7240__), .dinb(new_new_n10399__), .dout(new_new_n7243__));
  and1  g4145(.dina(new_new_n10436__), .dinb(new_new_n10422__), .dout(new_new_n7244__));
  or1   g4146(.dina(new_new_n7244__), .dinb(new_new_n10465__), .dout(new_new_n7245__));
  and1  g4147(.dina(new_new_n10437__), .dinb(new_new_n10423__), .dout(new_new_n7246__));
  or1   g4148(.dina(new_new_n7215__), .dinb(new_new_n10424__), .dout(new_new_n7247__));
  and1  g4149(.dina(new_new_n7203__), .dinb(new_new_n6348__), .dout(new_new_n7248__));
  or1   g4150(.dina(new_new_n10403__), .dinb(new_new_n10456__), .dout(new_new_n7249__));
  and1  g4151(.dina(new_new_n7248__), .dinb(new_new_n7211__), .dout(new_new_n7250__));
  or1   g4152(.dina(new_new_n7249__), .dinb(new_new_n10433__), .dout(new_new_n7251__));
  and1  g4153(.dina(new_new_n10467__), .dinb(new_new_n7247__), .dout(new_new_n7252__));
  or1   g4154(.dina(new_new_n10469__), .dinb(new_new_n7246__), .dout(new_new_n7253__));
  and1  g4155(.dina(new_new_n9786__), .dinb(new_new_n9789__), .dout(new_new_n7254__));
  or1   g4156(.dina(new_new_n9779__), .dinb(new_new_n9783__), .dout(new_new_n7255__));
  or1   g4157(.dina(new_new_n7254__), .dinb(new_new_n7252__), .dout(new_new_n7256__));
  or1   g4158(.dina(new_new_n7255__), .dinb(new_new_n7253__), .dout(new_new_n7257__));
  and1  g4159(.dina(new_new_n7257__), .dinb(new_new_n7256__), .dout(new_new_n7258__));
  and1  g4160(.dina(new_new_n10470__), .dinb(new_new_n10471__), .dout(new_new_n7259__));
  and1  g4161(.dina(new_new_n10463__), .dinb(new_new_n10464__), .dout(new_new_n7260__));
  or1   g4162(.dina(new_new_n10470__), .dinb(new_new_n10471__), .dout(new_new_n7261__));
  and1  g4163(.dina(new_new_n10472__), .dinb(new_new_n10474__), .dout(new_new_n7262__));
  and1  g4164(.dina(new_new_n10475__), .dinb(new_new_n10477__), .dout(new_new_n7263__));
  or1   g4165(.dina(new_new_n10478__), .dinb(new_new_n10479__), .dout(new_new_n7264__));
  or1   g4166(.dina(new_new_n7264__), .dinb(new_new_n10480__), .dout(new_new_n7265__));
  or1   g4167(.dina(new_new_n7265__), .dinb(new_new_n10481__), .dout(new_new_n7266__));
  and1  g4168(.dina(new_new_n10482__), .dinb(new_new_n10483__), .dout(new_new_n7267__));
  and1  g4169(.dina(new_new_n7267__), .dinb(new_new_n10484__), .dout(new_new_n7268__));
  and1  g4170(.dina(new_new_n7268__), .dinb(new_new_n10485__), .dout(new_new_n7269__));
  and1  g4171(.dina(new_new_n10474__), .dinb(new_new_n10486__), .dout(new_new_n7270__));
  or1   g4172(.dina(new_new_n7270__), .dinb(new_new_n10487__), .dout(new_new_n7271__));
  and1  g4173(.dina(new_new_n10477__), .dinb(new_new_n10488__), .dout(new_new_n7272__));
  or1   g4174(.dina(new_new_n7272__), .dinb(new_new_n10489__), .dout(new_new_n7273__));
  and1  g4175(.dina(new_new_n10467__), .dinb(new_new_n10427__), .dout(new_new_n7274__));
  or1   g4176(.dina(new_new_n10469__), .dinb(new_new_n10432__), .dout(new_new_n7275__));
  and1  g4177(.dina(new_new_n10468__), .dinb(new_new_n10432__), .dout(new_new_n7276__));
  or1   g4178(.dina(new_new_n10466__), .dinb(new_new_n10429__), .dout(new_new_n7277__));
  and1  g4179(.dina(new_new_n7277__), .dinb(new_new_n7275__), .dout(new_new_n7278__));
  or1   g4180(.dina(new_new_n7276__), .dinb(new_new_n7274__), .dout(new_new_n7279__));
  or1   g4181(.dina(new_new_n7279__), .dinb(new_new_n10465__), .dout(new_new_n7280__));
  or1   g4182(.dina(new_new_n7278__), .dinb(new_new_n7242__), .dout(new_new_n7281__));
  and1  g4183(.dina(new_new_n7281__), .dinb(new_new_n7280__), .dout(new_new_n7282__));
  and1  g4184(.dina(new_new_n10460__), .dinb(new_new_n10445__), .dout(new_new_n7283__));
  or1   g4185(.dina(new_new_n10490__), .dinb(new_new_n10449__), .dout(new_new_n7284__));
  and1  g4186(.dina(new_new_n10490__), .dinb(new_new_n10451__), .dout(new_new_n7285__));
  or1   g4187(.dina(new_new_n10459__), .dinb(new_new_n10445__), .dout(new_new_n7286__));
  and1  g4188(.dina(new_new_n7286__), .dinb(new_new_n7284__), .dout(new_new_n7287__));
  or1   g4189(.dina(new_new_n7285__), .dinb(new_new_n7283__), .dout(new_new_n7288__));
  and1  g4190(.dina(new_new_n7287__), .dinb(new_new_n7236__), .dout(new_new_n7289__));
  and1  g4191(.dina(new_new_n7288__), .dinb(new_new_n10462__), .dout(new_new_n7290__));
  or1   g4192(.dina(new_new_n7290__), .dinb(new_new_n7289__), .dout(new_new_n7291__));
  and1  g4193(.dina(new_new_n10491__), .dinb(new_new_n10494__), .dout(new_new_n7292__));
  and1  g4194(.dina(new_new_n10496__), .dinb(new_new_n10497__), .dout(new_new_n7293__));
  or1   g4195(.dina(new_new_n7293__), .dinb(new_new_n7292__), .dout(new_new_n7294__));
  and1  g4196(.dina(new_new_n10498__), .dinb(new_new_n10494__), .dout(new_new_n7295__));
  and1  g4197(.dina(new_new_n10499__), .dinb(new_new_n10497__), .dout(new_new_n7296__));
  or1   g4198(.dina(new_new_n7296__), .dinb(new_new_n7295__), .dout(new_new_n7297__));
  and1  g4199(.dina(new_new_n10502__), .dinb(new_new_n10505__), .dout(new_new_n7298__));
  and1  g4200(.dina(new_new_n10507__), .dinb(new_new_n2538__), .dout(new_new_n7299__));
  or1   g4201(.dina(new_new_n7299__), .dinb(new_new_n7298__), .dout(new_new_n7300__));
  and1  g4202(.dina(new_new_n10502__), .dinb(new_new_n10508__), .dout(new_new_n7301__));
  and1  g4203(.dina(new_new_n10507__), .dinb(new_new_n2542__), .dout(new_new_n7302__));
  or1   g4204(.dina(new_new_n7302__), .dinb(new_new_n7301__), .dout(new_new_n7303__));
  and1  g4205(.dina(new_new_n10503__), .dinb(new_new_n10509__), .dout(new_new_n7304__));
  and1  g4206(.dina(new_new_n10506__), .dinb(new_new_n2546__), .dout(new_new_n7305__));
  or1   g4207(.dina(new_new_n7305__), .dinb(new_new_n7304__), .dout(new_new_n7306__));
  buf1  g4208(.din(new_new_n8486__), .dout(G5193));
  buf1  g4209(.din(new_new_n8501__), .dout(G5194));
  buf1  g4210(.din(new_new_n8445__), .dout(G5195));
  buf1  g4211(.din(new_new_n10511__), .dout(G5196));
  buf1  g4212(.din(new_new_n3511__), .dout(G5197));
  buf1  g4213(.din(new_new_n3519__), .dout(G5198));
  buf1  g4214(.din(new_new_n4710__), .dout(G5199));
  buf1  g4215(.din(new_new_n3619__), .dout(G5200));
  buf1  g4216(.din(G5196), .dout(G5201));
  buf1  g4217(.din(new_new_n10510__), .dout(G5202));
  buf1  g4218(.din(new_new_n3507__), .dout(G5203));
  buf1  g4219(.din(new_new_n3515__), .dout(G5204));
  buf1  g4220(.din(new_new_n4711__), .dout(G5205));
  buf1  g4221(.din(new_new_n9477__), .dout(G5206));
  buf1  g4222(.din(new_new_n9471__), .dout(G5207));
  buf1  g4223(.din(new_new_n9473__), .dout(G5208));
  buf1  g4224(.din(new_new_n9470__), .dout(G5209));
  buf1  g4225(.din(new_new_n4712__), .dout(G5210));
  buf1  g4226(.din(new_new_n4713__), .dout(G5211));
  buf1  g4227(.din(new_new_n4714__), .dout(G5212));
  buf1  g4228(.din(new_new_n4715__), .dout(G5213));
  buf1  g4229(.din(new_new_n9331__), .dout(G5214));
  buf1  g4230(.din(new_new_n8443__), .dout(G5215));
  buf1  g4231(.din(new_new_n8444__), .dout(G5216));
  buf1  g4232(.din(new_new_n10512__), .dout(G5217));
  buf1  g4233(.din(new_new_n3474__), .dout(G5218));
  buf1  g4234(.din(G5217), .dout(G5219));
  buf1  g4235(.din(new_new_n4718__), .dout(G5220));
  buf1  g4236(.din(new_new_n8460__), .dout(G5221));
  buf1  g4237(.din(new_new_n10514__), .dout(G5222));
  buf1  g4238(.din(G5222), .dout(G5223));
  buf1  g4239(.din(new_new_n10515__), .dout(G5224));
  buf1  g4240(.din(G5224), .dout(G5225));
  buf1  g4241(.din(new_new_n10516__), .dout(G5226));
  buf1  g4242(.din(G5226), .dout(G5227));
  buf1  g4243(.din(new_new_n4722__), .dout(G5228));
  buf1  g4244(.din(new_new_n10517__), .dout(G5229));
  buf1  g4245(.din(G5229), .dout(G5230));
  buf1  g4246(.din(new_new_n4730__), .dout(G5231));
  not1  g4247(.din(new_new_n4740__), .dout(G5232));
  not1  g4248(.din(new_new_n4748__), .dout(G5233));
  not1  g4249(.din(new_new_n4756__), .dout(G5234));
  not1  g4250(.din(new_new_n4764__), .dout(G5235));
  not1  g4251(.din(new_new_n4834__), .dout(G5236));
  not1  g4252(.din(new_new_n4922__), .dout(G5237));
  not1  g4253(.din(new_new_n4926__), .dout(G5238));
  not1  g4254(.din(new_new_n4938__), .dout(G5239));
  not1  g4255(.din(new_new_n4942__), .dout(G5240));
  not1  g4256(.din(new_new_n4954__), .dout(G5241));
  not1  g4257(.din(new_new_n9475__), .dout(G5242));
  not1  g4258(.din(new_new_n9476__), .dout(G5243));
  not1  g4259(.din(new_new_n5060__), .dout(G5244));
  not1  g4260(.din(new_new_n5101__), .dout(G5245));
  not1  g4261(.din(new_new_n5142__), .dout(G5246));
  not1  g4262(.din(new_new_n5153__), .dout(G5247));
  not1  g4263(.din(new_new_n8992__), .dout(G5248));
  not1  g4264(.din(new_new_n9441__), .dout(G5249));
  not1  g4265(.din(new_new_n9034__), .dout(G5250));
  buf1  g4266(.din(new_new_n9468__), .dout(G5251));
  buf1  g4267(.din(new_new_n5232__), .dout(G5252));
  not1  g4268(.din(new_new_n9411__), .dout(G5253));
  not1  g4269(.din(new_new_n9421__), .dout(G5254));
  not1  g4270(.din(new_new_n9431__), .dout(G5255));
  buf1  g4271(.din(new_new_n5314__), .dout(G5256));
  not1  g4272(.din(new_new_n9415__), .dout(G5257));
  not1  g4273(.din(new_new_n9425__), .dout(G5258));
  not1  g4274(.din(new_new_n9435__), .dout(G5259));
  not1  g4275(.din(new_new_n9445__), .dout(G5260));
  not1  g4276(.din(new_new_n9472__), .dout(G5261));
  not1  g4277(.din(new_new_n9474__), .dout(G5262));
  not1  g4278(.din(new_new_n5546__), .dout(G5263));
  not1  g4279(.din(new_new_n5579__), .dout(G5264));
  buf1  g4280(.din(new_new_n5591__), .dout(G5265));
  buf1  g4281(.din(new_new_n5603__), .dout(G5266));
  buf1  g4282(.din(new_new_n5614__), .dout(G5267));
  buf1  g4283(.din(new_new_n5625__), .dout(G5268));
  buf1  g4284(.din(new_new_n5636__), .dout(G5269));
  buf1  g4285(.din(new_new_n5647__), .dout(G5270));
  buf1  g4286(.din(new_new_n5658__), .dout(G5271));
  buf1  g4287(.din(new_new_n5669__), .dout(G5272));
  buf1  g4288(.din(new_new_n5680__), .dout(G5273));
  buf1  g4289(.din(new_new_n5691__), .dout(G5274));
  buf1  g4290(.din(new_new_n5703__), .dout(G5275));
  buf1  g4291(.din(new_new_n5715__), .dout(G5276));
  buf1  g4292(.din(new_new_n5727__), .dout(G5277));
  buf1  g4293(.din(new_new_n5739__), .dout(G5278));
  buf1  g4294(.din(new_new_n5751__), .dout(G5279));
  buf1  g4295(.din(new_new_n5763__), .dout(G5280));
  buf1  g4296(.din(new_new_n5775__), .dout(G5281));
  buf1  g4297(.din(new_new_n5787__), .dout(G5282));
  buf1  g4298(.din(new_new_n5808__), .dout(G5283));
  buf1  g4299(.din(new_new_n5812__), .dout(G5284));
  not1  g4300(.din(new_new_n9483__), .dout(G5285));
  not1  g4301(.din(new_new_n9493__), .dout(G5286));
  not1  g4302(.din(new_new_n9503__), .dout(G5287));
  not1  g4303(.din(new_new_n9513__), .dout(G5288));
  not1  g4304(.din(new_new_n5853__), .dout(G5289));
  not1  g4305(.din(new_new_n9487__), .dout(G5290));
  not1  g4306(.din(new_new_n9497__), .dout(G5291));
  not1  g4307(.din(new_new_n9507__), .dout(G5292));
  not1  g4308(.din(new_new_n9517__), .dout(G5293));
  buf1  g4309(.din(new_new_n5906__), .dout(G5294));
  buf1  g4310(.din(new_new_n5917__), .dout(G5295));
  buf1  g4311(.din(new_new_n5928__), .dout(G5296));
  buf1  g4312(.din(new_new_n5939__), .dout(G5297));
  buf1  g4313(.din(new_new_n5950__), .dout(G5298));
  buf1  g4314(.din(new_new_n5961__), .dout(G5299));
  buf1  g4315(.din(new_new_n5972__), .dout(G5300));
  buf1  g4316(.din(new_new_n5983__), .dout(G5301));
  buf1  g4317(.din(new_new_n5995__), .dout(G5302));
  buf1  g4318(.din(new_new_n6007__), .dout(G5303));
  buf1  g4319(.din(new_new_n6019__), .dout(G5304));
  buf1  g4320(.din(new_new_n6031__), .dout(G5305));
  buf1  g4321(.din(new_new_n6043__), .dout(G5306));
  buf1  g4322(.din(new_new_n6055__), .dout(G5307));
  buf1  g4323(.din(new_new_n6067__), .dout(G5308));
  buf1  g4324(.din(new_new_n6079__), .dout(G5309));
  not1  g4325(.din(new_new_n6095__), .dout(G5310));
  not1  g4326(.din(new_new_n6110__), .dout(G5311));
  buf1  g4327(.din(new_new_n6133__), .dout(G5312));
  buf1  g4328(.din(new_new_n6144__), .dout(G5313));
  not1  g4329(.din(new_new_n6156__), .dout(G5314));
  not1  g4330(.din(new_new_n6168__), .dout(G5315));
  buf1  g4331(.din(new_new_n2328__), .dout(n16425));
  buf1  g4332(.din(new_new_n2684__), .dout(n16428));
  buf1  g4333(.din(new_new_n2686__), .dout(n16431));
  buf1  g4334(.din(new_new_n2688__), .dout(n16434));
  buf1  g4335(.din(new_new_n2330__), .dout(n16437));
  buf1  g4336(.din(new_new_n2692__), .dout(n16440));
  buf1  g4337(.din(new_new_n2694__), .dout(n16443));
  buf1  g4338(.din(new_new_n2696__), .dout(n16446));
  buf1  g4339(.din(new_new_n2332__), .dout(n16449));
  buf1  g4340(.din(new_new_n2700__), .dout(n16452));
  buf1  g4341(.din(new_new_n2702__), .dout(n16455));
  buf1  g4342(.din(new_new_n2704__), .dout(n16458));
  buf1  g4343(.din(new_new_n2334__), .dout(n16461));
  buf1  g4344(.din(new_new_n2708__), .dout(n16464));
  buf1  g4345(.din(new_new_n2710__), .dout(n16467));
  buf1  g4346(.din(new_new_n2712__), .dout(n16470));
  buf1  g4347(.din(new_new_n2336__), .dout(n16473));
  buf1  g4348(.din(new_new_n2716__), .dout(n16476));
  buf1  g4349(.din(new_new_n2718__), .dout(n16479));
  buf1  g4350(.din(new_new_n2720__), .dout(n16482));
  buf1  g4351(.din(new_new_n2338__), .dout(n16485));
  buf1  g4352(.din(new_new_n2724__), .dout(n16488));
  buf1  g4353(.din(new_new_n2726__), .dout(n16491));
  buf1  g4354(.din(new_new_n2728__), .dout(n16494));
  buf1  g4355(.din(new_new_n2340__), .dout(n16497));
  buf1  g4356(.din(new_new_n2732__), .dout(n16500));
  buf1  g4357(.din(new_new_n2734__), .dout(n16503));
  buf1  g4358(.din(new_new_n2736__), .dout(n16506));
  buf1  g4359(.din(new_new_n2342__), .dout(n16509));
  buf1  g4360(.din(new_new_n2740__), .dout(n16512));
  buf1  g4361(.din(new_new_n2742__), .dout(n16515));
  buf1  g4362(.din(new_new_n2744__), .dout(n16518));
  buf1  g4363(.din(new_new_n2344__), .dout(n16521));
  buf1  g4364(.din(new_new_n2748__), .dout(n16524));
  buf1  g4365(.din(new_new_n2750__), .dout(n16527));
  buf1  g4366(.din(new_new_n2752__), .dout(n16530));
  buf1  g4367(.din(new_new_n2346__), .dout(n16533));
  buf1  g4368(.din(new_new_n2756__), .dout(n16536));
  buf1  g4369(.din(new_new_n2758__), .dout(n16539));
  buf1  g4370(.din(new_new_n2760__), .dout(n16542));
  buf1  g4371(.din(new_new_n2348__), .dout(n16545));
  buf1  g4372(.din(new_new_n2764__), .dout(n16548));
  buf1  g4373(.din(new_new_n2766__), .dout(n16551));
  buf1  g4374(.din(new_new_n2768__), .dout(n16554));
  buf1  g4375(.din(new_new_n2350__), .dout(n16557));
  buf1  g4376(.din(new_new_n2772__), .dout(n16560));
  buf1  g4377(.din(new_new_n2774__), .dout(n16563));
  buf1  g4378(.din(new_new_n2776__), .dout(n16566));
  buf1  g4379(.din(new_new_n2352__), .dout(n16569));
  buf1  g4380(.din(new_new_n2780__), .dout(n16572));
  buf1  g4381(.din(new_new_n2782__), .dout(n16575));
  buf1  g4382(.din(new_new_n2784__), .dout(n16578));
  buf1  g4383(.din(new_new_n2354__), .dout(n16581));
  buf1  g4384(.din(new_new_n2788__), .dout(n16584));
  buf1  g4385(.din(new_new_n2790__), .dout(n16587));
  buf1  g4386(.din(new_new_n2792__), .dout(n16590));
  buf1  g4387(.din(new_new_n2356__), .dout(n16593));
  buf1  g4388(.din(new_new_n2796__), .dout(n16596));
  buf1  g4389(.din(new_new_n2798__), .dout(n16599));
  buf1  g4390(.din(new_new_n2800__), .dout(n16602));
  buf1  g4391(.din(new_new_n2358__), .dout(n16605));
  buf1  g4392(.din(new_new_n2804__), .dout(n16608));
  buf1  g4393(.din(new_new_n2806__), .dout(n16611));
  buf1  g4394(.din(new_new_n2808__), .dout(n16614));
  buf1  g4395(.din(new_new_n2360__), .dout(n16617));
  buf1  g4396(.din(new_new_n2812__), .dout(n16620));
  buf1  g4397(.din(new_new_n2814__), .dout(n16623));
  buf1  g4398(.din(new_new_n2816__), .dout(n16626));
  buf1  g4399(.din(new_new_n2362__), .dout(n16629));
  buf1  g4400(.din(new_new_n2820__), .dout(n16632));
  buf1  g4401(.din(new_new_n2822__), .dout(n16635));
  buf1  g4402(.din(new_new_n2824__), .dout(n16638));
  buf1  g4403(.din(new_new_n2364__), .dout(n16641));
  buf1  g4404(.din(new_new_n2828__), .dout(n16644));
  buf1  g4405(.din(new_new_n2830__), .dout(n16647));
  buf1  g4406(.din(new_new_n2832__), .dout(n16650));
  buf1  g4407(.din(new_new_n2366__), .dout(n16653));
  buf1  g4408(.din(new_new_n2836__), .dout(n16656));
  buf1  g4409(.din(new_new_n2838__), .dout(n16659));
  buf1  g4410(.din(new_new_n2840__), .dout(n16662));
  buf1  g4411(.din(new_new_n2368__), .dout(n16665));
  buf1  g4412(.din(new_new_n2844__), .dout(n16668));
  buf1  g4413(.din(new_new_n2846__), .dout(n16671));
  buf1  g4414(.din(new_new_n2848__), .dout(n16674));
  buf1  g4415(.din(new_new_n2370__), .dout(n16677));
  buf1  g4416(.din(new_new_n2852__), .dout(n16680));
  buf1  g4417(.din(new_new_n2854__), .dout(n16683));
  buf1  g4418(.din(new_new_n2856__), .dout(n16686));
  buf1  g4419(.din(new_new_n2372__), .dout(n16689));
  buf1  g4420(.din(new_new_n2860__), .dout(n16692));
  buf1  g4421(.din(new_new_n2862__), .dout(n16695));
  buf1  g4422(.din(new_new_n2864__), .dout(n16698));
  buf1  g4423(.din(new_new_n2374__), .dout(n16701));
  buf1  g4424(.din(new_new_n2868__), .dout(n16704));
  buf1  g4425(.din(new_new_n2870__), .dout(n16707));
  buf1  g4426(.din(new_new_n2872__), .dout(n16710));
  buf1  g4427(.din(new_new_n2376__), .dout(n16713));
  buf1  g4428(.din(new_new_n2876__), .dout(n16716));
  buf1  g4429(.din(new_new_n2878__), .dout(n16719));
  buf1  g4430(.din(new_new_n2880__), .dout(n16722));
  buf1  g4431(.din(new_new_n2378__), .dout(n16725));
  buf1  g4432(.din(new_new_n2884__), .dout(n16728));
  buf1  g4433(.din(new_new_n2886__), .dout(n16731));
  buf1  g4434(.din(new_new_n2888__), .dout(n16734));
  buf1  g4435(.din(new_new_n2380__), .dout(n16737));
  buf1  g4436(.din(new_new_n2892__), .dout(n16740));
  buf1  g4437(.din(new_new_n2894__), .dout(n16743));
  buf1  g4438(.din(new_new_n2896__), .dout(n16746));
  buf1  g4439(.din(new_new_n2382__), .dout(n16749));
  buf1  g4440(.din(new_new_n2900__), .dout(n16752));
  buf1  g4441(.din(new_new_n2902__), .dout(n16755));
  buf1  g4442(.din(new_new_n2904__), .dout(n16758));
  buf1  g4443(.din(new_new_n2384__), .dout(n16761));
  buf1  g4444(.din(new_new_n2908__), .dout(n16764));
  buf1  g4445(.din(new_new_n2910__), .dout(n16767));
  buf1  g4446(.din(new_new_n2912__), .dout(n16770));
  buf1  g4447(.din(new_new_n2386__), .dout(n16773));
  buf1  g4448(.din(new_new_n2916__), .dout(n16776));
  buf1  g4449(.din(new_new_n2918__), .dout(n16779));
  buf1  g4450(.din(new_new_n2920__), .dout(n16782));
  buf1  g4451(.din(new_new_n2388__), .dout(n16785));
  buf1  g4452(.din(new_new_n2924__), .dout(n16788));
  buf1  g4453(.din(new_new_n2926__), .dout(n16791));
  buf1  g4454(.din(new_new_n2928__), .dout(n16794));
  buf1  g4455(.din(new_new_n2390__), .dout(n16797));
  buf1  g4456(.din(new_new_n2932__), .dout(n16800));
  buf1  g4457(.din(new_new_n2934__), .dout(n16803));
  buf1  g4458(.din(new_new_n2936__), .dout(n16806));
  buf1  g4459(.din(new_new_n2392__), .dout(n16809));
  buf1  g4460(.din(new_new_n2940__), .dout(n16812));
  buf1  g4461(.din(new_new_n2942__), .dout(n16815));
  buf1  g4462(.din(new_new_n2944__), .dout(n16818));
  buf1  g4463(.din(new_new_n2394__), .dout(n16821));
  buf1  g4464(.din(new_new_n2948__), .dout(n16824));
  buf1  g4465(.din(new_new_n2950__), .dout(n16827));
  buf1  g4466(.din(new_new_n2952__), .dout(n16830));
  buf1  g4467(.din(new_new_n2396__), .dout(n16833));
  buf1  g4468(.din(new_new_n2956__), .dout(n16836));
  buf1  g4469(.din(new_new_n2958__), .dout(n16839));
  buf1  g4470(.din(new_new_n2960__), .dout(n16842));
  buf1  g4471(.din(new_new_n2398__), .dout(n16845));
  buf1  g4472(.din(new_new_n2964__), .dout(n16848));
  buf1  g4473(.din(new_new_n2966__), .dout(n16851));
  buf1  g4474(.din(new_new_n2968__), .dout(n16854));
  buf1  g4475(.din(new_new_n2400__), .dout(n16857));
  buf1  g4476(.din(new_new_n2972__), .dout(n16860));
  buf1  g4477(.din(new_new_n2974__), .dout(n16863));
  buf1  g4478(.din(new_new_n2976__), .dout(n16866));
  buf1  g4479(.din(new_new_n2402__), .dout(n16869));
  buf1  g4480(.din(new_new_n2980__), .dout(n16872));
  buf1  g4481(.din(new_new_n2982__), .dout(n16875));
  buf1  g4482(.din(new_new_n2984__), .dout(n16878));
  buf1  g4483(.din(new_new_n2404__), .dout(n16881));
  buf1  g4484(.din(new_new_n2988__), .dout(n16884));
  buf1  g4485(.din(new_new_n2990__), .dout(n16887));
  buf1  g4486(.din(new_new_n2992__), .dout(n16890));
  buf1  g4487(.din(new_new_n2406__), .dout(n16893));
  buf1  g4488(.din(new_new_n2996__), .dout(n16896));
  buf1  g4489(.din(new_new_n2998__), .dout(n16899));
  buf1  g4490(.din(new_new_n3000__), .dout(n16902));
  buf1  g4491(.din(new_new_n2408__), .dout(n16905));
  buf1  g4492(.din(new_new_n3004__), .dout(n16908));
  buf1  g4493(.din(new_new_n3006__), .dout(n16911));
  buf1  g4494(.din(new_new_n3008__), .dout(n16914));
  buf1  g4495(.din(new_new_n2410__), .dout(n16917));
  buf1  g4496(.din(new_new_n3012__), .dout(n16920));
  buf1  g4497(.din(new_new_n3014__), .dout(n16923));
  buf1  g4498(.din(new_new_n3016__), .dout(n16926));
  buf1  g4499(.din(new_new_n2412__), .dout(n16929));
  buf1  g4500(.din(new_new_n3020__), .dout(n16932));
  buf1  g4501(.din(new_new_n3022__), .dout(n16935));
  buf1  g4502(.din(new_new_n3024__), .dout(n16938));
  buf1  g4503(.din(new_new_n2414__), .dout(n16941));
  buf1  g4504(.din(new_new_n3028__), .dout(n16944));
  buf1  g4505(.din(new_new_n3030__), .dout(n16947));
  buf1  g4506(.din(new_new_n3032__), .dout(n16950));
  buf1  g4507(.din(new_new_n2416__), .dout(n16953));
  buf1  g4508(.din(new_new_n3036__), .dout(n16956));
  buf1  g4509(.din(new_new_n3038__), .dout(n16959));
  buf1  g4510(.din(new_new_n3040__), .dout(n16962));
  buf1  g4511(.din(new_new_n2418__), .dout(n16965));
  buf1  g4512(.din(new_new_n3044__), .dout(n16968));
  buf1  g4513(.din(new_new_n3046__), .dout(n16971));
  buf1  g4514(.din(new_new_n3048__), .dout(n16974));
  buf1  g4515(.din(new_new_n2420__), .dout(n16977));
  buf1  g4516(.din(new_new_n3052__), .dout(n16980));
  buf1  g4517(.din(new_new_n3054__), .dout(n16983));
  buf1  g4518(.din(new_new_n3056__), .dout(n16986));
  buf1  g4519(.din(new_new_n2422__), .dout(n16989));
  buf1  g4520(.din(new_new_n3060__), .dout(n16992));
  buf1  g4521(.din(new_new_n3062__), .dout(n16995));
  buf1  g4522(.din(new_new_n3064__), .dout(n16998));
  buf1  g4523(.din(new_new_n2424__), .dout(n17001));
  buf1  g4524(.din(new_new_n3068__), .dout(n17004));
  buf1  g4525(.din(new_new_n3070__), .dout(n17007));
  buf1  g4526(.din(new_new_n3072__), .dout(n17010));
  buf1  g4527(.din(new_new_n2426__), .dout(n17013));
  buf1  g4528(.din(new_new_n3076__), .dout(n17016));
  buf1  g4529(.din(new_new_n3078__), .dout(n17019));
  buf1  g4530(.din(new_new_n3080__), .dout(n17022));
  buf1  g4531(.din(new_new_n2428__), .dout(n17025));
  buf1  g4532(.din(new_new_n3084__), .dout(n17028));
  buf1  g4533(.din(new_new_n3086__), .dout(n17031));
  buf1  g4534(.din(new_new_n3088__), .dout(n17034));
  buf1  g4535(.din(new_new_n2430__), .dout(n17037));
  buf1  g4536(.din(new_new_n3092__), .dout(n17040));
  buf1  g4537(.din(new_new_n3094__), .dout(n17043));
  buf1  g4538(.din(new_new_n3096__), .dout(n17046));
  buf1  g4539(.din(new_new_n2432__), .dout(n17049));
  buf1  g4540(.din(new_new_n3100__), .dout(n17052));
  buf1  g4541(.din(new_new_n3102__), .dout(n17055));
  buf1  g4542(.din(new_new_n3104__), .dout(n17058));
  buf1  g4543(.din(new_new_n2434__), .dout(n17061));
  buf1  g4544(.din(new_new_n3108__), .dout(n17064));
  buf1  g4545(.din(new_new_n3110__), .dout(n17067));
  buf1  g4546(.din(new_new_n3112__), .dout(n17070));
  buf1  g4547(.din(new_new_n2436__), .dout(n17073));
  buf1  g4548(.din(new_new_n3116__), .dout(n17076));
  buf1  g4549(.din(new_new_n3118__), .dout(n17079));
  buf1  g4550(.din(new_new_n3120__), .dout(n17082));
  buf1  g4551(.din(new_new_n2438__), .dout(n17085));
  buf1  g4552(.din(new_new_n3124__), .dout(n17088));
  buf1  g4553(.din(new_new_n3126__), .dout(n17091));
  buf1  g4554(.din(new_new_n3128__), .dout(n17094));
  buf1  g4555(.din(new_new_n2440__), .dout(n17097));
  buf1  g4556(.din(new_new_n3132__), .dout(n17100));
  buf1  g4557(.din(new_new_n3134__), .dout(n17103));
  buf1  g4558(.din(new_new_n3136__), .dout(n17106));
  buf1  g4559(.din(new_new_n2442__), .dout(n17109));
  buf1  g4560(.din(new_new_n3140__), .dout(n17112));
  buf1  g4561(.din(new_new_n3142__), .dout(n17115));
  buf1  g4562(.din(new_new_n3144__), .dout(n17118));
  buf1  g4563(.din(new_new_n2444__), .dout(n17121));
  buf1  g4564(.din(new_new_n3148__), .dout(n17124));
  buf1  g4565(.din(new_new_n3150__), .dout(n17127));
  buf1  g4566(.din(new_new_n3152__), .dout(n17130));
  buf1  g4567(.din(new_new_n2446__), .dout(n17133));
  buf1  g4568(.din(new_new_n3156__), .dout(n17136));
  buf1  g4569(.din(new_new_n3158__), .dout(n17139));
  buf1  g4570(.din(new_new_n3160__), .dout(n17142));
  buf1  g4571(.din(new_new_n2448__), .dout(n17145));
  buf1  g4572(.din(new_new_n3164__), .dout(n17148));
  buf1  g4573(.din(new_new_n3166__), .dout(n17151));
  buf1  g4574(.din(new_new_n3168__), .dout(n17154));
  buf1  g4575(.din(new_new_n2450__), .dout(n17157));
  buf1  g4576(.din(new_new_n3172__), .dout(n17160));
  buf1  g4577(.din(new_new_n3174__), .dout(n17163));
  buf1  g4578(.din(new_new_n3176__), .dout(n17166));
  buf1  g4579(.din(new_new_n2452__), .dout(n17169));
  buf1  g4580(.din(new_new_n3180__), .dout(n17172));
  buf1  g4581(.din(new_new_n3182__), .dout(n17175));
  buf1  g4582(.din(new_new_n3184__), .dout(n17178));
  buf1  g4583(.din(new_new_n2454__), .dout(n17181));
  buf1  g4584(.din(new_new_n3188__), .dout(n17184));
  buf1  g4585(.din(new_new_n3190__), .dout(n17187));
  buf1  g4586(.din(new_new_n3192__), .dout(n17190));
  buf1  g4587(.din(new_new_n2456__), .dout(n17193));
  buf1  g4588(.din(new_new_n3196__), .dout(n17196));
  buf1  g4589(.din(new_new_n3198__), .dout(n17199));
  buf1  g4590(.din(new_new_n3200__), .dout(n17202));
  buf1  g4591(.din(new_new_n2458__), .dout(n17205));
  buf1  g4592(.din(new_new_n3204__), .dout(n17208));
  buf1  g4593(.din(new_new_n3206__), .dout(n17211));
  buf1  g4594(.din(new_new_n3208__), .dout(n17214));
  buf1  g4595(.din(new_new_n2460__), .dout(n17217));
  buf1  g4596(.din(new_new_n3212__), .dout(n17220));
  buf1  g4597(.din(new_new_n3214__), .dout(n17223));
  buf1  g4598(.din(new_new_n3216__), .dout(n17226));
  buf1  g4599(.din(new_new_n2462__), .dout(n17229));
  buf1  g4600(.din(new_new_n3220__), .dout(n17232));
  buf1  g4601(.din(new_new_n3222__), .dout(n17235));
  buf1  g4602(.din(new_new_n3224__), .dout(n17238));
  buf1  g4603(.din(new_new_n2464__), .dout(n17241));
  buf1  g4604(.din(new_new_n3228__), .dout(n17244));
  buf1  g4605(.din(new_new_n3230__), .dout(n17247));
  buf1  g4606(.din(new_new_n3232__), .dout(n17250));
  buf1  g4607(.din(new_new_n2466__), .dout(n17253));
  buf1  g4608(.din(new_new_n3236__), .dout(n17256));
  buf1  g4609(.din(new_new_n3238__), .dout(n17259));
  buf1  g4610(.din(new_new_n3240__), .dout(n17262));
  buf1  g4611(.din(new_new_n2468__), .dout(n17265));
  buf1  g4612(.din(new_new_n3244__), .dout(n17268));
  buf1  g4613(.din(new_new_n3246__), .dout(n17271));
  buf1  g4614(.din(new_new_n3248__), .dout(n17274));
  buf1  g4615(.din(new_new_n2470__), .dout(n17277));
  buf1  g4616(.din(new_new_n3252__), .dout(n17280));
  buf1  g4617(.din(new_new_n3254__), .dout(n17283));
  buf1  g4618(.din(new_new_n3256__), .dout(n17286));
  buf1  g4619(.din(new_new_n2472__), .dout(n17289));
  buf1  g4620(.din(new_new_n3260__), .dout(n17292));
  buf1  g4621(.din(new_new_n3262__), .dout(n17295));
  buf1  g4622(.din(new_new_n3264__), .dout(n17298));
  buf1  g4623(.din(new_new_n2474__), .dout(n17301));
  buf1  g4624(.din(new_new_n3268__), .dout(n17304));
  buf1  g4625(.din(new_new_n3270__), .dout(n17307));
  buf1  g4626(.din(new_new_n3272__), .dout(n17310));
  buf1  g4627(.din(new_new_n2476__), .dout(n17313));
  buf1  g4628(.din(new_new_n3276__), .dout(n17316));
  buf1  g4629(.din(new_new_n3278__), .dout(n17319));
  buf1  g4630(.din(new_new_n3280__), .dout(n17322));
  buf1  g4631(.din(new_new_n2478__), .dout(n17325));
  buf1  g4632(.din(new_new_n3284__), .dout(n17328));
  buf1  g4633(.din(new_new_n3286__), .dout(n17331));
  buf1  g4634(.din(new_new_n3288__), .dout(n17334));
  buf1  g4635(.din(new_new_n2480__), .dout(n17337));
  buf1  g4636(.din(new_new_n3292__), .dout(n17340));
  buf1  g4637(.din(new_new_n3294__), .dout(n17343));
  buf1  g4638(.din(new_new_n3296__), .dout(n17346));
  buf1  g4639(.din(new_new_n2482__), .dout(n17349));
  buf1  g4640(.din(new_new_n3300__), .dout(n17352));
  buf1  g4641(.din(new_new_n3302__), .dout(n17355));
  buf1  g4642(.din(new_new_n3304__), .dout(n17358));
  buf1  g4643(.din(new_new_n2484__), .dout(n17361));
  buf1  g4644(.din(new_new_n3308__), .dout(n17364));
  buf1  g4645(.din(new_new_n3310__), .dout(n17367));
  buf1  g4646(.din(new_new_n3312__), .dout(n17370));
  buf1  g4647(.din(new_new_n2486__), .dout(n17373));
  buf1  g4648(.din(new_new_n3316__), .dout(n17376));
  buf1  g4649(.din(new_new_n3318__), .dout(n17379));
  buf1  g4650(.din(new_new_n3320__), .dout(n17382));
  buf1  g4651(.din(new_new_n2488__), .dout(n17385));
  buf1  g4652(.din(new_new_n3324__), .dout(n17388));
  buf1  g4653(.din(new_new_n3326__), .dout(n17391));
  buf1  g4654(.din(new_new_n3328__), .dout(n17394));
  buf1  g4655(.din(new_new_n2490__), .dout(n17397));
  buf1  g4656(.din(new_new_n3332__), .dout(n17400));
  buf1  g4657(.din(new_new_n3334__), .dout(n17403));
  buf1  g4658(.din(new_new_n3336__), .dout(n17406));
  buf1  g4659(.din(new_new_n2492__), .dout(n17409));
  buf1  g4660(.din(new_new_n3340__), .dout(n17412));
  buf1  g4661(.din(new_new_n3342__), .dout(n17415));
  buf1  g4662(.din(new_new_n3344__), .dout(n17418));
  buf1  g4663(.din(new_new_n2494__), .dout(n17421));
  buf1  g4664(.din(new_new_n3348__), .dout(n17424));
  buf1  g4665(.din(new_new_n3350__), .dout(n17427));
  buf1  g4666(.din(new_new_n3352__), .dout(n17430));
  buf1  g4667(.din(new_new_n2496__), .dout(n17433));
  buf1  g4668(.din(new_new_n3356__), .dout(n17436));
  buf1  g4669(.din(new_new_n3358__), .dout(n17439));
  buf1  g4670(.din(new_new_n3360__), .dout(n17442));
  buf1  g4671(.din(new_new_n2498__), .dout(n17445));
  buf1  g4672(.din(new_new_n3364__), .dout(n17448));
  buf1  g4673(.din(new_new_n3366__), .dout(n17451));
  buf1  g4674(.din(new_new_n3368__), .dout(n17454));
  buf1  g4675(.din(new_new_n2500__), .dout(n17457));
  buf1  g4676(.din(new_new_n3372__), .dout(n17460));
  buf1  g4677(.din(new_new_n3374__), .dout(n17463));
  buf1  g4678(.din(new_new_n3376__), .dout(n17466));
  buf1  g4679(.din(new_new_n2502__), .dout(n17469));
  buf1  g4680(.din(new_new_n3380__), .dout(n17472));
  buf1  g4681(.din(new_new_n2504__), .dout(n17475));
  buf1  g4682(.din(new_new_n3384__), .dout(n17478));
  buf1  g4683(.din(new_new_n2506__), .dout(n17481));
  buf1  g4684(.din(new_new_n10128__), .dout(n17484));
  buf1  g4685(.din(new_new_n2508__), .dout(n17487));
  buf1  g4686(.din(new_new_n2510__), .dout(n17490));
  buf1  g4687(.din(new_new_n10117__), .dout(n17493));
  buf1  g4688(.din(new_new_n2512__), .dout(n17496));
  buf1  g4689(.din(new_new_n2514__), .dout(n17499));
  buf1  g4690(.din(new_new_n10095__), .dout(n17502));
  buf1  g4691(.din(new_new_n2516__), .dout(n17505));
  buf1  g4692(.din(new_new_n2518__), .dout(n17508));
  buf1  g4693(.din(new_new_n3406__), .dout(n17511));
  buf1  g4694(.din(new_new_n10033__), .dout(n17514));
  buf1  g4695(.din(new_new_n2520__), .dout(n17517));
  buf1  g4696(.din(new_new_n3412__), .dout(n17520));
  buf1  g4697(.din(new_new_n2522__), .dout(n17523));
  buf1  g4698(.din(new_new_n3416__), .dout(n17526));
  buf1  g4699(.din(new_new_n2524__), .dout(n17529));
  buf1  g4700(.din(new_new_n3420__), .dout(n17532));
  buf1  g4701(.din(new_new_n3422__), .dout(n17535));
  buf1  g4702(.din(new_new_n3424__), .dout(n17538));
  buf1  g4703(.din(new_new_n2526__), .dout(n17541));
  buf1  g4704(.din(new_new_n3428__), .dout(n17544));
  buf1  g4705(.din(new_new_n2528__), .dout(n17547));
  buf1  g4706(.din(new_new_n3432__), .dout(n17550));
  buf1  g4707(.din(new_new_n2530__), .dout(n17553));
  buf1  g4708(.din(new_new_n3436__), .dout(n17556));
  buf1  g4709(.din(new_new_n2532__), .dout(n17559));
  buf1  g4710(.din(new_new_n10034__), .dout(n17562));
  buf1  g4711(.din(new_new_n2534__), .dout(n17565));
  buf1  g4712(.din(new_new_n9977__), .dout(n17568));
  buf1  g4713(.din(new_new_n9976__), .dout(n17571));
  buf1  g4714(.din(new_new_n9987__), .dout(n17574));
  buf1  g4715(.din(new_new_n2548__), .dout(n17577));
  buf1  g4716(.din(new_new_n3452__), .dout(n17580));
  buf1  g4717(.din(new_new_n3454__), .dout(n17583));
  buf1  g4718(.din(new_new_n2550__), .dout(n17586));
  buf1  g4719(.din(new_new_n3458__), .dout(n17589));
  buf1  g4720(.din(new_new_n3460__), .dout(n17592));
  buf1  g4721(.din(new_new_n2552__), .dout(n17595));
  buf1  g4722(.din(new_new_n3464__), .dout(n17598));
  buf1  g4723(.din(new_new_n10161__), .dout(n17601));
  buf1  g4724(.din(new_new_n2554__), .dout(n17604));
  buf1  g4725(.din(new_new_n3470__), .dout(n17607));
  buf1  g4726(.din(new_new_n4244__), .dout(n17610));
  buf1  g4727(.din(new_new_n2556__), .dout(n17613));
  buf1  g4728(.din(new_new_n10156__), .dout(n17616));
  buf1  g4729(.din(new_new_n2558__), .dout(n17619));
  buf1  g4730(.din(new_new_n2560__), .dout(n17622));
  buf1  g4731(.din(new_new_n10147__), .dout(n17625));
  buf1  g4732(.din(new_new_n2562__), .dout(n17628));
  buf1  g4733(.din(new_new_n2564__), .dout(n17631));
  buf1  g4734(.din(new_new_n10140__), .dout(n17634));
  buf1  g4735(.din(new_new_n2566__), .dout(n17637));
  buf1  g4736(.din(new_new_n2568__), .dout(n17640));
  buf1  g4737(.din(new_new_n3494__), .dout(n17643));
  buf1  g4738(.din(new_new_n10518__), .dout(n17646));
  buf1  g4739(.din(new_new_n2570__), .dout(n17649));
  buf1  g4740(.din(new_new_n3500__), .dout(n17652));
  buf1  g4741(.din(new_new_n2576__), .dout(n17655));
  buf1  g4742(.din(new_new_n3932__), .dout(n17658));
  buf1  g4743(.din(new_new_n9990__), .dout(n17661));
  buf1  g4744(.din(new_new_n3874__), .dout(n17664));
  buf1  g4745(.din(new_new_n9989__), .dout(n17667));
  buf1  g4746(.din(new_new_n3878__), .dout(n17670));
  buf1  g4747(.din(new_new_n9696__), .dout(n17673));
  buf1  g4748(.din(new_new_n3914__), .dout(n17676));
  buf1  g4749(.din(new_new_n2590__), .dout(n17679));
  buf1  g4750(.din(new_new_n3520__), .dout(n17682));
  buf1  g4751(.din(new_new_n3522__), .dout(n17685));
  buf1  g4752(.din(new_new_n2592__), .dout(n17688));
  buf1  g4753(.din(new_new_n3526__), .dout(n17691));
  buf1  g4754(.din(new_new_n3528__), .dout(n17694));
  buf1  g4755(.din(new_new_n2594__), .dout(n17697));
  buf1  g4756(.din(new_new_n3532__), .dout(n17700));
  buf1  g4757(.din(new_new_n3534__), .dout(n17703));
  buf1  g4758(.din(new_new_n3536__), .dout(n17706));
  buf1  g4759(.din(new_new_n9933__), .dout(n17709));
  buf1  g4760(.din(new_new_n2598__), .dout(n17712));
  buf1  g4761(.din(new_new_n3542__), .dout(n17715));
  buf1  g4762(.din(new_new_n3544__), .dout(n17718));
  buf1  g4763(.din(new_new_n3546__), .dout(n17721));
  buf1  g4764(.din(new_new_n2600__), .dout(n17724));
  buf1  g4765(.din(new_new_n9939__), .dout(n17727));
  buf1  g4766(.din(new_new_n9947__), .dout(n17730));
  buf1  g4767(.din(new_new_n9955__), .dout(n17733));
  buf1  g4768(.din(new_new_n2606__), .dout(n17736));
  buf1  g4769(.din(new_new_n9728__), .dout(n17739));
  buf1  g4770(.din(new_new_n2608__), .dout(n17742));
  buf1  g4771(.din(new_new_n3562__), .dout(n17745));
  buf1  g4772(.din(new_new_n9677__), .dout(n17748));
  buf1  g4773(.din(new_new_n2610__), .dout(n17751));
  buf1  g4774(.din(new_new_n3568__), .dout(n17754));
  buf1  g4775(.din(new_new_n9553__), .dout(n17757));
  buf1  g4776(.din(new_new_n2612__), .dout(n17760));
  buf1  g4777(.din(new_new_n9763__), .dout(n17763));
  buf1  g4778(.din(new_new_n2614__), .dout(n17766));
  buf1  g4779(.din(new_new_n9736__), .dout(n17769));
  buf1  g4780(.din(new_new_n2616__), .dout(n17772));
  buf1  g4781(.din(new_new_n9775__), .dout(n17775));
  buf1  g4782(.din(new_new_n2618__), .dout(n17778));
  buf1  g4783(.din(new_new_n9911__), .dout(n17781));
  buf1  g4784(.din(new_new_n2620__), .dout(n17784));
  buf1  g4785(.din(new_new_n3590__), .dout(n17787));
  buf1  g4786(.din(new_new_n9687__), .dout(n17790));
  buf1  g4787(.din(new_new_n2622__), .dout(n17793));
  buf1  g4788(.din(new_new_n9961__), .dout(n17796));
  buf1  g4789(.din(new_new_n9968__), .dout(n17799));
  buf1  g4790(.din(new_new_n9975__), .dout(n17802));
  buf1  g4791(.din(new_new_n2628__), .dout(n17805));
  buf1  g4792(.din(new_new_n3604__), .dout(n17808));
  buf1  g4793(.din(new_new_n3606__), .dout(n17811));
  buf1  g4794(.din(new_new_n3608__), .dout(n17814));
  buf1  g4795(.din(new_new_n2630__), .dout(n17817));
  buf1  g4796(.din(new_new_n3612__), .dout(n17820));
  buf1  g4797(.din(new_new_n3614__), .dout(n17823));
  buf1  g4798(.din(new_new_n3616__), .dout(n17826));
  buf1  g4799(.din(new_new_n2632__), .dout(n17829));
  buf1  g4800(.din(new_new_n3620__), .dout(n17832));
  buf1  g4801(.din(new_new_n3622__), .dout(n17835));
  buf1  g4802(.din(new_new_n3624__), .dout(n17838));
  buf1  g4803(.din(new_new_n2634__), .dout(n17841));
  buf1  g4804(.din(new_new_n3628__), .dout(n17844));
  buf1  g4805(.din(new_new_n3630__), .dout(n17847));
  buf1  g4806(.din(new_new_n3632__), .dout(n17850));
  buf1  g4807(.din(new_new_n2636__), .dout(n17853));
  buf1  g4808(.din(new_new_n3636__), .dout(n17856));
  buf1  g4809(.din(new_new_n3638__), .dout(n17859));
  buf1  g4810(.din(new_new_n3640__), .dout(n17862));
  buf1  g4811(.din(new_new_n2638__), .dout(n17865));
  buf1  g4812(.din(new_new_n3644__), .dout(n17868));
  buf1  g4813(.din(new_new_n3646__), .dout(n17871));
  buf1  g4814(.din(new_new_n3648__), .dout(n17874));
  buf1  g4815(.din(new_new_n2640__), .dout(n17877));
  buf1  g4816(.din(new_new_n3652__), .dout(n17880));
  buf1  g4817(.din(new_new_n3654__), .dout(n17883));
  buf1  g4818(.din(new_new_n2642__), .dout(n17886));
  buf1  g4819(.din(new_new_n3658__), .dout(n17889));
  buf1  g4820(.din(new_new_n3660__), .dout(n17892));
  buf1  g4821(.din(new_new_n3662__), .dout(n17895));
  buf1  g4822(.din(new_new_n2644__), .dout(n17898));
  buf1  g4823(.din(new_new_n3666__), .dout(n17901));
  buf1  g4824(.din(new_new_n3668__), .dout(n17904));
  buf1  g4825(.din(new_new_n3670__), .dout(n17907));
  buf1  g4826(.din(new_new_n2646__), .dout(n17910));
  buf1  g4827(.din(new_new_n3674__), .dout(n17913));
  buf1  g4828(.din(new_new_n3676__), .dout(n17916));
  buf1  g4829(.din(new_new_n3678__), .dout(n17919));
  buf1  g4830(.din(new_new_n2648__), .dout(n17922));
  buf1  g4831(.din(new_new_n3682__), .dout(n17925));
  buf1  g4832(.din(new_new_n3684__), .dout(n17928));
  buf1  g4833(.din(new_new_n3686__), .dout(n17931));
  buf1  g4834(.din(new_new_n2650__), .dout(n17934));
  buf1  g4835(.din(new_new_n3690__), .dout(n17937));
  buf1  g4836(.din(new_new_n3692__), .dout(n17940));
  buf1  g4837(.din(new_new_n2652__), .dout(n17943));
  buf1  g4838(.din(new_new_n3696__), .dout(n17946));
  buf1  g4839(.din(new_new_n3698__), .dout(n17949));
  buf1  g4840(.din(new_new_n3700__), .dout(n17952));
  buf1  g4841(.din(new_new_n2654__), .dout(n17955));
  buf1  g4842(.din(new_new_n3704__), .dout(n17958));
  buf1  g4843(.din(new_new_n3706__), .dout(n17961));
  buf1  g4844(.din(new_new_n3708__), .dout(n17964));
  buf1  g4845(.din(new_new_n2656__), .dout(n17967));
  buf1  g4846(.din(new_new_n3712__), .dout(n17970));
  buf1  g4847(.din(new_new_n3714__), .dout(n17973));
  buf1  g4848(.din(new_new_n3716__), .dout(n17976));
  buf1  g4849(.din(new_new_n2658__), .dout(n17979));
  buf1  g4850(.din(new_new_n3720__), .dout(n17982));
  buf1  g4851(.din(new_new_n3722__), .dout(n17985));
  buf1  g4852(.din(new_new_n3724__), .dout(n17988));
  buf1  g4853(.din(new_new_n2660__), .dout(n17991));
  buf1  g4854(.din(new_new_n3728__), .dout(n17994));
  buf1  g4855(.din(new_new_n3730__), .dout(n17997));
  buf1  g4856(.din(new_new_n3732__), .dout(n18000));
  buf1  g4857(.din(new_new_n2662__), .dout(n18003));
  buf1  g4858(.din(new_new_n3736__), .dout(n18006));
  buf1  g4859(.din(new_new_n3738__), .dout(n18009));
  buf1  g4860(.din(new_new_n3740__), .dout(n18012));
  buf1  g4861(.din(new_new_n2664__), .dout(n18015));
  buf1  g4862(.din(new_new_n3744__), .dout(n18018));
  buf1  g4863(.din(new_new_n3746__), .dout(n18021));
  buf1  g4864(.din(new_new_n3748__), .dout(n18024));
  buf1  g4865(.din(new_new_n2666__), .dout(n18027));
  buf1  g4866(.din(new_new_n3752__), .dout(n18030));
  buf1  g4867(.din(new_new_n3754__), .dout(n18033));
  buf1  g4868(.din(new_new_n3756__), .dout(n18036));
  buf1  g4869(.din(new_new_n2668__), .dout(n18039));
  buf1  g4870(.din(new_new_n3760__), .dout(n18042));
  buf1  g4871(.din(new_new_n3762__), .dout(n18045));
  buf1  g4872(.din(new_new_n3764__), .dout(n18048));
  buf1  g4873(.din(new_new_n2670__), .dout(n18051));
  buf1  g4874(.din(new_new_n3768__), .dout(n18054));
  buf1  g4875(.din(new_new_n3770__), .dout(n18057));
  buf1  g4876(.din(new_new_n3772__), .dout(n18060));
  buf1  g4877(.din(new_new_n2672__), .dout(n18063));
  buf1  g4878(.din(new_new_n3776__), .dout(n18066));
  buf1  g4879(.din(new_new_n3778__), .dout(n18069));
  buf1  g4880(.din(new_new_n3780__), .dout(n18072));
  buf1  g4881(.din(new_new_n2674__), .dout(n18075));
  buf1  g4882(.din(new_new_n3784__), .dout(n18078));
  buf1  g4883(.din(new_new_n3786__), .dout(n18081));
  buf1  g4884(.din(new_new_n3788__), .dout(n18084));
  buf1  g4885(.din(new_new_n2676__), .dout(n18087));
  buf1  g4886(.din(new_new_n3792__), .dout(n18090));
  buf1  g4887(.din(new_new_n3794__), .dout(n18093));
  buf1  g4888(.din(new_new_n3796__), .dout(n18096));
  buf1  g4889(.din(new_new_n2678__), .dout(n18099));
  buf1  g4890(.din(new_new_n3800__), .dout(n18102));
  buf1  g4891(.din(new_new_n3802__), .dout(n18105));
  buf1  g4892(.din(new_new_n3804__), .dout(n18108));
  buf1  g4893(.din(new_new_n2680__), .dout(n18111));
  buf1  g4894(.din(new_new_n3808__), .dout(n18114));
  buf1  g4895(.din(new_new_n3810__), .dout(n18117));
  buf1  g4896(.din(new_new_n3812__), .dout(n18120));
  buf1  g4897(.din(new_new_n2682__), .dout(n18123));
  buf1  g4898(.din(new_new_n3816__), .dout(n18126));
  buf1  g4899(.din(new_new_n3818__), .dout(n18129));
  buf1  g4900(.din(new_new_n3820__), .dout(n18132));
  buf1  g4901(.din(new_new_n3996__), .dout(n18135));
  buf1  g4902(.din(new_new_n3998__), .dout(n18138));
  buf1  g4903(.din(new_new_n4008__), .dout(n18141));
  buf1  g4904(.din(new_new_n4010__), .dout(n18144));
  buf1  g4905(.din(new_new_n4018__), .dout(n18147));
  buf1  g4906(.din(new_new_n4020__), .dout(n18150));
  buf1  g4907(.din(new_new_n4024__), .dout(n18153));
  buf1  g4908(.din(new_new_n4026__), .dout(n18156));
  buf1  g4909(.din(new_new_n9845__), .dout(n18159));
  buf1  g4910(.din(new_new_n9878__), .dout(n18162));
  buf1  g4911(.din(new_new_n4060__), .dout(n18165));
  buf1  g4912(.din(new_new_n4062__), .dout(n18168));
  buf1  g4913(.din(new_new_n9674__), .dout(n18171));
  buf1  g4914(.din(new_new_n9684__), .dout(n18174));
  buf1  g4915(.din(new_new_n9901__), .dout(n18177));
  buf1  g4916(.din(new_new_n10520__), .dout(n18180));
  buf1  g4917(.din(new_new_n4032__), .dout(n18183));
  buf1  g4918(.din(new_new_n4034__), .dout(n18186));
  buf1  g4919(.din(new_new_n10063__), .dout(n18189));
  buf1  g4920(.din(new_new_n9561__), .dout(n18192));
  buf1  g4921(.din(new_new_n10076__), .dout(n18195));
  buf1  g4922(.din(new_new_n9577__), .dout(n18198));
  buf1  g4923(.din(new_new_n10522__), .dout(n18201));
  buf1  g4924(.din(new_new_n10525__), .dout(n18204));
  buf1  g4925(.din(new_new_n10528__), .dout(n18207));
  buf1  g4926(.din(new_new_n4050__), .dout(n18210));
  buf1  g4927(.din(new_new_n10531__), .dout(n18213));
  buf1  g4928(.din(new_new_n4054__), .dout(n18216));
  buf1  g4929(.din(new_new_n4056__), .dout(n18219));
  buf1  g4930(.din(new_new_n4058__), .dout(n18222));
  buf1  g4931(.din(new_new_n4064__), .dout(n18225));
  buf1  g4932(.din(new_new_n10093__), .dout(n18228));
  buf1  g4933(.din(new_new_n9593__), .dout(n18231));
  buf1  g4934(.din(new_new_n9607__), .dout(n18234));
  buf1  g4935(.din(new_new_n10112__), .dout(n18237));
  buf1  g4936(.din(new_new_n4066__), .dout(n18240));
  buf1  g4937(.din(new_new_n4068__), .dout(n18243));
  buf1  g4938(.din(new_new_n4070__), .dout(n18246));
  buf1  g4939(.din(new_new_n4072__), .dout(n18249));
  buf1  g4940(.din(new_new_n9870__), .dout(n18252));
  buf1  g4941(.din(new_new_n4074__), .dout(n18255));
  buf1  g4942(.din(new_new_n4076__), .dout(n18258));
  buf1  g4943(.din(new_new_n4078__), .dout(n18261));
  buf1  g4944(.din(new_new_n4080__), .dout(n18264));
  buf1  g4945(.din(new_new_n4090__), .dout(n18267));
  buf1  g4946(.din(new_new_n4092__), .dout(n18270));
  buf1  g4947(.din(new_new_n4094__), .dout(n18273));
  buf1  g4948(.din(new_new_n4096__), .dout(n18276));
  buf1  g4949(.din(new_new_n9844__), .dout(n18279));
  buf1  g4950(.din(n18252), .dout(n18282));
  buf1  g4951(.din(new_new_n4102__), .dout(n18285));
  buf1  g4952(.din(new_new_n10533__), .dout(n18288));
  buf1  g4953(.din(new_new_n10366__), .dout(n18291));
  buf1  g4954(.din(new_new_n10534__), .dout(n18294));
  buf1  g4955(.din(new_new_n4132__), .dout(n18297));
  buf1  g4956(.din(new_new_n4114__), .dout(n18300));
  buf1  g4957(.din(new_new_n4116__), .dout(n18303));
  buf1  g4958(.din(new_new_n4124__), .dout(n18306));
  buf1  g4959(.din(new_new_n4138__), .dout(n18309));
  buf1  g4960(.din(new_new_n10227__), .dout(n18312));
  buf1  g4961(.din(new_new_n4142__), .dout(n18315));
  buf1  g4962(.din(new_new_n10244__), .dout(n18318));
  buf1  g4963(.din(new_new_n4146__), .dout(n18321));
  buf1  g4964(.din(new_new_n10535__), .dout(n18324));
  buf1  g4965(.din(new_new_n10536__), .dout(n18327));
  buf1  g4966(.din(new_new_n4148__), .dout(n18330));
  buf1  g4967(.din(new_new_n4150__), .dout(n18333));
  buf1  g4968(.din(new_new_n10226__), .dout(n18336));
  buf1  g4969(.din(new_new_n10359__), .dout(n18339));
  buf1  g4970(.din(new_new_n4162__), .dout(n18342));
  buf1  g4971(.din(new_new_n4164__), .dout(n18345));
  buf1  g4972(.din(new_new_n4166__), .dout(n18348));
  buf1  g4973(.din(new_new_n4158__), .dout(n18351));
  buf1  g4974(.din(new_new_n4168__), .dout(n18354));
  buf1  g4975(.din(new_new_n4170__), .dout(n18357));
  buf1  g4976(.din(new_new_n4172__), .dout(n18360));
  buf1  g4977(.din(new_new_n10280__), .dout(n18363));
  buf1  g4978(.din(new_new_n10327__), .dout(n18366));
  buf1  g4979(.din(new_new_n10326__), .dout(n18369));
  buf1  g4980(.din(new_new_n10279__), .dout(n18372));
  buf1  g4981(.din(new_new_n10537__), .dout(n18375));
  buf1  g4982(.din(new_new_n10239__), .dout(n18378));
  buf1  g4983(.din(new_new_n10134__), .dout(n18381));
  buf1  g4984(.din(new_new_n9698__), .dout(n18384));
  buf1  g4985(.din(new_new_n9857__), .dout(n18387));
  buf1  g4986(.din(new_new_n9890__), .dout(n18390));
  buf1  g4987(.din(new_new_n10261__), .dout(n18393));
  buf1  g4988(.din(new_new_n10309__), .dout(n18396));
  buf1  g4989(.din(new_new_n9849__), .dout(n18399));
  buf1  g4990(.din(new_new_n9888__), .dout(n18402));
  buf1  g4991(.din(new_new_n9697__), .dout(n18405));
  buf1  g4992(.din(new_new_n4486__), .dout(n18408));
  buf1  g4993(.din(new_new_n10256__), .dout(n18411));
  buf1  g4994(.din(new_new_n10304__), .dout(n18414));
  buf1  g4995(.din(new_new_n4484__), .dout(n18417));
  buf1  g4996(.din(new_new_n4568__), .dout(n18420));
  buf1  g4997(.din(new_new_n10213__), .dout(n18423));
  buf1  g4998(.din(new_new_n10250__), .dout(n18426));
  buf1  g4999(.din(new_new_n10294__), .dout(n18429));
  buf1  g5000(.din(new_new_n10230__), .dout(n18432));
  buf1  g5001(.din(new_new_n10267__), .dout(n18435));
  buf1  g5002(.din(new_new_n10315__), .dout(n18438));
  buf1  g5003(.din(new_new_n10201__), .dout(n18441));
  buf1  g5004(.din(new_new_n10300__), .dout(n18444));
  buf1  g5005(.din(new_new_n9719__), .dout(n18447));
  buf1  g5006(.din(new_new_n9813__), .dout(n18450));
  buf1  g5007(.din(new_new_n9708__), .dout(n18453));
  buf1  g5008(.din(new_new_n9701__), .dout(n18456));
  buf1  g5009(.din(new_new_n10249__), .dout(n18459));
  buf1  g5010(.din(n18444), .dout(n18462));
  buf1  g5011(.din(new_new_n4492__), .dout(n18465));
  buf1  g5012(.din(new_new_n4494__), .dout(n18468));
  buf1  g5013(.din(new_new_n4496__), .dout(n18471));
  buf1  g5014(.din(new_new_n4498__), .dout(n18474));
  buf1  g5015(.din(new_new_n4500__), .dout(n18477));
  buf1  g5016(.din(new_new_n4502__), .dout(n18480));
  buf1  g5017(.din(new_new_n9714__), .dout(n18483));
  buf1  g5018(.din(new_new_n9811__), .dout(n18486));
  buf1  g5019(.din(new_new_n10270__), .dout(n18489));
  buf1  g5020(.din(new_new_n10299__), .dout(n18492));
  buf1  g5021(.din(new_new_n4620__), .dout(n18495));
  buf1  g5022(.din(new_new_n9806__), .dout(n18498));
  buf1  g5023(.din(new_new_n9749__), .dout(n18501));
  buf1  g5024(.din(new_new_n9808__), .dout(n18504));
  buf1  g5025(.din(new_new_n9751__), .dout(n18507));
  buf1  g5026(.din(new_new_n9809__), .dout(n18510));
  buf1  g5027(.din(new_new_n9752__), .dout(n18513));
  buf1  g5028(.din(new_new_n9807__), .dout(n18516));
  buf1  g5029(.din(new_new_n9750__), .dout(n18519));
  buf1  g5030(.din(new_new_n9918__), .dout(n18522));
  buf1  g5031(.din(new_new_n9922__), .dout(n18525));
  buf1  g5032(.din(new_new_n9923__), .dout(n18528));
  buf1  g5033(.din(new_new_n9919__), .dout(n18531));
  buf1  g5034(.din(new_new_n9713__), .dout(n18534));
  buf1  g5035(.din(new_new_n9717__), .dout(n18537));
  buf1  g5036(.din(new_new_n9779__), .dout(n18540));
  buf1  g5037(.din(new_new_n9783__), .dout(n18543));
  buf1  g5038(.din(new_new_n9819__), .dout(n18546));
  buf1  g5039(.din(new_new_n9830__), .dout(n18549));
  buf1  g5040(.din(new_new_n10451__), .dout(n18552));
  buf1  g5041(.din(new_new_n9995__), .dout(n18555));
  buf1  g5042(.din(new_new_n10002__), .dout(n18558));
  not1  g5043(.din(new_new_n10004__), .dout(n18561));
  not1  g5044(.din(new_new_n10013__), .dout(n18564));
  buf1  g5045(.din(new_new_n10009__), .dout(n18567));
  buf1  g5046(.din(new_new_n10398__), .dout(n18570));
  buf1  g5047(.din(new_new_n10410__), .dout(n18573));
  buf1  g5048(.din(new_new_n10001__), .dout(n18576));
  buf1  g5049(.din(new_new_n9994__), .dout(n18579));
  buf1  g5050(.din(new_new_n10024__), .dout(n18582));
  buf1  g5051(.din(new_new_n10429__), .dout(n18585));
  buf1  g5052(.din(new_new_n9831__), .dout(n18588));
  buf1  g5053(.din(new_new_n9812__), .dout(n18591));
  buf1  g5054(.din(new_new_n9820__), .dout(n18594));
  buf1  g5055(.din(new_new_n9810__), .dout(n18597));
  buf1  g5056(.din(new_new_n9818__), .dout(n18600));
  buf1  g5057(.din(new_new_n9829__), .dout(n18603));
  buf1  g5058(.din(new_new_n10397__), .dout(n18606));
  buf1  g5059(.din(new_new_n10423__), .dout(n18609));
  buf1  g5060(.din(new_new_n10408__), .dout(n18612));
  buf1  g5061(.din(new_new_n10438__), .dout(n18615));
  buf1  g5062(.din(new_new_n10452__), .dout(n18618));
  buf1  g5063(.din(new_new_n10455__), .dout(n18621));
  buf1  g5064(.din(new_new_n10458__), .dout(n18624));
  buf1  g5065(.din(new_new_n9925__), .dout(n18627));
  buf1  g5066(.din(new_new_n9924__), .dout(n18630));
  buf1  g5067(.din(new_new_n10435__), .dout(n18633));
  buf1  g5068(.din(new_new_n10343__), .dout(n18636));
  buf1  g5069(.din(new_new_n10347__), .dout(n18639));
  buf1  g5070(.din(new_new_n10351__), .dout(n18642));
  buf1  g5071(.din(new_new_n10355__), .dout(n18645));
  buf1  g5072(.din(new_new_n10341__), .dout(n18648));
  buf1  g5073(.din(new_new_n10349__), .dout(n18651));
  buf1  g5074(.din(new_new_n10357__), .dout(n18654));
  buf1  g5075(.din(new_new_n10353__), .dout(n18657));
  buf1  g5076(.din(new_new_n10130__), .dout(n18660));
  buf1  g5077(.din(new_new_n10119__), .dout(n18663));
  buf1  g5078(.din(new_new_n10097__), .dout(n18666));
  buf1  g5079(.din(new_new_n10163__), .dout(n18669));
  buf1  g5080(.din(new_new_n10158__), .dout(n18672));
  buf1  g5081(.din(new_new_n10149__), .dout(n18675));
  buf1  g5082(.din(new_new_n10142__), .dout(n18678));
  buf1  g5083(.din(new_new_n3570__), .dout(n18681));
  buf1  g5084(.din(new_new_n10029__), .dout(n18684));
  buf1  g5085(.din(new_new_n9942__), .dout(n18687));
  buf1  g5086(.din(new_new_n9950__), .dout(n18690));
  buf1  g5087(.din(new_new_n9928__), .dout(n18693));
  buf1  g5088(.din(new_new_n9936__), .dout(n18696));
  buf1  g5089(.din(new_new_n9770__), .dout(n18699));
  buf1  g5090(.din(new_new_n9906__), .dout(n18702));
  buf1  g5091(.din(new_new_n10011__), .dout(n18705));
  buf1  g5092(.din(n18705), .dout(n18708));
  buf1  g5093(.din(n18180), .dout(n18711));
  buf1  g5094(.din(new_new_n9872__), .dout(n18714));
  buf1  g5095(.din(n18714), .dout(n18717));
  buf1  g5096(.din(new_new_n10538__), .dout(n18720));
  buf1  g5097(.din(new_new_n10539__), .dout(n18723));
  buf1  g5098(.din(new_new_n10540__), .dout(n18726));
  buf1  g5099(.din(new_new_n10541__), .dout(n18729));
  buf1  g5100(.din(new_new_n10026__), .dout(n18732));
  buf1  g5101(.din(new_new_n10542__), .dout(n18735));
  buf1  g5102(.din(new_new_n10022__), .dout(n18738));
  buf1  g5103(.din(new_new_n10368__), .dout(n18741));
  buf1  g5104(.din(new_new_n10379__), .dout(n18744));
  buf1  g5105(.din(new_new_n10390__), .dout(n18747));
  buf1  g5106(.din(new_new_n10207__), .dout(n18750));
  buf1  g5107(.din(new_new_n10211__), .dout(n18753));
  buf1  g5108(.din(new_new_n10209__), .dout(n18756));
  buf1  g5109(.din(new_new_n10205__), .dout(n18759));
  buf1  g5110(.din(new_new_n10393__), .dout(n18762));
  buf1  g5111(.din(new_new_n10394__), .dout(n18765));
  buf1  g5112(.din(n18618), .dout(n18768));
  buf1  g5113(.din(new_new_n9914__), .dout(n18771));
  buf1  g5114(.din(new_new_n10338__), .dout(n18774));
  buf1  g5115(.din(new_new_n10493__), .dout(n18777));
  buf1  g5116(.din(new_new_n10503__), .dout(n18780));
  buf1  g5117(.din(new_new_n10495__), .dout(n18783));
  buf1  g5118(.din(new_new_n10504__), .dout(n18786));
  buf1  g5119(.din(n17646), .dout(n18789));
  buf1  g5120(.din(new_new_n6554__), .dout(n18792));
  buf1  g5121(.din(new_new_n6555__), .dout(n18795));
  buf1  g5122(.din(new_new_n6556__), .dout(n18798));
  buf1  g5123(.din(new_new_n6557__), .dout(n18801));
  buf1  g5124(.din(new_new_n6558__), .dout(n18804));
  buf1  g5125(.din(new_new_n6559__), .dout(n18807));
  buf1  g5126(.din(new_new_n6560__), .dout(n18810));
  buf1  g5127(.din(new_new_n6561__), .dout(n18813));
  buf1  g5128(.din(new_new_n6562__), .dout(n18816));
  buf1  g5129(.din(new_new_n10021__), .dout(n18819));
  buf1  g5130(.din(n18819), .dout(n18822));
  buf1  g5131(.din(n18201), .dout(n18825));
  buf1  g5132(.din(n18204), .dout(n18828));
  buf1  g5133(.din(n18207), .dout(n18831));
  buf1  g5134(.din(n18213), .dout(n18834));
  buf1  g5135(.din(new_new_n10367__), .dout(n18837));
  buf1  g5136(.din(n18411), .dout(n18840));
  buf1  g5137(.din(new_new_n10258__), .dout(n18843));
  buf1  g5138(.din(n18414), .dout(n18846));
  buf1  g5139(.din(new_new_n10306__), .dout(n18849));
  buf1  g5140(.din(new_new_n9710__), .dout(n18852));
  buf1  g5141(.din(new_new_n9703__), .dout(n18855));
  buf1  g5142(.din(new_new_n6563__), .dout(n18858));
  buf1  g5143(.din(new_new_n6564__), .dout(n18861));
  buf1  g5144(.din(new_new_n6565__), .dout(n18864));
  buf1  g5145(.din(new_new_n6566__), .dout(n18867));
  buf1  g5146(.din(new_new_n6567__), .dout(n18870));
  buf1  g5147(.din(new_new_n6568__), .dout(n18873));
  buf1  g5148(.din(new_new_n6569__), .dout(n18876));
  buf1  g5149(.din(new_new_n6570__), .dout(n18879));
  buf1  g5150(.din(new_new_n10030__), .dout(n18882));
  buf1  g5151(.din(new_new_n9996__), .dout(n18885));
  buf1  g5152(.din(new_new_n10028__), .dout(n18888));
  buf1  g5153(.din(new_new_n6574__), .dout(n18891));
  not1  g5154(.din(new_new_n10031__), .dout(n18894));
  not1  g5155(.din(new_new_n6577__), .dout(n18897));
  not1  g5156(.din(new_new_n10032__), .dout(n18900));
  not1  g5157(.din(new_new_n10014__), .dout(n18903));
  buf1  g5158(.din(new_new_n6579__), .dout(n18906));
  buf1  g5159(.din(new_new_n6580__), .dout(n18909));
  buf1  g5160(.din(new_new_n6584__), .dout(n18912));
  buf1  g5161(.din(new_new_n6585__), .dout(n18915));
  buf1  g5162(.din(new_new_n6586__), .dout(n18918));
  buf1  g5163(.din(new_new_n6587__), .dout(n18921));
  buf1  g5164(.din(new_new_n10012__), .dout(n18924));
  buf1  g5165(.din(new_new_n6589__), .dout(n18927));
  buf1  g5166(.din(new_new_n6590__), .dout(n18930));
  buf1  g5167(.din(new_new_n6591__), .dout(n18933));
  buf1  g5168(.din(new_new_n6593__), .dout(n18936));
  buf1  g5169(.din(n18576), .dout(n18939));
  buf1  g5170(.din(new_new_n10027__), .dout(n18942));
  buf1  g5171(.din(n18579), .dout(n18945));
  buf1  g5172(.din(new_new_n10025__), .dout(n18948));
  buf1  g5173(.din(new_new_n10023__), .dout(n18951));
  buf1  g5174(.din(n18660), .dout(n18954));
  buf1  g5175(.din(n18663), .dout(n18957));
  buf1  g5176(.din(n18666), .dout(n18960));
  buf1  g5177(.din(n18669), .dout(n18963));
  buf1  g5178(.din(n18672), .dout(n18966));
  buf1  g5179(.din(n18675), .dout(n18969));
  buf1  g5180(.din(n18678), .dout(n18972));
  buf1  g5181(.din(new_new_n6595__), .dout(n18975));
  buf1  g5182(.din(n18687), .dout(n18978));
  buf1  g5183(.din(n18690), .dout(n18981));
  buf1  g5184(.din(n18693), .dout(n18984));
  buf1  g5185(.din(n18696), .dout(n18987));
  buf1  g5186(.din(n18699), .dout(n18990));
  buf1  g5187(.din(n18702), .dout(n18993));
  buf1  g5188(.din(new_new_n6597__), .dout(n18996));
  buf1  g5189(.din(n18924), .dout(n18999));
  buf1  g5190(.din(new_new_n10519__), .dout(n19002));
  buf1  g5191(.din(new_new_n9873__), .dout(n19005));
  buf1  g5192(.din(n19005), .dout(n19008));
  buf1  g5193(.din(new_new_n6600__), .dout(n19011));
  buf1  g5194(.din(new_new_n6603__), .dout(n19014));
  buf1  g5195(.din(new_new_n6606__), .dout(n19017));
  buf1  g5196(.din(new_new_n6609__), .dout(n19020));
  buf1  g5197(.din(new_new_n6612__), .dout(n19023));
  buf1  g5198(.din(new_new_n6615__), .dout(n19026));
  buf1  g5199(.din(new_new_n6618__), .dout(n19029));
  buf1  g5200(.din(new_new_n6621__), .dout(n19032));
  buf1  g5201(.din(new_new_n6624__), .dout(n19035));
  buf1  g5202(.din(new_new_n6627__), .dout(n19038));
  buf1  g5203(.din(new_new_n6630__), .dout(n19041));
  buf1  g5204(.din(new_new_n6639__), .dout(n19044));
  buf1  g5205(.din(new_new_n6714__), .dout(n19047));
  buf1  g5206(.din(new_new_n6781__), .dout(n19050));
  buf1  g5207(.din(n18720), .dout(n19053));
  buf1  g5208(.din(n18723), .dout(n19056));
  buf1  g5209(.din(n18726), .dout(n19059));
  buf1  g5210(.din(n18729), .dout(n19062));
  buf1  g5211(.din(n18735), .dout(n19065));
  buf1  g5212(.din(new_new_n6888__), .dout(n19068));
  buf1  g5213(.din(new_new_n6969__), .dout(n19071));
  buf1  g5214(.din(new_new_n10381__), .dout(n19074));
  buf1  g5215(.din(new_new_n10392__), .dout(n19077));
  buf1  g5216(.din(new_new_n10486__), .dout(n19080));
  buf1  g5217(.din(new_new_n10488__), .dout(n19083));
  buf1  g5218(.din(new_new_n10543__), .dout(n19086));
  buf1  g5219(.din(n19086), .dout(n19089));
  buf1  g5220(.din(new_new_n10544__), .dout(n19092));
  buf1  g5221(.din(n19092), .dout(n19095));
  buf1  g5222(.din(new_new_n9913__), .dout(n19098));
  buf1  g5223(.din(new_new_n10545__), .dout(n19101));
  buf1  g5224(.din(new_new_n10546__), .dout(n19104));
  buf1  g5225(.din(new_new_n10547__), .dout(n19107));
  buf1  g5226(.din(new_new_n10548__), .dout(n19110));
  buf1  g5227(.din(new_new_n10549__), .dout(n19113));
  buf1  g5228(.din(new_new_n10550__), .dout(n19116));
  buf1  g5229(.din(new_new_n10552__), .dout(n19119));
  buf1  g5230(.din(new_new_n10554__), .dout(n19122));
  buf1  g5231(.din(new_new_n7130__), .dout(n19125));
  buf1  g5232(.din(new_new_n10407__), .dout(n19128));
  buf1  g5233(.din(new_new_n10473__), .dout(n19131));
  buf1  g5234(.din(new_new_n10476__), .dout(n19134));
  buf1  g5235(.din(new_new_n10505__), .dout(n19137));
  buf1  g5236(.din(new_new_n10508__), .dout(n19140));
  buf1  g5237(.din(new_new_n10491__), .dout(n19143));
  buf1  g5238(.din(new_new_n10496__), .dout(n19146));
  buf1  g5239(.din(new_new_n10498__), .dout(n19149));
  buf1  g5240(.din(new_new_n10499__), .dout(n19152));
  buf1  g5241(.din(n18783), .dout(n19155));
  buf1  g5242(.din(n18786), .dout(n19158));
  buf1  g5243(.din(new_new_n10523__), .dout(n19161));
  buf1  g5244(.din(new_new_n10526__), .dout(n19164));
  buf1  g5245(.din(new_new_n10529__), .dout(n19167));
  buf1  g5246(.din(new_new_n10532__), .dout(n19170));
  buf1  g5247(.din(n18288), .dout(n19173));
  buf1  g5248(.din(n18294), .dout(n19176));
  buf1  g5249(.din(n18324), .dout(n19179));
  buf1  g5250(.din(n18327), .dout(n19182));
  buf1  g5251(.din(new_new_n7141__), .dout(n19185));
  buf1  g5252(.din(new_new_n7143__), .dout(n19188));
  buf1  g5253(.din(n18375), .dout(n19191));
  buf1  g5254(.din(new_new_n7145__), .dout(n19194));
  buf1  g5255(.din(new_new_n7147__), .dout(n19197));
  buf1  g5256(.din(new_new_n7149__), .dout(n19200));
  buf1  g5257(.din(new_new_n7151__), .dout(n19203));
  not1  g5258(.din(new_new_n10483__), .dout(n19206));
  buf1  g5259(.din(new_new_n10479__), .dout(n19209));
  buf1  g5260(.din(new_new_n10487__), .dout(n19212));
  buf1  g5261(.din(new_new_n10489__), .dout(n19215));
  buf1  g5262(.din(new_new_n9915__), .dout(n19218));
  buf1  g5263(.din(new_new_n7156__), .dout(n19221));
  buf1  g5264(.din(new_new_n7172__), .dout(n19224));
  buf1  g5265(.din(new_new_n7188__), .dout(n19227));
  not1  g5266(.din(new_new_n7189__), .dout(n19230));
  buf1  g5267(.din(new_new_n7190__), .dout(n19233));
  buf1  g5268(.din(new_new_n7191__), .dout(n19236));
  buf1  g5269(.din(new_new_n10555__), .dout(n19239));
  buf1  g5270(.din(n19239), .dout(n19242));
  buf1  g5271(.din(new_new_n10556__), .dout(n19245));
  buf1  g5272(.din(n19245), .dout(n19248));
  buf1  g5273(.din(new_new_n10434__), .dout(n19251));
  buf1  g5274(.din(n19161), .dout(n19254));
  buf1  g5275(.din(n19164), .dout(n19257));
  buf1  g5276(.din(n19167), .dout(n19260));
  buf1  g5277(.din(n19170), .dout(n19263));
  buf1  g5278(.din(new_new_n7194__), .dout(n19266));
  buf1  g5279(.din(n18837), .dout(n19269));
  buf1  g5280(.din(n18843), .dout(n19272));
  buf1  g5281(.din(new_new_n10257__), .dout(n19275));
  buf1  g5282(.din(n18849), .dout(n19278));
  buf1  g5283(.din(new_new_n10305__), .dout(n19281));
  buf1  g5284(.din(n18852), .dout(n19284));
  buf1  g5285(.din(n18855), .dout(n19287));
  buf1  g5286(.din(n19074), .dout(n19290));
  buf1  g5287(.din(n19077), .dout(n19293));
  buf1  g5288(.din(n19218), .dout(n19296));
  buf1  g5289(.din(n19101), .dout(n19299));
  buf1  g5290(.din(n19104), .dout(n19302));
  buf1  g5291(.din(n19107), .dout(n19305));
  buf1  g5292(.din(n19110), .dout(n19308));
  buf1  g5293(.din(n19113), .dout(n19311));
  buf1  g5294(.din(n19116), .dout(n19314));
  buf1  g5295(.din(new_new_n10472__), .dout(n19317));
  buf1  g5296(.din(new_new_n10475__), .dout(n19320));
  buf1  g5297(.din(n19119), .dout(n19323));
  buf1  g5298(.din(n19122), .dout(n19326));
  buf1  g5299(.din(new_new_n10509__), .dout(n19329));
  buf1  g5300(.din(new_new_n7201__), .dout(n19332));
  buf1  g5301(.din(new_new_n10480__), .dout(n19335));
  not1  g5302(.din(new_new_n10484__), .dout(n19338));
  buf1  g5303(.din(new_new_n10481__), .dout(n19341));
  buf1  g5304(.din(new_new_n7213__), .dout(n19344));
  buf1  g5305(.din(new_new_n7217__), .dout(n19347));
  not1  g5306(.din(new_new_n10485__), .dout(n19350));
  not1  g5307(.din(new_new_n7225__), .dout(n19353));
  buf1  g5308(.din(new_new_n10478__), .dout(n19356));
  not1  g5309(.din(new_new_n10482__), .dout(n19359));
  not1  g5310(.din(new_new_n7239__), .dout(n19362));
  buf1  g5311(.din(new_new_n7259__), .dout(n19365));
  buf1  g5312(.din(new_new_n7260__), .dout(n19368));
  buf1  g5313(.din(new_new_n7261__), .dout(n19371));
  buf1  g5314(.din(new_new_n7262__), .dout(n19374));
  buf1  g5315(.din(new_new_n7263__), .dout(n19377));
  buf1  g5316(.din(new_new_n7266__), .dout(n19380));
  not1  g5317(.din(new_new_n7269__), .dout(n19383));
  buf1  g5318(.din(new_new_n7271__), .dout(n19386));
  buf1  g5319(.din(new_new_n7273__), .dout(n19389));
  buf1  g5320(.din(new_new_n7282__), .dout(n19392));
  buf1  g5321(.din(new_new_n7291__), .dout(n19395));
  buf1  g5322(.din(new_new_n10557__), .dout(n19398));
  buf1  g5323(.din(new_new_n10558__), .dout(n19401));
  buf1  g5324(.din(new_new_n10559__), .dout(n19404));
  buf1  g5325(.din(new_new_n10560__), .dout(n19407));
  buf1  g5326(.din(new_new_n10561__), .dout(n19410));
  buf1  g5327(.din(new_new_n10562__), .dout(n19413));
  buf1  g5328(.din(new_new_n10563__), .dout(n19416));
  buf1  g5329(.din(new_new_n10564__), .dout(n19419));
  buf1  g5330(.din(new_new_n10551__), .dout(n19422));
  buf1  g5331(.din(new_new_n10553__), .dout(n19425));
  buf1  g5332(.din(new_new_n7306__), .dout(n19428));
  buf1  g5333(.din(new_new_n2586__), .dout(n19431));
  buf1  g5334(.din(new_new_n2588__), .dout(n19434));
  buf1  g5335(.din(new_new_n2596__), .dout(n19437));
  buf1  g5336(.din(n19398), .dout(n19440));
  buf1  g5337(.din(n19401), .dout(n19443));
  buf1  g5338(.din(n19404), .dout(n19446));
  buf1  g5339(.din(n19407), .dout(n19449));
  buf1  g5340(.din(n19410), .dout(n19452));
  buf1  g5341(.din(n19413), .dout(n19455));
  buf1  g5342(.din(n19416), .dout(n19458));
  buf1  g5343(.din(n19419), .dout(n19461));
  buf1  g5344(.din(new_new_n3210__), .dout(new_new_n8443__));
  buf1  g5345(.din(new_new_n2690__), .dout(new_new_n8444__));
  buf1  g5346(.din(new_new_n3719__), .dout(new_new_n8445__));
  buf1  g5347(.din(new_new_n2771__), .dout(new_new_n8446__));
  buf1  g5348(.din(new_new_n3635__), .dout(new_new_n8447__));
  buf1  g5349(.din(new_new_n3549__), .dout(new_new_n8448__));
  buf1  g5350(.din(new_new_n4717__), .dout(new_new_n8449__));
  buf1  g5351(.din(new_new_n8449__), .dout(new_new_n8450__));
  buf1  g5352(.din(new_new_n8450__), .dout(new_new_n8451__));
  buf1  g5353(.din(new_new_n8451__), .dout(new_new_n8452__));
  buf1  g5354(.din(new_new_n8451__), .dout(new_new_n8453__));
  buf1  g5355(.din(new_new_n8450__), .dout(new_new_n8454__));
  buf1  g5356(.din(new_new_n8454__), .dout(new_new_n8455__));
  buf1  g5357(.din(new_new_n8454__), .dout(new_new_n8456__));
  buf1  g5358(.din(new_new_n8449__), .dout(new_new_n8457__));
  buf1  g5359(.din(new_new_n8457__), .dout(new_new_n8458__));
  buf1  g5360(.din(new_new_n8458__), .dout(new_new_n8459__));
  buf1  g5361(.din(new_new_n8457__), .dout(new_new_n8460__));
  buf1  g5362(.din(new_new_n3703__), .dout(new_new_n8461__));
  buf1  g5363(.din(new_new_n8461__), .dout(new_new_n8462__));
  buf1  g5364(.din(new_new_n8462__), .dout(new_new_n8463__));
  buf1  g5365(.din(new_new_n8462__), .dout(new_new_n8464__));
  buf1  g5366(.din(new_new_n8461__), .dout(new_new_n8465__));
  buf1  g5367(.din(new_new_n8465__), .dout(new_new_n8466__));
  buf1  g5368(.din(new_new_n8465__), .dout(new_new_n8467__));
  buf1  g5369(.din(new_new_n3702__), .dout(new_new_n8468__));
  buf1  g5370(.din(new_new_n8468__), .dout(new_new_n8469__));
  buf1  g5371(.din(new_new_n8469__), .dout(new_new_n8470__));
  buf1  g5372(.din(new_new_n8469__), .dout(new_new_n8471__));
  buf1  g5373(.din(new_new_n8468__), .dout(new_new_n8472__));
  buf1  g5374(.din(new_new_n8472__), .dout(new_new_n8473__));
  buf1  g5375(.din(new_new_n8472__), .dout(new_new_n8474__));
  buf1  g5376(.din(new_new_n2939__), .dout(new_new_n8475__));
  buf1  g5377(.din(new_new_n4716__), .dout(new_new_n8476__));
  buf1  g5378(.din(new_new_n4735__), .dout(new_new_n8477__));
  buf1  g5379(.din(new_new_n8477__), .dout(new_new_n8478__));
  buf1  g5380(.din(new_new_n8477__), .dout(new_new_n8479__));
  buf1  g5381(.din(new_new_n4736__), .dout(new_new_n8480__));
  buf1  g5382(.din(new_new_n8480__), .dout(new_new_n8481__));
  buf1  g5383(.din(new_new_n8480__), .dout(new_new_n8482__));
  buf1  g5384(.din(new_new_n3211__), .dout(new_new_n8483__));
  buf1  g5385(.din(new_new_n8483__), .dout(new_new_n8484__));
  buf1  g5386(.din(new_new_n8484__), .dout(new_new_n8485__));
  buf1  g5387(.din(new_new_n8483__), .dout(new_new_n8486__));
  buf1  g5388(.din(new_new_n3860__), .dout(new_new_n8487__));
  buf1  g5389(.din(new_new_n8487__), .dout(new_new_n8488__));
  buf1  g5390(.din(new_new_n3589__), .dout(new_new_n8489__));
  buf1  g5391(.din(new_new_n3490__), .dout(new_new_n8490__));
  buf1  g5392(.din(new_new_n3864__), .dout(new_new_n8491__));
  buf1  g5393(.din(new_new_n8491__), .dout(new_new_n8492__));
  buf1  g5394(.din(new_new_n3491__), .dout(new_new_n8493__));
  buf1  g5395(.din(new_new_n3887__), .dout(new_new_n8494__));
  buf1  g5396(.din(new_new_n8494__), .dout(new_new_n8495__));
  buf1  g5397(.din(new_new_n3893__), .dout(new_new_n8496__));
  buf1  g5398(.din(new_new_n8496__), .dout(new_new_n8497__));
  buf1  g5399(.din(new_new_n3585__), .dout(new_new_n8498__));
  buf1  g5400(.din(new_new_n3484__), .dout(new_new_n8499__));
  buf1  g5401(.din(new_new_n3485__), .dout(new_new_n8500__));
  buf1  g5402(.din(new_new_n3469__), .dout(new_new_n8501__));
  buf1  g5403(.din(new_new_n8501__), .dout(new_new_n8502__));
  buf1  g5404(.din(new_new_n3468__), .dout(new_new_n8503__));
  buf1  g5405(.din(new_new_n4784__), .dout(new_new_n8504__));
  buf1  g5406(.din(new_new_n4774__), .dout(new_new_n8505__));
  buf1  g5407(.din(new_new_n4787__), .dout(new_new_n8506__));
  buf1  g5408(.din(new_new_n3750__), .dout(new_new_n8507__));
  buf1  g5409(.din(new_new_n8507__), .dout(new_new_n8508__));
  buf1  g5410(.din(new_new_n8508__), .dout(new_new_n8509__));
  buf1  g5411(.din(new_new_n8509__), .dout(new_new_n8510__));
  buf1  g5412(.din(new_new_n8509__), .dout(new_new_n8511__));
  buf1  g5413(.din(new_new_n8508__), .dout(new_new_n8512__));
  buf1  g5414(.din(new_new_n8512__), .dout(new_new_n8513__));
  buf1  g5415(.din(new_new_n8512__), .dout(new_new_n8514__));
  buf1  g5416(.din(new_new_n8507__), .dout(new_new_n8515__));
  buf1  g5417(.din(new_new_n8515__), .dout(new_new_n8516__));
  buf1  g5418(.din(new_new_n8515__), .dout(new_new_n8517__));
  buf1  g5419(.din(new_new_n3603__), .dout(new_new_n8518__));
  buf1  g5420(.din(new_new_n3512__), .dout(new_new_n8519__));
  buf1  g5421(.din(new_new_n3742__), .dout(new_new_n8520__));
  buf1  g5422(.din(new_new_n8520__), .dout(new_new_n8521__));
  buf1  g5423(.din(new_new_n8521__), .dout(new_new_n8522__));
  buf1  g5424(.din(new_new_n8522__), .dout(new_new_n8523__));
  buf1  g5425(.din(new_new_n8522__), .dout(new_new_n8524__));
  buf1  g5426(.din(new_new_n8521__), .dout(new_new_n8525__));
  buf1  g5427(.din(new_new_n8525__), .dout(new_new_n8526__));
  buf1  g5428(.din(new_new_n8520__), .dout(new_new_n8527__));
  buf1  g5429(.din(new_new_n8527__), .dout(new_new_n8528__));
  buf1  g5430(.din(new_new_n8527__), .dout(new_new_n8529__));
  buf1  g5431(.din(new_new_n3513__), .dout(new_new_n8530__));
  buf1  g5432(.din(new_new_n3727__), .dout(new_new_n8531__));
  buf1  g5433(.din(new_new_n8531__), .dout(new_new_n8532__));
  buf1  g5434(.din(new_new_n8532__), .dout(new_new_n8533__));
  buf1  g5435(.din(new_new_n8533__), .dout(new_new_n8534__));
  buf1  g5436(.din(new_new_n8533__), .dout(new_new_n8535__));
  buf1  g5437(.din(new_new_n8532__), .dout(new_new_n8536__));
  buf1  g5438(.din(new_new_n8536__), .dout(new_new_n8537__));
  buf1  g5439(.din(new_new_n8536__), .dout(new_new_n8538__));
  buf1  g5440(.din(new_new_n8531__), .dout(new_new_n8539__));
  buf1  g5441(.din(new_new_n8539__), .dout(new_new_n8540__));
  buf1  g5442(.din(new_new_n8539__), .dout(new_new_n8541__));
  buf1  g5443(.din(new_new_n3735__), .dout(new_new_n8542__));
  buf1  g5444(.din(new_new_n8542__), .dout(new_new_n8543__));
  buf1  g5445(.din(new_new_n8543__), .dout(new_new_n8544__));
  buf1  g5446(.din(new_new_n8544__), .dout(new_new_n8545__));
  buf1  g5447(.din(new_new_n8544__), .dout(new_new_n8546__));
  buf1  g5448(.din(new_new_n8543__), .dout(new_new_n8547__));
  buf1  g5449(.din(new_new_n8547__), .dout(new_new_n8548__));
  buf1  g5450(.din(new_new_n8542__), .dout(new_new_n8549__));
  buf1  g5451(.din(new_new_n8549__), .dout(new_new_n8550__));
  buf1  g5452(.din(new_new_n8549__), .dout(new_new_n8551__));
  buf1  g5453(.din(new_new_n3601__), .dout(new_new_n8552__));
  buf1  g5454(.din(new_new_n3508__), .dout(new_new_n8553__));
  buf1  g5455(.din(new_new_n3509__), .dout(new_new_n8554__));
  buf1  g5456(.din(new_new_n3595__), .dout(new_new_n8555__));
  buf1  g5457(.din(new_new_n8555__), .dout(new_new_n8556__));
  buf1  g5458(.din(new_new_n3498__), .dout(new_new_n8557__));
  buf1  g5459(.din(new_new_n3499__), .dout(new_new_n8558__));
  buf1  g5460(.din(new_new_n3594__), .dout(new_new_n8559__));
  buf1  g5461(.din(new_new_n4816__), .dout(new_new_n8560__));
  buf1  g5462(.din(new_new_n4806__), .dout(new_new_n8561__));
  buf1  g5463(.din(new_new_n4819__), .dout(new_new_n8562__));
  buf1  g5464(.din(new_new_n4829__), .dout(new_new_n8563__));
  buf1  g5465(.din(new_new_n3567__), .dout(new_new_n8564__));
  buf1  g5466(.din(new_new_n8564__), .dout(new_new_n8565__));
  buf1  g5467(.din(new_new_n3410__), .dout(new_new_n8566__));
  buf1  g5468(.din(new_new_n3411__), .dout(new_new_n8567__));
  buf1  g5469(.din(new_new_n3566__), .dout(new_new_n8568__));
  buf1  g5470(.din(new_new_n3561__), .dout(new_new_n8569__));
  buf1  g5471(.din(new_new_n3402__), .dout(new_new_n8570__));
  buf1  g5472(.din(new_new_n3403__), .dout(new_new_n8571__));
  buf1  g5473(.din(new_new_n3581__), .dout(new_new_n8572__));
  buf1  g5474(.din(new_new_n3396__), .dout(new_new_n8573__));
  buf1  g5475(.din(new_new_n3397__), .dout(new_new_n8574__));
  buf1  g5476(.din(new_new_n3577__), .dout(new_new_n8575__));
  buf1  g5477(.din(new_new_n3390__), .dout(new_new_n8576__));
  buf1  g5478(.din(new_new_n3391__), .dout(new_new_n8577__));
  buf1  g5479(.din(new_new_n4854__), .dout(new_new_n8578__));
  buf1  g5480(.din(new_new_n4844__), .dout(new_new_n8579__));
  buf1  g5481(.din(new_new_n4864__), .dout(new_new_n8580__));
  buf1  g5482(.din(new_new_n4874__), .dout(new_new_n8581__));
  buf1  g5483(.din(new_new_n3541__), .dout(new_new_n8582__));
  buf1  g5484(.din(new_new_n3450__), .dout(new_new_n8583__));
  buf1  g5485(.din(new_new_n3451__), .dout(new_new_n8584__));
  buf1  g5486(.din(new_new_n3557__), .dout(new_new_n8585__));
  buf1  g5487(.din(new_new_n3448__), .dout(new_new_n8586__));
  buf1  g5488(.din(new_new_n3449__), .dout(new_new_n8587__));
  buf1  g5489(.din(new_new_n3555__), .dout(new_new_n8588__));
  buf1  g5490(.din(new_new_n3446__), .dout(new_new_n8589__));
  buf1  g5491(.din(new_new_n3447__), .dout(new_new_n8590__));
  buf1  g5492(.din(new_new_n3553__), .dout(new_new_n8591__));
  buf1  g5493(.din(new_new_n3442__), .dout(new_new_n8592__));
  buf1  g5494(.din(new_new_n3443__), .dout(new_new_n8593__));
  buf1  g5495(.din(new_new_n4897__), .dout(new_new_n8594__));
  buf1  g5496(.din(new_new_n4887__), .dout(new_new_n8595__));
  buf1  g5497(.din(new_new_n4907__), .dout(new_new_n8596__));
  buf1  g5498(.din(new_new_n4917__), .dout(new_new_n8597__));
  buf1  g5499(.din(new_new_n3829__), .dout(new_new_n8598__));
  buf1  g5500(.din(new_new_n3841__), .dout(new_new_n8599__));
  buf1  g5501(.din(new_new_n8599__), .dout(new_new_n8600__));
  buf1  g5502(.din(new_new_n3921__), .dout(new_new_n8601__));
  buf1  g5503(.din(new_new_n8601__), .dout(new_new_n8602__));
  buf1  g5504(.din(new_new_n8601__), .dout(new_new_n8603__));
  buf1  g5505(.din(new_new_n4925__), .dout(new_new_n8604__));
  buf1  g5506(.din(new_new_n4227__), .dout(new_new_n8605__));
  buf1  g5507(.din(new_new_n4112__), .dout(new_new_n8606__));
  buf1  g5508(.din(new_new_n8606__), .dout(new_new_n8607__));
  buf1  g5509(.din(new_new_n8606__), .dout(new_new_n8608__));
  buf1  g5510(.din(new_new_n4123__), .dout(new_new_n8609__));
  buf1  g5511(.din(new_new_n8609__), .dout(new_new_n8610__));
  buf1  g5512(.din(new_new_n4210__), .dout(new_new_n8611__));
  buf1  g5513(.din(new_new_n8611__), .dout(new_new_n8612__));
  buf1  g5514(.din(new_new_n8612__), .dout(new_new_n8613__));
  buf1  g5515(.din(new_new_n8612__), .dout(new_new_n8614__));
  buf1  g5516(.din(new_new_n8611__), .dout(new_new_n8615__));
  buf1  g5517(.din(new_new_n4422__), .dout(new_new_n8616__));
  buf1  g5518(.din(new_new_n8616__), .dout(new_new_n8617__));
  buf1  g5519(.din(new_new_n8617__), .dout(new_new_n8618__));
  buf1  g5520(.din(new_new_n8618__), .dout(new_new_n8619__));
  buf1  g5521(.din(new_new_n8617__), .dout(new_new_n8620__));
  buf1  g5522(.din(new_new_n8616__), .dout(new_new_n8621__));
  buf1  g5523(.din(new_new_n8621__), .dout(new_new_n8622__));
  buf1  g5524(.din(new_new_n8621__), .dout(new_new_n8623__));
  buf1  g5525(.din(new_new_n4281__), .dout(new_new_n8624__));
  buf1  g5526(.din(new_new_n8624__), .dout(new_new_n8625__));
  buf1  g5527(.din(new_new_n4423__), .dout(new_new_n8626__));
  buf1  g5528(.din(new_new_n8626__), .dout(new_new_n8627__));
  buf1  g5529(.din(new_new_n8627__), .dout(new_new_n8628__));
  buf1  g5530(.din(new_new_n8628__), .dout(new_new_n8629__));
  buf1  g5531(.din(new_new_n8627__), .dout(new_new_n8630__));
  buf1  g5532(.din(new_new_n8626__), .dout(new_new_n8631__));
  buf1  g5533(.din(new_new_n8631__), .dout(new_new_n8632__));
  buf1  g5534(.din(new_new_n8631__), .dout(new_new_n8633__));
  buf1  g5535(.din(new_new_n4280__), .dout(new_new_n8634__));
  buf1  g5536(.din(new_new_n8634__), .dout(new_new_n8635__));
  buf1  g5537(.din(new_new_n4424__), .dout(new_new_n8636__));
  buf1  g5538(.din(new_new_n8636__), .dout(new_new_n8637__));
  buf1  g5539(.din(new_new_n8637__), .dout(new_new_n8638__));
  buf1  g5540(.din(new_new_n8637__), .dout(new_new_n8639__));
  buf1  g5541(.din(new_new_n8636__), .dout(new_new_n8640__));
  buf1  g5542(.din(new_new_n4425__), .dout(new_new_n8641__));
  buf1  g5543(.din(new_new_n8641__), .dout(new_new_n8642__));
  buf1  g5544(.din(new_new_n8642__), .dout(new_new_n8643__));
  buf1  g5545(.din(new_new_n8642__), .dout(new_new_n8644__));
  buf1  g5546(.din(new_new_n8641__), .dout(new_new_n8645__));
  buf1  g5547(.din(new_new_n4420__), .dout(new_new_n8646__));
  buf1  g5548(.din(new_new_n8646__), .dout(new_new_n8647__));
  buf1  g5549(.din(new_new_n8647__), .dout(new_new_n8648__));
  buf1  g5550(.din(new_new_n8647__), .dout(new_new_n8649__));
  buf1  g5551(.din(new_new_n8646__), .dout(new_new_n8650__));
  buf1  g5552(.din(new_new_n4421__), .dout(new_new_n8651__));
  buf1  g5553(.din(new_new_n8651__), .dout(new_new_n8652__));
  buf1  g5554(.din(new_new_n8652__), .dout(new_new_n8653__));
  buf1  g5555(.din(new_new_n8652__), .dout(new_new_n8654__));
  buf1  g5556(.din(new_new_n8651__), .dout(new_new_n8655__));
  buf1  g5557(.din(new_new_n4426__), .dout(new_new_n8656__));
  buf1  g5558(.din(new_new_n8656__), .dout(new_new_n8657__));
  buf1  g5559(.din(new_new_n8657__), .dout(new_new_n8658__));
  buf1  g5560(.din(new_new_n8657__), .dout(new_new_n8659__));
  buf1  g5561(.din(new_new_n8656__), .dout(new_new_n8660__));
  buf1  g5562(.din(new_new_n4427__), .dout(new_new_n8661__));
  buf1  g5563(.din(new_new_n8661__), .dout(new_new_n8662__));
  buf1  g5564(.din(new_new_n8662__), .dout(new_new_n8663__));
  buf1  g5565(.din(new_new_n8662__), .dout(new_new_n8664__));
  buf1  g5566(.din(new_new_n8661__), .dout(new_new_n8665__));
  buf1  g5567(.din(new_new_n4937__), .dout(new_new_n8666__));
  buf1  g5568(.din(new_new_n4929__), .dout(new_new_n8667__));
  buf1  g5569(.din(new_new_n3831__), .dout(new_new_n8668__));
  buf1  g5570(.din(new_new_n3842__), .dout(new_new_n8669__));
  buf1  g5571(.din(new_new_n8669__), .dout(new_new_n8670__));
  buf1  g5572(.din(new_new_n3922__), .dout(new_new_n8671__));
  buf1  g5573(.din(new_new_n8671__), .dout(new_new_n8672__));
  buf1  g5574(.din(new_new_n8671__), .dout(new_new_n8673__));
  buf1  g5575(.din(new_new_n4941__), .dout(new_new_n8674__));
  buf1  g5576(.din(new_new_n4223__), .dout(new_new_n8675__));
  buf1  g5577(.din(new_new_n4119__), .dout(new_new_n8676__));
  buf1  g5578(.din(new_new_n8676__), .dout(new_new_n8677__));
  buf1  g5579(.din(new_new_n8676__), .dout(new_new_n8678__));
  buf1  g5580(.din(new_new_n4121__), .dout(new_new_n8679__));
  buf1  g5581(.din(new_new_n8679__), .dout(new_new_n8680__));
  buf1  g5582(.din(new_new_n4225__), .dout(new_new_n8681__));
  buf1  g5583(.din(new_new_n8681__), .dout(new_new_n8682__));
  buf1  g5584(.din(new_new_n8682__), .dout(new_new_n8683__));
  buf1  g5585(.din(new_new_n8681__), .dout(new_new_n8684__));
  buf1  g5586(.din(new_new_n4412__), .dout(new_new_n8685__));
  buf1  g5587(.din(new_new_n8685__), .dout(new_new_n8686__));
  buf1  g5588(.din(new_new_n8686__), .dout(new_new_n8687__));
  buf1  g5589(.din(new_new_n8687__), .dout(new_new_n8688__));
  buf1  g5590(.din(new_new_n8686__), .dout(new_new_n8689__));
  buf1  g5591(.din(new_new_n8685__), .dout(new_new_n8690__));
  buf1  g5592(.din(new_new_n8690__), .dout(new_new_n8691__));
  buf1  g5593(.din(new_new_n8690__), .dout(new_new_n8692__));
  buf1  g5594(.din(new_new_n4410__), .dout(new_new_n8693__));
  buf1  g5595(.din(new_new_n8693__), .dout(new_new_n8694__));
  buf1  g5596(.din(new_new_n4413__), .dout(new_new_n8695__));
  buf1  g5597(.din(new_new_n8695__), .dout(new_new_n8696__));
  buf1  g5598(.din(new_new_n8696__), .dout(new_new_n8697__));
  buf1  g5599(.din(new_new_n8697__), .dout(new_new_n8698__));
  buf1  g5600(.din(new_new_n8696__), .dout(new_new_n8699__));
  buf1  g5601(.din(new_new_n8695__), .dout(new_new_n8700__));
  buf1  g5602(.din(new_new_n8700__), .dout(new_new_n8701__));
  buf1  g5603(.din(new_new_n8700__), .dout(new_new_n8702__));
  buf1  g5604(.din(new_new_n4411__), .dout(new_new_n8703__));
  buf1  g5605(.din(new_new_n8703__), .dout(new_new_n8704__));
  buf1  g5606(.din(new_new_n4414__), .dout(new_new_n8705__));
  buf1  g5607(.din(new_new_n8705__), .dout(new_new_n8706__));
  buf1  g5608(.din(new_new_n8706__), .dout(new_new_n8707__));
  buf1  g5609(.din(new_new_n8706__), .dout(new_new_n8708__));
  buf1  g5610(.din(new_new_n8705__), .dout(new_new_n8709__));
  buf1  g5611(.din(new_new_n4415__), .dout(new_new_n8710__));
  buf1  g5612(.din(new_new_n8710__), .dout(new_new_n8711__));
  buf1  g5613(.din(new_new_n8711__), .dout(new_new_n8712__));
  buf1  g5614(.din(new_new_n8711__), .dout(new_new_n8713__));
  buf1  g5615(.din(new_new_n8710__), .dout(new_new_n8714__));
  buf1  g5616(.din(new_new_n4418__), .dout(new_new_n8715__));
  buf1  g5617(.din(new_new_n8715__), .dout(new_new_n8716__));
  buf1  g5618(.din(new_new_n8716__), .dout(new_new_n8717__));
  buf1  g5619(.din(new_new_n8716__), .dout(new_new_n8718__));
  buf1  g5620(.din(new_new_n8715__), .dout(new_new_n8719__));
  buf1  g5621(.din(new_new_n4419__), .dout(new_new_n8720__));
  buf1  g5622(.din(new_new_n8720__), .dout(new_new_n8721__));
  buf1  g5623(.din(new_new_n8721__), .dout(new_new_n8722__));
  buf1  g5624(.din(new_new_n8721__), .dout(new_new_n8723__));
  buf1  g5625(.din(new_new_n8720__), .dout(new_new_n8724__));
  buf1  g5626(.din(new_new_n4416__), .dout(new_new_n8725__));
  buf1  g5627(.din(new_new_n8725__), .dout(new_new_n8726__));
  buf1  g5628(.din(new_new_n8726__), .dout(new_new_n8727__));
  buf1  g5629(.din(new_new_n8726__), .dout(new_new_n8728__));
  buf1  g5630(.din(new_new_n8725__), .dout(new_new_n8729__));
  buf1  g5631(.din(new_new_n4417__), .dout(new_new_n8730__));
  buf1  g5632(.din(new_new_n8730__), .dout(new_new_n8731__));
  buf1  g5633(.din(new_new_n8731__), .dout(new_new_n8732__));
  buf1  g5634(.din(new_new_n8731__), .dout(new_new_n8733__));
  buf1  g5635(.din(new_new_n8730__), .dout(new_new_n8734__));
  buf1  g5636(.din(new_new_n4953__), .dout(new_new_n8735__));
  buf1  g5637(.din(new_new_n4945__), .dout(new_new_n8736__));
  buf1  g5638(.din(new_new_n4965__), .dout(new_new_n8737__));
  buf1  g5639(.din(new_new_n4960__), .dout(new_new_n8738__));
  buf1  g5640(.din(new_new_n4966__), .dout(new_new_n8739__));
  buf1  g5641(.din(new_new_n4959__), .dout(new_new_n8740__));
  buf1  g5642(.din(new_new_n4975__), .dout(new_new_n8741__));
  buf1  g5643(.din(new_new_n8741__), .dout(new_new_n8742__));
  buf1  g5644(.din(new_new_n8741__), .dout(new_new_n8743__));
  buf1  g5645(.din(new_new_n4974__), .dout(new_new_n8744__));
  buf1  g5646(.din(new_new_n8744__), .dout(new_new_n8745__));
  buf1  g5647(.din(new_new_n8744__), .dout(new_new_n8746__));
  buf1  g5648(.din(new_new_n4976__), .dout(new_new_n8747__));
  buf1  g5649(.din(new_new_n8747__), .dout(new_new_n8748__));
  buf1  g5650(.din(new_new_n8747__), .dout(new_new_n8749__));
  buf1  g5651(.din(new_new_n4973__), .dout(new_new_n8750__));
  buf1  g5652(.din(new_new_n8750__), .dout(new_new_n8751__));
  buf1  g5653(.din(new_new_n8750__), .dout(new_new_n8752__));
  buf1  g5654(.din(new_new_n4261__), .dout(new_new_n8753__));
  buf1  g5655(.din(new_new_n8753__), .dout(new_new_n8754__));
  buf1  g5656(.din(new_new_n8753__), .dout(new_new_n8755__));
  buf1  g5657(.din(new_new_n4260__), .dout(new_new_n8756__));
  buf1  g5658(.din(new_new_n8756__), .dout(new_new_n8757__));
  buf1  g5659(.din(new_new_n8756__), .dout(new_new_n8758__));
  buf1  g5660(.din(new_new_n5012__), .dout(new_new_n8759__));
  buf1  g5661(.din(new_new_n5007__), .dout(new_new_n8760__));
  buf1  g5662(.din(new_new_n5013__), .dout(new_new_n8761__));
  buf1  g5663(.din(new_new_n5006__), .dout(new_new_n8762__));
  buf1  g5664(.din(new_new_n5022__), .dout(new_new_n8763__));
  buf1  g5665(.din(new_new_n8763__), .dout(new_new_n8764__));
  buf1  g5666(.din(new_new_n8763__), .dout(new_new_n8765__));
  buf1  g5667(.din(new_new_n5021__), .dout(new_new_n8766__));
  buf1  g5668(.din(new_new_n8766__), .dout(new_new_n8767__));
  buf1  g5669(.din(new_new_n8766__), .dout(new_new_n8768__));
  buf1  g5670(.din(new_new_n5023__), .dout(new_new_n8769__));
  buf1  g5671(.din(new_new_n8769__), .dout(new_new_n8770__));
  buf1  g5672(.din(new_new_n8769__), .dout(new_new_n8771__));
  buf1  g5673(.din(new_new_n5020__), .dout(new_new_n8772__));
  buf1  g5674(.din(new_new_n8772__), .dout(new_new_n8773__));
  buf1  g5675(.din(new_new_n8772__), .dout(new_new_n8774__));
  buf1  g5676(.din(new_new_n4408__), .dout(new_new_n8775__));
  buf1  g5677(.din(new_new_n8775__), .dout(new_new_n8776__));
  buf1  g5678(.din(new_new_n8775__), .dout(new_new_n8777__));
  buf1  g5679(.din(new_new_n4409__), .dout(new_new_n8778__));
  buf1  g5680(.din(new_new_n8778__), .dout(new_new_n8779__));
  buf1  g5681(.din(new_new_n8778__), .dout(new_new_n8780__));
  buf1  g5682(.din(new_new_n3573__), .dout(new_new_n8781__));
  buf1  g5683(.din(new_new_n8781__), .dout(new_new_n8782__));
  buf1  g5684(.din(new_new_n5049__), .dout(new_new_n8783__));
  buf1  g5685(.din(new_new_n4204__), .dout(new_new_n8784__));
  buf1  g5686(.din(new_new_n4109__), .dout(new_new_n8785__));
  buf1  g5687(.din(new_new_n4111__), .dout(new_new_n8786__));
  buf1  g5688(.din(new_new_n3903__), .dout(new_new_n8787__));
  buf1  g5689(.din(new_new_n8787__), .dout(new_new_n8788__));
  buf1  g5690(.din(new_new_n8787__), .dout(new_new_n8789__));
  buf1  g5691(.din(new_new_n4274__), .dout(new_new_n8790__));
  buf1  g5692(.din(new_new_n4275__), .dout(new_new_n8791__));
  buf1  g5693(.din(new_new_n4276__), .dout(new_new_n8792__));
  buf1  g5694(.din(new_new_n8792__), .dout(new_new_n8793__));
  buf1  g5695(.din(new_new_n4277__), .dout(new_new_n8794__));
  buf1  g5696(.din(new_new_n8794__), .dout(new_new_n8795__));
  buf1  g5697(.din(new_new_n4278__), .dout(new_new_n8796__));
  buf1  g5698(.din(new_new_n8796__), .dout(new_new_n8797__));
  buf1  g5699(.din(new_new_n4279__), .dout(new_new_n8798__));
  buf1  g5700(.din(new_new_n8798__), .dout(new_new_n8799__));
  buf1  g5701(.din(new_new_n5084__), .dout(new_new_n8800__));
  buf1  g5702(.din(new_new_n5085__), .dout(new_new_n8801__));
  buf1  g5703(.din(new_new_n4283__), .dout(new_new_n8802__));
  buf1  g5704(.din(new_new_n8802__), .dout(new_new_n8803__));
  buf1  g5705(.din(new_new_n8802__), .dout(new_new_n8804__));
  buf1  g5706(.din(new_new_n4282__), .dout(new_new_n8805__));
  buf1  g5707(.din(new_new_n8805__), .dout(new_new_n8806__));
  buf1  g5708(.din(new_new_n8805__), .dout(new_new_n8807__));
  buf1  g5709(.din(new_new_n5098__), .dout(new_new_n8808__));
  buf1  g5710(.din(new_new_n4191__), .dout(new_new_n8809__));
  buf1  g5711(.din(new_new_n4107__), .dout(new_new_n8810__));
  buf1  g5712(.din(new_new_n4105__), .dout(new_new_n8811__));
  buf1  g5713(.din(new_new_n4264__), .dout(new_new_n8812__));
  buf1  g5714(.din(new_new_n4265__), .dout(new_new_n8813__));
  buf1  g5715(.din(new_new_n4266__), .dout(new_new_n8814__));
  buf1  g5716(.din(new_new_n8814__), .dout(new_new_n8815__));
  buf1  g5717(.din(new_new_n4267__), .dout(new_new_n8816__));
  buf1  g5718(.din(new_new_n8816__), .dout(new_new_n8817__));
  buf1  g5719(.din(new_new_n4268__), .dout(new_new_n8818__));
  buf1  g5720(.din(new_new_n8818__), .dout(new_new_n8819__));
  buf1  g5721(.din(new_new_n4269__), .dout(new_new_n8820__));
  buf1  g5722(.din(new_new_n8820__), .dout(new_new_n8821__));
  buf1  g5723(.din(new_new_n5125__), .dout(new_new_n8822__));
  buf1  g5724(.din(new_new_n5126__), .dout(new_new_n8823__));
  buf1  g5725(.din(new_new_n4262__), .dout(new_new_n8824__));
  buf1  g5726(.din(new_new_n8824__), .dout(new_new_n8825__));
  buf1  g5727(.din(new_new_n8824__), .dout(new_new_n8826__));
  buf1  g5728(.din(new_new_n4263__), .dout(new_new_n8827__));
  buf1  g5729(.din(new_new_n8827__), .dout(new_new_n8828__));
  buf1  g5730(.din(new_new_n8827__), .dout(new_new_n8829__));
  buf1  g5731(.din(new_new_n5139__), .dout(new_new_n8830__));
  buf1  g5732(.din(new_new_n3862__), .dout(new_new_n8831__));
  buf1  g5733(.din(new_new_n3866__), .dout(new_new_n8832__));
  buf1  g5734(.din(new_new_n3806__), .dout(new_new_n8833__));
  buf1  g5735(.din(new_new_n8833__), .dout(new_new_n8834__));
  buf1  g5736(.din(new_new_n8834__), .dout(new_new_n8835__));
  buf1  g5737(.din(new_new_n8835__), .dout(new_new_n8836__));
  buf1  g5738(.din(new_new_n8836__), .dout(new_new_n8837__));
  buf1  g5739(.din(new_new_n8837__), .dout(new_new_n8838__));
  buf1  g5740(.din(new_new_n8837__), .dout(new_new_n8839__));
  buf1  g5741(.din(new_new_n8836__), .dout(new_new_n8840__));
  buf1  g5742(.din(new_new_n8840__), .dout(new_new_n8841__));
  buf1  g5743(.din(new_new_n8840__), .dout(new_new_n8842__));
  buf1  g5744(.din(new_new_n8835__), .dout(new_new_n8843__));
  buf1  g5745(.din(new_new_n8843__), .dout(new_new_n8844__));
  buf1  g5746(.din(new_new_n8844__), .dout(new_new_n8845__));
  buf1  g5747(.din(new_new_n8844__), .dout(new_new_n8846__));
  buf1  g5748(.din(new_new_n8843__), .dout(new_new_n8847__));
  buf1  g5749(.din(new_new_n8847__), .dout(new_new_n8848__));
  buf1  g5750(.din(new_new_n8847__), .dout(new_new_n8849__));
  buf1  g5751(.din(new_new_n8834__), .dout(new_new_n8850__));
  buf1  g5752(.din(new_new_n8850__), .dout(new_new_n8851__));
  buf1  g5753(.din(new_new_n8851__), .dout(new_new_n8852__));
  buf1  g5754(.din(new_new_n8852__), .dout(new_new_n8853__));
  buf1  g5755(.din(new_new_n8851__), .dout(new_new_n8854__));
  buf1  g5756(.din(new_new_n8850__), .dout(new_new_n8855__));
  buf1  g5757(.din(new_new_n8855__), .dout(new_new_n8856__));
  buf1  g5758(.din(new_new_n8855__), .dout(new_new_n8857__));
  buf1  g5759(.din(new_new_n8833__), .dout(new_new_n8858__));
  buf1  g5760(.din(new_new_n8858__), .dout(new_new_n8859__));
  buf1  g5761(.din(new_new_n8859__), .dout(new_new_n8860__));
  buf1  g5762(.din(new_new_n8860__), .dout(new_new_n8861__));
  buf1  g5763(.din(new_new_n8860__), .dout(new_new_n8862__));
  buf1  g5764(.din(new_new_n8859__), .dout(new_new_n8863__));
  buf1  g5765(.din(new_new_n8863__), .dout(new_new_n8864__));
  buf1  g5766(.din(new_new_n8863__), .dout(new_new_n8865__));
  buf1  g5767(.din(new_new_n8858__), .dout(new_new_n8866__));
  buf1  g5768(.din(new_new_n8866__), .dout(new_new_n8867__));
  buf1  g5769(.din(new_new_n8867__), .dout(new_new_n8868__));
  buf1  g5770(.din(new_new_n8867__), .dout(new_new_n8869__));
  buf1  g5771(.din(new_new_n8866__), .dout(new_new_n8870__));
  buf1  g5772(.din(new_new_n8870__), .dout(new_new_n8871__));
  buf1  g5773(.din(new_new_n8870__), .dout(new_new_n8872__));
  buf1  g5774(.din(new_new_n3814__), .dout(new_new_n8873__));
  buf1  g5775(.din(new_new_n8873__), .dout(new_new_n8874__));
  buf1  g5776(.din(new_new_n8874__), .dout(new_new_n8875__));
  buf1  g5777(.din(new_new_n8875__), .dout(new_new_n8876__));
  buf1  g5778(.din(new_new_n8876__), .dout(new_new_n8877__));
  buf1  g5779(.din(new_new_n8877__), .dout(new_new_n8878__));
  buf1  g5780(.din(new_new_n8877__), .dout(new_new_n8879__));
  buf1  g5781(.din(new_new_n8876__), .dout(new_new_n8880__));
  buf1  g5782(.din(new_new_n8880__), .dout(new_new_n8881__));
  buf1  g5783(.din(new_new_n8880__), .dout(new_new_n8882__));
  buf1  g5784(.din(new_new_n8875__), .dout(new_new_n8883__));
  buf1  g5785(.din(new_new_n8883__), .dout(new_new_n8884__));
  buf1  g5786(.din(new_new_n8884__), .dout(new_new_n8885__));
  buf1  g5787(.din(new_new_n8884__), .dout(new_new_n8886__));
  buf1  g5788(.din(new_new_n8883__), .dout(new_new_n8887__));
  buf1  g5789(.din(new_new_n8887__), .dout(new_new_n8888__));
  buf1  g5790(.din(new_new_n8887__), .dout(new_new_n8889__));
  buf1  g5791(.din(new_new_n8874__), .dout(new_new_n8890__));
  buf1  g5792(.din(new_new_n8890__), .dout(new_new_n8891__));
  buf1  g5793(.din(new_new_n8891__), .dout(new_new_n8892__));
  buf1  g5794(.din(new_new_n8892__), .dout(new_new_n8893__));
  buf1  g5795(.din(new_new_n8891__), .dout(new_new_n8894__));
  buf1  g5796(.din(new_new_n8890__), .dout(new_new_n8895__));
  buf1  g5797(.din(new_new_n8895__), .dout(new_new_n8896__));
  buf1  g5798(.din(new_new_n8895__), .dout(new_new_n8897__));
  buf1  g5799(.din(new_new_n8873__), .dout(new_new_n8898__));
  buf1  g5800(.din(new_new_n8898__), .dout(new_new_n8899__));
  buf1  g5801(.din(new_new_n8899__), .dout(new_new_n8900__));
  buf1  g5802(.din(new_new_n8900__), .dout(new_new_n8901__));
  buf1  g5803(.din(new_new_n8900__), .dout(new_new_n8902__));
  buf1  g5804(.din(new_new_n8899__), .dout(new_new_n8903__));
  buf1  g5805(.din(new_new_n8903__), .dout(new_new_n8904__));
  buf1  g5806(.din(new_new_n8903__), .dout(new_new_n8905__));
  buf1  g5807(.din(new_new_n8898__), .dout(new_new_n8906__));
  buf1  g5808(.din(new_new_n8906__), .dout(new_new_n8907__));
  buf1  g5809(.din(new_new_n8907__), .dout(new_new_n8908__));
  buf1  g5810(.din(new_new_n8907__), .dout(new_new_n8909__));
  buf1  g5811(.din(new_new_n8906__), .dout(new_new_n8910__));
  buf1  g5812(.din(new_new_n8910__), .dout(new_new_n8911__));
  buf1  g5813(.din(new_new_n8910__), .dout(new_new_n8912__));
  buf1  g5814(.din(new_new_n2850__), .dout(new_new_n8913__));
  buf1  g5815(.din(new_new_n8913__), .dout(new_new_n8914__));
  buf1  g5816(.din(new_new_n2851__), .dout(new_new_n8915__));
  buf1  g5817(.din(new_new_n8915__), .dout(new_new_n8916__));
  buf1  g5818(.din(new_new_n5161__), .dout(new_new_n8917__));
  buf1  g5819(.din(new_new_n3807__), .dout(new_new_n8918__));
  buf1  g5820(.din(new_new_n8918__), .dout(new_new_n8919__));
  buf1  g5821(.din(new_new_n8919__), .dout(new_new_n8920__));
  buf1  g5822(.din(new_new_n8920__), .dout(new_new_n8921__));
  buf1  g5823(.din(new_new_n8921__), .dout(new_new_n8922__));
  buf1  g5824(.din(new_new_n8921__), .dout(new_new_n8923__));
  buf1  g5825(.din(new_new_n8920__), .dout(new_new_n8924__));
  buf1  g5826(.din(new_new_n8924__), .dout(new_new_n8925__));
  buf1  g5827(.din(new_new_n8924__), .dout(new_new_n8926__));
  buf1  g5828(.din(new_new_n8919__), .dout(new_new_n8927__));
  buf1  g5829(.din(new_new_n8927__), .dout(new_new_n8928__));
  buf1  g5830(.din(new_new_n8928__), .dout(new_new_n8929__));
  buf1  g5831(.din(new_new_n8928__), .dout(new_new_n8930__));
  buf1  g5832(.din(new_new_n8927__), .dout(new_new_n8931__));
  buf1  g5833(.din(new_new_n8931__), .dout(new_new_n8932__));
  buf1  g5834(.din(new_new_n8931__), .dout(new_new_n8933__));
  buf1  g5835(.din(new_new_n8918__), .dout(new_new_n8934__));
  buf1  g5836(.din(new_new_n8934__), .dout(new_new_n8935__));
  buf1  g5837(.din(new_new_n8935__), .dout(new_new_n8936__));
  buf1  g5838(.din(new_new_n8935__), .dout(new_new_n8937__));
  buf1  g5839(.din(new_new_n8934__), .dout(new_new_n8938__));
  buf1  g5840(.din(new_new_n8938__), .dout(new_new_n8939__));
  buf1  g5841(.din(new_new_n8938__), .dout(new_new_n8940__));
  buf1  g5842(.din(new_new_n3815__), .dout(new_new_n8941__));
  buf1  g5843(.din(new_new_n8941__), .dout(new_new_n8942__));
  buf1  g5844(.din(new_new_n8942__), .dout(new_new_n8943__));
  buf1  g5845(.din(new_new_n8943__), .dout(new_new_n8944__));
  buf1  g5846(.din(new_new_n8944__), .dout(new_new_n8945__));
  buf1  g5847(.din(new_new_n8944__), .dout(new_new_n8946__));
  buf1  g5848(.din(new_new_n8943__), .dout(new_new_n8947__));
  buf1  g5849(.din(new_new_n8947__), .dout(new_new_n8948__));
  buf1  g5850(.din(new_new_n8947__), .dout(new_new_n8949__));
  buf1  g5851(.din(new_new_n8942__), .dout(new_new_n8950__));
  buf1  g5852(.din(new_new_n8950__), .dout(new_new_n8951__));
  buf1  g5853(.din(new_new_n8951__), .dout(new_new_n8952__));
  buf1  g5854(.din(new_new_n8951__), .dout(new_new_n8953__));
  buf1  g5855(.din(new_new_n8950__), .dout(new_new_n8954__));
  buf1  g5856(.din(new_new_n8954__), .dout(new_new_n8955__));
  buf1  g5857(.din(new_new_n8954__), .dout(new_new_n8956__));
  buf1  g5858(.din(new_new_n8941__), .dout(new_new_n8957__));
  buf1  g5859(.din(new_new_n8957__), .dout(new_new_n8958__));
  buf1  g5860(.din(new_new_n8958__), .dout(new_new_n8959__));
  buf1  g5861(.din(new_new_n8958__), .dout(new_new_n8960__));
  buf1  g5862(.din(new_new_n8957__), .dout(new_new_n8961__));
  buf1  g5863(.din(new_new_n8961__), .dout(new_new_n8962__));
  buf1  g5864(.din(new_new_n8961__), .dout(new_new_n8963__));
  buf1  g5865(.din(new_new_n5171__), .dout(new_new_n8964__));
  buf1  g5866(.din(new_new_n8964__), .dout(new_new_n8965__));
  buf1  g5867(.din(new_new_n5170__), .dout(new_new_n8966__));
  buf1  g5868(.din(new_new_n8966__), .dout(new_new_n8967__));
  buf1  g5869(.din(new_new_n5176__), .dout(new_new_n8968__));
  buf1  g5870(.din(new_new_n2698__), .dout(new_new_n8969__));
  buf1  g5871(.din(new_new_n8969__), .dout(new_new_n8970__));
  buf1  g5872(.din(new_new_n2699__), .dout(new_new_n8971__));
  buf1  g5873(.din(new_new_n8971__), .dout(new_new_n8972__));
  buf1  g5874(.din(new_new_n5187__), .dout(new_new_n8973__));
  buf1  g5875(.din(new_new_n4404__), .dout(new_new_n8974__));
  buf1  g5876(.din(new_new_n4399__), .dout(new_new_n8975__));
  buf1  g5877(.din(new_new_n4405__), .dout(new_new_n8976__));
  buf1  g5878(.din(new_new_n4398__), .dout(new_new_n8977__));
  buf1  g5879(.din(new_new_n5202__), .dout(new_new_n8978__));
  buf1  g5880(.din(new_new_n8978__), .dout(new_new_n8979__));
  buf1  g5881(.din(new_new_n8979__), .dout(new_new_n8980__));
  buf1  g5882(.din(new_new_n8978__), .dout(new_new_n8981__));
  buf1  g5883(.din(new_new_n5203__), .dout(new_new_n8982__));
  buf1  g5884(.din(new_new_n8982__), .dout(new_new_n8983__));
  buf1  g5885(.din(new_new_n8983__), .dout(new_new_n8984__));
  buf1  g5886(.din(new_new_n8982__), .dout(new_new_n8985__));
  buf1  g5887(.din(new_new_n5210__), .dout(new_new_n8986__));
  buf1  g5888(.din(new_new_n5211__), .dout(new_new_n8987__));
  buf1  g5889(.din(new_new_n4211__), .dout(new_new_n8988__));
  buf1  g5890(.din(new_new_n5167__), .dout(new_new_n8989__));
  buf1  g5891(.din(new_new_n8989__), .dout(new_new_n8990__));
  buf1  g5892(.din(new_new_n8990__), .dout(new_new_n8991__));
  buf1  g5893(.din(new_new_n8989__), .dout(new_new_n8992__));
  buf1  g5894(.din(new_new_n3782__), .dout(new_new_n8993__));
  buf1  g5895(.din(new_new_n8993__), .dout(new_new_n8994__));
  buf1  g5896(.din(new_new_n8994__), .dout(new_new_n8995__));
  buf1  g5897(.din(new_new_n8995__), .dout(new_new_n8996__));
  buf1  g5898(.din(new_new_n8996__), .dout(new_new_n8997__));
  buf1  g5899(.din(new_new_n8996__), .dout(new_new_n8998__));
  buf1  g5900(.din(new_new_n8995__), .dout(new_new_n8999__));
  buf1  g5901(.din(new_new_n8999__), .dout(new_new_n9000__));
  buf1  g5902(.din(new_new_n8999__), .dout(new_new_n9001__));
  buf1  g5903(.din(new_new_n8994__), .dout(new_new_n9002__));
  buf1  g5904(.din(new_new_n9002__), .dout(new_new_n9003__));
  buf1  g5905(.din(new_new_n9002__), .dout(new_new_n9004__));
  buf1  g5906(.din(new_new_n8993__), .dout(new_new_n9005__));
  buf1  g5907(.din(new_new_n9005__), .dout(new_new_n9006__));
  buf1  g5908(.din(new_new_n9006__), .dout(new_new_n9007__));
  buf1  g5909(.din(new_new_n9006__), .dout(new_new_n9008__));
  buf1  g5910(.din(new_new_n9005__), .dout(new_new_n9009__));
  buf1  g5911(.din(new_new_n9009__), .dout(new_new_n9010__));
  buf1  g5912(.din(new_new_n9009__), .dout(new_new_n9011__));
  buf1  g5913(.din(new_new_n3774__), .dout(new_new_n9012__));
  buf1  g5914(.din(new_new_n9012__), .dout(new_new_n9013__));
  buf1  g5915(.din(new_new_n9013__), .dout(new_new_n9014__));
  buf1  g5916(.din(new_new_n9014__), .dout(new_new_n9015__));
  buf1  g5917(.din(new_new_n9015__), .dout(new_new_n9016__));
  buf1  g5918(.din(new_new_n9015__), .dout(new_new_n9017__));
  buf1  g5919(.din(new_new_n9014__), .dout(new_new_n9018__));
  buf1  g5920(.din(new_new_n9018__), .dout(new_new_n9019__));
  buf1  g5921(.din(new_new_n9018__), .dout(new_new_n9020__));
  buf1  g5922(.din(new_new_n9013__), .dout(new_new_n9021__));
  buf1  g5923(.din(new_new_n9021__), .dout(new_new_n9022__));
  buf1  g5924(.din(new_new_n9021__), .dout(new_new_n9023__));
  buf1  g5925(.din(new_new_n9012__), .dout(new_new_n9024__));
  buf1  g5926(.din(new_new_n9024__), .dout(new_new_n9025__));
  buf1  g5927(.din(new_new_n9025__), .dout(new_new_n9026__));
  buf1  g5928(.din(new_new_n9025__), .dout(new_new_n9027__));
  buf1  g5929(.din(new_new_n9024__), .dout(new_new_n9028__));
  buf1  g5930(.din(new_new_n9028__), .dout(new_new_n9029__));
  buf1  g5931(.din(new_new_n9028__), .dout(new_new_n9030__));
  buf1  g5932(.din(new_new_n5193__), .dout(new_new_n9031__));
  buf1  g5933(.din(new_new_n9031__), .dout(new_new_n9032__));
  buf1  g5934(.din(new_new_n9032__), .dout(new_new_n9033__));
  buf1  g5935(.din(new_new_n9031__), .dout(new_new_n9034__));
  buf1  g5936(.din(new_new_n3783__), .dout(new_new_n9035__));
  buf1  g5937(.din(new_new_n9035__), .dout(new_new_n9036__));
  buf1  g5938(.din(new_new_n9036__), .dout(new_new_n9037__));
  buf1  g5939(.din(new_new_n9037__), .dout(new_new_n9038__));
  buf1  g5940(.din(new_new_n9038__), .dout(new_new_n9039__));
  buf1  g5941(.din(new_new_n9038__), .dout(new_new_n9040__));
  buf1  g5942(.din(new_new_n9037__), .dout(new_new_n9041__));
  buf1  g5943(.din(new_new_n9041__), .dout(new_new_n9042__));
  buf1  g5944(.din(new_new_n9041__), .dout(new_new_n9043__));
  buf1  g5945(.din(new_new_n9036__), .dout(new_new_n9044__));
  buf1  g5946(.din(new_new_n9044__), .dout(new_new_n9045__));
  buf1  g5947(.din(new_new_n9044__), .dout(new_new_n9046__));
  buf1  g5948(.din(new_new_n9035__), .dout(new_new_n9047__));
  buf1  g5949(.din(new_new_n9047__), .dout(new_new_n9048__));
  buf1  g5950(.din(new_new_n9048__), .dout(new_new_n9049__));
  buf1  g5951(.din(new_new_n9048__), .dout(new_new_n9050__));
  buf1  g5952(.din(new_new_n9047__), .dout(new_new_n9051__));
  buf1  g5953(.din(new_new_n9051__), .dout(new_new_n9052__));
  buf1  g5954(.din(new_new_n9051__), .dout(new_new_n9053__));
  buf1  g5955(.din(new_new_n2706__), .dout(new_new_n9054__));
  buf1  g5956(.din(new_new_n3775__), .dout(new_new_n9055__));
  buf1  g5957(.din(new_new_n9055__), .dout(new_new_n9056__));
  buf1  g5958(.din(new_new_n9056__), .dout(new_new_n9057__));
  buf1  g5959(.din(new_new_n9057__), .dout(new_new_n9058__));
  buf1  g5960(.din(new_new_n9058__), .dout(new_new_n9059__));
  buf1  g5961(.din(new_new_n9058__), .dout(new_new_n9060__));
  buf1  g5962(.din(new_new_n9057__), .dout(new_new_n9061__));
  buf1  g5963(.din(new_new_n9061__), .dout(new_new_n9062__));
  buf1  g5964(.din(new_new_n9061__), .dout(new_new_n9063__));
  buf1  g5965(.din(new_new_n9056__), .dout(new_new_n9064__));
  buf1  g5966(.din(new_new_n9064__), .dout(new_new_n9065__));
  buf1  g5967(.din(new_new_n9064__), .dout(new_new_n9066__));
  buf1  g5968(.din(new_new_n9055__), .dout(new_new_n9067__));
  buf1  g5969(.din(new_new_n9067__), .dout(new_new_n9068__));
  buf1  g5970(.din(new_new_n9068__), .dout(new_new_n9069__));
  buf1  g5971(.din(new_new_n9068__), .dout(new_new_n9070__));
  buf1  g5972(.din(new_new_n9067__), .dout(new_new_n9071__));
  buf1  g5973(.din(new_new_n9071__), .dout(new_new_n9072__));
  buf1  g5974(.din(new_new_n9071__), .dout(new_new_n9073__));
  buf1  g5975(.din(new_new_n2858__), .dout(new_new_n9074__));
  buf1  g5976(.din(new_new_n5237__), .dout(new_new_n9075__));
  buf1  g5977(.din(new_new_n5238__), .dout(new_new_n9076__));
  buf1  g5978(.din(new_new_n5241__), .dout(new_new_n9077__));
  buf1  g5979(.din(new_new_n5242__), .dout(new_new_n9078__));
  buf1  g5980(.din(new_new_n5247__), .dout(new_new_n9079__));
  buf1  g5981(.din(new_new_n5248__), .dout(new_new_n9080__));
  buf1  g5982(.din(new_new_n5261__), .dout(new_new_n9081__));
  buf1  g5983(.din(new_new_n5278__), .dout(new_new_n9082__));
  buf1  g5984(.din(new_new_n5297__), .dout(new_new_n9083__));
  buf1  g5985(.din(new_new_n3790__), .dout(new_new_n9084__));
  buf1  g5986(.din(new_new_n9084__), .dout(new_new_n9085__));
  buf1  g5987(.din(new_new_n9085__), .dout(new_new_n9086__));
  buf1  g5988(.din(new_new_n9086__), .dout(new_new_n9087__));
  buf1  g5989(.din(new_new_n9087__), .dout(new_new_n9088__));
  buf1  g5990(.din(new_new_n9087__), .dout(new_new_n9089__));
  buf1  g5991(.din(new_new_n9086__), .dout(new_new_n9090__));
  buf1  g5992(.din(new_new_n9090__), .dout(new_new_n9091__));
  buf1  g5993(.din(new_new_n9090__), .dout(new_new_n9092__));
  buf1  g5994(.din(new_new_n9085__), .dout(new_new_n9093__));
  buf1  g5995(.din(new_new_n9093__), .dout(new_new_n9094__));
  buf1  g5996(.din(new_new_n9093__), .dout(new_new_n9095__));
  buf1  g5997(.din(new_new_n9084__), .dout(new_new_n9096__));
  buf1  g5998(.din(new_new_n9096__), .dout(new_new_n9097__));
  buf1  g5999(.din(new_new_n9097__), .dout(new_new_n9098__));
  buf1  g6000(.din(new_new_n9097__), .dout(new_new_n9099__));
  buf1  g6001(.din(new_new_n9096__), .dout(new_new_n9100__));
  buf1  g6002(.din(new_new_n9100__), .dout(new_new_n9101__));
  buf1  g6003(.din(new_new_n9100__), .dout(new_new_n9102__));
  buf1  g6004(.din(new_new_n3798__), .dout(new_new_n9103__));
  buf1  g6005(.din(new_new_n9103__), .dout(new_new_n9104__));
  buf1  g6006(.din(new_new_n9104__), .dout(new_new_n9105__));
  buf1  g6007(.din(new_new_n9105__), .dout(new_new_n9106__));
  buf1  g6008(.din(new_new_n9106__), .dout(new_new_n9107__));
  buf1  g6009(.din(new_new_n9106__), .dout(new_new_n9108__));
  buf1  g6010(.din(new_new_n9105__), .dout(new_new_n9109__));
  buf1  g6011(.din(new_new_n9109__), .dout(new_new_n9110__));
  buf1  g6012(.din(new_new_n9109__), .dout(new_new_n9111__));
  buf1  g6013(.din(new_new_n9104__), .dout(new_new_n9112__));
  buf1  g6014(.din(new_new_n9112__), .dout(new_new_n9113__));
  buf1  g6015(.din(new_new_n9112__), .dout(new_new_n9114__));
  buf1  g6016(.din(new_new_n9103__), .dout(new_new_n9115__));
  buf1  g6017(.din(new_new_n9115__), .dout(new_new_n9116__));
  buf1  g6018(.din(new_new_n9116__), .dout(new_new_n9117__));
  buf1  g6019(.din(new_new_n9116__), .dout(new_new_n9118__));
  buf1  g6020(.din(new_new_n9115__), .dout(new_new_n9119__));
  buf1  g6021(.din(new_new_n9119__), .dout(new_new_n9120__));
  buf1  g6022(.din(new_new_n9119__), .dout(new_new_n9121__));
  buf1  g6023(.din(new_new_n3791__), .dout(new_new_n9122__));
  buf1  g6024(.din(new_new_n9122__), .dout(new_new_n9123__));
  buf1  g6025(.din(new_new_n9123__), .dout(new_new_n9124__));
  buf1  g6026(.din(new_new_n9124__), .dout(new_new_n9125__));
  buf1  g6027(.din(new_new_n9125__), .dout(new_new_n9126__));
  buf1  g6028(.din(new_new_n9125__), .dout(new_new_n9127__));
  buf1  g6029(.din(new_new_n9124__), .dout(new_new_n9128__));
  buf1  g6030(.din(new_new_n9128__), .dout(new_new_n9129__));
  buf1  g6031(.din(new_new_n9128__), .dout(new_new_n9130__));
  buf1  g6032(.din(new_new_n9123__), .dout(new_new_n9131__));
  buf1  g6033(.din(new_new_n9131__), .dout(new_new_n9132__));
  buf1  g6034(.din(new_new_n9131__), .dout(new_new_n9133__));
  buf1  g6035(.din(new_new_n9122__), .dout(new_new_n9134__));
  buf1  g6036(.din(new_new_n9134__), .dout(new_new_n9135__));
  buf1  g6037(.din(new_new_n9135__), .dout(new_new_n9136__));
  buf1  g6038(.din(new_new_n9135__), .dout(new_new_n9137__));
  buf1  g6039(.din(new_new_n9134__), .dout(new_new_n9138__));
  buf1  g6040(.din(new_new_n9138__), .dout(new_new_n9139__));
  buf1  g6041(.din(new_new_n9138__), .dout(new_new_n9140__));
  buf1  g6042(.din(new_new_n3799__), .dout(new_new_n9141__));
  buf1  g6043(.din(new_new_n9141__), .dout(new_new_n9142__));
  buf1  g6044(.din(new_new_n9142__), .dout(new_new_n9143__));
  buf1  g6045(.din(new_new_n9143__), .dout(new_new_n9144__));
  buf1  g6046(.din(new_new_n9144__), .dout(new_new_n9145__));
  buf1  g6047(.din(new_new_n9144__), .dout(new_new_n9146__));
  buf1  g6048(.din(new_new_n9143__), .dout(new_new_n9147__));
  buf1  g6049(.din(new_new_n9147__), .dout(new_new_n9148__));
  buf1  g6050(.din(new_new_n9147__), .dout(new_new_n9149__));
  buf1  g6051(.din(new_new_n9142__), .dout(new_new_n9150__));
  buf1  g6052(.din(new_new_n9150__), .dout(new_new_n9151__));
  buf1  g6053(.din(new_new_n9150__), .dout(new_new_n9152__));
  buf1  g6054(.din(new_new_n9141__), .dout(new_new_n9153__));
  buf1  g6055(.din(new_new_n9153__), .dout(new_new_n9154__));
  buf1  g6056(.din(new_new_n9154__), .dout(new_new_n9155__));
  buf1  g6057(.din(new_new_n9154__), .dout(new_new_n9156__));
  buf1  g6058(.din(new_new_n9153__), .dout(new_new_n9157__));
  buf1  g6059(.din(new_new_n9157__), .dout(new_new_n9158__));
  buf1  g6060(.din(new_new_n9157__), .dout(new_new_n9159__));
  buf1  g6061(.din(new_new_n5319__), .dout(new_new_n9160__));
  buf1  g6062(.din(new_new_n5320__), .dout(new_new_n9161__));
  buf1  g6063(.din(new_new_n5323__), .dout(new_new_n9162__));
  buf1  g6064(.din(new_new_n5324__), .dout(new_new_n9163__));
  buf1  g6065(.din(new_new_n5327__), .dout(new_new_n9164__));
  buf1  g6066(.din(new_new_n9164__), .dout(new_new_n9165__));
  buf1  g6067(.din(new_new_n5328__), .dout(new_new_n9166__));
  buf1  g6068(.din(new_new_n9166__), .dout(new_new_n9167__));
  buf1  g6069(.din(new_new_n5331__), .dout(new_new_n9168__));
  buf1  g6070(.din(new_new_n5332__), .dout(new_new_n9169__));
  buf1  g6071(.din(new_new_n5345__), .dout(new_new_n9170__));
  buf1  g6072(.din(new_new_n5362__), .dout(new_new_n9171__));
  buf1  g6073(.din(new_new_n5381__), .dout(new_new_n9172__));
  buf1  g6074(.din(new_new_n5394__), .dout(new_new_n9173__));
  buf1  g6075(.din(new_new_n5411__), .dout(new_new_n9174__));
  buf1  g6076(.din(new_new_n5406__), .dout(new_new_n9175__));
  buf1  g6077(.din(new_new_n5412__), .dout(new_new_n9176__));
  buf1  g6078(.din(new_new_n5405__), .dout(new_new_n9177__));
  buf1  g6079(.din(new_new_n5421__), .dout(new_new_n9178__));
  buf1  g6080(.din(new_new_n9178__), .dout(new_new_n9179__));
  buf1  g6081(.din(new_new_n9178__), .dout(new_new_n9180__));
  buf1  g6082(.din(new_new_n5420__), .dout(new_new_n9181__));
  buf1  g6083(.din(new_new_n9181__), .dout(new_new_n9182__));
  buf1  g6084(.din(new_new_n9181__), .dout(new_new_n9183__));
  buf1  g6085(.din(new_new_n5422__), .dout(new_new_n9184__));
  buf1  g6086(.din(new_new_n9184__), .dout(new_new_n9185__));
  buf1  g6087(.din(new_new_n9184__), .dout(new_new_n9186__));
  buf1  g6088(.din(new_new_n5419__), .dout(new_new_n9187__));
  buf1  g6089(.din(new_new_n9187__), .dout(new_new_n9188__));
  buf1  g6090(.din(new_new_n9187__), .dout(new_new_n9189__));
  buf1  g6091(.din(new_new_n4428__), .dout(new_new_n9190__));
  buf1  g6092(.din(new_new_n9190__), .dout(new_new_n9191__));
  buf1  g6093(.din(new_new_n9190__), .dout(new_new_n9192__));
  buf1  g6094(.din(new_new_n4429__), .dout(new_new_n9193__));
  buf1  g6095(.din(new_new_n9193__), .dout(new_new_n9194__));
  buf1  g6096(.din(new_new_n9193__), .dout(new_new_n9195__));
  buf1  g6097(.din(new_new_n5458__), .dout(new_new_n9196__));
  buf1  g6098(.din(new_new_n5453__), .dout(new_new_n9197__));
  buf1  g6099(.din(new_new_n5459__), .dout(new_new_n9198__));
  buf1  g6100(.din(new_new_n5452__), .dout(new_new_n9199__));
  buf1  g6101(.din(new_new_n5468__), .dout(new_new_n9200__));
  buf1  g6102(.din(new_new_n9200__), .dout(new_new_n9201__));
  buf1  g6103(.din(new_new_n9200__), .dout(new_new_n9202__));
  buf1  g6104(.din(new_new_n5467__), .dout(new_new_n9203__));
  buf1  g6105(.din(new_new_n9203__), .dout(new_new_n9204__));
  buf1  g6106(.din(new_new_n9203__), .dout(new_new_n9205__));
  buf1  g6107(.din(new_new_n5469__), .dout(new_new_n9206__));
  buf1  g6108(.din(new_new_n9206__), .dout(new_new_n9207__));
  buf1  g6109(.din(new_new_n9206__), .dout(new_new_n9208__));
  buf1  g6110(.din(new_new_n5466__), .dout(new_new_n9209__));
  buf1  g6111(.din(new_new_n9209__), .dout(new_new_n9210__));
  buf1  g6112(.din(new_new_n9209__), .dout(new_new_n9211__));
  buf1  g6113(.din(new_new_n4431__), .dout(new_new_n9212__));
  buf1  g6114(.din(new_new_n9212__), .dout(new_new_n9213__));
  buf1  g6115(.din(new_new_n9212__), .dout(new_new_n9214__));
  buf1  g6116(.din(new_new_n4430__), .dout(new_new_n9215__));
  buf1  g6117(.din(new_new_n9215__), .dout(new_new_n9216__));
  buf1  g6118(.din(new_new_n9215__), .dout(new_new_n9217__));
  buf1  g6119(.din(new_new_n5497__), .dout(new_new_n9218__));
  buf1  g6120(.din(new_new_n9218__), .dout(new_new_n9219__));
  buf1  g6121(.din(new_new_n9218__), .dout(new_new_n9220__));
  buf1  g6122(.din(new_new_n5498__), .dout(new_new_n9221__));
  buf1  g6123(.din(new_new_n9221__), .dout(new_new_n9222__));
  buf1  g6124(.din(new_new_n9221__), .dout(new_new_n9223__));
  buf1  g6125(.din(new_new_n5501__), .dout(new_new_n9224__));
  buf1  g6126(.din(new_new_n5510__), .dout(new_new_n9225__));
  buf1  g6127(.din(new_new_n5523__), .dout(new_new_n9226__));
  buf1  g6128(.din(new_new_n5538__), .dout(new_new_n9227__));
  buf1  g6129(.din(new_new_n5549__), .dout(new_new_n9228__));
  buf1  g6130(.din(new_new_n5558__), .dout(new_new_n9229__));
  buf1  g6131(.din(new_new_n5571__), .dout(new_new_n9230__));
  buf1  g6132(.din(new_new_n5221__), .dout(new_new_n9231__));
  buf1  g6133(.din(new_new_n9231__), .dout(new_new_n9232__));
  buf1  g6134(.din(new_new_n9231__), .dout(new_new_n9233__));
  buf1  g6135(.din(new_new_n3664__), .dout(new_new_n9234__));
  buf1  g6136(.din(new_new_n9234__), .dout(new_new_n9235__));
  buf1  g6137(.din(new_new_n9235__), .dout(new_new_n9236__));
  buf1  g6138(.din(new_new_n9236__), .dout(new_new_n9237__));
  buf1  g6139(.din(new_new_n9237__), .dout(new_new_n9238__));
  buf1  g6140(.din(new_new_n9237__), .dout(new_new_n9239__));
  buf1  g6141(.din(new_new_n9236__), .dout(new_new_n9240__));
  buf1  g6142(.din(new_new_n9240__), .dout(new_new_n9241__));
  buf1  g6143(.din(new_new_n9240__), .dout(new_new_n9242__));
  buf1  g6144(.din(new_new_n9235__), .dout(new_new_n9243__));
  buf1  g6145(.din(new_new_n9243__), .dout(new_new_n9244__));
  buf1  g6146(.din(new_new_n9243__), .dout(new_new_n9245__));
  buf1  g6147(.din(new_new_n9234__), .dout(new_new_n9246__));
  buf1  g6148(.din(new_new_n9246__), .dout(new_new_n9247__));
  buf1  g6149(.din(new_new_n9247__), .dout(new_new_n9248__));
  buf1  g6150(.din(new_new_n9247__), .dout(new_new_n9249__));
  buf1  g6151(.din(new_new_n9246__), .dout(new_new_n9250__));
  buf1  g6152(.din(new_new_n9250__), .dout(new_new_n9251__));
  buf1  g6153(.din(new_new_n9250__), .dout(new_new_n9252__));
  buf1  g6154(.din(new_new_n3672__), .dout(new_new_n9253__));
  buf1  g6155(.din(new_new_n9253__), .dout(new_new_n9254__));
  buf1  g6156(.din(new_new_n9254__), .dout(new_new_n9255__));
  buf1  g6157(.din(new_new_n9255__), .dout(new_new_n9256__));
  buf1  g6158(.din(new_new_n9256__), .dout(new_new_n9257__));
  buf1  g6159(.din(new_new_n9256__), .dout(new_new_n9258__));
  buf1  g6160(.din(new_new_n9255__), .dout(new_new_n9259__));
  buf1  g6161(.din(new_new_n9259__), .dout(new_new_n9260__));
  buf1  g6162(.din(new_new_n9259__), .dout(new_new_n9261__));
  buf1  g6163(.din(new_new_n9254__), .dout(new_new_n9262__));
  buf1  g6164(.din(new_new_n9262__), .dout(new_new_n9263__));
  buf1  g6165(.din(new_new_n9262__), .dout(new_new_n9264__));
  buf1  g6166(.din(new_new_n9253__), .dout(new_new_n9265__));
  buf1  g6167(.din(new_new_n9265__), .dout(new_new_n9266__));
  buf1  g6168(.din(new_new_n9266__), .dout(new_new_n9267__));
  buf1  g6169(.din(new_new_n9266__), .dout(new_new_n9268__));
  buf1  g6170(.din(new_new_n9265__), .dout(new_new_n9269__));
  buf1  g6171(.din(new_new_n9269__), .dout(new_new_n9270__));
  buf1  g6172(.din(new_new_n9269__), .dout(new_new_n9271__));
  buf1  g6173(.din(new_new_n3665__), .dout(new_new_n9272__));
  buf1  g6174(.din(new_new_n9272__), .dout(new_new_n9273__));
  buf1  g6175(.din(new_new_n9273__), .dout(new_new_n9274__));
  buf1  g6176(.din(new_new_n9274__), .dout(new_new_n9275__));
  buf1  g6177(.din(new_new_n9275__), .dout(new_new_n9276__));
  buf1  g6178(.din(new_new_n9275__), .dout(new_new_n9277__));
  buf1  g6179(.din(new_new_n9274__), .dout(new_new_n9278__));
  buf1  g6180(.din(new_new_n9278__), .dout(new_new_n9279__));
  buf1  g6181(.din(new_new_n9278__), .dout(new_new_n9280__));
  buf1  g6182(.din(new_new_n9273__), .dout(new_new_n9281__));
  buf1  g6183(.din(new_new_n9281__), .dout(new_new_n9282__));
  buf1  g6184(.din(new_new_n9281__), .dout(new_new_n9283__));
  buf1  g6185(.din(new_new_n9272__), .dout(new_new_n9284__));
  buf1  g6186(.din(new_new_n9284__), .dout(new_new_n9285__));
  buf1  g6187(.din(new_new_n9285__), .dout(new_new_n9286__));
  buf1  g6188(.din(new_new_n9285__), .dout(new_new_n9287__));
  buf1  g6189(.din(new_new_n9284__), .dout(new_new_n9288__));
  buf1  g6190(.din(new_new_n9288__), .dout(new_new_n9289__));
  buf1  g6191(.din(new_new_n9288__), .dout(new_new_n9290__));
  buf1  g6192(.din(new_new_n3322__), .dout(new_new_n9291__));
  buf1  g6193(.din(new_new_n3673__), .dout(new_new_n9292__));
  buf1  g6194(.din(new_new_n9292__), .dout(new_new_n9293__));
  buf1  g6195(.din(new_new_n9293__), .dout(new_new_n9294__));
  buf1  g6196(.din(new_new_n9294__), .dout(new_new_n9295__));
  buf1  g6197(.din(new_new_n9295__), .dout(new_new_n9296__));
  buf1  g6198(.din(new_new_n9295__), .dout(new_new_n9297__));
  buf1  g6199(.din(new_new_n9294__), .dout(new_new_n9298__));
  buf1  g6200(.din(new_new_n9298__), .dout(new_new_n9299__));
  buf1  g6201(.din(new_new_n9298__), .dout(new_new_n9300__));
  buf1  g6202(.din(new_new_n9293__), .dout(new_new_n9301__));
  buf1  g6203(.din(new_new_n9301__), .dout(new_new_n9302__));
  buf1  g6204(.din(new_new_n9301__), .dout(new_new_n9303__));
  buf1  g6205(.din(new_new_n9292__), .dout(new_new_n9304__));
  buf1  g6206(.din(new_new_n9304__), .dout(new_new_n9305__));
  buf1  g6207(.din(new_new_n9305__), .dout(new_new_n9306__));
  buf1  g6208(.din(new_new_n9305__), .dout(new_new_n9307__));
  buf1  g6209(.din(new_new_n9304__), .dout(new_new_n9308__));
  buf1  g6210(.din(new_new_n9308__), .dout(new_new_n9309__));
  buf1  g6211(.din(new_new_n9308__), .dout(new_new_n9310__));
  buf1  g6212(.din(new_new_n3330__), .dout(new_new_n9311__));
  buf1  g6213(.din(new_new_n3194__), .dout(new_new_n9312__));
  buf1  g6214(.din(new_new_n9312__), .dout(new_new_n9313__));
  buf1  g6215(.din(new_new_n9313__), .dout(new_new_n9314__));
  buf1  g6216(.din(new_new_n9314__), .dout(new_new_n9315__));
  buf1  g6217(.din(new_new_n9315__), .dout(new_new_n9316__));
  buf1  g6218(.din(new_new_n9315__), .dout(new_new_n9317__));
  buf1  g6219(.din(new_new_n9314__), .dout(new_new_n9318__));
  buf1  g6220(.din(new_new_n9318__), .dout(new_new_n9319__));
  buf1  g6221(.din(new_new_n9318__), .dout(new_new_n9320__));
  buf1  g6222(.din(new_new_n9313__), .dout(new_new_n9321__));
  buf1  g6223(.din(new_new_n9321__), .dout(new_new_n9322__));
  buf1  g6224(.din(new_new_n9322__), .dout(new_new_n9323__));
  buf1  g6225(.din(new_new_n9321__), .dout(new_new_n9324__));
  buf1  g6226(.din(new_new_n9312__), .dout(new_new_n9325__));
  buf1  g6227(.din(new_new_n9325__), .dout(new_new_n9326__));
  buf1  g6228(.din(new_new_n9326__), .dout(new_new_n9327__));
  buf1  g6229(.din(new_new_n9326__), .dout(new_new_n9328__));
  buf1  g6230(.din(new_new_n9325__), .dout(new_new_n9329__));
  buf1  g6231(.din(new_new_n9329__), .dout(new_new_n9330__));
  buf1  g6232(.din(new_new_n9329__), .dout(new_new_n9331__));
  buf1  g6233(.din(new_new_n3680__), .dout(new_new_n9332__));
  buf1  g6234(.din(new_new_n9332__), .dout(new_new_n9333__));
  buf1  g6235(.din(new_new_n9333__), .dout(new_new_n9334__));
  buf1  g6236(.din(new_new_n9334__), .dout(new_new_n9335__));
  buf1  g6237(.din(new_new_n9335__), .dout(new_new_n9336__));
  buf1  g6238(.din(new_new_n9335__), .dout(new_new_n9337__));
  buf1  g6239(.din(new_new_n9334__), .dout(new_new_n9338__));
  buf1  g6240(.din(new_new_n9338__), .dout(new_new_n9339__));
  buf1  g6241(.din(new_new_n9338__), .dout(new_new_n9340__));
  buf1  g6242(.din(new_new_n9333__), .dout(new_new_n9341__));
  buf1  g6243(.din(new_new_n9341__), .dout(new_new_n9342__));
  buf1  g6244(.din(new_new_n9341__), .dout(new_new_n9343__));
  buf1  g6245(.din(new_new_n9332__), .dout(new_new_n9344__));
  buf1  g6246(.din(new_new_n9344__), .dout(new_new_n9345__));
  buf1  g6247(.din(new_new_n9345__), .dout(new_new_n9346__));
  buf1  g6248(.din(new_new_n9345__), .dout(new_new_n9347__));
  buf1  g6249(.din(new_new_n9344__), .dout(new_new_n9348__));
  buf1  g6250(.din(new_new_n9348__), .dout(new_new_n9349__));
  buf1  g6251(.din(new_new_n9348__), .dout(new_new_n9350__));
  buf1  g6252(.din(new_new_n3688__), .dout(new_new_n9351__));
  buf1  g6253(.din(new_new_n9351__), .dout(new_new_n9352__));
  buf1  g6254(.din(new_new_n9352__), .dout(new_new_n9353__));
  buf1  g6255(.din(new_new_n9353__), .dout(new_new_n9354__));
  buf1  g6256(.din(new_new_n9354__), .dout(new_new_n9355__));
  buf1  g6257(.din(new_new_n9354__), .dout(new_new_n9356__));
  buf1  g6258(.din(new_new_n9353__), .dout(new_new_n9357__));
  buf1  g6259(.din(new_new_n9357__), .dout(new_new_n9358__));
  buf1  g6260(.din(new_new_n9357__), .dout(new_new_n9359__));
  buf1  g6261(.din(new_new_n9352__), .dout(new_new_n9360__));
  buf1  g6262(.din(new_new_n9360__), .dout(new_new_n9361__));
  buf1  g6263(.din(new_new_n9360__), .dout(new_new_n9362__));
  buf1  g6264(.din(new_new_n9351__), .dout(new_new_n9363__));
  buf1  g6265(.din(new_new_n9363__), .dout(new_new_n9364__));
  buf1  g6266(.din(new_new_n9364__), .dout(new_new_n9365__));
  buf1  g6267(.din(new_new_n9364__), .dout(new_new_n9366__));
  buf1  g6268(.din(new_new_n9363__), .dout(new_new_n9367__));
  buf1  g6269(.din(new_new_n9367__), .dout(new_new_n9368__));
  buf1  g6270(.din(new_new_n9367__), .dout(new_new_n9369__));
  buf1  g6271(.din(new_new_n3681__), .dout(new_new_n9370__));
  buf1  g6272(.din(new_new_n9370__), .dout(new_new_n9371__));
  buf1  g6273(.din(new_new_n9371__), .dout(new_new_n9372__));
  buf1  g6274(.din(new_new_n9372__), .dout(new_new_n9373__));
  buf1  g6275(.din(new_new_n9373__), .dout(new_new_n9374__));
  buf1  g6276(.din(new_new_n9373__), .dout(new_new_n9375__));
  buf1  g6277(.din(new_new_n9372__), .dout(new_new_n9376__));
  buf1  g6278(.din(new_new_n9376__), .dout(new_new_n9377__));
  buf1  g6279(.din(new_new_n9376__), .dout(new_new_n9378__));
  buf1  g6280(.din(new_new_n9371__), .dout(new_new_n9379__));
  buf1  g6281(.din(new_new_n9379__), .dout(new_new_n9380__));
  buf1  g6282(.din(new_new_n9379__), .dout(new_new_n9381__));
  buf1  g6283(.din(new_new_n9370__), .dout(new_new_n9382__));
  buf1  g6284(.din(new_new_n9382__), .dout(new_new_n9383__));
  buf1  g6285(.din(new_new_n9383__), .dout(new_new_n9384__));
  buf1  g6286(.din(new_new_n9383__), .dout(new_new_n9385__));
  buf1  g6287(.din(new_new_n9382__), .dout(new_new_n9386__));
  buf1  g6288(.din(new_new_n9386__), .dout(new_new_n9387__));
  buf1  g6289(.din(new_new_n9386__), .dout(new_new_n9388__));
  buf1  g6290(.din(new_new_n3689__), .dout(new_new_n9389__));
  buf1  g6291(.din(new_new_n9389__), .dout(new_new_n9390__));
  buf1  g6292(.din(new_new_n9390__), .dout(new_new_n9391__));
  buf1  g6293(.din(new_new_n9391__), .dout(new_new_n9392__));
  buf1  g6294(.din(new_new_n9392__), .dout(new_new_n9393__));
  buf1  g6295(.din(new_new_n9392__), .dout(new_new_n9394__));
  buf1  g6296(.din(new_new_n9391__), .dout(new_new_n9395__));
  buf1  g6297(.din(new_new_n9395__), .dout(new_new_n9396__));
  buf1  g6298(.din(new_new_n9395__), .dout(new_new_n9397__));
  buf1  g6299(.din(new_new_n9390__), .dout(new_new_n9398__));
  buf1  g6300(.din(new_new_n9398__), .dout(new_new_n9399__));
  buf1  g6301(.din(new_new_n9398__), .dout(new_new_n9400__));
  buf1  g6302(.din(new_new_n9389__), .dout(new_new_n9401__));
  buf1  g6303(.din(new_new_n9401__), .dout(new_new_n9402__));
  buf1  g6304(.din(new_new_n9402__), .dout(new_new_n9403__));
  buf1  g6305(.din(new_new_n9402__), .dout(new_new_n9404__));
  buf1  g6306(.din(new_new_n9401__), .dout(new_new_n9405__));
  buf1  g6307(.din(new_new_n9405__), .dout(new_new_n9406__));
  buf1  g6308(.din(new_new_n9405__), .dout(new_new_n9407__));
  buf1  g6309(.din(new_new_n5267__), .dout(new_new_n9408__));
  buf1  g6310(.din(new_new_n9408__), .dout(new_new_n9409__));
  buf1  g6311(.din(new_new_n9409__), .dout(new_new_n9410__));
  buf1  g6312(.din(new_new_n9408__), .dout(new_new_n9411__));
  buf1  g6313(.din(new_new_n5351__), .dout(new_new_n9412__));
  buf1  g6314(.din(new_new_n9412__), .dout(new_new_n9413__));
  buf1  g6315(.din(new_new_n9413__), .dout(new_new_n9414__));
  buf1  g6316(.din(new_new_n9412__), .dout(new_new_n9415__));
  buf1  g6317(.din(new_new_n2810__), .dout(new_new_n9416__));
  buf1  g6318(.din(new_new_n2794__), .dout(new_new_n9417__));
  buf1  g6319(.din(new_new_n5284__), .dout(new_new_n9418__));
  buf1  g6320(.din(new_new_n9418__), .dout(new_new_n9419__));
  buf1  g6321(.din(new_new_n9419__), .dout(new_new_n9420__));
  buf1  g6322(.din(new_new_n9418__), .dout(new_new_n9421__));
  buf1  g6323(.din(new_new_n5368__), .dout(new_new_n9422__));
  buf1  g6324(.din(new_new_n9422__), .dout(new_new_n9423__));
  buf1  g6325(.din(new_new_n9423__), .dout(new_new_n9424__));
  buf1  g6326(.din(new_new_n9422__), .dout(new_new_n9425__));
  buf1  g6327(.din(new_new_n2898__), .dout(new_new_n9426__));
  buf1  g6328(.din(new_new_n2730__), .dout(new_new_n9427__));
  buf1  g6329(.din(new_new_n5303__), .dout(new_new_n9428__));
  buf1  g6330(.din(new_new_n9428__), .dout(new_new_n9429__));
  buf1  g6331(.din(new_new_n9429__), .dout(new_new_n9430__));
  buf1  g6332(.din(new_new_n9428__), .dout(new_new_n9431__));
  buf1  g6333(.din(new_new_n5387__), .dout(new_new_n9432__));
  buf1  g6334(.din(new_new_n9432__), .dout(new_new_n9433__));
  buf1  g6335(.din(new_new_n9433__), .dout(new_new_n9434__));
  buf1  g6336(.din(new_new_n9432__), .dout(new_new_n9435__));
  buf1  g6337(.din(new_new_n2890__), .dout(new_new_n9436__));
  buf1  g6338(.din(new_new_n2722__), .dout(new_new_n9437__));
  buf1  g6339(.din(new_new_n5182__), .dout(new_new_n9438__));
  buf1  g6340(.din(new_new_n9438__), .dout(new_new_n9439__));
  buf1  g6341(.din(new_new_n9439__), .dout(new_new_n9440__));
  buf1  g6342(.din(new_new_n9438__), .dout(new_new_n9441__));
  buf1  g6343(.din(new_new_n5400__), .dout(new_new_n9442__));
  buf1  g6344(.din(new_new_n9442__), .dout(new_new_n9443__));
  buf1  g6345(.din(new_new_n9443__), .dout(new_new_n9444__));
  buf1  g6346(.din(new_new_n9442__), .dout(new_new_n9445__));
  buf1  g6347(.din(new_new_n2874__), .dout(new_new_n9446__));
  buf1  g6348(.din(new_new_n2882__), .dout(new_new_n9447__));
  buf1  g6349(.din(new_new_n3370__), .dout(new_new_n9448__));
  buf1  g6350(.din(new_new_n3290__), .dout(new_new_n9449__));
  buf1  g6351(.din(new_new_n3338__), .dout(new_new_n9450__));
  buf1  g6352(.din(new_new_n3258__), .dout(new_new_n9451__));
  buf1  g6353(.din(new_new_n3250__), .dout(new_new_n9452__));
  buf1  g6354(.din(new_new_n3242__), .dout(new_new_n9453__));
  buf1  g6355(.din(new_new_n3234__), .dout(new_new_n9454__));
  buf1  g6356(.din(new_new_n3226__), .dout(new_new_n9455__));
  buf1  g6357(.din(new_new_n4792__), .dout(new_new_n9456__));
  buf1  g6358(.din(new_new_n3767__), .dout(new_new_n9457__));
  buf1  g6359(.din(new_new_n3759__), .dout(new_new_n9458__));
  buf1  g6360(.din(new_new_n3902__), .dout(new_new_n9459__));
  buf1  g6361(.din(new_new_n3170__), .dout(new_new_n9460__));
  buf1  g6362(.din(new_new_n3171__), .dout(new_new_n9461__));
  buf1  g6363(.din(new_new_n5792__), .dout(new_new_n9462__));
  buf1  g6364(.din(new_new_n5791__), .dout(new_new_n9463__));
  buf1  g6365(.din(new_new_n5798__), .dout(new_new_n9464__));
  buf1  g6366(.din(new_new_n3766__), .dout(new_new_n9465__));
  buf1  g6367(.din(new_new_n3114__), .dout(new_new_n9466__));
  buf1  g6368(.din(new_new_n3758__), .dout(new_new_n9467__));
  buf1  g6369(.din(new_new_n5220__), .dout(new_new_n9468__));
  buf1  g6370(.din(new_new_n5809__), .dout(new_new_n9469__));
  buf1  g6371(.din(new_new_n3643__), .dout(new_new_n9470__));
  buf1  g6372(.din(new_new_n3627__), .dout(new_new_n9471__));
  buf1  g6373(.din(new_new_n5447__), .dout(new_new_n9472__));
  buf1  g6374(.din(new_new_n3651__), .dout(new_new_n9473__));
  buf1  g6375(.din(new_new_n5494__), .dout(new_new_n9474__));
  buf1  g6376(.din(new_new_n5001__), .dout(new_new_n9475__));
  buf1  g6377(.din(new_new_n5048__), .dout(new_new_n9476__));
  buf1  g6378(.din(new_new_n3427__), .dout(new_new_n9477__));
  buf1  g6379(.din(new_new_n3855__), .dout(new_new_n9478__));
  buf1  g6380(.din(new_new_n3854__), .dout(new_new_n9479__));
  buf1  g6381(.din(new_new_n5820__), .dout(new_new_n9480__));
  buf1  g6382(.din(new_new_n9480__), .dout(new_new_n9481__));
  buf1  g6383(.din(new_new_n9481__), .dout(new_new_n9482__));
  buf1  g6384(.din(new_new_n9480__), .dout(new_new_n9483__));
  buf1  g6385(.din(new_new_n5871__), .dout(new_new_n9484__));
  buf1  g6386(.din(new_new_n9484__), .dout(new_new_n9485__));
  buf1  g6387(.din(new_new_n9485__), .dout(new_new_n9486__));
  buf1  g6388(.din(new_new_n9484__), .dout(new_new_n9487__));
  buf1  g6389(.din(new_new_n3018__), .dout(new_new_n9488__));
  buf1  g6390(.din(new_new_n3010__), .dout(new_new_n9489__));
  buf1  g6391(.din(new_new_n5828__), .dout(new_new_n9490__));
  buf1  g6392(.din(new_new_n9490__), .dout(new_new_n9491__));
  buf1  g6393(.din(new_new_n9491__), .dout(new_new_n9492__));
  buf1  g6394(.din(new_new_n9490__), .dout(new_new_n9493__));
  buf1  g6395(.din(new_new_n5879__), .dout(new_new_n9494__));
  buf1  g6396(.din(new_new_n9494__), .dout(new_new_n9495__));
  buf1  g6397(.din(new_new_n9495__), .dout(new_new_n9496__));
  buf1  g6398(.din(new_new_n9494__), .dout(new_new_n9497__));
  buf1  g6399(.din(new_new_n2818__), .dout(new_new_n9498__));
  buf1  g6400(.din(new_new_n2826__), .dout(new_new_n9499__));
  buf1  g6401(.din(new_new_n5836__), .dout(new_new_n9500__));
  buf1  g6402(.din(new_new_n9500__), .dout(new_new_n9501__));
  buf1  g6403(.din(new_new_n9501__), .dout(new_new_n9502__));
  buf1  g6404(.din(new_new_n9500__), .dout(new_new_n9503__));
  buf1  g6405(.din(new_new_n5887__), .dout(new_new_n9504__));
  buf1  g6406(.din(new_new_n9504__), .dout(new_new_n9505__));
  buf1  g6407(.din(new_new_n9505__), .dout(new_new_n9506__));
  buf1  g6408(.din(new_new_n9504__), .dout(new_new_n9507__));
  buf1  g6409(.din(new_new_n2994__), .dout(new_new_n9508__));
  buf1  g6410(.din(new_new_n3002__), .dout(new_new_n9509__));
  buf1  g6411(.din(new_new_n5844__), .dout(new_new_n9510__));
  buf1  g6412(.din(new_new_n9510__), .dout(new_new_n9511__));
  buf1  g6413(.din(new_new_n9511__), .dout(new_new_n9512__));
  buf1  g6414(.din(new_new_n9510__), .dout(new_new_n9513__));
  buf1  g6415(.din(new_new_n5895__), .dout(new_new_n9514__));
  buf1  g6416(.din(new_new_n9514__), .dout(new_new_n9515__));
  buf1  g6417(.din(new_new_n9515__), .dout(new_new_n9516__));
  buf1  g6418(.din(new_new_n9514__), .dout(new_new_n9517__));
  buf1  g6419(.din(new_new_n2970__), .dout(new_new_n9518__));
  buf1  g6420(.din(new_new_n2802__), .dout(new_new_n9519__));
  buf1  g6421(.din(new_new_n3378__), .dout(new_new_n9520__));
  buf1  g6422(.din(new_new_n3298__), .dout(new_new_n9521__));
  buf1  g6423(.din(new_new_n3362__), .dout(new_new_n9522__));
  buf1  g6424(.din(new_new_n3282__), .dout(new_new_n9523__));
  buf1  g6425(.din(new_new_n3354__), .dout(new_new_n9524__));
  buf1  g6426(.din(new_new_n3274__), .dout(new_new_n9525__));
  buf1  g6427(.din(new_new_n3346__), .dout(new_new_n9526__));
  buf1  g6428(.din(new_new_n3266__), .dout(new_new_n9527__));
  buf1  g6429(.din(new_new_n6082__), .dout(new_new_n9528__));
  buf1  g6430(.din(new_new_n6087__), .dout(new_new_n9529__));
  buf1  g6431(.din(new_new_n6092__), .dout(new_new_n9530__));
  buf1  g6432(.din(new_new_n6098__), .dout(new_new_n9531__));
  buf1  g6433(.din(new_new_n6103__), .dout(new_new_n9532__));
  buf1  g6434(.din(new_new_n6116__), .dout(new_new_n9533__));
  buf1  g6435(.din(new_new_n9533__), .dout(new_new_n9534__));
  buf1  g6436(.din(new_new_n9533__), .dout(new_new_n9535__));
  buf1  g6437(.din(new_new_n6124__), .dout(new_new_n9536__));
  buf1  g6438(.din(new_new_n9536__), .dout(new_new_n9537__));
  buf1  g6439(.din(new_new_n9536__), .dout(new_new_n9538__));
  buf1  g6440(.din(new_new_n2714__), .dout(new_new_n9539__));
  buf1  g6441(.din(new_new_n2866__), .dout(new_new_n9540__));
  buf1  g6442(.din(new_new_n3306__), .dout(new_new_n9541__));
  buf1  g6443(.din(new_new_n3314__), .dout(new_new_n9542__));
  buf1  g6444(.din(new_new_n4461__), .dout(new_new_n9543__));
  buf1  g6445(.din(new_new_n9543__), .dout(new_new_n9544__));
  buf1  g6446(.din(new_new_n9544__), .dout(new_new_n9545__));
  buf1  g6447(.din(new_new_n9544__), .dout(new_new_n9546__));
  buf1  g6448(.din(new_new_n9543__), .dout(new_new_n9547__));
  buf1  g6449(.din(new_new_n9547__), .dout(new_new_n9548__));
  buf1  g6450(.din(new_new_n9547__), .dout(new_new_n9549__));
  buf1  g6451(.din(new_new_n4188__), .dout(new_new_n9550__));
  buf1  g6452(.din(new_new_n9550__), .dout(new_new_n9551__));
  buf1  g6453(.din(new_new_n9551__), .dout(new_new_n9552__));
  buf1  g6454(.din(new_new_n9550__), .dout(new_new_n9553__));
  buf1  g6455(.din(new_new_n4460__), .dout(new_new_n9554__));
  buf1  g6456(.din(new_new_n9554__), .dout(new_new_n9555__));
  buf1  g6457(.din(new_new_n9555__), .dout(new_new_n9556__));
  buf1  g6458(.din(new_new_n9556__), .dout(new_new_n9557__));
  buf1  g6459(.din(new_new_n9555__), .dout(new_new_n9558__));
  buf1  g6460(.din(new_new_n9554__), .dout(new_new_n9559__));
  buf1  g6461(.din(new_new_n9559__), .dout(new_new_n9560__));
  buf1  g6462(.din(new_new_n9559__), .dout(new_new_n9561__));
  buf1  g6463(.din(new_new_n4189__), .dout(new_new_n9562__));
  buf1  g6464(.din(new_new_n9562__), .dout(new_new_n9563__));
  buf1  g6465(.din(new_new_n9562__), .dout(new_new_n9564__));
  buf1  g6466(.din(new_new_n4465__), .dout(new_new_n9565__));
  buf1  g6467(.din(new_new_n9565__), .dout(new_new_n9566__));
  buf1  g6468(.din(new_new_n9566__), .dout(new_new_n9567__));
  buf1  g6469(.din(new_new_n9566__), .dout(new_new_n9568__));
  buf1  g6470(.din(new_new_n9565__), .dout(new_new_n9569__));
  buf1  g6471(.din(new_new_n9569__), .dout(new_new_n9570__));
  buf1  g6472(.din(new_new_n4464__), .dout(new_new_n9571__));
  buf1  g6473(.din(new_new_n9571__), .dout(new_new_n9572__));
  buf1  g6474(.din(new_new_n9572__), .dout(new_new_n9573__));
  buf1  g6475(.din(new_new_n9572__), .dout(new_new_n9574__));
  buf1  g6476(.din(new_new_n9571__), .dout(new_new_n9575__));
  buf1  g6477(.din(new_new_n9575__), .dout(new_new_n9576__));
  buf1  g6478(.din(new_new_n9575__), .dout(new_new_n9577__));
  buf1  g6479(.din(new_new_n4563__), .dout(new_new_n9578__));
  buf1  g6480(.din(new_new_n9578__), .dout(new_new_n9579__));
  buf1  g6481(.din(new_new_n9579__), .dout(new_new_n9580__));
  buf1  g6482(.din(new_new_n9579__), .dout(new_new_n9581__));
  buf1  g6483(.din(new_new_n9578__), .dout(new_new_n9582__));
  buf1  g6484(.din(new_new_n9582__), .dout(new_new_n9583__));
  buf1  g6485(.din(new_new_n9582__), .dout(new_new_n9584__));
  buf1  g6486(.din(new_new_n4546__), .dout(new_new_n9585__));
  buf1  g6487(.din(new_new_n4562__), .dout(new_new_n9586__));
  buf1  g6488(.din(new_new_n9586__), .dout(new_new_n9587__));
  buf1  g6489(.din(new_new_n9587__), .dout(new_new_n9588__));
  buf1  g6490(.din(new_new_n9588__), .dout(new_new_n9589__));
  buf1  g6491(.din(new_new_n9587__), .dout(new_new_n9590__));
  buf1  g6492(.din(new_new_n9586__), .dout(new_new_n9591__));
  buf1  g6493(.din(new_new_n9591__), .dout(new_new_n9592__));
  buf1  g6494(.din(new_new_n9591__), .dout(new_new_n9593__));
  buf1  g6495(.din(new_new_n4547__), .dout(new_new_n9594__));
  buf1  g6496(.din(new_new_n4565__), .dout(new_new_n9595__));
  buf1  g6497(.din(new_new_n9595__), .dout(new_new_n9596__));
  buf1  g6498(.din(new_new_n9596__), .dout(new_new_n9597__));
  buf1  g6499(.din(new_new_n9596__), .dout(new_new_n9598__));
  buf1  g6500(.din(new_new_n9595__), .dout(new_new_n9599__));
  buf1  g6501(.din(new_new_n9599__), .dout(new_new_n9600__));
  buf1  g6502(.din(new_new_n4564__), .dout(new_new_n9601__));
  buf1  g6503(.din(new_new_n9601__), .dout(new_new_n9602__));
  buf1  g6504(.din(new_new_n9602__), .dout(new_new_n9603__));
  buf1  g6505(.din(new_new_n9602__), .dout(new_new_n9604__));
  buf1  g6506(.din(new_new_n9601__), .dout(new_new_n9605__));
  buf1  g6507(.din(new_new_n9605__), .dout(new_new_n9606__));
  buf1  g6508(.din(new_new_n9605__), .dout(new_new_n9607__));
  buf1  g6509(.din(new_new_n3942__), .dout(new_new_n9608__));
  buf1  g6510(.din(new_new_n3943__), .dout(new_new_n9609__));
  buf1  g6511(.din(new_new_n3940__), .dout(new_new_n9610__));
  buf1  g6512(.din(new_new_n9610__), .dout(new_new_n9611__));
  buf1  g6513(.din(new_new_n9611__), .dout(new_new_n9612__));
  buf1  g6514(.din(new_new_n9611__), .dout(new_new_n9613__));
  buf1  g6515(.din(new_new_n9610__), .dout(new_new_n9614__));
  buf1  g6516(.din(new_new_n9614__), .dout(new_new_n9615__));
  buf1  g6517(.din(new_new_n3941__), .dout(new_new_n9616__));
  buf1  g6518(.din(new_new_n9616__), .dout(new_new_n9617__));
  buf1  g6519(.din(new_new_n9617__), .dout(new_new_n9618__));
  buf1  g6520(.din(new_new_n9617__), .dout(new_new_n9619__));
  buf1  g6521(.din(new_new_n9616__), .dout(new_new_n9620__));
  buf1  g6522(.din(new_new_n9620__), .dout(new_new_n9621__));
  buf1  g6523(.din(new_new_n4006__), .dout(new_new_n9622__));
  buf1  g6524(.din(new_new_n9622__), .dout(new_new_n9623__));
  buf1  g6525(.din(new_new_n9623__), .dout(new_new_n9624__));
  buf1  g6526(.din(new_new_n9623__), .dout(new_new_n9625__));
  buf1  g6527(.din(new_new_n9622__), .dout(new_new_n9626__));
  buf1  g6528(.din(new_new_n4007__), .dout(new_new_n9627__));
  buf1  g6529(.din(new_new_n9627__), .dout(new_new_n9628__));
  buf1  g6530(.din(new_new_n9628__), .dout(new_new_n9629__));
  buf1  g6531(.din(new_new_n9628__), .dout(new_new_n9630__));
  buf1  g6532(.din(new_new_n9627__), .dout(new_new_n9631__));
  buf1  g6533(.din(new_new_n4230__), .dout(new_new_n9632__));
  buf1  g6534(.din(new_new_n9632__), .dout(new_new_n9633__));
  buf1  g6535(.din(new_new_n9633__), .dout(new_new_n9634__));
  buf1  g6536(.din(new_new_n9632__), .dout(new_new_n9635__));
  buf1  g6537(.din(new_new_n4231__), .dout(new_new_n9636__));
  buf1  g6538(.din(new_new_n9636__), .dout(new_new_n9637__));
  buf1  g6539(.din(new_new_n9637__), .dout(new_new_n9638__));
  buf1  g6540(.din(new_new_n9636__), .dout(new_new_n9639__));
  buf1  g6541(.din(new_new_n3946__), .dout(new_new_n9640__));
  buf1  g6542(.din(new_new_n3947__), .dout(new_new_n9641__));
  buf1  g6543(.din(new_new_n3944__), .dout(new_new_n9642__));
  buf1  g6544(.din(new_new_n9642__), .dout(new_new_n9643__));
  buf1  g6545(.din(new_new_n9643__), .dout(new_new_n9644__));
  buf1  g6546(.din(new_new_n9643__), .dout(new_new_n9645__));
  buf1  g6547(.din(new_new_n9642__), .dout(new_new_n9646__));
  buf1  g6548(.din(new_new_n9646__), .dout(new_new_n9647__));
  buf1  g6549(.din(new_new_n3945__), .dout(new_new_n9648__));
  buf1  g6550(.din(new_new_n9648__), .dout(new_new_n9649__));
  buf1  g6551(.din(new_new_n9649__), .dout(new_new_n9650__));
  buf1  g6552(.din(new_new_n9649__), .dout(new_new_n9651__));
  buf1  g6553(.din(new_new_n9648__), .dout(new_new_n9652__));
  buf1  g6554(.din(new_new_n9652__), .dout(new_new_n9653__));
  buf1  g6555(.din(new_new_n4012__), .dout(new_new_n9654__));
  buf1  g6556(.din(new_new_n9654__), .dout(new_new_n9655__));
  buf1  g6557(.din(new_new_n9655__), .dout(new_new_n9656__));
  buf1  g6558(.din(new_new_n9655__), .dout(new_new_n9657__));
  buf1  g6559(.din(new_new_n9654__), .dout(new_new_n9658__));
  buf1  g6560(.din(new_new_n4013__), .dout(new_new_n9659__));
  buf1  g6561(.din(new_new_n9659__), .dout(new_new_n9660__));
  buf1  g6562(.din(new_new_n9660__), .dout(new_new_n9661__));
  buf1  g6563(.din(new_new_n9660__), .dout(new_new_n9662__));
  buf1  g6564(.din(new_new_n9659__), .dout(new_new_n9663__));
  buf1  g6565(.din(new_new_n4232__), .dout(new_new_n9664__));
  buf1  g6566(.din(new_new_n9664__), .dout(new_new_n9665__));
  buf1  g6567(.din(new_new_n9665__), .dout(new_new_n9666__));
  buf1  g6568(.din(new_new_n9664__), .dout(new_new_n9667__));
  buf1  g6569(.din(new_new_n4233__), .dout(new_new_n9668__));
  buf1  g6570(.din(new_new_n9668__), .dout(new_new_n9669__));
  buf1  g6571(.din(new_new_n9669__), .dout(new_new_n9670__));
  buf1  g6572(.din(new_new_n9668__), .dout(new_new_n9671__));
  buf1  g6573(.din(new_new_n4088__), .dout(new_new_n9672__));
  buf1  g6574(.din(new_new_n9672__), .dout(new_new_n9673__));
  buf1  g6575(.din(new_new_n9672__), .dout(new_new_n9674__));
  buf1  g6576(.din(new_new_n4082__), .dout(new_new_n9675__));
  buf1  g6577(.din(new_new_n9675__), .dout(new_new_n9676__));
  buf1  g6578(.din(new_new_n9675__), .dout(new_new_n9677__));
  buf1  g6579(.din(new_new_n4089__), .dout(new_new_n9678__));
  buf1  g6580(.din(new_new_n9678__), .dout(new_new_n9679__));
  buf1  g6581(.din(new_new_n4083__), .dout(new_new_n9680__));
  buf1  g6582(.din(new_new_n9680__), .dout(new_new_n9681__));
  buf1  g6583(.din(new_new_n4086__), .dout(new_new_n9682__));
  buf1  g6584(.din(new_new_n9682__), .dout(new_new_n9683__));
  buf1  g6585(.din(new_new_n9682__), .dout(new_new_n9684__));
  buf1  g6586(.din(new_new_n4084__), .dout(new_new_n9685__));
  buf1  g6587(.din(new_new_n9685__), .dout(new_new_n9686__));
  buf1  g6588(.din(new_new_n9685__), .dout(new_new_n9687__));
  buf1  g6589(.din(new_new_n4087__), .dout(new_new_n9688__));
  buf1  g6590(.din(new_new_n9688__), .dout(new_new_n9689__));
  buf1  g6591(.din(new_new_n4085__), .dout(new_new_n9690__));
  buf1  g6592(.din(new_new_n9690__), .dout(new_new_n9691__));
  buf1  g6593(.din(new_new_n3913__), .dout(new_new_n9692__));
  buf1  g6594(.din(new_new_n9692__), .dout(new_new_n9693__));
  buf1  g6595(.din(new_new_n3912__), .dout(new_new_n9694__));
  buf1  g6596(.din(new_new_n9694__), .dout(new_new_n9695__));
  buf1  g6597(.din(new_new_n9694__), .dout(new_new_n9696__));
  buf1  g6598(.din(new_new_n4482__), .dout(new_new_n9697__));
  buf1  g6599(.din(new_new_n4480__), .dout(new_new_n9698__));
  buf1  g6600(.din(new_new_n4134__), .dout(new_new_n9699__));
  buf1  g6601(.din(new_new_n3496__), .dout(new_new_n9700__));
  buf1  g6602(.din(new_new_n9700__), .dout(new_new_n9701__));
  buf1  g6603(.din(new_new_n9701__), .dout(new_new_n9702__));
  buf1  g6604(.din(new_new_n9700__), .dout(new_new_n9703__));
  buf1  g6605(.din(new_new_n3497__), .dout(new_new_n9704__));
  buf1  g6606(.din(new_new_n4099__), .dout(new_new_n9705__));
  buf1  g6607(.din(new_new_n4136__), .dout(new_new_n9706__));
  buf1  g6608(.din(new_new_n3408__), .dout(new_new_n9707__));
  buf1  g6609(.din(new_new_n9707__), .dout(new_new_n9708__));
  buf1  g6610(.din(new_new_n9708__), .dout(new_new_n9709__));
  buf1  g6611(.din(new_new_n9707__), .dout(new_new_n9710__));
  buf1  g6612(.din(new_new_n3409__), .dout(new_new_n9711__));
  buf1  g6613(.din(new_new_n4101__), .dout(new_new_n9712__));
  buf1  g6614(.din(new_new_n4688__), .dout(new_new_n9713__));
  buf1  g6615(.din(new_new_n4504__), .dout(new_new_n9714__));
  buf1  g6616(.din(new_new_n9714__), .dout(new_new_n9715__));
  buf1  g6617(.din(new_new_n4505__), .dout(new_new_n9716__));
  buf1  g6618(.din(new_new_n4690__), .dout(new_new_n9717__));
  buf1  g6619(.din(new_new_n4257__), .dout(new_new_n9718__));
  buf1  g6620(.din(new_new_n4256__), .dout(new_new_n9719__));
  buf1  g6621(.din(new_new_n9719__), .dout(new_new_n9720__));
  buf1  g6622(.din(new_new_n3982__), .dout(new_new_n9721__));
  buf1  g6623(.din(new_new_n9721__), .dout(new_new_n9722__));
  buf1  g6624(.din(new_new_n9721__), .dout(new_new_n9723__));
  buf1  g6625(.din(new_new_n3976__), .dout(new_new_n9724__));
  buf1  g6626(.din(new_new_n9724__), .dout(new_new_n9725__));
  buf1  g6627(.din(new_new_n9725__), .dout(new_new_n9726__));
  buf1  g6628(.din(new_new_n9725__), .dout(new_new_n9727__));
  buf1  g6629(.din(new_new_n9724__), .dout(new_new_n9728__));
  buf1  g6630(.din(new_new_n9728__), .dout(new_new_n9729__));
  buf1  g6631(.din(new_new_n3974__), .dout(new_new_n9730__));
  buf1  g6632(.din(new_new_n9730__), .dout(new_new_n9731__));
  buf1  g6633(.din(new_new_n3962__), .dout(new_new_n9732__));
  buf1  g6634(.din(new_new_n9732__), .dout(new_new_n9733__));
  buf1  g6635(.din(new_new_n9733__), .dout(new_new_n9734__));
  buf1  g6636(.din(new_new_n9733__), .dout(new_new_n9735__));
  buf1  g6637(.din(new_new_n9732__), .dout(new_new_n9736__));
  buf1  g6638(.din(new_new_n3973__), .dout(new_new_n9737__));
  buf1  g6639(.din(new_new_n9737__), .dout(new_new_n9738__));
  buf1  g6640(.din(new_new_n3965__), .dout(new_new_n9739__));
  buf1  g6641(.din(new_new_n9739__), .dout(new_new_n9740__));
  buf1  g6642(.din(new_new_n9740__), .dout(new_new_n9741__));
  buf1  g6643(.din(new_new_n9740__), .dout(new_new_n9742__));
  buf1  g6644(.din(new_new_n9739__), .dout(new_new_n9743__));
  buf1  g6645(.din(new_new_n3981__), .dout(new_new_n9744__));
  buf1  g6646(.din(new_new_n3979__), .dout(new_new_n9745__));
  buf1  g6647(.din(new_new_n9745__), .dout(new_new_n9746__));
  buf1  g6648(.din(new_new_n9746__), .dout(new_new_n9747__));
  buf1  g6649(.din(new_new_n9745__), .dout(new_new_n9748__));
  buf1  g6650(.din(new_new_n4676__), .dout(new_new_n9749__));
  buf1  g6651(.din(new_new_n4672__), .dout(new_new_n9750__));
  buf1  g6652(.din(new_new_n4680__), .dout(new_new_n9751__));
  buf1  g6653(.din(new_new_n4668__), .dout(new_new_n9752__));
  buf1  g6654(.din(new_new_n4004__), .dout(new_new_n9753__));
  buf1  g6655(.din(new_new_n9753__), .dout(new_new_n9754__));
  buf1  g6656(.din(new_new_n3991__), .dout(new_new_n9755__));
  buf1  g6657(.din(new_new_n9755__), .dout(new_new_n9756__));
  buf1  g6658(.din(new_new_n9755__), .dout(new_new_n9757__));
  buf1  g6659(.din(new_new_n4005__), .dout(new_new_n9758__));
  buf1  g6660(.din(new_new_n3990__), .dout(new_new_n9759__));
  buf1  g6661(.din(new_new_n9759__), .dout(new_new_n9760__));
  buf1  g6662(.din(new_new_n9760__), .dout(new_new_n9761__));
  buf1  g6663(.din(new_new_n9760__), .dout(new_new_n9762__));
  buf1  g6664(.din(new_new_n9759__), .dout(new_new_n9763__));
  buf1  g6665(.din(new_new_n3963__), .dout(new_new_n9764__));
  buf1  g6666(.din(new_new_n9764__), .dout(new_new_n9765__));
  buf1  g6667(.din(new_new_n9764__), .dout(new_new_n9766__));
  buf1  g6668(.din(new_new_n3975__), .dout(new_new_n9767__));
  buf1  g6669(.din(new_new_n3972__), .dout(new_new_n9768__));
  buf1  g6670(.din(new_new_n9768__), .dout(new_new_n9769__));
  buf1  g6671(.din(new_new_n9768__), .dout(new_new_n9770__));
  buf1  g6672(.din(new_new_n3964__), .dout(new_new_n9771__));
  buf1  g6673(.din(new_new_n9771__), .dout(new_new_n9772__));
  buf1  g6674(.din(new_new_n9772__), .dout(new_new_n9773__));
  buf1  g6675(.din(new_new_n9772__), .dout(new_new_n9774__));
  buf1  g6676(.din(new_new_n9771__), .dout(new_new_n9775__));
  buf1  g6677(.din(new_new_n4692__), .dout(new_new_n9776__));
  buf1  g6678(.din(new_new_n9776__), .dout(new_new_n9777__));
  buf1  g6679(.din(new_new_n9777__), .dout(new_new_n9778__));
  buf1  g6680(.din(new_new_n9776__), .dout(new_new_n9779__));
  buf1  g6681(.din(new_new_n4686__), .dout(new_new_n9780__));
  buf1  g6682(.din(new_new_n9780__), .dout(new_new_n9781__));
  buf1  g6683(.din(new_new_n9781__), .dout(new_new_n9782__));
  buf1  g6684(.din(new_new_n9780__), .dout(new_new_n9783__));
  buf1  g6685(.din(new_new_n4693__), .dout(new_new_n9784__));
  buf1  g6686(.din(new_new_n9784__), .dout(new_new_n9785__));
  buf1  g6687(.din(new_new_n9784__), .dout(new_new_n9786__));
  buf1  g6688(.din(new_new_n4687__), .dout(new_new_n9787__));
  buf1  g6689(.din(new_new_n9787__), .dout(new_new_n9788__));
  buf1  g6690(.din(new_new_n9787__), .dout(new_new_n9789__));
  buf1  g6691(.din(new_new_n4702__), .dout(new_new_n9790__));
  buf1  g6692(.din(new_new_n4699__), .dout(new_new_n9791__));
  buf1  g6693(.din(new_new_n4703__), .dout(new_new_n9792__));
  buf1  g6694(.din(new_new_n4698__), .dout(new_new_n9793__));
  buf1  g6695(.din(new_new_n4704__), .dout(new_new_n9794__));
  buf1  g6696(.din(new_new_n4701__), .dout(new_new_n9795__));
  buf1  g6697(.din(new_new_n4705__), .dout(new_new_n9796__));
  buf1  g6698(.din(new_new_n4700__), .dout(new_new_n9797__));
  buf1  g6699(.din(new_new_n4706__), .dout(new_new_n9798__));
  buf1  g6700(.din(new_new_n4695__), .dout(new_new_n9799__));
  buf1  g6701(.din(new_new_n4707__), .dout(new_new_n9800__));
  buf1  g6702(.din(new_new_n4694__), .dout(new_new_n9801__));
  buf1  g6703(.din(new_new_n4708__), .dout(new_new_n9802__));
  buf1  g6704(.din(new_new_n4697__), .dout(new_new_n9803__));
  buf1  g6705(.din(new_new_n4709__), .dout(new_new_n9804__));
  buf1  g6706(.din(new_new_n4696__), .dout(new_new_n9805__));
  buf1  g6707(.din(new_new_n4674__), .dout(new_new_n9806__));
  buf1  g6708(.din(new_new_n4670__), .dout(new_new_n9807__));
  buf1  g6709(.din(new_new_n4678__), .dout(new_new_n9808__));
  buf1  g6710(.din(new_new_n4666__), .dout(new_new_n9809__));
  buf1  g6711(.din(new_new_n3504__), .dout(new_new_n9810__));
  buf1  g6712(.din(new_new_n4506__), .dout(new_new_n9811__));
  buf1  g6713(.din(new_new_n3440__), .dout(new_new_n9812__));
  buf1  g6714(.din(new_new_n4258__), .dout(new_new_n9813__));
  buf1  g6715(.din(new_new_n4252__), .dout(new_new_n9814__));
  buf1  g6716(.din(new_new_n9814__), .dout(new_new_n9815__));
  buf1  g6717(.din(new_new_n9815__), .dout(new_new_n9816__));
  buf1  g6718(.din(new_new_n9815__), .dout(new_new_n9817__));
  buf1  g6719(.din(new_new_n9814__), .dout(new_new_n9818__));
  buf1  g6720(.din(new_new_n9818__), .dout(new_new_n9819__));
  buf1  g6721(.din(new_new_n3482__), .dout(new_new_n9820__));
  buf1  g6722(.din(new_new_n4253__), .dout(new_new_n9821__));
  buf1  g6723(.din(new_new_n9821__), .dout(new_new_n9822__));
  buf1  g6724(.din(new_new_n9822__), .dout(new_new_n9823__));
  buf1  g6725(.din(new_new_n9821__), .dout(new_new_n9824__));
  buf1  g6726(.din(new_new_n4254__), .dout(new_new_n9825__));
  buf1  g6727(.din(new_new_n9825__), .dout(new_new_n9826__));
  buf1  g6728(.din(new_new_n9826__), .dout(new_new_n9827__));
  buf1  g6729(.din(new_new_n9826__), .dout(new_new_n9828__));
  buf1  g6730(.din(new_new_n9825__), .dout(new_new_n9829__));
  buf1  g6731(.din(new_new_n9829__), .dout(new_new_n9830__));
  buf1  g6732(.din(new_new_n3394__), .dout(new_new_n9831__));
  buf1  g6733(.din(new_new_n4255__), .dout(new_new_n9832__));
  buf1  g6734(.din(new_new_n9832__), .dout(new_new_n9833__));
  buf1  g6735(.din(new_new_n9833__), .dout(new_new_n9834__));
  buf1  g6736(.din(new_new_n9832__), .dout(new_new_n9835__));
  buf1  g6737(.din(new_new_n6384__), .dout(new_new_n9836__));
  buf1  g6738(.din(new_new_n6169__), .dout(new_new_n9837__));
  buf1  g6739(.din(new_new_n9837__), .dout(new_new_n9838__));
  buf1  g6740(.din(new_new_n9837__), .dout(new_new_n9839__));
  buf1  g6741(.din(new_new_n6385__), .dout(new_new_n9840__));
  buf1  g6742(.din(new_new_n6170__), .dout(new_new_n9841__));
  buf1  g6743(.din(new_new_n9841__), .dout(new_new_n9842__));
  buf1  g6744(.din(new_new_n9842__), .dout(new_new_n9843__));
  buf1  g6745(.din(new_new_n9841__), .dout(new_new_n9844__));
  buf1  g6746(.din(new_new_n4040__), .dout(new_new_n9845__));
  buf1  g6747(.din(new_new_n9845__), .dout(new_new_n9846__));
  buf1  g6748(.din(new_new_n4041__), .dout(new_new_n9847__));
  buf1  g6749(.din(new_new_n6394__), .dout(new_new_n9848__));
  buf1  g6750(.din(new_new_n6236__), .dout(new_new_n9849__));
  buf1  g6751(.din(new_new_n9849__), .dout(new_new_n9850__));
  buf1  g6752(.din(new_new_n3656__), .dout(new_new_n9851__));
  buf1  g6753(.din(new_new_n9851__), .dout(new_new_n9852__));
  buf1  g6754(.din(new_new_n6401__), .dout(new_new_n9853__));
  buf1  g6755(.din(new_new_n6402__), .dout(new_new_n9854__));
  buf1  g6756(.din(new_new_n6411__), .dout(new_new_n9855__));
  buf1  g6757(.din(new_new_n6235__), .dout(new_new_n9856__));
  buf1  g6758(.din(new_new_n6197__), .dout(new_new_n9857__));
  buf1  g6759(.din(new_new_n3657__), .dout(new_new_n9858__));
  buf1  g6760(.din(new_new_n9858__), .dout(new_new_n9859__));
  buf1  g6761(.din(new_new_n6423__), .dout(new_new_n9860__));
  buf1  g6762(.din(new_new_n6424__), .dout(new_new_n9861__));
  buf1  g6763(.din(new_new_n6439__), .dout(new_new_n9862__));
  buf1  g6764(.din(new_new_n6440__), .dout(new_new_n9863__));
  buf1  g6765(.din(new_new_n6456__), .dout(new_new_n9864__));
  buf1  g6766(.din(new_new_n4578__), .dout(new_new_n9865__));
  buf1  g6767(.din(new_new_n9865__), .dout(new_new_n9866__));
  buf1  g6768(.din(new_new_n9866__), .dout(new_new_n9867__));
  buf1  g6769(.din(new_new_n9867__), .dout(new_new_n9868__));
  buf1  g6770(.din(new_new_n9867__), .dout(new_new_n9869__));
  buf1  g6771(.din(new_new_n9866__), .dout(new_new_n9870__));
  buf1  g6772(.din(new_new_n9865__), .dout(new_new_n9871__));
  buf1  g6773(.din(new_new_n9871__), .dout(new_new_n9872__));
  buf1  g6774(.din(new_new_n9871__), .dout(new_new_n9873__));
  buf1  g6775(.din(new_new_n6457__), .dout(new_new_n9874__));
  buf1  g6776(.din(new_new_n4579__), .dout(new_new_n9875__));
  buf1  g6777(.din(new_new_n9875__), .dout(new_new_n9876__));
  buf1  g6778(.din(new_new_n9875__), .dout(new_new_n9877__));
  buf1  g6779(.din(new_new_n4042__), .dout(new_new_n9878__));
  buf1  g6780(.din(new_new_n9878__), .dout(new_new_n9879__));
  buf1  g6781(.din(new_new_n4043__), .dout(new_new_n9880__));
  buf1  g6782(.din(new_new_n6466__), .dout(new_new_n9881__));
  buf1  g6783(.din(new_new_n6265__), .dout(new_new_n9882__));
  buf1  g6784(.din(new_new_n3695__), .dout(new_new_n9883__));
  buf1  g6785(.din(new_new_n9883__), .dout(new_new_n9884__));
  buf1  g6786(.din(new_new_n6473__), .dout(new_new_n9885__));
  buf1  g6787(.din(new_new_n6474__), .dout(new_new_n9886__));
  buf1  g6788(.din(new_new_n6483__), .dout(new_new_n9887__));
  buf1  g6789(.din(new_new_n6266__), .dout(new_new_n9888__));
  buf1  g6790(.din(new_new_n9888__), .dout(new_new_n9889__));
  buf1  g6791(.din(new_new_n6205__), .dout(new_new_n9890__));
  buf1  g6792(.din(new_new_n3694__), .dout(new_new_n9891__));
  buf1  g6793(.din(new_new_n9891__), .dout(new_new_n9892__));
  buf1  g6794(.din(new_new_n6495__), .dout(new_new_n9893__));
  buf1  g6795(.din(new_new_n6496__), .dout(new_new_n9894__));
  buf1  g6796(.din(new_new_n6511__), .dout(new_new_n9895__));
  buf1  g6797(.din(new_new_n6512__), .dout(new_new_n9896__));
  buf1  g6798(.din(new_new_n3977__), .dout(new_new_n9897__));
  buf1  g6799(.din(new_new_n9897__), .dout(new_new_n9898__));
  buf1  g6800(.din(new_new_n9897__), .dout(new_new_n9899__));
  buf1  g6801(.din(new_new_n3983__), .dout(new_new_n9900__));
  buf1  g6802(.din(new_new_n4228__), .dout(new_new_n9901__));
  buf1  g6803(.din(new_new_n9901__), .dout(new_new_n9902__));
  buf1  g6804(.din(new_new_n4229__), .dout(new_new_n9903__));
  buf1  g6805(.din(new_new_n3980__), .dout(new_new_n9904__));
  buf1  g6806(.din(new_new_n9904__), .dout(new_new_n9905__));
  buf1  g6807(.din(new_new_n9904__), .dout(new_new_n9906__));
  buf1  g6808(.din(new_new_n3978__), .dout(new_new_n9907__));
  buf1  g6809(.din(new_new_n9907__), .dout(new_new_n9908__));
  buf1  g6810(.din(new_new_n9908__), .dout(new_new_n9909__));
  buf1  g6811(.din(new_new_n9908__), .dout(new_new_n9910__));
  buf1  g6812(.din(new_new_n9907__), .dout(new_new_n9911__));
  buf1  g6813(.din(new_new_n3382__), .dout(new_new_n9912__));
  buf1  g6814(.din(new_new_n9912__), .dout(new_new_n9913__));
  buf1  g6815(.din(new_new_n9913__), .dout(new_new_n9914__));
  buf1  g6816(.din(new_new_n9912__), .dout(new_new_n9915__));
  buf1  g6817(.din(new_new_n3564__), .dout(new_new_n9916__));
  buf1  g6818(.din(new_new_n9916__), .dout(new_new_n9917__));
  buf1  g6819(.din(new_new_n9916__), .dout(new_new_n9918__));
  buf1  g6820(.din(new_new_n6294__), .dout(new_new_n9919__));
  buf1  g6821(.din(new_new_n3592__), .dout(new_new_n9920__));
  buf1  g6822(.din(new_new_n9920__), .dout(new_new_n9921__));
  buf1  g6823(.din(new_new_n9920__), .dout(new_new_n9922__));
  buf1  g6824(.din(new_new_n6288__), .dout(new_new_n9923__));
  buf1  g6825(.din(new_new_n3488__), .dout(new_new_n9924__));
  buf1  g6826(.din(new_new_n3400__), .dout(new_new_n9925__));
  buf1  g6827(.din(new_new_n3918__), .dout(new_new_n9926__));
  buf1  g6828(.din(new_new_n9926__), .dout(new_new_n9927__));
  buf1  g6829(.din(new_new_n9926__), .dout(new_new_n9928__));
  buf1  g6830(.din(new_new_n3916__), .dout(new_new_n9929__));
  buf1  g6831(.din(new_new_n9929__), .dout(new_new_n9930__));
  buf1  g6832(.din(new_new_n9930__), .dout(new_new_n9931__));
  buf1  g6833(.din(new_new_n9930__), .dout(new_new_n9932__));
  buf1  g6834(.din(new_new_n9929__), .dout(new_new_n9933__));
  buf1  g6835(.din(new_new_n3970__), .dout(new_new_n9934__));
  buf1  g6836(.din(new_new_n9934__), .dout(new_new_n9935__));
  buf1  g6837(.din(new_new_n9934__), .dout(new_new_n9936__));
  buf1  g6838(.din(new_new_n3960__), .dout(new_new_n9937__));
  buf1  g6839(.din(new_new_n9937__), .dout(new_new_n9938__));
  buf1  g6840(.din(new_new_n9937__), .dout(new_new_n9939__));
  buf1  g6841(.din(new_new_n3908__), .dout(new_new_n9940__));
  buf1  g6842(.din(new_new_n9940__), .dout(new_new_n9941__));
  buf1  g6843(.din(new_new_n9940__), .dout(new_new_n9942__));
  buf1  g6844(.din(new_new_n3894__), .dout(new_new_n9943__));
  buf1  g6845(.din(new_new_n9943__), .dout(new_new_n9944__));
  buf1  g6846(.din(new_new_n9944__), .dout(new_new_n9945__));
  buf1  g6847(.din(new_new_n9944__), .dout(new_new_n9946__));
  buf1  g6848(.din(new_new_n9943__), .dout(new_new_n9947__));
  buf1  g6849(.din(new_new_n3910__), .dout(new_new_n9948__));
  buf1  g6850(.din(new_new_n9948__), .dout(new_new_n9949__));
  buf1  g6851(.din(new_new_n9948__), .dout(new_new_n9950__));
  buf1  g6852(.din(new_new_n3896__), .dout(new_new_n9951__));
  buf1  g6853(.din(new_new_n9951__), .dout(new_new_n9952__));
  buf1  g6854(.din(new_new_n9952__), .dout(new_new_n9953__));
  buf1  g6855(.din(new_new_n9952__), .dout(new_new_n9954__));
  buf1  g6856(.din(new_new_n9951__), .dout(new_new_n9955__));
  buf1  g6857(.din(new_new_n3968__), .dout(new_new_n9956__));
  buf1  g6858(.din(new_new_n9956__), .dout(new_new_n9957__));
  buf1  g6859(.din(new_new_n3966__), .dout(new_new_n9958__));
  buf1  g6860(.din(new_new_n9958__), .dout(new_new_n9959__));
  buf1  g6861(.din(new_new_n9959__), .dout(new_new_n9960__));
  buf1  g6862(.din(new_new_n9958__), .dout(new_new_n9961__));
  buf1  g6863(.din(new_new_n3904__), .dout(new_new_n9962__));
  buf1  g6864(.din(new_new_n9962__), .dout(new_new_n9963__));
  buf1  g6865(.din(new_new_n3898__), .dout(new_new_n9964__));
  buf1  g6866(.din(new_new_n9964__), .dout(new_new_n9965__));
  buf1  g6867(.din(new_new_n9965__), .dout(new_new_n9966__));
  buf1  g6868(.din(new_new_n9965__), .dout(new_new_n9967__));
  buf1  g6869(.din(new_new_n9964__), .dout(new_new_n9968__));
  buf1  g6870(.din(new_new_n3906__), .dout(new_new_n9969__));
  buf1  g6871(.din(new_new_n9969__), .dout(new_new_n9970__));
  buf1  g6872(.din(new_new_n3900__), .dout(new_new_n9971__));
  buf1  g6873(.din(new_new_n9971__), .dout(new_new_n9972__));
  buf1  g6874(.din(new_new_n9972__), .dout(new_new_n9973__));
  buf1  g6875(.din(new_new_n9972__), .dout(new_new_n9974__));
  buf1  g6876(.din(new_new_n9971__), .dout(new_new_n9975__));
  buf1  g6877(.din(new_new_n3870__), .dout(new_new_n9976__));
  buf1  g6878(.din(new_new_n3868__), .dout(new_new_n9977__));
  buf1  g6879(.din(new_new_n3885__), .dout(new_new_n9978__));
  buf1  g6880(.din(new_new_n9978__), .dout(new_new_n9979__));
  buf1  g6881(.din(new_new_n9979__), .dout(new_new_n9980__));
  buf1  g6882(.din(new_new_n9978__), .dout(new_new_n9981__));
  buf1  g6883(.din(new_new_n3456__), .dout(new_new_n9982__));
  buf1  g6884(.din(new_new_n3884__), .dout(new_new_n9983__));
  buf1  g6885(.din(new_new_n9983__), .dout(new_new_n9984__));
  buf1  g6886(.din(new_new_n9984__), .dout(new_new_n9985__));
  buf1  g6887(.din(new_new_n9984__), .dout(new_new_n9986__));
  buf1  g6888(.din(new_new_n9983__), .dout(new_new_n9987__));
  buf1  g6889(.din(new_new_n3457__), .dout(new_new_n9988__));
  buf1  g6890(.din(new_new_n3876__), .dout(new_new_n9989__));
  buf1  g6891(.din(new_new_n3872__), .dout(new_new_n9990__));
  buf1  g6892(.din(new_new_n3524__), .dout(new_new_n9991__));
  buf1  g6893(.din(new_new_n6314__), .dout(new_new_n9992__));
  buf1  g6894(.din(new_new_n9992__), .dout(new_new_n9993__));
  buf1  g6895(.din(new_new_n9992__), .dout(new_new_n9994__));
  buf1  g6896(.din(new_new_n6301__), .dout(new_new_n9995__));
  buf1  g6897(.din(new_new_n6571__), .dout(new_new_n9996__));
  buf1  g6898(.din(new_new_n9996__), .dout(new_new_n9997__));
  buf1  g6899(.din(new_new_n6311__), .dout(new_new_n9998__));
  buf1  g6900(.din(new_new_n9998__), .dout(new_new_n9999__));
  buf1  g6901(.din(new_new_n9999__), .dout(new_new_n10000__));
  buf1  g6902(.din(new_new_n9998__), .dout(new_new_n10001__));
  buf1  g6903(.din(new_new_n6302__), .dout(new_new_n10002__));
  buf1  g6904(.din(new_new_n10002__), .dout(new_new_n10003__));
  buf1  g6905(.din(new_new_n6303__), .dout(new_new_n10004__));
  buf1  g6906(.din(new_new_n10004__), .dout(new_new_n10005__));
  buf1  g6907(.din(new_new_n4030__), .dout(new_new_n10006__));
  buf1  g6908(.din(new_new_n10006__), .dout(new_new_n10007__));
  buf1  g6909(.din(new_new_n10007__), .dout(new_new_n10008__));
  buf1  g6910(.din(new_new_n10007__), .dout(new_new_n10009__));
  buf1  g6911(.din(new_new_n10006__), .dout(new_new_n10010__));
  buf1  g6912(.din(new_new_n10010__), .dout(new_new_n10011__));
  buf1  g6913(.din(new_new_n10010__), .dout(new_new_n10012__));
  buf1  g6914(.din(new_new_n6304__), .dout(new_new_n10013__));
  buf1  g6915(.din(new_new_n6576__), .dout(new_new_n10014__));
  buf1  g6916(.din(new_new_n10014__), .dout(new_new_n10015__));
  buf1  g6917(.din(new_new_n3905__), .dout(new_new_n10016__));
  buf1  g6918(.din(new_new_n3907__), .dout(new_new_n10017__));
  buf1  g6919(.din(new_new_n6583__), .dout(new_new_n10018__));
  buf1  g6920(.din(new_new_n3924__), .dout(new_new_n10019__));
  buf1  g6921(.din(new_new_n10019__), .dout(new_new_n10020__));
  buf1  g6922(.din(new_new_n10019__), .dout(new_new_n10021__));
  buf1  g6923(.din(new_new_n6532__), .dout(new_new_n10022__));
  buf1  g6924(.din(new_new_n6320__), .dout(new_new_n10023__));
  buf1  g6925(.din(new_new_n10023__), .dout(new_new_n10024__));
  buf1  g6926(.din(new_new_n6588__), .dout(new_new_n10025__));
  buf1  g6927(.din(new_new_n6526__), .dout(new_new_n10026__));
  buf1  g6928(.din(new_new_n6592__), .dout(new_new_n10027__));
  buf1  g6929(.din(new_new_n6573__), .dout(new_new_n10028__));
  buf1  g6930(.din(new_new_n6379__), .dout(new_new_n10029__));
  buf1  g6931(.din(new_new_n6572__), .dout(new_new_n10030__));
  buf1  g6932(.din(new_new_n6575__), .dout(new_new_n10031__));
  buf1  g6933(.din(new_new_n6578__), .dout(new_new_n10032__));
  buf1  g6934(.din(new_new_n4036__), .dout(new_new_n10033__));
  buf1  g6935(.din(new_new_n3928__), .dout(new_new_n10034__));
  buf1  g6936(.din(new_new_n3917__), .dout(new_new_n10035__));
  buf1  g6937(.din(new_new_n10035__), .dout(new_new_n10036__));
  buf1  g6938(.din(new_new_n10035__), .dout(new_new_n10037__));
  buf1  g6939(.din(new_new_n3961__), .dout(new_new_n10038__));
  buf1  g6940(.din(new_new_n3895__), .dout(new_new_n10039__));
  buf1  g6941(.din(new_new_n10039__), .dout(new_new_n10040__));
  buf1  g6942(.din(new_new_n10039__), .dout(new_new_n10041__));
  buf1  g6943(.din(new_new_n3897__), .dout(new_new_n10042__));
  buf1  g6944(.din(new_new_n10042__), .dout(new_new_n10043__));
  buf1  g6945(.din(new_new_n10042__), .dout(new_new_n10044__));
  buf1  g6946(.din(new_new_n3967__), .dout(new_new_n10045__));
  buf1  g6947(.din(new_new_n10045__), .dout(new_new_n10046__));
  buf1  g6948(.din(new_new_n3969__), .dout(new_new_n10047__));
  buf1  g6949(.din(new_new_n3899__), .dout(new_new_n10048__));
  buf1  g6950(.din(new_new_n10048__), .dout(new_new_n10049__));
  buf1  g6951(.din(new_new_n10048__), .dout(new_new_n10050__));
  buf1  g6952(.din(new_new_n3901__), .dout(new_new_n10051__));
  buf1  g6953(.din(new_new_n10051__), .dout(new_new_n10052__));
  buf1  g6954(.din(new_new_n10051__), .dout(new_new_n10053__));
  buf1  g6955(.din(new_new_n4459__), .dout(new_new_n10054__));
  buf1  g6956(.din(new_new_n10054__), .dout(new_new_n10055__));
  buf1  g6957(.din(new_new_n10055__), .dout(new_new_n10056__));
  buf1  g6958(.din(new_new_n10055__), .dout(new_new_n10057__));
  buf1  g6959(.din(new_new_n10054__), .dout(new_new_n10058__));
  buf1  g6960(.din(new_new_n4458__), .dout(new_new_n10059__));
  buf1  g6961(.din(new_new_n10059__), .dout(new_new_n10060__));
  buf1  g6962(.din(new_new_n10060__), .dout(new_new_n10061__));
  buf1  g6963(.din(new_new_n10060__), .dout(new_new_n10062__));
  buf1  g6964(.din(new_new_n10059__), .dout(new_new_n10063__));
  buf1  g6965(.din(new_new_n10063__), .dout(new_new_n10064__));
  buf1  g6966(.din(new_new_n4521__), .dout(new_new_n10065__));
  buf1  g6967(.din(new_new_n4520__), .dout(new_new_n10066__));
  buf1  g6968(.din(new_new_n4463__), .dout(new_new_n10067__));
  buf1  g6969(.din(new_new_n10067__), .dout(new_new_n10068__));
  buf1  g6970(.din(new_new_n10068__), .dout(new_new_n10069__));
  buf1  g6971(.din(new_new_n10068__), .dout(new_new_n10070__));
  buf1  g6972(.din(new_new_n10067__), .dout(new_new_n10071__));
  buf1  g6973(.din(new_new_n4462__), .dout(new_new_n10072__));
  buf1  g6974(.din(new_new_n10072__), .dout(new_new_n10073__));
  buf1  g6975(.din(new_new_n10073__), .dout(new_new_n10074__));
  buf1  g6976(.din(new_new_n10073__), .dout(new_new_n10075__));
  buf1  g6977(.din(new_new_n10072__), .dout(new_new_n10076__));
  buf1  g6978(.din(new_new_n10076__), .dout(new_new_n10077__));
  buf1  g6979(.din(new_new_n4561__), .dout(new_new_n10078__));
  buf1  g6980(.din(new_new_n10078__), .dout(new_new_n10079__));
  buf1  g6981(.din(new_new_n10079__), .dout(new_new_n10080__));
  buf1  g6982(.din(new_new_n10079__), .dout(new_new_n10081__));
  buf1  g6983(.din(new_new_n10078__), .dout(new_new_n10082__));
  buf1  g6984(.din(new_new_n10082__), .dout(new_new_n10083__));
  buf1  g6985(.din(new_new_n10082__), .dout(new_new_n10084__));
  buf1  g6986(.din(new_new_n3951__), .dout(new_new_n10085__));
  buf1  g6987(.din(new_new_n4560__), .dout(new_new_n10086__));
  buf1  g6988(.din(new_new_n10086__), .dout(new_new_n10087__));
  buf1  g6989(.din(new_new_n10087__), .dout(new_new_n10088__));
  buf1  g6990(.din(new_new_n10088__), .dout(new_new_n10089__));
  buf1  g6991(.din(new_new_n10087__), .dout(new_new_n10090__));
  buf1  g6992(.din(new_new_n10086__), .dout(new_new_n10091__));
  buf1  g6993(.din(new_new_n10091__), .dout(new_new_n10092__));
  buf1  g6994(.din(new_new_n10091__), .dout(new_new_n10093__));
  buf1  g6995(.din(new_new_n3950__), .dout(new_new_n10094__));
  buf1  g6996(.din(new_new_n10094__), .dout(new_new_n10095__));
  buf1  g6997(.din(new_new_n10095__), .dout(new_new_n10096__));
  buf1  g6998(.din(new_new_n10094__), .dout(new_new_n10097__));
  buf1  g6999(.din(new_new_n4567__), .dout(new_new_n10098__));
  buf1  g7000(.din(new_new_n10098__), .dout(new_new_n10099__));
  buf1  g7001(.din(new_new_n10099__), .dout(new_new_n10100__));
  buf1  g7002(.din(new_new_n10099__), .dout(new_new_n10101__));
  buf1  g7003(.din(new_new_n10098__), .dout(new_new_n10102__));
  buf1  g7004(.din(new_new_n10102__), .dout(new_new_n10103__));
  buf1  g7005(.din(new_new_n10102__), .dout(new_new_n10104__));
  buf1  g7006(.din(new_new_n4566__), .dout(new_new_n10105__));
  buf1  g7007(.din(new_new_n10105__), .dout(new_new_n10106__));
  buf1  g7008(.din(new_new_n10106__), .dout(new_new_n10107__));
  buf1  g7009(.din(new_new_n10107__), .dout(new_new_n10108__));
  buf1  g7010(.din(new_new_n10106__), .dout(new_new_n10109__));
  buf1  g7011(.din(new_new_n10105__), .dout(new_new_n10110__));
  buf1  g7012(.din(new_new_n10110__), .dout(new_new_n10111__));
  buf1  g7013(.din(new_new_n10110__), .dout(new_new_n10112__));
  buf1  g7014(.din(new_new_n4517__), .dout(new_new_n10113__));
  buf1  g7015(.din(new_new_n4516__), .dout(new_new_n10114__));
  buf1  g7016(.din(new_new_n3927__), .dout(new_new_n10115__));
  buf1  g7017(.din(new_new_n3926__), .dout(new_new_n10116__));
  buf1  g7018(.din(new_new_n10116__), .dout(new_new_n10117__));
  buf1  g7019(.din(new_new_n10117__), .dout(new_new_n10118__));
  buf1  g7020(.din(new_new_n10116__), .dout(new_new_n10119__));
  buf1  g7021(.din(new_new_n6679__), .dout(new_new_n10120__));
  buf1  g7022(.din(new_new_n6658__), .dout(new_new_n10121__));
  buf1  g7023(.din(new_new_n6678__), .dout(new_new_n10122__));
  buf1  g7024(.din(new_new_n6659__), .dout(new_new_n10123__));
  buf1  g7025(.din(new_new_n4529__), .dout(new_new_n10124__));
  buf1  g7026(.din(new_new_n4528__), .dout(new_new_n10125__));
  buf1  g7027(.din(new_new_n3985__), .dout(new_new_n10126__));
  buf1  g7028(.din(new_new_n3984__), .dout(new_new_n10127__));
  buf1  g7029(.din(new_new_n10127__), .dout(new_new_n10128__));
  buf1  g7030(.din(new_new_n10128__), .dout(new_new_n10129__));
  buf1  g7031(.din(new_new_n10127__), .dout(new_new_n10130__));
  buf1  g7032(.din(new_new_n6704__), .dout(new_new_n10131__));
  buf1  g7033(.din(new_new_n6189__), .dout(new_new_n10132__));
  buf1  g7034(.din(new_new_n6705__), .dout(new_new_n10133__));
  buf1  g7035(.din(new_new_n6190__), .dout(new_new_n10134__));
  buf1  g7036(.din(new_new_n10134__), .dout(new_new_n10135__));
  buf1  g7037(.din(new_new_n4523__), .dout(new_new_n10136__));
  buf1  g7038(.din(new_new_n4522__), .dout(new_new_n10137__));
  buf1  g7039(.din(new_new_n3953__), .dout(new_new_n10138__));
  buf1  g7040(.din(new_new_n3952__), .dout(new_new_n10139__));
  buf1  g7041(.din(new_new_n10139__), .dout(new_new_n10140__));
  buf1  g7042(.din(new_new_n10140__), .dout(new_new_n10141__));
  buf1  g7043(.din(new_new_n10139__), .dout(new_new_n10142__));
  buf1  g7044(.din(new_new_n4519__), .dout(new_new_n10143__));
  buf1  g7045(.din(new_new_n4518__), .dout(new_new_n10144__));
  buf1  g7046(.din(new_new_n3931__), .dout(new_new_n10145__));
  buf1  g7047(.din(new_new_n3930__), .dout(new_new_n10146__));
  buf1  g7048(.din(new_new_n10146__), .dout(new_new_n10147__));
  buf1  g7049(.din(new_new_n10147__), .dout(new_new_n10148__));
  buf1  g7050(.din(new_new_n10146__), .dout(new_new_n10149__));
  buf1  g7051(.din(new_new_n6754__), .dout(new_new_n10150__));
  buf1  g7052(.din(new_new_n6733__), .dout(new_new_n10151__));
  buf1  g7053(.din(new_new_n6753__), .dout(new_new_n10152__));
  buf1  g7054(.din(new_new_n6734__), .dout(new_new_n10153__));
  buf1  g7055(.din(new_new_n4015__), .dout(new_new_n10154__));
  buf1  g7056(.din(new_new_n4014__), .dout(new_new_n10155__));
  buf1  g7057(.din(new_new_n10155__), .dout(new_new_n10156__));
  buf1  g7058(.din(new_new_n10156__), .dout(new_new_n10157__));
  buf1  g7059(.din(new_new_n10155__), .dout(new_new_n10158__));
  buf1  g7060(.din(new_new_n4243__), .dout(new_new_n10159__));
  buf1  g7061(.din(new_new_n4242__), .dout(new_new_n10160__));
  buf1  g7062(.din(new_new_n10160__), .dout(new_new_n10161__));
  buf1  g7063(.din(new_new_n10161__), .dout(new_new_n10162__));
  buf1  g7064(.din(new_new_n10160__), .dout(new_new_n10163__));
  buf1  g7065(.din(new_new_n6771__), .dout(new_new_n10164__));
  buf1  g7066(.din(new_new_n6765__), .dout(new_new_n10165__));
  buf1  g7067(.din(new_new_n6772__), .dout(new_new_n10166__));
  buf1  g7068(.din(new_new_n6766__), .dout(new_new_n10167__));
  buf1  g7069(.din(new_new_n4511__), .dout(new_new_n10168__));
  buf1  g7070(.din(new_new_n4510__), .dout(new_new_n10169__));
  buf1  g7071(.din(new_new_n4509__), .dout(new_new_n10170__));
  buf1  g7072(.din(new_new_n4508__), .dout(new_new_n10171__));
  buf1  g7073(.din(new_new_n6841__), .dout(new_new_n10172__));
  buf1  g7074(.din(new_new_n6820__), .dout(new_new_n10173__));
  buf1  g7075(.din(new_new_n6840__), .dout(new_new_n10174__));
  buf1  g7076(.din(new_new_n6821__), .dout(new_new_n10175__));
  buf1  g7077(.din(new_new_n6871__), .dout(new_new_n10176__));
  buf1  g7078(.din(new_new_n6858__), .dout(new_new_n10177__));
  buf1  g7079(.din(new_new_n6870__), .dout(new_new_n10178__));
  buf1  g7080(.din(new_new_n6859__), .dout(new_new_n10179__));
  buf1  g7081(.din(new_new_n6847__), .dout(new_new_n10180__));
  buf1  g7082(.din(new_new_n6800__), .dout(new_new_n10181__));
  buf1  g7083(.din(new_new_n6876__), .dout(new_new_n10182__));
  buf1  g7084(.din(new_new_n6801__), .dout(new_new_n10183__));
  buf1  g7085(.din(new_new_n6877__), .dout(new_new_n10184__));
  buf1  g7086(.din(new_new_n6846__), .dout(new_new_n10185__));
  buf1  g7087(.din(new_new_n4515__), .dout(new_new_n10186__));
  buf1  g7088(.din(new_new_n4514__), .dout(new_new_n10187__));
  buf1  g7089(.din(new_new_n4513__), .dout(new_new_n10188__));
  buf1  g7090(.din(new_new_n4512__), .dout(new_new_n10189__));
  buf1  g7091(.din(new_new_n6928__), .dout(new_new_n10190__));
  buf1  g7092(.din(new_new_n6907__), .dout(new_new_n10191__));
  buf1  g7093(.din(new_new_n6927__), .dout(new_new_n10192__));
  buf1  g7094(.din(new_new_n6908__), .dout(new_new_n10193__));
  buf1  g7095(.din(new_new_n6952__), .dout(new_new_n10194__));
  buf1  g7096(.din(new_new_n6939__), .dout(new_new_n10195__));
  buf1  g7097(.din(new_new_n6951__), .dout(new_new_n10196__));
  buf1  g7098(.din(new_new_n6940__), .dout(new_new_n10197__));
  buf1  g7099(.din(new_new_n6933__), .dout(new_new_n10198__));
  buf1  g7100(.din(new_new_n6272__), .dout(new_new_n10199__));
  buf1  g7101(.din(new_new_n6958__), .dout(new_new_n10200__));
  buf1  g7102(.din(new_new_n6271__), .dout(new_new_n10201__));
  buf1  g7103(.din(new_new_n10201__), .dout(new_new_n10202__));
  buf1  g7104(.din(new_new_n6957__), .dout(new_new_n10203__));
  buf1  g7105(.din(new_new_n6934__), .dout(new_new_n10204__));
  buf1  g7106(.din(new_new_n6553__), .dout(new_new_n10205__));
  buf1  g7107(.din(new_new_n10205__), .dout(new_new_n10206__));
  buf1  g7108(.din(new_new_n3558__), .dout(new_new_n10207__));
  buf1  g7109(.din(new_new_n10207__), .dout(new_new_n10208__));
  buf1  g7110(.din(new_new_n6547__), .dout(new_new_n10209__));
  buf1  g7111(.din(new_new_n10209__), .dout(new_new_n10210__));
  buf1  g7112(.din(new_new_n3586__), .dout(new_new_n10211__));
  buf1  g7113(.din(new_new_n10211__), .dout(new_new_n10212__));
  buf1  g7114(.din(new_new_n4540__), .dout(new_new_n10213__));
  buf1  g7115(.din(new_new_n6980__), .dout(new_new_n10214__));
  buf1  g7116(.din(new_new_n6979__), .dout(new_new_n10215__));
  buf1  g7117(.din(new_new_n6981__), .dout(new_new_n10216__));
  buf1  g7118(.din(new_new_n6978__), .dout(new_new_n10217__));
  buf1  g7119(.din(new_new_n6986__), .dout(new_new_n10218__));
  buf1  g7120(.din(new_new_n4157__), .dout(new_new_n10219__));
  buf1  g7121(.din(new_new_n10219__), .dout(new_new_n10220__));
  buf1  g7122(.din(new_new_n10219__), .dout(new_new_n10221__));
  buf1  g7123(.din(new_new_n6987__), .dout(new_new_n10222__));
  buf1  g7124(.din(new_new_n4156__), .dout(new_new_n10223__));
  buf1  g7125(.din(new_new_n10223__), .dout(new_new_n10224__));
  buf1  g7126(.din(new_new_n10224__), .dout(new_new_n10225__));
  buf1  g7127(.din(new_new_n10223__), .dout(new_new_n10226__));
  buf1  g7128(.din(new_new_n4140__), .dout(new_new_n10227__));
  buf1  g7129(.din(new_new_n10227__), .dout(new_new_n10228__));
  buf1  g7130(.din(new_new_n4141__), .dout(new_new_n10229__));
  buf1  g7131(.din(new_new_n4538__), .dout(new_new_n10230__));
  buf1  g7132(.din(new_new_n7005__), .dout(new_new_n10231__));
  buf1  g7133(.din(new_new_n7004__), .dout(new_new_n10232__));
  buf1  g7134(.din(new_new_n7006__), .dout(new_new_n10233__));
  buf1  g7135(.din(new_new_n7003__), .dout(new_new_n10234__));
  buf1  g7136(.din(new_new_n7011__), .dout(new_new_n10235__));
  buf1  g7137(.din(new_new_n4246__), .dout(new_new_n10236__));
  buf1  g7138(.din(new_new_n10236__), .dout(new_new_n10237__));
  buf1  g7139(.din(new_new_n10237__), .dout(new_new_n10238__));
  buf1  g7140(.din(new_new_n10236__), .dout(new_new_n10239__));
  buf1  g7141(.din(new_new_n7012__), .dout(new_new_n10240__));
  buf1  g7142(.din(new_new_n4247__), .dout(new_new_n10241__));
  buf1  g7143(.din(new_new_n10241__), .dout(new_new_n10242__));
  buf1  g7144(.din(new_new_n10241__), .dout(new_new_n10243__));
  buf1  g7145(.din(new_new_n4144__), .dout(new_new_n10244__));
  buf1  g7146(.din(new_new_n10244__), .dout(new_new_n10245__));
  buf1  g7147(.din(new_new_n4145__), .dout(new_new_n10246__));
  buf1  g7148(.din(new_new_n6280__), .dout(new_new_n10247__));
  buf1  g7149(.din(new_new_n10247__), .dout(new_new_n10248__));
  buf1  g7150(.din(new_new_n10247__), .dout(new_new_n10249__));
  buf1  g7151(.din(new_new_n4542__), .dout(new_new_n10250__));
  buf1  g7152(.din(new_new_n6279__), .dout(new_new_n10251__));
  buf1  g7153(.din(new_new_n10251__), .dout(new_new_n10252__));
  buf1  g7154(.din(new_new_n4488__), .dout(new_new_n10253__));
  buf1  g7155(.din(new_new_n10253__), .dout(new_new_n10254__));
  buf1  g7156(.din(new_new_n10254__), .dout(new_new_n10255__));
  buf1  g7157(.din(new_new_n10254__), .dout(new_new_n10256__));
  buf1  g7158(.din(new_new_n10253__), .dout(new_new_n10257__));
  buf1  g7159(.din(new_new_n10257__), .dout(new_new_n10258__));
  buf1  g7160(.din(new_new_n4454__), .dout(new_new_n10259__));
  buf1  g7161(.din(new_new_n10259__), .dout(new_new_n10260__));
  buf1  g7162(.din(new_new_n10259__), .dout(new_new_n10261__));
  buf1  g7163(.din(new_new_n4489__), .dout(new_new_n10262__));
  buf1  g7164(.din(new_new_n4455__), .dout(new_new_n10263__));
  buf1  g7165(.din(new_new_n10263__), .dout(new_new_n10264__));
  buf1  g7166(.din(new_new_n4612__), .dout(new_new_n10265__));
  buf1  g7167(.din(new_new_n10265__), .dout(new_new_n10266__));
  buf1  g7168(.din(new_new_n10265__), .dout(new_new_n10267__));
  buf1  g7169(.din(new_new_n4613__), .dout(new_new_n10268__));
  buf1  g7170(.din(new_new_n10268__), .dout(new_new_n10269__));
  buf1  g7171(.din(new_new_n6281__), .dout(new_new_n10270__));
  buf1  g7172(.din(new_new_n7034__), .dout(new_new_n10271__));
  buf1  g7173(.din(new_new_n10271__), .dout(new_new_n10272__));
  buf1  g7174(.din(new_new_n7035__), .dout(new_new_n10273__));
  buf1  g7175(.din(new_new_n10273__), .dout(new_new_n10274__));
  buf1  g7176(.din(new_new_n4659__), .dout(new_new_n10275__));
  buf1  g7177(.din(new_new_n10275__), .dout(new_new_n10276__));
  buf1  g7178(.din(new_new_n4658__), .dout(new_new_n10277__));
  buf1  g7179(.din(new_new_n10277__), .dout(new_new_n10278__));
  buf1  g7180(.din(new_new_n4240__), .dout(new_new_n10279__));
  buf1  g7181(.din(new_new_n4234__), .dout(new_new_n10280__));
  buf1  g7182(.din(new_new_n7041__), .dout(new_new_n10281__));
  buf1  g7183(.din(new_new_n7039__), .dout(new_new_n10282__));
  buf1  g7184(.din(new_new_n7040__), .dout(new_new_n10283__));
  buf1  g7185(.din(new_new_n7038__), .dout(new_new_n10284__));
  buf1  g7186(.din(new_new_n7046__), .dout(new_new_n10285__));
  buf1  g7187(.din(new_new_n7037__), .dout(new_new_n10286__));
  buf1  g7188(.din(new_new_n7047__), .dout(new_new_n10287__));
  buf1  g7189(.din(new_new_n7036__), .dout(new_new_n10288__));
  buf1  g7190(.din(new_new_n7061__), .dout(new_new_n10289__));
  buf1  g7191(.din(new_new_n7062__), .dout(new_new_n10290__));
  buf1  g7192(.din(new_new_n6273__), .dout(new_new_n10291__));
  buf1  g7193(.din(new_new_n10291__), .dout(new_new_n10292__));
  buf1  g7194(.din(new_new_n10291__), .dout(new_new_n10293__));
  buf1  g7195(.din(new_new_n4544__), .dout(new_new_n10294__));
  buf1  g7196(.din(new_new_n6274__), .dout(new_new_n10295__));
  buf1  g7197(.din(new_new_n10295__), .dout(new_new_n10296__));
  buf1  g7198(.din(new_new_n10296__), .dout(new_new_n10297__));
  buf1  g7199(.din(new_new_n10296__), .dout(new_new_n10298__));
  buf1  g7200(.din(new_new_n10295__), .dout(new_new_n10299__));
  buf1  g7201(.din(new_new_n10299__), .dout(new_new_n10300__));
  buf1  g7202(.din(new_new_n4490__), .dout(new_new_n10301__));
  buf1  g7203(.din(new_new_n10301__), .dout(new_new_n10302__));
  buf1  g7204(.din(new_new_n10302__), .dout(new_new_n10303__));
  buf1  g7205(.din(new_new_n10302__), .dout(new_new_n10304__));
  buf1  g7206(.din(new_new_n10301__), .dout(new_new_n10305__));
  buf1  g7207(.din(new_new_n10305__), .dout(new_new_n10306__));
  buf1  g7208(.din(new_new_n4456__), .dout(new_new_n10307__));
  buf1  g7209(.din(new_new_n10307__), .dout(new_new_n10308__));
  buf1  g7210(.din(new_new_n10307__), .dout(new_new_n10309__));
  buf1  g7211(.din(new_new_n4491__), .dout(new_new_n10310__));
  buf1  g7212(.din(new_new_n4457__), .dout(new_new_n10311__));
  buf1  g7213(.din(new_new_n10311__), .dout(new_new_n10312__));
  buf1  g7214(.din(new_new_n4614__), .dout(new_new_n10313__));
  buf1  g7215(.din(new_new_n10313__), .dout(new_new_n10314__));
  buf1  g7216(.din(new_new_n10313__), .dout(new_new_n10315__));
  buf1  g7217(.din(new_new_n4615__), .dout(new_new_n10316__));
  buf1  g7218(.din(new_new_n10316__), .dout(new_new_n10317__));
  buf1  g7219(.din(new_new_n7084__), .dout(new_new_n10318__));
  buf1  g7220(.din(new_new_n10318__), .dout(new_new_n10319__));
  buf1  g7221(.din(new_new_n7085__), .dout(new_new_n10320__));
  buf1  g7222(.din(new_new_n10320__), .dout(new_new_n10321__));
  buf1  g7223(.din(new_new_n4661__), .dout(new_new_n10322__));
  buf1  g7224(.din(new_new_n10322__), .dout(new_new_n10323__));
  buf1  g7225(.din(new_new_n4660__), .dout(new_new_n10324__));
  buf1  g7226(.din(new_new_n10324__), .dout(new_new_n10325__));
  buf1  g7227(.din(new_new_n4238__), .dout(new_new_n10326__));
  buf1  g7228(.din(new_new_n4236__), .dout(new_new_n10327__));
  buf1  g7229(.din(new_new_n7091__), .dout(new_new_n10328__));
  buf1  g7230(.din(new_new_n7089__), .dout(new_new_n10329__));
  buf1  g7231(.din(new_new_n7090__), .dout(new_new_n10330__));
  buf1  g7232(.din(new_new_n7088__), .dout(new_new_n10331__));
  buf1  g7233(.din(new_new_n7096__), .dout(new_new_n10332__));
  buf1  g7234(.din(new_new_n7087__), .dout(new_new_n10333__));
  buf1  g7235(.din(new_new_n7097__), .dout(new_new_n10334__));
  buf1  g7236(.din(new_new_n7086__), .dout(new_new_n10335__));
  buf1  g7237(.din(new_new_n7111__), .dout(new_new_n10336__));
  buf1  g7238(.din(new_new_n7112__), .dout(new_new_n10337__));
  buf1  g7239(.din(new_new_n3388__), .dout(new_new_n10338__));
  buf1  g7240(.din(new_new_n6359__), .dout(new_new_n10339__));
  buf1  g7241(.din(new_new_n10339__), .dout(new_new_n10340__));
  buf1  g7242(.din(new_new_n3596__), .dout(new_new_n10341__));
  buf1  g7243(.din(new_new_n10341__), .dout(new_new_n10342__));
  buf1  g7244(.din(new_new_n6360__), .dout(new_new_n10343__));
  buf1  g7245(.din(new_new_n10343__), .dout(new_new_n10344__));
  buf1  g7246(.din(new_new_n3597__), .dout(new_new_n10345__));
  buf1  g7247(.din(new_new_n10345__), .dout(new_new_n10346__));
  buf1  g7248(.din(new_new_n3550__), .dout(new_new_n10347__));
  buf1  g7249(.din(new_new_n10347__), .dout(new_new_n10348__));
  buf1  g7250(.din(new_new_n6366__), .dout(new_new_n10349__));
  buf1  g7251(.din(new_new_n10349__), .dout(new_new_n10350__));
  buf1  g7252(.din(new_new_n3578__), .dout(new_new_n10351__));
  buf1  g7253(.din(new_new_n10351__), .dout(new_new_n10352__));
  buf1  g7254(.din(new_new_n6378__), .dout(new_new_n10353__));
  buf1  g7255(.din(new_new_n10353__), .dout(new_new_n10354__));
  buf1  g7256(.din(new_new_n3582__), .dout(new_new_n10355__));
  buf1  g7257(.din(new_new_n10355__), .dout(new_new_n10356__));
  buf1  g7258(.din(new_new_n6372__), .dout(new_new_n10357__));
  buf1  g7259(.din(new_new_n10357__), .dout(new_new_n10358__));
  buf1  g7260(.din(new_new_n4160__), .dout(new_new_n10359__));
  buf1  g7261(.din(new_new_n10359__), .dout(new_new_n10360__));
  buf1  g7262(.din(new_new_n3431__), .dout(new_new_n10361__));
  buf1  g7263(.din(new_new_n10361__), .dout(new_new_n10362__));
  buf1  g7264(.din(new_new_n3435__), .dout(new_new_n10363__));
  buf1  g7265(.din(new_new_n10363__), .dout(new_new_n10364__));
  buf1  g7266(.din(new_new_n4128__), .dout(new_new_n10365__));
  buf1  g7267(.din(new_new_n10365__), .dout(new_new_n10366__));
  buf1  g7268(.din(new_new_n10365__), .dout(new_new_n10367__));
  buf1  g7269(.din(new_new_n6535__), .dout(new_new_n10368__));
  buf1  g7270(.din(new_new_n10368__), .dout(new_new_n10369__));
  buf1  g7271(.din(new_new_n3571__), .dout(new_new_n10370__));
  buf1  g7272(.din(new_new_n4662__), .dout(new_new_n10371__));
  buf1  g7273(.din(new_new_n4655__), .dout(new_new_n10372__));
  buf1  g7274(.din(new_new_n4663__), .dout(new_new_n10373__));
  buf1  g7275(.din(new_new_n4654__), .dout(new_new_n10374__));
  buf1  g7276(.din(new_new_n7161__), .dout(new_new_n10375__));
  buf1  g7277(.din(new_new_n7162__), .dout(new_new_n10376__));
  buf1  g7278(.din(new_new_n7171__), .dout(new_new_n10377__));
  buf1  g7279(.din(new_new_n6538__), .dout(new_new_n10378__));
  buf1  g7280(.din(new_new_n10378__), .dout(new_new_n10379__));
  buf1  g7281(.din(new_new_n10379__), .dout(new_new_n10380__));
  buf1  g7282(.din(new_new_n10378__), .dout(new_new_n10381__));
  buf1  g7283(.din(new_new_n4665__), .dout(new_new_n10382__));
  buf1  g7284(.din(new_new_n4657__), .dout(new_new_n10383__));
  buf1  g7285(.din(new_new_n4664__), .dout(new_new_n10384__));
  buf1  g7286(.din(new_new_n4656__), .dout(new_new_n10385__));
  buf1  g7287(.din(new_new_n7177__), .dout(new_new_n10386__));
  buf1  g7288(.din(new_new_n7178__), .dout(new_new_n10387__));
  buf1  g7289(.din(new_new_n7187__), .dout(new_new_n10388__));
  buf1  g7290(.din(new_new_n6541__), .dout(new_new_n10389__));
  buf1  g7291(.din(new_new_n10389__), .dout(new_new_n10390__));
  buf1  g7292(.din(new_new_n10390__), .dout(new_new_n10391__));
  buf1  g7293(.din(new_new_n10389__), .dout(new_new_n10392__));
  buf1  g7294(.din(new_new_n3466__), .dout(new_new_n10393__));
  buf1  g7295(.din(new_new_n3472__), .dout(new_new_n10394__));
  buf1  g7296(.din(new_new_n6328__), .dout(new_new_n10395__));
  buf1  g7297(.din(new_new_n10395__), .dout(new_new_n10396__));
  buf1  g7298(.din(new_new_n10395__), .dout(new_new_n10397__));
  buf1  g7299(.din(new_new_n6305__), .dout(new_new_n10398__));
  buf1  g7300(.din(new_new_n10398__), .dout(new_new_n10399__));
  buf1  g7301(.din(new_new_n6327__), .dout(new_new_n10400__));
  buf1  g7302(.din(new_new_n10400__), .dout(new_new_n10401__));
  buf1  g7303(.din(new_new_n6306__), .dout(new_new_n10402__));
  buf1  g7304(.din(new_new_n7202__), .dout(new_new_n10403__));
  buf1  g7305(.din(new_new_n7133__), .dout(new_new_n10404__));
  buf1  g7306(.din(new_new_n10404__), .dout(new_new_n10405__));
  buf1  g7307(.din(new_new_n10405__), .dout(new_new_n10406__));
  buf1  g7308(.din(new_new_n10404__), .dout(new_new_n10407__));
  buf1  g7309(.din(new_new_n6340__), .dout(new_new_n10408__));
  buf1  g7310(.din(new_new_n10408__), .dout(new_new_n10409__));
  buf1  g7311(.din(new_new_n6307__), .dout(new_new_n10410__));
  buf1  g7312(.din(new_new_n10410__), .dout(new_new_n10411__));
  buf1  g7313(.din(new_new_n6339__), .dout(new_new_n10412__));
  buf1  g7314(.din(new_new_n10412__), .dout(new_new_n10413__));
  buf1  g7315(.din(new_new_n6308__), .dout(new_new_n10414__));
  buf1  g7316(.din(new_new_n7206__), .dout(new_new_n10415__));
  buf1  g7317(.din(new_new_n7129__), .dout(new_new_n10416__));
  buf1  g7318(.din(new_new_n10416__), .dout(new_new_n10417__));
  buf1  g7319(.din(new_new_n10416__), .dout(new_new_n10418__));
  buf1  g7320(.din(new_new_n6334__), .dout(new_new_n10419__));
  buf1  g7321(.din(new_new_n10419__), .dout(new_new_n10420__));
  buf1  g7322(.din(new_new_n10420__), .dout(new_new_n10421__));
  buf1  g7323(.din(new_new_n10420__), .dout(new_new_n10422__));
  buf1  g7324(.din(new_new_n10419__), .dout(new_new_n10423__));
  buf1  g7325(.din(new_new_n6333__), .dout(new_new_n10424__));
  buf1  g7326(.din(new_new_n10424__), .dout(new_new_n10425__));
  buf1  g7327(.din(new_new_n6321__), .dout(new_new_n10426__));
  buf1  g7328(.din(new_new_n10426__), .dout(new_new_n10427__));
  buf1  g7329(.din(new_new_n10427__), .dout(new_new_n10428__));
  buf1  g7330(.din(new_new_n10426__), .dout(new_new_n10429__));
  buf1  g7331(.din(new_new_n6322__), .dout(new_new_n10430__));
  buf1  g7332(.din(new_new_n10430__), .dout(new_new_n10431__));
  buf1  g7333(.din(new_new_n10430__), .dout(new_new_n10432__));
  buf1  g7334(.din(new_new_n7210__), .dout(new_new_n10433__));
  buf1  g7335(.din(new_new_n3476__), .dout(new_new_n10434__));
  buf1  g7336(.din(new_new_n6356__), .dout(new_new_n10435__));
  buf1  g7337(.din(new_new_n10435__), .dout(new_new_n10436__));
  buf1  g7338(.din(new_new_n7214__), .dout(new_new_n10437__));
  buf1  g7339(.din(new_new_n6346__), .dout(new_new_n10438__));
  buf1  g7340(.din(new_new_n10438__), .dout(new_new_n10439__));
  buf1  g7341(.din(new_new_n6345__), .dout(new_new_n10440__));
  buf1  g7342(.din(new_new_n10440__), .dout(new_new_n10441__));
  buf1  g7343(.din(new_new_n10440__), .dout(new_new_n10442__));
  buf1  g7344(.din(new_new_n6299__), .dout(new_new_n10443__));
  buf1  g7345(.din(new_new_n10443__), .dout(new_new_n10444__));
  buf1  g7346(.din(new_new_n10443__), .dout(new_new_n10445__));
  buf1  g7347(.din(new_new_n6300__), .dout(new_new_n10446__));
  buf1  g7348(.din(new_new_n10446__), .dout(new_new_n10447__));
  buf1  g7349(.din(new_new_n10447__), .dout(new_new_n10448__));
  buf1  g7350(.din(new_new_n10447__), .dout(new_new_n10449__));
  buf1  g7351(.din(new_new_n10446__), .dout(new_new_n10450__));
  buf1  g7352(.din(new_new_n10450__), .dout(new_new_n10451__));
  buf1  g7353(.din(new_new_n10450__), .dout(new_new_n10452__));
  buf1  g7354(.din(new_new_n7221__), .dout(new_new_n10453__));
  buf1  g7355(.din(new_new_n7223__), .dout(new_new_n10454__));
  buf1  g7356(.din(new_new_n6347__), .dout(new_new_n10455__));
  buf1  g7357(.din(new_new_n10455__), .dout(new_new_n10456__));
  buf1  g7358(.din(new_new_n6350__), .dout(new_new_n10457__));
  buf1  g7359(.din(new_new_n6349__), .dout(new_new_n10458__));
  buf1  g7360(.din(new_new_n7231__), .dout(new_new_n10459__));
  buf1  g7361(.din(new_new_n10459__), .dout(new_new_n10460__));
  buf1  g7362(.din(new_new_n7234__), .dout(new_new_n10461__));
  buf1  g7363(.din(new_new_n7237__), .dout(new_new_n10462__));
  buf1  g7364(.din(new_new_n7238__), .dout(new_new_n10463__));
  buf1  g7365(.din(new_new_n7233__), .dout(new_new_n10464__));
  buf1  g7366(.din(new_new_n7243__), .dout(new_new_n10465__));
  buf1  g7367(.din(new_new_n7250__), .dout(new_new_n10466__));
  buf1  g7368(.din(new_new_n10466__), .dout(new_new_n10467__));
  buf1  g7369(.din(new_new_n7251__), .dout(new_new_n10468__));
  buf1  g7370(.din(new_new_n10468__), .dout(new_new_n10469__));
  buf1  g7371(.din(new_new_n7258__), .dout(new_new_n10470__));
  buf1  g7372(.din(new_new_n7245__), .dout(new_new_n10471__));
  buf1  g7373(.din(new_new_n7197__), .dout(new_new_n10472__));
  buf1  g7374(.din(new_new_n7136__), .dout(new_new_n10473__));
  buf1  g7375(.din(new_new_n10473__), .dout(new_new_n10474__));
  buf1  g7376(.din(new_new_n7200__), .dout(new_new_n10475__));
  buf1  g7377(.din(new_new_n7139__), .dout(new_new_n10476__));
  buf1  g7378(.din(new_new_n10476__), .dout(new_new_n10477__));
  buf1  g7379(.din(new_new_n7226__), .dout(new_new_n10478__));
  buf1  g7380(.din(new_new_n7153__), .dout(new_new_n10479__));
  buf1  g7381(.din(new_new_n7204__), .dout(new_new_n10480__));
  buf1  g7382(.din(new_new_n7212__), .dout(new_new_n10481__));
  buf1  g7383(.din(new_new_n7227__), .dout(new_new_n10482__));
  buf1  g7384(.din(new_new_n7152__), .dout(new_new_n10483__));
  buf1  g7385(.din(new_new_n7207__), .dout(new_new_n10484__));
  buf1  g7386(.din(new_new_n7222__), .dout(new_new_n10485__));
  buf1  g7387(.din(new_new_n6970__), .dout(new_new_n10486__));
  buf1  g7388(.din(new_new_n7154__), .dout(new_new_n10487__));
  buf1  g7389(.din(new_new_n6971__), .dout(new_new_n10488__));
  buf1  g7390(.din(new_new_n7155__), .dout(new_new_n10489__));
  buf1  g7391(.din(new_new_n7232__), .dout(new_new_n10490__));
  buf1  g7392(.din(new_new_n2578__), .dout(new_new_n10491__));
  buf1  g7393(.din(new_new_n2572__), .dout(new_new_n10492__));
  buf1  g7394(.din(new_new_n10492__), .dout(new_new_n10493__));
  buf1  g7395(.din(new_new_n10493__), .dout(new_new_n10494__));
  buf1  g7396(.din(new_new_n10492__), .dout(new_new_n10495__));
  buf1  g7397(.din(new_new_n2580__), .dout(new_new_n10496__));
  buf1  g7398(.din(new_new_n2573__), .dout(new_new_n10497__));
  buf1  g7399(.din(new_new_n2582__), .dout(new_new_n10498__));
  buf1  g7400(.din(new_new_n2584__), .dout(new_new_n10499__));
  buf1  g7401(.din(new_new_n2574__), .dout(new_new_n10500__));
  buf1  g7402(.din(new_new_n10500__), .dout(new_new_n10501__));
  buf1  g7403(.din(new_new_n10501__), .dout(new_new_n10502__));
  buf1  g7404(.din(new_new_n10501__), .dout(new_new_n10503__));
  buf1  g7405(.din(new_new_n10500__), .dout(new_new_n10504__));
  buf1  g7406(.din(new_new_n2536__), .dout(new_new_n10505__));
  buf1  g7407(.din(new_new_n2575__), .dout(new_new_n10506__));
  buf1  g7408(.din(new_new_n10506__), .dout(new_new_n10507__));
  buf1  g7409(.din(new_new_n2540__), .dout(new_new_n10508__));
  buf1  g7410(.din(new_new_n2544__), .dout(new_new_n10509__));
  buf1  g7411(.din(new_new_n3611__), .dout(new_new_n10510__));
  buf1  g7412(.din(new_new_n10510__), .dout(new_new_n10511__));
  buf1  g7413(.din(new_new_n3618__), .dout(new_new_n10512__));
  buf1  g7414(.din(new_new_n2691__), .dout(new_new_n10513__));
  buf1  g7415(.din(new_new_n10513__), .dout(new_new_n10514__));
  buf1  g7416(.din(new_new_n10513__), .dout(new_new_n10515__));
  buf1  g7417(.din(new_new_n3475__), .dout(new_new_n10516__));
  buf1  g7418(.din(new_new_n4726__), .dout(new_new_n10517__));
  buf1  g7419(.din(new_new_n4038__), .dout(new_new_n10518__));
  buf1  g7420(.din(new_new_n4248__), .dout(new_new_n10519__));
  buf1  g7421(.din(new_new_n10519__), .dout(new_new_n10520__));
  buf1  g7422(.din(new_new_n4044__), .dout(new_new_n10521__));
  buf1  g7423(.din(new_new_n10521__), .dout(new_new_n10522__));
  buf1  g7424(.din(new_new_n10521__), .dout(new_new_n10523__));
  buf1  g7425(.din(new_new_n4046__), .dout(new_new_n10524__));
  buf1  g7426(.din(new_new_n10524__), .dout(new_new_n10525__));
  buf1  g7427(.din(new_new_n10524__), .dout(new_new_n10526__));
  buf1  g7428(.din(new_new_n4048__), .dout(new_new_n10527__));
  buf1  g7429(.din(new_new_n10527__), .dout(new_new_n10528__));
  buf1  g7430(.din(new_new_n10527__), .dout(new_new_n10529__));
  buf1  g7431(.din(new_new_n4052__), .dout(new_new_n10530__));
  buf1  g7432(.din(new_new_n10530__), .dout(new_new_n10531__));
  buf1  g7433(.din(new_new_n10530__), .dout(new_new_n10532__));
  buf1  g7434(.din(new_new_n4126__), .dout(new_new_n10533__));
  buf1  g7435(.din(new_new_n4130__), .dout(new_new_n10534__));
  buf1  g7436(.din(new_new_n4152__), .dout(new_new_n10535__));
  buf1  g7437(.din(new_new_n4154__), .dout(new_new_n10536__));
  buf1  g7438(.din(new_new_n4250__), .dout(new_new_n10537__));
  buf1  g7439(.din(new_new_n6422__), .dout(new_new_n10538__));
  buf1  g7440(.din(new_new_n6451__), .dout(new_new_n10539__));
  buf1  g7441(.din(new_new_n6494__), .dout(new_new_n10540__));
  buf1  g7442(.din(new_new_n6523__), .dout(new_new_n10541__));
  buf1  g7443(.din(new_new_n6529__), .dout(new_new_n10542__));
  buf1  g7444(.din(new_new_n3430__), .dout(new_new_n10543__));
  buf1  g7445(.din(new_new_n3434__), .dout(new_new_n10544__));
  buf1  g7446(.din(new_new_n6996__), .dout(new_new_n10545__));
  buf1  g7447(.din(new_new_n7021__), .dout(new_new_n10546__));
  buf1  g7448(.din(new_new_n7056__), .dout(new_new_n10547__));
  buf1  g7449(.din(new_new_n7071__), .dout(new_new_n10548__));
  buf1  g7450(.din(new_new_n7106__), .dout(new_new_n10549__));
  buf1  g7451(.din(new_new_n7121__), .dout(new_new_n10550__));
  buf1  g7452(.din(new_new_n3574__), .dout(new_new_n10551__));
  buf1  g7453(.din(new_new_n10551__), .dout(new_new_n10552__));
  buf1  g7454(.din(new_new_n7124__), .dout(new_new_n10553__));
  buf1  g7455(.din(new_new_n10553__), .dout(new_new_n10554__));
  buf1  g7456(.din(new_new_n3418__), .dout(new_new_n10555__));
  buf1  g7457(.din(new_new_n3438__), .dout(new_new_n10556__));
  buf1  g7458(.din(new_new_n7294__), .dout(new_new_n10557__));
  buf1  g7459(.din(new_new_n7297__), .dout(new_new_n10558__));
  buf1  g7460(.din(new_new_n7300__), .dout(new_new_n10559__));
  buf1  g7461(.din(new_new_n7303__), .dout(new_new_n10560__));
  buf1  g7462(.din(new_new_n2602__), .dout(new_new_n10561__));
  buf1  g7463(.din(new_new_n2604__), .dout(new_new_n10562__));
  buf1  g7464(.din(new_new_n2624__), .dout(new_new_n10563__));
  buf1  g7465(.din(new_new_n2626__), .dout(new_new_n10564__));
  always @ (posedge clock) begin
    n2610_lo <= n16425;
    n2613_lo <= n16428;
    n2616_lo <= n16431;
    n2619_lo <= n16434;
    n2622_lo <= n16437;
    n2625_lo <= n16440;
    n2628_lo <= n16443;
    n2631_lo <= n16446;
    n2634_lo <= n16449;
    n2637_lo <= n16452;
    n2640_lo <= n16455;
    n2643_lo <= n16458;
    n2646_lo <= n16461;
    n2649_lo <= n16464;
    n2652_lo <= n16467;
    n2655_lo <= n16470;
    n2658_lo <= n16473;
    n2661_lo <= n16476;
    n2664_lo <= n16479;
    n2667_lo <= n16482;
    n2670_lo <= n16485;
    n2673_lo <= n16488;
    n2676_lo <= n16491;
    n2679_lo <= n16494;
    n2682_lo <= n16497;
    n2685_lo <= n16500;
    n2688_lo <= n16503;
    n2691_lo <= n16506;
    n2694_lo <= n16509;
    n2697_lo <= n16512;
    n2700_lo <= n16515;
    n2703_lo <= n16518;
    n2706_lo <= n16521;
    n2709_lo <= n16524;
    n2712_lo <= n16527;
    n2715_lo <= n16530;
    n2718_lo <= n16533;
    n2721_lo <= n16536;
    n2724_lo <= n16539;
    n2727_lo <= n16542;
    n2730_lo <= n16545;
    n2733_lo <= n16548;
    n2736_lo <= n16551;
    n2739_lo <= n16554;
    n2742_lo <= n16557;
    n2745_lo <= n16560;
    n2748_lo <= n16563;
    n2751_lo <= n16566;
    n2754_lo <= n16569;
    n2757_lo <= n16572;
    n2760_lo <= n16575;
    n2763_lo <= n16578;
    n2766_lo <= n16581;
    n2769_lo <= n16584;
    n2772_lo <= n16587;
    n2775_lo <= n16590;
    n2778_lo <= n16593;
    n2781_lo <= n16596;
    n2784_lo <= n16599;
    n2787_lo <= n16602;
    n2790_lo <= n16605;
    n2793_lo <= n16608;
    n2796_lo <= n16611;
    n2799_lo <= n16614;
    n2802_lo <= n16617;
    n2805_lo <= n16620;
    n2808_lo <= n16623;
    n2811_lo <= n16626;
    n2814_lo <= n16629;
    n2817_lo <= n16632;
    n2820_lo <= n16635;
    n2823_lo <= n16638;
    n2826_lo <= n16641;
    n2829_lo <= n16644;
    n2832_lo <= n16647;
    n2835_lo <= n16650;
    n2838_lo <= n16653;
    n2841_lo <= n16656;
    n2844_lo <= n16659;
    n2847_lo <= n16662;
    n2850_lo <= n16665;
    n2853_lo <= n16668;
    n2856_lo <= n16671;
    n2859_lo <= n16674;
    n2862_lo <= n16677;
    n2865_lo <= n16680;
    n2868_lo <= n16683;
    n2871_lo <= n16686;
    n2874_lo <= n16689;
    n2877_lo <= n16692;
    n2880_lo <= n16695;
    n2883_lo <= n16698;
    n2886_lo <= n16701;
    n2889_lo <= n16704;
    n2892_lo <= n16707;
    n2895_lo <= n16710;
    n2898_lo <= n16713;
    n2901_lo <= n16716;
    n2904_lo <= n16719;
    n2907_lo <= n16722;
    n2910_lo <= n16725;
    n2913_lo <= n16728;
    n2916_lo <= n16731;
    n2919_lo <= n16734;
    n2922_lo <= n16737;
    n2925_lo <= n16740;
    n2928_lo <= n16743;
    n2931_lo <= n16746;
    n2934_lo <= n16749;
    n2937_lo <= n16752;
    n2940_lo <= n16755;
    n2943_lo <= n16758;
    n2946_lo <= n16761;
    n2949_lo <= n16764;
    n2952_lo <= n16767;
    n2955_lo <= n16770;
    n2958_lo <= n16773;
    n2961_lo <= n16776;
    n2964_lo <= n16779;
    n2967_lo <= n16782;
    n2970_lo <= n16785;
    n2973_lo <= n16788;
    n2976_lo <= n16791;
    n2979_lo <= n16794;
    n2982_lo <= n16797;
    n2985_lo <= n16800;
    n2988_lo <= n16803;
    n2991_lo <= n16806;
    n2994_lo <= n16809;
    n2997_lo <= n16812;
    n3000_lo <= n16815;
    n3003_lo <= n16818;
    n3006_lo <= n16821;
    n3009_lo <= n16824;
    n3012_lo <= n16827;
    n3015_lo <= n16830;
    n3018_lo <= n16833;
    n3021_lo <= n16836;
    n3024_lo <= n16839;
    n3027_lo <= n16842;
    n3030_lo <= n16845;
    n3033_lo <= n16848;
    n3036_lo <= n16851;
    n3039_lo <= n16854;
    n3042_lo <= n16857;
    n3045_lo <= n16860;
    n3048_lo <= n16863;
    n3051_lo <= n16866;
    n3054_lo <= n16869;
    n3057_lo <= n16872;
    n3060_lo <= n16875;
    n3063_lo <= n16878;
    n3066_lo <= n16881;
    n3069_lo <= n16884;
    n3072_lo <= n16887;
    n3075_lo <= n16890;
    n3078_lo <= n16893;
    n3081_lo <= n16896;
    n3084_lo <= n16899;
    n3087_lo <= n16902;
    n3090_lo <= n16905;
    n3093_lo <= n16908;
    n3096_lo <= n16911;
    n3099_lo <= n16914;
    n3102_lo <= n16917;
    n3105_lo <= n16920;
    n3108_lo <= n16923;
    n3111_lo <= n16926;
    n3114_lo <= n16929;
    n3117_lo <= n16932;
    n3120_lo <= n16935;
    n3123_lo <= n16938;
    n3126_lo <= n16941;
    n3129_lo <= n16944;
    n3132_lo <= n16947;
    n3135_lo <= n16950;
    n3138_lo <= n16953;
    n3141_lo <= n16956;
    n3144_lo <= n16959;
    n3147_lo <= n16962;
    n3150_lo <= n16965;
    n3153_lo <= n16968;
    n3156_lo <= n16971;
    n3159_lo <= n16974;
    n3162_lo <= n16977;
    n3165_lo <= n16980;
    n3168_lo <= n16983;
    n3171_lo <= n16986;
    n3174_lo <= n16989;
    n3177_lo <= n16992;
    n3180_lo <= n16995;
    n3183_lo <= n16998;
    n3186_lo <= n17001;
    n3189_lo <= n17004;
    n3192_lo <= n17007;
    n3195_lo <= n17010;
    n3198_lo <= n17013;
    n3201_lo <= n17016;
    n3204_lo <= n17019;
    n3207_lo <= n17022;
    n3210_lo <= n17025;
    n3213_lo <= n17028;
    n3216_lo <= n17031;
    n3219_lo <= n17034;
    n3222_lo <= n17037;
    n3225_lo <= n17040;
    n3228_lo <= n17043;
    n3231_lo <= n17046;
    n3234_lo <= n17049;
    n3237_lo <= n17052;
    n3240_lo <= n17055;
    n3243_lo <= n17058;
    n3246_lo <= n17061;
    n3249_lo <= n17064;
    n3252_lo <= n17067;
    n3255_lo <= n17070;
    n3258_lo <= n17073;
    n3261_lo <= n17076;
    n3264_lo <= n17079;
    n3267_lo <= n17082;
    n3270_lo <= n17085;
    n3273_lo <= n17088;
    n3276_lo <= n17091;
    n3279_lo <= n17094;
    n3282_lo <= n17097;
    n3285_lo <= n17100;
    n3288_lo <= n17103;
    n3291_lo <= n17106;
    n3294_lo <= n17109;
    n3297_lo <= n17112;
    n3300_lo <= n17115;
    n3303_lo <= n17118;
    n3306_lo <= n17121;
    n3309_lo <= n17124;
    n3312_lo <= n17127;
    n3315_lo <= n17130;
    n3318_lo <= n17133;
    n3321_lo <= n17136;
    n3324_lo <= n17139;
    n3327_lo <= n17142;
    n3330_lo <= n17145;
    n3333_lo <= n17148;
    n3336_lo <= n17151;
    n3339_lo <= n17154;
    n3342_lo <= n17157;
    n3345_lo <= n17160;
    n3348_lo <= n17163;
    n3351_lo <= n17166;
    n3354_lo <= n17169;
    n3357_lo <= n17172;
    n3360_lo <= n17175;
    n3363_lo <= n17178;
    n3366_lo <= n17181;
    n3369_lo <= n17184;
    n3372_lo <= n17187;
    n3375_lo <= n17190;
    n3378_lo <= n17193;
    n3381_lo <= n17196;
    n3384_lo <= n17199;
    n3387_lo <= n17202;
    n3390_lo <= n17205;
    n3393_lo <= n17208;
    n3396_lo <= n17211;
    n3399_lo <= n17214;
    n3402_lo <= n17217;
    n3405_lo <= n17220;
    n3408_lo <= n17223;
    n3411_lo <= n17226;
    n3414_lo <= n17229;
    n3417_lo <= n17232;
    n3420_lo <= n17235;
    n3423_lo <= n17238;
    n3426_lo <= n17241;
    n3429_lo <= n17244;
    n3432_lo <= n17247;
    n3435_lo <= n17250;
    n3438_lo <= n17253;
    n3441_lo <= n17256;
    n3444_lo <= n17259;
    n3447_lo <= n17262;
    n3450_lo <= n17265;
    n3453_lo <= n17268;
    n3456_lo <= n17271;
    n3459_lo <= n17274;
    n3462_lo <= n17277;
    n3465_lo <= n17280;
    n3468_lo <= n17283;
    n3471_lo <= n17286;
    n3474_lo <= n17289;
    n3477_lo <= n17292;
    n3480_lo <= n17295;
    n3483_lo <= n17298;
    n3486_lo <= n17301;
    n3489_lo <= n17304;
    n3492_lo <= n17307;
    n3495_lo <= n17310;
    n3498_lo <= n17313;
    n3501_lo <= n17316;
    n3504_lo <= n17319;
    n3507_lo <= n17322;
    n3510_lo <= n17325;
    n3513_lo <= n17328;
    n3516_lo <= n17331;
    n3519_lo <= n17334;
    n3522_lo <= n17337;
    n3525_lo <= n17340;
    n3528_lo <= n17343;
    n3531_lo <= n17346;
    n3534_lo <= n17349;
    n3537_lo <= n17352;
    n3540_lo <= n17355;
    n3543_lo <= n17358;
    n3546_lo <= n17361;
    n3549_lo <= n17364;
    n3552_lo <= n17367;
    n3555_lo <= n17370;
    n3558_lo <= n17373;
    n3561_lo <= n17376;
    n3564_lo <= n17379;
    n3567_lo <= n17382;
    n3570_lo <= n17385;
    n3573_lo <= n17388;
    n3576_lo <= n17391;
    n3579_lo <= n17394;
    n3582_lo <= n17397;
    n3585_lo <= n17400;
    n3588_lo <= n17403;
    n3591_lo <= n17406;
    n3594_lo <= n17409;
    n3597_lo <= n17412;
    n3600_lo <= n17415;
    n3603_lo <= n17418;
    n3606_lo <= n17421;
    n3609_lo <= n17424;
    n3612_lo <= n17427;
    n3615_lo <= n17430;
    n3618_lo <= n17433;
    n3621_lo <= n17436;
    n3624_lo <= n17439;
    n3627_lo <= n17442;
    n3630_lo <= n17445;
    n3633_lo <= n17448;
    n3636_lo <= n17451;
    n3639_lo <= n17454;
    n3642_lo <= n17457;
    n3645_lo <= n17460;
    n3648_lo <= n17463;
    n3651_lo <= n17466;
    n3654_lo <= n17469;
    n3657_lo <= n17472;
    n3666_lo <= n17475;
    n3669_lo <= n17478;
    n3678_lo <= n17481;
    n3687_lo <= n17484;
    n3690_lo <= n17487;
    n3702_lo <= n17490;
    n3711_lo <= n17493;
    n3714_lo <= n17496;
    n3726_lo <= n17499;
    n3735_lo <= n17502;
    n3738_lo <= n17505;
    n3750_lo <= n17508;
    n3753_lo <= n17511;
    n3759_lo <= n17514;
    n3762_lo <= n17517;
    n3765_lo <= n17520;
    n3774_lo <= n17523;
    n3777_lo <= n17526;
    n3786_lo <= n17529;
    n3789_lo <= n17532;
    n3792_lo <= n17535;
    n3795_lo <= n17538;
    n3798_lo <= n17541;
    n3801_lo <= n17544;
    n3810_lo <= n17547;
    n3813_lo <= n17550;
    n3822_lo <= n17553;
    n3825_lo <= n17556;
    n3834_lo <= n17559;
    n3843_lo <= n17562;
    n3846_lo <= n17565;
    n3867_lo <= n17568;
    n3891_lo <= n17571;
    n3915_lo <= n17574;
    n3930_lo <= n17577;
    n3933_lo <= n17580;
    n3936_lo <= n17583;
    n3942_lo <= n17586;
    n3945_lo <= n17589;
    n3948_lo <= n17592;
    n3954_lo <= n17595;
    n3957_lo <= n17598;
    n3963_lo <= n17601;
    n3966_lo <= n17604;
    n3969_lo <= n17607;
    n3975_lo <= n17610;
    n3978_lo <= n17613;
    n3987_lo <= n17616;
    n3990_lo <= n17619;
    n4002_lo <= n17622;
    n4011_lo <= n17625;
    n4014_lo <= n17628;
    n4026_lo <= n17631;
    n4035_lo <= n17634;
    n4038_lo <= n17637;
    n4050_lo <= n17640;
    n4053_lo <= n17643;
    n4059_lo <= n17646;
    n4062_lo <= n17649;
    n4065_lo <= n17652;
    n4098_lo <= n17655;
    n4107_lo <= n17658;
    n4119_lo <= n17661;
    n4131_lo <= n17664;
    n4143_lo <= n17667;
    n4155_lo <= n17670;
    n4167_lo <= n17673;
    n4179_lo <= n17676;
    n4182_lo <= n17679;
    n4185_lo <= n17682;
    n4188_lo <= n17685;
    n4194_lo <= n17688;
    n4197_lo <= n17691;
    n4200_lo <= n17694;
    n4206_lo <= n17697;
    n4209_lo <= n17700;
    n4212_lo <= n17703;
    n4215_lo <= n17706;
    n4227_lo <= n17709;
    n4230_lo <= n17712;
    n4233_lo <= n17715;
    n4236_lo <= n17718;
    n4239_lo <= n17721;
    n4242_lo <= n17724;
    n4251_lo <= n17727;
    n4263_lo <= n17730;
    n4275_lo <= n17733;
    n4278_lo <= n17736;
    n4287_lo <= n17739;
    n4290_lo <= n17742;
    n4293_lo <= n17745;
    n4299_lo <= n17748;
    n4302_lo <= n17751;
    n4305_lo <= n17754;
    n4311_lo <= n17757;
    n4314_lo <= n17760;
    n4323_lo <= n17763;
    n4326_lo <= n17766;
    n4335_lo <= n17769;
    n4338_lo <= n17772;
    n4347_lo <= n17775;
    n4350_lo <= n17778;
    n4359_lo <= n17781;
    n4362_lo <= n17784;
    n4365_lo <= n17787;
    n4371_lo <= n17790;
    n4374_lo <= n17793;
    n4383_lo <= n17796;
    n4395_lo <= n17799;
    n4407_lo <= n17802;
    n4410_lo <= n17805;
    n4413_lo <= n17808;
    n4416_lo <= n17811;
    n4419_lo <= n17814;
    n4422_lo <= n17817;
    n4425_lo <= n17820;
    n4428_lo <= n17823;
    n4431_lo <= n17826;
    n4434_lo <= n17829;
    n4437_lo <= n17832;
    n4440_lo <= n17835;
    n4443_lo <= n17838;
    n4446_lo <= n17841;
    n4449_lo <= n17844;
    n4452_lo <= n17847;
    n4455_lo <= n17850;
    n4458_lo <= n17853;
    n4461_lo <= n17856;
    n4464_lo <= n17859;
    n4467_lo <= n17862;
    n4470_lo <= n17865;
    n4473_lo <= n17868;
    n4476_lo <= n17871;
    n4479_lo <= n17874;
    n4482_lo <= n17877;
    n4485_lo <= n17880;
    n4488_lo <= n17883;
    n4494_lo <= n17886;
    n4497_lo <= n17889;
    n4500_lo <= n17892;
    n4503_lo <= n17895;
    n4506_lo <= n17898;
    n4509_lo <= n17901;
    n4512_lo <= n17904;
    n4515_lo <= n17907;
    n4518_lo <= n17910;
    n4521_lo <= n17913;
    n4524_lo <= n17916;
    n4527_lo <= n17919;
    n4530_lo <= n17922;
    n4533_lo <= n17925;
    n4536_lo <= n17928;
    n4539_lo <= n17931;
    n4542_lo <= n17934;
    n4545_lo <= n17937;
    n4548_lo <= n17940;
    n4554_lo <= n17943;
    n4557_lo <= n17946;
    n4560_lo <= n17949;
    n4563_lo <= n17952;
    n4566_lo <= n17955;
    n4569_lo <= n17958;
    n4572_lo <= n17961;
    n4575_lo <= n17964;
    n4578_lo <= n17967;
    n4581_lo <= n17970;
    n4584_lo <= n17973;
    n4587_lo <= n17976;
    n4590_lo <= n17979;
    n4593_lo <= n17982;
    n4596_lo <= n17985;
    n4599_lo <= n17988;
    n4602_lo <= n17991;
    n4605_lo <= n17994;
    n4608_lo <= n17997;
    n4611_lo <= n18000;
    n4614_lo <= n18003;
    n4617_lo <= n18006;
    n4620_lo <= n18009;
    n4623_lo <= n18012;
    n4626_lo <= n18015;
    n4629_lo <= n18018;
    n4632_lo <= n18021;
    n4635_lo <= n18024;
    n4638_lo <= n18027;
    n4641_lo <= n18030;
    n4644_lo <= n18033;
    n4647_lo <= n18036;
    n4650_lo <= n18039;
    n4653_lo <= n18042;
    n4656_lo <= n18045;
    n4659_lo <= n18048;
    n4662_lo <= n18051;
    n4665_lo <= n18054;
    n4668_lo <= n18057;
    n4671_lo <= n18060;
    n4674_lo <= n18063;
    n4677_lo <= n18066;
    n4680_lo <= n18069;
    n4683_lo <= n18072;
    n4686_lo <= n18075;
    n4689_lo <= n18078;
    n4692_lo <= n18081;
    n4695_lo <= n18084;
    n4698_lo <= n18087;
    n4701_lo <= n18090;
    n4704_lo <= n18093;
    n4707_lo <= n18096;
    n4710_lo <= n18099;
    n4713_lo <= n18102;
    n4716_lo <= n18105;
    n4719_lo <= n18108;
    n4722_lo <= n18111;
    n4725_lo <= n18114;
    n4728_lo <= n18117;
    n4731_lo <= n18120;
    n4734_lo <= n18123;
    n4737_lo <= n18126;
    n4740_lo <= n18129;
    n4743_lo <= n18132;
    n6382_o2 <= n18135;
    n6383_o2 <= n18138;
    n6419_o2 <= n18141;
    n6420_o2 <= n18144;
    n6435_o2 <= n18147;
    n6436_o2 <= n18150;
    n6448_o2 <= n18153;
    n6449_o2 <= n18156;
    n6613_o2 <= n18159;
    n6614_o2 <= n18162;
    n6641_o2 <= n18165;
    n6658_o2 <= n18168;
    n6757_o2 <= n18171;
    n6756_o2 <= n18174;
    n7116_o2 <= n18177;
    n7156_o2 <= n18180;
    n6549_o2 <= n18183;
    n6550_o2 <= n18186;
    n7357_o2 <= n18189;
    n7358_o2 <= n18192;
    n7359_o2 <= n18195;
    n7360_o2 <= n18198;
    n6621_o2 <= n18201;
    n6623_o2 <= n18204;
    n6625_o2 <= n18207;
    n6626_o2 <= n18210;
    n6627_o2 <= n18213;
    n6628_o2 <= n18216;
    n6629_o2 <= n18219;
    n6630_o2 <= n18222;
    n6669_o2 <= n18225;
    n7449_o2 <= n18228;
    n7450_o2 <= n18231;
    n7451_o2 <= n18234;
    n7452_o2 <= n18237;
    n6682_o2 <= n18240;
    n6683_o2 <= n18243;
    n6684_o2 <= n18246;
    n6685_o2 <= n18249;
    n7463_o2 <= n18252;
    n6686_o2 <= n18255;
    n6687_o2 <= n18258;
    n6688_o2 <= n18261;
    n6689_o2 <= n18264;
    n6772_o2 <= n18267;
    n6773_o2 <= n18270;
    n6774_o2 <= n18273;
    n6775_o2 <= n18276;
    G3467_o2 <= n18279;
    G2810_o2 <= n18282;
    n6833_o2 <= n18285;
    n6945_o2 <= n18288;
    n6947_o2 <= n18291;
    n6949_o2 <= n18294;
    n6951_o2 <= n18297;
    n6888_o2 <= n18300;
    n6889_o2 <= n18303;
    n6936_o2 <= n18306;
    n6954_o2 <= n18309;
    n6955_o2 <= n18312;
    n6956_o2 <= n18315;
    n6957_o2 <= n18318;
    n6958_o2 <= n18321;
    n6982_o2 <= n18324;
    n6984_o2 <= n18327;
    n6974_o2 <= n18330;
    n6975_o2 <= n18333;
    n6999_o2 <= n18336;
    n7015_o2 <= n18339;
    n7016_o2 <= n18342;
    n7017_o2 <= n18345;
    n7018_o2 <= n18348;
    n7005_o2 <= n18351;
    n7019_o2 <= n18354;
    n7022_o2 <= n18357;
    n7023_o2 <= n18360;
    n7132_o2 <= n18363;
    n7133_o2 <= n18366;
    n7135_o2 <= n18369;
    n7136_o2 <= n18372;
    n7175_o2 <= n18375;
    n7155_o2 <= n18378;
    G3060_o2 <= n18381;
    n7383_o2 <= n18384;
    G3802_o2 <= n18387;
    G3859_o2 <= n18390;
    n7355_o2 <= n18393;
    n7356_o2 <= n18396;
    G4054_o2 <= n18399;
    G4068_o2 <= n18402;
    n7384_o2 <= n18405;
    n7387_o2 <= n18408;
    n7388_o2 <= n18411;
    n7389_o2 <= n18414;
    n7386_o2 <= n18417;
    n7453_o2 <= n18420;
    n7431_o2 <= n18423;
    n7432_o2 <= n18426;
    n7433_o2 <= n18429;
    n7430_o2 <= n18432;
    n7485_o2 <= n18435;
    n7486_o2 <= n18438;
    G2508_o2 <= n18441;
    G2486_o2 <= n18444;
    n2326_inv <= n18447;
    n2329_inv <= n18450;
    n3756_lo_buf_o2 <= n18453;
    n4056_lo_buf_o2 <= n18456;
    G3474_o2 <= n18459;
    n2341_inv <= n18462;
    n7396_o2 <= n18465;
    n7398_o2 <= n18468;
    n7400_o2 <= n18471;
    n7401_o2 <= n18474;
    n7402_o2 <= n18477;
    n7403_o2 <= n18480;
    n7404_o2 <= n18483;
    n7405_o2 <= n18486;
    G2711_o2 <= n18489;
    n2371_inv <= n18492;
    n7490_o2 <= n18495;
    n7527_o2 <= n18498;
    n7528_o2 <= n18501;
    n7529_o2 <= n18504;
    n7530_o2 <= n18507;
    n7523_o2 <= n18510;
    n7524_o2 <= n18513;
    n7525_o2 <= n18516;
    n7526_o2 <= n18519;
    n4296_lo_buf_o2 <= n18522;
    n4368_lo_buf_o2 <= n18525;
    G2466_o2 <= n18528;
    G2404_o2 <= n18531;
    n7534_o2 <= n18534;
    n7535_o2 <= n18537;
    n7536_o2 <= n18540;
    n7533_o2 <= n18543;
    G1060_o2 <= n18546;
    G963_o2 <= n18549;
    G2448_o2 <= n18552;
    G2685_o2 <= n18555;
    G2679_o2 <= n18558;
    G2774_o2 <= n18561;
    G2780_o2 <= n18564;
    G2759_o2 <= n18567;
    G2737_o2 <= n18570;
    G2850_o2 <= n18573;
    G3393_o2 <= n18576;
    G3404_o2 <= n18579;
    G3559_o2 <= n18582;
    G2744_o2 <= n18585;
    n3708_lo_buf_o2 <= n18588;
    n3840_lo_buf_o2 <= n18591;
    n4008_lo_buf_o2 <= n18594;
    n4104_lo_buf_o2 <= n18597;
    G1821_o2 <= n18600;
    G1734_o2 <= n18603;
    G3517_o2 <= n18606;
    G3533_o2 <= n18609;
    G3629_o2 <= n18612;
    G3645_o2 <= n18615;
    n2497_inv <= n18618;
    G2731_o2 <= n18621;
    G2844_o2 <= n18624;
    n3732_lo_buf_o2 <= n18627;
    n4032_lo_buf_o2 <= n18630;
    G3552_o2 <= n18633;
    G2271_o2 <= n18636;
    n4248_lo_buf_o2 <= n18639;
    n4332_lo_buf_o2 <= n18642;
    n4344_lo_buf_o2 <= n18645;
    n4380_lo_buf_o2 <= n18648;
    G2398_o2 <= n18651;
    G2480_o2 <= n18654;
    G2418_o2 <= n18657;
    G1455_o2 <= n18660;
    G1449_o2 <= n18663;
    G1452_o2 <= n18666;
    G1425_o2 <= n18669;
    G1428_o2 <= n18672;
    G1419_o2 <= n18675;
    G1422_o2 <= n18678;
    n4308_lo_buf_o2 <= n18681;
    G2675_o2 <= n18684;
    G3035_o2 <= n18687;
    G3026_o2 <= n18690;
    G3029_o2 <= n18693;
    G3032_o2 <= n18696;
    G2999_o2 <= n18699;
    G3002_o2 <= n18702;
    G2770_o2 <= n18705;
    G3008_o2 <= n18708;
    G2073_o2 <= n18711;
    G2752_o2 <= n18714;
    G3005_o2 <= n18717;
    G5108_o2 <= n18720;
    G5135_o2 <= n18723;
    G5111_o2 <= n18726;
    G5138_o2 <= n18729;
    G3415_o2 <= n18732;
    G3386_o2 <= n18735;
    G3570_o2 <= n18738;
    G2430_o2 <= n18741;
    G3495_o2 <= n18744;
    G3621_o2 <= n18747;
    n4284_lo_buf_o2 <= n18750;
    n4356_lo_buf_o2 <= n18753;
    G2472_o2 <= n18756;
    G2410_o2 <= n18759;
    n3960_lo_buf_o2 <= n18762;
    n3972_lo_buf_o2 <= n18765;
    n2647_inv <= n18768;
    n2650_inv <= n18771;
    n3684_lo_buf_o2 <= n18774;
    n4080_lo_buf_o2 <= n18777;
    n4092_lo_buf_o2 <= n18780;
    n2662_inv <= n18783;
    n2665_inv <= n18786;
    G1147_o2 <= n18789;
    G2705_o2 <= n18792;
    G2693_o2 <= n18795;
    G2696_o2 <= n18798;
    G2700_o2 <= n18801;
    G2915_o2 <= n18804;
    G2966_o2 <= n18807;
    G2540_o2 <= n18810;
    G2788_o2 <= n18813;
    G2792_o2 <= n18816;
    G2797_o2 <= n18819;
    G2804_o2 <= n18822;
    G1038_o2 <= n18825;
    G1044_o2 <= n18828;
    G1090_o2 <= n18831;
    G1096_o2 <= n18834;
    G1029_o2 <= n18837;
    G3942_o2 <= n18840;
    G3954_o2 <= n18843;
    G4011_o2 <= n18846;
    G4017_o2 <= n18849;
    G1141_o2 <= n18852;
    G1081_o2 <= n18855;
    G2146_o2 <= n18858;
    G2145_o2 <= n18861;
    G2144_o2 <= n18864;
    G2143_o2 <= n18867;
    G2142_o2 <= n18870;
    G2141_o2 <= n18873;
    G2140_o2 <= n18876;
    G2139_o2 <= n18879;
    G3769_o2 <= n18882;
    G3773_o2 <= n18885;
    G3768_o2 <= n18888;
    G4101_o2 <= n18891;
    G3161_o2 <= n18894;
    G4143_o2 <= n18897;
    G3828_o2 <= n18900;
    G3831_o2 <= n18903;
    G3334_o2 <= n18906;
    G3335_o2 <= n18909;
    G3180_o2 <= n18912;
    G3340_o2 <= n18915;
    G3339_o2 <= n18918;
    G3341_o2 <= n18921;
    G3234_o2 <= n18924;
    G3829_o2 <= n18927;
    G3338_o2 <= n18930;
    G3336_o2 <= n18933;
    G3770_o2 <= n18936;
    G3918_o2 <= n18939;
    G3774_o2 <= n18942;
    G3921_o2 <= n18945;
    G3832_o2 <= n18948;
    G3993_o2 <= n18951;
    G2076_o2 <= n18954;
    G2071_o2 <= n18957;
    G2072_o2 <= n18960;
    G2069_o2 <= n18963;
    G2070_o2 <= n18966;
    G2067_o2 <= n18969;
    G2068_o2 <= n18972;
    G4095_o2 <= n18975;
    G3272_o2 <= n18978;
    G3269_o2 <= n18981;
    G3270_o2 <= n18984;
    G3271_o2 <= n18987;
    G3265_o2 <= n18990;
    G3266_o2 <= n18993;
    G4137_o2 <= n18996;
    G3268_o2 <= n18999;
    G2361_o2 <= n19002;
    G3228_o2 <= n19005;
    G3267_o2 <= n19008;
    G2336_o2 <= n19011;
    G3459_o2 <= n19014;
    G3428_o2 <= n19017;
    G3438_o2 <= n19020;
    G3449_o2 <= n19023;
    G3421_o2 <= n19026;
    G3576_o2 <= n19029;
    G3303_o2 <= n19032;
    G3583_o2 <= n19035;
    G3594_o2 <= n19038;
    G3674_o2 <= n19041;
    G3685_o2 <= n19044;
    G4504_o2 <= n19047;
    G4180_o2 <= n19050;
    G5123_o2 <= n19053;
    G5142_o2 <= n19056;
    G5126_o2 <= n19059;
    G5144_o2 <= n19062;
    G3912_o2 <= n19065;
    G4417_o2 <= n19068;
    G4420_o2 <= n19071;
    G3969_o2 <= n19074;
    G4023_o2 <= n19077;
    G2720_o2 <= n19080;
    G2837_o2 <= n19083;
    n2965_inv <= n19086;
    n2968_inv <= n19089;
    n2971_inv <= n19092;
    n2974_inv <= n19095;
    G1876_o2 <= n19098;
    G4996_o2 <= n19101;
    G4984_o2 <= n19104;
    G4920_o2 <= n19107;
    G4923_o2 <= n19110;
    G4930_o2 <= n19113;
    G4933_o2 <= n19116;
    n4320_lo_buf_o2 <= n19119;
    G2424_o2 <= n19122;
    G3317_o2 <= n19125;
    G3503_o2 <= n19128;
    G3485_o2 <= n19131;
    G3611_o2 <= n19134;
    n3864_lo_buf_o2 <= n19137;
    n3888_lo_buf_o2 <= n19140;
    n4116_lo_buf_o2 <= n19143;
    n4128_lo_buf_o2 <= n19146;
    n4140_lo_buf_o2 <= n19149;
    n4152_lo_buf_o2 <= n19152;
    G1815_o2 <= n19155;
    G1728_o2 <= n19158;
    G1035_o2 <= n19161;
    G1041_o2 <= n19164;
    G1087_o2 <= n19167;
    G1093_o2 <= n19170;
    G1132_o2 <= n19173;
    G1108_o2 <= n19176;
    G1138_o2 <= n19179;
    G1114_o2 <= n19182;
    G1807_o2 <= n19185;
    G2108_o2 <= n19188;
    G1126_o2 <= n19191;
    G1899_o2 <= n19194;
    G2134_o2 <= n19197;
    G1852_o2 <= n19200;
    G2116_o2 <= n19203;
    G2543_o2 <= n19206;
    G2727_o2 <= n19209;
    G2715_o2 <= n19212;
    G2832_o2 <= n19215;
    G1873_o2 <= n19218;
    G3291_o2 <= n19221;
    G5025_o2 <= n19224;
    G5036_o2 <= n19227;
    G3132_o2 <= n19230;
    G5038_o2 <= n19233;
    G5039_o2 <= n19236;
    n3118_inv <= n19239;
    n3121_inv <= n19242;
    n3124_inv <= n19245;
    n3127_inv <= n19248;
    n3984_lo_buf_o2 <= n19251;
    G1802_o2 <= n19254;
    G1804_o2 <= n19257;
    G1849_o2 <= n19260;
    G1851_o2 <= n19263;
    G2492_o2 <= n19266;
    G1799_o2 <= n19269;
    G4231_o2 <= n19272;
    G4234_o2 <= n19275;
    G4245_o2 <= n19278;
    G4247_o2 <= n19281;
    G1894_o2 <= n19284;
    G1846_o2 <= n19287;
    G4238_o2 <= n19290;
    G4249_o2 <= n19293;
    G2293_o2 <= n19296;
    G5022_o2 <= n19299;
    G5006_o2 <= n19302;
    G4944_o2 <= n19305;
    G4946_o2 <= n19308;
    G4954_o2 <= n19311;
    G4956_o2 <= n19314;
    G3546_o2 <= n19317;
    G3658_o2 <= n19320;
    G1344_o2 <= n19323;
    G2921_o2 <= n19326;
    n3912_lo_buf_o2 <= n19329;
    G1835_o2 <= n19332;
    G3810_o2 <= n19335;
    G3866_o2 <= n19338;
    G3811_o2 <= n19341;
    G2269_o2 <= n19344;
    G3812_o2 <= n19347;
    G3867_o2 <= n19350;
    G3868_o2 <= n19353;
    G3809_o2 <= n19356;
    G3716_o2 <= n19359;
    G4529_o2 <= n19362;
    G4670_o2 <= n19365;
    G4493_o2 <= n19368;
    G4580_o2 <= n19371;
    G3822_o2 <= n19374;
    G3877_o2 <= n19377;
    G4131_o2 <= n19380;
    G4170_o2 <= n19383;
    G4051_o2 <= n19386;
    G4065_o2 <= n19389;
    G4697_o2 <= n19392;
    G4706_o2 <= n19395;
    G2460_o2 <= n19398;
    G2454_o2 <= n19401;
    G2392_o2 <= n19404;
    G2386_o2 <= n19407;
    n4260_lo_buf_o2 <= n19410;
    n4272_lo_buf_o2 <= n19413;
    n4392_lo_buf_o2 <= n19416;
    n4404_lo_buf_o2 <= n19419;
    G1512_o2 <= n19422;
    G3135_o2 <= n19425;
    G2379_o2 <= n19428;
    n4164_lo_buf_o2 <= n19431;
    n4176_lo_buf_o2 <= n19434;
    n4224_lo_buf_o2 <= n19437;
    G2975_o2 <= n19440;
    G2978_o2 <= n19443;
    G2933_o2 <= n19446;
    G2936_o2 <= n19449;
    G1356_o2 <= n19452;
    G1359_o2 <= n19455;
    G1398_o2 <= n19458;
    G1401_o2 <= n19461;
  end
  initial begin
    n2610_lo <= 1'b0;
    n2613_lo <= 1'b0;
    n2616_lo <= 1'b0;
    n2619_lo <= 1'b0;
    n2622_lo <= 1'b0;
    n2625_lo <= 1'b0;
    n2628_lo <= 1'b0;
    n2631_lo <= 1'b0;
    n2634_lo <= 1'b0;
    n2637_lo <= 1'b0;
    n2640_lo <= 1'b0;
    n2643_lo <= 1'b0;
    n2646_lo <= 1'b0;
    n2649_lo <= 1'b0;
    n2652_lo <= 1'b0;
    n2655_lo <= 1'b0;
    n2658_lo <= 1'b0;
    n2661_lo <= 1'b0;
    n2664_lo <= 1'b0;
    n2667_lo <= 1'b0;
    n2670_lo <= 1'b0;
    n2673_lo <= 1'b0;
    n2676_lo <= 1'b0;
    n2679_lo <= 1'b0;
    n2682_lo <= 1'b0;
    n2685_lo <= 1'b0;
    n2688_lo <= 1'b0;
    n2691_lo <= 1'b0;
    n2694_lo <= 1'b0;
    n2697_lo <= 1'b0;
    n2700_lo <= 1'b0;
    n2703_lo <= 1'b0;
    n2706_lo <= 1'b0;
    n2709_lo <= 1'b0;
    n2712_lo <= 1'b0;
    n2715_lo <= 1'b0;
    n2718_lo <= 1'b0;
    n2721_lo <= 1'b0;
    n2724_lo <= 1'b0;
    n2727_lo <= 1'b0;
    n2730_lo <= 1'b0;
    n2733_lo <= 1'b0;
    n2736_lo <= 1'b0;
    n2739_lo <= 1'b0;
    n2742_lo <= 1'b0;
    n2745_lo <= 1'b0;
    n2748_lo <= 1'b0;
    n2751_lo <= 1'b0;
    n2754_lo <= 1'b0;
    n2757_lo <= 1'b0;
    n2760_lo <= 1'b0;
    n2763_lo <= 1'b0;
    n2766_lo <= 1'b0;
    n2769_lo <= 1'b0;
    n2772_lo <= 1'b0;
    n2775_lo <= 1'b0;
    n2778_lo <= 1'b0;
    n2781_lo <= 1'b0;
    n2784_lo <= 1'b0;
    n2787_lo <= 1'b0;
    n2790_lo <= 1'b0;
    n2793_lo <= 1'b0;
    n2796_lo <= 1'b0;
    n2799_lo <= 1'b0;
    n2802_lo <= 1'b0;
    n2805_lo <= 1'b0;
    n2808_lo <= 1'b0;
    n2811_lo <= 1'b0;
    n2814_lo <= 1'b0;
    n2817_lo <= 1'b0;
    n2820_lo <= 1'b0;
    n2823_lo <= 1'b0;
    n2826_lo <= 1'b0;
    n2829_lo <= 1'b0;
    n2832_lo <= 1'b0;
    n2835_lo <= 1'b0;
    n2838_lo <= 1'b0;
    n2841_lo <= 1'b0;
    n2844_lo <= 1'b0;
    n2847_lo <= 1'b0;
    n2850_lo <= 1'b0;
    n2853_lo <= 1'b0;
    n2856_lo <= 1'b0;
    n2859_lo <= 1'b0;
    n2862_lo <= 1'b0;
    n2865_lo <= 1'b0;
    n2868_lo <= 1'b0;
    n2871_lo <= 1'b0;
    n2874_lo <= 1'b0;
    n2877_lo <= 1'b0;
    n2880_lo <= 1'b0;
    n2883_lo <= 1'b0;
    n2886_lo <= 1'b0;
    n2889_lo <= 1'b0;
    n2892_lo <= 1'b0;
    n2895_lo <= 1'b0;
    n2898_lo <= 1'b0;
    n2901_lo <= 1'b0;
    n2904_lo <= 1'b0;
    n2907_lo <= 1'b0;
    n2910_lo <= 1'b0;
    n2913_lo <= 1'b0;
    n2916_lo <= 1'b0;
    n2919_lo <= 1'b0;
    n2922_lo <= 1'b0;
    n2925_lo <= 1'b0;
    n2928_lo <= 1'b0;
    n2931_lo <= 1'b0;
    n2934_lo <= 1'b0;
    n2937_lo <= 1'b0;
    n2940_lo <= 1'b0;
    n2943_lo <= 1'b0;
    n2946_lo <= 1'b0;
    n2949_lo <= 1'b0;
    n2952_lo <= 1'b0;
    n2955_lo <= 1'b0;
    n2958_lo <= 1'b0;
    n2961_lo <= 1'b0;
    n2964_lo <= 1'b0;
    n2967_lo <= 1'b0;
    n2970_lo <= 1'b0;
    n2973_lo <= 1'b0;
    n2976_lo <= 1'b0;
    n2979_lo <= 1'b0;
    n2982_lo <= 1'b0;
    n2985_lo <= 1'b0;
    n2988_lo <= 1'b0;
    n2991_lo <= 1'b0;
    n2994_lo <= 1'b0;
    n2997_lo <= 1'b0;
    n3000_lo <= 1'b0;
    n3003_lo <= 1'b0;
    n3006_lo <= 1'b0;
    n3009_lo <= 1'b0;
    n3012_lo <= 1'b0;
    n3015_lo <= 1'b0;
    n3018_lo <= 1'b0;
    n3021_lo <= 1'b0;
    n3024_lo <= 1'b0;
    n3027_lo <= 1'b0;
    n3030_lo <= 1'b0;
    n3033_lo <= 1'b0;
    n3036_lo <= 1'b0;
    n3039_lo <= 1'b0;
    n3042_lo <= 1'b0;
    n3045_lo <= 1'b0;
    n3048_lo <= 1'b0;
    n3051_lo <= 1'b0;
    n3054_lo <= 1'b0;
    n3057_lo <= 1'b0;
    n3060_lo <= 1'b0;
    n3063_lo <= 1'b0;
    n3066_lo <= 1'b0;
    n3069_lo <= 1'b0;
    n3072_lo <= 1'b0;
    n3075_lo <= 1'b0;
    n3078_lo <= 1'b0;
    n3081_lo <= 1'b0;
    n3084_lo <= 1'b0;
    n3087_lo <= 1'b0;
    n3090_lo <= 1'b0;
    n3093_lo <= 1'b0;
    n3096_lo <= 1'b0;
    n3099_lo <= 1'b0;
    n3102_lo <= 1'b0;
    n3105_lo <= 1'b0;
    n3108_lo <= 1'b0;
    n3111_lo <= 1'b0;
    n3114_lo <= 1'b0;
    n3117_lo <= 1'b0;
    n3120_lo <= 1'b0;
    n3123_lo <= 1'b0;
    n3126_lo <= 1'b0;
    n3129_lo <= 1'b0;
    n3132_lo <= 1'b0;
    n3135_lo <= 1'b0;
    n3138_lo <= 1'b0;
    n3141_lo <= 1'b0;
    n3144_lo <= 1'b0;
    n3147_lo <= 1'b0;
    n3150_lo <= 1'b0;
    n3153_lo <= 1'b0;
    n3156_lo <= 1'b0;
    n3159_lo <= 1'b0;
    n3162_lo <= 1'b0;
    n3165_lo <= 1'b0;
    n3168_lo <= 1'b0;
    n3171_lo <= 1'b0;
    n3174_lo <= 1'b0;
    n3177_lo <= 1'b0;
    n3180_lo <= 1'b0;
    n3183_lo <= 1'b0;
    n3186_lo <= 1'b0;
    n3189_lo <= 1'b0;
    n3192_lo <= 1'b0;
    n3195_lo <= 1'b0;
    n3198_lo <= 1'b0;
    n3201_lo <= 1'b0;
    n3204_lo <= 1'b0;
    n3207_lo <= 1'b0;
    n3210_lo <= 1'b0;
    n3213_lo <= 1'b0;
    n3216_lo <= 1'b0;
    n3219_lo <= 1'b0;
    n3222_lo <= 1'b0;
    n3225_lo <= 1'b0;
    n3228_lo <= 1'b0;
    n3231_lo <= 1'b0;
    n3234_lo <= 1'b0;
    n3237_lo <= 1'b0;
    n3240_lo <= 1'b0;
    n3243_lo <= 1'b0;
    n3246_lo <= 1'b0;
    n3249_lo <= 1'b0;
    n3252_lo <= 1'b0;
    n3255_lo <= 1'b0;
    n3258_lo <= 1'b0;
    n3261_lo <= 1'b0;
    n3264_lo <= 1'b0;
    n3267_lo <= 1'b0;
    n3270_lo <= 1'b0;
    n3273_lo <= 1'b0;
    n3276_lo <= 1'b0;
    n3279_lo <= 1'b0;
    n3282_lo <= 1'b0;
    n3285_lo <= 1'b0;
    n3288_lo <= 1'b0;
    n3291_lo <= 1'b0;
    n3294_lo <= 1'b0;
    n3297_lo <= 1'b0;
    n3300_lo <= 1'b0;
    n3303_lo <= 1'b0;
    n3306_lo <= 1'b0;
    n3309_lo <= 1'b0;
    n3312_lo <= 1'b0;
    n3315_lo <= 1'b0;
    n3318_lo <= 1'b0;
    n3321_lo <= 1'b0;
    n3324_lo <= 1'b0;
    n3327_lo <= 1'b0;
    n3330_lo <= 1'b0;
    n3333_lo <= 1'b0;
    n3336_lo <= 1'b0;
    n3339_lo <= 1'b0;
    n3342_lo <= 1'b0;
    n3345_lo <= 1'b0;
    n3348_lo <= 1'b0;
    n3351_lo <= 1'b0;
    n3354_lo <= 1'b0;
    n3357_lo <= 1'b0;
    n3360_lo <= 1'b0;
    n3363_lo <= 1'b0;
    n3366_lo <= 1'b0;
    n3369_lo <= 1'b0;
    n3372_lo <= 1'b0;
    n3375_lo <= 1'b0;
    n3378_lo <= 1'b0;
    n3381_lo <= 1'b0;
    n3384_lo <= 1'b0;
    n3387_lo <= 1'b0;
    n3390_lo <= 1'b0;
    n3393_lo <= 1'b0;
    n3396_lo <= 1'b0;
    n3399_lo <= 1'b0;
    n3402_lo <= 1'b0;
    n3405_lo <= 1'b0;
    n3408_lo <= 1'b0;
    n3411_lo <= 1'b0;
    n3414_lo <= 1'b0;
    n3417_lo <= 1'b0;
    n3420_lo <= 1'b0;
    n3423_lo <= 1'b0;
    n3426_lo <= 1'b0;
    n3429_lo <= 1'b0;
    n3432_lo <= 1'b0;
    n3435_lo <= 1'b0;
    n3438_lo <= 1'b0;
    n3441_lo <= 1'b0;
    n3444_lo <= 1'b0;
    n3447_lo <= 1'b0;
    n3450_lo <= 1'b0;
    n3453_lo <= 1'b0;
    n3456_lo <= 1'b0;
    n3459_lo <= 1'b0;
    n3462_lo <= 1'b0;
    n3465_lo <= 1'b0;
    n3468_lo <= 1'b0;
    n3471_lo <= 1'b0;
    n3474_lo <= 1'b0;
    n3477_lo <= 1'b0;
    n3480_lo <= 1'b0;
    n3483_lo <= 1'b0;
    n3486_lo <= 1'b0;
    n3489_lo <= 1'b0;
    n3492_lo <= 1'b0;
    n3495_lo <= 1'b0;
    n3498_lo <= 1'b0;
    n3501_lo <= 1'b0;
    n3504_lo <= 1'b0;
    n3507_lo <= 1'b0;
    n3510_lo <= 1'b0;
    n3513_lo <= 1'b0;
    n3516_lo <= 1'b0;
    n3519_lo <= 1'b0;
    n3522_lo <= 1'b0;
    n3525_lo <= 1'b0;
    n3528_lo <= 1'b0;
    n3531_lo <= 1'b0;
    n3534_lo <= 1'b0;
    n3537_lo <= 1'b0;
    n3540_lo <= 1'b0;
    n3543_lo <= 1'b0;
    n3546_lo <= 1'b0;
    n3549_lo <= 1'b0;
    n3552_lo <= 1'b0;
    n3555_lo <= 1'b0;
    n3558_lo <= 1'b0;
    n3561_lo <= 1'b0;
    n3564_lo <= 1'b0;
    n3567_lo <= 1'b0;
    n3570_lo <= 1'b0;
    n3573_lo <= 1'b0;
    n3576_lo <= 1'b0;
    n3579_lo <= 1'b0;
    n3582_lo <= 1'b0;
    n3585_lo <= 1'b0;
    n3588_lo <= 1'b0;
    n3591_lo <= 1'b0;
    n3594_lo <= 1'b0;
    n3597_lo <= 1'b0;
    n3600_lo <= 1'b0;
    n3603_lo <= 1'b0;
    n3606_lo <= 1'b0;
    n3609_lo <= 1'b0;
    n3612_lo <= 1'b0;
    n3615_lo <= 1'b0;
    n3618_lo <= 1'b0;
    n3621_lo <= 1'b0;
    n3624_lo <= 1'b0;
    n3627_lo <= 1'b0;
    n3630_lo <= 1'b0;
    n3633_lo <= 1'b0;
    n3636_lo <= 1'b0;
    n3639_lo <= 1'b0;
    n3642_lo <= 1'b0;
    n3645_lo <= 1'b0;
    n3648_lo <= 1'b0;
    n3651_lo <= 1'b0;
    n3654_lo <= 1'b0;
    n3657_lo <= 1'b0;
    n3666_lo <= 1'b0;
    n3669_lo <= 1'b0;
    n3678_lo <= 1'b0;
    n3687_lo <= 1'b0;
    n3690_lo <= 1'b0;
    n3702_lo <= 1'b0;
    n3711_lo <= 1'b0;
    n3714_lo <= 1'b0;
    n3726_lo <= 1'b0;
    n3735_lo <= 1'b0;
    n3738_lo <= 1'b0;
    n3750_lo <= 1'b0;
    n3753_lo <= 1'b0;
    n3759_lo <= 1'b0;
    n3762_lo <= 1'b0;
    n3765_lo <= 1'b0;
    n3774_lo <= 1'b0;
    n3777_lo <= 1'b0;
    n3786_lo <= 1'b0;
    n3789_lo <= 1'b0;
    n3792_lo <= 1'b0;
    n3795_lo <= 1'b0;
    n3798_lo <= 1'b0;
    n3801_lo <= 1'b0;
    n3810_lo <= 1'b0;
    n3813_lo <= 1'b0;
    n3822_lo <= 1'b0;
    n3825_lo <= 1'b0;
    n3834_lo <= 1'b0;
    n3843_lo <= 1'b0;
    n3846_lo <= 1'b0;
    n3867_lo <= 1'b0;
    n3891_lo <= 1'b0;
    n3915_lo <= 1'b0;
    n3930_lo <= 1'b0;
    n3933_lo <= 1'b0;
    n3936_lo <= 1'b0;
    n3942_lo <= 1'b0;
    n3945_lo <= 1'b0;
    n3948_lo <= 1'b0;
    n3954_lo <= 1'b0;
    n3957_lo <= 1'b0;
    n3963_lo <= 1'b0;
    n3966_lo <= 1'b0;
    n3969_lo <= 1'b0;
    n3975_lo <= 1'b0;
    n3978_lo <= 1'b0;
    n3987_lo <= 1'b0;
    n3990_lo <= 1'b0;
    n4002_lo <= 1'b0;
    n4011_lo <= 1'b0;
    n4014_lo <= 1'b0;
    n4026_lo <= 1'b0;
    n4035_lo <= 1'b0;
    n4038_lo <= 1'b0;
    n4050_lo <= 1'b0;
    n4053_lo <= 1'b0;
    n4059_lo <= 1'b0;
    n4062_lo <= 1'b0;
    n4065_lo <= 1'b0;
    n4098_lo <= 1'b0;
    n4107_lo <= 1'b0;
    n4119_lo <= 1'b0;
    n4131_lo <= 1'b0;
    n4143_lo <= 1'b0;
    n4155_lo <= 1'b0;
    n4167_lo <= 1'b0;
    n4179_lo <= 1'b0;
    n4182_lo <= 1'b0;
    n4185_lo <= 1'b0;
    n4188_lo <= 1'b0;
    n4194_lo <= 1'b0;
    n4197_lo <= 1'b0;
    n4200_lo <= 1'b0;
    n4206_lo <= 1'b0;
    n4209_lo <= 1'b0;
    n4212_lo <= 1'b0;
    n4215_lo <= 1'b0;
    n4227_lo <= 1'b0;
    n4230_lo <= 1'b0;
    n4233_lo <= 1'b0;
    n4236_lo <= 1'b0;
    n4239_lo <= 1'b0;
    n4242_lo <= 1'b0;
    n4251_lo <= 1'b0;
    n4263_lo <= 1'b0;
    n4275_lo <= 1'b0;
    n4278_lo <= 1'b0;
    n4287_lo <= 1'b0;
    n4290_lo <= 1'b0;
    n4293_lo <= 1'b0;
    n4299_lo <= 1'b0;
    n4302_lo <= 1'b0;
    n4305_lo <= 1'b0;
    n4311_lo <= 1'b0;
    n4314_lo <= 1'b0;
    n4323_lo <= 1'b0;
    n4326_lo <= 1'b0;
    n4335_lo <= 1'b0;
    n4338_lo <= 1'b0;
    n4347_lo <= 1'b0;
    n4350_lo <= 1'b0;
    n4359_lo <= 1'b0;
    n4362_lo <= 1'b0;
    n4365_lo <= 1'b0;
    n4371_lo <= 1'b0;
    n4374_lo <= 1'b0;
    n4383_lo <= 1'b0;
    n4395_lo <= 1'b0;
    n4407_lo <= 1'b0;
    n4410_lo <= 1'b0;
    n4413_lo <= 1'b0;
    n4416_lo <= 1'b0;
    n4419_lo <= 1'b0;
    n4422_lo <= 1'b0;
    n4425_lo <= 1'b0;
    n4428_lo <= 1'b0;
    n4431_lo <= 1'b0;
    n4434_lo <= 1'b0;
    n4437_lo <= 1'b0;
    n4440_lo <= 1'b0;
    n4443_lo <= 1'b0;
    n4446_lo <= 1'b0;
    n4449_lo <= 1'b0;
    n4452_lo <= 1'b0;
    n4455_lo <= 1'b0;
    n4458_lo <= 1'b0;
    n4461_lo <= 1'b0;
    n4464_lo <= 1'b0;
    n4467_lo <= 1'b0;
    n4470_lo <= 1'b0;
    n4473_lo <= 1'b0;
    n4476_lo <= 1'b0;
    n4479_lo <= 1'b0;
    n4482_lo <= 1'b0;
    n4485_lo <= 1'b0;
    n4488_lo <= 1'b0;
    n4494_lo <= 1'b0;
    n4497_lo <= 1'b0;
    n4500_lo <= 1'b0;
    n4503_lo <= 1'b0;
    n4506_lo <= 1'b0;
    n4509_lo <= 1'b0;
    n4512_lo <= 1'b0;
    n4515_lo <= 1'b0;
    n4518_lo <= 1'b0;
    n4521_lo <= 1'b0;
    n4524_lo <= 1'b0;
    n4527_lo <= 1'b0;
    n4530_lo <= 1'b0;
    n4533_lo <= 1'b0;
    n4536_lo <= 1'b0;
    n4539_lo <= 1'b0;
    n4542_lo <= 1'b0;
    n4545_lo <= 1'b0;
    n4548_lo <= 1'b0;
    n4554_lo <= 1'b0;
    n4557_lo <= 1'b0;
    n4560_lo <= 1'b0;
    n4563_lo <= 1'b0;
    n4566_lo <= 1'b0;
    n4569_lo <= 1'b0;
    n4572_lo <= 1'b0;
    n4575_lo <= 1'b0;
    n4578_lo <= 1'b0;
    n4581_lo <= 1'b0;
    n4584_lo <= 1'b0;
    n4587_lo <= 1'b0;
    n4590_lo <= 1'b0;
    n4593_lo <= 1'b0;
    n4596_lo <= 1'b0;
    n4599_lo <= 1'b0;
    n4602_lo <= 1'b0;
    n4605_lo <= 1'b0;
    n4608_lo <= 1'b0;
    n4611_lo <= 1'b0;
    n4614_lo <= 1'b0;
    n4617_lo <= 1'b0;
    n4620_lo <= 1'b0;
    n4623_lo <= 1'b0;
    n4626_lo <= 1'b0;
    n4629_lo <= 1'b0;
    n4632_lo <= 1'b0;
    n4635_lo <= 1'b0;
    n4638_lo <= 1'b0;
    n4641_lo <= 1'b0;
    n4644_lo <= 1'b0;
    n4647_lo <= 1'b0;
    n4650_lo <= 1'b0;
    n4653_lo <= 1'b0;
    n4656_lo <= 1'b0;
    n4659_lo <= 1'b0;
    n4662_lo <= 1'b0;
    n4665_lo <= 1'b0;
    n4668_lo <= 1'b0;
    n4671_lo <= 1'b0;
    n4674_lo <= 1'b0;
    n4677_lo <= 1'b0;
    n4680_lo <= 1'b0;
    n4683_lo <= 1'b0;
    n4686_lo <= 1'b0;
    n4689_lo <= 1'b0;
    n4692_lo <= 1'b0;
    n4695_lo <= 1'b0;
    n4698_lo <= 1'b0;
    n4701_lo <= 1'b0;
    n4704_lo <= 1'b0;
    n4707_lo <= 1'b0;
    n4710_lo <= 1'b0;
    n4713_lo <= 1'b0;
    n4716_lo <= 1'b0;
    n4719_lo <= 1'b0;
    n4722_lo <= 1'b0;
    n4725_lo <= 1'b0;
    n4728_lo <= 1'b0;
    n4731_lo <= 1'b0;
    n4734_lo <= 1'b0;
    n4737_lo <= 1'b0;
    n4740_lo <= 1'b0;
    n4743_lo <= 1'b0;
    n6382_o2 <= 1'b0;
    n6383_o2 <= 1'b0;
    n6419_o2 <= 1'b0;
    n6420_o2 <= 1'b0;
    n6435_o2 <= 1'b0;
    n6436_o2 <= 1'b0;
    n6448_o2 <= 1'b0;
    n6449_o2 <= 1'b0;
    n6613_o2 <= 1'b0;
    n6614_o2 <= 1'b0;
    n6641_o2 <= 1'b0;
    n6658_o2 <= 1'b0;
    n6757_o2 <= 1'b0;
    n6756_o2 <= 1'b0;
    n7116_o2 <= 1'b0;
    n7156_o2 <= 1'b0;
    n6549_o2 <= 1'b0;
    n6550_o2 <= 1'b0;
    n7357_o2 <= 1'b0;
    n7358_o2 <= 1'b0;
    n7359_o2 <= 1'b0;
    n7360_o2 <= 1'b0;
    n6621_o2 <= 1'b0;
    n6623_o2 <= 1'b0;
    n6625_o2 <= 1'b0;
    n6626_o2 <= 1'b0;
    n6627_o2 <= 1'b0;
    n6628_o2 <= 1'b0;
    n6629_o2 <= 1'b0;
    n6630_o2 <= 1'b0;
    n6669_o2 <= 1'b0;
    n7449_o2 <= 1'b0;
    n7450_o2 <= 1'b0;
    n7451_o2 <= 1'b0;
    n7452_o2 <= 1'b0;
    n6682_o2 <= 1'b0;
    n6683_o2 <= 1'b0;
    n6684_o2 <= 1'b0;
    n6685_o2 <= 1'b0;
    n7463_o2 <= 1'b0;
    n6686_o2 <= 1'b0;
    n6687_o2 <= 1'b0;
    n6688_o2 <= 1'b0;
    n6689_o2 <= 1'b0;
    n6772_o2 <= 1'b0;
    n6773_o2 <= 1'b0;
    n6774_o2 <= 1'b0;
    n6775_o2 <= 1'b0;
    G3467_o2 <= 1'b0;
    G2810_o2 <= 1'b0;
    n6833_o2 <= 1'b0;
    n6945_o2 <= 1'b0;
    n6947_o2 <= 1'b0;
    n6949_o2 <= 1'b0;
    n6951_o2 <= 1'b0;
    n6888_o2 <= 1'b0;
    n6889_o2 <= 1'b0;
    n6936_o2 <= 1'b0;
    n6954_o2 <= 1'b0;
    n6955_o2 <= 1'b0;
    n6956_o2 <= 1'b0;
    n6957_o2 <= 1'b0;
    n6958_o2 <= 1'b0;
    n6982_o2 <= 1'b0;
    n6984_o2 <= 1'b0;
    n6974_o2 <= 1'b0;
    n6975_o2 <= 1'b0;
    n6999_o2 <= 1'b0;
    n7015_o2 <= 1'b0;
    n7016_o2 <= 1'b0;
    n7017_o2 <= 1'b0;
    n7018_o2 <= 1'b0;
    n7005_o2 <= 1'b0;
    n7019_o2 <= 1'b0;
    n7022_o2 <= 1'b0;
    n7023_o2 <= 1'b0;
    n7132_o2 <= 1'b0;
    n7133_o2 <= 1'b0;
    n7135_o2 <= 1'b0;
    n7136_o2 <= 1'b0;
    n7175_o2 <= 1'b0;
    n7155_o2 <= 1'b0;
    G3060_o2 <= 1'b0;
    n7383_o2 <= 1'b0;
    G3802_o2 <= 1'b0;
    G3859_o2 <= 1'b0;
    n7355_o2 <= 1'b0;
    n7356_o2 <= 1'b0;
    G4054_o2 <= 1'b0;
    G4068_o2 <= 1'b0;
    n7384_o2 <= 1'b0;
    n7387_o2 <= 1'b0;
    n7388_o2 <= 1'b0;
    n7389_o2 <= 1'b0;
    n7386_o2 <= 1'b0;
    n7453_o2 <= 1'b0;
    n7431_o2 <= 1'b0;
    n7432_o2 <= 1'b0;
    n7433_o2 <= 1'b0;
    n7430_o2 <= 1'b0;
    n7485_o2 <= 1'b0;
    n7486_o2 <= 1'b0;
    G2508_o2 <= 1'b0;
    G2486_o2 <= 1'b0;
    n2326_inv <= 1'b0;
    n2329_inv <= 1'b0;
    n3756_lo_buf_o2 <= 1'b0;
    n4056_lo_buf_o2 <= 1'b0;
    G3474_o2 <= 1'b0;
    n2341_inv <= 1'b0;
    n7396_o2 <= 1'b0;
    n7398_o2 <= 1'b0;
    n7400_o2 <= 1'b0;
    n7401_o2 <= 1'b0;
    n7402_o2 <= 1'b0;
    n7403_o2 <= 1'b0;
    n7404_o2 <= 1'b0;
    n7405_o2 <= 1'b0;
    G2711_o2 <= 1'b0;
    n2371_inv <= 1'b0;
    n7490_o2 <= 1'b0;
    n7527_o2 <= 1'b0;
    n7528_o2 <= 1'b0;
    n7529_o2 <= 1'b0;
    n7530_o2 <= 1'b0;
    n7523_o2 <= 1'b0;
    n7524_o2 <= 1'b0;
    n7525_o2 <= 1'b0;
    n7526_o2 <= 1'b0;
    n4296_lo_buf_o2 <= 1'b0;
    n4368_lo_buf_o2 <= 1'b0;
    G2466_o2 <= 1'b0;
    G2404_o2 <= 1'b0;
    n7534_o2 <= 1'b0;
    n7535_o2 <= 1'b0;
    n7536_o2 <= 1'b0;
    n7533_o2 <= 1'b0;
    G1060_o2 <= 1'b0;
    G963_o2 <= 1'b0;
    G2448_o2 <= 1'b0;
    G2685_o2 <= 1'b0;
    G2679_o2 <= 1'b0;
    G2774_o2 <= 1'b0;
    G2780_o2 <= 1'b0;
    G2759_o2 <= 1'b0;
    G2737_o2 <= 1'b0;
    G2850_o2 <= 1'b0;
    G3393_o2 <= 1'b0;
    G3404_o2 <= 1'b0;
    G3559_o2 <= 1'b0;
    G2744_o2 <= 1'b0;
    n3708_lo_buf_o2 <= 1'b0;
    n3840_lo_buf_o2 <= 1'b0;
    n4008_lo_buf_o2 <= 1'b0;
    n4104_lo_buf_o2 <= 1'b0;
    G1821_o2 <= 1'b0;
    G1734_o2 <= 1'b0;
    G3517_o2 <= 1'b0;
    G3533_o2 <= 1'b0;
    G3629_o2 <= 1'b0;
    G3645_o2 <= 1'b0;
    n2497_inv <= 1'b0;
    G2731_o2 <= 1'b0;
    G2844_o2 <= 1'b0;
    n3732_lo_buf_o2 <= 1'b0;
    n4032_lo_buf_o2 <= 1'b0;
    G3552_o2 <= 1'b0;
    G2271_o2 <= 1'b0;
    n4248_lo_buf_o2 <= 1'b0;
    n4332_lo_buf_o2 <= 1'b0;
    n4344_lo_buf_o2 <= 1'b0;
    n4380_lo_buf_o2 <= 1'b0;
    G2398_o2 <= 1'b0;
    G2480_o2 <= 1'b0;
    G2418_o2 <= 1'b0;
    G1455_o2 <= 1'b0;
    G1449_o2 <= 1'b0;
    G1452_o2 <= 1'b0;
    G1425_o2 <= 1'b0;
    G1428_o2 <= 1'b0;
    G1419_o2 <= 1'b0;
    G1422_o2 <= 1'b0;
    n4308_lo_buf_o2 <= 1'b0;
    G2675_o2 <= 1'b0;
    G3035_o2 <= 1'b0;
    G3026_o2 <= 1'b0;
    G3029_o2 <= 1'b0;
    G3032_o2 <= 1'b0;
    G2999_o2 <= 1'b0;
    G3002_o2 <= 1'b0;
    G2770_o2 <= 1'b0;
    G3008_o2 <= 1'b0;
    G2073_o2 <= 1'b0;
    G2752_o2 <= 1'b0;
    G3005_o2 <= 1'b0;
    G5108_o2 <= 1'b0;
    G5135_o2 <= 1'b0;
    G5111_o2 <= 1'b0;
    G5138_o2 <= 1'b0;
    G3415_o2 <= 1'b0;
    G3386_o2 <= 1'b0;
    G3570_o2 <= 1'b0;
    G2430_o2 <= 1'b0;
    G3495_o2 <= 1'b0;
    G3621_o2 <= 1'b0;
    n4284_lo_buf_o2 <= 1'b0;
    n4356_lo_buf_o2 <= 1'b0;
    G2472_o2 <= 1'b0;
    G2410_o2 <= 1'b0;
    n3960_lo_buf_o2 <= 1'b0;
    n3972_lo_buf_o2 <= 1'b0;
    n2647_inv <= 1'b0;
    n2650_inv <= 1'b0;
    n3684_lo_buf_o2 <= 1'b0;
    n4080_lo_buf_o2 <= 1'b0;
    n4092_lo_buf_o2 <= 1'b0;
    n2662_inv <= 1'b0;
    n2665_inv <= 1'b0;
    G1147_o2 <= 1'b0;
    G2705_o2 <= 1'b0;
    G2693_o2 <= 1'b0;
    G2696_o2 <= 1'b0;
    G2700_o2 <= 1'b0;
    G2915_o2 <= 1'b0;
    G2966_o2 <= 1'b0;
    G2540_o2 <= 1'b0;
    G2788_o2 <= 1'b0;
    G2792_o2 <= 1'b0;
    G2797_o2 <= 1'b0;
    G2804_o2 <= 1'b0;
    G1038_o2 <= 1'b0;
    G1044_o2 <= 1'b0;
    G1090_o2 <= 1'b0;
    G1096_o2 <= 1'b0;
    G1029_o2 <= 1'b0;
    G3942_o2 <= 1'b0;
    G3954_o2 <= 1'b0;
    G4011_o2 <= 1'b0;
    G4017_o2 <= 1'b0;
    G1141_o2 <= 1'b0;
    G1081_o2 <= 1'b0;
    G2146_o2 <= 1'b0;
    G2145_o2 <= 1'b0;
    G2144_o2 <= 1'b0;
    G2143_o2 <= 1'b0;
    G2142_o2 <= 1'b0;
    G2141_o2 <= 1'b0;
    G2140_o2 <= 1'b0;
    G2139_o2 <= 1'b0;
    G3769_o2 <= 1'b0;
    G3773_o2 <= 1'b0;
    G3768_o2 <= 1'b0;
    G4101_o2 <= 1'b0;
    G3161_o2 <= 1'b0;
    G4143_o2 <= 1'b0;
    G3828_o2 <= 1'b0;
    G3831_o2 <= 1'b0;
    G3334_o2 <= 1'b0;
    G3335_o2 <= 1'b0;
    G3180_o2 <= 1'b0;
    G3340_o2 <= 1'b0;
    G3339_o2 <= 1'b0;
    G3341_o2 <= 1'b0;
    G3234_o2 <= 1'b0;
    G3829_o2 <= 1'b0;
    G3338_o2 <= 1'b0;
    G3336_o2 <= 1'b0;
    G3770_o2 <= 1'b0;
    G3918_o2 <= 1'b0;
    G3774_o2 <= 1'b0;
    G3921_o2 <= 1'b0;
    G3832_o2 <= 1'b0;
    G3993_o2 <= 1'b0;
    G2076_o2 <= 1'b0;
    G2071_o2 <= 1'b0;
    G2072_o2 <= 1'b0;
    G2069_o2 <= 1'b0;
    G2070_o2 <= 1'b0;
    G2067_o2 <= 1'b0;
    G2068_o2 <= 1'b0;
    G4095_o2 <= 1'b0;
    G3272_o2 <= 1'b0;
    G3269_o2 <= 1'b0;
    G3270_o2 <= 1'b0;
    G3271_o2 <= 1'b0;
    G3265_o2 <= 1'b0;
    G3266_o2 <= 1'b0;
    G4137_o2 <= 1'b0;
    G3268_o2 <= 1'b0;
    G2361_o2 <= 1'b0;
    G3228_o2 <= 1'b0;
    G3267_o2 <= 1'b0;
    G2336_o2 <= 1'b0;
    G3459_o2 <= 1'b0;
    G3428_o2 <= 1'b0;
    G3438_o2 <= 1'b0;
    G3449_o2 <= 1'b0;
    G3421_o2 <= 1'b0;
    G3576_o2 <= 1'b0;
    G3303_o2 <= 1'b0;
    G3583_o2 <= 1'b0;
    G3594_o2 <= 1'b0;
    G3674_o2 <= 1'b0;
    G3685_o2 <= 1'b0;
    G4504_o2 <= 1'b0;
    G4180_o2 <= 1'b0;
    G5123_o2 <= 1'b0;
    G5142_o2 <= 1'b0;
    G5126_o2 <= 1'b0;
    G5144_o2 <= 1'b0;
    G3912_o2 <= 1'b0;
    G4417_o2 <= 1'b0;
    G4420_o2 <= 1'b0;
    G3969_o2 <= 1'b0;
    G4023_o2 <= 1'b0;
    G2720_o2 <= 1'b0;
    G2837_o2 <= 1'b0;
    n2965_inv <= 1'b0;
    n2968_inv <= 1'b0;
    n2971_inv <= 1'b0;
    n2974_inv <= 1'b0;
    G1876_o2 <= 1'b0;
    G4996_o2 <= 1'b0;
    G4984_o2 <= 1'b0;
    G4920_o2 <= 1'b0;
    G4923_o2 <= 1'b0;
    G4930_o2 <= 1'b0;
    G4933_o2 <= 1'b0;
    n4320_lo_buf_o2 <= 1'b0;
    G2424_o2 <= 1'b0;
    G3317_o2 <= 1'b0;
    G3503_o2 <= 1'b0;
    G3485_o2 <= 1'b0;
    G3611_o2 <= 1'b0;
    n3864_lo_buf_o2 <= 1'b0;
    n3888_lo_buf_o2 <= 1'b0;
    n4116_lo_buf_o2 <= 1'b0;
    n4128_lo_buf_o2 <= 1'b0;
    n4140_lo_buf_o2 <= 1'b0;
    n4152_lo_buf_o2 <= 1'b0;
    G1815_o2 <= 1'b0;
    G1728_o2 <= 1'b0;
    G1035_o2 <= 1'b0;
    G1041_o2 <= 1'b0;
    G1087_o2 <= 1'b0;
    G1093_o2 <= 1'b0;
    G1132_o2 <= 1'b0;
    G1108_o2 <= 1'b0;
    G1138_o2 <= 1'b0;
    G1114_o2 <= 1'b0;
    G1807_o2 <= 1'b0;
    G2108_o2 <= 1'b0;
    G1126_o2 <= 1'b0;
    G1899_o2 <= 1'b0;
    G2134_o2 <= 1'b0;
    G1852_o2 <= 1'b0;
    G2116_o2 <= 1'b0;
    G2543_o2 <= 1'b0;
    G2727_o2 <= 1'b0;
    G2715_o2 <= 1'b0;
    G2832_o2 <= 1'b0;
    G1873_o2 <= 1'b0;
    G3291_o2 <= 1'b0;
    G5025_o2 <= 1'b0;
    G5036_o2 <= 1'b0;
    G3132_o2 <= 1'b0;
    G5038_o2 <= 1'b0;
    G5039_o2 <= 1'b0;
    n3118_inv <= 1'b0;
    n3121_inv <= 1'b0;
    n3124_inv <= 1'b0;
    n3127_inv <= 1'b0;
    n3984_lo_buf_o2 <= 1'b0;
    G1802_o2 <= 1'b0;
    G1804_o2 <= 1'b0;
    G1849_o2 <= 1'b0;
    G1851_o2 <= 1'b0;
    G2492_o2 <= 1'b0;
    G1799_o2 <= 1'b0;
    G4231_o2 <= 1'b0;
    G4234_o2 <= 1'b0;
    G4245_o2 <= 1'b0;
    G4247_o2 <= 1'b0;
    G1894_o2 <= 1'b0;
    G1846_o2 <= 1'b0;
    G4238_o2 <= 1'b0;
    G4249_o2 <= 1'b0;
    G2293_o2 <= 1'b0;
    G5022_o2 <= 1'b0;
    G5006_o2 <= 1'b0;
    G4944_o2 <= 1'b0;
    G4946_o2 <= 1'b0;
    G4954_o2 <= 1'b0;
    G4956_o2 <= 1'b0;
    G3546_o2 <= 1'b0;
    G3658_o2 <= 1'b0;
    G1344_o2 <= 1'b0;
    G2921_o2 <= 1'b0;
    n3912_lo_buf_o2 <= 1'b0;
    G1835_o2 <= 1'b0;
    G3810_o2 <= 1'b0;
    G3866_o2 <= 1'b0;
    G3811_o2 <= 1'b0;
    G2269_o2 <= 1'b0;
    G3812_o2 <= 1'b0;
    G3867_o2 <= 1'b0;
    G3868_o2 <= 1'b0;
    G3809_o2 <= 1'b0;
    G3716_o2 <= 1'b0;
    G4529_o2 <= 1'b0;
    G4670_o2 <= 1'b0;
    G4493_o2 <= 1'b0;
    G4580_o2 <= 1'b0;
    G3822_o2 <= 1'b0;
    G3877_o2 <= 1'b0;
    G4131_o2 <= 1'b0;
    G4170_o2 <= 1'b0;
    G4051_o2 <= 1'b0;
    G4065_o2 <= 1'b0;
    G4697_o2 <= 1'b0;
    G4706_o2 <= 1'b0;
    G2460_o2 <= 1'b0;
    G2454_o2 <= 1'b0;
    G2392_o2 <= 1'b0;
    G2386_o2 <= 1'b0;
    n4260_lo_buf_o2 <= 1'b0;
    n4272_lo_buf_o2 <= 1'b0;
    n4392_lo_buf_o2 <= 1'b0;
    n4404_lo_buf_o2 <= 1'b0;
    G1512_o2 <= 1'b0;
    G3135_o2 <= 1'b0;
    G2379_o2 <= 1'b0;
    n4164_lo_buf_o2 <= 1'b0;
    n4176_lo_buf_o2 <= 1'b0;
    n4224_lo_buf_o2 <= 1'b0;
    G2975_o2 <= 1'b0;
    G2978_o2 <= 1'b0;
    G2933_o2 <= 1'b0;
    G2936_o2 <= 1'b0;
    G1356_o2 <= 1'b0;
    G1359_o2 <= 1'b0;
    G1398_o2 <= 1'b0;
    G1401_o2 <= 1'b0;
  end
endmodule


