// Benchmark "c6288" written by ABC on Sun Oct 29 22:18:03 2023

module c6288 ( 
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32,
    G6257, G6258, G6259, G6260, G6261, G6262, G6263, G6264, G6265, G6266,
    G6267, G6268, G6269, G6270, G6271, G6272, G6273, G6274, G6275, G6276,
    G6277, G6278, G6279, G6280, G6281, G6282, G6283, G6284, G6285, G6286,
    G6287, G6288  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32;
  output G6257, G6258, G6259, G6260, G6261, G6262, G6263, G6264, G6265, G6266,
    G6267, G6268, G6269, G6270, G6271, G6272, G6273, G6274, G6275, G6276,
    G6277, G6278, G6279, G6280, G6281, G6282, G6283, G6284, G6285, G6286,
    G6287, G6288;
  wire new_n66_, new_n67_, new_n68_, new_n69_, new_n71_, new_n72_, new_n73_,
    new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_,
    new_n81_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_,
    new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_,
    new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n131_, new_n132_, new_n133_,
    new_n134_, new_n135_, new_n136_, new_n137_, new_n138_, new_n139_,
    new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_,
    new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_,
    new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_,
    new_n164_, new_n165_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_,
    new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_,
    new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1081_,
    new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_,
    new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_,
    new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_,
    new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_,
    new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_,
    new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_,
    new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_,
    new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_,
    new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_,
    new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_,
    new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_,
    new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_,
    new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_,
    new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_,
    new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_,
    new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_,
    new_n1190_, new_n1191_, new_n1193_, new_n1194_, new_n1195_, new_n1196_,
    new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_,
    new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_,
    new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_,
    new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_,
    new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_,
    new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_,
    new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_,
    new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_,
    new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_,
    new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_,
    new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_,
    new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_,
    new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_,
    new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_,
    new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_,
    new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_,
    new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_,
    new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_,
    new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_,
    new_n1481_, new_n1482_, new_n1484_, new_n1485_, new_n1486_, new_n1487_,
    new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_,
    new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_,
    new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_,
    new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1638_, new_n1639_,
    new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_,
    new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_,
    new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_,
    new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_,
    new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_,
    new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_,
    new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_,
    new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_,
    new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_,
    new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_,
    new_n1700_, new_n1701_, new_n1703_, new_n1704_, new_n1705_, new_n1706_,
    new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_,
    new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_,
    new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_,
    new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_,
    new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_,
    new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_,
    new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_,
    new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1760_, new_n1761_,
    new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_,
    new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_,
    new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_,
    new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_,
    new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_,
    new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_,
    new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_,
    new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1809_, new_n1810_,
    new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_,
    new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_,
    new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_,
    new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_,
    new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_,
    new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_,
    new_n1847_, new_n1848_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_,
    new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_,
    new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_,
    new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_,
    new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1908_, new_n1909_,
    new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_,
    new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_,
    new_n1922_, new_n1923_, new_n1925_, new_n1926_, new_n1927_, new_n1928_,
    new_n1929_, new_n1930_, new_n1931_, new_n1933_;
  and1 g0000(.dina(G1), .dinb(G17), .dout(G6257));
  nor2 g0001(.dina(G2), .dinb(G17), .dout(new_n66_));
  and1 g0002(.dina(G1), .dinb(G18), .dout(new_n67_));
  anb2 g0003(.dina(new_n66_), .dinb(new_n67_), .dout(new_n68_));
  anb1 g0004(.dina(new_n66_), .dinb(new_n67_), .dout(new_n69_));
  anb1 g0005(.dina(new_n68_), .dinb(new_n69_), .dout(G6258));
  nor2 g0006(.dina(G1), .dinb(G19), .dout(new_n71_));
  nor2 g0007(.dina(G3), .dinb(G17), .dout(new_n72_));
  and1 g0008(.dina(G2), .dinb(G18), .dout(new_n73_));
  anb2 g0009(.dina(new_n72_), .dinb(new_n73_), .dout(new_n74_));
  anb1 g0010(.dina(new_n72_), .dinb(new_n73_), .dout(new_n75_));
  anb1 g0011(.dina(new_n74_), .dinb(new_n75_), .dout(new_n76_));
  anb1 g0012(.dina(new_n68_), .dinb(new_n76_), .dout(new_n77_));
  anb2 g0013(.dina(new_n68_), .dinb(new_n76_), .dout(new_n78_));
  anb2 g0014(.dina(new_n77_), .dinb(new_n78_), .dout(new_n79_));
  anb1 g0015(.dina(new_n71_), .dinb(new_n79_), .dout(new_n80_));
  anb2 g0016(.dina(new_n71_), .dinb(new_n79_), .dout(new_n81_));
  anb2 g0017(.dina(new_n80_), .dinb(new_n81_), .dout(G6259));
  nor2 g0018(.dina(G1), .dinb(G20), .dout(new_n83_));
  and2 g0019(.dina(new_n77_), .dinb(new_n80_), .dout(new_n84_));
  nor2 g0020(.dina(G2), .dinb(G19), .dout(new_n85_));
  nor2 g0021(.dina(G4), .dinb(G17), .dout(new_n86_));
  and1 g0022(.dina(G3), .dinb(G18), .dout(new_n87_));
  anb2 g0023(.dina(new_n86_), .dinb(new_n87_), .dout(new_n88_));
  anb1 g0024(.dina(new_n86_), .dinb(new_n87_), .dout(new_n89_));
  anb1 g0025(.dina(new_n88_), .dinb(new_n89_), .dout(new_n90_));
  anb1 g0026(.dina(new_n74_), .dinb(new_n90_), .dout(new_n91_));
  anb2 g0027(.dina(new_n74_), .dinb(new_n90_), .dout(new_n92_));
  anb2 g0028(.dina(new_n91_), .dinb(new_n92_), .dout(new_n93_));
  anb1 g0029(.dina(new_n85_), .dinb(new_n93_), .dout(new_n94_));
  anb2 g0030(.dina(new_n85_), .dinb(new_n93_), .dout(new_n95_));
  anb2 g0031(.dina(new_n94_), .dinb(new_n95_), .dout(new_n96_));
  anb1 g0032(.dina(new_n84_), .dinb(new_n96_), .dout(new_n97_));
  anb2 g0033(.dina(new_n84_), .dinb(new_n96_), .dout(new_n98_));
  anb2 g0034(.dina(new_n97_), .dinb(new_n98_), .dout(new_n99_));
  anb1 g0035(.dina(new_n83_), .dinb(new_n99_), .dout(new_n100_));
  anb2 g0036(.dina(new_n83_), .dinb(new_n99_), .dout(new_n101_));
  anb2 g0037(.dina(new_n100_), .dinb(new_n101_), .dout(G6260));
  nor2 g0038(.dina(G1), .dinb(G21), .dout(new_n103_));
  and2 g0039(.dina(new_n97_), .dinb(new_n100_), .dout(new_n104_));
  nor2 g0040(.dina(G2), .dinb(G20), .dout(new_n105_));
  and2 g0041(.dina(new_n91_), .dinb(new_n94_), .dout(new_n106_));
  nor2 g0042(.dina(G3), .dinb(G19), .dout(new_n107_));
  and1 g0043(.dina(G5), .dinb(G17), .dout(new_n108_));
  nor2 g0044(.dina(G4), .dinb(G18), .dout(new_n109_));
  anb1 g0045(.dina(new_n108_), .dinb(new_n109_), .dout(new_n110_));
  anb2 g0046(.dina(new_n108_), .dinb(new_n109_), .dout(new_n111_));
  nab1 g0047(.dina(new_n110_), .dinb(new_n111_), .dout(new_n112_));
  anb1 g0048(.dina(new_n88_), .dinb(new_n112_), .dout(new_n113_));
  anb2 g0049(.dina(new_n88_), .dinb(new_n112_), .dout(new_n114_));
  anb2 g0050(.dina(new_n113_), .dinb(new_n114_), .dout(new_n115_));
  anb1 g0051(.dina(new_n107_), .dinb(new_n115_), .dout(new_n116_));
  anb2 g0052(.dina(new_n107_), .dinb(new_n115_), .dout(new_n117_));
  anb2 g0053(.dina(new_n116_), .dinb(new_n117_), .dout(new_n118_));
  anb1 g0054(.dina(new_n106_), .dinb(new_n118_), .dout(new_n119_));
  anb2 g0055(.dina(new_n106_), .dinb(new_n118_), .dout(new_n120_));
  anb2 g0056(.dina(new_n119_), .dinb(new_n120_), .dout(new_n121_));
  anb1 g0057(.dina(new_n105_), .dinb(new_n121_), .dout(new_n122_));
  anb2 g0058(.dina(new_n105_), .dinb(new_n121_), .dout(new_n123_));
  anb2 g0059(.dina(new_n122_), .dinb(new_n123_), .dout(new_n124_));
  anb1 g0060(.dina(new_n104_), .dinb(new_n124_), .dout(new_n125_));
  anb2 g0061(.dina(new_n104_), .dinb(new_n124_), .dout(new_n126_));
  anb2 g0062(.dina(new_n125_), .dinb(new_n126_), .dout(new_n127_));
  anb1 g0063(.dina(new_n103_), .dinb(new_n127_), .dout(new_n128_));
  anb2 g0064(.dina(new_n103_), .dinb(new_n127_), .dout(new_n129_));
  anb2 g0065(.dina(new_n128_), .dinb(new_n129_), .dout(G6261));
  nor2 g0066(.dina(G1), .dinb(G22), .dout(new_n131_));
  and2 g0067(.dina(new_n125_), .dinb(new_n128_), .dout(new_n132_));
  nor2 g0068(.dina(G2), .dinb(G21), .dout(new_n133_));
  and2 g0069(.dina(new_n119_), .dinb(new_n122_), .dout(new_n134_));
  nor2 g0070(.dina(G3), .dinb(G20), .dout(new_n135_));
  and2 g0071(.dina(new_n113_), .dinb(new_n116_), .dout(new_n136_));
  nor2 g0072(.dina(G4), .dinb(G19), .dout(new_n137_));
  nor2 g0073(.dina(G6), .dinb(G17), .dout(new_n138_));
  and1 g0074(.dina(G5), .dinb(G18), .dout(new_n139_));
  anb2 g0075(.dina(new_n138_), .dinb(new_n139_), .dout(new_n140_));
  anb1 g0076(.dina(new_n138_), .dinb(new_n139_), .dout(new_n141_));
  nab2 g0077(.dina(new_n140_), .dinb(new_n141_), .dout(new_n142_));
  anb2 g0078(.dina(new_n110_), .dinb(new_n142_), .dout(new_n143_));
  anb1 g0079(.dina(new_n110_), .dinb(new_n142_), .dout(new_n144_));
  nab2 g0080(.dina(new_n143_), .dinb(new_n144_), .dout(new_n145_));
  anb1 g0081(.dina(new_n137_), .dinb(new_n145_), .dout(new_n146_));
  anb2 g0082(.dina(new_n137_), .dinb(new_n145_), .dout(new_n147_));
  anb2 g0083(.dina(new_n146_), .dinb(new_n147_), .dout(new_n148_));
  anb1 g0084(.dina(new_n136_), .dinb(new_n148_), .dout(new_n149_));
  anb2 g0085(.dina(new_n136_), .dinb(new_n148_), .dout(new_n150_));
  anb2 g0086(.dina(new_n149_), .dinb(new_n150_), .dout(new_n151_));
  anb1 g0087(.dina(new_n135_), .dinb(new_n151_), .dout(new_n152_));
  anb2 g0088(.dina(new_n135_), .dinb(new_n151_), .dout(new_n153_));
  anb2 g0089(.dina(new_n152_), .dinb(new_n153_), .dout(new_n154_));
  anb1 g0090(.dina(new_n134_), .dinb(new_n154_), .dout(new_n155_));
  anb2 g0091(.dina(new_n134_), .dinb(new_n154_), .dout(new_n156_));
  anb2 g0092(.dina(new_n155_), .dinb(new_n156_), .dout(new_n157_));
  anb1 g0093(.dina(new_n133_), .dinb(new_n157_), .dout(new_n158_));
  anb2 g0094(.dina(new_n133_), .dinb(new_n157_), .dout(new_n159_));
  anb2 g0095(.dina(new_n158_), .dinb(new_n159_), .dout(new_n160_));
  anb1 g0096(.dina(new_n132_), .dinb(new_n160_), .dout(new_n161_));
  anb2 g0097(.dina(new_n132_), .dinb(new_n160_), .dout(new_n162_));
  anb2 g0098(.dina(new_n161_), .dinb(new_n162_), .dout(new_n163_));
  anb1 g0099(.dina(new_n131_), .dinb(new_n163_), .dout(new_n164_));
  anb2 g0100(.dina(new_n131_), .dinb(new_n163_), .dout(new_n165_));
  anb2 g0101(.dina(new_n164_), .dinb(new_n165_), .dout(G6262));
  nor2 g0102(.dina(G1), .dinb(G23), .dout(new_n167_));
  and2 g0103(.dina(new_n161_), .dinb(new_n164_), .dout(new_n168_));
  nor2 g0104(.dina(G2), .dinb(G22), .dout(new_n169_));
  and2 g0105(.dina(new_n155_), .dinb(new_n158_), .dout(new_n170_));
  nor2 g0106(.dina(G3), .dinb(G21), .dout(new_n171_));
  and2 g0107(.dina(new_n149_), .dinb(new_n152_), .dout(new_n172_));
  nor2 g0108(.dina(G4), .dinb(G20), .dout(new_n173_));
  anb1 g0109(.dina(new_n143_), .dinb(new_n146_), .dout(new_n174_));
  and1 g0110(.dina(G5), .dinb(G19), .dout(new_n175_));
  nor2 g0111(.dina(G7), .dinb(G17), .dout(new_n176_));
  and1 g0112(.dina(G6), .dinb(G18), .dout(new_n177_));
  anb2 g0113(.dina(new_n176_), .dinb(new_n177_), .dout(new_n178_));
  anb1 g0114(.dina(new_n176_), .dinb(new_n177_), .dout(new_n179_));
  anb1 g0115(.dina(new_n178_), .dinb(new_n179_), .dout(new_n180_));
  anb1 g0116(.dina(new_n140_), .dinb(new_n180_), .dout(new_n181_));
  anb2 g0117(.dina(new_n140_), .dinb(new_n180_), .dout(new_n182_));
  nab1 g0118(.dina(new_n181_), .dinb(new_n182_), .dout(new_n183_));
  anb2 g0119(.dina(new_n175_), .dinb(new_n183_), .dout(new_n184_));
  anb1 g0120(.dina(new_n175_), .dinb(new_n183_), .dout(new_n185_));
  anb1 g0121(.dina(new_n184_), .dinb(new_n185_), .dout(new_n186_));
  anb2 g0122(.dina(new_n174_), .dinb(new_n186_), .dout(new_n187_));
  anb1 g0123(.dina(new_n174_), .dinb(new_n186_), .dout(new_n188_));
  nab2 g0124(.dina(new_n187_), .dinb(new_n188_), .dout(new_n189_));
  anb1 g0125(.dina(new_n173_), .dinb(new_n189_), .dout(new_n190_));
  anb2 g0126(.dina(new_n173_), .dinb(new_n189_), .dout(new_n191_));
  anb2 g0127(.dina(new_n190_), .dinb(new_n191_), .dout(new_n192_));
  anb1 g0128(.dina(new_n172_), .dinb(new_n192_), .dout(new_n193_));
  anb2 g0129(.dina(new_n172_), .dinb(new_n192_), .dout(new_n194_));
  anb2 g0130(.dina(new_n193_), .dinb(new_n194_), .dout(new_n195_));
  anb1 g0131(.dina(new_n171_), .dinb(new_n195_), .dout(new_n196_));
  anb2 g0132(.dina(new_n171_), .dinb(new_n195_), .dout(new_n197_));
  anb2 g0133(.dina(new_n196_), .dinb(new_n197_), .dout(new_n198_));
  anb1 g0134(.dina(new_n170_), .dinb(new_n198_), .dout(new_n199_));
  anb2 g0135(.dina(new_n170_), .dinb(new_n198_), .dout(new_n200_));
  anb2 g0136(.dina(new_n199_), .dinb(new_n200_), .dout(new_n201_));
  anb1 g0137(.dina(new_n169_), .dinb(new_n201_), .dout(new_n202_));
  anb2 g0138(.dina(new_n169_), .dinb(new_n201_), .dout(new_n203_));
  anb2 g0139(.dina(new_n202_), .dinb(new_n203_), .dout(new_n204_));
  anb1 g0140(.dina(new_n168_), .dinb(new_n204_), .dout(new_n205_));
  anb2 g0141(.dina(new_n168_), .dinb(new_n204_), .dout(new_n206_));
  anb2 g0142(.dina(new_n205_), .dinb(new_n206_), .dout(new_n207_));
  anb1 g0143(.dina(new_n167_), .dinb(new_n207_), .dout(new_n208_));
  anb2 g0144(.dina(new_n167_), .dinb(new_n207_), .dout(new_n209_));
  anb2 g0145(.dina(new_n208_), .dinb(new_n209_), .dout(G6263));
  nor2 g0146(.dina(G1), .dinb(G24), .dout(new_n211_));
  and2 g0147(.dina(new_n205_), .dinb(new_n208_), .dout(new_n212_));
  nor2 g0148(.dina(G2), .dinb(G23), .dout(new_n213_));
  and2 g0149(.dina(new_n199_), .dinb(new_n202_), .dout(new_n214_));
  nor2 g0150(.dina(G3), .dinb(G22), .dout(new_n215_));
  and2 g0151(.dina(new_n193_), .dinb(new_n196_), .dout(new_n216_));
  nor2 g0152(.dina(G4), .dinb(G21), .dout(new_n217_));
  anb1 g0153(.dina(new_n187_), .dinb(new_n190_), .dout(new_n218_));
  and1 g0154(.dina(G5), .dinb(G20), .dout(new_n219_));
  anb2 g0155(.dina(new_n181_), .dinb(new_n184_), .dout(new_n220_));
  and1 g0156(.dina(G6), .dinb(G19), .dout(new_n221_));
  nor2 g0157(.dina(G8), .dinb(G17), .dout(new_n222_));
  and1 g0158(.dina(G7), .dinb(G18), .dout(new_n223_));
  anb2 g0159(.dina(new_n222_), .dinb(new_n223_), .dout(new_n224_));
  anb1 g0160(.dina(new_n222_), .dinb(new_n223_), .dout(new_n225_));
  anb1 g0161(.dina(new_n224_), .dinb(new_n225_), .dout(new_n226_));
  anb1 g0162(.dina(new_n178_), .dinb(new_n226_), .dout(new_n227_));
  anb2 g0163(.dina(new_n178_), .dinb(new_n226_), .dout(new_n228_));
  nab1 g0164(.dina(new_n227_), .dinb(new_n228_), .dout(new_n229_));
  anb2 g0165(.dina(new_n221_), .dinb(new_n229_), .dout(new_n230_));
  anb1 g0166(.dina(new_n221_), .dinb(new_n229_), .dout(new_n231_));
  nab2 g0167(.dina(new_n230_), .dinb(new_n231_), .dout(new_n232_));
  anb1 g0168(.dina(new_n220_), .dinb(new_n232_), .dout(new_n233_));
  anb2 g0169(.dina(new_n220_), .dinb(new_n232_), .dout(new_n234_));
  nab1 g0170(.dina(new_n233_), .dinb(new_n234_), .dout(new_n235_));
  anb2 g0171(.dina(new_n219_), .dinb(new_n235_), .dout(new_n236_));
  anb1 g0172(.dina(new_n219_), .dinb(new_n235_), .dout(new_n237_));
  anb1 g0173(.dina(new_n236_), .dinb(new_n237_), .dout(new_n238_));
  anb2 g0174(.dina(new_n218_), .dinb(new_n238_), .dout(new_n239_));
  anb1 g0175(.dina(new_n218_), .dinb(new_n238_), .dout(new_n240_));
  nab2 g0176(.dina(new_n239_), .dinb(new_n240_), .dout(new_n241_));
  anb1 g0177(.dina(new_n217_), .dinb(new_n241_), .dout(new_n242_));
  anb2 g0178(.dina(new_n217_), .dinb(new_n241_), .dout(new_n243_));
  anb2 g0179(.dina(new_n242_), .dinb(new_n243_), .dout(new_n244_));
  anb1 g0180(.dina(new_n216_), .dinb(new_n244_), .dout(new_n245_));
  anb2 g0181(.dina(new_n216_), .dinb(new_n244_), .dout(new_n246_));
  anb2 g0182(.dina(new_n245_), .dinb(new_n246_), .dout(new_n247_));
  anb1 g0183(.dina(new_n215_), .dinb(new_n247_), .dout(new_n248_));
  anb2 g0184(.dina(new_n215_), .dinb(new_n247_), .dout(new_n249_));
  anb2 g0185(.dina(new_n248_), .dinb(new_n249_), .dout(new_n250_));
  anb1 g0186(.dina(new_n214_), .dinb(new_n250_), .dout(new_n251_));
  anb2 g0187(.dina(new_n214_), .dinb(new_n250_), .dout(new_n252_));
  anb2 g0188(.dina(new_n251_), .dinb(new_n252_), .dout(new_n253_));
  anb1 g0189(.dina(new_n213_), .dinb(new_n253_), .dout(new_n254_));
  anb2 g0190(.dina(new_n213_), .dinb(new_n253_), .dout(new_n255_));
  anb2 g0191(.dina(new_n254_), .dinb(new_n255_), .dout(new_n256_));
  anb1 g0192(.dina(new_n212_), .dinb(new_n256_), .dout(new_n257_));
  anb2 g0193(.dina(new_n212_), .dinb(new_n256_), .dout(new_n258_));
  anb2 g0194(.dina(new_n257_), .dinb(new_n258_), .dout(new_n259_));
  anb1 g0195(.dina(new_n211_), .dinb(new_n259_), .dout(new_n260_));
  anb2 g0196(.dina(new_n211_), .dinb(new_n259_), .dout(new_n261_));
  anb2 g0197(.dina(new_n260_), .dinb(new_n261_), .dout(G6264));
  nor2 g0198(.dina(G1), .dinb(G25), .dout(new_n263_));
  and2 g0199(.dina(new_n257_), .dinb(new_n260_), .dout(new_n264_));
  nor2 g0200(.dina(G2), .dinb(G24), .dout(new_n265_));
  and2 g0201(.dina(new_n251_), .dinb(new_n254_), .dout(new_n266_));
  nor2 g0202(.dina(G3), .dinb(G23), .dout(new_n267_));
  and2 g0203(.dina(new_n245_), .dinb(new_n248_), .dout(new_n268_));
  nor2 g0204(.dina(G4), .dinb(G22), .dout(new_n269_));
  anb1 g0205(.dina(new_n239_), .dinb(new_n242_), .dout(new_n270_));
  and1 g0206(.dina(G5), .dinb(G21), .dout(new_n271_));
  anb2 g0207(.dina(new_n233_), .dinb(new_n236_), .dout(new_n272_));
  and1 g0208(.dina(G6), .dinb(G20), .dout(new_n273_));
  anb2 g0209(.dina(new_n227_), .dinb(new_n230_), .dout(new_n274_));
  and1 g0210(.dina(G7), .dinb(G19), .dout(new_n275_));
  nor2 g0211(.dina(G9), .dinb(G17), .dout(new_n276_));
  and1 g0212(.dina(G8), .dinb(G18), .dout(new_n277_));
  anb2 g0213(.dina(new_n276_), .dinb(new_n277_), .dout(new_n278_));
  anb1 g0214(.dina(new_n276_), .dinb(new_n277_), .dout(new_n279_));
  anb1 g0215(.dina(new_n278_), .dinb(new_n279_), .dout(new_n280_));
  anb1 g0216(.dina(new_n224_), .dinb(new_n280_), .dout(new_n281_));
  anb2 g0217(.dina(new_n224_), .dinb(new_n280_), .dout(new_n282_));
  nab1 g0218(.dina(new_n281_), .dinb(new_n282_), .dout(new_n283_));
  anb2 g0219(.dina(new_n275_), .dinb(new_n283_), .dout(new_n284_));
  anb1 g0220(.dina(new_n275_), .dinb(new_n283_), .dout(new_n285_));
  nab2 g0221(.dina(new_n284_), .dinb(new_n285_), .dout(new_n286_));
  anb1 g0222(.dina(new_n274_), .dinb(new_n286_), .dout(new_n287_));
  anb2 g0223(.dina(new_n274_), .dinb(new_n286_), .dout(new_n288_));
  nab1 g0224(.dina(new_n287_), .dinb(new_n288_), .dout(new_n289_));
  anb2 g0225(.dina(new_n273_), .dinb(new_n289_), .dout(new_n290_));
  anb1 g0226(.dina(new_n273_), .dinb(new_n289_), .dout(new_n291_));
  nab2 g0227(.dina(new_n290_), .dinb(new_n291_), .dout(new_n292_));
  anb1 g0228(.dina(new_n272_), .dinb(new_n292_), .dout(new_n293_));
  anb2 g0229(.dina(new_n272_), .dinb(new_n292_), .dout(new_n294_));
  nab1 g0230(.dina(new_n293_), .dinb(new_n294_), .dout(new_n295_));
  anb2 g0231(.dina(new_n271_), .dinb(new_n295_), .dout(new_n296_));
  anb1 g0232(.dina(new_n271_), .dinb(new_n295_), .dout(new_n297_));
  anb1 g0233(.dina(new_n296_), .dinb(new_n297_), .dout(new_n298_));
  anb2 g0234(.dina(new_n270_), .dinb(new_n298_), .dout(new_n299_));
  anb1 g0235(.dina(new_n270_), .dinb(new_n298_), .dout(new_n300_));
  nab2 g0236(.dina(new_n299_), .dinb(new_n300_), .dout(new_n301_));
  anb1 g0237(.dina(new_n269_), .dinb(new_n301_), .dout(new_n302_));
  anb2 g0238(.dina(new_n269_), .dinb(new_n301_), .dout(new_n303_));
  anb2 g0239(.dina(new_n302_), .dinb(new_n303_), .dout(new_n304_));
  anb1 g0240(.dina(new_n268_), .dinb(new_n304_), .dout(new_n305_));
  anb2 g0241(.dina(new_n268_), .dinb(new_n304_), .dout(new_n306_));
  anb2 g0242(.dina(new_n305_), .dinb(new_n306_), .dout(new_n307_));
  anb1 g0243(.dina(new_n267_), .dinb(new_n307_), .dout(new_n308_));
  anb2 g0244(.dina(new_n267_), .dinb(new_n307_), .dout(new_n309_));
  anb2 g0245(.dina(new_n308_), .dinb(new_n309_), .dout(new_n310_));
  anb1 g0246(.dina(new_n266_), .dinb(new_n310_), .dout(new_n311_));
  anb2 g0247(.dina(new_n266_), .dinb(new_n310_), .dout(new_n312_));
  anb2 g0248(.dina(new_n311_), .dinb(new_n312_), .dout(new_n313_));
  anb1 g0249(.dina(new_n265_), .dinb(new_n313_), .dout(new_n314_));
  anb2 g0250(.dina(new_n265_), .dinb(new_n313_), .dout(new_n315_));
  anb2 g0251(.dina(new_n314_), .dinb(new_n315_), .dout(new_n316_));
  anb1 g0252(.dina(new_n264_), .dinb(new_n316_), .dout(new_n317_));
  anb2 g0253(.dina(new_n264_), .dinb(new_n316_), .dout(new_n318_));
  anb2 g0254(.dina(new_n317_), .dinb(new_n318_), .dout(new_n319_));
  anb1 g0255(.dina(new_n263_), .dinb(new_n319_), .dout(new_n320_));
  anb2 g0256(.dina(new_n263_), .dinb(new_n319_), .dout(new_n321_));
  anb2 g0257(.dina(new_n320_), .dinb(new_n321_), .dout(G6265));
  nor2 g0258(.dina(G1), .dinb(G26), .dout(new_n323_));
  and2 g0259(.dina(new_n317_), .dinb(new_n320_), .dout(new_n324_));
  nor2 g0260(.dina(G2), .dinb(G25), .dout(new_n325_));
  and2 g0261(.dina(new_n311_), .dinb(new_n314_), .dout(new_n326_));
  nor2 g0262(.dina(G3), .dinb(G24), .dout(new_n327_));
  and2 g0263(.dina(new_n305_), .dinb(new_n308_), .dout(new_n328_));
  nor2 g0264(.dina(G4), .dinb(G23), .dout(new_n329_));
  anb1 g0265(.dina(new_n299_), .dinb(new_n302_), .dout(new_n330_));
  and1 g0266(.dina(G5), .dinb(G22), .dout(new_n331_));
  anb2 g0267(.dina(new_n293_), .dinb(new_n296_), .dout(new_n332_));
  and1 g0268(.dina(G6), .dinb(G21), .dout(new_n333_));
  anb2 g0269(.dina(new_n287_), .dinb(new_n290_), .dout(new_n334_));
  and1 g0270(.dina(G7), .dinb(G20), .dout(new_n335_));
  anb2 g0271(.dina(new_n281_), .dinb(new_n284_), .dout(new_n336_));
  and1 g0272(.dina(G8), .dinb(G19), .dout(new_n337_));
  nor2 g0273(.dina(G10), .dinb(G17), .dout(new_n338_));
  and1 g0274(.dina(G9), .dinb(G18), .dout(new_n339_));
  anb2 g0275(.dina(new_n338_), .dinb(new_n339_), .dout(new_n340_));
  anb1 g0276(.dina(new_n338_), .dinb(new_n339_), .dout(new_n341_));
  anb1 g0277(.dina(new_n340_), .dinb(new_n341_), .dout(new_n342_));
  anb1 g0278(.dina(new_n278_), .dinb(new_n342_), .dout(new_n343_));
  anb2 g0279(.dina(new_n278_), .dinb(new_n342_), .dout(new_n344_));
  nab1 g0280(.dina(new_n343_), .dinb(new_n344_), .dout(new_n345_));
  anb2 g0281(.dina(new_n337_), .dinb(new_n345_), .dout(new_n346_));
  anb1 g0282(.dina(new_n337_), .dinb(new_n345_), .dout(new_n347_));
  nab2 g0283(.dina(new_n346_), .dinb(new_n347_), .dout(new_n348_));
  anb1 g0284(.dina(new_n336_), .dinb(new_n348_), .dout(new_n349_));
  anb2 g0285(.dina(new_n336_), .dinb(new_n348_), .dout(new_n350_));
  nab1 g0286(.dina(new_n349_), .dinb(new_n350_), .dout(new_n351_));
  anb2 g0287(.dina(new_n335_), .dinb(new_n351_), .dout(new_n352_));
  anb1 g0288(.dina(new_n335_), .dinb(new_n351_), .dout(new_n353_));
  nab2 g0289(.dina(new_n352_), .dinb(new_n353_), .dout(new_n354_));
  anb1 g0290(.dina(new_n334_), .dinb(new_n354_), .dout(new_n355_));
  anb2 g0291(.dina(new_n334_), .dinb(new_n354_), .dout(new_n356_));
  nab1 g0292(.dina(new_n355_), .dinb(new_n356_), .dout(new_n357_));
  anb2 g0293(.dina(new_n333_), .dinb(new_n357_), .dout(new_n358_));
  anb1 g0294(.dina(new_n333_), .dinb(new_n357_), .dout(new_n359_));
  nab2 g0295(.dina(new_n358_), .dinb(new_n359_), .dout(new_n360_));
  anb1 g0296(.dina(new_n332_), .dinb(new_n360_), .dout(new_n361_));
  anb2 g0297(.dina(new_n332_), .dinb(new_n360_), .dout(new_n362_));
  nab1 g0298(.dina(new_n361_), .dinb(new_n362_), .dout(new_n363_));
  anb2 g0299(.dina(new_n331_), .dinb(new_n363_), .dout(new_n364_));
  anb1 g0300(.dina(new_n331_), .dinb(new_n363_), .dout(new_n365_));
  anb1 g0301(.dina(new_n364_), .dinb(new_n365_), .dout(new_n366_));
  anb2 g0302(.dina(new_n330_), .dinb(new_n366_), .dout(new_n367_));
  anb1 g0303(.dina(new_n330_), .dinb(new_n366_), .dout(new_n368_));
  nab2 g0304(.dina(new_n367_), .dinb(new_n368_), .dout(new_n369_));
  anb1 g0305(.dina(new_n329_), .dinb(new_n369_), .dout(new_n370_));
  anb2 g0306(.dina(new_n329_), .dinb(new_n369_), .dout(new_n371_));
  anb2 g0307(.dina(new_n370_), .dinb(new_n371_), .dout(new_n372_));
  anb1 g0308(.dina(new_n328_), .dinb(new_n372_), .dout(new_n373_));
  anb2 g0309(.dina(new_n328_), .dinb(new_n372_), .dout(new_n374_));
  anb2 g0310(.dina(new_n373_), .dinb(new_n374_), .dout(new_n375_));
  anb1 g0311(.dina(new_n327_), .dinb(new_n375_), .dout(new_n376_));
  anb2 g0312(.dina(new_n327_), .dinb(new_n375_), .dout(new_n377_));
  anb2 g0313(.dina(new_n376_), .dinb(new_n377_), .dout(new_n378_));
  anb1 g0314(.dina(new_n326_), .dinb(new_n378_), .dout(new_n379_));
  anb2 g0315(.dina(new_n326_), .dinb(new_n378_), .dout(new_n380_));
  anb2 g0316(.dina(new_n379_), .dinb(new_n380_), .dout(new_n381_));
  anb1 g0317(.dina(new_n325_), .dinb(new_n381_), .dout(new_n382_));
  anb2 g0318(.dina(new_n325_), .dinb(new_n381_), .dout(new_n383_));
  anb2 g0319(.dina(new_n382_), .dinb(new_n383_), .dout(new_n384_));
  anb1 g0320(.dina(new_n324_), .dinb(new_n384_), .dout(new_n385_));
  anb2 g0321(.dina(new_n324_), .dinb(new_n384_), .dout(new_n386_));
  anb2 g0322(.dina(new_n385_), .dinb(new_n386_), .dout(new_n387_));
  anb1 g0323(.dina(new_n323_), .dinb(new_n387_), .dout(new_n388_));
  anb2 g0324(.dina(new_n323_), .dinb(new_n387_), .dout(new_n389_));
  anb2 g0325(.dina(new_n388_), .dinb(new_n389_), .dout(G6266));
  nor2 g0326(.dina(G1), .dinb(G27), .dout(new_n391_));
  and2 g0327(.dina(new_n385_), .dinb(new_n388_), .dout(new_n392_));
  nor2 g0328(.dina(G2), .dinb(G26), .dout(new_n393_));
  and2 g0329(.dina(new_n379_), .dinb(new_n382_), .dout(new_n394_));
  nor2 g0330(.dina(G3), .dinb(G25), .dout(new_n395_));
  and2 g0331(.dina(new_n373_), .dinb(new_n376_), .dout(new_n396_));
  nor2 g0332(.dina(G4), .dinb(G24), .dout(new_n397_));
  anb1 g0333(.dina(new_n367_), .dinb(new_n370_), .dout(new_n398_));
  and1 g0334(.dina(G5), .dinb(G23), .dout(new_n399_));
  anb2 g0335(.dina(new_n361_), .dinb(new_n364_), .dout(new_n400_));
  and1 g0336(.dina(G6), .dinb(G22), .dout(new_n401_));
  anb2 g0337(.dina(new_n355_), .dinb(new_n358_), .dout(new_n402_));
  and1 g0338(.dina(G7), .dinb(G21), .dout(new_n403_));
  anb2 g0339(.dina(new_n349_), .dinb(new_n352_), .dout(new_n404_));
  and1 g0340(.dina(G8), .dinb(G20), .dout(new_n405_));
  anb2 g0341(.dina(new_n343_), .dinb(new_n346_), .dout(new_n406_));
  and1 g0342(.dina(G9), .dinb(G19), .dout(new_n407_));
  nor2 g0343(.dina(G11), .dinb(G17), .dout(new_n408_));
  and1 g0344(.dina(G10), .dinb(G18), .dout(new_n409_));
  anb2 g0345(.dina(new_n408_), .dinb(new_n409_), .dout(new_n410_));
  anb1 g0346(.dina(new_n408_), .dinb(new_n409_), .dout(new_n411_));
  anb1 g0347(.dina(new_n410_), .dinb(new_n411_), .dout(new_n412_));
  anb1 g0348(.dina(new_n340_), .dinb(new_n412_), .dout(new_n413_));
  anb2 g0349(.dina(new_n340_), .dinb(new_n412_), .dout(new_n414_));
  nab1 g0350(.dina(new_n413_), .dinb(new_n414_), .dout(new_n415_));
  anb2 g0351(.dina(new_n407_), .dinb(new_n415_), .dout(new_n416_));
  anb1 g0352(.dina(new_n407_), .dinb(new_n415_), .dout(new_n417_));
  nab2 g0353(.dina(new_n416_), .dinb(new_n417_), .dout(new_n418_));
  anb1 g0354(.dina(new_n406_), .dinb(new_n418_), .dout(new_n419_));
  anb2 g0355(.dina(new_n406_), .dinb(new_n418_), .dout(new_n420_));
  nab1 g0356(.dina(new_n419_), .dinb(new_n420_), .dout(new_n421_));
  anb2 g0357(.dina(new_n405_), .dinb(new_n421_), .dout(new_n422_));
  anb1 g0358(.dina(new_n405_), .dinb(new_n421_), .dout(new_n423_));
  nab2 g0359(.dina(new_n422_), .dinb(new_n423_), .dout(new_n424_));
  anb1 g0360(.dina(new_n404_), .dinb(new_n424_), .dout(new_n425_));
  anb2 g0361(.dina(new_n404_), .dinb(new_n424_), .dout(new_n426_));
  nab1 g0362(.dina(new_n425_), .dinb(new_n426_), .dout(new_n427_));
  anb2 g0363(.dina(new_n403_), .dinb(new_n427_), .dout(new_n428_));
  anb1 g0364(.dina(new_n403_), .dinb(new_n427_), .dout(new_n429_));
  nab2 g0365(.dina(new_n428_), .dinb(new_n429_), .dout(new_n430_));
  anb1 g0366(.dina(new_n402_), .dinb(new_n430_), .dout(new_n431_));
  anb2 g0367(.dina(new_n402_), .dinb(new_n430_), .dout(new_n432_));
  nab1 g0368(.dina(new_n431_), .dinb(new_n432_), .dout(new_n433_));
  anb2 g0369(.dina(new_n401_), .dinb(new_n433_), .dout(new_n434_));
  anb1 g0370(.dina(new_n401_), .dinb(new_n433_), .dout(new_n435_));
  nab2 g0371(.dina(new_n434_), .dinb(new_n435_), .dout(new_n436_));
  anb1 g0372(.dina(new_n400_), .dinb(new_n436_), .dout(new_n437_));
  anb2 g0373(.dina(new_n400_), .dinb(new_n436_), .dout(new_n438_));
  nab1 g0374(.dina(new_n437_), .dinb(new_n438_), .dout(new_n439_));
  anb2 g0375(.dina(new_n399_), .dinb(new_n439_), .dout(new_n440_));
  anb1 g0376(.dina(new_n399_), .dinb(new_n439_), .dout(new_n441_));
  anb1 g0377(.dina(new_n440_), .dinb(new_n441_), .dout(new_n442_));
  anb2 g0378(.dina(new_n398_), .dinb(new_n442_), .dout(new_n443_));
  anb1 g0379(.dina(new_n398_), .dinb(new_n442_), .dout(new_n444_));
  nab2 g0380(.dina(new_n443_), .dinb(new_n444_), .dout(new_n445_));
  anb1 g0381(.dina(new_n397_), .dinb(new_n445_), .dout(new_n446_));
  anb2 g0382(.dina(new_n397_), .dinb(new_n445_), .dout(new_n447_));
  anb2 g0383(.dina(new_n446_), .dinb(new_n447_), .dout(new_n448_));
  anb1 g0384(.dina(new_n396_), .dinb(new_n448_), .dout(new_n449_));
  anb2 g0385(.dina(new_n396_), .dinb(new_n448_), .dout(new_n450_));
  anb2 g0386(.dina(new_n449_), .dinb(new_n450_), .dout(new_n451_));
  anb1 g0387(.dina(new_n395_), .dinb(new_n451_), .dout(new_n452_));
  anb2 g0388(.dina(new_n395_), .dinb(new_n451_), .dout(new_n453_));
  anb2 g0389(.dina(new_n452_), .dinb(new_n453_), .dout(new_n454_));
  anb1 g0390(.dina(new_n394_), .dinb(new_n454_), .dout(new_n455_));
  anb2 g0391(.dina(new_n394_), .dinb(new_n454_), .dout(new_n456_));
  anb2 g0392(.dina(new_n455_), .dinb(new_n456_), .dout(new_n457_));
  anb1 g0393(.dina(new_n393_), .dinb(new_n457_), .dout(new_n458_));
  anb2 g0394(.dina(new_n393_), .dinb(new_n457_), .dout(new_n459_));
  anb2 g0395(.dina(new_n458_), .dinb(new_n459_), .dout(new_n460_));
  anb1 g0396(.dina(new_n392_), .dinb(new_n460_), .dout(new_n461_));
  anb2 g0397(.dina(new_n392_), .dinb(new_n460_), .dout(new_n462_));
  anb2 g0398(.dina(new_n461_), .dinb(new_n462_), .dout(new_n463_));
  anb1 g0399(.dina(new_n391_), .dinb(new_n463_), .dout(new_n464_));
  anb2 g0400(.dina(new_n391_), .dinb(new_n463_), .dout(new_n465_));
  anb2 g0401(.dina(new_n464_), .dinb(new_n465_), .dout(G6267));
  nor2 g0402(.dina(G1), .dinb(G28), .dout(new_n467_));
  and2 g0403(.dina(new_n461_), .dinb(new_n464_), .dout(new_n468_));
  nor2 g0404(.dina(G2), .dinb(G27), .dout(new_n469_));
  and2 g0405(.dina(new_n455_), .dinb(new_n458_), .dout(new_n470_));
  nor2 g0406(.dina(G3), .dinb(G26), .dout(new_n471_));
  and2 g0407(.dina(new_n449_), .dinb(new_n452_), .dout(new_n472_));
  nor2 g0408(.dina(G4), .dinb(G25), .dout(new_n473_));
  anb1 g0409(.dina(new_n443_), .dinb(new_n446_), .dout(new_n474_));
  and1 g0410(.dina(G5), .dinb(G24), .dout(new_n475_));
  anb2 g0411(.dina(new_n437_), .dinb(new_n440_), .dout(new_n476_));
  and1 g0412(.dina(G6), .dinb(G23), .dout(new_n477_));
  anb2 g0413(.dina(new_n431_), .dinb(new_n434_), .dout(new_n478_));
  and1 g0414(.dina(G7), .dinb(G22), .dout(new_n479_));
  anb2 g0415(.dina(new_n425_), .dinb(new_n428_), .dout(new_n480_));
  and1 g0416(.dina(G8), .dinb(G21), .dout(new_n481_));
  anb2 g0417(.dina(new_n419_), .dinb(new_n422_), .dout(new_n482_));
  and1 g0418(.dina(G9), .dinb(G20), .dout(new_n483_));
  anb2 g0419(.dina(new_n413_), .dinb(new_n416_), .dout(new_n484_));
  and1 g0420(.dina(G10), .dinb(G19), .dout(new_n485_));
  nor2 g0421(.dina(G12), .dinb(G17), .dout(new_n486_));
  and1 g0422(.dina(G11), .dinb(G18), .dout(new_n487_));
  anb2 g0423(.dina(new_n486_), .dinb(new_n487_), .dout(new_n488_));
  anb1 g0424(.dina(new_n486_), .dinb(new_n487_), .dout(new_n489_));
  anb1 g0425(.dina(new_n488_), .dinb(new_n489_), .dout(new_n490_));
  anb1 g0426(.dina(new_n410_), .dinb(new_n490_), .dout(new_n491_));
  anb2 g0427(.dina(new_n410_), .dinb(new_n490_), .dout(new_n492_));
  nab1 g0428(.dina(new_n491_), .dinb(new_n492_), .dout(new_n493_));
  anb2 g0429(.dina(new_n485_), .dinb(new_n493_), .dout(new_n494_));
  anb1 g0430(.dina(new_n485_), .dinb(new_n493_), .dout(new_n495_));
  nab2 g0431(.dina(new_n494_), .dinb(new_n495_), .dout(new_n496_));
  anb1 g0432(.dina(new_n484_), .dinb(new_n496_), .dout(new_n497_));
  anb2 g0433(.dina(new_n484_), .dinb(new_n496_), .dout(new_n498_));
  nab1 g0434(.dina(new_n497_), .dinb(new_n498_), .dout(new_n499_));
  anb2 g0435(.dina(new_n483_), .dinb(new_n499_), .dout(new_n500_));
  anb1 g0436(.dina(new_n483_), .dinb(new_n499_), .dout(new_n501_));
  nab2 g0437(.dina(new_n500_), .dinb(new_n501_), .dout(new_n502_));
  anb1 g0438(.dina(new_n482_), .dinb(new_n502_), .dout(new_n503_));
  anb2 g0439(.dina(new_n482_), .dinb(new_n502_), .dout(new_n504_));
  nab1 g0440(.dina(new_n503_), .dinb(new_n504_), .dout(new_n505_));
  anb2 g0441(.dina(new_n481_), .dinb(new_n505_), .dout(new_n506_));
  anb1 g0442(.dina(new_n481_), .dinb(new_n505_), .dout(new_n507_));
  nab2 g0443(.dina(new_n506_), .dinb(new_n507_), .dout(new_n508_));
  anb1 g0444(.dina(new_n480_), .dinb(new_n508_), .dout(new_n509_));
  anb2 g0445(.dina(new_n480_), .dinb(new_n508_), .dout(new_n510_));
  nab1 g0446(.dina(new_n509_), .dinb(new_n510_), .dout(new_n511_));
  anb2 g0447(.dina(new_n479_), .dinb(new_n511_), .dout(new_n512_));
  anb1 g0448(.dina(new_n479_), .dinb(new_n511_), .dout(new_n513_));
  nab2 g0449(.dina(new_n512_), .dinb(new_n513_), .dout(new_n514_));
  anb1 g0450(.dina(new_n478_), .dinb(new_n514_), .dout(new_n515_));
  anb2 g0451(.dina(new_n478_), .dinb(new_n514_), .dout(new_n516_));
  nab1 g0452(.dina(new_n515_), .dinb(new_n516_), .dout(new_n517_));
  anb2 g0453(.dina(new_n477_), .dinb(new_n517_), .dout(new_n518_));
  anb1 g0454(.dina(new_n477_), .dinb(new_n517_), .dout(new_n519_));
  nab2 g0455(.dina(new_n518_), .dinb(new_n519_), .dout(new_n520_));
  anb1 g0456(.dina(new_n476_), .dinb(new_n520_), .dout(new_n521_));
  anb2 g0457(.dina(new_n476_), .dinb(new_n520_), .dout(new_n522_));
  nab1 g0458(.dina(new_n521_), .dinb(new_n522_), .dout(new_n523_));
  anb2 g0459(.dina(new_n475_), .dinb(new_n523_), .dout(new_n524_));
  anb1 g0460(.dina(new_n475_), .dinb(new_n523_), .dout(new_n525_));
  anb1 g0461(.dina(new_n524_), .dinb(new_n525_), .dout(new_n526_));
  anb2 g0462(.dina(new_n474_), .dinb(new_n526_), .dout(new_n527_));
  anb1 g0463(.dina(new_n474_), .dinb(new_n526_), .dout(new_n528_));
  nab2 g0464(.dina(new_n527_), .dinb(new_n528_), .dout(new_n529_));
  anb1 g0465(.dina(new_n473_), .dinb(new_n529_), .dout(new_n530_));
  anb2 g0466(.dina(new_n473_), .dinb(new_n529_), .dout(new_n531_));
  anb2 g0467(.dina(new_n530_), .dinb(new_n531_), .dout(new_n532_));
  anb1 g0468(.dina(new_n472_), .dinb(new_n532_), .dout(new_n533_));
  anb2 g0469(.dina(new_n472_), .dinb(new_n532_), .dout(new_n534_));
  anb2 g0470(.dina(new_n533_), .dinb(new_n534_), .dout(new_n535_));
  anb1 g0471(.dina(new_n471_), .dinb(new_n535_), .dout(new_n536_));
  anb2 g0472(.dina(new_n471_), .dinb(new_n535_), .dout(new_n537_));
  anb2 g0473(.dina(new_n536_), .dinb(new_n537_), .dout(new_n538_));
  anb1 g0474(.dina(new_n470_), .dinb(new_n538_), .dout(new_n539_));
  anb2 g0475(.dina(new_n470_), .dinb(new_n538_), .dout(new_n540_));
  anb2 g0476(.dina(new_n539_), .dinb(new_n540_), .dout(new_n541_));
  anb1 g0477(.dina(new_n469_), .dinb(new_n541_), .dout(new_n542_));
  anb2 g0478(.dina(new_n469_), .dinb(new_n541_), .dout(new_n543_));
  anb2 g0479(.dina(new_n542_), .dinb(new_n543_), .dout(new_n544_));
  anb1 g0480(.dina(new_n468_), .dinb(new_n544_), .dout(new_n545_));
  anb2 g0481(.dina(new_n468_), .dinb(new_n544_), .dout(new_n546_));
  anb2 g0482(.dina(new_n545_), .dinb(new_n546_), .dout(new_n547_));
  anb1 g0483(.dina(new_n467_), .dinb(new_n547_), .dout(new_n548_));
  anb2 g0484(.dina(new_n467_), .dinb(new_n547_), .dout(new_n549_));
  anb2 g0485(.dina(new_n548_), .dinb(new_n549_), .dout(G6268));
  nor2 g0486(.dina(G1), .dinb(G29), .dout(new_n551_));
  and2 g0487(.dina(new_n545_), .dinb(new_n548_), .dout(new_n552_));
  nor2 g0488(.dina(G2), .dinb(G28), .dout(new_n553_));
  and2 g0489(.dina(new_n539_), .dinb(new_n542_), .dout(new_n554_));
  nor2 g0490(.dina(G3), .dinb(G27), .dout(new_n555_));
  and2 g0491(.dina(new_n533_), .dinb(new_n536_), .dout(new_n556_));
  nor2 g0492(.dina(G4), .dinb(G26), .dout(new_n557_));
  anb1 g0493(.dina(new_n527_), .dinb(new_n530_), .dout(new_n558_));
  and1 g0494(.dina(G5), .dinb(G25), .dout(new_n559_));
  anb2 g0495(.dina(new_n521_), .dinb(new_n524_), .dout(new_n560_));
  and1 g0496(.dina(G6), .dinb(G24), .dout(new_n561_));
  anb2 g0497(.dina(new_n515_), .dinb(new_n518_), .dout(new_n562_));
  and1 g0498(.dina(G7), .dinb(G23), .dout(new_n563_));
  anb2 g0499(.dina(new_n509_), .dinb(new_n512_), .dout(new_n564_));
  and1 g0500(.dina(G8), .dinb(G22), .dout(new_n565_));
  anb2 g0501(.dina(new_n503_), .dinb(new_n506_), .dout(new_n566_));
  and1 g0502(.dina(G9), .dinb(G21), .dout(new_n567_));
  anb2 g0503(.dina(new_n497_), .dinb(new_n500_), .dout(new_n568_));
  and1 g0504(.dina(G10), .dinb(G20), .dout(new_n569_));
  anb2 g0505(.dina(new_n491_), .dinb(new_n494_), .dout(new_n570_));
  and1 g0506(.dina(G11), .dinb(G19), .dout(new_n571_));
  nor2 g0507(.dina(G13), .dinb(G17), .dout(new_n572_));
  and1 g0508(.dina(G12), .dinb(G18), .dout(new_n573_));
  anb2 g0509(.dina(new_n572_), .dinb(new_n573_), .dout(new_n574_));
  anb1 g0510(.dina(new_n572_), .dinb(new_n573_), .dout(new_n575_));
  anb1 g0511(.dina(new_n574_), .dinb(new_n575_), .dout(new_n576_));
  anb1 g0512(.dina(new_n488_), .dinb(new_n576_), .dout(new_n577_));
  anb2 g0513(.dina(new_n488_), .dinb(new_n576_), .dout(new_n578_));
  nab1 g0514(.dina(new_n577_), .dinb(new_n578_), .dout(new_n579_));
  anb2 g0515(.dina(new_n571_), .dinb(new_n579_), .dout(new_n580_));
  anb1 g0516(.dina(new_n571_), .dinb(new_n579_), .dout(new_n581_));
  nab2 g0517(.dina(new_n580_), .dinb(new_n581_), .dout(new_n582_));
  anb1 g0518(.dina(new_n570_), .dinb(new_n582_), .dout(new_n583_));
  anb2 g0519(.dina(new_n570_), .dinb(new_n582_), .dout(new_n584_));
  nab1 g0520(.dina(new_n583_), .dinb(new_n584_), .dout(new_n585_));
  anb2 g0521(.dina(new_n569_), .dinb(new_n585_), .dout(new_n586_));
  anb1 g0522(.dina(new_n569_), .dinb(new_n585_), .dout(new_n587_));
  nab2 g0523(.dina(new_n586_), .dinb(new_n587_), .dout(new_n588_));
  anb1 g0524(.dina(new_n568_), .dinb(new_n588_), .dout(new_n589_));
  anb2 g0525(.dina(new_n568_), .dinb(new_n588_), .dout(new_n590_));
  nab1 g0526(.dina(new_n589_), .dinb(new_n590_), .dout(new_n591_));
  anb2 g0527(.dina(new_n567_), .dinb(new_n591_), .dout(new_n592_));
  anb1 g0528(.dina(new_n567_), .dinb(new_n591_), .dout(new_n593_));
  nab2 g0529(.dina(new_n592_), .dinb(new_n593_), .dout(new_n594_));
  anb1 g0530(.dina(new_n566_), .dinb(new_n594_), .dout(new_n595_));
  anb2 g0531(.dina(new_n566_), .dinb(new_n594_), .dout(new_n596_));
  nab1 g0532(.dina(new_n595_), .dinb(new_n596_), .dout(new_n597_));
  anb2 g0533(.dina(new_n565_), .dinb(new_n597_), .dout(new_n598_));
  anb1 g0534(.dina(new_n565_), .dinb(new_n597_), .dout(new_n599_));
  nab2 g0535(.dina(new_n598_), .dinb(new_n599_), .dout(new_n600_));
  anb1 g0536(.dina(new_n564_), .dinb(new_n600_), .dout(new_n601_));
  anb2 g0537(.dina(new_n564_), .dinb(new_n600_), .dout(new_n602_));
  nab1 g0538(.dina(new_n601_), .dinb(new_n602_), .dout(new_n603_));
  anb2 g0539(.dina(new_n563_), .dinb(new_n603_), .dout(new_n604_));
  anb1 g0540(.dina(new_n563_), .dinb(new_n603_), .dout(new_n605_));
  nab2 g0541(.dina(new_n604_), .dinb(new_n605_), .dout(new_n606_));
  anb1 g0542(.dina(new_n562_), .dinb(new_n606_), .dout(new_n607_));
  anb2 g0543(.dina(new_n562_), .dinb(new_n606_), .dout(new_n608_));
  nab1 g0544(.dina(new_n607_), .dinb(new_n608_), .dout(new_n609_));
  anb2 g0545(.dina(new_n561_), .dinb(new_n609_), .dout(new_n610_));
  anb1 g0546(.dina(new_n561_), .dinb(new_n609_), .dout(new_n611_));
  nab2 g0547(.dina(new_n610_), .dinb(new_n611_), .dout(new_n612_));
  anb1 g0548(.dina(new_n560_), .dinb(new_n612_), .dout(new_n613_));
  anb2 g0549(.dina(new_n560_), .dinb(new_n612_), .dout(new_n614_));
  nab1 g0550(.dina(new_n613_), .dinb(new_n614_), .dout(new_n615_));
  anb2 g0551(.dina(new_n559_), .dinb(new_n615_), .dout(new_n616_));
  anb1 g0552(.dina(new_n559_), .dinb(new_n615_), .dout(new_n617_));
  anb1 g0553(.dina(new_n616_), .dinb(new_n617_), .dout(new_n618_));
  anb2 g0554(.dina(new_n558_), .dinb(new_n618_), .dout(new_n619_));
  anb1 g0555(.dina(new_n558_), .dinb(new_n618_), .dout(new_n620_));
  nab2 g0556(.dina(new_n619_), .dinb(new_n620_), .dout(new_n621_));
  anb1 g0557(.dina(new_n557_), .dinb(new_n621_), .dout(new_n622_));
  anb2 g0558(.dina(new_n557_), .dinb(new_n621_), .dout(new_n623_));
  anb2 g0559(.dina(new_n622_), .dinb(new_n623_), .dout(new_n624_));
  anb1 g0560(.dina(new_n556_), .dinb(new_n624_), .dout(new_n625_));
  anb2 g0561(.dina(new_n556_), .dinb(new_n624_), .dout(new_n626_));
  anb2 g0562(.dina(new_n625_), .dinb(new_n626_), .dout(new_n627_));
  anb1 g0563(.dina(new_n555_), .dinb(new_n627_), .dout(new_n628_));
  anb2 g0564(.dina(new_n555_), .dinb(new_n627_), .dout(new_n629_));
  anb2 g0565(.dina(new_n628_), .dinb(new_n629_), .dout(new_n630_));
  anb1 g0566(.dina(new_n554_), .dinb(new_n630_), .dout(new_n631_));
  anb2 g0567(.dina(new_n554_), .dinb(new_n630_), .dout(new_n632_));
  anb2 g0568(.dina(new_n631_), .dinb(new_n632_), .dout(new_n633_));
  anb1 g0569(.dina(new_n553_), .dinb(new_n633_), .dout(new_n634_));
  anb2 g0570(.dina(new_n553_), .dinb(new_n633_), .dout(new_n635_));
  anb2 g0571(.dina(new_n634_), .dinb(new_n635_), .dout(new_n636_));
  anb1 g0572(.dina(new_n552_), .dinb(new_n636_), .dout(new_n637_));
  anb2 g0573(.dina(new_n552_), .dinb(new_n636_), .dout(new_n638_));
  anb2 g0574(.dina(new_n637_), .dinb(new_n638_), .dout(new_n639_));
  anb1 g0575(.dina(new_n551_), .dinb(new_n639_), .dout(new_n640_));
  anb2 g0576(.dina(new_n551_), .dinb(new_n639_), .dout(new_n641_));
  anb2 g0577(.dina(new_n640_), .dinb(new_n641_), .dout(G6269));
  nor2 g0578(.dina(G1), .dinb(G30), .dout(new_n643_));
  and2 g0579(.dina(new_n637_), .dinb(new_n640_), .dout(new_n644_));
  nor2 g0580(.dina(G2), .dinb(G29), .dout(new_n645_));
  and2 g0581(.dina(new_n631_), .dinb(new_n634_), .dout(new_n646_));
  nor2 g0582(.dina(G3), .dinb(G28), .dout(new_n647_));
  and2 g0583(.dina(new_n625_), .dinb(new_n628_), .dout(new_n648_));
  nor2 g0584(.dina(G4), .dinb(G27), .dout(new_n649_));
  anb1 g0585(.dina(new_n619_), .dinb(new_n622_), .dout(new_n650_));
  and1 g0586(.dina(G5), .dinb(G26), .dout(new_n651_));
  anb2 g0587(.dina(new_n613_), .dinb(new_n616_), .dout(new_n652_));
  and1 g0588(.dina(G6), .dinb(G25), .dout(new_n653_));
  anb2 g0589(.dina(new_n607_), .dinb(new_n610_), .dout(new_n654_));
  and1 g0590(.dina(G7), .dinb(G24), .dout(new_n655_));
  anb2 g0591(.dina(new_n601_), .dinb(new_n604_), .dout(new_n656_));
  and1 g0592(.dina(G8), .dinb(G23), .dout(new_n657_));
  anb2 g0593(.dina(new_n595_), .dinb(new_n598_), .dout(new_n658_));
  and1 g0594(.dina(G9), .dinb(G22), .dout(new_n659_));
  anb2 g0595(.dina(new_n589_), .dinb(new_n592_), .dout(new_n660_));
  and1 g0596(.dina(G10), .dinb(G21), .dout(new_n661_));
  anb2 g0597(.dina(new_n583_), .dinb(new_n586_), .dout(new_n662_));
  and1 g0598(.dina(G11), .dinb(G20), .dout(new_n663_));
  anb2 g0599(.dina(new_n577_), .dinb(new_n580_), .dout(new_n664_));
  and1 g0600(.dina(G12), .dinb(G19), .dout(new_n665_));
  nor2 g0601(.dina(G14), .dinb(G17), .dout(new_n666_));
  and1 g0602(.dina(G13), .dinb(G18), .dout(new_n667_));
  anb2 g0603(.dina(new_n666_), .dinb(new_n667_), .dout(new_n668_));
  anb1 g0604(.dina(new_n666_), .dinb(new_n667_), .dout(new_n669_));
  anb1 g0605(.dina(new_n668_), .dinb(new_n669_), .dout(new_n670_));
  anb1 g0606(.dina(new_n574_), .dinb(new_n670_), .dout(new_n671_));
  anb2 g0607(.dina(new_n574_), .dinb(new_n670_), .dout(new_n672_));
  nab1 g0608(.dina(new_n671_), .dinb(new_n672_), .dout(new_n673_));
  anb2 g0609(.dina(new_n665_), .dinb(new_n673_), .dout(new_n674_));
  anb1 g0610(.dina(new_n665_), .dinb(new_n673_), .dout(new_n675_));
  nab2 g0611(.dina(new_n674_), .dinb(new_n675_), .dout(new_n676_));
  anb1 g0612(.dina(new_n664_), .dinb(new_n676_), .dout(new_n677_));
  anb2 g0613(.dina(new_n664_), .dinb(new_n676_), .dout(new_n678_));
  nab1 g0614(.dina(new_n677_), .dinb(new_n678_), .dout(new_n679_));
  anb2 g0615(.dina(new_n663_), .dinb(new_n679_), .dout(new_n680_));
  anb1 g0616(.dina(new_n663_), .dinb(new_n679_), .dout(new_n681_));
  nab2 g0617(.dina(new_n680_), .dinb(new_n681_), .dout(new_n682_));
  anb1 g0618(.dina(new_n662_), .dinb(new_n682_), .dout(new_n683_));
  anb2 g0619(.dina(new_n662_), .dinb(new_n682_), .dout(new_n684_));
  nab1 g0620(.dina(new_n683_), .dinb(new_n684_), .dout(new_n685_));
  anb2 g0621(.dina(new_n661_), .dinb(new_n685_), .dout(new_n686_));
  anb1 g0622(.dina(new_n661_), .dinb(new_n685_), .dout(new_n687_));
  nab2 g0623(.dina(new_n686_), .dinb(new_n687_), .dout(new_n688_));
  anb1 g0624(.dina(new_n660_), .dinb(new_n688_), .dout(new_n689_));
  anb2 g0625(.dina(new_n660_), .dinb(new_n688_), .dout(new_n690_));
  nab1 g0626(.dina(new_n689_), .dinb(new_n690_), .dout(new_n691_));
  anb2 g0627(.dina(new_n659_), .dinb(new_n691_), .dout(new_n692_));
  anb1 g0628(.dina(new_n659_), .dinb(new_n691_), .dout(new_n693_));
  nab2 g0629(.dina(new_n692_), .dinb(new_n693_), .dout(new_n694_));
  anb1 g0630(.dina(new_n658_), .dinb(new_n694_), .dout(new_n695_));
  anb2 g0631(.dina(new_n658_), .dinb(new_n694_), .dout(new_n696_));
  nab1 g0632(.dina(new_n695_), .dinb(new_n696_), .dout(new_n697_));
  anb2 g0633(.dina(new_n657_), .dinb(new_n697_), .dout(new_n698_));
  anb1 g0634(.dina(new_n657_), .dinb(new_n697_), .dout(new_n699_));
  nab2 g0635(.dina(new_n698_), .dinb(new_n699_), .dout(new_n700_));
  anb1 g0636(.dina(new_n656_), .dinb(new_n700_), .dout(new_n701_));
  anb2 g0637(.dina(new_n656_), .dinb(new_n700_), .dout(new_n702_));
  nab1 g0638(.dina(new_n701_), .dinb(new_n702_), .dout(new_n703_));
  anb2 g0639(.dina(new_n655_), .dinb(new_n703_), .dout(new_n704_));
  anb1 g0640(.dina(new_n655_), .dinb(new_n703_), .dout(new_n705_));
  nab2 g0641(.dina(new_n704_), .dinb(new_n705_), .dout(new_n706_));
  anb1 g0642(.dina(new_n654_), .dinb(new_n706_), .dout(new_n707_));
  anb2 g0643(.dina(new_n654_), .dinb(new_n706_), .dout(new_n708_));
  nab1 g0644(.dina(new_n707_), .dinb(new_n708_), .dout(new_n709_));
  anb2 g0645(.dina(new_n653_), .dinb(new_n709_), .dout(new_n710_));
  anb1 g0646(.dina(new_n653_), .dinb(new_n709_), .dout(new_n711_));
  nab2 g0647(.dina(new_n710_), .dinb(new_n711_), .dout(new_n712_));
  anb1 g0648(.dina(new_n652_), .dinb(new_n712_), .dout(new_n713_));
  anb2 g0649(.dina(new_n652_), .dinb(new_n712_), .dout(new_n714_));
  nab1 g0650(.dina(new_n713_), .dinb(new_n714_), .dout(new_n715_));
  anb2 g0651(.dina(new_n651_), .dinb(new_n715_), .dout(new_n716_));
  anb1 g0652(.dina(new_n651_), .dinb(new_n715_), .dout(new_n717_));
  anb1 g0653(.dina(new_n716_), .dinb(new_n717_), .dout(new_n718_));
  anb2 g0654(.dina(new_n650_), .dinb(new_n718_), .dout(new_n719_));
  anb1 g0655(.dina(new_n650_), .dinb(new_n718_), .dout(new_n720_));
  nab2 g0656(.dina(new_n719_), .dinb(new_n720_), .dout(new_n721_));
  anb1 g0657(.dina(new_n649_), .dinb(new_n721_), .dout(new_n722_));
  anb2 g0658(.dina(new_n649_), .dinb(new_n721_), .dout(new_n723_));
  anb2 g0659(.dina(new_n722_), .dinb(new_n723_), .dout(new_n724_));
  anb1 g0660(.dina(new_n648_), .dinb(new_n724_), .dout(new_n725_));
  anb2 g0661(.dina(new_n648_), .dinb(new_n724_), .dout(new_n726_));
  anb2 g0662(.dina(new_n725_), .dinb(new_n726_), .dout(new_n727_));
  anb1 g0663(.dina(new_n647_), .dinb(new_n727_), .dout(new_n728_));
  anb2 g0664(.dina(new_n647_), .dinb(new_n727_), .dout(new_n729_));
  anb2 g0665(.dina(new_n728_), .dinb(new_n729_), .dout(new_n730_));
  anb1 g0666(.dina(new_n646_), .dinb(new_n730_), .dout(new_n731_));
  anb2 g0667(.dina(new_n646_), .dinb(new_n730_), .dout(new_n732_));
  anb2 g0668(.dina(new_n731_), .dinb(new_n732_), .dout(new_n733_));
  anb1 g0669(.dina(new_n645_), .dinb(new_n733_), .dout(new_n734_));
  anb2 g0670(.dina(new_n645_), .dinb(new_n733_), .dout(new_n735_));
  anb2 g0671(.dina(new_n734_), .dinb(new_n735_), .dout(new_n736_));
  anb1 g0672(.dina(new_n644_), .dinb(new_n736_), .dout(new_n737_));
  anb2 g0673(.dina(new_n644_), .dinb(new_n736_), .dout(new_n738_));
  anb2 g0674(.dina(new_n737_), .dinb(new_n738_), .dout(new_n739_));
  anb1 g0675(.dina(new_n643_), .dinb(new_n739_), .dout(new_n740_));
  anb2 g0676(.dina(new_n643_), .dinb(new_n739_), .dout(new_n741_));
  anb2 g0677(.dina(new_n740_), .dinb(new_n741_), .dout(G6270));
  nor2 g0678(.dina(G1), .dinb(G31), .dout(new_n743_));
  and2 g0679(.dina(new_n737_), .dinb(new_n740_), .dout(new_n744_));
  nor2 g0680(.dina(G2), .dinb(G30), .dout(new_n745_));
  and2 g0681(.dina(new_n731_), .dinb(new_n734_), .dout(new_n746_));
  nor2 g0682(.dina(G3), .dinb(G29), .dout(new_n747_));
  and2 g0683(.dina(new_n725_), .dinb(new_n728_), .dout(new_n748_));
  nor2 g0684(.dina(G4), .dinb(G28), .dout(new_n749_));
  anb1 g0685(.dina(new_n719_), .dinb(new_n722_), .dout(new_n750_));
  and1 g0686(.dina(G5), .dinb(G27), .dout(new_n751_));
  anb2 g0687(.dina(new_n713_), .dinb(new_n716_), .dout(new_n752_));
  and1 g0688(.dina(G6), .dinb(G26), .dout(new_n753_));
  anb2 g0689(.dina(new_n707_), .dinb(new_n710_), .dout(new_n754_));
  and1 g0690(.dina(G7), .dinb(G25), .dout(new_n755_));
  anb2 g0691(.dina(new_n701_), .dinb(new_n704_), .dout(new_n756_));
  and1 g0692(.dina(G8), .dinb(G24), .dout(new_n757_));
  anb2 g0693(.dina(new_n695_), .dinb(new_n698_), .dout(new_n758_));
  and1 g0694(.dina(G9), .dinb(G23), .dout(new_n759_));
  anb2 g0695(.dina(new_n689_), .dinb(new_n692_), .dout(new_n760_));
  and1 g0696(.dina(G10), .dinb(G22), .dout(new_n761_));
  anb2 g0697(.dina(new_n683_), .dinb(new_n686_), .dout(new_n762_));
  and1 g0698(.dina(G11), .dinb(G21), .dout(new_n763_));
  anb2 g0699(.dina(new_n677_), .dinb(new_n680_), .dout(new_n764_));
  and1 g0700(.dina(G12), .dinb(G20), .dout(new_n765_));
  anb2 g0701(.dina(new_n671_), .dinb(new_n674_), .dout(new_n766_));
  and1 g0702(.dina(G13), .dinb(G19), .dout(new_n767_));
  nor2 g0703(.dina(G15), .dinb(G17), .dout(new_n768_));
  and1 g0704(.dina(G14), .dinb(G18), .dout(new_n769_));
  anb2 g0705(.dina(new_n768_), .dinb(new_n769_), .dout(new_n770_));
  anb1 g0706(.dina(new_n768_), .dinb(new_n769_), .dout(new_n771_));
  anb1 g0707(.dina(new_n770_), .dinb(new_n771_), .dout(new_n772_));
  anb1 g0708(.dina(new_n668_), .dinb(new_n772_), .dout(new_n773_));
  anb2 g0709(.dina(new_n668_), .dinb(new_n772_), .dout(new_n774_));
  nab1 g0710(.dina(new_n773_), .dinb(new_n774_), .dout(new_n775_));
  anb2 g0711(.dina(new_n767_), .dinb(new_n775_), .dout(new_n776_));
  anb1 g0712(.dina(new_n767_), .dinb(new_n775_), .dout(new_n777_));
  nab2 g0713(.dina(new_n776_), .dinb(new_n777_), .dout(new_n778_));
  anb1 g0714(.dina(new_n766_), .dinb(new_n778_), .dout(new_n779_));
  anb2 g0715(.dina(new_n766_), .dinb(new_n778_), .dout(new_n780_));
  nab1 g0716(.dina(new_n779_), .dinb(new_n780_), .dout(new_n781_));
  anb2 g0717(.dina(new_n765_), .dinb(new_n781_), .dout(new_n782_));
  anb1 g0718(.dina(new_n765_), .dinb(new_n781_), .dout(new_n783_));
  nab2 g0719(.dina(new_n782_), .dinb(new_n783_), .dout(new_n784_));
  anb1 g0720(.dina(new_n764_), .dinb(new_n784_), .dout(new_n785_));
  anb2 g0721(.dina(new_n764_), .dinb(new_n784_), .dout(new_n786_));
  nab1 g0722(.dina(new_n785_), .dinb(new_n786_), .dout(new_n787_));
  anb2 g0723(.dina(new_n763_), .dinb(new_n787_), .dout(new_n788_));
  anb1 g0724(.dina(new_n763_), .dinb(new_n787_), .dout(new_n789_));
  nab2 g0725(.dina(new_n788_), .dinb(new_n789_), .dout(new_n790_));
  anb1 g0726(.dina(new_n762_), .dinb(new_n790_), .dout(new_n791_));
  anb2 g0727(.dina(new_n762_), .dinb(new_n790_), .dout(new_n792_));
  nab1 g0728(.dina(new_n791_), .dinb(new_n792_), .dout(new_n793_));
  anb2 g0729(.dina(new_n761_), .dinb(new_n793_), .dout(new_n794_));
  anb1 g0730(.dina(new_n761_), .dinb(new_n793_), .dout(new_n795_));
  nab2 g0731(.dina(new_n794_), .dinb(new_n795_), .dout(new_n796_));
  anb1 g0732(.dina(new_n760_), .dinb(new_n796_), .dout(new_n797_));
  anb2 g0733(.dina(new_n760_), .dinb(new_n796_), .dout(new_n798_));
  nab1 g0734(.dina(new_n797_), .dinb(new_n798_), .dout(new_n799_));
  anb2 g0735(.dina(new_n759_), .dinb(new_n799_), .dout(new_n800_));
  anb1 g0736(.dina(new_n759_), .dinb(new_n799_), .dout(new_n801_));
  nab2 g0737(.dina(new_n800_), .dinb(new_n801_), .dout(new_n802_));
  anb1 g0738(.dina(new_n758_), .dinb(new_n802_), .dout(new_n803_));
  anb2 g0739(.dina(new_n758_), .dinb(new_n802_), .dout(new_n804_));
  nab1 g0740(.dina(new_n803_), .dinb(new_n804_), .dout(new_n805_));
  anb2 g0741(.dina(new_n757_), .dinb(new_n805_), .dout(new_n806_));
  anb1 g0742(.dina(new_n757_), .dinb(new_n805_), .dout(new_n807_));
  nab2 g0743(.dina(new_n806_), .dinb(new_n807_), .dout(new_n808_));
  anb1 g0744(.dina(new_n756_), .dinb(new_n808_), .dout(new_n809_));
  anb2 g0745(.dina(new_n756_), .dinb(new_n808_), .dout(new_n810_));
  nab1 g0746(.dina(new_n809_), .dinb(new_n810_), .dout(new_n811_));
  anb2 g0747(.dina(new_n755_), .dinb(new_n811_), .dout(new_n812_));
  anb1 g0748(.dina(new_n755_), .dinb(new_n811_), .dout(new_n813_));
  nab2 g0749(.dina(new_n812_), .dinb(new_n813_), .dout(new_n814_));
  anb1 g0750(.dina(new_n754_), .dinb(new_n814_), .dout(new_n815_));
  anb2 g0751(.dina(new_n754_), .dinb(new_n814_), .dout(new_n816_));
  nab1 g0752(.dina(new_n815_), .dinb(new_n816_), .dout(new_n817_));
  anb2 g0753(.dina(new_n753_), .dinb(new_n817_), .dout(new_n818_));
  anb1 g0754(.dina(new_n753_), .dinb(new_n817_), .dout(new_n819_));
  nab2 g0755(.dina(new_n818_), .dinb(new_n819_), .dout(new_n820_));
  anb1 g0756(.dina(new_n752_), .dinb(new_n820_), .dout(new_n821_));
  anb2 g0757(.dina(new_n752_), .dinb(new_n820_), .dout(new_n822_));
  nab1 g0758(.dina(new_n821_), .dinb(new_n822_), .dout(new_n823_));
  anb2 g0759(.dina(new_n751_), .dinb(new_n823_), .dout(new_n824_));
  anb1 g0760(.dina(new_n751_), .dinb(new_n823_), .dout(new_n825_));
  anb1 g0761(.dina(new_n824_), .dinb(new_n825_), .dout(new_n826_));
  anb2 g0762(.dina(new_n750_), .dinb(new_n826_), .dout(new_n827_));
  anb1 g0763(.dina(new_n750_), .dinb(new_n826_), .dout(new_n828_));
  nab2 g0764(.dina(new_n827_), .dinb(new_n828_), .dout(new_n829_));
  anb1 g0765(.dina(new_n749_), .dinb(new_n829_), .dout(new_n830_));
  anb2 g0766(.dina(new_n749_), .dinb(new_n829_), .dout(new_n831_));
  anb2 g0767(.dina(new_n830_), .dinb(new_n831_), .dout(new_n832_));
  anb1 g0768(.dina(new_n748_), .dinb(new_n832_), .dout(new_n833_));
  anb2 g0769(.dina(new_n748_), .dinb(new_n832_), .dout(new_n834_));
  anb2 g0770(.dina(new_n833_), .dinb(new_n834_), .dout(new_n835_));
  anb1 g0771(.dina(new_n747_), .dinb(new_n835_), .dout(new_n836_));
  anb2 g0772(.dina(new_n747_), .dinb(new_n835_), .dout(new_n837_));
  anb2 g0773(.dina(new_n836_), .dinb(new_n837_), .dout(new_n838_));
  anb1 g0774(.dina(new_n746_), .dinb(new_n838_), .dout(new_n839_));
  anb2 g0775(.dina(new_n746_), .dinb(new_n838_), .dout(new_n840_));
  anb2 g0776(.dina(new_n839_), .dinb(new_n840_), .dout(new_n841_));
  anb1 g0777(.dina(new_n745_), .dinb(new_n841_), .dout(new_n842_));
  anb2 g0778(.dina(new_n745_), .dinb(new_n841_), .dout(new_n843_));
  anb2 g0779(.dina(new_n842_), .dinb(new_n843_), .dout(new_n844_));
  anb1 g0780(.dina(new_n744_), .dinb(new_n844_), .dout(new_n845_));
  anb2 g0781(.dina(new_n744_), .dinb(new_n844_), .dout(new_n846_));
  anb2 g0782(.dina(new_n845_), .dinb(new_n846_), .dout(new_n847_));
  anb1 g0783(.dina(new_n743_), .dinb(new_n847_), .dout(new_n848_));
  anb2 g0784(.dina(new_n743_), .dinb(new_n847_), .dout(new_n849_));
  anb2 g0785(.dina(new_n848_), .dinb(new_n849_), .dout(G6271));
  nor2 g0786(.dina(G1), .dinb(G32), .dout(new_n851_));
  and2 g0787(.dina(new_n845_), .dinb(new_n848_), .dout(new_n852_));
  nor2 g0788(.dina(G2), .dinb(G31), .dout(new_n853_));
  and2 g0789(.dina(new_n839_), .dinb(new_n842_), .dout(new_n854_));
  nor2 g0790(.dina(G3), .dinb(G30), .dout(new_n855_));
  and2 g0791(.dina(new_n833_), .dinb(new_n836_), .dout(new_n856_));
  nor2 g0792(.dina(G4), .dinb(G29), .dout(new_n857_));
  anb1 g0793(.dina(new_n827_), .dinb(new_n830_), .dout(new_n858_));
  and1 g0794(.dina(G5), .dinb(G28), .dout(new_n859_));
  anb2 g0795(.dina(new_n821_), .dinb(new_n824_), .dout(new_n860_));
  and1 g0796(.dina(G6), .dinb(G27), .dout(new_n861_));
  anb2 g0797(.dina(new_n815_), .dinb(new_n818_), .dout(new_n862_));
  and1 g0798(.dina(G7), .dinb(G26), .dout(new_n863_));
  anb2 g0799(.dina(new_n809_), .dinb(new_n812_), .dout(new_n864_));
  and1 g0800(.dina(G8), .dinb(G25), .dout(new_n865_));
  anb2 g0801(.dina(new_n803_), .dinb(new_n806_), .dout(new_n866_));
  and1 g0802(.dina(G9), .dinb(G24), .dout(new_n867_));
  anb2 g0803(.dina(new_n797_), .dinb(new_n800_), .dout(new_n868_));
  and1 g0804(.dina(G10), .dinb(G23), .dout(new_n869_));
  anb2 g0805(.dina(new_n791_), .dinb(new_n794_), .dout(new_n870_));
  and1 g0806(.dina(G11), .dinb(G22), .dout(new_n871_));
  anb2 g0807(.dina(new_n785_), .dinb(new_n788_), .dout(new_n872_));
  and1 g0808(.dina(G12), .dinb(G21), .dout(new_n873_));
  anb2 g0809(.dina(new_n779_), .dinb(new_n782_), .dout(new_n874_));
  and1 g0810(.dina(G13), .dinb(G20), .dout(new_n875_));
  anb2 g0811(.dina(new_n773_), .dinb(new_n776_), .dout(new_n876_));
  and1 g0812(.dina(G14), .dinb(G19), .dout(new_n877_));
  and1 g0813(.dina(G16), .dinb(G17), .dout(new_n878_));
  nor2 g0814(.dina(G15), .dinb(G18), .dout(new_n879_));
  anb1 g0815(.dina(new_n878_), .dinb(new_n879_), .dout(new_n880_));
  anb2 g0816(.dina(new_n878_), .dinb(new_n879_), .dout(new_n881_));
  nab1 g0817(.dina(new_n880_), .dinb(new_n881_), .dout(new_n882_));
  anb1 g0818(.dina(new_n770_), .dinb(new_n882_), .dout(new_n883_));
  anb2 g0819(.dina(new_n770_), .dinb(new_n882_), .dout(new_n884_));
  nab1 g0820(.dina(new_n883_), .dinb(new_n884_), .dout(new_n885_));
  anb2 g0821(.dina(new_n877_), .dinb(new_n885_), .dout(new_n886_));
  anb1 g0822(.dina(new_n877_), .dinb(new_n885_), .dout(new_n887_));
  nab2 g0823(.dina(new_n886_), .dinb(new_n887_), .dout(new_n888_));
  anb1 g0824(.dina(new_n876_), .dinb(new_n888_), .dout(new_n889_));
  anb2 g0825(.dina(new_n876_), .dinb(new_n888_), .dout(new_n890_));
  nab1 g0826(.dina(new_n889_), .dinb(new_n890_), .dout(new_n891_));
  anb2 g0827(.dina(new_n875_), .dinb(new_n891_), .dout(new_n892_));
  anb1 g0828(.dina(new_n875_), .dinb(new_n891_), .dout(new_n893_));
  nab2 g0829(.dina(new_n892_), .dinb(new_n893_), .dout(new_n894_));
  anb1 g0830(.dina(new_n874_), .dinb(new_n894_), .dout(new_n895_));
  anb2 g0831(.dina(new_n874_), .dinb(new_n894_), .dout(new_n896_));
  nab1 g0832(.dina(new_n895_), .dinb(new_n896_), .dout(new_n897_));
  anb2 g0833(.dina(new_n873_), .dinb(new_n897_), .dout(new_n898_));
  anb1 g0834(.dina(new_n873_), .dinb(new_n897_), .dout(new_n899_));
  nab2 g0835(.dina(new_n898_), .dinb(new_n899_), .dout(new_n900_));
  anb1 g0836(.dina(new_n872_), .dinb(new_n900_), .dout(new_n901_));
  anb2 g0837(.dina(new_n872_), .dinb(new_n900_), .dout(new_n902_));
  nab1 g0838(.dina(new_n901_), .dinb(new_n902_), .dout(new_n903_));
  anb2 g0839(.dina(new_n871_), .dinb(new_n903_), .dout(new_n904_));
  anb1 g0840(.dina(new_n871_), .dinb(new_n903_), .dout(new_n905_));
  nab2 g0841(.dina(new_n904_), .dinb(new_n905_), .dout(new_n906_));
  anb1 g0842(.dina(new_n870_), .dinb(new_n906_), .dout(new_n907_));
  anb2 g0843(.dina(new_n870_), .dinb(new_n906_), .dout(new_n908_));
  nab1 g0844(.dina(new_n907_), .dinb(new_n908_), .dout(new_n909_));
  anb2 g0845(.dina(new_n869_), .dinb(new_n909_), .dout(new_n910_));
  anb1 g0846(.dina(new_n869_), .dinb(new_n909_), .dout(new_n911_));
  nab2 g0847(.dina(new_n910_), .dinb(new_n911_), .dout(new_n912_));
  anb1 g0848(.dina(new_n868_), .dinb(new_n912_), .dout(new_n913_));
  anb2 g0849(.dina(new_n868_), .dinb(new_n912_), .dout(new_n914_));
  nab1 g0850(.dina(new_n913_), .dinb(new_n914_), .dout(new_n915_));
  anb2 g0851(.dina(new_n867_), .dinb(new_n915_), .dout(new_n916_));
  anb1 g0852(.dina(new_n867_), .dinb(new_n915_), .dout(new_n917_));
  nab2 g0853(.dina(new_n916_), .dinb(new_n917_), .dout(new_n918_));
  anb1 g0854(.dina(new_n866_), .dinb(new_n918_), .dout(new_n919_));
  anb2 g0855(.dina(new_n866_), .dinb(new_n918_), .dout(new_n920_));
  nab1 g0856(.dina(new_n919_), .dinb(new_n920_), .dout(new_n921_));
  anb2 g0857(.dina(new_n865_), .dinb(new_n921_), .dout(new_n922_));
  anb1 g0858(.dina(new_n865_), .dinb(new_n921_), .dout(new_n923_));
  nab2 g0859(.dina(new_n922_), .dinb(new_n923_), .dout(new_n924_));
  anb1 g0860(.dina(new_n864_), .dinb(new_n924_), .dout(new_n925_));
  anb2 g0861(.dina(new_n864_), .dinb(new_n924_), .dout(new_n926_));
  nab1 g0862(.dina(new_n925_), .dinb(new_n926_), .dout(new_n927_));
  anb2 g0863(.dina(new_n863_), .dinb(new_n927_), .dout(new_n928_));
  anb1 g0864(.dina(new_n863_), .dinb(new_n927_), .dout(new_n929_));
  nab2 g0865(.dina(new_n928_), .dinb(new_n929_), .dout(new_n930_));
  anb1 g0866(.dina(new_n862_), .dinb(new_n930_), .dout(new_n931_));
  anb2 g0867(.dina(new_n862_), .dinb(new_n930_), .dout(new_n932_));
  nab1 g0868(.dina(new_n931_), .dinb(new_n932_), .dout(new_n933_));
  anb2 g0869(.dina(new_n861_), .dinb(new_n933_), .dout(new_n934_));
  anb1 g0870(.dina(new_n861_), .dinb(new_n933_), .dout(new_n935_));
  nab2 g0871(.dina(new_n934_), .dinb(new_n935_), .dout(new_n936_));
  anb1 g0872(.dina(new_n860_), .dinb(new_n936_), .dout(new_n937_));
  anb2 g0873(.dina(new_n860_), .dinb(new_n936_), .dout(new_n938_));
  nab1 g0874(.dina(new_n937_), .dinb(new_n938_), .dout(new_n939_));
  anb2 g0875(.dina(new_n859_), .dinb(new_n939_), .dout(new_n940_));
  anb1 g0876(.dina(new_n859_), .dinb(new_n939_), .dout(new_n941_));
  anb1 g0877(.dina(new_n940_), .dinb(new_n941_), .dout(new_n942_));
  anb2 g0878(.dina(new_n858_), .dinb(new_n942_), .dout(new_n943_));
  anb1 g0879(.dina(new_n858_), .dinb(new_n942_), .dout(new_n944_));
  nab2 g0880(.dina(new_n943_), .dinb(new_n944_), .dout(new_n945_));
  anb1 g0881(.dina(new_n857_), .dinb(new_n945_), .dout(new_n946_));
  anb2 g0882(.dina(new_n857_), .dinb(new_n945_), .dout(new_n947_));
  anb2 g0883(.dina(new_n946_), .dinb(new_n947_), .dout(new_n948_));
  anb1 g0884(.dina(new_n856_), .dinb(new_n948_), .dout(new_n949_));
  anb2 g0885(.dina(new_n856_), .dinb(new_n948_), .dout(new_n950_));
  anb2 g0886(.dina(new_n949_), .dinb(new_n950_), .dout(new_n951_));
  anb1 g0887(.dina(new_n855_), .dinb(new_n951_), .dout(new_n952_));
  anb2 g0888(.dina(new_n855_), .dinb(new_n951_), .dout(new_n953_));
  anb2 g0889(.dina(new_n952_), .dinb(new_n953_), .dout(new_n954_));
  anb1 g0890(.dina(new_n854_), .dinb(new_n954_), .dout(new_n955_));
  anb2 g0891(.dina(new_n854_), .dinb(new_n954_), .dout(new_n956_));
  anb2 g0892(.dina(new_n955_), .dinb(new_n956_), .dout(new_n957_));
  anb1 g0893(.dina(new_n853_), .dinb(new_n957_), .dout(new_n958_));
  anb2 g0894(.dina(new_n853_), .dinb(new_n957_), .dout(new_n959_));
  anb2 g0895(.dina(new_n958_), .dinb(new_n959_), .dout(new_n960_));
  anb1 g0896(.dina(new_n852_), .dinb(new_n960_), .dout(new_n961_));
  anb2 g0897(.dina(new_n852_), .dinb(new_n960_), .dout(new_n962_));
  anb2 g0898(.dina(new_n961_), .dinb(new_n962_), .dout(new_n963_));
  anb1 g0899(.dina(new_n851_), .dinb(new_n963_), .dout(new_n964_));
  anb2 g0900(.dina(new_n851_), .dinb(new_n963_), .dout(new_n965_));
  anb2 g0901(.dina(new_n964_), .dinb(new_n965_), .dout(G6272));
  nor1 g0902(.dina(new_n961_), .dinb(new_n964_), .dout(new_n967_));
  and1 g0903(.dina(G2), .dinb(G32), .dout(new_n968_));
  nor1 g0904(.dina(new_n955_), .dinb(new_n958_), .dout(new_n969_));
  and1 g0905(.dina(G3), .dinb(G31), .dout(new_n970_));
  nor1 g0906(.dina(new_n949_), .dinb(new_n952_), .dout(new_n971_));
  and1 g0907(.dina(G4), .dinb(G30), .dout(new_n972_));
  anb1 g0908(.dina(new_n943_), .dinb(new_n946_), .dout(new_n973_));
  and1 g0909(.dina(G5), .dinb(G29), .dout(new_n974_));
  anb2 g0910(.dina(new_n937_), .dinb(new_n940_), .dout(new_n975_));
  and1 g0911(.dina(G6), .dinb(G28), .dout(new_n976_));
  anb2 g0912(.dina(new_n931_), .dinb(new_n934_), .dout(new_n977_));
  and1 g0913(.dina(G7), .dinb(G27), .dout(new_n978_));
  anb2 g0914(.dina(new_n925_), .dinb(new_n928_), .dout(new_n979_));
  and1 g0915(.dina(G8), .dinb(G26), .dout(new_n980_));
  anb2 g0916(.dina(new_n919_), .dinb(new_n922_), .dout(new_n981_));
  and1 g0917(.dina(G9), .dinb(G25), .dout(new_n982_));
  anb2 g0918(.dina(new_n913_), .dinb(new_n916_), .dout(new_n983_));
  and1 g0919(.dina(G10), .dinb(G24), .dout(new_n984_));
  anb2 g0920(.dina(new_n907_), .dinb(new_n910_), .dout(new_n985_));
  and1 g0921(.dina(G11), .dinb(G23), .dout(new_n986_));
  anb2 g0922(.dina(new_n901_), .dinb(new_n904_), .dout(new_n987_));
  and1 g0923(.dina(G12), .dinb(G22), .dout(new_n988_));
  anb2 g0924(.dina(new_n895_), .dinb(new_n898_), .dout(new_n989_));
  and1 g0925(.dina(G13), .dinb(G21), .dout(new_n990_));
  anb2 g0926(.dina(new_n889_), .dinb(new_n892_), .dout(new_n991_));
  and1 g0927(.dina(G14), .dinb(G20), .dout(new_n992_));
  anb2 g0928(.dina(new_n883_), .dinb(new_n886_), .dout(new_n993_));
  and1 g0929(.dina(G16), .dinb(G18), .dout(new_n994_));
  anb1 g0930(.dina(new_n994_), .dinb(new_n880_), .dout(new_n995_));
  and1 g0931(.dina(G15), .dinb(G19), .dout(new_n996_));
  anb1 g0932(.dina(new_n995_), .dinb(new_n996_), .dout(new_n997_));
  anb2 g0933(.dina(new_n995_), .dinb(new_n996_), .dout(new_n998_));
  anb2 g0934(.dina(new_n997_), .dinb(new_n998_), .dout(new_n999_));
  anb1 g0935(.dina(new_n993_), .dinb(new_n999_), .dout(new_n1000_));
  anb2 g0936(.dina(new_n993_), .dinb(new_n999_), .dout(new_n1001_));
  nab1 g0937(.dina(new_n1000_), .dinb(new_n1001_), .dout(new_n1002_));
  anb2 g0938(.dina(new_n992_), .dinb(new_n1002_), .dout(new_n1003_));
  anb1 g0939(.dina(new_n992_), .dinb(new_n1002_), .dout(new_n1004_));
  nab2 g0940(.dina(new_n1003_), .dinb(new_n1004_), .dout(new_n1005_));
  anb1 g0941(.dina(new_n991_), .dinb(new_n1005_), .dout(new_n1006_));
  anb2 g0942(.dina(new_n991_), .dinb(new_n1005_), .dout(new_n1007_));
  nab1 g0943(.dina(new_n1006_), .dinb(new_n1007_), .dout(new_n1008_));
  anb2 g0944(.dina(new_n990_), .dinb(new_n1008_), .dout(new_n1009_));
  anb1 g0945(.dina(new_n990_), .dinb(new_n1008_), .dout(new_n1010_));
  nab2 g0946(.dina(new_n1009_), .dinb(new_n1010_), .dout(new_n1011_));
  anb1 g0947(.dina(new_n989_), .dinb(new_n1011_), .dout(new_n1012_));
  anb2 g0948(.dina(new_n989_), .dinb(new_n1011_), .dout(new_n1013_));
  nab1 g0949(.dina(new_n1012_), .dinb(new_n1013_), .dout(new_n1014_));
  anb2 g0950(.dina(new_n988_), .dinb(new_n1014_), .dout(new_n1015_));
  anb1 g0951(.dina(new_n988_), .dinb(new_n1014_), .dout(new_n1016_));
  nab2 g0952(.dina(new_n1015_), .dinb(new_n1016_), .dout(new_n1017_));
  anb1 g0953(.dina(new_n987_), .dinb(new_n1017_), .dout(new_n1018_));
  anb2 g0954(.dina(new_n987_), .dinb(new_n1017_), .dout(new_n1019_));
  nab1 g0955(.dina(new_n1018_), .dinb(new_n1019_), .dout(new_n1020_));
  anb2 g0956(.dina(new_n986_), .dinb(new_n1020_), .dout(new_n1021_));
  anb1 g0957(.dina(new_n986_), .dinb(new_n1020_), .dout(new_n1022_));
  nab2 g0958(.dina(new_n1021_), .dinb(new_n1022_), .dout(new_n1023_));
  anb1 g0959(.dina(new_n985_), .dinb(new_n1023_), .dout(new_n1024_));
  anb2 g0960(.dina(new_n985_), .dinb(new_n1023_), .dout(new_n1025_));
  nab1 g0961(.dina(new_n1024_), .dinb(new_n1025_), .dout(new_n1026_));
  anb2 g0962(.dina(new_n984_), .dinb(new_n1026_), .dout(new_n1027_));
  anb1 g0963(.dina(new_n984_), .dinb(new_n1026_), .dout(new_n1028_));
  nab2 g0964(.dina(new_n1027_), .dinb(new_n1028_), .dout(new_n1029_));
  anb1 g0965(.dina(new_n983_), .dinb(new_n1029_), .dout(new_n1030_));
  anb2 g0966(.dina(new_n983_), .dinb(new_n1029_), .dout(new_n1031_));
  nab1 g0967(.dina(new_n1030_), .dinb(new_n1031_), .dout(new_n1032_));
  anb2 g0968(.dina(new_n982_), .dinb(new_n1032_), .dout(new_n1033_));
  anb1 g0969(.dina(new_n982_), .dinb(new_n1032_), .dout(new_n1034_));
  nab2 g0970(.dina(new_n1033_), .dinb(new_n1034_), .dout(new_n1035_));
  anb1 g0971(.dina(new_n981_), .dinb(new_n1035_), .dout(new_n1036_));
  anb2 g0972(.dina(new_n981_), .dinb(new_n1035_), .dout(new_n1037_));
  nab1 g0973(.dina(new_n1036_), .dinb(new_n1037_), .dout(new_n1038_));
  anb2 g0974(.dina(new_n980_), .dinb(new_n1038_), .dout(new_n1039_));
  anb1 g0975(.dina(new_n980_), .dinb(new_n1038_), .dout(new_n1040_));
  nab2 g0976(.dina(new_n1039_), .dinb(new_n1040_), .dout(new_n1041_));
  anb1 g0977(.dina(new_n979_), .dinb(new_n1041_), .dout(new_n1042_));
  anb2 g0978(.dina(new_n979_), .dinb(new_n1041_), .dout(new_n1043_));
  nab1 g0979(.dina(new_n1042_), .dinb(new_n1043_), .dout(new_n1044_));
  anb2 g0980(.dina(new_n978_), .dinb(new_n1044_), .dout(new_n1045_));
  anb1 g0981(.dina(new_n978_), .dinb(new_n1044_), .dout(new_n1046_));
  nab2 g0982(.dina(new_n1045_), .dinb(new_n1046_), .dout(new_n1047_));
  anb1 g0983(.dina(new_n977_), .dinb(new_n1047_), .dout(new_n1048_));
  anb2 g0984(.dina(new_n977_), .dinb(new_n1047_), .dout(new_n1049_));
  nab1 g0985(.dina(new_n1048_), .dinb(new_n1049_), .dout(new_n1050_));
  anb2 g0986(.dina(new_n976_), .dinb(new_n1050_), .dout(new_n1051_));
  anb1 g0987(.dina(new_n976_), .dinb(new_n1050_), .dout(new_n1052_));
  nab2 g0988(.dina(new_n1051_), .dinb(new_n1052_), .dout(new_n1053_));
  anb1 g0989(.dina(new_n975_), .dinb(new_n1053_), .dout(new_n1054_));
  anb2 g0990(.dina(new_n975_), .dinb(new_n1053_), .dout(new_n1055_));
  nab1 g0991(.dina(new_n1054_), .dinb(new_n1055_), .dout(new_n1056_));
  anb2 g0992(.dina(new_n974_), .dinb(new_n1056_), .dout(new_n1057_));
  anb1 g0993(.dina(new_n974_), .dinb(new_n1056_), .dout(new_n1058_));
  anb1 g0994(.dina(new_n1057_), .dinb(new_n1058_), .dout(new_n1059_));
  anb2 g0995(.dina(new_n973_), .dinb(new_n1059_), .dout(new_n1060_));
  anb1 g0996(.dina(new_n973_), .dinb(new_n1059_), .dout(new_n1061_));
  anb1 g0997(.dina(new_n1060_), .dinb(new_n1061_), .dout(new_n1062_));
  anb2 g0998(.dina(new_n972_), .dinb(new_n1062_), .dout(new_n1063_));
  anb1 g0999(.dina(new_n972_), .dinb(new_n1062_), .dout(new_n1064_));
  anb1 g1000(.dina(new_n1063_), .dinb(new_n1064_), .dout(new_n1065_));
  anb2 g1001(.dina(new_n971_), .dinb(new_n1065_), .dout(new_n1066_));
  anb1 g1002(.dina(new_n971_), .dinb(new_n1065_), .dout(new_n1067_));
  anb1 g1003(.dina(new_n1066_), .dinb(new_n1067_), .dout(new_n1068_));
  anb2 g1004(.dina(new_n970_), .dinb(new_n1068_), .dout(new_n1069_));
  anb1 g1005(.dina(new_n970_), .dinb(new_n1068_), .dout(new_n1070_));
  anb1 g1006(.dina(new_n1069_), .dinb(new_n1070_), .dout(new_n1071_));
  anb2 g1007(.dina(new_n969_), .dinb(new_n1071_), .dout(new_n1072_));
  anb1 g1008(.dina(new_n969_), .dinb(new_n1071_), .dout(new_n1073_));
  anb1 g1009(.dina(new_n1072_), .dinb(new_n1073_), .dout(new_n1074_));
  anb2 g1010(.dina(new_n968_), .dinb(new_n1074_), .dout(new_n1075_));
  anb1 g1011(.dina(new_n968_), .dinb(new_n1074_), .dout(new_n1076_));
  anb1 g1012(.dina(new_n1075_), .dinb(new_n1076_), .dout(new_n1077_));
  anb2 g1013(.dina(new_n967_), .dinb(new_n1077_), .dout(new_n1078_));
  anb2 g1014(.dina(new_n1077_), .dinb(new_n967_), .dout(new_n1079_));
  and1 g1015(.dina(new_n1078_), .dinb(new_n1079_), .dout(G6273));
  nor2 g1016(.dina(new_n1072_), .dinb(new_n1075_), .dout(new_n1081_));
  nor2 g1017(.dina(G3), .dinb(G32), .dout(new_n1082_));
  nor2 g1018(.dina(new_n1066_), .dinb(new_n1069_), .dout(new_n1083_));
  nor2 g1019(.dina(G4), .dinb(G31), .dout(new_n1084_));
  nor2 g1020(.dina(new_n1060_), .dinb(new_n1063_), .dout(new_n1085_));
  nor2 g1021(.dina(G5), .dinb(G30), .dout(new_n1086_));
  anb2 g1022(.dina(new_n1054_), .dinb(new_n1057_), .dout(new_n1087_));
  and1 g1023(.dina(G6), .dinb(G29), .dout(new_n1088_));
  anb2 g1024(.dina(new_n1048_), .dinb(new_n1051_), .dout(new_n1089_));
  and1 g1025(.dina(G7), .dinb(G28), .dout(new_n1090_));
  anb2 g1026(.dina(new_n1042_), .dinb(new_n1045_), .dout(new_n1091_));
  and1 g1027(.dina(G8), .dinb(G27), .dout(new_n1092_));
  anb2 g1028(.dina(new_n1036_), .dinb(new_n1039_), .dout(new_n1093_));
  and1 g1029(.dina(G9), .dinb(G26), .dout(new_n1094_));
  anb2 g1030(.dina(new_n1030_), .dinb(new_n1033_), .dout(new_n1095_));
  and1 g1031(.dina(G10), .dinb(G25), .dout(new_n1096_));
  anb2 g1032(.dina(new_n1024_), .dinb(new_n1027_), .dout(new_n1097_));
  and1 g1033(.dina(G11), .dinb(G24), .dout(new_n1098_));
  anb2 g1034(.dina(new_n1018_), .dinb(new_n1021_), .dout(new_n1099_));
  and1 g1035(.dina(G12), .dinb(G23), .dout(new_n1100_));
  anb2 g1036(.dina(new_n1012_), .dinb(new_n1015_), .dout(new_n1101_));
  and1 g1037(.dina(G13), .dinb(G22), .dout(new_n1102_));
  anb2 g1038(.dina(new_n1006_), .dinb(new_n1009_), .dout(new_n1103_));
  and1 g1039(.dina(G14), .dinb(G21), .dout(new_n1104_));
  anb2 g1040(.dina(new_n1000_), .dinb(new_n1003_), .dout(new_n1105_));
  and1 g1041(.dina(G15), .dinb(G20), .dout(new_n1106_));
  nor2 g1042(.dina(G16), .dinb(G19), .dout(new_n1107_));
  anb1 g1043(.dina(new_n994_), .dinb(new_n997_), .dout(new_n1108_));
  anb1 g1044(.dina(new_n1107_), .dinb(new_n1108_), .dout(new_n1109_));
  anb2 g1045(.dina(new_n1107_), .dinb(new_n1108_), .dout(new_n1110_));
  nab1 g1046(.dina(new_n1109_), .dinb(new_n1110_), .dout(new_n1111_));
  anb2 g1047(.dina(new_n1106_), .dinb(new_n1111_), .dout(new_n1112_));
  anb1 g1048(.dina(new_n1106_), .dinb(new_n1111_), .dout(new_n1113_));
  nab2 g1049(.dina(new_n1112_), .dinb(new_n1113_), .dout(new_n1114_));
  anb1 g1050(.dina(new_n1105_), .dinb(new_n1114_), .dout(new_n1115_));
  anb2 g1051(.dina(new_n1105_), .dinb(new_n1114_), .dout(new_n1116_));
  nab1 g1052(.dina(new_n1115_), .dinb(new_n1116_), .dout(new_n1117_));
  anb2 g1053(.dina(new_n1104_), .dinb(new_n1117_), .dout(new_n1118_));
  anb1 g1054(.dina(new_n1104_), .dinb(new_n1117_), .dout(new_n1119_));
  nab2 g1055(.dina(new_n1118_), .dinb(new_n1119_), .dout(new_n1120_));
  anb1 g1056(.dina(new_n1103_), .dinb(new_n1120_), .dout(new_n1121_));
  anb2 g1057(.dina(new_n1103_), .dinb(new_n1120_), .dout(new_n1122_));
  nab1 g1058(.dina(new_n1121_), .dinb(new_n1122_), .dout(new_n1123_));
  anb2 g1059(.dina(new_n1102_), .dinb(new_n1123_), .dout(new_n1124_));
  anb1 g1060(.dina(new_n1102_), .dinb(new_n1123_), .dout(new_n1125_));
  nab2 g1061(.dina(new_n1124_), .dinb(new_n1125_), .dout(new_n1126_));
  anb1 g1062(.dina(new_n1101_), .dinb(new_n1126_), .dout(new_n1127_));
  anb2 g1063(.dina(new_n1101_), .dinb(new_n1126_), .dout(new_n1128_));
  nab1 g1064(.dina(new_n1127_), .dinb(new_n1128_), .dout(new_n1129_));
  anb2 g1065(.dina(new_n1100_), .dinb(new_n1129_), .dout(new_n1130_));
  anb1 g1066(.dina(new_n1100_), .dinb(new_n1129_), .dout(new_n1131_));
  nab2 g1067(.dina(new_n1130_), .dinb(new_n1131_), .dout(new_n1132_));
  anb1 g1068(.dina(new_n1099_), .dinb(new_n1132_), .dout(new_n1133_));
  anb2 g1069(.dina(new_n1099_), .dinb(new_n1132_), .dout(new_n1134_));
  nab1 g1070(.dina(new_n1133_), .dinb(new_n1134_), .dout(new_n1135_));
  anb2 g1071(.dina(new_n1098_), .dinb(new_n1135_), .dout(new_n1136_));
  anb1 g1072(.dina(new_n1098_), .dinb(new_n1135_), .dout(new_n1137_));
  nab2 g1073(.dina(new_n1136_), .dinb(new_n1137_), .dout(new_n1138_));
  anb1 g1074(.dina(new_n1097_), .dinb(new_n1138_), .dout(new_n1139_));
  anb2 g1075(.dina(new_n1097_), .dinb(new_n1138_), .dout(new_n1140_));
  nab1 g1076(.dina(new_n1139_), .dinb(new_n1140_), .dout(new_n1141_));
  anb2 g1077(.dina(new_n1096_), .dinb(new_n1141_), .dout(new_n1142_));
  anb1 g1078(.dina(new_n1096_), .dinb(new_n1141_), .dout(new_n1143_));
  nab2 g1079(.dina(new_n1142_), .dinb(new_n1143_), .dout(new_n1144_));
  anb1 g1080(.dina(new_n1095_), .dinb(new_n1144_), .dout(new_n1145_));
  anb2 g1081(.dina(new_n1095_), .dinb(new_n1144_), .dout(new_n1146_));
  nab1 g1082(.dina(new_n1145_), .dinb(new_n1146_), .dout(new_n1147_));
  anb2 g1083(.dina(new_n1094_), .dinb(new_n1147_), .dout(new_n1148_));
  anb1 g1084(.dina(new_n1094_), .dinb(new_n1147_), .dout(new_n1149_));
  nab2 g1085(.dina(new_n1148_), .dinb(new_n1149_), .dout(new_n1150_));
  anb1 g1086(.dina(new_n1093_), .dinb(new_n1150_), .dout(new_n1151_));
  anb2 g1087(.dina(new_n1093_), .dinb(new_n1150_), .dout(new_n1152_));
  nab1 g1088(.dina(new_n1151_), .dinb(new_n1152_), .dout(new_n1153_));
  anb2 g1089(.dina(new_n1092_), .dinb(new_n1153_), .dout(new_n1154_));
  anb1 g1090(.dina(new_n1092_), .dinb(new_n1153_), .dout(new_n1155_));
  nab2 g1091(.dina(new_n1154_), .dinb(new_n1155_), .dout(new_n1156_));
  anb1 g1092(.dina(new_n1091_), .dinb(new_n1156_), .dout(new_n1157_));
  anb2 g1093(.dina(new_n1091_), .dinb(new_n1156_), .dout(new_n1158_));
  nab1 g1094(.dina(new_n1157_), .dinb(new_n1158_), .dout(new_n1159_));
  anb2 g1095(.dina(new_n1090_), .dinb(new_n1159_), .dout(new_n1160_));
  anb1 g1096(.dina(new_n1090_), .dinb(new_n1159_), .dout(new_n1161_));
  nab2 g1097(.dina(new_n1160_), .dinb(new_n1161_), .dout(new_n1162_));
  anb1 g1098(.dina(new_n1089_), .dinb(new_n1162_), .dout(new_n1163_));
  anb2 g1099(.dina(new_n1089_), .dinb(new_n1162_), .dout(new_n1164_));
  nab1 g1100(.dina(new_n1163_), .dinb(new_n1164_), .dout(new_n1165_));
  anb2 g1101(.dina(new_n1088_), .dinb(new_n1165_), .dout(new_n1166_));
  anb1 g1102(.dina(new_n1088_), .dinb(new_n1165_), .dout(new_n1167_));
  nab2 g1103(.dina(new_n1166_), .dinb(new_n1167_), .dout(new_n1168_));
  anb1 g1104(.dina(new_n1087_), .dinb(new_n1168_), .dout(new_n1169_));
  anb2 g1105(.dina(new_n1087_), .dinb(new_n1168_), .dout(new_n1170_));
  anb2 g1106(.dina(new_n1169_), .dinb(new_n1170_), .dout(new_n1171_));
  anb1 g1107(.dina(new_n1086_), .dinb(new_n1171_), .dout(new_n1172_));
  anb2 g1108(.dina(new_n1086_), .dinb(new_n1171_), .dout(new_n1173_));
  anb2 g1109(.dina(new_n1172_), .dinb(new_n1173_), .dout(new_n1174_));
  anb1 g1110(.dina(new_n1085_), .dinb(new_n1174_), .dout(new_n1175_));
  anb2 g1111(.dina(new_n1085_), .dinb(new_n1174_), .dout(new_n1176_));
  anb2 g1112(.dina(new_n1175_), .dinb(new_n1176_), .dout(new_n1177_));
  anb1 g1113(.dina(new_n1084_), .dinb(new_n1177_), .dout(new_n1178_));
  anb2 g1114(.dina(new_n1084_), .dinb(new_n1177_), .dout(new_n1179_));
  anb2 g1115(.dina(new_n1178_), .dinb(new_n1179_), .dout(new_n1180_));
  anb1 g1116(.dina(new_n1083_), .dinb(new_n1180_), .dout(new_n1181_));
  anb2 g1117(.dina(new_n1083_), .dinb(new_n1180_), .dout(new_n1182_));
  anb2 g1118(.dina(new_n1181_), .dinb(new_n1182_), .dout(new_n1183_));
  anb1 g1119(.dina(new_n1082_), .dinb(new_n1183_), .dout(new_n1184_));
  anb2 g1120(.dina(new_n1082_), .dinb(new_n1183_), .dout(new_n1185_));
  anb2 g1121(.dina(new_n1184_), .dinb(new_n1185_), .dout(new_n1186_));
  anb1 g1122(.dina(new_n1081_), .dinb(new_n1186_), .dout(new_n1187_));
  anb2 g1123(.dina(new_n1081_), .dinb(new_n1186_), .dout(new_n1188_));
  anb2 g1124(.dina(new_n1187_), .dinb(new_n1188_), .dout(new_n1189_));
  anb1 g1125(.dina(new_n1079_), .dinb(new_n1189_), .dout(new_n1190_));
  anb2 g1126(.dina(new_n1079_), .dinb(new_n1189_), .dout(new_n1191_));
  anb2 g1127(.dina(new_n1190_), .dinb(new_n1191_), .dout(G6274));
  and2 g1128(.dina(new_n1187_), .dinb(new_n1190_), .dout(new_n1193_));
  and2 g1129(.dina(new_n1181_), .dinb(new_n1184_), .dout(new_n1194_));
  nor2 g1130(.dina(G4), .dinb(G32), .dout(new_n1195_));
  and2 g1131(.dina(new_n1175_), .dinb(new_n1178_), .dout(new_n1196_));
  nor2 g1132(.dina(G5), .dinb(G31), .dout(new_n1197_));
  and2 g1133(.dina(new_n1169_), .dinb(new_n1172_), .dout(new_n1198_));
  nor2 g1134(.dina(G6), .dinb(G30), .dout(new_n1199_));
  anb2 g1135(.dina(new_n1163_), .dinb(new_n1166_), .dout(new_n1200_));
  and1 g1136(.dina(G7), .dinb(G29), .dout(new_n1201_));
  anb2 g1137(.dina(new_n1157_), .dinb(new_n1160_), .dout(new_n1202_));
  and1 g1138(.dina(G8), .dinb(G28), .dout(new_n1203_));
  anb2 g1139(.dina(new_n1151_), .dinb(new_n1154_), .dout(new_n1204_));
  and1 g1140(.dina(G9), .dinb(G27), .dout(new_n1205_));
  anb2 g1141(.dina(new_n1145_), .dinb(new_n1148_), .dout(new_n1206_));
  and1 g1142(.dina(G10), .dinb(G26), .dout(new_n1207_));
  anb2 g1143(.dina(new_n1139_), .dinb(new_n1142_), .dout(new_n1208_));
  and1 g1144(.dina(G11), .dinb(G25), .dout(new_n1209_));
  anb2 g1145(.dina(new_n1133_), .dinb(new_n1136_), .dout(new_n1210_));
  and1 g1146(.dina(G12), .dinb(G24), .dout(new_n1211_));
  anb2 g1147(.dina(new_n1127_), .dinb(new_n1130_), .dout(new_n1212_));
  and1 g1148(.dina(G13), .dinb(G23), .dout(new_n1213_));
  anb2 g1149(.dina(new_n1121_), .dinb(new_n1124_), .dout(new_n1214_));
  and1 g1150(.dina(G14), .dinb(G22), .dout(new_n1215_));
  anb2 g1151(.dina(new_n1115_), .dinb(new_n1118_), .dout(new_n1216_));
  nor2 g1152(.dina(G15), .dinb(G21), .dout(new_n1217_));
  and1 g1153(.dina(G16), .dinb(G20), .dout(new_n1218_));
  anb2 g1154(.dina(new_n1109_), .dinb(new_n1112_), .dout(new_n1219_));
  anb2 g1155(.dina(new_n1218_), .dinb(new_n1219_), .dout(new_n1220_));
  anb1 g1156(.dina(new_n1218_), .dinb(new_n1219_), .dout(new_n1221_));
  nab2 g1157(.dina(new_n1220_), .dinb(new_n1221_), .dout(new_n1222_));
  anb1 g1158(.dina(new_n1217_), .dinb(new_n1222_), .dout(new_n1223_));
  anb2 g1159(.dina(new_n1217_), .dinb(new_n1222_), .dout(new_n1224_));
  anb2 g1160(.dina(new_n1223_), .dinb(new_n1224_), .dout(new_n1225_));
  anb1 g1161(.dina(new_n1216_), .dinb(new_n1225_), .dout(new_n1226_));
  anb2 g1162(.dina(new_n1216_), .dinb(new_n1225_), .dout(new_n1227_));
  nab1 g1163(.dina(new_n1226_), .dinb(new_n1227_), .dout(new_n1228_));
  anb2 g1164(.dina(new_n1215_), .dinb(new_n1228_), .dout(new_n1229_));
  anb1 g1165(.dina(new_n1215_), .dinb(new_n1228_), .dout(new_n1230_));
  nab2 g1166(.dina(new_n1229_), .dinb(new_n1230_), .dout(new_n1231_));
  anb1 g1167(.dina(new_n1214_), .dinb(new_n1231_), .dout(new_n1232_));
  anb2 g1168(.dina(new_n1214_), .dinb(new_n1231_), .dout(new_n1233_));
  nab1 g1169(.dina(new_n1232_), .dinb(new_n1233_), .dout(new_n1234_));
  anb2 g1170(.dina(new_n1213_), .dinb(new_n1234_), .dout(new_n1235_));
  anb1 g1171(.dina(new_n1213_), .dinb(new_n1234_), .dout(new_n1236_));
  nab2 g1172(.dina(new_n1235_), .dinb(new_n1236_), .dout(new_n1237_));
  anb1 g1173(.dina(new_n1212_), .dinb(new_n1237_), .dout(new_n1238_));
  anb2 g1174(.dina(new_n1212_), .dinb(new_n1237_), .dout(new_n1239_));
  nab1 g1175(.dina(new_n1238_), .dinb(new_n1239_), .dout(new_n1240_));
  anb2 g1176(.dina(new_n1211_), .dinb(new_n1240_), .dout(new_n1241_));
  anb1 g1177(.dina(new_n1211_), .dinb(new_n1240_), .dout(new_n1242_));
  nab2 g1178(.dina(new_n1241_), .dinb(new_n1242_), .dout(new_n1243_));
  anb1 g1179(.dina(new_n1210_), .dinb(new_n1243_), .dout(new_n1244_));
  anb2 g1180(.dina(new_n1210_), .dinb(new_n1243_), .dout(new_n1245_));
  nab1 g1181(.dina(new_n1244_), .dinb(new_n1245_), .dout(new_n1246_));
  anb2 g1182(.dina(new_n1209_), .dinb(new_n1246_), .dout(new_n1247_));
  anb1 g1183(.dina(new_n1209_), .dinb(new_n1246_), .dout(new_n1248_));
  nab2 g1184(.dina(new_n1247_), .dinb(new_n1248_), .dout(new_n1249_));
  anb1 g1185(.dina(new_n1208_), .dinb(new_n1249_), .dout(new_n1250_));
  anb2 g1186(.dina(new_n1208_), .dinb(new_n1249_), .dout(new_n1251_));
  nab1 g1187(.dina(new_n1250_), .dinb(new_n1251_), .dout(new_n1252_));
  anb2 g1188(.dina(new_n1207_), .dinb(new_n1252_), .dout(new_n1253_));
  anb1 g1189(.dina(new_n1207_), .dinb(new_n1252_), .dout(new_n1254_));
  nab2 g1190(.dina(new_n1253_), .dinb(new_n1254_), .dout(new_n1255_));
  anb1 g1191(.dina(new_n1206_), .dinb(new_n1255_), .dout(new_n1256_));
  anb2 g1192(.dina(new_n1206_), .dinb(new_n1255_), .dout(new_n1257_));
  nab1 g1193(.dina(new_n1256_), .dinb(new_n1257_), .dout(new_n1258_));
  anb2 g1194(.dina(new_n1205_), .dinb(new_n1258_), .dout(new_n1259_));
  anb1 g1195(.dina(new_n1205_), .dinb(new_n1258_), .dout(new_n1260_));
  nab2 g1196(.dina(new_n1259_), .dinb(new_n1260_), .dout(new_n1261_));
  anb1 g1197(.dina(new_n1204_), .dinb(new_n1261_), .dout(new_n1262_));
  anb2 g1198(.dina(new_n1204_), .dinb(new_n1261_), .dout(new_n1263_));
  nab1 g1199(.dina(new_n1262_), .dinb(new_n1263_), .dout(new_n1264_));
  anb2 g1200(.dina(new_n1203_), .dinb(new_n1264_), .dout(new_n1265_));
  anb1 g1201(.dina(new_n1203_), .dinb(new_n1264_), .dout(new_n1266_));
  nab2 g1202(.dina(new_n1265_), .dinb(new_n1266_), .dout(new_n1267_));
  anb1 g1203(.dina(new_n1202_), .dinb(new_n1267_), .dout(new_n1268_));
  anb2 g1204(.dina(new_n1202_), .dinb(new_n1267_), .dout(new_n1269_));
  nab1 g1205(.dina(new_n1268_), .dinb(new_n1269_), .dout(new_n1270_));
  anb2 g1206(.dina(new_n1201_), .dinb(new_n1270_), .dout(new_n1271_));
  anb1 g1207(.dina(new_n1201_), .dinb(new_n1270_), .dout(new_n1272_));
  nab2 g1208(.dina(new_n1271_), .dinb(new_n1272_), .dout(new_n1273_));
  anb1 g1209(.dina(new_n1200_), .dinb(new_n1273_), .dout(new_n1274_));
  anb2 g1210(.dina(new_n1200_), .dinb(new_n1273_), .dout(new_n1275_));
  anb2 g1211(.dina(new_n1274_), .dinb(new_n1275_), .dout(new_n1276_));
  anb1 g1212(.dina(new_n1199_), .dinb(new_n1276_), .dout(new_n1277_));
  anb2 g1213(.dina(new_n1199_), .dinb(new_n1276_), .dout(new_n1278_));
  anb2 g1214(.dina(new_n1277_), .dinb(new_n1278_), .dout(new_n1279_));
  anb1 g1215(.dina(new_n1198_), .dinb(new_n1279_), .dout(new_n1280_));
  anb2 g1216(.dina(new_n1198_), .dinb(new_n1279_), .dout(new_n1281_));
  anb2 g1217(.dina(new_n1280_), .dinb(new_n1281_), .dout(new_n1282_));
  anb1 g1218(.dina(new_n1197_), .dinb(new_n1282_), .dout(new_n1283_));
  anb2 g1219(.dina(new_n1197_), .dinb(new_n1282_), .dout(new_n1284_));
  anb2 g1220(.dina(new_n1283_), .dinb(new_n1284_), .dout(new_n1285_));
  anb1 g1221(.dina(new_n1196_), .dinb(new_n1285_), .dout(new_n1286_));
  anb2 g1222(.dina(new_n1196_), .dinb(new_n1285_), .dout(new_n1287_));
  anb2 g1223(.dina(new_n1286_), .dinb(new_n1287_), .dout(new_n1288_));
  anb1 g1224(.dina(new_n1195_), .dinb(new_n1288_), .dout(new_n1289_));
  anb2 g1225(.dina(new_n1195_), .dinb(new_n1288_), .dout(new_n1290_));
  anb2 g1226(.dina(new_n1289_), .dinb(new_n1290_), .dout(new_n1291_));
  anb1 g1227(.dina(new_n1194_), .dinb(new_n1291_), .dout(new_n1292_));
  anb2 g1228(.dina(new_n1194_), .dinb(new_n1291_), .dout(new_n1293_));
  anb2 g1229(.dina(new_n1292_), .dinb(new_n1293_), .dout(new_n1294_));
  anb1 g1230(.dina(new_n1193_), .dinb(new_n1294_), .dout(new_n1295_));
  anb2 g1231(.dina(new_n1193_), .dinb(new_n1294_), .dout(new_n1296_));
  anb2 g1232(.dina(new_n1295_), .dinb(new_n1296_), .dout(G6275));
  and2 g1233(.dina(new_n1292_), .dinb(new_n1295_), .dout(new_n1298_));
  and2 g1234(.dina(new_n1286_), .dinb(new_n1289_), .dout(new_n1299_));
  nor2 g1235(.dina(G5), .dinb(G32), .dout(new_n1300_));
  and2 g1236(.dina(new_n1280_), .dinb(new_n1283_), .dout(new_n1301_));
  nor2 g1237(.dina(G6), .dinb(G31), .dout(new_n1302_));
  and2 g1238(.dina(new_n1274_), .dinb(new_n1277_), .dout(new_n1303_));
  nor2 g1239(.dina(G7), .dinb(G30), .dout(new_n1304_));
  anb2 g1240(.dina(new_n1268_), .dinb(new_n1271_), .dout(new_n1305_));
  and1 g1241(.dina(G8), .dinb(G29), .dout(new_n1306_));
  anb2 g1242(.dina(new_n1262_), .dinb(new_n1265_), .dout(new_n1307_));
  and1 g1243(.dina(G9), .dinb(G28), .dout(new_n1308_));
  anb2 g1244(.dina(new_n1256_), .dinb(new_n1259_), .dout(new_n1309_));
  and1 g1245(.dina(G10), .dinb(G27), .dout(new_n1310_));
  anb2 g1246(.dina(new_n1250_), .dinb(new_n1253_), .dout(new_n1311_));
  and1 g1247(.dina(G11), .dinb(G26), .dout(new_n1312_));
  anb2 g1248(.dina(new_n1244_), .dinb(new_n1247_), .dout(new_n1313_));
  and1 g1249(.dina(G12), .dinb(G25), .dout(new_n1314_));
  anb2 g1250(.dina(new_n1238_), .dinb(new_n1241_), .dout(new_n1315_));
  and1 g1251(.dina(G13), .dinb(G24), .dout(new_n1316_));
  anb2 g1252(.dina(new_n1232_), .dinb(new_n1235_), .dout(new_n1317_));
  and1 g1253(.dina(G14), .dinb(G23), .dout(new_n1318_));
  anb2 g1254(.dina(new_n1226_), .dinb(new_n1229_), .dout(new_n1319_));
  and1 g1255(.dina(G15), .dinb(G22), .dout(new_n1320_));
  nor2 g1256(.dina(G16), .dinb(G21), .dout(new_n1321_));
  anb1 g1257(.dina(new_n1220_), .dinb(new_n1223_), .dout(new_n1322_));
  anb1 g1258(.dina(new_n1321_), .dinb(new_n1322_), .dout(new_n1323_));
  anb2 g1259(.dina(new_n1321_), .dinb(new_n1322_), .dout(new_n1324_));
  nab1 g1260(.dina(new_n1323_), .dinb(new_n1324_), .dout(new_n1325_));
  anb2 g1261(.dina(new_n1320_), .dinb(new_n1325_), .dout(new_n1326_));
  anb1 g1262(.dina(new_n1320_), .dinb(new_n1325_), .dout(new_n1327_));
  nab2 g1263(.dina(new_n1326_), .dinb(new_n1327_), .dout(new_n1328_));
  anb1 g1264(.dina(new_n1319_), .dinb(new_n1328_), .dout(new_n1329_));
  anb2 g1265(.dina(new_n1319_), .dinb(new_n1328_), .dout(new_n1330_));
  nab1 g1266(.dina(new_n1329_), .dinb(new_n1330_), .dout(new_n1331_));
  anb2 g1267(.dina(new_n1318_), .dinb(new_n1331_), .dout(new_n1332_));
  anb1 g1268(.dina(new_n1318_), .dinb(new_n1331_), .dout(new_n1333_));
  nab2 g1269(.dina(new_n1332_), .dinb(new_n1333_), .dout(new_n1334_));
  anb1 g1270(.dina(new_n1317_), .dinb(new_n1334_), .dout(new_n1335_));
  anb2 g1271(.dina(new_n1317_), .dinb(new_n1334_), .dout(new_n1336_));
  nab1 g1272(.dina(new_n1335_), .dinb(new_n1336_), .dout(new_n1337_));
  anb2 g1273(.dina(new_n1316_), .dinb(new_n1337_), .dout(new_n1338_));
  anb1 g1274(.dina(new_n1316_), .dinb(new_n1337_), .dout(new_n1339_));
  nab2 g1275(.dina(new_n1338_), .dinb(new_n1339_), .dout(new_n1340_));
  anb1 g1276(.dina(new_n1315_), .dinb(new_n1340_), .dout(new_n1341_));
  anb2 g1277(.dina(new_n1315_), .dinb(new_n1340_), .dout(new_n1342_));
  nab1 g1278(.dina(new_n1341_), .dinb(new_n1342_), .dout(new_n1343_));
  anb2 g1279(.dina(new_n1314_), .dinb(new_n1343_), .dout(new_n1344_));
  anb1 g1280(.dina(new_n1314_), .dinb(new_n1343_), .dout(new_n1345_));
  nab2 g1281(.dina(new_n1344_), .dinb(new_n1345_), .dout(new_n1346_));
  anb1 g1282(.dina(new_n1313_), .dinb(new_n1346_), .dout(new_n1347_));
  anb2 g1283(.dina(new_n1313_), .dinb(new_n1346_), .dout(new_n1348_));
  nab1 g1284(.dina(new_n1347_), .dinb(new_n1348_), .dout(new_n1349_));
  anb2 g1285(.dina(new_n1312_), .dinb(new_n1349_), .dout(new_n1350_));
  anb1 g1286(.dina(new_n1312_), .dinb(new_n1349_), .dout(new_n1351_));
  nab2 g1287(.dina(new_n1350_), .dinb(new_n1351_), .dout(new_n1352_));
  anb1 g1288(.dina(new_n1311_), .dinb(new_n1352_), .dout(new_n1353_));
  anb2 g1289(.dina(new_n1311_), .dinb(new_n1352_), .dout(new_n1354_));
  nab1 g1290(.dina(new_n1353_), .dinb(new_n1354_), .dout(new_n1355_));
  anb2 g1291(.dina(new_n1310_), .dinb(new_n1355_), .dout(new_n1356_));
  anb1 g1292(.dina(new_n1310_), .dinb(new_n1355_), .dout(new_n1357_));
  nab2 g1293(.dina(new_n1356_), .dinb(new_n1357_), .dout(new_n1358_));
  anb1 g1294(.dina(new_n1309_), .dinb(new_n1358_), .dout(new_n1359_));
  anb2 g1295(.dina(new_n1309_), .dinb(new_n1358_), .dout(new_n1360_));
  nab1 g1296(.dina(new_n1359_), .dinb(new_n1360_), .dout(new_n1361_));
  anb2 g1297(.dina(new_n1308_), .dinb(new_n1361_), .dout(new_n1362_));
  anb1 g1298(.dina(new_n1308_), .dinb(new_n1361_), .dout(new_n1363_));
  nab2 g1299(.dina(new_n1362_), .dinb(new_n1363_), .dout(new_n1364_));
  anb1 g1300(.dina(new_n1307_), .dinb(new_n1364_), .dout(new_n1365_));
  anb2 g1301(.dina(new_n1307_), .dinb(new_n1364_), .dout(new_n1366_));
  nab1 g1302(.dina(new_n1365_), .dinb(new_n1366_), .dout(new_n1367_));
  anb2 g1303(.dina(new_n1306_), .dinb(new_n1367_), .dout(new_n1368_));
  anb1 g1304(.dina(new_n1306_), .dinb(new_n1367_), .dout(new_n1369_));
  nab2 g1305(.dina(new_n1368_), .dinb(new_n1369_), .dout(new_n1370_));
  anb1 g1306(.dina(new_n1305_), .dinb(new_n1370_), .dout(new_n1371_));
  anb2 g1307(.dina(new_n1305_), .dinb(new_n1370_), .dout(new_n1372_));
  anb2 g1308(.dina(new_n1371_), .dinb(new_n1372_), .dout(new_n1373_));
  anb1 g1309(.dina(new_n1304_), .dinb(new_n1373_), .dout(new_n1374_));
  anb2 g1310(.dina(new_n1304_), .dinb(new_n1373_), .dout(new_n1375_));
  anb2 g1311(.dina(new_n1374_), .dinb(new_n1375_), .dout(new_n1376_));
  anb1 g1312(.dina(new_n1303_), .dinb(new_n1376_), .dout(new_n1377_));
  anb2 g1313(.dina(new_n1303_), .dinb(new_n1376_), .dout(new_n1378_));
  anb2 g1314(.dina(new_n1377_), .dinb(new_n1378_), .dout(new_n1379_));
  anb1 g1315(.dina(new_n1302_), .dinb(new_n1379_), .dout(new_n1380_));
  anb2 g1316(.dina(new_n1302_), .dinb(new_n1379_), .dout(new_n1381_));
  anb2 g1317(.dina(new_n1380_), .dinb(new_n1381_), .dout(new_n1382_));
  anb1 g1318(.dina(new_n1301_), .dinb(new_n1382_), .dout(new_n1383_));
  anb2 g1319(.dina(new_n1301_), .dinb(new_n1382_), .dout(new_n1384_));
  anb2 g1320(.dina(new_n1383_), .dinb(new_n1384_), .dout(new_n1385_));
  anb1 g1321(.dina(new_n1300_), .dinb(new_n1385_), .dout(new_n1386_));
  anb2 g1322(.dina(new_n1300_), .dinb(new_n1385_), .dout(new_n1387_));
  anb2 g1323(.dina(new_n1386_), .dinb(new_n1387_), .dout(new_n1388_));
  anb1 g1324(.dina(new_n1299_), .dinb(new_n1388_), .dout(new_n1389_));
  anb2 g1325(.dina(new_n1299_), .dinb(new_n1388_), .dout(new_n1390_));
  anb2 g1326(.dina(new_n1389_), .dinb(new_n1390_), .dout(new_n1391_));
  anb1 g1327(.dina(new_n1298_), .dinb(new_n1391_), .dout(new_n1392_));
  anb2 g1328(.dina(new_n1298_), .dinb(new_n1391_), .dout(new_n1393_));
  anb2 g1329(.dina(new_n1392_), .dinb(new_n1393_), .dout(G6276));
  and2 g1330(.dina(new_n1389_), .dinb(new_n1392_), .dout(new_n1395_));
  and2 g1331(.dina(new_n1383_), .dinb(new_n1386_), .dout(new_n1396_));
  nor2 g1332(.dina(G6), .dinb(G32), .dout(new_n1397_));
  and2 g1333(.dina(new_n1377_), .dinb(new_n1380_), .dout(new_n1398_));
  nor2 g1334(.dina(G7), .dinb(G31), .dout(new_n1399_));
  and2 g1335(.dina(new_n1371_), .dinb(new_n1374_), .dout(new_n1400_));
  nor2 g1336(.dina(G8), .dinb(G30), .dout(new_n1401_));
  anb2 g1337(.dina(new_n1365_), .dinb(new_n1368_), .dout(new_n1402_));
  and1 g1338(.dina(G9), .dinb(G29), .dout(new_n1403_));
  anb2 g1339(.dina(new_n1359_), .dinb(new_n1362_), .dout(new_n1404_));
  and1 g1340(.dina(G10), .dinb(G28), .dout(new_n1405_));
  anb2 g1341(.dina(new_n1353_), .dinb(new_n1356_), .dout(new_n1406_));
  and1 g1342(.dina(G11), .dinb(G27), .dout(new_n1407_));
  anb2 g1343(.dina(new_n1347_), .dinb(new_n1350_), .dout(new_n1408_));
  and1 g1344(.dina(G12), .dinb(G26), .dout(new_n1409_));
  anb2 g1345(.dina(new_n1341_), .dinb(new_n1344_), .dout(new_n1410_));
  and1 g1346(.dina(G13), .dinb(G25), .dout(new_n1411_));
  anb2 g1347(.dina(new_n1335_), .dinb(new_n1338_), .dout(new_n1412_));
  and1 g1348(.dina(G14), .dinb(G24), .dout(new_n1413_));
  anb2 g1349(.dina(new_n1329_), .dinb(new_n1332_), .dout(new_n1414_));
  nor2 g1350(.dina(G15), .dinb(G23), .dout(new_n1415_));
  and1 g1351(.dina(G16), .dinb(G22), .dout(new_n1416_));
  anb2 g1352(.dina(new_n1323_), .dinb(new_n1326_), .dout(new_n1417_));
  anb2 g1353(.dina(new_n1416_), .dinb(new_n1417_), .dout(new_n1418_));
  anb1 g1354(.dina(new_n1416_), .dinb(new_n1417_), .dout(new_n1419_));
  nab2 g1355(.dina(new_n1418_), .dinb(new_n1419_), .dout(new_n1420_));
  anb1 g1356(.dina(new_n1415_), .dinb(new_n1420_), .dout(new_n1421_));
  anb2 g1357(.dina(new_n1415_), .dinb(new_n1420_), .dout(new_n1422_));
  anb2 g1358(.dina(new_n1421_), .dinb(new_n1422_), .dout(new_n1423_));
  anb1 g1359(.dina(new_n1414_), .dinb(new_n1423_), .dout(new_n1424_));
  anb2 g1360(.dina(new_n1414_), .dinb(new_n1423_), .dout(new_n1425_));
  nab1 g1361(.dina(new_n1424_), .dinb(new_n1425_), .dout(new_n1426_));
  anb2 g1362(.dina(new_n1413_), .dinb(new_n1426_), .dout(new_n1427_));
  anb1 g1363(.dina(new_n1413_), .dinb(new_n1426_), .dout(new_n1428_));
  nab2 g1364(.dina(new_n1427_), .dinb(new_n1428_), .dout(new_n1429_));
  anb1 g1365(.dina(new_n1412_), .dinb(new_n1429_), .dout(new_n1430_));
  anb2 g1366(.dina(new_n1412_), .dinb(new_n1429_), .dout(new_n1431_));
  nab1 g1367(.dina(new_n1430_), .dinb(new_n1431_), .dout(new_n1432_));
  anb2 g1368(.dina(new_n1411_), .dinb(new_n1432_), .dout(new_n1433_));
  anb1 g1369(.dina(new_n1411_), .dinb(new_n1432_), .dout(new_n1434_));
  nab2 g1370(.dina(new_n1433_), .dinb(new_n1434_), .dout(new_n1435_));
  anb1 g1371(.dina(new_n1410_), .dinb(new_n1435_), .dout(new_n1436_));
  anb2 g1372(.dina(new_n1410_), .dinb(new_n1435_), .dout(new_n1437_));
  nab1 g1373(.dina(new_n1436_), .dinb(new_n1437_), .dout(new_n1438_));
  anb2 g1374(.dina(new_n1409_), .dinb(new_n1438_), .dout(new_n1439_));
  anb1 g1375(.dina(new_n1409_), .dinb(new_n1438_), .dout(new_n1440_));
  nab2 g1376(.dina(new_n1439_), .dinb(new_n1440_), .dout(new_n1441_));
  anb1 g1377(.dina(new_n1408_), .dinb(new_n1441_), .dout(new_n1442_));
  anb2 g1378(.dina(new_n1408_), .dinb(new_n1441_), .dout(new_n1443_));
  nab1 g1379(.dina(new_n1442_), .dinb(new_n1443_), .dout(new_n1444_));
  anb2 g1380(.dina(new_n1407_), .dinb(new_n1444_), .dout(new_n1445_));
  anb1 g1381(.dina(new_n1407_), .dinb(new_n1444_), .dout(new_n1446_));
  nab2 g1382(.dina(new_n1445_), .dinb(new_n1446_), .dout(new_n1447_));
  anb1 g1383(.dina(new_n1406_), .dinb(new_n1447_), .dout(new_n1448_));
  anb2 g1384(.dina(new_n1406_), .dinb(new_n1447_), .dout(new_n1449_));
  nab1 g1385(.dina(new_n1448_), .dinb(new_n1449_), .dout(new_n1450_));
  anb2 g1386(.dina(new_n1405_), .dinb(new_n1450_), .dout(new_n1451_));
  anb1 g1387(.dina(new_n1405_), .dinb(new_n1450_), .dout(new_n1452_));
  nab2 g1388(.dina(new_n1451_), .dinb(new_n1452_), .dout(new_n1453_));
  anb1 g1389(.dina(new_n1404_), .dinb(new_n1453_), .dout(new_n1454_));
  anb2 g1390(.dina(new_n1404_), .dinb(new_n1453_), .dout(new_n1455_));
  nab1 g1391(.dina(new_n1454_), .dinb(new_n1455_), .dout(new_n1456_));
  anb2 g1392(.dina(new_n1403_), .dinb(new_n1456_), .dout(new_n1457_));
  anb1 g1393(.dina(new_n1403_), .dinb(new_n1456_), .dout(new_n1458_));
  nab2 g1394(.dina(new_n1457_), .dinb(new_n1458_), .dout(new_n1459_));
  anb1 g1395(.dina(new_n1402_), .dinb(new_n1459_), .dout(new_n1460_));
  anb2 g1396(.dina(new_n1402_), .dinb(new_n1459_), .dout(new_n1461_));
  anb2 g1397(.dina(new_n1460_), .dinb(new_n1461_), .dout(new_n1462_));
  anb1 g1398(.dina(new_n1401_), .dinb(new_n1462_), .dout(new_n1463_));
  anb2 g1399(.dina(new_n1401_), .dinb(new_n1462_), .dout(new_n1464_));
  anb2 g1400(.dina(new_n1463_), .dinb(new_n1464_), .dout(new_n1465_));
  anb1 g1401(.dina(new_n1400_), .dinb(new_n1465_), .dout(new_n1466_));
  anb2 g1402(.dina(new_n1400_), .dinb(new_n1465_), .dout(new_n1467_));
  anb2 g1403(.dina(new_n1466_), .dinb(new_n1467_), .dout(new_n1468_));
  anb1 g1404(.dina(new_n1399_), .dinb(new_n1468_), .dout(new_n1469_));
  anb2 g1405(.dina(new_n1399_), .dinb(new_n1468_), .dout(new_n1470_));
  anb2 g1406(.dina(new_n1469_), .dinb(new_n1470_), .dout(new_n1471_));
  anb1 g1407(.dina(new_n1398_), .dinb(new_n1471_), .dout(new_n1472_));
  anb2 g1408(.dina(new_n1398_), .dinb(new_n1471_), .dout(new_n1473_));
  anb2 g1409(.dina(new_n1472_), .dinb(new_n1473_), .dout(new_n1474_));
  anb1 g1410(.dina(new_n1397_), .dinb(new_n1474_), .dout(new_n1475_));
  anb2 g1411(.dina(new_n1397_), .dinb(new_n1474_), .dout(new_n1476_));
  anb2 g1412(.dina(new_n1475_), .dinb(new_n1476_), .dout(new_n1477_));
  anb1 g1413(.dina(new_n1396_), .dinb(new_n1477_), .dout(new_n1478_));
  anb2 g1414(.dina(new_n1396_), .dinb(new_n1477_), .dout(new_n1479_));
  anb2 g1415(.dina(new_n1478_), .dinb(new_n1479_), .dout(new_n1480_));
  anb1 g1416(.dina(new_n1395_), .dinb(new_n1480_), .dout(new_n1481_));
  anb2 g1417(.dina(new_n1395_), .dinb(new_n1480_), .dout(new_n1482_));
  anb2 g1418(.dina(new_n1481_), .dinb(new_n1482_), .dout(G6277));
  and2 g1419(.dina(new_n1478_), .dinb(new_n1481_), .dout(new_n1484_));
  and2 g1420(.dina(new_n1472_), .dinb(new_n1475_), .dout(new_n1485_));
  nor2 g1421(.dina(G7), .dinb(G32), .dout(new_n1486_));
  and2 g1422(.dina(new_n1466_), .dinb(new_n1469_), .dout(new_n1487_));
  nor2 g1423(.dina(G8), .dinb(G31), .dout(new_n1488_));
  and2 g1424(.dina(new_n1460_), .dinb(new_n1463_), .dout(new_n1489_));
  nor2 g1425(.dina(G9), .dinb(G30), .dout(new_n1490_));
  anb2 g1426(.dina(new_n1454_), .dinb(new_n1457_), .dout(new_n1491_));
  and1 g1427(.dina(G10), .dinb(G29), .dout(new_n1492_));
  anb2 g1428(.dina(new_n1448_), .dinb(new_n1451_), .dout(new_n1493_));
  and1 g1429(.dina(G11), .dinb(G28), .dout(new_n1494_));
  anb2 g1430(.dina(new_n1442_), .dinb(new_n1445_), .dout(new_n1495_));
  and1 g1431(.dina(G12), .dinb(G27), .dout(new_n1496_));
  anb2 g1432(.dina(new_n1436_), .dinb(new_n1439_), .dout(new_n1497_));
  and1 g1433(.dina(G13), .dinb(G26), .dout(new_n1498_));
  anb2 g1434(.dina(new_n1430_), .dinb(new_n1433_), .dout(new_n1499_));
  and1 g1435(.dina(G14), .dinb(G25), .dout(new_n1500_));
  anb2 g1436(.dina(new_n1424_), .dinb(new_n1427_), .dout(new_n1501_));
  and1 g1437(.dina(G15), .dinb(G24), .dout(new_n1502_));
  nor2 g1438(.dina(G16), .dinb(G23), .dout(new_n1503_));
  anb1 g1439(.dina(new_n1418_), .dinb(new_n1421_), .dout(new_n1504_));
  anb1 g1440(.dina(new_n1503_), .dinb(new_n1504_), .dout(new_n1505_));
  anb2 g1441(.dina(new_n1503_), .dinb(new_n1504_), .dout(new_n1506_));
  nab1 g1442(.dina(new_n1505_), .dinb(new_n1506_), .dout(new_n1507_));
  anb2 g1443(.dina(new_n1502_), .dinb(new_n1507_), .dout(new_n1508_));
  anb1 g1444(.dina(new_n1502_), .dinb(new_n1507_), .dout(new_n1509_));
  nab2 g1445(.dina(new_n1508_), .dinb(new_n1509_), .dout(new_n1510_));
  anb1 g1446(.dina(new_n1501_), .dinb(new_n1510_), .dout(new_n1511_));
  anb2 g1447(.dina(new_n1501_), .dinb(new_n1510_), .dout(new_n1512_));
  nab1 g1448(.dina(new_n1511_), .dinb(new_n1512_), .dout(new_n1513_));
  anb2 g1449(.dina(new_n1500_), .dinb(new_n1513_), .dout(new_n1514_));
  anb1 g1450(.dina(new_n1500_), .dinb(new_n1513_), .dout(new_n1515_));
  nab2 g1451(.dina(new_n1514_), .dinb(new_n1515_), .dout(new_n1516_));
  anb1 g1452(.dina(new_n1499_), .dinb(new_n1516_), .dout(new_n1517_));
  anb2 g1453(.dina(new_n1499_), .dinb(new_n1516_), .dout(new_n1518_));
  nab1 g1454(.dina(new_n1517_), .dinb(new_n1518_), .dout(new_n1519_));
  anb2 g1455(.dina(new_n1498_), .dinb(new_n1519_), .dout(new_n1520_));
  anb1 g1456(.dina(new_n1498_), .dinb(new_n1519_), .dout(new_n1521_));
  nab2 g1457(.dina(new_n1520_), .dinb(new_n1521_), .dout(new_n1522_));
  anb1 g1458(.dina(new_n1497_), .dinb(new_n1522_), .dout(new_n1523_));
  anb2 g1459(.dina(new_n1497_), .dinb(new_n1522_), .dout(new_n1524_));
  nab1 g1460(.dina(new_n1523_), .dinb(new_n1524_), .dout(new_n1525_));
  anb2 g1461(.dina(new_n1496_), .dinb(new_n1525_), .dout(new_n1526_));
  anb1 g1462(.dina(new_n1496_), .dinb(new_n1525_), .dout(new_n1527_));
  nab2 g1463(.dina(new_n1526_), .dinb(new_n1527_), .dout(new_n1528_));
  anb1 g1464(.dina(new_n1495_), .dinb(new_n1528_), .dout(new_n1529_));
  anb2 g1465(.dina(new_n1495_), .dinb(new_n1528_), .dout(new_n1530_));
  nab1 g1466(.dina(new_n1529_), .dinb(new_n1530_), .dout(new_n1531_));
  anb2 g1467(.dina(new_n1494_), .dinb(new_n1531_), .dout(new_n1532_));
  anb1 g1468(.dina(new_n1494_), .dinb(new_n1531_), .dout(new_n1533_));
  nab2 g1469(.dina(new_n1532_), .dinb(new_n1533_), .dout(new_n1534_));
  anb1 g1470(.dina(new_n1493_), .dinb(new_n1534_), .dout(new_n1535_));
  anb2 g1471(.dina(new_n1493_), .dinb(new_n1534_), .dout(new_n1536_));
  nab1 g1472(.dina(new_n1535_), .dinb(new_n1536_), .dout(new_n1537_));
  anb2 g1473(.dina(new_n1492_), .dinb(new_n1537_), .dout(new_n1538_));
  anb1 g1474(.dina(new_n1492_), .dinb(new_n1537_), .dout(new_n1539_));
  nab2 g1475(.dina(new_n1538_), .dinb(new_n1539_), .dout(new_n1540_));
  anb1 g1476(.dina(new_n1491_), .dinb(new_n1540_), .dout(new_n1541_));
  anb2 g1477(.dina(new_n1491_), .dinb(new_n1540_), .dout(new_n1542_));
  anb2 g1478(.dina(new_n1541_), .dinb(new_n1542_), .dout(new_n1543_));
  anb1 g1479(.dina(new_n1490_), .dinb(new_n1543_), .dout(new_n1544_));
  anb2 g1480(.dina(new_n1490_), .dinb(new_n1543_), .dout(new_n1545_));
  anb2 g1481(.dina(new_n1544_), .dinb(new_n1545_), .dout(new_n1546_));
  anb1 g1482(.dina(new_n1489_), .dinb(new_n1546_), .dout(new_n1547_));
  anb2 g1483(.dina(new_n1489_), .dinb(new_n1546_), .dout(new_n1548_));
  anb2 g1484(.dina(new_n1547_), .dinb(new_n1548_), .dout(new_n1549_));
  anb1 g1485(.dina(new_n1488_), .dinb(new_n1549_), .dout(new_n1550_));
  anb2 g1486(.dina(new_n1488_), .dinb(new_n1549_), .dout(new_n1551_));
  anb2 g1487(.dina(new_n1550_), .dinb(new_n1551_), .dout(new_n1552_));
  anb1 g1488(.dina(new_n1487_), .dinb(new_n1552_), .dout(new_n1553_));
  anb2 g1489(.dina(new_n1487_), .dinb(new_n1552_), .dout(new_n1554_));
  anb2 g1490(.dina(new_n1553_), .dinb(new_n1554_), .dout(new_n1555_));
  anb1 g1491(.dina(new_n1486_), .dinb(new_n1555_), .dout(new_n1556_));
  anb2 g1492(.dina(new_n1486_), .dinb(new_n1555_), .dout(new_n1557_));
  anb2 g1493(.dina(new_n1556_), .dinb(new_n1557_), .dout(new_n1558_));
  anb1 g1494(.dina(new_n1485_), .dinb(new_n1558_), .dout(new_n1559_));
  anb2 g1495(.dina(new_n1485_), .dinb(new_n1558_), .dout(new_n1560_));
  anb2 g1496(.dina(new_n1559_), .dinb(new_n1560_), .dout(new_n1561_));
  anb1 g1497(.dina(new_n1484_), .dinb(new_n1561_), .dout(new_n1562_));
  anb2 g1498(.dina(new_n1484_), .dinb(new_n1561_), .dout(new_n1563_));
  anb2 g1499(.dina(new_n1562_), .dinb(new_n1563_), .dout(G6278));
  and2 g1500(.dina(new_n1559_), .dinb(new_n1562_), .dout(new_n1565_));
  and2 g1501(.dina(new_n1553_), .dinb(new_n1556_), .dout(new_n1566_));
  nor2 g1502(.dina(G8), .dinb(G32), .dout(new_n1567_));
  and2 g1503(.dina(new_n1547_), .dinb(new_n1550_), .dout(new_n1568_));
  nor2 g1504(.dina(G9), .dinb(G31), .dout(new_n1569_));
  and2 g1505(.dina(new_n1541_), .dinb(new_n1544_), .dout(new_n1570_));
  nor2 g1506(.dina(G10), .dinb(G30), .dout(new_n1571_));
  anb2 g1507(.dina(new_n1535_), .dinb(new_n1538_), .dout(new_n1572_));
  and1 g1508(.dina(G11), .dinb(G29), .dout(new_n1573_));
  anb2 g1509(.dina(new_n1529_), .dinb(new_n1532_), .dout(new_n1574_));
  and1 g1510(.dina(G12), .dinb(G28), .dout(new_n1575_));
  anb2 g1511(.dina(new_n1523_), .dinb(new_n1526_), .dout(new_n1576_));
  and1 g1512(.dina(G13), .dinb(G27), .dout(new_n1577_));
  anb2 g1513(.dina(new_n1517_), .dinb(new_n1520_), .dout(new_n1578_));
  and1 g1514(.dina(G14), .dinb(G26), .dout(new_n1579_));
  anb2 g1515(.dina(new_n1511_), .dinb(new_n1514_), .dout(new_n1580_));
  nor2 g1516(.dina(G15), .dinb(G25), .dout(new_n1581_));
  and1 g1517(.dina(G16), .dinb(G24), .dout(new_n1582_));
  anb2 g1518(.dina(new_n1505_), .dinb(new_n1508_), .dout(new_n1583_));
  anb2 g1519(.dina(new_n1582_), .dinb(new_n1583_), .dout(new_n1584_));
  anb1 g1520(.dina(new_n1582_), .dinb(new_n1583_), .dout(new_n1585_));
  nab2 g1521(.dina(new_n1584_), .dinb(new_n1585_), .dout(new_n1586_));
  anb1 g1522(.dina(new_n1581_), .dinb(new_n1586_), .dout(new_n1587_));
  anb2 g1523(.dina(new_n1581_), .dinb(new_n1586_), .dout(new_n1588_));
  anb2 g1524(.dina(new_n1587_), .dinb(new_n1588_), .dout(new_n1589_));
  anb1 g1525(.dina(new_n1580_), .dinb(new_n1589_), .dout(new_n1590_));
  anb2 g1526(.dina(new_n1580_), .dinb(new_n1589_), .dout(new_n1591_));
  nab1 g1527(.dina(new_n1590_), .dinb(new_n1591_), .dout(new_n1592_));
  anb2 g1528(.dina(new_n1579_), .dinb(new_n1592_), .dout(new_n1593_));
  anb1 g1529(.dina(new_n1579_), .dinb(new_n1592_), .dout(new_n1594_));
  nab2 g1530(.dina(new_n1593_), .dinb(new_n1594_), .dout(new_n1595_));
  anb1 g1531(.dina(new_n1578_), .dinb(new_n1595_), .dout(new_n1596_));
  anb2 g1532(.dina(new_n1578_), .dinb(new_n1595_), .dout(new_n1597_));
  nab1 g1533(.dina(new_n1596_), .dinb(new_n1597_), .dout(new_n1598_));
  anb2 g1534(.dina(new_n1577_), .dinb(new_n1598_), .dout(new_n1599_));
  anb1 g1535(.dina(new_n1577_), .dinb(new_n1598_), .dout(new_n1600_));
  nab2 g1536(.dina(new_n1599_), .dinb(new_n1600_), .dout(new_n1601_));
  anb1 g1537(.dina(new_n1576_), .dinb(new_n1601_), .dout(new_n1602_));
  anb2 g1538(.dina(new_n1576_), .dinb(new_n1601_), .dout(new_n1603_));
  nab1 g1539(.dina(new_n1602_), .dinb(new_n1603_), .dout(new_n1604_));
  anb2 g1540(.dina(new_n1575_), .dinb(new_n1604_), .dout(new_n1605_));
  anb1 g1541(.dina(new_n1575_), .dinb(new_n1604_), .dout(new_n1606_));
  nab2 g1542(.dina(new_n1605_), .dinb(new_n1606_), .dout(new_n1607_));
  anb1 g1543(.dina(new_n1574_), .dinb(new_n1607_), .dout(new_n1608_));
  anb2 g1544(.dina(new_n1574_), .dinb(new_n1607_), .dout(new_n1609_));
  nab1 g1545(.dina(new_n1608_), .dinb(new_n1609_), .dout(new_n1610_));
  anb2 g1546(.dina(new_n1573_), .dinb(new_n1610_), .dout(new_n1611_));
  anb1 g1547(.dina(new_n1573_), .dinb(new_n1610_), .dout(new_n1612_));
  nab2 g1548(.dina(new_n1611_), .dinb(new_n1612_), .dout(new_n1613_));
  anb1 g1549(.dina(new_n1572_), .dinb(new_n1613_), .dout(new_n1614_));
  anb2 g1550(.dina(new_n1572_), .dinb(new_n1613_), .dout(new_n1615_));
  anb2 g1551(.dina(new_n1614_), .dinb(new_n1615_), .dout(new_n1616_));
  anb1 g1552(.dina(new_n1571_), .dinb(new_n1616_), .dout(new_n1617_));
  anb2 g1553(.dina(new_n1571_), .dinb(new_n1616_), .dout(new_n1618_));
  anb2 g1554(.dina(new_n1617_), .dinb(new_n1618_), .dout(new_n1619_));
  anb1 g1555(.dina(new_n1570_), .dinb(new_n1619_), .dout(new_n1620_));
  anb2 g1556(.dina(new_n1570_), .dinb(new_n1619_), .dout(new_n1621_));
  anb2 g1557(.dina(new_n1620_), .dinb(new_n1621_), .dout(new_n1622_));
  anb1 g1558(.dina(new_n1569_), .dinb(new_n1622_), .dout(new_n1623_));
  anb2 g1559(.dina(new_n1569_), .dinb(new_n1622_), .dout(new_n1624_));
  anb2 g1560(.dina(new_n1623_), .dinb(new_n1624_), .dout(new_n1625_));
  anb1 g1561(.dina(new_n1568_), .dinb(new_n1625_), .dout(new_n1626_));
  anb2 g1562(.dina(new_n1568_), .dinb(new_n1625_), .dout(new_n1627_));
  anb2 g1563(.dina(new_n1626_), .dinb(new_n1627_), .dout(new_n1628_));
  anb1 g1564(.dina(new_n1567_), .dinb(new_n1628_), .dout(new_n1629_));
  anb2 g1565(.dina(new_n1567_), .dinb(new_n1628_), .dout(new_n1630_));
  anb2 g1566(.dina(new_n1629_), .dinb(new_n1630_), .dout(new_n1631_));
  anb1 g1567(.dina(new_n1566_), .dinb(new_n1631_), .dout(new_n1632_));
  anb2 g1568(.dina(new_n1566_), .dinb(new_n1631_), .dout(new_n1633_));
  anb2 g1569(.dina(new_n1632_), .dinb(new_n1633_), .dout(new_n1634_));
  anb1 g1570(.dina(new_n1565_), .dinb(new_n1634_), .dout(new_n1635_));
  anb2 g1571(.dina(new_n1565_), .dinb(new_n1634_), .dout(new_n1636_));
  anb2 g1572(.dina(new_n1635_), .dinb(new_n1636_), .dout(G6279));
  and2 g1573(.dina(new_n1632_), .dinb(new_n1635_), .dout(new_n1638_));
  and2 g1574(.dina(new_n1626_), .dinb(new_n1629_), .dout(new_n1639_));
  nor2 g1575(.dina(G9), .dinb(G32), .dout(new_n1640_));
  and2 g1576(.dina(new_n1620_), .dinb(new_n1623_), .dout(new_n1641_));
  nor2 g1577(.dina(G10), .dinb(G31), .dout(new_n1642_));
  and2 g1578(.dina(new_n1614_), .dinb(new_n1617_), .dout(new_n1643_));
  nor2 g1579(.dina(G11), .dinb(G30), .dout(new_n1644_));
  anb2 g1580(.dina(new_n1608_), .dinb(new_n1611_), .dout(new_n1645_));
  and1 g1581(.dina(G12), .dinb(G29), .dout(new_n1646_));
  anb2 g1582(.dina(new_n1602_), .dinb(new_n1605_), .dout(new_n1647_));
  and1 g1583(.dina(G13), .dinb(G28), .dout(new_n1648_));
  anb2 g1584(.dina(new_n1596_), .dinb(new_n1599_), .dout(new_n1649_));
  and1 g1585(.dina(G14), .dinb(G27), .dout(new_n1650_));
  anb2 g1586(.dina(new_n1590_), .dinb(new_n1593_), .dout(new_n1651_));
  and1 g1587(.dina(G15), .dinb(G26), .dout(new_n1652_));
  nor2 g1588(.dina(G16), .dinb(G25), .dout(new_n1653_));
  anb1 g1589(.dina(new_n1584_), .dinb(new_n1587_), .dout(new_n1654_));
  anb1 g1590(.dina(new_n1653_), .dinb(new_n1654_), .dout(new_n1655_));
  anb2 g1591(.dina(new_n1653_), .dinb(new_n1654_), .dout(new_n1656_));
  nab1 g1592(.dina(new_n1655_), .dinb(new_n1656_), .dout(new_n1657_));
  anb2 g1593(.dina(new_n1652_), .dinb(new_n1657_), .dout(new_n1658_));
  anb1 g1594(.dina(new_n1652_), .dinb(new_n1657_), .dout(new_n1659_));
  nab2 g1595(.dina(new_n1658_), .dinb(new_n1659_), .dout(new_n1660_));
  anb1 g1596(.dina(new_n1651_), .dinb(new_n1660_), .dout(new_n1661_));
  anb2 g1597(.dina(new_n1651_), .dinb(new_n1660_), .dout(new_n1662_));
  nab1 g1598(.dina(new_n1661_), .dinb(new_n1662_), .dout(new_n1663_));
  anb2 g1599(.dina(new_n1650_), .dinb(new_n1663_), .dout(new_n1664_));
  anb1 g1600(.dina(new_n1650_), .dinb(new_n1663_), .dout(new_n1665_));
  nab2 g1601(.dina(new_n1664_), .dinb(new_n1665_), .dout(new_n1666_));
  anb1 g1602(.dina(new_n1649_), .dinb(new_n1666_), .dout(new_n1667_));
  anb2 g1603(.dina(new_n1649_), .dinb(new_n1666_), .dout(new_n1668_));
  nab1 g1604(.dina(new_n1667_), .dinb(new_n1668_), .dout(new_n1669_));
  anb2 g1605(.dina(new_n1648_), .dinb(new_n1669_), .dout(new_n1670_));
  anb1 g1606(.dina(new_n1648_), .dinb(new_n1669_), .dout(new_n1671_));
  nab2 g1607(.dina(new_n1670_), .dinb(new_n1671_), .dout(new_n1672_));
  anb1 g1608(.dina(new_n1647_), .dinb(new_n1672_), .dout(new_n1673_));
  anb2 g1609(.dina(new_n1647_), .dinb(new_n1672_), .dout(new_n1674_));
  nab1 g1610(.dina(new_n1673_), .dinb(new_n1674_), .dout(new_n1675_));
  anb2 g1611(.dina(new_n1646_), .dinb(new_n1675_), .dout(new_n1676_));
  anb1 g1612(.dina(new_n1646_), .dinb(new_n1675_), .dout(new_n1677_));
  nab2 g1613(.dina(new_n1676_), .dinb(new_n1677_), .dout(new_n1678_));
  anb1 g1614(.dina(new_n1645_), .dinb(new_n1678_), .dout(new_n1679_));
  anb2 g1615(.dina(new_n1645_), .dinb(new_n1678_), .dout(new_n1680_));
  anb2 g1616(.dina(new_n1679_), .dinb(new_n1680_), .dout(new_n1681_));
  anb1 g1617(.dina(new_n1644_), .dinb(new_n1681_), .dout(new_n1682_));
  anb2 g1618(.dina(new_n1644_), .dinb(new_n1681_), .dout(new_n1683_));
  anb2 g1619(.dina(new_n1682_), .dinb(new_n1683_), .dout(new_n1684_));
  anb1 g1620(.dina(new_n1643_), .dinb(new_n1684_), .dout(new_n1685_));
  anb2 g1621(.dina(new_n1643_), .dinb(new_n1684_), .dout(new_n1686_));
  anb2 g1622(.dina(new_n1685_), .dinb(new_n1686_), .dout(new_n1687_));
  anb1 g1623(.dina(new_n1642_), .dinb(new_n1687_), .dout(new_n1688_));
  anb2 g1624(.dina(new_n1642_), .dinb(new_n1687_), .dout(new_n1689_));
  anb2 g1625(.dina(new_n1688_), .dinb(new_n1689_), .dout(new_n1690_));
  anb1 g1626(.dina(new_n1641_), .dinb(new_n1690_), .dout(new_n1691_));
  anb2 g1627(.dina(new_n1641_), .dinb(new_n1690_), .dout(new_n1692_));
  anb2 g1628(.dina(new_n1691_), .dinb(new_n1692_), .dout(new_n1693_));
  anb1 g1629(.dina(new_n1640_), .dinb(new_n1693_), .dout(new_n1694_));
  anb2 g1630(.dina(new_n1640_), .dinb(new_n1693_), .dout(new_n1695_));
  anb2 g1631(.dina(new_n1694_), .dinb(new_n1695_), .dout(new_n1696_));
  anb1 g1632(.dina(new_n1639_), .dinb(new_n1696_), .dout(new_n1697_));
  anb2 g1633(.dina(new_n1639_), .dinb(new_n1696_), .dout(new_n1698_));
  anb2 g1634(.dina(new_n1697_), .dinb(new_n1698_), .dout(new_n1699_));
  anb1 g1635(.dina(new_n1638_), .dinb(new_n1699_), .dout(new_n1700_));
  anb2 g1636(.dina(new_n1638_), .dinb(new_n1699_), .dout(new_n1701_));
  anb2 g1637(.dina(new_n1700_), .dinb(new_n1701_), .dout(G6280));
  and2 g1638(.dina(new_n1697_), .dinb(new_n1700_), .dout(new_n1703_));
  and2 g1639(.dina(new_n1691_), .dinb(new_n1694_), .dout(new_n1704_));
  nor2 g1640(.dina(G10), .dinb(G32), .dout(new_n1705_));
  and2 g1641(.dina(new_n1685_), .dinb(new_n1688_), .dout(new_n1706_));
  nor2 g1642(.dina(G11), .dinb(G31), .dout(new_n1707_));
  and2 g1643(.dina(new_n1679_), .dinb(new_n1682_), .dout(new_n1708_));
  nor2 g1644(.dina(G12), .dinb(G30), .dout(new_n1709_));
  anb2 g1645(.dina(new_n1673_), .dinb(new_n1676_), .dout(new_n1710_));
  and1 g1646(.dina(G13), .dinb(G29), .dout(new_n1711_));
  anb2 g1647(.dina(new_n1667_), .dinb(new_n1670_), .dout(new_n1712_));
  and1 g1648(.dina(G14), .dinb(G28), .dout(new_n1713_));
  anb2 g1649(.dina(new_n1661_), .dinb(new_n1664_), .dout(new_n1714_));
  nor2 g1650(.dina(G15), .dinb(G27), .dout(new_n1715_));
  and1 g1651(.dina(G16), .dinb(G26), .dout(new_n1716_));
  anb2 g1652(.dina(new_n1655_), .dinb(new_n1658_), .dout(new_n1717_));
  anb2 g1653(.dina(new_n1716_), .dinb(new_n1717_), .dout(new_n1718_));
  anb1 g1654(.dina(new_n1716_), .dinb(new_n1717_), .dout(new_n1719_));
  nab2 g1655(.dina(new_n1718_), .dinb(new_n1719_), .dout(new_n1720_));
  anb1 g1656(.dina(new_n1715_), .dinb(new_n1720_), .dout(new_n1721_));
  anb2 g1657(.dina(new_n1715_), .dinb(new_n1720_), .dout(new_n1722_));
  anb2 g1658(.dina(new_n1721_), .dinb(new_n1722_), .dout(new_n1723_));
  anb1 g1659(.dina(new_n1714_), .dinb(new_n1723_), .dout(new_n1724_));
  anb2 g1660(.dina(new_n1714_), .dinb(new_n1723_), .dout(new_n1725_));
  nab1 g1661(.dina(new_n1724_), .dinb(new_n1725_), .dout(new_n1726_));
  anb2 g1662(.dina(new_n1713_), .dinb(new_n1726_), .dout(new_n1727_));
  anb1 g1663(.dina(new_n1713_), .dinb(new_n1726_), .dout(new_n1728_));
  nab2 g1664(.dina(new_n1727_), .dinb(new_n1728_), .dout(new_n1729_));
  anb1 g1665(.dina(new_n1712_), .dinb(new_n1729_), .dout(new_n1730_));
  anb2 g1666(.dina(new_n1712_), .dinb(new_n1729_), .dout(new_n1731_));
  nab1 g1667(.dina(new_n1730_), .dinb(new_n1731_), .dout(new_n1732_));
  anb2 g1668(.dina(new_n1711_), .dinb(new_n1732_), .dout(new_n1733_));
  anb1 g1669(.dina(new_n1711_), .dinb(new_n1732_), .dout(new_n1734_));
  nab2 g1670(.dina(new_n1733_), .dinb(new_n1734_), .dout(new_n1735_));
  anb1 g1671(.dina(new_n1710_), .dinb(new_n1735_), .dout(new_n1736_));
  anb2 g1672(.dina(new_n1710_), .dinb(new_n1735_), .dout(new_n1737_));
  anb2 g1673(.dina(new_n1736_), .dinb(new_n1737_), .dout(new_n1738_));
  anb1 g1674(.dina(new_n1709_), .dinb(new_n1738_), .dout(new_n1739_));
  anb2 g1675(.dina(new_n1709_), .dinb(new_n1738_), .dout(new_n1740_));
  anb2 g1676(.dina(new_n1739_), .dinb(new_n1740_), .dout(new_n1741_));
  anb1 g1677(.dina(new_n1708_), .dinb(new_n1741_), .dout(new_n1742_));
  anb2 g1678(.dina(new_n1708_), .dinb(new_n1741_), .dout(new_n1743_));
  anb2 g1679(.dina(new_n1742_), .dinb(new_n1743_), .dout(new_n1744_));
  anb1 g1680(.dina(new_n1707_), .dinb(new_n1744_), .dout(new_n1745_));
  anb2 g1681(.dina(new_n1707_), .dinb(new_n1744_), .dout(new_n1746_));
  anb2 g1682(.dina(new_n1745_), .dinb(new_n1746_), .dout(new_n1747_));
  anb1 g1683(.dina(new_n1706_), .dinb(new_n1747_), .dout(new_n1748_));
  anb2 g1684(.dina(new_n1706_), .dinb(new_n1747_), .dout(new_n1749_));
  anb2 g1685(.dina(new_n1748_), .dinb(new_n1749_), .dout(new_n1750_));
  anb1 g1686(.dina(new_n1705_), .dinb(new_n1750_), .dout(new_n1751_));
  anb2 g1687(.dina(new_n1705_), .dinb(new_n1750_), .dout(new_n1752_));
  anb2 g1688(.dina(new_n1751_), .dinb(new_n1752_), .dout(new_n1753_));
  anb1 g1689(.dina(new_n1704_), .dinb(new_n1753_), .dout(new_n1754_));
  anb2 g1690(.dina(new_n1704_), .dinb(new_n1753_), .dout(new_n1755_));
  anb2 g1691(.dina(new_n1754_), .dinb(new_n1755_), .dout(new_n1756_));
  anb1 g1692(.dina(new_n1703_), .dinb(new_n1756_), .dout(new_n1757_));
  anb2 g1693(.dina(new_n1703_), .dinb(new_n1756_), .dout(new_n1758_));
  anb2 g1694(.dina(new_n1757_), .dinb(new_n1758_), .dout(G6281));
  and2 g1695(.dina(new_n1754_), .dinb(new_n1757_), .dout(new_n1760_));
  and2 g1696(.dina(new_n1748_), .dinb(new_n1751_), .dout(new_n1761_));
  nor2 g1697(.dina(G11), .dinb(G32), .dout(new_n1762_));
  and2 g1698(.dina(new_n1742_), .dinb(new_n1745_), .dout(new_n1763_));
  nor2 g1699(.dina(G12), .dinb(G31), .dout(new_n1764_));
  and2 g1700(.dina(new_n1736_), .dinb(new_n1739_), .dout(new_n1765_));
  nor2 g1701(.dina(G13), .dinb(G30), .dout(new_n1766_));
  anb2 g1702(.dina(new_n1730_), .dinb(new_n1733_), .dout(new_n1767_));
  and1 g1703(.dina(G14), .dinb(G29), .dout(new_n1768_));
  anb2 g1704(.dina(new_n1724_), .dinb(new_n1727_), .dout(new_n1769_));
  and1 g1705(.dina(G15), .dinb(G28), .dout(new_n1770_));
  nor2 g1706(.dina(G16), .dinb(G27), .dout(new_n1771_));
  anb1 g1707(.dina(new_n1718_), .dinb(new_n1721_), .dout(new_n1772_));
  anb1 g1708(.dina(new_n1771_), .dinb(new_n1772_), .dout(new_n1773_));
  anb2 g1709(.dina(new_n1771_), .dinb(new_n1772_), .dout(new_n1774_));
  nab1 g1710(.dina(new_n1773_), .dinb(new_n1774_), .dout(new_n1775_));
  anb2 g1711(.dina(new_n1770_), .dinb(new_n1775_), .dout(new_n1776_));
  anb1 g1712(.dina(new_n1770_), .dinb(new_n1775_), .dout(new_n1777_));
  nab2 g1713(.dina(new_n1776_), .dinb(new_n1777_), .dout(new_n1778_));
  anb1 g1714(.dina(new_n1769_), .dinb(new_n1778_), .dout(new_n1779_));
  anb2 g1715(.dina(new_n1769_), .dinb(new_n1778_), .dout(new_n1780_));
  nab1 g1716(.dina(new_n1779_), .dinb(new_n1780_), .dout(new_n1781_));
  anb2 g1717(.dina(new_n1768_), .dinb(new_n1781_), .dout(new_n1782_));
  anb1 g1718(.dina(new_n1768_), .dinb(new_n1781_), .dout(new_n1783_));
  nab2 g1719(.dina(new_n1782_), .dinb(new_n1783_), .dout(new_n1784_));
  anb1 g1720(.dina(new_n1767_), .dinb(new_n1784_), .dout(new_n1785_));
  anb2 g1721(.dina(new_n1767_), .dinb(new_n1784_), .dout(new_n1786_));
  anb2 g1722(.dina(new_n1785_), .dinb(new_n1786_), .dout(new_n1787_));
  anb1 g1723(.dina(new_n1766_), .dinb(new_n1787_), .dout(new_n1788_));
  anb2 g1724(.dina(new_n1766_), .dinb(new_n1787_), .dout(new_n1789_));
  anb2 g1725(.dina(new_n1788_), .dinb(new_n1789_), .dout(new_n1790_));
  anb1 g1726(.dina(new_n1765_), .dinb(new_n1790_), .dout(new_n1791_));
  anb2 g1727(.dina(new_n1765_), .dinb(new_n1790_), .dout(new_n1792_));
  anb2 g1728(.dina(new_n1791_), .dinb(new_n1792_), .dout(new_n1793_));
  anb1 g1729(.dina(new_n1764_), .dinb(new_n1793_), .dout(new_n1794_));
  anb2 g1730(.dina(new_n1764_), .dinb(new_n1793_), .dout(new_n1795_));
  anb2 g1731(.dina(new_n1794_), .dinb(new_n1795_), .dout(new_n1796_));
  anb1 g1732(.dina(new_n1763_), .dinb(new_n1796_), .dout(new_n1797_));
  anb2 g1733(.dina(new_n1763_), .dinb(new_n1796_), .dout(new_n1798_));
  anb2 g1734(.dina(new_n1797_), .dinb(new_n1798_), .dout(new_n1799_));
  anb1 g1735(.dina(new_n1762_), .dinb(new_n1799_), .dout(new_n1800_));
  anb2 g1736(.dina(new_n1762_), .dinb(new_n1799_), .dout(new_n1801_));
  anb2 g1737(.dina(new_n1800_), .dinb(new_n1801_), .dout(new_n1802_));
  anb1 g1738(.dina(new_n1761_), .dinb(new_n1802_), .dout(new_n1803_));
  anb2 g1739(.dina(new_n1761_), .dinb(new_n1802_), .dout(new_n1804_));
  anb2 g1740(.dina(new_n1803_), .dinb(new_n1804_), .dout(new_n1805_));
  anb1 g1741(.dina(new_n1760_), .dinb(new_n1805_), .dout(new_n1806_));
  anb2 g1742(.dina(new_n1760_), .dinb(new_n1805_), .dout(new_n1807_));
  anb2 g1743(.dina(new_n1806_), .dinb(new_n1807_), .dout(G6282));
  and2 g1744(.dina(new_n1803_), .dinb(new_n1806_), .dout(new_n1809_));
  and2 g1745(.dina(new_n1797_), .dinb(new_n1800_), .dout(new_n1810_));
  nor2 g1746(.dina(G12), .dinb(G32), .dout(new_n1811_));
  and2 g1747(.dina(new_n1791_), .dinb(new_n1794_), .dout(new_n1812_));
  nor2 g1748(.dina(G13), .dinb(G31), .dout(new_n1813_));
  and2 g1749(.dina(new_n1785_), .dinb(new_n1788_), .dout(new_n1814_));
  nor2 g1750(.dina(G14), .dinb(G30), .dout(new_n1815_));
  anb2 g1751(.dina(new_n1779_), .dinb(new_n1782_), .dout(new_n1816_));
  nor2 g1752(.dina(G15), .dinb(G29), .dout(new_n1817_));
  and1 g1753(.dina(G16), .dinb(G28), .dout(new_n1818_));
  anb2 g1754(.dina(new_n1773_), .dinb(new_n1776_), .dout(new_n1819_));
  anb2 g1755(.dina(new_n1818_), .dinb(new_n1819_), .dout(new_n1820_));
  anb1 g1756(.dina(new_n1818_), .dinb(new_n1819_), .dout(new_n1821_));
  nab2 g1757(.dina(new_n1820_), .dinb(new_n1821_), .dout(new_n1822_));
  anb1 g1758(.dina(new_n1817_), .dinb(new_n1822_), .dout(new_n1823_));
  anb2 g1759(.dina(new_n1817_), .dinb(new_n1822_), .dout(new_n1824_));
  anb2 g1760(.dina(new_n1823_), .dinb(new_n1824_), .dout(new_n1825_));
  anb1 g1761(.dina(new_n1816_), .dinb(new_n1825_), .dout(new_n1826_));
  anb2 g1762(.dina(new_n1816_), .dinb(new_n1825_), .dout(new_n1827_));
  anb2 g1763(.dina(new_n1826_), .dinb(new_n1827_), .dout(new_n1828_));
  anb1 g1764(.dina(new_n1815_), .dinb(new_n1828_), .dout(new_n1829_));
  anb2 g1765(.dina(new_n1815_), .dinb(new_n1828_), .dout(new_n1830_));
  anb2 g1766(.dina(new_n1829_), .dinb(new_n1830_), .dout(new_n1831_));
  anb1 g1767(.dina(new_n1814_), .dinb(new_n1831_), .dout(new_n1832_));
  anb2 g1768(.dina(new_n1814_), .dinb(new_n1831_), .dout(new_n1833_));
  anb2 g1769(.dina(new_n1832_), .dinb(new_n1833_), .dout(new_n1834_));
  anb1 g1770(.dina(new_n1813_), .dinb(new_n1834_), .dout(new_n1835_));
  anb2 g1771(.dina(new_n1813_), .dinb(new_n1834_), .dout(new_n1836_));
  anb2 g1772(.dina(new_n1835_), .dinb(new_n1836_), .dout(new_n1837_));
  anb1 g1773(.dina(new_n1812_), .dinb(new_n1837_), .dout(new_n1838_));
  anb2 g1774(.dina(new_n1812_), .dinb(new_n1837_), .dout(new_n1839_));
  anb2 g1775(.dina(new_n1838_), .dinb(new_n1839_), .dout(new_n1840_));
  anb1 g1776(.dina(new_n1811_), .dinb(new_n1840_), .dout(new_n1841_));
  anb2 g1777(.dina(new_n1811_), .dinb(new_n1840_), .dout(new_n1842_));
  anb2 g1778(.dina(new_n1841_), .dinb(new_n1842_), .dout(new_n1843_));
  anb1 g1779(.dina(new_n1810_), .dinb(new_n1843_), .dout(new_n1844_));
  anb2 g1780(.dina(new_n1810_), .dinb(new_n1843_), .dout(new_n1845_));
  anb2 g1781(.dina(new_n1844_), .dinb(new_n1845_), .dout(new_n1846_));
  anb1 g1782(.dina(new_n1809_), .dinb(new_n1846_), .dout(new_n1847_));
  anb2 g1783(.dina(new_n1809_), .dinb(new_n1846_), .dout(new_n1848_));
  anb2 g1784(.dina(new_n1847_), .dinb(new_n1848_), .dout(G6283));
  and2 g1785(.dina(new_n1844_), .dinb(new_n1847_), .dout(new_n1850_));
  and2 g1786(.dina(new_n1838_), .dinb(new_n1841_), .dout(new_n1851_));
  nor2 g1787(.dina(G13), .dinb(G32), .dout(new_n1852_));
  and2 g1788(.dina(new_n1832_), .dinb(new_n1835_), .dout(new_n1853_));
  nor2 g1789(.dina(G14), .dinb(G31), .dout(new_n1854_));
  and2 g1790(.dina(new_n1826_), .dinb(new_n1829_), .dout(new_n1855_));
  nor2 g1791(.dina(G15), .dinb(G30), .dout(new_n1856_));
  nor2 g1792(.dina(G16), .dinb(G29), .dout(new_n1857_));
  anb1 g1793(.dina(new_n1820_), .dinb(new_n1823_), .dout(new_n1858_));
  anb1 g1794(.dina(new_n1857_), .dinb(new_n1858_), .dout(new_n1859_));
  anb2 g1795(.dina(new_n1857_), .dinb(new_n1858_), .dout(new_n1860_));
  anb2 g1796(.dina(new_n1859_), .dinb(new_n1860_), .dout(new_n1861_));
  anb1 g1797(.dina(new_n1856_), .dinb(new_n1861_), .dout(new_n1862_));
  anb2 g1798(.dina(new_n1856_), .dinb(new_n1861_), .dout(new_n1863_));
  anb2 g1799(.dina(new_n1862_), .dinb(new_n1863_), .dout(new_n1864_));
  anb1 g1800(.dina(new_n1855_), .dinb(new_n1864_), .dout(new_n1865_));
  anb2 g1801(.dina(new_n1855_), .dinb(new_n1864_), .dout(new_n1866_));
  anb2 g1802(.dina(new_n1865_), .dinb(new_n1866_), .dout(new_n1867_));
  anb1 g1803(.dina(new_n1854_), .dinb(new_n1867_), .dout(new_n1868_));
  anb2 g1804(.dina(new_n1854_), .dinb(new_n1867_), .dout(new_n1869_));
  anb2 g1805(.dina(new_n1868_), .dinb(new_n1869_), .dout(new_n1870_));
  anb1 g1806(.dina(new_n1853_), .dinb(new_n1870_), .dout(new_n1871_));
  anb2 g1807(.dina(new_n1853_), .dinb(new_n1870_), .dout(new_n1872_));
  anb2 g1808(.dina(new_n1871_), .dinb(new_n1872_), .dout(new_n1873_));
  anb1 g1809(.dina(new_n1852_), .dinb(new_n1873_), .dout(new_n1874_));
  anb2 g1810(.dina(new_n1852_), .dinb(new_n1873_), .dout(new_n1875_));
  anb2 g1811(.dina(new_n1874_), .dinb(new_n1875_), .dout(new_n1876_));
  anb1 g1812(.dina(new_n1851_), .dinb(new_n1876_), .dout(new_n1877_));
  anb2 g1813(.dina(new_n1851_), .dinb(new_n1876_), .dout(new_n1878_));
  anb2 g1814(.dina(new_n1877_), .dinb(new_n1878_), .dout(new_n1879_));
  anb1 g1815(.dina(new_n1850_), .dinb(new_n1879_), .dout(new_n1880_));
  anb2 g1816(.dina(new_n1850_), .dinb(new_n1879_), .dout(new_n1881_));
  anb2 g1817(.dina(new_n1880_), .dinb(new_n1881_), .dout(G6284));
  and2 g1818(.dina(new_n1877_), .dinb(new_n1880_), .dout(new_n1883_));
  and2 g1819(.dina(new_n1871_), .dinb(new_n1874_), .dout(new_n1884_));
  nor2 g1820(.dina(G14), .dinb(G32), .dout(new_n1885_));
  and2 g1821(.dina(new_n1865_), .dinb(new_n1868_), .dout(new_n1886_));
  nor2 g1822(.dina(G15), .dinb(G31), .dout(new_n1887_));
  nor2 g1823(.dina(G16), .dinb(G30), .dout(new_n1888_));
  nor1 g1824(.dina(new_n1859_), .dinb(new_n1862_), .dout(new_n1889_));
  anb1 g1825(.dina(new_n1888_), .dinb(new_n1889_), .dout(new_n1890_));
  anb2 g1826(.dina(new_n1888_), .dinb(new_n1889_), .dout(new_n1891_));
  anb2 g1827(.dina(new_n1890_), .dinb(new_n1891_), .dout(new_n1892_));
  anb1 g1828(.dina(new_n1887_), .dinb(new_n1892_), .dout(new_n1893_));
  anb2 g1829(.dina(new_n1887_), .dinb(new_n1892_), .dout(new_n1894_));
  anb2 g1830(.dina(new_n1893_), .dinb(new_n1894_), .dout(new_n1895_));
  anb1 g1831(.dina(new_n1886_), .dinb(new_n1895_), .dout(new_n1896_));
  anb2 g1832(.dina(new_n1886_), .dinb(new_n1895_), .dout(new_n1897_));
  anb2 g1833(.dina(new_n1896_), .dinb(new_n1897_), .dout(new_n1898_));
  anb1 g1834(.dina(new_n1885_), .dinb(new_n1898_), .dout(new_n1899_));
  anb2 g1835(.dina(new_n1885_), .dinb(new_n1898_), .dout(new_n1900_));
  anb2 g1836(.dina(new_n1899_), .dinb(new_n1900_), .dout(new_n1901_));
  anb1 g1837(.dina(new_n1884_), .dinb(new_n1901_), .dout(new_n1902_));
  anb2 g1838(.dina(new_n1884_), .dinb(new_n1901_), .dout(new_n1903_));
  anb2 g1839(.dina(new_n1902_), .dinb(new_n1903_), .dout(new_n1904_));
  anb1 g1840(.dina(new_n1883_), .dinb(new_n1904_), .dout(new_n1905_));
  anb2 g1841(.dina(new_n1883_), .dinb(new_n1904_), .dout(new_n1906_));
  anb2 g1842(.dina(new_n1905_), .dinb(new_n1906_), .dout(G6285));
  and2 g1843(.dina(new_n1902_), .dinb(new_n1905_), .dout(new_n1908_));
  and2 g1844(.dina(new_n1896_), .dinb(new_n1899_), .dout(new_n1909_));
  nor2 g1845(.dina(G15), .dinb(G32), .dout(new_n1910_));
  nor2 g1846(.dina(G16), .dinb(G31), .dout(new_n1911_));
  nor1 g1847(.dina(new_n1890_), .dinb(new_n1893_), .dout(new_n1912_));
  anb1 g1848(.dina(new_n1911_), .dinb(new_n1912_), .dout(new_n1913_));
  anb2 g1849(.dina(new_n1911_), .dinb(new_n1912_), .dout(new_n1914_));
  anb2 g1850(.dina(new_n1913_), .dinb(new_n1914_), .dout(new_n1915_));
  anb1 g1851(.dina(new_n1910_), .dinb(new_n1915_), .dout(new_n1916_));
  anb2 g1852(.dina(new_n1910_), .dinb(new_n1915_), .dout(new_n1917_));
  anb2 g1853(.dina(new_n1916_), .dinb(new_n1917_), .dout(new_n1918_));
  anb1 g1854(.dina(new_n1909_), .dinb(new_n1918_), .dout(new_n1919_));
  anb2 g1855(.dina(new_n1909_), .dinb(new_n1918_), .dout(new_n1920_));
  anb2 g1856(.dina(new_n1919_), .dinb(new_n1920_), .dout(new_n1921_));
  anb1 g1857(.dina(new_n1908_), .dinb(new_n1921_), .dout(new_n1922_));
  anb2 g1858(.dina(new_n1908_), .dinb(new_n1921_), .dout(new_n1923_));
  anb2 g1859(.dina(new_n1922_), .dinb(new_n1923_), .dout(G6286));
  nor2 g1860(.dina(G16), .dinb(G32), .dout(new_n1925_));
  nor1 g1861(.dina(new_n1913_), .dinb(new_n1916_), .dout(new_n1926_));
  anb1 g1862(.dina(new_n1925_), .dinb(new_n1926_), .dout(new_n1927_));
  and2 g1863(.dina(new_n1919_), .dinb(new_n1922_), .dout(new_n1928_));
  anb2 g1864(.dina(new_n1925_), .dinb(new_n1926_), .dout(new_n1929_));
  anb2 g1865(.dina(new_n1927_), .dinb(new_n1929_), .dout(new_n1930_));
  anb1 g1866(.dina(new_n1928_), .dinb(new_n1930_), .dout(new_n1931_));
  nor1 g1867(.dina(new_n1927_), .dinb(new_n1931_), .dout(G6287));
  anb2 g1868(.dina(new_n1928_), .dinb(new_n1930_), .dout(new_n1933_));
  anb2 g1869(.dina(new_n1931_), .dinb(new_n1933_), .dout(G6288));
endmodule


