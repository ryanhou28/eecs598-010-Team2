// Benchmark "mymod" written by ABC on Sun Oct 29 19:31:53 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33,
    G1884, G1885, G1886, G1887, G1888, G1889, G1890, G1891, G1892, G1893,
    G1894, G1895, G1896, G1897, G1898, G1899, G1900, G1901, G1902, G1903,
    G1904, G1905, G1906, G1907, G1908  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33;
  output G1884, G1885, G1886, G1887, G1888, G1889, G1890, G1891, G1892, G1893,
    G1894, G1895, G1896, G1897, G1898, G1899, G1900, G1901, G1902, G1903,
    G1904, G1905, G1906, G1907, G1908;
  reg n949_lo, n961_lo, n973_lo, n976_lo, n985_lo, n997_lo, n1009_lo,
    n1021_lo, n1024_lo, n1033_lo, n1036_lo, n1045_lo, n1057_lo, n1069_lo,
    n1081_lo, n1093_lo, n1105_lo, n1117_lo, n1129_lo, n1132_lo, n1141_lo,
    n1144_lo, n1156_lo, n1159_lo, n1165_lo, n1168_lo, n1180_lo, n1189_lo,
    n1192_lo, n1201_lo, n1204_lo, n1216_lo, n1228_lo, n1231_lo, n1237_lo,
    n1240_lo, n1243_lo, n1249_lo, n1252_lo, n1255_lo, n1261_lo, n1264_lo,
    n1267_lo, n1273_lo, n1276_lo, n1279_lo, n1282_lo, n1285_lo, n1288_lo,
    n1291_lo, n1294_lo, n1297_lo, n1300_lo, n1303_lo, n1309_lo, n1312_lo,
    n1315_lo, n1318_lo, n1321_lo, n1324_lo, n1333_lo, n1874_o2, n2180_o2,
    n2372_o2, n2190_o2, n2191_o2, n2212_o2, n2213_o2, n2214_o2, n2215_o2,
    n2275_o2, n2276_o2, n2290_o2, n2291_o2, n2681_o2, n2680_o2, n2683_o2,
    n2684_o2, n2686_o2, n2319_o2, n2320_o2, n304_inv, G554_o2, G557_o2,
    G185_o2, G188_o2, G191_o2, G194_o2, G1182_o2, G1222_o2, G1247_o2,
    G1371_o2, G1383_o2, G1386_o2, n2416_o2, n2428_o2, n2438_o2, n2439_o2,
    n2440_o2, n2444_o2, n2497_o2, n2498_o2, n2503_o2, n2505_o2, n2529_o2,
    n2562_o2, n2570_o2, n2571_o2, n2574_o2, n2575_o2, G546_o2, G550_o2,
    n2633_o2, n2639_o2, n2642_o2, n2645_o2, n2679_o2, n2662_o2, n2724_o2,
    G382_o2, G199_o2, G202_o2, G225_o2, G248_o2, G260_o2, n2716_o2,
    n2737_o2, n1174_lo_buf_o2, n1198_lo_buf_o2, G371_o2, G1059_o2,
    n2586_o2, n2587_o2, n460_inv, n2648_o2, n2649_o2, n2650_o2, n2651_o2,
    n2652_o2, G365_o2, G1496_o2, G1502_o2, n2700_o2, n2701_o2, n2733_o2,
    n2734_o2, n2744_o2, n2747_o2, n2754_o2, n2755_o2, n511_inv, G1609_o2,
    G1625_o2, G738_o2, G755_o2, G1511_o2, G1522_o2, G1538_o2, G1549_o2,
    G1563_o2, G1584_o2, G1576_o2, G1598_o2, G1395_o2, G1410_o2, G1420_o2,
    G1434_o2, n562_inv, n1162_lo_buf_o2, n1102_lo_buf_o2, G359_o2,
    n982_lo_buf_o2, n1030_lo_buf_o2, n1042_lo_buf_o2, n583_inv, G606_o2,
    G1118_o2, G1069_o2, G1145_o2, G1209_o2, G1189_o2, G1699_o2, G1702_o2,
    G1705_o2, G1708_o2, G1684_o2, G1687_o2, G1690_o2, G1693_o2, G1696_o2,
    G1642_o2, G1645_o2, G1648_o2, G1651_o2, G1654_o2, G1657_o2, G1660_o2,
    n1222_lo_buf_o2, n1330_lo_buf_o2, n658_inv, n661_inv, n1306_lo_buf_o2,
    n1150_lo_buf_o2, G175_o2, G241_o2, G356_o2, G989_o2, G984_o2, n685_inv,
    n688_inv, n958_lo_buf_o2, n1114_lo_buf_o2, G182_o2, G1215_o2, G971_o2,
    G938_o2, G1198_o2, G1203_o2, G1218_o2, G785_o2, G1168_o2, G1130_o2,
    G1185_o2, G1250_o2, G1225_o2, G1791_o2, G1788_o2, G981_o2, n745_inv,
    n748_inv, G1062_o2, n970_lo_buf_o2, n1006_lo_buf_o2, n1078_lo_buf_o2,
    n1126_lo_buf_o2, n766_inv, G165_o2, n1234_lo_buf_o2, n1246_lo_buf_o2,
    n1258_lo_buf_o2, n1270_lo_buf_o2, G368_o2, G428_o2, G212_o2, G841_o2,
    G788_o2, n1186_lo_buf_o2, G391_o2, G387_o2, G645_o2, G1140_o2,
    G1178_o2, G1370_o2, n820_inv, G1357_o2, G816_o2, G1369_o2, G901_o2,
    G1056_o2, G1107_o2, G1087_o2, G1135_o2, n1018_lo_buf_o2,
    n1090_lo_buf_o2, n853_inv, G131_o2, n859_inv, n862_inv, G338_o2,
    n1171_lo_buf_o2, n1195_lo_buf_o2, G419_o2, G425_o2, G497_o2, G416_o2,
    G491_o2, G500_o2, G353_o2, G641_o2, G1117_o2, G1096_o2, G1143_o2,
    G1112_o2, n1138_lo_buf_o2, n1210_lo_buf_o2, G687_o2, G541_o2, G802_o2,
    G813_o2, G810_o2, G987_o2, G898_o2, n946_lo_buf_o2, n1054_lo_buf_o2,
    G728_o2, G856_o2, n949_1_inv, G942_o2, G1099_o2, G1154_o2, G1131_o2,
    G1169_o2, G134_o2, n970_inv, G470_o2, G344_o2, G362_o2, G482_o2,
    G660_o2, G672_o2, n1096_lo_buf_o2, G479_o2, G669_o2, n994_lo_buf_o2,
    n1066_lo_buf_o2, n1006_inv, G147_o2, G473_o2, G488_o2, G589_o2,
    G663_o2, G684_o2, G605_o2, G774_o2, G782_o2;
  wire new_new_n709__, new_new_n711__, new_new_n713__, new_new_n715__,
    new_new_n717__, new_new_n719__, new_new_n721__, new_new_n723__,
    new_new_n725__, new_new_n727__, new_new_n729__, new_new_n731__,
    new_new_n733__, new_new_n735__, new_new_n737__, new_new_n739__,
    new_new_n741__, new_new_n743__, new_new_n745__, new_new_n747__,
    new_new_n749__, new_new_n751__, new_new_n753__, new_new_n755__,
    new_new_n757__, new_new_n759__, new_new_n761__, new_new_n763__,
    new_new_n765__, new_new_n767__, new_new_n769__, new_new_n771__,
    new_new_n773__, new_new_n775__, new_new_n776__, new_new_n777__,
    new_new_n778__, new_new_n779__, new_new_n780__, new_new_n781__,
    new_new_n782__, new_new_n783__, new_new_n784__, new_new_n785__,
    new_new_n786__, new_new_n787__, new_new_n788__, new_new_n789__,
    new_new_n790__, new_new_n791__, new_new_n792__, new_new_n793__,
    new_new_n794__, new_new_n795__, new_new_n796__, new_new_n797__,
    new_new_n798__, new_new_n799__, new_new_n800__, new_new_n801__,
    new_new_n802__, new_new_n803__, new_new_n804__, new_new_n805__,
    new_new_n806__, new_new_n807__, new_new_n808__, new_new_n809__,
    new_new_n810__, new_new_n811__, new_new_n812__, new_new_n813__,
    new_new_n815__, new_new_n816__, new_new_n817__, new_new_n818__,
    new_new_n819__, new_new_n821__, new_new_n822__, new_new_n823__,
    new_new_n824__, new_new_n825__, new_new_n827__, new_new_n829__,
    new_new_n830__, new_new_n831__, new_new_n833__, new_new_n834__,
    new_new_n835__, new_new_n837__, new_new_n838__, new_new_n839__,
    new_new_n841__, new_new_n843__, new_new_n844__, new_new_n845__,
    new_new_n847__, new_new_n849__, new_new_n850__, new_new_n851__,
    new_new_n853__, new_new_n855__, new_new_n856__, new_new_n857__,
    new_new_n859__, new_new_n861__, new_new_n862__, new_new_n863__,
    new_new_n865__, new_new_n867__, new_new_n868__, new_new_n869__,
    new_new_n870__, new_new_n871__, new_new_n873__, new_new_n875__,
    new_new_n876__, new_new_n877__, new_new_n878__, new_new_n879__,
    new_new_n881__, new_new_n883__, new_new_n884__, new_new_n885__,
    new_new_n887__, new_new_n889__, new_new_n890__, new_new_n891__,
    new_new_n892__, new_new_n893__, new_new_n894__, new_new_n895__,
    new_new_n896__, new_new_n897__, new_new_n898__, new_new_n899__,
    new_new_n900__, new_new_n901__, new_new_n902__, new_new_n903__,
    new_new_n905__, new_new_n907__, new_new_n909__, new_new_n911__,
    new_new_n913__, new_new_n915__, new_new_n917__, new_new_n919__,
    new_new_n921__, new_new_n923__, new_new_n924__, new_new_n925__,
    new_new_n926__, new_new_n927__, new_new_n928__, new_new_n929__,
    new_new_n930__, new_new_n931__, new_new_n932__, new_new_n933__,
    new_new_n935__, new_new_n937__, new_new_n939__, new_new_n940__,
    new_new_n941__, new_new_n942__, new_new_n943__, new_new_n944__,
    new_new_n945__, new_new_n946__, new_new_n947__, new_new_n948__,
    new_new_n949__, new_new_n950__, new_new_n951__, new_new_n952__,
    new_new_n953__, new_new_n954__, new_new_n955__, new_new_n956__,
    new_new_n957__, new_new_n958__, new_new_n959__, new_new_n960__,
    new_new_n961__, new_new_n962__, new_new_n963__, new_new_n965__,
    new_new_n966__, new_new_n967__, new_new_n969__, new_new_n971__,
    new_new_n973__, new_new_n974__, new_new_n976__, new_new_n977__,
    new_new_n978__, new_new_n979__, new_new_n980__, new_new_n981__,
    new_new_n982__, new_new_n983__, new_new_n984__, new_new_n985__,
    new_new_n986__, new_new_n987__, new_new_n988__, new_new_n989__,
    new_new_n990__, new_new_n991__, new_new_n992__, new_new_n993__,
    new_new_n994__, new_new_n995__, new_new_n996__, new_new_n997__,
    new_new_n998__, new_new_n999__, new_new_n1000__, new_new_n1001__,
    new_new_n1002__, new_new_n1003__, new_new_n1004__, new_new_n1005__,
    new_new_n1006__, new_new_n1007__, new_new_n1009__, new_new_n1010__,
    new_new_n1011__, new_new_n1012__, new_new_n1014__, new_new_n1015__,
    new_new_n1016__, new_new_n1017__, new_new_n1018__, new_new_n1020__,
    new_new_n1021__, new_new_n1022__, new_new_n1023__, new_new_n1024__,
    new_new_n1025__, new_new_n1028__, new_new_n1029__, new_new_n1030__,
    new_new_n1031__, new_new_n1033__, new_new_n1035__, new_new_n1037__,
    new_new_n1039__, new_new_n1041__, new_new_n1043__, new_new_n1045__,
    new_new_n1047__, new_new_n1049__, new_new_n1051__, new_new_n1052__,
    new_new_n1053__, new_new_n1055__, new_new_n1058__, new_new_n1059__,
    new_new_n1061__, new_new_n1063__, new_new_n1065__, new_new_n1067__,
    new_new_n1068__, new_new_n1069__, new_new_n1071__, new_new_n1073__,
    new_new_n1075__, new_new_n1076__, new_new_n1077__, new_new_n1078__,
    new_new_n1079__, new_new_n1080__, new_new_n1081__, new_new_n1082__,
    new_new_n1083__, new_new_n1084__, new_new_n1085__, new_new_n1086__,
    new_new_n1087__, new_new_n1088__, new_new_n1089__, new_new_n1090__,
    new_new_n1091__, new_new_n1092__, new_new_n1093__, new_new_n1094__,
    new_new_n1095__, new_new_n1096__, new_new_n1097__, new_new_n1098__,
    new_new_n1099__, new_new_n1100__, new_new_n1101__, new_new_n1102__,
    new_new_n1103__, new_new_n1104__, new_new_n1105__, new_new_n1106__,
    new_new_n1107__, new_new_n1108__, new_new_n1109__, new_new_n1111__,
    new_new_n1112__, new_new_n1113__, new_new_n1115__, new_new_n1117__,
    new_new_n1119__, new_new_n1121__, new_new_n1123__, new_new_n1125__,
    new_new_n1126__, new_new_n1127__, new_new_n1128__, new_new_n1129__,
    new_new_n1130__, new_new_n1131__, new_new_n1132__, new_new_n1133__,
    new_new_n1134__, new_new_n1135__, new_new_n1136__, new_new_n1137__,
    new_new_n1138__, new_new_n1139__, new_new_n1140__, new_new_n1141__,
    new_new_n1142__, new_new_n1143__, new_new_n1144__, new_new_n1145__,
    new_new_n1146__, new_new_n1147__, new_new_n1148__, new_new_n1149__,
    new_new_n1150__, new_new_n1151__, new_new_n1152__, new_new_n1153__,
    new_new_n1154__, new_new_n1155__, new_new_n1156__, new_new_n1157__,
    new_new_n1158__, new_new_n1159__, new_new_n1160__, new_new_n1161__,
    new_new_n1162__, new_new_n1163__, new_new_n1164__, new_new_n1165__,
    new_new_n1166__, new_new_n1167__, new_new_n1168__, new_new_n1169__,
    new_new_n1171__, new_new_n1173__, new_new_n1175__, new_new_n1177__,
    new_new_n1178__, new_new_n1179__, new_new_n1181__, new_new_n1182__,
    new_new_n1183__, new_new_n1184__, new_new_n1185__, new_new_n1187__,
    new_new_n1189__, new_new_n1191__, new_new_n1193__, new_new_n1195__,
    new_new_n1197__, new_new_n1199__, new_new_n1201__, new_new_n1202__,
    new_new_n1203__, new_new_n1204__, new_new_n1205__, new_new_n1206__,
    new_new_n1207__, new_new_n1208__, new_new_n1209__, new_new_n1210__,
    new_new_n1211__, new_new_n1212__, new_new_n1213__, new_new_n1214__,
    new_new_n1215__, new_new_n1216__, new_new_n1217__, new_new_n1218__,
    new_new_n1219__, new_new_n1220__, new_new_n1221__, new_new_n1222__,
    new_new_n1223__, new_new_n1224__, new_new_n1225__, new_new_n1226__,
    new_new_n1227__, new_new_n1228__, new_new_n1229__, new_new_n1231__,
    new_new_n1233__, new_new_n1234__, new_new_n1235__, new_new_n1237__,
    new_new_n1239__, new_new_n1241__, new_new_n1243__, new_new_n1245__,
    new_new_n1247__, new_new_n1248__, new_new_n1249__, new_new_n1250__,
    new_new_n1251__, new_new_n1252__, new_new_n1253__, new_new_n1254__,
    new_new_n1255__, new_new_n1256__, new_new_n1257__, new_new_n1259__,
    new_new_n1260__, new_new_n1261__, new_new_n1262__, new_new_n1263__,
    new_new_n1264__, new_new_n1265__, new_new_n1266__, new_new_n1267__,
    new_new_n1269__, new_new_n1270__, new_new_n1271__, new_new_n1272__,
    new_new_n1273__, new_new_n1274__, new_new_n1275__, new_new_n1276__,
    new_new_n1277__, new_new_n1278__, new_new_n1279__, new_new_n1280__,
    new_new_n1281__, new_new_n1282__, new_new_n1283__, new_new_n1284__,
    new_new_n1285__, new_new_n1286__, new_new_n1287__, new_new_n1288__,
    new_new_n1289__, new_new_n1290__, new_new_n1291__, new_new_n1292__,
    new_new_n1293__, new_new_n1294__, new_new_n1295__, new_new_n1296__,
    new_new_n1297__, new_new_n1298__, new_new_n1299__, new_new_n1301__,
    new_new_n1303__, new_new_n1304__, new_new_n1305__, new_new_n1306__,
    new_new_n1307__, new_new_n1309__, new_new_n1311__, new_new_n1312__,
    new_new_n1313__, new_new_n1314__, new_new_n1315__, new_new_n1316__,
    new_new_n1317__, new_new_n1318__, new_new_n1319__, new_new_n1320__,
    new_new_n1321__, new_new_n1322__, new_new_n1323__, new_new_n1324__,
    new_new_n1325__, new_new_n1326__, new_new_n1327__, new_new_n1328__,
    new_new_n1329__, new_new_n1330__, new_new_n1331__, new_new_n1332__,
    new_new_n1333__, new_new_n1334__, new_new_n1335__, new_new_n1336__,
    new_new_n1337__, new_new_n1338__, new_new_n1339__, new_new_n1340__,
    new_new_n1341__, new_new_n1342__, new_new_n1343__, new_new_n1344__,
    new_new_n1345__, new_new_n1346__, new_new_n1347__, new_new_n1348__,
    new_new_n1349__, new_new_n1350__, new_new_n1351__, new_new_n1352__,
    new_new_n1353__, new_new_n1354__, new_new_n1355__, new_new_n1356__,
    new_new_n1357__, new_new_n1358__, new_new_n1359__, new_new_n1361__,
    new_new_n1363__, new_new_n1364__, new_new_n1365__, new_new_n1366__,
    new_new_n1367__, new_new_n1368__, new_new_n1369__, new_new_n1370__,
    new_new_n1371__, new_new_n1372__, new_new_n1373__, new_new_n1374__,
    new_new_n1375__, new_new_n1376__, new_new_n1377__, new_new_n1378__,
    new_new_n1379__, new_new_n1380__, new_new_n1381__, new_new_n1383__,
    new_new_n1384__, new_new_n1385__, new_new_n1386__, new_new_n1387__,
    new_new_n1389__, new_new_n1390__, new_new_n1391__, new_new_n1392__,
    new_new_n1393__, new_new_n1394__, new_new_n1395__, new_new_n1396__,
    new_new_n1397__, new_new_n1398__, new_new_n1399__, new_new_n1400__,
    new_new_n1401__, new_new_n1402__, new_new_n1403__, new_new_n1404__,
    new_new_n1405__, new_new_n1406__, new_new_n1407__, new_new_n1408__,
    new_new_n1409__, new_new_n1410__, new_new_n1411__, new_new_n1412__,
    new_new_n1413__, new_new_n1414__, new_new_n1415__, new_new_n1416__,
    new_new_n1417__, new_new_n1418__, new_new_n1419__, new_new_n1420__,
    new_new_n1421__, new_new_n1422__, new_new_n1423__, new_new_n1424__,
    new_new_n1425__, new_new_n1426__, new_new_n1427__, new_new_n1428__,
    new_new_n1429__, new_new_n1430__, new_new_n1431__, new_new_n1432__,
    new_new_n1433__, new_new_n1434__, new_new_n1435__, new_new_n1436__,
    new_new_n1437__, new_new_n1438__, new_new_n1439__, new_new_n1440__,
    new_new_n1441__, new_new_n1442__, new_new_n1443__, new_new_n1444__,
    new_new_n1445__, new_new_n1446__, new_new_n1447__, new_new_n1448__,
    new_new_n1449__, new_new_n1450__, new_new_n1451__, new_new_n1452__,
    new_new_n1453__, new_new_n1454__, new_new_n1455__, new_new_n1456__,
    new_new_n1457__, new_new_n1458__, new_new_n1459__, new_new_n1460__,
    new_new_n1461__, new_new_n1462__, new_new_n1463__, new_new_n1464__,
    new_new_n1465__, new_new_n1466__, new_new_n1467__, new_new_n1468__,
    new_new_n1469__, new_new_n1470__, new_new_n1471__, new_new_n1472__,
    new_new_n1473__, new_new_n1474__, new_new_n1475__, new_new_n1476__,
    new_new_n1477__, new_new_n1478__, new_new_n1479__, new_new_n1480__,
    new_new_n1481__, new_new_n1482__, new_new_n1483__, new_new_n1484__,
    new_new_n1485__, new_new_n1486__, new_new_n1487__, new_new_n1488__,
    new_new_n1489__, new_new_n1490__, new_new_n1491__, new_new_n1492__,
    new_new_n1493__, new_new_n1494__, new_new_n1495__, new_new_n1496__,
    new_new_n1497__, new_new_n1498__, new_new_n1499__, new_new_n1500__,
    new_new_n1501__, new_new_n1502__, new_new_n1503__, new_new_n1504__,
    new_new_n1505__, new_new_n1506__, new_new_n1507__, new_new_n1508__,
    new_new_n1509__, new_new_n1510__, new_new_n1511__, new_new_n1512__,
    new_new_n1513__, new_new_n1514__, new_new_n1515__, new_new_n1516__,
    new_new_n1517__, new_new_n1518__, new_new_n1519__, new_new_n1520__,
    new_new_n1521__, new_new_n1522__, new_new_n1523__, new_new_n1524__,
    new_new_n1525__, new_new_n1526__, new_new_n1527__, new_new_n1528__,
    new_new_n1529__, new_new_n1530__, new_new_n1531__, new_new_n1532__,
    new_new_n1533__, new_new_n1534__, new_new_n1535__, new_new_n1536__,
    new_new_n1537__, new_new_n1538__, new_new_n1539__, new_new_n1540__,
    new_new_n1541__, new_new_n1542__, new_new_n1543__, new_new_n1544__,
    new_new_n1545__, new_new_n1546__, new_new_n1547__, new_new_n1548__,
    new_new_n1549__, new_new_n1550__, new_new_n1551__, new_new_n1552__,
    new_new_n1553__, new_new_n1554__, new_new_n1555__, new_new_n1556__,
    new_new_n1557__, new_new_n1558__, new_new_n1559__, new_new_n1560__,
    new_new_n1561__, new_new_n1562__, new_new_n1563__, new_new_n1564__,
    new_new_n1565__, new_new_n1566__, new_new_n1567__, new_new_n1568__,
    new_new_n1569__, new_new_n1570__, new_new_n1571__, new_new_n1572__,
    new_new_n1573__, new_new_n1574__, new_new_n1575__, new_new_n1576__,
    new_new_n1577__, new_new_n1578__, new_new_n1579__, new_new_n1580__,
    new_new_n1581__, new_new_n1582__, new_new_n1583__, new_new_n1584__,
    new_new_n1585__, new_new_n1586__, new_new_n1587__, new_new_n1588__,
    new_new_n1589__, new_new_n1590__, new_new_n1591__, new_new_n1592__,
    new_new_n1593__, new_new_n1594__, new_new_n1595__, new_new_n1596__,
    new_new_n1597__, new_new_n1598__, new_new_n1599__, new_new_n1600__,
    new_new_n1601__, new_new_n1602__, new_new_n1603__, new_new_n1604__,
    new_new_n1605__, new_new_n1606__, new_new_n1607__, new_new_n1608__,
    new_new_n1609__, new_new_n1610__, new_new_n1611__, new_new_n1612__,
    new_new_n1613__, new_new_n1614__, new_new_n1615__, new_new_n1616__,
    new_new_n1617__, new_new_n1618__, new_new_n1619__, new_new_n1620__,
    new_new_n1621__, new_new_n1622__, new_new_n1623__, new_new_n1624__,
    new_new_n1625__, new_new_n1626__, new_new_n1627__, new_new_n1628__,
    new_new_n1629__, new_new_n1630__, new_new_n1631__, new_new_n1632__,
    new_new_n1633__, new_new_n1634__, new_new_n1635__, new_new_n1636__,
    new_new_n1637__, new_new_n1638__, new_new_n1639__, new_new_n1640__,
    new_new_n1641__, new_new_n1642__, new_new_n1643__, new_new_n1644__,
    new_new_n1645__, new_new_n1646__, new_new_n1647__, new_new_n1648__,
    new_new_n1649__, new_new_n1650__, new_new_n1651__, new_new_n1652__,
    new_new_n1653__, new_new_n1654__, new_new_n1655__, new_new_n1656__,
    new_new_n1657__, new_new_n1658__, new_new_n1659__, new_new_n1660__,
    new_new_n1661__, new_new_n1662__, new_new_n1663__, new_new_n1664__,
    new_new_n1665__, new_new_n1666__, new_new_n1667__, new_new_n1668__,
    new_new_n1669__, new_new_n1670__, new_new_n1671__, new_new_n1672__,
    new_new_n1673__, new_new_n1674__, new_new_n1675__, new_new_n1676__,
    new_new_n1677__, new_new_n1678__, new_new_n1679__, new_new_n1680__,
    new_new_n1681__, new_new_n1682__, new_new_n1683__, new_new_n1684__,
    new_new_n1685__, new_new_n1686__, new_new_n1687__, new_new_n1688__,
    new_new_n1689__, new_new_n1690__, new_new_n1691__, new_new_n1692__,
    new_new_n1693__, new_new_n1694__, new_new_n1695__, new_new_n1696__,
    new_new_n1697__, new_new_n1698__, new_new_n1699__, new_new_n1700__,
    new_new_n1701__, new_new_n1702__, new_new_n1703__, new_new_n1704__,
    new_new_n1705__, new_new_n1706__, new_new_n1707__, new_new_n1708__,
    new_new_n1709__, new_new_n1710__, new_new_n1711__, new_new_n1712__,
    new_new_n1713__, new_new_n1714__, new_new_n1715__, new_new_n1716__,
    new_new_n1717__, new_new_n1718__, new_new_n1719__, new_new_n1720__,
    new_new_n1721__, new_new_n1722__, new_new_n1723__, new_new_n1724__,
    new_new_n1725__, new_new_n1726__, new_new_n1727__, new_new_n1728__,
    new_new_n1729__, new_new_n1730__, new_new_n1731__, new_new_n1732__,
    new_new_n1733__, new_new_n1734__, new_new_n1735__, new_new_n1736__,
    new_new_n1737__, new_new_n1738__, new_new_n1739__, new_new_n1740__,
    new_new_n1741__, new_new_n1742__, new_new_n1743__, new_new_n1744__,
    new_new_n1745__, new_new_n1746__, new_new_n1747__, new_new_n1748__,
    new_new_n1749__, new_new_n1750__, new_new_n1751__, new_new_n1752__,
    new_new_n1753__, new_new_n1754__, new_new_n1755__, new_new_n1756__,
    new_new_n1757__, new_new_n1758__, new_new_n1759__, new_new_n1760__,
    new_new_n1761__, new_new_n1762__, new_new_n1763__, new_new_n1764__,
    new_new_n1765__, new_new_n1766__, new_new_n1767__, new_new_n1768__,
    new_new_n1769__, new_new_n1770__, new_new_n1771__, new_new_n1772__,
    new_new_n1773__, new_new_n1774__, new_new_n1775__, new_new_n1776__,
    new_new_n1777__, new_new_n1778__, new_new_n1779__, new_new_n1780__,
    new_new_n1781__, new_new_n1782__, new_new_n1783__, new_new_n1784__,
    new_new_n1785__, new_new_n1786__, new_new_n1787__, new_new_n1788__,
    new_new_n1789__, new_new_n1790__, new_new_n1791__, new_new_n1792__,
    new_new_n1793__, new_new_n1794__, new_new_n1795__, new_new_n1796__,
    new_new_n1797__, new_new_n1798__, new_new_n1799__, new_new_n1800__,
    new_new_n1801__, new_new_n1802__, new_new_n1803__, new_new_n1804__,
    new_new_n1805__, new_new_n1806__, new_new_n1807__, new_new_n1808__,
    new_new_n1809__, new_new_n1810__, new_new_n1811__, new_new_n1812__,
    new_new_n1813__, new_new_n1814__, new_new_n1815__, new_new_n1816__,
    new_new_n1817__, new_new_n1818__, new_new_n1819__, new_new_n1820__,
    new_new_n1821__, new_new_n1822__, new_new_n1823__, new_new_n1824__,
    new_new_n1825__, new_new_n1826__, new_new_n1827__, new_new_n1828__,
    new_new_n1829__, new_new_n1830__, new_new_n1831__, new_new_n1832__,
    new_new_n1833__, new_new_n1834__, new_new_n1835__, new_new_n1836__,
    new_new_n1837__, new_new_n1838__, new_new_n1839__, new_new_n1840__,
    new_new_n1841__, new_new_n1842__, new_new_n1843__, new_new_n1844__,
    new_new_n1845__, new_new_n1846__, new_new_n1847__, new_new_n1848__,
    new_new_n1849__, new_new_n1850__, new_new_n1851__, new_new_n1852__,
    new_new_n1853__, new_new_n1854__, new_new_n1855__, new_new_n1856__,
    new_new_n1857__, new_new_n1858__, new_new_n1859__, new_new_n1860__,
    new_new_n1861__, new_new_n1862__, new_new_n1863__, new_new_n1864__,
    new_new_n1865__, new_new_n1866__, new_new_n1867__, new_new_n1868__,
    new_new_n1869__, new_new_n1870__, new_new_n1871__, new_new_n1872__,
    new_new_n1873__, new_new_n1874__, new_new_n1875__, new_new_n1876__,
    new_new_n1877__, new_new_n1878__, new_new_n1879__, new_new_n1880__,
    new_new_n1881__, new_new_n1882__, new_new_n1883__, new_new_n1884__,
    new_new_n1885__, new_new_n1886__, new_new_n1887__, new_new_n1888__,
    new_new_n1889__, new_new_n1890__, new_new_n1891__, new_new_n1892__,
    new_new_n1893__, new_new_n1894__, new_new_n1895__, new_new_n1896__,
    new_new_n1897__, new_new_n1898__, new_new_n1899__, new_new_n1900__,
    new_new_n1901__, new_new_n1902__, new_new_n1903__, new_new_n1904__,
    new_new_n1905__, new_new_n1906__, new_new_n1907__, new_new_n1908__,
    new_new_n1909__, new_new_n1910__, new_new_n1911__, new_new_n1912__,
    new_new_n1913__, new_new_n1914__, new_new_n1915__, new_new_n1916__,
    new_new_n1917__, new_new_n1918__, new_new_n1919__, new_new_n1920__,
    new_new_n1921__, new_new_n1922__, new_new_n1923__, new_new_n1924__,
    new_new_n1925__, new_new_n1926__, new_new_n1927__, new_new_n1928__,
    new_new_n1929__, new_new_n1930__, new_new_n1931__, new_new_n1932__,
    new_new_n1933__, new_new_n1934__, new_new_n1935__, new_new_n1936__,
    new_new_n1937__, new_new_n1938__, new_new_n1939__, new_new_n1940__,
    new_new_n1941__, new_new_n1942__, new_new_n1943__, new_new_n1944__,
    new_new_n1945__, new_new_n1946__, new_new_n1947__, new_new_n1948__,
    new_new_n1949__, new_new_n1950__, new_new_n1951__, new_new_n1952__,
    new_new_n1953__, new_new_n1954__, new_new_n1955__, new_new_n1956__,
    new_new_n1957__, new_new_n1958__, new_new_n1959__, new_new_n1960__,
    new_new_n1961__, new_new_n1962__, new_new_n1963__, new_new_n1964__,
    new_new_n1965__, new_new_n1966__, new_new_n1967__, new_new_n1968__,
    new_new_n1969__, new_new_n1970__, new_new_n1971__, new_new_n1972__,
    new_new_n1973__, new_new_n1974__, new_new_n1975__, new_new_n1976__,
    new_new_n1977__, new_new_n1978__, new_new_n1979__, new_new_n1980__,
    new_new_n1981__, new_new_n1982__, new_new_n1983__, new_new_n1984__,
    new_new_n1985__, new_new_n1986__, new_new_n1987__, new_new_n1988__,
    new_new_n1989__, new_new_n1990__, new_new_n1991__, new_new_n1992__,
    new_new_n1993__, new_new_n1994__, new_new_n1995__, new_new_n1996__,
    new_new_n1997__, new_new_n1998__, new_new_n1999__, new_new_n2000__,
    new_new_n2001__, new_new_n2002__, new_new_n2003__, new_new_n2004__,
    new_new_n2005__, new_new_n2006__, new_new_n2007__, new_new_n2008__,
    new_new_n2009__, new_new_n2010__, new_new_n2011__, new_new_n2012__,
    new_new_n2013__, new_new_n2014__, new_new_n2015__, new_new_n2016__,
    new_new_n2017__, new_new_n2018__, new_new_n2019__, new_new_n2020__,
    new_new_n2021__, new_new_n2022__, new_new_n2023__, new_new_n2024__,
    new_new_n2025__, new_new_n2026__, new_new_n2027__, new_new_n2028__,
    new_new_n2029__, new_new_n2030__, new_new_n2031__, new_new_n2032__,
    new_new_n2033__, new_new_n2034__, new_new_n2035__, new_new_n2036__,
    new_new_n2037__, new_new_n2038__, new_new_n2039__, new_new_n2040__,
    new_new_n2041__, new_new_n2042__, new_new_n2043__, new_new_n2044__,
    new_new_n2045__, new_new_n2046__, new_new_n2047__, new_new_n2048__,
    new_new_n2049__, new_new_n2050__, new_new_n2051__, new_new_n2052__,
    new_new_n2053__, new_new_n2054__, new_new_n2055__, new_new_n2056__,
    new_new_n2057__, new_new_n2058__, new_new_n2059__, new_new_n2060__,
    new_new_n2061__, new_new_n2062__, new_new_n2063__, new_new_n2064__,
    new_new_n2065__, new_new_n2066__, new_new_n2067__, new_new_n2068__,
    new_new_n2069__, new_new_n2070__, new_new_n2071__, new_new_n2072__,
    new_new_n2073__, new_new_n2074__, new_new_n2075__, new_new_n2076__,
    new_new_n2077__, new_new_n2078__, new_new_n2079__, new_new_n2080__,
    new_new_n2081__, new_new_n2082__, new_new_n2083__, new_new_n2084__,
    new_new_n2085__, new_new_n2086__, new_new_n2087__, new_new_n2088__,
    new_new_n2089__, new_new_n2090__, new_new_n2091__, new_new_n2092__,
    new_new_n2093__, new_new_n2094__, new_new_n2095__, new_new_n2096__,
    new_new_n2097__, new_new_n2098__, new_new_n2099__, new_new_n2100__,
    new_new_n2101__, new_new_n2102__, new_new_n2103__, new_new_n2104__,
    new_new_n2105__, new_new_n2106__, new_new_n2107__, new_new_n2108__,
    new_new_n2109__, new_new_n2110__, new_new_n2111__, new_new_n2112__,
    new_new_n2113__, new_new_n2114__, new_new_n2115__, new_new_n2116__,
    new_new_n2117__, new_new_n2118__, new_new_n2119__, new_new_n2120__,
    new_new_n2121__, new_new_n2122__, new_new_n2123__, new_new_n2124__,
    new_new_n2125__, new_new_n2126__, new_new_n2127__, new_new_n2128__,
    new_new_n2129__, new_new_n2130__, new_new_n2131__, new_new_n2132__,
    new_new_n2133__, new_new_n2134__, new_new_n2135__, new_new_n2136__,
    new_new_n2137__, new_new_n2138__, new_new_n2139__, new_new_n2140__,
    new_new_n2141__, new_new_n2142__, new_new_n2143__, new_new_n2144__,
    new_new_n2145__, new_new_n2146__, new_new_n2147__, new_new_n2148__,
    new_new_n2149__, new_new_n2150__, new_new_n2151__, new_new_n2152__,
    new_new_n2153__, new_new_n2154__, new_new_n2155__, new_new_n2156__,
    new_new_n2157__, new_new_n2158__, new_new_n2159__, new_new_n2160__,
    new_new_n2161__, new_new_n2162__, new_new_n2163__, new_new_n2164__,
    new_new_n2165__, new_new_n2166__, new_new_n2167__, new_new_n2168__,
    new_new_n2169__, new_new_n2170__, new_new_n2171__, new_new_n2172__,
    new_new_n2173__, new_new_n2174__, new_new_n2175__, new_new_n2176__,
    new_new_n2177__, new_new_n2178__, new_new_n2179__, new_new_n2180__,
    new_new_n2181__, new_new_n2182__, new_new_n2183__, new_new_n2184__,
    new_new_n2535__, new_new_n2536__, new_new_n2537__, new_new_n2538__,
    new_new_n2539__, new_new_n2540__, new_new_n2541__, new_new_n2542__,
    new_new_n2543__, new_new_n2544__, new_new_n2545__, new_new_n2546__,
    new_new_n2547__, new_new_n2548__, new_new_n2549__, new_new_n2550__,
    new_new_n2551__, new_new_n2552__, new_new_n2553__, new_new_n2554__,
    new_new_n2555__, new_new_n2556__, new_new_n2557__, new_new_n2558__,
    new_new_n2559__, new_new_n2560__, new_new_n2561__, new_new_n2562__,
    new_new_n2563__, new_new_n2564__, new_new_n2565__, new_new_n2566__,
    new_new_n2567__, new_new_n2568__, new_new_n2569__, new_new_n2570__,
    new_new_n2571__, new_new_n2572__, new_new_n2573__, new_new_n2574__,
    new_new_n2575__, new_new_n2576__, new_new_n2577__, new_new_n2578__,
    new_new_n2579__, new_new_n2580__, new_new_n2581__, new_new_n2582__,
    new_new_n2583__, new_new_n2584__, new_new_n2585__, new_new_n2586__,
    new_new_n2587__, new_new_n2588__, new_new_n2589__, new_new_n2590__,
    new_new_n2591__, new_new_n2592__, new_new_n2593__, new_new_n2594__,
    new_new_n2595__, new_new_n2596__, new_new_n2597__, new_new_n2598__,
    new_new_n2599__, new_new_n2600__, new_new_n2601__, new_new_n2602__,
    new_new_n2603__, new_new_n2604__, new_new_n2605__, new_new_n2606__,
    new_new_n2607__, new_new_n2608__, new_new_n2609__, new_new_n2610__,
    new_new_n2611__, new_new_n2612__, new_new_n2613__, new_new_n2614__,
    new_new_n2615__, new_new_n2616__, new_new_n2617__, new_new_n2618__,
    new_new_n2619__, new_new_n2620__, new_new_n2621__, new_new_n2622__,
    new_new_n2623__, new_new_n2624__, new_new_n2625__, new_new_n2626__,
    new_new_n2627__, new_new_n2628__, new_new_n2629__, new_new_n2630__,
    new_new_n2631__, new_new_n2632__, new_new_n2633__, new_new_n2634__,
    new_new_n2635__, new_new_n2636__, new_new_n2637__, new_new_n2638__,
    new_new_n2639__, new_new_n2640__, new_new_n2641__, new_new_n2642__,
    new_new_n2643__, new_new_n2644__, new_new_n2645__, new_new_n2646__,
    new_new_n2647__, new_new_n2648__, new_new_n2649__, new_new_n2650__,
    new_new_n2651__, new_new_n2652__, new_new_n2653__, new_new_n2654__,
    new_new_n2655__, new_new_n2656__, new_new_n2657__, new_new_n2658__,
    new_new_n2659__, new_new_n2660__, new_new_n2661__, new_new_n2662__,
    new_new_n2663__, new_new_n2664__, new_new_n2665__, new_new_n2666__,
    new_new_n2667__, new_new_n2668__, new_new_n2669__, new_new_n2670__,
    new_new_n2671__, new_new_n2672__, new_new_n2673__, new_new_n2674__,
    new_new_n2675__, new_new_n2676__, new_new_n2677__, new_new_n2678__,
    new_new_n2679__, new_new_n2680__, new_new_n2681__, new_new_n2682__,
    new_new_n2683__, new_new_n2684__, new_new_n2685__, new_new_n2686__,
    new_new_n2687__, new_new_n2688__, new_new_n2689__, new_new_n2690__,
    new_new_n2691__, new_new_n2692__, new_new_n2693__, new_new_n2694__,
    new_new_n2695__, new_new_n2696__, new_new_n2697__, new_new_n2698__,
    new_new_n2699__, new_new_n2700__, new_new_n2701__, new_new_n2702__,
    new_new_n2703__, new_new_n2704__, new_new_n2705__, new_new_n2706__,
    new_new_n2707__, new_new_n2708__, new_new_n2709__, new_new_n2710__,
    new_new_n2711__, new_new_n2712__, new_new_n2713__, new_new_n2714__,
    new_new_n2715__, new_new_n2716__, new_new_n2717__, new_new_n2718__,
    new_new_n2719__, new_new_n2720__, new_new_n2721__, new_new_n2722__,
    new_new_n2723__, new_new_n2724__, new_new_n2725__, new_new_n2726__,
    new_new_n2727__, new_new_n2728__, new_new_n2729__, new_new_n2730__,
    new_new_n2731__, new_new_n2732__, new_new_n2733__, new_new_n2734__,
    new_new_n2735__, new_new_n2736__, new_new_n2737__, new_new_n2738__,
    new_new_n2739__, new_new_n2740__, new_new_n2741__, new_new_n2742__,
    new_new_n2743__, new_new_n2744__, new_new_n2745__, new_new_n2746__,
    new_new_n2747__, new_new_n2748__, new_new_n2749__, new_new_n2750__,
    new_new_n2751__, new_new_n2752__, new_new_n2753__, new_new_n2754__,
    new_new_n2755__, new_new_n2756__, new_new_n2757__, new_new_n2758__,
    new_new_n2759__, new_new_n2760__, new_new_n2761__, new_new_n2762__,
    new_new_n2763__, new_new_n2764__, new_new_n2765__, new_new_n2766__,
    new_new_n2767__, new_new_n2768__, new_new_n2769__, new_new_n2770__,
    new_new_n2771__, new_new_n2772__, new_new_n2773__, new_new_n2774__,
    new_new_n2775__, new_new_n2776__, new_new_n2777__, new_new_n2778__,
    new_new_n2779__, new_new_n2780__, new_new_n2781__, new_new_n2782__,
    new_new_n2783__, new_new_n2784__, new_new_n2785__, new_new_n2786__,
    new_new_n2787__, new_new_n2788__, new_new_n2789__, new_new_n2790__,
    new_new_n2791__, new_new_n2792__, new_new_n2793__, new_new_n2794__,
    new_new_n2795__, new_new_n2796__, new_new_n2797__, new_new_n2798__,
    new_new_n2799__, new_new_n2800__, new_new_n2801__, new_new_n2802__,
    new_new_n2803__, new_new_n2804__, new_new_n2805__, new_new_n2806__,
    new_new_n2807__, new_new_n2808__, new_new_n2809__, new_new_n2810__,
    new_new_n2811__, new_new_n2812__, new_new_n2813__, new_new_n2814__,
    new_new_n2815__, new_new_n2816__, new_new_n2817__, new_new_n2818__,
    new_new_n2819__, new_new_n2820__, new_new_n2821__, new_new_n2822__,
    new_new_n2823__, new_new_n2824__, new_new_n2825__, new_new_n2826__,
    new_new_n2827__, new_new_n2828__, new_new_n2829__, new_new_n2830__,
    new_new_n2831__, new_new_n2832__, new_new_n2833__, new_new_n2834__,
    new_new_n2835__, new_new_n2836__, new_new_n2837__, new_new_n2838__,
    new_new_n2839__, new_new_n2840__, new_new_n2841__, new_new_n2842__,
    new_new_n2843__, new_new_n2844__, new_new_n2845__, new_new_n2846__,
    new_new_n2847__, new_new_n2848__, new_new_n2849__, new_new_n2850__,
    new_new_n2851__, new_new_n2852__, new_new_n2853__, new_new_n2854__,
    new_new_n2855__, new_new_n2856__, new_new_n2857__, new_new_n2858__,
    new_new_n2859__, new_new_n2860__, new_new_n2861__, new_new_n2862__,
    new_new_n2863__, new_new_n2864__, new_new_n2865__, new_new_n2866__,
    new_new_n2867__, new_new_n2868__, new_new_n2869__, new_new_n2870__,
    new_new_n2871__, new_new_n2872__, new_new_n2873__, new_new_n2874__,
    new_new_n2875__, new_new_n2876__, new_new_n2877__, new_new_n2878__,
    new_new_n2879__, new_new_n2880__, new_new_n2881__, new_new_n2882__,
    new_new_n2883__, new_new_n2884__, new_new_n2885__, new_new_n2886__,
    new_new_n2887__, new_new_n2888__, new_new_n2889__, new_new_n2890__,
    new_new_n2891__, new_new_n2892__, new_new_n2893__, new_new_n2894__,
    new_new_n2895__, new_new_n2896__, new_new_n2897__, new_new_n2898__,
    new_new_n2899__, new_new_n2900__, new_new_n2901__, new_new_n2902__,
    new_new_n2903__, new_new_n2904__, new_new_n2905__, new_new_n2906__,
    new_new_n2907__, new_new_n2908__, new_new_n2909__, new_new_n2910__,
    new_new_n2911__, new_new_n2912__, new_new_n2913__, new_new_n2914__,
    new_new_n2915__, new_new_n2916__, new_new_n2917__, new_new_n2918__,
    new_new_n2919__, new_new_n2920__, new_new_n2921__, new_new_n2922__,
    new_new_n2923__, new_new_n2924__, new_new_n2925__, new_new_n2926__,
    new_new_n2927__, new_new_n2928__, new_new_n2929__, new_new_n2930__,
    new_new_n2931__, new_new_n2932__, new_new_n2933__, new_new_n2934__,
    new_new_n2935__, new_new_n2936__, new_new_n2937__, new_new_n2938__,
    new_new_n2939__, new_new_n2940__, new_new_n2941__, new_new_n2942__,
    new_new_n2943__, new_new_n2944__, new_new_n2945__, new_new_n2946__,
    new_new_n2947__, new_new_n2948__, new_new_n2949__, new_new_n2950__,
    new_new_n2951__, new_new_n2952__, new_new_n2953__, new_new_n2954__,
    new_new_n2955__, new_new_n2956__, new_new_n2957__, new_new_n2958__,
    new_new_n2959__, new_new_n2960__, new_new_n2961__, new_new_n2962__,
    new_new_n2963__, new_new_n2964__, new_new_n2965__, new_new_n2966__,
    new_new_n2967__, new_new_n2968__, new_new_n2969__, new_new_n2970__,
    new_new_n2971__, new_new_n2972__, new_new_n2973__, new_new_n2974__,
    new_new_n2975__, new_new_n2976__, new_new_n2977__, new_new_n2978__,
    new_new_n2979__, new_new_n2980__, new_new_n2981__, new_new_n2982__,
    new_new_n2983__, new_new_n2984__, new_new_n2985__, new_new_n2986__,
    new_new_n2987__, new_new_n2988__, new_new_n2989__, new_new_n2990__,
    new_new_n2991__, new_new_n2992__, new_new_n2993__, new_new_n2994__,
    new_new_n2995__, new_new_n2996__, new_new_n2997__, new_new_n2998__,
    new_new_n2999__, new_new_n3000__, new_new_n3001__, new_new_n3002__,
    new_new_n3003__, new_new_n3004__, new_new_n3005__, new_new_n3006__,
    new_new_n3007__, new_new_n3008__, new_new_n3009__, new_new_n3010__,
    new_new_n3011__, new_new_n3012__, new_new_n3013__, new_new_n3014__,
    new_new_n3015__, new_new_n3016__, new_new_n3017__, new_new_n3018__,
    new_new_n3019__, new_new_n3020__, new_new_n3021__, new_new_n3022__,
    new_new_n3023__, new_new_n3024__, new_new_n3025__, new_new_n3026__,
    new_new_n3027__, new_new_n3028__, new_new_n3029__, new_new_n3030__,
    new_new_n3031__, new_new_n3032__, new_new_n3033__, new_new_n3034__,
    new_new_n3035__, new_new_n3036__, new_new_n3037__, new_new_n3038__,
    new_new_n3039__, new_new_n3040__, new_new_n3041__, new_new_n3042__,
    new_new_n3043__, new_new_n3044__, new_new_n3045__, new_new_n3046__,
    new_new_n3047__, new_new_n3048__, new_new_n3049__, new_new_n3050__,
    new_new_n3051__, new_new_n3052__, new_new_n3053__, new_new_n3054__,
    new_new_n3055__, new_new_n3056__, new_new_n3057__, new_new_n3058__,
    new_new_n3059__, new_new_n3060__, new_new_n3061__, new_new_n3062__,
    new_new_n3063__, new_new_n3064__, n4857, n4860, n4863, n4866, n4869,
    n4872, n4875, n4878, n4881, n4884, n4887, n4890, n4893, n4896, n4899,
    n4902, n4905, n4908, n4911, n4914, n4917, n4920, n4923, n4926, n4929,
    n4932, n4935, n4938, n4941, n4944, n4947, n4950, n4953, n4956, n4959,
    n4962, n4965, n4968, n4971, n4974, n4977, n4980, n4983, n4986, n4989,
    n4992, n4995, n4998, n5001, n5004, n5007, n5010, n5013, n5016, n5019,
    n5022, n5025, n5028, n5031, n5034, n5037, n5040, n5043, n5046, n5049,
    n5052, n5055, n5058, n5061, n5064, n5067, n5070, n5073, n5076, n5079,
    n5082, n5085, n5088, n5091, n5094, n5097, n5100, n5103, n5106, n5109,
    n5112, n5115, n5118, n5121, n5124, n5127, n5130, n5133, n5136, n5139,
    n5142, n5145, n5148, n5151, n5154, n5157, n5160, n5163, n5166, n5169,
    n5172, n5175, n5178, n5181, n5184, n5187, n5190, n5193, n5196, n5199,
    n5202, n5205, n5208, n5211, n5214, n5217, n5220, n5223, n5226, n5229,
    n5232, n5235, n5238, n5241, n5244, n5247, n5250, n5253, n5256, n5259,
    n5262, n5265, n5268, n5271, n5274, n5277, n5280, n5283, n5286, n5289,
    n5292, n5295, n5298, n5301, n5304, n5307, n5310, n5313, n5316, n5319,
    n5322, n5325, n5328, n5331, n5334, n5337, n5340, n5343, n5346, n5349,
    n5352, n5355, n5358, n5361, n5364, n5367, n5370, n5373, n5376, n5379,
    n5382, n5385, n5388, n5391, n5394, n5397, n5400, n5403, n5406, n5409,
    n5412, n5415, n5418, n5421, n5424, n5427, n5430, n5433, n5436, n5439,
    n5442, n5445, n5448, n5451, n5454, n5457, n5460, n5463, n5466, n5469,
    n5472, n5475, n5478, n5481, n5484, n5487, n5490, n5493, n5496, n5499,
    n5502, n5505, n5508, n5511, n5514, n5517, n5520, n5523, n5526, n5529,
    n5532, n5535, n5538, n5541, n5544, n5547, n5550, n5553, n5556, n5559,
    n5562, n5565, n5568, n5571, n5574, n5577, n5580, n5583, n5586, n5589,
    n5592, n5595, n5598, n5601, n5604, n5607, n5610, n5613, n5616, n5619,
    n5622, n5625, n5628, n5631, n5634, n5637, n5640, n5643, n5646, n5649,
    n5652, n5655, n5658, n5661, n5664, n5667, n5670, n5673, n5676, n5679,
    n5682, n5685, n5688, n5691, n5694, n5697, n5700, n5703, n5706, n5709,
    n5712, n5715, n5718, n5721, n5724, n5727, n5730, n5733, n5736, n5739,
    n5742, n5745, n5748, n5751, n5754, n5757, n5760, n5763, n5766, n5769,
    n5772, n5775, n5778, n5781, n5784, n5787, n5790, n5793, n5796, n5799,
    n5802, n5805, n5808, n5811, n5814, n5817, n5820, n5823, n5826, n5829;
  buf1  g0000(.din(G1), .dout(new_new_n709__));
  buf1  g0001(.din(G2), .dout(new_new_n711__));
  buf1  g0002(.din(G3), .dout(new_new_n713__));
  buf1  g0003(.din(G4), .dout(new_new_n715__));
  buf1  g0004(.din(G5), .dout(new_new_n717__));
  buf1  g0005(.din(G6), .dout(new_new_n719__));
  buf1  g0006(.din(G7), .dout(new_new_n721__));
  buf1  g0007(.din(G8), .dout(new_new_n723__));
  buf1  g0008(.din(G9), .dout(new_new_n725__));
  buf1  g0009(.din(G10), .dout(new_new_n727__));
  buf1  g0010(.din(G11), .dout(new_new_n729__));
  buf1  g0011(.din(G12), .dout(new_new_n731__));
  buf1  g0012(.din(G13), .dout(new_new_n733__));
  buf1  g0013(.din(G14), .dout(new_new_n735__));
  buf1  g0014(.din(G15), .dout(new_new_n737__));
  buf1  g0015(.din(G16), .dout(new_new_n739__));
  buf1  g0016(.din(G17), .dout(new_new_n741__));
  buf1  g0017(.din(G18), .dout(new_new_n743__));
  buf1  g0018(.din(G19), .dout(new_new_n745__));
  buf1  g0019(.din(G20), .dout(new_new_n747__));
  buf1  g0020(.din(G21), .dout(new_new_n749__));
  buf1  g0021(.din(G22), .dout(new_new_n751__));
  buf1  g0022(.din(G23), .dout(new_new_n753__));
  buf1  g0023(.din(G24), .dout(new_new_n755__));
  buf1  g0024(.din(G25), .dout(new_new_n757__));
  buf1  g0025(.din(G26), .dout(new_new_n759__));
  buf1  g0026(.din(G27), .dout(new_new_n761__));
  buf1  g0027(.din(G28), .dout(new_new_n763__));
  buf1  g0028(.din(G29), .dout(new_new_n765__));
  buf1  g0029(.din(G30), .dout(new_new_n767__));
  buf1  g0030(.din(G31), .dout(new_new_n769__));
  buf1  g0031(.din(G32), .dout(new_new_n771__));
  buf1  g0032(.din(G33), .dout(new_new_n773__));
  buf1  g0033(.din(n949_lo), .dout(new_new_n775__));
  not1  g0034(.din(n949_lo), .dout(new_new_n776__));
  buf1  g0035(.din(n961_lo), .dout(new_new_n777__));
  not1  g0036(.din(n961_lo), .dout(new_new_n778__));
  buf1  g0037(.din(n973_lo), .dout(new_new_n779__));
  not1  g0038(.din(n973_lo), .dout(new_new_n780__));
  buf1  g0039(.din(n976_lo), .dout(new_new_n781__));
  not1  g0040(.din(n976_lo), .dout(new_new_n782__));
  buf1  g0041(.din(n985_lo), .dout(new_new_n783__));
  not1  g0042(.din(n985_lo), .dout(new_new_n784__));
  buf1  g0043(.din(n997_lo), .dout(new_new_n785__));
  not1  g0044(.din(n997_lo), .dout(new_new_n786__));
  buf1  g0045(.din(n1009_lo), .dout(new_new_n787__));
  not1  g0046(.din(n1009_lo), .dout(new_new_n788__));
  buf1  g0047(.din(n1021_lo), .dout(new_new_n789__));
  not1  g0048(.din(n1021_lo), .dout(new_new_n790__));
  buf1  g0049(.din(n1024_lo), .dout(new_new_n791__));
  not1  g0050(.din(n1024_lo), .dout(new_new_n792__));
  buf1  g0051(.din(n1033_lo), .dout(new_new_n793__));
  not1  g0052(.din(n1033_lo), .dout(new_new_n794__));
  buf1  g0053(.din(n1036_lo), .dout(new_new_n795__));
  not1  g0054(.din(n1036_lo), .dout(new_new_n796__));
  buf1  g0055(.din(n1045_lo), .dout(new_new_n797__));
  not1  g0056(.din(n1045_lo), .dout(new_new_n798__));
  buf1  g0057(.din(n1057_lo), .dout(new_new_n799__));
  not1  g0058(.din(n1057_lo), .dout(new_new_n800__));
  buf1  g0059(.din(n1069_lo), .dout(new_new_n801__));
  not1  g0060(.din(n1069_lo), .dout(new_new_n802__));
  buf1  g0061(.din(n1081_lo), .dout(new_new_n803__));
  not1  g0062(.din(n1081_lo), .dout(new_new_n804__));
  buf1  g0063(.din(n1093_lo), .dout(new_new_n805__));
  not1  g0064(.din(n1093_lo), .dout(new_new_n806__));
  buf1  g0065(.din(n1105_lo), .dout(new_new_n807__));
  not1  g0066(.din(n1105_lo), .dout(new_new_n808__));
  buf1  g0067(.din(n1117_lo), .dout(new_new_n809__));
  not1  g0068(.din(n1117_lo), .dout(new_new_n810__));
  buf1  g0069(.din(n1129_lo), .dout(new_new_n811__));
  not1  g0070(.din(n1129_lo), .dout(new_new_n812__));
  buf1  g0071(.din(n1132_lo), .dout(new_new_n813__));
  buf1  g0072(.din(n1141_lo), .dout(new_new_n815__));
  not1  g0073(.din(n1141_lo), .dout(new_new_n816__));
  buf1  g0074(.din(n1144_lo), .dout(new_new_n817__));
  not1  g0075(.din(n1144_lo), .dout(new_new_n818__));
  buf1  g0076(.din(n1156_lo), .dout(new_new_n819__));
  buf1  g0077(.din(n1159_lo), .dout(new_new_n821__));
  not1  g0078(.din(n1159_lo), .dout(new_new_n822__));
  buf1  g0079(.din(n1165_lo), .dout(new_new_n823__));
  not1  g0080(.din(n1165_lo), .dout(new_new_n824__));
  buf1  g0081(.din(n1168_lo), .dout(new_new_n825__));
  buf1  g0082(.din(n1180_lo), .dout(new_new_n827__));
  buf1  g0083(.din(n1189_lo), .dout(new_new_n829__));
  not1  g0084(.din(n1189_lo), .dout(new_new_n830__));
  buf1  g0085(.din(n1192_lo), .dout(new_new_n831__));
  buf1  g0086(.din(n1201_lo), .dout(new_new_n833__));
  not1  g0087(.din(n1201_lo), .dout(new_new_n834__));
  buf1  g0088(.din(n1204_lo), .dout(new_new_n835__));
  buf1  g0089(.din(n1216_lo), .dout(new_new_n837__));
  not1  g0090(.din(n1216_lo), .dout(new_new_n838__));
  buf1  g0091(.din(n1228_lo), .dout(new_new_n839__));
  buf1  g0092(.din(n1231_lo), .dout(new_new_n841__));
  buf1  g0093(.din(n1237_lo), .dout(new_new_n843__));
  not1  g0094(.din(n1237_lo), .dout(new_new_n844__));
  buf1  g0095(.din(n1240_lo), .dout(new_new_n845__));
  buf1  g0096(.din(n1243_lo), .dout(new_new_n847__));
  buf1  g0097(.din(n1249_lo), .dout(new_new_n849__));
  not1  g0098(.din(n1249_lo), .dout(new_new_n850__));
  buf1  g0099(.din(n1252_lo), .dout(new_new_n851__));
  buf1  g0100(.din(n1255_lo), .dout(new_new_n853__));
  buf1  g0101(.din(n1261_lo), .dout(new_new_n855__));
  not1  g0102(.din(n1261_lo), .dout(new_new_n856__));
  buf1  g0103(.din(n1264_lo), .dout(new_new_n857__));
  buf1  g0104(.din(n1267_lo), .dout(new_new_n859__));
  buf1  g0105(.din(n1273_lo), .dout(new_new_n861__));
  not1  g0106(.din(n1273_lo), .dout(new_new_n862__));
  buf1  g0107(.din(n1276_lo), .dout(new_new_n863__));
  buf1  g0108(.din(n1279_lo), .dout(new_new_n865__));
  buf1  g0109(.din(n1282_lo), .dout(new_new_n867__));
  not1  g0110(.din(n1282_lo), .dout(new_new_n868__));
  buf1  g0111(.din(n1285_lo), .dout(new_new_n869__));
  not1  g0112(.din(n1285_lo), .dout(new_new_n870__));
  buf1  g0113(.din(n1288_lo), .dout(new_new_n871__));
  buf1  g0114(.din(n1291_lo), .dout(new_new_n873__));
  buf1  g0115(.din(n1294_lo), .dout(new_new_n875__));
  not1  g0116(.din(n1294_lo), .dout(new_new_n876__));
  buf1  g0117(.din(n1297_lo), .dout(new_new_n877__));
  not1  g0118(.din(n1297_lo), .dout(new_new_n878__));
  buf1  g0119(.din(n1300_lo), .dout(new_new_n879__));
  buf1  g0120(.din(n1303_lo), .dout(new_new_n881__));
  buf1  g0121(.din(n1309_lo), .dout(new_new_n883__));
  not1  g0122(.din(n1309_lo), .dout(new_new_n884__));
  buf1  g0123(.din(n1312_lo), .dout(new_new_n885__));
  buf1  g0124(.din(n1315_lo), .dout(new_new_n887__));
  buf1  g0125(.din(n1318_lo), .dout(new_new_n889__));
  not1  g0126(.din(n1318_lo), .dout(new_new_n890__));
  buf1  g0127(.din(n1321_lo), .dout(new_new_n891__));
  not1  g0128(.din(n1321_lo), .dout(new_new_n892__));
  buf1  g0129(.din(n1324_lo), .dout(new_new_n893__));
  not1  g0130(.din(n1324_lo), .dout(new_new_n894__));
  buf1  g0131(.din(n1333_lo), .dout(new_new_n895__));
  not1  g0132(.din(n1333_lo), .dout(new_new_n896__));
  buf1  g0133(.din(n1874_o2), .dout(new_new_n897__));
  not1  g0134(.din(n1874_o2), .dout(new_new_n898__));
  buf1  g0135(.din(n2180_o2), .dout(new_new_n899__));
  not1  g0136(.din(n2180_o2), .dout(new_new_n900__));
  buf1  g0137(.din(n2372_o2), .dout(new_new_n901__));
  not1  g0138(.din(n2372_o2), .dout(new_new_n902__));
  buf1  g0139(.din(n2190_o2), .dout(new_new_n903__));
  buf1  g0140(.din(n2191_o2), .dout(new_new_n905__));
  buf1  g0141(.din(n2212_o2), .dout(new_new_n907__));
  buf1  g0142(.din(n2213_o2), .dout(new_new_n909__));
  buf1  g0143(.din(n2214_o2), .dout(new_new_n911__));
  buf1  g0144(.din(n2215_o2), .dout(new_new_n913__));
  buf1  g0145(.din(n2275_o2), .dout(new_new_n915__));
  buf1  g0146(.din(n2276_o2), .dout(new_new_n917__));
  buf1  g0147(.din(n2290_o2), .dout(new_new_n919__));
  buf1  g0148(.din(n2291_o2), .dout(new_new_n921__));
  buf1  g0149(.din(n2681_o2), .dout(new_new_n923__));
  not1  g0150(.din(n2681_o2), .dout(new_new_n924__));
  buf1  g0151(.din(n2680_o2), .dout(new_new_n925__));
  not1  g0152(.din(n2680_o2), .dout(new_new_n926__));
  buf1  g0153(.din(n2683_o2), .dout(new_new_n927__));
  not1  g0154(.din(n2683_o2), .dout(new_new_n928__));
  buf1  g0155(.din(n2684_o2), .dout(new_new_n929__));
  not1  g0156(.din(n2684_o2), .dout(new_new_n930__));
  buf1  g0157(.din(n2686_o2), .dout(new_new_n931__));
  not1  g0158(.din(n2686_o2), .dout(new_new_n932__));
  buf1  g0159(.din(n2319_o2), .dout(new_new_n933__));
  buf1  g0160(.din(n2320_o2), .dout(new_new_n935__));
  buf1  g0161(.din(n304_inv), .dout(new_new_n937__));
  buf1  g0162(.din(G554_o2), .dout(new_new_n939__));
  not1  g0163(.din(G554_o2), .dout(new_new_n940__));
  buf1  g0164(.din(G557_o2), .dout(new_new_n941__));
  not1  g0165(.din(G557_o2), .dout(new_new_n942__));
  buf1  g0166(.din(G185_o2), .dout(new_new_n943__));
  not1  g0167(.din(G185_o2), .dout(new_new_n944__));
  buf1  g0168(.din(G188_o2), .dout(new_new_n945__));
  not1  g0169(.din(G188_o2), .dout(new_new_n946__));
  buf1  g0170(.din(G191_o2), .dout(new_new_n947__));
  not1  g0171(.din(G191_o2), .dout(new_new_n948__));
  buf1  g0172(.din(G194_o2), .dout(new_new_n949__));
  not1  g0173(.din(G194_o2), .dout(new_new_n950__));
  buf1  g0174(.din(G1182_o2), .dout(new_new_n951__));
  not1  g0175(.din(G1182_o2), .dout(new_new_n952__));
  buf1  g0176(.din(G1222_o2), .dout(new_new_n953__));
  not1  g0177(.din(G1222_o2), .dout(new_new_n954__));
  buf1  g0178(.din(G1247_o2), .dout(new_new_n955__));
  not1  g0179(.din(G1247_o2), .dout(new_new_n956__));
  buf1  g0180(.din(G1371_o2), .dout(new_new_n957__));
  not1  g0181(.din(G1371_o2), .dout(new_new_n958__));
  buf1  g0182(.din(G1383_o2), .dout(new_new_n959__));
  not1  g0183(.din(G1383_o2), .dout(new_new_n960__));
  buf1  g0184(.din(G1386_o2), .dout(new_new_n961__));
  not1  g0185(.din(G1386_o2), .dout(new_new_n962__));
  buf1  g0186(.din(n2416_o2), .dout(new_new_n963__));
  buf1  g0187(.din(n2428_o2), .dout(new_new_n965__));
  not1  g0188(.din(n2428_o2), .dout(new_new_n966__));
  buf1  g0189(.din(n2438_o2), .dout(new_new_n967__));
  buf1  g0190(.din(n2439_o2), .dout(new_new_n969__));
  buf1  g0191(.din(n2440_o2), .dout(new_new_n971__));
  buf1  g0192(.din(n2444_o2), .dout(new_new_n973__));
  not1  g0193(.din(n2444_o2), .dout(new_new_n974__));
  not1  g0194(.din(n2497_o2), .dout(new_new_n976__));
  buf1  g0195(.din(n2498_o2), .dout(new_new_n977__));
  not1  g0196(.din(n2498_o2), .dout(new_new_n978__));
  buf1  g0197(.din(n2503_o2), .dout(new_new_n979__));
  not1  g0198(.din(n2503_o2), .dout(new_new_n980__));
  buf1  g0199(.din(n2505_o2), .dout(new_new_n981__));
  not1  g0200(.din(n2505_o2), .dout(new_new_n982__));
  buf1  g0201(.din(n2529_o2), .dout(new_new_n983__));
  not1  g0202(.din(n2529_o2), .dout(new_new_n984__));
  buf1  g0203(.din(n2562_o2), .dout(new_new_n985__));
  not1  g0204(.din(n2562_o2), .dout(new_new_n986__));
  buf1  g0205(.din(n2570_o2), .dout(new_new_n987__));
  not1  g0206(.din(n2570_o2), .dout(new_new_n988__));
  buf1  g0207(.din(n2571_o2), .dout(new_new_n989__));
  not1  g0208(.din(n2571_o2), .dout(new_new_n990__));
  buf1  g0209(.din(n2574_o2), .dout(new_new_n991__));
  not1  g0210(.din(n2574_o2), .dout(new_new_n992__));
  buf1  g0211(.din(n2575_o2), .dout(new_new_n993__));
  not1  g0212(.din(n2575_o2), .dout(new_new_n994__));
  buf1  g0213(.din(G546_o2), .dout(new_new_n995__));
  not1  g0214(.din(G546_o2), .dout(new_new_n996__));
  buf1  g0215(.din(G550_o2), .dout(new_new_n997__));
  not1  g0216(.din(G550_o2), .dout(new_new_n998__));
  buf1  g0217(.din(n2633_o2), .dout(new_new_n999__));
  not1  g0218(.din(n2633_o2), .dout(new_new_n1000__));
  buf1  g0219(.din(n2639_o2), .dout(new_new_n1001__));
  not1  g0220(.din(n2639_o2), .dout(new_new_n1002__));
  buf1  g0221(.din(n2642_o2), .dout(new_new_n1003__));
  not1  g0222(.din(n2642_o2), .dout(new_new_n1004__));
  buf1  g0223(.din(n2645_o2), .dout(new_new_n1005__));
  not1  g0224(.din(n2645_o2), .dout(new_new_n1006__));
  buf1  g0225(.din(n2679_o2), .dout(new_new_n1007__));
  buf1  g0226(.din(n2662_o2), .dout(new_new_n1009__));
  not1  g0227(.din(n2662_o2), .dout(new_new_n1010__));
  buf1  g0228(.din(n2724_o2), .dout(new_new_n1011__));
  not1  g0229(.din(n2724_o2), .dout(new_new_n1012__));
  not1  g0230(.din(G382_o2), .dout(new_new_n1014__));
  buf1  g0231(.din(G199_o2), .dout(new_new_n1015__));
  not1  g0232(.din(G199_o2), .dout(new_new_n1016__));
  buf1  g0233(.din(G202_o2), .dout(new_new_n1017__));
  not1  g0234(.din(G202_o2), .dout(new_new_n1018__));
  not1  g0235(.din(G225_o2), .dout(new_new_n1020__));
  buf1  g0236(.din(G248_o2), .dout(new_new_n1021__));
  not1  g0237(.din(G248_o2), .dout(new_new_n1022__));
  buf1  g0238(.din(G260_o2), .dout(new_new_n1023__));
  not1  g0239(.din(G260_o2), .dout(new_new_n1024__));
  buf1  g0240(.din(n2716_o2), .dout(new_new_n1025__));
  not1  g0241(.din(n2737_o2), .dout(new_new_n1028__));
  buf1  g0242(.din(n1174_lo_buf_o2), .dout(new_new_n1029__));
  not1  g0243(.din(n1174_lo_buf_o2), .dout(new_new_n1030__));
  buf1  g0244(.din(n1198_lo_buf_o2), .dout(new_new_n1031__));
  buf1  g0245(.din(G371_o2), .dout(new_new_n1033__));
  buf1  g0246(.din(G1059_o2), .dout(new_new_n1035__));
  buf1  g0247(.din(n2586_o2), .dout(new_new_n1037__));
  buf1  g0248(.din(n2587_o2), .dout(new_new_n1039__));
  buf1  g0249(.din(n460_inv), .dout(new_new_n1041__));
  buf1  g0250(.din(n2648_o2), .dout(new_new_n1043__));
  buf1  g0251(.din(n2649_o2), .dout(new_new_n1045__));
  buf1  g0252(.din(n2650_o2), .dout(new_new_n1047__));
  buf1  g0253(.din(n2651_o2), .dout(new_new_n1049__));
  buf1  g0254(.din(n2652_o2), .dout(new_new_n1051__));
  not1  g0255(.din(n2652_o2), .dout(new_new_n1052__));
  buf1  g0256(.din(G365_o2), .dout(new_new_n1053__));
  buf1  g0257(.din(G1496_o2), .dout(new_new_n1055__));
  not1  g0258(.din(G1502_o2), .dout(new_new_n1058__));
  buf1  g0259(.din(n2700_o2), .dout(new_new_n1059__));
  buf1  g0260(.din(n2701_o2), .dout(new_new_n1061__));
  buf1  g0261(.din(n2733_o2), .dout(new_new_n1063__));
  buf1  g0262(.din(n2734_o2), .dout(new_new_n1065__));
  buf1  g0263(.din(n2744_o2), .dout(new_new_n1067__));
  not1  g0264(.din(n2744_o2), .dout(new_new_n1068__));
  buf1  g0265(.din(n2747_o2), .dout(new_new_n1069__));
  buf1  g0266(.din(n2754_o2), .dout(new_new_n1071__));
  buf1  g0267(.din(n2755_o2), .dout(new_new_n1073__));
  buf1  g0268(.din(n511_inv), .dout(new_new_n1075__));
  not1  g0269(.din(n511_inv), .dout(new_new_n1076__));
  buf1  g0270(.din(G1609_o2), .dout(new_new_n1077__));
  not1  g0271(.din(G1609_o2), .dout(new_new_n1078__));
  buf1  g0272(.din(G1625_o2), .dout(new_new_n1079__));
  not1  g0273(.din(G1625_o2), .dout(new_new_n1080__));
  buf1  g0274(.din(G738_o2), .dout(new_new_n1081__));
  not1  g0275(.din(G738_o2), .dout(new_new_n1082__));
  buf1  g0276(.din(G755_o2), .dout(new_new_n1083__));
  not1  g0277(.din(G755_o2), .dout(new_new_n1084__));
  buf1  g0278(.din(G1511_o2), .dout(new_new_n1085__));
  not1  g0279(.din(G1511_o2), .dout(new_new_n1086__));
  buf1  g0280(.din(G1522_o2), .dout(new_new_n1087__));
  not1  g0281(.din(G1522_o2), .dout(new_new_n1088__));
  buf1  g0282(.din(G1538_o2), .dout(new_new_n1089__));
  not1  g0283(.din(G1538_o2), .dout(new_new_n1090__));
  buf1  g0284(.din(G1549_o2), .dout(new_new_n1091__));
  not1  g0285(.din(G1549_o2), .dout(new_new_n1092__));
  buf1  g0286(.din(G1563_o2), .dout(new_new_n1093__));
  not1  g0287(.din(G1563_o2), .dout(new_new_n1094__));
  buf1  g0288(.din(G1584_o2), .dout(new_new_n1095__));
  not1  g0289(.din(G1584_o2), .dout(new_new_n1096__));
  buf1  g0290(.din(G1576_o2), .dout(new_new_n1097__));
  not1  g0291(.din(G1576_o2), .dout(new_new_n1098__));
  buf1  g0292(.din(G1598_o2), .dout(new_new_n1099__));
  not1  g0293(.din(G1598_o2), .dout(new_new_n1100__));
  buf1  g0294(.din(G1395_o2), .dout(new_new_n1101__));
  not1  g0295(.din(G1395_o2), .dout(new_new_n1102__));
  buf1  g0296(.din(G1410_o2), .dout(new_new_n1103__));
  not1  g0297(.din(G1410_o2), .dout(new_new_n1104__));
  buf1  g0298(.din(G1420_o2), .dout(new_new_n1105__));
  not1  g0299(.din(G1420_o2), .dout(new_new_n1106__));
  buf1  g0300(.din(G1434_o2), .dout(new_new_n1107__));
  not1  g0301(.din(G1434_o2), .dout(new_new_n1108__));
  buf1  g0302(.din(n562_inv), .dout(new_new_n1109__));
  buf1  g0303(.din(n1162_lo_buf_o2), .dout(new_new_n1111__));
  not1  g0304(.din(n1162_lo_buf_o2), .dout(new_new_n1112__));
  buf1  g0305(.din(n1102_lo_buf_o2), .dout(new_new_n1113__));
  buf1  g0306(.din(G359_o2), .dout(new_new_n1115__));
  buf1  g0307(.din(n982_lo_buf_o2), .dout(new_new_n1117__));
  buf1  g0308(.din(n1030_lo_buf_o2), .dout(new_new_n1119__));
  buf1  g0309(.din(n1042_lo_buf_o2), .dout(new_new_n1121__));
  buf1  g0310(.din(n583_inv), .dout(new_new_n1123__));
  buf1  g0311(.din(G606_o2), .dout(new_new_n1125__));
  not1  g0312(.din(G606_o2), .dout(new_new_n1126__));
  buf1  g0313(.din(G1118_o2), .dout(new_new_n1127__));
  not1  g0314(.din(G1118_o2), .dout(new_new_n1128__));
  buf1  g0315(.din(G1069_o2), .dout(new_new_n1129__));
  not1  g0316(.din(G1069_o2), .dout(new_new_n1130__));
  buf1  g0317(.din(G1145_o2), .dout(new_new_n1131__));
  not1  g0318(.din(G1145_o2), .dout(new_new_n1132__));
  buf1  g0319(.din(G1209_o2), .dout(new_new_n1133__));
  not1  g0320(.din(G1209_o2), .dout(new_new_n1134__));
  buf1  g0321(.din(G1189_o2), .dout(new_new_n1135__));
  not1  g0322(.din(G1189_o2), .dout(new_new_n1136__));
  buf1  g0323(.din(G1699_o2), .dout(new_new_n1137__));
  not1  g0324(.din(G1699_o2), .dout(new_new_n1138__));
  buf1  g0325(.din(G1702_o2), .dout(new_new_n1139__));
  not1  g0326(.din(G1702_o2), .dout(new_new_n1140__));
  buf1  g0327(.din(G1705_o2), .dout(new_new_n1141__));
  not1  g0328(.din(G1705_o2), .dout(new_new_n1142__));
  buf1  g0329(.din(G1708_o2), .dout(new_new_n1143__));
  not1  g0330(.din(G1708_o2), .dout(new_new_n1144__));
  buf1  g0331(.din(G1684_o2), .dout(new_new_n1145__));
  not1  g0332(.din(G1684_o2), .dout(new_new_n1146__));
  buf1  g0333(.din(G1687_o2), .dout(new_new_n1147__));
  not1  g0334(.din(G1687_o2), .dout(new_new_n1148__));
  buf1  g0335(.din(G1690_o2), .dout(new_new_n1149__));
  not1  g0336(.din(G1690_o2), .dout(new_new_n1150__));
  buf1  g0337(.din(G1693_o2), .dout(new_new_n1151__));
  not1  g0338(.din(G1693_o2), .dout(new_new_n1152__));
  buf1  g0339(.din(G1696_o2), .dout(new_new_n1153__));
  not1  g0340(.din(G1696_o2), .dout(new_new_n1154__));
  buf1  g0341(.din(G1642_o2), .dout(new_new_n1155__));
  not1  g0342(.din(G1642_o2), .dout(new_new_n1156__));
  buf1  g0343(.din(G1645_o2), .dout(new_new_n1157__));
  not1  g0344(.din(G1645_o2), .dout(new_new_n1158__));
  buf1  g0345(.din(G1648_o2), .dout(new_new_n1159__));
  not1  g0346(.din(G1648_o2), .dout(new_new_n1160__));
  buf1  g0347(.din(G1651_o2), .dout(new_new_n1161__));
  not1  g0348(.din(G1651_o2), .dout(new_new_n1162__));
  buf1  g0349(.din(G1654_o2), .dout(new_new_n1163__));
  not1  g0350(.din(G1654_o2), .dout(new_new_n1164__));
  buf1  g0351(.din(G1657_o2), .dout(new_new_n1165__));
  not1  g0352(.din(G1657_o2), .dout(new_new_n1166__));
  buf1  g0353(.din(G1660_o2), .dout(new_new_n1167__));
  not1  g0354(.din(G1660_o2), .dout(new_new_n1168__));
  buf1  g0355(.din(n1222_lo_buf_o2), .dout(new_new_n1169__));
  buf1  g0356(.din(n1330_lo_buf_o2), .dout(new_new_n1171__));
  buf1  g0357(.din(n658_inv), .dout(new_new_n1173__));
  buf1  g0358(.din(n661_inv), .dout(new_new_n1175__));
  buf1  g0359(.din(n1306_lo_buf_o2), .dout(new_new_n1177__));
  not1  g0360(.din(n1306_lo_buf_o2), .dout(new_new_n1178__));
  buf1  g0361(.din(n1150_lo_buf_o2), .dout(new_new_n1179__));
  buf1  g0362(.din(G175_o2), .dout(new_new_n1181__));
  not1  g0363(.din(G175_o2), .dout(new_new_n1182__));
  buf1  g0364(.din(G241_o2), .dout(new_new_n1183__));
  not1  g0365(.din(G241_o2), .dout(new_new_n1184__));
  buf1  g0366(.din(G356_o2), .dout(new_new_n1185__));
  buf1  g0367(.din(G989_o2), .dout(new_new_n1187__));
  buf1  g0368(.din(G984_o2), .dout(new_new_n1189__));
  buf1  g0369(.din(n685_inv), .dout(new_new_n1191__));
  buf1  g0370(.din(n688_inv), .dout(new_new_n1193__));
  buf1  g0371(.din(n958_lo_buf_o2), .dout(new_new_n1195__));
  buf1  g0372(.din(n1114_lo_buf_o2), .dout(new_new_n1197__));
  buf1  g0373(.din(G182_o2), .dout(new_new_n1199__));
  buf1  g0374(.din(G1215_o2), .dout(new_new_n1201__));
  not1  g0375(.din(G1215_o2), .dout(new_new_n1202__));
  buf1  g0376(.din(G971_o2), .dout(new_new_n1203__));
  not1  g0377(.din(G971_o2), .dout(new_new_n1204__));
  buf1  g0378(.din(G938_o2), .dout(new_new_n1205__));
  not1  g0379(.din(G938_o2), .dout(new_new_n1206__));
  buf1  g0380(.din(G1198_o2), .dout(new_new_n1207__));
  not1  g0381(.din(G1198_o2), .dout(new_new_n1208__));
  buf1  g0382(.din(G1203_o2), .dout(new_new_n1209__));
  not1  g0383(.din(G1203_o2), .dout(new_new_n1210__));
  buf1  g0384(.din(G1218_o2), .dout(new_new_n1211__));
  not1  g0385(.din(G1218_o2), .dout(new_new_n1212__));
  buf1  g0386(.din(G785_o2), .dout(new_new_n1213__));
  not1  g0387(.din(G785_o2), .dout(new_new_n1214__));
  buf1  g0388(.din(G1168_o2), .dout(new_new_n1215__));
  not1  g0389(.din(G1168_o2), .dout(new_new_n1216__));
  buf1  g0390(.din(G1130_o2), .dout(new_new_n1217__));
  not1  g0391(.din(G1130_o2), .dout(new_new_n1218__));
  buf1  g0392(.din(G1185_o2), .dout(new_new_n1219__));
  not1  g0393(.din(G1185_o2), .dout(new_new_n1220__));
  buf1  g0394(.din(G1250_o2), .dout(new_new_n1221__));
  not1  g0395(.din(G1250_o2), .dout(new_new_n1222__));
  buf1  g0396(.din(G1225_o2), .dout(new_new_n1223__));
  not1  g0397(.din(G1225_o2), .dout(new_new_n1224__));
  buf1  g0398(.din(G1791_o2), .dout(new_new_n1225__));
  not1  g0399(.din(G1791_o2), .dout(new_new_n1226__));
  buf1  g0400(.din(G1788_o2), .dout(new_new_n1227__));
  not1  g0401(.din(G1788_o2), .dout(new_new_n1228__));
  buf1  g0402(.din(G981_o2), .dout(new_new_n1229__));
  buf1  g0403(.din(n745_inv), .dout(new_new_n1231__));
  buf1  g0404(.din(n748_inv), .dout(new_new_n1233__));
  not1  g0405(.din(n748_inv), .dout(new_new_n1234__));
  buf1  g0406(.din(G1062_o2), .dout(new_new_n1235__));
  buf1  g0407(.din(n970_lo_buf_o2), .dout(new_new_n1237__));
  buf1  g0408(.din(n1006_lo_buf_o2), .dout(new_new_n1239__));
  buf1  g0409(.din(n1078_lo_buf_o2), .dout(new_new_n1241__));
  buf1  g0410(.din(n1126_lo_buf_o2), .dout(new_new_n1243__));
  buf1  g0411(.din(n766_inv), .dout(new_new_n1245__));
  buf1  g0412(.din(G165_o2), .dout(new_new_n1247__));
  not1  g0413(.din(G165_o2), .dout(new_new_n1248__));
  buf1  g0414(.din(n1234_lo_buf_o2), .dout(new_new_n1249__));
  not1  g0415(.din(n1234_lo_buf_o2), .dout(new_new_n1250__));
  buf1  g0416(.din(n1246_lo_buf_o2), .dout(new_new_n1251__));
  not1  g0417(.din(n1246_lo_buf_o2), .dout(new_new_n1252__));
  buf1  g0418(.din(n1258_lo_buf_o2), .dout(new_new_n1253__));
  not1  g0419(.din(n1258_lo_buf_o2), .dout(new_new_n1254__));
  buf1  g0420(.din(n1270_lo_buf_o2), .dout(new_new_n1255__));
  not1  g0421(.din(n1270_lo_buf_o2), .dout(new_new_n1256__));
  buf1  g0422(.din(G368_o2), .dout(new_new_n1257__));
  buf1  g0423(.din(G428_o2), .dout(new_new_n1259__));
  not1  g0424(.din(G428_o2), .dout(new_new_n1260__));
  buf1  g0425(.din(G212_o2), .dout(new_new_n1261__));
  not1  g0426(.din(G212_o2), .dout(new_new_n1262__));
  buf1  g0427(.din(G841_o2), .dout(new_new_n1263__));
  not1  g0428(.din(G841_o2), .dout(new_new_n1264__));
  buf1  g0429(.din(G788_o2), .dout(new_new_n1265__));
  not1  g0430(.din(G788_o2), .dout(new_new_n1266__));
  buf1  g0431(.din(n1186_lo_buf_o2), .dout(new_new_n1267__));
  buf1  g0432(.din(G391_o2), .dout(new_new_n1269__));
  not1  g0433(.din(G391_o2), .dout(new_new_n1270__));
  buf1  g0434(.din(G387_o2), .dout(new_new_n1271__));
  not1  g0435(.din(G387_o2), .dout(new_new_n1272__));
  buf1  g0436(.din(G645_o2), .dout(new_new_n1273__));
  not1  g0437(.din(G645_o2), .dout(new_new_n1274__));
  buf1  g0438(.din(G1140_o2), .dout(new_new_n1275__));
  not1  g0439(.din(G1140_o2), .dout(new_new_n1276__));
  buf1  g0440(.din(G1178_o2), .dout(new_new_n1277__));
  not1  g0441(.din(G1178_o2), .dout(new_new_n1278__));
  buf1  g0442(.din(G1370_o2), .dout(new_new_n1279__));
  not1  g0443(.din(G1370_o2), .dout(new_new_n1280__));
  buf1  g0444(.din(n820_inv), .dout(new_new_n1281__));
  not1  g0445(.din(n820_inv), .dout(new_new_n1282__));
  buf1  g0446(.din(G1357_o2), .dout(new_new_n1283__));
  not1  g0447(.din(G1357_o2), .dout(new_new_n1284__));
  buf1  g0448(.din(G816_o2), .dout(new_new_n1285__));
  not1  g0449(.din(G816_o2), .dout(new_new_n1286__));
  buf1  g0450(.din(G1369_o2), .dout(new_new_n1287__));
  not1  g0451(.din(G1369_o2), .dout(new_new_n1288__));
  buf1  g0452(.din(G901_o2), .dout(new_new_n1289__));
  not1  g0453(.din(G901_o2), .dout(new_new_n1290__));
  buf1  g0454(.din(G1056_o2), .dout(new_new_n1291__));
  not1  g0455(.din(G1056_o2), .dout(new_new_n1292__));
  buf1  g0456(.din(G1107_o2), .dout(new_new_n1293__));
  not1  g0457(.din(G1107_o2), .dout(new_new_n1294__));
  buf1  g0458(.din(G1087_o2), .dout(new_new_n1295__));
  not1  g0459(.din(G1087_o2), .dout(new_new_n1296__));
  buf1  g0460(.din(G1135_o2), .dout(new_new_n1297__));
  not1  g0461(.din(G1135_o2), .dout(new_new_n1298__));
  buf1  g0462(.din(n1018_lo_buf_o2), .dout(new_new_n1299__));
  buf1  g0463(.din(n1090_lo_buf_o2), .dout(new_new_n1301__));
  buf1  g0464(.din(n853_inv), .dout(new_new_n1303__));
  not1  g0465(.din(n853_inv), .dout(new_new_n1304__));
  buf1  g0466(.din(G131_o2), .dout(new_new_n1305__));
  not1  g0467(.din(G131_o2), .dout(new_new_n1306__));
  buf1  g0468(.din(n859_inv), .dout(new_new_n1307__));
  buf1  g0469(.din(n862_inv), .dout(new_new_n1309__));
  buf1  g0470(.din(G338_o2), .dout(new_new_n1311__));
  not1  g0471(.din(G338_o2), .dout(new_new_n1312__));
  buf1  g0472(.din(n1171_lo_buf_o2), .dout(new_new_n1313__));
  not1  g0473(.din(n1171_lo_buf_o2), .dout(new_new_n1314__));
  buf1  g0474(.din(n1195_lo_buf_o2), .dout(new_new_n1315__));
  not1  g0475(.din(n1195_lo_buf_o2), .dout(new_new_n1316__));
  buf1  g0476(.din(G419_o2), .dout(new_new_n1317__));
  not1  g0477(.din(G419_o2), .dout(new_new_n1318__));
  buf1  g0478(.din(G425_o2), .dout(new_new_n1319__));
  not1  g0479(.din(G425_o2), .dout(new_new_n1320__));
  buf1  g0480(.din(G497_o2), .dout(new_new_n1321__));
  not1  g0481(.din(G497_o2), .dout(new_new_n1322__));
  buf1  g0482(.din(G416_o2), .dout(new_new_n1323__));
  not1  g0483(.din(G416_o2), .dout(new_new_n1324__));
  buf1  g0484(.din(G491_o2), .dout(new_new_n1325__));
  not1  g0485(.din(G491_o2), .dout(new_new_n1326__));
  buf1  g0486(.din(G500_o2), .dout(new_new_n1327__));
  not1  g0487(.din(G500_o2), .dout(new_new_n1328__));
  buf1  g0488(.din(G353_o2), .dout(new_new_n1329__));
  not1  g0489(.din(G353_o2), .dout(new_new_n1330__));
  buf1  g0490(.din(G641_o2), .dout(new_new_n1331__));
  not1  g0491(.din(G641_o2), .dout(new_new_n1332__));
  buf1  g0492(.din(G1117_o2), .dout(new_new_n1333__));
  not1  g0493(.din(G1117_o2), .dout(new_new_n1334__));
  buf1  g0494(.din(G1096_o2), .dout(new_new_n1335__));
  not1  g0495(.din(G1096_o2), .dout(new_new_n1336__));
  buf1  g0496(.din(G1143_o2), .dout(new_new_n1337__));
  not1  g0497(.din(G1143_o2), .dout(new_new_n1338__));
  buf1  g0498(.din(G1112_o2), .dout(new_new_n1339__));
  not1  g0499(.din(G1112_o2), .dout(new_new_n1340__));
  buf1  g0500(.din(n1138_lo_buf_o2), .dout(new_new_n1341__));
  not1  g0501(.din(n1138_lo_buf_o2), .dout(new_new_n1342__));
  buf1  g0502(.din(n1210_lo_buf_o2), .dout(new_new_n1343__));
  not1  g0503(.din(n1210_lo_buf_o2), .dout(new_new_n1344__));
  buf1  g0504(.din(G687_o2), .dout(new_new_n1345__));
  not1  g0505(.din(G687_o2), .dout(new_new_n1346__));
  buf1  g0506(.din(G541_o2), .dout(new_new_n1347__));
  not1  g0507(.din(G541_o2), .dout(new_new_n1348__));
  buf1  g0508(.din(G802_o2), .dout(new_new_n1349__));
  not1  g0509(.din(G802_o2), .dout(new_new_n1350__));
  buf1  g0510(.din(G813_o2), .dout(new_new_n1351__));
  not1  g0511(.din(G813_o2), .dout(new_new_n1352__));
  buf1  g0512(.din(G810_o2), .dout(new_new_n1353__));
  not1  g0513(.din(G810_o2), .dout(new_new_n1354__));
  buf1  g0514(.din(G987_o2), .dout(new_new_n1355__));
  not1  g0515(.din(G987_o2), .dout(new_new_n1356__));
  buf1  g0516(.din(G898_o2), .dout(new_new_n1357__));
  not1  g0517(.din(G898_o2), .dout(new_new_n1358__));
  buf1  g0518(.din(n946_lo_buf_o2), .dout(new_new_n1359__));
  buf1  g0519(.din(n1054_lo_buf_o2), .dout(new_new_n1361__));
  buf1  g0520(.din(G728_o2), .dout(new_new_n1363__));
  not1  g0521(.din(G728_o2), .dout(new_new_n1364__));
  buf1  g0522(.din(G856_o2), .dout(new_new_n1365__));
  not1  g0523(.din(G856_o2), .dout(new_new_n1366__));
  buf1  g0524(.din(n949_1_inv), .dout(new_new_n1367__));
  not1  g0525(.din(n949_1_inv), .dout(new_new_n1368__));
  buf1  g0526(.din(G942_o2), .dout(new_new_n1369__));
  not1  g0527(.din(G942_o2), .dout(new_new_n1370__));
  buf1  g0528(.din(G1099_o2), .dout(new_new_n1371__));
  not1  g0529(.din(G1099_o2), .dout(new_new_n1372__));
  buf1  g0530(.din(G1154_o2), .dout(new_new_n1373__));
  not1  g0531(.din(G1154_o2), .dout(new_new_n1374__));
  buf1  g0532(.din(G1131_o2), .dout(new_new_n1375__));
  not1  g0533(.din(G1131_o2), .dout(new_new_n1376__));
  buf1  g0534(.din(G1169_o2), .dout(new_new_n1377__));
  not1  g0535(.din(G1169_o2), .dout(new_new_n1378__));
  buf1  g0536(.din(G134_o2), .dout(new_new_n1379__));
  not1  g0537(.din(G134_o2), .dout(new_new_n1380__));
  buf1  g0538(.din(n970_inv), .dout(new_new_n1381__));
  buf1  g0539(.din(G470_o2), .dout(new_new_n1383__));
  not1  g0540(.din(G470_o2), .dout(new_new_n1384__));
  buf1  g0541(.din(G344_o2), .dout(new_new_n1385__));
  not1  g0542(.din(G344_o2), .dout(new_new_n1386__));
  buf1  g0543(.din(G362_o2), .dout(new_new_n1387__));
  buf1  g0544(.din(G482_o2), .dout(new_new_n1389__));
  not1  g0545(.din(G482_o2), .dout(new_new_n1390__));
  buf1  g0546(.din(G660_o2), .dout(new_new_n1391__));
  not1  g0547(.din(G660_o2), .dout(new_new_n1392__));
  buf1  g0548(.din(G672_o2), .dout(new_new_n1393__));
  not1  g0549(.din(G672_o2), .dout(new_new_n1394__));
  buf1  g0550(.din(n1096_lo_buf_o2), .dout(new_new_n1395__));
  not1  g0551(.din(n1096_lo_buf_o2), .dout(new_new_n1396__));
  buf1  g0552(.din(G479_o2), .dout(new_new_n1397__));
  not1  g0553(.din(G479_o2), .dout(new_new_n1398__));
  buf1  g0554(.din(G669_o2), .dout(new_new_n1399__));
  not1  g0555(.din(G669_o2), .dout(new_new_n1400__));
  buf1  g0556(.din(n994_lo_buf_o2), .dout(new_new_n1401__));
  not1  g0557(.din(n994_lo_buf_o2), .dout(new_new_n1402__));
  buf1  g0558(.din(n1066_lo_buf_o2), .dout(new_new_n1403__));
  not1  g0559(.din(n1066_lo_buf_o2), .dout(new_new_n1404__));
  buf1  g0560(.din(n1006_inv), .dout(new_new_n1405__));
  not1  g0561(.din(n1006_inv), .dout(new_new_n1406__));
  buf1  g0562(.din(G147_o2), .dout(new_new_n1407__));
  not1  g0563(.din(G147_o2), .dout(new_new_n1408__));
  buf1  g0564(.din(G473_o2), .dout(new_new_n1409__));
  not1  g0565(.din(G473_o2), .dout(new_new_n1410__));
  buf1  g0566(.din(G488_o2), .dout(new_new_n1411__));
  not1  g0567(.din(G488_o2), .dout(new_new_n1412__));
  buf1  g0568(.din(G589_o2), .dout(new_new_n1413__));
  not1  g0569(.din(G589_o2), .dout(new_new_n1414__));
  buf1  g0570(.din(G663_o2), .dout(new_new_n1415__));
  not1  g0571(.din(G663_o2), .dout(new_new_n1416__));
  buf1  g0572(.din(G684_o2), .dout(new_new_n1417__));
  not1  g0573(.din(G684_o2), .dout(new_new_n1418__));
  buf1  g0574(.din(G605_o2), .dout(new_new_n1419__));
  not1  g0575(.din(G605_o2), .dout(new_new_n1420__));
  buf1  g0576(.din(G774_o2), .dout(new_new_n1421__));
  not1  g0577(.din(G774_o2), .dout(new_new_n1422__));
  buf1  g0578(.din(G782_o2), .dout(new_new_n1423__));
  not1  g0579(.din(G782_o2), .dout(new_new_n1424__));
  and1  g0580(.dina(new_new_n2535__), .dinb(new_new_n2536__), .dout(new_new_n1425__));
  or1   g0581(.dina(new_new_n2537__), .dinb(new_new_n2538__), .dout(new_new_n1426__));
  and1  g0582(.dina(new_new_n2540__), .dinb(new_new_n2543__), .dout(new_new_n1427__));
  or1   g0583(.dina(new_new_n2547__), .dinb(new_new_n2550__), .dout(new_new_n1428__));
  and1  g0584(.dina(new_new_n1427__), .dinb(new_new_n2555__), .dout(new_new_n1429__));
  or1   g0585(.dina(new_new_n1428__), .dinb(new_new_n2562__), .dout(new_new_n1430__));
  and1  g0586(.dina(new_new_n1429__), .dinb(new_new_n2566__), .dout(new_new_n1431__));
  or1   g0587(.dina(new_new_n1430__), .dinb(new_new_n2573__), .dout(new_new_n1432__));
  and1  g0588(.dina(new_new_n1431__), .dinb(new_new_n775__), .dout(new_new_n1433__));
  and1  g0589(.dina(new_new_n1432__), .dinb(new_new_n776__), .dout(new_new_n1434__));
  or1   g0590(.dina(new_new_n1434__), .dinb(new_new_n1433__), .dout(new_new_n1435__));
  and1  g0591(.dina(new_new_n2540__), .dinb(new_new_n2580__), .dout(new_new_n1436__));
  or1   g0592(.dina(new_new_n2547__), .dinb(new_new_n2583__), .dout(new_new_n1437__));
  and1  g0593(.dina(new_new_n2584__), .dinb(new_new_n2587__), .dout(new_new_n1438__));
  or1   g0594(.dina(new_new_n2591__), .dinb(new_new_n2594__), .dout(new_new_n1439__));
  and1  g0595(.dina(new_new_n1438__), .dinb(new_new_n2566__), .dout(new_new_n1440__));
  or1   g0596(.dina(new_new_n1439__), .dinb(new_new_n2573__), .dout(new_new_n1441__));
  and1  g0597(.dina(new_new_n1440__), .dinb(new_new_n777__), .dout(new_new_n1442__));
  and1  g0598(.dina(new_new_n1441__), .dinb(new_new_n778__), .dout(new_new_n1443__));
  or1   g0599(.dina(new_new_n1443__), .dinb(new_new_n1442__), .dout(new_new_n1444__));
  and1  g0600(.dina(new_new_n2584__), .dinb(new_new_n2599__), .dout(new_new_n1445__));
  or1   g0601(.dina(new_new_n2591__), .dinb(new_new_n2602__), .dout(new_new_n1446__));
  and1  g0602(.dina(new_new_n1445__), .dinb(new_new_n2567__), .dout(new_new_n1447__));
  or1   g0603(.dina(new_new_n1446__), .dinb(new_new_n2574__), .dout(new_new_n1448__));
  and1  g0604(.dina(new_new_n1447__), .dinb(new_new_n779__), .dout(new_new_n1449__));
  and1  g0605(.dina(new_new_n1448__), .dinb(new_new_n780__), .dout(new_new_n1450__));
  or1   g0606(.dina(new_new_n1450__), .dinb(new_new_n1449__), .dout(new_new_n1451__));
  and1  g0607(.dina(new_new_n2539__), .dinb(new_new_n2605__), .dout(new_new_n1452__));
  or1   g0608(.dina(new_new_n2546__), .dinb(new_new_n2608__), .dout(new_new_n1453__));
  and1  g0609(.dina(new_new_n1452__), .dinb(new_new_n2555__), .dout(new_new_n1454__));
  or1   g0610(.dina(new_new_n1453__), .dinb(new_new_n2562__), .dout(new_new_n1455__));
  and1  g0611(.dina(new_new_n1454__), .dinb(new_new_n2567__), .dout(new_new_n1456__));
  or1   g0612(.dina(new_new_n1455__), .dinb(new_new_n2574__), .dout(new_new_n1457__));
  and1  g0613(.dina(new_new_n1456__), .dinb(new_new_n783__), .dout(new_new_n1458__));
  and1  g0614(.dina(new_new_n1457__), .dinb(new_new_n784__), .dout(new_new_n1459__));
  or1   g0615(.dina(new_new_n1459__), .dinb(new_new_n1458__), .dout(new_new_n1460__));
  and1  g0616(.dina(new_new_n2535__), .dinb(new_new_n2610__), .dout(new_new_n1461__));
  or1   g0617(.dina(new_new_n2537__), .dinb(new_new_n2612__), .dout(new_new_n1462__));
  and1  g0618(.dina(new_new_n1461__), .dinb(new_new_n2614__), .dout(new_new_n1463__));
  or1   g0619(.dina(new_new_n1462__), .dinb(new_new_n2617__), .dout(new_new_n1464__));
  and1  g0620(.dina(new_new_n1463__), .dinb(new_new_n2599__), .dout(new_new_n1465__));
  or1   g0621(.dina(new_new_n1464__), .dinb(new_new_n2602__), .dout(new_new_n1466__));
  and1  g0622(.dina(new_new_n1465__), .dinb(new_new_n2621__), .dout(new_new_n1467__));
  or1   g0623(.dina(new_new_n1466__), .dinb(new_new_n2628__), .dout(new_new_n1468__));
  and1  g0624(.dina(new_new_n1467__), .dinb(new_new_n799__), .dout(new_new_n1469__));
  and1  g0625(.dina(new_new_n1468__), .dinb(new_new_n800__), .dout(new_new_n1470__));
  or1   g0626(.dina(new_new_n1470__), .dinb(new_new_n1469__), .dout(new_new_n1471__));
  and1  g0627(.dina(new_new_n2633__), .dinb(new_new_n2610__), .dout(new_new_n1472__));
  or1   g0628(.dina(new_new_n2634__), .dinb(new_new_n2612__), .dout(new_new_n1473__));
  and1  g0629(.dina(new_new_n2635__), .dinb(new_new_n2543__), .dout(new_new_n1474__));
  or1   g0630(.dina(new_new_n2636__), .dinb(new_new_n2550__), .dout(new_new_n1475__));
  and1  g0631(.dina(new_new_n1474__), .dinb(new_new_n2637__), .dout(new_new_n1476__));
  or1   g0632(.dina(new_new_n1475__), .dinb(new_new_n2638__), .dout(new_new_n1477__));
  and1  g0633(.dina(new_new_n1476__), .dinb(new_new_n2621__), .dout(new_new_n1478__));
  or1   g0634(.dina(new_new_n1477__), .dinb(new_new_n2628__), .dout(new_new_n1479__));
  and1  g0635(.dina(new_new_n1478__), .dinb(new_new_n809__), .dout(new_new_n1480__));
  and1  g0636(.dina(new_new_n1479__), .dinb(new_new_n810__), .dout(new_new_n1481__));
  or1   g0637(.dina(new_new_n1481__), .dinb(new_new_n1480__), .dout(new_new_n1482__));
  and1  g0638(.dina(new_new_n2635__), .dinb(new_new_n2614__), .dout(new_new_n1483__));
  or1   g0639(.dina(new_new_n2636__), .dinb(new_new_n2617__), .dout(new_new_n1484__));
  and1  g0640(.dina(new_new_n1483__), .dinb(new_new_n2587__), .dout(new_new_n1485__));
  or1   g0641(.dina(new_new_n1484__), .dinb(new_new_n2594__), .dout(new_new_n1486__));
  and1  g0642(.dina(new_new_n1485__), .dinb(new_new_n2622__), .dout(new_new_n1487__));
  or1   g0643(.dina(new_new_n1486__), .dinb(new_new_n2629__), .dout(new_new_n1488__));
  and1  g0644(.dina(new_new_n1487__), .dinb(new_new_n811__), .dout(new_new_n1489__));
  and1  g0645(.dina(new_new_n1488__), .dinb(new_new_n812__), .dout(new_new_n1490__));
  or1   g0646(.dina(new_new_n1490__), .dinb(new_new_n1489__), .dout(new_new_n1491__));
  and1  g0647(.dina(new_new_n2536__), .dinb(new_new_n2640__), .dout(new_new_n1492__));
  or1   g0648(.dina(new_new_n2538__), .dinb(new_new_n2642__), .dout(new_new_n1493__));
  and1  g0649(.dina(new_new_n1492__), .dinb(new_new_n2544__), .dout(new_new_n1494__));
  or1   g0650(.dina(new_new_n1493__), .dinb(new_new_n2549__), .dout(new_new_n1495__));
  and1  g0651(.dina(new_new_n1494__), .dinb(new_new_n2588__), .dout(new_new_n1496__));
  or1   g0652(.dina(new_new_n1495__), .dinb(new_new_n2595__), .dout(new_new_n1497__));
  and1  g0653(.dina(new_new_n1496__), .dinb(new_new_n2569__), .dout(new_new_n1498__));
  or1   g0654(.dina(new_new_n1497__), .dinb(new_new_n2576__), .dout(new_new_n1499__));
  and1  g0655(.dina(new_new_n1498__), .dinb(new_new_n785__), .dout(new_new_n1500__));
  and1  g0656(.dina(new_new_n1499__), .dinb(new_new_n786__), .dout(new_new_n1501__));
  or1   g0657(.dina(new_new_n1501__), .dinb(new_new_n1500__), .dout(new_new_n1502__));
  and1  g0658(.dina(new_new_n2609__), .dinb(new_new_n2640__), .dout(new_new_n1503__));
  or1   g0659(.dina(new_new_n2611__), .dinb(new_new_n2642__), .dout(new_new_n1504__));
  and1  g0660(.dina(new_new_n2644__), .dinb(new_new_n2544__), .dout(new_new_n1505__));
  or1   g0661(.dina(new_new_n2647__), .dinb(new_new_n2551__), .dout(new_new_n1506__));
  and1  g0662(.dina(new_new_n1505__), .dinb(new_new_n2598__), .dout(new_new_n1507__));
  or1   g0663(.dina(new_new_n1506__), .dinb(new_new_n2603__), .dout(new_new_n1508__));
  and1  g0664(.dina(new_new_n1507__), .dinb(new_new_n2569__), .dout(new_new_n1509__));
  or1   g0665(.dina(new_new_n1508__), .dinb(new_new_n2576__), .dout(new_new_n1510__));
  and1  g0666(.dina(new_new_n1509__), .dinb(new_new_n787__), .dout(new_new_n1511__));
  and1  g0667(.dina(new_new_n1510__), .dinb(new_new_n788__), .dout(new_new_n1512__));
  or1   g0668(.dina(new_new_n1512__), .dinb(new_new_n1511__), .dout(new_new_n1513__));
  and1  g0669(.dina(new_new_n2644__), .dinb(new_new_n2615__), .dout(new_new_n1514__));
  or1   g0670(.dina(new_new_n2647__), .dinb(new_new_n2618__), .dout(new_new_n1515__));
  and1  g0671(.dina(new_new_n1514__), .dinb(new_new_n2556__), .dout(new_new_n1516__));
  or1   g0672(.dina(new_new_n1515__), .dinb(new_new_n2563__), .dout(new_new_n1517__));
  and1  g0673(.dina(new_new_n1516__), .dinb(new_new_n2570__), .dout(new_new_n1518__));
  or1   g0674(.dina(new_new_n1517__), .dinb(new_new_n2577__), .dout(new_new_n1519__));
  and1  g0675(.dina(new_new_n1518__), .dinb(new_new_n789__), .dout(new_new_n1520__));
  and1  g0676(.dina(new_new_n1519__), .dinb(new_new_n790__), .dout(new_new_n1521__));
  or1   g0677(.dina(new_new_n1521__), .dinb(new_new_n1520__), .dout(new_new_n1522__));
  and1  g0678(.dina(new_new_n2645__), .dinb(new_new_n2580__), .dout(new_new_n1523__));
  or1   g0679(.dina(new_new_n2648__), .dinb(new_new_n2583__), .dout(new_new_n1524__));
  and1  g0680(.dina(new_new_n2649__), .dinb(new_new_n2637__), .dout(new_new_n1525__));
  or1   g0681(.dina(new_new_n1524__), .dinb(new_new_n2638__), .dout(new_new_n1526__));
  and1  g0682(.dina(new_new_n1525__), .dinb(new_new_n2570__), .dout(new_new_n1527__));
  or1   g0683(.dina(new_new_n1526__), .dinb(new_new_n2577__), .dout(new_new_n1528__));
  and1  g0684(.dina(new_new_n1527__), .dinb(new_new_n793__), .dout(new_new_n1529__));
  and1  g0685(.dina(new_new_n1528__), .dinb(new_new_n794__), .dout(new_new_n1530__));
  or1   g0686(.dina(new_new_n1530__), .dinb(new_new_n1529__), .dout(new_new_n1531__));
  and1  g0687(.dina(new_new_n2645__), .dinb(new_new_n2605__), .dout(new_new_n1532__));
  or1   g0688(.dina(new_new_n2648__), .dinb(new_new_n2608__), .dout(new_new_n1533__));
  and1  g0689(.dina(new_new_n1532__), .dinb(new_new_n2588__), .dout(new_new_n1534__));
  or1   g0690(.dina(new_new_n1533__), .dinb(new_new_n2595__), .dout(new_new_n1535__));
  and1  g0691(.dina(new_new_n1534__), .dinb(new_new_n2622__), .dout(new_new_n1536__));
  or1   g0692(.dina(new_new_n1535__), .dinb(new_new_n2629__), .dout(new_new_n1537__));
  and1  g0693(.dina(new_new_n1536__), .dinb(new_new_n797__), .dout(new_new_n1538__));
  and1  g0694(.dina(new_new_n1537__), .dinb(new_new_n798__), .dout(new_new_n1539__));
  or1   g0695(.dina(new_new_n1539__), .dinb(new_new_n1538__), .dout(new_new_n1540__));
  and1  g0696(.dina(new_new_n2633__), .dinb(new_new_n2651__), .dout(new_new_n1541__));
  or1   g0697(.dina(new_new_n2634__), .dinb(new_new_n1078__), .dout(new_new_n1542__));
  and1  g0698(.dina(new_new_n2653__), .dinb(new_new_n2545__), .dout(new_new_n1543__));
  or1   g0699(.dina(new_new_n2656__), .dinb(new_new_n2551__), .dout(new_new_n1544__));
  and1  g0700(.dina(new_new_n2657__), .dinb(new_new_n2590__), .dout(new_new_n1545__));
  or1   g0701(.dina(new_new_n2658__), .dinb(new_new_n2596__), .dout(new_new_n1546__));
  and1  g0702(.dina(new_new_n1545__), .dinb(new_new_n2624__), .dout(new_new_n1547__));
  or1   g0703(.dina(new_new_n1546__), .dinb(new_new_n2631__), .dout(new_new_n1548__));
  and1  g0704(.dina(new_new_n1547__), .dinb(new_new_n801__), .dout(new_new_n1549__));
  and1  g0705(.dina(new_new_n1548__), .dinb(new_new_n802__), .dout(new_new_n1550__));
  or1   g0706(.dina(new_new_n1550__), .dinb(new_new_n1549__), .dout(new_new_n1551__));
  and1  g0707(.dina(new_new_n2657__), .dinb(new_new_n2600__), .dout(new_new_n1552__));
  or1   g0708(.dina(new_new_n2658__), .dinb(new_new_n2603__), .dout(new_new_n1553__));
  and1  g0709(.dina(new_new_n1552__), .dinb(new_new_n2624__), .dout(new_new_n1554__));
  or1   g0710(.dina(new_new_n1553__), .dinb(new_new_n2631__), .dout(new_new_n1555__));
  and1  g0711(.dina(new_new_n1554__), .dinb(new_new_n803__), .dout(new_new_n1556__));
  and1  g0712(.dina(new_new_n1555__), .dinb(new_new_n804__), .dout(new_new_n1557__));
  or1   g0713(.dina(new_new_n1557__), .dinb(new_new_n1556__), .dout(new_new_n1558__));
  and1  g0714(.dina(new_new_n2653__), .dinb(new_new_n2615__), .dout(new_new_n1559__));
  or1   g0715(.dina(new_new_n2656__), .dinb(new_new_n2618__), .dout(new_new_n1560__));
  and1  g0716(.dina(new_new_n1559__), .dinb(new_new_n2556__), .dout(new_new_n1561__));
  or1   g0717(.dina(new_new_n1560__), .dinb(new_new_n2563__), .dout(new_new_n1562__));
  and1  g0718(.dina(new_new_n1561__), .dinb(new_new_n2625__), .dout(new_new_n1563__));
  or1   g0719(.dina(new_new_n1562__), .dinb(new_new_n2632__), .dout(new_new_n1564__));
  and1  g0720(.dina(new_new_n1563__), .dinb(new_new_n805__), .dout(new_new_n1565__));
  and1  g0721(.dina(new_new_n1564__), .dinb(new_new_n806__), .dout(new_new_n1566__));
  or1   g0722(.dina(new_new_n1566__), .dinb(new_new_n1565__), .dout(new_new_n1567__));
  and1  g0723(.dina(new_new_n2654__), .dinb(new_new_n2606__), .dout(new_new_n1568__));
  or1   g0724(.dina(new_new_n2655__), .dinb(new_new_n2607__), .dout(new_new_n1569__));
  and1  g0725(.dina(new_new_n1568__), .dinb(new_new_n2590__), .dout(new_new_n1570__));
  or1   g0726(.dina(new_new_n1569__), .dinb(new_new_n2596__), .dout(new_new_n1571__));
  and1  g0727(.dina(new_new_n1570__), .dinb(new_new_n2625__), .dout(new_new_n1572__));
  or1   g0728(.dina(new_new_n1571__), .dinb(new_new_n2632__), .dout(new_new_n1573__));
  and1  g0729(.dina(new_new_n1572__), .dinb(new_new_n807__), .dout(new_new_n1574__));
  and1  g0730(.dina(new_new_n1573__), .dinb(new_new_n808__), .dout(new_new_n1575__));
  or1   g0731(.dina(new_new_n1575__), .dinb(new_new_n1574__), .dout(new_new_n1576__));
  or1   g0732(.dina(new_new_n955__), .dinb(new_new_n941__), .dout(new_new_n1577__));
  or1   g0733(.dina(new_new_n956__), .dinb(new_new_n942__), .dout(new_new_n1578__));
  and1  g0734(.dina(new_new_n1578__), .dinb(new_new_n1577__), .dout(new_new_n1579__));
  or1   g0735(.dina(new_new_n952__), .dinb(new_new_n949__), .dout(new_new_n1580__));
  or1   g0736(.dina(new_new_n951__), .dinb(new_new_n950__), .dout(new_new_n1581__));
  and1  g0737(.dina(new_new_n1581__), .dinb(new_new_n1580__), .dout(new_new_n1582__));
  or1   g0738(.dina(new_new_n954__), .dinb(new_new_n947__), .dout(new_new_n1583__));
  or1   g0739(.dina(new_new_n953__), .dinb(new_new_n948__), .dout(new_new_n1584__));
  and1  g0740(.dina(new_new_n1584__), .dinb(new_new_n1583__), .dout(new_new_n1585__));
  or1   g0741(.dina(new_new_n957__), .dinb(new_new_n945__), .dout(new_new_n1586__));
  or1   g0742(.dina(new_new_n958__), .dinb(new_new_n946__), .dout(new_new_n1587__));
  and1  g0743(.dina(new_new_n1587__), .dinb(new_new_n1586__), .dout(new_new_n1588__));
  or1   g0744(.dina(new_new_n962__), .dinb(new_new_n943__), .dout(new_new_n1589__));
  or1   g0745(.dina(new_new_n961__), .dinb(new_new_n944__), .dout(new_new_n1590__));
  and1  g0746(.dina(new_new_n1590__), .dinb(new_new_n1589__), .dout(new_new_n1591__));
  or1   g0747(.dina(new_new_n959__), .dinb(new_new_n939__), .dout(new_new_n1592__));
  or1   g0748(.dina(new_new_n960__), .dinb(new_new_n940__), .dout(new_new_n1593__));
  and1  g0749(.dina(new_new_n1593__), .dinb(new_new_n1592__), .dout(new_new_n1594__));
  and1  g0750(.dina(new_new_n1582__), .dinb(new_new_n1579__), .dout(new_new_n1595__));
  and1  g0751(.dina(new_new_n1595__), .dinb(new_new_n1585__), .dout(new_new_n1596__));
  and1  g0752(.dina(new_new_n1596__), .dinb(new_new_n1588__), .dout(new_new_n1597__));
  and1  g0753(.dina(new_new_n1597__), .dinb(new_new_n996__), .dout(new_new_n1598__));
  and1  g0754(.dina(new_new_n1598__), .dinb(new_new_n1591__), .dout(new_new_n1599__));
  and1  g0755(.dina(new_new_n1599__), .dinb(new_new_n1594__), .dout(new_new_n1600__));
  and1  g0756(.dina(new_new_n1600__), .dinb(new_new_n998__), .dout(new_new_n1601__));
  or1   g0757(.dina(new_new_n1601__), .dinb(new_new_n1023__), .dout(new_new_n1602__));
  or1   g0758(.dina(new_new_n2659__), .dinb(new_new_n2661__), .dout(new_new_n1603__));
  or1   g0759(.dina(new_new_n1603__), .dinb(new_new_n2661__), .dout(new_new_n1604__));
  and1  g0760(.dina(new_new_n1024__), .dinb(new_new_n1020__), .dout(new_new_n1605__));
  and1  g0761(.dina(new_new_n1605__), .dinb(new_new_n1014__), .dout(new_new_n1606__));
  and1  g0762(.dina(new_new_n2649__), .dinb(new_new_n2557__), .dout(new_new_n1607__));
  and1  g0763(.dina(new_new_n1607__), .dinb(new_new_n2664__), .dout(new_new_n1608__));
  and1  g0764(.dina(new_new_n2654__), .dinb(new_new_n2581__), .dout(new_new_n1609__));
  and1  g0765(.dina(new_new_n1609__), .dinb(new_new_n2557__), .dout(new_new_n1610__));
  and1  g0766(.dina(new_new_n1610__), .dinb(new_new_n2664__), .dout(new_new_n1611__));
  and1  g0767(.dina(new_new_n2641__), .dinb(new_new_n2651__), .dout(new_new_n1612__));
  and1  g0768(.dina(new_new_n2670__), .dinb(new_new_n2545__), .dout(new_new_n1613__));
  and1  g0769(.dina(new_new_n1613__), .dinb(new_new_n2559__), .dout(new_new_n1614__));
  and1  g0770(.dina(new_new_n1614__), .dinb(new_new_n2665__), .dout(new_new_n1615__));
  and1  g0771(.dina(new_new_n2670__), .dinb(new_new_n2581__), .dout(new_new_n1616__));
  and1  g0772(.dina(new_new_n2671__), .dinb(new_new_n2589__), .dout(new_new_n1617__));
  and1  g0773(.dina(new_new_n1617__), .dinb(new_new_n2665__), .dout(new_new_n1618__));
  and1  g0774(.dina(new_new_n2671__), .dinb(new_new_n2600__), .dout(new_new_n1619__));
  and1  g0775(.dina(new_new_n1619__), .dinb(new_new_n2667__), .dout(new_new_n1620__));
  and1  g0776(.dina(new_new_n2669__), .dinb(new_new_n2606__), .dout(new_new_n1621__));
  and1  g0777(.dina(new_new_n1621__), .dinb(new_new_n2559__), .dout(new_new_n1622__));
  and1  g0778(.dina(new_new_n1622__), .dinb(new_new_n2667__), .dout(new_new_n1623__));
  and1  g0779(.dina(new_new_n1058__), .dinb(new_new_n997__), .dout(new_new_n1624__));
  and1  g0780(.dina(new_new_n1624__), .dinb(new_new_n2650__), .dout(new_new_n1625__));
  and1  g0781(.dina(new_new_n1625__), .dinb(new_new_n2582__), .dout(new_new_n1626__));
  and1  g0782(.dina(new_new_n1626__), .dinb(new_new_n2560__), .dout(new_new_n1627__));
  and1  g0783(.dina(new_new_n1627__), .dinb(new_new_n2668__), .dout(new_new_n1628__));
  and1  g0784(.dina(new_new_n1055__), .dinb(new_new_n995__), .dout(new_new_n1629__));
  and1  g0785(.dina(new_new_n1629__), .dinb(new_new_n2641__), .dout(new_new_n1630__));
  and1  g0786(.dina(new_new_n1630__), .dinb(new_new_n2582__), .dout(new_new_n1631__));
  and1  g0787(.dina(new_new_n1631__), .dinb(new_new_n2560__), .dout(new_new_n1632__));
  and1  g0788(.dina(new_new_n1632__), .dinb(new_new_n2668__), .dout(new_new_n1633__));
  or1   g0789(.dina(new_new_n1611__), .dinb(new_new_n1608__), .dout(new_new_n1634__));
  or1   g0790(.dina(new_new_n1634__), .dinb(new_new_n1615__), .dout(new_new_n1635__));
  or1   g0791(.dina(new_new_n1635__), .dinb(new_new_n1618__), .dout(new_new_n1636__));
  or1   g0792(.dina(new_new_n1636__), .dinb(new_new_n1620__), .dout(new_new_n1637__));
  or1   g0793(.dina(new_new_n1637__), .dinb(new_new_n1623__), .dout(new_new_n1638__));
  or1   g0794(.dina(new_new_n1638__), .dinb(new_new_n1628__), .dout(new_new_n1639__));
  or1   g0795(.dina(new_new_n1639__), .dinb(new_new_n1633__), .dout(new_new_n1640__));
  and1  g0796(.dina(new_new_n1228__), .dinb(new_new_n1226__), .dout(new_new_n1641__));
  or1   g0797(.dina(new_new_n1227__), .dinb(new_new_n1225__), .dout(new_new_n1642__));
  or1   g0798(.dina(new_new_n2674__), .dinb(new_new_n1640__), .dout(new_new_n1643__));
  or1   g0799(.dina(new_new_n2659__), .dinb(new_new_n892__), .dout(new_new_n1644__));
  or1   g0800(.dina(new_new_n1644__), .dinb(new_new_n1643__), .dout(new_new_n1645__));
  and1  g0801(.dina(new_new_n1645__), .dinb(new_new_n1604__), .dout(new_new_n1646__));
  and1  g0802(.dina(new_new_n1213__), .dinb(new_new_n1131__), .dout(new_new_n1647__));
  or1   g0803(.dina(new_new_n1214__), .dinb(new_new_n1132__), .dout(new_new_n1648__));
  and1  g0804(.dina(new_new_n1220__), .dinb(new_new_n1126__), .dout(new_new_n1649__));
  or1   g0805(.dina(new_new_n1219__), .dinb(new_new_n1125__), .dout(new_new_n1650__));
  and1  g0806(.dina(new_new_n1650__), .dinb(new_new_n1648__), .dout(new_new_n1651__));
  or1   g0807(.dina(new_new_n1649__), .dinb(new_new_n1647__), .dout(new_new_n1652__));
  and1  g0808(.dina(new_new_n2678__), .dinb(new_new_n2679__), .dout(new_new_n1653__));
  or1   g0809(.dina(new_new_n2680__), .dinb(new_new_n2681__), .dout(new_new_n1654__));
  and1  g0810(.dina(new_new_n2680__), .dinb(new_new_n2681__), .dout(new_new_n1655__));
  or1   g0811(.dina(new_new_n2678__), .dinb(new_new_n2679__), .dout(new_new_n1656__));
  and1  g0812(.dina(new_new_n1656__), .dinb(new_new_n1654__), .dout(new_new_n1657__));
  or1   g0813(.dina(new_new_n1655__), .dinb(new_new_n1653__), .dout(new_new_n1658__));
  and1  g0814(.dina(new_new_n925__), .dinb(new_new_n815__), .dout(new_new_n1659__));
  or1   g0815(.dina(new_new_n926__), .dinb(new_new_n816__), .dout(new_new_n1660__));
  and1  g0816(.dina(new_new_n1659__), .dinb(new_new_n2684__), .dout(new_new_n1661__));
  or1   g0817(.dina(new_new_n1660__), .dinb(new_new_n2689__), .dout(new_new_n1662__));
  and1  g0818(.dina(new_new_n1661__), .dinb(new_new_n2674__), .dout(new_new_n1663__));
  or1   g0819(.dina(new_new_n1662__), .dinb(new_new_n2694__), .dout(new_new_n1664__));
  and1  g0820(.dina(new_new_n1664__), .dinb(new_new_n1658__), .dout(new_new_n1665__));
  and1  g0821(.dina(new_new_n1663__), .dinb(new_new_n1657__), .dout(new_new_n1666__));
  or1   g0822(.dina(new_new_n1666__), .dinb(new_new_n1665__), .dout(new_new_n1667__));
  or1   g0823(.dina(new_new_n2699__), .dinb(new_new_n2660__), .dout(new_new_n1668__));
  and1  g0824(.dina(new_new_n2703__), .dinb(new_new_n1667__), .dout(new_new_n1669__));
  and1  g0825(.dina(new_new_n1206__), .dinb(new_new_n1204__), .dout(new_new_n1670__));
  or1   g0826(.dina(new_new_n1205__), .dinb(new_new_n1203__), .dout(new_new_n1671__));
  and1  g0827(.dina(new_new_n1215__), .dinb(new_new_n1133__), .dout(new_new_n1672__));
  or1   g0828(.dina(new_new_n1216__), .dinb(new_new_n1134__), .dout(new_new_n1673__));
  and1  g0829(.dina(new_new_n1222__), .dinb(new_new_n1128__), .dout(new_new_n1674__));
  or1   g0830(.dina(new_new_n1221__), .dinb(new_new_n1127__), .dout(new_new_n1675__));
  and1  g0831(.dina(new_new_n1675__), .dinb(new_new_n1673__), .dout(new_new_n1676__));
  or1   g0832(.dina(new_new_n1674__), .dinb(new_new_n1672__), .dout(new_new_n1677__));
  and1  g0833(.dina(new_new_n2706__), .dinb(new_new_n2707__), .dout(new_new_n1678__));
  or1   g0834(.dina(new_new_n2708__), .dinb(new_new_n2709__), .dout(new_new_n1679__));
  and1  g0835(.dina(new_new_n2708__), .dinb(new_new_n2709__), .dout(new_new_n1680__));
  or1   g0836(.dina(new_new_n2706__), .dinb(new_new_n2707__), .dout(new_new_n1681__));
  and1  g0837(.dina(new_new_n1681__), .dinb(new_new_n1679__), .dout(new_new_n1682__));
  or1   g0838(.dina(new_new_n1680__), .dinb(new_new_n1678__), .dout(new_new_n1683__));
  and1  g0839(.dina(new_new_n2684__), .dinb(new_new_n843__), .dout(new_new_n1684__));
  or1   g0840(.dina(new_new_n2689__), .dinb(new_new_n844__), .dout(new_new_n1685__));
  and1  g0841(.dina(new_new_n1684__), .dinb(new_new_n2675__), .dout(new_new_n1686__));
  or1   g0842(.dina(new_new_n1685__), .dinb(new_new_n2694__), .dout(new_new_n1687__));
  and1  g0843(.dina(new_new_n1687__), .dinb(new_new_n1683__), .dout(new_new_n1688__));
  and1  g0844(.dina(new_new_n1686__), .dinb(new_new_n1682__), .dout(new_new_n1689__));
  or1   g0845(.dina(new_new_n1689__), .dinb(new_new_n1688__), .dout(new_new_n1690__));
  and1  g0846(.dina(new_new_n1690__), .dinb(new_new_n2703__), .dout(new_new_n1691__));
  and1  g0847(.dina(new_new_n2685__), .dinb(new_new_n855__), .dout(new_new_n1692__));
  or1   g0848(.dina(new_new_n2690__), .dinb(new_new_n856__), .dout(new_new_n1693__));
  and1  g0849(.dina(new_new_n1692__), .dinb(new_new_n2675__), .dout(new_new_n1694__));
  or1   g0850(.dina(new_new_n1693__), .dinb(new_new_n2695__), .dout(new_new_n1695__));
  and1  g0851(.dina(new_new_n1695__), .dinb(new_new_n930__), .dout(new_new_n1696__));
  and1  g0852(.dina(new_new_n1694__), .dinb(new_new_n929__), .dout(new_new_n1697__));
  or1   g0853(.dina(new_new_n1697__), .dinb(new_new_n1696__), .dout(new_new_n1698__));
  and1  g0854(.dina(new_new_n1698__), .dinb(new_new_n2704__), .dout(new_new_n1699__));
  and1  g0855(.dina(new_new_n2685__), .dinb(new_new_n861__), .dout(new_new_n1700__));
  or1   g0856(.dina(new_new_n2690__), .dinb(new_new_n862__), .dout(new_new_n1701__));
  and1  g0857(.dina(new_new_n1700__), .dinb(new_new_n2677__), .dout(new_new_n1702__));
  or1   g0858(.dina(new_new_n1701__), .dinb(new_new_n2695__), .dout(new_new_n1703__));
  and1  g0859(.dina(new_new_n1703__), .dinb(new_new_n928__), .dout(new_new_n1704__));
  and1  g0860(.dina(new_new_n1702__), .dinb(new_new_n927__), .dout(new_new_n1705__));
  or1   g0861(.dina(new_new_n1705__), .dinb(new_new_n1704__), .dout(new_new_n1706__));
  and1  g0862(.dina(new_new_n1706__), .dinb(new_new_n2704__), .dout(new_new_n1707__));
  and1  g0863(.dina(new_new_n923__), .dinb(new_new_n823__), .dout(new_new_n1708__));
  or1   g0864(.dina(new_new_n924__), .dinb(new_new_n824__), .dout(new_new_n1709__));
  and1  g0865(.dina(new_new_n1708__), .dinb(new_new_n2686__), .dout(new_new_n1710__));
  or1   g0866(.dina(new_new_n1709__), .dinb(new_new_n2691__), .dout(new_new_n1711__));
  and1  g0867(.dina(new_new_n1710__), .dinb(new_new_n2677__), .dout(new_new_n1712__));
  or1   g0868(.dina(new_new_n1711__), .dinb(new_new_n2696__), .dout(new_new_n1713__));
  and1  g0869(.dina(new_new_n1713__), .dinb(new_new_n931__), .dout(new_new_n1714__));
  and1  g0870(.dina(new_new_n1712__), .dinb(new_new_n932__), .dout(new_new_n1715__));
  or1   g0871(.dina(new_new_n1715__), .dinb(new_new_n1714__), .dout(new_new_n1716__));
  and1  g0872(.dina(new_new_n1716__), .dinb(new_new_n2705__), .dout(new_new_n1717__));
  and1  g0873(.dina(new_new_n1158__), .dinb(new_new_n1156__), .dout(new_new_n1718__));
  or1   g0874(.dina(new_new_n1157__), .dinb(new_new_n1155__), .dout(new_new_n1719__));
  and1  g0875(.dina(new_new_n1718__), .dinb(new_new_n1160__), .dout(new_new_n1720__));
  or1   g0876(.dina(new_new_n1719__), .dinb(new_new_n1159__), .dout(new_new_n1721__));
  and1  g0877(.dina(new_new_n1720__), .dinb(new_new_n1162__), .dout(new_new_n1722__));
  or1   g0878(.dina(new_new_n1721__), .dinb(new_new_n1161__), .dout(new_new_n1723__));
  and1  g0879(.dina(new_new_n1722__), .dinb(new_new_n1146__), .dout(new_new_n1724__));
  or1   g0880(.dina(new_new_n1723__), .dinb(new_new_n1145__), .dout(new_new_n1725__));
  and1  g0881(.dina(new_new_n1724__), .dinb(new_new_n1148__), .dout(new_new_n1726__));
  or1   g0882(.dina(new_new_n1725__), .dinb(new_new_n1147__), .dout(new_new_n1727__));
  and1  g0883(.dina(new_new_n1726__), .dinb(new_new_n1150__), .dout(new_new_n1728__));
  or1   g0884(.dina(new_new_n1727__), .dinb(new_new_n1149__), .dout(new_new_n1729__));
  and1  g0885(.dina(new_new_n1728__), .dinb(new_new_n1152__), .dout(new_new_n1730__));
  or1   g0886(.dina(new_new_n1729__), .dinb(new_new_n1151__), .dout(new_new_n1731__));
  and1  g0887(.dina(new_new_n1731__), .dinb(new_new_n2711__), .dout(new_new_n1732__));
  or1   g0888(.dina(new_new_n1730__), .dinb(new_new_n2699__), .dout(new_new_n1733__));
  and1  g0889(.dina(new_new_n1207__), .dinb(new_new_n1202__), .dout(new_new_n1734__));
  or1   g0890(.dina(new_new_n1208__), .dinb(new_new_n1201__), .dout(new_new_n1735__));
  and1  g0891(.dina(new_new_n2713__), .dinb(new_new_n1016__), .dout(new_new_n1736__));
  or1   g0892(.dina(new_new_n2714__), .dinb(new_new_n1015__), .dout(new_new_n1737__));
  and1  g0893(.dina(new_new_n1737__), .dinb(new_new_n1734__), .dout(new_new_n1738__));
  or1   g0894(.dina(new_new_n1736__), .dinb(new_new_n1735__), .dout(new_new_n1739__));
  and1  g0895(.dina(new_new_n2715__), .dinb(new_new_n2716__), .dout(new_new_n1740__));
  or1   g0896(.dina(new_new_n2717__), .dinb(new_new_n2718__), .dout(new_new_n1741__));
  and1  g0897(.dina(new_new_n2717__), .dinb(new_new_n2718__), .dout(new_new_n1742__));
  or1   g0898(.dina(new_new_n2715__), .dinb(new_new_n2716__), .dout(new_new_n1743__));
  and1  g0899(.dina(new_new_n1743__), .dinb(new_new_n1741__), .dout(new_new_n1744__));
  or1   g0900(.dina(new_new_n1742__), .dinb(new_new_n1740__), .dout(new_new_n1745__));
  and1  g0901(.dina(new_new_n869__), .dinb(new_new_n829__), .dout(new_new_n1746__));
  or1   g0902(.dina(new_new_n870__), .dinb(new_new_n830__), .dout(new_new_n1747__));
  and1  g0903(.dina(new_new_n1747__), .dinb(new_new_n2711__), .dout(new_new_n1748__));
  or1   g0904(.dina(new_new_n1746__), .dinb(new_new_n2698__), .dout(new_new_n1749__));
  and1  g0905(.dina(new_new_n1749__), .dinb(new_new_n1745__), .dout(new_new_n1750__));
  and1  g0906(.dina(new_new_n1748__), .dinb(new_new_n1744__), .dout(new_new_n1751__));
  or1   g0907(.dina(new_new_n1751__), .dinb(new_new_n1750__), .dout(new_new_n1752__));
  and1  g0908(.dina(new_new_n1164__), .dinb(new_new_n1154__), .dout(new_new_n1753__));
  or1   g0909(.dina(new_new_n1163__), .dinb(new_new_n1153__), .dout(new_new_n1754__));
  and1  g0910(.dina(new_new_n1753__), .dinb(new_new_n1138__), .dout(new_new_n1755__));
  or1   g0911(.dina(new_new_n1754__), .dinb(new_new_n1137__), .dout(new_new_n1756__));
  and1  g0912(.dina(new_new_n1755__), .dinb(new_new_n1140__), .dout(new_new_n1757__));
  or1   g0913(.dina(new_new_n1756__), .dinb(new_new_n1139__), .dout(new_new_n1758__));
  and1  g0914(.dina(new_new_n1757__), .dinb(new_new_n1142__), .dout(new_new_n1759__));
  or1   g0915(.dina(new_new_n1758__), .dinb(new_new_n1141__), .dout(new_new_n1760__));
  and1  g0916(.dina(new_new_n1759__), .dinb(new_new_n1144__), .dout(new_new_n1761__));
  or1   g0917(.dina(new_new_n1760__), .dinb(new_new_n1143__), .dout(new_new_n1762__));
  and1  g0918(.dina(new_new_n1761__), .dinb(new_new_n1166__), .dout(new_new_n1763__));
  or1   g0919(.dina(new_new_n1762__), .dinb(new_new_n1165__), .dout(new_new_n1764__));
  and1  g0920(.dina(new_new_n1763__), .dinb(new_new_n1168__), .dout(new_new_n1765__));
  or1   g0921(.dina(new_new_n1764__), .dinb(new_new_n1167__), .dout(new_new_n1766__));
  and1  g0922(.dina(new_new_n1766__), .dinb(new_new_n2712__), .dout(new_new_n1767__));
  or1   g0923(.dina(new_new_n1765__), .dinb(new_new_n2700__), .dout(new_new_n1768__));
  and1  g0924(.dina(new_new_n2713__), .dinb(new_new_n1018__), .dout(new_new_n1769__));
  or1   g0925(.dina(new_new_n2714__), .dinb(new_new_n1017__), .dout(new_new_n1770__));
  and1  g0926(.dina(new_new_n1211__), .dinb(new_new_n1210__), .dout(new_new_n1771__));
  or1   g0927(.dina(new_new_n1212__), .dinb(new_new_n1209__), .dout(new_new_n1772__));
  and1  g0928(.dina(new_new_n1771__), .dinb(new_new_n1770__), .dout(new_new_n1773__));
  or1   g0929(.dina(new_new_n1772__), .dinb(new_new_n1769__), .dout(new_new_n1774__));
  and1  g0930(.dina(new_new_n2719__), .dinb(new_new_n2720__), .dout(new_new_n1775__));
  or1   g0931(.dina(new_new_n2721__), .dinb(new_new_n2722__), .dout(new_new_n1776__));
  and1  g0932(.dina(new_new_n2721__), .dinb(new_new_n2722__), .dout(new_new_n1777__));
  or1   g0933(.dina(new_new_n2719__), .dinb(new_new_n2720__), .dout(new_new_n1778__));
  and1  g0934(.dina(new_new_n1778__), .dinb(new_new_n1776__), .dout(new_new_n1779__));
  or1   g0935(.dina(new_new_n1777__), .dinb(new_new_n1775__), .dout(new_new_n1780__));
  and1  g0936(.dina(new_new_n877__), .dinb(new_new_n833__), .dout(new_new_n1781__));
  or1   g0937(.dina(new_new_n878__), .dinb(new_new_n834__), .dout(new_new_n1782__));
  and1  g0938(.dina(new_new_n1782__), .dinb(new_new_n2712__), .dout(new_new_n1783__));
  or1   g0939(.dina(new_new_n1781__), .dinb(new_new_n2700__), .dout(new_new_n1784__));
  and1  g0940(.dina(new_new_n1784__), .dinb(new_new_n1780__), .dout(new_new_n1785__));
  and1  g0941(.dina(new_new_n1783__), .dinb(new_new_n1779__), .dout(new_new_n1786__));
  or1   g0942(.dina(new_new_n1786__), .dinb(new_new_n1785__), .dout(new_new_n1787__));
  and1  g0943(.dina(new_new_n1218__), .dinb(new_new_n1135__), .dout(new_new_n1788__));
  or1   g0944(.dina(new_new_n1217__), .dinb(new_new_n1136__), .dout(new_new_n1789__));
  and1  g0945(.dina(new_new_n1224__), .dinb(new_new_n1129__), .dout(new_new_n1790__));
  or1   g0946(.dina(new_new_n1223__), .dinb(new_new_n1130__), .dout(new_new_n1791__));
  and1  g0947(.dina(new_new_n1791__), .dinb(new_new_n1789__), .dout(new_new_n1792__));
  or1   g0948(.dina(new_new_n1790__), .dinb(new_new_n1788__), .dout(new_new_n1793__));
  and1  g0949(.dina(new_new_n2686__), .dinb(new_new_n849__), .dout(new_new_n1794__));
  or1   g0950(.dina(new_new_n2691__), .dinb(new_new_n850__), .dout(new_new_n1795__));
  and1  g0951(.dina(new_new_n1794__), .dinb(new_new_n2676__), .dout(new_new_n1796__));
  or1   g0952(.dina(new_new_n1795__), .dinb(new_new_n2696__), .dout(new_new_n1797__));
  and1  g0953(.dina(new_new_n2723__), .dinb(new_new_n2724__), .dout(new_new_n1798__));
  or1   g0954(.dina(new_new_n2725__), .dinb(new_new_n2726__), .dout(new_new_n1799__));
  and1  g0955(.dina(new_new_n2725__), .dinb(new_new_n2726__), .dout(new_new_n1800__));
  or1   g0956(.dina(new_new_n2723__), .dinb(new_new_n2724__), .dout(new_new_n1801__));
  and1  g0957(.dina(new_new_n1801__), .dinb(new_new_n1799__), .dout(new_new_n1802__));
  or1   g0958(.dina(new_new_n1800__), .dinb(new_new_n1798__), .dout(new_new_n1803__));
  and1  g0959(.dina(new_new_n2727__), .dinb(new_new_n2728__), .dout(new_new_n1804__));
  or1   g0960(.dina(new_new_n2729__), .dinb(new_new_n2730__), .dout(new_new_n1805__));
  and1  g0961(.dina(new_new_n2729__), .dinb(new_new_n2730__), .dout(new_new_n1806__));
  or1   g0962(.dina(new_new_n2727__), .dinb(new_new_n2728__), .dout(new_new_n1807__));
  and1  g0963(.dina(new_new_n1807__), .dinb(new_new_n1805__), .dout(new_new_n1808__));
  or1   g0964(.dina(new_new_n1806__), .dinb(new_new_n1804__), .dout(new_new_n1809__));
  and1  g0965(.dina(new_new_n1808__), .dinb(new_new_n1803__), .dout(new_new_n1810__));
  and1  g0966(.dina(new_new_n1809__), .dinb(new_new_n1802__), .dout(new_new_n1811__));
  or1   g0967(.dina(new_new_n1811__), .dinb(new_new_n1810__), .dout(new_new_n1812__));
  and1  g0968(.dina(new_new_n1812__), .dinb(new_new_n2705__), .dout(new_new_n1813__));
  and1  g0969(.dina(new_new_n2732__), .dinb(new_new_n2733__), .dout(new_new_n1814__));
  or1   g0970(.dina(new_new_n2734__), .dinb(new_new_n1012__), .dout(new_new_n1815__));
  and1  g0971(.dina(new_new_n2736__), .dinb(new_new_n2737__), .dout(new_new_n1816__));
  or1   g0972(.dina(new_new_n2738__), .dinb(new_new_n1112__), .dout(new_new_n1817__));
  and1  g0973(.dina(new_new_n2739__), .dinb(new_new_n2742__), .dout(new_new_n1818__));
  or1   g0974(.dina(new_new_n1276__), .dinb(new_new_n2747__), .dout(new_new_n1819__));
  and1  g0975(.dina(new_new_n2750__), .dinb(new_new_n2742__), .dout(new_new_n1820__));
  or1   g0976(.dina(new_new_n1278__), .dinb(new_new_n2747__), .dout(new_new_n1821__));
  and1  g0977(.dina(new_new_n1282__), .dinb(new_new_n2743__), .dout(new_new_n1822__));
  or1   g0978(.dina(new_new_n2751__), .dinb(new_new_n2748__), .dout(new_new_n1823__));
  and1  g0979(.dina(new_new_n1284__), .dinb(new_new_n2743__), .dout(new_new_n1824__));
  or1   g0980(.dina(new_new_n1283__), .dinb(new_new_n2748__), .dout(new_new_n1825__));
  and1  g0981(.dina(new_new_n1288__), .dinb(new_new_n2744__), .dout(new_new_n1826__));
  or1   g0982(.dina(new_new_n1287__), .dinb(new_new_n2749__), .dout(new_new_n1827__));
  and1  g0983(.dina(new_new_n1279__), .dinb(new_new_n2744__), .dout(new_new_n1828__));
  or1   g0984(.dina(new_new_n1280__), .dinb(new_new_n2749__), .dout(new_new_n1829__));
  and1  g0985(.dina(new_new_n2732__), .dinb(new_new_n983__), .dout(new_new_n1830__));
  or1   g0986(.dina(new_new_n2734__), .dinb(new_new_n984__), .dout(new_new_n1831__));
  and1  g0987(.dina(new_new_n2736__), .dinb(new_new_n1029__), .dout(new_new_n1832__));
  or1   g0988(.dina(new_new_n2738__), .dinb(new_new_n1030__), .dout(new_new_n1833__));
  or1   g0989(.dina(new_new_n1199__), .dinb(new_new_n976__), .dout(new_new_n1834__));
  and1  g0990(.dina(new_new_n2752__), .dinb(new_new_n1182__), .dout(new_new_n1835__));
  or1   g0991(.dina(new_new_n1342__), .dinb(new_new_n1181__), .dout(new_new_n1836__));
  and1  g0992(.dina(new_new_n1835__), .dinb(new_new_n2754__), .dout(new_new_n1837__));
  or1   g0993(.dina(new_new_n1836__), .dinb(new_new_n2757__), .dout(new_new_n1838__));
  and1  g0994(.dina(new_new_n2759__), .dinb(new_new_n2754__), .dout(new_new_n1839__));
  or1   g0995(.dina(new_new_n1316__), .dinb(new_new_n2757__), .dout(new_new_n1840__));
  or1   g0996(.dina(new_new_n2760__), .dinb(new_new_n2761__), .dout(new_new_n1841__));
  or1   g0997(.dina(new_new_n1826__), .dinb(new_new_n1815__), .dout(new_new_n1842__));
  and1  g0998(.dina(new_new_n1842__), .dinb(new_new_n1841__), .dout(new_new_n1843__));
  or1   g0999(.dina(new_new_n1829__), .dinb(new_new_n2763__), .dout(new_new_n1844__));
  or1   g1000(.dina(new_new_n2764__), .dinb(new_new_n1250__), .dout(new_new_n1845__));
  and1  g1001(.dina(new_new_n1845__), .dinb(new_new_n1844__), .dout(new_new_n1846__));
  and1  g1002(.dina(new_new_n2766__), .dinb(new_new_n2767__), .dout(new_new_n1847__));
  and1  g1003(.dina(new_new_n2769__), .dinb(new_new_n2770__), .dout(new_new_n1848__));
  and1  g1004(.dina(new_new_n2771__), .dinb(new_new_n868__), .dout(new_new_n1849__));
  and1  g1005(.dina(new_new_n1849__), .dinb(new_new_n2773__), .dout(new_new_n1850__));
  and1  g1006(.dina(new_new_n1850__), .dinb(new_new_n2775__), .dout(new_new_n1851__));
  and1  g1007(.dina(new_new_n2773__), .dinb(new_new_n890__), .dout(new_new_n1852__));
  and1  g1008(.dina(new_new_n1852__), .dinb(new_new_n2775__), .dout(new_new_n1853__));
  or1   g1009(.dina(new_new_n2777__), .dinb(new_new_n1851__), .dout(new_new_n1854__));
  and1  g1010(.dina(new_new_n2771__), .dinb(new_new_n876__), .dout(new_new_n1855__));
  and1  g1011(.dina(new_new_n1855__), .dinb(new_new_n2772__), .dout(new_new_n1856__));
  and1  g1012(.dina(new_new_n1856__), .dinb(new_new_n2776__), .dout(new_new_n1857__));
  or1   g1013(.dina(new_new_n1857__), .dinb(new_new_n2777__), .dout(new_new_n1858__));
  or1   g1014(.dina(new_new_n2766__), .dinb(new_new_n1831__), .dout(new_new_n1859__));
  or1   g1015(.dina(new_new_n2769__), .dinb(new_new_n1833__), .dout(new_new_n1860__));
  or1   g1016(.dina(new_new_n2778__), .dinb(new_new_n2779__), .dout(new_new_n1861__));
  or1   g1017(.dina(new_new_n1822__), .dinb(new_new_n1817__), .dout(new_new_n1862__));
  and1  g1018(.dina(new_new_n1862__), .dinb(new_new_n1861__), .dout(new_new_n1863__));
  or1   g1019(.dina(new_new_n2780__), .dinb(new_new_n2782__), .dout(new_new_n1864__));
  or1   g1020(.dina(new_new_n1824__), .dinb(new_new_n1252__), .dout(new_new_n1865__));
  and1  g1021(.dina(new_new_n1865__), .dinb(new_new_n1864__), .dout(new_new_n1866__));
  and1  g1022(.dina(new_new_n1866__), .dinb(new_new_n1863__), .dout(new_new_n1867__));
  or1   g1023(.dina(new_new_n1819__), .dinb(new_new_n2784__), .dout(new_new_n1868__));
  or1   g1024(.dina(new_new_n2785__), .dinb(new_new_n1256__), .dout(new_new_n1869__));
  and1  g1025(.dina(new_new_n1869__), .dinb(new_new_n1868__), .dout(new_new_n1870__));
  or1   g1026(.dina(new_new_n1821__), .dinb(new_new_n2787__), .dout(new_new_n1871__));
  or1   g1027(.dina(new_new_n2788__), .dinb(new_new_n1254__), .dout(new_new_n1872__));
  and1  g1028(.dina(new_new_n1872__), .dinb(new_new_n1871__), .dout(new_new_n1873__));
  and1  g1029(.dina(new_new_n1873__), .dinb(new_new_n1870__), .dout(new_new_n1874__));
  and1  g1030(.dina(new_new_n1340__), .dinb(new_new_n1337__), .dout(new_new_n1875__));
  or1   g1031(.dina(new_new_n1339__), .dinb(new_new_n1338__), .dout(new_new_n1876__));
  and1  g1032(.dina(new_new_n2789__), .dinb(new_new_n2790__), .dout(new_new_n1877__));
  or1   g1033(.dina(new_new_n2791__), .dinb(new_new_n2793__), .dout(new_new_n1878__));
  and1  g1034(.dina(new_new_n2791__), .dinb(new_new_n2793__), .dout(new_new_n1879__));
  or1   g1035(.dina(new_new_n2789__), .dinb(new_new_n2790__), .dout(new_new_n1880__));
  and1  g1036(.dina(new_new_n1880__), .dinb(new_new_n1878__), .dout(new_new_n1881__));
  or1   g1037(.dina(new_new_n1879__), .dinb(new_new_n1877__), .dout(new_new_n1882__));
  and1  g1038(.dina(new_new_n988__), .dinb(new_new_n985__), .dout(new_new_n1883__));
  and1  g1039(.dina(new_new_n987__), .dinb(new_new_n986__), .dout(new_new_n1884__));
  or1   g1040(.dina(new_new_n1884__), .dinb(new_new_n1883__), .dout(new_new_n1885__));
  and1  g1041(.dina(new_new_n1005__), .dinb(new_new_n1000__), .dout(new_new_n1886__));
  and1  g1042(.dina(new_new_n1006__), .dinb(new_new_n999__), .dout(new_new_n1887__));
  or1   g1043(.dina(new_new_n1887__), .dinb(new_new_n1886__), .dout(new_new_n1888__));
  and1  g1044(.dina(new_new_n1003__), .dinb(new_new_n1002__), .dout(new_new_n1889__));
  and1  g1045(.dina(new_new_n1004__), .dinb(new_new_n1001__), .dout(new_new_n1890__));
  or1   g1046(.dina(new_new_n1890__), .dinb(new_new_n1889__), .dout(new_new_n1891__));
  and1  g1047(.dina(new_new_n2795__), .dinb(new_new_n2797__), .dout(new_new_n1892__));
  and1  g1048(.dina(new_new_n1892__), .dinb(new_new_n2800__), .dout(new_new_n1893__));
  and1  g1049(.dina(new_new_n1893__), .dinb(new_new_n2806__), .dout(new_new_n1894__));
  and1  g1050(.dina(new_new_n1894__), .dinb(new_new_n2811__), .dout(new_new_n1895__));
  and1  g1051(.dina(new_new_n2814__), .dinb(new_new_n2816__), .dout(new_new_n1896__));
  and1  g1052(.dina(new_new_n1896__), .dinb(new_new_n2800__), .dout(new_new_n1897__));
  and1  g1053(.dina(new_new_n1897__), .dinb(new_new_n2806__), .dout(new_new_n1898__));
  and1  g1054(.dina(new_new_n2817__), .dinb(new_new_n2819__), .dout(new_new_n1899__));
  and1  g1055(.dina(new_new_n2817__), .dinb(new_new_n2811__), .dout(new_new_n1900__));
  and1  g1056(.dina(new_new_n2795__), .dinb(new_new_n2814__), .dout(new_new_n1901__));
  and1  g1057(.dina(new_new_n1901__), .dinb(new_new_n2801__), .dout(new_new_n1902__));
  and1  g1058(.dina(new_new_n1902__), .dinb(new_new_n2807__), .dout(new_new_n1903__));
  and1  g1059(.dina(new_new_n2820__), .dinb(new_new_n2819__), .dout(new_new_n1904__));
  and1  g1060(.dina(new_new_n2820__), .dinb(new_new_n2812__), .dout(new_new_n1905__));
  and1  g1061(.dina(new_new_n2821__), .dinb(new_new_n2822__), .dout(new_new_n1906__));
  or1   g1062(.dina(new_new_n2823__), .dinb(new_new_n2824__), .dout(new_new_n1907__));
  and1  g1063(.dina(new_new_n2823__), .dinb(new_new_n2824__), .dout(new_new_n1908__));
  or1   g1064(.dina(new_new_n2821__), .dinb(new_new_n2822__), .dout(new_new_n1909__));
  and1  g1065(.dina(new_new_n1909__), .dinb(new_new_n1907__), .dout(new_new_n1910__));
  or1   g1066(.dina(new_new_n1908__), .dinb(new_new_n1906__), .dout(new_new_n1911__));
  and1  g1067(.dina(new_new_n1911__), .dinb(new_new_n2826__), .dout(new_new_n1912__));
  and1  g1068(.dina(new_new_n1910__), .dinb(new_new_n2829__), .dout(new_new_n1913__));
  or1   g1069(.dina(new_new_n1913__), .dinb(new_new_n1912__), .dout(new_new_n1914__));
  and1  g1070(.dina(new_new_n2831__), .dinb(new_new_n2832__), .dout(new_new_n1915__));
  or1   g1071(.dina(new_new_n2833__), .dinb(new_new_n2834__), .dout(new_new_n1916__));
  and1  g1072(.dina(new_new_n2833__), .dinb(new_new_n2834__), .dout(new_new_n1917__));
  or1   g1073(.dina(new_new_n2831__), .dinb(new_new_n2832__), .dout(new_new_n1918__));
  and1  g1074(.dina(new_new_n1918__), .dinb(new_new_n1916__), .dout(new_new_n1919__));
  or1   g1075(.dina(new_new_n1917__), .dinb(new_new_n1915__), .dout(new_new_n1920__));
  and1  g1076(.dina(new_new_n1920__), .dinb(new_new_n2836__), .dout(new_new_n1921__));
  and1  g1077(.dina(new_new_n1919__), .dinb(new_new_n2838__), .dout(new_new_n1922__));
  or1   g1078(.dina(new_new_n1922__), .dinb(new_new_n1921__), .dout(new_new_n1923__));
  and1  g1079(.dina(new_new_n1421__), .dinb(new_new_n1383__), .dout(new_new_n1924__));
  or1   g1080(.dina(new_new_n1422__), .dinb(new_new_n1384__), .dout(new_new_n1925__));
  and1  g1081(.dina(new_new_n1414__), .dinb(new_new_n1392__), .dout(new_new_n1926__));
  or1   g1082(.dina(new_new_n1413__), .dinb(new_new_n1391__), .dout(new_new_n1927__));
  and1  g1083(.dina(new_new_n1927__), .dinb(new_new_n1925__), .dout(new_new_n1928__));
  or1   g1084(.dina(new_new_n1926__), .dinb(new_new_n1924__), .dout(new_new_n1929__));
  and1  g1085(.dina(new_new_n1929__), .dinb(new_new_n2840__), .dout(new_new_n1930__));
  and1  g1086(.dina(new_new_n1928__), .dinb(new_new_n2841__), .dout(new_new_n1931__));
  or1   g1087(.dina(new_new_n1931__), .dinb(new_new_n1930__), .dout(new_new_n1932__));
  and1  g1088(.dina(new_new_n1423__), .dinb(new_new_n1389__), .dout(new_new_n1933__));
  or1   g1089(.dina(new_new_n1424__), .dinb(new_new_n1390__), .dout(new_new_n1934__));
  and1  g1090(.dina(new_new_n1420__), .dinb(new_new_n1394__), .dout(new_new_n1935__));
  or1   g1091(.dina(new_new_n1419__), .dinb(new_new_n1393__), .dout(new_new_n1936__));
  and1  g1092(.dina(new_new_n1936__), .dinb(new_new_n1934__), .dout(new_new_n1937__));
  or1   g1093(.dina(new_new_n1935__), .dinb(new_new_n1933__), .dout(new_new_n1938__));
  and1  g1094(.dina(new_new_n1938__), .dinb(new_new_n2826__), .dout(new_new_n1939__));
  and1  g1095(.dina(new_new_n1937__), .dinb(new_new_n2829__), .dout(new_new_n1940__));
  or1   g1096(.dina(new_new_n1940__), .dinb(new_new_n1939__), .dout(new_new_n1941__));
  and1  g1097(.dina(new_new_n991__), .dinb(new_new_n989__), .dout(new_new_n1942__));
  and1  g1098(.dina(new_new_n992__), .dinb(new_new_n990__), .dout(new_new_n1943__));
  or1   g1099(.dina(new_new_n1943__), .dinb(new_new_n1942__), .dout(new_new_n1944__));
  or1   g1100(.dina(new_new_n2842__), .dinb(new_new_n2843__), .dout(new_new_n1945__));
  and1  g1101(.dina(new_new_n1009__), .dinb(new_new_n979__), .dout(new_new_n1946__));
  and1  g1102(.dina(new_new_n1010__), .dinb(new_new_n980__), .dout(new_new_n1947__));
  or1   g1103(.dina(new_new_n1947__), .dinb(new_new_n1946__), .dout(new_new_n1948__));
  or1   g1104(.dina(new_new_n2844__), .dinb(new_new_n2845__), .dout(new_new_n1949__));
  and1  g1105(.dina(new_new_n2844__), .dinb(new_new_n2845__), .dout(new_new_n1950__));
  and1  g1106(.dina(new_new_n2842__), .dinb(new_new_n2843__), .dout(new_new_n1951__));
  and1  g1107(.dina(new_new_n1265__), .dinb(new_new_n1264__), .dout(new_new_n1952__));
  or1   g1108(.dina(new_new_n1266__), .dinb(new_new_n1263__), .dout(new_new_n1953__));
  and1  g1109(.dina(new_new_n2846__), .dinb(new_new_n2847__), .dout(new_new_n1954__));
  or1   g1110(.dina(new_new_n2848__), .dinb(new_new_n2849__), .dout(new_new_n1955__));
  and1  g1111(.dina(new_new_n2848__), .dinb(new_new_n2849__), .dout(new_new_n1956__));
  or1   g1112(.dina(new_new_n2846__), .dinb(new_new_n2847__), .dout(new_new_n1957__));
  and1  g1113(.dina(new_new_n1957__), .dinb(new_new_n1955__), .dout(new_new_n1958__));
  or1   g1114(.dina(new_new_n1956__), .dinb(new_new_n1954__), .dout(new_new_n1959__));
  and1  g1115(.dina(new_new_n1958__), .dinb(new_new_n993__), .dout(new_new_n1960__));
  and1  g1116(.dina(new_new_n1959__), .dinb(new_new_n994__), .dout(new_new_n1961__));
  or1   g1117(.dina(new_new_n1961__), .dinb(new_new_n1960__), .dout(new_new_n1962__));
  and1  g1118(.dina(new_new_n982__), .dinb(new_new_n973__), .dout(new_new_n1963__));
  and1  g1119(.dina(new_new_n981__), .dinb(new_new_n974__), .dout(new_new_n1964__));
  or1   g1120(.dina(new_new_n1964__), .dinb(new_new_n1963__), .dout(new_new_n1965__));
  and1  g1121(.dina(new_new_n2850__), .dinb(new_new_n2851__), .dout(new_new_n1966__));
  or1   g1122(.dina(new_new_n2850__), .dinb(new_new_n2851__), .dout(new_new_n1967__));
  or1   g1123(.dina(new_new_n2854__), .dinb(new_new_n2857__), .dout(new_new_n1968__));
  or1   g1124(.dina(new_new_n1968__), .dinb(new_new_n2860__), .dout(new_new_n1969__));
  or1   g1125(.dina(new_new_n1969__), .dinb(new_new_n2860__), .dout(new_new_n1970__));
  or1   g1126(.dina(new_new_n1970__), .dinb(new_new_n2861__), .dout(new_new_n1971__));
  or1   g1127(.dina(new_new_n1971__), .dinb(new_new_n2861__), .dout(new_new_n1972__));
  or1   g1128(.dina(new_new_n1972__), .dinb(new_new_n2854__), .dout(new_new_n1973__));
  or1   g1129(.dina(new_new_n1973__), .dinb(new_new_n2855__), .dout(new_new_n1974__));
  or1   g1130(.dina(new_new_n2867__), .dinb(new_new_n2871__), .dout(new_new_n1975__));
  or1   g1131(.dina(new_new_n1975__), .dinb(new_new_n2871__), .dout(new_new_n1976__));
  or1   g1132(.dina(new_new_n1976__), .dinb(new_new_n2872__), .dout(new_new_n1977__));
  or1   g1133(.dina(new_new_n1977__), .dinb(new_new_n2872__), .dout(new_new_n1978__));
  and1  g1134(.dina(new_new_n2876__), .dinb(new_new_n2878__), .dout(new_new_n1979__));
  or1   g1135(.dina(new_new_n2879__), .dinb(new_new_n2880__), .dout(new_new_n1980__));
  and1  g1136(.dina(new_new_n2879__), .dinb(new_new_n2880__), .dout(new_new_n1981__));
  or1   g1137(.dina(new_new_n2876__), .dinb(new_new_n2878__), .dout(new_new_n1982__));
  and1  g1138(.dina(new_new_n1982__), .dinb(new_new_n1980__), .dout(new_new_n1983__));
  or1   g1139(.dina(new_new_n1981__), .dinb(new_new_n1979__), .dout(new_new_n1984__));
  and1  g1140(.dina(new_new_n1984__), .dinb(new_new_n2840__), .dout(new_new_n1985__));
  and1  g1141(.dina(new_new_n1983__), .dinb(new_new_n2841__), .dout(new_new_n1986__));
  or1   g1142(.dina(new_new_n1986__), .dinb(new_new_n1985__), .dout(new_new_n1987__));
  and1  g1143(.dina(new_new_n2881__), .dinb(new_new_n2882__), .dout(new_new_n1988__));
  or1   g1144(.dina(new_new_n2883__), .dinb(new_new_n2884__), .dout(new_new_n1989__));
  and1  g1145(.dina(new_new_n2883__), .dinb(new_new_n2884__), .dout(new_new_n1990__));
  or1   g1146(.dina(new_new_n2881__), .dinb(new_new_n2882__), .dout(new_new_n1991__));
  and1  g1147(.dina(new_new_n1991__), .dinb(new_new_n1989__), .dout(new_new_n1992__));
  or1   g1148(.dina(new_new_n1990__), .dinb(new_new_n1988__), .dout(new_new_n1993__));
  and1  g1149(.dina(new_new_n1993__), .dinb(new_new_n2886__), .dout(new_new_n1994__));
  and1  g1150(.dina(new_new_n1992__), .dinb(new_new_n1404__), .dout(new_new_n1995__));
  or1   g1151(.dina(new_new_n1995__), .dinb(new_new_n1994__), .dout(new_new_n1996__));
  and1  g1152(.dina(new_new_n2888__), .dinb(new_new_n2890__), .dout(new_new_n1997__));
  or1   g1153(.dina(new_new_n2888__), .dinb(new_new_n2890__), .dout(new_new_n1998__));
  or1   g1154(.dina(new_new_n2892__), .dinb(new_new_n2894__), .dout(new_new_n1999__));
  or1   g1155(.dina(new_new_n2897__), .dinb(new_new_n2894__), .dout(new_new_n2000__));
  and1  g1156(.dina(new_new_n2899__), .dinb(new_new_n2900__), .dout(new_new_n2001__));
  or1   g1157(.dina(new_new_n2901__), .dinb(new_new_n2902__), .dout(new_new_n2002__));
  and1  g1158(.dina(new_new_n2901__), .dinb(new_new_n2902__), .dout(new_new_n2003__));
  or1   g1159(.dina(new_new_n2899__), .dinb(new_new_n2900__), .dout(new_new_n2004__));
  and1  g1160(.dina(new_new_n2004__), .dinb(new_new_n2002__), .dout(new_new_n2005__));
  or1   g1161(.dina(new_new_n2003__), .dinb(new_new_n2001__), .dout(new_new_n2006__));
  and1  g1162(.dina(new_new_n2903__), .dinb(new_new_n2904__), .dout(new_new_n2007__));
  or1   g1163(.dina(new_new_n2905__), .dinb(new_new_n2906__), .dout(new_new_n2008__));
  and1  g1164(.dina(new_new_n2905__), .dinb(new_new_n2906__), .dout(new_new_n2009__));
  or1   g1165(.dina(new_new_n2903__), .dinb(new_new_n2904__), .dout(new_new_n2010__));
  and1  g1166(.dina(new_new_n2010__), .dinb(new_new_n2008__), .dout(new_new_n2011__));
  or1   g1167(.dina(new_new_n2009__), .dinb(new_new_n2007__), .dout(new_new_n2012__));
  and1  g1168(.dina(new_new_n2907__), .dinb(new_new_n2908__), .dout(new_new_n2013__));
  or1   g1169(.dina(new_new_n2909__), .dinb(new_new_n2910__), .dout(new_new_n2014__));
  and1  g1170(.dina(new_new_n2909__), .dinb(new_new_n2910__), .dout(new_new_n2015__));
  or1   g1171(.dina(new_new_n2907__), .dinb(new_new_n2908__), .dout(new_new_n2016__));
  and1  g1172(.dina(new_new_n2016__), .dinb(new_new_n2014__), .dout(new_new_n2017__));
  or1   g1173(.dina(new_new_n2015__), .dinb(new_new_n2013__), .dout(new_new_n2018__));
  and1  g1174(.dina(new_new_n2911__), .dinb(new_new_n2912__), .dout(new_new_n2019__));
  or1   g1175(.dina(new_new_n2897__), .dinb(new_new_n822__), .dout(new_new_n2020__));
  and1  g1176(.dina(new_new_n2019__), .dinb(new_new_n2755__), .dout(new_new_n2021__));
  or1   g1177(.dina(new_new_n2020__), .dinb(new_new_n2758__), .dout(new_new_n2022__));
  and1  g1178(.dina(new_new_n2022__), .dinb(new_new_n2018__), .dout(new_new_n2023__));
  and1  g1179(.dina(new_new_n2021__), .dinb(new_new_n2017__), .dout(new_new_n2024__));
  or1   g1180(.dina(new_new_n2024__), .dinb(new_new_n2023__), .dout(new_new_n2025__));
  and1  g1181(.dina(new_new_n2913__), .dinb(new_new_n2914__), .dout(new_new_n2026__));
  or1   g1182(.dina(new_new_n2915__), .dinb(new_new_n2916__), .dout(new_new_n2027__));
  and1  g1183(.dina(new_new_n2915__), .dinb(new_new_n2916__), .dout(new_new_n2028__));
  or1   g1184(.dina(new_new_n2913__), .dinb(new_new_n2914__), .dout(new_new_n2029__));
  and1  g1185(.dina(new_new_n2029__), .dinb(new_new_n2027__), .dout(new_new_n2030__));
  or1   g1186(.dina(new_new_n2028__), .dinb(new_new_n2026__), .dout(new_new_n2031__));
  and1  g1187(.dina(new_new_n2917__), .dinb(new_new_n2918__), .dout(new_new_n2032__));
  or1   g1188(.dina(new_new_n2919__), .dinb(new_new_n2920__), .dout(new_new_n2033__));
  and1  g1189(.dina(new_new_n2919__), .dinb(new_new_n2920__), .dout(new_new_n2034__));
  or1   g1190(.dina(new_new_n2917__), .dinb(new_new_n2918__), .dout(new_new_n2035__));
  and1  g1191(.dina(new_new_n2035__), .dinb(new_new_n2033__), .dout(new_new_n2036__));
  or1   g1192(.dina(new_new_n2034__), .dinb(new_new_n2032__), .dout(new_new_n2037__));
  and1  g1193(.dina(new_new_n2921__), .dinb(new_new_n2922__), .dout(new_new_n2038__));
  or1   g1194(.dina(new_new_n2923__), .dinb(new_new_n2924__), .dout(new_new_n2039__));
  and1  g1195(.dina(new_new_n2923__), .dinb(new_new_n2924__), .dout(new_new_n2040__));
  or1   g1196(.dina(new_new_n2921__), .dinb(new_new_n2922__), .dout(new_new_n2041__));
  and1  g1197(.dina(new_new_n2041__), .dinb(new_new_n2039__), .dout(new_new_n2042__));
  or1   g1198(.dina(new_new_n2040__), .dinb(new_new_n2038__), .dout(new_new_n2043__));
  and1  g1199(.dina(new_new_n2925__), .dinb(new_new_n2926__), .dout(new_new_n2044__));
  or1   g1200(.dina(new_new_n2927__), .dinb(new_new_n2928__), .dout(new_new_n2045__));
  and1  g1201(.dina(new_new_n2927__), .dinb(new_new_n2928__), .dout(new_new_n2046__));
  or1   g1202(.dina(new_new_n2925__), .dinb(new_new_n2926__), .dout(new_new_n2047__));
  and1  g1203(.dina(new_new_n2047__), .dinb(new_new_n2045__), .dout(new_new_n2048__));
  or1   g1204(.dina(new_new_n2046__), .dinb(new_new_n2044__), .dout(new_new_n2049__));
  and1  g1205(.dina(new_new_n2929__), .dinb(new_new_n2930__), .dout(new_new_n2050__));
  or1   g1206(.dina(new_new_n2931__), .dinb(new_new_n2932__), .dout(new_new_n2051__));
  and1  g1207(.dina(new_new_n2931__), .dinb(new_new_n2932__), .dout(new_new_n2052__));
  or1   g1208(.dina(new_new_n2929__), .dinb(new_new_n2930__), .dout(new_new_n2053__));
  and1  g1209(.dina(new_new_n2053__), .dinb(new_new_n2051__), .dout(new_new_n2054__));
  or1   g1210(.dina(new_new_n2052__), .dinb(new_new_n2050__), .dout(new_new_n2055__));
  and1  g1211(.dina(new_new_n2054__), .dinb(new_new_n2043__), .dout(new_new_n2056__));
  and1  g1212(.dina(new_new_n2055__), .dinb(new_new_n2042__), .dout(new_new_n2057__));
  or1   g1213(.dina(new_new_n2057__), .dinb(new_new_n2056__), .dout(new_new_n2058__));
  and1  g1214(.dina(new_new_n2933__), .dinb(new_new_n2934__), .dout(new_new_n2059__));
  or1   g1215(.dina(new_new_n2935__), .dinb(new_new_n2936__), .dout(new_new_n2060__));
  and1  g1216(.dina(new_new_n2935__), .dinb(new_new_n2936__), .dout(new_new_n2061__));
  or1   g1217(.dina(new_new_n2933__), .dinb(new_new_n2934__), .dout(new_new_n2062__));
  and1  g1218(.dina(new_new_n2062__), .dinb(new_new_n2060__), .dout(new_new_n2063__));
  or1   g1219(.dina(new_new_n2061__), .dinb(new_new_n2059__), .dout(new_new_n2064__));
  and1  g1220(.dina(new_new_n2937__), .dinb(new_new_n2939__), .dout(new_new_n2065__));
  or1   g1221(.dina(new_new_n2940__), .dinb(new_new_n2941__), .dout(new_new_n2066__));
  and1  g1222(.dina(new_new_n2940__), .dinb(new_new_n2941__), .dout(new_new_n2067__));
  or1   g1223(.dina(new_new_n2937__), .dinb(new_new_n2939__), .dout(new_new_n2068__));
  and1  g1224(.dina(new_new_n2068__), .dinb(new_new_n2066__), .dout(new_new_n2069__));
  or1   g1225(.dina(new_new_n2067__), .dinb(new_new_n2065__), .dout(new_new_n2070__));
  and1  g1226(.dina(new_new_n1377__), .dinb(new_new_n1292__), .dout(new_new_n2071__));
  or1   g1227(.dina(new_new_n1378__), .dinb(new_new_n1291__), .dout(new_new_n2072__));
  and1  g1228(.dina(new_new_n1371__), .dinb(new_new_n1298__), .dout(new_new_n2073__));
  or1   g1229(.dina(new_new_n1372__), .dinb(new_new_n1297__), .dout(new_new_n2074__));
  and1  g1230(.dina(new_new_n2074__), .dinb(new_new_n2072__), .dout(new_new_n2075__));
  or1   g1231(.dina(new_new_n2073__), .dinb(new_new_n2071__), .dout(new_new_n2076__));
  and1  g1232(.dina(new_new_n2942__), .dinb(new_new_n2944__), .dout(new_new_n2077__));
  or1   g1233(.dina(new_new_n2946__), .dinb(new_new_n2947__), .dout(new_new_n2078__));
  and1  g1234(.dina(new_new_n2946__), .dinb(new_new_n2947__), .dout(new_new_n2079__));
  or1   g1235(.dina(new_new_n2942__), .dinb(new_new_n2944__), .dout(new_new_n2080__));
  and1  g1236(.dina(new_new_n2080__), .dinb(new_new_n2078__), .dout(new_new_n2081__));
  or1   g1237(.dina(new_new_n2079__), .dinb(new_new_n2077__), .dout(new_new_n2082__));
  and1  g1238(.dina(new_new_n2082__), .dinb(new_new_n2070__), .dout(new_new_n2083__));
  and1  g1239(.dina(new_new_n2081__), .dinb(new_new_n2069__), .dout(new_new_n2084__));
  or1   g1240(.dina(new_new_n2084__), .dinb(new_new_n2083__), .dout(new_new_n2085__));
  and1  g1241(.dina(new_new_n1363__), .dinb(new_new_n1290__), .dout(new_new_n2086__));
  or1   g1242(.dina(new_new_n1364__), .dinb(new_new_n1289__), .dout(new_new_n2087__));
  and1  g1243(.dina(new_new_n1369__), .dinb(new_new_n1274__), .dout(new_new_n2088__));
  or1   g1244(.dina(new_new_n1370__), .dinb(new_new_n1273__), .dout(new_new_n2089__));
  and1  g1245(.dina(new_new_n2089__), .dinb(new_new_n2087__), .dout(new_new_n2090__));
  or1   g1246(.dina(new_new_n2088__), .dinb(new_new_n2086__), .dout(new_new_n2091__));
  and1  g1247(.dina(new_new_n1348__), .dinb(new_new_n1285__), .dout(new_new_n2092__));
  or1   g1248(.dina(new_new_n1347__), .dinb(new_new_n1286__), .dout(new_new_n2093__));
  and1  g1249(.dina(new_new_n1366__), .dinb(new_new_n1259__), .dout(new_new_n2094__));
  or1   g1250(.dina(new_new_n1365__), .dinb(new_new_n1260__), .dout(new_new_n2095__));
  and1  g1251(.dina(new_new_n2095__), .dinb(new_new_n2093__), .dout(new_new_n2096__));
  or1   g1252(.dina(new_new_n2094__), .dinb(new_new_n2092__), .dout(new_new_n2097__));
  and1  g1253(.dina(new_new_n2948__), .dinb(new_new_n2949__), .dout(new_new_n2098__));
  or1   g1254(.dina(new_new_n2950__), .dinb(new_new_n2951__), .dout(new_new_n2099__));
  and1  g1255(.dina(new_new_n2950__), .dinb(new_new_n2951__), .dout(new_new_n2100__));
  or1   g1256(.dina(new_new_n2948__), .dinb(new_new_n2949__), .dout(new_new_n2101__));
  and1  g1257(.dina(new_new_n2101__), .dinb(new_new_n2099__), .dout(new_new_n2102__));
  or1   g1258(.dina(new_new_n2100__), .dinb(new_new_n2098__), .dout(new_new_n2103__));
  and1  g1259(.dina(new_new_n2911__), .dinb(new_new_n2952__), .dout(new_new_n2104__));
  or1   g1260(.dina(new_new_n2898__), .dinb(new_new_n1314__), .dout(new_new_n2105__));
  and1  g1261(.dina(new_new_n2104__), .dinb(new_new_n2755__), .dout(new_new_n2106__));
  or1   g1262(.dina(new_new_n2105__), .dinb(new_new_n2758__), .dout(new_new_n2107__));
  and1  g1263(.dina(new_new_n2953__), .dinb(new_new_n2954__), .dout(new_new_n2108__));
  or1   g1264(.dina(new_new_n2955__), .dinb(new_new_n2891__), .dout(new_new_n2109__));
  and1  g1265(.dina(new_new_n2955__), .dinb(new_new_n2891__), .dout(new_new_n2110__));
  or1   g1266(.dina(new_new_n2953__), .dinb(new_new_n2954__), .dout(new_new_n2111__));
  and1  g1267(.dina(new_new_n2111__), .dinb(new_new_n2109__), .dout(new_new_n2112__));
  or1   g1268(.dina(new_new_n2110__), .dinb(new_new_n2108__), .dout(new_new_n2113__));
  or1   g1269(.dina(new_new_n2112__), .dinb(new_new_n2102__), .dout(new_new_n2114__));
  or1   g1270(.dina(new_new_n2113__), .dinb(new_new_n2103__), .dout(new_new_n2115__));
  and1  g1271(.dina(new_new_n2115__), .dinb(new_new_n2114__), .dout(new_new_n2116__));
  and1  g1272(.dina(new_new_n2957__), .dinb(new_new_n2959__), .dout(new_new_n2117__));
  or1   g1273(.dina(new_new_n2960__), .dinb(new_new_n2961__), .dout(new_new_n2118__));
  and1  g1274(.dina(new_new_n2960__), .dinb(new_new_n2961__), .dout(new_new_n2119__));
  or1   g1275(.dina(new_new_n2957__), .dinb(new_new_n2959__), .dout(new_new_n2120__));
  and1  g1276(.dina(new_new_n2120__), .dinb(new_new_n2118__), .dout(new_new_n2121__));
  or1   g1277(.dina(new_new_n2119__), .dinb(new_new_n2117__), .dout(new_new_n2122__));
  and1  g1278(.dina(new_new_n1374__), .dinb(new_new_n1295__), .dout(new_new_n2123__));
  or1   g1279(.dina(new_new_n1373__), .dinb(new_new_n1296__), .dout(new_new_n2124__));
  and1  g1280(.dina(new_new_n1376__), .dinb(new_new_n1293__), .dout(new_new_n2125__));
  or1   g1281(.dina(new_new_n1375__), .dinb(new_new_n1294__), .dout(new_new_n2126__));
  and1  g1282(.dina(new_new_n2126__), .dinb(new_new_n2124__), .dout(new_new_n2127__));
  or1   g1283(.dina(new_new_n2125__), .dinb(new_new_n2123__), .dout(new_new_n2128__));
  and1  g1284(.dina(new_new_n2962__), .dinb(new_new_n2963__), .dout(new_new_n2129__));
  or1   g1285(.dina(new_new_n2964__), .dinb(new_new_n2966__), .dout(new_new_n2130__));
  and1  g1286(.dina(new_new_n2964__), .dinb(new_new_n2966__), .dout(new_new_n2131__));
  or1   g1287(.dina(new_new_n2962__), .dinb(new_new_n2963__), .dout(new_new_n2132__));
  and1  g1288(.dina(new_new_n2132__), .dinb(new_new_n2130__), .dout(new_new_n2133__));
  or1   g1289(.dina(new_new_n2131__), .dinb(new_new_n2129__), .dout(new_new_n2134__));
  or1   g1290(.dina(new_new_n2133__), .dinb(new_new_n2122__), .dout(new_new_n2135__));
  or1   g1291(.dina(new_new_n2134__), .dinb(new_new_n2121__), .dout(new_new_n2136__));
  and1  g1292(.dina(new_new_n2136__), .dinb(new_new_n2135__), .dout(new_new_n2137__));
  and1  g1293(.dina(new_new_n2827__), .dinb(new_new_n2968__), .dout(new_new_n2138__));
  and1  g1294(.dina(new_new_n2830__), .dinb(new_new_n2970__), .dout(new_new_n2139__));
  or1   g1295(.dina(new_new_n2139__), .dinb(new_new_n2138__), .dout(new_new_n2140__));
  and1  g1296(.dina(new_new_n1336__), .dinb(new_new_n1334__), .dout(new_new_n2141__));
  or1   g1297(.dina(new_new_n1335__), .dinb(new_new_n1333__), .dout(new_new_n2142__));
  and1  g1298(.dina(new_new_n2971__), .dinb(new_new_n2973__), .dout(new_new_n2143__));
  or1   g1299(.dina(new_new_n2974__), .dinb(new_new_n2975__), .dout(new_new_n2144__));
  and1  g1300(.dina(new_new_n2974__), .dinb(new_new_n2975__), .dout(new_new_n2145__));
  or1   g1301(.dina(new_new_n2971__), .dinb(new_new_n2973__), .dout(new_new_n2146__));
  and1  g1302(.dina(new_new_n2146__), .dinb(new_new_n2144__), .dout(new_new_n2147__));
  or1   g1303(.dina(new_new_n2145__), .dinb(new_new_n2143__), .dout(new_new_n2148__));
  and1  g1304(.dina(new_new_n2147__), .dinb(new_new_n1882__), .dout(new_new_n2149__));
  and1  g1305(.dina(new_new_n2148__), .dinb(new_new_n2976__), .dout(new_new_n2150__));
  or1   g1306(.dina(new_new_n2150__), .dinb(new_new_n2149__), .dout(new_new_n2151__));
  or1   g1307(.dina(new_new_n1396__), .dinb(new_new_n2978__), .dout(new_new_n2152__));
  or1   g1308(.dina(new_new_n2981__), .dinb(new_new_n2984__), .dout(new_new_n2153__));
  and1  g1309(.dina(new_new_n2153__), .dinb(new_new_n2152__), .dout(new_new_n2154__));
  and1  g1310(.dina(new_new_n2986__), .dinb(new_new_n2987__), .dout(new_new_n2155__));
  and1  g1311(.dina(new_new_n2990__), .dinb(new_new_n2978__), .dout(new_new_n2156__));
  or1   g1312(.dina(new_new_n2990__), .dinb(new_new_n2977__), .dout(new_new_n2157__));
  or1   g1313(.dina(new_new_n2994__), .dinb(new_new_n2996__), .dout(new_new_n2158__));
  and1  g1314(.dina(new_new_n2994__), .dinb(new_new_n2996__), .dout(new_new_n2159__));
  and1  g1315(.dina(new_new_n838__), .dinb(new_new_n2997__), .dout(new_new_n2160__));
  or1   g1316(.dina(new_new_n2999__), .dinb(new_new_n818__), .dout(new_new_n2161__));
  and1  g1317(.dina(new_new_n2160__), .dinb(new_new_n2986__), .dout(new_new_n2162__));
  or1   g1318(.dina(new_new_n2161__), .dinb(new_new_n3001__), .dout(new_new_n2163__));
  and1  g1319(.dina(new_new_n2163__), .dinb(new_new_n3002__), .dout(new_new_n2164__));
  and1  g1320(.dina(new_new_n2162__), .dinb(new_new_n3003__), .dout(new_new_n2165__));
  or1   g1321(.dina(new_new_n2165__), .dinb(new_new_n2164__), .dout(new_new_n2166__));
  and1  g1322(.dina(new_new_n2830__), .dinb(new_new_n3002__), .dout(new_new_n2167__));
  and1  g1323(.dina(new_new_n2827__), .dinb(new_new_n3003__), .dout(new_new_n2168__));
  or1   g1324(.dina(new_new_n2168__), .dinb(new_new_n2167__), .dout(new_new_n2169__));
  and1  g1325(.dina(new_new_n1306__), .dinb(new_new_n3005__), .dout(new_new_n2170__));
  and1  g1326(.dina(new_new_n1305__), .dinb(new_new_n3007__), .dout(new_new_n2171__));
  or1   g1327(.dina(new_new_n2171__), .dinb(new_new_n2170__), .dout(new_new_n2172__));
  and1  g1328(.dina(new_new_n3008__), .dinb(new_new_n2970__), .dout(new_new_n2173__));
  or1   g1329(.dina(new_new_n3009__), .dinb(new_new_n2968__), .dout(new_new_n2174__));
  and1  g1330(.dina(new_new_n3009__), .dinb(new_new_n2967__), .dout(new_new_n2175__));
  or1   g1331(.dina(new_new_n3008__), .dinb(new_new_n2969__), .dout(new_new_n2176__));
  and1  g1332(.dina(new_new_n2176__), .dinb(new_new_n2174__), .dout(new_new_n2177__));
  or1   g1333(.dina(new_new_n2175__), .dinb(new_new_n2173__), .dout(new_new_n2178__));
  and1  g1334(.dina(new_new_n2178__), .dinb(new_new_n2836__), .dout(new_new_n2179__));
  and1  g1335(.dina(new_new_n2177__), .dinb(new_new_n2838__), .dout(new_new_n2180__));
  or1   g1336(.dina(new_new_n2180__), .dinb(new_new_n2179__), .dout(new_new_n2181__));
  and1  g1337(.dina(new_new_n3005__), .dinb(new_new_n782__), .dout(new_new_n2182__));
  and1  g1338(.dina(new_new_n3007__), .dinb(new_new_n3012__), .dout(new_new_n2183__));
  or1   g1339(.dina(new_new_n2183__), .dinb(new_new_n2182__), .dout(new_new_n2184__));
  buf1  g1340(.din(new_new_n1435__), .dout(G1884));
  buf1  g1341(.din(new_new_n1444__), .dout(G1885));
  buf1  g1342(.din(new_new_n1451__), .dout(G1886));
  buf1  g1343(.din(new_new_n1460__), .dout(G1887));
  buf1  g1344(.din(new_new_n1471__), .dout(G1888));
  buf1  g1345(.din(new_new_n1482__), .dout(G1889));
  buf1  g1346(.din(new_new_n1491__), .dout(G1890));
  buf1  g1347(.din(new_new_n1502__), .dout(G1891));
  buf1  g1348(.din(new_new_n1513__), .dout(G1892));
  buf1  g1349(.din(new_new_n1522__), .dout(G1893));
  buf1  g1350(.din(new_new_n1531__), .dout(G1894));
  buf1  g1351(.din(new_new_n1540__), .dout(G1895));
  buf1  g1352(.din(new_new_n1551__), .dout(G1896));
  buf1  g1353(.din(new_new_n1558__), .dout(G1897));
  buf1  g1354(.din(new_new_n1567__), .dout(G1898));
  buf1  g1355(.din(new_new_n1576__), .dout(G1899));
  buf1  g1356(.din(new_new_n1646__), .dout(G1900));
  buf1  g1357(.din(new_new_n1669__), .dout(G1901));
  buf1  g1358(.din(new_new_n1691__), .dout(G1902));
  buf1  g1359(.din(new_new_n1699__), .dout(G1903));
  buf1  g1360(.din(new_new_n1707__), .dout(G1904));
  buf1  g1361(.din(new_new_n1717__), .dout(G1905));
  buf1  g1362(.din(new_new_n1752__), .dout(G1906));
  buf1  g1363(.din(new_new_n1787__), .dout(G1907));
  buf1  g1364(.din(new_new_n1813__), .dout(G1908));
  buf1  g1365(.din(new_new_n919__), .dout(n4857));
  buf1  g1366(.din(new_new_n903__), .dout(n4860));
  buf1  g1367(.din(new_new_n907__), .dout(n4863));
  buf1  g1368(.din(new_new_n715__), .dout(n4866));
  buf1  g1369(.din(new_new_n967__), .dout(n4869));
  buf1  g1370(.din(new_new_n933__), .dout(n4872));
  buf1  g1371(.din(new_new_n909__), .dout(n4875));
  buf1  g1372(.din(new_new_n915__), .dout(n4878));
  buf1  g1373(.din(new_new_n723__), .dout(n4881));
  buf1  g1374(.din(new_new_n969__), .dout(n4884));
  buf1  g1375(.din(new_new_n725__), .dout(n4887));
  buf1  g1376(.din(new_new_n971__), .dout(n4890));
  buf1  g1377(.din(new_new_n921__), .dout(n4893));
  buf1  g1378(.din(new_new_n935__), .dout(n4896));
  buf1  g1379(.din(new_new_n911__), .dout(n4899));
  buf1  g1380(.din(new_new_n917__), .dout(n4902));
  buf1  g1381(.din(new_new_n963__), .dout(n4905));
  buf1  g1382(.din(new_new_n905__), .dout(n4908));
  buf1  g1383(.din(new_new_n913__), .dout(n4911));
  buf1  g1384(.din(new_new_n741__), .dout(n4914));
  buf1  g1385(.din(new_new_n2733__), .dout(n4917));
  buf1  g1386(.din(new_new_n743__), .dout(n4920));
  buf1  g1387(.din(new_new_n745__), .dout(n4923));
  buf1  g1388(.din(new_new_n819__), .dout(n4926));
  buf1  g1389(.din(new_new_n2737__), .dout(n4929));
  buf1  g1390(.din(new_new_n747__), .dout(n4932));
  buf1  g1391(.din(new_new_n749__), .dout(n4935));
  buf1  g1392(.din(new_new_n1007__), .dout(n4938));
  buf1  g1393(.din(new_new_n751__), .dout(n4941));
  buf1  g1394(.din(new_new_n1031__), .dout(n4944));
  buf1  g1395(.din(new_new_n753__), .dout(n4947));
  buf1  g1396(.din(new_new_n755__), .dout(n4950));
  buf1  g1397(.din(new_new_n757__), .dout(n4953));
  buf1  g1398(.din(new_new_n839__), .dout(n4956));
  buf1  g1399(.din(new_new_n2763__), .dout(n4959));
  buf1  g1400(.din(new_new_n759__), .dout(n4962));
  buf1  g1401(.din(new_new_n845__), .dout(n4965));
  buf1  g1402(.din(new_new_n2782__), .dout(n4968));
  buf1  g1403(.din(new_new_n761__), .dout(n4971));
  buf1  g1404(.din(new_new_n851__), .dout(n4974));
  buf1  g1405(.din(new_new_n2787__), .dout(n4977));
  buf1  g1406(.din(new_new_n763__), .dout(n4980));
  buf1  g1407(.din(new_new_n857__), .dout(n4983));
  buf1  g1408(.din(new_new_n2784__), .dout(n4986));
  buf1  g1409(.din(new_new_n765__), .dout(n4989));
  buf1  g1410(.din(new_new_n863__), .dout(n4992));
  buf1  g1411(.din(new_new_n865__), .dout(n4995));
  buf1  g1412(.din(new_new_n3015__), .dout(n4998));
  buf1  g1413(.din(new_new_n767__), .dout(n5001));
  buf1  g1414(.din(new_new_n871__), .dout(n5004));
  buf1  g1415(.din(new_new_n873__), .dout(n5007));
  buf1  g1416(.din(new_new_n3016__), .dout(n5010));
  buf1  g1417(.din(new_new_n769__), .dout(n5013));
  buf1  g1418(.din(new_new_n879__), .dout(n5016));
  buf1  g1419(.din(new_new_n1177__), .dout(n5019));
  buf1  g1420(.din(new_new_n771__), .dout(n5022));
  buf1  g1421(.din(new_new_n885__), .dout(n5025));
  buf1  g1422(.din(new_new_n887__), .dout(n5028));
  buf1  g1423(.din(new_new_n3017__), .dout(n5031));
  buf1  g1424(.din(new_new_n773__), .dout(n5034));
  buf1  g1425(.din(new_new_n3019__), .dout(n5037));
  buf1  g1426(.din(new_new_n937__), .dout(n5040));
  buf1  g1427(.din(new_new_n1033__), .dout(n5043));
  buf1  g1428(.din(new_new_n1109__), .dout(n5046));
  buf1  g1429(.din(new_new_n1037__), .dout(n5049));
  buf1  g1430(.din(new_new_n1039__), .dout(n5052));
  buf1  g1431(.din(new_new_n1043__), .dout(n5055));
  buf1  g1432(.din(new_new_n1045__), .dout(n5058));
  buf1  g1433(.din(new_new_n1047__), .dout(n5061));
  buf1  g1434(.din(new_new_n1049__), .dout(n5064));
  buf1  g1435(.din(new_new_n1059__), .dout(n5067));
  buf1  g1436(.din(new_new_n1061__), .dout(n5070));
  buf1  g1437(.din(new_new_n1063__), .dout(n5073));
  buf1  g1438(.din(new_new_n1065__), .dout(n5076));
  buf1  g1439(.din(new_new_n2735__), .dout(n5079));
  buf1  g1440(.din(new_new_n2731__), .dout(n5082));
  buf1  g1441(.din(new_new_n2739__), .dout(n5085));
  buf1  g1442(.din(new_new_n2750__), .dout(n5088));
  buf1  g1443(.din(new_new_n2751__), .dout(n5091));
  buf1  g1444(.din(new_new_n1071__), .dout(n5094));
  buf1  g1445(.din(new_new_n1073__), .dout(n5097));
  buf1  g1446(.din(new_new_n2958__), .dout(n5100));
  buf1  g1447(.din(new_new_n2761__), .dout(n5103));
  buf1  g1448(.din(new_new_n2779__), .dout(n5106));
  buf1  g1449(.din(new_new_n2762__), .dout(n5109));
  buf1  g1450(.din(new_new_n2781__), .dout(n5112));
  buf1  g1451(.din(new_new_n2786__), .dout(n5115));
  buf1  g1452(.din(new_new_n2783__), .dout(n5118));
  buf1  g1453(.din(new_new_n2785__), .dout(n5121));
  buf1  g1454(.din(new_new_n2788__), .dout(n5124));
  buf1  g1455(.din(new_new_n2778__), .dout(n5127));
  buf1  g1456(.din(new_new_n2780__), .dout(n5130));
  buf1  g1457(.din(new_new_n2760__), .dout(n5133));
  buf1  g1458(.din(new_new_n2764__), .dout(n5136));
  buf1  g1459(.din(new_new_n1113__), .dout(n5139));
  buf1  g1460(.din(new_new_n1115__), .dout(n5142));
  buf1  g1461(.din(new_new_n1117__), .dout(n5145));
  buf1  g1462(.din(new_new_n1119__), .dout(n5148));
  buf1  g1463(.din(new_new_n1121__), .dout(n5151));
  buf1  g1464(.din(new_new_n1123__), .dout(n5154));
  buf1  g1465(.din(new_new_n2892__), .dout(n5157));
  buf1  g1466(.din(new_new_n1171__), .dout(n5160));
  buf1  g1467(.din(new_new_n1173__), .dout(n5163));
  buf1  g1468(.din(new_new_n1175__), .dout(n5166));
  buf1  g1469(.din(new_new_n1179__), .dout(n5169));
  buf1  g1470(.din(new_new_n1185__), .dout(n5172));
  buf1  g1471(.din(new_new_n1187__), .dout(n5175));
  buf1  g1472(.din(new_new_n1189__), .dout(n5178));
  buf1  g1473(.din(new_new_n1191__), .dout(n5181));
  buf1  g1474(.din(new_new_n1193__), .dout(n5184));
  buf1  g1475(.din(new_new_n2767__), .dout(n5187));
  buf1  g1476(.din(new_new_n2770__), .dout(n5190));
  buf1  g1477(.din(new_new_n1229__), .dout(n5193));
  buf1  g1478(.din(new_new_n1231__), .dout(n5196));
  buf1  g1479(.din(new_new_n2945__), .dout(n5199));
  buf1  g1480(.din(new_new_n1235__), .dout(n5202));
  buf1  g1481(.din(new_new_n1267__), .dout(n5205));
  buf1  g1482(.din(new_new_n1257__), .dout(n5208));
  buf1  g1483(.din(new_new_n2752__), .dout(n5211));
  not1  g1484(.din(new_new_n2776__), .dout(n5214));
  buf1  g1485(.din(n4998), .dout(n5217));
  buf1  g1486(.din(n5010), .dout(n5220));
  buf1  g1487(.din(n5031), .dout(n5223));
  buf1  g1488(.din(n5037), .dout(n5226));
  buf1  g1489(.din(new_new_n3018__), .dout(n5229));
  buf1  g1490(.din(new_new_n2972__), .dout(n5232));
  buf1  g1491(.din(new_new_n2792__), .dout(n5235));
  buf1  g1492(.din(new_new_n2952__), .dout(n5238));
  buf1  g1493(.din(new_new_n2759__), .dout(n5241));
  buf1  g1494(.din(new_new_n2956__), .dout(n5244));
  buf1  g1495(.din(n5199), .dout(n5247));
  buf1  g1496(.din(new_new_n1195__), .dout(n5250));
  buf1  g1497(.din(new_new_n1197__), .dout(n5253));
  buf1  g1498(.din(new_new_n2965__), .dout(n5256));
  buf1  g1499(.din(new_new_n1237__), .dout(n5259));
  buf1  g1500(.din(new_new_n1239__), .dout(n5262));
  buf1  g1501(.din(new_new_n1241__), .dout(n5265));
  buf1  g1502(.din(new_new_n1243__), .dout(n5268));
  buf1  g1503(.din(new_new_n1245__), .dout(n5271));
  buf1  g1504(.din(new_new_n2938__), .dout(n5274));
  buf1  g1505(.din(new_new_n2765__), .dout(n5277));
  not1  g1506(.din(new_new_n2768__), .dout(n5280));
  buf1  g1507(.din(new_new_n1299__), .dout(n5283));
  buf1  g1508(.din(new_new_n1301__), .dout(n5286));
  buf1  g1509(.din(new_new_n1359__), .dout(n5289));
  buf1  g1510(.din(new_new_n1361__), .dout(n5292));
  buf1  g1511(.din(new_new_n1381__), .dout(n5295));
  buf1  g1512(.din(new_new_n1387__), .dout(n5298));
  buf1  g1513(.din(new_new_n2837__), .dout(n5301));
  buf1  g1514(.din(new_new_n2886__), .dout(n5304));
  buf1  g1515(.din(new_new_n2839__), .dout(n5307));
  buf1  g1516(.din(new_new_n2797__), .dout(n5310));
  buf1  g1517(.din(new_new_n2816__), .dout(n5313));
  not1  g1518(.din(new_new_n2818__), .dout(n5316));
  not1  g1519(.din(new_new_n2812__), .dout(n5319));
  not1  g1520(.din(new_new_n2815__), .dout(n5322));
  buf1  g1521(.din(n5322), .dout(n5325));
  not1  g1522(.din(new_new_n2796__), .dout(n5328));
  buf1  g1523(.din(n5328), .dout(n5331));
  buf1  g1524(.din(new_new_n2801__), .dout(n5334));
  buf1  g1525(.din(new_new_n2803__), .dout(n5337));
  buf1  g1526(.din(n5337), .dout(n5340));
  buf1  g1527(.din(new_new_n2802__), .dout(n5343));
  not1  g1528(.din(new_new_n2807__), .dout(n5346));
  not1  g1529(.din(new_new_n2809__), .dout(n5349));
  buf1  g1530(.din(n5349), .dout(n5352));
  not1  g1531(.din(new_new_n2808__), .dout(n5355));
  buf1  g1532(.din(new_new_n2976__), .dout(n5358));
  buf1  g1533(.din(new_new_n2912__), .dout(n5361));
  buf1  g1534(.din(new_new_n2981__), .dout(n5364));
  buf1  g1535(.din(new_new_n2887__), .dout(n5367));
  buf1  g1536(.din(new_new_n3012__), .dout(n5370));
  buf1  g1537(.din(new_new_n3006__), .dout(n5373));
  buf1  g1538(.din(new_new_n2984__), .dout(n5376));
  buf1  g1539(.din(new_new_n2980__), .dout(n5379));
  buf1  g1540(.din(new_new_n3020__), .dout(n5382));
  buf1  g1541(.din(new_new_n3021__), .dout(n5385));
  buf1  g1542(.din(new_new_n3022__), .dout(n5388));
  buf1  g1543(.din(new_new_n3023__), .dout(n5391));
  buf1  g1544(.din(new_new_n3024__), .dout(n5394));
  buf1  g1545(.din(new_new_n3025__), .dout(n5397));
  buf1  g1546(.din(new_new_n2863__), .dout(n5400));
  buf1  g1547(.din(n5400), .dout(n5403));
  buf1  g1548(.din(new_new_n2864__), .dout(n5406));
  buf1  g1549(.din(n5406), .dout(n5409));
  buf1  g1550(.din(new_new_n2874__), .dout(n5412));
  buf1  g1551(.din(n5412), .dout(n5415));
  buf1  g1552(.din(new_new_n2875__), .dout(n5418));
  buf1  g1553(.din(n5418), .dout(n5421));
  buf1  g1554(.din(new_new_n2857__), .dout(n5424));
  buf1  g1555(.din(new_new_n2867__), .dout(n5427));
  buf1  g1556(.din(new_new_n2866__), .dout(n5430));
  buf1  g1557(.din(new_new_n2868__), .dout(n5433));
  buf1  g1558(.din(n5433), .dout(n5436));
  buf1  g1559(.din(new_new_n2855__), .dout(n5439));
  buf1  g1560(.din(new_new_n2856__), .dout(n5442));
  buf1  g1561(.din(n5442), .dout(n5445));
  buf1  g1562(.din(new_new_n2999__), .dout(n5448));
  buf1  g1563(.din(new_new_n3001__), .dout(n5451));
  buf1  g1564(.din(new_new_n3013__), .dout(n5454));
  buf1  g1565(.din(new_new_n2985__), .dout(n5457));
  buf1  g1566(.din(new_new_n2895__), .dout(n5460));
  buf1  g1567(.din(new_new_n2997__), .dout(n5463));
  buf1  g1568(.din(new_new_n2998__), .dout(n5466));
  buf1  g1569(.din(new_new_n3000__), .dout(n5469));
  buf1  g1570(.din(n5457), .dout(n5472));
  buf1  g1571(.din(new_new_n2991__), .dout(n5475));
  buf1  g1572(.din(new_new_n2995__), .dout(n5478));
  buf1  g1573(.din(new_new_n2993__), .dout(n5481));
  buf1  g1574(.din(new_new_n3027__), .dout(n5484));
  buf1  g1575(.din(new_new_n3031__), .dout(n5487));
  buf1  g1576(.din(new_new_n3035__), .dout(n5490));
  buf1  g1577(.din(new_new_n2898__), .dout(n5493));
  not1  g1578(.din(new_new_n1945__), .dout(n5496));
  not1  g1579(.din(new_new_n1949__), .dout(n5499));
  buf1  g1580(.din(new_new_n1950__), .dout(n5502));
  not1  g1581(.din(new_new_n1951__), .dout(n5505));
  buf1  g1582(.din(new_new_n1966__), .dout(n5508));
  buf1  g1583(.din(new_new_n1967__), .dout(n5511));
  buf1  g1584(.din(n5382), .dout(n5514));
  buf1  g1585(.din(n5385), .dout(n5517));
  buf1  g1586(.din(n5388), .dout(n5520));
  buf1  g1587(.din(n5391), .dout(n5523));
  buf1  g1588(.din(n5394), .dout(n5526));
  buf1  g1589(.din(n5397), .dout(n5529));
  buf1  g1590(.din(new_new_n1974__), .dout(n5532));
  buf1  g1591(.din(new_new_n1978__), .dout(n5535));
  buf1  g1592(.din(new_new_n3038__), .dout(n5538));
  buf1  g1593(.din(n5475), .dout(n5541));
  buf1  g1594(.din(new_new_n3040__), .dout(n5544));
  buf1  g1595(.din(n5484), .dout(n5547));
  buf1  g1596(.din(new_new_n3042__), .dout(n5550));
  buf1  g1597(.din(new_new_n3045__), .dout(n5553));
  buf1  g1598(.din(new_new_n3048__), .dout(n5556));
  buf1  g1599(.din(new_new_n3052__), .dout(n5559));
  buf1  g1600(.din(n5487), .dout(n5562));
  buf1  g1601(.din(n5490), .dout(n5565));
  buf1  g1602(.din(new_new_n841__), .dout(n5568));
  buf1  g1603(.din(new_new_n847__), .dout(n5571));
  buf1  g1604(.din(new_new_n853__), .dout(n5574));
  buf1  g1605(.din(new_new_n859__), .dout(n5577));
  buf1  g1606(.din(new_new_n2982__), .dout(n5580));
  buf1  g1607(.din(n5454), .dout(n5583));
  buf1  g1608(.din(n5460), .dout(n5586));
  buf1  g1609(.din(new_new_n1997__), .dout(n5589));
  buf1  g1610(.din(new_new_n1998__), .dout(n5592));
  buf1  g1611(.din(new_new_n2987__), .dout(n5595));
  buf1  g1612(.din(new_new_n1999__), .dout(n5598));
  buf1  g1613(.din(new_new_n2000__), .dout(n5601));
  buf1  g1614(.din(new_new_n3055__), .dout(n5604));
  buf1  g1615(.din(new_new_n2025__), .dout(n5607));
  buf1  g1616(.din(new_new_n2058__), .dout(n5610));
  buf1  g1617(.din(new_new_n2085__), .dout(n5613));
  buf1  g1618(.din(new_new_n2116__), .dout(n5616));
  buf1  g1619(.din(new_new_n2137__), .dout(n5619));
  buf1  g1620(.din(new_new_n3056__), .dout(n5622));
  buf1  g1621(.din(new_new_n2151__), .dout(n5625));
  buf1  g1622(.din(new_new_n3058__), .dout(n5628));
  buf1  g1623(.din(n5538), .dout(n5631));
  buf1  g1624(.din(new_new_n2992__), .dout(n5634));
  buf1  g1625(.din(n5544), .dout(n5637));
  buf1  g1626(.din(new_new_n3028__), .dout(n5640));
  buf1  g1627(.din(new_new_n3060__), .dout(n5643));
  buf1  g1628(.din(new_new_n3062__), .dout(n5646));
  buf1  g1629(.din(n5550), .dout(n5649));
  buf1  g1630(.din(n5553), .dout(n5652));
  buf1  g1631(.din(n5556), .dout(n5655));
  buf1  g1632(.din(n5559), .dout(n5658));
  buf1  g1633(.din(new_new_n3030__), .dout(n5661));
  buf1  g1634(.din(new_new_n825__), .dout(n5664));
  buf1  g1635(.din(new_new_n831__), .dout(n5667));
  buf1  g1636(.din(new_new_n2877__), .dout(n5670));
  buf1  g1637(.din(new_new_n1307__), .dout(n5673));
  buf1  g1638(.din(n5301), .dout(n5676));
  buf1  g1639(.din(n5367), .dout(n5679));
  buf1  g1640(.din(new_new_n3014__), .dout(n5682));
  buf1  g1641(.din(n5373), .dout(n5685));
  buf1  g1642(.din(new_new_n2155__), .dout(n5688));
  buf1  g1643(.din(n5604), .dout(n5691));
  buf1  g1644(.din(new_new_n2156__), .dout(n5694));
  not1  g1645(.din(new_new_n2157__), .dout(n5697));
  buf1  g1646(.din(new_new_n2158__), .dout(n5700));
  buf1  g1647(.din(new_new_n2159__), .dout(n5703));
  buf1  g1648(.din(new_new_n813__), .dout(n5706));
  buf1  g1649(.din(new_new_n835__), .dout(n5709));
  buf1  g1650(.din(n5580), .dout(n5712));
  buf1  g1651(.din(n5682), .dout(n5715));
  buf1  g1652(.din(new_new_n2166__), .dout(n5718));
  buf1  g1653(.din(new_new_n2169__), .dout(n5721));
  buf1  g1654(.din(new_new_n2172__), .dout(n5724));
  buf1  g1655(.din(new_new_n2181__), .dout(n5727));
  buf1  g1656(.din(n5628), .dout(n5730));
  buf1  g1657(.din(new_new_n3063__), .dout(n5733));
  buf1  g1658(.din(new_new_n3064__), .dout(n5736));
  buf1  g1659(.din(new_new_n3054__), .dout(n5739));
  buf1  g1660(.din(n5622), .dout(n5742));
  buf1  g1661(.din(new_new_n2184__), .dout(n5745));
  buf1  g1662(.din(new_new_n3057__), .dout(n5748));
  buf1  g1663(.din(new_new_n3037__), .dout(n5751));
  buf1  g1664(.din(n5634), .dout(n5754));
  buf1  g1665(.din(new_new_n3039__), .dout(n5757));
  buf1  g1666(.din(n5640), .dout(n5760));
  buf1  g1667(.din(n5643), .dout(n5763));
  buf1  g1668(.din(n5646), .dout(n5766));
  buf1  g1669(.din(new_new_n3043__), .dout(n5769));
  buf1  g1670(.din(new_new_n3046__), .dout(n5772));
  buf1  g1671(.din(new_new_n3049__), .dout(n5775));
  buf1  g1672(.din(new_new_n3051__), .dout(n5778));
  buf1  g1673(.din(new_new_n3032__), .dout(n5781));
  buf1  g1674(.din(new_new_n3034__), .dout(n5784));
  buf1  g1675(.din(new_new_n735__), .dout(n5787));
  buf1  g1676(.din(new_new_n3053__), .dout(n5790));
  buf1  g1677(.din(new_new_n3036__), .dout(n5793));
  buf1  g1678(.din(new_new_n717__), .dout(n5796));
  buf1  g1679(.din(new_new_n729__), .dout(n5799));
  buf1  g1680(.din(n5733), .dout(n5802));
  buf1  g1681(.din(n5736), .dout(n5805));
  buf1  g1682(.din(new_new_n3059__), .dout(n5808));
  buf1  g1683(.din(new_new_n3061__), .dout(n5811));
  buf1  g1684(.din(n5769), .dout(n5814));
  buf1  g1685(.din(n5772), .dout(n5817));
  buf1  g1686(.din(n5775), .dout(n5820));
  buf1  g1687(.din(n5790), .dout(n5823));
  buf1  g1688(.din(n5781), .dout(n5826));
  buf1  g1689(.din(n5793), .dout(n5829));
  buf1  g1690(.din(new_new_n1090__), .dout(new_new_n2535__));
  buf1  g1691(.din(new_new_n1086__), .dout(new_new_n2536__));
  buf1  g1692(.din(new_new_n1089__), .dout(new_new_n2537__));
  buf1  g1693(.din(new_new_n1085__), .dout(new_new_n2538__));
  buf1  g1694(.din(new_new_n1425__), .dout(new_new_n2539__));
  buf1  g1695(.din(new_new_n2539__), .dout(new_new_n2540__));
  buf1  g1696(.din(new_new_n1095__), .dout(new_new_n2541__));
  buf1  g1697(.din(new_new_n2541__), .dout(new_new_n2542__));
  buf1  g1698(.din(new_new_n2542__), .dout(new_new_n2543__));
  buf1  g1699(.din(new_new_n2542__), .dout(new_new_n2544__));
  buf1  g1700(.din(new_new_n2541__), .dout(new_new_n2545__));
  buf1  g1701(.din(new_new_n1426__), .dout(new_new_n2546__));
  buf1  g1702(.din(new_new_n2546__), .dout(new_new_n2547__));
  buf1  g1703(.din(new_new_n1096__), .dout(new_new_n2548__));
  buf1  g1704(.din(new_new_n2548__), .dout(new_new_n2549__));
  buf1  g1705(.din(new_new_n2549__), .dout(new_new_n2550__));
  buf1  g1706(.din(new_new_n2548__), .dout(new_new_n2551__));
  buf1  g1707(.din(new_new_n1102__), .dout(new_new_n2552__));
  buf1  g1708(.din(new_new_n2552__), .dout(new_new_n2553__));
  buf1  g1709(.din(new_new_n2553__), .dout(new_new_n2554__));
  buf1  g1710(.din(new_new_n2554__), .dout(new_new_n2555__));
  buf1  g1711(.din(new_new_n2554__), .dout(new_new_n2556__));
  buf1  g1712(.din(new_new_n2553__), .dout(new_new_n2557__));
  buf1  g1713(.din(new_new_n2552__), .dout(new_new_n2558__));
  buf1  g1714(.din(new_new_n2558__), .dout(new_new_n2559__));
  buf1  g1715(.din(new_new_n2558__), .dout(new_new_n2560__));
  buf1  g1716(.din(new_new_n1101__), .dout(new_new_n2561__));
  buf1  g1717(.din(new_new_n2561__), .dout(new_new_n2562__));
  buf1  g1718(.din(new_new_n2561__), .dout(new_new_n2563__));
  buf1  g1719(.din(new_new_n1082__), .dout(new_new_n2564__));
  buf1  g1720(.din(new_new_n2564__), .dout(new_new_n2565__));
  buf1  g1721(.din(new_new_n2565__), .dout(new_new_n2566__));
  buf1  g1722(.din(new_new_n2565__), .dout(new_new_n2567__));
  buf1  g1723(.din(new_new_n2564__), .dout(new_new_n2568__));
  buf1  g1724(.din(new_new_n2568__), .dout(new_new_n2569__));
  buf1  g1725(.din(new_new_n2568__), .dout(new_new_n2570__));
  buf1  g1726(.din(new_new_n1081__), .dout(new_new_n2571__));
  buf1  g1727(.din(new_new_n2571__), .dout(new_new_n2572__));
  buf1  g1728(.din(new_new_n2572__), .dout(new_new_n2573__));
  buf1  g1729(.din(new_new_n2572__), .dout(new_new_n2574__));
  buf1  g1730(.din(new_new_n2571__), .dout(new_new_n2575__));
  buf1  g1731(.din(new_new_n2575__), .dout(new_new_n2576__));
  buf1  g1732(.din(new_new_n2575__), .dout(new_new_n2577__));
  buf1  g1733(.din(new_new_n1093__), .dout(new_new_n2578__));
  buf1  g1734(.din(new_new_n2578__), .dout(new_new_n2579__));
  buf1  g1735(.din(new_new_n2579__), .dout(new_new_n2580__));
  buf1  g1736(.din(new_new_n2579__), .dout(new_new_n2581__));
  buf1  g1737(.din(new_new_n2578__), .dout(new_new_n2582__));
  buf1  g1738(.din(new_new_n1094__), .dout(new_new_n2583__));
  buf1  g1739(.din(new_new_n1436__), .dout(new_new_n2584__));
  buf1  g1740(.din(new_new_n1106__), .dout(new_new_n2585__));
  buf1  g1741(.din(new_new_n2585__), .dout(new_new_n2586__));
  buf1  g1742(.din(new_new_n2586__), .dout(new_new_n2587__));
  buf1  g1743(.din(new_new_n2586__), .dout(new_new_n2588__));
  buf1  g1744(.din(new_new_n2585__), .dout(new_new_n2589__));
  buf1  g1745(.din(new_new_n2589__), .dout(new_new_n2590__));
  buf1  g1746(.din(new_new_n1437__), .dout(new_new_n2591__));
  buf1  g1747(.din(new_new_n1105__), .dout(new_new_n2592__));
  buf1  g1748(.din(new_new_n2592__), .dout(new_new_n2593__));
  buf1  g1749(.din(new_new_n2593__), .dout(new_new_n2594__));
  buf1  g1750(.din(new_new_n2593__), .dout(new_new_n2595__));
  buf1  g1751(.din(new_new_n2592__), .dout(new_new_n2596__));
  buf1  g1752(.din(new_new_n1104__), .dout(new_new_n2597__));
  buf1  g1753(.din(new_new_n2597__), .dout(new_new_n2598__));
  buf1  g1754(.din(new_new_n2598__), .dout(new_new_n2599__));
  buf1  g1755(.din(new_new_n2597__), .dout(new_new_n2600__));
  buf1  g1756(.din(new_new_n1103__), .dout(new_new_n2601__));
  buf1  g1757(.din(new_new_n2601__), .dout(new_new_n2602__));
  buf1  g1758(.din(new_new_n2601__), .dout(new_new_n2603__));
  buf1  g1759(.din(new_new_n1097__), .dout(new_new_n2604__));
  buf1  g1760(.din(new_new_n2604__), .dout(new_new_n2605__));
  buf1  g1761(.din(new_new_n2604__), .dout(new_new_n2606__));
  buf1  g1762(.din(new_new_n1098__), .dout(new_new_n2607__));
  buf1  g1763(.din(new_new_n2607__), .dout(new_new_n2608__));
  buf1  g1764(.din(new_new_n1088__), .dout(new_new_n2609__));
  buf1  g1765(.din(new_new_n2609__), .dout(new_new_n2610__));
  buf1  g1766(.din(new_new_n1087__), .dout(new_new_n2611__));
  buf1  g1767(.din(new_new_n2611__), .dout(new_new_n2612__));
  buf1  g1768(.din(new_new_n1099__), .dout(new_new_n2613__));
  buf1  g1769(.din(new_new_n2613__), .dout(new_new_n2614__));
  buf1  g1770(.din(new_new_n2613__), .dout(new_new_n2615__));
  buf1  g1771(.din(new_new_n1100__), .dout(new_new_n2616__));
  buf1  g1772(.din(new_new_n2616__), .dout(new_new_n2617__));
  buf1  g1773(.din(new_new_n2616__), .dout(new_new_n2618__));
  buf1  g1774(.din(new_new_n1084__), .dout(new_new_n2619__));
  buf1  g1775(.din(new_new_n2619__), .dout(new_new_n2620__));
  buf1  g1776(.din(new_new_n2620__), .dout(new_new_n2621__));
  buf1  g1777(.din(new_new_n2620__), .dout(new_new_n2622__));
  buf1  g1778(.din(new_new_n2619__), .dout(new_new_n2623__));
  buf1  g1779(.din(new_new_n2623__), .dout(new_new_n2624__));
  buf1  g1780(.din(new_new_n2623__), .dout(new_new_n2625__));
  buf1  g1781(.din(new_new_n1083__), .dout(new_new_n2626__));
  buf1  g1782(.din(new_new_n2626__), .dout(new_new_n2627__));
  buf1  g1783(.din(new_new_n2627__), .dout(new_new_n2628__));
  buf1  g1784(.din(new_new_n2627__), .dout(new_new_n2629__));
  buf1  g1785(.din(new_new_n2626__), .dout(new_new_n2630__));
  buf1  g1786(.din(new_new_n2630__), .dout(new_new_n2631__));
  buf1  g1787(.din(new_new_n2630__), .dout(new_new_n2632__));
  buf1  g1788(.din(new_new_n1092__), .dout(new_new_n2633__));
  buf1  g1789(.din(new_new_n1091__), .dout(new_new_n2634__));
  buf1  g1790(.din(new_new_n1472__), .dout(new_new_n2635__));
  buf1  g1791(.din(new_new_n1473__), .dout(new_new_n2636__));
  buf1  g1792(.din(new_new_n1108__), .dout(new_new_n2637__));
  buf1  g1793(.din(new_new_n1107__), .dout(new_new_n2638__));
  buf1  g1794(.din(new_new_n1079__), .dout(new_new_n2639__));
  buf1  g1795(.din(new_new_n2639__), .dout(new_new_n2640__));
  buf1  g1796(.din(new_new_n2639__), .dout(new_new_n2641__));
  buf1  g1797(.din(new_new_n1080__), .dout(new_new_n2642__));
  buf1  g1798(.din(new_new_n1503__), .dout(new_new_n2643__));
  buf1  g1799(.din(new_new_n2643__), .dout(new_new_n2644__));
  buf1  g1800(.din(new_new_n2643__), .dout(new_new_n2645__));
  buf1  g1801(.din(new_new_n1504__), .dout(new_new_n2646__));
  buf1  g1802(.din(new_new_n2646__), .dout(new_new_n2647__));
  buf1  g1803(.din(new_new_n2646__), .dout(new_new_n2648__));
  buf1  g1804(.din(new_new_n1523__), .dout(new_new_n2649__));
  buf1  g1805(.din(new_new_n1077__), .dout(new_new_n2650__));
  buf1  g1806(.din(new_new_n2650__), .dout(new_new_n2651__));
  buf1  g1807(.din(new_new_n1541__), .dout(new_new_n2652__));
  buf1  g1808(.din(new_new_n2652__), .dout(new_new_n2653__));
  buf1  g1809(.din(new_new_n2652__), .dout(new_new_n2654__));
  buf1  g1810(.din(new_new_n1542__), .dout(new_new_n2655__));
  buf1  g1811(.din(new_new_n2655__), .dout(new_new_n2656__));
  buf1  g1812(.din(new_new_n1543__), .dout(new_new_n2657__));
  buf1  g1813(.din(new_new_n1544__), .dout(new_new_n2658__));
  buf1  g1814(.din(new_new_n1602__), .dout(new_new_n2659__));
  buf1  g1815(.din(new_new_n891__), .dout(new_new_n2660__));
  buf1  g1816(.din(new_new_n2660__), .dout(new_new_n2661__));
  buf1  g1817(.din(new_new_n1606__), .dout(new_new_n2662__));
  buf1  g1818(.din(new_new_n2662__), .dout(new_new_n2663__));
  buf1  g1819(.din(new_new_n2663__), .dout(new_new_n2664__));
  buf1  g1820(.din(new_new_n2663__), .dout(new_new_n2665__));
  buf1  g1821(.din(new_new_n2662__), .dout(new_new_n2666__));
  buf1  g1822(.din(new_new_n2666__), .dout(new_new_n2667__));
  buf1  g1823(.din(new_new_n2666__), .dout(new_new_n2668__));
  buf1  g1824(.din(new_new_n1612__), .dout(new_new_n2669__));
  buf1  g1825(.din(new_new_n2669__), .dout(new_new_n2670__));
  buf1  g1826(.din(new_new_n1616__), .dout(new_new_n2671__));
  buf1  g1827(.din(new_new_n1642__), .dout(new_new_n2672__));
  buf1  g1828(.din(new_new_n2672__), .dout(new_new_n2673__));
  buf1  g1829(.din(new_new_n2673__), .dout(new_new_n2674__));
  buf1  g1830(.din(new_new_n2673__), .dout(new_new_n2675__));
  buf1  g1831(.din(new_new_n2672__), .dout(new_new_n2676__));
  buf1  g1832(.din(new_new_n2676__), .dout(new_new_n2677__));
  buf1  g1833(.din(new_new_n1652__), .dout(new_new_n2678__));
  buf1  g1834(.din(new_new_n902__), .dout(new_new_n2679__));
  buf1  g1835(.din(new_new_n1651__), .dout(new_new_n2680__));
  buf1  g1836(.din(new_new_n901__), .dout(new_new_n2681__));
  buf1  g1837(.din(new_new_n884__), .dout(new_new_n2682__));
  buf1  g1838(.din(new_new_n2682__), .dout(new_new_n2683__));
  buf1  g1839(.din(new_new_n2683__), .dout(new_new_n2684__));
  buf1  g1840(.din(new_new_n2683__), .dout(new_new_n2685__));
  buf1  g1841(.din(new_new_n2682__), .dout(new_new_n2686__));
  buf1  g1842(.din(new_new_n883__), .dout(new_new_n2687__));
  buf1  g1843(.din(new_new_n2687__), .dout(new_new_n2688__));
  buf1  g1844(.din(new_new_n2688__), .dout(new_new_n2689__));
  buf1  g1845(.din(new_new_n2688__), .dout(new_new_n2690__));
  buf1  g1846(.din(new_new_n2687__), .dout(new_new_n2691__));
  buf1  g1847(.din(new_new_n1641__), .dout(new_new_n2692__));
  buf1  g1848(.din(new_new_n2692__), .dout(new_new_n2693__));
  buf1  g1849(.din(new_new_n2693__), .dout(new_new_n2694__));
  buf1  g1850(.din(new_new_n2693__), .dout(new_new_n2695__));
  buf1  g1851(.din(new_new_n2692__), .dout(new_new_n2696__));
  buf1  g1852(.din(new_new_n895__), .dout(new_new_n2697__));
  buf1  g1853(.din(new_new_n2697__), .dout(new_new_n2698__));
  buf1  g1854(.din(new_new_n2698__), .dout(new_new_n2699__));
  buf1  g1855(.din(new_new_n2697__), .dout(new_new_n2700__));
  buf1  g1856(.din(new_new_n1668__), .dout(new_new_n2701__));
  buf1  g1857(.din(new_new_n2701__), .dout(new_new_n2702__));
  buf1  g1858(.din(new_new_n2702__), .dout(new_new_n2703__));
  buf1  g1859(.din(new_new_n2702__), .dout(new_new_n2704__));
  buf1  g1860(.din(new_new_n2701__), .dout(new_new_n2705__));
  buf1  g1861(.din(new_new_n1676__), .dout(new_new_n2706__));
  buf1  g1862(.din(new_new_n1670__), .dout(new_new_n2707__));
  buf1  g1863(.din(new_new_n1677__), .dout(new_new_n2708__));
  buf1  g1864(.din(new_new_n1671__), .dout(new_new_n2709__));
  buf1  g1865(.din(new_new_n896__), .dout(new_new_n2710__));
  buf1  g1866(.din(new_new_n2710__), .dout(new_new_n2711__));
  buf1  g1867(.din(new_new_n2710__), .dout(new_new_n2712__));
  buf1  g1868(.din(new_new_n1022__), .dout(new_new_n2713__));
  buf1  g1869(.din(new_new_n1021__), .dout(new_new_n2714__));
  buf1  g1870(.din(new_new_n1739__), .dout(new_new_n2715__));
  buf1  g1871(.din(new_new_n1732__), .dout(new_new_n2716__));
  buf1  g1872(.din(new_new_n1738__), .dout(new_new_n2717__));
  buf1  g1873(.din(new_new_n1733__), .dout(new_new_n2718__));
  buf1  g1874(.din(new_new_n1774__), .dout(new_new_n2719__));
  buf1  g1875(.din(new_new_n1767__), .dout(new_new_n2720__));
  buf1  g1876(.din(new_new_n1773__), .dout(new_new_n2721__));
  buf1  g1877(.din(new_new_n1768__), .dout(new_new_n2722__));
  buf1  g1878(.din(new_new_n1797__), .dout(new_new_n2723__));
  buf1  g1879(.din(new_new_n1793__), .dout(new_new_n2724__));
  buf1  g1880(.din(new_new_n1796__), .dout(new_new_n2725__));
  buf1  g1881(.din(new_new_n1792__), .dout(new_new_n2726__));
  buf1  g1882(.din(new_new_n899__), .dout(new_new_n2727__));
  buf1  g1883(.din(new_new_n897__), .dout(new_new_n2728__));
  buf1  g1884(.din(new_new_n900__), .dout(new_new_n2729__));
  buf1  g1885(.din(new_new_n898__), .dout(new_new_n2730__));
  buf1  g1886(.din(new_new_n1269__), .dout(new_new_n2731__));
  buf1  g1887(.din(new_new_n2731__), .dout(new_new_n2732__));
  buf1  g1888(.din(new_new_n1011__), .dout(new_new_n2733__));
  buf1  g1889(.din(new_new_n1270__), .dout(new_new_n2734__));
  buf1  g1890(.din(new_new_n1271__), .dout(new_new_n2735__));
  buf1  g1891(.din(new_new_n2735__), .dout(new_new_n2736__));
  buf1  g1892(.din(new_new_n1111__), .dout(new_new_n2737__));
  buf1  g1893(.din(new_new_n1272__), .dout(new_new_n2738__));
  buf1  g1894(.din(new_new_n1275__), .dout(new_new_n2739__));
  buf1  g1895(.din(new_new_n1262__), .dout(new_new_n2740__));
  buf1  g1896(.din(new_new_n2740__), .dout(new_new_n2741__));
  buf1  g1897(.din(new_new_n2741__), .dout(new_new_n2742__));
  buf1  g1898(.din(new_new_n2741__), .dout(new_new_n2743__));
  buf1  g1899(.din(new_new_n2740__), .dout(new_new_n2744__));
  buf1  g1900(.din(new_new_n1261__), .dout(new_new_n2745__));
  buf1  g1901(.din(new_new_n2745__), .dout(new_new_n2746__));
  buf1  g1902(.din(new_new_n2746__), .dout(new_new_n2747__));
  buf1  g1903(.din(new_new_n2746__), .dout(new_new_n2748__));
  buf1  g1904(.din(new_new_n2745__), .dout(new_new_n2749__));
  buf1  g1905(.din(new_new_n1277__), .dout(new_new_n2750__));
  buf1  g1906(.din(new_new_n1281__), .dout(new_new_n2751__));
  buf1  g1907(.din(new_new_n1341__), .dout(new_new_n2752__));
  buf1  g1908(.din(new_new_n1184__), .dout(new_new_n2753__));
  buf1  g1909(.din(new_new_n2753__), .dout(new_new_n2754__));
  buf1  g1910(.din(new_new_n2753__), .dout(new_new_n2755__));
  buf1  g1911(.din(new_new_n1183__), .dout(new_new_n2756__));
  buf1  g1912(.din(new_new_n2756__), .dout(new_new_n2757__));
  buf1  g1913(.din(new_new_n2756__), .dout(new_new_n2758__));
  buf1  g1914(.din(new_new_n1315__), .dout(new_new_n2759__));
  buf1  g1915(.din(new_new_n1827__), .dout(new_new_n2760__));
  buf1  g1916(.din(new_new_n1814__), .dout(new_new_n2761__));
  buf1  g1917(.din(new_new_n1249__), .dout(new_new_n2762__));
  buf1  g1918(.din(new_new_n2762__), .dout(new_new_n2763__));
  buf1  g1919(.din(new_new_n1828__), .dout(new_new_n2764__));
  buf1  g1920(.din(new_new_n1843__), .dout(new_new_n2765__));
  buf1  g1921(.din(new_new_n2765__), .dout(new_new_n2766__));
  buf1  g1922(.din(new_new_n1830__), .dout(new_new_n2767__));
  buf1  g1923(.din(new_new_n1846__), .dout(new_new_n2768__));
  buf1  g1924(.din(new_new_n2768__), .dout(new_new_n2769__));
  buf1  g1925(.din(new_new_n1832__), .dout(new_new_n2770__));
  buf1  g1926(.din(new_new_n1178__), .dout(new_new_n2771__));
  buf1  g1927(.din(new_new_n978__), .dout(new_new_n2772__));
  buf1  g1928(.din(new_new_n2772__), .dout(new_new_n2773__));
  buf1  g1929(.din(new_new_n1834__), .dout(new_new_n2774__));
  buf1  g1930(.din(new_new_n2774__), .dout(new_new_n2775__));
  buf1  g1931(.din(new_new_n2774__), .dout(new_new_n2776__));
  buf1  g1932(.din(new_new_n1853__), .dout(new_new_n2777__));
  buf1  g1933(.din(new_new_n1823__), .dout(new_new_n2778__));
  buf1  g1934(.din(new_new_n1816__), .dout(new_new_n2779__));
  buf1  g1935(.din(new_new_n1825__), .dout(new_new_n2780__));
  buf1  g1936(.din(new_new_n1251__), .dout(new_new_n2781__));
  buf1  g1937(.din(new_new_n2781__), .dout(new_new_n2782__));
  buf1  g1938(.din(new_new_n1255__), .dout(new_new_n2783__));
  buf1  g1939(.din(new_new_n2783__), .dout(new_new_n2784__));
  buf1  g1940(.din(new_new_n1818__), .dout(new_new_n2785__));
  buf1  g1941(.din(new_new_n1253__), .dout(new_new_n2786__));
  buf1  g1942(.din(new_new_n2786__), .dout(new_new_n2787__));
  buf1  g1943(.din(new_new_n1820__), .dout(new_new_n2788__));
  buf1  g1944(.din(new_new_n1876__), .dout(new_new_n2789__));
  buf1  g1945(.din(new_new_n1368__), .dout(new_new_n2790__));
  buf1  g1946(.din(new_new_n1875__), .dout(new_new_n2791__));
  buf1  g1947(.din(new_new_n1367__), .dout(new_new_n2792__));
  buf1  g1948(.din(new_new_n2792__), .dout(new_new_n2793__));
  buf1  g1949(.din(new_new_n1860__), .dout(new_new_n2794__));
  buf1  g1950(.din(new_new_n2794__), .dout(new_new_n2795__));
  buf1  g1951(.din(new_new_n2794__), .dout(new_new_n2796__));
  buf1  g1952(.din(new_new_n1847__), .dout(new_new_n2797__));
  buf1  g1953(.din(new_new_n1867__), .dout(new_new_n2798__));
  buf1  g1954(.din(new_new_n2798__), .dout(new_new_n2799__));
  buf1  g1955(.din(new_new_n2799__), .dout(new_new_n2800__));
  buf1  g1956(.din(new_new_n2799__), .dout(new_new_n2801__));
  buf1  g1957(.din(new_new_n2798__), .dout(new_new_n2802__));
  buf1  g1958(.din(new_new_n2802__), .dout(new_new_n2803__));
  buf1  g1959(.din(new_new_n1874__), .dout(new_new_n2804__));
  buf1  g1960(.din(new_new_n2804__), .dout(new_new_n2805__));
  buf1  g1961(.din(new_new_n2805__), .dout(new_new_n2806__));
  buf1  g1962(.din(new_new_n2805__), .dout(new_new_n2807__));
  buf1  g1963(.din(new_new_n2804__), .dout(new_new_n2808__));
  buf1  g1964(.din(new_new_n2808__), .dout(new_new_n2809__));
  buf1  g1965(.din(new_new_n1858__), .dout(new_new_n2810__));
  buf1  g1966(.din(new_new_n2810__), .dout(new_new_n2811__));
  buf1  g1967(.din(new_new_n2810__), .dout(new_new_n2812__));
  buf1  g1968(.din(new_new_n1859__), .dout(new_new_n2813__));
  buf1  g1969(.din(new_new_n2813__), .dout(new_new_n2814__));
  buf1  g1970(.din(new_new_n2813__), .dout(new_new_n2815__));
  buf1  g1971(.din(new_new_n1848__), .dout(new_new_n2816__));
  buf1  g1972(.din(new_new_n1898__), .dout(new_new_n2817__));
  buf1  g1973(.din(new_new_n1854__), .dout(new_new_n2818__));
  buf1  g1974(.din(new_new_n2818__), .dout(new_new_n2819__));
  buf1  g1975(.din(new_new_n1903__), .dout(new_new_n2820__));
  buf1  g1976(.din(new_new_n1399__), .dout(new_new_n2821__));
  buf1  g1977(.din(new_new_n1397__), .dout(new_new_n2822__));
  buf1  g1978(.din(new_new_n1400__), .dout(new_new_n2823__));
  buf1  g1979(.din(new_new_n1398__), .dout(new_new_n2824__));
  buf1  g1980(.din(new_new_n1407__), .dout(new_new_n2825__));
  buf1  g1981(.din(new_new_n2825__), .dout(new_new_n2826__));
  buf1  g1982(.din(new_new_n2825__), .dout(new_new_n2827__));
  buf1  g1983(.din(new_new_n1408__), .dout(new_new_n2828__));
  buf1  g1984(.din(new_new_n2828__), .dout(new_new_n2829__));
  buf1  g1985(.din(new_new_n2828__), .dout(new_new_n2830__));
  buf1  g1986(.din(new_new_n1415__), .dout(new_new_n2831__));
  buf1  g1987(.din(new_new_n1409__), .dout(new_new_n2832__));
  buf1  g1988(.din(new_new_n1416__), .dout(new_new_n2833__));
  buf1  g1989(.din(new_new_n1410__), .dout(new_new_n2834__));
  buf1  g1990(.din(new_new_n1401__), .dout(new_new_n2835__));
  buf1  g1991(.din(new_new_n2835__), .dout(new_new_n2836__));
  buf1  g1992(.din(new_new_n2835__), .dout(new_new_n2837__));
  buf1  g1993(.din(new_new_n1402__), .dout(new_new_n2838__));
  buf1  g1994(.din(new_new_n1405__), .dout(new_new_n2839__));
  buf1  g1995(.din(new_new_n2839__), .dout(new_new_n2840__));
  buf1  g1996(.din(new_new_n1406__), .dout(new_new_n2841__));
  buf1  g1997(.din(new_new_n1944__), .dout(new_new_n2842__));
  buf1  g1998(.din(new_new_n1028__), .dout(new_new_n2843__));
  buf1  g1999(.din(new_new_n1948__), .dout(new_new_n2844__));
  buf1  g2000(.din(new_new_n1053__), .dout(new_new_n2845__));
  buf1  g2001(.din(new_new_n1953__), .dout(new_new_n2846__));
  buf1  g2002(.din(new_new_n965__), .dout(new_new_n2847__));
  buf1  g2003(.din(new_new_n1952__), .dout(new_new_n2848__));
  buf1  g2004(.din(new_new_n966__), .dout(new_new_n2849__));
  buf1  g2005(.din(new_new_n1965__), .dout(new_new_n2850__));
  buf1  g2006(.din(new_new_n1962__), .dout(new_new_n2851__));
  buf1  g2007(.din(new_new_n1905__), .dout(new_new_n2852__));
  buf1  g2008(.din(new_new_n2852__), .dout(new_new_n2853__));
  buf1  g2009(.din(new_new_n2853__), .dout(new_new_n2854__));
  buf1  g2010(.din(new_new_n2853__), .dout(new_new_n2855__));
  buf1  g2011(.din(new_new_n2852__), .dout(new_new_n2856__));
  buf1  g2012(.din(new_new_n1900__), .dout(new_new_n2857__));
  buf1  g2013(.din(new_new_n1895__), .dout(new_new_n2858__));
  buf1  g2014(.din(new_new_n2858__), .dout(new_new_n2859__));
  buf1  g2015(.din(new_new_n2859__), .dout(new_new_n2860__));
  buf1  g2016(.din(new_new_n2859__), .dout(new_new_n2861__));
  buf1  g2017(.din(new_new_n2858__), .dout(new_new_n2862__));
  buf1  g2018(.din(new_new_n2862__), .dout(new_new_n2863__));
  buf1  g2019(.din(new_new_n2862__), .dout(new_new_n2864__));
  buf1  g2020(.din(new_new_n1904__), .dout(new_new_n2865__));
  buf1  g2021(.din(new_new_n2865__), .dout(new_new_n2866__));
  buf1  g2022(.din(new_new_n2866__), .dout(new_new_n2867__));
  buf1  g2023(.din(new_new_n2865__), .dout(new_new_n2868__));
  buf1  g2024(.din(new_new_n1899__), .dout(new_new_n2869__));
  buf1  g2025(.din(new_new_n2869__), .dout(new_new_n2870__));
  buf1  g2026(.din(new_new_n2870__), .dout(new_new_n2871__));
  buf1  g2027(.din(new_new_n2870__), .dout(new_new_n2872__));
  buf1  g2028(.din(new_new_n2869__), .dout(new_new_n2873__));
  buf1  g2029(.din(new_new_n2873__), .dout(new_new_n2874__));
  buf1  g2030(.din(new_new_n2873__), .dout(new_new_n2875__));
  buf1  g2031(.din(new_new_n1311__), .dout(new_new_n2876__));
  buf1  g2032(.din(new_new_n1303__), .dout(new_new_n2877__));
  buf1  g2033(.din(new_new_n2877__), .dout(new_new_n2878__));
  buf1  g2034(.din(new_new_n1312__), .dout(new_new_n2879__));
  buf1  g2035(.din(new_new_n1304__), .dout(new_new_n2880__));
  buf1  g2036(.din(new_new_n1417__), .dout(new_new_n2881__));
  buf1  g2037(.din(new_new_n1411__), .dout(new_new_n2882__));
  buf1  g2038(.din(new_new_n1418__), .dout(new_new_n2883__));
  buf1  g2039(.din(new_new_n1412__), .dout(new_new_n2884__));
  buf1  g2040(.din(new_new_n1403__), .dout(new_new_n2885__));
  buf1  g2041(.din(new_new_n2885__), .dout(new_new_n2886__));
  buf1  g2042(.din(new_new_n2885__), .dout(new_new_n2887__));
  buf1  g2043(.din(new_new_n1069__), .dout(new_new_n2888__));
  buf1  g2044(.din(new_new_n1067__), .dout(new_new_n2889__));
  buf1  g2045(.din(new_new_n2889__), .dout(new_new_n2890__));
  buf1  g2046(.din(new_new_n2889__), .dout(new_new_n2891__));
  buf1  g2047(.din(new_new_n1169__), .dout(new_new_n2892__));
  buf1  g2048(.din(new_new_n881__), .dout(new_new_n2893__));
  buf1  g2049(.din(new_new_n2893__), .dout(new_new_n2894__));
  buf1  g2050(.din(new_new_n2893__), .dout(new_new_n2895__));
  buf1  g2051(.din(new_new_n1343__), .dout(new_new_n2896__));
  buf1  g2052(.din(new_new_n2896__), .dout(new_new_n2897__));
  buf1  g2053(.din(new_new_n2896__), .dout(new_new_n2898__));
  buf1  g2054(.din(new_new_n1353__), .dout(new_new_n2899__));
  buf1  g2055(.din(new_new_n1318__), .dout(new_new_n2900__));
  buf1  g2056(.din(new_new_n1354__), .dout(new_new_n2901__));
  buf1  g2057(.din(new_new_n1317__), .dout(new_new_n2902__));
  buf1  g2058(.din(new_new_n1351__), .dout(new_new_n2903__));
  buf1  g2059(.din(new_new_n1320__), .dout(new_new_n2904__));
  buf1  g2060(.din(new_new_n1352__), .dout(new_new_n2905__));
  buf1  g2061(.din(new_new_n1319__), .dout(new_new_n2906__));
  buf1  g2062(.din(new_new_n2011__), .dout(new_new_n2907__));
  buf1  g2063(.din(new_new_n2006__), .dout(new_new_n2908__));
  buf1  g2064(.din(new_new_n2012__), .dout(new_new_n2909__));
  buf1  g2065(.din(new_new_n2005__), .dout(new_new_n2910__));
  buf1  g2066(.din(new_new_n1344__), .dout(new_new_n2911__));
  buf1  g2067(.din(new_new_n821__), .dout(new_new_n2912__));
  buf1  g2068(.din(new_new_n1358__), .dout(new_new_n2913__));
  buf1  g2069(.din(new_new_n1331__), .dout(new_new_n2914__));
  buf1  g2070(.din(new_new_n1357__), .dout(new_new_n2915__));
  buf1  g2071(.din(new_new_n1332__), .dout(new_new_n2916__));
  buf1  g2072(.din(new_new_n1349__), .dout(new_new_n2917__));
  buf1  g2073(.din(new_new_n1324__), .dout(new_new_n2918__));
  buf1  g2074(.din(new_new_n1350__), .dout(new_new_n2919__));
  buf1  g2075(.din(new_new_n1323__), .dout(new_new_n2920__));
  buf1  g2076(.din(new_new_n2036__), .dout(new_new_n2921__));
  buf1  g2077(.din(new_new_n2031__), .dout(new_new_n2922__));
  buf1  g2078(.din(new_new_n2037__), .dout(new_new_n2923__));
  buf1  g2079(.din(new_new_n2030__), .dout(new_new_n2924__));
  buf1  g2080(.din(new_new_n1327__), .dout(new_new_n2925__));
  buf1  g2081(.din(new_new_n1322__), .dout(new_new_n2926__));
  buf1  g2082(.din(new_new_n1328__), .dout(new_new_n2927__));
  buf1  g2083(.din(new_new_n1321__), .dout(new_new_n2928__));
  buf1  g2084(.din(new_new_n2049__), .dout(new_new_n2929__));
  buf1  g2085(.din(new_new_n1052__), .dout(new_new_n2930__));
  buf1  g2086(.din(new_new_n2048__), .dout(new_new_n2931__));
  buf1  g2087(.din(new_new_n1051__), .dout(new_new_n2932__));
  buf1  g2088(.din(new_new_n1345__), .dout(new_new_n2933__));
  buf1  g2089(.din(new_new_n1325__), .dout(new_new_n2934__));
  buf1  g2090(.din(new_new_n1346__), .dout(new_new_n2935__));
  buf1  g2091(.din(new_new_n1326__), .dout(new_new_n2936__));
  buf1  g2092(.din(new_new_n2064__), .dout(new_new_n2937__));
  buf1  g2093(.din(new_new_n1839__), .dout(new_new_n2938__));
  buf1  g2094(.din(new_new_n2938__), .dout(new_new_n2939__));
  buf1  g2095(.din(new_new_n2063__), .dout(new_new_n2940__));
  buf1  g2096(.din(new_new_n1840__), .dout(new_new_n2941__));
  buf1  g2097(.din(new_new_n2076__), .dout(new_new_n2942__));
  buf1  g2098(.din(new_new_n1233__), .dout(new_new_n2943__));
  buf1  g2099(.din(new_new_n2943__), .dout(new_new_n2944__));
  buf1  g2100(.din(new_new_n2943__), .dout(new_new_n2945__));
  buf1  g2101(.din(new_new_n2075__), .dout(new_new_n2946__));
  buf1  g2102(.din(new_new_n1234__), .dout(new_new_n2947__));
  buf1  g2103(.din(new_new_n2097__), .dout(new_new_n2948__));
  buf1  g2104(.din(new_new_n2090__), .dout(new_new_n2949__));
  buf1  g2105(.din(new_new_n2096__), .dout(new_new_n2950__));
  buf1  g2106(.din(new_new_n2091__), .dout(new_new_n2951__));
  buf1  g2107(.din(new_new_n1313__), .dout(new_new_n2952__));
  buf1  g2108(.din(new_new_n2106__), .dout(new_new_n2953__));
  buf1  g2109(.din(new_new_n1068__), .dout(new_new_n2954__));
  buf1  g2110(.din(new_new_n2107__), .dout(new_new_n2955__));
  buf1  g2111(.din(new_new_n1837__), .dout(new_new_n2956__));
  buf1  g2112(.din(new_new_n2956__), .dout(new_new_n2957__));
  buf1  g2113(.din(new_new_n1075__), .dout(new_new_n2958__));
  buf1  g2114(.din(new_new_n2958__), .dout(new_new_n2959__));
  buf1  g2115(.din(new_new_n1838__), .dout(new_new_n2960__));
  buf1  g2116(.din(new_new_n1076__), .dout(new_new_n2961__));
  buf1  g2117(.din(new_new_n2128__), .dout(new_new_n2962__));
  buf1  g2118(.din(new_new_n1356__), .dout(new_new_n2963__));
  buf1  g2119(.din(new_new_n2127__), .dout(new_new_n2964__));
  buf1  g2120(.din(new_new_n1355__), .dout(new_new_n2965__));
  buf1  g2121(.din(new_new_n2965__), .dout(new_new_n2966__));
  buf1  g2122(.din(new_new_n1380__), .dout(new_new_n2967__));
  buf1  g2123(.din(new_new_n2967__), .dout(new_new_n2968__));
  buf1  g2124(.din(new_new_n1379__), .dout(new_new_n2969__));
  buf1  g2125(.din(new_new_n2969__), .dout(new_new_n2970__));
  buf1  g2126(.din(new_new_n2142__), .dout(new_new_n2971__));
  buf1  g2127(.din(new_new_n1329__), .dout(new_new_n2972__));
  buf1  g2128(.din(new_new_n2972__), .dout(new_new_n2973__));
  buf1  g2129(.din(new_new_n2141__), .dout(new_new_n2974__));
  buf1  g2130(.din(new_new_n1330__), .dout(new_new_n2975__));
  buf1  g2131(.din(new_new_n1881__), .dout(new_new_n2976__));
  buf1  g2132(.din(new_new_n796__), .dout(new_new_n2977__));
  buf1  g2133(.din(new_new_n2977__), .dout(new_new_n2978__));
  buf1  g2134(.din(new_new_n1395__), .dout(new_new_n2979__));
  buf1  g2135(.din(new_new_n2979__), .dout(new_new_n2980__));
  buf1  g2136(.din(new_new_n2980__), .dout(new_new_n2981__));
  buf1  g2137(.din(new_new_n2979__), .dout(new_new_n2982__));
  buf1  g2138(.din(new_new_n795__), .dout(new_new_n2983__));
  buf1  g2139(.din(new_new_n2983__), .dout(new_new_n2984__));
  buf1  g2140(.din(new_new_n2983__), .dout(new_new_n2985__));
  buf1  g2141(.din(new_new_n894__), .dout(new_new_n2986__));
  buf1  g2142(.din(new_new_n827__), .dout(new_new_n2987__));
  buf1  g2143(.din(new_new_n1914__), .dout(new_new_n2988__));
  buf1  g2144(.din(new_new_n2988__), .dout(new_new_n2989__));
  buf1  g2145(.din(new_new_n2989__), .dout(new_new_n2990__));
  buf1  g2146(.din(new_new_n2989__), .dout(new_new_n2991__));
  buf1  g2147(.din(new_new_n2988__), .dout(new_new_n2992__));
  buf1  g2148(.din(new_new_n1932__), .dout(new_new_n2993__));
  buf1  g2149(.din(new_new_n2993__), .dout(new_new_n2994__));
  buf1  g2150(.din(new_new_n1923__), .dout(new_new_n2995__));
  buf1  g2151(.din(new_new_n2995__), .dout(new_new_n2996__));
  buf1  g2152(.din(new_new_n817__), .dout(new_new_n2997__));
  buf1  g2153(.din(new_new_n837__), .dout(new_new_n2998__));
  buf1  g2154(.din(new_new_n2998__), .dout(new_new_n2999__));
  buf1  g2155(.din(new_new_n893__), .dout(new_new_n3000__));
  buf1  g2156(.din(new_new_n3000__), .dout(new_new_n3001__));
  buf1  g2157(.din(new_new_n1247__), .dout(new_new_n3002__));
  buf1  g2158(.din(new_new_n1248__), .dout(new_new_n3003__));
  buf1  g2159(.din(new_new_n791__), .dout(new_new_n3004__));
  buf1  g2160(.din(new_new_n3004__), .dout(new_new_n3005__));
  buf1  g2161(.din(new_new_n3004__), .dout(new_new_n3006__));
  buf1  g2162(.din(new_new_n792__), .dout(new_new_n3007__));
  buf1  g2163(.din(new_new_n1385__), .dout(new_new_n3008__));
  buf1  g2164(.din(new_new_n1386__), .dout(new_new_n3009__));
  buf1  g2165(.din(new_new_n781__), .dout(new_new_n3010__));
  buf1  g2166(.din(new_new_n3010__), .dout(new_new_n3011__));
  buf1  g2167(.din(new_new_n3011__), .dout(new_new_n3012__));
  buf1  g2168(.din(new_new_n3011__), .dout(new_new_n3013__));
  buf1  g2169(.din(new_new_n3010__), .dout(new_new_n3014__));
  buf1  g2170(.din(new_new_n867__), .dout(new_new_n3015__));
  buf1  g2171(.din(new_new_n875__), .dout(new_new_n3016__));
  buf1  g2172(.din(new_new_n889__), .dout(new_new_n3017__));
  buf1  g2173(.din(new_new_n977__), .dout(new_new_n3018__));
  buf1  g2174(.din(new_new_n3018__), .dout(new_new_n3019__));
  buf1  g2175(.din(new_new_n1025__), .dout(new_new_n3020__));
  buf1  g2176(.din(new_new_n1035__), .dout(new_new_n3021__));
  buf1  g2177(.din(new_new_n1041__), .dout(new_new_n3022__));
  buf1  g2178(.din(new_new_n1885__), .dout(new_new_n3023__));
  buf1  g2179(.din(new_new_n1888__), .dout(new_new_n3024__));
  buf1  g2180(.din(new_new_n1891__), .dout(new_new_n3025__));
  buf1  g2181(.din(new_new_n1941__), .dout(new_new_n3026__));
  buf1  g2182(.din(new_new_n3026__), .dout(new_new_n3027__));
  buf1  g2183(.din(new_new_n3026__), .dout(new_new_n3028__));
  buf1  g2184(.din(new_new_n711__), .dout(new_new_n3029__));
  buf1  g2185(.din(new_new_n3029__), .dout(new_new_n3030__));
  buf1  g2186(.din(new_new_n3030__), .dout(new_new_n3031__));
  buf1  g2187(.din(new_new_n3029__), .dout(new_new_n3032__));
  buf1  g2188(.din(new_new_n737__), .dout(new_new_n3033__));
  buf1  g2189(.din(new_new_n3033__), .dout(new_new_n3034__));
  buf1  g2190(.din(new_new_n3034__), .dout(new_new_n3035__));
  buf1  g2191(.din(new_new_n3033__), .dout(new_new_n3036__));
  buf1  g2192(.din(new_new_n1987__), .dout(new_new_n3037__));
  buf1  g2193(.din(new_new_n3037__), .dout(new_new_n3038__));
  buf1  g2194(.din(new_new_n1996__), .dout(new_new_n3039__));
  buf1  g2195(.din(new_new_n3039__), .dout(new_new_n3040__));
  buf1  g2196(.din(new_new_n713__), .dout(new_new_n3041__));
  buf1  g2197(.din(new_new_n3041__), .dout(new_new_n3042__));
  buf1  g2198(.din(new_new_n3041__), .dout(new_new_n3043__));
  buf1  g2199(.din(new_new_n719__), .dout(new_new_n3044__));
  buf1  g2200(.din(new_new_n3044__), .dout(new_new_n3045__));
  buf1  g2201(.din(new_new_n3044__), .dout(new_new_n3046__));
  buf1  g2202(.din(new_new_n731__), .dout(new_new_n3047__));
  buf1  g2203(.din(new_new_n3047__), .dout(new_new_n3048__));
  buf1  g2204(.din(new_new_n3047__), .dout(new_new_n3049__));
  buf1  g2205(.din(new_new_n739__), .dout(new_new_n3050__));
  buf1  g2206(.din(new_new_n3050__), .dout(new_new_n3051__));
  buf1  g2207(.din(new_new_n3051__), .dout(new_new_n3052__));
  buf1  g2208(.din(new_new_n3050__), .dout(new_new_n3053__));
  buf1  g2209(.din(new_new_n1309__), .dout(new_new_n3054__));
  buf1  g2210(.din(new_new_n3054__), .dout(new_new_n3055__));
  buf1  g2211(.din(new_new_n2140__), .dout(new_new_n3056__));
  buf1  g2212(.din(new_new_n2154__), .dout(new_new_n3057__));
  buf1  g2213(.din(new_new_n3057__), .dout(new_new_n3058__));
  buf1  g2214(.din(new_new_n721__), .dout(new_new_n3059__));
  buf1  g2215(.din(new_new_n3059__), .dout(new_new_n3060__));
  buf1  g2216(.din(new_new_n733__), .dout(new_new_n3061__));
  buf1  g2217(.din(new_new_n3061__), .dout(new_new_n3062__));
  buf1  g2218(.din(new_new_n709__), .dout(new_new_n3063__));
  buf1  g2219(.din(new_new_n727__), .dout(new_new_n3064__));
  always @ (posedge clock) begin
    n949_lo <= n4857;
    n961_lo <= n4860;
    n973_lo <= n4863;
    n976_lo <= n4866;
    n985_lo <= n4869;
    n997_lo <= n4872;
    n1009_lo <= n4875;
    n1021_lo <= n4878;
    n1024_lo <= n4881;
    n1033_lo <= n4884;
    n1036_lo <= n4887;
    n1045_lo <= n4890;
    n1057_lo <= n4893;
    n1069_lo <= n4896;
    n1081_lo <= n4899;
    n1093_lo <= n4902;
    n1105_lo <= n4905;
    n1117_lo <= n4908;
    n1129_lo <= n4911;
    n1132_lo <= n4914;
    n1141_lo <= n4917;
    n1144_lo <= n4920;
    n1156_lo <= n4923;
    n1159_lo <= n4926;
    n1165_lo <= n4929;
    n1168_lo <= n4932;
    n1180_lo <= n4935;
    n1189_lo <= n4938;
    n1192_lo <= n4941;
    n1201_lo <= n4944;
    n1204_lo <= n4947;
    n1216_lo <= n4950;
    n1228_lo <= n4953;
    n1231_lo <= n4956;
    n1237_lo <= n4959;
    n1240_lo <= n4962;
    n1243_lo <= n4965;
    n1249_lo <= n4968;
    n1252_lo <= n4971;
    n1255_lo <= n4974;
    n1261_lo <= n4977;
    n1264_lo <= n4980;
    n1267_lo <= n4983;
    n1273_lo <= n4986;
    n1276_lo <= n4989;
    n1279_lo <= n4992;
    n1282_lo <= n4995;
    n1285_lo <= n4998;
    n1288_lo <= n5001;
    n1291_lo <= n5004;
    n1294_lo <= n5007;
    n1297_lo <= n5010;
    n1300_lo <= n5013;
    n1303_lo <= n5016;
    n1309_lo <= n5019;
    n1312_lo <= n5022;
    n1315_lo <= n5025;
    n1318_lo <= n5028;
    n1321_lo <= n5031;
    n1324_lo <= n5034;
    n1333_lo <= n5037;
    n1874_o2 <= n5040;
    n2180_o2 <= n5043;
    n2372_o2 <= n5046;
    n2190_o2 <= n5049;
    n2191_o2 <= n5052;
    n2212_o2 <= n5055;
    n2213_o2 <= n5058;
    n2214_o2 <= n5061;
    n2215_o2 <= n5064;
    n2275_o2 <= n5067;
    n2276_o2 <= n5070;
    n2290_o2 <= n5073;
    n2291_o2 <= n5076;
    n2681_o2 <= n5079;
    n2680_o2 <= n5082;
    n2683_o2 <= n5085;
    n2684_o2 <= n5088;
    n2686_o2 <= n5091;
    n2319_o2 <= n5094;
    n2320_o2 <= n5097;
    n304_inv <= n5100;
    G554_o2 <= n5103;
    G557_o2 <= n5106;
    G185_o2 <= n5109;
    G188_o2 <= n5112;
    G191_o2 <= n5115;
    G194_o2 <= n5118;
    G1182_o2 <= n5121;
    G1222_o2 <= n5124;
    G1247_o2 <= n5127;
    G1371_o2 <= n5130;
    G1383_o2 <= n5133;
    G1386_o2 <= n5136;
    n2416_o2 <= n5139;
    n2428_o2 <= n5142;
    n2438_o2 <= n5145;
    n2439_o2 <= n5148;
    n2440_o2 <= n5151;
    n2444_o2 <= n5154;
    n2497_o2 <= n5157;
    n2498_o2 <= n5160;
    n2503_o2 <= n5163;
    n2505_o2 <= n5166;
    n2529_o2 <= n5169;
    n2562_o2 <= n5172;
    n2570_o2 <= n5175;
    n2571_o2 <= n5178;
    n2574_o2 <= n5181;
    n2575_o2 <= n5184;
    G546_o2 <= n5187;
    G550_o2 <= n5190;
    n2633_o2 <= n5193;
    n2639_o2 <= n5196;
    n2642_o2 <= n5199;
    n2645_o2 <= n5202;
    n2679_o2 <= n5205;
    n2662_o2 <= n5208;
    n2724_o2 <= n5211;
    G382_o2 <= n5214;
    G199_o2 <= n5217;
    G202_o2 <= n5220;
    G225_o2 <= n5223;
    G248_o2 <= n5226;
    G260_o2 <= n5229;
    n2716_o2 <= n5232;
    n2737_o2 <= n5235;
    n1174_lo_buf_o2 <= n5238;
    n1198_lo_buf_o2 <= n5241;
    G371_o2 <= n5244;
    G1059_o2 <= n5247;
    n2586_o2 <= n5250;
    n2587_o2 <= n5253;
    n460_inv <= n5256;
    n2648_o2 <= n5259;
    n2649_o2 <= n5262;
    n2650_o2 <= n5265;
    n2651_o2 <= n5268;
    n2652_o2 <= n5271;
    G365_o2 <= n5274;
    G1496_o2 <= n5277;
    G1502_o2 <= n5280;
    n2700_o2 <= n5283;
    n2701_o2 <= n5286;
    n2733_o2 <= n5289;
    n2734_o2 <= n5292;
    n2744_o2 <= n5295;
    n2747_o2 <= n5298;
    n2754_o2 <= n5301;
    n2755_o2 <= n5304;
    n511_inv <= n5307;
    G1609_o2 <= n5310;
    G1625_o2 <= n5313;
    G738_o2 <= n5316;
    G755_o2 <= n5319;
    G1511_o2 <= n5322;
    G1522_o2 <= n5325;
    G1538_o2 <= n5328;
    G1549_o2 <= n5331;
    G1563_o2 <= n5334;
    G1584_o2 <= n5337;
    G1576_o2 <= n5340;
    G1598_o2 <= n5343;
    G1395_o2 <= n5346;
    G1410_o2 <= n5349;
    G1420_o2 <= n5352;
    G1434_o2 <= n5355;
    n562_inv <= n5358;
    n1162_lo_buf_o2 <= n5361;
    n1102_lo_buf_o2 <= n5364;
    G359_o2 <= n5367;
    n982_lo_buf_o2 <= n5370;
    n1030_lo_buf_o2 <= n5373;
    n1042_lo_buf_o2 <= n5376;
    n583_inv <= n5379;
    G606_o2 <= n5382;
    G1118_o2 <= n5385;
    G1069_o2 <= n5388;
    G1145_o2 <= n5391;
    G1209_o2 <= n5394;
    G1189_o2 <= n5397;
    G1699_o2 <= n5400;
    G1702_o2 <= n5403;
    G1705_o2 <= n5406;
    G1708_o2 <= n5409;
    G1684_o2 <= n5412;
    G1687_o2 <= n5415;
    G1690_o2 <= n5418;
    G1693_o2 <= n5421;
    G1696_o2 <= n5424;
    G1642_o2 <= n5427;
    G1645_o2 <= n5430;
    G1648_o2 <= n5433;
    G1651_o2 <= n5436;
    G1654_o2 <= n5439;
    G1657_o2 <= n5442;
    G1660_o2 <= n5445;
    n1222_lo_buf_o2 <= n5448;
    n1330_lo_buf_o2 <= n5451;
    n658_inv <= n5454;
    n661_inv <= n5457;
    n1306_lo_buf_o2 <= n5460;
    n1150_lo_buf_o2 <= n5463;
    G175_o2 <= n5466;
    G241_o2 <= n5469;
    G356_o2 <= n5472;
    G989_o2 <= n5475;
    G984_o2 <= n5478;
    n685_inv <= n5481;
    n688_inv <= n5484;
    n958_lo_buf_o2 <= n5487;
    n1114_lo_buf_o2 <= n5490;
    G182_o2 <= n5493;
    G1215_o2 <= n5496;
    G971_o2 <= n5499;
    G938_o2 <= n5502;
    G1198_o2 <= n5505;
    G1203_o2 <= n5508;
    G1218_o2 <= n5511;
    G785_o2 <= n5514;
    G1168_o2 <= n5517;
    G1130_o2 <= n5520;
    G1185_o2 <= n5523;
    G1250_o2 <= n5526;
    G1225_o2 <= n5529;
    G1791_o2 <= n5532;
    G1788_o2 <= n5535;
    G981_o2 <= n5538;
    n745_inv <= n5541;
    n748_inv <= n5544;
    G1062_o2 <= n5547;
    n970_lo_buf_o2 <= n5550;
    n1006_lo_buf_o2 <= n5553;
    n1078_lo_buf_o2 <= n5556;
    n1126_lo_buf_o2 <= n5559;
    n766_inv <= n5562;
    G165_o2 <= n5565;
    n1234_lo_buf_o2 <= n5568;
    n1246_lo_buf_o2 <= n5571;
    n1258_lo_buf_o2 <= n5574;
    n1270_lo_buf_o2 <= n5577;
    G368_o2 <= n5580;
    G428_o2 <= n5583;
    G212_o2 <= n5586;
    G841_o2 <= n5589;
    G788_o2 <= n5592;
    n1186_lo_buf_o2 <= n5595;
    G391_o2 <= n5598;
    G387_o2 <= n5601;
    G645_o2 <= n5604;
    G1140_o2 <= n5607;
    G1178_o2 <= n5610;
    G1370_o2 <= n5613;
    n820_inv <= n5616;
    G1357_o2 <= n5619;
    G816_o2 <= n5622;
    G1369_o2 <= n5625;
    G901_o2 <= n5628;
    G1056_o2 <= n5631;
    G1107_o2 <= n5634;
    G1087_o2 <= n5637;
    G1135_o2 <= n5640;
    n1018_lo_buf_o2 <= n5643;
    n1090_lo_buf_o2 <= n5646;
    n853_inv <= n5649;
    G131_o2 <= n5652;
    n859_inv <= n5655;
    n862_inv <= n5658;
    G338_o2 <= n5661;
    n1171_lo_buf_o2 <= n5664;
    n1195_lo_buf_o2 <= n5667;
    G419_o2 <= n5670;
    G425_o2 <= n5673;
    G497_o2 <= n5676;
    G416_o2 <= n5679;
    G491_o2 <= n5682;
    G500_o2 <= n5685;
    G353_o2 <= n5688;
    G641_o2 <= n5691;
    G1117_o2 <= n5694;
    G1096_o2 <= n5697;
    G1143_o2 <= n5700;
    G1112_o2 <= n5703;
    n1138_lo_buf_o2 <= n5706;
    n1210_lo_buf_o2 <= n5709;
    G687_o2 <= n5712;
    G541_o2 <= n5715;
    G802_o2 <= n5718;
    G813_o2 <= n5721;
    G810_o2 <= n5724;
    G987_o2 <= n5727;
    G898_o2 <= n5730;
    n946_lo_buf_o2 <= n5733;
    n1054_lo_buf_o2 <= n5736;
    G728_o2 <= n5739;
    G856_o2 <= n5742;
    n949_1_inv <= n5745;
    G942_o2 <= n5748;
    G1099_o2 <= n5751;
    G1154_o2 <= n5754;
    G1131_o2 <= n5757;
    G1169_o2 <= n5760;
    G134_o2 <= n5763;
    n970_inv <= n5766;
    G470_o2 <= n5769;
    G344_o2 <= n5772;
    G362_o2 <= n5775;
    G482_o2 <= n5778;
    G660_o2 <= n5781;
    G672_o2 <= n5784;
    n1096_lo_buf_o2 <= n5787;
    G479_o2 <= n5790;
    G669_o2 <= n5793;
    n994_lo_buf_o2 <= n5796;
    n1066_lo_buf_o2 <= n5799;
    n1006_inv <= n5802;
    G147_o2 <= n5805;
    G473_o2 <= n5808;
    G488_o2 <= n5811;
    G589_o2 <= n5814;
    G663_o2 <= n5817;
    G684_o2 <= n5820;
    G605_o2 <= n5823;
    G774_o2 <= n5826;
    G782_o2 <= n5829;
  end
  initial begin
    n949_lo <= 1'b0;
    n961_lo <= 1'b0;
    n973_lo <= 1'b0;
    n976_lo <= 1'b0;
    n985_lo <= 1'b0;
    n997_lo <= 1'b0;
    n1009_lo <= 1'b0;
    n1021_lo <= 1'b0;
    n1024_lo <= 1'b0;
    n1033_lo <= 1'b0;
    n1036_lo <= 1'b0;
    n1045_lo <= 1'b0;
    n1057_lo <= 1'b0;
    n1069_lo <= 1'b0;
    n1081_lo <= 1'b0;
    n1093_lo <= 1'b0;
    n1105_lo <= 1'b0;
    n1117_lo <= 1'b0;
    n1129_lo <= 1'b0;
    n1132_lo <= 1'b0;
    n1141_lo <= 1'b0;
    n1144_lo <= 1'b0;
    n1156_lo <= 1'b0;
    n1159_lo <= 1'b0;
    n1165_lo <= 1'b0;
    n1168_lo <= 1'b0;
    n1180_lo <= 1'b0;
    n1189_lo <= 1'b0;
    n1192_lo <= 1'b0;
    n1201_lo <= 1'b0;
    n1204_lo <= 1'b0;
    n1216_lo <= 1'b0;
    n1228_lo <= 1'b0;
    n1231_lo <= 1'b0;
    n1237_lo <= 1'b0;
    n1240_lo <= 1'b0;
    n1243_lo <= 1'b0;
    n1249_lo <= 1'b0;
    n1252_lo <= 1'b0;
    n1255_lo <= 1'b0;
    n1261_lo <= 1'b0;
    n1264_lo <= 1'b0;
    n1267_lo <= 1'b0;
    n1273_lo <= 1'b0;
    n1276_lo <= 1'b0;
    n1279_lo <= 1'b0;
    n1282_lo <= 1'b0;
    n1285_lo <= 1'b0;
    n1288_lo <= 1'b0;
    n1291_lo <= 1'b0;
    n1294_lo <= 1'b0;
    n1297_lo <= 1'b0;
    n1300_lo <= 1'b0;
    n1303_lo <= 1'b0;
    n1309_lo <= 1'b0;
    n1312_lo <= 1'b0;
    n1315_lo <= 1'b0;
    n1318_lo <= 1'b0;
    n1321_lo <= 1'b0;
    n1324_lo <= 1'b0;
    n1333_lo <= 1'b0;
    n1874_o2 <= 1'b0;
    n2180_o2 <= 1'b0;
    n2372_o2 <= 1'b0;
    n2190_o2 <= 1'b0;
    n2191_o2 <= 1'b0;
    n2212_o2 <= 1'b0;
    n2213_o2 <= 1'b0;
    n2214_o2 <= 1'b0;
    n2215_o2 <= 1'b0;
    n2275_o2 <= 1'b0;
    n2276_o2 <= 1'b0;
    n2290_o2 <= 1'b0;
    n2291_o2 <= 1'b0;
    n2681_o2 <= 1'b0;
    n2680_o2 <= 1'b0;
    n2683_o2 <= 1'b0;
    n2684_o2 <= 1'b0;
    n2686_o2 <= 1'b0;
    n2319_o2 <= 1'b0;
    n2320_o2 <= 1'b0;
    n304_inv <= 1'b0;
    G554_o2 <= 1'b0;
    G557_o2 <= 1'b0;
    G185_o2 <= 1'b0;
    G188_o2 <= 1'b0;
    G191_o2 <= 1'b0;
    G194_o2 <= 1'b0;
    G1182_o2 <= 1'b0;
    G1222_o2 <= 1'b0;
    G1247_o2 <= 1'b0;
    G1371_o2 <= 1'b0;
    G1383_o2 <= 1'b0;
    G1386_o2 <= 1'b0;
    n2416_o2 <= 1'b0;
    n2428_o2 <= 1'b0;
    n2438_o2 <= 1'b0;
    n2439_o2 <= 1'b0;
    n2440_o2 <= 1'b0;
    n2444_o2 <= 1'b0;
    n2497_o2 <= 1'b0;
    n2498_o2 <= 1'b0;
    n2503_o2 <= 1'b0;
    n2505_o2 <= 1'b0;
    n2529_o2 <= 1'b0;
    n2562_o2 <= 1'b0;
    n2570_o2 <= 1'b0;
    n2571_o2 <= 1'b0;
    n2574_o2 <= 1'b0;
    n2575_o2 <= 1'b0;
    G546_o2 <= 1'b0;
    G550_o2 <= 1'b0;
    n2633_o2 <= 1'b0;
    n2639_o2 <= 1'b0;
    n2642_o2 <= 1'b0;
    n2645_o2 <= 1'b0;
    n2679_o2 <= 1'b0;
    n2662_o2 <= 1'b0;
    n2724_o2 <= 1'b0;
    G382_o2 <= 1'b0;
    G199_o2 <= 1'b0;
    G202_o2 <= 1'b0;
    G225_o2 <= 1'b0;
    G248_o2 <= 1'b0;
    G260_o2 <= 1'b0;
    n2716_o2 <= 1'b0;
    n2737_o2 <= 1'b0;
    n1174_lo_buf_o2 <= 1'b0;
    n1198_lo_buf_o2 <= 1'b0;
    G371_o2 <= 1'b0;
    G1059_o2 <= 1'b0;
    n2586_o2 <= 1'b0;
    n2587_o2 <= 1'b0;
    n460_inv <= 1'b0;
    n2648_o2 <= 1'b0;
    n2649_o2 <= 1'b0;
    n2650_o2 <= 1'b0;
    n2651_o2 <= 1'b0;
    n2652_o2 <= 1'b0;
    G365_o2 <= 1'b0;
    G1496_o2 <= 1'b0;
    G1502_o2 <= 1'b0;
    n2700_o2 <= 1'b0;
    n2701_o2 <= 1'b0;
    n2733_o2 <= 1'b0;
    n2734_o2 <= 1'b0;
    n2744_o2 <= 1'b0;
    n2747_o2 <= 1'b0;
    n2754_o2 <= 1'b0;
    n2755_o2 <= 1'b0;
    n511_inv <= 1'b0;
    G1609_o2 <= 1'b0;
    G1625_o2 <= 1'b0;
    G738_o2 <= 1'b0;
    G755_o2 <= 1'b0;
    G1511_o2 <= 1'b0;
    G1522_o2 <= 1'b0;
    G1538_o2 <= 1'b0;
    G1549_o2 <= 1'b0;
    G1563_o2 <= 1'b0;
    G1584_o2 <= 1'b0;
    G1576_o2 <= 1'b0;
    G1598_o2 <= 1'b0;
    G1395_o2 <= 1'b0;
    G1410_o2 <= 1'b0;
    G1420_o2 <= 1'b0;
    G1434_o2 <= 1'b0;
    n562_inv <= 1'b0;
    n1162_lo_buf_o2 <= 1'b0;
    n1102_lo_buf_o2 <= 1'b0;
    G359_o2 <= 1'b0;
    n982_lo_buf_o2 <= 1'b0;
    n1030_lo_buf_o2 <= 1'b0;
    n1042_lo_buf_o2 <= 1'b0;
    n583_inv <= 1'b0;
    G606_o2 <= 1'b0;
    G1118_o2 <= 1'b0;
    G1069_o2 <= 1'b0;
    G1145_o2 <= 1'b0;
    G1209_o2 <= 1'b0;
    G1189_o2 <= 1'b0;
    G1699_o2 <= 1'b0;
    G1702_o2 <= 1'b0;
    G1705_o2 <= 1'b0;
    G1708_o2 <= 1'b0;
    G1684_o2 <= 1'b0;
    G1687_o2 <= 1'b0;
    G1690_o2 <= 1'b0;
    G1693_o2 <= 1'b0;
    G1696_o2 <= 1'b0;
    G1642_o2 <= 1'b0;
    G1645_o2 <= 1'b0;
    G1648_o2 <= 1'b0;
    G1651_o2 <= 1'b0;
    G1654_o2 <= 1'b0;
    G1657_o2 <= 1'b0;
    G1660_o2 <= 1'b0;
    n1222_lo_buf_o2 <= 1'b0;
    n1330_lo_buf_o2 <= 1'b0;
    n658_inv <= 1'b0;
    n661_inv <= 1'b0;
    n1306_lo_buf_o2 <= 1'b0;
    n1150_lo_buf_o2 <= 1'b0;
    G175_o2 <= 1'b0;
    G241_o2 <= 1'b0;
    G356_o2 <= 1'b0;
    G989_o2 <= 1'b0;
    G984_o2 <= 1'b0;
    n685_inv <= 1'b0;
    n688_inv <= 1'b0;
    n958_lo_buf_o2 <= 1'b0;
    n1114_lo_buf_o2 <= 1'b0;
    G182_o2 <= 1'b0;
    G1215_o2 <= 1'b0;
    G971_o2 <= 1'b0;
    G938_o2 <= 1'b0;
    G1198_o2 <= 1'b0;
    G1203_o2 <= 1'b0;
    G1218_o2 <= 1'b0;
    G785_o2 <= 1'b0;
    G1168_o2 <= 1'b0;
    G1130_o2 <= 1'b0;
    G1185_o2 <= 1'b0;
    G1250_o2 <= 1'b0;
    G1225_o2 <= 1'b0;
    G1791_o2 <= 1'b0;
    G1788_o2 <= 1'b0;
    G981_o2 <= 1'b0;
    n745_inv <= 1'b0;
    n748_inv <= 1'b0;
    G1062_o2 <= 1'b0;
    n970_lo_buf_o2 <= 1'b0;
    n1006_lo_buf_o2 <= 1'b0;
    n1078_lo_buf_o2 <= 1'b0;
    n1126_lo_buf_o2 <= 1'b0;
    n766_inv <= 1'b0;
    G165_o2 <= 1'b0;
    n1234_lo_buf_o2 <= 1'b0;
    n1246_lo_buf_o2 <= 1'b0;
    n1258_lo_buf_o2 <= 1'b0;
    n1270_lo_buf_o2 <= 1'b0;
    G368_o2 <= 1'b0;
    G428_o2 <= 1'b0;
    G212_o2 <= 1'b0;
    G841_o2 <= 1'b0;
    G788_o2 <= 1'b0;
    n1186_lo_buf_o2 <= 1'b0;
    G391_o2 <= 1'b0;
    G387_o2 <= 1'b0;
    G645_o2 <= 1'b0;
    G1140_o2 <= 1'b0;
    G1178_o2 <= 1'b0;
    G1370_o2 <= 1'b0;
    n820_inv <= 1'b0;
    G1357_o2 <= 1'b0;
    G816_o2 <= 1'b0;
    G1369_o2 <= 1'b0;
    G901_o2 <= 1'b0;
    G1056_o2 <= 1'b0;
    G1107_o2 <= 1'b0;
    G1087_o2 <= 1'b0;
    G1135_o2 <= 1'b0;
    n1018_lo_buf_o2 <= 1'b0;
    n1090_lo_buf_o2 <= 1'b0;
    n853_inv <= 1'b0;
    G131_o2 <= 1'b0;
    n859_inv <= 1'b0;
    n862_inv <= 1'b0;
    G338_o2 <= 1'b0;
    n1171_lo_buf_o2 <= 1'b0;
    n1195_lo_buf_o2 <= 1'b0;
    G419_o2 <= 1'b0;
    G425_o2 <= 1'b0;
    G497_o2 <= 1'b0;
    G416_o2 <= 1'b0;
    G491_o2 <= 1'b0;
    G500_o2 <= 1'b0;
    G353_o2 <= 1'b0;
    G641_o2 <= 1'b0;
    G1117_o2 <= 1'b0;
    G1096_o2 <= 1'b0;
    G1143_o2 <= 1'b0;
    G1112_o2 <= 1'b0;
    n1138_lo_buf_o2 <= 1'b0;
    n1210_lo_buf_o2 <= 1'b0;
    G687_o2 <= 1'b0;
    G541_o2 <= 1'b0;
    G802_o2 <= 1'b0;
    G813_o2 <= 1'b0;
    G810_o2 <= 1'b0;
    G987_o2 <= 1'b0;
    G898_o2 <= 1'b0;
    n946_lo_buf_o2 <= 1'b0;
    n1054_lo_buf_o2 <= 1'b0;
    G728_o2 <= 1'b0;
    G856_o2 <= 1'b0;
    n949_1_inv <= 1'b0;
    G942_o2 <= 1'b0;
    G1099_o2 <= 1'b0;
    G1154_o2 <= 1'b0;
    G1131_o2 <= 1'b0;
    G1169_o2 <= 1'b0;
    G134_o2 <= 1'b0;
    n970_inv <= 1'b0;
    G470_o2 <= 1'b0;
    G344_o2 <= 1'b0;
    G362_o2 <= 1'b0;
    G482_o2 <= 1'b0;
    G660_o2 <= 1'b0;
    G672_o2 <= 1'b0;
    n1096_lo_buf_o2 <= 1'b0;
    G479_o2 <= 1'b0;
    G669_o2 <= 1'b0;
    n994_lo_buf_o2 <= 1'b0;
    n1066_lo_buf_o2 <= 1'b0;
    n1006_inv <= 1'b0;
    G147_o2 <= 1'b0;
    G473_o2 <= 1'b0;
    G488_o2 <= 1'b0;
    G589_o2 <= 1'b0;
    G663_o2 <= 1'b0;
    G684_o2 <= 1'b0;
    G605_o2 <= 1'b0;
    G774_o2 <= 1'b0;
    G782_o2 <= 1'b0;
  end
endmodule


