// Benchmark "mymod" written by ABC on Sun Oct 29 23:44:48 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58,
    G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70, G71, G72,
    G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86,
    G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G109, G110, G111, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G124,
    G125, G126, G127, G128, G129, G130, G131, G132, G133, G134, G135, G136,
    G137, G138, G139, G140, G141, G142, G143, G144, G145, G146, G147, G148,
    G149, G150, G151, G152, G153, G154, G155, G156, G157, G158, G159, G160,
    G161, G162, G163, G164, G165, G166, G167, G168, G169, G170, G171, G172,
    G173, G174, G175, G176, G177, G178,
    G5193, G5194, G5195, G5196, G5197, G5198, G5199, G5200, G5201, G5202,
    G5203, G5204, G5205, G5206, G5207, G5208, G5209, G5210, G5211, G5212,
    G5213, G5214, G5215, G5216, G5217, G5218, G5219, G5220, G5221, G5222,
    G5223, G5224, G5225, G5226, G5227, G5228, G5229, G5230, G5231, G5232,
    G5233, G5234, G5235, G5236, G5237, G5238, G5239, G5240, G5241, G5242,
    G5243, G5244, G5245, G5246, G5247, G5248, G5249, G5250, G5251, G5252,
    G5253, G5254, G5255, G5256, G5257, G5258, G5259, G5260, G5261, G5262,
    G5263, G5264, G5265, G5266, G5267, G5268, G5269, G5270, G5271, G5272,
    G5273, G5274, G5275, G5276, G5277, G5278, G5279, G5280, G5281, G5282,
    G5283, G5284, G5285, G5286, G5287, G5288, G5289, G5290, G5291, G5292,
    G5293, G5294, G5295, G5296, G5297, G5298, G5299, G5300, G5301, G5302,
    G5303, G5304, G5305, G5306, G5307, G5308, G5309, G5310, G5311, G5312,
    G5313, G5314, G5315  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70,
    G71, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98,
    G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G110,
    G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G133, G134,
    G135, G136, G137, G138, G139, G140, G141, G142, G143, G144, G145, G146,
    G147, G148, G149, G150, G151, G152, G153, G154, G155, G156, G157, G158,
    G159, G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G170,
    G171, G172, G173, G174, G175, G176, G177, G178;
  output G5193, G5194, G5195, G5196, G5197, G5198, G5199, G5200, G5201, G5202,
    G5203, G5204, G5205, G5206, G5207, G5208, G5209, G5210, G5211, G5212,
    G5213, G5214, G5215, G5216, G5217, G5218, G5219, G5220, G5221, G5222,
    G5223, G5224, G5225, G5226, G5227, G5228, G5229, G5230, G5231, G5232,
    G5233, G5234, G5235, G5236, G5237, G5238, G5239, G5240, G5241, G5242,
    G5243, G5244, G5245, G5246, G5247, G5248, G5249, G5250, G5251, G5252,
    G5253, G5254, G5255, G5256, G5257, G5258, G5259, G5260, G5261, G5262,
    G5263, G5264, G5265, G5266, G5267, G5268, G5269, G5270, G5271, G5272,
    G5273, G5274, G5275, G5276, G5277, G5278, G5279, G5280, G5281, G5282,
    G5283, G5284, G5285, G5286, G5287, G5288, G5289, G5290, G5291, G5292,
    G5293, G5294, G5295, G5296, G5297, G5298, G5299, G5300, G5301, G5302,
    G5303, G5304, G5305, G5306, G5307, G5308, G5309, G5310, G5311, G5312,
    G5313, G5314, G5315;
  reg n2610_lo, n2613_lo, n2616_lo, n2619_lo, n2622_lo, n2625_lo, n2628_lo,
    n2634_lo, n2637_lo, n2640_lo, n2643_lo, n2646_lo, n2649_lo, n2652_lo,
    n2655_lo, n2658_lo, n2661_lo, n2664_lo, n2667_lo, n2670_lo, n2673_lo,
    n2676_lo, n2679_lo, n2682_lo, n2685_lo, n2688_lo, n2691_lo, n2694_lo,
    n2697_lo, n2700_lo, n2703_lo, n2706_lo, n2709_lo, n2712_lo, n2715_lo,
    n2718_lo, n2721_lo, n2724_lo, n2727_lo, n2730_lo, n2733_lo, n2736_lo,
    n2739_lo, n2742_lo, n2745_lo, n2748_lo, n2751_lo, n2754_lo, n2757_lo,
    n2760_lo, n2763_lo, n2766_lo, n2769_lo, n2772_lo, n2775_lo, n2778_lo,
    n2781_lo, n2784_lo, n2787_lo, n2790_lo, n2793_lo, n2796_lo, n2799_lo,
    n2802_lo, n2805_lo, n2808_lo, n2811_lo, n2814_lo, n2817_lo, n2820_lo,
    n2823_lo, n2826_lo, n2829_lo, n2832_lo, n2838_lo, n2841_lo, n2844_lo,
    n2847_lo, n2850_lo, n2853_lo, n2856_lo, n2862_lo, n2865_lo, n2868_lo,
    n2871_lo, n2874_lo, n2877_lo, n2880_lo, n2883_lo, n2886_lo, n2889_lo,
    n2892_lo, n2895_lo, n2898_lo, n2901_lo, n2904_lo, n2907_lo, n2910_lo,
    n2913_lo, n2916_lo, n2919_lo, n2922_lo, n2925_lo, n2928_lo, n2931_lo,
    n2934_lo, n2937_lo, n2940_lo, n2943_lo, n2946_lo, n2949_lo, n2952_lo,
    n2955_lo, n2958_lo, n2961_lo, n2964_lo, n2967_lo, n2970_lo, n2973_lo,
    n2976_lo, n2979_lo, n2982_lo, n2985_lo, n2988_lo, n2991_lo, n2994_lo,
    n2997_lo, n3000_lo, n3003_lo, n3006_lo, n3009_lo, n3012_lo, n3015_lo,
    n3018_lo, n3021_lo, n3024_lo, n3027_lo, n3030_lo, n3033_lo, n3036_lo,
    n3039_lo, n3042_lo, n3045_lo, n3048_lo, n3051_lo, n3054_lo, n3057_lo,
    n3060_lo, n3063_lo, n3066_lo, n3069_lo, n3072_lo, n3075_lo, n3078_lo,
    n3081_lo, n3084_lo, n3087_lo, n3090_lo, n3093_lo, n3096_lo, n3099_lo,
    n3102_lo, n3105_lo, n3108_lo, n3111_lo, n3114_lo, n3117_lo, n3120_lo,
    n3126_lo, n3129_lo, n3132_lo, n3138_lo, n3141_lo, n3144_lo, n3147_lo,
    n3150_lo, n3153_lo, n3156_lo, n3162_lo, n3165_lo, n3168_lo, n3174_lo,
    n3177_lo, n3180_lo, n3186_lo, n3189_lo, n3192_lo, n3195_lo, n3198_lo,
    n3201_lo, n3204_lo, n3210_lo, n3213_lo, n3216_lo, n3219_lo, n3222_lo,
    n3225_lo, n3228_lo, n3234_lo, n3237_lo, n3240_lo, n3243_lo, n3246_lo,
    n3249_lo, n3252_lo, n3255_lo, n3258_lo, n3261_lo, n3264_lo, n3267_lo,
    n3270_lo, n3273_lo, n3276_lo, n3279_lo, n3282_lo, n3285_lo, n3288_lo,
    n3294_lo, n3297_lo, n3300_lo, n3306_lo, n3309_lo, n3312_lo, n3318_lo,
    n3321_lo, n3324_lo, n3330_lo, n3333_lo, n3336_lo, n3339_lo, n3342_lo,
    n3345_lo, n3348_lo, n3351_lo, n3354_lo, n3357_lo, n3360_lo, n3363_lo,
    n3366_lo, n3369_lo, n3372_lo, n3375_lo, n3378_lo, n3381_lo, n3384_lo,
    n3387_lo, n3390_lo, n3393_lo, n3396_lo, n3399_lo, n3402_lo, n3405_lo,
    n3408_lo, n3411_lo, n3414_lo, n3417_lo, n3420_lo, n3423_lo, n3426_lo,
    n3429_lo, n3432_lo, n3435_lo, n3438_lo, n3441_lo, n3444_lo, n3447_lo,
    n3450_lo, n3453_lo, n3456_lo, n3459_lo, n3462_lo, n3465_lo, n3468_lo,
    n3471_lo, n3474_lo, n3477_lo, n3480_lo, n3483_lo, n3486_lo, n3489_lo,
    n3492_lo, n3495_lo, n3498_lo, n3501_lo, n3504_lo, n3507_lo, n3510_lo,
    n3513_lo, n3516_lo, n3519_lo, n3522_lo, n3525_lo, n3528_lo, n3531_lo,
    n3534_lo, n3537_lo, n3540_lo, n3543_lo, n3546_lo, n3549_lo, n3552_lo,
    n3555_lo, n3558_lo, n3561_lo, n3564_lo, n3567_lo, n3570_lo, n3573_lo,
    n3576_lo, n3579_lo, n3582_lo, n3585_lo, n3588_lo, n3591_lo, n3594_lo,
    n3597_lo, n3600_lo, n3603_lo, n3606_lo, n3609_lo, n3612_lo, n3615_lo,
    n3618_lo, n3621_lo, n3624_lo, n3627_lo, n3630_lo, n3633_lo, n3636_lo,
    n3639_lo, n3642_lo, n3645_lo, n3648_lo, n3651_lo, n3654_lo, n3666_lo,
    n3750_lo, n3762_lo, n3774_lo, n3786_lo, n3789_lo, n3792_lo, n3795_lo,
    n3798_lo, n3810_lo, n3822_lo, n3834_lo, n3846_lo, n3930_lo, n3933_lo,
    n3936_lo, n3942_lo, n3945_lo, n3948_lo, n3954_lo, n3957_lo, n3963_lo,
    n3966_lo, n3969_lo, n3975_lo, n3978_lo, n3990_lo, n4050_lo, n4062_lo,
    n4098_lo, n4107_lo, n4110_lo, n4122_lo, n4131_lo, n4155_lo, n4158_lo,
    n4170_lo, n4179_lo, n4182_lo, n4185_lo, n4188_lo, n4194_lo, n4197_lo,
    n4200_lo, n4206_lo, n4209_lo, n4212_lo, n4215_lo, n4230_lo, n4233_lo,
    n4236_lo, n4239_lo, n4242_lo, n4254_lo, n4290_lo, n4293_lo, n4302_lo,
    n4314_lo, n4350_lo, n4362_lo, n4374_lo, n4386_lo, n4398_lo, n4410_lo,
    n4413_lo, n4416_lo, n4419_lo, n4422_lo, n4425_lo, n4428_lo, n4431_lo,
    n4434_lo, n4437_lo, n4440_lo, n4443_lo, n4446_lo, n4449_lo, n4452_lo,
    n4455_lo, n4458_lo, n4461_lo, n4464_lo, n4467_lo, n4470_lo, n4473_lo,
    n4476_lo, n4479_lo, n4482_lo, n4485_lo, n4488_lo, n4494_lo, n4497_lo,
    n4500_lo, n4503_lo, n4506_lo, n4509_lo, n4512_lo, n4515_lo, n4518_lo,
    n4521_lo, n4524_lo, n4527_lo, n4530_lo, n4533_lo, n4536_lo, n4539_lo,
    n4542_lo, n4545_lo, n4554_lo, n4557_lo, n4560_lo, n4563_lo, n4566_lo,
    n4569_lo, n4572_lo, n4575_lo, n4578_lo, n4581_lo, n4584_lo, n4587_lo,
    n4590_lo, n4593_lo, n4596_lo, n4602_lo, n4605_lo, n4608_lo, n4614_lo,
    n4617_lo, n4620_lo, n4626_lo, n4629_lo, n4632_lo, n4638_lo, n4641_lo,
    n4644_lo, n4647_lo, n4650_lo, n4653_lo, n4656_lo, n4659_lo, n4662_lo,
    n4665_lo, n4668_lo, n4671_lo, n4674_lo, n4677_lo, n4680_lo, n4683_lo,
    n4686_lo, n4689_lo, n4692_lo, n4695_lo, n4698_lo, n4701_lo, n4704_lo,
    n4707_lo, n4710_lo, n4713_lo, n4716_lo, n4719_lo, n4722_lo, n4725_lo,
    n4728_lo, n4731_lo, n4734_lo, n4737_lo, n4740_lo, n4743_lo, n4970_o2,
    n4972_o2, n4989_o2, n5024_o2, n5025_o2, n5029_o2, n5042_o2, n5048_o2,
    n5093_o2, n5096_o2, n5193_o2, n5199_o2, n5203_o2, n5214_o2, n5221_o2,
    n5222_o2, n5273_o2, n5365_o2, n5385_o2, n5553_o2, n5636_o2, n5782_o2,
    n5778_o2, n5323_o2, n5325_o2, n5327_o2, n5329_o2, n5816_o2, n5817_o2,
    n5837_o2, n5844_o2, n5859_o2, n5857_o2, n5369_o2, n5371_o2, n5373_o2,
    n5400_o2, n5402_o2, n5404_o2, n5406_o2, n5407_o2, n5408_o2, n2722_o2,
    n1942_inv, n5412_o2, n1948_inv, n5557_o2, n5558_o2, n5559_o2, n5564_o2,
    n5565_o2, n1966_inv, n5568_o2, n5598_o2, n5600_o2, n5601_o2, n5602_o2,
    n5603_o2, n2853_o2, n5637_o2, n1993_inv, n1996_inv, n5635_o2, n5640_o2,
    n5641_o2, n5642_o2, n5650_o2, n5652_o2, n5653_o2, n5654_o2, n5655_o2,
    n5657_o2, n2029_inv, n5661_o2, n5656_o2, n5663_o2, n2041_inv, n5795_o2,
    n5796_o2, n5797_o2, n5739_o2, n5773_o2, n2059_inv, n5799_o2, n5802_o2,
    n2068_inv, n5831_o2, n5833_o2, n5820_o2, n5823_o2, n5824_o2, n5869_o2,
    n5848_o2, n5849_o2, n5856_o2, n5896_o2, n2754_o2, n2908_o2, n5892_o2,
    n5915_o2, n5919_o2, n5918_o2, n5920_o2, n5917_o2, lo586_buf_o2,
    n2818_o2, n2863_o2, n2134_inv, n2725_o2, n3016_o2, n3013_o2, n2655_o2,
    n2149_inv, lo562_buf_o2, n2155_inv, n2531_o2, n2700_o2, n5908_o2,
    n5910_o2, n5912_o2, n5914_o2, n2753_o2, n2878_o2, n2182_inv, n5934_o2,
    n5936_o2, n5938_o2, n2728_o2, lo358_buf_o2, lo418_buf_o2, lo474_buf_o2,
    lo554_buf_o2, lo558_buf_o2, lo574_buf_o2, n2215_inv, n2218_inv,
    n2221_inv, lo450_buf_o2, n2910_o2, n2683_o2, n2828_o2, n2582_o2,
    n2600_o2, n2542_o2, n2703_o2, lo510_buf_o2, lo514_buf_o2, lo538_buf_o2,
    lo578_buf_o2, n2260_inv, n2666_o2, n2667_o2, n2660_o2, n2272_inv,
    lo454_buf_o2, n3593_o2, n3048_o2, lo410_buf_o2, lo502_buf_o2,
    lo506_buf_o2, lo550_buf_o2, lo570_buf_o2, lo582_buf_o2, n2302_inv,
    n2305_inv, n3499_o2, n2311_inv, n2870_o2, n2317_inv, n2689_o2,
    n2323_inv, n2662_o2, lo350_buf_o2, lo498_buf_o2, lo518_buf_o2,
    lo522_buf_o2, lo598_buf_o2, n2344_inv, n2347_inv, n2350_inv, n2353_inv,
    n2356_inv, n2359_inv, n2872_o2, n3313_o2, n3273_o2, n2848_o2, n2893_o2,
    n3267_o2, n2925_o2, n2839_o2, n2831_o2, n2558_o2, n2562_o2, n2825_o2,
    n3263_o2, n3517_o2, n2873_o2, n2926_o2, n3261_o2, n3268_o2, n3274_o2,
    n3314_o2, n3571_o2, n2950_o2, n2951_o2, n3022_o2, n3023_o2, n3057_o2,
    n3058_o2, n2931_o2, n2911_o2, n2959_o2, n2960_o2, n2922_o2, n2888_o2,
    n2889_o2, n3051_o2, n3052_o2, n3063_o2, n2845_o2, n2476_inv, n3281_o2,
    n3294_o2, n2885_o2, n2786_o2, n2783_o2, n2801_o2, n2572_o2, n2628_o2,
    n2609_o2, n2618_o2, n2637_o2, n2525_o2, n2551_o2, n3759_o2, n2994_o2,
    n3040_o2, n2943_o2, n2991_o2, n3034_o2, n2881_o2, n3021_o2, n3062_o2,
    n2763_o2, n2764_o2, n2775_o2, n2776_o2, n2968_o2, n2969_o2, n2798_o2,
    n3661_o2, n2694_o2, n2572_inv, n2817_o2, n2514_o2, n2501_o2, n2584_inv,
    n2505_o2, n2492_o2, lo546_buf_o2, lo590_buf_o2, lo594_buf_o2,
    n2602_inv, n2605_inv, n2709_o2, n2611_inv, n2614_inv, n2617_inv,
    n2620_inv, n3590_o2, n3591_o2, n2629_inv, n3638_o2, n3639_o2,
    n2638_inv, n2641_inv, lo458_buf_o2, lo482_buf_o2, lo566_buf_o2,
    n2718_o2, n3707_o2, n3671_o2, n3680_o2, n3749_o2, n3716_o2, n3692_o2,
    n2591_o2, n3478_o2, n3610_o2, n3611_o2, n2686_inv, n2689_inv, n2738_o2,
    n3616_o2, n3617_o2, n3031_o2, n2704_inv, n3562_o2, n2502_o2, n3560_o2,
    n3554_o2, n3555_o2, n3536_o2, n3537_o2, n3508_o2, n3650_o2, n3740_o2,
    n3484_o2, n2740_inv, n2734_o2, n2735_o2, n2711_o2, lo585_buf_o2,
    n2719_o2, n2720_o2, n2723_o2, n2724_o2, n3624_o2, n3625_o2, n3015_o2,
    n3491_o2, n2779_inv, n2811_o2, n3010_o2, n3012_o2, lo382_buf_o2,
    lo386_buf_o2, lo390_buf_o2, lo398_buf_o2, lo402_buf_o2, lo406_buf_o2,
    n3492_o2, lo366_buf_o2, lo374_buf_o2, lo426_buf_o2, lo494_buf_o2,
    n2653_o2, n2654_o2, n2715_o2, n2740_o2, n2682_o2, n2736_o2,
    lo508_buf_o2, lo512_buf_o2, lo536_buf_o2, lo576_buf_o2, lo357_buf_o2,
    lo361_buf_o2, lo417_buf_o2, lo421_buf_o2, lo473_buf_o2, lo477_buf_o2,
    lo553_buf_o2, lo557_buf_o2, lo573_buf_o2, lo434_buf_o2, lo438_buf_o2,
    lo466_buf_o2, lo470_buf_o2, lo490_buf_o2, n2657_o2, n2658_o2, n2663_o2,
    n2664_o2, n2684_o2, n2685_o2;
  wire new_n2042_, new_n2044_, new_n2046_, new_n2048_, new_n2050_,
    new_n2052_, new_n2054_, new_n2056_, new_n2058_, new_n2060_, new_n2062_,
    new_n2064_, new_n2066_, new_n2068_, new_n2070_, new_n2072_, new_n2074_,
    new_n2076_, new_n2078_, new_n2080_, new_n2082_, new_n2084_, new_n2086_,
    new_n2088_, new_n2090_, new_n2092_, new_n2094_, new_n2096_, new_n2098_,
    new_n2100_, new_n2102_, new_n2104_, new_n2106_, new_n2108_, new_n2110_,
    new_n2112_, new_n2114_, new_n2116_, new_n2118_, new_n2120_, new_n2122_,
    new_n2124_, new_n2126_, new_n2128_, new_n2130_, new_n2132_, new_n2134_,
    new_n2136_, new_n2138_, new_n2140_, new_n2142_, new_n2144_, new_n2146_,
    new_n2148_, new_n2150_, new_n2152_, new_n2154_, new_n2156_, new_n2158_,
    new_n2160_, new_n2162_, new_n2164_, new_n2166_, new_n2168_, new_n2170_,
    new_n2172_, new_n2174_, new_n2176_, new_n2178_, new_n2180_, new_n2182_,
    new_n2184_, new_n2186_, new_n2188_, new_n2190_, new_n2192_, new_n2194_,
    new_n2196_, new_n2198_, new_n2200_, new_n2202_, new_n2204_, new_n2206_,
    new_n2208_, new_n2210_, new_n2212_, new_n2214_, new_n2216_, new_n2218_,
    new_n2220_, new_n2222_, new_n2224_, new_n2226_, new_n2228_, new_n2230_,
    new_n2232_, new_n2234_, new_n2236_, new_n2238_, new_n2240_, new_n2242_,
    new_n2244_, new_n2246_, new_n2248_, new_n2250_, new_n2252_, new_n2254_,
    new_n2256_, new_n2258_, new_n2260_, new_n2262_, new_n2264_, new_n2266_,
    new_n2268_, new_n2270_, new_n2272_, new_n2274_, new_n2276_, new_n2278_,
    new_n2280_, new_n2282_, new_n2284_, new_n2286_, new_n2288_, new_n2289_,
    new_n2290_, new_n2292_, new_n2294_, new_n2296_, new_n2298_, new_n2300_,
    new_n2302_, new_n2304_, new_n2306_, new_n2308_, new_n2310_, new_n2312_,
    new_n2314_, new_n2316_, new_n2318_, new_n2320_, new_n2322_, new_n2324_,
    new_n2326_, new_n2328_, new_n2330_, new_n2332_, new_n2334_, new_n2336_,
    new_n2338_, new_n2340_, new_n2342_, new_n2344_, new_n2346_, new_n2348_,
    new_n2350_, new_n2352_, new_n2354_, new_n2356_, new_n2358_, new_n2360_,
    new_n2362_, new_n2364_, new_n2366_, new_n2368_, new_n2370_, new_n2372_,
    new_n2374_, new_n2376_, new_n2378_, new_n2380_, new_n2382_, new_n2384_,
    new_n2386_, new_n2388_, new_n2390_, new_n2392_, new_n2394_, new_n2396_,
    new_n2398_, new_n2400_, new_n2402_, new_n2404_, new_n2405_, new_n2406_,
    new_n2408_, new_n2410_, new_n2411_, new_n2412_, new_n2414_, new_n2416_,
    new_n2418_, new_n2420_, new_n2422_, new_n2424_, new_n2427_, new_n2428_,
    new_n2430_, new_n2432_, new_n2434_, new_n2436_, new_n2438_, new_n2440_,
    new_n2442_, new_n2444_, new_n2446_, new_n2448_, new_n2450_, new_n2452_,
    new_n2454_, new_n2456_, new_n2458_, new_n2460_, new_n2462_, new_n2464_,
    new_n2466_, new_n2468_, new_n2470_, new_n2472_, new_n2474_, new_n2476_,
    new_n2478_, new_n2480_, new_n2483_, new_n2484_, new_n2486_, new_n2488_,
    new_n2491_, new_n2492_, new_n2494_, new_n2496_, new_n2499_, new_n2500_,
    new_n2502_, new_n2504_, new_n2506_, new_n2508_, new_n2510_, new_n2512_,
    new_n2514_, new_n2516_, new_n2518_, new_n2520_, new_n2522_, new_n2524_,
    new_n2526_, new_n2528_, new_n2530_, new_n2532_, new_n2534_, new_n2536_,
    new_n2538_, new_n2540_, new_n2542_, new_n2544_, new_n2546_, new_n2548_,
    new_n2550_, new_n2552_, new_n2554_, new_n2556_, new_n2558_, new_n2559_,
    new_n2560_, new_n2562_, new_n2564_, new_n2566_, new_n2568_, new_n2570_,
    new_n2572_, new_n2575_, new_n2576_, new_n2578_, new_n2580_, new_n2583_,
    new_n2584_, new_n2586_, new_n2588_, new_n2591_, new_n2592_, new_n2594_,
    new_n2596_, new_n2598_, new_n2600_, new_n2602_, new_n2604_, new_n2606_,
    new_n2608_, new_n2610_, new_n2612_, new_n2614_, new_n2616_, new_n2618_,
    new_n2620_, new_n2622_, new_n2624_, new_n2626_, new_n2628_, new_n2630_,
    new_n2632_, new_n2634_, new_n2636_, new_n2638_, new_n2640_, new_n2642_,
    new_n2644_, new_n2647_, new_n2648_, new_n2650_, new_n2652_, new_n2655_,
    new_n2656_, new_n2658_, new_n2660_, new_n2663_, new_n2664_, new_n2666_,
    new_n2668_, new_n2671_, new_n2672_, new_n2674_, new_n2676_, new_n2678_,
    new_n2680_, new_n2682_, new_n2684_, new_n2687_, new_n2688_, new_n2690_,
    new_n2692_, new_n2695_, new_n2696_, new_n2698_, new_n2700_, new_n2702_,
    new_n2704_, new_n2706_, new_n2708_, new_n2710_, new_n2712_, new_n2714_,
    new_n2716_, new_n2718_, new_n2720_, new_n2722_, new_n2724_, new_n2726_,
    new_n2728_, new_n2730_, new_n2732_, new_n2734_, new_n2736_, new_n2738_,
    new_n2740_, new_n2742_, new_n2744_, new_n2746_, new_n2748_, new_n2750_,
    new_n2752_, new_n2754_, new_n2756_, new_n2758_, new_n2760_, new_n2762_,
    new_n2764_, new_n2766_, new_n2768_, new_n2770_, new_n2772_, new_n2774_,
    new_n2776_, new_n2778_, new_n2780_, new_n2782_, new_n2784_, new_n2786_,
    new_n2788_, new_n2790_, new_n2792_, new_n2794_, new_n2796_, new_n2798_,
    new_n2800_, new_n2802_, new_n2804_, new_n2806_, new_n2808_, new_n2810_,
    new_n2812_, new_n2814_, new_n2817_, new_n2818_, new_n2820_, new_n2822_,
    new_n2824_, new_n2826_, new_n2828_, new_n2830_, new_n2832_, new_n2834_,
    new_n2836_, new_n2838_, new_n2840_, new_n2843_, new_n2844_, new_n2846_,
    new_n2848_, new_n2850_, new_n2852_, new_n2854_, new_n2856_, new_n2857_,
    new_n2858_, new_n2860_, new_n2862_, new_n2865_, new_n2866_, new_n2868_,
    new_n2870_, new_n2872_, new_n2874_, new_n2876_, new_n2878_, new_n2880_,
    new_n2881_, new_n2882_, new_n2884_, new_n2886_, new_n2889_, new_n2890_,
    new_n2892_, new_n2894_, new_n2896_, new_n2897_, new_n2898_, new_n2900_,
    new_n2902_, new_n2904_, new_n2906_, new_n2908_, new_n2910_, new_n2912_,
    new_n2914_, new_n2916_, new_n2918_, new_n2920_, new_n2922_, new_n2924_,
    new_n2926_, new_n2928_, new_n2930_, new_n2932_, new_n2934_, new_n2936_,
    new_n2938_, new_n2940_, new_n2942_, new_n2945_, new_n2946_, new_n2948_,
    new_n2950_, new_n2952_, new_n2954_, new_n2956_, new_n2958_, new_n2960_,
    new_n2962_, new_n2964_, new_n2966_, new_n2968_, new_n2970_, new_n2972_,
    new_n2974_, new_n2976_, new_n2978_, new_n2980_, new_n2982_, new_n2984_,
    new_n2986_, new_n2988_, new_n2990_, new_n2993_, new_n2994_, new_n2996_,
    new_n2998_, new_n3001_, new_n3002_, new_n3004_, new_n3006_, new_n3008_,
    new_n3010_, new_n3012_, new_n3014_, new_n3016_, new_n3018_, new_n3020_,
    new_n3022_, new_n3025_, new_n3026_, new_n3028_, new_n3030_, new_n3032_,
    new_n3034_, new_n3036_, new_n3038_, new_n3040_, new_n3042_, new_n3044_,
    new_n3046_, new_n3048_, new_n3050_, new_n3052_, new_n3054_, new_n3056_,
    new_n3058_, new_n3060_, new_n3062_, new_n3064_, new_n3066_, new_n3068_,
    new_n3070_, new_n3072_, new_n3074_, new_n3076_, new_n3078_, new_n3080_,
    new_n3083_, new_n3084_, new_n3086_, new_n3088_, new_n3090_, new_n3091_,
    new_n3092_, new_n3093_, new_n3094_, new_n3096_, new_n3098_, new_n3099_,
    new_n3100_, new_n3102_, new_n3104_, new_n3105_, new_n3106_, new_n3108_,
    new_n3109_, new_n3111_, new_n3112_, new_n3114_, new_n3116_, new_n3117_,
    new_n3118_, new_n3120_, new_n3122_, new_n3124_, new_n3126_, new_n3127_,
    new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3135_,
    new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3143_,
    new_n3144_, new_n3146_, new_n3148_, new_n3149_, new_n3150_, new_n3152_,
    new_n3154_, new_n3156_, new_n3158_, new_n3160_, new_n3162_, new_n3164_,
    new_n3166_, new_n3168_, new_n3171_, new_n3172_, new_n3173_, new_n3174_,
    new_n3175_, new_n3176_, new_n3178_, new_n3179_, new_n3180_, new_n3182_,
    new_n3183_, new_n3184_, new_n3186_, new_n3188_, new_n3189_, new_n3190_,
    new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3196_, new_n3198_,
    new_n3201_, new_n3202_, new_n3204_, new_n3206_, new_n3208_, new_n3209_,
    new_n3210_, new_n3212_, new_n3214_, new_n3217_, new_n3218_, new_n3220_,
    new_n3222_, new_n3225_, new_n3226_, new_n3228_, new_n3230_, new_n3233_,
    new_n3234_, new_n3236_, new_n3238_, new_n3241_, new_n3242_, new_n3244_,
    new_n3246_, new_n3247_, new_n3248_, new_n3250_, new_n3252_, new_n3254_,
    new_n3255_, new_n3256_, new_n3258_, new_n3260_, new_n3262_, new_n3263_,
    new_n3264_, new_n3266_, new_n3268_, new_n3270_, new_n3271_, new_n3272_,
    new_n3274_, new_n3276_, new_n3278_, new_n3279_, new_n3280_, new_n3282_,
    new_n3283_, new_n3284_, new_n3286_, new_n3288_, new_n3290_, new_n3291_,
    new_n3292_, new_n3294_, new_n3296_, new_n3298_, new_n3300_, new_n3302_,
    new_n3304_, new_n3307_, new_n3308_, new_n3310_, new_n3312_, new_n3314_,
    new_n3316_, new_n3318_, new_n3320_, new_n3322_, new_n3325_, new_n3326_,
    new_n3328_, new_n3331_, new_n3332_, new_n3334_, new_n3336_, new_n3338_,
    new_n3339_, new_n3340_, new_n3342_, new_n3344_, new_n3346_, new_n3347_,
    new_n3348_, new_n3350_, new_n3352_, new_n3354_, new_n3355_, new_n3356_,
    new_n3358_, new_n3360_, new_n3362_, new_n3363_, new_n3364_, new_n3366_,
    new_n3368_, new_n3370_, new_n3371_, new_n3372_, new_n3374_, new_n3376_,
    new_n3378_, new_n3379_, new_n3380_, new_n3382_, new_n3384_, new_n3385_,
    new_n3386_, new_n3387_, new_n3388_, new_n3390_, new_n3392_, new_n3393_,
    new_n3394_, new_n3395_, new_n3396_, new_n3398_, new_n3400_, new_n3403_,
    new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_,
    new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_,
    new_n3417_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_,
    new_n3425_, new_n3426_, new_n3429_, new_n3431_, new_n3433_, new_n3434_,
    new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3442_, new_n3443_,
    new_n3445_, new_n3446_, new_n3448_, new_n3449_, new_n3450_, new_n3451_,
    new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_,
    new_n3459_, new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3466_,
    new_n3468_, new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_,
    new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_,
    new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_,
    new_n3487_, new_n3489_, new_n3490_, new_n3492_, new_n3493_, new_n3494_,
    new_n3496_, new_n3497_, new_n3498_, new_n3500_, new_n3501_, new_n3502_,
    new_n3505_, new_n3506_, new_n3508_, new_n3509_, new_n3510_, new_n3511_,
    new_n3512_, new_n3513_, new_n3514_, new_n3516_, new_n3517_, new_n3518_,
    new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_,
    new_n3526_, new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_,
    new_n3533_, new_n3534_, new_n3536_, new_n3537_, new_n3538_, new_n3540_,
    new_n3541_, new_n3542_, new_n3544_, new_n3545_, new_n3546_, new_n3548_,
    new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_,
    new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_,
    new_n3564_, new_n3565_, new_n3566_, new_n3568_, new_n3570_, new_n3571_,
    new_n3572_, new_n3574_, new_n3576_, new_n3577_, new_n3578_, new_n3579_,
    new_n3580_, new_n3582_, new_n3583_, new_n3585_, new_n3586_, new_n3588_,
    new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3594_, new_n3595_,
    new_n3596_, new_n3598_, new_n3600_, new_n3602_, new_n3604_, new_n3606_,
    new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3612_, new_n3613_,
    new_n3614_, new_n3616_, new_n3618_, new_n3619_, new_n3620_, new_n3621_,
    new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_,
    new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3634_,
    new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_,
    new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_,
    new_n3648_, new_n3649_, new_n3650_, new_n3652_, new_n3653_, new_n3654_,
    new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3660_, new_n3661_,
    new_n3662_, new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_,
    new_n3668_, new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3674_,
    new_n3676_, new_n3678_, new_n3679_, new_n3680_, new_n3682_, new_n3683_,
    new_n3685_, new_n3686_, new_n3688_, new_n3690_, new_n3692_, new_n3694_,
    new_n3695_, new_n3696_, new_n3698_, new_n3699_, new_n3700_, new_n3701_,
    new_n3702_, new_n3704_, new_n3706_, new_n3708_, new_n3709_, new_n3710_,
    new_n3712_, new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_,
    new_n3719_, new_n3720_, new_n3721_, new_n3722_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3732_,
    new_n3734_, new_n3735_, new_n3736_, new_n3738_, new_n3740_, new_n3741_,
    new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_,
    new_n3748_, new_n3749_, new_n3750_, new_n3752_, new_n3753_, new_n3754_,
    new_n3756_, new_n3757_, new_n3758_, new_n3760_, new_n3762_, new_n3764_,
    new_n3765_, new_n3766_, new_n3768_, new_n3770_, new_n3772_, new_n3774_,
    new_n3776_, new_n3778_, new_n3780_, new_n3782_, new_n3785_, new_n3786_,
    new_n3788_, new_n3790_, new_n3792_, new_n3793_, new_n3794_, new_n3796_,
    new_n3798_, new_n3800_, new_n3803_, new_n3804_, new_n3806_, new_n3808_,
    new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_,
    new_n3818_, new_n3821_, new_n3822_, new_n3825_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3833_, new_n3834_,
    new_n3837_, new_n3838_, new_n3841_, new_n3843_, new_n3844_, new_n3846_,
    new_n3848_, new_n3850_, new_n3852_, new_n3854_, new_n3855_, new_n3856_,
    new_n3857_, new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_,
    new_n3863_, new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_,
    new_n3869_, new_n3870_, new_n3871_, new_n3872_, new_n3874_, new_n3876_,
    new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_, new_n3882_,
    new_n3883_, new_n3884_, new_n3885_, new_n3887_, new_n3889_, new_n3890_,
    new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_,
    new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_, new_n3903_,
    new_n3904_, new_n3905_, new_n3907_, new_n3908_, new_n3909_, new_n3910_,
    new_n3911_, new_n3912_, new_n3913_, new_n3915_, new_n3917_, new_n3918_,
    new_n3920_, new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_,
    new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3932_, new_n3934_,
    new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_,
    new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_,
    new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_,
    new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_,
    new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_,
    new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_,
    new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_,
    new_n3977_, new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_,
    new_n3983_, new_n3984_, new_n3985_, new_n3986_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3996_, new_n3998_, new_n3999_, new_n4000_, new_n4001_, new_n4002_,
    new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_, new_n4008_,
    new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_, new_n4014_,
    new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_, new_n4020_,
    new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_, new_n4026_,
    new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_, new_n4032_,
    new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_, new_n4038_,
    new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_,
    new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_,
    new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_, new_n4056_,
    new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_,
    new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_,
    new_n4069_, new_n4070_, new_n4072_, new_n4074_, new_n4076_, new_n4077_,
    new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_, new_n4083_,
    new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_, new_n4089_,
    new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_, new_n4095_,
    new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_, new_n4101_,
    new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_, new_n4108_,
    new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_,
    new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_,
    new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_,
    new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_,
    new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_,
    new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_,
    new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_,
    new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_,
    new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_,
    new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_,
    new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_,
    new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_,
    new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_,
    new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_,
    new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_,
    new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_,
    new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_,
    new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_,
    new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_,
    new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_,
    new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_,
    new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_,
    new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_,
    new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_,
    new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_,
    new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_,
    new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_,
    new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_,
    new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_,
    new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_,
    new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_,
    new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_,
    new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_,
    new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_,
    new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_,
    new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_,
    new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_,
    new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_,
    new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_,
    new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_,
    new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_,
    new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_,
    new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_,
    new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_,
    new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_,
    new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_,
    new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_,
    new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_,
    new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_,
    new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_,
    new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_,
    new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_,
    new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_,
    new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_,
    new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_,
    new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_,
    new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_,
    new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_,
    new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_,
    new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_,
    new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_,
    new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_,
    new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_,
    new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_,
    new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_,
    new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_,
    new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_,
    new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_,
    new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_,
    new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_,
    new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_,
    new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_,
    new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_,
    new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_,
    new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_,
    new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_,
    new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_,
    new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_,
    new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_,
    new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_,
    new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_,
    new_n4614_, new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_,
    new_n4620_, new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_,
    new_n4626_, new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_,
    new_n4632_, new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_,
    new_n4638_, new_n4639_, new_n4640_, new_n4641_, new_n4642_, new_n4643_,
    new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_,
    new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_,
    new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4661_,
    new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_,
    new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_, new_n4673_,
    new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_, new_n4679_,
    new_n4680_, new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_,
    new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_,
    new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_, new_n4697_,
    new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_, new_n4703_,
    new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_, new_n4709_,
    new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_, new_n4715_,
    new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_,
    new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_, new_n4727_,
    new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_, new_n4733_,
    new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_, new_n4739_,
    new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_,
    new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_,
    new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_,
    new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_,
    new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_,
    new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_,
    new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_,
    new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_,
    new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_,
    new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_,
    new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_,
    new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_,
    new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_,
    new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_,
    new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_,
    new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_,
    new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_,
    new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4847_,
    new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_,
    new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_,
    new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_,
    new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_,
    new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_,
    new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_,
    new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_,
    new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_,
    new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_,
    new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_,
    new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_,
    new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_,
    new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4925_,
    new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_,
    new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_,
    new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_,
    new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_,
    new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_,
    new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_,
    new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_,
    new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_,
    new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_,
    new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_,
    new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_,
    new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_,
    new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_,
    new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_,
    new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_,
    new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_,
    new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_,
    new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_,
    new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_,
    new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_,
    new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_,
    new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_,
    new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_,
    new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_,
    new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_,
    new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_,
    new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_,
    new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_,
    new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_,
    new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_,
    new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_,
    new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_,
    new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_,
    new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_,
    new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_,
    new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_,
    new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_,
    new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_,
    new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_,
    new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_,
    new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_,
    new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_,
    new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_,
    new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_,
    new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_,
    new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_,
    new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_,
    new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_,
    new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_,
    new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_,
    new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_,
    new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_,
    new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_,
    new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_,
    new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_,
    new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_,
    new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_,
    new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_,
    new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_,
    new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_,
    new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_,
    new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_,
    new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_,
    new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_,
    new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_,
    new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_,
    new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_,
    new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_,
    new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_,
    new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_,
    new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_,
    new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_,
    new_n5364_, new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_,
    new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_,
    new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_,
    new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_,
    new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_,
    new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_,
    new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_,
    new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_,
    new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_,
    new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_,
    new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_,
    new_n5430_, new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_,
    new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_,
    new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_,
    new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_,
    new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_,
    new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_,
    new_n5466_, new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_,
    new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_,
    new_n5478_, new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_,
    new_n5484_, new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_,
    new_n5490_, new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_,
    new_n5496_, new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_,
    new_n5502_, new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_,
    new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_,
    new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_,
    new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_,
    new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_,
    new_n5532_, new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_,
    new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_,
    new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_,
    new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_,
    new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_,
    new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_,
    new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_, new_n5573_,
    new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_, new_n5579_,
    new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_, new_n5585_,
    new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_, new_n5591_,
    new_n5592_, new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_,
    new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_,
    new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_,
    new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_, new_n5615_,
    new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_,
    new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_,
    new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_,
    new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_,
    new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_,
    new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_,
    new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_,
    new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_,
    new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_,
    new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_,
    new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_,
    new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_,
    new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_,
    new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_,
    new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_,
    new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_,
    new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_,
    new_n5718_, new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_,
    new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_,
    new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_,
    new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_,
    new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_,
    new_n6741_, new_n6742_, new_n6743_, new_n6744_, new_n6745_, new_n6746_,
    new_n6747_, new_n6748_, new_n6749_, new_n6750_, new_n6751_, new_n6752_,
    new_n6753_, new_n6754_, new_n6755_, new_n6756_, new_n6757_, new_n6758_,
    new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_, new_n6764_,
    new_n6765_, new_n6766_, new_n6767_, new_n6768_, new_n6769_, new_n6770_,
    new_n6771_, new_n6772_, new_n6773_, new_n6774_, new_n6775_, new_n6776_,
    new_n6777_, new_n6778_, new_n6779_, new_n6780_, new_n6781_, new_n6782_,
    new_n6783_, new_n6784_, new_n6785_, new_n6786_, new_n6787_, new_n6788_,
    new_n6789_, new_n6790_, new_n6791_, new_n6792_, new_n6793_, new_n6794_,
    new_n6795_, new_n6796_, new_n6797_, new_n6798_, new_n6799_, new_n6800_,
    new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_, new_n6806_,
    new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_, new_n6812_,
    new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_, new_n6818_,
    new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_, new_n6824_,
    new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_, new_n6830_,
    new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_, new_n6836_,
    new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_, new_n6842_,
    new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_, new_n6848_,
    new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_, new_n6854_,
    new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_, new_n6860_,
    new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_, new_n6866_,
    new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_, new_n6872_,
    new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_, new_n6878_,
    new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_, new_n6884_,
    new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_, new_n6890_,
    new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_, new_n6896_,
    new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_, new_n6902_,
    new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_, new_n6908_,
    new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_, new_n6914_,
    new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_, new_n6920_,
    new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_, new_n6926_,
    new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_, new_n6932_,
    new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_, new_n6938_,
    new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_, new_n6944_,
    new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_, new_n6950_,
    new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_, new_n6956_,
    new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_, new_n6962_,
    new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_, new_n6968_,
    new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_, new_n6974_,
    new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_, new_n6980_,
    new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_, new_n6986_,
    new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_, new_n6992_,
    new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_, new_n6998_,
    new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_, new_n7004_,
    new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_, new_n7010_,
    new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_, new_n7016_,
    new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_, new_n7022_,
    new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_, new_n7028_,
    new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_, new_n7034_,
    new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_, new_n7040_,
    new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_, new_n7046_,
    new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_, new_n7052_,
    new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_, new_n7058_,
    new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_, new_n7064_,
    new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_, new_n7070_,
    new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_, new_n7076_,
    new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_, new_n7082_,
    new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_, new_n7088_,
    new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_, new_n7094_,
    new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_, new_n7100_,
    new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_, new_n7106_,
    new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_, new_n7112_,
    new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_, new_n7118_,
    new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_, new_n7124_,
    new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_, new_n7130_,
    new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_, new_n7136_,
    new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_, new_n7142_,
    new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_, new_n7148_,
    new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_, new_n7154_,
    new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_, new_n7160_,
    new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_, new_n7166_,
    new_n7167_, new_n7168_, new_n7169_, new_n7170_, new_n7171_, new_n7172_,
    new_n7173_, new_n7174_, new_n7175_, new_n7176_, new_n7177_, new_n7178_,
    new_n7179_, new_n7180_, new_n7181_, new_n7182_, new_n7183_, new_n7184_,
    new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_, new_n7190_,
    new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_, new_n7196_,
    new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_, new_n7202_,
    new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7207_, new_n7208_,
    new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_, new_n7214_,
    new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_, new_n7220_,
    new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_, new_n7226_,
    new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_, new_n7232_,
    new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_, new_n7238_,
    new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_, new_n7244_,
    new_n7245_, new_n7246_, new_n7247_, new_n7248_, new_n7249_, new_n7250_,
    new_n7251_, new_n7252_, new_n7253_, new_n7254_, new_n7255_, new_n7256_,
    new_n7257_, new_n7258_, new_n7259_, new_n7260_, new_n7261_, new_n7262_,
    new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_, new_n7268_,
    new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_, new_n7274_,
    new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_, new_n7280_,
    new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_, new_n7286_,
    new_n7287_, new_n7288_, new_n7289_, new_n7290_, new_n7291_, new_n7292_,
    new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_, new_n7298_,
    new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_, new_n7304_,
    new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_, new_n7310_,
    new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_, new_n7316_,
    new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_, new_n7322_,
    new_n7323_, new_n7324_, new_n7325_, new_n7326_, new_n7327_, new_n7328_,
    new_n7329_, new_n7330_, new_n7331_, new_n7332_, new_n7333_, new_n7334_,
    new_n7335_, new_n7336_, new_n7337_, new_n7338_, new_n7339_, new_n7340_,
    new_n7341_, new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_,
    new_n7347_, new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_,
    new_n7353_, new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_,
    new_n7359_, new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_,
    new_n7365_, new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_,
    new_n7371_, new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_,
    new_n7377_, new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_,
    new_n7383_, new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_,
    new_n7389_, new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_,
    new_n7395_, new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_,
    new_n7401_, new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_,
    new_n7407_, new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_,
    new_n7413_, new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_,
    new_n7419_, new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_,
    new_n7425_, new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_,
    new_n7431_, new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_,
    new_n7437_, new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_,
    new_n7443_, new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_,
    new_n7449_, new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_,
    new_n7455_, new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_,
    new_n7461_, new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_,
    new_n7467_, new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_,
    new_n7473_, new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_,
    new_n7479_, new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_,
    new_n7485_, new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_,
    new_n7491_, new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_,
    new_n7497_, new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_,
    new_n7503_, new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_,
    new_n7509_, new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_,
    new_n7515_, new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_,
    new_n7521_, new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_,
    new_n7527_, new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_,
    new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_,
    new_n7539_, new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7544_,
    new_n7545_, new_n7546_, new_n7547_, new_n7548_, new_n7549_, new_n7550_,
    new_n7551_, new_n7552_, new_n7553_, new_n7554_, new_n7555_, new_n7556_,
    new_n7557_, new_n7558_, new_n7559_, new_n7560_, new_n7561_, new_n7562_,
    new_n7563_, new_n7564_, new_n7565_, new_n7566_, new_n7567_, new_n7568_,
    new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_, new_n7574_,
    new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_, new_n7580_,
    new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_, new_n7586_,
    new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_, new_n7592_,
    new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_, new_n7598_,
    new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_, new_n7604_,
    new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_, new_n7610_,
    new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_, new_n7616_,
    new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_, new_n7622_,
    new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_, new_n7628_,
    new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_, new_n7634_,
    new_n7635_, new_n7636_, new_n7637_, new_n7638_, new_n7639_, new_n7640_,
    new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_,
    new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_, new_n7652_,
    new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_, new_n7658_,
    new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_, new_n7664_,
    new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_, new_n7670_,
    new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_, new_n7676_,
    new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7681_, new_n7682_,
    new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_, new_n7688_,
    new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_, new_n7694_,
    new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_, new_n7700_,
    new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_, new_n7706_,
    new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_, new_n7712_,
    new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_, new_n7718_,
    new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_,
    new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7729_, new_n7730_,
    new_n7731_, new_n7732_, new_n7733_, new_n7734_, new_n7735_, new_n7736_,
    new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_,
    new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_,
    new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_,
    new_n7755_, new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_,
    new_n7761_, new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_,
    new_n7767_, new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_,
    new_n7773_, new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_,
    new_n7779_, new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_,
    new_n7785_, new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_,
    new_n7791_, new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_,
    new_n7797_, new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_,
    new_n7803_, new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_,
    new_n7809_, new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_,
    new_n7815_, new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_,
    new_n7821_, new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_,
    new_n7827_, new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_,
    new_n7833_, new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_,
    new_n7839_, new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_,
    new_n7845_, new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_,
    new_n7851_, new_n7852_, new_n7853_, new_n7854_, new_n7855_, new_n7856_,
    new_n7857_, new_n7858_, new_n7859_, new_n7860_, new_n7861_, new_n7862_,
    new_n7863_, new_n7864_, new_n7865_, new_n7866_, new_n7867_, new_n7868_,
    new_n7869_, new_n7870_, new_n7871_, new_n7872_, new_n7873_, new_n7874_,
    new_n7875_, new_n7876_, new_n7877_, new_n7878_, new_n7879_, new_n7880_,
    new_n7881_, new_n7882_, new_n7883_, new_n7884_, new_n7885_, new_n7886_,
    new_n7887_, new_n7888_, new_n7889_, new_n7890_, new_n7891_, new_n7892_,
    new_n7893_, new_n7894_, new_n7895_, new_n7896_, new_n7897_, new_n7898_,
    new_n7899_, new_n7900_, new_n7901_, new_n7902_, new_n7903_, new_n7904_,
    new_n7905_, new_n7906_, new_n7907_, new_n7908_, new_n7909_, new_n7910_,
    new_n7911_, new_n7912_, new_n7913_, new_n7914_, new_n7915_, new_n7916_,
    new_n7917_, new_n7918_, new_n7919_, new_n7920_, new_n7921_, new_n7922_,
    new_n7923_, new_n7924_, new_n7925_, new_n7926_, new_n7927_, new_n7928_,
    new_n7929_, new_n7930_, new_n7931_, new_n7932_, new_n7933_, new_n7934_,
    new_n7935_, new_n7936_, new_n7937_, new_n7938_, new_n7939_, new_n7940_,
    new_n7941_, new_n7942_, new_n7943_, new_n7944_, new_n7945_, new_n7946_,
    new_n7947_, new_n7948_, new_n7949_, new_n7950_, new_n7951_, new_n7952_,
    new_n7953_, new_n7954_, new_n7955_, new_n7956_, new_n7957_, new_n7958_,
    new_n7959_, new_n7960_, new_n7961_, new_n7962_, new_n7963_, new_n7964_,
    new_n7965_, new_n7966_, new_n7967_, new_n7968_, new_n7969_, new_n7970_,
    new_n7971_, new_n7972_, new_n7973_, new_n7974_, new_n7975_, new_n7976_,
    new_n7977_, new_n7978_, new_n7979_, new_n7980_, new_n7981_, new_n7982_,
    new_n7983_, new_n7984_, new_n7985_, new_n7986_, new_n7987_, new_n7988_,
    new_n7989_, new_n7990_, new_n7991_, new_n7992_, new_n7993_, new_n7994_,
    new_n7995_, new_n7996_, new_n7997_, new_n7998_, new_n7999_, new_n8000_,
    new_n8001_, new_n8002_, new_n8003_, new_n8004_, new_n8005_, new_n8006_,
    new_n8007_, new_n8008_, new_n8009_, new_n8010_, new_n8011_, new_n8012_,
    new_n8013_, new_n8014_, new_n8015_, new_n8016_, new_n8017_, new_n8018_,
    new_n8019_, new_n8020_, n7230_li000_li000, n7233_li001_li001,
    n7236_li002_li002, n7239_li003_li003, n7242_li004_li004,
    n7245_li005_li005, n7248_li006_li006, n7254_li008_li008,
    n7257_li009_li009, n7260_li010_li010, n7263_li011_li011,
    n7266_li012_li012, n7269_li013_li013, n7272_li014_li014,
    n7275_li015_li015, n7278_li016_li016, n7281_li017_li017,
    n7284_li018_li018, n7287_li019_li019, n7290_li020_li020,
    n7293_li021_li021, n7296_li022_li022, n7299_li023_li023,
    n7302_li024_li024, n7305_li025_li025, n7308_li026_li026,
    n7311_li027_li027, n7314_li028_li028, n7317_li029_li029,
    n7320_li030_li030, n7323_li031_li031, n7326_li032_li032,
    n7329_li033_li033, n7332_li034_li034, n7335_li035_li035,
    n7338_li036_li036, n7341_li037_li037, n7344_li038_li038,
    n7347_li039_li039, n7350_li040_li040, n7353_li041_li041,
    n7356_li042_li042, n7359_li043_li043, n7362_li044_li044,
    n7365_li045_li045, n7368_li046_li046, n7371_li047_li047,
    n7374_li048_li048, n7377_li049_li049, n7380_li050_li050,
    n7383_li051_li051, n7386_li052_li052, n7389_li053_li053,
    n7392_li054_li054, n7395_li055_li055, n7398_li056_li056,
    n7401_li057_li057, n7404_li058_li058, n7407_li059_li059,
    n7410_li060_li060, n7413_li061_li061, n7416_li062_li062,
    n7419_li063_li063, n7422_li064_li064, n7425_li065_li065,
    n7428_li066_li066, n7431_li067_li067, n7434_li068_li068,
    n7437_li069_li069, n7440_li070_li070, n7443_li071_li071,
    n7446_li072_li072, n7449_li073_li073, n7452_li074_li074,
    n7458_li076_li076, n7461_li077_li077, n7464_li078_li078,
    n7467_li079_li079, n7470_li080_li080, n7473_li081_li081,
    n7476_li082_li082, n7482_li084_li084, n7485_li085_li085,
    n7488_li086_li086, n7491_li087_li087, n7494_li088_li088,
    n7497_li089_li089, n7500_li090_li090, n7503_li091_li091,
    n7506_li092_li092, n7509_li093_li093, n7512_li094_li094,
    n7515_li095_li095, n7518_li096_li096, n7521_li097_li097,
    n7524_li098_li098, n7527_li099_li099, n7530_li100_li100,
    n7533_li101_li101, n7536_li102_li102, n7539_li103_li103,
    n7542_li104_li104, n7545_li105_li105, n7548_li106_li106,
    n7551_li107_li107, n7554_li108_li108, n7557_li109_li109,
    n7560_li110_li110, n7563_li111_li111, n7566_li112_li112,
    n7569_li113_li113, n7572_li114_li114, n7575_li115_li115,
    n7578_li116_li116, n7581_li117_li117, n7584_li118_li118,
    n7587_li119_li119, n7590_li120_li120, n7593_li121_li121,
    n7596_li122_li122, n7599_li123_li123, n7602_li124_li124,
    n7605_li125_li125, n7608_li126_li126, n7611_li127_li127,
    n7614_li128_li128, n7617_li129_li129, n7620_li130_li130,
    n7623_li131_li131, n7626_li132_li132, n7629_li133_li133,
    n7632_li134_li134, n7635_li135_li135, n7638_li136_li136,
    n7641_li137_li137, n7644_li138_li138, n7647_li139_li139,
    n7650_li140_li140, n7653_li141_li141, n7656_li142_li142,
    n7659_li143_li143, n7662_li144_li144, n7665_li145_li145,
    n7668_li146_li146, n7671_li147_li147, n7674_li148_li148,
    n7677_li149_li149, n7680_li150_li150, n7683_li151_li151,
    n7686_li152_li152, n7689_li153_li153, n7692_li154_li154,
    n7695_li155_li155, n7698_li156_li156, n7701_li157_li157,
    n7704_li158_li158, n7707_li159_li159, n7710_li160_li160,
    n7713_li161_li161, n7716_li162_li162, n7719_li163_li163,
    n7722_li164_li164, n7725_li165_li165, n7728_li166_li166,
    n7731_li167_li167, n7734_li168_li168, n7737_li169_li169,
    n7740_li170_li170, n7746_li172_li172, n7749_li173_li173,
    n7752_li174_li174, n7758_li176_li176, n7761_li177_li177,
    n7764_li178_li178, n7767_li179_li179, n7770_li180_li180,
    n7773_li181_li181, n7776_li182_li182, n7782_li184_li184,
    n7785_li185_li185, n7788_li186_li186, n7794_li188_li188,
    n7797_li189_li189, n7800_li190_li190, n7806_li192_li192,
    n7809_li193_li193, n7812_li194_li194, n7815_li195_li195,
    n7818_li196_li196, n7821_li197_li197, n7824_li198_li198,
    n7830_li200_li200, n7833_li201_li201, n7836_li202_li202,
    n7839_li203_li203, n7842_li204_li204, n7845_li205_li205,
    n7848_li206_li206, n7854_li208_li208, n7857_li209_li209,
    n7860_li210_li210, n7863_li211_li211, n7866_li212_li212,
    n7869_li213_li213, n7872_li214_li214, n7875_li215_li215,
    n7878_li216_li216, n7881_li217_li217, n7884_li218_li218,
    n7887_li219_li219, n7890_li220_li220, n7893_li221_li221,
    n7896_li222_li222, n7899_li223_li223, n7902_li224_li224,
    n7905_li225_li225, n7908_li226_li226, n7914_li228_li228,
    n7917_li229_li229, n7920_li230_li230, n7926_li232_li232,
    n7929_li233_li233, n7932_li234_li234, n7938_li236_li236,
    n7941_li237_li237, n7944_li238_li238, n7950_li240_li240,
    n7953_li241_li241, n7956_li242_li242, n7959_li243_li243,
    n7962_li244_li244, n7965_li245_li245, n7968_li246_li246,
    n7971_li247_li247, n7974_li248_li248, n7977_li249_li249,
    n7980_li250_li250, n7983_li251_li251, n7986_li252_li252,
    n7989_li253_li253, n7992_li254_li254, n7995_li255_li255,
    n7998_li256_li256, n8001_li257_li257, n8004_li258_li258,
    n8007_li259_li259, n8010_li260_li260, n8013_li261_li261,
    n8016_li262_li262, n8019_li263_li263, n8022_li264_li264,
    n8025_li265_li265, n8028_li266_li266, n8031_li267_li267,
    n8034_li268_li268, n8037_li269_li269, n8040_li270_li270,
    n8043_li271_li271, n8046_li272_li272, n8049_li273_li273,
    n8052_li274_li274, n8055_li275_li275, n8058_li276_li276,
    n8061_li277_li277, n8064_li278_li278, n8067_li279_li279,
    n8070_li280_li280, n8073_li281_li281, n8076_li282_li282,
    n8079_li283_li283, n8082_li284_li284, n8085_li285_li285,
    n8088_li286_li286, n8091_li287_li287, n8094_li288_li288,
    n8097_li289_li289, n8100_li290_li290, n8103_li291_li291,
    n8106_li292_li292, n8109_li293_li293, n8112_li294_li294,
    n8115_li295_li295, n8118_li296_li296, n8121_li297_li297,
    n8124_li298_li298, n8127_li299_li299, n8130_li300_li300,
    n8133_li301_li301, n8136_li302_li302, n8139_li303_li303,
    n8142_li304_li304, n8145_li305_li305, n8148_li306_li306,
    n8151_li307_li307, n8154_li308_li308, n8157_li309_li309,
    n8160_li310_li310, n8163_li311_li311, n8166_li312_li312,
    n8169_li313_li313, n8172_li314_li314, n8175_li315_li315,
    n8178_li316_li316, n8181_li317_li317, n8184_li318_li318,
    n8187_li319_li319, n8190_li320_li320, n8193_li321_li321,
    n8196_li322_li322, n8199_li323_li323, n8202_li324_li324,
    n8205_li325_li325, n8208_li326_li326, n8211_li327_li327,
    n8214_li328_li328, n8217_li329_li329, n8220_li330_li330,
    n8223_li331_li331, n8226_li332_li332, n8229_li333_li333,
    n8232_li334_li334, n8235_li335_li335, n8238_li336_li336,
    n8241_li337_li337, n8244_li338_li338, n8247_li339_li339,
    n8250_li340_li340, n8253_li341_li341, n8256_li342_li342,
    n8259_li343_li343, n8262_li344_li344, n8265_li345_li345,
    n8268_li346_li346, n8271_li347_li347, n8274_li348_li348,
    n8286_li352_li352, n8370_li380_li380, n8382_li384_li384,
    n8394_li388_li388, n8406_li392_li392, n8409_li393_li393,
    n8412_li394_li394, n8415_li395_li395, n8418_li396_li396,
    n8430_li400_li400, n8442_li404_li404, n8454_li408_li408,
    n8466_li412_li412, n8550_li440_li440, n8553_li441_li441,
    n8556_li442_li442, n8562_li444_li444, n8565_li445_li445,
    n8568_li446_li446, n8574_li448_li448, n8577_li449_li449,
    n8583_li451_li451, n8586_li452_li452, n8589_li453_li453,
    n8595_li455_li455, n8598_li456_li456, n8610_li460_li460,
    n8670_li480_li480, n8682_li484_li484, n8718_li496_li496,
    n8727_li499_li499, n8730_li500_li500, n8742_li504_li504,
    n8751_li507_li507, n8775_li515_li515, n8778_li516_li516,
    n8790_li520_li520, n8799_li523_li523, n8802_li524_li524,
    n8805_li525_li525, n8808_li526_li526, n8814_li528_li528,
    n8817_li529_li529, n8820_li530_li530, n8826_li532_li532,
    n8829_li533_li533, n8832_li534_li534, n8835_li535_li535,
    n8850_li540_li540, n8853_li541_li541, n8856_li542_li542,
    n8859_li543_li543, n8862_li544_li544, n8874_li548_li548,
    n8910_li560_li560, n8913_li561_li561, n8922_li564_li564,
    n8934_li568_li568, n8970_li580_li580, n8982_li584_li584,
    n8994_li588_li588, n9006_li592_li592, n9018_li596_li596,
    n9030_li600_li600, n9033_li601_li601, n9036_li602_li602,
    n9039_li603_li603, n9042_li604_li604, n9045_li605_li605,
    n9048_li606_li606, n9051_li607_li607, n9054_li608_li608,
    n9057_li609_li609, n9060_li610_li610, n9063_li611_li611,
    n9066_li612_li612, n9069_li613_li613, n9072_li614_li614,
    n9075_li615_li615, n9078_li616_li616, n9081_li617_li617,
    n9084_li618_li618, n9087_li619_li619, n9090_li620_li620,
    n9093_li621_li621, n9096_li622_li622, n9099_li623_li623,
    n9102_li624_li624, n9105_li625_li625, n9108_li626_li626,
    n9114_li628_li628, n9117_li629_li629, n9120_li630_li630,
    n9123_li631_li631, n9126_li632_li632, n9129_li633_li633,
    n9132_li634_li634, n9135_li635_li635, n9138_li636_li636,
    n9141_li637_li637, n9144_li638_li638, n9147_li639_li639,
    n9150_li640_li640, n9153_li641_li641, n9156_li642_li642,
    n9159_li643_li643, n9162_li644_li644, n9165_li645_li645,
    n9174_li648_li648, n9177_li649_li649, n9180_li650_li650,
    n9183_li651_li651, n9186_li652_li652, n9189_li653_li653,
    n9192_li654_li654, n9195_li655_li655, n9198_li656_li656,
    n9201_li657_li657, n9204_li658_li658, n9207_li659_li659,
    n9210_li660_li660, n9213_li661_li661, n9216_li662_li662,
    n9222_li664_li664, n9225_li665_li665, n9228_li666_li666,
    n9234_li668_li668, n9237_li669_li669, n9240_li670_li670,
    n9246_li672_li672, n9249_li673_li673, n9252_li674_li674,
    n9258_li676_li676, n9261_li677_li677, n9264_li678_li678,
    n9267_li679_li679, n9270_li680_li680, n9273_li681_li681,
    n9276_li682_li682, n9279_li683_li683, n9282_li684_li684,
    n9285_li685_li685, n9288_li686_li686, n9291_li687_li687,
    n9294_li688_li688, n9297_li689_li689, n9300_li690_li690,
    n9303_li691_li691, n9306_li692_li692, n9309_li693_li693,
    n9312_li694_li694, n9315_li695_li695, n9318_li696_li696,
    n9321_li697_li697, n9324_li698_li698, n9327_li699_li699,
    n9330_li700_li700, n9333_li701_li701, n9336_li702_li702,
    n9339_li703_li703, n9342_li704_li704, n9345_li705_li705,
    n9348_li706_li706, n9351_li707_li707, n9354_li708_li708,
    n9357_li709_li709, n9360_li710_li710, n9363_li711_li711, n4970_i2,
    n4972_i2, n4989_i2, n5024_i2, n5025_i2, n5029_i2, n5042_i2, n5048_i2,
    n5093_i2, n5096_i2, n5193_i2, n5199_i2, n5203_i2, n5214_i2, n5221_i2,
    n5222_i2, n5273_i2, n5365_i2, n5385_i2, n5553_i2, n5636_i2, n5782_i2,
    n5778_i2, n5323_i2, n5325_i2, n5327_i2, n5329_i2, n5816_i2, n5817_i2,
    n5837_i2, n5844_i2, n5859_i2, n5857_i2, n5369_i2, n5371_i2, n5373_i2,
    n5400_i2, n5402_i2, n5404_i2, n5406_i2, n5407_i2, n5408_i2, n2722_i2,
    n5411_i2, n5412_i2, n5413_i2, n5557_i2, n5558_i2, n5559_i2, n5564_i2,
    n5565_i2, n5561_i2, n5568_i2, n5598_i2, n5600_i2, n5601_i2, n5602_i2,
    n5603_i2, n2853_i2, n5637_i2, n5627_i2, n5628_i2, n5635_i2, n5640_i2,
    n5641_i2, n5642_i2, n5650_i2, n5652_i2, n5653_i2, n5654_i2, n5655_i2,
    n5657_i2, n5659_i2, n5661_i2, n5656_i2, n5663_i2, n5664_i2, n5795_i2,
    n5796_i2, n5797_i2, n5739_i2, n5773_i2, n5798_i2, n5799_i2, n5802_i2,
    n5803_i2, n5831_i2, n5833_i2, n5820_i2, n5823_i2, n5824_i2, n5869_i2,
    n5848_i2, n5849_i2, n5856_i2, n5896_i2, n2754_i2, n2908_i2, n5892_i2,
    n5915_i2, n5919_i2, n5918_i2, n5920_i2, n5917_i2, lo586_buf_i2,
    n2818_i2, n2863_i2, n2721_i2, n2725_i2, n3016_i2, n3013_i2, n2655_i2,
    n2741_i2, lo562_buf_i2, n2656_i2, n2531_i2, n2700_i2, n5908_i2,
    n5910_i2, n5912_i2, n5914_i2, n2753_i2, n2878_i2, n2836_i2, n5934_i2,
    n5936_i2, n5938_i2, n2728_i2, lo358_buf_i2, lo418_buf_i2, lo474_buf_i2,
    lo554_buf_i2, lo558_buf_i2, lo574_buf_i2, n2659_i2, n2665_i2, n2686_i2,
    lo450_buf_i2, n2910_i2, n2683_i2, n2828_i2, n2582_i2, n2600_i2,
    n2542_i2, n2703_i2, lo510_buf_i2, lo514_buf_i2, lo538_buf_i2,
    lo578_buf_i2, n2692_i2, n2666_i2, n2667_i2, n2660_i2, n2744_i2,
    lo454_buf_i2, n3593_i2, n3048_i2, lo410_buf_i2, lo502_buf_i2,
    lo506_buf_i2, lo550_buf_i2, lo570_buf_i2, lo582_buf_i2, n2646_i2,
    n2673_i2, n3499_i2, n2750_i2, n2870_i2, n2693_i2, n2689_i2, n2668_i2,
    n2662_i2, lo350_buf_i2, lo498_buf_i2, lo518_buf_i2, lo522_buf_i2,
    lo598_buf_i2, n2708_i2, n2674_i2, n2647_i2, n2751_i2, n2747_i2,
    n2669_i2, n2872_i2, n3313_i2, n3273_i2, n2848_i2, n2893_i2, n3267_i2,
    n2925_i2, n2839_i2, n2831_i2, n2558_i2, n2562_i2, n2825_i2, n3263_i2,
    n3517_i2, n2873_i2, n2926_i2, n3261_i2, n3268_i2, n3274_i2, n3314_i2,
    n3571_i2, n2950_i2, n2951_i2, n3022_i2, n3023_i2, n3057_i2, n3058_i2,
    n2931_i2, n2911_i2, n2959_i2, n2960_i2, n2922_i2, n2888_i2, n2889_i2,
    n3051_i2, n3052_i2, n3063_i2, n2845_i2, n2737_i2, n3281_i2, n3294_i2,
    n2885_i2, n2786_i2, n2783_i2, n2801_i2, n2572_i2, n2628_i2, n2609_i2,
    n2618_i2, n2637_i2, n2525_i2, n2551_i2, n3759_i2, n2994_i2, n3040_i2,
    n2943_i2, n2991_i2, n3034_i2, n2881_i2, n3021_i2, n3062_i2, n2763_i2,
    n2764_i2, n2775_i2, n2776_i2, n2968_i2, n2969_i2, n2798_i2, n3661_i2,
    n2694_i2, n2809_i2, n2817_i2, n2514_i2, n2501_i2, n2528_i2, n2505_i2,
    n2492_i2, lo546_buf_i2, lo590_buf_i2, lo594_buf_i2, n2679_i2, n2733_i2,
    n2709_i2, n2676_i2, n2649_i2, n2815_i2, n2704_i2, n3590_i2, n3591_i2,
    n2752_i2, n3638_i2, n3639_i2, n2695_i2, n3047_i2, lo458_buf_i2,
    lo482_buf_i2, lo566_buf_i2, n2718_i2, n3707_i2, n3671_i2, n3680_i2,
    n3749_i2, n3716_i2, n3692_i2, n2591_i2, n3478_i2, n3610_i2, n3611_i2,
    n2652_i2, n2714_i2, n2738_i2, n3616_i2, n3617_i2, n3031_i2, n2515_i2,
    n3562_i2, n2502_i2, n3560_i2, n3554_i2, n3555_i2, n3536_i2, n3537_i2,
    n3508_i2, n3650_i2, n3740_i2, n3484_i2, n2680_i2, n2734_i2, n2735_i2,
    n2711_i2, lo585_buf_i2, n2719_i2, n2720_i2, n2723_i2, n2724_i2,
    n3624_i2, n3625_i2, n3015_i2, n3491_i2, n2696_i2, n2811_i2, n3010_i2,
    n3012_i2, lo382_buf_i2, lo386_buf_i2, lo390_buf_i2, lo398_buf_i2,
    lo402_buf_i2, lo406_buf_i2, n3492_i2, lo366_buf_i2, lo374_buf_i2,
    lo426_buf_i2, lo494_buf_i2, n2653_i2, n2654_i2, n2715_i2, n2740_i2,
    n2682_i2, n2736_i2, lo508_buf_i2, lo512_buf_i2, lo536_buf_i2,
    lo576_buf_i2, lo357_buf_i2, lo361_buf_i2, lo417_buf_i2, lo421_buf_i2,
    lo473_buf_i2, lo477_buf_i2, lo553_buf_i2, lo557_buf_i2, lo573_buf_i2,
    lo434_buf_i2, lo438_buf_i2, lo466_buf_i2, lo470_buf_i2, lo490_buf_i2,
    n2657_i2, n2658_i2, n2663_i2, n2664_i2, n2684_i2, n2685_i2;
  assign new_n2042_ = G1;
  assign new_n2044_ = G2;
  assign new_n2046_ = G3;
  assign new_n2048_ = G4;
  assign new_n2050_ = G5;
  assign new_n2052_ = G6;
  assign new_n2054_ = G7;
  assign new_n2056_ = G8;
  assign new_n2058_ = G9;
  assign new_n2060_ = G10;
  assign new_n2062_ = G11;
  assign new_n2064_ = G12;
  assign new_n2066_ = G13;
  assign new_n2068_ = G14;
  assign new_n2070_ = G15;
  assign new_n2072_ = G16;
  assign new_n2074_ = G17;
  assign new_n2076_ = G18;
  assign new_n2078_ = G19;
  assign new_n2080_ = G20;
  assign new_n2082_ = G21;
  assign new_n2084_ = G22;
  assign new_n2086_ = G23;
  assign new_n2088_ = G24;
  assign new_n2090_ = G25;
  assign new_n2092_ = G26;
  assign new_n2094_ = G27;
  assign new_n2096_ = G28;
  assign new_n2098_ = G29;
  assign new_n2100_ = G30;
  assign new_n2102_ = G31;
  assign new_n2104_ = G32;
  assign new_n2106_ = G33;
  assign new_n2108_ = G34;
  assign new_n2110_ = G35;
  assign new_n2112_ = G36;
  assign new_n2114_ = G37;
  assign new_n2116_ = G38;
  assign new_n2118_ = G39;
  assign new_n2120_ = G40;
  assign new_n2122_ = G41;
  assign new_n2124_ = G42;
  assign new_n2126_ = G43;
  assign new_n2128_ = G44;
  assign new_n2130_ = G45;
  assign new_n2132_ = G46;
  assign new_n2134_ = G47;
  assign new_n2136_ = G48;
  assign new_n2138_ = G49;
  assign new_n2140_ = G50;
  assign new_n2142_ = G51;
  assign new_n2144_ = G52;
  assign new_n2146_ = G53;
  assign new_n2148_ = G54;
  assign new_n2150_ = G55;
  assign new_n2152_ = G56;
  assign new_n2154_ = G57;
  assign new_n2156_ = G58;
  assign new_n2158_ = G59;
  assign new_n2160_ = G60;
  assign new_n2162_ = G61;
  assign new_n2164_ = G62;
  assign new_n2166_ = G63;
  assign new_n2168_ = G64;
  assign new_n2170_ = G65;
  assign new_n2172_ = G66;
  assign new_n2174_ = G67;
  assign new_n2176_ = G68;
  assign new_n2178_ = G69;
  assign new_n2180_ = G70;
  assign new_n2182_ = G71;
  assign new_n2184_ = G72;
  assign new_n2186_ = G73;
  assign new_n2188_ = G74;
  assign new_n2190_ = G75;
  assign new_n2192_ = G76;
  assign new_n2194_ = G77;
  assign new_n2196_ = G78;
  assign new_n2198_ = G79;
  assign new_n2200_ = G80;
  assign new_n2202_ = G81;
  assign new_n2204_ = G82;
  assign new_n2206_ = G83;
  assign new_n2208_ = G84;
  assign new_n2210_ = G85;
  assign new_n2212_ = G86;
  assign new_n2214_ = G87;
  assign new_n2216_ = G88;
  assign new_n2218_ = G89;
  assign new_n2220_ = G90;
  assign new_n2222_ = G91;
  assign new_n2224_ = G92;
  assign new_n2226_ = G93;
  assign new_n2228_ = G94;
  assign new_n2230_ = G95;
  assign new_n2232_ = G96;
  assign new_n2234_ = G97;
  assign new_n2236_ = G98;
  assign new_n2238_ = G99;
  assign new_n2240_ = G100;
  assign new_n2242_ = G101;
  assign new_n2244_ = G102;
  assign new_n2246_ = G103;
  assign new_n2248_ = G104;
  assign new_n2250_ = G105;
  assign new_n2252_ = G106;
  assign new_n2254_ = G107;
  assign new_n2256_ = G108;
  assign new_n2258_ = G109;
  assign new_n2260_ = G110;
  assign new_n2262_ = G111;
  assign new_n2264_ = G112;
  assign new_n2266_ = G113;
  assign new_n2268_ = G114;
  assign new_n2270_ = G115;
  assign new_n2272_ = G116;
  assign new_n2274_ = G117;
  assign new_n2276_ = G118;
  assign new_n2278_ = G119;
  assign new_n2280_ = G120;
  assign new_n2282_ = G121;
  assign new_n2284_ = G122;
  assign new_n2286_ = G123;
  assign new_n2288_ = G124;
  assign new_n2289_ = ~G124;
  assign new_n2290_ = G125;
  assign new_n2292_ = G126;
  assign new_n2294_ = G127;
  assign new_n2296_ = G128;
  assign new_n2298_ = G129;
  assign new_n2300_ = G130;
  assign new_n2302_ = G131;
  assign new_n2304_ = G132;
  assign new_n2306_ = G133;
  assign new_n2308_ = G134;
  assign new_n2310_ = G135;
  assign new_n2312_ = G136;
  assign new_n2314_ = G137;
  assign new_n2316_ = G138;
  assign new_n2318_ = G139;
  assign new_n2320_ = G140;
  assign new_n2322_ = G141;
  assign new_n2324_ = G142;
  assign new_n2326_ = G143;
  assign new_n2328_ = G144;
  assign new_n2330_ = G145;
  assign new_n2332_ = G146;
  assign new_n2334_ = G147;
  assign new_n2336_ = G148;
  assign new_n2338_ = G149;
  assign new_n2340_ = G150;
  assign new_n2342_ = G151;
  assign new_n2344_ = G152;
  assign new_n2346_ = G153;
  assign new_n2348_ = G154;
  assign new_n2350_ = G155;
  assign new_n2352_ = G156;
  assign new_n2354_ = G157;
  assign new_n2356_ = G158;
  assign new_n2358_ = G159;
  assign new_n2360_ = G160;
  assign new_n2362_ = G161;
  assign new_n2364_ = G162;
  assign new_n2366_ = G163;
  assign new_n2368_ = G164;
  assign new_n2370_ = G165;
  assign new_n2372_ = G166;
  assign new_n2374_ = G167;
  assign new_n2376_ = G168;
  assign new_n2378_ = G169;
  assign new_n2380_ = G170;
  assign new_n2382_ = G171;
  assign new_n2384_ = G172;
  assign new_n2386_ = G173;
  assign new_n2388_ = G174;
  assign new_n2390_ = G175;
  assign new_n2392_ = G176;
  assign new_n2394_ = G177;
  assign new_n2396_ = G178;
  assign new_n2398_ = n2610_lo;
  assign new_n2400_ = n2613_lo;
  assign new_n2402_ = n2616_lo;
  assign new_n2404_ = n2619_lo;
  assign new_n2405_ = ~n2619_lo;
  assign new_n2406_ = n2622_lo;
  assign new_n2408_ = n2625_lo;
  assign new_n2410_ = n2628_lo;
  assign new_n2411_ = ~n2628_lo;
  assign new_n2412_ = n2634_lo;
  assign new_n2414_ = n2637_lo;
  assign new_n2416_ = n2640_lo;
  assign new_n2418_ = n2643_lo;
  assign new_n2420_ = n2646_lo;
  assign new_n2422_ = n2649_lo;
  assign new_n2424_ = n2652_lo;
  assign new_n2427_ = ~n2655_lo;
  assign new_n2428_ = n2658_lo;
  assign new_n2430_ = n2661_lo;
  assign new_n2432_ = n2664_lo;
  assign new_n2434_ = n2667_lo;
  assign new_n2436_ = n2670_lo;
  assign new_n2438_ = n2673_lo;
  assign new_n2440_ = n2676_lo;
  assign new_n2442_ = n2679_lo;
  assign new_n2444_ = n2682_lo;
  assign new_n2446_ = n2685_lo;
  assign new_n2448_ = n2688_lo;
  assign new_n2450_ = n2691_lo;
  assign new_n2452_ = n2694_lo;
  assign new_n2454_ = n2697_lo;
  assign new_n2456_ = n2700_lo;
  assign new_n2458_ = n2703_lo;
  assign new_n2460_ = n2706_lo;
  assign new_n2462_ = n2709_lo;
  assign new_n2464_ = n2712_lo;
  assign new_n2466_ = n2715_lo;
  assign new_n2468_ = n2718_lo;
  assign new_n2470_ = n2721_lo;
  assign new_n2472_ = n2724_lo;
  assign new_n2474_ = n2727_lo;
  assign new_n2476_ = n2730_lo;
  assign new_n2478_ = n2733_lo;
  assign new_n2480_ = n2736_lo;
  assign new_n2483_ = ~n2739_lo;
  assign new_n2484_ = n2742_lo;
  assign new_n2486_ = n2745_lo;
  assign new_n2488_ = n2748_lo;
  assign new_n2491_ = ~n2751_lo;
  assign new_n2492_ = n2754_lo;
  assign new_n2494_ = n2757_lo;
  assign new_n2496_ = n2760_lo;
  assign new_n2499_ = ~n2763_lo;
  assign new_n2500_ = n2766_lo;
  assign new_n2502_ = n2769_lo;
  assign new_n2504_ = n2772_lo;
  assign new_n2506_ = n2775_lo;
  assign new_n2508_ = n2778_lo;
  assign new_n2510_ = n2781_lo;
  assign new_n2512_ = n2784_lo;
  assign new_n2514_ = n2787_lo;
  assign new_n2516_ = n2790_lo;
  assign new_n2518_ = n2793_lo;
  assign new_n2520_ = n2796_lo;
  assign new_n2522_ = n2799_lo;
  assign new_n2524_ = n2802_lo;
  assign new_n2526_ = n2805_lo;
  assign new_n2528_ = n2808_lo;
  assign new_n2530_ = n2811_lo;
  assign new_n2532_ = n2814_lo;
  assign new_n2534_ = n2817_lo;
  assign new_n2536_ = n2820_lo;
  assign new_n2538_ = n2823_lo;
  assign new_n2540_ = n2826_lo;
  assign new_n2542_ = n2829_lo;
  assign new_n2544_ = n2832_lo;
  assign new_n2546_ = n2838_lo;
  assign new_n2548_ = n2841_lo;
  assign new_n2550_ = n2844_lo;
  assign new_n2552_ = n2847_lo;
  assign new_n2554_ = n2850_lo;
  assign new_n2556_ = n2853_lo;
  assign new_n2558_ = n2856_lo;
  assign new_n2559_ = ~n2856_lo;
  assign new_n2560_ = n2862_lo;
  assign new_n2562_ = n2865_lo;
  assign new_n2564_ = n2868_lo;
  assign new_n2566_ = n2871_lo;
  assign new_n2568_ = n2874_lo;
  assign new_n2570_ = n2877_lo;
  assign new_n2572_ = n2880_lo;
  assign new_n2575_ = ~n2883_lo;
  assign new_n2576_ = n2886_lo;
  assign new_n2578_ = n2889_lo;
  assign new_n2580_ = n2892_lo;
  assign new_n2583_ = ~n2895_lo;
  assign new_n2584_ = n2898_lo;
  assign new_n2586_ = n2901_lo;
  assign new_n2588_ = n2904_lo;
  assign new_n2591_ = ~n2907_lo;
  assign new_n2592_ = n2910_lo;
  assign new_n2594_ = n2913_lo;
  assign new_n2596_ = n2916_lo;
  assign new_n2598_ = n2919_lo;
  assign new_n2600_ = n2922_lo;
  assign new_n2602_ = n2925_lo;
  assign new_n2604_ = n2928_lo;
  assign new_n2606_ = n2931_lo;
  assign new_n2608_ = n2934_lo;
  assign new_n2610_ = n2937_lo;
  assign new_n2612_ = n2940_lo;
  assign new_n2614_ = n2943_lo;
  assign new_n2616_ = n2946_lo;
  assign new_n2618_ = n2949_lo;
  assign new_n2620_ = n2952_lo;
  assign new_n2622_ = n2955_lo;
  assign new_n2624_ = n2958_lo;
  assign new_n2626_ = n2961_lo;
  assign new_n2628_ = n2964_lo;
  assign new_n2630_ = n2967_lo;
  assign new_n2632_ = n2970_lo;
  assign new_n2634_ = n2973_lo;
  assign new_n2636_ = n2976_lo;
  assign new_n2638_ = n2979_lo;
  assign new_n2640_ = n2982_lo;
  assign new_n2642_ = n2985_lo;
  assign new_n2644_ = n2988_lo;
  assign new_n2647_ = ~n2991_lo;
  assign new_n2648_ = n2994_lo;
  assign new_n2650_ = n2997_lo;
  assign new_n2652_ = n3000_lo;
  assign new_n2655_ = ~n3003_lo;
  assign new_n2656_ = n3006_lo;
  assign new_n2658_ = n3009_lo;
  assign new_n2660_ = n3012_lo;
  assign new_n2663_ = ~n3015_lo;
  assign new_n2664_ = n3018_lo;
  assign new_n2666_ = n3021_lo;
  assign new_n2668_ = n3024_lo;
  assign new_n2671_ = ~n3027_lo;
  assign new_n2672_ = n3030_lo;
  assign new_n2674_ = n3033_lo;
  assign new_n2676_ = n3036_lo;
  assign new_n2678_ = n3039_lo;
  assign new_n2680_ = n3042_lo;
  assign new_n2682_ = n3045_lo;
  assign new_n2684_ = n3048_lo;
  assign new_n2687_ = ~n3051_lo;
  assign new_n2688_ = n3054_lo;
  assign new_n2690_ = n3057_lo;
  assign new_n2692_ = n3060_lo;
  assign new_n2695_ = ~n3063_lo;
  assign new_n2696_ = n3066_lo;
  assign new_n2698_ = n3069_lo;
  assign new_n2700_ = n3072_lo;
  assign new_n2702_ = n3075_lo;
  assign new_n2704_ = n3078_lo;
  assign new_n2706_ = n3081_lo;
  assign new_n2708_ = n3084_lo;
  assign new_n2710_ = n3087_lo;
  assign new_n2712_ = n3090_lo;
  assign new_n2714_ = n3093_lo;
  assign new_n2716_ = n3096_lo;
  assign new_n2718_ = n3099_lo;
  assign new_n2720_ = n3102_lo;
  assign new_n2722_ = n3105_lo;
  assign new_n2724_ = n3108_lo;
  assign new_n2726_ = n3111_lo;
  assign new_n2728_ = n3114_lo;
  assign new_n2730_ = n3117_lo;
  assign new_n2732_ = n3120_lo;
  assign new_n2734_ = n3126_lo;
  assign new_n2736_ = n3129_lo;
  assign new_n2738_ = n3132_lo;
  assign new_n2740_ = n3138_lo;
  assign new_n2742_ = n3141_lo;
  assign new_n2744_ = n3144_lo;
  assign new_n2746_ = n3147_lo;
  assign new_n2748_ = n3150_lo;
  assign new_n2750_ = n3153_lo;
  assign new_n2752_ = n3156_lo;
  assign new_n2754_ = n3162_lo;
  assign new_n2756_ = n3165_lo;
  assign new_n2758_ = n3168_lo;
  assign new_n2760_ = n3174_lo;
  assign new_n2762_ = n3177_lo;
  assign new_n2764_ = n3180_lo;
  assign new_n2766_ = n3186_lo;
  assign new_n2768_ = n3189_lo;
  assign new_n2770_ = n3192_lo;
  assign new_n2772_ = n3195_lo;
  assign new_n2774_ = n3198_lo;
  assign new_n2776_ = n3201_lo;
  assign new_n2778_ = n3204_lo;
  assign new_n2780_ = n3210_lo;
  assign new_n2782_ = n3213_lo;
  assign new_n2784_ = n3216_lo;
  assign new_n2786_ = n3219_lo;
  assign new_n2788_ = n3222_lo;
  assign new_n2790_ = n3225_lo;
  assign new_n2792_ = n3228_lo;
  assign new_n2794_ = n3234_lo;
  assign new_n2796_ = n3237_lo;
  assign new_n2798_ = n3240_lo;
  assign new_n2800_ = n3243_lo;
  assign new_n2802_ = n3246_lo;
  assign new_n2804_ = n3249_lo;
  assign new_n2806_ = n3252_lo;
  assign new_n2808_ = n3255_lo;
  assign new_n2810_ = n3258_lo;
  assign new_n2812_ = n3261_lo;
  assign new_n2814_ = n3264_lo;
  assign new_n2817_ = ~n3267_lo;
  assign new_n2818_ = n3270_lo;
  assign new_n2820_ = n3273_lo;
  assign new_n2822_ = n3276_lo;
  assign new_n2824_ = n3279_lo;
  assign new_n2826_ = n3282_lo;
  assign new_n2828_ = n3285_lo;
  assign new_n2830_ = n3288_lo;
  assign new_n2832_ = n3294_lo;
  assign new_n2834_ = n3297_lo;
  assign new_n2836_ = n3300_lo;
  assign new_n2838_ = n3306_lo;
  assign new_n2840_ = n3309_lo;
  assign new_n2843_ = ~n3312_lo;
  assign new_n2844_ = n3318_lo;
  assign new_n2846_ = n3321_lo;
  assign new_n2848_ = n3324_lo;
  assign new_n2850_ = n3330_lo;
  assign new_n2852_ = n3333_lo;
  assign new_n2854_ = n3336_lo;
  assign new_n2856_ = n3339_lo;
  assign new_n2857_ = ~n3339_lo;
  assign new_n2858_ = n3342_lo;
  assign new_n2860_ = n3345_lo;
  assign new_n2862_ = n3348_lo;
  assign new_n2865_ = ~n3351_lo;
  assign new_n2866_ = n3354_lo;
  assign new_n2868_ = n3357_lo;
  assign new_n2870_ = n3360_lo;
  assign new_n2872_ = n3363_lo;
  assign new_n2874_ = n3366_lo;
  assign new_n2876_ = n3369_lo;
  assign new_n2878_ = n3372_lo;
  assign new_n2880_ = n3375_lo;
  assign new_n2881_ = ~n3375_lo;
  assign new_n2882_ = n3378_lo;
  assign new_n2884_ = n3381_lo;
  assign new_n2886_ = n3384_lo;
  assign new_n2889_ = ~n3387_lo;
  assign new_n2890_ = n3390_lo;
  assign new_n2892_ = n3393_lo;
  assign new_n2894_ = n3396_lo;
  assign new_n2896_ = n3399_lo;
  assign new_n2897_ = ~n3399_lo;
  assign new_n2898_ = n3402_lo;
  assign new_n2900_ = n3405_lo;
  assign new_n2902_ = n3408_lo;
  assign new_n2904_ = n3411_lo;
  assign new_n2906_ = n3414_lo;
  assign new_n2908_ = n3417_lo;
  assign new_n2910_ = n3420_lo;
  assign new_n2912_ = n3423_lo;
  assign new_n2914_ = n3426_lo;
  assign new_n2916_ = n3429_lo;
  assign new_n2918_ = n3432_lo;
  assign new_n2920_ = n3435_lo;
  assign new_n2922_ = n3438_lo;
  assign new_n2924_ = n3441_lo;
  assign new_n2926_ = n3444_lo;
  assign new_n2928_ = n3447_lo;
  assign new_n2930_ = n3450_lo;
  assign new_n2932_ = n3453_lo;
  assign new_n2934_ = n3456_lo;
  assign new_n2936_ = n3459_lo;
  assign new_n2938_ = n3462_lo;
  assign new_n2940_ = n3465_lo;
  assign new_n2942_ = n3468_lo;
  assign new_n2945_ = ~n3471_lo;
  assign new_n2946_ = n3474_lo;
  assign new_n2948_ = n3477_lo;
  assign new_n2950_ = n3480_lo;
  assign new_n2952_ = n3483_lo;
  assign new_n2954_ = n3486_lo;
  assign new_n2956_ = n3489_lo;
  assign new_n2958_ = n3492_lo;
  assign new_n2960_ = n3495_lo;
  assign new_n2962_ = n3498_lo;
  assign new_n2964_ = n3501_lo;
  assign new_n2966_ = n3504_lo;
  assign new_n2968_ = n3507_lo;
  assign new_n2970_ = n3510_lo;
  assign new_n2972_ = n3513_lo;
  assign new_n2974_ = n3516_lo;
  assign new_n2976_ = n3519_lo;
  assign new_n2978_ = n3522_lo;
  assign new_n2980_ = n3525_lo;
  assign new_n2982_ = n3528_lo;
  assign new_n2984_ = n3531_lo;
  assign new_n2986_ = n3534_lo;
  assign new_n2988_ = n3537_lo;
  assign new_n2990_ = n3540_lo;
  assign new_n2993_ = ~n3543_lo;
  assign new_n2994_ = n3546_lo;
  assign new_n2996_ = n3549_lo;
  assign new_n2998_ = n3552_lo;
  assign new_n3001_ = ~n3555_lo;
  assign new_n3002_ = n3558_lo;
  assign new_n3004_ = n3561_lo;
  assign new_n3006_ = n3564_lo;
  assign new_n3008_ = n3567_lo;
  assign new_n3010_ = n3570_lo;
  assign new_n3012_ = n3573_lo;
  assign new_n3014_ = n3576_lo;
  assign new_n3016_ = n3579_lo;
  assign new_n3018_ = n3582_lo;
  assign new_n3020_ = n3585_lo;
  assign new_n3022_ = n3588_lo;
  assign new_n3025_ = ~n3591_lo;
  assign new_n3026_ = n3594_lo;
  assign new_n3028_ = n3597_lo;
  assign new_n3030_ = n3600_lo;
  assign new_n3032_ = n3603_lo;
  assign new_n3034_ = n3606_lo;
  assign new_n3036_ = n3609_lo;
  assign new_n3038_ = n3612_lo;
  assign new_n3040_ = n3615_lo;
  assign new_n3042_ = n3618_lo;
  assign new_n3044_ = n3621_lo;
  assign new_n3046_ = n3624_lo;
  assign new_n3048_ = n3627_lo;
  assign new_n3050_ = n3630_lo;
  assign new_n3052_ = n3633_lo;
  assign new_n3054_ = n3636_lo;
  assign new_n3056_ = n3639_lo;
  assign new_n3058_ = n3642_lo;
  assign new_n3060_ = n3645_lo;
  assign new_n3062_ = n3648_lo;
  assign new_n3064_ = n3651_lo;
  assign new_n3066_ = n3654_lo;
  assign new_n3068_ = n3666_lo;
  assign new_n3070_ = n3750_lo;
  assign new_n3072_ = n3762_lo;
  assign new_n3074_ = n3774_lo;
  assign new_n3076_ = n3786_lo;
  assign new_n3078_ = n3789_lo;
  assign new_n3080_ = n3792_lo;
  assign new_n3083_ = ~n3795_lo;
  assign new_n3084_ = n3798_lo;
  assign new_n3086_ = n3810_lo;
  assign new_n3088_ = n3822_lo;
  assign new_n3090_ = n3834_lo;
  assign new_n3091_ = ~n3834_lo;
  assign new_n3092_ = n3846_lo;
  assign new_n3093_ = ~n3846_lo;
  assign new_n3094_ = n3930_lo;
  assign new_n3096_ = n3933_lo;
  assign new_n3098_ = n3936_lo;
  assign new_n3099_ = ~n3936_lo;
  assign new_n3100_ = n3942_lo;
  assign new_n3102_ = n3945_lo;
  assign new_n3104_ = n3948_lo;
  assign new_n3105_ = ~n3948_lo;
  assign new_n3106_ = n3954_lo;
  assign new_n3108_ = n3957_lo;
  assign new_n3109_ = ~n3957_lo;
  assign new_n3111_ = ~n3963_lo;
  assign new_n3112_ = n3966_lo;
  assign new_n3114_ = n3969_lo;
  assign new_n3116_ = n3975_lo;
  assign new_n3117_ = ~n3975_lo;
  assign new_n3118_ = n3978_lo;
  assign new_n3120_ = n3990_lo;
  assign new_n3122_ = n4050_lo;
  assign new_n3124_ = n4062_lo;
  assign new_n3126_ = n4098_lo;
  assign new_n3127_ = ~n4098_lo;
  assign new_n3129_ = ~n4107_lo;
  assign new_n3130_ = n4110_lo;
  assign new_n3131_ = ~n4110_lo;
  assign new_n3132_ = n4122_lo;
  assign new_n3133_ = ~n4122_lo;
  assign new_n3135_ = ~n4131_lo;
  assign new_n3137_ = ~n4155_lo;
  assign new_n3138_ = n4158_lo;
  assign new_n3139_ = ~n4158_lo;
  assign new_n3140_ = n4170_lo;
  assign new_n3141_ = ~n4170_lo;
  assign new_n3143_ = ~n4179_lo;
  assign new_n3144_ = n4182_lo;
  assign new_n3146_ = n4185_lo;
  assign new_n3148_ = n4188_lo;
  assign new_n3149_ = ~n4188_lo;
  assign new_n3150_ = n4194_lo;
  assign new_n3152_ = n4197_lo;
  assign new_n3154_ = n4200_lo;
  assign new_n3156_ = n4206_lo;
  assign new_n3158_ = n4209_lo;
  assign new_n3160_ = n4212_lo;
  assign new_n3162_ = n4215_lo;
  assign new_n3164_ = n4230_lo;
  assign new_n3166_ = n4233_lo;
  assign new_n3168_ = n4236_lo;
  assign new_n3171_ = ~n4239_lo;
  assign new_n3172_ = n4242_lo;
  assign new_n3173_ = ~n4242_lo;
  assign new_n3174_ = n4254_lo;
  assign new_n3175_ = ~n4254_lo;
  assign new_n3176_ = n4290_lo;
  assign new_n3178_ = n4293_lo;
  assign new_n3179_ = ~n4293_lo;
  assign new_n3180_ = n4302_lo;
  assign new_n3182_ = n4314_lo;
  assign new_n3183_ = ~n4314_lo;
  assign new_n3184_ = n4350_lo;
  assign new_n3186_ = n4362_lo;
  assign new_n3188_ = n4374_lo;
  assign new_n3189_ = ~n4374_lo;
  assign new_n3190_ = n4386_lo;
  assign new_n3191_ = ~n4386_lo;
  assign new_n3192_ = n4398_lo;
  assign new_n3193_ = ~n4398_lo;
  assign new_n3194_ = n4410_lo;
  assign new_n3196_ = n4413_lo;
  assign new_n3198_ = n4416_lo;
  assign new_n3201_ = ~n4419_lo;
  assign new_n3202_ = n4422_lo;
  assign new_n3204_ = n4425_lo;
  assign new_n3206_ = n4428_lo;
  assign new_n3208_ = n4431_lo;
  assign new_n3209_ = ~n4431_lo;
  assign new_n3210_ = n4434_lo;
  assign new_n3212_ = n4437_lo;
  assign new_n3214_ = n4440_lo;
  assign new_n3217_ = ~n4443_lo;
  assign new_n3218_ = n4446_lo;
  assign new_n3220_ = n4449_lo;
  assign new_n3222_ = n4452_lo;
  assign new_n3225_ = ~n4455_lo;
  assign new_n3226_ = n4458_lo;
  assign new_n3228_ = n4461_lo;
  assign new_n3230_ = n4464_lo;
  assign new_n3233_ = ~n4467_lo;
  assign new_n3234_ = n4470_lo;
  assign new_n3236_ = n4473_lo;
  assign new_n3238_ = n4476_lo;
  assign new_n3241_ = ~n4479_lo;
  assign new_n3242_ = n4482_lo;
  assign new_n3244_ = n4485_lo;
  assign new_n3246_ = n4488_lo;
  assign new_n3247_ = ~n4488_lo;
  assign new_n3248_ = n4494_lo;
  assign new_n3250_ = n4497_lo;
  assign new_n3252_ = n4500_lo;
  assign new_n3254_ = n4503_lo;
  assign new_n3255_ = ~n4503_lo;
  assign new_n3256_ = n4506_lo;
  assign new_n3258_ = n4509_lo;
  assign new_n3260_ = n4512_lo;
  assign new_n3262_ = n4515_lo;
  assign new_n3263_ = ~n4515_lo;
  assign new_n3264_ = n4518_lo;
  assign new_n3266_ = n4521_lo;
  assign new_n3268_ = n4524_lo;
  assign new_n3270_ = n4527_lo;
  assign new_n3271_ = ~n4527_lo;
  assign new_n3272_ = n4530_lo;
  assign new_n3274_ = n4533_lo;
  assign new_n3276_ = n4536_lo;
  assign new_n3278_ = n4539_lo;
  assign new_n3279_ = ~n4539_lo;
  assign new_n3280_ = n4542_lo;
  assign new_n3282_ = n4545_lo;
  assign new_n3283_ = ~n4545_lo;
  assign new_n3284_ = n4554_lo;
  assign new_n3286_ = n4557_lo;
  assign new_n3288_ = n4560_lo;
  assign new_n3290_ = n4563_lo;
  assign new_n3291_ = ~n4563_lo;
  assign new_n3292_ = n4566_lo;
  assign new_n3294_ = n4569_lo;
  assign new_n3296_ = n4572_lo;
  assign new_n3298_ = n4575_lo;
  assign new_n3300_ = n4578_lo;
  assign new_n3302_ = n4581_lo;
  assign new_n3304_ = n4584_lo;
  assign new_n3307_ = ~n4587_lo;
  assign new_n3308_ = n4590_lo;
  assign new_n3310_ = n4593_lo;
  assign new_n3312_ = n4596_lo;
  assign new_n3314_ = n4602_lo;
  assign new_n3316_ = n4605_lo;
  assign new_n3318_ = n4608_lo;
  assign new_n3320_ = n4614_lo;
  assign new_n3322_ = n4617_lo;
  assign new_n3325_ = ~n4620_lo;
  assign new_n3326_ = n4626_lo;
  assign new_n3328_ = n4629_lo;
  assign new_n3331_ = ~n4632_lo;
  assign new_n3332_ = n4638_lo;
  assign new_n3334_ = n4641_lo;
  assign new_n3336_ = n4644_lo;
  assign new_n3338_ = n4647_lo;
  assign new_n3339_ = ~n4647_lo;
  assign new_n3340_ = n4650_lo;
  assign new_n3342_ = n4653_lo;
  assign new_n3344_ = n4656_lo;
  assign new_n3346_ = n4659_lo;
  assign new_n3347_ = ~n4659_lo;
  assign new_n3348_ = n4662_lo;
  assign new_n3350_ = n4665_lo;
  assign new_n3352_ = n4668_lo;
  assign new_n3354_ = n4671_lo;
  assign new_n3355_ = ~n4671_lo;
  assign new_n3356_ = n4674_lo;
  assign new_n3358_ = n4677_lo;
  assign new_n3360_ = n4680_lo;
  assign new_n3362_ = n4683_lo;
  assign new_n3363_ = ~n4683_lo;
  assign new_n3364_ = n4686_lo;
  assign new_n3366_ = n4689_lo;
  assign new_n3368_ = n4692_lo;
  assign new_n3370_ = n4695_lo;
  assign new_n3371_ = ~n4695_lo;
  assign new_n3372_ = n4698_lo;
  assign new_n3374_ = n4701_lo;
  assign new_n3376_ = n4704_lo;
  assign new_n3378_ = n4707_lo;
  assign new_n3379_ = ~n4707_lo;
  assign new_n3380_ = n4710_lo;
  assign new_n3382_ = n4713_lo;
  assign new_n3384_ = n4716_lo;
  assign new_n3385_ = ~n4716_lo;
  assign new_n3386_ = n4719_lo;
  assign new_n3387_ = ~n4719_lo;
  assign new_n3388_ = n4722_lo;
  assign new_n3390_ = n4725_lo;
  assign new_n3392_ = n4728_lo;
  assign new_n3393_ = ~n4728_lo;
  assign new_n3394_ = n4731_lo;
  assign new_n3395_ = ~n4731_lo;
  assign new_n3396_ = n4734_lo;
  assign new_n3398_ = n4737_lo;
  assign new_n3400_ = n4740_lo;
  assign new_n3403_ = ~n4743_lo;
  assign new_n3404_ = n4970_o2;
  assign new_n3405_ = ~n4970_o2;
  assign new_n3406_ = n4972_o2;
  assign new_n3407_ = ~n4972_o2;
  assign new_n3408_ = n4989_o2;
  assign new_n3409_ = ~n4989_o2;
  assign new_n3410_ = n5024_o2;
  assign new_n3411_ = ~n5024_o2;
  assign new_n3412_ = n5025_o2;
  assign new_n3413_ = ~n5025_o2;
  assign new_n3414_ = n5029_o2;
  assign new_n3415_ = ~n5029_o2;
  assign new_n3417_ = ~n5042_o2;
  assign new_n3419_ = ~n5048_o2;
  assign new_n3420_ = n5093_o2;
  assign new_n3421_ = ~n5093_o2;
  assign new_n3422_ = n5096_o2;
  assign new_n3423_ = ~n5096_o2;
  assign new_n3425_ = ~n5193_o2;
  assign new_n3426_ = n5199_o2;
  assign new_n3429_ = ~n5203_o2;
  assign new_n3431_ = ~n5214_o2;
  assign new_n3433_ = ~n5221_o2;
  assign new_n3434_ = n5222_o2;
  assign new_n3437_ = ~n5273_o2;
  assign new_n3438_ = n5365_o2;
  assign new_n3439_ = ~n5365_o2;
  assign new_n3440_ = n5385_o2;
  assign new_n3442_ = n5553_o2;
  assign new_n3443_ = ~n5553_o2;
  assign new_n3445_ = ~n5636_o2;
  assign new_n3446_ = n5782_o2;
  assign new_n3448_ = n5778_o2;
  assign new_n3449_ = ~n5778_o2;
  assign new_n3450_ = n5323_o2;
  assign new_n3451_ = ~n5323_o2;
  assign new_n3452_ = n5325_o2;
  assign new_n3453_ = ~n5325_o2;
  assign new_n3454_ = n5327_o2;
  assign new_n3455_ = ~n5327_o2;
  assign new_n3456_ = n5329_o2;
  assign new_n3457_ = ~n5329_o2;
  assign new_n3459_ = ~n5816_o2;
  assign new_n3461_ = ~n5817_o2;
  assign new_n3462_ = n5837_o2;
  assign new_n3463_ = ~n5837_o2;
  assign new_n3464_ = n5844_o2;
  assign new_n3466_ = n5859_o2;
  assign new_n3468_ = n5857_o2;
  assign new_n3470_ = n5369_o2;
  assign new_n3471_ = ~n5369_o2;
  assign new_n3472_ = n5371_o2;
  assign new_n3473_ = ~n5371_o2;
  assign new_n3474_ = n5373_o2;
  assign new_n3475_ = ~n5373_o2;
  assign new_n3476_ = n5400_o2;
  assign new_n3477_ = ~n5400_o2;
  assign new_n3478_ = n5402_o2;
  assign new_n3479_ = ~n5402_o2;
  assign new_n3480_ = n5404_o2;
  assign new_n3481_ = ~n5404_o2;
  assign new_n3482_ = n5406_o2;
  assign new_n3483_ = ~n5406_o2;
  assign new_n3484_ = n5407_o2;
  assign new_n3485_ = ~n5407_o2;
  assign new_n3486_ = n5408_o2;
  assign new_n3487_ = ~n5408_o2;
  assign new_n3489_ = ~n2722_o2;
  assign new_n3490_ = n1942_inv;
  assign new_n3492_ = n5412_o2;
  assign new_n3493_ = ~n5412_o2;
  assign new_n3494_ = n1948_inv;
  assign new_n3496_ = n5557_o2;
  assign new_n3497_ = ~n5557_o2;
  assign new_n3498_ = n5558_o2;
  assign new_n3500_ = n5559_o2;
  assign new_n3501_ = ~n5559_o2;
  assign new_n3502_ = n5564_o2;
  assign new_n3505_ = ~n5565_o2;
  assign new_n3506_ = n1966_inv;
  assign new_n3508_ = n5568_o2;
  assign new_n3509_ = ~n5568_o2;
  assign new_n3510_ = n5598_o2;
  assign new_n3511_ = ~n5598_o2;
  assign new_n3512_ = n5600_o2;
  assign new_n3513_ = ~n5600_o2;
  assign new_n3514_ = n5601_o2;
  assign new_n3516_ = n5602_o2;
  assign new_n3517_ = ~n5602_o2;
  assign new_n3518_ = n5603_o2;
  assign new_n3519_ = ~n5603_o2;
  assign new_n3520_ = n2853_o2;
  assign new_n3521_ = ~n2853_o2;
  assign new_n3522_ = n5637_o2;
  assign new_n3523_ = ~n5637_o2;
  assign new_n3524_ = n1993_inv;
  assign new_n3526_ = n1996_inv;
  assign new_n3528_ = n5635_o2;
  assign new_n3529_ = ~n5635_o2;
  assign new_n3530_ = n5640_o2;
  assign new_n3531_ = ~n5640_o2;
  assign new_n3532_ = n5641_o2;
  assign new_n3533_ = ~n5641_o2;
  assign new_n3534_ = n5642_o2;
  assign new_n3536_ = n5650_o2;
  assign new_n3537_ = ~n5650_o2;
  assign new_n3538_ = n5652_o2;
  assign new_n3540_ = n5653_o2;
  assign new_n3541_ = ~n5653_o2;
  assign new_n3542_ = n5654_o2;
  assign new_n3544_ = n5655_o2;
  assign new_n3545_ = ~n5655_o2;
  assign new_n3546_ = n5657_o2;
  assign new_n3548_ = n2029_inv;
  assign new_n3551_ = ~n5661_o2;
  assign new_n3552_ = n5656_o2;
  assign new_n3553_ = ~n5656_o2;
  assign new_n3554_ = n5663_o2;
  assign new_n3555_ = ~n5663_o2;
  assign new_n3556_ = n2041_inv;
  assign new_n3558_ = n5795_o2;
  assign new_n3559_ = ~n5795_o2;
  assign new_n3560_ = n5796_o2;
  assign new_n3561_ = ~n5796_o2;
  assign new_n3562_ = n5797_o2;
  assign new_n3563_ = ~n5797_o2;
  assign new_n3564_ = n5739_o2;
  assign new_n3565_ = ~n5739_o2;
  assign new_n3566_ = n5773_o2;
  assign new_n3568_ = n2059_inv;
  assign new_n3570_ = n5799_o2;
  assign new_n3571_ = ~n5799_o2;
  assign new_n3572_ = n5802_o2;
  assign new_n3574_ = n2068_inv;
  assign new_n3576_ = n5831_o2;
  assign new_n3577_ = ~n5831_o2;
  assign new_n3578_ = n5833_o2;
  assign new_n3579_ = ~n5833_o2;
  assign new_n3580_ = n5820_o2;
  assign new_n3582_ = n5823_o2;
  assign new_n3583_ = ~n5823_o2;
  assign new_n3585_ = ~n5824_o2;
  assign new_n3586_ = n5869_o2;
  assign new_n3588_ = n5848_o2;
  assign new_n3589_ = ~n5848_o2;
  assign new_n3590_ = n5849_o2;
  assign new_n3591_ = ~n5849_o2;
  assign new_n3592_ = n5856_o2;
  assign new_n3594_ = n5896_o2;
  assign new_n3595_ = ~n5896_o2;
  assign new_n3596_ = n2754_o2;
  assign new_n3598_ = n2908_o2;
  assign new_n3600_ = n5892_o2;
  assign new_n3602_ = n5915_o2;
  assign new_n3604_ = n5919_o2;
  assign new_n3606_ = n5918_o2;
  assign new_n3607_ = ~n5918_o2;
  assign new_n3608_ = n5920_o2;
  assign new_n3609_ = ~n5920_o2;
  assign new_n3610_ = n5917_o2;
  assign new_n3612_ = lo586_buf_o2;
  assign new_n3613_ = ~lo586_buf_o2;
  assign new_n3614_ = n2818_o2;
  assign new_n3616_ = n2863_o2;
  assign new_n3618_ = n2134_inv;
  assign new_n3619_ = ~n2134_inv;
  assign new_n3620_ = n2725_o2;
  assign new_n3621_ = ~n2725_o2;
  assign new_n3622_ = n3016_o2;
  assign new_n3623_ = ~n3016_o2;
  assign new_n3624_ = n3013_o2;
  assign new_n3625_ = ~n3013_o2;
  assign new_n3626_ = n2655_o2;
  assign new_n3627_ = ~n2655_o2;
  assign new_n3628_ = n2149_inv;
  assign new_n3629_ = ~n2149_inv;
  assign new_n3630_ = lo562_buf_o2;
  assign new_n3631_ = ~lo562_buf_o2;
  assign new_n3632_ = n2155_inv;
  assign new_n3634_ = n2531_o2;
  assign new_n3636_ = n2700_o2;
  assign new_n3637_ = ~n2700_o2;
  assign new_n3638_ = n5908_o2;
  assign new_n3639_ = ~n5908_o2;
  assign new_n3640_ = n5910_o2;
  assign new_n3641_ = ~n5910_o2;
  assign new_n3642_ = n5912_o2;
  assign new_n3643_ = ~n5912_o2;
  assign new_n3644_ = n5914_o2;
  assign new_n3645_ = ~n5914_o2;
  assign new_n3646_ = n2753_o2;
  assign new_n3647_ = ~n2753_o2;
  assign new_n3648_ = n2878_o2;
  assign new_n3649_ = ~n2878_o2;
  assign new_n3650_ = n2182_inv;
  assign new_n3652_ = n5934_o2;
  assign new_n3653_ = ~n5934_o2;
  assign new_n3654_ = n5936_o2;
  assign new_n3655_ = ~n5936_o2;
  assign new_n3656_ = n5938_o2;
  assign new_n3657_ = ~n5938_o2;
  assign new_n3658_ = n2728_o2;
  assign new_n3660_ = lo358_buf_o2;
  assign new_n3661_ = ~lo358_buf_o2;
  assign new_n3662_ = lo418_buf_o2;
  assign new_n3663_ = ~lo418_buf_o2;
  assign new_n3664_ = lo474_buf_o2;
  assign new_n3665_ = ~lo474_buf_o2;
  assign new_n3666_ = lo554_buf_o2;
  assign new_n3667_ = ~lo554_buf_o2;
  assign new_n3668_ = lo558_buf_o2;
  assign new_n3669_ = ~lo558_buf_o2;
  assign new_n3670_ = lo574_buf_o2;
  assign new_n3671_ = ~lo574_buf_o2;
  assign new_n3672_ = n2215_inv;
  assign new_n3674_ = n2218_inv;
  assign new_n3676_ = n2221_inv;
  assign new_n3678_ = lo450_buf_o2;
  assign new_n3679_ = ~lo450_buf_o2;
  assign new_n3680_ = n2910_o2;
  assign new_n3682_ = n2683_o2;
  assign new_n3683_ = ~n2683_o2;
  assign new_n3685_ = ~n2828_o2;
  assign new_n3686_ = n2582_o2;
  assign new_n3688_ = n2600_o2;
  assign new_n3690_ = n2542_o2;
  assign new_n3692_ = n2703_o2;
  assign new_n3694_ = lo510_buf_o2;
  assign new_n3695_ = ~lo510_buf_o2;
  assign new_n3696_ = lo514_buf_o2;
  assign new_n3698_ = lo538_buf_o2;
  assign new_n3699_ = ~lo538_buf_o2;
  assign new_n3700_ = lo578_buf_o2;
  assign new_n3701_ = ~lo578_buf_o2;
  assign new_n3702_ = n2260_inv;
  assign new_n3704_ = n2666_o2;
  assign new_n3706_ = n2667_o2;
  assign new_n3708_ = n2660_o2;
  assign new_n3709_ = ~n2660_o2;
  assign new_n3710_ = n2272_inv;
  assign new_n3712_ = lo454_buf_o2;
  assign new_n3714_ = n3593_o2;
  assign new_n3715_ = ~n3593_o2;
  assign new_n3716_ = n3048_o2;
  assign new_n3717_ = ~n3048_o2;
  assign new_n3718_ = lo410_buf_o2;
  assign new_n3719_ = ~lo410_buf_o2;
  assign new_n3720_ = lo502_buf_o2;
  assign new_n3721_ = ~lo502_buf_o2;
  assign new_n3722_ = lo506_buf_o2;
  assign new_n3724_ = lo550_buf_o2;
  assign new_n3725_ = ~lo550_buf_o2;
  assign new_n3726_ = lo570_buf_o2;
  assign new_n3727_ = ~lo570_buf_o2;
  assign new_n3728_ = lo582_buf_o2;
  assign new_n3729_ = ~lo582_buf_o2;
  assign new_n3730_ = n2302_inv;
  assign new_n3732_ = n2305_inv;
  assign new_n3734_ = n3499_o2;
  assign new_n3735_ = ~n3499_o2;
  assign new_n3736_ = n2311_inv;
  assign new_n3738_ = n2870_o2;
  assign new_n3740_ = n2317_inv;
  assign new_n3741_ = ~n2317_inv;
  assign new_n3742_ = n2689_o2;
  assign new_n3743_ = ~n2689_o2;
  assign new_n3744_ = n2323_inv;
  assign new_n3745_ = ~n2323_inv;
  assign new_n3746_ = n2662_o2;
  assign new_n3747_ = ~n2662_o2;
  assign new_n3748_ = lo350_buf_o2;
  assign new_n3749_ = ~lo350_buf_o2;
  assign new_n3750_ = lo498_buf_o2;
  assign new_n3752_ = lo518_buf_o2;
  assign new_n3753_ = ~lo518_buf_o2;
  assign new_n3754_ = lo522_buf_o2;
  assign new_n3756_ = lo598_buf_o2;
  assign new_n3757_ = ~lo598_buf_o2;
  assign new_n3758_ = n2344_inv;
  assign new_n3760_ = n2347_inv;
  assign new_n3762_ = n2350_inv;
  assign new_n3764_ = n2353_inv;
  assign new_n3765_ = ~n2353_inv;
  assign new_n3766_ = n2356_inv;
  assign new_n3768_ = n2359_inv;
  assign new_n3770_ = n2872_o2;
  assign new_n3772_ = n3313_o2;
  assign new_n3774_ = n3273_o2;
  assign new_n3776_ = n2848_o2;
  assign new_n3778_ = n2893_o2;
  assign new_n3780_ = n3267_o2;
  assign new_n3782_ = n2925_o2;
  assign new_n3785_ = ~n2839_o2;
  assign new_n3786_ = n2831_o2;
  assign new_n3788_ = n2558_o2;
  assign new_n3790_ = n2562_o2;
  assign new_n3792_ = n2825_o2;
  assign new_n3793_ = ~n2825_o2;
  assign new_n3794_ = n3263_o2;
  assign new_n3796_ = n3517_o2;
  assign new_n3798_ = n2873_o2;
  assign new_n3800_ = n2926_o2;
  assign new_n3803_ = ~n3261_o2;
  assign new_n3804_ = n3268_o2;
  assign new_n3806_ = n3274_o2;
  assign new_n3808_ = n3314_o2;
  assign new_n3811_ = ~n3571_o2;
  assign new_n3812_ = n2950_o2;
  assign new_n3813_ = ~n2950_o2;
  assign new_n3814_ = n2951_o2;
  assign new_n3815_ = ~n2951_o2;
  assign new_n3816_ = n3022_o2;
  assign new_n3818_ = n3023_o2;
  assign new_n3821_ = ~n3057_o2;
  assign new_n3822_ = n3058_o2;
  assign new_n3825_ = ~n2931_o2;
  assign new_n3826_ = n2911_o2;
  assign new_n3827_ = ~n2911_o2;
  assign new_n3828_ = n2959_o2;
  assign new_n3829_ = ~n2959_o2;
  assign new_n3830_ = n2960_o2;
  assign new_n3831_ = ~n2960_o2;
  assign new_n3833_ = ~n2922_o2;
  assign new_n3834_ = n2888_o2;
  assign new_n3837_ = ~n2889_o2;
  assign new_n3838_ = n3051_o2;
  assign new_n3841_ = ~n3052_o2;
  assign new_n3843_ = ~n3063_o2;
  assign new_n3844_ = n2845_o2;
  assign new_n3846_ = n2476_inv;
  assign new_n3848_ = n3281_o2;
  assign new_n3850_ = n3294_o2;
  assign new_n3852_ = n2885_o2;
  assign new_n3854_ = n2786_o2;
  assign new_n3855_ = ~n2786_o2;
  assign new_n3856_ = n2783_o2;
  assign new_n3857_ = ~n2783_o2;
  assign new_n3858_ = n2801_o2;
  assign new_n3859_ = ~n2801_o2;
  assign new_n3860_ = n2572_o2;
  assign new_n3861_ = ~n2572_o2;
  assign new_n3862_ = n2628_o2;
  assign new_n3863_ = ~n2628_o2;
  assign new_n3864_ = n2609_o2;
  assign new_n3865_ = ~n2609_o2;
  assign new_n3866_ = n2618_o2;
  assign new_n3867_ = ~n2618_o2;
  assign new_n3868_ = n2637_o2;
  assign new_n3869_ = ~n2637_o2;
  assign new_n3870_ = n2525_o2;
  assign new_n3871_ = ~n2525_o2;
  assign new_n3872_ = n2551_o2;
  assign new_n3874_ = n3759_o2;
  assign new_n3876_ = n2994_o2;
  assign new_n3877_ = ~n2994_o2;
  assign new_n3878_ = n3040_o2;
  assign new_n3879_ = ~n3040_o2;
  assign new_n3880_ = n2943_o2;
  assign new_n3881_ = ~n2943_o2;
  assign new_n3882_ = n2991_o2;
  assign new_n3883_ = ~n2991_o2;
  assign new_n3884_ = n3034_o2;
  assign new_n3885_ = ~n3034_o2;
  assign new_n3887_ = ~n2881_o2;
  assign new_n3889_ = ~n3021_o2;
  assign new_n3890_ = n3062_o2;
  assign new_n3892_ = n2763_o2;
  assign new_n3893_ = ~n2763_o2;
  assign new_n3894_ = n2764_o2;
  assign new_n3895_ = ~n2764_o2;
  assign new_n3896_ = n2775_o2;
  assign new_n3897_ = ~n2775_o2;
  assign new_n3898_ = n2776_o2;
  assign new_n3899_ = ~n2776_o2;
  assign new_n3900_ = n2968_o2;
  assign new_n3901_ = ~n2968_o2;
  assign new_n3902_ = n2969_o2;
  assign new_n3903_ = ~n2969_o2;
  assign new_n3904_ = n2798_o2;
  assign new_n3905_ = ~n2798_o2;
  assign new_n3907_ = ~n3661_o2;
  assign new_n3908_ = n2694_o2;
  assign new_n3909_ = ~n2694_o2;
  assign new_n3910_ = n2572_inv;
  assign new_n3911_ = ~n2572_inv;
  assign new_n3912_ = n2817_o2;
  assign new_n3913_ = ~n2817_o2;
  assign new_n3915_ = ~n2514_o2;
  assign new_n3917_ = ~n2501_o2;
  assign new_n3918_ = n2584_inv;
  assign new_n3920_ = n2505_o2;
  assign new_n3922_ = n2492_o2;
  assign new_n3923_ = ~n2492_o2;
  assign new_n3924_ = lo546_buf_o2;
  assign new_n3925_ = ~lo546_buf_o2;
  assign new_n3926_ = lo590_buf_o2;
  assign new_n3927_ = ~lo590_buf_o2;
  assign new_n3928_ = lo594_buf_o2;
  assign new_n3929_ = ~lo594_buf_o2;
  assign new_n3930_ = n2602_inv;
  assign new_n3932_ = n2605_inv;
  assign new_n3934_ = n2709_o2;
  assign new_n3935_ = ~n2709_o2;
  assign new_n3936_ = n2611_inv;
  assign new_n3937_ = ~n2611_inv;
  assign new_n3938_ = n2614_inv;
  assign new_n3939_ = ~n2614_inv;
  assign new_n3940_ = n2617_inv;
  assign new_n3941_ = ~n2617_inv;
  assign new_n3942_ = n2620_inv;
  assign new_n3943_ = ~n2620_inv;
  assign new_n3944_ = n3590_o2;
  assign new_n3945_ = ~n3590_o2;
  assign new_n3946_ = n3591_o2;
  assign new_n3947_ = ~n3591_o2;
  assign new_n3948_ = n2629_inv;
  assign new_n3949_ = ~n2629_inv;
  assign new_n3950_ = n3638_o2;
  assign new_n3951_ = ~n3638_o2;
  assign new_n3952_ = n3639_o2;
  assign new_n3953_ = ~n3639_o2;
  assign new_n3954_ = n2638_inv;
  assign new_n3955_ = ~n2638_inv;
  assign new_n3956_ = n2641_inv;
  assign new_n3957_ = ~n2641_inv;
  assign new_n3958_ = lo458_buf_o2;
  assign new_n3959_ = ~lo458_buf_o2;
  assign new_n3960_ = lo482_buf_o2;
  assign new_n3961_ = ~lo482_buf_o2;
  assign new_n3962_ = lo566_buf_o2;
  assign new_n3963_ = ~lo566_buf_o2;
  assign new_n3964_ = n2718_o2;
  assign new_n3965_ = ~n2718_o2;
  assign new_n3966_ = n3707_o2;
  assign new_n3967_ = ~n3707_o2;
  assign new_n3968_ = n3671_o2;
  assign new_n3969_ = ~n3671_o2;
  assign new_n3970_ = n3680_o2;
  assign new_n3971_ = ~n3680_o2;
  assign new_n3972_ = n3749_o2;
  assign new_n3973_ = ~n3749_o2;
  assign new_n3974_ = n3716_o2;
  assign new_n3975_ = ~n3716_o2;
  assign new_n3976_ = n3692_o2;
  assign new_n3977_ = ~n3692_o2;
  assign new_n3978_ = n2591_o2;
  assign new_n3979_ = ~n2591_o2;
  assign new_n3980_ = n3478_o2;
  assign new_n3981_ = ~n3478_o2;
  assign new_n3982_ = n3610_o2;
  assign new_n3983_ = ~n3610_o2;
  assign new_n3984_ = n3611_o2;
  assign new_n3985_ = ~n3611_o2;
  assign new_n3986_ = n2686_inv;
  assign new_n3988_ = n2689_inv;
  assign new_n3989_ = ~n2689_inv;
  assign new_n3990_ = n2738_o2;
  assign new_n3991_ = ~n2738_o2;
  assign new_n3992_ = n3616_o2;
  assign new_n3993_ = ~n3616_o2;
  assign new_n3994_ = n3617_o2;
  assign new_n3995_ = ~n3617_o2;
  assign new_n3996_ = n3031_o2;
  assign new_n3998_ = n2704_inv;
  assign new_n3999_ = ~n2704_inv;
  assign new_n4000_ = n3562_o2;
  assign new_n4001_ = ~n3562_o2;
  assign new_n4002_ = n2502_o2;
  assign new_n4003_ = ~n2502_o2;
  assign new_n4004_ = n3560_o2;
  assign new_n4005_ = ~n3560_o2;
  assign new_n4006_ = n3554_o2;
  assign new_n4007_ = ~n3554_o2;
  assign new_n4008_ = n3555_o2;
  assign new_n4009_ = ~n3555_o2;
  assign new_n4010_ = n3536_o2;
  assign new_n4011_ = ~n3536_o2;
  assign new_n4012_ = n3537_o2;
  assign new_n4013_ = ~n3537_o2;
  assign new_n4014_ = n3508_o2;
  assign new_n4015_ = ~n3508_o2;
  assign new_n4016_ = n3650_o2;
  assign new_n4017_ = ~n3650_o2;
  assign new_n4018_ = n3740_o2;
  assign new_n4019_ = ~n3740_o2;
  assign new_n4020_ = n3484_o2;
  assign new_n4021_ = ~n3484_o2;
  assign new_n4022_ = n2740_inv;
  assign new_n4023_ = ~n2740_inv;
  assign new_n4024_ = n2734_o2;
  assign new_n4025_ = ~n2734_o2;
  assign new_n4026_ = n2735_o2;
  assign new_n4027_ = ~n2735_o2;
  assign new_n4028_ = n2711_o2;
  assign new_n4029_ = ~n2711_o2;
  assign new_n4030_ = lo585_buf_o2;
  assign new_n4031_ = ~lo585_buf_o2;
  assign new_n4032_ = n2719_o2;
  assign new_n4033_ = ~n2719_o2;
  assign new_n4034_ = n2720_o2;
  assign new_n4035_ = ~n2720_o2;
  assign new_n4036_ = n2723_o2;
  assign new_n4037_ = ~n2723_o2;
  assign new_n4038_ = n2724_o2;
  assign new_n4039_ = ~n2724_o2;
  assign new_n4040_ = n3624_o2;
  assign new_n4041_ = ~n3624_o2;
  assign new_n4042_ = n3625_o2;
  assign new_n4043_ = ~n3625_o2;
  assign new_n4044_ = n3015_o2;
  assign new_n4045_ = ~n3015_o2;
  assign new_n4046_ = n3491_o2;
  assign new_n4047_ = ~n3491_o2;
  assign new_n4048_ = n2779_inv;
  assign new_n4049_ = ~n2779_inv;
  assign new_n4050_ = n2811_o2;
  assign new_n4051_ = ~n2811_o2;
  assign new_n4052_ = n3010_o2;
  assign new_n4053_ = ~n3010_o2;
  assign new_n4054_ = n3012_o2;
  assign new_n4055_ = ~n3012_o2;
  assign new_n4056_ = lo382_buf_o2;
  assign new_n4057_ = ~lo382_buf_o2;
  assign new_n4058_ = lo386_buf_o2;
  assign new_n4059_ = ~lo386_buf_o2;
  assign new_n4060_ = lo390_buf_o2;
  assign new_n4061_ = ~lo390_buf_o2;
  assign new_n4062_ = lo398_buf_o2;
  assign new_n4063_ = ~lo398_buf_o2;
  assign new_n4064_ = lo402_buf_o2;
  assign new_n4065_ = ~lo402_buf_o2;
  assign new_n4066_ = lo406_buf_o2;
  assign new_n4067_ = ~lo406_buf_o2;
  assign new_n4068_ = n3492_o2;
  assign new_n4069_ = ~n3492_o2;
  assign new_n4070_ = lo366_buf_o2;
  assign new_n4072_ = lo374_buf_o2;
  assign new_n4074_ = lo426_buf_o2;
  assign new_n4076_ = lo494_buf_o2;
  assign new_n4077_ = ~lo494_buf_o2;
  assign new_n4078_ = n2653_o2;
  assign new_n4079_ = ~n2653_o2;
  assign new_n4080_ = n2654_o2;
  assign new_n4081_ = ~n2654_o2;
  assign new_n4082_ = n2715_o2;
  assign new_n4083_ = ~n2715_o2;
  assign new_n4084_ = n2740_o2;
  assign new_n4085_ = ~n2740_o2;
  assign new_n4086_ = n2682_o2;
  assign new_n4087_ = ~n2682_o2;
  assign new_n4088_ = n2736_o2;
  assign new_n4089_ = ~n2736_o2;
  assign new_n4090_ = lo508_buf_o2;
  assign new_n4091_ = ~lo508_buf_o2;
  assign new_n4092_ = lo512_buf_o2;
  assign new_n4093_ = ~lo512_buf_o2;
  assign new_n4094_ = lo536_buf_o2;
  assign new_n4095_ = ~lo536_buf_o2;
  assign new_n4096_ = lo576_buf_o2;
  assign new_n4097_ = ~lo576_buf_o2;
  assign new_n4098_ = lo357_buf_o2;
  assign new_n4099_ = ~lo357_buf_o2;
  assign new_n4100_ = lo361_buf_o2;
  assign new_n4101_ = ~lo361_buf_o2;
  assign new_n4102_ = lo417_buf_o2;
  assign new_n4103_ = ~lo417_buf_o2;
  assign new_n4104_ = lo421_buf_o2;
  assign new_n4105_ = ~lo421_buf_o2;
  assign new_n4106_ = lo473_buf_o2;
  assign new_n4108_ = lo477_buf_o2;
  assign new_n4110_ = lo553_buf_o2;
  assign new_n4111_ = ~lo553_buf_o2;
  assign new_n4112_ = lo557_buf_o2;
  assign new_n4113_ = ~lo557_buf_o2;
  assign new_n4114_ = lo573_buf_o2;
  assign new_n4115_ = ~lo573_buf_o2;
  assign new_n4116_ = lo434_buf_o2;
  assign new_n4117_ = ~lo434_buf_o2;
  assign new_n4118_ = lo438_buf_o2;
  assign new_n4119_ = ~lo438_buf_o2;
  assign new_n4120_ = lo466_buf_o2;
  assign new_n4121_ = ~lo466_buf_o2;
  assign new_n4122_ = lo470_buf_o2;
  assign new_n4123_ = ~lo470_buf_o2;
  assign new_n4124_ = lo490_buf_o2;
  assign new_n4125_ = ~lo490_buf_o2;
  assign new_n4126_ = n2657_o2;
  assign new_n4127_ = ~n2657_o2;
  assign new_n4128_ = n2658_o2;
  assign new_n4129_ = ~n2658_o2;
  assign new_n4130_ = n2663_o2;
  assign new_n4131_ = ~n2663_o2;
  assign new_n4132_ = n2664_o2;
  assign new_n4133_ = ~n2664_o2;
  assign new_n4134_ = n2684_o2;
  assign new_n4135_ = ~n2684_o2;
  assign new_n4136_ = n2685_o2;
  assign new_n4137_ = ~n2685_o2;
  assign new_n4138_ = new_n6741_ | new_n6742_;
  assign new_n4139_ = new_n2904_ & new_n6745_;
  assign new_n4140_ = new_n3162_ & new_n6748_;
  assign new_n4141_ = new_n6749_ & new_n2872_;
  assign new_n4142_ = new_n3298_ | new_n6750_;
  assign new_n4143_ = new_n3225_ | new_n3171_;
  assign new_n4144_ = new_n2491_ | new_n6750_;
  assign new_n4145_ = new_n6754_ | new_n2889_;
  assign new_n4146_ = new_n6761_ | new_n2663_;
  assign new_n4147_ = new_n6766_ | new_n2655_;
  assign new_n4148_ = new_n4147_ & new_n4146_;
  assign new_n4149_ = new_n4148_ | new_n6754_;
  assign new_n4150_ = new_n6761_ | new_n2499_;
  assign new_n4151_ = new_n6766_ | new_n2671_;
  assign new_n4152_ = new_n4151_ & new_n4150_;
  assign new_n4153_ = new_n4152_ | new_n6753_;
  assign new_n4154_ = new_n6755_ | new_n2647_;
  assign new_n4155_ = new_n6762_ & new_n2466_;
  assign new_n4156_ = new_n6767_ & new_n2458_;
  assign new_n4157_ = new_n4156_ | new_n6755_;
  assign new_n4158_ = new_n4157_ | new_n4155_;
  assign new_n4159_ = new_n4158_ & new_n6745_;
  assign new_n4160_ = new_n6762_ & new_n2630_;
  assign new_n4161_ = new_n6767_ & new_n2474_;
  assign new_n4162_ = new_n4161_ | new_n6757_;
  assign new_n4163_ = new_n4162_ | new_n4160_;
  assign new_n4164_ = new_n4163_ & new_n6746_;
  assign new_n4165_ = new_n6763_ & new_n2450_;
  assign new_n4166_ = new_n6768_ & new_n2614_;
  assign new_n4167_ = new_n4166_ | new_n6757_;
  assign new_n4168_ = new_n4167_ | new_n4165_;
  assign new_n4169_ = new_n4168_ & new_n6746_;
  assign new_n4170_ = new_n6763_ & new_n2622_;
  assign new_n4171_ = new_n6768_ & new_n2638_;
  assign new_n4172_ = new_n4171_ | new_n6758_;
  assign new_n4173_ = new_n4172_ | new_n4170_;
  assign new_n4174_ = new_n4173_ & new_n6747_;
  assign new_n4175_ = new_n3468_ & new_n3466_;
  assign new_n4176_ = new_n3634_ & new_n3449_;
  assign new_n4177_ = new_n4176_ & new_n3870_;
  assign new_n4178_ = new_n6769_ & new_n3690_;
  assign new_n4179_ = new_n4178_ & new_n4177_;
  assign new_n4180_ = new_n4179_ & new_n4175_;
  assign new_n4181_ = new_n3866_ & new_n3864_;
  assign new_n4182_ = new_n4181_ & new_n3862_;
  assign new_n4183_ = new_n3790_ | new_n3788_;
  assign new_n4184_ = new_n6770_ & new_n3860_;
  assign new_n4185_ = new_n3686_ & new_n3464_;
  assign new_n4186_ = new_n3868_ & new_n3688_;
  assign new_n4187_ = new_n4186_ & new_n4185_;
  assign new_n4188_ = new_n4187_ & new_n4184_;
  assign new_n4189_ = new_n4188_ & new_n4182_;
  assign new_n4190_ = new_n6771_ | new_n3419_;
  assign new_n4191_ = new_n6772_ | new_n3461_;
  assign new_n4192_ = new_n3489_ & new_n3440_;
  assign new_n4193_ = new_n4192_ & new_n3426_;
  assign new_n4194_ = new_n3596_ & new_n3434_;
  assign new_n4195_ = new_n4194_ & new_n4193_;
  assign new_n4196_ = new_n3895_ & new_n3893_;
  assign new_n4197_ = new_n3894_ | new_n3892_;
  assign new_n4198_ = new_n3899_ & new_n3897_;
  assign new_n4199_ = new_n3898_ | new_n3896_;
  assign new_n4200_ = new_n4198_ & new_n4197_;
  assign new_n4201_ = new_n4199_ & new_n4196_;
  assign new_n4202_ = new_n4201_ | new_n4200_;
  assign new_n4203_ = new_n6773_ & new_n6774_;
  assign new_n4204_ = new_n6775_ | new_n6776_;
  assign new_n4205_ = new_n6775_ & new_n6776_;
  assign new_n4206_ = new_n6773_ | new_n6774_;
  assign new_n4207_ = new_n4206_ & new_n4204_;
  assign new_n4208_ = new_n4205_ | new_n4203_;
  assign new_n4209_ = new_n6777_ & new_n6778_;
  assign new_n4210_ = new_n6779_ | new_n6780_;
  assign new_n4211_ = new_n6779_ & new_n6780_;
  assign new_n4212_ = new_n6777_ | new_n6778_;
  assign new_n4213_ = new_n4212_ & new_n4210_;
  assign new_n4214_ = new_n4211_ | new_n4209_;
  assign new_n4215_ = new_n4213_ & new_n4208_;
  assign new_n4216_ = new_n4214_ & new_n4207_;
  assign new_n4217_ = new_n4216_ | new_n4215_;
  assign new_n4218_ = new_n6772_ | new_n3459_;
  assign new_n4219_ = new_n6771_ | new_n3429_;
  assign new_n4220_ = new_n3433_ | new_n3417_;
  assign new_n4221_ = new_n4220_ & new_n3425_;
  assign new_n4222_ = new_n4221_ & new_n4219_;
  assign new_n4223_ = new_n4222_ & new_n4218_;
  assign new_n4224_ = new_n6782_ | new_n3431_;
  assign new_n4225_ = new_n6786_ & new_n3685_;
  assign new_n4226_ = new_n3448_ | new_n6801_;
  assign new_n4227_ = new_n3786_ & new_n6809_;
  assign new_n4228_ = new_n4227_ & new_n4226_;
  assign new_n4229_ = new_n4228_ | new_n4225_;
  assign new_n4230_ = new_n6820_ | new_n3439_;
  assign new_n4231_ = new_n6769_ & new_n6824_;
  assign new_n4232_ = new_n3785_ | new_n6830_;
  assign new_n4233_ = new_n4232_ | new_n4231_;
  assign new_n4234_ = new_n4233_ & new_n4230_;
  assign new_n4235_ = new_n6832_ & new_n6786_;
  assign new_n4236_ = new_n3861_ | new_n6801_;
  assign new_n4237_ = new_n3776_ & new_n6809_;
  assign new_n4238_ = new_n4237_ & new_n4236_;
  assign new_n4239_ = new_n4238_ | new_n4235_;
  assign new_n4240_ = new_n6835_ | new_n6841_;
  assign new_n4241_ = new_n6858_ | new_n6864_;
  assign new_n4242_ = new_n4241_ & new_n4240_;
  assign new_n4243_ = new_n4242_ & new_n6882_;
  assign new_n4244_ = new_n6841_ | new_n6888_;
  assign new_n4245_ = new_n6864_ | new_n6889_;
  assign new_n4246_ = new_n4245_ & new_n4244_;
  assign new_n4247_ = new_n4246_ & new_n6893_;
  assign new_n4248_ = new_n4247_ | new_n4243_;
  assign new_n4249_ = new_n6787_ & new_n6899_;
  assign new_n4250_ = new_n3798_ | new_n3770_;
  assign new_n4251_ = new_n4250_ & new_n6810_;
  assign new_n4252_ = new_n4251_ | new_n4249_;
  assign new_n4253_ = new_n6900_ & new_n6787_;
  assign new_n4254_ = new_n3852_ & new_n6810_;
  assign new_n4255_ = new_n4254_ | new_n4253_;
  assign new_n4256_ = new_n3837_ | new_n3834_;
  assign new_n4257_ = new_n6901_ & new_n6789_;
  assign new_n4258_ = new_n3871_ | new_n6800_;
  assign new_n4259_ = new_n3778_ & new_n6812_;
  assign new_n4260_ = new_n4259_ & new_n4258_;
  assign new_n4261_ = new_n4260_ | new_n4257_;
  assign new_n4262_ = new_n6835_ | new_n6906_;
  assign new_n4263_ = new_n6858_ | new_n6925_;
  assign new_n4264_ = new_n4263_ & new_n4262_;
  assign new_n4265_ = new_n4264_ & new_n6943_;
  assign new_n4266_ = new_n6906_ | new_n6888_;
  assign new_n4267_ = new_n6925_ | new_n6889_;
  assign new_n4268_ = new_n4267_ & new_n4266_;
  assign new_n4269_ = new_n4268_ & new_n6952_;
  assign new_n4270_ = new_n4269_ | new_n4265_;
  assign new_n4271_ = new_n3827_ & new_n3443_;
  assign new_n4272_ = new_n3826_ & new_n3442_;
  assign new_n4273_ = new_n4272_ | new_n4271_;
  assign new_n4274_ = new_n6958_ & new_n6789_;
  assign new_n4275_ = new_n6802_ & new_n2800_;
  assign new_n4276_ = new_n3865_ & new_n6824_;
  assign new_n4277_ = new_n4276_ | new_n4275_;
  assign new_n4278_ = new_n4277_ & new_n6812_;
  assign new_n4279_ = new_n4278_ | new_n4274_;
  assign new_n4280_ = new_n3833_ | new_n3680_;
  assign new_n4281_ = new_n6959_ & new_n6790_;
  assign new_n4282_ = new_n3800_ | new_n3782_;
  assign new_n4283_ = new_n4282_ & new_n6813_;
  assign new_n4284_ = new_n4283_ | new_n4281_;
  assign new_n4285_ = new_n3825_ | new_n3598_;
  assign new_n4286_ = new_n6960_ & new_n6790_;
  assign new_n4287_ = new_n6802_ & new_n2824_;
  assign new_n4288_ = new_n3863_ & new_n6823_;
  assign new_n4289_ = new_n4288_ | new_n4287_;
  assign new_n4290_ = new_n4289_ & new_n6813_;
  assign new_n4291_ = new_n4290_ | new_n4286_;
  assign new_n4292_ = new_n3880_ | new_n6820_;
  assign new_n4293_ = new_n6770_ & new_n6825_;
  assign new_n4294_ = new_n6804_ & new_n2817_;
  assign new_n4295_ = new_n4294_ | new_n6830_;
  assign new_n4296_ = new_n4295_ | new_n4293_;
  assign new_n4297_ = new_n4296_ & new_n4292_;
  assign new_n4298_ = new_n3815_ & new_n3813_;
  assign new_n4299_ = new_n3814_ | new_n3812_;
  assign new_n4300_ = new_n6961_ & new_n6964_;
  assign new_n4301_ = new_n6966_ | new_n6968_;
  assign new_n4302_ = new_n6966_ & new_n6968_;
  assign new_n4303_ = new_n6961_ | new_n6964_;
  assign new_n4304_ = new_n4303_ & new_n4301_;
  assign new_n4305_ = new_n4302_ | new_n4300_;
  assign new_n4306_ = new_n3831_ & new_n3828_;
  assign new_n4307_ = new_n3830_ | new_n3829_;
  assign new_n4308_ = new_n3903_ & new_n3900_;
  assign new_n4309_ = new_n3902_ | new_n3901_;
  assign new_n4310_ = new_n6970_ & new_n6971_;
  assign new_n4311_ = new_n6972_ | new_n6973_;
  assign new_n4312_ = new_n6972_ & new_n6973_;
  assign new_n4313_ = new_n6970_ | new_n6971_;
  assign new_n4314_ = new_n4313_ & new_n4311_;
  assign new_n4315_ = new_n4312_ | new_n4310_;
  assign new_n4316_ = new_n4314_ & new_n4305_;
  assign new_n4317_ = new_n4315_ & new_n4304_;
  assign new_n4318_ = new_n4317_ | new_n4316_;
  assign new_n4319_ = new_n6974_ & new_n6975_;
  assign new_n4320_ = new_n6976_ | new_n6977_;
  assign new_n4321_ = new_n6976_ & new_n6977_;
  assign new_n4322_ = new_n6974_ | new_n6975_;
  assign new_n4323_ = new_n4322_ & new_n4320_;
  assign new_n4324_ = new_n4321_ | new_n4319_;
  assign new_n4325_ = new_n6978_ & new_n6979_;
  assign new_n4326_ = new_n6980_ | new_n6981_;
  assign new_n4327_ = new_n6980_ & new_n6981_;
  assign new_n4328_ = new_n6978_ | new_n6979_;
  assign new_n4329_ = new_n4328_ & new_n4326_;
  assign new_n4330_ = new_n4327_ | new_n4325_;
  assign new_n4331_ = new_n6982_ & new_n6983_;
  assign new_n4332_ = new_n6984_ | new_n6985_;
  assign new_n4333_ = new_n6984_ & new_n6985_;
  assign new_n4334_ = new_n6982_ | new_n6983_;
  assign new_n4335_ = new_n4334_ & new_n4332_;
  assign new_n4336_ = new_n4333_ | new_n4331_;
  assign new_n4337_ = new_n6986_ & new_n6987_;
  assign new_n4338_ = new_n6988_ | new_n6989_;
  assign new_n4339_ = new_n6988_ & new_n6989_;
  assign new_n4340_ = new_n6986_ | new_n6987_;
  assign new_n4341_ = new_n4340_ & new_n4338_;
  assign new_n4342_ = new_n4339_ | new_n4337_;
  assign new_n4343_ = new_n6990_ & new_n6991_;
  assign new_n4344_ = new_n6992_ | new_n6993_;
  assign new_n4345_ = new_n6992_ & new_n6993_;
  assign new_n4346_ = new_n6990_ | new_n6991_;
  assign new_n4347_ = new_n4346_ & new_n4344_;
  assign new_n4348_ = new_n4345_ | new_n4343_;
  assign new_n4349_ = new_n6994_ & new_n6995_;
  assign new_n4350_ = new_n6996_ | new_n6997_;
  assign new_n4351_ = new_n6996_ & new_n6997_;
  assign new_n4352_ = new_n6994_ | new_n6995_;
  assign new_n4353_ = new_n4352_ & new_n4350_;
  assign new_n4354_ = new_n4351_ | new_n4349_;
  assign new_n4355_ = new_n4353_ & new_n4336_;
  assign new_n4356_ = new_n4354_ & new_n4335_;
  assign new_n4357_ = new_n4356_ | new_n4355_;
  assign new_n4358_ = new_n3818_ | new_n3816_;
  assign new_n4359_ = new_n3881_ | new_n6832_;
  assign new_n4360_ = new_n4359_ | new_n6960_;
  assign new_n4361_ = new_n4360_ | new_n6959_;
  assign new_n4362_ = new_n4361_ | new_n6958_;
  assign new_n4363_ = new_n4362_ | new_n6998_;
  assign new_n4364_ = new_n4363_ | new_n6999_;
  assign new_n4365_ = new_n3884_ | new_n3423_;
  assign new_n4366_ = new_n3885_ | new_n3422_;
  assign new_n4367_ = new_n4366_ & new_n4365_;
  assign new_n4368_ = new_n3879_ | new_n3415_;
  assign new_n4369_ = new_n3878_ | new_n3414_;
  assign new_n4370_ = new_n4369_ & new_n4368_;
  assign new_n4371_ = new_n7000_ | new_n7001_;
  assign new_n4372_ = new_n4371_ | new_n4364_;
  assign new_n4373_ = new_n3841_ & new_n3838_;
  assign new_n4374_ = new_n3822_ & new_n3821_;
  assign new_n4375_ = new_n3843_ | new_n3438_;
  assign new_n4376_ = new_n4375_ | new_n6901_;
  assign new_n4377_ = new_n4376_ | new_n6899_;
  assign new_n4378_ = new_n4377_ | new_n6900_;
  assign new_n4379_ = new_n4378_ | new_n7002_;
  assign new_n4380_ = new_n4379_ | new_n7003_;
  assign new_n4381_ = new_n4380_ | new_n7004_;
  assign new_n4382_ = new_n6857_ & new_n7009_;
  assign new_n4383_ = new_n6834_ & new_n7028_;
  assign new_n4384_ = new_n4383_ | new_n7046_;
  assign new_n4385_ = new_n4384_ | new_n4382_;
  assign new_n4386_ = new_n7009_ & new_n7052_;
  assign new_n4387_ = new_n7028_ & new_n7053_;
  assign new_n4388_ = new_n4387_ | new_n7057_;
  assign new_n4389_ = new_n4388_ | new_n4386_;
  assign new_n4390_ = new_n4389_ & new_n7067_;
  assign new_n4391_ = new_n4390_ & new_n4385_;
  assign new_n4392_ = new_n6859_ & new_n7083_;
  assign new_n4393_ = new_n6836_ & new_n7102_;
  assign new_n4394_ = new_n4393_ | new_n7120_;
  assign new_n4395_ = new_n4394_ | new_n4392_;
  assign new_n4396_ = new_n7083_ & new_n7052_;
  assign new_n4397_ = new_n7102_ & new_n7053_;
  assign new_n4398_ = new_n4397_ | new_n7129_;
  assign new_n4399_ = new_n4398_ | new_n4396_;
  assign new_n4400_ = new_n4399_ & new_n7067_;
  assign new_n4401_ = new_n4400_ & new_n4395_;
  assign new_n4402_ = new_n6865_ | new_n7135_;
  assign new_n4403_ = new_n6842_ | new_n7136_;
  assign new_n4404_ = new_n4403_ & new_n4402_;
  assign new_n4405_ = new_n4404_ | new_n6882_;
  assign new_n4406_ = new_n7139_ & new_n6842_;
  assign new_n4407_ = new_n7143_ & new_n6865_;
  assign new_n4408_ = new_n4407_ | new_n6893_;
  assign new_n4409_ = new_n4408_ | new_n4406_;
  assign new_n4410_ = new_n4409_ & new_n4405_;
  assign new_n4411_ = new_n6867_ | new_n7145_;
  assign new_n4412_ = new_n6844_ | new_n7146_;
  assign new_n4413_ = new_n4412_ & new_n4411_;
  assign new_n4414_ = new_n4413_ | new_n6883_;
  assign new_n4415_ = new_n7149_ & new_n6844_;
  assign new_n4416_ = new_n7153_ & new_n6867_;
  assign new_n4417_ = new_n4416_ | new_n6894_;
  assign new_n4418_ = new_n4417_ | new_n4415_;
  assign new_n4419_ = new_n4418_ & new_n4414_;
  assign new_n4420_ = new_n6868_ | new_n7155_;
  assign new_n4421_ = new_n6845_ | new_n7156_;
  assign new_n4422_ = new_n4421_ & new_n4420_;
  assign new_n4423_ = new_n4422_ | new_n6883_;
  assign new_n4424_ = new_n7159_ & new_n6845_;
  assign new_n4425_ = new_n7163_ & new_n6868_;
  assign new_n4426_ = new_n4425_ | new_n6894_;
  assign new_n4427_ = new_n4426_ | new_n4424_;
  assign new_n4428_ = new_n4427_ & new_n4423_;
  assign new_n4429_ = new_n6870_ | new_n7165_;
  assign new_n4430_ = new_n6847_ | new_n7166_;
  assign new_n4431_ = new_n4430_ & new_n4429_;
  assign new_n4432_ = new_n4431_ | new_n6884_;
  assign new_n4433_ = new_n7169_ & new_n6847_;
  assign new_n4434_ = new_n7173_ & new_n6870_;
  assign new_n4435_ = new_n4434_ | new_n6895_;
  assign new_n4436_ = new_n4435_ | new_n4433_;
  assign new_n4437_ = new_n4436_ & new_n4432_;
  assign new_n4438_ = new_n6926_ | new_n7135_;
  assign new_n4439_ = new_n6907_ | new_n7136_;
  assign new_n4440_ = new_n4439_ & new_n4438_;
  assign new_n4441_ = new_n4440_ | new_n6943_;
  assign new_n4442_ = new_n7139_ & new_n6907_;
  assign new_n4443_ = new_n7143_ & new_n6926_;
  assign new_n4444_ = new_n4443_ | new_n6952_;
  assign new_n4445_ = new_n4444_ | new_n4442_;
  assign new_n4446_ = new_n4445_ & new_n4441_;
  assign new_n4447_ = new_n6928_ | new_n7145_;
  assign new_n4448_ = new_n6909_ | new_n7146_;
  assign new_n4449_ = new_n4448_ & new_n4447_;
  assign new_n4450_ = new_n4449_ | new_n6944_;
  assign new_n4451_ = new_n7149_ & new_n6909_;
  assign new_n4452_ = new_n7153_ & new_n6928_;
  assign new_n4453_ = new_n4452_ | new_n6953_;
  assign new_n4454_ = new_n4453_ | new_n4451_;
  assign new_n4455_ = new_n4454_ & new_n4450_;
  assign new_n4456_ = new_n6929_ | new_n7155_;
  assign new_n4457_ = new_n6910_ | new_n7156_;
  assign new_n4458_ = new_n4457_ & new_n4456_;
  assign new_n4459_ = new_n4458_ | new_n6944_;
  assign new_n4460_ = new_n7159_ & new_n6910_;
  assign new_n4461_ = new_n7163_ & new_n6929_;
  assign new_n4462_ = new_n4461_ | new_n6953_;
  assign new_n4463_ = new_n4462_ | new_n4460_;
  assign new_n4464_ = new_n4463_ & new_n4459_;
  assign new_n4465_ = new_n6931_ | new_n7165_;
  assign new_n4466_ = new_n6912_ | new_n7166_;
  assign new_n4467_ = new_n4466_ & new_n4465_;
  assign new_n4468_ = new_n4467_ | new_n6945_;
  assign new_n4469_ = new_n7169_ & new_n6912_;
  assign new_n4470_ = new_n7173_ & new_n6931_;
  assign new_n4471_ = new_n4470_ | new_n6954_;
  assign new_n4472_ = new_n4471_ | new_n4469_;
  assign new_n4473_ = new_n4472_ & new_n4468_;
  assign new_n4474_ = new_n7138_ & new_n7010_;
  assign new_n4475_ = new_n7142_ & new_n7029_;
  assign new_n4476_ = new_n4475_ | new_n7046_;
  assign new_n4477_ = new_n4476_ | new_n4474_;
  assign new_n4478_ = new_n7010_ & new_n7175_;
  assign new_n4479_ = new_n7029_ & new_n7176_;
  assign new_n4480_ = new_n4479_ | new_n7057_;
  assign new_n4481_ = new_n4480_ | new_n4478_;
  assign new_n4482_ = new_n4481_ & new_n7066_;
  assign new_n4483_ = new_n4482_ & new_n4477_;
  assign new_n4484_ = new_n7168_ | new_n7031_;
  assign new_n4485_ = new_n7172_ | new_n7012_;
  assign new_n4486_ = new_n4485_ & new_n7058_;
  assign new_n4487_ = new_n4486_ & new_n4484_;
  assign new_n4488_ = new_n7031_ | new_n7177_;
  assign new_n4489_ = new_n7012_ | new_n7178_;
  assign new_n4490_ = new_n4489_ & new_n7047_;
  assign new_n4491_ = new_n4490_ & new_n4488_;
  assign new_n4492_ = new_n4491_ | new_n7180_;
  assign new_n4493_ = new_n4492_ | new_n4487_;
  assign new_n4494_ = new_n7158_ & new_n7013_;
  assign new_n4495_ = new_n7162_ & new_n7032_;
  assign new_n4496_ = new_n4495_ | new_n7047_;
  assign new_n4497_ = new_n4496_ | new_n4494_;
  assign new_n4498_ = new_n7013_ & new_n7182_;
  assign new_n4499_ = new_n7032_ & new_n7183_;
  assign new_n4500_ = new_n4499_ | new_n7058_;
  assign new_n4501_ = new_n4500_ | new_n4498_;
  assign new_n4502_ = new_n4501_ & new_n7068_;
  assign new_n4503_ = new_n4502_ & new_n4497_;
  assign new_n4504_ = new_n7148_ & new_n7015_;
  assign new_n4505_ = new_n7152_ & new_n7034_;
  assign new_n4506_ = new_n4505_ | new_n7048_;
  assign new_n4507_ = new_n4506_ | new_n4504_;
  assign new_n4508_ = new_n7015_ & new_n7184_;
  assign new_n4509_ = new_n7034_ & new_n7185_;
  assign new_n4510_ = new_n4509_ | new_n7059_;
  assign new_n4511_ = new_n4510_ | new_n4508_;
  assign new_n4512_ = new_n4511_ & new_n7068_;
  assign new_n4513_ = new_n4512_ & new_n4507_;
  assign new_n4514_ = new_n7140_ & new_n7084_;
  assign new_n4515_ = new_n7144_ & new_n7103_;
  assign new_n4516_ = new_n4515_ | new_n7120_;
  assign new_n4517_ = new_n4516_ | new_n4514_;
  assign new_n4518_ = new_n7084_ & new_n7175_;
  assign new_n4519_ = new_n7103_ & new_n7176_;
  assign new_n4520_ = new_n4519_ | new_n7129_;
  assign new_n4521_ = new_n4520_ | new_n4518_;
  assign new_n4522_ = new_n4521_ & new_n7070_;
  assign new_n4523_ = new_n4522_ & new_n4517_;
  assign new_n4524_ = new_n7170_ | new_n7105_;
  assign new_n4525_ = new_n7174_ | new_n7086_;
  assign new_n4526_ = new_n4525_ & new_n7130_;
  assign new_n4527_ = new_n4526_ & new_n4524_;
  assign new_n4528_ = new_n7105_ | new_n7177_;
  assign new_n4529_ = new_n7086_ | new_n7178_;
  assign new_n4530_ = new_n4529_ & new_n7121_;
  assign new_n4531_ = new_n4530_ & new_n4528_;
  assign new_n4532_ = new_n4531_ | new_n7180_;
  assign new_n4533_ = new_n4532_ | new_n4527_;
  assign new_n4534_ = new_n7160_ & new_n7087_;
  assign new_n4535_ = new_n7164_ & new_n7106_;
  assign new_n4536_ = new_n4535_ | new_n7121_;
  assign new_n4537_ = new_n4536_ | new_n4534_;
  assign new_n4538_ = new_n7087_ & new_n7182_;
  assign new_n4539_ = new_n7106_ & new_n7183_;
  assign new_n4540_ = new_n4539_ | new_n7130_;
  assign new_n4541_ = new_n4540_ | new_n4538_;
  assign new_n4542_ = new_n4541_ & new_n7070_;
  assign new_n4543_ = new_n4542_ & new_n4537_;
  assign new_n4544_ = new_n7089_ & new_n7184_;
  assign new_n4545_ = new_n7108_ & new_n7185_;
  assign new_n4546_ = new_n4545_ | new_n4544_;
  assign new_n4547_ = new_n4546_ & new_n7122_;
  assign new_n4548_ = new_n7150_ | new_n7108_;
  assign new_n4549_ = new_n7154_ | new_n7089_;
  assign new_n4550_ = new_n4549_ & new_n7131_;
  assign new_n4551_ = new_n4550_ & new_n4548_;
  assign new_n4552_ = new_n4551_ | new_n4547_;
  assign new_n4553_ = new_n4552_ & new_n7071_;
  assign new_n4554_ = new_n3403_ | new_n2865_;
  assign new_n4555_ = new_n7186_ & new_n2808_;
  assign new_n4556_ = new_n6963_ & new_n7187_;
  assign new_n4557_ = new_n4556_ | new_n4555_;
  assign new_n4558_ = new_n4557_ & new_n3338_;
  assign new_n4559_ = new_n6782_ & new_n7188_;
  assign new_n4560_ = new_n7189_ | new_n7190_;
  assign new_n4561_ = new_n7189_ & new_n7190_;
  assign new_n4562_ = new_n6781_ | new_n7188_;
  assign new_n4563_ = new_n4562_ & new_n4560_;
  assign new_n4564_ = new_n4561_ | new_n4559_;
  assign new_n4565_ = new_n7191_ & new_n7187_;
  assign new_n4566_ = new_n3446_ & new_n7186_;
  assign new_n4567_ = new_n4566_ | new_n4565_;
  assign new_n4568_ = new_n4567_ & new_n3339_;
  assign new_n4569_ = new_n4568_ | new_n4558_;
  assign new_n4570_ = new_n4569_ & new_n4554_;
  assign new_n4571_ = new_n4563_ | new_n6969_;
  assign new_n4572_ = new_n7191_ | new_n6965_;
  assign new_n4573_ = new_n4572_ & new_n4571_;
  assign new_n4574_ = new_n6793_ & new_n6965_;
  assign new_n4575_ = new_n3803_ & new_n3794_;
  assign new_n4576_ = new_n4575_ | new_n4574_;
  assign new_n4577_ = new_n7004_ & new_n6793_;
  assign new_n4578_ = new_n3804_ | new_n3780_;
  assign new_n4579_ = new_n4578_ & new_n6816_;
  assign new_n4580_ = new_n4579_ | new_n4577_;
  assign new_n4581_ = new_n7003_ & new_n6794_;
  assign new_n4582_ = new_n3806_ | new_n3774_;
  assign new_n4583_ = new_n4582_ & new_n6816_;
  assign new_n4584_ = new_n4583_ | new_n4581_;
  assign new_n4585_ = new_n7002_ & new_n6794_;
  assign new_n4586_ = new_n3848_ & new_n6817_;
  assign new_n4587_ = new_n4586_ | new_n4585_;
  assign new_n4588_ = new_n7192_ | new_n7193_;
  assign new_n4589_ = new_n4588_ | new_n7194_;
  assign new_n4590_ = new_n4589_ | new_n7195_;
  assign new_n4591_ = new_n4590_ | new_n7196_;
  assign new_n4592_ = new_n4591_ | new_n7197_;
  assign new_n4593_ = new_n4592_ | new_n7198_;
  assign new_n4594_ = new_n4593_ | new_n7199_;
  assign new_n4595_ = new_n6999_ & new_n6796_;
  assign new_n4596_ = new_n3850_ & new_n6817_;
  assign new_n4597_ = new_n4596_ | new_n4595_;
  assign new_n4598_ = new_n7001_ & new_n6796_;
  assign new_n4599_ = new_n6804_ & new_n2746_;
  assign new_n4600_ = new_n3867_ & new_n6825_;
  assign new_n4601_ = new_n4600_ | new_n4599_;
  assign new_n4602_ = new_n4601_ & new_n6819_;
  assign new_n4603_ = new_n4602_ | new_n4598_;
  assign new_n4604_ = new_n7000_ & new_n6797_;
  assign new_n4605_ = new_n6805_ & new_n2552_;
  assign new_n4606_ = new_n3869_ & new_n6827_;
  assign new_n4607_ = new_n4606_ | new_n4605_;
  assign new_n4608_ = new_n4607_ & new_n6819_;
  assign new_n4609_ = new_n4608_ | new_n4604_;
  assign new_n4610_ = new_n6998_ & new_n6797_;
  assign new_n4611_ = new_n3808_ | new_n3772_;
  assign new_n4612_ = new_n4611_ & new_n6818_;
  assign new_n4613_ = new_n4612_ | new_n4610_;
  assign new_n4614_ = new_n6913_ & new_n7200_;
  assign new_n4615_ = new_n6932_ & new_n7201_;
  assign new_n4616_ = new_n4615_ | new_n4614_;
  assign new_n4617_ = new_n4616_ & new_n6954_;
  assign new_n4618_ = new_n7204_ & new_n6913_;
  assign new_n4619_ = new_n7208_ & new_n6932_;
  assign new_n4620_ = new_n4619_ | new_n4618_;
  assign new_n4621_ = new_n4620_ & new_n6945_;
  assign new_n4622_ = new_n4621_ | new_n4617_;
  assign new_n4623_ = new_n7204_ & new_n6848_;
  assign new_n4624_ = new_n7208_ & new_n6871_;
  assign new_n4625_ = new_n4624_ | new_n6895_;
  assign new_n4626_ = new_n4625_ | new_n4623_;
  assign new_n4627_ = new_n6871_ | new_n7200_;
  assign new_n4628_ = new_n6848_ | new_n7201_;
  assign new_n4629_ = new_n4628_ & new_n4627_;
  assign new_n4630_ = new_n4629_ | new_n6884_;
  assign new_n4631_ = new_n4630_ & new_n4626_;
  assign new_n4632_ = new_n6874_ | new_n7210_;
  assign new_n4633_ = new_n6851_ | new_n7211_;
  assign new_n4634_ = new_n4633_ & new_n4632_;
  assign new_n4635_ = new_n4634_ | new_n6886_;
  assign new_n4636_ = new_n7214_ & new_n6851_;
  assign new_n4637_ = new_n7218_ & new_n6874_;
  assign new_n4638_ = new_n4637_ | new_n6897_;
  assign new_n4639_ = new_n4638_ | new_n4636_;
  assign new_n4640_ = new_n4639_ & new_n4635_;
  assign new_n4641_ = new_n6875_ | new_n7220_;
  assign new_n4642_ = new_n6852_ | new_n7221_;
  assign new_n4643_ = new_n4642_ & new_n4641_;
  assign new_n4644_ = new_n4643_ | new_n6886_;
  assign new_n4645_ = new_n7224_ & new_n6852_;
  assign new_n4646_ = new_n7228_ & new_n6875_;
  assign new_n4647_ = new_n4646_ | new_n6897_;
  assign new_n4648_ = new_n4647_ | new_n4645_;
  assign new_n4649_ = new_n4648_ & new_n4644_;
  assign new_n4650_ = new_n6877_ | new_n7230_;
  assign new_n4651_ = new_n6854_ | new_n7231_;
  assign new_n4652_ = new_n4651_ & new_n4650_;
  assign new_n4653_ = new_n4652_ | new_n6887_;
  assign new_n4654_ = new_n7234_ & new_n6854_;
  assign new_n4655_ = new_n7238_ & new_n6877_;
  assign new_n4656_ = new_n4655_ | new_n6898_;
  assign new_n4657_ = new_n4656_ | new_n4654_;
  assign new_n4658_ = new_n4657_ & new_n4653_;
  assign new_n4659_ = new_n6935_ | new_n7210_;
  assign new_n4660_ = new_n6916_ | new_n7211_;
  assign new_n4661_ = new_n4660_ & new_n4659_;
  assign new_n4662_ = new_n4661_ | new_n6947_;
  assign new_n4663_ = new_n7214_ & new_n6916_;
  assign new_n4664_ = new_n7218_ & new_n6935_;
  assign new_n4665_ = new_n4664_ | new_n6956_;
  assign new_n4666_ = new_n4665_ | new_n4663_;
  assign new_n4667_ = new_n4666_ & new_n4662_;
  assign new_n4668_ = new_n6936_ | new_n7220_;
  assign new_n4669_ = new_n6917_ | new_n7221_;
  assign new_n4670_ = new_n4669_ & new_n4668_;
  assign new_n4671_ = new_n4670_ | new_n6947_;
  assign new_n4672_ = new_n7224_ & new_n6917_;
  assign new_n4673_ = new_n7228_ & new_n6936_;
  assign new_n4674_ = new_n4673_ | new_n6956_;
  assign new_n4675_ = new_n4674_ | new_n4672_;
  assign new_n4676_ = new_n4675_ & new_n4671_;
  assign new_n4677_ = new_n6938_ | new_n7230_;
  assign new_n4678_ = new_n6919_ | new_n7231_;
  assign new_n4679_ = new_n4678_ & new_n4677_;
  assign new_n4680_ = new_n4679_ | new_n6948_;
  assign new_n4681_ = new_n7234_ & new_n6919_;
  assign new_n4682_ = new_n7238_ & new_n6938_;
  assign new_n4683_ = new_n4682_ | new_n6957_;
  assign new_n4684_ = new_n4683_ | new_n4681_;
  assign new_n4685_ = new_n4684_ & new_n4680_;
  assign new_n4686_ = new_n7233_ & new_n7016_;
  assign new_n4687_ = new_n7237_ & new_n7035_;
  assign new_n4688_ = new_n4687_ | new_n7048_;
  assign new_n4689_ = new_n4688_ | new_n4686_;
  assign new_n4690_ = new_n7016_ & new_n7240_;
  assign new_n4691_ = new_n7035_ & new_n7241_;
  assign new_n4692_ = new_n4691_ | new_n7059_;
  assign new_n4693_ = new_n4692_ | new_n4690_;
  assign new_n4694_ = new_n4693_ & new_n7071_;
  assign new_n4695_ = new_n4694_ & new_n4689_;
  assign new_n4696_ = new_n7223_ & new_n7019_;
  assign new_n4697_ = new_n7227_ & new_n7038_;
  assign new_n4698_ = new_n4697_ | new_n7050_;
  assign new_n4699_ = new_n4698_ | new_n4696_;
  assign new_n4700_ = new_n7019_ & new_n7242_;
  assign new_n4701_ = new_n7038_ & new_n7243_;
  assign new_n4702_ = new_n4701_ | new_n7061_;
  assign new_n4703_ = new_n4702_ | new_n4700_;
  assign new_n4704_ = new_n4703_ & new_n7074_;
  assign new_n4705_ = new_n4704_ & new_n4699_;
  assign new_n4706_ = new_n7213_ & new_n7020_;
  assign new_n4707_ = new_n7217_ & new_n7039_;
  assign new_n4708_ = new_n4707_ | new_n7050_;
  assign new_n4709_ = new_n4708_ | new_n4706_;
  assign new_n4710_ = new_n7020_ & new_n7244_;
  assign new_n4711_ = new_n7039_ & new_n7245_;
  assign new_n4712_ = new_n4711_ | new_n7061_;
  assign new_n4713_ = new_n4712_ | new_n4710_;
  assign new_n4714_ = new_n4713_ & new_n7074_;
  assign new_n4715_ = new_n4714_ & new_n4709_;
  assign new_n4716_ = new_n7022_ & new_n7246_;
  assign new_n4717_ = new_n7041_ & new_n7247_;
  assign new_n4718_ = new_n4717_ | new_n4716_;
  assign new_n4719_ = new_n4718_ & new_n7051_;
  assign new_n4720_ = new_n7203_ & new_n7022_;
  assign new_n4721_ = new_n7207_ & new_n7041_;
  assign new_n4722_ = new_n4721_ | new_n4720_;
  assign new_n4723_ = new_n4722_ & new_n7062_;
  assign new_n4724_ = new_n4723_ | new_n4719_;
  assign new_n4725_ = new_n4724_ & new_n7075_;
  assign new_n4726_ = new_n7090_ & new_n7240_;
  assign new_n4727_ = new_n7109_ & new_n7241_;
  assign new_n4728_ = new_n4727_ | new_n4726_;
  assign new_n4729_ = new_n4728_ & new_n7122_;
  assign new_n4730_ = new_n7235_ | new_n7109_;
  assign new_n4731_ = new_n7239_ | new_n7090_;
  assign new_n4732_ = new_n4731_ & new_n7131_;
  assign new_n4733_ = new_n4732_ & new_n4730_;
  assign new_n4734_ = new_n4733_ | new_n4729_;
  assign new_n4735_ = new_n4734_ & new_n7075_;
  assign new_n4736_ = new_n7225_ & new_n7093_;
  assign new_n4737_ = new_n7229_ & new_n7112_;
  assign new_n4738_ = new_n4737_ | new_n7124_;
  assign new_n4739_ = new_n4738_ | new_n4736_;
  assign new_n4740_ = new_n7093_ & new_n7242_;
  assign new_n4741_ = new_n7112_ & new_n7243_;
  assign new_n4742_ = new_n4741_ | new_n7133_;
  assign new_n4743_ = new_n4742_ | new_n4740_;
  assign new_n4744_ = new_n4743_ & new_n7077_;
  assign new_n4745_ = new_n4744_ & new_n4739_;
  assign new_n4746_ = new_n7215_ & new_n7094_;
  assign new_n4747_ = new_n7219_ & new_n7113_;
  assign new_n4748_ = new_n4747_ | new_n7124_;
  assign new_n4749_ = new_n4748_ | new_n4746_;
  assign new_n4750_ = new_n7094_ & new_n7244_;
  assign new_n4751_ = new_n7113_ & new_n7245_;
  assign new_n4752_ = new_n4751_ | new_n7133_;
  assign new_n4753_ = new_n4752_ | new_n4750_;
  assign new_n4754_ = new_n4753_ & new_n7077_;
  assign new_n4755_ = new_n4754_ & new_n4749_;
  assign new_n4756_ = new_n7205_ & new_n7096_;
  assign new_n4757_ = new_n7209_ & new_n7115_;
  assign new_n4758_ = new_n4757_ | new_n7125_;
  assign new_n4759_ = new_n4758_ | new_n4756_;
  assign new_n4760_ = new_n7096_ & new_n7246_;
  assign new_n4761_ = new_n7115_ & new_n7247_;
  assign new_n4762_ = new_n4761_ | new_n7134_;
  assign new_n4763_ = new_n4762_ | new_n4760_;
  assign new_n4764_ = new_n4763_ & new_n7078_;
  assign new_n4765_ = new_n4764_ & new_n4759_;
  assign new_n4766_ = new_n3811_ | new_n3796_;
  assign new_n4767_ = new_n6827_ | new_n6831_;
  assign new_n4768_ = new_n7248_ | new_n2786_;
  assign new_n4769_ = new_n4768_ & new_n7249_;
  assign new_n4770_ = new_n3907_ & new_n6831_;
  assign new_n4771_ = new_n3874_ | new_n6805_;
  assign new_n4772_ = new_n4771_ | new_n4770_;
  assign new_n4773_ = new_n7248_ | new_n2772_;
  assign new_n4774_ = new_n4773_ & new_n7250_;
  assign new_n4775_ = new_n6855_ & new_n7251_;
  assign new_n4776_ = new_n6878_ & new_n7252_;
  assign new_n4777_ = new_n4776_ | new_n4775_;
  assign new_n4778_ = new_n4777_ & new_n6898_;
  assign new_n4779_ = new_n6828_ | new_n2695_;
  assign new_n4780_ = new_n4779_ & new_n7250_;
  assign new_n4781_ = new_n7254_ | new_n6878_;
  assign new_n4782_ = new_n6828_ | new_n2687_;
  assign new_n4783_ = new_n4782_ & new_n7249_;
  assign new_n4784_ = new_n7257_ | new_n6855_;
  assign new_n4785_ = new_n4784_ & new_n6887_;
  assign new_n4786_ = new_n4785_ & new_n4781_;
  assign new_n4787_ = new_n4786_ | new_n4778_;
  assign new_n4788_ = new_n6920_ & new_n7251_;
  assign new_n4789_ = new_n6939_ & new_n7252_;
  assign new_n4790_ = new_n4789_ | new_n4788_;
  assign new_n4791_ = new_n4790_ & new_n6957_;
  assign new_n4792_ = new_n7254_ | new_n6939_;
  assign new_n4793_ = new_n7257_ | new_n6920_;
  assign new_n4794_ = new_n4793_ & new_n6948_;
  assign new_n4795_ = new_n4794_ & new_n4792_;
  assign new_n4796_ = new_n4795_ | new_n4791_;
  assign new_n4797_ = new_n7255_ | new_n7042_;
  assign new_n4798_ = new_n7258_ | new_n7023_;
  assign new_n4799_ = new_n4798_ & new_n7062_;
  assign new_n4800_ = new_n4799_ & new_n4797_;
  assign new_n4801_ = new_n7042_ | new_n7259_;
  assign new_n4802_ = new_n7023_ | new_n7260_;
  assign new_n4803_ = new_n4802_ & new_n7051_;
  assign new_n4804_ = new_n4803_ & new_n4801_;
  assign new_n4805_ = new_n4804_ | new_n7181_;
  assign new_n4806_ = new_n4805_ | new_n4800_;
  assign new_n4807_ = new_n7116_ | new_n7259_;
  assign new_n4808_ = new_n7097_ | new_n7260_;
  assign new_n4809_ = new_n4808_ & new_n4807_;
  assign new_n4810_ = new_n4809_ | new_n7134_;
  assign new_n4811_ = new_n7255_ & new_n7097_;
  assign new_n4812_ = new_n7258_ & new_n7116_;
  assign new_n4813_ = new_n4812_ | new_n7125_;
  assign new_n4814_ = new_n4813_ | new_n4811_;
  assign new_n4815_ = new_n4814_ & new_n4810_;
  assign new_n4816_ = new_n4815_ | new_n7181_;
  assign new_n4817_ = new_n7261_ & new_n7263_;
  assign new_n4818_ = new_n7266_ | new_n7268_;
  assign new_n4819_ = new_n7266_ & new_n7268_;
  assign new_n4820_ = new_n7261_ | new_n7263_;
  assign new_n4821_ = new_n4820_ & new_n7269_;
  assign new_n4822_ = new_n4819_ | new_n4817_;
  assign new_n4823_ = new_n7270_ | new_n7273_;
  assign new_n4824_ = new_n3600_ & new_n7276_;
  assign new_n4825_ = new_n4824_ | new_n3566_;
  assign new_n4826_ = new_n7278_ & new_n7279_;
  assign new_n4827_ = new_n3913_ & new_n3709_;
  assign new_n4828_ = new_n3912_ | new_n3708_;
  assign new_n4829_ = new_n7280_ & new_n3935_;
  assign new_n4830_ = new_n7282_ | new_n3934_;
  assign new_n4831_ = new_n4035_ & new_n4033_;
  assign new_n4832_ = new_n4034_ | new_n4032_;
  assign new_n4833_ = new_n4039_ & new_n4037_;
  assign new_n4834_ = new_n4038_ | new_n4036_;
  assign new_n4835_ = new_n7283_ & new_n4045_;
  assign new_n4836_ = new_n7284_ | new_n4044_;
  assign new_n4837_ = new_n4055_ & new_n7283_;
  assign new_n4838_ = new_n4054_ | new_n7284_;
  assign new_n4839_ = new_n4080_ & new_n4079_;
  assign new_n4840_ = new_n4081_ | new_n7285_;
  assign new_n4841_ = new_n7286_ & new_n7288_;
  assign new_n4842_ = new_n4089_ | new_n7289_;
  assign new_n4843_ = new_n7291_ & new_n7293_;
  assign new_n4844_ = new_n7294_ | new_n7295_;
  assign new_n4845_ = new_n3560_ & new_n7299_;
  assign new_n4846_ = new_n3561_ & new_n7310_;
  assign new_n4847_ = new_n4846_ | new_n4845_;
  assign new_n4848_ = new_n7320_ & new_n7324_;
  assign new_n4849_ = new_n7327_ | new_n7329_;
  assign new_n4850_ = new_n4058_ & new_n7329_;
  assign new_n4851_ = new_n4059_ | new_n7324_;
  assign new_n4852_ = new_n4851_ & new_n4849_;
  assign new_n4853_ = new_n4850_ | new_n4848_;
  assign new_n4854_ = new_n7330_ & new_n3765_;
  assign new_n4855_ = new_n3949_ | new_n7331_;
  assign new_n4856_ = new_n7333_ & new_n4026_;
  assign new_n4857_ = new_n7336_ | new_n4027_;
  assign new_n4858_ = new_n4857_ & new_n7337_;
  assign new_n4859_ = new_n4856_ | new_n7338_;
  assign new_n4860_ = new_n7339_ & new_n7341_;
  assign new_n4861_ = new_n7343_ | new_n7345_;
  assign new_n4862_ = new_n4861_ & new_n7280_;
  assign new_n4863_ = new_n4860_ | new_n7282_;
  assign new_n4864_ = new_n7347_ & new_n7350_;
  assign new_n4865_ = new_n7352_ | new_n7354_;
  assign new_n4866_ = new_n7352_ & new_n7354_;
  assign new_n4867_ = new_n7347_ | new_n7350_;
  assign new_n4868_ = new_n4867_ & new_n7356_;
  assign new_n4869_ = new_n4866_ | new_n7357_;
  assign new_n4870_ = new_n4129_ & new_n4127_;
  assign new_n4871_ = new_n4128_ | new_n4126_;
  assign new_n4872_ = new_n4133_ & new_n4131_;
  assign new_n4873_ = new_n4132_ | new_n4130_;
  assign new_n4874_ = new_n4137_ & new_n4135_;
  assign new_n4875_ = new_n4136_ | new_n4134_;
  assign new_n4876_ = new_n7358_ | new_n3546_;
  assign new_n4877_ = new_n7359_ & new_n7360_;
  assign new_n4878_ = new_n7362_ & new_n7365_;
  assign new_n4879_ = new_n7367_ | new_n7368_;
  assign new_n4880_ = new_n7370_ & new_n2558_;
  assign new_n4881_ = new_n3591_ & new_n2559_;
  assign new_n4882_ = new_n4881_ | new_n4880_;
  assign new_n4883_ = new_n7372_ & new_n7299_;
  assign new_n4884_ = new_n7375_ & new_n7380_;
  assign new_n4885_ = new_n4884_ | new_n4883_;
  assign new_n4886_ = new_n4885_ & new_n3558_;
  assign new_n4887_ = new_n7375_ & new_n7390_;
  assign new_n4888_ = new_n7372_ & new_n7310_;
  assign new_n4889_ = new_n4888_ | new_n4887_;
  assign new_n4890_ = new_n4889_ & new_n3559_;
  assign new_n4891_ = new_n4890_ | new_n4886_;
  assign new_n4892_ = new_n7398_ & new_n7300_;
  assign new_n4893_ = new_n7400_ & new_n7380_;
  assign new_n4894_ = new_n4893_ | new_n4892_;
  assign new_n4895_ = new_n4894_ & new_n3484_;
  assign new_n4896_ = new_n7400_ & new_n7390_;
  assign new_n4897_ = new_n7398_ & new_n7311_;
  assign new_n4898_ = new_n4897_ | new_n4896_;
  assign new_n4899_ = new_n4898_ & new_n3485_;
  assign new_n4900_ = new_n4899_ | new_n4895_;
  assign new_n4901_ = new_n7402_ & new_n7300_;
  assign new_n4902_ = new_n7404_ & new_n7381_;
  assign new_n4903_ = new_n4902_ | new_n4901_;
  assign new_n4904_ = new_n4903_ & new_n3612_;
  assign new_n4905_ = new_n7404_ & new_n7391_;
  assign new_n4906_ = new_n7402_ & new_n7311_;
  assign new_n4907_ = new_n4906_ | new_n4905_;
  assign new_n4908_ = new_n4907_ & new_n3613_;
  assign new_n4909_ = new_n4908_ | new_n4904_;
  assign new_n4910_ = new_n7406_ & new_n7409_;
  assign new_n4911_ = new_n7411_ | new_n7413_;
  assign new_n4912_ = new_n7411_ & new_n7413_;
  assign new_n4913_ = new_n7406_ | new_n7409_;
  assign new_n4914_ = new_n4913_ & new_n4911_;
  assign new_n4915_ = new_n4912_ | new_n7415_;
  assign new_n4916_ = new_n7416_ & new_n7420_;
  assign new_n4917_ = new_n4117_ | new_n7429_;
  assign new_n4918_ = new_n4118_ & new_n7429_;
  assign new_n4919_ = new_n4119_ | new_n7420_;
  assign new_n4920_ = new_n4919_ & new_n4917_;
  assign new_n4921_ = new_n4918_ | new_n4916_;
  assign new_n4922_ = new_n7435_ & new_n7437_;
  assign new_n4923_ = new_n4872_ | new_n4113_;
  assign new_n4924_ = new_n7435_ | new_n7437_;
  assign new_n4925_ = new_n7439_ & new_n7441_;
  assign new_n4926_ = new_n4870_ | new_n4115_;
  assign new_n4927_ = new_n7445_ & new_n7453_;
  assign new_n4928_ = new_n7457_ | new_n4121_;
  assign new_n4929_ = new_n7457_ & new_n4122_;
  assign new_n4930_ = new_n7445_ | new_n4123_;
  assign new_n4931_ = new_n4930_ & new_n4928_;
  assign new_n4932_ = new_n4929_ | new_n4927_;
  assign new_n4933_ = new_n7362_ | new_n7365_;
  assign new_n4934_ = new_n7464_ & new_n7333_;
  assign new_n4935_ = new_n4842_ | new_n7336_;
  assign new_n4936_ = new_n7288_ & new_n7338_;
  assign new_n4937_ = new_n7289_ | new_n7337_;
  assign new_n4938_ = new_n4937_ & new_n3991_;
  assign new_n4939_ = new_n4936_ | new_n3990_;
  assign new_n4940_ = new_n4938_ & new_n4935_;
  assign new_n4941_ = new_n4939_ | new_n4934_;
  assign new_n4942_ = new_n7465_ & new_n7467_;
  assign new_n4943_ = new_n7468_ | new_n7469_;
  assign new_n4944_ = new_n7470_ & new_n7356_;
  assign new_n4945_ = new_n7471_ | new_n7357_;
  assign new_n4946_ = new_n7472_ & new_n7421_;
  assign new_n4947_ = new_n4099_ | new_n7428_;
  assign new_n4948_ = new_n4100_ & new_n7430_;
  assign new_n4949_ = new_n4101_ | new_n7421_;
  assign new_n4950_ = new_n4949_ & new_n4947_;
  assign new_n4951_ = new_n4948_ | new_n4946_;
  assign new_n4952_ = new_n7473_ & new_n7422_;
  assign new_n4953_ = new_n4103_ | new_n7430_;
  assign new_n4954_ = new_n4104_ & new_n7432_;
  assign new_n4955_ = new_n4105_ | new_n7422_;
  assign new_n4956_ = new_n4955_ & new_n4953_;
  assign new_n4957_ = new_n4954_ | new_n4952_;
  assign new_n4958_ = new_n4068_ & new_n4047_;
  assign new_n4959_ = new_n4069_ | new_n4046_;
  assign new_n4960_ = new_n7474_ & new_n7476_;
  assign new_n4961_ = new_n7477_ | new_n7479_;
  assign new_n4962_ = new_n7477_ & new_n7479_;
  assign new_n4963_ = new_n7474_ | new_n7476_;
  assign new_n4964_ = new_n4963_ & new_n4961_;
  assign new_n4965_ = new_n4962_ | new_n4960_;
  assign new_n4966_ = new_n4964_ & new_n4855_;
  assign new_n4967_ = new_n4965_ & new_n7482_;
  assign new_n4968_ = new_n4967_ | new_n7483_;
  assign new_n4969_ = new_n7446_ & new_n7484_;
  assign new_n4970_ = new_n7458_ & new_n4108_;
  assign new_n4971_ = new_n4970_ | new_n4969_;
  assign new_n4972_ = new_n7468_ & new_n7469_;
  assign new_n4973_ = new_n7465_ | new_n7467_;
  assign new_n4974_ = new_n4973_ & new_n7470_;
  assign new_n4975_ = new_n4972_ | new_n7471_;
  assign new_n4976_ = new_n7486_ & new_n7488_;
  assign new_n4977_ = new_n4920_ | new_n4095_;
  assign new_n4978_ = new_n7490_ & new_n7492_;
  assign new_n4979_ = new_n4874_ | new_n4111_;
  assign new_n4980_ = new_n7490_ | new_n7492_;
  assign new_n4981_ = new_n4980_ & new_n4979_;
  assign new_n4982_ = new_n7494_ & new_n4923_;
  assign new_n4983_ = new_n7439_ | new_n7441_;
  assign new_n4984_ = new_n4983_ & new_n4926_;
  assign new_n4985_ = new_n7446_ & new_n7496_;
  assign new_n4986_ = new_n7458_ | new_n4091_;
  assign new_n4987_ = new_n7460_ & new_n7497_;
  assign new_n4988_ = new_n7448_ | new_n4093_;
  assign new_n4989_ = new_n4988_ & new_n4986_;
  assign new_n4990_ = new_n4987_ | new_n4985_;
  assign new_n4991_ = new_n7499_ & new_n7501_;
  assign new_n4992_ = new_n4956_ | new_n3175_;
  assign new_n4993_ = new_n7503_ & new_n7505_;
  assign new_n4994_ = new_n4950_ | new_n3183_;
  assign new_n4995_ = new_n7507_ & new_n7509_;
  assign new_n4996_ = new_n7511_ & new_n7513_;
  assign new_n4997_ = new_n4931_ | new_n4097_;
  assign new_n4998_ = new_n7511_ | new_n7513_;
  assign new_n4999_ = new_n7514_ & new_n4997_;
  assign new_n5000_ = new_n7516_ & new_n7517_;
  assign new_n5001_ = new_n7521_ & new_n2544_;
  assign new_n5002_ = new_n7521_ & new_n2738_;
  assign new_n5003_ = new_n7522_ & new_n2758_;
  assign new_n5004_ = new_n7531_ | new_n2764_;
  assign new_n5005_ = new_n7531_ | new_n2778_;
  assign new_n5006_ = new_n7522_ & new_n2792_;
  assign new_n5007_ = new_n7524_ & new_n2830_;
  assign new_n5008_ = new_n7532_ | new_n2836_;
  assign new_n5009_ = new_n7532_ | new_n2848_;
  assign new_n5010_ = new_n7542_ & new_n7302_;
  assign new_n5011_ = new_n7544_ & new_n7381_;
  assign new_n5012_ = new_n5011_ | new_n5010_;
  assign new_n5013_ = new_n5012_ & new_n3482_;
  assign new_n5014_ = new_n7544_ & new_n7391_;
  assign new_n5015_ = new_n7542_ & new_n7313_;
  assign new_n5016_ = new_n5015_ | new_n5014_;
  assign new_n5017_ = new_n5016_ & new_n3483_;
  assign new_n5018_ = new_n7534_ & new_n7546_;
  assign new_n5019_ = new_n7534_ | new_n7547_;
  assign new_n5020_ = new_n5019_ & new_n7549_;
  assign new_n5021_ = new_n3609_ & new_n7550_;
  assign new_n5022_ = new_n7552_ | new_n7553_;
  assign new_n5023_ = new_n5022_ & new_n3629_;
  assign new_n5024_ = new_n5021_ | new_n7554_;
  assign new_n5025_ = new_n7555_ & new_n7556_;
  assign new_n5026_ = new_n7557_ | new_n7558_;
  assign new_n5027_ = new_n7557_ & new_n7558_;
  assign new_n5028_ = new_n7555_ | new_n7556_;
  assign new_n5029_ = new_n5028_ & new_n5026_;
  assign new_n5030_ = new_n5027_ | new_n5025_;
  assign new_n5031_ = new_n7559_ & new_n7560_;
  assign new_n5032_ = new_n7561_ | new_n7562_;
  assign new_n5033_ = new_n7561_ & new_n7562_;
  assign new_n5034_ = new_n7559_ | new_n7560_;
  assign new_n5035_ = new_n5034_ & new_n5032_;
  assign new_n5036_ = new_n5033_ | new_n5031_;
  assign new_n5037_ = new_n3734_ & new_n7563_;
  assign new_n5038_ = new_n3735_ | new_n7273_;
  assign new_n5039_ = new_n4015_ & new_n7272_;
  assign new_n5040_ = new_n4014_ | new_n7563_;
  assign new_n5041_ = new_n5040_ & new_n5038_;
  assign new_n5042_ = new_n5039_ | new_n5037_;
  assign new_n5043_ = new_n7564_ & new_n7566_;
  assign new_n5044_ = new_n7567_ | new_n7569_;
  assign new_n5045_ = new_n7567_ & new_n7569_;
  assign new_n5046_ = new_n7564_ | new_n7566_;
  assign new_n5047_ = new_n5046_ & new_n5044_;
  assign new_n5048_ = new_n5045_ | new_n5043_;
  assign new_n5049_ = new_n5047_ & new_n5036_;
  assign new_n5050_ = new_n5048_ & new_n5035_;
  assign new_n5051_ = new_n5050_ | new_n5049_;
  assign new_n5052_ = new_n5051_ & new_n7546_;
  assign new_n5053_ = new_n7570_ | new_n7524_;
  assign new_n5054_ = new_n7571_ | new_n7523_;
  assign new_n5055_ = new_n3923_ & new_n7535_;
  assign new_n5056_ = new_n3920_ & new_n7535_;
  assign new_n5057_ = new_n3915_ & new_n7538_;
  assign new_n5058_ = new_n7572_ | new_n7526_;
  assign new_n5059_ = new_n4013_ & new_n4011_;
  assign new_n5060_ = new_n4012_ | new_n4010_;
  assign new_n5061_ = new_n4009_ & new_n4007_;
  assign new_n5062_ = new_n4008_ | new_n4006_;
  assign new_n5063_ = new_n7573_ & new_n7574_;
  assign new_n5064_ = new_n7575_ | new_n7576_;
  assign new_n5065_ = new_n7575_ & new_n7576_;
  assign new_n5066_ = new_n7573_ | new_n7574_;
  assign new_n5067_ = new_n5066_ & new_n5064_;
  assign new_n5068_ = new_n5065_ | new_n5063_;
  assign new_n5069_ = new_n4004_ & new_n4003_;
  assign new_n5070_ = new_n4005_ | new_n7577_;
  assign new_n5071_ = new_n4001_ & new_n3999_;
  assign new_n5072_ = new_n4000_ | new_n7578_;
  assign new_n5073_ = new_n7579_ & new_n7580_;
  assign new_n5074_ = new_n7581_ | new_n7582_;
  assign new_n5075_ = new_n7581_ & new_n7582_;
  assign new_n5076_ = new_n7579_ | new_n7580_;
  assign new_n5077_ = new_n5076_ & new_n5074_;
  assign new_n5078_ = new_n5075_ | new_n5073_;
  assign new_n5079_ = new_n5077_ & new_n5067_;
  assign new_n5080_ = new_n5078_ & new_n5068_;
  assign new_n5081_ = new_n5080_ | new_n7545_;
  assign new_n5082_ = new_n5081_ | new_n5079_;
  assign new_n5083_ = new_n5082_ & new_n7538_;
  assign new_n5084_ = new_n3528_ & new_n3509_;
  assign new_n5085_ = new_n3529_ & new_n3508_;
  assign new_n5086_ = new_n7584_ & new_n7276_;
  assign new_n5087_ = new_n7587_ | new_n7588_;
  assign new_n5088_ = new_n5087_ & new_n7590_;
  assign new_n5089_ = new_n5086_ | new_n7594_;
  assign new_n5090_ = new_n7598_ & new_n3533_;
  assign new_n5091_ = new_n7602_ & new_n3532_;
  assign new_n5092_ = new_n7604_ & new_n3580_;
  assign new_n5093_ = new_n7606_ & new_n3551_;
  assign new_n5094_ = new_n5093_ | new_n5092_;
  assign new_n5095_ = new_n7607_ | new_n7274_;
  assign new_n5096_ = new_n7607_ & new_n7274_;
  assign new_n5097_ = new_n7278_ | new_n7279_;
  assign new_n5098_ = new_n7608_ | new_n3586_;
  assign new_n5099_ = new_n3474_ & new_n7610_;
  assign new_n5100_ = new_n3475_ & new_n3154_;
  assign new_n5101_ = new_n5100_ | new_n5099_;
  assign new_n5102_ = new_n7611_ | new_n7370_;
  assign new_n5103_ = new_n7611_ & new_n7369_;
  assign new_n5104_ = new_n7359_ | new_n7360_;
  assign new_n5105_ = new_n7612_ & new_n7552_;
  assign new_n5106_ = new_n7612_ | new_n7551_;
  assign new_n5107_ = new_n7613_ | new_n7606_;
  assign new_n5108_ = new_n5107_ & new_n3585_;
  assign new_n5109_ = new_n7614_ & new_n7264_;
  assign new_n5110_ = new_n7614_ | new_n7264_;
  assign new_n5111_ = new_n7615_ | new_n7568_;
  assign new_n5112_ = new_n7616_ & new_n7277_;
  assign new_n5113_ = new_n3583_ | new_n7588_;
  assign new_n5114_ = new_n7616_ | new_n7277_;
  assign new_n5115_ = new_n5114_ & new_n7617_;
  assign new_n5116_ = new_n7460_ & new_n3127_;
  assign new_n5117_ = new_n7448_ | new_n7618_;
  assign new_n5118_ = new_n7526_ & new_n2732_;
  assign new_n5119_ = new_n3917_ & new_n7539_;
  assign new_n5120_ = new_n5119_ | new_n5118_;
  assign new_n5121_ = new_n7527_ & new_n2752_;
  assign new_n5122_ = new_n7620_ & new_n7539_;
  assign new_n5123_ = new_n5122_ | new_n5121_;
  assign new_n5124_ = new_n7540_ | new_n2843_;
  assign new_n5125_ = new_n7621_ | new_n7527_;
  assign new_n5126_ = new_n5125_ & new_n5124_;
  assign new_n5127_ = new_n3536_ | new_n7623_;
  assign new_n5128_ = new_n3537_ | new_n7625_;
  assign new_n5129_ = new_n5128_ & new_n5127_;
  assign new_n5130_ = new_n7397_ & new_n7627_;
  assign new_n5131_ = new_n7399_ & new_n7629_;
  assign new_n5132_ = new_n5131_ | new_n5130_;
  assign new_n5133_ = new_n7631_ & new_n7541_;
  assign new_n5134_ = new_n7633_ & new_n7543_;
  assign new_n5135_ = new_n5134_ | new_n5133_;
  assign new_n5136_ = new_n7635_ & new_n7302_;
  assign new_n5137_ = new_n7638_ & new_n7383_;
  assign new_n5138_ = new_n5137_ | new_n5136_;
  assign new_n5139_ = new_n5138_ & new_n3500_;
  assign new_n5140_ = new_n7638_ & new_n7393_;
  assign new_n5141_ = new_n7635_ & new_n7313_;
  assign new_n5142_ = new_n5141_ | new_n5140_;
  assign new_n5143_ = new_n5142_ & new_n3501_;
  assign new_n5144_ = new_n5143_ | new_n5139_;
  assign new_n5145_ = new_n7633_ & new_n7303_;
  assign new_n5146_ = new_n7631_ & new_n7383_;
  assign new_n5147_ = new_n5146_ | new_n5145_;
  assign new_n5148_ = new_n5147_ & new_n3516_;
  assign new_n5149_ = new_n7630_ & new_n7393_;
  assign new_n5150_ = new_n7632_ & new_n7314_;
  assign new_n5151_ = new_n5150_ | new_n5149_;
  assign new_n5152_ = new_n5151_ & new_n3517_;
  assign new_n5153_ = new_n5152_ | new_n5148_;
  assign new_n5154_ = new_n7641_ & new_n7303_;
  assign new_n5155_ = new_n7644_ & new_n7382_;
  assign new_n5156_ = new_n5155_ | new_n5154_;
  assign new_n5157_ = new_n5156_ & new_n3630_;
  assign new_n5158_ = new_n7644_ & new_n7392_;
  assign new_n5159_ = new_n7641_ & new_n7314_;
  assign new_n5160_ = new_n5159_ | new_n5158_;
  assign new_n5161_ = new_n5160_ & new_n3631_;
  assign new_n5162_ = new_n5161_ | new_n5157_;
  assign new_n5163_ = new_n7625_ & new_n7305_;
  assign new_n5164_ = new_n7623_ & new_n7385_;
  assign new_n5165_ = new_n5164_ | new_n5163_;
  assign new_n5166_ = new_n5165_ & new_n3518_;
  assign new_n5167_ = new_n7622_ & new_n7395_;
  assign new_n5168_ = new_n7624_ & new_n7316_;
  assign new_n5169_ = new_n5168_ | new_n5167_;
  assign new_n5170_ = new_n5169_ & new_n3519_;
  assign new_n5171_ = new_n5170_ | new_n5166_;
  assign new_n5172_ = new_n7629_ & new_n7305_;
  assign new_n5173_ = new_n7627_ & new_n7385_;
  assign new_n5174_ = new_n5173_ | new_n5172_;
  assign new_n5175_ = new_n5174_ & new_n3486_;
  assign new_n5176_ = new_n7626_ & new_n7395_;
  assign new_n5177_ = new_n7628_ & new_n7316_;
  assign new_n5178_ = new_n5177_ | new_n5176_;
  assign new_n5179_ = new_n5178_ & new_n3487_;
  assign new_n5180_ = new_n5179_ | new_n5175_;
  assign new_n5181_ = new_n7647_ & new_n7306_;
  assign new_n5182_ = new_n7649_ & new_n7386_;
  assign new_n5183_ = new_n5182_ | new_n5181_;
  assign new_n5184_ = new_n5183_ & new_n3562_;
  assign new_n5185_ = new_n7649_ & new_n7396_;
  assign new_n5186_ = new_n7647_ & new_n7317_;
  assign new_n5187_ = new_n5186_ | new_n5185_;
  assign new_n5188_ = new_n5187_ & new_n3563_;
  assign new_n5189_ = new_n5188_ | new_n5184_;
  assign new_n5190_ = new_n7651_ & new_n7306_;
  assign new_n5191_ = new_n7653_ & new_n7386_;
  assign new_n5192_ = new_n5191_ | new_n5190_;
  assign new_n5193_ = new_n5192_ & new_n3544_;
  assign new_n5194_ = new_n7653_ & new_n7396_;
  assign new_n5195_ = new_n7651_ & new_n7317_;
  assign new_n5196_ = new_n5195_ | new_n5194_;
  assign new_n5197_ = new_n5196_ & new_n3545_;
  assign new_n5198_ = new_n5197_ | new_n5193_;
  assign new_n5199_ = new_n7654_ & new_n7655_;
  assign new_n5200_ = new_n7656_ | new_n7657_;
  assign new_n5201_ = new_n7656_ & new_n7657_;
  assign new_n5202_ = new_n7654_ | new_n7655_;
  assign new_n5203_ = new_n5202_ & new_n5200_;
  assign new_n5204_ = new_n5201_ | new_n5199_;
  assign new_n5205_ = new_n7620_ & new_n7658_;
  assign new_n5206_ = new_n7660_ | new_n7661_;
  assign new_n5207_ = new_n7660_ & new_n7661_;
  assign new_n5208_ = new_n7619_ | new_n7658_;
  assign new_n5209_ = new_n5208_ & new_n5206_;
  assign new_n5210_ = new_n5207_ | new_n5205_;
  assign new_n5211_ = new_n7662_ & new_n7663_;
  assign new_n5212_ = new_n7664_ | new_n7665_;
  assign new_n5213_ = new_n7664_ & new_n7665_;
  assign new_n5214_ = new_n7662_ | new_n7663_;
  assign new_n5215_ = new_n5214_ & new_n5212_;
  assign new_n5216_ = new_n5213_ | new_n5211_;
  assign new_n5217_ = new_n7666_ & new_n7667_;
  assign new_n5218_ = new_n7668_ | new_n7669_;
  assign new_n5219_ = new_n7668_ & new_n7669_;
  assign new_n5220_ = new_n7666_ | new_n7667_;
  assign new_n5221_ = new_n5220_ & new_n5218_;
  assign new_n5222_ = new_n5219_ | new_n5217_;
  assign new_n5223_ = new_n7670_ & new_n7671_;
  assign new_n5224_ = new_n7672_ | new_n7673_;
  assign new_n5225_ = new_n7672_ & new_n7673_;
  assign new_n5226_ = new_n7670_ | new_n7671_;
  assign new_n5227_ = new_n5226_ & new_n5224_;
  assign new_n5228_ = new_n5225_ | new_n5223_;
  assign new_n5229_ = new_n7674_ & new_n7675_;
  assign new_n5230_ = new_n7676_ | new_n7677_;
  assign new_n5231_ = new_n7676_ & new_n7677_;
  assign new_n5232_ = new_n7674_ | new_n7675_;
  assign new_n5233_ = new_n5232_ & new_n5230_;
  assign new_n5234_ = new_n5231_ | new_n5229_;
  assign new_n5235_ = new_n5234_ | new_n5215_;
  assign new_n5236_ = new_n5233_ | new_n5216_;
  assign new_n5237_ = new_n5236_ & new_n7549_;
  assign new_n5238_ = new_n5237_ & new_n5235_;
  assign new_n5239_ = new_n3636_ & new_n3493_;
  assign new_n5240_ = new_n3637_ & new_n3492_;
  assign new_n5241_ = new_n5240_ | new_n5239_;
  assign new_n5242_ = new_n7602_ | new_n3505_;
  assign new_n5243_ = new_n7598_ | new_n3502_;
  assign new_n5244_ = new_n5243_ & new_n5242_;
  assign new_n5245_ = new_n7617_ & new_n3523_;
  assign new_n5246_ = new_n5112_ | new_n3522_;
  assign new_n5247_ = new_n5246_ | new_n3530_;
  assign new_n5248_ = new_n5245_ | new_n3531_;
  assign new_n5249_ = new_n5248_ & new_n5247_;
  assign new_n5250_ = new_n7678_ & new_n7680_;
  assign new_n5251_ = new_n7681_ | new_n7683_;
  assign new_n5252_ = new_n7681_ & new_n3104_;
  assign new_n5253_ = new_n7678_ | new_n3105_;
  assign new_n5254_ = new_n5253_ & new_n5251_;
  assign new_n5255_ = new_n5252_ | new_n5250_;
  assign new_n5256_ = new_n5255_ | new_n3588_;
  assign new_n5257_ = new_n5254_ | new_n3589_;
  assign new_n5258_ = new_n5257_ & new_n5256_;
  assign new_n5259_ = new_n7597_ & new_n3592_;
  assign new_n5260_ = new_n7601_ & new_n7684_;
  assign new_n5261_ = new_n5260_ | new_n5259_;
  assign new_n5262_ = new_n3649_ | new_n7550_;
  assign new_n5263_ = new_n3648_ | new_n7553_;
  assign new_n5264_ = new_n5263_ & new_n5262_;
  assign new_n5265_ = new_n7599_ & new_n3624_;
  assign new_n5266_ = new_n7603_ | new_n3625_;
  assign new_n5267_ = new_n7603_ & new_n3622_;
  assign new_n5268_ = new_n7599_ | new_n3623_;
  assign new_n5269_ = new_n5268_ & new_n5266_;
  assign new_n5270_ = new_n5267_ | new_n5265_;
  assign new_n5271_ = new_n5269_ & new_n7685_;
  assign new_n5272_ = new_n5270_ & new_n3627_;
  assign new_n5273_ = new_n5272_ | new_n5271_;
  assign new_n5274_ = new_n7604_ & new_n7270_;
  assign new_n5275_ = new_n7605_ & new_n3646_;
  assign new_n5276_ = new_n5275_ | new_n5274_;
  assign new_n5277_ = new_n3481_ & new_n3472_;
  assign new_n5278_ = new_n3480_ & new_n3473_;
  assign new_n5279_ = new_n5278_ | new_n5277_;
  assign new_n5280_ = new_n3679_ | new_n3576_;
  assign new_n5281_ = new_n7686_ | new_n3577_;
  assign new_n5282_ = new_n5281_ & new_n5280_;
  assign new_n5283_ = new_n7687_ & new_n7688_;
  assign new_n5284_ = new_n7687_ | new_n7688_;
  assign new_n5285_ = new_n7689_ & new_n7690_;
  assign new_n5286_ = new_n7691_ | new_n7610_;
  assign new_n5287_ = new_n7691_ & new_n7609_;
  assign new_n5288_ = new_n7689_ | new_n7690_;
  assign new_n5289_ = new_n5288_ & new_n5286_;
  assign new_n5290_ = new_n5287_ | new_n5285_;
  assign new_n5291_ = new_n5289_ & new_n7403_;
  assign new_n5292_ = new_n5290_ & new_n7401_;
  assign new_n5293_ = new_n5292_ | new_n5291_;
  assign new_n5294_ = new_n7646_ | new_n7652_;
  assign new_n5295_ = new_n7648_ | new_n7650_;
  assign new_n5296_ = new_n5295_ & new_n5294_;
  assign new_n5297_ = new_n7692_ & new_n7693_;
  assign new_n5298_ = new_n7692_ | new_n7693_;
  assign new_n5299_ = new_n3620_ & new_n3565_;
  assign new_n5300_ = new_n3621_ & new_n3564_;
  assign new_n5301_ = new_n5300_ | new_n5299_;
  assign new_n5302_ = new_n3570_ & new_n3553_;
  assign new_n5303_ = new_n3571_ & new_n3552_;
  assign new_n5304_ = new_n5303_ | new_n5302_;
  assign new_n5305_ = new_n7694_ | new_n7695_;
  assign new_n5306_ = new_n7694_ & new_n7695_;
  assign new_n5307_ = new_n7645_ & new_n7373_;
  assign new_n5308_ = new_n7642_ | new_n7376_;
  assign new_n5309_ = new_n7642_ & new_n7376_;
  assign new_n5310_ = new_n7645_ | new_n7373_;
  assign new_n5311_ = new_n5310_ & new_n5308_;
  assign new_n5312_ = new_n5309_ | new_n5307_;
  assign new_n5313_ = new_n7639_ & new_n7683_;
  assign new_n5314_ = new_n7636_ | new_n7680_;
  assign new_n5315_ = new_n7636_ & new_n7679_;
  assign new_n5316_ = new_n7639_ | new_n7682_;
  assign new_n5317_ = new_n5316_ & new_n5314_;
  assign new_n5318_ = new_n5315_ | new_n5313_;
  assign new_n5319_ = new_n5318_ | new_n5312_;
  assign new_n5320_ = new_n5317_ | new_n5311_;
  assign new_n5321_ = new_n5320_ & new_n5319_;
  assign new_n5322_ = new_n3947_ & new_n3944_;
  assign new_n5323_ = new_n3946_ | new_n3945_;
  assign new_n5324_ = new_n3714_ & new_n3683_;
  assign new_n5325_ = new_n3715_ | new_n3682_;
  assign new_n5326_ = new_n7696_ & new_n7697_;
  assign new_n5327_ = new_n7698_ | new_n7699_;
  assign new_n5328_ = new_n7698_ & new_n7699_;
  assign new_n5329_ = new_n7696_ | new_n7697_;
  assign new_n5330_ = new_n5329_ & new_n5327_;
  assign new_n5331_ = new_n5328_ | new_n5326_;
  assign new_n5332_ = new_n5331_ & new_n7701_;
  assign new_n5333_ = new_n5330_ | new_n7704_;
  assign new_n5334_ = new_n3984_ & new_n3983_;
  assign new_n5335_ = new_n3985_ | new_n3982_;
  assign new_n5336_ = new_n3995_ & new_n3992_;
  assign new_n5337_ = new_n3994_ | new_n3993_;
  assign new_n5338_ = new_n7706_ & new_n7707_;
  assign new_n5339_ = new_n7708_ | new_n7709_;
  assign new_n5340_ = new_n7708_ & new_n7709_;
  assign new_n5341_ = new_n7706_ | new_n7707_;
  assign new_n5342_ = new_n5341_ & new_n5339_;
  assign new_n5343_ = new_n5340_ | new_n5338_;
  assign new_n5344_ = new_n5342_ & new_n7704_;
  assign new_n5345_ = new_n5343_ | new_n7701_;
  assign new_n5346_ = new_n5345_ & new_n5333_;
  assign new_n5347_ = new_n5344_ | new_n5332_;
  assign new_n5348_ = new_n3952_ & new_n3951_;
  assign new_n5349_ = new_n3953_ | new_n3950_;
  assign new_n5350_ = new_n7587_ & new_n7590_;
  assign new_n5351_ = new_n7584_ | new_n7594_;
  assign new_n5352_ = new_n5351_ & new_n7710_;
  assign new_n5353_ = new_n5350_ | new_n7711_;
  assign new_n5354_ = new_n4017_ & new_n7591_;
  assign new_n5355_ = new_n4016_ | new_n7593_;
  assign new_n5356_ = new_n7712_ & new_n7586_;
  assign new_n5357_ = new_n7713_ | new_n7585_;
  assign new_n5358_ = new_n5357_ & new_n5353_;
  assign new_n5359_ = new_n5356_ | new_n5352_;
  assign new_n5360_ = new_n5359_ & new_n7705_;
  assign new_n5361_ = new_n5358_ | new_n7702_;
  assign new_n5362_ = new_n7710_ & new_n7595_;
  assign new_n5363_ = new_n7711_ | new_n7591_;
  assign new_n5364_ = new_n5363_ & new_n7713_;
  assign new_n5365_ = new_n5362_ | new_n7712_;
  assign new_n5366_ = new_n5365_ & new_n7702_;
  assign new_n5367_ = new_n5364_ | new_n7705_;
  assign new_n5368_ = new_n5367_ & new_n5361_;
  assign new_n5369_ = new_n5366_ | new_n5360_;
  assign new_n5370_ = new_n5369_ | new_n5346_;
  assign new_n5371_ = new_n5368_ | new_n5347_;
  assign new_n5372_ = new_n5371_ & new_n5370_;
  assign new_n5373_ = new_n7486_ | new_n7488_;
  assign new_n5374_ = new_n7715_ & new_n7716_;
  assign new_n5375_ = new_n5374_ | new_n4978_;
  assign new_n5376_ = new_n7516_ & new_n7717_;
  assign new_n5377_ = new_n7721_ & new_n7733_;
  assign new_n5378_ = new_n7737_ & new_n7749_;
  assign new_n5379_ = new_n5378_ | new_n5377_;
  assign new_n5380_ = new_n5379_ & new_n3700_;
  assign new_n5381_ = new_n7753_ & new_n7749_;
  assign new_n5382_ = new_n7766_ & new_n7733_;
  assign new_n5383_ = new_n5382_ | new_n5381_;
  assign new_n5384_ = new_n5383_ & new_n3701_;
  assign new_n5385_ = new_n5384_ | new_n5380_;
  assign new_n5386_ = new_n7721_ & new_n7777_;
  assign new_n5387_ = new_n7737_ & new_n7779_;
  assign new_n5388_ = new_n5387_ | new_n5386_;
  assign new_n5389_ = new_n5388_ & new_n3728_;
  assign new_n5390_ = new_n7753_ & new_n7779_;
  assign new_n5391_ = new_n7766_ & new_n7777_;
  assign new_n5392_ = new_n5391_ | new_n5390_;
  assign new_n5393_ = new_n5392_ & new_n3729_;
  assign new_n5394_ = new_n5393_ | new_n5389_;
  assign new_n5395_ = new_n7722_ & new_n3753_;
  assign new_n5396_ = new_n7738_ & new_n7780_;
  assign new_n5397_ = new_n5396_ | new_n5395_;
  assign new_n5398_ = new_n7722_ & new_n3959_;
  assign new_n5399_ = new_n7738_ & new_n7781_;
  assign new_n5400_ = new_n5399_ | new_n5398_;
  assign new_n5401_ = new_n7767_ | new_n7783_;
  assign new_n5402_ = new_n7754_ | new_n3109_;
  assign new_n5403_ = new_n5402_ & new_n5401_;
  assign new_n5404_ = new_n7424_ & new_n7784_;
  assign new_n5405_ = new_n7432_ | new_n3091_;
  assign new_n5406_ = new_n7433_ & new_n3092_;
  assign new_n5407_ = new_n7424_ | new_n3093_;
  assign new_n5408_ = new_n5407_ & new_n5405_;
  assign new_n5409_ = new_n5406_ | new_n5404_;
  assign new_n5410_ = new_n7449_ & new_n7785_;
  assign new_n5411_ = new_n7459_ | new_n3131_;
  assign new_n5412_ = new_n7462_ & new_n7786_;
  assign new_n5413_ = new_n7449_ | new_n3133_;
  assign new_n5414_ = new_n5413_ & new_n5411_;
  assign new_n5415_ = new_n5412_ | new_n5410_;
  assign new_n5416_ = new_n4989_ | new_n3193_;
  assign new_n5417_ = new_n7499_ | new_n7501_;
  assign new_n5418_ = new_n5417_ & new_n4992_;
  assign new_n5419_ = new_n7503_ | new_n7505_;
  assign new_n5420_ = new_n5419_ & new_n4994_;
  assign new_n5421_ = new_n7363_ & new_n7788_;
  assign new_n5422_ = new_n7367_ | new_n7791_;
  assign new_n5423_ = new_n5422_ & new_n4023_;
  assign new_n5424_ = new_n5421_ | new_n7793_;
  assign new_n5425_ = new_n7795_ & new_n7797_;
  assign new_n5426_ = new_n5425_ | new_n7415_;
  assign new_n5427_ = new_n7798_ | new_n7800_;
  assign new_n5428_ = new_n7802_ | new_n7804_;
  assign new_n5429_ = new_n7788_ & new_n7806_;
  assign new_n5430_ = new_n7791_ | new_n7808_;
  assign new_n5431_ = new_n7792_ & new_n7808_;
  assign new_n5432_ = new_n7789_ | new_n7806_;
  assign new_n5433_ = new_n5432_ & new_n5430_;
  assign new_n5434_ = new_n5431_ | new_n5429_;
  assign new_n5435_ = new_n7809_ & new_n7811_;
  assign new_n5436_ = new_n7812_ | new_n7814_;
  assign new_n5437_ = new_n7812_ & new_n7814_;
  assign new_n5438_ = new_n7809_ | new_n7811_;
  assign new_n5439_ = new_n5438_ & new_n5436_;
  assign new_n5440_ = new_n5437_ | new_n5435_;
  assign new_n5441_ = new_n3955_ & new_n3743_;
  assign new_n5442_ = new_n7816_ | new_n7817_;
  assign new_n5443_ = new_n5442_ & new_n7800_;
  assign new_n5444_ = new_n5441_ | new_n7819_;
  assign new_n5445_ = new_n7822_ & new_n7824_;
  assign new_n5446_ = new_n7826_ | new_n7795_;
  assign new_n5447_ = new_n7826_ & new_n7794_;
  assign new_n5448_ = new_n7822_ | new_n7824_;
  assign new_n5449_ = new_n5448_ & new_n5446_;
  assign new_n5450_ = new_n5447_ | new_n5445_;
  assign new_n5451_ = new_n5450_ & new_n5440_;
  assign new_n5452_ = new_n5449_ & new_n5439_;
  assign new_n5453_ = new_n5452_ | new_n5451_;
  assign new_n5454_ = new_n7827_ & new_n7804_;
  assign new_n5455_ = new_n7827_ | new_n7805_;
  assign new_n5456_ = new_n7507_ | new_n7509_;
  assign new_n5457_ = new_n4042_ & new_n4041_;
  assign new_n5458_ = new_n4043_ | new_n4040_;
  assign new_n5459_ = new_n7828_ & new_n7830_;
  assign new_n5460_ = new_n7831_ | new_n7832_;
  assign new_n5461_ = new_n7831_ & new_n7832_;
  assign new_n5462_ = new_n7828_ | new_n7830_;
  assign new_n5463_ = new_n5462_ & new_n5460_;
  assign new_n5464_ = new_n5461_ | new_n5459_;
  assign new_n5465_ = new_n5463_ & new_n7833_;
  assign new_n5466_ = new_n7834_ | new_n7836_;
  assign new_n5467_ = new_n7834_ & new_n7836_;
  assign new_n5468_ = new_n5467_ | new_n7838_;
  assign new_n5469_ = new_n7294_ & new_n7295_;
  assign new_n5470_ = new_n7291_ | new_n7293_;
  assign new_n5471_ = new_n5470_ & new_n4844_;
  assign new_n5472_ = new_n5469_ | new_n7839_;
  assign new_n5473_ = new_n7840_ & new_n7842_;
  assign new_n5474_ = new_n7843_ | new_n7844_;
  assign new_n5475_ = new_n7843_ & new_n7844_;
  assign new_n5476_ = new_n7840_ | new_n7842_;
  assign new_n5477_ = new_n5476_ & new_n5474_;
  assign new_n5478_ = new_n5475_ | new_n5473_;
  assign new_n5479_ = new_n7846_ & new_n7847_;
  assign new_n5480_ = new_n7846_ | new_n7847_;
  assign new_n5481_ = new_n7848_ & new_n4977_;
  assign new_n5482_ = new_n7849_ & new_n7850_;
  assign new_n5483_ = new_n5482_ | new_n4996_;
  assign new_n5484_ = new_n7851_ & new_n7783_;
  assign new_n5485_ = new_n3657_ & new_n7852_;
  assign new_n5486_ = new_n5485_ | new_n5484_;
  assign new_n5487_ = new_n7724_ & new_n7853_;
  assign new_n5488_ = new_n7740_ & new_n7855_;
  assign new_n5489_ = new_n5488_ | new_n5487_;
  assign new_n5490_ = new_n5489_ & new_n7856_;
  assign new_n5491_ = new_n7754_ & new_n7855_;
  assign new_n5492_ = new_n7767_ & new_n7853_;
  assign new_n5493_ = new_n5492_ | new_n5491_;
  assign new_n5494_ = new_n5493_ & new_n3667_;
  assign new_n5495_ = new_n5494_ | new_n5490_;
  assign new_n5496_ = new_n7724_ & new_n7857_;
  assign new_n5497_ = new_n7740_ & new_n7859_;
  assign new_n5498_ = new_n5497_ | new_n5496_;
  assign new_n5499_ = new_n5498_ & new_n7860_;
  assign new_n5500_ = new_n7756_ & new_n7859_;
  assign new_n5501_ = new_n7769_ & new_n7857_;
  assign new_n5502_ = new_n5501_ | new_n5500_;
  assign new_n5503_ = new_n5502_ & new_n3669_;
  assign new_n5504_ = new_n5503_ | new_n5499_;
  assign new_n5505_ = new_n7725_ & new_n7861_;
  assign new_n5506_ = new_n7741_ & new_n7863_;
  assign new_n5507_ = new_n5506_ | new_n5505_;
  assign new_n5508_ = new_n5507_ & new_n7864_;
  assign new_n5509_ = new_n7756_ & new_n7863_;
  assign new_n5510_ = new_n7769_ & new_n7861_;
  assign new_n5511_ = new_n5510_ | new_n5509_;
  assign new_n5512_ = new_n5511_ & new_n3671_;
  assign new_n5513_ = new_n5512_ | new_n5508_;
  assign new_n5514_ = new_n7725_ & new_n7865_;
  assign new_n5515_ = new_n7741_ & new_n7867_;
  assign new_n5516_ = new_n5515_ | new_n5514_;
  assign new_n5517_ = new_n5516_ & new_n7868_;
  assign new_n5518_ = new_n7757_ & new_n7867_;
  assign new_n5519_ = new_n7770_ & new_n7865_;
  assign new_n5520_ = new_n5519_ | new_n5518_;
  assign new_n5521_ = new_n5520_ & new_n3699_;
  assign new_n5522_ = new_n5521_ | new_n5517_;
  assign new_n5523_ = new_n7728_ & new_n7869_;
  assign new_n5524_ = new_n7744_ & new_n7871_;
  assign new_n5525_ = new_n5524_ | new_n5523_;
  assign new_n5526_ = new_n5525_ & new_n7872_;
  assign new_n5527_ = new_n7757_ & new_n7871_;
  assign new_n5528_ = new_n7770_ & new_n7869_;
  assign new_n5529_ = new_n5528_ | new_n5527_;
  assign new_n5530_ = new_n5529_ & new_n3725_;
  assign new_n5531_ = new_n5530_ | new_n5526_;
  assign new_n5532_ = new_n7728_ & new_n7873_;
  assign new_n5533_ = new_n7744_ & new_n7875_;
  assign new_n5534_ = new_n5533_ | new_n5532_;
  assign new_n5535_ = new_n5534_ & new_n7876_;
  assign new_n5536_ = new_n7760_ & new_n7875_;
  assign new_n5537_ = new_n7773_ & new_n7873_;
  assign new_n5538_ = new_n5537_ | new_n5536_;
  assign new_n5539_ = new_n5538_ & new_n3727_;
  assign new_n5540_ = new_n5539_ | new_n5535_;
  assign new_n5541_ = new_n7745_ & new_n7877_;
  assign new_n5542_ = new_n7729_ & new_n7879_;
  assign new_n5543_ = new_n5542_ | new_n5541_;
  assign new_n5544_ = new_n5543_ & new_n3962_;
  assign new_n5545_ = new_n7760_ & new_n7877_;
  assign new_n5546_ = new_n7773_ & new_n7879_;
  assign new_n5547_ = new_n5546_ | new_n5545_;
  assign new_n5548_ = new_n5547_ & new_n3963_;
  assign new_n5549_ = new_n5548_ | new_n5544_;
  assign new_n5550_ = new_n7881_ & new_n7345_;
  assign new_n5551_ = new_n7882_ | new_n7341_;
  assign new_n5552_ = new_n7882_ & new_n7342_;
  assign new_n5553_ = new_n7881_ | new_n7344_;
  assign new_n5554_ = new_n5553_ & new_n5551_;
  assign new_n5555_ = new_n5552_ | new_n5550_;
  assign new_n5556_ = new_n5555_ & new_n7335_;
  assign new_n5557_ = new_n5554_ & new_n7334_;
  assign new_n5558_ = new_n5557_ | new_n5556_;
  assign new_n5559_ = new_n7802_ & new_n7823_;
  assign new_n5560_ = new_n7801_ & new_n7810_;
  assign new_n5561_ = new_n7819_ | new_n7815_;
  assign new_n5562_ = new_n7820_ & new_n7366_;
  assign new_n5563_ = new_n7801_ | new_n7368_;
  assign new_n5564_ = new_n5563_ & new_n7792_;
  assign new_n5565_ = new_n5562_ | new_n7789_;
  assign new_n5566_ = new_n7883_ & new_n7884_;
  assign new_n5567_ = new_n7885_ | new_n7886_;
  assign new_n5568_ = new_n7885_ & new_n7886_;
  assign new_n5569_ = new_n7883_ | new_n7884_;
  assign new_n5570_ = new_n5569_ & new_n5567_;
  assign new_n5571_ = new_n5568_ | new_n5566_;
  assign new_n5572_ = new_n5570_ & new_n5561_;
  assign new_n5573_ = new_n5571_ & new_n5560_;
  assign new_n5574_ = new_n5573_ | new_n5572_;
  assign new_n5575_ = new_n7887_ | new_n7888_;
  assign new_n5576_ = new_n7887_ & new_n7888_;
  assign new_n5577_ = new_n7425_ & new_n7889_;
  assign new_n5578_ = new_n7433_ & new_n3068_;
  assign new_n5579_ = new_n5578_ | new_n5577_;
  assign new_n5580_ = new_n7462_ | new_n3139_;
  assign new_n5581_ = new_n7451_ | new_n3141_;
  assign new_n5582_ = new_n5581_ & new_n5580_;
  assign new_n5583_ = new_n5116_ | new_n3189_;
  assign new_n5584_ = new_n7890_ & new_n7798_;
  assign new_n5585_ = new_n7825_ | new_n7797_;
  assign new_n5586_ = new_n7821_ | new_n7805_;
  assign new_n5587_ = new_n5586_ & new_n5585_;
  assign new_n5588_ = new_n7891_ | new_n7892_;
  assign new_n5589_ = new_n7891_ & new_n7892_;
  assign new_n5590_ = new_n7893_ | new_n7895_;
  assign new_n5591_ = new_n7896_ | new_n7898_;
  assign new_n5592_ = new_n7900_ & new_n7902_;
  assign new_n5593_ = new_n7900_ | new_n7902_;
  assign new_n5594_ = new_n7904_ & new_n7906_;
  assign new_n5595_ = new_n7904_ | new_n7906_;
  assign new_n5596_ = new_n7729_ & new_n7908_;
  assign new_n5597_ = new_n7911_ | new_n7913_;
  assign new_n5598_ = new_n7774_ & new_n7913_;
  assign new_n5599_ = new_n7916_ | new_n7908_;
  assign new_n5600_ = new_n5599_ & new_n5597_;
  assign new_n5601_ = new_n5598_ | new_n5596_;
  assign new_n5602_ = new_n7731_ & new_n7919_;
  assign new_n5603_ = new_n7911_ | new_n7923_;
  assign new_n5604_ = new_n7745_ & new_n7923_;
  assign new_n5605_ = new_n7926_ | new_n7919_;
  assign new_n5606_ = new_n5605_ & new_n5603_;
  assign new_n5607_ = new_n5604_ | new_n5602_;
  assign new_n5608_ = new_n5607_ & new_n7349_;
  assign new_n5609_ = new_n5606_ | new_n7355_;
  assign new_n5610_ = new_n7761_ & new_n7922_;
  assign new_n5611_ = new_n7929_ | new_n7920_;
  assign new_n5612_ = new_n7774_ & new_n7920_;
  assign new_n5613_ = new_n7916_ | new_n7924_;
  assign new_n5614_ = new_n5613_ & new_n5611_;
  assign new_n5615_ = new_n5612_ | new_n5610_;
  assign new_n5616_ = new_n5615_ & new_n7355_;
  assign new_n5617_ = new_n5614_ | new_n7351_;
  assign new_n5618_ = new_n5617_ & new_n5609_;
  assign new_n5619_ = new_n5616_ | new_n5608_;
  assign new_n5620_ = new_n5619_ & new_n5600_;
  assign new_n5621_ = new_n5618_ & new_n5601_;
  assign new_n5622_ = new_n5621_ | new_n5620_;
  assign new_n5623_ = new_n7931_ | new_n7933_;
  assign new_n5624_ = new_n7931_ & new_n7933_;
  assign new_n5625_ = new_n7731_ & new_n7934_;
  assign new_n5626_ = new_n7747_ & new_n7936_;
  assign new_n5627_ = new_n5626_ | new_n5625_;
  assign new_n5628_ = new_n5627_ & new_n7937_;
  assign new_n5629_ = new_n7761_ & new_n7936_;
  assign new_n5630_ = new_n7776_ & new_n7934_;
  assign new_n5631_ = new_n5630_ | new_n5629_;
  assign new_n5632_ = new_n5631_ & new_n3757_;
  assign new_n5633_ = new_n5632_ | new_n5628_;
  assign new_n5634_ = new_n7910_ | new_n7939_;
  assign new_n5635_ = new_n7926_ | new_n7940_;
  assign new_n5636_ = new_n5635_ & new_n5634_;
  assign new_n5637_ = new_n5636_ | new_n3929_;
  assign new_n5638_ = new_n7929_ | new_n7940_;
  assign new_n5639_ = new_n7915_ | new_n7939_;
  assign new_n5640_ = new_n5639_ & new_n5638_;
  assign new_n5641_ = new_n5640_ | new_n7941_;
  assign new_n5642_ = new_n5641_ & new_n5637_;
  assign new_n5643_ = new_n7942_ | new_n7943_;
  assign new_n5644_ = new_n7942_ & new_n7943_;
  assign new_n5645_ = new_n7480_ & new_n3957_;
  assign new_n5646_ = new_n7475_ & new_n7944_;
  assign new_n5647_ = new_n5646_ | new_n5645_;
  assign new_n5648_ = new_n5647_ & new_n7482_;
  assign new_n5649_ = new_n5648_ | new_n7483_;
  assign new_n5650_ = new_n5649_ & new_n4944_;
  assign new_n5651_ = new_n7945_ & new_n7946_;
  assign new_n5652_ = new_n5651_ | new_n5650_;
  assign new_n5653_ = new_n7947_ & new_n7949_;
  assign new_n5654_ = new_n7951_ | new_n7952_;
  assign new_n5655_ = new_n7951_ & new_n7952_;
  assign new_n5656_ = new_n7947_ | new_n7949_;
  assign new_n5657_ = new_n5656_ & new_n7837_;
  assign new_n5658_ = new_n5655_ | new_n7833_;
  assign new_n5659_ = new_n5657_ & new_n5654_;
  assign new_n5660_ = new_n5658_ | new_n5653_;
  assign new_n5661_ = new_n5660_ & new_n5466_;
  assign new_n5662_ = new_n5659_ | new_n7838_;
  assign new_n5663_ = new_n5661_ | new_n5477_;
  assign new_n5664_ = new_n5662_ | new_n7845_;
  assign new_n5665_ = new_n5664_ & new_n5663_;
  assign new_n5666_ = new_n7732_ & new_n7954_;
  assign new_n5667_ = new_n7912_ | new_n7958_;
  assign new_n5668_ = new_n7747_ & new_n7958_;
  assign new_n5669_ = new_n7927_ | new_n7954_;
  assign new_n5670_ = new_n5669_ & new_n5667_;
  assign new_n5671_ = new_n5668_ | new_n5666_;
  assign new_n5672_ = new_n5671_ & new_n7961_;
  assign new_n5673_ = new_n5670_ | new_n7962_;
  assign new_n5674_ = new_n7762_ & new_n7957_;
  assign new_n5675_ = new_n7930_ | new_n7955_;
  assign new_n5676_ = new_n7776_ & new_n7955_;
  assign new_n5677_ = new_n7917_ | new_n7959_;
  assign new_n5678_ = new_n5677_ & new_n5675_;
  assign new_n5679_ = new_n5676_ | new_n5674_;
  assign new_n5680_ = new_n5679_ & new_n7962_;
  assign new_n5681_ = new_n5678_ | new_n7961_;
  assign new_n5682_ = new_n5681_ & new_n5673_;
  assign new_n5683_ = new_n5680_ | new_n5672_;
  assign new_n5684_ = new_n7732_ & new_n7327_;
  assign new_n5685_ = new_n7912_ | new_n7320_;
  assign new_n5686_ = new_n7746_ & new_n7321_;
  assign new_n5687_ = new_n7927_ | new_n7326_;
  assign new_n5688_ = new_n5687_ & new_n5685_;
  assign new_n5689_ = new_n5686_ | new_n5684_;
  assign new_n5690_ = new_n5689_ & new_n7408_;
  assign new_n5691_ = new_n5688_ | new_n7414_;
  assign new_n5692_ = new_n7762_ & new_n7321_;
  assign new_n5693_ = new_n7930_ | new_n7328_;
  assign new_n5694_ = new_n7775_ & new_n7328_;
  assign new_n5695_ = new_n7917_ | new_n7322_;
  assign new_n5696_ = new_n5695_ & new_n5693_;
  assign new_n5697_ = new_n5694_ | new_n5692_;
  assign new_n5698_ = new_n5697_ & new_n7414_;
  assign new_n5699_ = new_n5696_ | new_n7410_;
  assign new_n5700_ = new_n5699_ & new_n5691_;
  assign new_n5701_ = new_n5698_ | new_n5690_;
  assign new_n5702_ = new_n5701_ & new_n5682_;
  assign new_n5703_ = new_n5700_ & new_n5683_;
  assign new_n5704_ = new_n5703_ | new_n5702_;
  assign new_n5705_ = new_n4862_ & new_n7963_;
  assign new_n5706_ = new_n7964_ | new_n7965_;
  assign new_n5707_ = new_n7339_ & new_n7965_;
  assign new_n5708_ = new_n7343_ | new_n7963_;
  assign new_n5709_ = new_n5708_ & new_n5706_;
  assign new_n5710_ = new_n5707_ | new_n5705_;
  assign new_n5711_ = new_n5710_ & new_n7966_;
  assign new_n5712_ = new_n5709_ & new_n4975_;
  assign new_n5713_ = new_n5712_ | new_n5711_;
  assign new_n5714_ = new_n5408_ | new_n3173_;
  assign new_n5715_ = new_n5414_ | new_n3191_;
  assign new_n5716_ = new_n7967_ | new_n7968_;
  assign new_n5717_ = new_n7969_ | new_n7970_;
  assign new_n5718_ = new_n5717_ & new_n7971_;
  assign new_n5719_ = new_n7451_ & new_n7972_;
  assign new_n5720_ = new_n7463_ & new_n3120_;
  assign new_n5721_ = new_n7452_ & new_n7973_;
  assign new_n5722_ = new_n7463_ & new_n3124_;
  assign new_n5723_ = new_n7975_ & new_n7494_;
  assign new_n5724_ = new_n7975_ | new_n7495_;
  assign new_n5725_ = new_n7977_ & new_n7895_;
  assign new_n5726_ = new_n7980_ & new_n7514_;
  assign new_n5727_ = new_n7981_ & new_n7715_;
  assign new_n5728_ = new_n7982_ & new_n7983_;
  assign new_n5729_ = new_n5728_ | new_n7984_;
  assign new_n5730_ = new_n7977_ & new_n7898_;
  assign new_n5731_ = new_n5730_ | new_n7985_;
  assign new_n5732_ = new_n7896_ & new_n7978_;
  assign new_n5733_ = new_n7986_ | new_n7980_;
  assign new_n5734_ = new_n7988_ & new_n7990_;
  assign new_n5735_ = new_n7988_ | new_n7990_;
  assign new_n5736_ = new_n7991_ & new_n7992_;
  assign new_n5737_ = new_n7993_ | new_n7994_;
  assign new_n5738_ = new_n5737_ & new_n7995_;
  assign new_n5739_ = new_n7996_ | new_n7997_;
  assign new_n5740_ = new_n5739_ & new_n7998_;
  assign new_n5741_ = new_n7999_ & new_n8000_;
  assign new_n5742_ = new_n8002_ & new_n8004_;
  assign new_n5743_ = new_n8006_ & new_n2226_;
  assign new_n5744_ = new_n8002_ & new_n8007_;
  assign new_n5745_ = new_n8006_ & new_n2230_;
  assign new_n5746_ = new_n8003_ & new_n8008_;
  assign new_n5747_ = new_n8005_ & new_n2256_;
  assign G5193 = new_n2897_;
  assign G5194 = new_n3111_;
  assign G5195 = new_n6749_;
  assign G5196 = new_n8010_;
  assign G5197 = new_n3135_;
  assign G5198 = new_n3143_;
  assign G5199 = ~new_n7194_;
  assign G5200 = new_n3209_;
  assign G5201 = G5196;
  assign G5202 = new_n8009_;
  assign G5203 = new_n3129_;
  assign G5204 = new_n3137_;
  assign G5205 = new_n4139_;
  assign G5206 = new_n7193_;
  assign G5207 = new_n6742_;
  assign G5208 = new_n6741_;
  assign G5209 = new_n7192_;
  assign G5210 = new_n4140_;
  assign G5211 = new_n4141_;
  assign G5212 = new_n4142_;
  assign G5213 = new_n7195_;
  assign G5214 = new_n7078_;
  assign G5215 = new_n6747_;
  assign G5216 = new_n6748_;
  assign G5217 = new_n8011_;
  assign G5218 = new_n3116_;
  assign G5219 = G5217;
  assign G5220 = new_n4145_;
  assign G5221 = new_n6758_;
  assign G5222 = new_n8013_;
  assign G5223 = G5222;
  assign G5224 = new_n8014_;
  assign G5225 = G5224;
  assign G5226 = new_n8015_;
  assign G5227 = G5226;
  assign G5228 = new_n4149_;
  assign G5229 = new_n8016_;
  assign G5230 = G5229;
  assign G5231 = new_n4154_;
  assign G5232 = new_n4159_;
  assign G5233 = new_n4164_;
  assign G5234 = new_n4169_;
  assign G5235 = new_n4174_;
  assign G5236 = new_n4180_;
  assign G5237 = new_n4189_;
  assign G5238 = ~new_n8017_;
  assign G5239 = new_n8018_;
  assign G5240 = G5239;
  assign G5241 = G5238;
  assign G5242 = ~new_n7196_;
  assign G5243 = ~new_n7197_;
  assign G5244 = ~new_n8019_;
  assign G5245 = new_n8020_;
  assign G5246 = G5244;
  assign G5247 = G5245;
  assign G5248 = ~new_n6836_;
  assign G5249 = new_n7174_;
  assign G5250 = ~new_n6859_;
  assign G5251 = new_n6969_;
  assign G5252 = new_n4248_;
  assign G5253 = ~new_n7144_;
  assign G5254 = ~new_n7154_;
  assign G5255 = ~new_n7164_;
  assign G5256 = new_n4270_;
  assign G5257 = ~new_n7140_;
  assign G5258 = ~new_n7150_;
  assign G5259 = ~new_n7160_;
  assign G5260 = new_n7170_;
  assign G5261 = ~new_n7198_;
  assign G5262 = ~new_n7199_;
  assign G5263 = ~new_n4372_;
  assign G5264 = ~new_n4381_;
  assign G5265 = new_n4391_;
  assign G5266 = new_n4401_;
  assign G5267 = new_n4410_;
  assign G5268 = new_n4419_;
  assign G5269 = new_n4428_;
  assign G5270 = ~new_n4437_;
  assign G5271 = new_n4446_;
  assign G5272 = new_n4455_;
  assign G5273 = new_n4464_;
  assign G5274 = ~new_n4473_;
  assign G5275 = new_n4483_;
  assign G5276 = ~new_n4493_;
  assign G5277 = new_n4503_;
  assign G5278 = new_n4513_;
  assign G5279 = new_n4523_;
  assign G5280 = ~new_n4533_;
  assign G5281 = new_n4543_;
  assign G5282 = new_n4553_;
  assign G5283 = new_n4570_;
  assign G5284 = new_n4573_;
  assign G5285 = ~new_n7209_;
  assign G5286 = ~new_n7219_;
  assign G5287 = ~new_n7229_;
  assign G5288 = ~new_n7239_;
  assign G5289 = ~new_n4594_;
  assign G5290 = ~new_n7205_;
  assign G5291 = ~new_n7215_;
  assign G5292 = ~new_n7225_;
  assign G5293 = ~new_n7235_;
  assign G5294 = new_n4622_;
  assign G5295 = new_n4631_;
  assign G5296 = new_n4640_;
  assign G5297 = new_n4649_;
  assign G5298 = new_n4658_;
  assign G5299 = new_n4667_;
  assign G5300 = new_n4676_;
  assign G5301 = new_n4685_;
  assign G5302 = new_n4695_;
  assign G5303 = new_n4705_;
  assign G5304 = new_n4715_;
  assign G5305 = new_n4725_;
  assign G5306 = new_n4735_;
  assign G5307 = new_n4745_;
  assign G5308 = new_n4755_;
  assign G5309 = new_n4765_;
  assign G5310 = new_n4769_;
  assign G5311 = new_n4774_;
  assign G5312 = ~new_n4787_;
  assign G5313 = ~new_n4796_;
  assign G5314 = new_n4806_;
  assign G5315 = new_n4816_;
  assign n7230_li000_li000 = new_n2042_;
  assign n7233_li001_li001 = new_n2398_;
  assign n7236_li002_li002 = new_n2400_;
  assign n7239_li003_li003 = new_n2402_;
  assign n7242_li004_li004 = new_n2044_;
  assign n7245_li005_li005 = new_n2406_;
  assign n7248_li006_li006 = new_n2408_;
  assign n7254_li008_li008 = new_n2046_;
  assign n7257_li009_li009 = new_n2412_;
  assign n7260_li010_li010 = new_n2414_;
  assign n7263_li011_li011 = new_n2416_;
  assign n7266_li012_li012 = new_n2048_;
  assign n7269_li013_li013 = new_n2420_;
  assign n7272_li014_li014 = new_n2422_;
  assign n7275_li015_li015 = new_n2424_;
  assign n7278_li016_li016 = new_n2050_;
  assign n7281_li017_li017 = new_n2428_;
  assign n7284_li018_li018 = new_n2430_;
  assign n7287_li019_li019 = new_n2432_;
  assign n7290_li020_li020 = new_n2052_;
  assign n7293_li021_li021 = new_n2436_;
  assign n7296_li022_li022 = new_n2438_;
  assign n7299_li023_li023 = new_n2440_;
  assign n7302_li024_li024 = new_n2054_;
  assign n7305_li025_li025 = new_n2444_;
  assign n7308_li026_li026 = new_n2446_;
  assign n7311_li027_li027 = new_n2448_;
  assign n7314_li028_li028 = new_n2056_;
  assign n7317_li029_li029 = new_n2452_;
  assign n7320_li030_li030 = new_n2454_;
  assign n7323_li031_li031 = new_n2456_;
  assign n7326_li032_li032 = new_n2058_;
  assign n7329_li033_li033 = new_n2460_;
  assign n7332_li034_li034 = new_n2462_;
  assign n7335_li035_li035 = new_n2464_;
  assign n7338_li036_li036 = new_n2060_;
  assign n7341_li037_li037 = new_n2468_;
  assign n7344_li038_li038 = new_n2470_;
  assign n7347_li039_li039 = new_n2472_;
  assign n7350_li040_li040 = new_n2062_;
  assign n7353_li041_li041 = new_n2476_;
  assign n7356_li042_li042 = new_n2478_;
  assign n7359_li043_li043 = new_n2480_;
  assign n7362_li044_li044 = new_n2064_;
  assign n7365_li045_li045 = new_n2484_;
  assign n7368_li046_li046 = new_n2486_;
  assign n7371_li047_li047 = new_n2488_;
  assign n7374_li048_li048 = new_n2066_;
  assign n7377_li049_li049 = new_n2492_;
  assign n7380_li050_li050 = new_n2494_;
  assign n7383_li051_li051 = new_n2496_;
  assign n7386_li052_li052 = new_n2068_;
  assign n7389_li053_li053 = new_n2500_;
  assign n7392_li054_li054 = new_n2502_;
  assign n7395_li055_li055 = new_n2504_;
  assign n7398_li056_li056 = new_n2070_;
  assign n7401_li057_li057 = new_n2508_;
  assign n7404_li058_li058 = new_n2510_;
  assign n7407_li059_li059 = new_n2512_;
  assign n7410_li060_li060 = new_n2072_;
  assign n7413_li061_li061 = new_n2516_;
  assign n7416_li062_li062 = new_n2518_;
  assign n7419_li063_li063 = new_n2520_;
  assign n7422_li064_li064 = new_n2074_;
  assign n7425_li065_li065 = new_n2524_;
  assign n7428_li066_li066 = new_n2526_;
  assign n7431_li067_li067 = new_n2528_;
  assign n7434_li068_li068 = new_n2076_;
  assign n7437_li069_li069 = new_n2532_;
  assign n7440_li070_li070 = new_n2534_;
  assign n7443_li071_li071 = new_n2536_;
  assign n7446_li072_li072 = new_n2078_;
  assign n7449_li073_li073 = new_n2540_;
  assign n7452_li074_li074 = new_n2542_;
  assign n7458_li076_li076 = new_n2080_;
  assign n7461_li077_li077 = new_n2546_;
  assign n7464_li078_li078 = new_n2548_;
  assign n7467_li079_li079 = new_n2550_;
  assign n7470_li080_li080 = new_n2082_;
  assign n7473_li081_li081 = new_n2554_;
  assign n7476_li082_li082 = new_n2556_;
  assign n7482_li084_li084 = new_n2084_;
  assign n7485_li085_li085 = new_n2560_;
  assign n7488_li086_li086 = new_n2562_;
  assign n7491_li087_li087 = new_n2564_;
  assign n7494_li088_li088 = new_n2086_;
  assign n7497_li089_li089 = new_n2568_;
  assign n7500_li090_li090 = new_n2570_;
  assign n7503_li091_li091 = new_n2572_;
  assign n7506_li092_li092 = new_n2088_;
  assign n7509_li093_li093 = new_n2576_;
  assign n7512_li094_li094 = new_n2578_;
  assign n7515_li095_li095 = new_n2580_;
  assign n7518_li096_li096 = new_n2090_;
  assign n7521_li097_li097 = new_n2584_;
  assign n7524_li098_li098 = new_n2586_;
  assign n7527_li099_li099 = new_n2588_;
  assign n7530_li100_li100 = new_n2092_;
  assign n7533_li101_li101 = new_n2592_;
  assign n7536_li102_li102 = new_n2594_;
  assign n7539_li103_li103 = new_n2596_;
  assign n7542_li104_li104 = new_n2094_;
  assign n7545_li105_li105 = new_n2600_;
  assign n7548_li106_li106 = new_n2602_;
  assign n7551_li107_li107 = new_n2604_;
  assign n7554_li108_li108 = new_n2096_;
  assign n7557_li109_li109 = new_n2608_;
  assign n7560_li110_li110 = new_n2610_;
  assign n7563_li111_li111 = new_n2612_;
  assign n7566_li112_li112 = new_n2098_;
  assign n7569_li113_li113 = new_n2616_;
  assign n7572_li114_li114 = new_n2618_;
  assign n7575_li115_li115 = new_n2620_;
  assign n7578_li116_li116 = new_n2100_;
  assign n7581_li117_li117 = new_n2624_;
  assign n7584_li118_li118 = new_n2626_;
  assign n7587_li119_li119 = new_n2628_;
  assign n7590_li120_li120 = new_n2102_;
  assign n7593_li121_li121 = new_n2632_;
  assign n7596_li122_li122 = new_n2634_;
  assign n7599_li123_li123 = new_n2636_;
  assign n7602_li124_li124 = new_n2104_;
  assign n7605_li125_li125 = new_n2640_;
  assign n7608_li126_li126 = new_n2642_;
  assign n7611_li127_li127 = new_n2644_;
  assign n7614_li128_li128 = new_n2106_;
  assign n7617_li129_li129 = new_n2648_;
  assign n7620_li130_li130 = new_n2650_;
  assign n7623_li131_li131 = new_n2652_;
  assign n7626_li132_li132 = new_n2108_;
  assign n7629_li133_li133 = new_n2656_;
  assign n7632_li134_li134 = new_n2658_;
  assign n7635_li135_li135 = new_n2660_;
  assign n7638_li136_li136 = new_n2110_;
  assign n7641_li137_li137 = new_n2664_;
  assign n7644_li138_li138 = new_n2666_;
  assign n7647_li139_li139 = new_n2668_;
  assign n7650_li140_li140 = new_n2112_;
  assign n7653_li141_li141 = new_n2672_;
  assign n7656_li142_li142 = new_n2674_;
  assign n7659_li143_li143 = new_n2676_;
  assign n7662_li144_li144 = new_n2114_;
  assign n7665_li145_li145 = new_n2680_;
  assign n7668_li146_li146 = new_n2682_;
  assign n7671_li147_li147 = new_n2684_;
  assign n7674_li148_li148 = new_n2116_;
  assign n7677_li149_li149 = new_n2688_;
  assign n7680_li150_li150 = new_n2690_;
  assign n7683_li151_li151 = new_n2692_;
  assign n7686_li152_li152 = new_n2118_;
  assign n7689_li153_li153 = new_n2696_;
  assign n7692_li154_li154 = new_n2698_;
  assign n7695_li155_li155 = new_n2700_;
  assign n7698_li156_li156 = new_n2120_;
  assign n7701_li157_li157 = new_n2704_;
  assign n7704_li158_li158 = new_n2706_;
  assign n7707_li159_li159 = new_n2708_;
  assign n7710_li160_li160 = new_n2122_;
  assign n7713_li161_li161 = new_n2712_;
  assign n7716_li162_li162 = new_n2714_;
  assign n7719_li163_li163 = new_n2716_;
  assign n7722_li164_li164 = new_n2124_;
  assign n7725_li165_li165 = new_n2720_;
  assign n7728_li166_li166 = new_n2722_;
  assign n7731_li167_li167 = new_n2724_;
  assign n7734_li168_li168 = new_n2126_;
  assign n7737_li169_li169 = new_n2728_;
  assign n7740_li170_li170 = new_n2730_;
  assign n7746_li172_li172 = new_n2128_;
  assign n7749_li173_li173 = new_n2734_;
  assign n7752_li174_li174 = new_n2736_;
  assign n7758_li176_li176 = new_n2130_;
  assign n7761_li177_li177 = new_n2740_;
  assign n7764_li178_li178 = new_n2742_;
  assign n7767_li179_li179 = new_n2744_;
  assign n7770_li180_li180 = new_n2132_;
  assign n7773_li181_li181 = new_n2748_;
  assign n7776_li182_li182 = new_n2750_;
  assign n7782_li184_li184 = new_n2134_;
  assign n7785_li185_li185 = new_n2754_;
  assign n7788_li186_li186 = new_n2756_;
  assign n7794_li188_li188 = new_n2136_;
  assign n7797_li189_li189 = new_n2760_;
  assign n7800_li190_li190 = new_n2762_;
  assign n7806_li192_li192 = new_n2138_;
  assign n7809_li193_li193 = new_n2766_;
  assign n7812_li194_li194 = new_n2768_;
  assign n7815_li195_li195 = new_n2770_;
  assign n7818_li196_li196 = new_n2140_;
  assign n7821_li197_li197 = new_n2774_;
  assign n7824_li198_li198 = new_n2776_;
  assign n7830_li200_li200 = new_n2142_;
  assign n7833_li201_li201 = new_n2780_;
  assign n7836_li202_li202 = new_n2782_;
  assign n7839_li203_li203 = new_n2784_;
  assign n7842_li204_li204 = new_n2144_;
  assign n7845_li205_li205 = new_n2788_;
  assign n7848_li206_li206 = new_n2790_;
  assign n7854_li208_li208 = new_n2146_;
  assign n7857_li209_li209 = new_n2794_;
  assign n7860_li210_li210 = new_n2796_;
  assign n7863_li211_li211 = new_n2798_;
  assign n7866_li212_li212 = new_n2148_;
  assign n7869_li213_li213 = new_n2802_;
  assign n7872_li214_li214 = new_n2804_;
  assign n7875_li215_li215 = new_n7547_;
  assign n7878_li216_li216 = new_n2150_;
  assign n7881_li217_li217 = new_n2810_;
  assign n7884_li218_li218 = new_n2812_;
  assign n7887_li219_li219 = new_n2814_;
  assign n7890_li220_li220 = new_n2152_;
  assign n7893_li221_li221 = new_n2818_;
  assign n7896_li222_li222 = new_n2820_;
  assign n7899_li223_li223 = new_n2822_;
  assign n7902_li224_li224 = new_n2154_;
  assign n7905_li225_li225 = new_n2826_;
  assign n7908_li226_li226 = new_n2828_;
  assign n7914_li228_li228 = new_n2156_;
  assign n7917_li229_li229 = new_n2832_;
  assign n7920_li230_li230 = new_n2834_;
  assign n7926_li232_li232 = new_n2158_;
  assign n7929_li233_li233 = new_n2838_;
  assign n7932_li234_li234 = new_n2840_;
  assign n7938_li236_li236 = new_n2160_;
  assign n7941_li237_li237 = new_n2844_;
  assign n7944_li238_li238 = new_n2846_;
  assign n7950_li240_li240 = new_n2162_;
  assign n7953_li241_li241 = new_n2850_;
  assign n7956_li242_li242 = new_n2852_;
  assign n7959_li243_li243 = new_n2854_;
  assign n7962_li244_li244 = new_n2164_;
  assign n7965_li245_li245 = new_n2858_;
  assign n7968_li246_li246 = new_n2860_;
  assign n7971_li247_li247 = new_n2862_;
  assign n7974_li248_li248 = new_n2166_;
  assign n7977_li249_li249 = new_n2866_;
  assign n7980_li250_li250 = new_n2868_;
  assign n7983_li251_li251 = new_n2870_;
  assign n7986_li252_li252 = new_n2168_;
  assign n7989_li253_li253 = new_n2874_;
  assign n7992_li254_li254 = new_n2876_;
  assign n7995_li255_li255 = new_n2878_;
  assign n7998_li256_li256 = new_n2170_;
  assign n8001_li257_li257 = new_n2882_;
  assign n8004_li258_li258 = new_n2884_;
  assign n8007_li259_li259 = new_n2886_;
  assign n8010_li260_li260 = new_n2172_;
  assign n8013_li261_li261 = new_n2890_;
  assign n8016_li262_li262 = new_n2892_;
  assign n8019_li263_li263 = new_n2894_;
  assign n8022_li264_li264 = new_n2174_;
  assign n8025_li265_li265 = new_n2898_;
  assign n8028_li266_li266 = new_n2900_;
  assign n8031_li267_li267 = new_n2902_;
  assign n8034_li268_li268 = new_n2176_;
  assign n8037_li269_li269 = new_n2906_;
  assign n8040_li270_li270 = new_n2908_;
  assign n8043_li271_li271 = new_n2910_;
  assign n8046_li272_li272 = new_n2178_;
  assign n8049_li273_li273 = new_n2914_;
  assign n8052_li274_li274 = new_n2916_;
  assign n8055_li275_li275 = new_n2918_;
  assign n8058_li276_li276 = new_n2180_;
  assign n8061_li277_li277 = new_n2922_;
  assign n8064_li278_li278 = new_n2924_;
  assign n8067_li279_li279 = new_n2926_;
  assign n8070_li280_li280 = new_n2182_;
  assign n8073_li281_li281 = new_n2930_;
  assign n8076_li282_li282 = new_n2932_;
  assign n8079_li283_li283 = new_n2934_;
  assign n8082_li284_li284 = new_n2184_;
  assign n8085_li285_li285 = new_n2938_;
  assign n8088_li286_li286 = new_n2940_;
  assign n8091_li287_li287 = new_n2942_;
  assign n8094_li288_li288 = new_n2186_;
  assign n8097_li289_li289 = new_n2946_;
  assign n8100_li290_li290 = new_n2948_;
  assign n8103_li291_li291 = new_n2950_;
  assign n8106_li292_li292 = new_n2188_;
  assign n8109_li293_li293 = new_n2954_;
  assign n8112_li294_li294 = new_n2956_;
  assign n8115_li295_li295 = new_n2958_;
  assign n8118_li296_li296 = new_n2190_;
  assign n8121_li297_li297 = new_n2962_;
  assign n8124_li298_li298 = new_n2964_;
  assign n8127_li299_li299 = new_n2966_;
  assign n8130_li300_li300 = new_n2192_;
  assign n8133_li301_li301 = new_n2970_;
  assign n8136_li302_li302 = new_n2972_;
  assign n8139_li303_li303 = new_n2974_;
  assign n8142_li304_li304 = new_n2194_;
  assign n8145_li305_li305 = new_n2978_;
  assign n8148_li306_li306 = new_n2980_;
  assign n8151_li307_li307 = new_n2982_;
  assign n8154_li308_li308 = new_n2196_;
  assign n8157_li309_li309 = new_n2986_;
  assign n8160_li310_li310 = new_n2988_;
  assign n8163_li311_li311 = new_n2990_;
  assign n8166_li312_li312 = new_n2198_;
  assign n8169_li313_li313 = new_n2994_;
  assign n8172_li314_li314 = new_n2996_;
  assign n8175_li315_li315 = new_n2998_;
  assign n8178_li316_li316 = new_n2200_;
  assign n8181_li317_li317 = new_n3002_;
  assign n8184_li318_li318 = new_n3004_;
  assign n8187_li319_li319 = new_n3006_;
  assign n8190_li320_li320 = new_n2202_;
  assign n8193_li321_li321 = new_n3010_;
  assign n8196_li322_li322 = new_n3012_;
  assign n8199_li323_li323 = new_n3014_;
  assign n8202_li324_li324 = new_n2204_;
  assign n8205_li325_li325 = new_n3018_;
  assign n8208_li326_li326 = new_n3020_;
  assign n8211_li327_li327 = new_n3022_;
  assign n8214_li328_li328 = new_n2206_;
  assign n8217_li329_li329 = new_n3026_;
  assign n8220_li330_li330 = new_n3028_;
  assign n8223_li331_li331 = new_n3030_;
  assign n8226_li332_li332 = new_n2208_;
  assign n8229_li333_li333 = new_n3034_;
  assign n8232_li334_li334 = new_n3036_;
  assign n8235_li335_li335 = new_n3038_;
  assign n8238_li336_li336 = new_n2210_;
  assign n8241_li337_li337 = new_n3042_;
  assign n8244_li338_li338 = new_n3044_;
  assign n8247_li339_li339 = new_n3046_;
  assign n8250_li340_li340 = new_n2212_;
  assign n8253_li341_li341 = new_n3050_;
  assign n8256_li342_li342 = new_n3052_;
  assign n8259_li343_li343 = new_n3054_;
  assign n8262_li344_li344 = new_n2214_;
  assign n8265_li345_li345 = new_n3058_;
  assign n8268_li346_li346 = new_n3060_;
  assign n8271_li347_li347 = new_n3062_;
  assign n8274_li348_li348 = new_n2216_;
  assign n8286_li352_li352 = new_n2218_;
  assign n8370_li380_li380 = new_n2232_;
  assign n8382_li384_li384 = new_n2234_;
  assign n8394_li388_li388 = new_n2236_;
  assign n8406_li392_li392 = new_n2238_;
  assign n8409_li393_li393 = new_n3076_;
  assign n8412_li394_li394 = new_n3078_;
  assign n8415_li395_li395 = new_n3080_;
  assign n8418_li396_li396 = new_n2240_;
  assign n8430_li400_li400 = new_n2242_;
  assign n8442_li404_li404 = new_n2244_;
  assign n8454_li408_li408 = new_n2246_;
  assign n8466_li412_li412 = new_n2248_;
  assign n8550_li440_li440 = new_n2262_;
  assign n8553_li441_li441 = new_n3094_;
  assign n8556_li442_li442 = new_n3096_;
  assign n8562_li444_li444 = new_n2264_;
  assign n8565_li445_li445 = new_n3100_;
  assign n8568_li446_li446 = new_n3102_;
  assign n8574_li448_li448 = new_n2266_;
  assign n8577_li449_li449 = new_n3106_;
  assign n8583_li451_li451 = new_n7686_;
  assign n8586_li452_li452 = new_n2268_;
  assign n8589_li453_li453 = new_n3112_;
  assign n8595_li455_li455 = new_n3712_;
  assign n8598_li456_li456 = new_n2270_;
  assign n8610_li460_li460 = new_n2272_;
  assign n8670_li480_li480 = new_n2282_;
  assign n8682_li484_li484 = new_n2284_;
  assign n8718_li496_li496 = new_n2290_;
  assign n8727_li499_li499 = new_n3538_;
  assign n8730_li500_li500 = new_n2292_;
  assign n8742_li504_li504 = new_n2294_;
  assign n8751_li507_li507 = new_n3514_;
  assign n8775_li515_li515 = new_n3498_;
  assign n8778_li516_li516 = new_n2300_;
  assign n8790_li520_li520 = new_n2302_;
  assign n8799_li523_li523 = new_n3542_;
  assign n8802_li524_li524 = new_n2304_;
  assign n8805_li525_li525 = new_n3144_;
  assign n8808_li526_li526 = new_n3146_;
  assign n8814_li528_li528 = new_n2306_;
  assign n8817_li529_li529 = new_n3150_;
  assign n8820_li530_li530 = new_n3152_;
  assign n8826_li532_li532 = new_n2308_;
  assign n8829_li533_li533 = new_n3156_;
  assign n8832_li534_li534 = new_n3158_;
  assign n8835_li535_li535 = new_n3160_;
  assign n8850_li540_li540 = new_n2312_;
  assign n8853_li541_li541 = new_n3164_;
  assign n8856_li542_li542 = new_n3166_;
  assign n8859_li543_li543 = new_n3168_;
  assign n8862_li544_li544 = new_n2314_;
  assign n8874_li548_li548 = new_n2316_;
  assign n8910_li560_li560 = new_n2322_;
  assign n8913_li561_li561 = new_n3176_;
  assign n8922_li564_li564 = new_n2324_;
  assign n8934_li568_li568 = new_n2326_;
  assign n8970_li580_li580 = new_n2332_;
  assign n8982_li584_li584 = new_n2334_;
  assign n8994_li588_li588 = new_n2336_;
  assign n9006_li592_li592 = new_n2338_;
  assign n9018_li596_li596 = new_n2340_;
  assign n9030_li600_li600 = new_n2342_;
  assign n9033_li601_li601 = new_n3194_;
  assign n9036_li602_li602 = new_n3196_;
  assign n9039_li603_li603 = new_n3198_;
  assign n9042_li604_li604 = new_n2344_;
  assign n9045_li605_li605 = new_n3202_;
  assign n9048_li606_li606 = new_n3204_;
  assign n9051_li607_li607 = new_n3206_;
  assign n9054_li608_li608 = new_n2346_;
  assign n9057_li609_li609 = new_n3210_;
  assign n9060_li610_li610 = new_n3212_;
  assign n9063_li611_li611 = new_n3214_;
  assign n9066_li612_li612 = new_n2348_;
  assign n9069_li613_li613 = new_n3218_;
  assign n9072_li614_li614 = new_n3220_;
  assign n9075_li615_li615 = new_n3222_;
  assign n9078_li616_li616 = new_n2350_;
  assign n9081_li617_li617 = new_n3226_;
  assign n9084_li618_li618 = new_n3228_;
  assign n9087_li619_li619 = new_n3230_;
  assign n9090_li620_li620 = new_n2352_;
  assign n9093_li621_li621 = new_n3234_;
  assign n9096_li622_li622 = new_n3236_;
  assign n9099_li623_li623 = new_n3238_;
  assign n9102_li624_li624 = new_n2354_;
  assign n9105_li625_li625 = new_n3242_;
  assign n9108_li626_li626 = new_n3244_;
  assign n9114_li628_li628 = new_n2356_;
  assign n9117_li629_li629 = new_n3248_;
  assign n9120_li630_li630 = new_n3250_;
  assign n9123_li631_li631 = new_n3252_;
  assign n9126_li632_li632 = new_n2358_;
  assign n9129_li633_li633 = new_n3256_;
  assign n9132_li634_li634 = new_n3258_;
  assign n9135_li635_li635 = new_n3260_;
  assign n9138_li636_li636 = new_n2360_;
  assign n9141_li637_li637 = new_n3264_;
  assign n9144_li638_li638 = new_n3266_;
  assign n9147_li639_li639 = new_n3268_;
  assign n9150_li640_li640 = new_n2362_;
  assign n9153_li641_li641 = new_n3272_;
  assign n9156_li642_li642 = new_n3274_;
  assign n9159_li643_li643 = new_n3276_;
  assign n9162_li644_li644 = new_n2364_;
  assign n9165_li645_li645 = new_n3280_;
  assign n9174_li648_li648 = new_n2366_;
  assign n9177_li649_li649 = new_n3284_;
  assign n9180_li650_li650 = new_n3286_;
  assign n9183_li651_li651 = new_n3288_;
  assign n9186_li652_li652 = new_n2368_;
  assign n9189_li653_li653 = new_n3292_;
  assign n9192_li654_li654 = new_n3294_;
  assign n9195_li655_li655 = new_n3296_;
  assign n9198_li656_li656 = new_n2370_;
  assign n9201_li657_li657 = new_n3300_;
  assign n9204_li658_li658 = new_n3302_;
  assign n9207_li659_li659 = new_n3304_;
  assign n9210_li660_li660 = new_n2372_;
  assign n9213_li661_li661 = new_n3308_;
  assign n9216_li662_li662 = new_n3310_;
  assign n9222_li664_li664 = new_n2374_;
  assign n9225_li665_li665 = new_n3314_;
  assign n9228_li666_li666 = new_n3316_;
  assign n9234_li668_li668 = new_n2376_;
  assign n9237_li669_li669 = new_n3320_;
  assign n9240_li670_li670 = new_n3322_;
  assign n9246_li672_li672 = new_n2378_;
  assign n9249_li673_li673 = new_n3326_;
  assign n9252_li674_li674 = new_n3328_;
  assign n9258_li676_li676 = new_n2380_;
  assign n9261_li677_li677 = new_n3332_;
  assign n9264_li678_li678 = new_n3334_;
  assign n9267_li679_li679 = new_n3336_;
  assign n9270_li680_li680 = new_n2382_;
  assign n9273_li681_li681 = new_n3340_;
  assign n9276_li682_li682 = new_n3342_;
  assign n9279_li683_li683 = new_n3344_;
  assign n9282_li684_li684 = new_n2384_;
  assign n9285_li685_li685 = new_n3348_;
  assign n9288_li686_li686 = new_n3350_;
  assign n9291_li687_li687 = new_n3352_;
  assign n9294_li688_li688 = new_n2386_;
  assign n9297_li689_li689 = new_n3356_;
  assign n9300_li690_li690 = new_n3358_;
  assign n9303_li691_li691 = new_n3360_;
  assign n9306_li692_li692 = new_n2388_;
  assign n9309_li693_li693 = new_n3364_;
  assign n9312_li694_li694 = new_n3366_;
  assign n9315_li695_li695 = new_n3368_;
  assign n9318_li696_li696 = new_n2390_;
  assign n9321_li697_li697 = new_n3372_;
  assign n9324_li698_li698 = new_n3374_;
  assign n9327_li699_li699 = new_n3376_;
  assign n9330_li700_li700 = new_n2392_;
  assign n9333_li701_li701 = new_n3380_;
  assign n9336_li702_li702 = new_n3382_;
  assign n9339_li703_li703 = new_n7548_;
  assign n9342_li704_li704 = new_n2394_;
  assign n9345_li705_li705 = new_n3388_;
  assign n9348_li706_li706 = new_n3390_;
  assign n9351_li707_li707 = new_n7540_;
  assign n9354_li708_li708 = new_n2396_;
  assign n9357_li709_li709 = new_n3396_;
  assign n9360_li710_li710 = new_n3398_;
  assign n9363_li711_li711 = new_n3400_;
  assign n4970_i2 = new_n3490_;
  assign n4972_i2 = new_n3494_;
  assign n4989_i2 = new_n3506_;
  assign n5024_i2 = new_n3524_;
  assign n5025_i2 = new_n3526_;
  assign n5029_i2 = new_n3534_;
  assign n5042_i2 = new_n3548_;
  assign n5048_i2 = new_n3556_;
  assign n5093_i2 = new_n3568_;
  assign n5096_i2 = new_n3574_;
  assign n5193_i2 = new_n3602_;
  assign n5199_i2 = new_n3610_;
  assign n5203_i2 = new_n7684_;
  assign n5214_i2 = new_n7267_;
  assign n5221_i2 = new_n7685_;
  assign n5222_i2 = new_n7554_;
  assign n5273_i2 = new_n3632_;
  assign n5365_i2 = new_n3650_;
  assign n5385_i2 = new_n3658_;
  assign n5553_i2 = new_n3692_;
  assign n5636_i2 = new_n3738_;
  assign n5782_i2 = new_n3922_;
  assign n5778_i2 = new_n3918_;
  assign n5323_i2 = new_n7862_;
  assign n5325_i2 = new_n7858_;
  assign n5327_i2 = new_n7854_;
  assign n5329_i2 = new_n7323_;
  assign n5816_i2 = new_n7595_;
  assign n5817_i2 = new_n7585_;
  assign n5837_i2 = new_n7265_;
  assign n5844_i2 = new_n7659_;
  assign n5859_i2 = new_n7577_;
  assign n5857_i2 = new_n7578_;
  assign n5369_i2 = new_n7866_;
  assign n5371_i2 = new_n7748_;
  assign n5373_i2 = new_n7851_;
  assign n5400_i2 = new_n7874_;
  assign n5402_i2 = new_n7870_;
  assign n5404_i2 = new_n7778_;
  assign n5406_i2 = new_n7856_;
  assign n5407_i2 = new_n7860_;
  assign n5408_i2 = new_n7864_;
  assign n2722_i2 = new_n7269_;
  assign n5411_i2 = new_n3672_;
  assign n5412_i2 = new_n3674_;
  assign n5413_i2 = new_n3676_;
  assign n5557_i2 = new_n7935_;
  assign n5558_i2 = new_n3696_;
  assign n5559_i2 = new_n7868_;
  assign n5564_i2 = new_n3704_;
  assign n5565_i2 = new_n3706_;
  assign n5561_i2 = new_n3702_;
  assign n5568_i2 = new_n3710_;
  assign n5598_i2 = new_n7959_;
  assign n5600_i2 = new_n7938_;
  assign n5601_i2 = new_n3722_;
  assign n5602_i2 = new_n7872_;
  assign n5603_i2 = new_n7876_;
  assign n2853_i2 = new_n7565_;
  assign n5637_i2 = new_n7807_;
  assign n5627_i2 = new_n3730_;
  assign n5628_i2 = new_n3732_;
  assign n5635_i2 = new_n3736_;
  assign n5640_i2 = new_n7817_;
  assign n5641_i2 = new_n7837_;
  assign n5642_i2 = new_n7841_;
  assign n5650_i2 = new_n7878_;
  assign n5652_i2 = new_n3750_;
  assign n5653_i2 = new_n7780_;
  assign n5654_i2 = new_n3754_;
  assign n5655_i2 = new_n7937_;
  assign n5657_i2 = new_n3760_;
  assign n5659_i2 = new_n3762_;
  assign n5661_i2 = new_n7331_;
  assign n5656_i2 = new_n3758_;
  assign n5663_i2 = new_n3766_;
  assign n5664_i2 = new_n3768_;
  assign n5795_i2 = new_n7960_;
  assign n5796_i2 = new_n7907_;
  assign n5797_i2 = new_n7941_;
  assign n5739_i2 = new_n3846_;
  assign n5773_i2 = new_n7815_;
  assign n5798_i2 = new_n3930_;
  assign n5799_i2 = new_n3932_;
  assign n5802_i2 = new_n7366_;
  assign n5803_i2 = new_n7292_;
  assign n5831_i2 = new_n7781_;
  assign n5833_i2 = new_n7924_;
  assign n5820_i2 = new_n7330_;
  assign n5823_i2 = new_n7816_;
  assign n5824_i2 = new_n7944_;
  assign n5869_i2 = new_n7793_;
  assign n5848_i2 = new_n3986_;
  assign n5849_i2 = new_n7342_;
  assign n5856_i2 = new_n3996_;
  assign n5896_i2 = new_n7322_;
  assign n2754_i2 = ~new_n7613_;
  assign n2908_i2 = new_n7358_;
  assign n5892_i2 = new_n7820_;
  assign n5915_i2 = new_n7285_;
  assign n5919_i2 = new_n7363_;
  assign n5918_i2 = new_n7287_;
  assign n5920_i2 = new_n7286_;
  assign n5917_i2 = new_n7281_;
  assign lo586_buf_i2 = new_n7351_;
  assign n2818_i2 = new_n7948_;
  assign n2863_i2 = new_n7334_;
  assign n2721_i2 = new_n7480_;
  assign n2725_i2 = new_n7346_;
  assign n3016_i2 = new_n7950_;
  assign n3013_i2 = new_n7829_;
  assign n2655_i2 = new_n7290_;
  assign n2741_i2 = new_n7464_;
  assign lo562_buf_i2 = new_n7410_;
  assign n2656_i2 = new_n7839_;
  assign n2531_i2 = new_n7621_;
  assign n2700_i2 = new_n7405_;
  assign n5908_i2 = new_n4070_;
  assign n5910_i2 = new_n4072_;
  assign n5912_i2 = new_n4074_;
  assign n5914_i2 = new_n7425_;
  assign n2753_i2 = new_n7481_;
  assign n2878_i2 = new_n7880_;
  assign n2836_i2 = new_n7964_;
  assign n5934_i2 = new_n7416_;
  assign n5936_i2 = new_n7453_;
  assign n5938_i2 = new_n7452_;
  assign n2728_i2 = new_n7466_;
  assign lo358_buf_i2 = new_n7472_;
  assign lo418_buf_i2 = new_n7473_;
  assign lo474_buf_i2 = new_n7484_;
  assign lo554_buf_i2 = new_n7491_;
  assign lo558_buf_i2 = new_n7436_;
  assign lo574_buf_i2 = new_n7440_;
  assign n2659_i2 = new_n7438_;
  assign n2665_i2 = new_n7434_;
  assign n2686_i2 = new_n7489_;
  assign lo450_buf_i2 = new_n7782_;
  assign n2910_i2 = new_n7608_;
  assign n2683_i2 = new_n4878_;
  assign n2828_i2 = ~new_n7615_;
  assign n2582_i2 = new_n7571_;
  assign n2600_i2 = new_n7572_;
  assign n2542_i2 = new_n7570_;
  assign n2703_i2 = new_n7796_;
  assign lo510_buf_i2 = new_n7496_;
  assign lo514_buf_i2 = new_n7497_;
  assign lo538_buf_i2 = new_n7487_;
  assign lo578_buf_i2 = new_n7512_;
  assign n2692_i2 = new_n7485_;
  assign n2666_i2 = new_n7717_;
  assign n2667_i2 = new_n7495_;
  assign n2660_i2 = new_n7894_;
  assign n2744_i2 = new_n7510_;
  assign lo454_buf_i2 = new_n7852_;
  assign n3593_i2 = new_n7890_;
  assign n3048_i2 = new_n7946_;
  assign lo410_buf_i2 = new_n7784_;
  assign lo502_buf_i2 = new_n7785_;
  assign lo506_buf_i2 = new_n7786_;
  assign lo550_buf_i2 = new_n7500_;
  assign lo570_buf_i2 = new_n7504_;
  assign lo582_buf_i2 = new_n7508_;
  assign n2646_i2 = new_n7502_;
  assign n2673_i2 = new_n7498_;
  assign n3499_i2 = ~new_n7945_;
  assign n2750_i2 = new_n7506_;
  assign n2870_i2 = new_n7966_;
  assign n2693_i2 = new_n7716_;
  assign n2689_i2 = new_n7714_;
  assign n2668_i2 = new_n7517_;
  assign n2662_i2 = new_n7515_;
  assign lo350_buf_i2 = new_n7889_;
  assign lo498_buf_i2 = new_n7618_;
  assign lo518_buf_i2 = new_n3138_;
  assign lo522_buf_i2 = new_n3140_;
  assign lo598_buf_i2 = new_n7970_;
  assign n2708_i2 = new_n7969_;
  assign n2674_i2 = new_n7984_;
  assign n2647_i2 = new_n7985_;
  assign n2751_i2 = new_n7850_;
  assign n2747_i2 = new_n7849_;
  assign n2669_i2 = new_n7893_;
  assign n2872_i2 = new_n5001_;
  assign n3313_i2 = new_n5002_;
  assign n3273_i2 = new_n5003_;
  assign n2848_i2 = new_n5004_;
  assign n2893_i2 = new_n5005_;
  assign n3267_i2 = new_n5006_;
  assign n2925_i2 = new_n5007_;
  assign n2839_i2 = new_n5008_;
  assign n2831_i2 = new_n5009_;
  assign n2558_i2 = new_n5013_;
  assign n2562_i2 = new_n5017_;
  assign n2825_i2 = new_n5018_;
  assign n3263_i2 = new_n5020_;
  assign n3517_i2 = new_n5052_;
  assign n2873_i2 = ~new_n5053_;
  assign n2926_i2 = ~new_n5054_;
  assign n3261_i2 = new_n5055_;
  assign n3268_i2 = new_n5056_;
  assign n3274_i2 = new_n5057_;
  assign n3314_i2 = ~new_n5058_;
  assign n3571_i2 = new_n5083_;
  assign n2950_i2 = new_n5084_;
  assign n2951_i2 = new_n5085_;
  assign n3022_i2 = new_n5090_;
  assign n3023_i2 = new_n5091_;
  assign n3057_i2 = ~new_n5095_;
  assign n3058_i2 = ~new_n5096_;
  assign n2931_i2 = new_n5097_;
  assign n2911_i2 = new_n5098_;
  assign n2959_i2 = new_n5102_;
  assign n2960_i2 = new_n5103_;
  assign n2922_i2 = new_n5104_;
  assign n2888_i2 = new_n5105_;
  assign n2889_i2 = new_n5106_;
  assign n3051_i2 = ~new_n5109_;
  assign n3052_i2 = ~new_n5110_;
  assign n3063_i2 = ~new_n5111_;
  assign n2845_i2 = new_n5115_;
  assign n2737_i2 = new_n7993_;
  assign n3281_i2 = new_n5120_;
  assign n3294_i2 = new_n5123_;
  assign n2885_i2 = ~new_n5126_;
  assign n2786_i2 = new_n5129_;
  assign n2783_i2 = new_n5132_;
  assign n2801_i2 = new_n5135_;
  assign n2572_i2 = new_n5144_;
  assign n2628_i2 = new_n5153_;
  assign n2609_i2 = new_n5162_;
  assign n2618_i2 = new_n5171_;
  assign n2637_i2 = new_n5180_;
  assign n2525_i2 = new_n5189_;
  assign n2551_i2 = new_n5198_;
  assign n3759_i2 = new_n5238_;
  assign n2994_i2 = new_n5241_;
  assign n3040_i2 = new_n5244_;
  assign n2943_i2 = new_n5249_;
  assign n2991_i2 = new_n5258_;
  assign n3034_i2 = new_n5261_;
  assign n2881_i2 = new_n5264_;
  assign n3021_i2 = new_n5273_;
  assign n3062_i2 = new_n5276_;
  assign n2763_i2 = new_n5283_;
  assign n2764_i2 = ~new_n5284_;
  assign n2775_i2 = new_n5297_;
  assign n2776_i2 = ~new_n5298_;
  assign n2968_i2 = new_n5305_;
  assign n2969_i2 = new_n5306_;
  assign n2798_i2 = new_n5321_;
  assign n3661_i2 = new_n5372_;
  assign n2694_i2 = new_n7848_;
  assign n2809_i2 = new_n7983_;
  assign n2817_i2 = new_n7897_;
  assign n2514_i2 = new_n7901_;
  assign n2501_i2 = new_n7905_;
  assign n2528_i2 = ~new_n7932_;
  assign n2505_i2 = ~new_n7899_;
  assign n2492_i2 = new_n7903_;
  assign lo546_buf_i2 = new_n7997_;
  assign lo590_buf_i2 = new_n7994_;
  assign lo594_buf_i2 = new_n7968_;
  assign n2679_i2 = new_n7996_;
  assign n2733_i2 = new_n7967_;
  assign n2709_i2 = ~new_n7971_;
  assign n2676_i2 = new_n7982_;
  assign n2649_i2 = new_n7978_;
  assign n2815_i2 = new_n5426_;
  assign n2704_i2 = ~new_n5428_;
  assign n3590_i2 = ~new_n5454_;
  assign n3591_i2 = ~new_n5455_;
  assign n2752_i2 = new_n7979_;
  assign n3638_i2 = new_n5479_;
  assign n3639_i2 = new_n5480_;
  assign n2695_i2 = new_n7981_;
  assign n3047_i2 = new_n7986_;
  assign lo458_buf_i2 = new_n7972_;
  assign lo482_buf_i2 = new_n7973_;
  assign lo566_buf_i2 = new_n7989_;
  assign n2718_i2 = new_n5486_;
  assign n3707_i2 = new_n5495_;
  assign n3671_i2 = new_n5504_;
  assign n3680_i2 = new_n5513_;
  assign n3749_i2 = new_n5522_;
  assign n3716_i2 = new_n5531_;
  assign n3692_i2 = new_n5540_;
  assign n2591_i2 = new_n5549_;
  assign n3478_i2 = new_n5558_;
  assign n3610_i2 = ~new_n5575_;
  assign n3611_i2 = ~new_n5576_;
  assign n2652_i2 = new_n7987_;
  assign n2714_i2 = ~new_n7992_;
  assign n2738_i2 = ~new_n7995_;
  assign n3616_i2 = new_n5588_;
  assign n3617_i2 = new_n5589_;
  assign n3031_i2 = new_n7974_;
  assign n2515_i2 = new_n5592_;
  assign n3562_i2 = ~new_n5593_;
  assign n2502_i2 = new_n5594_;
  assign n3560_i2 = new_n5595_;
  assign n3554_i2 = ~new_n5623_;
  assign n3555_i2 = new_n5624_;
  assign n3536_i2 = ~new_n5643_;
  assign n3537_i2 = new_n5644_;
  assign n3508_i2 = ~new_n5652_;
  assign n3650_i2 = new_n5665_;
  assign n3740_i2 = new_n5704_;
  assign n3484_i2 = new_n5713_;
  assign n2680_i2 = ~new_n7998_;
  assign n2734_i2 = ~new_n8000_;
  assign n2735_i2 = new_n7999_;
  assign n2711_i2 = new_n7991_;
  assign lo585_buf_i2 = new_n3186_;
  assign n2719_i2 = new_n5719_;
  assign n2720_i2 = new_n5720_;
  assign n2723_i2 = new_n5721_;
  assign n2724_i2 = new_n5722_;
  assign n3624_i2 = new_n5723_;
  assign n3625_i2 = new_n5724_;
  assign n3015_i2 = new_n5725_;
  assign n3491_i2 = new_n5726_;
  assign n2696_i2 = new_n5727_;
  assign n2811_i2 = new_n5729_;
  assign n3010_i2 = new_n5731_;
  assign n3012_i2 = new_n5732_;
  assign lo382_buf_i2 = new_n3070_;
  assign lo386_buf_i2 = new_n3072_;
  assign lo390_buf_i2 = new_n3074_;
  assign lo398_buf_i2 = new_n3084_;
  assign lo402_buf_i2 = new_n3086_;
  assign lo406_buf_i2 = new_n3088_;
  assign n3492_i2 = new_n5733_;
  assign lo366_buf_i2 = new_n8004_;
  assign lo374_buf_i2 = new_n8007_;
  assign lo426_buf_i2 = new_n8008_;
  assign lo494_buf_i2 = new_n8003_;
  assign n2653_i2 = new_n5734_;
  assign n2654_i2 = new_n5735_;
  assign n2715_i2 = new_n5736_;
  assign n2740_i2 = new_n5738_;
  assign n2682_i2 = new_n5740_;
  assign n2736_i2 = new_n5741_;
  assign lo508_buf_i2 = new_n2296_;
  assign lo512_buf_i2 = new_n2298_;
  assign lo536_buf_i2 = new_n2310_;
  assign lo576_buf_i2 = new_n2330_;
  assign lo357_buf_i2 = new_n2220_;
  assign lo361_buf_i2 = new_n2222_;
  assign lo417_buf_i2 = new_n2250_;
  assign lo421_buf_i2 = new_n2252_;
  assign lo473_buf_i2 = new_n2278_;
  assign lo477_buf_i2 = new_n2280_;
  assign lo553_buf_i2 = new_n2318_;
  assign lo557_buf_i2 = new_n2320_;
  assign lo573_buf_i2 = new_n2328_;
  assign lo434_buf_i2 = new_n2258_;
  assign lo438_buf_i2 = new_n2260_;
  assign lo466_buf_i2 = new_n2274_;
  assign lo470_buf_i2 = new_n2276_;
  assign lo490_buf_i2 = new_n2286_;
  assign n2657_i2 = new_n5742_;
  assign n2658_i2 = new_n5743_;
  assign n2663_i2 = new_n5744_;
  assign n2664_i2 = new_n5745_;
  assign n2684_i2 = new_n5746_;
  assign n2685_i2 = new_n5747_;
  assign new_n6741_ = new_n3241_;
  assign new_n6742_ = new_n3217_;
  assign new_n6743_ = new_n2896_;
  assign new_n6744_ = new_n6743_;
  assign new_n6745_ = new_n6744_;
  assign new_n6746_ = new_n6744_;
  assign new_n6747_ = new_n6743_;
  assign new_n6748_ = new_n2404_;
  assign new_n6749_ = new_n3307_;
  assign new_n6750_ = new_n2483_;
  assign new_n6751_ = new_n4144_;
  assign new_n6752_ = new_n6751_;
  assign new_n6753_ = new_n6752_;
  assign new_n6754_ = new_n6753_;
  assign new_n6755_ = new_n6752_;
  assign new_n6756_ = new_n6751_;
  assign new_n6757_ = new_n6756_;
  assign new_n6758_ = new_n6756_;
  assign new_n6759_ = new_n3291_;
  assign new_n6760_ = new_n6759_;
  assign new_n6761_ = new_n6760_;
  assign new_n6762_ = new_n6760_;
  assign new_n6763_ = new_n6759_;
  assign new_n6764_ = new_n3290_;
  assign new_n6765_ = new_n6764_;
  assign new_n6766_ = new_n6765_;
  assign new_n6767_ = new_n6765_;
  assign new_n6768_ = new_n6764_;
  assign new_n6769_ = new_n3872_;
  assign new_n6770_ = new_n4183_;
  assign new_n6771_ = new_n3437_;
  assign new_n6772_ = new_n4190_;
  assign new_n6773_ = new_n3856_;
  assign new_n6774_ = new_n3854_;
  assign new_n6775_ = new_n3857_;
  assign new_n6776_ = new_n3855_;
  assign new_n6777_ = new_n3905_;
  assign new_n6778_ = new_n3859_;
  assign new_n6779_ = new_n3904_;
  assign new_n6780_ = new_n3858_;
  assign new_n6781_ = new_n3462_;
  assign new_n6782_ = new_n6781_;
  assign new_n6783_ = new_n3792_;
  assign new_n6784_ = new_n6783_;
  assign new_n6785_ = new_n6784_;
  assign new_n6786_ = new_n6785_;
  assign new_n6787_ = new_n6785_;
  assign new_n6788_ = new_n6784_;
  assign new_n6789_ = new_n6788_;
  assign new_n6790_ = new_n6788_;
  assign new_n6791_ = new_n6783_;
  assign new_n6792_ = new_n6791_;
  assign new_n6793_ = new_n6792_;
  assign new_n6794_ = new_n6792_;
  assign new_n6795_ = new_n6791_;
  assign new_n6796_ = new_n6795_;
  assign new_n6797_ = new_n6795_;
  assign new_n6798_ = new_n3395_;
  assign new_n6799_ = new_n6798_;
  assign new_n6800_ = new_n6799_;
  assign new_n6801_ = new_n6800_;
  assign new_n6802_ = new_n6799_;
  assign new_n6803_ = new_n6798_;
  assign new_n6804_ = new_n6803_;
  assign new_n6805_ = new_n6803_;
  assign new_n6806_ = new_n3386_;
  assign new_n6807_ = new_n6806_;
  assign new_n6808_ = new_n6807_;
  assign new_n6809_ = new_n6808_;
  assign new_n6810_ = new_n6808_;
  assign new_n6811_ = new_n6807_;
  assign new_n6812_ = new_n6811_;
  assign new_n6813_ = new_n6811_;
  assign new_n6814_ = new_n6806_;
  assign new_n6815_ = new_n6814_;
  assign new_n6816_ = new_n6815_;
  assign new_n6817_ = new_n6815_;
  assign new_n6818_ = new_n6814_;
  assign new_n6819_ = new_n6818_;
  assign new_n6820_ = new_n3793_;
  assign new_n6821_ = new_n3394_;
  assign new_n6822_ = new_n6821_;
  assign new_n6823_ = new_n6822_;
  assign new_n6824_ = new_n6823_;
  assign new_n6825_ = new_n6822_;
  assign new_n6826_ = new_n6821_;
  assign new_n6827_ = new_n6826_;
  assign new_n6828_ = new_n6826_;
  assign new_n6829_ = new_n3387_;
  assign new_n6830_ = new_n6829_;
  assign new_n6831_ = new_n6829_;
  assign new_n6832_ = new_n3844_;
  assign new_n6833_ = new_n4229_;
  assign new_n6834_ = new_n6833_;
  assign new_n6835_ = new_n6834_;
  assign new_n6836_ = new_n6833_;
  assign new_n6837_ = new_n3363_;
  assign new_n6838_ = new_n6837_;
  assign new_n6839_ = new_n6838_;
  assign new_n6840_ = new_n6839_;
  assign new_n6841_ = new_n6840_;
  assign new_n6842_ = new_n6840_;
  assign new_n6843_ = new_n6839_;
  assign new_n6844_ = new_n6843_;
  assign new_n6845_ = new_n6843_;
  assign new_n6846_ = new_n6838_;
  assign new_n6847_ = new_n6846_;
  assign new_n6848_ = new_n6846_;
  assign new_n6849_ = new_n6837_;
  assign new_n6850_ = new_n6849_;
  assign new_n6851_ = new_n6850_;
  assign new_n6852_ = new_n6850_;
  assign new_n6853_ = new_n6849_;
  assign new_n6854_ = new_n6853_;
  assign new_n6855_ = new_n6853_;
  assign new_n6856_ = new_n4239_;
  assign new_n6857_ = new_n6856_;
  assign new_n6858_ = new_n6857_;
  assign new_n6859_ = new_n6856_;
  assign new_n6860_ = new_n3362_;
  assign new_n6861_ = new_n6860_;
  assign new_n6862_ = new_n6861_;
  assign new_n6863_ = new_n6862_;
  assign new_n6864_ = new_n6863_;
  assign new_n6865_ = new_n6863_;
  assign new_n6866_ = new_n6862_;
  assign new_n6867_ = new_n6866_;
  assign new_n6868_ = new_n6866_;
  assign new_n6869_ = new_n6861_;
  assign new_n6870_ = new_n6869_;
  assign new_n6871_ = new_n6869_;
  assign new_n6872_ = new_n6860_;
  assign new_n6873_ = new_n6872_;
  assign new_n6874_ = new_n6873_;
  assign new_n6875_ = new_n6873_;
  assign new_n6876_ = new_n6872_;
  assign new_n6877_ = new_n6876_;
  assign new_n6878_ = new_n6876_;
  assign new_n6879_ = new_n3354_;
  assign new_n6880_ = new_n6879_;
  assign new_n6881_ = new_n6880_;
  assign new_n6882_ = new_n6881_;
  assign new_n6883_ = new_n6881_;
  assign new_n6884_ = new_n6880_;
  assign new_n6885_ = new_n6879_;
  assign new_n6886_ = new_n6885_;
  assign new_n6887_ = new_n6885_;
  assign new_n6888_ = new_n2418_;
  assign new_n6889_ = new_n2566_;
  assign new_n6890_ = new_n3355_;
  assign new_n6891_ = new_n6890_;
  assign new_n6892_ = new_n6891_;
  assign new_n6893_ = new_n6892_;
  assign new_n6894_ = new_n6892_;
  assign new_n6895_ = new_n6891_;
  assign new_n6896_ = new_n6890_;
  assign new_n6897_ = new_n6896_;
  assign new_n6898_ = new_n6896_;
  assign new_n6899_ = new_n3445_;
  assign new_n6900_ = new_n3887_;
  assign new_n6901_ = new_n4256_;
  assign new_n6902_ = new_n3371_;
  assign new_n6903_ = new_n6902_;
  assign new_n6904_ = new_n6903_;
  assign new_n6905_ = new_n6904_;
  assign new_n6906_ = new_n6905_;
  assign new_n6907_ = new_n6905_;
  assign new_n6908_ = new_n6904_;
  assign new_n6909_ = new_n6908_;
  assign new_n6910_ = new_n6908_;
  assign new_n6911_ = new_n6903_;
  assign new_n6912_ = new_n6911_;
  assign new_n6913_ = new_n6911_;
  assign new_n6914_ = new_n6902_;
  assign new_n6915_ = new_n6914_;
  assign new_n6916_ = new_n6915_;
  assign new_n6917_ = new_n6915_;
  assign new_n6918_ = new_n6914_;
  assign new_n6919_ = new_n6918_;
  assign new_n6920_ = new_n6918_;
  assign new_n6921_ = new_n3370_;
  assign new_n6922_ = new_n6921_;
  assign new_n6923_ = new_n6922_;
  assign new_n6924_ = new_n6923_;
  assign new_n6925_ = new_n6924_;
  assign new_n6926_ = new_n6924_;
  assign new_n6927_ = new_n6923_;
  assign new_n6928_ = new_n6927_;
  assign new_n6929_ = new_n6927_;
  assign new_n6930_ = new_n6922_;
  assign new_n6931_ = new_n6930_;
  assign new_n6932_ = new_n6930_;
  assign new_n6933_ = new_n6921_;
  assign new_n6934_ = new_n6933_;
  assign new_n6935_ = new_n6934_;
  assign new_n6936_ = new_n6934_;
  assign new_n6937_ = new_n6933_;
  assign new_n6938_ = new_n6937_;
  assign new_n6939_ = new_n6937_;
  assign new_n6940_ = new_n3378_;
  assign new_n6941_ = new_n6940_;
  assign new_n6942_ = new_n6941_;
  assign new_n6943_ = new_n6942_;
  assign new_n6944_ = new_n6942_;
  assign new_n6945_ = new_n6941_;
  assign new_n6946_ = new_n6940_;
  assign new_n6947_ = new_n6946_;
  assign new_n6948_ = new_n6946_;
  assign new_n6949_ = new_n3379_;
  assign new_n6950_ = new_n6949_;
  assign new_n6951_ = new_n6950_;
  assign new_n6952_ = new_n6951_;
  assign new_n6953_ = new_n6951_;
  assign new_n6954_ = new_n6950_;
  assign new_n6955_ = new_n6949_;
  assign new_n6956_ = new_n6955_;
  assign new_n6957_ = new_n6955_;
  assign new_n6958_ = new_n4273_;
  assign new_n6959_ = new_n4280_;
  assign new_n6960_ = new_n4285_;
  assign new_n6961_ = new_n4299_;
  assign new_n6962_ = new_n3521_;
  assign new_n6963_ = new_n6962_;
  assign new_n6964_ = new_n6963_;
  assign new_n6965_ = new_n6962_;
  assign new_n6966_ = new_n4298_;
  assign new_n6967_ = new_n3520_;
  assign new_n6968_ = new_n6967_;
  assign new_n6969_ = new_n6967_;
  assign new_n6970_ = new_n4309_;
  assign new_n6971_ = new_n4306_;
  assign new_n6972_ = new_n4308_;
  assign new_n6973_ = new_n4307_;
  assign new_n6974_ = new_n3408_;
  assign new_n6975_ = new_n3407_;
  assign new_n6976_ = new_n3409_;
  assign new_n6977_ = new_n3406_;
  assign new_n6978_ = new_n3420_;
  assign new_n6979_ = new_n3413_;
  assign new_n6980_ = new_n3421_;
  assign new_n6981_ = new_n3412_;
  assign new_n6982_ = new_n4329_;
  assign new_n6983_ = new_n4324_;
  assign new_n6984_ = new_n4330_;
  assign new_n6985_ = new_n4323_;
  assign new_n6986_ = new_n3882_;
  assign new_n6987_ = new_n3877_;
  assign new_n6988_ = new_n3883_;
  assign new_n6989_ = new_n3876_;
  assign new_n6990_ = new_n3411_;
  assign new_n6991_ = new_n3404_;
  assign new_n6992_ = new_n3410_;
  assign new_n6993_ = new_n3405_;
  assign new_n6994_ = new_n4347_;
  assign new_n6995_ = new_n4342_;
  assign new_n6996_ = new_n4348_;
  assign new_n6997_ = new_n4341_;
  assign new_n6998_ = new_n4358_;
  assign new_n6999_ = new_n3889_;
  assign new_n7000_ = new_n4370_;
  assign new_n7001_ = new_n4367_;
  assign new_n7002_ = new_n3890_;
  assign new_n7003_ = new_n4374_;
  assign new_n7004_ = new_n4373_;
  assign new_n7005_ = new_n3255_;
  assign new_n7006_ = new_n7005_;
  assign new_n7007_ = new_n7006_;
  assign new_n7008_ = new_n7007_;
  assign new_n7009_ = new_n7008_;
  assign new_n7010_ = new_n7008_;
  assign new_n7011_ = new_n7007_;
  assign new_n7012_ = new_n7011_;
  assign new_n7013_ = new_n7011_;
  assign new_n7014_ = new_n7006_;
  assign new_n7015_ = new_n7014_;
  assign new_n7016_ = new_n7014_;
  assign new_n7017_ = new_n7005_;
  assign new_n7018_ = new_n7017_;
  assign new_n7019_ = new_n7018_;
  assign new_n7020_ = new_n7018_;
  assign new_n7021_ = new_n7017_;
  assign new_n7022_ = new_n7021_;
  assign new_n7023_ = new_n7021_;
  assign new_n7024_ = new_n3254_;
  assign new_n7025_ = new_n7024_;
  assign new_n7026_ = new_n7025_;
  assign new_n7027_ = new_n7026_;
  assign new_n7028_ = new_n7027_;
  assign new_n7029_ = new_n7027_;
  assign new_n7030_ = new_n7026_;
  assign new_n7031_ = new_n7030_;
  assign new_n7032_ = new_n7030_;
  assign new_n7033_ = new_n7025_;
  assign new_n7034_ = new_n7033_;
  assign new_n7035_ = new_n7033_;
  assign new_n7036_ = new_n7024_;
  assign new_n7037_ = new_n7036_;
  assign new_n7038_ = new_n7037_;
  assign new_n7039_ = new_n7037_;
  assign new_n7040_ = new_n7036_;
  assign new_n7041_ = new_n7040_;
  assign new_n7042_ = new_n7040_;
  assign new_n7043_ = new_n3263_;
  assign new_n7044_ = new_n7043_;
  assign new_n7045_ = new_n7044_;
  assign new_n7046_ = new_n7045_;
  assign new_n7047_ = new_n7045_;
  assign new_n7048_ = new_n7044_;
  assign new_n7049_ = new_n7043_;
  assign new_n7050_ = new_n7049_;
  assign new_n7051_ = new_n7049_;
  assign new_n7052_ = new_n3016_;
  assign new_n7053_ = new_n3008_;
  assign new_n7054_ = new_n3262_;
  assign new_n7055_ = new_n7054_;
  assign new_n7056_ = new_n7055_;
  assign new_n7057_ = new_n7056_;
  assign new_n7058_ = new_n7056_;
  assign new_n7059_ = new_n7055_;
  assign new_n7060_ = new_n7054_;
  assign new_n7061_ = new_n7060_;
  assign new_n7062_ = new_n7060_;
  assign new_n7063_ = new_n2880_;
  assign new_n7064_ = new_n7063_;
  assign new_n7065_ = new_n7064_;
  assign new_n7066_ = new_n7065_;
  assign new_n7067_ = new_n7066_;
  assign new_n7068_ = new_n7065_;
  assign new_n7069_ = new_n7064_;
  assign new_n7070_ = new_n7069_;
  assign new_n7071_ = new_n7069_;
  assign new_n7072_ = new_n7063_;
  assign new_n7073_ = new_n7072_;
  assign new_n7074_ = new_n7073_;
  assign new_n7075_ = new_n7073_;
  assign new_n7076_ = new_n7072_;
  assign new_n7077_ = new_n7076_;
  assign new_n7078_ = new_n7076_;
  assign new_n7079_ = new_n3271_;
  assign new_n7080_ = new_n7079_;
  assign new_n7081_ = new_n7080_;
  assign new_n7082_ = new_n7081_;
  assign new_n7083_ = new_n7082_;
  assign new_n7084_ = new_n7082_;
  assign new_n7085_ = new_n7081_;
  assign new_n7086_ = new_n7085_;
  assign new_n7087_ = new_n7085_;
  assign new_n7088_ = new_n7080_;
  assign new_n7089_ = new_n7088_;
  assign new_n7090_ = new_n7088_;
  assign new_n7091_ = new_n7079_;
  assign new_n7092_ = new_n7091_;
  assign new_n7093_ = new_n7092_;
  assign new_n7094_ = new_n7092_;
  assign new_n7095_ = new_n7091_;
  assign new_n7096_ = new_n7095_;
  assign new_n7097_ = new_n7095_;
  assign new_n7098_ = new_n3270_;
  assign new_n7099_ = new_n7098_;
  assign new_n7100_ = new_n7099_;
  assign new_n7101_ = new_n7100_;
  assign new_n7102_ = new_n7101_;
  assign new_n7103_ = new_n7101_;
  assign new_n7104_ = new_n7100_;
  assign new_n7105_ = new_n7104_;
  assign new_n7106_ = new_n7104_;
  assign new_n7107_ = new_n7099_;
  assign new_n7108_ = new_n7107_;
  assign new_n7109_ = new_n7107_;
  assign new_n7110_ = new_n7098_;
  assign new_n7111_ = new_n7110_;
  assign new_n7112_ = new_n7111_;
  assign new_n7113_ = new_n7111_;
  assign new_n7114_ = new_n7110_;
  assign new_n7115_ = new_n7114_;
  assign new_n7116_ = new_n7114_;
  assign new_n7117_ = new_n3279_;
  assign new_n7118_ = new_n7117_;
  assign new_n7119_ = new_n7118_;
  assign new_n7120_ = new_n7119_;
  assign new_n7121_ = new_n7119_;
  assign new_n7122_ = new_n7118_;
  assign new_n7123_ = new_n7117_;
  assign new_n7124_ = new_n7123_;
  assign new_n7125_ = new_n7123_;
  assign new_n7126_ = new_n3278_;
  assign new_n7127_ = new_n7126_;
  assign new_n7128_ = new_n7127_;
  assign new_n7129_ = new_n7128_;
  assign new_n7130_ = new_n7128_;
  assign new_n7131_ = new_n7127_;
  assign new_n7132_ = new_n7126_;
  assign new_n7133_ = new_n7132_;
  assign new_n7134_ = new_n7132_;
  assign new_n7135_ = new_n2506_;
  assign new_n7136_ = new_n2522_;
  assign new_n7137_ = new_n4279_;
  assign new_n7138_ = new_n7137_;
  assign new_n7139_ = new_n7138_;
  assign new_n7140_ = new_n7137_;
  assign new_n7141_ = new_n4252_;
  assign new_n7142_ = new_n7141_;
  assign new_n7143_ = new_n7142_;
  assign new_n7144_ = new_n7141_;
  assign new_n7145_ = new_n2442_;
  assign new_n7146_ = new_n2606_;
  assign new_n7147_ = new_n4284_;
  assign new_n7148_ = new_n7147_;
  assign new_n7149_ = new_n7148_;
  assign new_n7150_ = new_n7147_;
  assign new_n7151_ = new_n4255_;
  assign new_n7152_ = new_n7151_;
  assign new_n7153_ = new_n7152_;
  assign new_n7154_ = new_n7151_;
  assign new_n7155_ = new_n2434_;
  assign new_n7156_ = new_n2598_;
  assign new_n7157_ = new_n4291_;
  assign new_n7158_ = new_n7157_;
  assign new_n7159_ = new_n7158_;
  assign new_n7160_ = new_n7157_;
  assign new_n7161_ = new_n4261_;
  assign new_n7162_ = new_n7161_;
  assign new_n7163_ = new_n7162_;
  assign new_n7164_ = new_n7161_;
  assign new_n7165_ = new_n2591_;
  assign new_n7166_ = new_n2583_;
  assign new_n7167_ = new_n4297_;
  assign new_n7168_ = new_n7167_;
  assign new_n7169_ = new_n7168_;
  assign new_n7170_ = new_n7167_;
  assign new_n7171_ = new_n4234_;
  assign new_n7172_ = new_n7171_;
  assign new_n7173_ = new_n7172_;
  assign new_n7174_ = new_n7171_;
  assign new_n7175_ = new_n2976_;
  assign new_n7176_ = new_n3056_;
  assign new_n7177_ = new_n2945_;
  assign new_n7178_ = new_n3025_;
  assign new_n7179_ = new_n2881_;
  assign new_n7180_ = new_n7179_;
  assign new_n7181_ = new_n7179_;
  assign new_n7182_ = new_n2928_;
  assign new_n7183_ = new_n2936_;
  assign new_n7184_ = new_n2912_;
  assign new_n7185_ = new_n2920_;
  assign new_n7186_ = new_n3347_;
  assign new_n7187_ = new_n3346_;
  assign new_n7188_ = new_n2857_;
  assign new_n7189_ = new_n3463_;
  assign new_n7190_ = new_n2856_;
  assign new_n7191_ = new_n4564_;
  assign new_n7192_ = new_n3233_;
  assign new_n7193_ = new_n3083_;
  assign new_n7194_ = new_n4138_;
  assign new_n7195_ = new_n4143_;
  assign new_n7196_ = new_n4202_;
  assign new_n7197_ = new_n4217_;
  assign new_n7198_ = new_n4318_;
  assign new_n7199_ = new_n4357_;
  assign new_n7200_ = new_n2718_;
  assign new_n7201_ = new_n2726_;
  assign new_n7202_ = new_n4597_;
  assign new_n7203_ = new_n7202_;
  assign new_n7204_ = new_n7203_;
  assign new_n7205_ = new_n7202_;
  assign new_n7206_ = new_n4576_;
  assign new_n7207_ = new_n7206_;
  assign new_n7208_ = new_n7207_;
  assign new_n7209_ = new_n7206_;
  assign new_n7210_ = new_n2538_;
  assign new_n7211_ = new_n2530_;
  assign new_n7212_ = new_n4603_;
  assign new_n7213_ = new_n7212_;
  assign new_n7214_ = new_n7213_;
  assign new_n7215_ = new_n7212_;
  assign new_n7216_ = new_n4580_;
  assign new_n7217_ = new_n7216_;
  assign new_n7218_ = new_n7217_;
  assign new_n7219_ = new_n7216_;
  assign new_n7220_ = new_n2710_;
  assign new_n7221_ = new_n2702_;
  assign new_n7222_ = new_n4609_;
  assign new_n7223_ = new_n7222_;
  assign new_n7224_ = new_n7223_;
  assign new_n7225_ = new_n7222_;
  assign new_n7226_ = new_n4584_;
  assign new_n7227_ = new_n7226_;
  assign new_n7228_ = new_n7227_;
  assign new_n7229_ = new_n7226_;
  assign new_n7230_ = new_n2514_;
  assign new_n7231_ = new_n2678_;
  assign new_n7232_ = new_n4613_;
  assign new_n7233_ = new_n7232_;
  assign new_n7234_ = new_n7233_;
  assign new_n7235_ = new_n7232_;
  assign new_n7236_ = new_n4587_;
  assign new_n7237_ = new_n7236_;
  assign new_n7238_ = new_n7237_;
  assign new_n7239_ = new_n7236_;
  assign new_n7240_ = new_n2984_;
  assign new_n7241_ = new_n3064_;
  assign new_n7242_ = new_n2968_;
  assign new_n7243_ = new_n3048_;
  assign new_n7244_ = new_n2960_;
  assign new_n7245_ = new_n3040_;
  assign new_n7246_ = new_n2952_;
  assign new_n7247_ = new_n3032_;
  assign new_n7248_ = new_n4767_;
  assign new_n7249_ = new_n4766_;
  assign new_n7250_ = new_n4772_;
  assign new_n7251_ = new_n2575_;
  assign new_n7252_ = new_n2427_;
  assign new_n7253_ = new_n4780_;
  assign new_n7254_ = new_n7253_;
  assign new_n7255_ = new_n7253_;
  assign new_n7256_ = new_n4783_;
  assign new_n7257_ = new_n7256_;
  assign new_n7258_ = new_n7256_;
  assign new_n7259_ = new_n3001_;
  assign new_n7260_ = new_n2993_;
  assign new_n7261_ = new_n3965_;
  assign new_n7262_ = new_n3619_;
  assign new_n7263_ = new_n7262_;
  assign new_n7264_ = new_n7262_;
  assign new_n7265_ = new_n3964_;
  assign new_n7266_ = new_n7265_;
  assign new_n7267_ = new_n3618_;
  assign new_n7268_ = new_n7267_;
  assign new_n7269_ = new_n4818_;
  assign new_n7270_ = new_n3647_;
  assign new_n7271_ = new_n3555_;
  assign new_n7272_ = new_n7271_;
  assign new_n7273_ = new_n7272_;
  assign new_n7274_ = new_n7271_;
  assign new_n7275_ = new_n2410_;
  assign new_n7276_ = new_n7275_;
  assign new_n7277_ = new_n7275_;
  assign new_n7278_ = new_n4825_;
  assign new_n7279_ = new_n3572_;
  assign new_n7280_ = new_n4083_;
  assign new_n7281_ = new_n4082_;
  assign new_n7282_ = new_n7281_;
  assign new_n7283_ = new_n4053_;
  assign new_n7284_ = new_n4052_;
  assign new_n7285_ = new_n4078_;
  assign new_n7286_ = new_n4088_;
  assign new_n7287_ = new_n4084_;
  assign new_n7288_ = new_n7287_;
  assign new_n7289_ = new_n4085_;
  assign new_n7290_ = new_n4839_;
  assign new_n7291_ = new_n7290_;
  assign new_n7292_ = new_n3938_;
  assign new_n7293_ = new_n7292_;
  assign new_n7294_ = new_n4840_;
  assign new_n7295_ = new_n3939_;
  assign new_n7296_ = new_n3331_;
  assign new_n7297_ = new_n7296_;
  assign new_n7298_ = new_n7297_;
  assign new_n7299_ = new_n7298_;
  assign new_n7300_ = new_n7298_;
  assign new_n7301_ = new_n7297_;
  assign new_n7302_ = new_n7301_;
  assign new_n7303_ = new_n7301_;
  assign new_n7304_ = new_n7296_;
  assign new_n7305_ = new_n7304_;
  assign new_n7306_ = new_n7304_;
  assign new_n7307_ = new_n3312_;
  assign new_n7308_ = new_n7307_;
  assign new_n7309_ = new_n7308_;
  assign new_n7310_ = new_n7309_;
  assign new_n7311_ = new_n7309_;
  assign new_n7312_ = new_n7308_;
  assign new_n7313_ = new_n7312_;
  assign new_n7314_ = new_n7312_;
  assign new_n7315_ = new_n7307_;
  assign new_n7316_ = new_n7315_;
  assign new_n7317_ = new_n7315_;
  assign new_n7318_ = new_n4056_;
  assign new_n7319_ = new_n7318_;
  assign new_n7320_ = new_n7319_;
  assign new_n7321_ = new_n7319_;
  assign new_n7322_ = new_n7318_;
  assign new_n7323_ = new_n3644_;
  assign new_n7324_ = new_n7323_;
  assign new_n7325_ = new_n4057_;
  assign new_n7326_ = new_n7325_;
  assign new_n7327_ = new_n7326_;
  assign new_n7328_ = new_n7325_;
  assign new_n7329_ = new_n3645_;
  assign new_n7330_ = new_n3948_;
  assign new_n7331_ = new_n3764_;
  assign new_n7332_ = new_n4830_;
  assign new_n7333_ = new_n7332_;
  assign new_n7334_ = new_n7332_;
  assign new_n7335_ = new_n4829_;
  assign new_n7336_ = new_n7335_;
  assign new_n7337_ = new_n4025_;
  assign new_n7338_ = new_n4024_;
  assign new_n7339_ = new_n4029_;
  assign new_n7340_ = new_n3988_;
  assign new_n7341_ = new_n7340_;
  assign new_n7342_ = new_n7340_;
  assign new_n7343_ = new_n4028_;
  assign new_n7344_ = new_n3989_;
  assign new_n7345_ = new_n7344_;
  assign new_n7346_ = new_n4834_;
  assign new_n7347_ = new_n7346_;
  assign new_n7348_ = new_n4030_;
  assign new_n7349_ = new_n7348_;
  assign new_n7350_ = new_n7349_;
  assign new_n7351_ = new_n7348_;
  assign new_n7352_ = new_n4833_;
  assign new_n7353_ = new_n4031_;
  assign new_n7354_ = new_n7353_;
  assign new_n7355_ = new_n7353_;
  assign new_n7356_ = new_n4865_;
  assign new_n7357_ = new_n4864_;
  assign new_n7358_ = new_n4826_;
  assign new_n7359_ = new_n4876_;
  assign new_n7360_ = new_n3604_;
  assign new_n7361_ = new_n4086_;
  assign new_n7362_ = new_n7361_;
  assign new_n7363_ = new_n7361_;
  assign new_n7364_ = new_n3936_;
  assign new_n7365_ = new_n7364_;
  assign new_n7366_ = new_n7364_;
  assign new_n7367_ = new_n4087_;
  assign new_n7368_ = new_n3937_;
  assign new_n7369_ = new_n3590_;
  assign new_n7370_ = new_n7369_;
  assign new_n7371_ = new_n3511_;
  assign new_n7372_ = new_n7371_;
  assign new_n7373_ = new_n7371_;
  assign new_n7374_ = new_n3510_;
  assign new_n7375_ = new_n7374_;
  assign new_n7376_ = new_n7374_;
  assign new_n7377_ = new_n3325_;
  assign new_n7378_ = new_n7377_;
  assign new_n7379_ = new_n7378_;
  assign new_n7380_ = new_n7379_;
  assign new_n7381_ = new_n7379_;
  assign new_n7382_ = new_n7378_;
  assign new_n7383_ = new_n7382_;
  assign new_n7384_ = new_n7377_;
  assign new_n7385_ = new_n7384_;
  assign new_n7386_ = new_n7384_;
  assign new_n7387_ = new_n3318_;
  assign new_n7388_ = new_n7387_;
  assign new_n7389_ = new_n7388_;
  assign new_n7390_ = new_n7389_;
  assign new_n7391_ = new_n7389_;
  assign new_n7392_ = new_n7388_;
  assign new_n7393_ = new_n7392_;
  assign new_n7394_ = new_n7387_;
  assign new_n7395_ = new_n7394_;
  assign new_n7396_ = new_n7394_;
  assign new_n7397_ = new_n3453_;
  assign new_n7398_ = new_n7397_;
  assign new_n7399_ = new_n3452_;
  assign new_n7400_ = new_n7399_;
  assign new_n7401_ = new_n3579_;
  assign new_n7402_ = new_n7401_;
  assign new_n7403_ = new_n3578_;
  assign new_n7404_ = new_n7403_;
  assign new_n7405_ = new_n4853_;
  assign new_n7406_ = new_n7405_;
  assign new_n7407_ = new_n3178_;
  assign new_n7408_ = new_n7407_;
  assign new_n7409_ = new_n7408_;
  assign new_n7410_ = new_n7407_;
  assign new_n7411_ = new_n4852_;
  assign new_n7412_ = new_n3179_;
  assign new_n7413_ = new_n7412_;
  assign new_n7414_ = new_n7412_;
  assign new_n7415_ = new_n4910_;
  assign new_n7416_ = new_n4116_;
  assign new_n7417_ = new_n4076_;
  assign new_n7418_ = new_n7417_;
  assign new_n7419_ = new_n7418_;
  assign new_n7420_ = new_n7419_;
  assign new_n7421_ = new_n7419_;
  assign new_n7422_ = new_n7418_;
  assign new_n7423_ = new_n7417_;
  assign new_n7424_ = new_n7423_;
  assign new_n7425_ = new_n7423_;
  assign new_n7426_ = new_n4077_;
  assign new_n7427_ = new_n7426_;
  assign new_n7428_ = new_n7427_;
  assign new_n7429_ = new_n7428_;
  assign new_n7430_ = new_n7427_;
  assign new_n7431_ = new_n7426_;
  assign new_n7432_ = new_n7431_;
  assign new_n7433_ = new_n7431_;
  assign new_n7434_ = new_n4873_;
  assign new_n7435_ = new_n7434_;
  assign new_n7436_ = new_n4112_;
  assign new_n7437_ = new_n7436_;
  assign new_n7438_ = new_n4871_;
  assign new_n7439_ = new_n7438_;
  assign new_n7440_ = new_n4114_;
  assign new_n7441_ = new_n7440_;
  assign new_n7442_ = new_n4124_;
  assign new_n7443_ = new_n7442_;
  assign new_n7444_ = new_n7443_;
  assign new_n7445_ = new_n7444_;
  assign new_n7446_ = new_n7444_;
  assign new_n7447_ = new_n7443_;
  assign new_n7448_ = new_n7447_;
  assign new_n7449_ = new_n7447_;
  assign new_n7450_ = new_n7442_;
  assign new_n7451_ = new_n7450_;
  assign new_n7452_ = new_n7450_;
  assign new_n7453_ = new_n4120_;
  assign new_n7454_ = new_n4125_;
  assign new_n7455_ = new_n7454_;
  assign new_n7456_ = new_n7455_;
  assign new_n7457_ = new_n7456_;
  assign new_n7458_ = new_n7456_;
  assign new_n7459_ = new_n7455_;
  assign new_n7460_ = new_n7459_;
  assign new_n7461_ = new_n7454_;
  assign new_n7462_ = new_n7461_;
  assign new_n7463_ = new_n7461_;
  assign new_n7464_ = new_n4841_;
  assign new_n7465_ = new_n4941_;
  assign new_n7466_ = new_n4868_;
  assign new_n7467_ = new_n7466_;
  assign new_n7468_ = new_n4940_;
  assign new_n7469_ = new_n4869_;
  assign new_n7470_ = new_n4943_;
  assign new_n7471_ = new_n4942_;
  assign new_n7472_ = new_n4098_;
  assign new_n7473_ = new_n4102_;
  assign new_n7474_ = new_n4958_;
  assign new_n7475_ = new_n4831_;
  assign new_n7476_ = new_n7475_;
  assign new_n7477_ = new_n4959_;
  assign new_n7478_ = new_n4832_;
  assign new_n7479_ = new_n7478_;
  assign new_n7480_ = new_n7478_;
  assign new_n7481_ = new_n4854_;
  assign new_n7482_ = new_n7481_;
  assign new_n7483_ = new_n4966_;
  assign new_n7484_ = new_n4106_;
  assign new_n7485_ = new_n4921_;
  assign new_n7486_ = new_n7485_;
  assign new_n7487_ = new_n4094_;
  assign new_n7488_ = new_n7487_;
  assign new_n7489_ = new_n4875_;
  assign new_n7490_ = new_n7489_;
  assign new_n7491_ = new_n4110_;
  assign new_n7492_ = new_n7491_;
  assign new_n7493_ = new_n4924_;
  assign new_n7494_ = new_n7493_;
  assign new_n7495_ = new_n7493_;
  assign new_n7496_ = new_n4090_;
  assign new_n7497_ = new_n4092_;
  assign new_n7498_ = new_n4957_;
  assign new_n7499_ = new_n7498_;
  assign new_n7500_ = new_n3174_;
  assign new_n7501_ = new_n7500_;
  assign new_n7502_ = new_n4951_;
  assign new_n7503_ = new_n7502_;
  assign new_n7504_ = new_n3182_;
  assign new_n7505_ = new_n7504_;
  assign new_n7506_ = new_n4971_;
  assign new_n7507_ = new_n7506_;
  assign new_n7508_ = new_n3184_;
  assign new_n7509_ = new_n7508_;
  assign new_n7510_ = new_n4932_;
  assign new_n7511_ = new_n7510_;
  assign new_n7512_ = new_n4096_;
  assign new_n7513_ = new_n7512_;
  assign new_n7514_ = new_n4998_;
  assign new_n7515_ = new_n4984_;
  assign new_n7516_ = new_n7515_;
  assign new_n7517_ = new_n4982_;
  assign new_n7518_ = new_n3393_;
  assign new_n7519_ = new_n7518_;
  assign new_n7520_ = new_n7519_;
  assign new_n7521_ = new_n7520_;
  assign new_n7522_ = new_n7520_;
  assign new_n7523_ = new_n7519_;
  assign new_n7524_ = new_n7523_;
  assign new_n7525_ = new_n7518_;
  assign new_n7526_ = new_n7525_;
  assign new_n7527_ = new_n7525_;
  assign new_n7528_ = new_n3392_;
  assign new_n7529_ = new_n7528_;
  assign new_n7530_ = new_n7529_;
  assign new_n7531_ = new_n7530_;
  assign new_n7532_ = new_n7530_;
  assign new_n7533_ = new_n7529_;
  assign new_n7534_ = new_n7533_;
  assign new_n7535_ = new_n7533_;
  assign new_n7536_ = new_n7528_;
  assign new_n7537_ = new_n7536_;
  assign new_n7538_ = new_n7537_;
  assign new_n7539_ = new_n7537_;
  assign new_n7540_ = new_n7536_;
  assign new_n7541_ = new_n3455_;
  assign new_n7542_ = new_n7541_;
  assign new_n7543_ = new_n3454_;
  assign new_n7544_ = new_n7543_;
  assign new_n7545_ = new_n3385_;
  assign new_n7546_ = new_n7545_;
  assign new_n7547_ = new_n2806_;
  assign new_n7548_ = new_n3384_;
  assign new_n7549_ = new_n7548_;
  assign new_n7550_ = new_n3607_;
  assign new_n7551_ = new_n3608_;
  assign new_n7552_ = new_n7551_;
  assign new_n7553_ = new_n3606_;
  assign new_n7554_ = new_n3628_;
  assign new_n7555_ = new_n4020_;
  assign new_n7556_ = new_n3980_;
  assign new_n7557_ = new_n4021_;
  assign new_n7558_ = new_n3981_;
  assign new_n7559_ = new_n5030_;
  assign new_n7560_ = new_n5023_;
  assign new_n7561_ = new_n5029_;
  assign new_n7562_ = new_n5024_;
  assign new_n7563_ = new_n3554_;
  assign new_n7564_ = new_n5042_;
  assign new_n7565_ = new_n4821_;
  assign new_n7566_ = new_n7565_;
  assign new_n7567_ = new_n5041_;
  assign new_n7568_ = new_n4822_;
  assign new_n7569_ = new_n7568_;
  assign new_n7570_ = new_n4909_;
  assign new_n7571_ = new_n4891_;
  assign new_n7572_ = new_n4900_;
  assign new_n7573_ = new_n5062_;
  assign new_n7574_ = new_n5059_;
  assign new_n7575_ = new_n5061_;
  assign new_n7576_ = new_n5060_;
  assign new_n7577_ = new_n4002_;
  assign new_n7578_ = new_n3998_;
  assign new_n7579_ = new_n5071_;
  assign new_n7580_ = new_n5069_;
  assign new_n7581_ = new_n5072_;
  assign new_n7582_ = new_n5070_;
  assign new_n7583_ = new_n3942_;
  assign new_n7584_ = new_n7583_;
  assign new_n7585_ = new_n7583_;
  assign new_n7586_ = new_n3943_;
  assign new_n7587_ = new_n7586_;
  assign new_n7588_ = new_n2411_;
  assign new_n7589_ = new_n3941_;
  assign new_n7590_ = new_n7589_;
  assign new_n7591_ = new_n7589_;
  assign new_n7592_ = new_n3940_;
  assign new_n7593_ = new_n7592_;
  assign new_n7594_ = new_n7593_;
  assign new_n7595_ = new_n7592_;
  assign new_n7596_ = new_n5089_;
  assign new_n7597_ = new_n7596_;
  assign new_n7598_ = new_n7597_;
  assign new_n7599_ = new_n7596_;
  assign new_n7600_ = new_n5088_;
  assign new_n7601_ = new_n7600_;
  assign new_n7602_ = new_n7601_;
  assign new_n7603_ = new_n7600_;
  assign new_n7604_ = new_n3716_;
  assign new_n7605_ = new_n3717_;
  assign new_n7606_ = new_n7605_;
  assign new_n7607_ = new_n5094_;
  assign new_n7608_ = new_n4877_;
  assign new_n7609_ = new_n3148_;
  assign new_n7610_ = new_n7609_;
  assign new_n7611_ = new_n5101_;
  assign new_n7612_ = new_n3616_;
  assign new_n7613_ = new_n4823_;
  assign new_n7614_ = new_n5108_;
  assign new_n7615_ = new_n4882_;
  assign new_n7616_ = new_n3582_;
  assign new_n7617_ = new_n5113_;
  assign new_n7618_ = new_n3126_;
  assign new_n7619_ = new_n3979_;
  assign new_n7620_ = new_n7619_;
  assign new_n7621_ = new_n4847_;
  assign new_n7622_ = new_n3476_;
  assign new_n7623_ = new_n7622_;
  assign new_n7624_ = new_n3477_;
  assign new_n7625_ = new_n7624_;
  assign new_n7626_ = new_n3450_;
  assign new_n7627_ = new_n7626_;
  assign new_n7628_ = new_n3451_;
  assign new_n7629_ = new_n7628_;
  assign new_n7630_ = new_n3478_;
  assign new_n7631_ = new_n7630_;
  assign new_n7632_ = new_n3479_;
  assign new_n7633_ = new_n7632_;
  assign new_n7634_ = new_n3471_;
  assign new_n7635_ = new_n7634_;
  assign new_n7636_ = new_n7634_;
  assign new_n7637_ = new_n3470_;
  assign new_n7638_ = new_n7637_;
  assign new_n7639_ = new_n7637_;
  assign new_n7640_ = new_n3595_;
  assign new_n7641_ = new_n7640_;
  assign new_n7642_ = new_n7640_;
  assign new_n7643_ = new_n3594_;
  assign new_n7644_ = new_n7643_;
  assign new_n7645_ = new_n7643_;
  assign new_n7646_ = new_n3513_;
  assign new_n7647_ = new_n7646_;
  assign new_n7648_ = new_n3512_;
  assign new_n7649_ = new_n7648_;
  assign new_n7650_ = new_n3497_;
  assign new_n7651_ = new_n7650_;
  assign new_n7652_ = new_n3496_;
  assign new_n7653_ = new_n7652_;
  assign new_n7654_ = new_n3970_;
  assign new_n7655_ = new_n3969_;
  assign new_n7656_ = new_n3971_;
  assign new_n7657_ = new_n3968_;
  assign new_n7658_ = new_n3977_;
  assign new_n7659_ = new_n3978_;
  assign new_n7660_ = new_n7659_;
  assign new_n7661_ = new_n3976_;
  assign new_n7662_ = new_n5209_;
  assign new_n7663_ = new_n5204_;
  assign new_n7664_ = new_n5210_;
  assign new_n7665_ = new_n5203_;
  assign new_n7666_ = new_n3974_;
  assign new_n7667_ = new_n3967_;
  assign new_n7668_ = new_n3975_;
  assign new_n7669_ = new_n3966_;
  assign new_n7670_ = new_n4019_;
  assign new_n7671_ = new_n3973_;
  assign new_n7672_ = new_n4018_;
  assign new_n7673_ = new_n3972_;
  assign new_n7674_ = new_n5228_;
  assign new_n7675_ = new_n5221_;
  assign new_n7676_ = new_n5227_;
  assign new_n7677_ = new_n5222_;
  assign new_n7678_ = new_n3456_;
  assign new_n7679_ = new_n3098_;
  assign new_n7680_ = new_n7679_;
  assign new_n7681_ = new_n3457_;
  assign new_n7682_ = new_n3099_;
  assign new_n7683_ = new_n7682_;
  assign new_n7684_ = new_n3614_;
  assign new_n7685_ = new_n3626_;
  assign new_n7686_ = new_n3678_;
  assign new_n7687_ = new_n5282_;
  assign new_n7688_ = new_n5279_;
  assign new_n7689_ = new_n3540_;
  assign new_n7690_ = new_n3149_;
  assign new_n7691_ = new_n3541_;
  assign new_n7692_ = new_n5296_;
  assign new_n7693_ = new_n5293_;
  assign new_n7694_ = new_n5304_;
  assign new_n7695_ = new_n5301_;
  assign new_n7696_ = new_n5325_;
  assign new_n7697_ = new_n5322_;
  assign new_n7698_ = new_n5324_;
  assign new_n7699_ = new_n5323_;
  assign new_n7700_ = new_n3247_;
  assign new_n7701_ = new_n7700_;
  assign new_n7702_ = new_n7700_;
  assign new_n7703_ = new_n3246_;
  assign new_n7704_ = new_n7703_;
  assign new_n7705_ = new_n7703_;
  assign new_n7706_ = new_n5336_;
  assign new_n7707_ = new_n5334_;
  assign new_n7708_ = new_n5337_;
  assign new_n7709_ = new_n5335_;
  assign new_n7710_ = new_n5349_;
  assign new_n7711_ = new_n5348_;
  assign new_n7712_ = new_n5354_;
  assign new_n7713_ = new_n5355_;
  assign new_n7714_ = new_n4981_;
  assign new_n7715_ = new_n7714_;
  assign new_n7716_ = new_n4976_;
  assign new_n7717_ = new_n4922_;
  assign new_n7718_ = new_n4063_;
  assign new_n7719_ = new_n7718_;
  assign new_n7720_ = new_n7719_;
  assign new_n7721_ = new_n7720_;
  assign new_n7722_ = new_n7720_;
  assign new_n7723_ = new_n7719_;
  assign new_n7724_ = new_n7723_;
  assign new_n7725_ = new_n7723_;
  assign new_n7726_ = new_n7718_;
  assign new_n7727_ = new_n7726_;
  assign new_n7728_ = new_n7727_;
  assign new_n7729_ = new_n7727_;
  assign new_n7730_ = new_n7726_;
  assign new_n7731_ = new_n7730_;
  assign new_n7732_ = new_n7730_;
  assign new_n7733_ = new_n3655_;
  assign new_n7734_ = new_n4065_;
  assign new_n7735_ = new_n7734_;
  assign new_n7736_ = new_n7735_;
  assign new_n7737_ = new_n7736_;
  assign new_n7738_ = new_n7736_;
  assign new_n7739_ = new_n7735_;
  assign new_n7740_ = new_n7739_;
  assign new_n7741_ = new_n7739_;
  assign new_n7742_ = new_n7734_;
  assign new_n7743_ = new_n7742_;
  assign new_n7744_ = new_n7743_;
  assign new_n7745_ = new_n7743_;
  assign new_n7746_ = new_n7742_;
  assign new_n7747_ = new_n7746_;
  assign new_n7748_ = new_n3654_;
  assign new_n7749_ = new_n7748_;
  assign new_n7750_ = new_n4066_;
  assign new_n7751_ = new_n7750_;
  assign new_n7752_ = new_n7751_;
  assign new_n7753_ = new_n7752_;
  assign new_n7754_ = new_n7752_;
  assign new_n7755_ = new_n7751_;
  assign new_n7756_ = new_n7755_;
  assign new_n7757_ = new_n7755_;
  assign new_n7758_ = new_n7750_;
  assign new_n7759_ = new_n7758_;
  assign new_n7760_ = new_n7759_;
  assign new_n7761_ = new_n7759_;
  assign new_n7762_ = new_n7758_;
  assign new_n7763_ = new_n4060_;
  assign new_n7764_ = new_n7763_;
  assign new_n7765_ = new_n7764_;
  assign new_n7766_ = new_n7765_;
  assign new_n7767_ = new_n7765_;
  assign new_n7768_ = new_n7764_;
  assign new_n7769_ = new_n7768_;
  assign new_n7770_ = new_n7768_;
  assign new_n7771_ = new_n7763_;
  assign new_n7772_ = new_n7771_;
  assign new_n7773_ = new_n7772_;
  assign new_n7774_ = new_n7772_;
  assign new_n7775_ = new_n7771_;
  assign new_n7776_ = new_n7775_;
  assign new_n7777_ = new_n3665_;
  assign new_n7778_ = new_n3664_;
  assign new_n7779_ = new_n7778_;
  assign new_n7780_ = new_n3752_;
  assign new_n7781_ = new_n3958_;
  assign new_n7782_ = new_n3108_;
  assign new_n7783_ = new_n7782_;
  assign new_n7784_ = new_n3090_;
  assign new_n7785_ = new_n3130_;
  assign new_n7786_ = new_n3132_;
  assign new_n7787_ = new_n4050_;
  assign new_n7788_ = new_n7787_;
  assign new_n7789_ = new_n7787_;
  assign new_n7790_ = new_n4051_;
  assign new_n7791_ = new_n7790_;
  assign new_n7792_ = new_n7790_;
  assign new_n7793_ = new_n4022_;
  assign new_n7794_ = new_n5424_;
  assign new_n7795_ = new_n7794_;
  assign new_n7796_ = new_n4914_;
  assign new_n7797_ = new_n7796_;
  assign new_n7798_ = new_n4879_;
  assign new_n7799_ = new_n4049_;
  assign new_n7800_ = new_n7799_;
  assign new_n7801_ = new_n7799_;
  assign new_n7802_ = new_n5427_;
  assign new_n7803_ = new_n4915_;
  assign new_n7804_ = new_n7803_;
  assign new_n7805_ = new_n7803_;
  assign new_n7806_ = new_n3741_;
  assign new_n7807_ = new_n3740_;
  assign new_n7808_ = new_n7807_;
  assign new_n7809_ = new_n5433_;
  assign new_n7810_ = new_n3911_;
  assign new_n7811_ = new_n7810_;
  assign new_n7812_ = new_n5434_;
  assign new_n7813_ = new_n3910_;
  assign new_n7814_ = new_n7813_;
  assign new_n7815_ = new_n7813_;
  assign new_n7816_ = new_n3954_;
  assign new_n7817_ = new_n3742_;
  assign new_n7818_ = new_n4048_;
  assign new_n7819_ = new_n7818_;
  assign new_n7820_ = new_n7818_;
  assign new_n7821_ = new_n5444_;
  assign new_n7822_ = new_n7821_;
  assign new_n7823_ = new_n5423_;
  assign new_n7824_ = new_n7823_;
  assign new_n7825_ = new_n5443_;
  assign new_n7826_ = new_n7825_;
  assign new_n7827_ = new_n5453_;
  assign new_n7828_ = new_n5457_;
  assign new_n7829_ = new_n4838_;
  assign new_n7830_ = new_n7829_;
  assign new_n7831_ = new_n5458_;
  assign new_n7832_ = new_n4837_;
  assign new_n7833_ = new_n3745_;
  assign new_n7834_ = new_n5464_;
  assign new_n7835_ = new_n3744_;
  assign new_n7836_ = new_n7835_;
  assign new_n7837_ = new_n7835_;
  assign new_n7838_ = new_n5465_;
  assign new_n7839_ = new_n4843_;
  assign new_n7840_ = new_n5472_;
  assign new_n7841_ = new_n3746_;
  assign new_n7842_ = new_n7841_;
  assign new_n7843_ = new_n5471_;
  assign new_n7844_ = new_n3747_;
  assign new_n7845_ = new_n5478_;
  assign new_n7846_ = new_n7845_;
  assign new_n7847_ = new_n5468_;
  assign new_n7848_ = new_n5373_;
  assign new_n7849_ = new_n4999_;
  assign new_n7850_ = new_n4995_;
  assign new_n7851_ = new_n3656_;
  assign new_n7852_ = new_n3114_;
  assign new_n7853_ = new_n3643_;
  assign new_n7854_ = new_n3642_;
  assign new_n7855_ = new_n7854_;
  assign new_n7856_ = new_n3666_;
  assign new_n7857_ = new_n3641_;
  assign new_n7858_ = new_n3640_;
  assign new_n7859_ = new_n7858_;
  assign new_n7860_ = new_n3668_;
  assign new_n7861_ = new_n3639_;
  assign new_n7862_ = new_n3638_;
  assign new_n7863_ = new_n7862_;
  assign new_n7864_ = new_n3670_;
  assign new_n7865_ = new_n3653_;
  assign new_n7866_ = new_n3652_;
  assign new_n7867_ = new_n7866_;
  assign new_n7868_ = new_n3698_;
  assign new_n7869_ = new_n3663_;
  assign new_n7870_ = new_n3662_;
  assign new_n7871_ = new_n7870_;
  assign new_n7872_ = new_n3724_;
  assign new_n7873_ = new_n3661_;
  assign new_n7874_ = new_n3660_;
  assign new_n7875_ = new_n7874_;
  assign new_n7876_ = new_n3726_;
  assign new_n7877_ = new_n3749_;
  assign new_n7878_ = new_n3748_;
  assign new_n7879_ = new_n7878_;
  assign new_n7880_ = new_n4859_;
  assign new_n7881_ = new_n7880_;
  assign new_n7882_ = new_n4858_;
  assign new_n7883_ = new_n5565_;
  assign new_n7884_ = new_n3908_;
  assign new_n7885_ = new_n5564_;
  assign new_n7886_ = new_n3909_;
  assign new_n7887_ = new_n5574_;
  assign new_n7888_ = new_n5559_;
  assign new_n7889_ = new_n3066_;
  assign new_n7890_ = new_n4933_;
  assign new_n7891_ = new_n5587_;
  assign new_n7892_ = new_n5584_;
  assign new_n7893_ = new_n5000_;
  assign new_n7894_ = new_n4925_;
  assign new_n7895_ = new_n7894_;
  assign new_n7896_ = new_n5590_;
  assign new_n7897_ = new_n5376_;
  assign new_n7898_ = new_n7897_;
  assign new_n7899_ = new_n5400_;
  assign new_n7900_ = new_n7899_;
  assign new_n7901_ = new_n5385_;
  assign new_n7902_ = new_n7901_;
  assign new_n7903_ = new_n5403_;
  assign new_n7904_ = new_n7903_;
  assign new_n7905_ = new_n5394_;
  assign new_n7906_ = new_n7905_;
  assign new_n7907_ = new_n3926_;
  assign new_n7908_ = new_n7907_;
  assign new_n7909_ = new_n4062_;
  assign new_n7910_ = new_n7909_;
  assign new_n7911_ = new_n7910_;
  assign new_n7912_ = new_n7909_;
  assign new_n7913_ = new_n3927_;
  assign new_n7914_ = new_n4061_;
  assign new_n7915_ = new_n7914_;
  assign new_n7916_ = new_n7915_;
  assign new_n7917_ = new_n7914_;
  assign new_n7918_ = new_n3961_;
  assign new_n7919_ = new_n7918_;
  assign new_n7920_ = new_n7918_;
  assign new_n7921_ = new_n3960_;
  assign new_n7922_ = new_n7921_;
  assign new_n7923_ = new_n7922_;
  assign new_n7924_ = new_n7921_;
  assign new_n7925_ = new_n4064_;
  assign new_n7926_ = new_n7925_;
  assign new_n7927_ = new_n7925_;
  assign new_n7928_ = new_n4067_;
  assign new_n7929_ = new_n7928_;
  assign new_n7930_ = new_n7928_;
  assign new_n7931_ = new_n5622_;
  assign new_n7932_ = new_n5397_;
  assign new_n7933_ = new_n7932_;
  assign new_n7934_ = new_n3695_;
  assign new_n7935_ = new_n3694_;
  assign new_n7936_ = new_n7935_;
  assign new_n7937_ = new_n3756_;
  assign new_n7938_ = new_n3720_;
  assign new_n7939_ = new_n7938_;
  assign new_n7940_ = new_n3721_;
  assign new_n7941_ = new_n3928_;
  assign new_n7942_ = new_n5642_;
  assign new_n7943_ = new_n5633_;
  assign new_n7944_ = new_n3956_;
  assign new_n7945_ = new_n4968_;
  assign new_n7946_ = new_n4945_;
  assign new_n7947_ = new_n4835_;
  assign new_n7948_ = new_n4828_;
  assign new_n7949_ = new_n7948_;
  assign new_n7950_ = new_n4836_;
  assign new_n7951_ = new_n7950_;
  assign new_n7952_ = new_n4827_;
  assign new_n7953_ = new_n3719_;
  assign new_n7954_ = new_n7953_;
  assign new_n7955_ = new_n7953_;
  assign new_n7956_ = new_n3718_;
  assign new_n7957_ = new_n7956_;
  assign new_n7958_ = new_n7957_;
  assign new_n7959_ = new_n7956_;
  assign new_n7960_ = new_n3924_;
  assign new_n7961_ = new_n7960_;
  assign new_n7962_ = new_n3925_;
  assign new_n7963_ = new_n3283_;
  assign new_n7964_ = new_n4863_;
  assign new_n7965_ = new_n3282_;
  assign new_n7966_ = new_n4974_;
  assign new_n7967_ = new_n5415_;
  assign new_n7968_ = new_n3190_;
  assign new_n7969_ = new_n4990_;
  assign new_n7970_ = new_n3192_;
  assign new_n7971_ = new_n5416_;
  assign new_n7972_ = new_n3118_;
  assign new_n7973_ = new_n3122_;
  assign new_n7974_ = new_n5591_;
  assign new_n7975_ = new_n7974_;
  assign new_n7976_ = new_n5420_;
  assign new_n7977_ = new_n7976_;
  assign new_n7978_ = new_n7976_;
  assign new_n7979_ = new_n5456_;
  assign new_n7980_ = new_n7979_;
  assign new_n7981_ = new_n5481_;
  assign new_n7982_ = new_n5418_;
  assign new_n7983_ = new_n5375_;
  assign new_n7984_ = new_n4991_;
  assign new_n7985_ = new_n4993_;
  assign new_n7986_ = new_n5483_;
  assign new_n7987_ = new_n5579_;
  assign new_n7988_ = new_n7987_;
  assign new_n7989_ = new_n3180_;
  assign new_n7990_ = new_n7989_;
  assign new_n7991_ = new_n5718_;
  assign new_n7992_ = new_n5582_;
  assign new_n7993_ = new_n5117_;
  assign new_n7994_ = new_n3188_;
  assign new_n7995_ = new_n5583_;
  assign new_n7996_ = new_n5409_;
  assign new_n7997_ = new_n3172_;
  assign new_n7998_ = new_n5714_;
  assign new_n7999_ = new_n5716_;
  assign new_n8000_ = new_n5715_;
  assign new_n8001_ = new_n2288_;
  assign new_n8002_ = new_n8001_;
  assign new_n8003_ = new_n8001_;
  assign new_n8004_ = new_n2224_;
  assign new_n8005_ = new_n2289_;
  assign new_n8006_ = new_n8005_;
  assign new_n8007_ = new_n2228_;
  assign new_n8008_ = new_n2254_;
  assign new_n8009_ = new_n3201_;
  assign new_n8010_ = new_n8009_;
  assign new_n8011_ = new_n3208_;
  assign new_n8012_ = new_n2405_;
  assign new_n8013_ = new_n8012_;
  assign new_n8014_ = new_n8012_;
  assign new_n8015_ = new_n3117_;
  assign new_n8016_ = new_n4153_;
  assign new_n8017_ = new_n4191_;
  assign new_n8018_ = new_n4195_;
  assign new_n8019_ = new_n4223_;
  assign new_n8020_ = new_n4224_;
  always @ (posedge clock) begin
    n2610_lo <= n7230_li000_li000;
    n2613_lo <= n7233_li001_li001;
    n2616_lo <= n7236_li002_li002;
    n2619_lo <= n7239_li003_li003;
    n2622_lo <= n7242_li004_li004;
    n2625_lo <= n7245_li005_li005;
    n2628_lo <= n7248_li006_li006;
    n2634_lo <= n7254_li008_li008;
    n2637_lo <= n7257_li009_li009;
    n2640_lo <= n7260_li010_li010;
    n2643_lo <= n7263_li011_li011;
    n2646_lo <= n7266_li012_li012;
    n2649_lo <= n7269_li013_li013;
    n2652_lo <= n7272_li014_li014;
    n2655_lo <= n7275_li015_li015;
    n2658_lo <= n7278_li016_li016;
    n2661_lo <= n7281_li017_li017;
    n2664_lo <= n7284_li018_li018;
    n2667_lo <= n7287_li019_li019;
    n2670_lo <= n7290_li020_li020;
    n2673_lo <= n7293_li021_li021;
    n2676_lo <= n7296_li022_li022;
    n2679_lo <= n7299_li023_li023;
    n2682_lo <= n7302_li024_li024;
    n2685_lo <= n7305_li025_li025;
    n2688_lo <= n7308_li026_li026;
    n2691_lo <= n7311_li027_li027;
    n2694_lo <= n7314_li028_li028;
    n2697_lo <= n7317_li029_li029;
    n2700_lo <= n7320_li030_li030;
    n2703_lo <= n7323_li031_li031;
    n2706_lo <= n7326_li032_li032;
    n2709_lo <= n7329_li033_li033;
    n2712_lo <= n7332_li034_li034;
    n2715_lo <= n7335_li035_li035;
    n2718_lo <= n7338_li036_li036;
    n2721_lo <= n7341_li037_li037;
    n2724_lo <= n7344_li038_li038;
    n2727_lo <= n7347_li039_li039;
    n2730_lo <= n7350_li040_li040;
    n2733_lo <= n7353_li041_li041;
    n2736_lo <= n7356_li042_li042;
    n2739_lo <= n7359_li043_li043;
    n2742_lo <= n7362_li044_li044;
    n2745_lo <= n7365_li045_li045;
    n2748_lo <= n7368_li046_li046;
    n2751_lo <= n7371_li047_li047;
    n2754_lo <= n7374_li048_li048;
    n2757_lo <= n7377_li049_li049;
    n2760_lo <= n7380_li050_li050;
    n2763_lo <= n7383_li051_li051;
    n2766_lo <= n7386_li052_li052;
    n2769_lo <= n7389_li053_li053;
    n2772_lo <= n7392_li054_li054;
    n2775_lo <= n7395_li055_li055;
    n2778_lo <= n7398_li056_li056;
    n2781_lo <= n7401_li057_li057;
    n2784_lo <= n7404_li058_li058;
    n2787_lo <= n7407_li059_li059;
    n2790_lo <= n7410_li060_li060;
    n2793_lo <= n7413_li061_li061;
    n2796_lo <= n7416_li062_li062;
    n2799_lo <= n7419_li063_li063;
    n2802_lo <= n7422_li064_li064;
    n2805_lo <= n7425_li065_li065;
    n2808_lo <= n7428_li066_li066;
    n2811_lo <= n7431_li067_li067;
    n2814_lo <= n7434_li068_li068;
    n2817_lo <= n7437_li069_li069;
    n2820_lo <= n7440_li070_li070;
    n2823_lo <= n7443_li071_li071;
    n2826_lo <= n7446_li072_li072;
    n2829_lo <= n7449_li073_li073;
    n2832_lo <= n7452_li074_li074;
    n2838_lo <= n7458_li076_li076;
    n2841_lo <= n7461_li077_li077;
    n2844_lo <= n7464_li078_li078;
    n2847_lo <= n7467_li079_li079;
    n2850_lo <= n7470_li080_li080;
    n2853_lo <= n7473_li081_li081;
    n2856_lo <= n7476_li082_li082;
    n2862_lo <= n7482_li084_li084;
    n2865_lo <= n7485_li085_li085;
    n2868_lo <= n7488_li086_li086;
    n2871_lo <= n7491_li087_li087;
    n2874_lo <= n7494_li088_li088;
    n2877_lo <= n7497_li089_li089;
    n2880_lo <= n7500_li090_li090;
    n2883_lo <= n7503_li091_li091;
    n2886_lo <= n7506_li092_li092;
    n2889_lo <= n7509_li093_li093;
    n2892_lo <= n7512_li094_li094;
    n2895_lo <= n7515_li095_li095;
    n2898_lo <= n7518_li096_li096;
    n2901_lo <= n7521_li097_li097;
    n2904_lo <= n7524_li098_li098;
    n2907_lo <= n7527_li099_li099;
    n2910_lo <= n7530_li100_li100;
    n2913_lo <= n7533_li101_li101;
    n2916_lo <= n7536_li102_li102;
    n2919_lo <= n7539_li103_li103;
    n2922_lo <= n7542_li104_li104;
    n2925_lo <= n7545_li105_li105;
    n2928_lo <= n7548_li106_li106;
    n2931_lo <= n7551_li107_li107;
    n2934_lo <= n7554_li108_li108;
    n2937_lo <= n7557_li109_li109;
    n2940_lo <= n7560_li110_li110;
    n2943_lo <= n7563_li111_li111;
    n2946_lo <= n7566_li112_li112;
    n2949_lo <= n7569_li113_li113;
    n2952_lo <= n7572_li114_li114;
    n2955_lo <= n7575_li115_li115;
    n2958_lo <= n7578_li116_li116;
    n2961_lo <= n7581_li117_li117;
    n2964_lo <= n7584_li118_li118;
    n2967_lo <= n7587_li119_li119;
    n2970_lo <= n7590_li120_li120;
    n2973_lo <= n7593_li121_li121;
    n2976_lo <= n7596_li122_li122;
    n2979_lo <= n7599_li123_li123;
    n2982_lo <= n7602_li124_li124;
    n2985_lo <= n7605_li125_li125;
    n2988_lo <= n7608_li126_li126;
    n2991_lo <= n7611_li127_li127;
    n2994_lo <= n7614_li128_li128;
    n2997_lo <= n7617_li129_li129;
    n3000_lo <= n7620_li130_li130;
    n3003_lo <= n7623_li131_li131;
    n3006_lo <= n7626_li132_li132;
    n3009_lo <= n7629_li133_li133;
    n3012_lo <= n7632_li134_li134;
    n3015_lo <= n7635_li135_li135;
    n3018_lo <= n7638_li136_li136;
    n3021_lo <= n7641_li137_li137;
    n3024_lo <= n7644_li138_li138;
    n3027_lo <= n7647_li139_li139;
    n3030_lo <= n7650_li140_li140;
    n3033_lo <= n7653_li141_li141;
    n3036_lo <= n7656_li142_li142;
    n3039_lo <= n7659_li143_li143;
    n3042_lo <= n7662_li144_li144;
    n3045_lo <= n7665_li145_li145;
    n3048_lo <= n7668_li146_li146;
    n3051_lo <= n7671_li147_li147;
    n3054_lo <= n7674_li148_li148;
    n3057_lo <= n7677_li149_li149;
    n3060_lo <= n7680_li150_li150;
    n3063_lo <= n7683_li151_li151;
    n3066_lo <= n7686_li152_li152;
    n3069_lo <= n7689_li153_li153;
    n3072_lo <= n7692_li154_li154;
    n3075_lo <= n7695_li155_li155;
    n3078_lo <= n7698_li156_li156;
    n3081_lo <= n7701_li157_li157;
    n3084_lo <= n7704_li158_li158;
    n3087_lo <= n7707_li159_li159;
    n3090_lo <= n7710_li160_li160;
    n3093_lo <= n7713_li161_li161;
    n3096_lo <= n7716_li162_li162;
    n3099_lo <= n7719_li163_li163;
    n3102_lo <= n7722_li164_li164;
    n3105_lo <= n7725_li165_li165;
    n3108_lo <= n7728_li166_li166;
    n3111_lo <= n7731_li167_li167;
    n3114_lo <= n7734_li168_li168;
    n3117_lo <= n7737_li169_li169;
    n3120_lo <= n7740_li170_li170;
    n3126_lo <= n7746_li172_li172;
    n3129_lo <= n7749_li173_li173;
    n3132_lo <= n7752_li174_li174;
    n3138_lo <= n7758_li176_li176;
    n3141_lo <= n7761_li177_li177;
    n3144_lo <= n7764_li178_li178;
    n3147_lo <= n7767_li179_li179;
    n3150_lo <= n7770_li180_li180;
    n3153_lo <= n7773_li181_li181;
    n3156_lo <= n7776_li182_li182;
    n3162_lo <= n7782_li184_li184;
    n3165_lo <= n7785_li185_li185;
    n3168_lo <= n7788_li186_li186;
    n3174_lo <= n7794_li188_li188;
    n3177_lo <= n7797_li189_li189;
    n3180_lo <= n7800_li190_li190;
    n3186_lo <= n7806_li192_li192;
    n3189_lo <= n7809_li193_li193;
    n3192_lo <= n7812_li194_li194;
    n3195_lo <= n7815_li195_li195;
    n3198_lo <= n7818_li196_li196;
    n3201_lo <= n7821_li197_li197;
    n3204_lo <= n7824_li198_li198;
    n3210_lo <= n7830_li200_li200;
    n3213_lo <= n7833_li201_li201;
    n3216_lo <= n7836_li202_li202;
    n3219_lo <= n7839_li203_li203;
    n3222_lo <= n7842_li204_li204;
    n3225_lo <= n7845_li205_li205;
    n3228_lo <= n7848_li206_li206;
    n3234_lo <= n7854_li208_li208;
    n3237_lo <= n7857_li209_li209;
    n3240_lo <= n7860_li210_li210;
    n3243_lo <= n7863_li211_li211;
    n3246_lo <= n7866_li212_li212;
    n3249_lo <= n7869_li213_li213;
    n3252_lo <= n7872_li214_li214;
    n3255_lo <= n7875_li215_li215;
    n3258_lo <= n7878_li216_li216;
    n3261_lo <= n7881_li217_li217;
    n3264_lo <= n7884_li218_li218;
    n3267_lo <= n7887_li219_li219;
    n3270_lo <= n7890_li220_li220;
    n3273_lo <= n7893_li221_li221;
    n3276_lo <= n7896_li222_li222;
    n3279_lo <= n7899_li223_li223;
    n3282_lo <= n7902_li224_li224;
    n3285_lo <= n7905_li225_li225;
    n3288_lo <= n7908_li226_li226;
    n3294_lo <= n7914_li228_li228;
    n3297_lo <= n7917_li229_li229;
    n3300_lo <= n7920_li230_li230;
    n3306_lo <= n7926_li232_li232;
    n3309_lo <= n7929_li233_li233;
    n3312_lo <= n7932_li234_li234;
    n3318_lo <= n7938_li236_li236;
    n3321_lo <= n7941_li237_li237;
    n3324_lo <= n7944_li238_li238;
    n3330_lo <= n7950_li240_li240;
    n3333_lo <= n7953_li241_li241;
    n3336_lo <= n7956_li242_li242;
    n3339_lo <= n7959_li243_li243;
    n3342_lo <= n7962_li244_li244;
    n3345_lo <= n7965_li245_li245;
    n3348_lo <= n7968_li246_li246;
    n3351_lo <= n7971_li247_li247;
    n3354_lo <= n7974_li248_li248;
    n3357_lo <= n7977_li249_li249;
    n3360_lo <= n7980_li250_li250;
    n3363_lo <= n7983_li251_li251;
    n3366_lo <= n7986_li252_li252;
    n3369_lo <= n7989_li253_li253;
    n3372_lo <= n7992_li254_li254;
    n3375_lo <= n7995_li255_li255;
    n3378_lo <= n7998_li256_li256;
    n3381_lo <= n8001_li257_li257;
    n3384_lo <= n8004_li258_li258;
    n3387_lo <= n8007_li259_li259;
    n3390_lo <= n8010_li260_li260;
    n3393_lo <= n8013_li261_li261;
    n3396_lo <= n8016_li262_li262;
    n3399_lo <= n8019_li263_li263;
    n3402_lo <= n8022_li264_li264;
    n3405_lo <= n8025_li265_li265;
    n3408_lo <= n8028_li266_li266;
    n3411_lo <= n8031_li267_li267;
    n3414_lo <= n8034_li268_li268;
    n3417_lo <= n8037_li269_li269;
    n3420_lo <= n8040_li270_li270;
    n3423_lo <= n8043_li271_li271;
    n3426_lo <= n8046_li272_li272;
    n3429_lo <= n8049_li273_li273;
    n3432_lo <= n8052_li274_li274;
    n3435_lo <= n8055_li275_li275;
    n3438_lo <= n8058_li276_li276;
    n3441_lo <= n8061_li277_li277;
    n3444_lo <= n8064_li278_li278;
    n3447_lo <= n8067_li279_li279;
    n3450_lo <= n8070_li280_li280;
    n3453_lo <= n8073_li281_li281;
    n3456_lo <= n8076_li282_li282;
    n3459_lo <= n8079_li283_li283;
    n3462_lo <= n8082_li284_li284;
    n3465_lo <= n8085_li285_li285;
    n3468_lo <= n8088_li286_li286;
    n3471_lo <= n8091_li287_li287;
    n3474_lo <= n8094_li288_li288;
    n3477_lo <= n8097_li289_li289;
    n3480_lo <= n8100_li290_li290;
    n3483_lo <= n8103_li291_li291;
    n3486_lo <= n8106_li292_li292;
    n3489_lo <= n8109_li293_li293;
    n3492_lo <= n8112_li294_li294;
    n3495_lo <= n8115_li295_li295;
    n3498_lo <= n8118_li296_li296;
    n3501_lo <= n8121_li297_li297;
    n3504_lo <= n8124_li298_li298;
    n3507_lo <= n8127_li299_li299;
    n3510_lo <= n8130_li300_li300;
    n3513_lo <= n8133_li301_li301;
    n3516_lo <= n8136_li302_li302;
    n3519_lo <= n8139_li303_li303;
    n3522_lo <= n8142_li304_li304;
    n3525_lo <= n8145_li305_li305;
    n3528_lo <= n8148_li306_li306;
    n3531_lo <= n8151_li307_li307;
    n3534_lo <= n8154_li308_li308;
    n3537_lo <= n8157_li309_li309;
    n3540_lo <= n8160_li310_li310;
    n3543_lo <= n8163_li311_li311;
    n3546_lo <= n8166_li312_li312;
    n3549_lo <= n8169_li313_li313;
    n3552_lo <= n8172_li314_li314;
    n3555_lo <= n8175_li315_li315;
    n3558_lo <= n8178_li316_li316;
    n3561_lo <= n8181_li317_li317;
    n3564_lo <= n8184_li318_li318;
    n3567_lo <= n8187_li319_li319;
    n3570_lo <= n8190_li320_li320;
    n3573_lo <= n8193_li321_li321;
    n3576_lo <= n8196_li322_li322;
    n3579_lo <= n8199_li323_li323;
    n3582_lo <= n8202_li324_li324;
    n3585_lo <= n8205_li325_li325;
    n3588_lo <= n8208_li326_li326;
    n3591_lo <= n8211_li327_li327;
    n3594_lo <= n8214_li328_li328;
    n3597_lo <= n8217_li329_li329;
    n3600_lo <= n8220_li330_li330;
    n3603_lo <= n8223_li331_li331;
    n3606_lo <= n8226_li332_li332;
    n3609_lo <= n8229_li333_li333;
    n3612_lo <= n8232_li334_li334;
    n3615_lo <= n8235_li335_li335;
    n3618_lo <= n8238_li336_li336;
    n3621_lo <= n8241_li337_li337;
    n3624_lo <= n8244_li338_li338;
    n3627_lo <= n8247_li339_li339;
    n3630_lo <= n8250_li340_li340;
    n3633_lo <= n8253_li341_li341;
    n3636_lo <= n8256_li342_li342;
    n3639_lo <= n8259_li343_li343;
    n3642_lo <= n8262_li344_li344;
    n3645_lo <= n8265_li345_li345;
    n3648_lo <= n8268_li346_li346;
    n3651_lo <= n8271_li347_li347;
    n3654_lo <= n8274_li348_li348;
    n3666_lo <= n8286_li352_li352;
    n3750_lo <= n8370_li380_li380;
    n3762_lo <= n8382_li384_li384;
    n3774_lo <= n8394_li388_li388;
    n3786_lo <= n8406_li392_li392;
    n3789_lo <= n8409_li393_li393;
    n3792_lo <= n8412_li394_li394;
    n3795_lo <= n8415_li395_li395;
    n3798_lo <= n8418_li396_li396;
    n3810_lo <= n8430_li400_li400;
    n3822_lo <= n8442_li404_li404;
    n3834_lo <= n8454_li408_li408;
    n3846_lo <= n8466_li412_li412;
    n3930_lo <= n8550_li440_li440;
    n3933_lo <= n8553_li441_li441;
    n3936_lo <= n8556_li442_li442;
    n3942_lo <= n8562_li444_li444;
    n3945_lo <= n8565_li445_li445;
    n3948_lo <= n8568_li446_li446;
    n3954_lo <= n8574_li448_li448;
    n3957_lo <= n8577_li449_li449;
    n3963_lo <= n8583_li451_li451;
    n3966_lo <= n8586_li452_li452;
    n3969_lo <= n8589_li453_li453;
    n3975_lo <= n8595_li455_li455;
    n3978_lo <= n8598_li456_li456;
    n3990_lo <= n8610_li460_li460;
    n4050_lo <= n8670_li480_li480;
    n4062_lo <= n8682_li484_li484;
    n4098_lo <= n8718_li496_li496;
    n4107_lo <= n8727_li499_li499;
    n4110_lo <= n8730_li500_li500;
    n4122_lo <= n8742_li504_li504;
    n4131_lo <= n8751_li507_li507;
    n4155_lo <= n8775_li515_li515;
    n4158_lo <= n8778_li516_li516;
    n4170_lo <= n8790_li520_li520;
    n4179_lo <= n8799_li523_li523;
    n4182_lo <= n8802_li524_li524;
    n4185_lo <= n8805_li525_li525;
    n4188_lo <= n8808_li526_li526;
    n4194_lo <= n8814_li528_li528;
    n4197_lo <= n8817_li529_li529;
    n4200_lo <= n8820_li530_li530;
    n4206_lo <= n8826_li532_li532;
    n4209_lo <= n8829_li533_li533;
    n4212_lo <= n8832_li534_li534;
    n4215_lo <= n8835_li535_li535;
    n4230_lo <= n8850_li540_li540;
    n4233_lo <= n8853_li541_li541;
    n4236_lo <= n8856_li542_li542;
    n4239_lo <= n8859_li543_li543;
    n4242_lo <= n8862_li544_li544;
    n4254_lo <= n8874_li548_li548;
    n4290_lo <= n8910_li560_li560;
    n4293_lo <= n8913_li561_li561;
    n4302_lo <= n8922_li564_li564;
    n4314_lo <= n8934_li568_li568;
    n4350_lo <= n8970_li580_li580;
    n4362_lo <= n8982_li584_li584;
    n4374_lo <= n8994_li588_li588;
    n4386_lo <= n9006_li592_li592;
    n4398_lo <= n9018_li596_li596;
    n4410_lo <= n9030_li600_li600;
    n4413_lo <= n9033_li601_li601;
    n4416_lo <= n9036_li602_li602;
    n4419_lo <= n9039_li603_li603;
    n4422_lo <= n9042_li604_li604;
    n4425_lo <= n9045_li605_li605;
    n4428_lo <= n9048_li606_li606;
    n4431_lo <= n9051_li607_li607;
    n4434_lo <= n9054_li608_li608;
    n4437_lo <= n9057_li609_li609;
    n4440_lo <= n9060_li610_li610;
    n4443_lo <= n9063_li611_li611;
    n4446_lo <= n9066_li612_li612;
    n4449_lo <= n9069_li613_li613;
    n4452_lo <= n9072_li614_li614;
    n4455_lo <= n9075_li615_li615;
    n4458_lo <= n9078_li616_li616;
    n4461_lo <= n9081_li617_li617;
    n4464_lo <= n9084_li618_li618;
    n4467_lo <= n9087_li619_li619;
    n4470_lo <= n9090_li620_li620;
    n4473_lo <= n9093_li621_li621;
    n4476_lo <= n9096_li622_li622;
    n4479_lo <= n9099_li623_li623;
    n4482_lo <= n9102_li624_li624;
    n4485_lo <= n9105_li625_li625;
    n4488_lo <= n9108_li626_li626;
    n4494_lo <= n9114_li628_li628;
    n4497_lo <= n9117_li629_li629;
    n4500_lo <= n9120_li630_li630;
    n4503_lo <= n9123_li631_li631;
    n4506_lo <= n9126_li632_li632;
    n4509_lo <= n9129_li633_li633;
    n4512_lo <= n9132_li634_li634;
    n4515_lo <= n9135_li635_li635;
    n4518_lo <= n9138_li636_li636;
    n4521_lo <= n9141_li637_li637;
    n4524_lo <= n9144_li638_li638;
    n4527_lo <= n9147_li639_li639;
    n4530_lo <= n9150_li640_li640;
    n4533_lo <= n9153_li641_li641;
    n4536_lo <= n9156_li642_li642;
    n4539_lo <= n9159_li643_li643;
    n4542_lo <= n9162_li644_li644;
    n4545_lo <= n9165_li645_li645;
    n4554_lo <= n9174_li648_li648;
    n4557_lo <= n9177_li649_li649;
    n4560_lo <= n9180_li650_li650;
    n4563_lo <= n9183_li651_li651;
    n4566_lo <= n9186_li652_li652;
    n4569_lo <= n9189_li653_li653;
    n4572_lo <= n9192_li654_li654;
    n4575_lo <= n9195_li655_li655;
    n4578_lo <= n9198_li656_li656;
    n4581_lo <= n9201_li657_li657;
    n4584_lo <= n9204_li658_li658;
    n4587_lo <= n9207_li659_li659;
    n4590_lo <= n9210_li660_li660;
    n4593_lo <= n9213_li661_li661;
    n4596_lo <= n9216_li662_li662;
    n4602_lo <= n9222_li664_li664;
    n4605_lo <= n9225_li665_li665;
    n4608_lo <= n9228_li666_li666;
    n4614_lo <= n9234_li668_li668;
    n4617_lo <= n9237_li669_li669;
    n4620_lo <= n9240_li670_li670;
    n4626_lo <= n9246_li672_li672;
    n4629_lo <= n9249_li673_li673;
    n4632_lo <= n9252_li674_li674;
    n4638_lo <= n9258_li676_li676;
    n4641_lo <= n9261_li677_li677;
    n4644_lo <= n9264_li678_li678;
    n4647_lo <= n9267_li679_li679;
    n4650_lo <= n9270_li680_li680;
    n4653_lo <= n9273_li681_li681;
    n4656_lo <= n9276_li682_li682;
    n4659_lo <= n9279_li683_li683;
    n4662_lo <= n9282_li684_li684;
    n4665_lo <= n9285_li685_li685;
    n4668_lo <= n9288_li686_li686;
    n4671_lo <= n9291_li687_li687;
    n4674_lo <= n9294_li688_li688;
    n4677_lo <= n9297_li689_li689;
    n4680_lo <= n9300_li690_li690;
    n4683_lo <= n9303_li691_li691;
    n4686_lo <= n9306_li692_li692;
    n4689_lo <= n9309_li693_li693;
    n4692_lo <= n9312_li694_li694;
    n4695_lo <= n9315_li695_li695;
    n4698_lo <= n9318_li696_li696;
    n4701_lo <= n9321_li697_li697;
    n4704_lo <= n9324_li698_li698;
    n4707_lo <= n9327_li699_li699;
    n4710_lo <= n9330_li700_li700;
    n4713_lo <= n9333_li701_li701;
    n4716_lo <= n9336_li702_li702;
    n4719_lo <= n9339_li703_li703;
    n4722_lo <= n9342_li704_li704;
    n4725_lo <= n9345_li705_li705;
    n4728_lo <= n9348_li706_li706;
    n4731_lo <= n9351_li707_li707;
    n4734_lo <= n9354_li708_li708;
    n4737_lo <= n9357_li709_li709;
    n4740_lo <= n9360_li710_li710;
    n4743_lo <= n9363_li711_li711;
    n4970_o2 <= n4970_i2;
    n4972_o2 <= n4972_i2;
    n4989_o2 <= n4989_i2;
    n5024_o2 <= n5024_i2;
    n5025_o2 <= n5025_i2;
    n5029_o2 <= n5029_i2;
    n5042_o2 <= n5042_i2;
    n5048_o2 <= n5048_i2;
    n5093_o2 <= n5093_i2;
    n5096_o2 <= n5096_i2;
    n5193_o2 <= n5193_i2;
    n5199_o2 <= n5199_i2;
    n5203_o2 <= n5203_i2;
    n5214_o2 <= n5214_i2;
    n5221_o2 <= n5221_i2;
    n5222_o2 <= n5222_i2;
    n5273_o2 <= n5273_i2;
    n5365_o2 <= n5365_i2;
    n5385_o2 <= n5385_i2;
    n5553_o2 <= n5553_i2;
    n5636_o2 <= n5636_i2;
    n5782_o2 <= n5782_i2;
    n5778_o2 <= n5778_i2;
    n5323_o2 <= n5323_i2;
    n5325_o2 <= n5325_i2;
    n5327_o2 <= n5327_i2;
    n5329_o2 <= n5329_i2;
    n5816_o2 <= n5816_i2;
    n5817_o2 <= n5817_i2;
    n5837_o2 <= n5837_i2;
    n5844_o2 <= n5844_i2;
    n5859_o2 <= n5859_i2;
    n5857_o2 <= n5857_i2;
    n5369_o2 <= n5369_i2;
    n5371_o2 <= n5371_i2;
    n5373_o2 <= n5373_i2;
    n5400_o2 <= n5400_i2;
    n5402_o2 <= n5402_i2;
    n5404_o2 <= n5404_i2;
    n5406_o2 <= n5406_i2;
    n5407_o2 <= n5407_i2;
    n5408_o2 <= n5408_i2;
    n2722_o2 <= n2722_i2;
    n1942_inv <= n5411_i2;
    n5412_o2 <= n5412_i2;
    n1948_inv <= n5413_i2;
    n5557_o2 <= n5557_i2;
    n5558_o2 <= n5558_i2;
    n5559_o2 <= n5559_i2;
    n5564_o2 <= n5564_i2;
    n5565_o2 <= n5565_i2;
    n1966_inv <= n5561_i2;
    n5568_o2 <= n5568_i2;
    n5598_o2 <= n5598_i2;
    n5600_o2 <= n5600_i2;
    n5601_o2 <= n5601_i2;
    n5602_o2 <= n5602_i2;
    n5603_o2 <= n5603_i2;
    n2853_o2 <= n2853_i2;
    n5637_o2 <= n5637_i2;
    n1993_inv <= n5627_i2;
    n1996_inv <= n5628_i2;
    n5635_o2 <= n5635_i2;
    n5640_o2 <= n5640_i2;
    n5641_o2 <= n5641_i2;
    n5642_o2 <= n5642_i2;
    n5650_o2 <= n5650_i2;
    n5652_o2 <= n5652_i2;
    n5653_o2 <= n5653_i2;
    n5654_o2 <= n5654_i2;
    n5655_o2 <= n5655_i2;
    n5657_o2 <= n5657_i2;
    n2029_inv <= n5659_i2;
    n5661_o2 <= n5661_i2;
    n5656_o2 <= n5656_i2;
    n5663_o2 <= n5663_i2;
    n2041_inv <= n5664_i2;
    n5795_o2 <= n5795_i2;
    n5796_o2 <= n5796_i2;
    n5797_o2 <= n5797_i2;
    n5739_o2 <= n5739_i2;
    n5773_o2 <= n5773_i2;
    n2059_inv <= n5798_i2;
    n5799_o2 <= n5799_i2;
    n5802_o2 <= n5802_i2;
    n2068_inv <= n5803_i2;
    n5831_o2 <= n5831_i2;
    n5833_o2 <= n5833_i2;
    n5820_o2 <= n5820_i2;
    n5823_o2 <= n5823_i2;
    n5824_o2 <= n5824_i2;
    n5869_o2 <= n5869_i2;
    n5848_o2 <= n5848_i2;
    n5849_o2 <= n5849_i2;
    n5856_o2 <= n5856_i2;
    n5896_o2 <= n5896_i2;
    n2754_o2 <= n2754_i2;
    n2908_o2 <= n2908_i2;
    n5892_o2 <= n5892_i2;
    n5915_o2 <= n5915_i2;
    n5919_o2 <= n5919_i2;
    n5918_o2 <= n5918_i2;
    n5920_o2 <= n5920_i2;
    n5917_o2 <= n5917_i2;
    lo586_buf_o2 <= lo586_buf_i2;
    n2818_o2 <= n2818_i2;
    n2863_o2 <= n2863_i2;
    n2134_inv <= n2721_i2;
    n2725_o2 <= n2725_i2;
    n3016_o2 <= n3016_i2;
    n3013_o2 <= n3013_i2;
    n2655_o2 <= n2655_i2;
    n2149_inv <= n2741_i2;
    lo562_buf_o2 <= lo562_buf_i2;
    n2155_inv <= n2656_i2;
    n2531_o2 <= n2531_i2;
    n2700_o2 <= n2700_i2;
    n5908_o2 <= n5908_i2;
    n5910_o2 <= n5910_i2;
    n5912_o2 <= n5912_i2;
    n5914_o2 <= n5914_i2;
    n2753_o2 <= n2753_i2;
    n2878_o2 <= n2878_i2;
    n2182_inv <= n2836_i2;
    n5934_o2 <= n5934_i2;
    n5936_o2 <= n5936_i2;
    n5938_o2 <= n5938_i2;
    n2728_o2 <= n2728_i2;
    lo358_buf_o2 <= lo358_buf_i2;
    lo418_buf_o2 <= lo418_buf_i2;
    lo474_buf_o2 <= lo474_buf_i2;
    lo554_buf_o2 <= lo554_buf_i2;
    lo558_buf_o2 <= lo558_buf_i2;
    lo574_buf_o2 <= lo574_buf_i2;
    n2215_inv <= n2659_i2;
    n2218_inv <= n2665_i2;
    n2221_inv <= n2686_i2;
    lo450_buf_o2 <= lo450_buf_i2;
    n2910_o2 <= n2910_i2;
    n2683_o2 <= n2683_i2;
    n2828_o2 <= n2828_i2;
    n2582_o2 <= n2582_i2;
    n2600_o2 <= n2600_i2;
    n2542_o2 <= n2542_i2;
    n2703_o2 <= n2703_i2;
    lo510_buf_o2 <= lo510_buf_i2;
    lo514_buf_o2 <= lo514_buf_i2;
    lo538_buf_o2 <= lo538_buf_i2;
    lo578_buf_o2 <= lo578_buf_i2;
    n2260_inv <= n2692_i2;
    n2666_o2 <= n2666_i2;
    n2667_o2 <= n2667_i2;
    n2660_o2 <= n2660_i2;
    n2272_inv <= n2744_i2;
    lo454_buf_o2 <= lo454_buf_i2;
    n3593_o2 <= n3593_i2;
    n3048_o2 <= n3048_i2;
    lo410_buf_o2 <= lo410_buf_i2;
    lo502_buf_o2 <= lo502_buf_i2;
    lo506_buf_o2 <= lo506_buf_i2;
    lo550_buf_o2 <= lo550_buf_i2;
    lo570_buf_o2 <= lo570_buf_i2;
    lo582_buf_o2 <= lo582_buf_i2;
    n2302_inv <= n2646_i2;
    n2305_inv <= n2673_i2;
    n3499_o2 <= n3499_i2;
    n2311_inv <= n2750_i2;
    n2870_o2 <= n2870_i2;
    n2317_inv <= n2693_i2;
    n2689_o2 <= n2689_i2;
    n2323_inv <= n2668_i2;
    n2662_o2 <= n2662_i2;
    lo350_buf_o2 <= lo350_buf_i2;
    lo498_buf_o2 <= lo498_buf_i2;
    lo518_buf_o2 <= lo518_buf_i2;
    lo522_buf_o2 <= lo522_buf_i2;
    lo598_buf_o2 <= lo598_buf_i2;
    n2344_inv <= n2708_i2;
    n2347_inv <= n2674_i2;
    n2350_inv <= n2647_i2;
    n2353_inv <= n2751_i2;
    n2356_inv <= n2747_i2;
    n2359_inv <= n2669_i2;
    n2872_o2 <= n2872_i2;
    n3313_o2 <= n3313_i2;
    n3273_o2 <= n3273_i2;
    n2848_o2 <= n2848_i2;
    n2893_o2 <= n2893_i2;
    n3267_o2 <= n3267_i2;
    n2925_o2 <= n2925_i2;
    n2839_o2 <= n2839_i2;
    n2831_o2 <= n2831_i2;
    n2558_o2 <= n2558_i2;
    n2562_o2 <= n2562_i2;
    n2825_o2 <= n2825_i2;
    n3263_o2 <= n3263_i2;
    n3517_o2 <= n3517_i2;
    n2873_o2 <= n2873_i2;
    n2926_o2 <= n2926_i2;
    n3261_o2 <= n3261_i2;
    n3268_o2 <= n3268_i2;
    n3274_o2 <= n3274_i2;
    n3314_o2 <= n3314_i2;
    n3571_o2 <= n3571_i2;
    n2950_o2 <= n2950_i2;
    n2951_o2 <= n2951_i2;
    n3022_o2 <= n3022_i2;
    n3023_o2 <= n3023_i2;
    n3057_o2 <= n3057_i2;
    n3058_o2 <= n3058_i2;
    n2931_o2 <= n2931_i2;
    n2911_o2 <= n2911_i2;
    n2959_o2 <= n2959_i2;
    n2960_o2 <= n2960_i2;
    n2922_o2 <= n2922_i2;
    n2888_o2 <= n2888_i2;
    n2889_o2 <= n2889_i2;
    n3051_o2 <= n3051_i2;
    n3052_o2 <= n3052_i2;
    n3063_o2 <= n3063_i2;
    n2845_o2 <= n2845_i2;
    n2476_inv <= n2737_i2;
    n3281_o2 <= n3281_i2;
    n3294_o2 <= n3294_i2;
    n2885_o2 <= n2885_i2;
    n2786_o2 <= n2786_i2;
    n2783_o2 <= n2783_i2;
    n2801_o2 <= n2801_i2;
    n2572_o2 <= n2572_i2;
    n2628_o2 <= n2628_i2;
    n2609_o2 <= n2609_i2;
    n2618_o2 <= n2618_i2;
    n2637_o2 <= n2637_i2;
    n2525_o2 <= n2525_i2;
    n2551_o2 <= n2551_i2;
    n3759_o2 <= n3759_i2;
    n2994_o2 <= n2994_i2;
    n3040_o2 <= n3040_i2;
    n2943_o2 <= n2943_i2;
    n2991_o2 <= n2991_i2;
    n3034_o2 <= n3034_i2;
    n2881_o2 <= n2881_i2;
    n3021_o2 <= n3021_i2;
    n3062_o2 <= n3062_i2;
    n2763_o2 <= n2763_i2;
    n2764_o2 <= n2764_i2;
    n2775_o2 <= n2775_i2;
    n2776_o2 <= n2776_i2;
    n2968_o2 <= n2968_i2;
    n2969_o2 <= n2969_i2;
    n2798_o2 <= n2798_i2;
    n3661_o2 <= n3661_i2;
    n2694_o2 <= n2694_i2;
    n2572_inv <= n2809_i2;
    n2817_o2 <= n2817_i2;
    n2514_o2 <= n2514_i2;
    n2501_o2 <= n2501_i2;
    n2584_inv <= n2528_i2;
    n2505_o2 <= n2505_i2;
    n2492_o2 <= n2492_i2;
    lo546_buf_o2 <= lo546_buf_i2;
    lo590_buf_o2 <= lo590_buf_i2;
    lo594_buf_o2 <= lo594_buf_i2;
    n2602_inv <= n2679_i2;
    n2605_inv <= n2733_i2;
    n2709_o2 <= n2709_i2;
    n2611_inv <= n2676_i2;
    n2614_inv <= n2649_i2;
    n2617_inv <= n2815_i2;
    n2620_inv <= n2704_i2;
    n3590_o2 <= n3590_i2;
    n3591_o2 <= n3591_i2;
    n2629_inv <= n2752_i2;
    n3638_o2 <= n3638_i2;
    n3639_o2 <= n3639_i2;
    n2638_inv <= n2695_i2;
    n2641_inv <= n3047_i2;
    lo458_buf_o2 <= lo458_buf_i2;
    lo482_buf_o2 <= lo482_buf_i2;
    lo566_buf_o2 <= lo566_buf_i2;
    n2718_o2 <= n2718_i2;
    n3707_o2 <= n3707_i2;
    n3671_o2 <= n3671_i2;
    n3680_o2 <= n3680_i2;
    n3749_o2 <= n3749_i2;
    n3716_o2 <= n3716_i2;
    n3692_o2 <= n3692_i2;
    n2591_o2 <= n2591_i2;
    n3478_o2 <= n3478_i2;
    n3610_o2 <= n3610_i2;
    n3611_o2 <= n3611_i2;
    n2686_inv <= n2652_i2;
    n2689_inv <= n2714_i2;
    n2738_o2 <= n2738_i2;
    n3616_o2 <= n3616_i2;
    n3617_o2 <= n3617_i2;
    n3031_o2 <= n3031_i2;
    n2704_inv <= n2515_i2;
    n3562_o2 <= n3562_i2;
    n2502_o2 <= n2502_i2;
    n3560_o2 <= n3560_i2;
    n3554_o2 <= n3554_i2;
    n3555_o2 <= n3555_i2;
    n3536_o2 <= n3536_i2;
    n3537_o2 <= n3537_i2;
    n3508_o2 <= n3508_i2;
    n3650_o2 <= n3650_i2;
    n3740_o2 <= n3740_i2;
    n3484_o2 <= n3484_i2;
    n2740_inv <= n2680_i2;
    n2734_o2 <= n2734_i2;
    n2735_o2 <= n2735_i2;
    n2711_o2 <= n2711_i2;
    lo585_buf_o2 <= lo585_buf_i2;
    n2719_o2 <= n2719_i2;
    n2720_o2 <= n2720_i2;
    n2723_o2 <= n2723_i2;
    n2724_o2 <= n2724_i2;
    n3624_o2 <= n3624_i2;
    n3625_o2 <= n3625_i2;
    n3015_o2 <= n3015_i2;
    n3491_o2 <= n3491_i2;
    n2779_inv <= n2696_i2;
    n2811_o2 <= n2811_i2;
    n3010_o2 <= n3010_i2;
    n3012_o2 <= n3012_i2;
    lo382_buf_o2 <= lo382_buf_i2;
    lo386_buf_o2 <= lo386_buf_i2;
    lo390_buf_o2 <= lo390_buf_i2;
    lo398_buf_o2 <= lo398_buf_i2;
    lo402_buf_o2 <= lo402_buf_i2;
    lo406_buf_o2 <= lo406_buf_i2;
    n3492_o2 <= n3492_i2;
    lo366_buf_o2 <= lo366_buf_i2;
    lo374_buf_o2 <= lo374_buf_i2;
    lo426_buf_o2 <= lo426_buf_i2;
    lo494_buf_o2 <= lo494_buf_i2;
    n2653_o2 <= n2653_i2;
    n2654_o2 <= n2654_i2;
    n2715_o2 <= n2715_i2;
    n2740_o2 <= n2740_i2;
    n2682_o2 <= n2682_i2;
    n2736_o2 <= n2736_i2;
    lo508_buf_o2 <= lo508_buf_i2;
    lo512_buf_o2 <= lo512_buf_i2;
    lo536_buf_o2 <= lo536_buf_i2;
    lo576_buf_o2 <= lo576_buf_i2;
    lo357_buf_o2 <= lo357_buf_i2;
    lo361_buf_o2 <= lo361_buf_i2;
    lo417_buf_o2 <= lo417_buf_i2;
    lo421_buf_o2 <= lo421_buf_i2;
    lo473_buf_o2 <= lo473_buf_i2;
    lo477_buf_o2 <= lo477_buf_i2;
    lo553_buf_o2 <= lo553_buf_i2;
    lo557_buf_o2 <= lo557_buf_i2;
    lo573_buf_o2 <= lo573_buf_i2;
    lo434_buf_o2 <= lo434_buf_i2;
    lo438_buf_o2 <= lo438_buf_i2;
    lo466_buf_o2 <= lo466_buf_i2;
    lo470_buf_o2 <= lo470_buf_i2;
    lo490_buf_o2 <= lo490_buf_i2;
    n2657_o2 <= n2657_i2;
    n2658_o2 <= n2658_i2;
    n2663_o2 <= n2663_i2;
    n2664_o2 <= n2664_i2;
    n2684_o2 <= n2684_i2;
    n2685_o2 <= n2685_i2;
  end
  initial begin
    n2610_lo <= 1'b0;
    n2613_lo <= 1'b0;
    n2616_lo <= 1'b0;
    n2619_lo <= 1'b0;
    n2622_lo <= 1'b0;
    n2625_lo <= 1'b0;
    n2628_lo <= 1'b0;
    n2634_lo <= 1'b0;
    n2637_lo <= 1'b0;
    n2640_lo <= 1'b0;
    n2643_lo <= 1'b0;
    n2646_lo <= 1'b0;
    n2649_lo <= 1'b0;
    n2652_lo <= 1'b0;
    n2655_lo <= 1'b0;
    n2658_lo <= 1'b0;
    n2661_lo <= 1'b0;
    n2664_lo <= 1'b0;
    n2667_lo <= 1'b0;
    n2670_lo <= 1'b0;
    n2673_lo <= 1'b0;
    n2676_lo <= 1'b0;
    n2679_lo <= 1'b0;
    n2682_lo <= 1'b0;
    n2685_lo <= 1'b0;
    n2688_lo <= 1'b0;
    n2691_lo <= 1'b0;
    n2694_lo <= 1'b0;
    n2697_lo <= 1'b0;
    n2700_lo <= 1'b0;
    n2703_lo <= 1'b0;
    n2706_lo <= 1'b0;
    n2709_lo <= 1'b0;
    n2712_lo <= 1'b0;
    n2715_lo <= 1'b0;
    n2718_lo <= 1'b0;
    n2721_lo <= 1'b0;
    n2724_lo <= 1'b0;
    n2727_lo <= 1'b0;
    n2730_lo <= 1'b0;
    n2733_lo <= 1'b0;
    n2736_lo <= 1'b0;
    n2739_lo <= 1'b0;
    n2742_lo <= 1'b0;
    n2745_lo <= 1'b0;
    n2748_lo <= 1'b0;
    n2751_lo <= 1'b0;
    n2754_lo <= 1'b0;
    n2757_lo <= 1'b0;
    n2760_lo <= 1'b0;
    n2763_lo <= 1'b0;
    n2766_lo <= 1'b0;
    n2769_lo <= 1'b0;
    n2772_lo <= 1'b0;
    n2775_lo <= 1'b0;
    n2778_lo <= 1'b0;
    n2781_lo <= 1'b0;
    n2784_lo <= 1'b0;
    n2787_lo <= 1'b0;
    n2790_lo <= 1'b0;
    n2793_lo <= 1'b0;
    n2796_lo <= 1'b0;
    n2799_lo <= 1'b0;
    n2802_lo <= 1'b0;
    n2805_lo <= 1'b0;
    n2808_lo <= 1'b0;
    n2811_lo <= 1'b0;
    n2814_lo <= 1'b0;
    n2817_lo <= 1'b0;
    n2820_lo <= 1'b0;
    n2823_lo <= 1'b0;
    n2826_lo <= 1'b0;
    n2829_lo <= 1'b0;
    n2832_lo <= 1'b0;
    n2838_lo <= 1'b0;
    n2841_lo <= 1'b0;
    n2844_lo <= 1'b0;
    n2847_lo <= 1'b0;
    n2850_lo <= 1'b0;
    n2853_lo <= 1'b0;
    n2856_lo <= 1'b0;
    n2862_lo <= 1'b0;
    n2865_lo <= 1'b0;
    n2868_lo <= 1'b0;
    n2871_lo <= 1'b0;
    n2874_lo <= 1'b0;
    n2877_lo <= 1'b0;
    n2880_lo <= 1'b0;
    n2883_lo <= 1'b0;
    n2886_lo <= 1'b0;
    n2889_lo <= 1'b0;
    n2892_lo <= 1'b0;
    n2895_lo <= 1'b0;
    n2898_lo <= 1'b0;
    n2901_lo <= 1'b0;
    n2904_lo <= 1'b0;
    n2907_lo <= 1'b0;
    n2910_lo <= 1'b0;
    n2913_lo <= 1'b0;
    n2916_lo <= 1'b0;
    n2919_lo <= 1'b0;
    n2922_lo <= 1'b0;
    n2925_lo <= 1'b0;
    n2928_lo <= 1'b0;
    n2931_lo <= 1'b0;
    n2934_lo <= 1'b0;
    n2937_lo <= 1'b0;
    n2940_lo <= 1'b0;
    n2943_lo <= 1'b0;
    n2946_lo <= 1'b0;
    n2949_lo <= 1'b0;
    n2952_lo <= 1'b0;
    n2955_lo <= 1'b0;
    n2958_lo <= 1'b0;
    n2961_lo <= 1'b0;
    n2964_lo <= 1'b0;
    n2967_lo <= 1'b0;
    n2970_lo <= 1'b0;
    n2973_lo <= 1'b0;
    n2976_lo <= 1'b0;
    n2979_lo <= 1'b0;
    n2982_lo <= 1'b0;
    n2985_lo <= 1'b0;
    n2988_lo <= 1'b0;
    n2991_lo <= 1'b0;
    n2994_lo <= 1'b0;
    n2997_lo <= 1'b0;
    n3000_lo <= 1'b0;
    n3003_lo <= 1'b0;
    n3006_lo <= 1'b0;
    n3009_lo <= 1'b0;
    n3012_lo <= 1'b0;
    n3015_lo <= 1'b0;
    n3018_lo <= 1'b0;
    n3021_lo <= 1'b0;
    n3024_lo <= 1'b0;
    n3027_lo <= 1'b0;
    n3030_lo <= 1'b0;
    n3033_lo <= 1'b0;
    n3036_lo <= 1'b0;
    n3039_lo <= 1'b0;
    n3042_lo <= 1'b0;
    n3045_lo <= 1'b0;
    n3048_lo <= 1'b0;
    n3051_lo <= 1'b0;
    n3054_lo <= 1'b0;
    n3057_lo <= 1'b0;
    n3060_lo <= 1'b0;
    n3063_lo <= 1'b0;
    n3066_lo <= 1'b0;
    n3069_lo <= 1'b0;
    n3072_lo <= 1'b0;
    n3075_lo <= 1'b0;
    n3078_lo <= 1'b0;
    n3081_lo <= 1'b0;
    n3084_lo <= 1'b0;
    n3087_lo <= 1'b0;
    n3090_lo <= 1'b0;
    n3093_lo <= 1'b0;
    n3096_lo <= 1'b0;
    n3099_lo <= 1'b0;
    n3102_lo <= 1'b0;
    n3105_lo <= 1'b0;
    n3108_lo <= 1'b0;
    n3111_lo <= 1'b0;
    n3114_lo <= 1'b0;
    n3117_lo <= 1'b0;
    n3120_lo <= 1'b0;
    n3126_lo <= 1'b0;
    n3129_lo <= 1'b0;
    n3132_lo <= 1'b0;
    n3138_lo <= 1'b0;
    n3141_lo <= 1'b0;
    n3144_lo <= 1'b0;
    n3147_lo <= 1'b0;
    n3150_lo <= 1'b0;
    n3153_lo <= 1'b0;
    n3156_lo <= 1'b0;
    n3162_lo <= 1'b0;
    n3165_lo <= 1'b0;
    n3168_lo <= 1'b0;
    n3174_lo <= 1'b0;
    n3177_lo <= 1'b0;
    n3180_lo <= 1'b0;
    n3186_lo <= 1'b0;
    n3189_lo <= 1'b0;
    n3192_lo <= 1'b0;
    n3195_lo <= 1'b0;
    n3198_lo <= 1'b0;
    n3201_lo <= 1'b0;
    n3204_lo <= 1'b0;
    n3210_lo <= 1'b0;
    n3213_lo <= 1'b0;
    n3216_lo <= 1'b0;
    n3219_lo <= 1'b0;
    n3222_lo <= 1'b0;
    n3225_lo <= 1'b0;
    n3228_lo <= 1'b0;
    n3234_lo <= 1'b0;
    n3237_lo <= 1'b0;
    n3240_lo <= 1'b0;
    n3243_lo <= 1'b0;
    n3246_lo <= 1'b0;
    n3249_lo <= 1'b0;
    n3252_lo <= 1'b0;
    n3255_lo <= 1'b0;
    n3258_lo <= 1'b0;
    n3261_lo <= 1'b0;
    n3264_lo <= 1'b0;
    n3267_lo <= 1'b0;
    n3270_lo <= 1'b0;
    n3273_lo <= 1'b0;
    n3276_lo <= 1'b0;
    n3279_lo <= 1'b0;
    n3282_lo <= 1'b0;
    n3285_lo <= 1'b0;
    n3288_lo <= 1'b0;
    n3294_lo <= 1'b0;
    n3297_lo <= 1'b0;
    n3300_lo <= 1'b0;
    n3306_lo <= 1'b0;
    n3309_lo <= 1'b0;
    n3312_lo <= 1'b0;
    n3318_lo <= 1'b0;
    n3321_lo <= 1'b0;
    n3324_lo <= 1'b0;
    n3330_lo <= 1'b0;
    n3333_lo <= 1'b0;
    n3336_lo <= 1'b0;
    n3339_lo <= 1'b0;
    n3342_lo <= 1'b0;
    n3345_lo <= 1'b0;
    n3348_lo <= 1'b0;
    n3351_lo <= 1'b0;
    n3354_lo <= 1'b0;
    n3357_lo <= 1'b0;
    n3360_lo <= 1'b0;
    n3363_lo <= 1'b0;
    n3366_lo <= 1'b0;
    n3369_lo <= 1'b0;
    n3372_lo <= 1'b0;
    n3375_lo <= 1'b0;
    n3378_lo <= 1'b0;
    n3381_lo <= 1'b0;
    n3384_lo <= 1'b0;
    n3387_lo <= 1'b0;
    n3390_lo <= 1'b0;
    n3393_lo <= 1'b0;
    n3396_lo <= 1'b0;
    n3399_lo <= 1'b0;
    n3402_lo <= 1'b0;
    n3405_lo <= 1'b0;
    n3408_lo <= 1'b0;
    n3411_lo <= 1'b0;
    n3414_lo <= 1'b0;
    n3417_lo <= 1'b0;
    n3420_lo <= 1'b0;
    n3423_lo <= 1'b0;
    n3426_lo <= 1'b0;
    n3429_lo <= 1'b0;
    n3432_lo <= 1'b0;
    n3435_lo <= 1'b0;
    n3438_lo <= 1'b0;
    n3441_lo <= 1'b0;
    n3444_lo <= 1'b0;
    n3447_lo <= 1'b0;
    n3450_lo <= 1'b0;
    n3453_lo <= 1'b0;
    n3456_lo <= 1'b0;
    n3459_lo <= 1'b0;
    n3462_lo <= 1'b0;
    n3465_lo <= 1'b0;
    n3468_lo <= 1'b0;
    n3471_lo <= 1'b0;
    n3474_lo <= 1'b0;
    n3477_lo <= 1'b0;
    n3480_lo <= 1'b0;
    n3483_lo <= 1'b0;
    n3486_lo <= 1'b0;
    n3489_lo <= 1'b0;
    n3492_lo <= 1'b0;
    n3495_lo <= 1'b0;
    n3498_lo <= 1'b0;
    n3501_lo <= 1'b0;
    n3504_lo <= 1'b0;
    n3507_lo <= 1'b0;
    n3510_lo <= 1'b0;
    n3513_lo <= 1'b0;
    n3516_lo <= 1'b0;
    n3519_lo <= 1'b0;
    n3522_lo <= 1'b0;
    n3525_lo <= 1'b0;
    n3528_lo <= 1'b0;
    n3531_lo <= 1'b0;
    n3534_lo <= 1'b0;
    n3537_lo <= 1'b0;
    n3540_lo <= 1'b0;
    n3543_lo <= 1'b0;
    n3546_lo <= 1'b0;
    n3549_lo <= 1'b0;
    n3552_lo <= 1'b0;
    n3555_lo <= 1'b0;
    n3558_lo <= 1'b0;
    n3561_lo <= 1'b0;
    n3564_lo <= 1'b0;
    n3567_lo <= 1'b0;
    n3570_lo <= 1'b0;
    n3573_lo <= 1'b0;
    n3576_lo <= 1'b0;
    n3579_lo <= 1'b0;
    n3582_lo <= 1'b0;
    n3585_lo <= 1'b0;
    n3588_lo <= 1'b0;
    n3591_lo <= 1'b0;
    n3594_lo <= 1'b0;
    n3597_lo <= 1'b0;
    n3600_lo <= 1'b0;
    n3603_lo <= 1'b0;
    n3606_lo <= 1'b0;
    n3609_lo <= 1'b0;
    n3612_lo <= 1'b0;
    n3615_lo <= 1'b0;
    n3618_lo <= 1'b0;
    n3621_lo <= 1'b0;
    n3624_lo <= 1'b0;
    n3627_lo <= 1'b0;
    n3630_lo <= 1'b0;
    n3633_lo <= 1'b0;
    n3636_lo <= 1'b0;
    n3639_lo <= 1'b0;
    n3642_lo <= 1'b0;
    n3645_lo <= 1'b0;
    n3648_lo <= 1'b0;
    n3651_lo <= 1'b0;
    n3654_lo <= 1'b0;
    n3666_lo <= 1'b0;
    n3750_lo <= 1'b0;
    n3762_lo <= 1'b0;
    n3774_lo <= 1'b0;
    n3786_lo <= 1'b0;
    n3789_lo <= 1'b0;
    n3792_lo <= 1'b0;
    n3795_lo <= 1'b0;
    n3798_lo <= 1'b0;
    n3810_lo <= 1'b0;
    n3822_lo <= 1'b0;
    n3834_lo <= 1'b0;
    n3846_lo <= 1'b0;
    n3930_lo <= 1'b0;
    n3933_lo <= 1'b0;
    n3936_lo <= 1'b0;
    n3942_lo <= 1'b0;
    n3945_lo <= 1'b0;
    n3948_lo <= 1'b0;
    n3954_lo <= 1'b0;
    n3957_lo <= 1'b0;
    n3963_lo <= 1'b0;
    n3966_lo <= 1'b0;
    n3969_lo <= 1'b0;
    n3975_lo <= 1'b0;
    n3978_lo <= 1'b0;
    n3990_lo <= 1'b0;
    n4050_lo <= 1'b0;
    n4062_lo <= 1'b0;
    n4098_lo <= 1'b0;
    n4107_lo <= 1'b0;
    n4110_lo <= 1'b0;
    n4122_lo <= 1'b0;
    n4131_lo <= 1'b0;
    n4155_lo <= 1'b0;
    n4158_lo <= 1'b0;
    n4170_lo <= 1'b0;
    n4179_lo <= 1'b0;
    n4182_lo <= 1'b0;
    n4185_lo <= 1'b0;
    n4188_lo <= 1'b0;
    n4194_lo <= 1'b0;
    n4197_lo <= 1'b0;
    n4200_lo <= 1'b0;
    n4206_lo <= 1'b0;
    n4209_lo <= 1'b0;
    n4212_lo <= 1'b0;
    n4215_lo <= 1'b0;
    n4230_lo <= 1'b0;
    n4233_lo <= 1'b0;
    n4236_lo <= 1'b0;
    n4239_lo <= 1'b0;
    n4242_lo <= 1'b0;
    n4254_lo <= 1'b0;
    n4290_lo <= 1'b0;
    n4293_lo <= 1'b0;
    n4302_lo <= 1'b0;
    n4314_lo <= 1'b0;
    n4350_lo <= 1'b0;
    n4362_lo <= 1'b0;
    n4374_lo <= 1'b0;
    n4386_lo <= 1'b0;
    n4398_lo <= 1'b0;
    n4410_lo <= 1'b0;
    n4413_lo <= 1'b0;
    n4416_lo <= 1'b0;
    n4419_lo <= 1'b0;
    n4422_lo <= 1'b0;
    n4425_lo <= 1'b0;
    n4428_lo <= 1'b0;
    n4431_lo <= 1'b0;
    n4434_lo <= 1'b0;
    n4437_lo <= 1'b0;
    n4440_lo <= 1'b0;
    n4443_lo <= 1'b0;
    n4446_lo <= 1'b0;
    n4449_lo <= 1'b0;
    n4452_lo <= 1'b0;
    n4455_lo <= 1'b0;
    n4458_lo <= 1'b0;
    n4461_lo <= 1'b0;
    n4464_lo <= 1'b0;
    n4467_lo <= 1'b0;
    n4470_lo <= 1'b0;
    n4473_lo <= 1'b0;
    n4476_lo <= 1'b0;
    n4479_lo <= 1'b0;
    n4482_lo <= 1'b0;
    n4485_lo <= 1'b0;
    n4488_lo <= 1'b0;
    n4494_lo <= 1'b0;
    n4497_lo <= 1'b0;
    n4500_lo <= 1'b0;
    n4503_lo <= 1'b0;
    n4506_lo <= 1'b0;
    n4509_lo <= 1'b0;
    n4512_lo <= 1'b0;
    n4515_lo <= 1'b0;
    n4518_lo <= 1'b0;
    n4521_lo <= 1'b0;
    n4524_lo <= 1'b0;
    n4527_lo <= 1'b0;
    n4530_lo <= 1'b0;
    n4533_lo <= 1'b0;
    n4536_lo <= 1'b0;
    n4539_lo <= 1'b0;
    n4542_lo <= 1'b0;
    n4545_lo <= 1'b0;
    n4554_lo <= 1'b0;
    n4557_lo <= 1'b0;
    n4560_lo <= 1'b0;
    n4563_lo <= 1'b0;
    n4566_lo <= 1'b0;
    n4569_lo <= 1'b0;
    n4572_lo <= 1'b0;
    n4575_lo <= 1'b0;
    n4578_lo <= 1'b0;
    n4581_lo <= 1'b0;
    n4584_lo <= 1'b0;
    n4587_lo <= 1'b0;
    n4590_lo <= 1'b0;
    n4593_lo <= 1'b0;
    n4596_lo <= 1'b0;
    n4602_lo <= 1'b0;
    n4605_lo <= 1'b0;
    n4608_lo <= 1'b0;
    n4614_lo <= 1'b0;
    n4617_lo <= 1'b0;
    n4620_lo <= 1'b0;
    n4626_lo <= 1'b0;
    n4629_lo <= 1'b0;
    n4632_lo <= 1'b0;
    n4638_lo <= 1'b0;
    n4641_lo <= 1'b0;
    n4644_lo <= 1'b0;
    n4647_lo <= 1'b0;
    n4650_lo <= 1'b0;
    n4653_lo <= 1'b0;
    n4656_lo <= 1'b0;
    n4659_lo <= 1'b0;
    n4662_lo <= 1'b0;
    n4665_lo <= 1'b0;
    n4668_lo <= 1'b0;
    n4671_lo <= 1'b0;
    n4674_lo <= 1'b0;
    n4677_lo <= 1'b0;
    n4680_lo <= 1'b0;
    n4683_lo <= 1'b0;
    n4686_lo <= 1'b0;
    n4689_lo <= 1'b0;
    n4692_lo <= 1'b0;
    n4695_lo <= 1'b0;
    n4698_lo <= 1'b0;
    n4701_lo <= 1'b0;
    n4704_lo <= 1'b0;
    n4707_lo <= 1'b0;
    n4710_lo <= 1'b0;
    n4713_lo <= 1'b0;
    n4716_lo <= 1'b0;
    n4719_lo <= 1'b0;
    n4722_lo <= 1'b0;
    n4725_lo <= 1'b0;
    n4728_lo <= 1'b0;
    n4731_lo <= 1'b0;
    n4734_lo <= 1'b0;
    n4737_lo <= 1'b0;
    n4740_lo <= 1'b0;
    n4743_lo <= 1'b0;
    n4970_o2 <= 1'b0;
    n4972_o2 <= 1'b0;
    n4989_o2 <= 1'b0;
    n5024_o2 <= 1'b0;
    n5025_o2 <= 1'b0;
    n5029_o2 <= 1'b0;
    n5042_o2 <= 1'b0;
    n5048_o2 <= 1'b0;
    n5093_o2 <= 1'b0;
    n5096_o2 <= 1'b0;
    n5193_o2 <= 1'b0;
    n5199_o2 <= 1'b0;
    n5203_o2 <= 1'b0;
    n5214_o2 <= 1'b0;
    n5221_o2 <= 1'b0;
    n5222_o2 <= 1'b0;
    n5273_o2 <= 1'b0;
    n5365_o2 <= 1'b0;
    n5385_o2 <= 1'b0;
    n5553_o2 <= 1'b0;
    n5636_o2 <= 1'b0;
    n5782_o2 <= 1'b0;
    n5778_o2 <= 1'b0;
    n5323_o2 <= 1'b0;
    n5325_o2 <= 1'b0;
    n5327_o2 <= 1'b0;
    n5329_o2 <= 1'b0;
    n5816_o2 <= 1'b0;
    n5817_o2 <= 1'b0;
    n5837_o2 <= 1'b0;
    n5844_o2 <= 1'b0;
    n5859_o2 <= 1'b0;
    n5857_o2 <= 1'b0;
    n5369_o2 <= 1'b0;
    n5371_o2 <= 1'b0;
    n5373_o2 <= 1'b0;
    n5400_o2 <= 1'b0;
    n5402_o2 <= 1'b0;
    n5404_o2 <= 1'b0;
    n5406_o2 <= 1'b0;
    n5407_o2 <= 1'b0;
    n5408_o2 <= 1'b0;
    n2722_o2 <= 1'b0;
    n1942_inv <= 1'b0;
    n5412_o2 <= 1'b0;
    n1948_inv <= 1'b0;
    n5557_o2 <= 1'b0;
    n5558_o2 <= 1'b0;
    n5559_o2 <= 1'b0;
    n5564_o2 <= 1'b0;
    n5565_o2 <= 1'b0;
    n1966_inv <= 1'b0;
    n5568_o2 <= 1'b0;
    n5598_o2 <= 1'b0;
    n5600_o2 <= 1'b0;
    n5601_o2 <= 1'b0;
    n5602_o2 <= 1'b0;
    n5603_o2 <= 1'b0;
    n2853_o2 <= 1'b0;
    n5637_o2 <= 1'b0;
    n1993_inv <= 1'b0;
    n1996_inv <= 1'b0;
    n5635_o2 <= 1'b0;
    n5640_o2 <= 1'b0;
    n5641_o2 <= 1'b0;
    n5642_o2 <= 1'b0;
    n5650_o2 <= 1'b0;
    n5652_o2 <= 1'b0;
    n5653_o2 <= 1'b0;
    n5654_o2 <= 1'b0;
    n5655_o2 <= 1'b0;
    n5657_o2 <= 1'b0;
    n2029_inv <= 1'b0;
    n5661_o2 <= 1'b0;
    n5656_o2 <= 1'b0;
    n5663_o2 <= 1'b0;
    n2041_inv <= 1'b0;
    n5795_o2 <= 1'b0;
    n5796_o2 <= 1'b0;
    n5797_o2 <= 1'b0;
    n5739_o2 <= 1'b0;
    n5773_o2 <= 1'b0;
    n2059_inv <= 1'b0;
    n5799_o2 <= 1'b0;
    n5802_o2 <= 1'b0;
    n2068_inv <= 1'b0;
    n5831_o2 <= 1'b0;
    n5833_o2 <= 1'b0;
    n5820_o2 <= 1'b0;
    n5823_o2 <= 1'b0;
    n5824_o2 <= 1'b0;
    n5869_o2 <= 1'b0;
    n5848_o2 <= 1'b0;
    n5849_o2 <= 1'b0;
    n5856_o2 <= 1'b0;
    n5896_o2 <= 1'b0;
    n2754_o2 <= 1'b0;
    n2908_o2 <= 1'b0;
    n5892_o2 <= 1'b0;
    n5915_o2 <= 1'b0;
    n5919_o2 <= 1'b0;
    n5918_o2 <= 1'b0;
    n5920_o2 <= 1'b0;
    n5917_o2 <= 1'b0;
    lo586_buf_o2 <= 1'b0;
    n2818_o2 <= 1'b0;
    n2863_o2 <= 1'b0;
    n2134_inv <= 1'b0;
    n2725_o2 <= 1'b0;
    n3016_o2 <= 1'b0;
    n3013_o2 <= 1'b0;
    n2655_o2 <= 1'b0;
    n2149_inv <= 1'b0;
    lo562_buf_o2 <= 1'b0;
    n2155_inv <= 1'b0;
    n2531_o2 <= 1'b0;
    n2700_o2 <= 1'b0;
    n5908_o2 <= 1'b0;
    n5910_o2 <= 1'b0;
    n5912_o2 <= 1'b0;
    n5914_o2 <= 1'b0;
    n2753_o2 <= 1'b0;
    n2878_o2 <= 1'b0;
    n2182_inv <= 1'b0;
    n5934_o2 <= 1'b0;
    n5936_o2 <= 1'b0;
    n5938_o2 <= 1'b0;
    n2728_o2 <= 1'b0;
    lo358_buf_o2 <= 1'b0;
    lo418_buf_o2 <= 1'b0;
    lo474_buf_o2 <= 1'b0;
    lo554_buf_o2 <= 1'b0;
    lo558_buf_o2 <= 1'b0;
    lo574_buf_o2 <= 1'b0;
    n2215_inv <= 1'b0;
    n2218_inv <= 1'b0;
    n2221_inv <= 1'b0;
    lo450_buf_o2 <= 1'b0;
    n2910_o2 <= 1'b0;
    n2683_o2 <= 1'b0;
    n2828_o2 <= 1'b0;
    n2582_o2 <= 1'b0;
    n2600_o2 <= 1'b0;
    n2542_o2 <= 1'b0;
    n2703_o2 <= 1'b0;
    lo510_buf_o2 <= 1'b0;
    lo514_buf_o2 <= 1'b0;
    lo538_buf_o2 <= 1'b0;
    lo578_buf_o2 <= 1'b0;
    n2260_inv <= 1'b0;
    n2666_o2 <= 1'b0;
    n2667_o2 <= 1'b0;
    n2660_o2 <= 1'b0;
    n2272_inv <= 1'b0;
    lo454_buf_o2 <= 1'b0;
    n3593_o2 <= 1'b0;
    n3048_o2 <= 1'b0;
    lo410_buf_o2 <= 1'b0;
    lo502_buf_o2 <= 1'b0;
    lo506_buf_o2 <= 1'b0;
    lo550_buf_o2 <= 1'b0;
    lo570_buf_o2 <= 1'b0;
    lo582_buf_o2 <= 1'b0;
    n2302_inv <= 1'b0;
    n2305_inv <= 1'b0;
    n3499_o2 <= 1'b0;
    n2311_inv <= 1'b0;
    n2870_o2 <= 1'b0;
    n2317_inv <= 1'b0;
    n2689_o2 <= 1'b0;
    n2323_inv <= 1'b0;
    n2662_o2 <= 1'b0;
    lo350_buf_o2 <= 1'b0;
    lo498_buf_o2 <= 1'b0;
    lo518_buf_o2 <= 1'b0;
    lo522_buf_o2 <= 1'b0;
    lo598_buf_o2 <= 1'b0;
    n2344_inv <= 1'b0;
    n2347_inv <= 1'b0;
    n2350_inv <= 1'b0;
    n2353_inv <= 1'b0;
    n2356_inv <= 1'b0;
    n2359_inv <= 1'b0;
    n2872_o2 <= 1'b0;
    n3313_o2 <= 1'b0;
    n3273_o2 <= 1'b0;
    n2848_o2 <= 1'b0;
    n2893_o2 <= 1'b0;
    n3267_o2 <= 1'b0;
    n2925_o2 <= 1'b0;
    n2839_o2 <= 1'b0;
    n2831_o2 <= 1'b0;
    n2558_o2 <= 1'b0;
    n2562_o2 <= 1'b0;
    n2825_o2 <= 1'b0;
    n3263_o2 <= 1'b0;
    n3517_o2 <= 1'b0;
    n2873_o2 <= 1'b0;
    n2926_o2 <= 1'b0;
    n3261_o2 <= 1'b0;
    n3268_o2 <= 1'b0;
    n3274_o2 <= 1'b0;
    n3314_o2 <= 1'b0;
    n3571_o2 <= 1'b0;
    n2950_o2 <= 1'b0;
    n2951_o2 <= 1'b0;
    n3022_o2 <= 1'b0;
    n3023_o2 <= 1'b0;
    n3057_o2 <= 1'b0;
    n3058_o2 <= 1'b0;
    n2931_o2 <= 1'b0;
    n2911_o2 <= 1'b0;
    n2959_o2 <= 1'b0;
    n2960_o2 <= 1'b0;
    n2922_o2 <= 1'b0;
    n2888_o2 <= 1'b0;
    n2889_o2 <= 1'b0;
    n3051_o2 <= 1'b0;
    n3052_o2 <= 1'b0;
    n3063_o2 <= 1'b0;
    n2845_o2 <= 1'b0;
    n2476_inv <= 1'b0;
    n3281_o2 <= 1'b0;
    n3294_o2 <= 1'b0;
    n2885_o2 <= 1'b0;
    n2786_o2 <= 1'b0;
    n2783_o2 <= 1'b0;
    n2801_o2 <= 1'b0;
    n2572_o2 <= 1'b0;
    n2628_o2 <= 1'b0;
    n2609_o2 <= 1'b0;
    n2618_o2 <= 1'b0;
    n2637_o2 <= 1'b0;
    n2525_o2 <= 1'b0;
    n2551_o2 <= 1'b0;
    n3759_o2 <= 1'b0;
    n2994_o2 <= 1'b0;
    n3040_o2 <= 1'b0;
    n2943_o2 <= 1'b0;
    n2991_o2 <= 1'b0;
    n3034_o2 <= 1'b0;
    n2881_o2 <= 1'b0;
    n3021_o2 <= 1'b0;
    n3062_o2 <= 1'b0;
    n2763_o2 <= 1'b0;
    n2764_o2 <= 1'b0;
    n2775_o2 <= 1'b0;
    n2776_o2 <= 1'b0;
    n2968_o2 <= 1'b0;
    n2969_o2 <= 1'b0;
    n2798_o2 <= 1'b0;
    n3661_o2 <= 1'b0;
    n2694_o2 <= 1'b0;
    n2572_inv <= 1'b0;
    n2817_o2 <= 1'b0;
    n2514_o2 <= 1'b0;
    n2501_o2 <= 1'b0;
    n2584_inv <= 1'b0;
    n2505_o2 <= 1'b0;
    n2492_o2 <= 1'b0;
    lo546_buf_o2 <= 1'b0;
    lo590_buf_o2 <= 1'b0;
    lo594_buf_o2 <= 1'b0;
    n2602_inv <= 1'b0;
    n2605_inv <= 1'b0;
    n2709_o2 <= 1'b0;
    n2611_inv <= 1'b0;
    n2614_inv <= 1'b0;
    n2617_inv <= 1'b0;
    n2620_inv <= 1'b0;
    n3590_o2 <= 1'b0;
    n3591_o2 <= 1'b0;
    n2629_inv <= 1'b0;
    n3638_o2 <= 1'b0;
    n3639_o2 <= 1'b0;
    n2638_inv <= 1'b0;
    n2641_inv <= 1'b0;
    lo458_buf_o2 <= 1'b0;
    lo482_buf_o2 <= 1'b0;
    lo566_buf_o2 <= 1'b0;
    n2718_o2 <= 1'b0;
    n3707_o2 <= 1'b0;
    n3671_o2 <= 1'b0;
    n3680_o2 <= 1'b0;
    n3749_o2 <= 1'b0;
    n3716_o2 <= 1'b0;
    n3692_o2 <= 1'b0;
    n2591_o2 <= 1'b0;
    n3478_o2 <= 1'b0;
    n3610_o2 <= 1'b0;
    n3611_o2 <= 1'b0;
    n2686_inv <= 1'b0;
    n2689_inv <= 1'b0;
    n2738_o2 <= 1'b0;
    n3616_o2 <= 1'b0;
    n3617_o2 <= 1'b0;
    n3031_o2 <= 1'b0;
    n2704_inv <= 1'b0;
    n3562_o2 <= 1'b0;
    n2502_o2 <= 1'b0;
    n3560_o2 <= 1'b0;
    n3554_o2 <= 1'b0;
    n3555_o2 <= 1'b0;
    n3536_o2 <= 1'b0;
    n3537_o2 <= 1'b0;
    n3508_o2 <= 1'b0;
    n3650_o2 <= 1'b0;
    n3740_o2 <= 1'b0;
    n3484_o2 <= 1'b0;
    n2740_inv <= 1'b0;
    n2734_o2 <= 1'b0;
    n2735_o2 <= 1'b0;
    n2711_o2 <= 1'b0;
    lo585_buf_o2 <= 1'b0;
    n2719_o2 <= 1'b0;
    n2720_o2 <= 1'b0;
    n2723_o2 <= 1'b0;
    n2724_o2 <= 1'b0;
    n3624_o2 <= 1'b0;
    n3625_o2 <= 1'b0;
    n3015_o2 <= 1'b0;
    n3491_o2 <= 1'b0;
    n2779_inv <= 1'b0;
    n2811_o2 <= 1'b0;
    n3010_o2 <= 1'b0;
    n3012_o2 <= 1'b0;
    lo382_buf_o2 <= 1'b0;
    lo386_buf_o2 <= 1'b0;
    lo390_buf_o2 <= 1'b0;
    lo398_buf_o2 <= 1'b0;
    lo402_buf_o2 <= 1'b0;
    lo406_buf_o2 <= 1'b0;
    n3492_o2 <= 1'b0;
    lo366_buf_o2 <= 1'b0;
    lo374_buf_o2 <= 1'b0;
    lo426_buf_o2 <= 1'b0;
    lo494_buf_o2 <= 1'b0;
    n2653_o2 <= 1'b0;
    n2654_o2 <= 1'b0;
    n2715_o2 <= 1'b0;
    n2740_o2 <= 1'b0;
    n2682_o2 <= 1'b0;
    n2736_o2 <= 1'b0;
    lo508_buf_o2 <= 1'b0;
    lo512_buf_o2 <= 1'b0;
    lo536_buf_o2 <= 1'b0;
    lo576_buf_o2 <= 1'b0;
    lo357_buf_o2 <= 1'b0;
    lo361_buf_o2 <= 1'b0;
    lo417_buf_o2 <= 1'b0;
    lo421_buf_o2 <= 1'b0;
    lo473_buf_o2 <= 1'b0;
    lo477_buf_o2 <= 1'b0;
    lo553_buf_o2 <= 1'b0;
    lo557_buf_o2 <= 1'b0;
    lo573_buf_o2 <= 1'b0;
    lo434_buf_o2 <= 1'b0;
    lo438_buf_o2 <= 1'b0;
    lo466_buf_o2 <= 1'b0;
    lo470_buf_o2 <= 1'b0;
    lo490_buf_o2 <= 1'b0;
    n2657_o2 <= 1'b0;
    n2658_o2 <= 1'b0;
    n2663_o2 <= 1'b0;
    n2664_o2 <= 1'b0;
    n2684_o2 <= 1'b0;
    n2685_o2 <= 1'b0;
  end
endmodule


