
module mymod
(
  G1_p,
  G1_n,
  G2_p,
  G2_n,
  G3_p,
  G3_n,
  G4_p,
  G4_n,
  G5_p,
  G5_n,
  G6_p,
  G6_n,
  G7_p,
  G7_n,
  G8_p,
  G8_n,
  G9_p,
  G9_n,
  G10_p,
  G10_n,
  G11_p,
  G11_n,
  G12_p,
  G12_n,
  G13_p,
  G13_n,
  G14_p,
  G14_n,
  G15_p,
  G15_n,
  G16_p,
  G16_n,
  G17_p,
  G17_n,
  G18_p,
  G18_n,
  G19_p,
  G19_n,
  G20_p,
  G20_n,
  G21_p,
  G21_n,
  G22_p,
  G22_n,
  G23_p,
  G23_n,
  G24_p,
  G24_n,
  G25_p,
  G25_n,
  G26_p,
  G26_n,
  G27_p,
  G27_n,
  G28_p,
  G28_n,
  G29_p,
  G29_n,
  G30_p,
  G30_n,
  G31_p,
  G31_n,
  G32_p,
  G32_n,
  G33_p,
  G33_n,
  G34_p,
  G34_n,
  G35_p,
  G35_n,
  G36_p,
  G36_n,
  G426_p,
  G427_p,
  G428_p,
  G429_n,
  G430_n,
  G431_n,
  G432_n
);

  input G1_p;input G1_n;input G2_p;input G2_n;input G3_p;input G3_n;input G4_p;input G4_n;input G5_p;input G5_n;input G6_p;input G6_n;input G7_p;input G7_n;input G8_p;input G8_n;input G9_p;input G9_n;input G10_p;input G10_n;input G11_p;input G11_n;input G12_p;input G12_n;input G13_p;input G13_n;input G14_p;input G14_n;input G15_p;input G15_n;input G16_p;input G16_n;input G17_p;input G17_n;input G18_p;input G18_n;input G19_p;input G19_n;input G20_p;input G20_n;input G21_p;input G21_n;input G22_p;input G22_n;input G23_p;input G23_n;input G24_p;input G24_n;input G25_p;input G25_n;input G26_p;input G26_n;input G27_p;input G27_n;input G28_p;input G28_n;input G29_p;input G29_n;input G30_p;input G30_n;input G31_p;input G31_n;input G32_p;input G32_n;input G33_p;input G33_n;input G34_p;input G34_n;input G35_p;input G35_n;input G36_p;input G36_n;
  output G426_p;output G427_p;output G428_p;output G429_n;output G430_n;output G431_n;output G432_n;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire ffc_0_p;
  wire ffc_0_n;
  wire ffc_1_p;
  wire ffc_1_n;
  wire ffc_2_p;
  wire ffc_2_n;
  wire ffc_3_p;
  wire ffc_3_n;
  wire ffc_4_p;
  wire ffc_4_n;
  wire ffc_5_p;
  wire ffc_5_n;
  wire ffc_6_p;
  wire ffc_6_n;
  wire ffc_7_p;
  wire ffc_7_n;
  wire ffc_8_p;
  wire ffc_8_n;
  wire ffc_9_p;
  wire ffc_9_n;
  wire ffc_10_p;
  wire ffc_10_n;
  wire ffc_11_p;
  wire ffc_11_n;
  wire ffc_12_p;
  wire ffc_12_n;
  wire ffc_13_p;
  wire ffc_13_n;
  wire ffc_14_p;
  wire ffc_14_n;
  wire ffc_15_p;
  wire ffc_15_n;
  wire ffc_16_p;
  wire ffc_16_n;
  wire ffc_17_p;
  wire ffc_17_n;
  wire ffc_18_p;
  wire ffc_18_n;
  wire ffc_19_p;
  wire ffc_19_n;
  wire ffc_20_p;
  wire ffc_20_n;
  wire ffc_21_p;
  wire ffc_21_n;
  wire ffc_22_p;
  wire ffc_22_n;
  wire ffc_23_p;
  wire ffc_23_n;
  wire ffc_24_p;
  wire ffc_24_n;
  wire ffc_25_p;
  wire ffc_25_n;
  wire ffc_26_p;
  wire ffc_26_n;
  wire ffc_27_p;
  wire ffc_27_n;
  wire ffc_28_p;
  wire ffc_28_n;
  wire ffc_29_p;
  wire ffc_29_n;
  wire ffc_30_p;
  wire ffc_30_n;
  wire ffc_31_p;
  wire ffc_31_n;
  wire ffc_32_p;
  wire ffc_32_n;
  wire ffc_33_p;
  wire ffc_33_n;
  wire ffc_34_p;
  wire ffc_34_n;
  wire ffc_35_p;
  wire ffc_35_n;
  wire ffc_36_p;
  wire ffc_36_n;
  wire ffc_37_p;
  wire ffc_37_n;
  wire ffc_38_p;
  wire ffc_38_n;
  wire ffc_39_p;
  wire ffc_39_n;
  wire ffc_40_p;
  wire ffc_40_n;
  wire ffc_41_p;
  wire ffc_41_n;
  wire ffc_42_p;
  wire ffc_42_n;
  wire ffc_43_p;
  wire ffc_43_n;
  wire ffc_44_p;
  wire ffc_44_n;
  wire ffc_45_p;
  wire ffc_45_n;
  wire ffc_46_p;
  wire ffc_46_n;
  wire ffc_47_p;
  wire ffc_47_n;
  wire ffc_48_p;
  wire ffc_48_n;
  wire ffc_49_p;
  wire ffc_49_n;
  wire ffc_50_p;
  wire ffc_50_n;
  wire ffc_51_p;
  wire ffc_51_n;
  wire ffc_52_p;
  wire ffc_52_n;
  wire ffc_53_p;
  wire ffc_53_n;
  wire ffc_54_p;
  wire ffc_54_n;
  wire ffc_55_p;
  wire ffc_55_n;
  wire ffc_56_p;
  wire ffc_56_n;
  wire ffc_57_p;
  wire ffc_57_n;
  wire ffc_58_p;
  wire ffc_58_n;
  wire ffc_59_p;
  wire ffc_59_n;
  wire ffc_60_p;
  wire ffc_60_n;
  wire ffc_61_p;
  wire ffc_61_n;
  wire ffc_62_p;
  wire ffc_62_n;
  wire ffc_63_p;
  wire ffc_63_n;
  wire ffc_64_p;
  wire ffc_64_n;
  wire ffc_65_p;
  wire ffc_65_n;
  wire ffc_66_p;
  wire ffc_66_n;
  wire ffc_67_p;
  wire ffc_67_n;
  wire ffc_68_p;
  wire ffc_68_n;
  wire ffc_69_p;
  wire ffc_69_n;
  wire ffc_70_p;
  wire ffc_70_n;
  wire ffc_71_p;
  wire ffc_71_n;
  wire ffc_72_p;
  wire ffc_72_n;
  wire ffc_73_p;
  wire ffc_73_n;
  wire ffc_74_p;
  wire ffc_74_n;
  wire ffc_75_p;
  wire ffc_75_n;
  wire ffc_76_p;
  wire ffc_76_n;
  wire ffc_77_p;
  wire ffc_77_n;
  wire ffc_78_p;
  wire ffc_78_n;
  wire ffc_79_p;
  wire ffc_79_n;
  wire ffc_80_p;
  wire ffc_80_n;
  wire ffc_81_p;
  wire ffc_81_n;
  wire ffc_82_p;
  wire ffc_82_n;
  wire ffc_83_p;
  wire ffc_83_n;
  wire ffc_84_p;
  wire ffc_84_n;
  wire ffc_85_p;
  wire ffc_85_n;
  wire ffc_86_p;
  wire ffc_86_n;
  wire ffc_87_p;
  wire ffc_87_n;
  wire ffc_88_p;
  wire ffc_88_n;
  wire ffc_89_p;
  wire ffc_89_n;
  wire ffc_90_p;
  wire ffc_90_n;
  wire ffc_91_p;
  wire ffc_91_n;
  wire ffc_92_p;
  wire ffc_92_n;
  wire ffc_93_p;
  wire ffc_93_n;
  wire ffc_94_p;
  wire ffc_94_n;
  wire ffc_95_p;
  wire ffc_95_n;
  wire ffc_96_p;
  wire ffc_96_n;
  wire ffc_97_p;
  wire ffc_97_n;
  wire ffc_98_p;
  wire ffc_98_n;
  wire ffc_99_p;
  wire ffc_99_n;
  wire ffc_100_p;
  wire ffc_100_n;
  wire ffc_101_p;
  wire ffc_101_n;
  wire ffc_102_p;
  wire ffc_102_n;
  wire ffc_103_p;
  wire ffc_103_n;
  wire ffc_104_p;
  wire ffc_104_n;
  wire ffc_105_p;
  wire ffc_105_n;
  wire ffc_106_p;
  wire ffc_106_n;
  wire ffc_107_p;
  wire ffc_107_n;
  wire ffc_108_p;
  wire ffc_108_n;
  wire ffc_109_p;
  wire ffc_109_n;
  wire ffc_110_p;
  wire ffc_110_n;
  wire ffc_111_p;
  wire ffc_111_n;
  wire ffc_112_p;
  wire ffc_112_n;
  wire ffc_113_p;
  wire ffc_113_n;
  wire ffc_114_p;
  wire ffc_114_n;
  wire ffc_115_p;
  wire ffc_115_n;
  wire ffc_116_p;
  wire ffc_116_n;
  wire ffc_117_p;
  wire ffc_117_n;
  wire ffc_118_p;
  wire ffc_118_n;
  wire ffc_119_p;
  wire ffc_119_n;
  wire ffc_120_p;
  wire ffc_120_n;
  wire ffc_121_p;
  wire ffc_121_n;
  wire ffc_122_p;
  wire ffc_122_n;
  wire ffc_123_p;
  wire ffc_123_n;
  wire ffc_124_p;
  wire ffc_124_n;
  wire ffc_125_p;
  wire ffc_125_n;
  wire ffc_126_p;
  wire ffc_126_n;
  wire ffc_127_p;
  wire ffc_127_n;
  wire ffc_128_p;
  wire ffc_128_n;
  wire ffc_129_p;
  wire ffc_129_n;
  wire ffc_130_p;
  wire ffc_130_n;
  wire ffc_131_p;
  wire ffc_131_n;
  wire g169_p;
  wire g169_n;
  wire g170_p;
  wire g170_n;
  wire g171_p;
  wire g171_n;
  wire g172_p;
  wire g172_n;
  wire g173_p;
  wire g173_n;
  wire g174_p;
  wire g174_n;
  wire g175_p;
  wire g175_n;
  wire g176_p;
  wire g176_n;
  wire g177_p;
  wire g177_n;
  wire g178_p;
  wire g178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire ffc_87_n_spl_;
  wire ffc_87_n_spl_0;
  wire ffc_87_n_spl_00;
  wire ffc_87_n_spl_1;
  wire ffc_87_p_spl_;
  wire ffc_87_p_spl_0;
  wire ffc_87_p_spl_00;
  wire ffc_87_p_spl_01;
  wire ffc_87_p_spl_1;
  wire ffc_87_p_spl_10;
  wire ffc_87_p_spl_11;
  wire g175_n_spl_;
  wire g177_n_spl_;
  wire g180_n_spl_;
  wire g186_n_spl_;
  wire g186_p_spl_;
  wire g188_p_spl_;
  wire g191_n_spl_;
  wire g193_n_spl_;
  wire g195_p_spl_;
  wire g193_p_spl_;
  wire g200_p_spl_;
  wire ffc_88_p_spl_;
  wire ffc_88_p_spl_0;
  wire ffc_88_p_spl_00;
  wire ffc_88_p_spl_1;
  wire ffc_34_p_spl_;
  wire g222_n_spl_;
  wire ffc_39_p_spl_;
  wire g220_n_spl_;
  wire ffc_8_p_spl_;
  wire g214_n_spl_;
  wire ffc_23_p_spl_;
  wire g216_n_spl_;
  wire ffc_28_p_spl_;
  wire g218_n_spl_;
  wire ffc_3_p_spl_;
  wire g209_n_spl_;
  wire ffc_44_p_spl_;
  wire g212_n_spl_;
  wire ffc_18_p_spl_;
  wire g211_n_spl_;
  wire ffc_13_p_spl_;
  wire g210_n_spl_;
  wire ffc_31_p_spl_;
  wire g228_n_spl_;
  wire ffc_97_p_spl_;
  wire g226_n_spl_;
  wire ffc_94_p_spl_;
  wire g223_n_spl_;
  wire ffc_95_p_spl_;
  wire g224_n_spl_;
  wire ffc_96_p_spl_;
  wire g225_n_spl_;
  wire ffc_119_p_spl_;
  wire ffc_127_p_spl_;
  wire ffc_123_p_spl_;
  wire ffc_125_p_spl_;
  wire g233_p_spl_;
  wire g244_p_spl_;
  wire g249_p_spl_;
  wire g260_p_spl_;
  wire g265_n_spl_;
  wire g272_n_spl_;
  wire g274_p_spl_;
  wire g274_p_spl_0;
  wire g274_p_spl_00;
  wire g274_p_spl_1;
  wire g275_n_spl_;
  wire g275_n_spl_0;
  wire g275_n_spl_00;
  wire g275_n_spl_000;
  wire g275_n_spl_01;
  wire g275_n_spl_1;
  wire g275_n_spl_10;
  wire g275_n_spl_11;
  wire G6_p_spl_;
  wire G10_p_spl_;
  wire G14_p_spl_;
  wire G34_p_spl_;

  orX
  g_g169_n
  (
    .dout(g169_n),
    .din1(ffc_46_p),
    .din2(ffc_47_p)
  );


  orX
  g_g170_n
  (
    .dout(g170_n),
    .din1(ffc_48_p),
    .din2(ffc_49_p)
  );


  orX
  g_g171_n
  (
    .dout(g171_n),
    .din1(ffc_79_p),
    .din2(ffc_80_p)
  );


  orX
  g_g172_n
  (
    .dout(g172_n),
    .din1(ffc_4_n),
    .din2(ffc_87_n_spl_00)
  );


  andX
  g_g173_p
  (
    .dout(g173_p),
    .din1(ffc_50_p),
    .din2(g172_n)
  );


  andX
  g_g174_p
  (
    .dout(g174_p),
    .din1(ffc_40_p),
    .din2(ffc_87_p_spl_00)
  );


  orX
  g_g175_n
  (
    .dout(g175_n),
    .din1(ffc_57_n),
    .din2(g174_p)
  );


  andX
  g_g176_p
  (
    .dout(g176_p),
    .din1(ffc_35_p),
    .din2(ffc_87_p_spl_00)
  );


  orX
  g_g176_n
  (
    .dout(g176_n),
    .din1(ffc_35_n),
    .din2(ffc_87_n_spl_00)
  );


  andX
  g_g177_p
  (
    .dout(g177_p),
    .din1(ffc_60_p),
    .din2(g176_n)
  );


  orX
  g_g177_n
  (
    .dout(g177_n),
    .din1(ffc_60_n),
    .din2(g176_p)
  );


  andX
  g_g178_p
  (
    .dout(g178_p),
    .din1(g175_n_spl_),
    .din2(g177_n_spl_)
  );


  andX
  g_g179_p
  (
    .dout(g179_p),
    .din1(ffc_29_p),
    .din2(ffc_87_p_spl_01)
  );


  orX
  g_g180_n
  (
    .dout(g180_n),
    .din1(ffc_56_n),
    .din2(g179_p)
  );


  andX
  g_g181_p
  (
    .dout(g181_p),
    .din1(ffc_45_p),
    .din2(ffc_87_p_spl_01)
  );


  orX
  g_g182_n
  (
    .dout(g182_n),
    .din1(ffc_53_n),
    .din2(g181_p)
  );


  andX
  g_g183_p
  (
    .dout(g183_p),
    .din1(g180_n_spl_),
    .din2(g182_n)
  );


  andX
  g_g184_p
  (
    .dout(g184_p),
    .din1(g178_p),
    .din2(g183_p)
  );


  andX
  g_g185_p
  (
    .dout(g185_p),
    .din1(ffc_14_p),
    .din2(ffc_87_p_spl_10)
  );


  orX
  g_g185_n
  (
    .dout(g185_n),
    .din1(ffc_14_n),
    .din2(ffc_87_n_spl_0)
  );


  andX
  g_g186_p
  (
    .dout(g186_p),
    .din1(ffc_51_p),
    .din2(g185_n)
  );


  orX
  g_g186_n
  (
    .dout(g186_n),
    .din1(ffc_51_n),
    .din2(g185_p)
  );


  andX
  g_g187_p
  (
    .dout(g187_p),
    .din1(ffc_24_p),
    .din2(ffc_87_p_spl_10)
  );


  orX
  g_g187_n
  (
    .dout(g187_n),
    .din1(ffc_24_n),
    .din2(ffc_87_n_spl_1)
  );


  andX
  g_g188_p
  (
    .dout(g188_p),
    .din1(ffc_55_p),
    .din2(g187_n)
  );


  orX
  g_g188_n
  (
    .dout(g188_n),
    .din1(ffc_55_n),
    .din2(g187_p)
  );


  andX
  g_g189_p
  (
    .dout(g189_p),
    .din1(g186_n_spl_),
    .din2(g188_n)
  );


  orX
  g_g189_n
  (
    .dout(g189_n),
    .din1(g186_p_spl_),
    .din2(g188_p_spl_)
  );


  andX
  g_g190_p
  (
    .dout(g190_p),
    .din1(ffc_9_p),
    .din2(ffc_87_p_spl_11)
  );


  orX
  g_g191_n
  (
    .dout(g191_n),
    .din1(ffc_54_n),
    .din2(g190_p)
  );


  andX
  g_g192_p
  (
    .dout(g192_p),
    .din1(ffc_19_p),
    .din2(ffc_87_p_spl_11)
  );


  orX
  g_g192_n
  (
    .dout(g192_n),
    .din1(ffc_19_n),
    .din2(ffc_87_n_spl_1)
  );


  andX
  g_g193_p
  (
    .dout(g193_p),
    .din1(ffc_52_p),
    .din2(g192_n)
  );


  orX
  g_g193_n
  (
    .dout(g193_n),
    .din1(ffc_52_n),
    .din2(g192_p)
  );


  andX
  g_g194_p
  (
    .dout(g194_p),
    .din1(g191_n_spl_),
    .din2(g193_n_spl_)
  );


  andX
  g_g195_p
  (
    .dout(g195_p),
    .din1(g189_p),
    .din2(g194_p)
  );


  andX
  g_g196_p
  (
    .dout(g196_p),
    .din1(g184_p),
    .din2(g195_p_spl_)
  );


  orX
  g_g197_n
  (
    .dout(g197_n),
    .din1(g173_p),
    .din2(g196_p)
  );


  orX
  g_g198_n
  (
    .dout(g198_n),
    .din1(g180_n_spl_),
    .din2(g193_p_spl_)
  );


  orX
  g_g199_n
  (
    .dout(g199_n),
    .din1(g189_n),
    .din2(g198_n)
  );


  andX
  g_g200_p
  (
    .dout(g200_p),
    .din1(g191_n_spl_),
    .din2(g199_n)
  );


  orX
  g_g201_n
  (
    .dout(g201_n),
    .din1(g188_p_spl_),
    .din2(g193_p_spl_)
  );


  orX
  g_g202_n
  (
    .dout(g202_n),
    .din1(g177_n_spl_),
    .din2(g201_n)
  );


  andX
  g_g203_p
  (
    .dout(g203_p),
    .din1(g186_n_spl_),
    .din2(g202_n)
  );


  andX
  g_g204_p
  (
    .dout(g204_p),
    .din1(g200_p_spl_),
    .din2(g203_p)
  );


  orX
  g_g205_n
  (
    .dout(g205_n),
    .din1(g175_n_spl_),
    .din2(g177_p)
  );


  andX
  g_g206_p
  (
    .dout(g206_p),
    .din1(g193_n_spl_),
    .din2(g205_n)
  );


  orX
  g_g207_n
  (
    .dout(g207_n),
    .din1(g186_p_spl_),
    .din2(g206_p)
  );


  andX
  g_g208_p
  (
    .dout(g208_p),
    .din1(g200_p_spl_),
    .din2(g207_n)
  );


  orX
  g_g209_n
  (
    .dout(g209_n),
    .din1(ffc_64_n),
    .din2(ffc_90_p)
  );


  orX
  g_g210_n
  (
    .dout(g210_n),
    .din1(ffc_61_n),
    .din2(ffc_91_p)
  );


  orX
  g_g211_n
  (
    .dout(g211_n),
    .din1(ffc_62_n),
    .din2(ffc_92_p)
  );


  orX
  g_g212_n
  (
    .dout(g212_n),
    .din1(ffc_63_n),
    .din2(ffc_93_p)
  );


  andX
  g_g213_p
  (
    .dout(g213_p),
    .din1(ffc_65_p),
    .din2(ffc_88_p_spl_00)
  );


  orX
  g_g214_n
  (
    .dout(g214_n),
    .din1(ffc_69_n),
    .din2(g213_p)
  );


  andX
  g_g215_p
  (
    .dout(g215_p),
    .din1(ffc_66_p),
    .din2(ffc_88_p_spl_00)
  );


  orX
  g_g216_n
  (
    .dout(g216_n),
    .din1(ffc_70_n),
    .din2(g215_p)
  );


  andX
  g_g217_p
  (
    .dout(g217_p),
    .din1(ffc_67_p),
    .din2(ffc_88_p_spl_0)
  );


  orX
  g_g218_n
  (
    .dout(g218_n),
    .din1(ffc_71_n),
    .din2(g217_p)
  );


  andX
  g_g219_p
  (
    .dout(g219_p),
    .din1(ffc_68_p),
    .din2(ffc_88_p_spl_1)
  );


  orX
  g_g220_n
  (
    .dout(g220_n),
    .din1(ffc_72_n),
    .din2(g219_p)
  );


  andX
  g_g221_p
  (
    .dout(g221_p),
    .din1(ffc_73_p),
    .din2(ffc_88_p_spl_1)
  );


  orX
  g_g222_n
  (
    .dout(g222_n),
    .din1(ffc_74_n),
    .din2(g221_p)
  );


  orX
  g_g223_n
  (
    .dout(g223_n),
    .din1(ffc_75_n),
    .din2(ffc_98_p)
  );


  orX
  g_g224_n
  (
    .dout(g224_n),
    .din1(ffc_76_n),
    .din2(ffc_103_p)
  );


  orX
  g_g225_n
  (
    .dout(g225_n),
    .din1(ffc_77_n),
    .din2(ffc_104_p)
  );


  orX
  g_g226_n
  (
    .dout(g226_n),
    .din1(ffc_78_n),
    .din2(ffc_105_p)
  );


  andX
  g_g227_p
  (
    .dout(g227_p),
    .din1(ffc_81_p),
    .din2(ffc_89_p)
  );


  orX
  g_g228_n
  (
    .dout(g228_n),
    .din1(ffc_82_n),
    .din2(g227_p)
  );


  orX
  g_g229_n
  (
    .dout(g229_n),
    .din1(ffc_34_p_spl_),
    .din2(g222_n_spl_)
  );


  orX
  g_g230_n
  (
    .dout(g230_n),
    .din1(ffc_39_p_spl_),
    .din2(g220_n_spl_)
  );


  orX
  g_g231_n
  (
    .dout(g231_n),
    .din1(ffc_8_p_spl_),
    .din2(g214_n_spl_)
  );


  andX
  g_g232_p
  (
    .dout(g232_p),
    .din1(g230_n),
    .din2(g231_n)
  );


  andX
  g_g233_p
  (
    .dout(g233_p),
    .din1(g229_n),
    .din2(g232_p)
  );


  orX
  g_g234_n
  (
    .dout(g234_n),
    .din1(ffc_23_p_spl_),
    .din2(g216_n_spl_)
  );


  orX
  g_g235_n
  (
    .dout(g235_n),
    .din1(ffc_28_p_spl_),
    .din2(g218_n_spl_)
  );


  andX
  g_g236_p
  (
    .dout(g236_p),
    .din1(g234_n),
    .din2(g235_n)
  );


  orX
  g_g237_n
  (
    .dout(g237_n),
    .din1(ffc_3_p_spl_),
    .din2(g209_n_spl_)
  );


  orX
  g_g238_n
  (
    .dout(g238_n),
    .din1(ffc_44_p_spl_),
    .din2(g212_n_spl_)
  );


  andX
  g_g239_p
  (
    .dout(g239_p),
    .din1(g237_n),
    .din2(g238_n)
  );


  orX
  g_g240_n
  (
    .dout(g240_n),
    .din1(ffc_18_p_spl_),
    .din2(g211_n_spl_)
  );


  orX
  g_g241_n
  (
    .dout(g241_n),
    .din1(ffc_13_p_spl_),
    .din2(g210_n_spl_)
  );


  andX
  g_g242_p
  (
    .dout(g242_p),
    .din1(g240_n),
    .din2(g241_n)
  );


  andX
  g_g243_p
  (
    .dout(g243_p),
    .din1(g239_p),
    .din2(g242_p)
  );


  andX
  g_g244_p
  (
    .dout(g244_p),
    .din1(g236_p),
    .din2(g243_p)
  );


  orX
  g_g245_n
  (
    .dout(g245_n),
    .din1(ffc_31_p_spl_),
    .din2(g228_n_spl_)
  );


  orX
  g_g246_n
  (
    .dout(g246_n),
    .din1(ffc_97_p_spl_),
    .din2(g226_n_spl_)
  );


  orX
  g_g247_n
  (
    .dout(g247_n),
    .din1(ffc_94_p_spl_),
    .din2(g223_n_spl_)
  );


  andX
  g_g248_p
  (
    .dout(g248_p),
    .din1(g246_n),
    .din2(g247_n)
  );


  andX
  g_g249_p
  (
    .dout(g249_p),
    .din1(g245_n),
    .din2(g248_p)
  );


  orX
  g_g250_n
  (
    .dout(g250_n),
    .din1(ffc_95_p_spl_),
    .din2(g224_n_spl_)
  );


  orX
  g_g251_n
  (
    .dout(g251_n),
    .din1(ffc_96_p_spl_),
    .din2(g225_n_spl_)
  );


  andX
  g_g252_p
  (
    .dout(g252_p),
    .din1(g250_n),
    .din2(g251_n)
  );


  orX
  g_g253_n
  (
    .dout(g253_n),
    .din1(ffc_102_n),
    .din2(ffc_106_p)
  );


  orX
  g_g254_n
  (
    .dout(g254_n),
    .din1(ffc_101_n),
    .din2(ffc_109_p)
  );


  andX
  g_g255_p
  (
    .dout(g255_p),
    .din1(g253_n),
    .din2(g254_n)
  );


  orX
  g_g256_n
  (
    .dout(g256_n),
    .din1(ffc_100_n),
    .din2(ffc_108_p)
  );


  orX
  g_g257_n
  (
    .dout(g257_n),
    .din1(ffc_99_n),
    .din2(ffc_107_p)
  );


  andX
  g_g258_p
  (
    .dout(g258_p),
    .din1(g256_n),
    .din2(g257_n)
  );


  andX
  g_g259_p
  (
    .dout(g259_p),
    .din1(g255_p),
    .din2(g258_p)
  );


  andX
  g_g260_p
  (
    .dout(g260_p),
    .din1(g252_p),
    .din2(g259_p)
  );


  andX
  g_g261_p
  (
    .dout(g261_p),
    .din1(ffc_118_n),
    .din2(ffc_119_p_spl_)
  );


  andX
  g_g262_p
  (
    .dout(g262_p),
    .din1(ffc_126_n),
    .din2(ffc_127_p_spl_)
  );


  andX
  g_g263_p
  (
    .dout(g263_p),
    .din1(ffc_120_n),
    .din2(ffc_121_p)
  );


  orX
  g_g264_n
  (
    .dout(g264_n),
    .din1(g262_p),
    .din2(g263_p)
  );


  orX
  g_g265_n
  (
    .dout(g265_n),
    .din1(g261_p),
    .din2(g264_n)
  );


  andX
  g_g266_p
  (
    .dout(g266_p),
    .din1(ffc_122_n),
    .din2(ffc_123_p_spl_)
  );


  andX
  g_g267_p
  (
    .dout(g267_p),
    .din1(ffc_124_n),
    .din2(ffc_125_p_spl_)
  );


  orX
  g_g268_n
  (
    .dout(g268_n),
    .din1(g266_p),
    .din2(g267_p)
  );


  orX
  g_g269_n
  (
    .dout(g269_n),
    .din1(ffc_128_p),
    .din2(ffc_131_p)
  );


  orX
  g_g270_n
  (
    .dout(g270_n),
    .din1(ffc_129_p),
    .din2(ffc_130_p)
  );


  orX
  g_g271_n
  (
    .dout(g271_n),
    .din1(g269_n),
    .din2(g270_n)
  );


  orX
  g_g272_n
  (
    .dout(g272_n),
    .din1(g268_n),
    .din2(g271_n)
  );


  andX
  g_g273_p
  (
    .dout(g273_p),
    .din1(g233_p_spl_),
    .din2(g244_p_spl_)
  );


  andX
  g_g274_p
  (
    .dout(g274_p),
    .din1(g249_p_spl_),
    .din2(g260_p_spl_)
  );


  orX
  g_g275_n
  (
    .dout(g275_n),
    .din1(g265_n_spl_),
    .din2(g272_n_spl_)
  );


  orX
  g_g276_n
  (
    .dout(g276_n),
    .din1(ffc_106_n),
    .din2(g274_p_spl_00)
  );


  orX
  g_g277_n
  (
    .dout(g277_n),
    .din1(ffc_107_n),
    .din2(g274_p_spl_00)
  );


  orX
  g_g278_n
  (
    .dout(g278_n),
    .din1(ffc_108_n),
    .din2(g274_p_spl_0)
  );


  orX
  g_g279_n
  (
    .dout(g279_n),
    .din1(ffc_109_n),
    .din2(g274_p_spl_1)
  );


  andX
  g_g280_p
  (
    .dout(g280_p),
    .din1(ffc_110_p),
    .din2(g275_n_spl_000)
  );


  andX
  g_g281_p
  (
    .dout(g281_p),
    .din1(ffc_112_p),
    .din2(g275_n_spl_000)
  );


  orX
  g_g282_n
  (
    .dout(g282_n),
    .din1(ffc_113_n),
    .din2(g281_p)
  );


  andX
  g_g283_p
  (
    .dout(g283_p),
    .din1(ffc_114_p),
    .din2(g275_n_spl_00)
  );


  orX
  g_g284_n
  (
    .dout(g284_n),
    .din1(ffc_115_n),
    .din2(g283_p)
  );


  andX
  g_g285_p
  (
    .dout(g285_p),
    .din1(ffc_116_p),
    .din2(g275_n_spl_01)
  );


  orX
  g_g286_n
  (
    .dout(g286_n),
    .din1(ffc_117_n),
    .din2(g285_p)
  );


  andX
  g_g287_p
  (
    .dout(g287_p),
    .din1(ffc_120_p),
    .din2(g275_n_spl_01)
  );


  orX
  g_g288_n
  (
    .dout(g288_n),
    .din1(ffc_121_n),
    .din2(g287_p)
  );


  andX
  g_g289_p
  (
    .dout(g289_p),
    .din1(ffc_122_p),
    .din2(g275_n_spl_10)
  );


  andX
  g_g290_p
  (
    .dout(g290_p),
    .din1(ffc_124_p),
    .din2(g275_n_spl_10)
  );


  andX
  g_g291_p
  (
    .dout(g291_p),
    .din1(ffc_126_p),
    .din2(g275_n_spl_11)
  );


  andX
  g_g292_p
  (
    .dout(g292_p),
    .din1(G4_n),
    .din2(G6_p_spl_)
  );


  andX
  g_g293_p
  (
    .dout(g293_p),
    .din1(G8_n),
    .din2(G10_p_spl_)
  );


  andX
  g_g294_p
  (
    .dout(g294_p),
    .din1(G12_n),
    .din2(G14_p_spl_)
  );


  andX
  g_g295_p
  (
    .dout(g295_p),
    .din1(G32_n),
    .din2(G34_p_spl_)
  );


  buf

  (
    G426_p,
    g169_n
  );


  buf

  (
    G427_p,
    g170_n
  );


  buf

  (
    G428_p,
    g171_n
  );


  buf

  (
    G429_n,
    g197_n
  );


  buf

  (
    G430_n,
    g195_p_spl_
  );


  buf

  (
    G431_n,
    g204_p
  );


  buf

  (
    G432_n,
    g208_p
  );


  DROC
  ffc_0
  (
    .doutp(ffc_0_p),
    .doutn(ffc_0_n),
    .din(G3_p)
  );


  DROC
  ffc_1
  (
    .doutp(ffc_1_p),
    .doutn(ffc_1_n),
    .din(G5_p)
  );


  DROC
  ffc_2
  (
    .doutp(ffc_2_p),
    .doutn(ffc_2_n),
    .din(ffc_1_p)
  );


  DROC
  ffc_3
  (
    .doutp(ffc_3_p),
    .doutn(ffc_3_n),
    .din(ffc_2_p)
  );


  DROC
  ffc_4
  (
    .doutp(ffc_4_p),
    .doutn(ffc_4_n),
    .din(ffc_3_p_spl_)
  );


  DROC
  ffc_5
  (
    .doutp(ffc_5_p),
    .doutn(ffc_5_n),
    .din(G7_p)
  );


  DROC
  ffc_6
  (
    .doutp(ffc_6_p),
    .doutn(ffc_6_n),
    .din(G9_p)
  );


  DROC
  ffc_7
  (
    .doutp(ffc_7_p),
    .doutn(ffc_7_n),
    .din(ffc_6_p)
  );


  DROC
  ffc_8
  (
    .doutp(ffc_8_p),
    .doutn(ffc_8_n),
    .din(ffc_7_p)
  );


  DROC
  ffc_9
  (
    .doutp(ffc_9_p),
    .doutn(ffc_9_n),
    .din(ffc_8_p_spl_)
  );


  DROC
  ffc_10
  (
    .doutp(ffc_10_p),
    .doutn(ffc_10_n),
    .din(G11_p)
  );


  DROC
  ffc_11
  (
    .doutp(ffc_11_p),
    .doutn(ffc_11_n),
    .din(G13_p)
  );


  DROC
  ffc_12
  (
    .doutp(ffc_12_p),
    .doutn(ffc_12_n),
    .din(ffc_11_p)
  );


  DROC
  ffc_13
  (
    .doutp(ffc_13_p),
    .doutn(ffc_13_n),
    .din(ffc_12_p)
  );


  DROC
  ffc_14
  (
    .doutp(ffc_14_p),
    .doutn(ffc_14_n),
    .din(ffc_13_p_spl_)
  );


  DROC
  ffc_15
  (
    .doutp(ffc_15_p),
    .doutn(ffc_15_n),
    .din(G15_p)
  );


  DROC
  ffc_16
  (
    .doutp(ffc_16_p),
    .doutn(ffc_16_n),
    .din(G17_p)
  );


  DROC
  ffc_17
  (
    .doutp(ffc_17_p),
    .doutn(ffc_17_n),
    .din(ffc_16_p)
  );


  DROC
  ffc_18
  (
    .doutp(ffc_18_p),
    .doutn(ffc_18_n),
    .din(ffc_17_p)
  );


  DROC
  ffc_19
  (
    .doutp(ffc_19_p),
    .doutn(ffc_19_n),
    .din(ffc_18_p_spl_)
  );


  DROC
  ffc_20
  (
    .doutp(ffc_20_p),
    .doutn(ffc_20_n),
    .din(G19_p)
  );


  DROC
  ffc_21
  (
    .doutp(ffc_21_p),
    .doutn(ffc_21_n),
    .din(G21_p)
  );


  DROC
  ffc_22
  (
    .doutp(ffc_22_p),
    .doutn(ffc_22_n),
    .din(ffc_21_p)
  );


  DROC
  ffc_23
  (
    .doutp(ffc_23_p),
    .doutn(ffc_23_n),
    .din(ffc_22_p)
  );


  DROC
  ffc_24
  (
    .doutp(ffc_24_p),
    .doutn(ffc_24_n),
    .din(ffc_23_p_spl_)
  );


  DROC
  ffc_25
  (
    .doutp(ffc_25_p),
    .doutn(ffc_25_n),
    .din(G23_p)
  );


  DROC
  ffc_26
  (
    .doutp(ffc_26_p),
    .doutn(ffc_26_n),
    .din(G25_p)
  );


  DROC
  ffc_27
  (
    .doutp(ffc_27_p),
    .doutn(ffc_27_n),
    .din(ffc_26_p)
  );


  DROC
  ffc_28
  (
    .doutp(ffc_28_p),
    .doutn(ffc_28_n),
    .din(ffc_27_p)
  );


  DROC
  ffc_29
  (
    .doutp(ffc_29_p),
    .doutn(ffc_29_n),
    .din(ffc_28_p_spl_)
  );


  DROC
  ffc_30
  (
    .doutp(ffc_30_p),
    .doutn(ffc_30_n),
    .din(G27_p)
  );


  DROC
  ffc_31
  (
    .doutp(ffc_31_p),
    .doutn(ffc_31_n),
    .din(ffc_30_p)
  );


  DROC
  ffc_32
  (
    .doutp(ffc_32_p),
    .doutn(ffc_32_n),
    .din(G29_p)
  );


  DROC
  ffc_33
  (
    .doutp(ffc_33_p),
    .doutn(ffc_33_n),
    .din(ffc_32_p)
  );


  DROC
  ffc_34
  (
    .doutp(ffc_34_p),
    .doutn(ffc_34_n),
    .din(ffc_33_p)
  );


  DROC
  ffc_35
  (
    .doutp(ffc_35_p),
    .doutn(ffc_35_n),
    .din(ffc_34_p_spl_)
  );


  DROC
  ffc_36
  (
    .doutp(ffc_36_p),
    .doutn(ffc_36_n),
    .din(G31_p)
  );


  DROC
  ffc_37
  (
    .doutp(ffc_37_p),
    .doutn(ffc_37_n),
    .din(G33_p)
  );


  DROC
  ffc_38
  (
    .doutp(ffc_38_p),
    .doutn(ffc_38_n),
    .din(ffc_37_p)
  );


  DROC
  ffc_39
  (
    .doutp(ffc_39_p),
    .doutn(ffc_39_n),
    .din(ffc_38_p)
  );


  DROC
  ffc_40
  (
    .doutp(ffc_40_p),
    .doutn(ffc_40_n),
    .din(ffc_39_p_spl_)
  );


  DROC
  ffc_41
  (
    .doutp(ffc_41_p),
    .doutn(ffc_41_n),
    .din(G35_p)
  );


  DROC
  ffc_42
  (
    .doutp(ffc_42_p),
    .doutn(ffc_42_n),
    .din(G36_p)
  );


  DROC
  ffc_43
  (
    .doutp(ffc_43_p),
    .doutn(ffc_43_n),
    .din(ffc_42_p)
  );


  DROC
  ffc_44
  (
    .doutp(ffc_44_p),
    .doutn(ffc_44_n),
    .din(ffc_43_p)
  );


  DROC
  ffc_45
  (
    .doutp(ffc_45_p),
    .doutn(ffc_45_n),
    .din(ffc_44_p_spl_)
  );


  DROC
  ffc_46
  (
    .doutp(ffc_46_p),
    .doutn(ffc_46_n),
    .din(ffc_58_p)
  );


  DROC
  ffc_47
  (
    .doutp(ffc_47_p),
    .doutn(ffc_47_n),
    .din(ffc_59_p)
  );


  DROC
  ffc_48
  (
    .doutp(ffc_48_p),
    .doutn(ffc_48_n),
    .din(ffc_83_p)
  );


  DROC
  ffc_49
  (
    .doutp(ffc_49_p),
    .doutn(ffc_49_n),
    .din(ffc_84_p)
  );


  DROC
  ffc_50
  (
    .doutp(ffc_50_n),
    .doutn(ffc_50_p),
    .din(g209_n_spl_)
  );


  DROC
  ffc_51
  (
    .doutp(ffc_51_n),
    .doutn(ffc_51_p),
    .din(g210_n_spl_)
  );


  DROC
  ffc_52
  (
    .doutp(ffc_52_n),
    .doutn(ffc_52_p),
    .din(g211_n_spl_)
  );


  DROC
  ffc_53
  (
    .doutp(ffc_53_n),
    .doutn(ffc_53_p),
    .din(g212_n_spl_)
  );


  DROC
  ffc_54
  (
    .doutp(ffc_54_n),
    .doutn(ffc_54_p),
    .din(g214_n_spl_)
  );


  DROC
  ffc_55
  (
    .doutp(ffc_55_n),
    .doutn(ffc_55_p),
    .din(g216_n_spl_)
  );


  DROC
  ffc_56
  (
    .doutp(ffc_56_n),
    .doutn(ffc_56_p),
    .din(g218_n_spl_)
  );


  DROC
  ffc_57
  (
    .doutp(ffc_57_n),
    .doutn(ffc_57_p),
    .din(g220_n_spl_)
  );


  DROC
  ffc_58
  (
    .doutp(ffc_58_p),
    .doutn(ffc_58_n),
    .din(ffc_85_p)
  );


  DROC
  ffc_59
  (
    .doutp(ffc_59_p),
    .doutn(ffc_59_n),
    .din(ffc_86_p)
  );


  DROC
  ffc_60
  (
    .doutp(ffc_60_n),
    .doutn(ffc_60_p),
    .din(g222_n_spl_)
  );


  DROC
  ffc_61
  (
    .doutp(ffc_61_p),
    .doutn(ffc_61_n),
    .din(ffc_99_p)
  );


  DROC
  ffc_62
  (
    .doutp(ffc_62_p),
    .doutn(ffc_62_n),
    .din(ffc_100_p)
  );


  DROC
  ffc_63
  (
    .doutp(ffc_63_p),
    .doutn(ffc_63_n),
    .din(ffc_101_p)
  );


  DROC
  ffc_64
  (
    .doutp(ffc_64_p),
    .doutn(ffc_64_n),
    .din(ffc_102_p)
  );


  DROC
  ffc_65
  (
    .doutp(ffc_65_p),
    .doutn(ffc_65_n),
    .din(ffc_94_p_spl_)
  );


  DROC
  ffc_66
  (
    .doutp(ffc_66_p),
    .doutn(ffc_66_n),
    .din(ffc_95_p_spl_)
  );


  DROC
  ffc_67
  (
    .doutp(ffc_67_p),
    .doutn(ffc_67_n),
    .din(ffc_96_p_spl_)
  );


  DROC
  ffc_68
  (
    .doutp(ffc_68_p),
    .doutn(ffc_68_n),
    .din(ffc_97_p_spl_)
  );


  DROC
  ffc_69
  (
    .doutp(ffc_69_n),
    .doutn(ffc_69_p),
    .din(g223_n_spl_)
  );


  DROC
  ffc_70
  (
    .doutp(ffc_70_n),
    .doutn(ffc_70_p),
    .din(g224_n_spl_)
  );


  DROC
  ffc_71
  (
    .doutp(ffc_71_n),
    .doutn(ffc_71_p),
    .din(g225_n_spl_)
  );


  DROC
  ffc_72
  (
    .doutp(ffc_72_n),
    .doutn(ffc_72_p),
    .din(g226_n_spl_)
  );


  DROC
  ffc_73
  (
    .doutp(ffc_73_p),
    .doutn(ffc_73_n),
    .din(ffc_31_p_spl_)
  );


  DROC
  ffc_74
  (
    .doutp(ffc_74_n),
    .doutn(ffc_74_p),
    .din(g228_n_spl_)
  );


  DROC
  ffc_75
  (
    .doutp(ffc_75_p),
    .doutn(ffc_75_n),
    .din(ffc_111_p)
  );


  DROC
  ffc_76
  (
    .doutp(ffc_76_p),
    .doutn(ffc_76_n),
    .din(ffc_123_p_spl_)
  );


  DROC
  ffc_77
  (
    .doutp(ffc_77_p),
    .doutn(ffc_77_n),
    .din(ffc_125_p_spl_)
  );


  DROC
  ffc_78
  (
    .doutp(ffc_78_p),
    .doutn(ffc_78_n),
    .din(ffc_127_p_spl_)
  );


  DROC
  ffc_79
  (
    .doutp(ffc_79_n),
    .doutn(ffc_79_p),
    .din(g233_p_spl_)
  );


  DROC
  ffc_80
  (
    .doutp(ffc_80_n),
    .doutn(ffc_80_p),
    .din(g244_p_spl_)
  );


  DROC
  ffc_81
  (
    .doutp(ffc_81_p),
    .doutn(ffc_81_n),
    .din(ffc_118_p)
  );


  DROC
  ffc_82
  (
    .doutp(ffc_82_p),
    .doutn(ffc_82_n),
    .din(ffc_119_p_spl_)
  );


  DROC
  ffc_83
  (
    .doutp(ffc_83_n),
    .doutn(ffc_83_p),
    .din(g249_p_spl_)
  );


  DROC
  ffc_84
  (
    .doutp(ffc_84_n),
    .doutn(ffc_84_p),
    .din(g260_p_spl_)
  );


  DROC
  ffc_85
  (
    .doutp(ffc_85_p),
    .doutn(ffc_85_n),
    .din(g265_n_spl_)
  );


  DROC
  ffc_86
  (
    .doutp(ffc_86_p),
    .doutn(ffc_86_n),
    .din(g272_n_spl_)
  );


  DROC
  ffc_87
  (
    .doutp(ffc_87_n),
    .doutn(ffc_87_p),
    .din(g273_p)
  );


  DROC
  ffc_88
  (
    .doutp(ffc_88_n),
    .doutn(ffc_88_p),
    .din(g274_p_spl_1)
  );


  DROC
  ffc_89
  (
    .doutp(ffc_89_p),
    .doutn(ffc_89_n),
    .din(g275_n_spl_11)
  );


  DROC
  ffc_90
  (
    .doutp(ffc_90_n),
    .doutn(ffc_90_p),
    .din(g276_n)
  );


  DROC
  ffc_91
  (
    .doutp(ffc_91_n),
    .doutn(ffc_91_p),
    .din(g277_n)
  );


  DROC
  ffc_92
  (
    .doutp(ffc_92_n),
    .doutn(ffc_92_p),
    .din(g278_n)
  );


  DROC
  ffc_93
  (
    .doutp(ffc_93_n),
    .doutn(ffc_93_p),
    .din(g279_n)
  );


  DROC
  ffc_94
  (
    .doutp(ffc_94_p),
    .doutn(ffc_94_n),
    .din(ffc_5_p)
  );


  DROC
  ffc_95
  (
    .doutp(ffc_95_p),
    .doutn(ffc_95_n),
    .din(ffc_20_p)
  );


  DROC
  ffc_96
  (
    .doutp(ffc_96_p),
    .doutn(ffc_96_n),
    .din(ffc_25_p)
  );


  DROC
  ffc_97
  (
    .doutp(ffc_97_p),
    .doutn(ffc_97_n),
    .din(ffc_36_p)
  );


  DROC
  ffc_98
  (
    .doutp(ffc_98_p),
    .doutn(ffc_98_n),
    .din(g280_p)
  );


  DROC
  ffc_99
  (
    .doutp(ffc_99_n),
    .doutn(ffc_99_p),
    .din(g282_n)
  );


  DROC
  ffc_100
  (
    .doutp(ffc_100_n),
    .doutn(ffc_100_p),
    .din(g284_n)
  );


  DROC
  ffc_101
  (
    .doutp(ffc_101_n),
    .doutn(ffc_101_p),
    .din(g286_n)
  );


  DROC
  ffc_102
  (
    .doutp(ffc_102_n),
    .doutn(ffc_102_p),
    .din(g288_n)
  );


  DROC
  ffc_103
  (
    .doutp(ffc_103_p),
    .doutn(ffc_103_n),
    .din(g289_p)
  );


  DROC
  ffc_104
  (
    .doutp(ffc_104_p),
    .doutn(ffc_104_n),
    .din(g290_p)
  );


  DROC
  ffc_105
  (
    .doutp(ffc_105_p),
    .doutn(ffc_105_n),
    .din(g291_p)
  );


  DROC
  ffc_106
  (
    .doutp(ffc_106_p),
    .doutn(ffc_106_n),
    .din(ffc_0_p)
  );


  DROC
  ffc_107
  (
    .doutp(ffc_107_p),
    .doutn(ffc_107_n),
    .din(ffc_10_p)
  );


  DROC
  ffc_108
  (
    .doutp(ffc_108_p),
    .doutn(ffc_108_n),
    .din(ffc_15_p)
  );


  DROC
  ffc_109
  (
    .doutp(ffc_109_p),
    .doutn(ffc_109_n),
    .din(ffc_41_p)
  );


  DROC
  ffc_110
  (
    .doutp(ffc_110_p),
    .doutn(ffc_110_n),
    .din(G4_p)
  );


  DROC
  ffc_111
  (
    .doutp(ffc_111_p),
    .doutn(ffc_111_n),
    .din(G6_p_spl_)
  );


  DROC
  ffc_112
  (
    .doutp(ffc_112_p),
    .doutn(ffc_112_n),
    .din(G8_p)
  );


  DROC
  ffc_113
  (
    .doutp(ffc_113_p),
    .doutn(ffc_113_n),
    .din(G10_p_spl_)
  );


  DROC
  ffc_114
  (
    .doutp(ffc_114_p),
    .doutn(ffc_114_n),
    .din(G12_p)
  );


  DROC
  ffc_115
  (
    .doutp(ffc_115_p),
    .doutn(ffc_115_n),
    .din(G14_p_spl_)
  );


  DROC
  ffc_116
  (
    .doutp(ffc_116_p),
    .doutn(ffc_116_n),
    .din(G32_p)
  );


  DROC
  ffc_117
  (
    .doutp(ffc_117_p),
    .doutn(ffc_117_n),
    .din(G34_p_spl_)
  );


  DROC
  ffc_118
  (
    .doutp(ffc_118_p),
    .doutn(ffc_118_n),
    .din(G24_p)
  );


  DROC
  ffc_119
  (
    .doutp(ffc_119_p),
    .doutn(ffc_119_n),
    .din(G26_p)
  );


  DROC
  ffc_120
  (
    .doutp(ffc_120_p),
    .doutn(ffc_120_n),
    .din(G1_p)
  );


  DROC
  ffc_121
  (
    .doutp(ffc_121_p),
    .doutn(ffc_121_n),
    .din(G2_p)
  );


  DROC
  ffc_122
  (
    .doutp(ffc_122_p),
    .doutn(ffc_122_n),
    .din(G16_p)
  );


  DROC
  ffc_123
  (
    .doutp(ffc_123_p),
    .doutn(ffc_123_n),
    .din(G18_p)
  );


  DROC
  ffc_124
  (
    .doutp(ffc_124_p),
    .doutn(ffc_124_n),
    .din(G20_p)
  );


  DROC
  ffc_125
  (
    .doutp(ffc_125_p),
    .doutn(ffc_125_n),
    .din(G22_p)
  );


  DROC
  ffc_126
  (
    .doutp(ffc_126_p),
    .doutn(ffc_126_n),
    .din(G28_p)
  );


  DROC
  ffc_127
  (
    .doutp(ffc_127_p),
    .doutn(ffc_127_n),
    .din(G30_p)
  );


  DROC
  ffc_128
  (
    .doutp(ffc_128_p),
    .doutn(ffc_128_n),
    .din(g292_p)
  );


  DROC
  ffc_129
  (
    .doutp(ffc_129_p),
    .doutn(ffc_129_n),
    .din(g293_p)
  );


  DROC
  ffc_130
  (
    .doutp(ffc_130_p),
    .doutn(ffc_130_n),
    .din(g294_p)
  );


  DROC
  ffc_131
  (
    .doutp(ffc_131_p),
    .doutn(ffc_131_n),
    .din(g295_p)
  );


  buf

  (
    ffc_87_n_spl_,
    ffc_87_n
  );


  buf

  (
    ffc_87_n_spl_0,
    ffc_87_n_spl_
  );


  buf

  (
    ffc_87_n_spl_00,
    ffc_87_n_spl_0
  );


  buf

  (
    ffc_87_n_spl_1,
    ffc_87_n_spl_
  );


  buf

  (
    ffc_87_p_spl_,
    ffc_87_p
  );


  buf

  (
    ffc_87_p_spl_0,
    ffc_87_p_spl_
  );


  buf

  (
    ffc_87_p_spl_00,
    ffc_87_p_spl_0
  );


  buf

  (
    ffc_87_p_spl_01,
    ffc_87_p_spl_0
  );


  buf

  (
    ffc_87_p_spl_1,
    ffc_87_p_spl_
  );


  buf

  (
    ffc_87_p_spl_10,
    ffc_87_p_spl_1
  );


  buf

  (
    ffc_87_p_spl_11,
    ffc_87_p_spl_1
  );


  buf

  (
    g175_n_spl_,
    g175_n
  );


  buf

  (
    g177_n_spl_,
    g177_n
  );


  buf

  (
    g180_n_spl_,
    g180_n
  );


  buf

  (
    g186_n_spl_,
    g186_n
  );


  buf

  (
    g186_p_spl_,
    g186_p
  );


  buf

  (
    g188_p_spl_,
    g188_p
  );


  buf

  (
    g191_n_spl_,
    g191_n
  );


  buf

  (
    g193_n_spl_,
    g193_n
  );


  buf

  (
    g195_p_spl_,
    g195_p
  );


  buf

  (
    g193_p_spl_,
    g193_p
  );


  buf

  (
    g200_p_spl_,
    g200_p
  );


  buf

  (
    ffc_88_p_spl_,
    ffc_88_p
  );


  buf

  (
    ffc_88_p_spl_0,
    ffc_88_p_spl_
  );


  buf

  (
    ffc_88_p_spl_00,
    ffc_88_p_spl_0
  );


  buf

  (
    ffc_88_p_spl_1,
    ffc_88_p_spl_
  );


  buf

  (
    ffc_34_p_spl_,
    ffc_34_p
  );


  buf

  (
    g222_n_spl_,
    g222_n
  );


  buf

  (
    ffc_39_p_spl_,
    ffc_39_p
  );


  buf

  (
    g220_n_spl_,
    g220_n
  );


  buf

  (
    ffc_8_p_spl_,
    ffc_8_p
  );


  buf

  (
    g214_n_spl_,
    g214_n
  );


  buf

  (
    ffc_23_p_spl_,
    ffc_23_p
  );


  buf

  (
    g216_n_spl_,
    g216_n
  );


  buf

  (
    ffc_28_p_spl_,
    ffc_28_p
  );


  buf

  (
    g218_n_spl_,
    g218_n
  );


  buf

  (
    ffc_3_p_spl_,
    ffc_3_p
  );


  buf

  (
    g209_n_spl_,
    g209_n
  );


  buf

  (
    ffc_44_p_spl_,
    ffc_44_p
  );


  buf

  (
    g212_n_spl_,
    g212_n
  );


  buf

  (
    ffc_18_p_spl_,
    ffc_18_p
  );


  buf

  (
    g211_n_spl_,
    g211_n
  );


  buf

  (
    ffc_13_p_spl_,
    ffc_13_p
  );


  buf

  (
    g210_n_spl_,
    g210_n
  );


  buf

  (
    ffc_31_p_spl_,
    ffc_31_p
  );


  buf

  (
    g228_n_spl_,
    g228_n
  );


  buf

  (
    ffc_97_p_spl_,
    ffc_97_p
  );


  buf

  (
    g226_n_spl_,
    g226_n
  );


  buf

  (
    ffc_94_p_spl_,
    ffc_94_p
  );


  buf

  (
    g223_n_spl_,
    g223_n
  );


  buf

  (
    ffc_95_p_spl_,
    ffc_95_p
  );


  buf

  (
    g224_n_spl_,
    g224_n
  );


  buf

  (
    ffc_96_p_spl_,
    ffc_96_p
  );


  buf

  (
    g225_n_spl_,
    g225_n
  );


  buf

  (
    ffc_119_p_spl_,
    ffc_119_p
  );


  buf

  (
    ffc_127_p_spl_,
    ffc_127_p
  );


  buf

  (
    ffc_123_p_spl_,
    ffc_123_p
  );


  buf

  (
    ffc_125_p_spl_,
    ffc_125_p
  );


  buf

  (
    g233_p_spl_,
    g233_p
  );


  buf

  (
    g244_p_spl_,
    g244_p
  );


  buf

  (
    g249_p_spl_,
    g249_p
  );


  buf

  (
    g260_p_spl_,
    g260_p
  );


  buf

  (
    g265_n_spl_,
    g265_n
  );


  buf

  (
    g272_n_spl_,
    g272_n
  );


  buf

  (
    g274_p_spl_,
    g274_p
  );


  buf

  (
    g274_p_spl_0,
    g274_p_spl_
  );


  buf

  (
    g274_p_spl_00,
    g274_p_spl_0
  );


  buf

  (
    g274_p_spl_1,
    g274_p_spl_
  );


  buf

  (
    g275_n_spl_,
    g275_n
  );


  buf

  (
    g275_n_spl_0,
    g275_n_spl_
  );


  buf

  (
    g275_n_spl_00,
    g275_n_spl_0
  );


  buf

  (
    g275_n_spl_000,
    g275_n_spl_00
  );


  buf

  (
    g275_n_spl_01,
    g275_n_spl_0
  );


  buf

  (
    g275_n_spl_1,
    g275_n_spl_
  );


  buf

  (
    g275_n_spl_10,
    g275_n_spl_1
  );


  buf

  (
    g275_n_spl_11,
    g275_n_spl_1
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G10_p_spl_,
    G10_p
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G34_p_spl_,
    G34_p
  );


endmodule
