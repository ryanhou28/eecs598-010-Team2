// Benchmark "c880" written by ABC on Sun Oct 29 19:31:49 2023

module c880 (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58,
    G59, G60,
    G855, G856, G857, G858, G859, G860, G861, G862, G863, G864, G865, G866,
    G867, G868, G869, G870, G871, G872, G873, G874, G875, G876, G877, G878,
    G879, G880  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G58, G59, G60;
  output G855, G856, G857, G858, G859, G860, G861, G862, G863, G864, G865,
    G866, G867, G868, G869, G870, G871, G872, G873, G874, G875, G876, G877,
    G878, G879, G880;
  reg n471_lo, n474_lo, n477_lo, n480_lo, n483_lo, n486_lo, n489_lo,
    n492_lo, n495_lo, n498_lo, n501_lo, n504_lo, n507_lo, n510_lo, n513_lo,
    n516_lo, n519_lo, n522_lo, n525_lo, n528_lo, n531_lo, n534_lo, n537_lo,
    n540_lo, n543_lo, n546_lo, n549_lo, n552_lo, n555_lo, n558_lo, n561_lo,
    n564_lo, n567_lo, n570_lo, n573_lo, n576_lo, n579_lo, n582_lo, n585_lo,
    n588_lo, n591_lo, n594_lo, n597_lo, n600_lo, n603_lo, n606_lo, n609_lo,
    n612_lo, n615_lo, n618_lo, n621_lo, n624_lo, n627_lo, n630_lo, n633_lo,
    n636_lo, n639_lo, n642_lo, n645_lo, n648_lo, n651_lo, n654_lo, n657_lo,
    n660_lo, n663_lo, n666_lo, n669_lo, n672_lo, n675_lo, n678_lo, n681_lo,
    n684_lo, n687_lo, n690_lo, n693_lo, n696_lo, n699_lo, n702_lo, n705_lo,
    n708_lo, n711_lo, n714_lo, n717_lo, n720_lo, n723_lo, n726_lo, n729_lo,
    n732_lo, n735_lo, n738_lo, n741_lo, n744_lo, n747_lo, n750_lo, n753_lo,
    n756_lo, n759_lo, n762_lo, n765_lo, n768_lo, n771_lo, n774_lo, n777_lo,
    n780_lo, n783_lo, n786_lo, n789_lo, n792_lo, n795_lo, n798_lo, n801_lo,
    n804_lo, n807_lo, n810_lo, n813_lo, n816_lo, n819_lo, n822_lo, n825_lo,
    n828_lo, n831_lo, n834_lo, n837_lo, n840_lo, n843_lo, n846_lo, n849_lo,
    n852_lo, n855_lo, n858_lo, n861_lo, n864_lo, n867_lo, n870_lo, n873_lo,
    n876_lo, n879_lo, n882_lo, n885_lo, n888_lo, n891_lo, n894_lo, n897_lo,
    n900_lo, n903_lo, n906_lo, n909_lo, n912_lo, n915_lo, n918_lo, n921_lo,
    n924_lo, n927_lo, n930_lo, n933_lo, n936_lo, n939_lo, n942_lo, n945_lo,
    n948_lo, n951_lo, n954_lo, n957_lo, n960_lo, n963_lo, n966_lo, n969_lo,
    n972_lo, n975_lo, n978_lo, n981_lo, n984_lo, n987_lo, n990_lo, n993_lo,
    n996_lo, n999_lo, n1002_lo, n1005_lo, n1008_lo, n1011_lo, n1014_lo,
    n1017_lo, n1020_lo, n1023_lo, n1026_lo, n1029_lo, n1032_lo, n1035_lo,
    n1038_lo, n1041_lo, n1044_lo, n1047_lo, n1050_lo, n1053_lo, n1056_lo,
    n1059_lo, n1062_lo, n1065_lo, n1068_lo, n1071_lo, n1074_lo, n1077_lo,
    n1080_lo, n1083_lo, n1086_lo, n1089_lo, n1092_lo, n1095_lo, n1098_lo,
    n1101_lo, n1104_lo, n1107_lo, n1110_lo, n1113_lo, n1116_lo, n1119_lo,
    n1122_lo, n1125_lo, n1128_lo, n1131_lo, n1134_lo, n1137_lo, n1140_lo,
    n1143_lo, n1146_lo, n1149_lo, n1152_lo, n1155_lo, n1158_lo, n1161_lo,
    n1164_lo, n1167_lo, n1170_lo, n1173_lo, n1176_lo, n1179_lo, n1182_lo,
    n1185_lo, n1188_lo;
  wire new_G269_, new_G270_, new_G273_, new_G276_, new_G279_, new_G280_,
    new_G284_, new_G285_, new_G286_, new_G287_, new_G290_, new_G291_,
    new_G292_, new_G293_, new_G294_, new_G295_, new_G296_, new_G297_,
    new_G298_, new_G301_, new_G302_, new_G303_, new_G304_, new_G305_,
    new_G306_, new_G307_, new_G308_, new_G309_, new_G310_, new_G316_,
    new_G317_, new_G318_, new_G319_, new_G322_, new_G323_, new_G324_,
    new_G325_, new_G326_, new_G327_, new_G328_, new_G329_, new_G330_,
    new_G331_, new_G332_, new_G333_, new_G334_, new_G335_, new_G336_,
    new_G337_, new_G338_, new_G339_, new_G340_, new_G341_, new_G342_,
    new_G343_, new_G344_, new_G345_, new_G346_, new_G347_, new_G348_,
    new_G349_, new_G350_, new_G351_, new_G352_, new_G353_, new_G354_,
    new_G355_, new_G356_, new_G357_, new_G360_, new_G363_, new_G366_,
    new_G369_, new_G375_, new_G376_, new_G379_, new_G382_, new_G385_,
    new_G388_, new_G389_, new_G395_, new_G396_, new_G397_, new_G398_,
    new_G399_, new_G400_, new_G401_, new_G402_, new_G403_, new_G404_,
    new_G405_, new_G406_, new_G407_, new_G408_, new_G409_, new_G410_,
    new_G411_, new_G412_, new_G413_, new_G414_, new_G415_, new_G416_,
    new_G417_, new_G422_, new_G427_, new_G432_, new_G433_, new_G434_,
    new_G435_, new_G436_, new_G445_, new_G448_, new_G451_, new_G460_,
    new_G461_, new_G462_, new_G463_, new_G464_, new_G465_, new_G466_,
    new_G467_, new_G468_, new_G473_, new_G474_, new_G475_, new_G476_,
    new_G477_, new_G480_, new_G483_, new_G484_, new_G485_, new_G486_,
    new_G487_, new_G488_, new_G489_, new_G490_, new_G491_, new_G492_,
    new_G493_, new_G494_, new_G495_, new_G496_, new_G497_, new_G498_,
    new_G499_, new_G500_, new_G501_, new_G502_, new_G503_, new_G504_,
    new_G505_, new_G506_, new_G507_, new_G508_, new_G509_, new_G510_,
    new_G511_, new_G512_, new_G513_, new_G514_, new_G515_, new_G518_,
    new_G521_, new_G522_, new_G523_, new_G524_, new_G525_, new_G526_,
    new_G527_, new_G528_, new_G529_, new_G532_, new_G535_, new_G536_,
    new_G537_, new_G538_, new_G542_, new_G546_, new_G550_, new_G554_,
    new_G558_, new_G562_, new_G566_, new_G570_, new_G571_, new_G572_,
    new_G573_, new_G574_, new_G575_, new_G578_, new_G581_, new_G582_,
    new_G585_, new_G590_, new_G591_, new_G594_, new_G600_, new_G601_,
    new_G604_, new_G609_, new_G610_, new_G613_, new_G616_, new_G617_,
    new_G620_, new_G625_, new_G626_, new_G629_, new_G635_, new_G636_,
    new_G639_, new_G644_, new_G645_, new_G646_, new_G647_, new_G650_,
    new_G654_, new_G655_, new_G658_, new_G662_, new_G663_, new_G667_,
    new_G671_, new_G672_, new_G677_, new_G681_, new_G682_, new_G685_,
    new_G689_, new_G690_, new_G693_, new_G697_, new_G698_, new_G702_,
    new_G706_, new_G707_, new_G712_, new_G716_, new_G717_, new_G718_,
    new_G719_, new_G720_, new_G721_, new_G722_, new_G723_, new_G724_,
    new_G725_, new_G726_, new_G727_, new_G728_, new_G729_, new_G730_,
    new_G731_, new_G732_, new_G733_, new_G734_, new_G735_, new_G736_,
    new_G737_, new_G738_, new_G739_, new_G740_, new_G741_, new_G742_,
    new_G743_, new_G744_, new_G745_, new_G746_, new_G747_, new_G748_,
    new_G749_, new_G750_, new_G751_, new_G752_, new_G753_, new_G754_,
    new_G755_, new_G756_, new_G760_, new_G761_, new_G764_, new_G765_,
    new_G768_, new_G769_, new_G770_, new_G771_, new_G772_, new_G773_,
    new_G774_, new_G775_, new_G776_, new_G777_, new_G778_, new_G779_,
    new_G785_, new_G786_, new_G787_, new_G788_, new_G789_, new_G790_,
    new_G791_, new_G792_, new_G793_, new_G794_, new_G795_, new_G796_,
    new_G797_, new_G798_, new_G802_, new_G805_, new_G808_, new_G809_,
    new_G810_, new_G811_, new_G812_, new_G813_, new_G814_, new_G815_,
    new_G816_, new_G817_, new_G818_, new_G819_, new_G820_, new_G821_,
    new_G822_, new_G823_, new_G824_, new_G825_, new_G826_, new_G827_,
    new_G828_, new_G829_, new_G830_, new_G831_, new_G832_, new_G833_,
    new_G834_, new_G835_, new_G836_, new_G837_, new_G838_, new_G839_,
    new_G840_, new_G841_, new_G842_, new_G843_, new_G844_, new_G845_,
    new_G846_, new_G847_, new_G848_, new_G849_, new_G850_, new_G851_,
    new_G852_, new_G853_, new_G854_, n471_li, n474_li, n477_li, n480_li,
    n483_li, n486_li, n489_li, n492_li, n495_li, n498_li, n501_li, n504_li,
    n507_li, n510_li, n513_li, n516_li, n519_li, n522_li, n525_li, n528_li,
    n531_li, n534_li, n537_li, n540_li, n543_li, n546_li, n549_li, n552_li,
    n555_li, n558_li, n561_li, n564_li, n567_li, n570_li, n573_li, n576_li,
    n579_li, n582_li, n585_li, n588_li, n591_li, n594_li, n597_li, n600_li,
    n603_li, n606_li, n609_li, n612_li, n615_li, n618_li, n621_li, n624_li,
    n627_li, n630_li, n633_li, n636_li, n639_li, n642_li, n645_li, n648_li,
    n651_li, n654_li, n657_li, n660_li, n663_li, n666_li, n669_li, n672_li,
    n675_li, n678_li, n681_li, n684_li, n687_li, n690_li, n693_li, n696_li,
    n699_li, n702_li, n705_li, n708_li, n711_li, n714_li, n717_li, n720_li,
    n723_li, n726_li, n729_li, n732_li, n735_li, n738_li, n741_li, n744_li,
    n747_li, n750_li, n753_li, n756_li, n759_li, n762_li, n765_li, n768_li,
    n771_li, n774_li, n777_li, n780_li, n783_li, n786_li, n789_li, n792_li,
    n795_li, n798_li, n801_li, n804_li, n807_li, n810_li, n813_li, n816_li,
    n819_li, n822_li, n825_li, n828_li, n831_li, n834_li, n837_li, n840_li,
    n843_li, n846_li, n849_li, n852_li, n855_li, n858_li, n861_li, n864_li,
    n867_li, n870_li, n873_li, n876_li, n879_li, n882_li, n885_li, n888_li,
    n891_li, n894_li, n897_li, n900_li, n903_li, n906_li, n909_li, n912_li,
    n915_li, n918_li, n921_li, n924_li, n927_li, n930_li, n933_li, n936_li,
    n939_li, n942_li, n945_li, n948_li, n951_li, n954_li, n957_li, n960_li,
    n963_li, n966_li, n969_li, n972_li, n975_li, n978_li, n981_li, n984_li,
    n987_li, n990_li, n993_li, n996_li, n999_li, n1002_li, n1005_li,
    n1008_li, n1011_li, n1014_li, n1017_li, n1020_li, n1023_li, n1026_li,
    n1029_li, n1032_li, n1035_li, n1038_li, n1041_li, n1044_li, n1047_li,
    n1050_li, n1053_li, n1056_li, n1059_li, n1062_li, n1065_li, n1068_li,
    n1071_li, n1074_li, n1077_li, n1080_li, n1083_li, n1086_li, n1089_li,
    n1092_li, n1095_li, n1098_li, n1101_li, n1104_li, n1107_li, n1110_li,
    n1113_li, n1116_li, n1119_li, n1122_li, n1125_li, n1128_li, n1131_li,
    n1134_li, n1137_li, n1140_li, n1143_li, n1146_li, n1149_li, n1152_li,
    n1155_li, n1158_li, n1161_li, n1164_li, n1167_li, n1170_li, n1173_li,
    n1176_li, n1179_li, n1182_li, n1185_li, n1188_li;
  assign new_G269_ = ~n516_lo | ~n504_lo | ~n480_lo | ~n492_lo;
  assign new_G270_ = ~n516_lo | ~n504_lo | ~n480_lo | ~n528_lo;
  assign new_G273_ = n564_lo & n540_lo & n552_lo;
  assign new_G276_ = n576_lo & n480_lo & n528_lo;
  assign new_G279_ = ~n516_lo | ~n576_lo | ~n480_lo | ~n492_lo;
  assign new_G280_ = ~n588_lo | ~n504_lo | ~n480_lo | ~n492_lo;
  assign new_G284_ = ~n624_lo | ~n612_lo | ~n600_lo | ~n564_lo;
  assign new_G285_ = ~n540_lo | ~n612_lo;
  assign new_G286_ = ~n648_lo | ~n600_lo | ~n612_lo;
  assign new_G287_ = n672_lo & n540_lo & n660_lo;
  assign new_G290_ = n564_lo & n540_lo & n660_lo;
  assign new_G291_ = n672_lo & n540_lo & n552_lo;
  assign new_G292_ = n564_lo & n540_lo & n552_lo;
  assign new_G293_ = n672_lo & n600_lo & n660_lo;
  assign new_G294_ = n564_lo & n600_lo & n660_lo;
  assign new_G295_ = n672_lo & n600_lo & n552_lo;
  assign new_G296_ = n564_lo & n600_lo & n552_lo;
  assign new_G297_ = n684_lo & n696_lo;
  assign new_G298_ = n708_lo | n720_lo;
  assign new_G301_ = ~n756_lo | ~n768_lo;
  assign new_G302_ = n756_lo | n768_lo;
  assign new_G303_ = ~n780_lo | ~n792_lo;
  assign new_G304_ = n780_lo | n792_lo;
  assign new_G305_ = ~n804_lo | ~n816_lo;
  assign new_G306_ = n804_lo | n816_lo;
  assign new_G307_ = ~n828_lo | ~n840_lo;
  assign new_G308_ = n828_lo | n840_lo;
  assign new_G309_ = n492_lo & n876_lo;
  assign new_G310_ = ~n1188_lo;
  assign new_G316_ = n576_lo & n876_lo;
  assign new_G317_ = n516_lo & n876_lo;
  assign new_G318_ = n924_lo & n876_lo;
  assign new_G319_ = ~n600_lo | ~n948_lo;
  assign new_G322_ = ~n516_lo & ~n564_lo;
  assign new_G323_ = n516_lo & n564_lo;
  assign new_G324_ = ~n960_lo | ~n972_lo;
  assign new_G325_ = n960_lo | n972_lo;
  assign new_G326_ = ~n984_lo | ~n996_lo;
  assign new_G327_ = n984_lo | n996_lo;
  assign new_G328_ = ~n1008_lo | ~n1020_lo;
  assign new_G329_ = n1008_lo | n1020_lo;
  assign new_G330_ = ~n1032_lo | ~n1044_lo;
  assign new_G331_ = n1032_lo | n1044_lo;
  assign new_G332_ = n1068_lo & n756_lo;
  assign new_G333_ = n1068_lo & n768_lo;
  assign new_G334_ = n1068_lo & n780_lo;
  assign new_G335_ = n1068_lo & n792_lo;
  assign new_G336_ = n1068_lo & n804_lo;
  assign new_G337_ = n1128_lo & n1140_lo;
  assign new_G338_ = n1068_lo & n816_lo;
  assign new_G339_ = n1128_lo & n1152_lo;
  assign new_G340_ = n1068_lo & n828_lo;
  assign new_G341_ = n1128_lo & n1176_lo;
  assign new_G342_ = ~new_G269_;
  assign new_G343_ = ~new_G273_;
  assign new_G344_ = new_G270_ | new_G273_;
  assign new_G345_ = ~new_G276_;
  assign new_G346_ = ~new_G276_;
  assign new_G347_ = ~new_G279_;
  assign new_G348_ = ~new_G280_ & ~new_G284_;
  assign new_G349_ = new_G280_ | new_G285_;
  assign new_G350_ = new_G280_ | new_G286_;
  assign new_G351_ = ~new_G293_;
  assign new_G352_ = ~new_G294_;
  assign new_G353_ = ~new_G295_;
  assign new_G354_ = ~new_G296_;
  assign new_G355_ = ~n732_lo | ~new_G298_;
  assign new_G356_ = n744_lo & new_G298_;
  assign new_G357_ = ~new_G301_ | ~new_G302_;
  assign new_G360_ = ~new_G303_ | ~new_G304_;
  assign new_G363_ = ~new_G305_ | ~new_G306_;
  assign new_G366_ = ~new_G307_ | ~new_G308_;
  assign new_G369_ = ~new_G310_;
  assign new_G375_ = ~new_G322_ & ~new_G323_;
  assign new_G376_ = ~new_G324_ | ~new_G325_;
  assign new_G379_ = ~new_G326_ | ~new_G327_;
  assign new_G382_ = ~new_G328_ | ~new_G329_;
  assign new_G385_ = ~new_G330_ | ~new_G331_;
  assign new_G388_ = new_G270_ | new_G343_;
  assign new_G389_ = ~new_G345_;
  assign new_G395_ = ~new_G346_;
  assign new_G396_ = new_G348_ & n636_lo;
  assign new_G397_ = ~new_G349_;
  assign new_G398_ = ~new_G350_;
  assign new_G399_ = ~new_G355_;
  assign new_G400_ = ~new_G357_;
  assign new_G401_ = ~new_G360_;
  assign new_G402_ = new_G357_ & new_G360_;
  assign new_G403_ = ~new_G363_;
  assign new_G404_ = ~new_G366_;
  assign new_G405_ = new_G363_ & new_G366_;
  assign new_G406_ = ~new_G347_ | ~new_G352_;
  assign new_G407_ = ~new_G376_;
  assign new_G408_ = ~new_G379_;
  assign new_G409_ = new_G376_ & new_G379_;
  assign new_G410_ = ~new_G382_;
  assign new_G411_ = ~new_G385_;
  assign new_G412_ = new_G382_ & new_G385_;
  assign new_G413_ = n1068_lo & new_G369_;
  assign new_G414_ = ~new_G396_;
  assign new_G415_ = new_G400_ & new_G401_;
  assign new_G416_ = new_G403_ & new_G404_;
  assign new_G417_ = n588_lo & new_G319_ & new_G389_;
  assign new_G422_ = new_G287_ & new_G389_ & n516_lo;
  assign new_G427_ = ~n588_lo | ~new_G389_ | ~new_G287_;
  assign new_G432_ = ~new_G389_ | ~n948_lo | ~new_G375_ | ~n600_lo;
  assign new_G433_ = ~n516_lo | ~new_G389_ | ~new_G319_;
  assign new_G434_ = new_G407_ & new_G408_;
  assign new_G435_ = new_G410_ & new_G411_;
  assign new_G436_ = ~new_G414_;
  assign new_G445_ = ~new_G402_ & ~new_G415_;
  assign new_G448_ = ~new_G405_ & ~new_G416_;
  assign new_G451_ = ~new_G432_ | ~new_G406_;
  assign new_G460_ = n888_lo & new_G417_;
  assign new_G461_ = new_G310_ & new_G422_;
  assign new_G462_ = n900_lo & new_G417_;
  assign new_G463_ = new_G310_ & new_G422_;
  assign new_G464_ = n912_lo & new_G417_;
  assign new_G465_ = new_G310_ & new_G422_;
  assign new_G466_ = n936_lo & new_G417_;
  assign new_G467_ = new_G310_ & new_G422_;
  assign new_G468_ = ~new_G433_ | ~n480_lo;
  assign new_G473_ = new_G369_ | new_G427_;
  assign new_G474_ = new_G369_ | new_G427_;
  assign new_G475_ = new_G369_ | new_G427_;
  assign new_G476_ = new_G369_ | new_G427_;
  assign new_G477_ = ~new_G409_ & ~new_G434_;
  assign new_G480_ = ~new_G412_ & ~new_G435_;
  assign new_G483_ = ~n852_lo | ~new_G445_;
  assign new_G484_ = n852_lo | new_G445_;
  assign new_G485_ = ~new_G448_ | ~n864_lo;
  assign new_G486_ = new_G448_ | n864_lo;
  assign new_G487_ = n756_lo & new_G451_;
  assign new_G488_ = ~new_G460_ & ~new_G461_;
  assign new_G489_ = n768_lo & new_G451_;
  assign new_G490_ = ~new_G462_ & ~new_G463_;
  assign new_G491_ = n780_lo & new_G451_;
  assign new_G492_ = ~new_G464_ & ~new_G465_;
  assign new_G493_ = n792_lo & new_G451_;
  assign new_G494_ = ~new_G466_ & ~new_G467_;
  assign new_G495_ = n888_lo & new_G468_;
  assign new_G496_ = n804_lo & new_G451_;
  assign new_G497_ = n900_lo & new_G468_;
  assign new_G498_ = n816_lo & new_G451_;
  assign new_G499_ = n912_lo & new_G468_;
  assign new_G500_ = n828_lo & new_G451_;
  assign new_G501_ = n936_lo & new_G468_;
  assign new_G502_ = n840_lo & new_G451_;
  assign new_G503_ = ~n852_lo | ~new_G477_;
  assign new_G504_ = n852_lo | new_G477_;
  assign new_G505_ = ~new_G480_ | ~n1056_lo;
  assign new_G506_ = new_G480_ | n1056_lo;
  assign new_G507_ = new_G436_ & n960_lo;
  assign new_G508_ = new_G436_ & n972_lo;
  assign new_G509_ = new_G436_ & n984_lo;
  assign new_G510_ = new_G436_ & n996_lo;
  assign new_G511_ = new_G436_ & n1008_lo;
  assign new_G512_ = ~new_G436_ | ~n1020_lo;
  assign new_G513_ = ~new_G436_ | ~n1032_lo;
  assign new_G514_ = ~new_G436_ | ~n1044_lo;
  assign new_G515_ = ~new_G483_ | ~new_G484_;
  assign new_G518_ = ~new_G485_ | ~new_G486_;
  assign new_G521_ = ~new_G309_ & ~new_G487_;
  assign new_G522_ = ~new_G316_ & ~new_G489_;
  assign new_G523_ = ~new_G317_ & ~new_G491_;
  assign new_G524_ = ~new_G318_ & ~new_G493_;
  assign new_G525_ = ~new_G495_ & ~new_G496_;
  assign new_G526_ = ~new_G497_ & ~new_G498_;
  assign new_G527_ = ~new_G499_ & ~new_G500_;
  assign new_G528_ = ~new_G501_ & ~new_G502_;
  assign new_G529_ = ~new_G503_ | ~new_G504_;
  assign new_G532_ = ~new_G505_ | ~new_G506_;
  assign new_G535_ = ~new_G515_;
  assign new_G536_ = ~new_G518_;
  assign new_G537_ = new_G515_ & new_G518_;
  assign new_G538_ = ~new_G521_ | ~new_G488_;
  assign new_G542_ = ~new_G522_ | ~new_G490_;
  assign new_G546_ = ~new_G523_ | ~new_G492_;
  assign new_G550_ = ~new_G524_ | ~new_G494_;
  assign new_G554_ = ~new_G473_ | ~new_G525_;
  assign new_G558_ = ~new_G474_ | ~new_G526_;
  assign new_G562_ = ~new_G475_ | ~new_G527_;
  assign new_G566_ = ~new_G476_ | ~new_G528_;
  assign new_G570_ = ~new_G529_;
  assign new_G571_ = ~new_G532_;
  assign new_G572_ = new_G529_ & new_G532_;
  assign new_G573_ = new_G535_ & new_G536_;
  assign new_G574_ = new_G570_ & new_G571_;
  assign new_G575_ = ~new_G538_ | ~n960_lo;
  assign new_G578_ = new_G538_ | n960_lo;
  assign new_G581_ = n1116_lo & new_G538_;
  assign new_G582_ = ~new_G542_ | ~n972_lo;
  assign new_G585_ = new_G542_ | n972_lo;
  assign new_G590_ = n1116_lo & new_G542_;
  assign new_G591_ = ~new_G546_ | ~n984_lo;
  assign new_G594_ = new_G546_ | n984_lo;
  assign new_G600_ = n1116_lo & new_G546_;
  assign new_G601_ = ~new_G550_ | ~n996_lo;
  assign new_G604_ = new_G550_ | n996_lo;
  assign new_G609_ = n1116_lo & new_G550_;
  assign new_G610_ = ~new_G554_ | ~n1008_lo;
  assign new_G613_ = new_G554_ | n1008_lo;
  assign new_G616_ = n1116_lo & new_G554_;
  assign new_G617_ = ~new_G558_ | ~n1020_lo;
  assign new_G620_ = new_G558_ | n1020_lo;
  assign new_G625_ = n1116_lo & new_G558_;
  assign new_G626_ = ~new_G562_ | ~n1032_lo;
  assign new_G629_ = new_G562_ | n1032_lo;
  assign new_G635_ = n1116_lo & new_G562_;
  assign new_G636_ = ~new_G566_ | ~n1044_lo;
  assign new_G639_ = new_G566_ | n1044_lo;
  assign new_G644_ = n1116_lo & new_G566_;
  assign new_G645_ = ~new_G537_ & ~new_G573_;
  assign new_G646_ = ~new_G572_ & ~new_G574_;
  assign new_G647_ = ~new_G575_;
  assign new_G650_ = new_G578_ & new_G575_;
  assign new_G654_ = ~new_G581_ & ~new_G507_;
  assign new_G655_ = ~new_G582_;
  assign new_G658_ = new_G585_ & new_G582_;
  assign new_G662_ = ~new_G590_ & ~new_G508_;
  assign new_G663_ = ~new_G591_;
  assign new_G667_ = new_G594_ & new_G591_;
  assign new_G671_ = ~new_G600_ & ~new_G509_;
  assign new_G672_ = ~new_G601_;
  assign new_G677_ = new_G604_ & new_G601_;
  assign new_G681_ = ~new_G609_ & ~new_G510_;
  assign new_G682_ = ~new_G610_;
  assign new_G685_ = new_G613_ & new_G610_;
  assign new_G689_ = ~new_G616_ & ~new_G511_;
  assign new_G690_ = ~new_G617_;
  assign new_G693_ = new_G620_ & new_G617_;
  assign new_G697_ = ~new_G337_ & ~new_G625_;
  assign new_G698_ = ~new_G626_;
  assign new_G702_ = new_G629_ & new_G626_;
  assign new_G706_ = ~new_G339_ & ~new_G635_;
  assign new_G707_ = ~new_G636_;
  assign new_G712_ = new_G639_ & new_G636_;
  assign new_G716_ = ~new_G341_ & ~new_G644_;
  assign new_G717_ = ~new_G639_ | ~n1164_lo;
  assign new_G718_ = ~n1164_lo | ~new_G629_ | ~new_G639_;
  assign new_G719_ = ~n1164_lo | ~new_G639_ | ~new_G620_ | ~new_G629_;
  assign new_G720_ = ~new_G647_;
  assign new_G721_ = n1092_lo & new_G650_;
  assign new_G722_ = n1104_lo & new_G647_;
  assign new_G723_ = ~new_G655_;
  assign new_G724_ = n1092_lo & new_G658_;
  assign new_G725_ = n1104_lo & new_G655_;
  assign new_G726_ = ~new_G663_;
  assign new_G727_ = n1092_lo & new_G667_;
  assign new_G728_ = n1104_lo & new_G663_;
  assign new_G729_ = ~new_G672_;
  assign new_G730_ = n1092_lo & new_G677_;
  assign new_G731_ = n1104_lo & new_G672_;
  assign new_G732_ = ~new_G682_;
  assign new_G733_ = n1092_lo & new_G685_;
  assign new_G734_ = n1104_lo & new_G682_;
  assign new_G735_ = ~new_G690_;
  assign new_G736_ = n1092_lo & new_G693_;
  assign new_G737_ = n1104_lo & new_G690_;
  assign new_G738_ = ~new_G698_;
  assign new_G739_ = n1092_lo & new_G702_;
  assign new_G740_ = n1104_lo & new_G698_;
  assign new_G741_ = ~new_G707_;
  assign new_G742_ = ~new_G712_ & ~n1164_lo;
  assign new_G743_ = new_G712_ & n1164_lo;
  assign new_G744_ = n1092_lo & new_G712_;
  assign new_G745_ = n1104_lo & new_G707_;
  assign new_G746_ = ~new_G629_ | ~new_G707_;
  assign new_G747_ = ~new_G620_ | ~new_G698_;
  assign new_G748_ = ~new_G707_ | ~new_G620_ | ~new_G629_;
  assign new_G749_ = ~new_G594_ | ~new_G672_;
  assign new_G750_ = ~new_G585_ | ~new_G663_;
  assign new_G751_ = ~new_G672_ | ~new_G585_ | ~new_G594_;
  assign new_G752_ = ~new_G721_ & ~new_G722_;
  assign new_G753_ = ~new_G724_ & ~new_G725_;
  assign new_G754_ = ~new_G727_ & ~new_G728_;
  assign new_G755_ = ~new_G730_ & ~new_G731_;
  assign new_G756_ = ~new_G719_ | ~new_G748_ | ~new_G735_ | ~new_G747_;
  assign new_G760_ = ~new_G733_ & ~new_G734_;
  assign new_G761_ = ~new_G718_ | ~new_G738_ | ~new_G746_;
  assign new_G764_ = ~new_G736_ & ~new_G737_;
  assign new_G765_ = ~new_G741_ | ~new_G717_;
  assign new_G768_ = ~new_G739_ & ~new_G740_;
  assign new_G769_ = ~new_G742_ & ~new_G743_;
  assign new_G770_ = ~new_G744_ & ~new_G745_;
  assign new_G771_ = ~new_G685_ & ~new_G756_;
  assign new_G772_ = new_G685_ & new_G756_;
  assign new_G773_ = ~new_G693_ & ~new_G761_;
  assign new_G774_ = new_G693_ & new_G761_;
  assign new_G775_ = ~new_G702_ & ~new_G765_;
  assign new_G776_ = new_G702_ & new_G765_;
  assign new_G777_ = n1080_lo & new_G769_;
  assign new_G778_ = ~new_G613_ | ~new_G756_;
  assign new_G779_ = ~new_G778_ | ~new_G732_;
  assign new_G785_ = ~new_G771_ & ~new_G772_;
  assign new_G786_ = ~new_G773_ & ~new_G774_;
  assign new_G787_ = ~new_G775_ & ~new_G776_;
  assign new_G788_ = ~new_G340_ & ~new_G777_;
  assign new_G789_ = ~new_G677_ & ~new_G779_;
  assign new_G790_ = new_G677_ & new_G779_;
  assign new_G791_ = n1080_lo & new_G785_;
  assign new_G792_ = n1080_lo & new_G786_;
  assign new_G793_ = n1080_lo & new_G787_;
  assign new_G794_ = ~new_G514_ | ~new_G716_ | ~new_G788_ | ~new_G770_;
  assign new_G795_ = ~new_G604_ | ~new_G779_;
  assign new_G796_ = ~new_G779_ | ~new_G594_ | ~new_G604_;
  assign new_G797_ = ~new_G779_ | ~new_G604_ | ~new_G585_ | ~new_G594_;
  assign new_G798_ = ~new_G797_ | ~new_G751_ | ~new_G723_ | ~new_G750_;
  assign new_G802_ = ~new_G796_ | ~new_G726_ | ~new_G749_;
  assign new_G805_ = ~new_G729_ | ~new_G795_;
  assign new_G808_ = ~new_G789_ & ~new_G790_;
  assign new_G809_ = ~new_G335_ & ~new_G791_;
  assign new_G810_ = ~new_G336_ & ~new_G792_;
  assign new_G811_ = ~new_G338_ & ~new_G793_;
  assign new_G812_ = ~new_G794_;
  assign new_G813_ = ~new_G650_ & ~new_G798_;
  assign new_G814_ = new_G650_ & new_G798_;
  assign new_G815_ = ~new_G658_ & ~new_G802_;
  assign new_G816_ = new_G658_ & new_G802_;
  assign new_G817_ = ~new_G667_ & ~new_G805_;
  assign new_G818_ = new_G667_ & new_G805_;
  assign new_G819_ = n1080_lo & new_G808_;
  assign new_G820_ = ~new_G689_ | ~new_G809_ | ~new_G760_;
  assign new_G821_ = ~new_G512_ | ~new_G697_ | ~new_G810_ | ~new_G764_;
  assign new_G822_ = ~new_G513_ | ~new_G706_ | ~new_G811_ | ~new_G768_;
  assign new_G823_ = ~new_G812_;
  assign new_G824_ = ~new_G798_ | ~new_G578_;
  assign new_G825_ = ~new_G813_ & ~new_G814_;
  assign new_G826_ = ~new_G815_ & ~new_G816_;
  assign new_G827_ = ~new_G817_ & ~new_G818_;
  assign new_G828_ = ~new_G334_ & ~new_G819_;
  assign new_G829_ = ~new_G820_;
  assign new_G830_ = ~new_G821_;
  assign new_G831_ = ~new_G822_;
  assign new_G832_ = new_G720_ & new_G824_;
  assign new_G833_ = n1080_lo & new_G825_;
  assign new_G834_ = n1080_lo & new_G826_;
  assign new_G835_ = n1080_lo & new_G827_;
  assign new_G836_ = ~new_G681_ | ~new_G828_ | ~new_G755_;
  assign new_G837_ = ~new_G829_;
  assign new_G838_ = ~new_G830_;
  assign new_G839_ = ~new_G831_;
  assign new_G840_ = ~new_G832_;
  assign new_G841_ = ~new_G413_ & ~new_G833_;
  assign new_G842_ = ~new_G332_ & ~new_G834_;
  assign new_G843_ = ~new_G333_ & ~new_G835_;
  assign new_G844_ = ~new_G836_;
  assign new_G845_ = ~new_G654_ | ~new_G841_ | ~new_G752_;
  assign new_G846_ = ~new_G662_ | ~new_G842_ | ~new_G753_;
  assign new_G847_ = ~new_G671_ | ~new_G843_ | ~new_G754_;
  assign new_G848_ = ~new_G844_;
  assign new_G849_ = ~new_G845_;
  assign new_G850_ = ~new_G846_;
  assign new_G851_ = ~new_G847_;
  assign new_G852_ = ~new_G849_;
  assign new_G853_ = ~new_G850_;
  assign new_G854_ = ~new_G851_;
  assign G855 = ~new_G290_;
  assign G856 = ~new_G291_;
  assign G857 = ~new_G292_;
  assign G858 = ~new_G297_;
  assign G859 = ~new_G342_;
  assign G860 = ~new_G344_;
  assign G861 = ~new_G351_;
  assign G862 = ~new_G353_;
  assign G863 = ~new_G354_;
  assign G864 = ~new_G356_;
  assign G865 = ~new_G388_;
  assign G866 = ~new_G395_;
  assign G867 = ~new_G397_;
  assign G868 = ~new_G398_;
  assign G869 = ~new_G399_;
  assign G870 = ~new_G645_;
  assign G871 = ~new_G646_;
  assign G872 = ~new_G823_;
  assign G873 = ~new_G837_;
  assign G874 = ~new_G838_;
  assign G875 = ~new_G839_;
  assign G876 = ~new_G840_;
  assign G877 = ~new_G848_;
  assign G878 = ~new_G852_;
  assign G879 = ~new_G853_;
  assign G880 = ~new_G854_;
  assign n471_li = G1;
  assign n474_li = n471_lo;
  assign n477_li = n474_lo;
  assign n480_li = n477_lo;
  assign n483_li = G2;
  assign n486_li = n483_lo;
  assign n489_li = n486_lo;
  assign n492_li = n489_lo;
  assign n495_li = G3;
  assign n498_li = n495_lo;
  assign n501_li = n498_lo;
  assign n504_li = n501_lo;
  assign n507_li = G4;
  assign n510_li = n507_lo;
  assign n513_li = n510_lo;
  assign n516_li = n513_lo;
  assign n519_li = G5;
  assign n522_li = n519_lo;
  assign n525_li = n522_lo;
  assign n528_li = n525_lo;
  assign n531_li = G6;
  assign n534_li = n531_lo;
  assign n537_li = n534_lo;
  assign n540_li = n537_lo;
  assign n543_li = G7;
  assign n546_li = n543_lo;
  assign n549_li = n546_lo;
  assign n552_li = n549_lo;
  assign n555_li = G8;
  assign n558_li = n555_lo;
  assign n561_li = n558_lo;
  assign n564_li = n561_lo;
  assign n567_li = G9;
  assign n570_li = n567_lo;
  assign n573_li = n570_lo;
  assign n576_li = n573_lo;
  assign n579_li = G10;
  assign n582_li = n579_lo;
  assign n585_li = n582_lo;
  assign n588_li = n585_lo;
  assign n591_li = G11;
  assign n594_li = n591_lo;
  assign n597_li = n594_lo;
  assign n600_li = n597_lo;
  assign n603_li = G12;
  assign n606_li = n603_lo;
  assign n609_li = n606_lo;
  assign n612_li = n609_lo;
  assign n615_li = G13;
  assign n618_li = n615_lo;
  assign n621_li = n618_lo;
  assign n624_li = n621_lo;
  assign n627_li = G14;
  assign n630_li = n627_lo;
  assign n633_li = n630_lo;
  assign n636_li = n633_lo;
  assign n639_li = G15;
  assign n642_li = n639_lo;
  assign n645_li = n642_lo;
  assign n648_li = n645_lo;
  assign n651_li = G16;
  assign n654_li = n651_lo;
  assign n657_li = n654_lo;
  assign n660_li = n657_lo;
  assign n663_li = G17;
  assign n666_li = n663_lo;
  assign n669_li = n666_lo;
  assign n672_li = n669_lo;
  assign n675_li = G18;
  assign n678_li = n675_lo;
  assign n681_li = n678_lo;
  assign n684_li = n681_lo;
  assign n687_li = G19;
  assign n690_li = n687_lo;
  assign n693_li = n690_lo;
  assign n696_li = n693_lo;
  assign n699_li = G20;
  assign n702_li = n699_lo;
  assign n705_li = n702_lo;
  assign n708_li = n705_lo;
  assign n711_li = G21;
  assign n714_li = n711_lo;
  assign n717_li = n714_lo;
  assign n720_li = n717_lo;
  assign n723_li = G22;
  assign n726_li = n723_lo;
  assign n729_li = n726_lo;
  assign n732_li = n729_lo;
  assign n735_li = G23;
  assign n738_li = n735_lo;
  assign n741_li = n738_lo;
  assign n744_li = n741_lo;
  assign n747_li = G24;
  assign n750_li = n747_lo;
  assign n753_li = n750_lo;
  assign n756_li = n753_lo;
  assign n759_li = G25;
  assign n762_li = n759_lo;
  assign n765_li = n762_lo;
  assign n768_li = n765_lo;
  assign n771_li = G26;
  assign n774_li = n771_lo;
  assign n777_li = n774_lo;
  assign n780_li = n777_lo;
  assign n783_li = G27;
  assign n786_li = n783_lo;
  assign n789_li = n786_lo;
  assign n792_li = n789_lo;
  assign n795_li = G28;
  assign n798_li = n795_lo;
  assign n801_li = n798_lo;
  assign n804_li = n801_lo;
  assign n807_li = G29;
  assign n810_li = n807_lo;
  assign n813_li = n810_lo;
  assign n816_li = n813_lo;
  assign n819_li = G30;
  assign n822_li = n819_lo;
  assign n825_li = n822_lo;
  assign n828_li = n825_lo;
  assign n831_li = G31;
  assign n834_li = n831_lo;
  assign n837_li = n834_lo;
  assign n840_li = n837_lo;
  assign n843_li = G32;
  assign n846_li = n843_lo;
  assign n849_li = n846_lo;
  assign n852_li = n849_lo;
  assign n855_li = G33;
  assign n858_li = n855_lo;
  assign n861_li = n858_lo;
  assign n864_li = n861_lo;
  assign n867_li = G34;
  assign n870_li = n867_lo;
  assign n873_li = n870_lo;
  assign n876_li = n873_lo;
  assign n879_li = G35;
  assign n882_li = n879_lo;
  assign n885_li = n882_lo;
  assign n888_li = n885_lo;
  assign n891_li = G36;
  assign n894_li = n891_lo;
  assign n897_li = n894_lo;
  assign n900_li = n897_lo;
  assign n903_li = G37;
  assign n906_li = n903_lo;
  assign n909_li = n906_lo;
  assign n912_li = n909_lo;
  assign n915_li = G38;
  assign n918_li = n915_lo;
  assign n921_li = n918_lo;
  assign n924_li = n921_lo;
  assign n927_li = G39;
  assign n930_li = n927_lo;
  assign n933_li = n930_lo;
  assign n936_li = n933_lo;
  assign n939_li = G40;
  assign n942_li = n939_lo;
  assign n945_li = n942_lo;
  assign n948_li = n945_lo;
  assign n951_li = G41;
  assign n954_li = n951_lo;
  assign n957_li = n954_lo;
  assign n960_li = n957_lo;
  assign n963_li = G42;
  assign n966_li = n963_lo;
  assign n969_li = n966_lo;
  assign n972_li = n969_lo;
  assign n975_li = G43;
  assign n978_li = n975_lo;
  assign n981_li = n978_lo;
  assign n984_li = n981_lo;
  assign n987_li = G44;
  assign n990_li = n987_lo;
  assign n993_li = n990_lo;
  assign n996_li = n993_lo;
  assign n999_li = G45;
  assign n1002_li = n999_lo;
  assign n1005_li = n1002_lo;
  assign n1008_li = n1005_lo;
  assign n1011_li = G46;
  assign n1014_li = n1011_lo;
  assign n1017_li = n1014_lo;
  assign n1020_li = n1017_lo;
  assign n1023_li = G47;
  assign n1026_li = n1023_lo;
  assign n1029_li = n1026_lo;
  assign n1032_li = n1029_lo;
  assign n1035_li = G48;
  assign n1038_li = n1035_lo;
  assign n1041_li = n1038_lo;
  assign n1044_li = n1041_lo;
  assign n1047_li = G49;
  assign n1050_li = n1047_lo;
  assign n1053_li = n1050_lo;
  assign n1056_li = n1053_lo;
  assign n1059_li = G50;
  assign n1062_li = n1059_lo;
  assign n1065_li = n1062_lo;
  assign n1068_li = n1065_lo;
  assign n1071_li = G51;
  assign n1074_li = n1071_lo;
  assign n1077_li = n1074_lo;
  assign n1080_li = n1077_lo;
  assign n1083_li = G52;
  assign n1086_li = n1083_lo;
  assign n1089_li = n1086_lo;
  assign n1092_li = n1089_lo;
  assign n1095_li = G53;
  assign n1098_li = n1095_lo;
  assign n1101_li = n1098_lo;
  assign n1104_li = n1101_lo;
  assign n1107_li = G54;
  assign n1110_li = n1107_lo;
  assign n1113_li = n1110_lo;
  assign n1116_li = n1113_lo;
  assign n1119_li = G55;
  assign n1122_li = n1119_lo;
  assign n1125_li = n1122_lo;
  assign n1128_li = n1125_lo;
  assign n1131_li = G56;
  assign n1134_li = n1131_lo;
  assign n1137_li = n1134_lo;
  assign n1140_li = n1137_lo;
  assign n1143_li = G57;
  assign n1146_li = n1143_lo;
  assign n1149_li = n1146_lo;
  assign n1152_li = n1149_lo;
  assign n1155_li = G58;
  assign n1158_li = n1155_lo;
  assign n1161_li = n1158_lo;
  assign n1164_li = n1161_lo;
  assign n1167_li = G59;
  assign n1170_li = n1167_lo;
  assign n1173_li = n1170_lo;
  assign n1176_li = n1173_lo;
  assign n1179_li = G60;
  assign n1182_li = n1179_lo;
  assign n1185_li = n1182_lo;
  assign n1188_li = n1185_lo;
  always @ (posedge clock) begin
    n471_lo <= n471_li;
    n474_lo <= n474_li;
    n477_lo <= n477_li;
    n480_lo <= n480_li;
    n483_lo <= n483_li;
    n486_lo <= n486_li;
    n489_lo <= n489_li;
    n492_lo <= n492_li;
    n495_lo <= n495_li;
    n498_lo <= n498_li;
    n501_lo <= n501_li;
    n504_lo <= n504_li;
    n507_lo <= n507_li;
    n510_lo <= n510_li;
    n513_lo <= n513_li;
    n516_lo <= n516_li;
    n519_lo <= n519_li;
    n522_lo <= n522_li;
    n525_lo <= n525_li;
    n528_lo <= n528_li;
    n531_lo <= n531_li;
    n534_lo <= n534_li;
    n537_lo <= n537_li;
    n540_lo <= n540_li;
    n543_lo <= n543_li;
    n546_lo <= n546_li;
    n549_lo <= n549_li;
    n552_lo <= n552_li;
    n555_lo <= n555_li;
    n558_lo <= n558_li;
    n561_lo <= n561_li;
    n564_lo <= n564_li;
    n567_lo <= n567_li;
    n570_lo <= n570_li;
    n573_lo <= n573_li;
    n576_lo <= n576_li;
    n579_lo <= n579_li;
    n582_lo <= n582_li;
    n585_lo <= n585_li;
    n588_lo <= n588_li;
    n591_lo <= n591_li;
    n594_lo <= n594_li;
    n597_lo <= n597_li;
    n600_lo <= n600_li;
    n603_lo <= n603_li;
    n606_lo <= n606_li;
    n609_lo <= n609_li;
    n612_lo <= n612_li;
    n615_lo <= n615_li;
    n618_lo <= n618_li;
    n621_lo <= n621_li;
    n624_lo <= n624_li;
    n627_lo <= n627_li;
    n630_lo <= n630_li;
    n633_lo <= n633_li;
    n636_lo <= n636_li;
    n639_lo <= n639_li;
    n642_lo <= n642_li;
    n645_lo <= n645_li;
    n648_lo <= n648_li;
    n651_lo <= n651_li;
    n654_lo <= n654_li;
    n657_lo <= n657_li;
    n660_lo <= n660_li;
    n663_lo <= n663_li;
    n666_lo <= n666_li;
    n669_lo <= n669_li;
    n672_lo <= n672_li;
    n675_lo <= n675_li;
    n678_lo <= n678_li;
    n681_lo <= n681_li;
    n684_lo <= n684_li;
    n687_lo <= n687_li;
    n690_lo <= n690_li;
    n693_lo <= n693_li;
    n696_lo <= n696_li;
    n699_lo <= n699_li;
    n702_lo <= n702_li;
    n705_lo <= n705_li;
    n708_lo <= n708_li;
    n711_lo <= n711_li;
    n714_lo <= n714_li;
    n717_lo <= n717_li;
    n720_lo <= n720_li;
    n723_lo <= n723_li;
    n726_lo <= n726_li;
    n729_lo <= n729_li;
    n732_lo <= n732_li;
    n735_lo <= n735_li;
    n738_lo <= n738_li;
    n741_lo <= n741_li;
    n744_lo <= n744_li;
    n747_lo <= n747_li;
    n750_lo <= n750_li;
    n753_lo <= n753_li;
    n756_lo <= n756_li;
    n759_lo <= n759_li;
    n762_lo <= n762_li;
    n765_lo <= n765_li;
    n768_lo <= n768_li;
    n771_lo <= n771_li;
    n774_lo <= n774_li;
    n777_lo <= n777_li;
    n780_lo <= n780_li;
    n783_lo <= n783_li;
    n786_lo <= n786_li;
    n789_lo <= n789_li;
    n792_lo <= n792_li;
    n795_lo <= n795_li;
    n798_lo <= n798_li;
    n801_lo <= n801_li;
    n804_lo <= n804_li;
    n807_lo <= n807_li;
    n810_lo <= n810_li;
    n813_lo <= n813_li;
    n816_lo <= n816_li;
    n819_lo <= n819_li;
    n822_lo <= n822_li;
    n825_lo <= n825_li;
    n828_lo <= n828_li;
    n831_lo <= n831_li;
    n834_lo <= n834_li;
    n837_lo <= n837_li;
    n840_lo <= n840_li;
    n843_lo <= n843_li;
    n846_lo <= n846_li;
    n849_lo <= n849_li;
    n852_lo <= n852_li;
    n855_lo <= n855_li;
    n858_lo <= n858_li;
    n861_lo <= n861_li;
    n864_lo <= n864_li;
    n867_lo <= n867_li;
    n870_lo <= n870_li;
    n873_lo <= n873_li;
    n876_lo <= n876_li;
    n879_lo <= n879_li;
    n882_lo <= n882_li;
    n885_lo <= n885_li;
    n888_lo <= n888_li;
    n891_lo <= n891_li;
    n894_lo <= n894_li;
    n897_lo <= n897_li;
    n900_lo <= n900_li;
    n903_lo <= n903_li;
    n906_lo <= n906_li;
    n909_lo <= n909_li;
    n912_lo <= n912_li;
    n915_lo <= n915_li;
    n918_lo <= n918_li;
    n921_lo <= n921_li;
    n924_lo <= n924_li;
    n927_lo <= n927_li;
    n930_lo <= n930_li;
    n933_lo <= n933_li;
    n936_lo <= n936_li;
    n939_lo <= n939_li;
    n942_lo <= n942_li;
    n945_lo <= n945_li;
    n948_lo <= n948_li;
    n951_lo <= n951_li;
    n954_lo <= n954_li;
    n957_lo <= n957_li;
    n960_lo <= n960_li;
    n963_lo <= n963_li;
    n966_lo <= n966_li;
    n969_lo <= n969_li;
    n972_lo <= n972_li;
    n975_lo <= n975_li;
    n978_lo <= n978_li;
    n981_lo <= n981_li;
    n984_lo <= n984_li;
    n987_lo <= n987_li;
    n990_lo <= n990_li;
    n993_lo <= n993_li;
    n996_lo <= n996_li;
    n999_lo <= n999_li;
    n1002_lo <= n1002_li;
    n1005_lo <= n1005_li;
    n1008_lo <= n1008_li;
    n1011_lo <= n1011_li;
    n1014_lo <= n1014_li;
    n1017_lo <= n1017_li;
    n1020_lo <= n1020_li;
    n1023_lo <= n1023_li;
    n1026_lo <= n1026_li;
    n1029_lo <= n1029_li;
    n1032_lo <= n1032_li;
    n1035_lo <= n1035_li;
    n1038_lo <= n1038_li;
    n1041_lo <= n1041_li;
    n1044_lo <= n1044_li;
    n1047_lo <= n1047_li;
    n1050_lo <= n1050_li;
    n1053_lo <= n1053_li;
    n1056_lo <= n1056_li;
    n1059_lo <= n1059_li;
    n1062_lo <= n1062_li;
    n1065_lo <= n1065_li;
    n1068_lo <= n1068_li;
    n1071_lo <= n1071_li;
    n1074_lo <= n1074_li;
    n1077_lo <= n1077_li;
    n1080_lo <= n1080_li;
    n1083_lo <= n1083_li;
    n1086_lo <= n1086_li;
    n1089_lo <= n1089_li;
    n1092_lo <= n1092_li;
    n1095_lo <= n1095_li;
    n1098_lo <= n1098_li;
    n1101_lo <= n1101_li;
    n1104_lo <= n1104_li;
    n1107_lo <= n1107_li;
    n1110_lo <= n1110_li;
    n1113_lo <= n1113_li;
    n1116_lo <= n1116_li;
    n1119_lo <= n1119_li;
    n1122_lo <= n1122_li;
    n1125_lo <= n1125_li;
    n1128_lo <= n1128_li;
    n1131_lo <= n1131_li;
    n1134_lo <= n1134_li;
    n1137_lo <= n1137_li;
    n1140_lo <= n1140_li;
    n1143_lo <= n1143_li;
    n1146_lo <= n1146_li;
    n1149_lo <= n1149_li;
    n1152_lo <= n1152_li;
    n1155_lo <= n1155_li;
    n1158_lo <= n1158_li;
    n1161_lo <= n1161_li;
    n1164_lo <= n1164_li;
    n1167_lo <= n1167_li;
    n1170_lo <= n1170_li;
    n1173_lo <= n1173_li;
    n1176_lo <= n1176_li;
    n1179_lo <= n1179_li;
    n1182_lo <= n1182_li;
    n1185_lo <= n1185_li;
    n1188_lo <= n1188_li;
  end
  initial begin
    n471_lo <= 1'b0;
    n474_lo <= 1'b0;
    n477_lo <= 1'b0;
    n480_lo <= 1'b0;
    n483_lo <= 1'b0;
    n486_lo <= 1'b0;
    n489_lo <= 1'b0;
    n492_lo <= 1'b0;
    n495_lo <= 1'b0;
    n498_lo <= 1'b0;
    n501_lo <= 1'b0;
    n504_lo <= 1'b0;
    n507_lo <= 1'b0;
    n510_lo <= 1'b0;
    n513_lo <= 1'b0;
    n516_lo <= 1'b0;
    n519_lo <= 1'b0;
    n522_lo <= 1'b0;
    n525_lo <= 1'b0;
    n528_lo <= 1'b0;
    n531_lo <= 1'b0;
    n534_lo <= 1'b0;
    n537_lo <= 1'b0;
    n540_lo <= 1'b0;
    n543_lo <= 1'b0;
    n546_lo <= 1'b0;
    n549_lo <= 1'b0;
    n552_lo <= 1'b0;
    n555_lo <= 1'b0;
    n558_lo <= 1'b0;
    n561_lo <= 1'b0;
    n564_lo <= 1'b0;
    n567_lo <= 1'b0;
    n570_lo <= 1'b0;
    n573_lo <= 1'b0;
    n576_lo <= 1'b0;
    n579_lo <= 1'b0;
    n582_lo <= 1'b0;
    n585_lo <= 1'b0;
    n588_lo <= 1'b0;
    n591_lo <= 1'b0;
    n594_lo <= 1'b0;
    n597_lo <= 1'b0;
    n600_lo <= 1'b0;
    n603_lo <= 1'b0;
    n606_lo <= 1'b0;
    n609_lo <= 1'b0;
    n612_lo <= 1'b0;
    n615_lo <= 1'b0;
    n618_lo <= 1'b0;
    n621_lo <= 1'b0;
    n624_lo <= 1'b0;
    n627_lo <= 1'b0;
    n630_lo <= 1'b0;
    n633_lo <= 1'b0;
    n636_lo <= 1'b0;
    n639_lo <= 1'b0;
    n642_lo <= 1'b0;
    n645_lo <= 1'b0;
    n648_lo <= 1'b0;
    n651_lo <= 1'b0;
    n654_lo <= 1'b0;
    n657_lo <= 1'b0;
    n660_lo <= 1'b0;
    n663_lo <= 1'b0;
    n666_lo <= 1'b0;
    n669_lo <= 1'b0;
    n672_lo <= 1'b0;
    n675_lo <= 1'b0;
    n678_lo <= 1'b0;
    n681_lo <= 1'b0;
    n684_lo <= 1'b0;
    n687_lo <= 1'b0;
    n690_lo <= 1'b0;
    n693_lo <= 1'b0;
    n696_lo <= 1'b0;
    n699_lo <= 1'b0;
    n702_lo <= 1'b0;
    n705_lo <= 1'b0;
    n708_lo <= 1'b0;
    n711_lo <= 1'b0;
    n714_lo <= 1'b0;
    n717_lo <= 1'b0;
    n720_lo <= 1'b0;
    n723_lo <= 1'b0;
    n726_lo <= 1'b0;
    n729_lo <= 1'b0;
    n732_lo <= 1'b0;
    n735_lo <= 1'b0;
    n738_lo <= 1'b0;
    n741_lo <= 1'b0;
    n744_lo <= 1'b0;
    n747_lo <= 1'b0;
    n750_lo <= 1'b0;
    n753_lo <= 1'b0;
    n756_lo <= 1'b0;
    n759_lo <= 1'b0;
    n762_lo <= 1'b0;
    n765_lo <= 1'b0;
    n768_lo <= 1'b0;
    n771_lo <= 1'b0;
    n774_lo <= 1'b0;
    n777_lo <= 1'b0;
    n780_lo <= 1'b0;
    n783_lo <= 1'b0;
    n786_lo <= 1'b0;
    n789_lo <= 1'b0;
    n792_lo <= 1'b0;
    n795_lo <= 1'b0;
    n798_lo <= 1'b0;
    n801_lo <= 1'b0;
    n804_lo <= 1'b0;
    n807_lo <= 1'b0;
    n810_lo <= 1'b0;
    n813_lo <= 1'b0;
    n816_lo <= 1'b0;
    n819_lo <= 1'b0;
    n822_lo <= 1'b0;
    n825_lo <= 1'b0;
    n828_lo <= 1'b0;
    n831_lo <= 1'b0;
    n834_lo <= 1'b0;
    n837_lo <= 1'b0;
    n840_lo <= 1'b0;
    n843_lo <= 1'b0;
    n846_lo <= 1'b0;
    n849_lo <= 1'b0;
    n852_lo <= 1'b0;
    n855_lo <= 1'b0;
    n858_lo <= 1'b0;
    n861_lo <= 1'b0;
    n864_lo <= 1'b0;
    n867_lo <= 1'b0;
    n870_lo <= 1'b0;
    n873_lo <= 1'b0;
    n876_lo <= 1'b0;
    n879_lo <= 1'b0;
    n882_lo <= 1'b0;
    n885_lo <= 1'b0;
    n888_lo <= 1'b0;
    n891_lo <= 1'b0;
    n894_lo <= 1'b0;
    n897_lo <= 1'b0;
    n900_lo <= 1'b0;
    n903_lo <= 1'b0;
    n906_lo <= 1'b0;
    n909_lo <= 1'b0;
    n912_lo <= 1'b0;
    n915_lo <= 1'b0;
    n918_lo <= 1'b0;
    n921_lo <= 1'b0;
    n924_lo <= 1'b0;
    n927_lo <= 1'b0;
    n930_lo <= 1'b0;
    n933_lo <= 1'b0;
    n936_lo <= 1'b0;
    n939_lo <= 1'b0;
    n942_lo <= 1'b0;
    n945_lo <= 1'b0;
    n948_lo <= 1'b0;
    n951_lo <= 1'b0;
    n954_lo <= 1'b0;
    n957_lo <= 1'b0;
    n960_lo <= 1'b0;
    n963_lo <= 1'b0;
    n966_lo <= 1'b0;
    n969_lo <= 1'b0;
    n972_lo <= 1'b0;
    n975_lo <= 1'b0;
    n978_lo <= 1'b0;
    n981_lo <= 1'b0;
    n984_lo <= 1'b0;
    n987_lo <= 1'b0;
    n990_lo <= 1'b0;
    n993_lo <= 1'b0;
    n996_lo <= 1'b0;
    n999_lo <= 1'b0;
    n1002_lo <= 1'b0;
    n1005_lo <= 1'b0;
    n1008_lo <= 1'b0;
    n1011_lo <= 1'b0;
    n1014_lo <= 1'b0;
    n1017_lo <= 1'b0;
    n1020_lo <= 1'b0;
    n1023_lo <= 1'b0;
    n1026_lo <= 1'b0;
    n1029_lo <= 1'b0;
    n1032_lo <= 1'b0;
    n1035_lo <= 1'b0;
    n1038_lo <= 1'b0;
    n1041_lo <= 1'b0;
    n1044_lo <= 1'b0;
    n1047_lo <= 1'b0;
    n1050_lo <= 1'b0;
    n1053_lo <= 1'b0;
    n1056_lo <= 1'b0;
    n1059_lo <= 1'b0;
    n1062_lo <= 1'b0;
    n1065_lo <= 1'b0;
    n1068_lo <= 1'b0;
    n1071_lo <= 1'b0;
    n1074_lo <= 1'b0;
    n1077_lo <= 1'b0;
    n1080_lo <= 1'b0;
    n1083_lo <= 1'b0;
    n1086_lo <= 1'b0;
    n1089_lo <= 1'b0;
    n1092_lo <= 1'b0;
    n1095_lo <= 1'b0;
    n1098_lo <= 1'b0;
    n1101_lo <= 1'b0;
    n1104_lo <= 1'b0;
    n1107_lo <= 1'b0;
    n1110_lo <= 1'b0;
    n1113_lo <= 1'b0;
    n1116_lo <= 1'b0;
    n1119_lo <= 1'b0;
    n1122_lo <= 1'b0;
    n1125_lo <= 1'b0;
    n1128_lo <= 1'b0;
    n1131_lo <= 1'b0;
    n1134_lo <= 1'b0;
    n1137_lo <= 1'b0;
    n1140_lo <= 1'b0;
    n1143_lo <= 1'b0;
    n1146_lo <= 1'b0;
    n1149_lo <= 1'b0;
    n1152_lo <= 1'b0;
    n1155_lo <= 1'b0;
    n1158_lo <= 1'b0;
    n1161_lo <= 1'b0;
    n1164_lo <= 1'b0;
    n1167_lo <= 1'b0;
    n1170_lo <= 1'b0;
    n1173_lo <= 1'b0;
    n1176_lo <= 1'b0;
    n1179_lo <= 1'b0;
    n1182_lo <= 1'b0;
    n1185_lo <= 1'b0;
    n1188_lo <= 1'b0;
  end
endmodule


