// Benchmark "mymod" written by ABC on Sun Oct 29 23:44:44 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58,
    G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70, G71, G72,
    G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86,
    G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G109, G110, G111, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G124,
    G125, G126, G127, G128, G129, G130, G131, G132, G133, G134, G135, G136,
    G137, G138, G139, G140, G141, G142, G143, G144, G145, G146, G147, G148,
    G149, G150, G151, G152, G153, G154, G155, G156, G157,
    G2531, G2532, G2533, G2534, G2535, G2536, G2537, G2538, G2539, G2540,
    G2541, G2542, G2543, G2544, G2545, G2546, G2547, G2548, G2549, G2550,
    G2551, G2552, G2553, G2554, G2555, G2556, G2557, G2558, G2559, G2560,
    G2561, G2562, G2563, G2564, G2565, G2566, G2567, G2568, G2569, G2570,
    G2571, G2572, G2573, G2574, G2575, G2576, G2577, G2578, G2579, G2580,
    G2581, G2582, G2583, G2584, G2585, G2586, G2587, G2588, G2589, G2590,
    G2591, G2592, G2593, G2594  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70,
    G71, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98,
    G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G110,
    G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G133, G134,
    G135, G136, G137, G138, G139, G140, G141, G142, G143, G144, G145, G146,
    G147, G148, G149, G150, G151, G152, G153, G154, G155, G156, G157;
  output G2531, G2532, G2533, G2534, G2535, G2536, G2537, G2538, G2539, G2540,
    G2541, G2542, G2543, G2544, G2545, G2546, G2547, G2548, G2549, G2550,
    G2551, G2552, G2553, G2554, G2555, G2556, G2557, G2558, G2559, G2560,
    G2561, G2562, G2563, G2564, G2565, G2566, G2567, G2568, G2569, G2570,
    G2571, G2572, G2573, G2574, G2575, G2576, G2577, G2578, G2579, G2580,
    G2581, G2582, G2583, G2584, G2585, G2586, G2587, G2588, G2589, G2590,
    G2591, G2592, G2593, G2594;
  reg n1416_lo, n1419_lo, n1422_lo, n1425_lo, n1428_lo, n1431_lo, n1434_lo,
    n1437_lo, n1440_lo, n1443_lo, n1446_lo, n1449_lo, n1452_lo, n1455_lo,
    n1458_lo, n1464_lo, n1467_lo, n1470_lo, n1476_lo, n1479_lo, n1482_lo,
    n1488_lo, n1491_lo, n1494_lo, n1497_lo, n1500_lo, n1503_lo, n1512_lo,
    n1515_lo, n1518_lo, n1521_lo, n1524_lo, n1527_lo, n1530_lo, n1533_lo,
    n1536_lo, n1539_lo, n1542_lo, n1545_lo, n1548_lo, n1551_lo, n1554_lo,
    n1560_lo, n1563_lo, n1566_lo, n1572_lo, n1575_lo, n1578_lo, n1584_lo,
    n1587_lo, n1590_lo, n1596_lo, n1599_lo, n1602_lo, n1608_lo, n1611_lo,
    n1614_lo, n1620_lo, n1623_lo, n1626_lo, n1632_lo, n1635_lo, n1638_lo,
    n1644_lo, n1647_lo, n1650_lo, n1656_lo, n1659_lo, n1662_lo, n1668_lo,
    n1671_lo, n1674_lo, n1680_lo, n1683_lo, n1686_lo, n1692_lo, n1695_lo,
    n1698_lo, n1704_lo, n1707_lo, n1710_lo, n1716_lo, n1719_lo, n1722_lo,
    n1728_lo, n1731_lo, n1734_lo, n1740_lo, n1743_lo, n1746_lo, n1749_lo,
    n1752_lo, n1755_lo, n1758_lo, n1761_lo, n1764_lo, n1776_lo, n1788_lo,
    n1791_lo, n1794_lo, n1797_lo, n1800_lo, n1803_lo, n1812_lo, n1815_lo,
    n1824_lo, n1827_lo, n1836_lo, n1839_lo, n1848_lo, n1851_lo, n1860_lo,
    n1872_lo, n1875_lo, n1884_lo, n1896_lo, n1899_lo, n1908_lo, n1920_lo,
    n1923_lo, n1926_lo, n1929_lo, n1932_lo, n1935_lo, n1944_lo, n1947_lo,
    n1956_lo, n1959_lo, n1962_lo, n1968_lo, n1971_lo, n1980_lo, n1983_lo,
    n1992_lo, n1995_lo, n2004_lo, n2016_lo, n2019_lo, n2028_lo, n2040_lo,
    n2043_lo, n2046_lo, n2049_lo, n2052_lo, n2055_lo, n2064_lo, n2067_lo,
    n2076_lo, n2079_lo, n2088_lo, n2091_lo, n2100_lo, n2103_lo, n2112_lo,
    n2115_lo, n2124_lo, n2127_lo, n2136_lo, n2148_lo, n2151_lo, n2160_lo,
    n2172_lo, n2175_lo, n2178_lo, n2181_lo, n2184_lo, n2187_lo, n2196_lo,
    n2199_lo, n2208_lo, n2211_lo, n2220_lo, n2223_lo, n2232_lo, n2235_lo,
    n2244_lo, n2247_lo, n2256_lo, n2259_lo, n2268_lo, n2280_lo, n2283_lo,
    n2292_lo, n2295_lo, n2298_lo, n2301_lo, n2304_lo, n2307_lo, n2316_lo,
    n2319_lo, n2322_lo, n2325_lo, n2328_lo, n2331_lo, n2340_lo, n2343_lo,
    n2376_lo, n2379_lo, n2388_lo, n2391_lo, n2400_lo, n2403_lo, n2412_lo,
    n2415_lo, n2424_lo, n2427_lo, n2436_lo, n2439_lo, n2442_lo, n2445_lo,
    n2448_lo, n2451_lo, n2460_lo, n2463_lo, n2496_lo, n2499_lo, n2508_lo,
    n2511_lo, n2520_lo, n2523_lo, n2532_lo, n2535_lo, n2544_lo, n2547_lo,
    n2556_lo, n2559_lo, n2562_lo, n2565_lo, n2568_lo, n2571_lo, n2580_lo,
    n2583_lo, n2616_lo, n2619_lo, n2628_lo, n2631_lo, n2640_lo, n2643_lo,
    n2652_lo, n2655_lo, n2664_lo, n2667_lo, n2676_lo, n2679_lo, n2682_lo,
    n2685_lo, n2688_lo, n2691_lo, n2700_lo, n2703_lo, n2736_lo, n2739_lo,
    n2748_lo, n2751_lo, n2760_lo, n2763_lo, n2772_lo, n2775_lo, n2784_lo,
    n2787_lo, n2790_lo, n2793_lo, n2796_lo, n2799_lo, n2802_lo, n2805_lo,
    n2808_lo, n2820_lo, n2823_lo, n2826_lo, n2829_lo, n2832_lo, n2835_lo,
    n2838_lo, n2841_lo, n2844_lo, n2856_lo, n2859_lo, n2862_lo, n2865_lo,
    n2868_lo, n2871_lo, n2874_lo, n2877_lo, n2880_lo, n2883_lo, n2886_lo,
    n2889_lo, n2892_lo, n2895_lo, n2898_lo, n2901_lo, n2904_lo, n2907_lo,
    n2916_lo, n2919_lo, n2925_lo, n2928_lo, n2940_lo, n2943_lo, n2952_lo,
    n2955_lo, n2961_lo, n2964_lo, n2967_lo, n2970_lo, n2976_lo, n2979_lo,
    n2982_lo, n2988_lo, n2991_lo, n2994_lo, n2997_lo, n3000_lo, n3003_lo,
    n3006_lo, n3012_lo, n3015_lo, n3018_lo, n3021_lo, n3024_lo, n3027_lo,
    n3030_lo, n3033_lo, n3036_lo, n3039_lo, n3045_lo, n3048_lo, n3051_lo,
    n3054_lo, n3057_lo, n3060_lo, n3063_lo, n3069_lo, n3072_lo, n3075_lo,
    n3081_lo, n3084_lo, n3087_lo, n3093_lo, n3096_lo, n3099_lo, n3102_lo,
    n3105_lo, n3108_lo, n3111_lo, n3114_lo, n3117_lo, n3120_lo, n3123_lo,
    n3126_lo, n3129_lo, n3132_lo, n3135_lo, n3138_lo, n3141_lo, n3156_lo,
    n3168_lo, n3171_lo, n3174_lo, n3177_lo, n3180_lo, n3183_lo, n3192_lo,
    n3195_lo, n3204_lo, n3207_lo, n3210_lo, n3216_lo, n3219_lo, n3222_lo,
    n3228_lo, n3231_lo, n3240_lo, n3243_lo, n3252_lo, n3255_lo, n3258_lo,
    n3264_lo, n3267_lo, n3270_lo, n3276_lo, n3279_lo, n3282_lo, n3288_lo,
    n3291_lo, n3294_lo, n3603_o2, n3604_o2, n1391_inv, n3798_o2, n3846_o2,
    n4019_o2, n4017_o2, n2177_o2, n2150_o2, n2154_o2, n2184_o2, n2515_o2,
    n3837_o2, n2167_o2, n2118_o2, n2186_o2, n2174_o2, n3964_o2, n4005_o2,
    n4006_o2, n1445_inv, n2176_o2, n2227_o2, n2236_o2, n2245_o2, n2518_o2,
    n4023_o2, n1466_inv, n4038_o2, n4039_o2, n1475_inv, n2119_o2, n2275_o2,
    n2595_o2, n2594_o2, lo498_buf_o2, lo502_buf_o2, lo550_buf_o2, n2596_o2,
    n2593_o2, n2668_o2, lo542_buf_o2, n2667_o2, n2404_o2, n2410_o2,
    n2419_o2, n2392_o2, n2369_o2, n2397_o2, n2601_o2, n2658_o2, n2574_o2,
    n2205_o2, lo510_buf_o2, lo514_buf_o2, lo554_buf_o2, lo558_buf_o2,
    lo578_buf_o2, n2254_o2, n2421_o2, n2422_o2, n2130_o2, n2127_o2,
    n2131_o2, n2128_o2, n2264_o2, n2467_o2, n2471_o2, n2488_o2, n2478_o2,
    n2486_o2, n2485_o2, n2498_o2, n2495_o2, n2496_o2, n2458_o2, n2643_o2,
    n2462_o2, n2468_o2, n2639_o2, n2499_o2, n2472_o2, n2474_o2, n2489_o2,
    n2321_o2, n2322_o2, n2640_o2, n2642_o2, n2187_o2, n2373_o2, n2603_o2,
    n2388_o2, n2437_o2, n2356_o2, n2452_o2, n2347_o2, n2329_o2, n2669_o2,
    n2332_o2, n2664_o2, n2665_o2, n2653_o2, n2654_o2, n2636_o2, n2660_o2,
    n2318_o2, n2319_o2, n2586_o2, n2587_o2, n2288_o2, n2344_o2, n2530_o2,
    n2303_o2, n2566_o2, n2567_o2, n2554_o2, n2194_o2, lo582_buf_o2,
    lo030_buf_o2, lo174_buf_o2, lo178_buf_o2, lo186_buf_o2, lo266_buf_o2,
    lo306_buf_o2, lo346_buf_o2, lo386_buf_o2, lo426_buf_o2, lo590_buf_o2,
    lo594_buf_o2, lo606_buf_o2, lo610_buf_o2, n2238_o2, n2229_o2, n2242_o2,
    n2233_o2, n2168_o2, n2237_o2, n2228_o2, n2172_o2, n2223_o2, n2222_o2,
    n2170_o2, n2181_o2, n2510_o2, n2621_o2, lo466_buf_o2, lo478_buf_o2,
    n2149_o2, n2429_o2, n2444_o2, n2153_o2, n2433_o2, n2448_o2, n2367_o2,
    n2386_o2, n2539_o2, n2183_o2, n2220_o2, n2514_o2, n2196_o2, n2616_o2,
    n2612_o2, n2627_o2, n2140_o2, n1877_inv, lo149_buf_o2, lo197_buf_o2,
    lo118_buf_o2, lo158_buf_o2, lo166_buf_o2, lo242_buf_o2, lo286_buf_o2,
    lo506_buf_o2, n2198_o2, n2202_o2, n2197_o2, n1913_inv, n2146_o2,
    n1919_inv, lo312_buf_o2, lo316_buf_o2, lo352_buf_o2, lo356_buf_o2,
    lo392_buf_o2, lo396_buf_o2, lo432_buf_o2, lo436_buf_o2, lo576_buf_o2;
  wire new_new_n1372__, new_new_n1374__, new_new_n1376__, new_new_n1378__,
    new_new_n1380__, new_new_n1382__, new_new_n1384__, new_new_n1386__,
    new_new_n1388__, new_new_n1390__, new_new_n1392__, new_new_n1394__,
    new_new_n1396__, new_new_n1398__, new_new_n1400__, new_new_n1402__,
    new_new_n1404__, new_new_n1406__, new_new_n1408__, new_new_n1410__,
    new_new_n1412__, new_new_n1414__, new_new_n1416__, new_new_n1418__,
    new_new_n1420__, new_new_n1422__, new_new_n1424__, new_new_n1426__,
    new_new_n1428__, new_new_n1430__, new_new_n1432__, new_new_n1434__,
    new_new_n1436__, new_new_n1438__, new_new_n1440__, new_new_n1442__,
    new_new_n1444__, new_new_n1446__, new_new_n1448__, new_new_n1450__,
    new_new_n1452__, new_new_n1454__, new_new_n1456__, new_new_n1458__,
    new_new_n1460__, new_new_n1462__, new_new_n1464__, new_new_n1466__,
    new_new_n1468__, new_new_n1470__, new_new_n1472__, new_new_n1474__,
    new_new_n1476__, new_new_n1478__, new_new_n1480__, new_new_n1482__,
    new_new_n1484__, new_new_n1486__, new_new_n1488__, new_new_n1490__,
    new_new_n1492__, new_new_n1494__, new_new_n1496__, new_new_n1498__,
    new_new_n1500__, new_new_n1502__, new_new_n1504__, new_new_n1506__,
    new_new_n1508__, new_new_n1510__, new_new_n1512__, new_new_n1514__,
    new_new_n1516__, new_new_n1518__, new_new_n1520__, new_new_n1522__,
    new_new_n1524__, new_new_n1526__, new_new_n1528__, new_new_n1530__,
    new_new_n1532__, new_new_n1534__, new_new_n1536__, new_new_n1538__,
    new_new_n1540__, new_new_n1542__, new_new_n1544__, new_new_n1546__,
    new_new_n1548__, new_new_n1550__, new_new_n1552__, new_new_n1554__,
    new_new_n1556__, new_new_n1558__, new_new_n1560__, new_new_n1562__,
    new_new_n1564__, new_new_n1566__, new_new_n1568__, new_new_n1570__,
    new_new_n1572__, new_new_n1574__, new_new_n1576__, new_new_n1578__,
    new_new_n1580__, new_new_n1582__, new_new_n1584__, new_new_n1586__,
    new_new_n1588__, new_new_n1590__, new_new_n1592__, new_new_n1594__,
    new_new_n1596__, new_new_n1598__, new_new_n1600__, new_new_n1602__,
    new_new_n1604__, new_new_n1606__, new_new_n1608__, new_new_n1610__,
    new_new_n1612__, new_new_n1614__, new_new_n1616__, new_new_n1618__,
    new_new_n1620__, new_new_n1622__, new_new_n1624__, new_new_n1626__,
    new_new_n1628__, new_new_n1630__, new_new_n1632__, new_new_n1634__,
    new_new_n1636__, new_new_n1638__, new_new_n1640__, new_new_n1642__,
    new_new_n1644__, new_new_n1646__, new_new_n1648__, new_new_n1650__,
    new_new_n1652__, new_new_n1654__, new_new_n1656__, new_new_n1658__,
    new_new_n1660__, new_new_n1662__, new_new_n1664__, new_new_n1666__,
    new_new_n1668__, new_new_n1670__, new_new_n1672__, new_new_n1674__,
    new_new_n1676__, new_new_n1678__, new_new_n1680__, new_new_n1682__,
    new_new_n1684__, new_new_n1686__, new_new_n1688__, new_new_n1690__,
    new_new_n1692__, new_new_n1694__, new_new_n1696__, new_new_n1698__,
    new_new_n1701__, new_new_n1702__, new_new_n1704__, new_new_n1706__,
    new_new_n1708__, new_new_n1710__, new_new_n1712__, new_new_n1714__,
    new_new_n1716__, new_new_n1718__, new_new_n1720__, new_new_n1722__,
    new_new_n1724__, new_new_n1726__, new_new_n1728__, new_new_n1730__,
    new_new_n1732__, new_new_n1735__, new_new_n1736__, new_new_n1738__,
    new_new_n1740__, new_new_n1742__, new_new_n1744__, new_new_n1747__,
    new_new_n1748__, new_new_n1750__, new_new_n1752__, new_new_n1754__,
    new_new_n1756__, new_new_n1758__, new_new_n1760__, new_new_n1763__,
    new_new_n1764__, new_new_n1766__, new_new_n1768__, new_new_n1769__,
    new_new_n1770__, new_new_n1772__, new_new_n1774__, new_new_n1776__,
    new_new_n1778__, new_new_n1780__, new_new_n1782__, new_new_n1784__,
    new_new_n1786__, new_new_n1788__, new_new_n1790__, new_new_n1792__,
    new_new_n1794__, new_new_n1796__, new_new_n1798__, new_new_n1800__,
    new_new_n1802__, new_new_n1804__, new_new_n1806__, new_new_n1808__,
    new_new_n1810__, new_new_n1812__, new_new_n1814__, new_new_n1816__,
    new_new_n1818__, new_new_n1820__, new_new_n1822__, new_new_n1824__,
    new_new_n1826__, new_new_n1828__, new_new_n1830__, new_new_n1832__,
    new_new_n1834__, new_new_n1835__, new_new_n1836__, new_new_n1838__,
    new_new_n1840__, new_new_n1842__, new_new_n1844__, new_new_n1846__,
    new_new_n1848__, new_new_n1850__, new_new_n1852__, new_new_n1854__,
    new_new_n1856__, new_new_n1858__, new_new_n1860__, new_new_n1862__,
    new_new_n1864__, new_new_n1867__, new_new_n1868__, new_new_n1870__,
    new_new_n1872__, new_new_n1875__, new_new_n1876__, new_new_n1878__,
    new_new_n1880__, new_new_n1882__, new_new_n1884__, new_new_n1887__,
    new_new_n1888__, new_new_n1890__, new_new_n1892__, new_new_n1894__,
    new_new_n1896__, new_new_n1899__, new_new_n1900__, new_new_n1903__,
    new_new_n1904__, new_new_n1907__, new_new_n1908__, new_new_n1910__,
    new_new_n1912__, new_new_n1914__, new_new_n1916__, new_new_n1918__,
    new_new_n1920__, new_new_n1922__, new_new_n1924__, new_new_n1926__,
    new_new_n1929__, new_new_n1930__, new_new_n1932__, new_new_n1934__,
    new_new_n1936__, new_new_n1938__, new_new_n1940__, new_new_n1942__,
    new_new_n1943__, new_new_n1944__, new_new_n1946__, new_new_n1948__,
    new_new_n1951__, new_new_n1952__, new_new_n1954__, new_new_n1956__,
    new_new_n1958__, new_new_n1960__, new_new_n1962__, new_new_n1964__,
    new_new_n1966__, new_new_n1968__, new_new_n1971__, new_new_n1972__,
    new_new_n1974__, new_new_n1976__, new_new_n1978__, new_new_n1980__,
    new_new_n1982__, new_new_n1984__, new_new_n1986__, new_new_n1988__,
    new_new_n1990__, new_new_n1992__, new_new_n1995__, new_new_n1996__,
    new_new_n1998__, new_new_n2000__, new_new_n2002__, new_new_n2004__,
    new_new_n2006__, new_new_n2008__, new_new_n2010__, new_new_n2012__,
    new_new_n2015__, new_new_n2016__, new_new_n2018__, new_new_n2020__,
    new_new_n2022__, new_new_n2024__, new_new_n2026__, new_new_n2028__,
    new_new_n2031__, new_new_n2032__, new_new_n2035__, new_new_n2036__,
    new_new_n2039__, new_new_n2040__, new_new_n2042__, new_new_n2044__,
    new_new_n2046__, new_new_n2048__, new_new_n2050__, new_new_n2052__,
    new_new_n2054__, new_new_n2056__, new_new_n2058__, new_new_n2060__,
    new_new_n2062__, new_new_n2064__, new_new_n2066__, new_new_n2069__,
    new_new_n2070__, new_new_n2072__, new_new_n2074__, new_new_n2076__,
    new_new_n2078__, new_new_n2080__, new_new_n2082__, new_new_n2084__,
    new_new_n2086__, new_new_n2088__, new_new_n2090__, new_new_n2092__,
    new_new_n2094__, new_new_n2096__, new_new_n2098__, new_new_n2100__,
    new_new_n2102__, new_new_n2105__, new_new_n2106__, new_new_n2108__,
    new_new_n2110__, new_new_n2112__, new_new_n2114__, new_new_n2116__,
    new_new_n2118__, new_new_n2120__, new_new_n2122__, new_new_n2124__,
    new_new_n2126__, new_new_n2128__, new_new_n2130__, new_new_n2132__,
    new_new_n2134__, new_new_n2136__, new_new_n2138__, new_new_n2141__,
    new_new_n2142__, new_new_n2144__, new_new_n2146__, new_new_n2148__,
    new_new_n2150__, new_new_n2152__, new_new_n2154__, new_new_n2156__,
    new_new_n2158__, new_new_n2160__, new_new_n2162__, new_new_n2164__,
    new_new_n2166__, new_new_n2168__, new_new_n2170__, new_new_n2172__,
    new_new_n2174__, new_new_n2177__, new_new_n2178__, new_new_n2180__,
    new_new_n2182__, new_new_n2184__, new_new_n2186__, new_new_n2188__,
    new_new_n2190__, new_new_n2192__, new_new_n2194__, new_new_n2196__,
    new_new_n2198__, new_new_n2200__, new_new_n2202__, new_new_n2204__,
    new_new_n2206__, new_new_n2208__, new_new_n2209__, new_new_n2210__,
    new_new_n2212__, new_new_n2214__, new_new_n2217__, new_new_n2218__,
    new_new_n2219__, new_new_n2220__, new_new_n2222__, new_new_n2224__,
    new_new_n2226__, new_new_n2227__, new_new_n2228__, new_new_n2230__,
    new_new_n2232__, new_new_n2234__, new_new_n2235__, new_new_n2236__,
    new_new_n2237__, new_new_n2238__, new_new_n2240__, new_new_n2242__,
    new_new_n2244__, new_new_n2245__, new_new_n2246__, new_new_n2248__,
    new_new_n2250__, new_new_n2252__, new_new_n2253__, new_new_n2254__,
    new_new_n2256__, new_new_n2258__, new_new_n2260__, new_new_n2261__,
    new_new_n2262__, new_new_n2264__, new_new_n2266__, new_new_n2269__,
    new_new_n2270__, new_new_n2272__, new_new_n2274__, new_new_n2276__,
    new_new_n2279__, new_new_n2280__, new_new_n2282__, new_new_n2284__,
    new_new_n2286__, new_new_n2288__, new_new_n2290__, new_new_n2291__,
    new_new_n2292__, new_new_n2294__, new_new_n2296__, new_new_n2297__,
    new_new_n2298__, new_new_n2300__, new_new_n2302__, new_new_n2303__,
    new_new_n2304__, new_new_n2306__, new_new_n2308__, new_new_n2309__,
    new_new_n2310__, new_new_n2312__, new_new_n2314__, new_new_n2316__,
    new_new_n2317__, new_new_n2318__, new_new_n2320__, new_new_n2322__,
    new_new_n2323__, new_new_n2325__, new_new_n2326__, new_new_n2328__,
    new_new_n2330__, new_new_n2331__, new_new_n2332__, new_new_n2333__,
    new_new_n2334__, new_new_n2336__, new_new_n2338__, new_new_n2339__,
    new_new_n2340__, new_new_n2342__, new_new_n2344__, new_new_n2347__,
    new_new_n2348__, new_new_n2350__, new_new_n2352__, new_new_n2353__,
    new_new_n2354__, new_new_n2356__, new_new_n2358__, new_new_n2360__,
    new_new_n2362__, new_new_n2365__, new_new_n2366__, new_new_n2368__,
    new_new_n2370__, new_new_n2371__, new_new_n2372__, new_new_n2374__,
    new_new_n2376__, new_new_n2378__, new_new_n2379__, new_new_n2380__,
    new_new_n2381__, new_new_n2382__, new_new_n2384__, new_new_n2386__,
    new_new_n2387__, new_new_n2388__, new_new_n2389__, new_new_n2390__,
    new_new_n2392__, new_new_n2394__, new_new_n2395__, new_new_n2396__,
    new_new_n2398__, new_new_n2399__, new_new_n2400__, new_new_n2402__,
    new_new_n2404__, new_new_n2406__, new_new_n2407__, new_new_n2408__,
    new_new_n2410__, new_new_n2412__, new_new_n2414__, new_new_n2416__,
    new_new_n2418__, new_new_n2420__, new_new_n2421__, new_new_n2422__,
    new_new_n2424__, new_new_n2426__, new_new_n2427__, new_new_n2428__,
    new_new_n2430__, new_new_n2432__, new_new_n2434__, new_new_n2436__,
    new_new_n2438__, new_new_n2440__, new_new_n2441__, new_new_n2442__,
    new_new_n2444__, new_new_n2446__, new_new_n2447__, new_new_n2448__,
    new_new_n2450__, new_new_n2452__, new_new_n2453__, new_new_n2454__,
    new_new_n2456__, new_new_n2458__, new_new_n2459__, new_new_n2461__,
    new_new_n2463__, new_new_n2465__, new_new_n2466__, new_new_n2467__,
    new_new_n2468__, new_new_n2469__, new_new_n2470__, new_new_n2472__,
    new_new_n2473__, new_new_n2474__, new_new_n2477__, new_new_n2479__,
    new_new_n2480__, new_new_n2482__, new_new_n2484__, new_new_n2485__,
    new_new_n2487__, new_new_n2489__, new_new_n2490__, new_new_n2493__,
    new_new_n2494__, new_new_n2495__, new_new_n2496__, new_new_n2497__,
    new_new_n2498__, new_new_n2499__, new_new_n2501__, new_new_n2502__,
    new_new_n2504__, new_new_n2506__, new_new_n2508__, new_new_n2510__,
    new_new_n2511__, new_new_n2512__, new_new_n2514__, new_new_n2516__,
    new_new_n2517__, new_new_n2518__, new_new_n2519__, new_new_n2520__,
    new_new_n2521__, new_new_n2523__, new_new_n2524__, new_new_n2525__,
    new_new_n2526__, new_new_n2527__, new_new_n2528__, new_new_n2529__,
    new_new_n2530__, new_new_n2531__, new_new_n2532__, new_new_n2533__,
    new_new_n2534__, new_new_n2535__, new_new_n2536__, new_new_n2537__,
    new_new_n2538__, new_new_n2541__, new_new_n2542__, new_new_n2543__,
    new_new_n2544__, new_new_n2546__, new_new_n2548__, new_new_n2551__,
    new_new_n2552__, new_new_n2555__, new_new_n2557__, new_new_n2559__,
    new_new_n2561__, new_new_n2562__, new_new_n2563__, new_new_n2564__,
    new_new_n2565__, new_new_n2566__, new_new_n2567__, new_new_n2568__,
    new_new_n2569__, new_new_n2570__, new_new_n2571__, new_new_n2572__,
    new_new_n2573__, new_new_n2574__, new_new_n2575__, new_new_n2576__,
    new_new_n2577__, new_new_n2579__, new_new_n2581__, new_new_n2583__,
    new_new_n2585__, new_new_n2587__, new_new_n2589__, new_new_n2590__,
    new_new_n2591__, new_new_n2592__, new_new_n2594__, new_new_n2596__,
    new_new_n2598__, new_new_n2600__, new_new_n2602__, new_new_n2604__,
    new_new_n2606__, new_new_n2608__, new_new_n2610__, new_new_n2612__,
    new_new_n2613__, new_new_n2614__, new_new_n2616__, new_new_n2618__,
    new_new_n2619__, new_new_n2620__, new_new_n2622__, new_new_n2624__,
    new_new_n2626__, new_new_n2628__, new_new_n2629__, new_new_n2630__,
    new_new_n2631__, new_new_n2632__, new_new_n2634__, new_new_n2636__,
    new_new_n2637__, new_new_n2638__, new_new_n2639__, new_new_n2640__,
    new_new_n2642__, new_new_n2643__, new_new_n2644__, new_new_n2645__,
    new_new_n2646__, new_new_n2647__, new_new_n2648__, new_new_n2649__,
    new_new_n2650__, new_new_n2651__, new_new_n2652__, new_new_n2653__,
    new_new_n2654__, new_new_n2655__, new_new_n2656__, new_new_n2657__,
    new_new_n2658__, new_new_n2659__, new_new_n2660__, new_new_n2662__,
    new_new_n2663__, new_new_n2664__, new_new_n2666__, new_new_n2668__,
    new_new_n2670__, new_new_n2671__, new_new_n2672__, new_new_n2673__,
    new_new_n2674__, new_new_n2675__, new_new_n2676__, new_new_n2677__,
    new_new_n2678__, new_new_n2679__, new_new_n2680__, new_new_n2681__,
    new_new_n2682__, new_new_n2683__, new_new_n2684__, new_new_n2685__,
    new_new_n2686__, new_new_n2687__, new_new_n2688__, new_new_n2689__,
    new_new_n2690__, new_new_n2691__, new_new_n2692__, new_new_n2693__,
    new_new_n2694__, new_new_n2695__, new_new_n2696__, new_new_n2697__,
    new_new_n2698__, new_new_n2699__, new_new_n2700__, new_new_n2701__,
    new_new_n2702__, new_new_n2703__, new_new_n2704__, new_new_n2705__,
    new_new_n2706__, new_new_n2707__, new_new_n2708__, new_new_n2709__,
    new_new_n2710__, new_new_n2711__, new_new_n2712__, new_new_n2713__,
    new_new_n2714__, new_new_n2715__, new_new_n2716__, new_new_n2717__,
    new_new_n2718__, new_new_n2719__, new_new_n2720__, new_new_n2721__,
    new_new_n2722__, new_new_n2723__, new_new_n2724__, new_new_n2725__,
    new_new_n2726__, new_new_n2727__, new_new_n2728__, new_new_n2729__,
    new_new_n2730__, new_new_n2731__, new_new_n2732__, new_new_n2733__,
    new_new_n2734__, new_new_n2735__, new_new_n2736__, new_new_n2737__,
    new_new_n2738__, new_new_n2739__, new_new_n2740__, new_new_n2741__,
    new_new_n2742__, new_new_n2743__, new_new_n2744__, new_new_n2745__,
    new_new_n2746__, new_new_n2747__, new_new_n2749__, new_new_n2750__,
    new_new_n2751__, new_new_n2752__, new_new_n2753__, new_new_n2754__,
    new_new_n2755__, new_new_n2756__, new_new_n2757__, new_new_n2758__,
    new_new_n2759__, new_new_n2760__, new_new_n2761__, new_new_n2762__,
    new_new_n2763__, new_new_n2764__, new_new_n2765__, new_new_n2766__,
    new_new_n2767__, new_new_n2768__, new_new_n2769__, new_new_n2770__,
    new_new_n2771__, new_new_n2772__, new_new_n2773__, new_new_n2774__,
    new_new_n2775__, new_new_n2776__, new_new_n2777__, new_new_n2778__,
    new_new_n2781__, new_new_n2783__, new_new_n2785__, new_new_n2786__,
    new_new_n2788__, new_new_n2791__, new_new_n2792__, new_new_n2794__,
    new_new_n2795__, new_new_n2796__, new_new_n2798__, new_new_n2800__,
    new_new_n2802__, new_new_n2804__, new_new_n2805__, new_new_n2806__,
    new_new_n2808__, new_new_n2810__, new_new_n2812__, new_new_n2813__,
    new_new_n2814__, new_new_n2815__, new_new_n2816__, new_new_n2817__,
    new_new_n2819__, new_new_n2820__, new_new_n2823__, new_new_n2824__,
    new_new_n2827__, new_new_n2828__, new_new_n2831__, new_new_n2832__,
    new_new_n2834__, new_new_n2835__, new_new_n2836__, new_new_n2837__,
    new_new_n2838__, new_new_n2839__, new_new_n2840__, new_new_n2841__,
    new_new_n2842__, new_new_n2843__, new_new_n2844__, new_new_n2845__,
    new_new_n2846__, new_new_n2847__, new_new_n2848__, new_new_n2849__,
    new_new_n2850__, new_new_n2851__, new_new_n2852__, new_new_n2853__,
    new_new_n2854__, new_new_n2855__, new_new_n2856__, new_new_n2857__,
    new_new_n2858__, new_new_n2859__, new_new_n2860__, new_new_n2861__,
    new_new_n2862__, new_new_n2863__, new_new_n2864__, new_new_n2865__,
    new_new_n2866__, new_new_n2867__, new_new_n2868__, new_new_n2869__,
    new_new_n2870__, new_new_n2871__, new_new_n2872__, new_new_n2873__,
    new_new_n2874__, new_new_n2875__, new_new_n2876__, new_new_n2877__,
    new_new_n2878__, new_new_n2879__, new_new_n2880__, new_new_n2881__,
    new_new_n2882__, new_new_n2883__, new_new_n2884__, new_new_n2885__,
    new_new_n2886__, new_new_n2887__, new_new_n2888__, new_new_n2889__,
    new_new_n2890__, new_new_n2891__, new_new_n2892__, new_new_n2893__,
    new_new_n2894__, new_new_n2895__, new_new_n2896__, new_new_n2897__,
    new_new_n2898__, new_new_n2899__, new_new_n2900__, new_new_n2901__,
    new_new_n2902__, new_new_n2903__, new_new_n2904__, new_new_n2905__,
    new_new_n2906__, new_new_n2907__, new_new_n2908__, new_new_n2909__,
    new_new_n2910__, new_new_n2911__, new_new_n2912__, new_new_n2913__,
    new_new_n2914__, new_new_n2915__, new_new_n2916__, new_new_n2917__,
    new_new_n2918__, new_new_n2919__, new_new_n2920__, new_new_n2921__,
    new_new_n2922__, new_new_n2923__, new_new_n2924__, new_new_n2925__,
    new_new_n2926__, new_new_n2927__, new_new_n2928__, new_new_n2929__,
    new_new_n2930__, new_new_n2931__, new_new_n2932__, new_new_n2933__,
    new_new_n2934__, new_new_n2935__, new_new_n2936__, new_new_n2937__,
    new_new_n2938__, new_new_n2939__, new_new_n2940__, new_new_n2941__,
    new_new_n2942__, new_new_n2943__, new_new_n2944__, new_new_n2945__,
    new_new_n2946__, new_new_n2947__, new_new_n2948__, new_new_n2949__,
    new_new_n2950__, new_new_n2951__, new_new_n2952__, new_new_n2953__,
    new_new_n2954__, new_new_n2955__, new_new_n2956__, new_new_n2957__,
    new_new_n2958__, new_new_n2959__, new_new_n2960__, new_new_n2961__,
    new_new_n2962__, new_new_n2963__, new_new_n2964__, new_new_n2965__,
    new_new_n2966__, new_new_n2967__, new_new_n2968__, new_new_n2969__,
    new_new_n2970__, new_new_n2971__, new_new_n2972__, new_new_n2973__,
    new_new_n2974__, new_new_n2975__, new_new_n2976__, new_new_n2977__,
    new_new_n2978__, new_new_n2979__, new_new_n2980__, new_new_n2981__,
    new_new_n2982__, new_new_n2983__, new_new_n2984__, new_new_n2985__,
    new_new_n2986__, new_new_n2987__, new_new_n2988__, new_new_n2989__,
    new_new_n2990__, new_new_n2991__, new_new_n2992__, new_new_n2993__,
    new_new_n2994__, new_new_n2995__, new_new_n2996__, new_new_n2997__,
    new_new_n2998__, new_new_n2999__, new_new_n3000__, new_new_n3001__,
    new_new_n3002__, new_new_n3003__, new_new_n3004__, new_new_n3005__,
    new_new_n3006__, new_new_n3007__, new_new_n3008__, new_new_n3009__,
    new_new_n3010__, new_new_n3011__, new_new_n3012__, new_new_n3013__,
    new_new_n3014__, new_new_n3015__, new_new_n3016__, new_new_n3017__,
    new_new_n3018__, new_new_n3019__, new_new_n3020__, new_new_n3021__,
    new_new_n3022__, new_new_n3023__, new_new_n3024__, new_new_n3025__,
    new_new_n3026__, new_new_n3027__, new_new_n3028__, new_new_n3029__,
    new_new_n3030__, new_new_n3031__, new_new_n3032__, new_new_n3033__,
    new_new_n3034__, new_new_n3035__, new_new_n3036__, new_new_n3037__,
    new_new_n3038__, new_new_n3039__, new_new_n3040__, new_new_n3041__,
    new_new_n3042__, new_new_n3043__, new_new_n3044__, new_new_n3045__,
    new_new_n3046__, new_new_n3047__, new_new_n3048__, new_new_n3049__,
    new_new_n3050__, new_new_n3051__, new_new_n3052__, new_new_n3053__,
    new_new_n3054__, new_new_n3055__, new_new_n3056__, new_new_n3057__,
    new_new_n3058__, new_new_n3059__, new_new_n3060__, new_new_n3061__,
    new_new_n3062__, new_new_n3063__, new_new_n3064__, new_new_n3065__,
    new_new_n3066__, new_new_n3067__, new_new_n3068__, new_new_n3069__,
    new_new_n3070__, new_new_n3071__, new_new_n3072__, new_new_n3073__,
    new_new_n3074__, new_new_n3075__, new_new_n3076__, new_new_n3077__,
    new_new_n3078__, new_new_n3079__, new_new_n3080__, new_new_n3081__,
    new_new_n3082__, new_new_n3083__, new_new_n3084__, new_new_n3085__,
    new_new_n3086__, new_new_n3087__, new_new_n3088__, new_new_n3089__,
    new_new_n3090__, new_new_n3091__, new_new_n3092__, new_new_n3093__,
    new_new_n3094__, new_new_n3095__, new_new_n3096__, new_new_n3097__,
    new_new_n3098__, new_new_n3099__, new_new_n3100__, new_new_n3101__,
    new_new_n3102__, new_new_n3103__, new_new_n3104__, new_new_n3105__,
    new_new_n3106__, new_new_n3107__, new_new_n3108__, new_new_n3109__,
    new_new_n3110__, new_new_n3111__, new_new_n3112__, new_new_n3113__,
    new_new_n3114__, new_new_n3115__, new_new_n3116__, new_new_n3117__,
    new_new_n3118__, new_new_n3119__, new_new_n3120__, new_new_n3121__,
    new_new_n3122__, new_new_n3123__, new_new_n3124__, new_new_n3125__,
    new_new_n3126__, new_new_n3127__, new_new_n3128__, new_new_n3129__,
    new_new_n3130__, new_new_n3131__, new_new_n3132__, new_new_n3133__,
    new_new_n3134__, new_new_n3135__, new_new_n3136__, new_new_n3137__,
    new_new_n3138__, new_new_n3139__, new_new_n3140__, new_new_n3141__,
    new_new_n3142__, new_new_n3143__, new_new_n3144__, new_new_n3145__,
    new_new_n3146__, new_new_n3147__, new_new_n3148__, new_new_n3149__,
    new_new_n3150__, new_new_n3151__, new_new_n3152__, new_new_n3153__,
    new_new_n3154__, new_new_n3155__, new_new_n3156__, new_new_n3157__,
    new_new_n3158__, new_new_n3159__, new_new_n3160__, new_new_n3161__,
    new_new_n3162__, new_new_n3163__, new_new_n3164__, new_new_n3165__,
    new_new_n3166__, new_new_n3167__, new_new_n3168__, new_new_n3169__,
    new_new_n3170__, new_new_n3171__, new_new_n3172__, new_new_n3173__,
    new_new_n3174__, new_new_n3175__, new_new_n3176__, new_new_n3177__,
    new_new_n3178__, new_new_n3179__, new_new_n3180__, new_new_n3181__,
    new_new_n3182__, new_new_n3183__, new_new_n3184__, new_new_n3185__,
    new_new_n3186__, new_new_n3187__, new_new_n3188__, new_new_n3189__,
    new_new_n3190__, new_new_n3191__, new_new_n3192__, new_new_n3193__,
    new_new_n3194__, new_new_n3195__, new_new_n3196__, new_new_n3197__,
    new_new_n3198__, new_new_n3199__, new_new_n3200__, new_new_n3201__,
    new_new_n3202__, new_new_n3203__, new_new_n3204__, new_new_n3205__,
    new_new_n3206__, new_new_n3207__, new_new_n3208__, new_new_n3209__,
    new_new_n3210__, new_new_n3211__, new_new_n3212__, new_new_n3213__,
    new_new_n3214__, new_new_n3215__, new_new_n3216__, new_new_n3217__,
    new_new_n3218__, new_new_n3219__, new_new_n3220__, new_new_n3221__,
    new_new_n3222__, new_new_n3223__, new_new_n3224__, new_new_n3225__,
    new_new_n3226__, new_new_n3227__, new_new_n3228__, new_new_n3229__,
    new_new_n3230__, new_new_n3231__, new_new_n3232__, new_new_n3233__,
    new_new_n3234__, new_new_n3235__, new_new_n3236__, new_new_n3237__,
    new_new_n3238__, new_new_n3239__, new_new_n3240__, new_new_n3241__,
    new_new_n3242__, new_new_n3243__, new_new_n3244__, new_new_n3245__,
    new_new_n3246__, new_new_n3247__, new_new_n3248__, new_new_n3249__,
    new_new_n3250__, new_new_n3251__, new_new_n3252__, new_new_n3253__,
    new_new_n3254__, new_new_n3255__, new_new_n3256__, new_new_n3257__,
    new_new_n3258__, new_new_n3259__, new_new_n3260__, new_new_n3261__,
    new_new_n3262__, new_new_n3263__, new_new_n3264__, new_new_n3265__,
    new_new_n3266__, new_new_n3267__, new_new_n3268__, new_new_n3269__,
    new_new_n3270__, new_new_n3271__, new_new_n3272__, new_new_n3273__,
    new_new_n3274__, new_new_n3275__, new_new_n3276__, new_new_n3277__,
    new_new_n3278__, new_new_n3279__, new_new_n3280__, new_new_n3281__,
    new_new_n3282__, new_new_n3283__, new_new_n3284__, new_new_n3285__,
    new_new_n3286__, new_new_n3287__, new_new_n3288__, new_new_n3289__,
    new_new_n3290__, new_new_n3291__, new_new_n3292__, new_new_n3293__,
    new_new_n3294__, new_new_n3295__, new_new_n3296__, new_new_n3297__,
    new_new_n3298__, new_new_n3299__, new_new_n3300__, new_new_n3301__,
    new_new_n3302__, new_new_n3303__, new_new_n3304__, new_new_n3305__,
    new_new_n3306__, new_new_n3307__, new_new_n3308__, new_new_n3309__,
    new_new_n3310__, new_new_n3311__, new_new_n3312__, new_new_n3313__,
    new_new_n3314__, new_new_n3315__, new_new_n3316__, new_new_n3317__,
    new_new_n3318__, new_new_n3319__, new_new_n3320__, new_new_n3321__,
    new_new_n3322__, new_new_n3323__, new_new_n3324__, new_new_n3325__,
    new_new_n3326__, new_new_n3327__, new_new_n3328__, new_new_n3329__,
    new_new_n3330__, new_new_n3331__, new_new_n3332__, new_new_n3333__,
    new_new_n3334__, new_new_n3335__, new_new_n3336__, new_new_n3337__,
    new_new_n3338__, new_new_n3339__, new_new_n3340__, new_new_n3341__,
    new_new_n3342__, new_new_n3343__, new_new_n3344__, new_new_n3345__,
    new_new_n3346__, new_new_n3347__, new_new_n3348__, new_new_n3349__,
    new_new_n3350__, new_new_n3351__, new_new_n3352__, new_new_n3353__,
    new_new_n3354__, new_new_n3355__, new_new_n3356__, new_new_n3357__,
    new_new_n3358__, new_new_n3359__, new_new_n3360__, new_new_n3361__,
    new_new_n3362__, new_new_n3363__, new_new_n3364__, new_new_n3365__,
    new_new_n3366__, new_new_n3367__, new_new_n3368__, new_new_n3369__,
    new_new_n3370__, new_new_n3371__, new_new_n3372__, new_new_n3373__,
    new_new_n3374__, new_new_n3375__, new_new_n3376__, new_new_n3377__,
    new_new_n3378__, new_new_n3379__, new_new_n3380__, new_new_n3381__,
    new_new_n3382__, new_new_n3383__, new_new_n3384__, new_new_n3385__,
    new_new_n3386__, new_new_n3387__, new_new_n3388__, new_new_n3389__,
    new_new_n3390__, new_new_n3391__, new_new_n3392__, new_new_n3393__,
    new_new_n3394__, new_new_n3395__, new_new_n3396__, new_new_n3397__,
    new_new_n3398__, new_new_n3399__, new_new_n3400__, new_new_n3401__,
    new_new_n3402__, new_new_n3403__, new_new_n3404__, new_new_n3405__,
    new_new_n3406__, new_new_n3407__, new_new_n3408__, new_new_n3409__,
    new_new_n3410__, new_new_n3411__, new_new_n3412__, new_new_n3413__,
    new_new_n3414__, new_new_n3415__, new_new_n3416__, new_new_n3417__,
    new_new_n3418__, new_new_n3419__, new_new_n3420__, new_new_n3421__,
    new_new_n3422__, new_new_n3423__, new_new_n3424__, new_new_n3425__,
    new_new_n3426__, new_new_n3427__, new_new_n3428__, new_new_n3429__,
    new_new_n3430__, new_new_n3431__, new_new_n3432__, new_new_n3433__,
    new_new_n3434__, new_new_n3435__, new_new_n3436__, new_new_n3437__,
    new_new_n3438__, new_new_n3439__, new_new_n3440__, new_new_n3441__,
    new_new_n3442__, new_new_n3443__, new_new_n3444__, new_new_n3445__,
    new_new_n3446__, new_new_n3447__, new_new_n3448__, new_new_n3449__,
    new_new_n3450__, new_new_n3451__, new_new_n3452__, new_new_n3453__,
    new_new_n3454__, new_new_n3455__, new_new_n3456__, new_new_n3457__,
    new_new_n3458__, new_new_n3459__, new_new_n3460__, new_new_n3461__,
    new_new_n3462__, new_new_n3463__, new_new_n3464__, new_new_n3465__,
    new_new_n3466__, new_new_n3467__, new_new_n3468__, new_new_n3469__,
    new_new_n3470__, new_new_n3471__, new_new_n3472__, new_new_n3473__,
    new_new_n3474__, new_new_n3475__, new_new_n3476__, new_new_n3477__,
    new_new_n3478__, new_new_n3479__, new_new_n3480__, new_new_n3481__,
    new_new_n3482__, new_new_n3483__, new_new_n3484__, new_new_n3485__,
    new_new_n3486__, new_new_n3487__, new_new_n3488__, new_new_n3489__,
    new_new_n3490__, new_new_n3491__, new_new_n3492__, new_new_n3493__,
    new_new_n3494__, new_new_n3495__, new_new_n3496__, new_new_n3497__,
    new_new_n3498__, new_new_n3499__, new_new_n3500__, new_new_n3501__,
    new_new_n3502__, new_new_n3503__, new_new_n3504__, new_new_n3505__,
    new_new_n3506__, new_new_n3507__, new_new_n3508__, new_new_n3509__,
    new_new_n3510__, new_new_n3511__, new_new_n3512__, new_new_n3513__,
    new_new_n3514__, new_new_n3515__, new_new_n3516__, new_new_n3517__,
    new_new_n3518__, new_new_n3519__, new_new_n3520__, new_new_n3521__,
    new_new_n4161__, new_new_n4162__, new_new_n4163__, new_new_n4164__,
    new_new_n4165__, new_new_n4166__, new_new_n4167__, new_new_n4168__,
    new_new_n4169__, new_new_n4170__, new_new_n4171__, new_new_n4172__,
    new_new_n4173__, new_new_n4174__, new_new_n4175__, new_new_n4176__,
    new_new_n4177__, new_new_n4178__, new_new_n4179__, new_new_n4180__,
    new_new_n4181__, new_new_n4182__, new_new_n4183__, new_new_n4184__,
    new_new_n4185__, new_new_n4186__, new_new_n4187__, new_new_n4188__,
    new_new_n4189__, new_new_n4190__, new_new_n4191__, new_new_n4192__,
    new_new_n4193__, new_new_n4194__, new_new_n4195__, new_new_n4196__,
    new_new_n4197__, new_new_n4198__, new_new_n4199__, new_new_n4200__,
    new_new_n4201__, new_new_n4202__, new_new_n4203__, new_new_n4204__,
    new_new_n4205__, new_new_n4206__, new_new_n4207__, new_new_n4208__,
    new_new_n4209__, new_new_n4210__, new_new_n4211__, new_new_n4212__,
    new_new_n4213__, new_new_n4214__, new_new_n4215__, new_new_n4216__,
    new_new_n4217__, new_new_n4218__, new_new_n4219__, new_new_n4220__,
    new_new_n4221__, new_new_n4222__, new_new_n4223__, new_new_n4224__,
    new_new_n4225__, new_new_n4226__, new_new_n4227__, new_new_n4228__,
    new_new_n4229__, new_new_n4230__, new_new_n4231__, new_new_n4232__,
    new_new_n4233__, new_new_n4234__, new_new_n4235__, new_new_n4236__,
    new_new_n4237__, new_new_n4238__, new_new_n4239__, new_new_n4240__,
    new_new_n4241__, new_new_n4242__, new_new_n4243__, new_new_n4244__,
    new_new_n4245__, new_new_n4246__, new_new_n4247__, new_new_n4248__,
    new_new_n4249__, new_new_n4250__, new_new_n4251__, new_new_n4252__,
    new_new_n4253__, new_new_n4254__, new_new_n4255__, new_new_n4256__,
    new_new_n4257__, new_new_n4258__, new_new_n4259__, new_new_n4260__,
    new_new_n4261__, new_new_n4262__, new_new_n4263__, new_new_n4264__,
    new_new_n4265__, new_new_n4266__, new_new_n4267__, new_new_n4268__,
    new_new_n4269__, new_new_n4270__, new_new_n4271__, new_new_n4272__,
    new_new_n4273__, new_new_n4274__, new_new_n4275__, new_new_n4276__,
    new_new_n4277__, new_new_n4278__, new_new_n4279__, new_new_n4280__,
    new_new_n4281__, new_new_n4282__, new_new_n4283__, new_new_n4284__,
    new_new_n4285__, new_new_n4286__, new_new_n4287__, new_new_n4288__,
    new_new_n4289__, new_new_n4290__, new_new_n4291__, new_new_n4292__,
    new_new_n4293__, new_new_n4294__, new_new_n4295__, new_new_n4296__,
    new_new_n4297__, new_new_n4298__, new_new_n4299__, new_new_n4300__,
    new_new_n4301__, new_new_n4302__, new_new_n4303__, new_new_n4304__,
    new_new_n4305__, new_new_n4306__, new_new_n4307__, new_new_n4308__,
    new_new_n4309__, new_new_n4310__, new_new_n4311__, new_new_n4312__,
    new_new_n4313__, new_new_n4314__, new_new_n4315__, new_new_n4316__,
    new_new_n4317__, new_new_n4318__, new_new_n4319__, new_new_n4320__,
    new_new_n4321__, new_new_n4322__, new_new_n4323__, new_new_n4324__,
    new_new_n4325__, new_new_n4326__, new_new_n4327__, new_new_n4328__,
    new_new_n4329__, new_new_n4330__, new_new_n4331__, new_new_n4332__,
    new_new_n4333__, new_new_n4334__, new_new_n4335__, new_new_n4336__,
    new_new_n4337__, new_new_n4338__, new_new_n4339__, new_new_n4340__,
    new_new_n4341__, new_new_n4342__, new_new_n4343__, new_new_n4344__,
    new_new_n4345__, new_new_n4346__, new_new_n4347__, new_new_n4348__,
    new_new_n4349__, new_new_n4350__, new_new_n4351__, new_new_n4352__,
    new_new_n4353__, new_new_n4354__, new_new_n4355__, new_new_n4356__,
    new_new_n4357__, new_new_n4358__, new_new_n4359__, new_new_n4360__,
    new_new_n4361__, new_new_n4362__, new_new_n4363__, new_new_n4364__,
    new_new_n4365__, new_new_n4366__, new_new_n4367__, new_new_n4368__,
    new_new_n4369__, new_new_n4370__, new_new_n4371__, new_new_n4372__,
    new_new_n4373__, new_new_n4374__, new_new_n4375__, new_new_n4376__,
    new_new_n4377__, new_new_n4378__, new_new_n4379__, new_new_n4380__,
    new_new_n4381__, new_new_n4382__, new_new_n4383__, new_new_n4384__,
    new_new_n4385__, new_new_n4386__, new_new_n4387__, new_new_n4388__,
    new_new_n4389__, new_new_n4390__, new_new_n4391__, new_new_n4392__,
    new_new_n4393__, new_new_n4394__, new_new_n4395__, new_new_n4396__,
    new_new_n4397__, new_new_n4398__, new_new_n4399__, new_new_n4400__,
    new_new_n4401__, new_new_n4402__, new_new_n4403__, new_new_n4404__,
    new_new_n4405__, new_new_n4406__, new_new_n4407__, new_new_n4408__,
    new_new_n4409__, new_new_n4410__, new_new_n4411__, new_new_n4412__,
    new_new_n4413__, new_new_n4414__, new_new_n4415__, new_new_n4416__,
    new_new_n4417__, new_new_n4418__, new_new_n4419__, new_new_n4420__,
    new_new_n4421__, new_new_n4422__, new_new_n4423__, new_new_n4424__,
    new_new_n4425__, new_new_n4426__, new_new_n4427__, new_new_n4428__,
    new_new_n4429__, new_new_n4430__, new_new_n4431__, new_new_n4432__,
    new_new_n4433__, new_new_n4434__, new_new_n4435__, new_new_n4436__,
    new_new_n4437__, new_new_n4438__, new_new_n4439__, new_new_n4440__,
    new_new_n4441__, new_new_n4442__, new_new_n4443__, new_new_n4444__,
    new_new_n4445__, new_new_n4446__, new_new_n4447__, new_new_n4448__,
    new_new_n4449__, new_new_n4450__, new_new_n4451__, new_new_n4452__,
    new_new_n4453__, new_new_n4454__, new_new_n4455__, new_new_n4456__,
    new_new_n4457__, new_new_n4458__, new_new_n4459__, new_new_n4460__,
    new_new_n4461__, new_new_n4462__, new_new_n4463__, new_new_n4464__,
    new_new_n4465__, new_new_n4466__, new_new_n4467__, new_new_n4468__,
    new_new_n4469__, new_new_n4470__, new_new_n4471__, new_new_n4472__,
    new_new_n4473__, new_new_n4474__, new_new_n4475__, new_new_n4476__,
    new_new_n4477__, new_new_n4478__, new_new_n4479__, new_new_n4480__,
    new_new_n4481__, new_new_n4482__, new_new_n4483__, new_new_n4484__,
    new_new_n4485__, new_new_n4486__, new_new_n4487__, new_new_n4488__,
    new_new_n4489__, new_new_n4490__, new_new_n4491__, new_new_n4492__,
    new_new_n4493__, new_new_n4494__, new_new_n4495__, new_new_n4496__,
    new_new_n4497__, new_new_n4498__, new_new_n4499__, new_new_n4500__,
    new_new_n4501__, new_new_n4502__, new_new_n4503__, new_new_n4504__,
    new_new_n4505__, new_new_n4506__, new_new_n4507__, new_new_n4508__,
    new_new_n4509__, new_new_n4510__, new_new_n4511__, new_new_n4512__,
    new_new_n4513__, new_new_n4514__, new_new_n4515__, new_new_n4516__,
    new_new_n4517__, new_new_n4518__, new_new_n4519__, new_new_n4520__,
    new_new_n4521__, new_new_n4522__, new_new_n4523__, new_new_n4524__,
    new_new_n4525__, new_new_n4526__, new_new_n4527__, new_new_n4528__,
    new_new_n4529__, new_new_n4530__, new_new_n4531__, new_new_n4532__,
    new_new_n4533__, new_new_n4534__, new_new_n4535__, new_new_n4536__,
    new_new_n4537__, new_new_n4538__, new_new_n4539__, new_new_n4540__,
    new_new_n4541__, new_new_n4542__, new_new_n4543__, new_new_n4544__,
    new_new_n4545__, new_new_n4546__, new_new_n4547__, new_new_n4548__,
    new_new_n4549__, new_new_n4550__, new_new_n4551__, new_new_n4552__,
    new_new_n4553__, new_new_n4554__, new_new_n4555__, new_new_n4556__,
    new_new_n4557__, new_new_n4558__, new_new_n4559__, new_new_n4560__,
    new_new_n4561__, new_new_n4562__, new_new_n4563__, new_new_n4564__,
    new_new_n4565__, new_new_n4566__, new_new_n4567__, new_new_n4568__,
    new_new_n4569__, new_new_n4570__, new_new_n4571__, new_new_n4572__,
    new_new_n4573__, new_new_n4574__, new_new_n4575__, new_new_n4576__,
    new_new_n4577__, new_new_n4578__, new_new_n4579__, new_new_n4580__,
    new_new_n4581__, new_new_n4582__, new_new_n4583__, new_new_n4584__,
    new_new_n4585__, new_new_n4586__, new_new_n4587__, new_new_n4588__,
    new_new_n4589__, new_new_n4590__, new_new_n4591__, new_new_n4592__,
    new_new_n4593__, new_new_n4594__, new_new_n4595__, new_new_n4596__,
    new_new_n4597__, new_new_n4598__, new_new_n4599__, new_new_n4600__,
    new_new_n4601__, new_new_n4602__, new_new_n4603__, new_new_n4604__,
    new_new_n4605__, new_new_n4606__, new_new_n4607__, new_new_n4608__,
    new_new_n4609__, new_new_n4610__, new_new_n4611__, new_new_n4612__,
    new_new_n4613__, new_new_n4614__, new_new_n4615__, n6254, n6257, n6260,
    n6263, n6266, n6269, n6272, n6275, n6278, n6281, n6284, n6287, n6290,
    n6293, n6296, n6299, n6302, n6305, n6308, n6311, n6314, n6317, n6320,
    n6323, n6326, n6329, n6332, n6335, n6338, n6341, n6344, n6347, n6350,
    n6353, n6356, n6359, n6362, n6365, n6368, n6371, n6374, n6377, n6380,
    n6383, n6386, n6389, n6392, n6395, n6398, n6401, n6404, n6407, n6410,
    n6413, n6416, n6419, n6422, n6425, n6428, n6431, n6434, n6437, n6440,
    n6443, n6446, n6449, n6452, n6455, n6458, n6461, n6464, n6467, n6470,
    n6473, n6476, n6479, n6482, n6485, n6488, n6491, n6494, n6497, n6500,
    n6503, n6506, n6509, n6512, n6515, n6518, n6521, n6524, n6527, n6530,
    n6533, n6536, n6539, n6542, n6545, n6548, n6551, n6554, n6557, n6560,
    n6563, n6566, n6569, n6572, n6575, n6578, n6581, n6584, n6587, n6590,
    n6593, n6596, n6599, n6602, n6605, n6608, n6611, n6614, n6617, n6620,
    n6623, n6626, n6629, n6632, n6635, n6638, n6641, n6644, n6647, n6650,
    n6653, n6656, n6659, n6662, n6665, n6668, n6671, n6674, n6677, n6680,
    n6683, n6686, n6689, n6692, n6695, n6698, n6701, n6704, n6707, n6710,
    n6713, n6716, n6719, n6722, n6725, n6728, n6731, n6734, n6737, n6740,
    n6743, n6746, n6749, n6752, n6755, n6758, n6761, n6764, n6767, n6770,
    n6773, n6776, n6779, n6782, n6785, n6788, n6791, n6794, n6797, n6800,
    n6803, n6806, n6809, n6812, n6815, n6818, n6821, n6824, n6827, n6830,
    n6833, n6836, n6839, n6842, n6845, n6848, n6851, n6854, n6857, n6860,
    n6863, n6866, n6869, n6872, n6875, n6878, n6881, n6884, n6887, n6890,
    n6893, n6896, n6899, n6902, n6905, n6908, n6911, n6914, n6917, n6920,
    n6923, n6926, n6929, n6932, n6935, n6938, n6941, n6944, n6947, n6950,
    n6953, n6956, n6959, n6962, n6965, n6968, n6971, n6974, n6977, n6980,
    n6983, n6986, n6989, n6992, n6995, n6998, n7001, n7004, n7007, n7010,
    n7013, n7016, n7019, n7022, n7025, n7028, n7031, n7034, n7037, n7040,
    n7043, n7046, n7049, n7052, n7055, n7058, n7061, n7064, n7067, n7070,
    n7073, n7076, n7079, n7082, n7085, n7088, n7091, n7094, n7097, n7100,
    n7103, n7106, n7109, n7112, n7115, n7118, n7121, n7124, n7127, n7130,
    n7133, n7136, n7139, n7142, n7145, n7148, n7151, n7154, n7157, n7160,
    n7163, n7166, n7169, n7172, n7175, n7178, n7181, n7184, n7187, n7190,
    n7193, n7196, n7199, n7202, n7205, n7208, n7211, n7214, n7217, n7220,
    n7223, n7226, n7229, n7232, n7235, n7238, n7241, n7244, n7247, n7250,
    n7253, n7256, n7259, n7262, n7265, n7268, n7271, n7274, n7277, n7280,
    n7283, n7286, n7289, n7292, n7295, n7298, n7301, n7304, n7307, n7310,
    n7313, n7316, n7319, n7322, n7325, n7328, n7331, n7334, n7337, n7340,
    n7343, n7346, n7349, n7352, n7355, n7358, n7361, n7364, n7367, n7370,
    n7373, n7376, n7379, n7382, n7385, n7388, n7391, n7394, n7397, n7400,
    n7403, n7406, n7409, n7412, n7415, n7418, n7421, n7424, n7427, n7430,
    n7433, n7436, n7439, n7442, n7445, n7448, n7451, n7454, n7457, n7460,
    n7463, n7466, n7469, n7472, n7475, n7478, n7481, n7484, n7487, n7490,
    n7493, n7496, n7499, n7502, n7505, n7508, n7511, n7514, n7517, n7520,
    n7523, n7526, n7529, n7532, n7535, n7538, n7541, n7544, n7547, n7550,
    n7553, n7556, n7559, n7562, n7565, n7568, n7571, n7574, n7577, n7580,
    n7583, n7586, n7589, n7592, n7595, n7598, n7601, n7604, n7607, n7610,
    n7613, n7616, n7619, n7622, n7625, n7628, n7631, n7634, n7637, n7640,
    n7643, n7646, n7649, n7652, n7655, n7658, n7661, n7664, n7667, n7670,
    n7673, n7676, n7679, n7682, n7685, n7688, n7691, n7694, n7697, n7700,
    n7703, n7706, n7709, n7712, n7715, n7718, n7721, n7724, n7727, n7730,
    n7733, n7736, n7739, n7742, n7745, n7748, n7751, n7754, n7757, n7760,
    n7763, n7766, n7769, n7772, n7775, n7778, n7781, n7784, n7787, n7790,
    n7793, n7796, n7799, n7802, n7805, n7808, n7811, n7814, n7817, n7820,
    n7823, n7826, n7829, n7832, n7835, n7838, n7841, n7844, n7847, n7850,
    n7853, n7856, n7859, n7862, n7865, n7868, n7871, n7874, n7877, n7880,
    n7883, n7886, n7889, n7892, n7895, n7898, n7901, n7904, n7907, n7910,
    n7913, n7916, n7919, n7922, n7925, n7928, n7931, n7934, n7937, n7940,
    n7943, n7946, n7949, n7952, n7955, n7958, n7961, n7964, n7967, n7970,
    n7973, n7976;
  buf1  g0000(.din(G1), .dout(new_new_n1372__));
  buf1  g0001(.din(G2), .dout(new_new_n1374__));
  buf1  g0002(.din(G3), .dout(new_new_n1376__));
  buf1  g0003(.din(G4), .dout(new_new_n1378__));
  buf1  g0004(.din(G5), .dout(new_new_n1380__));
  buf1  g0005(.din(G6), .dout(new_new_n1382__));
  buf1  g0006(.din(G7), .dout(new_new_n1384__));
  buf1  g0007(.din(G8), .dout(new_new_n1386__));
  buf1  g0008(.din(G9), .dout(new_new_n1388__));
  buf1  g0009(.din(G10), .dout(new_new_n1390__));
  buf1  g0010(.din(G11), .dout(new_new_n1392__));
  buf1  g0011(.din(G12), .dout(new_new_n1394__));
  buf1  g0012(.din(G13), .dout(new_new_n1396__));
  buf1  g0013(.din(G14), .dout(new_new_n1398__));
  buf1  g0014(.din(G15), .dout(new_new_n1400__));
  buf1  g0015(.din(G16), .dout(new_new_n1402__));
  buf1  g0016(.din(G17), .dout(new_new_n1404__));
  buf1  g0017(.din(G18), .dout(new_new_n1406__));
  buf1  g0018(.din(G19), .dout(new_new_n1408__));
  buf1  g0019(.din(G20), .dout(new_new_n1410__));
  buf1  g0020(.din(G21), .dout(new_new_n1412__));
  buf1  g0021(.din(G22), .dout(new_new_n1414__));
  buf1  g0022(.din(G23), .dout(new_new_n1416__));
  buf1  g0023(.din(G24), .dout(new_new_n1418__));
  buf1  g0024(.din(G25), .dout(new_new_n1420__));
  buf1  g0025(.din(G26), .dout(new_new_n1422__));
  buf1  g0026(.din(G27), .dout(new_new_n1424__));
  buf1  g0027(.din(G28), .dout(new_new_n1426__));
  buf1  g0028(.din(G29), .dout(new_new_n1428__));
  buf1  g0029(.din(G30), .dout(new_new_n1430__));
  buf1  g0030(.din(G31), .dout(new_new_n1432__));
  buf1  g0031(.din(G32), .dout(new_new_n1434__));
  buf1  g0032(.din(G33), .dout(new_new_n1436__));
  buf1  g0033(.din(G34), .dout(new_new_n1438__));
  buf1  g0034(.din(G35), .dout(new_new_n1440__));
  buf1  g0035(.din(G36), .dout(new_new_n1442__));
  buf1  g0036(.din(G37), .dout(new_new_n1444__));
  buf1  g0037(.din(G38), .dout(new_new_n1446__));
  buf1  g0038(.din(G39), .dout(new_new_n1448__));
  buf1  g0039(.din(G40), .dout(new_new_n1450__));
  buf1  g0040(.din(G41), .dout(new_new_n1452__));
  buf1  g0041(.din(G42), .dout(new_new_n1454__));
  buf1  g0042(.din(G43), .dout(new_new_n1456__));
  buf1  g0043(.din(G44), .dout(new_new_n1458__));
  buf1  g0044(.din(G45), .dout(new_new_n1460__));
  buf1  g0045(.din(G46), .dout(new_new_n1462__));
  buf1  g0046(.din(G47), .dout(new_new_n1464__));
  buf1  g0047(.din(G48), .dout(new_new_n1466__));
  buf1  g0048(.din(G49), .dout(new_new_n1468__));
  buf1  g0049(.din(G50), .dout(new_new_n1470__));
  buf1  g0050(.din(G51), .dout(new_new_n1472__));
  buf1  g0051(.din(G52), .dout(new_new_n1474__));
  buf1  g0052(.din(G53), .dout(new_new_n1476__));
  buf1  g0053(.din(G54), .dout(new_new_n1478__));
  buf1  g0054(.din(G55), .dout(new_new_n1480__));
  buf1  g0055(.din(G56), .dout(new_new_n1482__));
  buf1  g0056(.din(G57), .dout(new_new_n1484__));
  buf1  g0057(.din(G58), .dout(new_new_n1486__));
  buf1  g0058(.din(G59), .dout(new_new_n1488__));
  buf1  g0059(.din(G60), .dout(new_new_n1490__));
  buf1  g0060(.din(G61), .dout(new_new_n1492__));
  buf1  g0061(.din(G62), .dout(new_new_n1494__));
  buf1  g0062(.din(G63), .dout(new_new_n1496__));
  buf1  g0063(.din(G64), .dout(new_new_n1498__));
  buf1  g0064(.din(G65), .dout(new_new_n1500__));
  buf1  g0065(.din(G66), .dout(new_new_n1502__));
  buf1  g0066(.din(G67), .dout(new_new_n1504__));
  buf1  g0067(.din(G68), .dout(new_new_n1506__));
  buf1  g0068(.din(G69), .dout(new_new_n1508__));
  buf1  g0069(.din(G70), .dout(new_new_n1510__));
  buf1  g0070(.din(G71), .dout(new_new_n1512__));
  buf1  g0071(.din(G72), .dout(new_new_n1514__));
  buf1  g0072(.din(G73), .dout(new_new_n1516__));
  buf1  g0073(.din(G74), .dout(new_new_n1518__));
  buf1  g0074(.din(G75), .dout(new_new_n1520__));
  buf1  g0075(.din(G76), .dout(new_new_n1522__));
  buf1  g0076(.din(G77), .dout(new_new_n1524__));
  buf1  g0077(.din(G78), .dout(new_new_n1526__));
  buf1  g0078(.din(G79), .dout(new_new_n1528__));
  buf1  g0079(.din(G80), .dout(new_new_n1530__));
  buf1  g0080(.din(G81), .dout(new_new_n1532__));
  buf1  g0081(.din(G82), .dout(new_new_n1534__));
  buf1  g0082(.din(G83), .dout(new_new_n1536__));
  buf1  g0083(.din(G84), .dout(new_new_n1538__));
  buf1  g0084(.din(G85), .dout(new_new_n1540__));
  buf1  g0085(.din(G86), .dout(new_new_n1542__));
  buf1  g0086(.din(G87), .dout(new_new_n1544__));
  buf1  g0087(.din(G88), .dout(new_new_n1546__));
  buf1  g0088(.din(G89), .dout(new_new_n1548__));
  buf1  g0089(.din(G90), .dout(new_new_n1550__));
  buf1  g0090(.din(G91), .dout(new_new_n1552__));
  buf1  g0091(.din(G92), .dout(new_new_n1554__));
  buf1  g0092(.din(G93), .dout(new_new_n1556__));
  buf1  g0093(.din(G94), .dout(new_new_n1558__));
  buf1  g0094(.din(G95), .dout(new_new_n1560__));
  buf1  g0095(.din(G96), .dout(new_new_n1562__));
  buf1  g0096(.din(G97), .dout(new_new_n1564__));
  buf1  g0097(.din(G98), .dout(new_new_n1566__));
  buf1  g0098(.din(G99), .dout(new_new_n1568__));
  buf1  g0099(.din(G100), .dout(new_new_n1570__));
  buf1  g0100(.din(G101), .dout(new_new_n1572__));
  buf1  g0101(.din(G102), .dout(new_new_n1574__));
  buf1  g0102(.din(G103), .dout(new_new_n1576__));
  buf1  g0103(.din(G104), .dout(new_new_n1578__));
  buf1  g0104(.din(G105), .dout(new_new_n1580__));
  buf1  g0105(.din(G106), .dout(new_new_n1582__));
  buf1  g0106(.din(G107), .dout(new_new_n1584__));
  buf1  g0107(.din(G108), .dout(new_new_n1586__));
  buf1  g0108(.din(G109), .dout(new_new_n1588__));
  buf1  g0109(.din(G110), .dout(new_new_n1590__));
  buf1  g0110(.din(G111), .dout(new_new_n1592__));
  buf1  g0111(.din(G112), .dout(new_new_n1594__));
  buf1  g0112(.din(G113), .dout(new_new_n1596__));
  buf1  g0113(.din(G114), .dout(new_new_n1598__));
  buf1  g0114(.din(G115), .dout(new_new_n1600__));
  buf1  g0115(.din(G116), .dout(new_new_n1602__));
  buf1  g0116(.din(G117), .dout(new_new_n1604__));
  buf1  g0117(.din(G118), .dout(new_new_n1606__));
  buf1  g0118(.din(G119), .dout(new_new_n1608__));
  buf1  g0119(.din(G120), .dout(new_new_n1610__));
  buf1  g0120(.din(G121), .dout(new_new_n1612__));
  buf1  g0121(.din(G122), .dout(new_new_n1614__));
  buf1  g0122(.din(G123), .dout(new_new_n1616__));
  buf1  g0123(.din(G124), .dout(new_new_n1618__));
  buf1  g0124(.din(G125), .dout(new_new_n1620__));
  buf1  g0125(.din(G126), .dout(new_new_n1622__));
  buf1  g0126(.din(G127), .dout(new_new_n1624__));
  buf1  g0127(.din(G128), .dout(new_new_n1626__));
  buf1  g0128(.din(G129), .dout(new_new_n1628__));
  buf1  g0129(.din(G130), .dout(new_new_n1630__));
  buf1  g0130(.din(G131), .dout(new_new_n1632__));
  buf1  g0131(.din(G132), .dout(new_new_n1634__));
  buf1  g0132(.din(G133), .dout(new_new_n1636__));
  buf1  g0133(.din(G134), .dout(new_new_n1638__));
  buf1  g0134(.din(G135), .dout(new_new_n1640__));
  buf1  g0135(.din(G136), .dout(new_new_n1642__));
  buf1  g0136(.din(G137), .dout(new_new_n1644__));
  buf1  g0137(.din(G138), .dout(new_new_n1646__));
  buf1  g0138(.din(G139), .dout(new_new_n1648__));
  buf1  g0139(.din(G140), .dout(new_new_n1650__));
  buf1  g0140(.din(G141), .dout(new_new_n1652__));
  buf1  g0141(.din(G142), .dout(new_new_n1654__));
  buf1  g0142(.din(G143), .dout(new_new_n1656__));
  buf1  g0143(.din(G144), .dout(new_new_n1658__));
  buf1  g0144(.din(G145), .dout(new_new_n1660__));
  buf1  g0145(.din(G146), .dout(new_new_n1662__));
  buf1  g0146(.din(G147), .dout(new_new_n1664__));
  buf1  g0147(.din(G148), .dout(new_new_n1666__));
  buf1  g0148(.din(G149), .dout(new_new_n1668__));
  buf1  g0149(.din(G150), .dout(new_new_n1670__));
  buf1  g0150(.din(G151), .dout(new_new_n1672__));
  buf1  g0151(.din(G152), .dout(new_new_n1674__));
  buf1  g0152(.din(G153), .dout(new_new_n1676__));
  buf1  g0153(.din(G154), .dout(new_new_n1678__));
  buf1  g0154(.din(G155), .dout(new_new_n1680__));
  buf1  g0155(.din(G156), .dout(new_new_n1682__));
  buf1  g0156(.din(G157), .dout(new_new_n1684__));
  buf1  g0157(.din(n1416_lo), .dout(new_new_n1686__));
  buf1  g0158(.din(n1419_lo), .dout(new_new_n1688__));
  buf1  g0159(.din(n1422_lo), .dout(new_new_n1690__));
  buf1  g0160(.din(n1425_lo), .dout(new_new_n1692__));
  buf1  g0161(.din(n1428_lo), .dout(new_new_n1694__));
  buf1  g0162(.din(n1431_lo), .dout(new_new_n1696__));
  buf1  g0163(.din(n1434_lo), .dout(new_new_n1698__));
  not1  g0164(.din(n1437_lo), .dout(new_new_n1701__));
  buf1  g0165(.din(n1440_lo), .dout(new_new_n1702__));
  buf1  g0166(.din(n1443_lo), .dout(new_new_n1704__));
  buf1  g0167(.din(n1446_lo), .dout(new_new_n1706__));
  buf1  g0168(.din(n1449_lo), .dout(new_new_n1708__));
  buf1  g0169(.din(n1452_lo), .dout(new_new_n1710__));
  buf1  g0170(.din(n1455_lo), .dout(new_new_n1712__));
  buf1  g0171(.din(n1458_lo), .dout(new_new_n1714__));
  buf1  g0172(.din(n1464_lo), .dout(new_new_n1716__));
  buf1  g0173(.din(n1467_lo), .dout(new_new_n1718__));
  buf1  g0174(.din(n1470_lo), .dout(new_new_n1720__));
  buf1  g0175(.din(n1476_lo), .dout(new_new_n1722__));
  buf1  g0176(.din(n1479_lo), .dout(new_new_n1724__));
  buf1  g0177(.din(n1482_lo), .dout(new_new_n1726__));
  buf1  g0178(.din(n1488_lo), .dout(new_new_n1728__));
  buf1  g0179(.din(n1491_lo), .dout(new_new_n1730__));
  buf1  g0180(.din(n1494_lo), .dout(new_new_n1732__));
  not1  g0181(.din(n1497_lo), .dout(new_new_n1735__));
  buf1  g0182(.din(n1500_lo), .dout(new_new_n1736__));
  buf1  g0183(.din(n1503_lo), .dout(new_new_n1738__));
  buf1  g0184(.din(n1512_lo), .dout(new_new_n1740__));
  buf1  g0185(.din(n1515_lo), .dout(new_new_n1742__));
  buf1  g0186(.din(n1518_lo), .dout(new_new_n1744__));
  not1  g0187(.din(n1521_lo), .dout(new_new_n1747__));
  buf1  g0188(.din(n1524_lo), .dout(new_new_n1748__));
  buf1  g0189(.din(n1527_lo), .dout(new_new_n1750__));
  buf1  g0190(.din(n1530_lo), .dout(new_new_n1752__));
  buf1  g0191(.din(n1533_lo), .dout(new_new_n1754__));
  buf1  g0192(.din(n1536_lo), .dout(new_new_n1756__));
  buf1  g0193(.din(n1539_lo), .dout(new_new_n1758__));
  buf1  g0194(.din(n1542_lo), .dout(new_new_n1760__));
  not1  g0195(.din(n1545_lo), .dout(new_new_n1763__));
  buf1  g0196(.din(n1548_lo), .dout(new_new_n1764__));
  buf1  g0197(.din(n1551_lo), .dout(new_new_n1766__));
  buf1  g0198(.din(n1554_lo), .dout(new_new_n1768__));
  not1  g0199(.din(n1554_lo), .dout(new_new_n1769__));
  buf1  g0200(.din(n1560_lo), .dout(new_new_n1770__));
  buf1  g0201(.din(n1563_lo), .dout(new_new_n1772__));
  buf1  g0202(.din(n1566_lo), .dout(new_new_n1774__));
  buf1  g0203(.din(n1572_lo), .dout(new_new_n1776__));
  buf1  g0204(.din(n1575_lo), .dout(new_new_n1778__));
  buf1  g0205(.din(n1578_lo), .dout(new_new_n1780__));
  buf1  g0206(.din(n1584_lo), .dout(new_new_n1782__));
  buf1  g0207(.din(n1587_lo), .dout(new_new_n1784__));
  buf1  g0208(.din(n1590_lo), .dout(new_new_n1786__));
  buf1  g0209(.din(n1596_lo), .dout(new_new_n1788__));
  buf1  g0210(.din(n1599_lo), .dout(new_new_n1790__));
  buf1  g0211(.din(n1602_lo), .dout(new_new_n1792__));
  buf1  g0212(.din(n1608_lo), .dout(new_new_n1794__));
  buf1  g0213(.din(n1611_lo), .dout(new_new_n1796__));
  buf1  g0214(.din(n1614_lo), .dout(new_new_n1798__));
  buf1  g0215(.din(n1620_lo), .dout(new_new_n1800__));
  buf1  g0216(.din(n1623_lo), .dout(new_new_n1802__));
  buf1  g0217(.din(n1626_lo), .dout(new_new_n1804__));
  buf1  g0218(.din(n1632_lo), .dout(new_new_n1806__));
  buf1  g0219(.din(n1635_lo), .dout(new_new_n1808__));
  buf1  g0220(.din(n1638_lo), .dout(new_new_n1810__));
  buf1  g0221(.din(n1644_lo), .dout(new_new_n1812__));
  buf1  g0222(.din(n1647_lo), .dout(new_new_n1814__));
  buf1  g0223(.din(n1650_lo), .dout(new_new_n1816__));
  buf1  g0224(.din(n1656_lo), .dout(new_new_n1818__));
  buf1  g0225(.din(n1659_lo), .dout(new_new_n1820__));
  buf1  g0226(.din(n1662_lo), .dout(new_new_n1822__));
  buf1  g0227(.din(n1668_lo), .dout(new_new_n1824__));
  buf1  g0228(.din(n1671_lo), .dout(new_new_n1826__));
  buf1  g0229(.din(n1674_lo), .dout(new_new_n1828__));
  buf1  g0230(.din(n1680_lo), .dout(new_new_n1830__));
  buf1  g0231(.din(n1683_lo), .dout(new_new_n1832__));
  buf1  g0232(.din(n1686_lo), .dout(new_new_n1834__));
  not1  g0233(.din(n1686_lo), .dout(new_new_n1835__));
  buf1  g0234(.din(n1692_lo), .dout(new_new_n1836__));
  buf1  g0235(.din(n1695_lo), .dout(new_new_n1838__));
  buf1  g0236(.din(n1698_lo), .dout(new_new_n1840__));
  buf1  g0237(.din(n1704_lo), .dout(new_new_n1842__));
  buf1  g0238(.din(n1707_lo), .dout(new_new_n1844__));
  buf1  g0239(.din(n1710_lo), .dout(new_new_n1846__));
  buf1  g0240(.din(n1716_lo), .dout(new_new_n1848__));
  buf1  g0241(.din(n1719_lo), .dout(new_new_n1850__));
  buf1  g0242(.din(n1722_lo), .dout(new_new_n1852__));
  buf1  g0243(.din(n1728_lo), .dout(new_new_n1854__));
  buf1  g0244(.din(n1731_lo), .dout(new_new_n1856__));
  buf1  g0245(.din(n1734_lo), .dout(new_new_n1858__));
  buf1  g0246(.din(n1740_lo), .dout(new_new_n1860__));
  buf1  g0247(.din(n1743_lo), .dout(new_new_n1862__));
  buf1  g0248(.din(n1746_lo), .dout(new_new_n1864__));
  not1  g0249(.din(n1749_lo), .dout(new_new_n1867__));
  buf1  g0250(.din(n1752_lo), .dout(new_new_n1868__));
  buf1  g0251(.din(n1755_lo), .dout(new_new_n1870__));
  buf1  g0252(.din(n1758_lo), .dout(new_new_n1872__));
  not1  g0253(.din(n1761_lo), .dout(new_new_n1875__));
  buf1  g0254(.din(n1764_lo), .dout(new_new_n1876__));
  buf1  g0255(.din(n1776_lo), .dout(new_new_n1878__));
  buf1  g0256(.din(n1788_lo), .dout(new_new_n1880__));
  buf1  g0257(.din(n1791_lo), .dout(new_new_n1882__));
  buf1  g0258(.din(n1794_lo), .dout(new_new_n1884__));
  not1  g0259(.din(n1797_lo), .dout(new_new_n1887__));
  buf1  g0260(.din(n1800_lo), .dout(new_new_n1888__));
  buf1  g0261(.din(n1803_lo), .dout(new_new_n1890__));
  buf1  g0262(.din(n1812_lo), .dout(new_new_n1892__));
  buf1  g0263(.din(n1815_lo), .dout(new_new_n1894__));
  buf1  g0264(.din(n1824_lo), .dout(new_new_n1896__));
  not1  g0265(.din(n1827_lo), .dout(new_new_n1899__));
  buf1  g0266(.din(n1836_lo), .dout(new_new_n1900__));
  not1  g0267(.din(n1839_lo), .dout(new_new_n1903__));
  buf1  g0268(.din(n1848_lo), .dout(new_new_n1904__));
  not1  g0269(.din(n1851_lo), .dout(new_new_n1907__));
  buf1  g0270(.din(n1860_lo), .dout(new_new_n1908__));
  buf1  g0271(.din(n1872_lo), .dout(new_new_n1910__));
  buf1  g0272(.din(n1875_lo), .dout(new_new_n1912__));
  buf1  g0273(.din(n1884_lo), .dout(new_new_n1914__));
  buf1  g0274(.din(n1896_lo), .dout(new_new_n1916__));
  buf1  g0275(.din(n1899_lo), .dout(new_new_n1918__));
  buf1  g0276(.din(n1908_lo), .dout(new_new_n1920__));
  buf1  g0277(.din(n1920_lo), .dout(new_new_n1922__));
  buf1  g0278(.din(n1923_lo), .dout(new_new_n1924__));
  buf1  g0279(.din(n1926_lo), .dout(new_new_n1926__));
  not1  g0280(.din(n1929_lo), .dout(new_new_n1929__));
  buf1  g0281(.din(n1932_lo), .dout(new_new_n1930__));
  buf1  g0282(.din(n1935_lo), .dout(new_new_n1932__));
  buf1  g0283(.din(n1944_lo), .dout(new_new_n1934__));
  buf1  g0284(.din(n1947_lo), .dout(new_new_n1936__));
  buf1  g0285(.din(n1956_lo), .dout(new_new_n1938__));
  buf1  g0286(.din(n1959_lo), .dout(new_new_n1940__));
  buf1  g0287(.din(n1962_lo), .dout(new_new_n1942__));
  not1  g0288(.din(n1962_lo), .dout(new_new_n1943__));
  buf1  g0289(.din(n1968_lo), .dout(new_new_n1944__));
  buf1  g0290(.din(n1971_lo), .dout(new_new_n1946__));
  buf1  g0291(.din(n1980_lo), .dout(new_new_n1948__));
  not1  g0292(.din(n1983_lo), .dout(new_new_n1951__));
  buf1  g0293(.din(n1992_lo), .dout(new_new_n1952__));
  buf1  g0294(.din(n1995_lo), .dout(new_new_n1954__));
  buf1  g0295(.din(n2004_lo), .dout(new_new_n1956__));
  buf1  g0296(.din(n2016_lo), .dout(new_new_n1958__));
  buf1  g0297(.din(n2019_lo), .dout(new_new_n1960__));
  buf1  g0298(.din(n2028_lo), .dout(new_new_n1962__));
  buf1  g0299(.din(n2040_lo), .dout(new_new_n1964__));
  buf1  g0300(.din(n2043_lo), .dout(new_new_n1966__));
  buf1  g0301(.din(n2046_lo), .dout(new_new_n1968__));
  not1  g0302(.din(n2049_lo), .dout(new_new_n1971__));
  buf1  g0303(.din(n2052_lo), .dout(new_new_n1972__));
  buf1  g0304(.din(n2055_lo), .dout(new_new_n1974__));
  buf1  g0305(.din(n2064_lo), .dout(new_new_n1976__));
  buf1  g0306(.din(n2067_lo), .dout(new_new_n1978__));
  buf1  g0307(.din(n2076_lo), .dout(new_new_n1980__));
  buf1  g0308(.din(n2079_lo), .dout(new_new_n1982__));
  buf1  g0309(.din(n2088_lo), .dout(new_new_n1984__));
  buf1  g0310(.din(n2091_lo), .dout(new_new_n1986__));
  buf1  g0311(.din(n2100_lo), .dout(new_new_n1988__));
  buf1  g0312(.din(n2103_lo), .dout(new_new_n1990__));
  buf1  g0313(.din(n2112_lo), .dout(new_new_n1992__));
  not1  g0314(.din(n2115_lo), .dout(new_new_n1995__));
  buf1  g0315(.din(n2124_lo), .dout(new_new_n1996__));
  buf1  g0316(.din(n2127_lo), .dout(new_new_n1998__));
  buf1  g0317(.din(n2136_lo), .dout(new_new_n2000__));
  buf1  g0318(.din(n2148_lo), .dout(new_new_n2002__));
  buf1  g0319(.din(n2151_lo), .dout(new_new_n2004__));
  buf1  g0320(.din(n2160_lo), .dout(new_new_n2006__));
  buf1  g0321(.din(n2172_lo), .dout(new_new_n2008__));
  buf1  g0322(.din(n2175_lo), .dout(new_new_n2010__));
  buf1  g0323(.din(n2178_lo), .dout(new_new_n2012__));
  not1  g0324(.din(n2181_lo), .dout(new_new_n2015__));
  buf1  g0325(.din(n2184_lo), .dout(new_new_n2016__));
  buf1  g0326(.din(n2187_lo), .dout(new_new_n2018__));
  buf1  g0327(.din(n2196_lo), .dout(new_new_n2020__));
  buf1  g0328(.din(n2199_lo), .dout(new_new_n2022__));
  buf1  g0329(.din(n2208_lo), .dout(new_new_n2024__));
  buf1  g0330(.din(n2211_lo), .dout(new_new_n2026__));
  buf1  g0331(.din(n2220_lo), .dout(new_new_n2028__));
  not1  g0332(.din(n2223_lo), .dout(new_new_n2031__));
  buf1  g0333(.din(n2232_lo), .dout(new_new_n2032__));
  not1  g0334(.din(n2235_lo), .dout(new_new_n2035__));
  buf1  g0335(.din(n2244_lo), .dout(new_new_n2036__));
  not1  g0336(.din(n2247_lo), .dout(new_new_n2039__));
  buf1  g0337(.din(n2256_lo), .dout(new_new_n2040__));
  buf1  g0338(.din(n2259_lo), .dout(new_new_n2042__));
  buf1  g0339(.din(n2268_lo), .dout(new_new_n2044__));
  buf1  g0340(.din(n2280_lo), .dout(new_new_n2046__));
  buf1  g0341(.din(n2283_lo), .dout(new_new_n2048__));
  buf1  g0342(.din(n2292_lo), .dout(new_new_n2050__));
  buf1  g0343(.din(n2295_lo), .dout(new_new_n2052__));
  buf1  g0344(.din(n2298_lo), .dout(new_new_n2054__));
  buf1  g0345(.din(n2301_lo), .dout(new_new_n2056__));
  buf1  g0346(.din(n2304_lo), .dout(new_new_n2058__));
  buf1  g0347(.din(n2307_lo), .dout(new_new_n2060__));
  buf1  g0348(.din(n2316_lo), .dout(new_new_n2062__));
  buf1  g0349(.din(n2319_lo), .dout(new_new_n2064__));
  buf1  g0350(.din(n2322_lo), .dout(new_new_n2066__));
  not1  g0351(.din(n2325_lo), .dout(new_new_n2069__));
  buf1  g0352(.din(n2328_lo), .dout(new_new_n2070__));
  buf1  g0353(.din(n2331_lo), .dout(new_new_n2072__));
  buf1  g0354(.din(n2340_lo), .dout(new_new_n2074__));
  buf1  g0355(.din(n2343_lo), .dout(new_new_n2076__));
  buf1  g0356(.din(n2376_lo), .dout(new_new_n2078__));
  buf1  g0357(.din(n2379_lo), .dout(new_new_n2080__));
  buf1  g0358(.din(n2388_lo), .dout(new_new_n2082__));
  buf1  g0359(.din(n2391_lo), .dout(new_new_n2084__));
  buf1  g0360(.din(n2400_lo), .dout(new_new_n2086__));
  buf1  g0361(.din(n2403_lo), .dout(new_new_n2088__));
  buf1  g0362(.din(n2412_lo), .dout(new_new_n2090__));
  buf1  g0363(.din(n2415_lo), .dout(new_new_n2092__));
  buf1  g0364(.din(n2424_lo), .dout(new_new_n2094__));
  buf1  g0365(.din(n2427_lo), .dout(new_new_n2096__));
  buf1  g0366(.din(n2436_lo), .dout(new_new_n2098__));
  buf1  g0367(.din(n2439_lo), .dout(new_new_n2100__));
  buf1  g0368(.din(n2442_lo), .dout(new_new_n2102__));
  not1  g0369(.din(n2445_lo), .dout(new_new_n2105__));
  buf1  g0370(.din(n2448_lo), .dout(new_new_n2106__));
  buf1  g0371(.din(n2451_lo), .dout(new_new_n2108__));
  buf1  g0372(.din(n2460_lo), .dout(new_new_n2110__));
  buf1  g0373(.din(n2463_lo), .dout(new_new_n2112__));
  buf1  g0374(.din(n2496_lo), .dout(new_new_n2114__));
  buf1  g0375(.din(n2499_lo), .dout(new_new_n2116__));
  buf1  g0376(.din(n2508_lo), .dout(new_new_n2118__));
  buf1  g0377(.din(n2511_lo), .dout(new_new_n2120__));
  buf1  g0378(.din(n2520_lo), .dout(new_new_n2122__));
  buf1  g0379(.din(n2523_lo), .dout(new_new_n2124__));
  buf1  g0380(.din(n2532_lo), .dout(new_new_n2126__));
  buf1  g0381(.din(n2535_lo), .dout(new_new_n2128__));
  buf1  g0382(.din(n2544_lo), .dout(new_new_n2130__));
  buf1  g0383(.din(n2547_lo), .dout(new_new_n2132__));
  buf1  g0384(.din(n2556_lo), .dout(new_new_n2134__));
  buf1  g0385(.din(n2559_lo), .dout(new_new_n2136__));
  buf1  g0386(.din(n2562_lo), .dout(new_new_n2138__));
  not1  g0387(.din(n2565_lo), .dout(new_new_n2141__));
  buf1  g0388(.din(n2568_lo), .dout(new_new_n2142__));
  buf1  g0389(.din(n2571_lo), .dout(new_new_n2144__));
  buf1  g0390(.din(n2580_lo), .dout(new_new_n2146__));
  buf1  g0391(.din(n2583_lo), .dout(new_new_n2148__));
  buf1  g0392(.din(n2616_lo), .dout(new_new_n2150__));
  buf1  g0393(.din(n2619_lo), .dout(new_new_n2152__));
  buf1  g0394(.din(n2628_lo), .dout(new_new_n2154__));
  buf1  g0395(.din(n2631_lo), .dout(new_new_n2156__));
  buf1  g0396(.din(n2640_lo), .dout(new_new_n2158__));
  buf1  g0397(.din(n2643_lo), .dout(new_new_n2160__));
  buf1  g0398(.din(n2652_lo), .dout(new_new_n2162__));
  buf1  g0399(.din(n2655_lo), .dout(new_new_n2164__));
  buf1  g0400(.din(n2664_lo), .dout(new_new_n2166__));
  buf1  g0401(.din(n2667_lo), .dout(new_new_n2168__));
  buf1  g0402(.din(n2676_lo), .dout(new_new_n2170__));
  buf1  g0403(.din(n2679_lo), .dout(new_new_n2172__));
  buf1  g0404(.din(n2682_lo), .dout(new_new_n2174__));
  not1  g0405(.din(n2685_lo), .dout(new_new_n2177__));
  buf1  g0406(.din(n2688_lo), .dout(new_new_n2178__));
  buf1  g0407(.din(n2691_lo), .dout(new_new_n2180__));
  buf1  g0408(.din(n2700_lo), .dout(new_new_n2182__));
  buf1  g0409(.din(n2703_lo), .dout(new_new_n2184__));
  buf1  g0410(.din(n2736_lo), .dout(new_new_n2186__));
  buf1  g0411(.din(n2739_lo), .dout(new_new_n2188__));
  buf1  g0412(.din(n2748_lo), .dout(new_new_n2190__));
  buf1  g0413(.din(n2751_lo), .dout(new_new_n2192__));
  buf1  g0414(.din(n2760_lo), .dout(new_new_n2194__));
  buf1  g0415(.din(n2763_lo), .dout(new_new_n2196__));
  buf1  g0416(.din(n2772_lo), .dout(new_new_n2198__));
  buf1  g0417(.din(n2775_lo), .dout(new_new_n2200__));
  buf1  g0418(.din(n2784_lo), .dout(new_new_n2202__));
  buf1  g0419(.din(n2787_lo), .dout(new_new_n2204__));
  buf1  g0420(.din(n2790_lo), .dout(new_new_n2206__));
  buf1  g0421(.din(n2793_lo), .dout(new_new_n2208__));
  not1  g0422(.din(n2793_lo), .dout(new_new_n2209__));
  buf1  g0423(.din(n2796_lo), .dout(new_new_n2210__));
  buf1  g0424(.din(n2799_lo), .dout(new_new_n2212__));
  buf1  g0425(.din(n2802_lo), .dout(new_new_n2214__));
  not1  g0426(.din(n2805_lo), .dout(new_new_n2217__));
  buf1  g0427(.din(n2808_lo), .dout(new_new_n2218__));
  not1  g0428(.din(n2808_lo), .dout(new_new_n2219__));
  buf1  g0429(.din(n2820_lo), .dout(new_new_n2220__));
  buf1  g0430(.din(n2823_lo), .dout(new_new_n2222__));
  buf1  g0431(.din(n2826_lo), .dout(new_new_n2224__));
  buf1  g0432(.din(n2829_lo), .dout(new_new_n2226__));
  not1  g0433(.din(n2829_lo), .dout(new_new_n2227__));
  buf1  g0434(.din(n2832_lo), .dout(new_new_n2228__));
  buf1  g0435(.din(n2835_lo), .dout(new_new_n2230__));
  buf1  g0436(.din(n2838_lo), .dout(new_new_n2232__));
  buf1  g0437(.din(n2841_lo), .dout(new_new_n2234__));
  not1  g0438(.din(n2841_lo), .dout(new_new_n2235__));
  buf1  g0439(.din(n2844_lo), .dout(new_new_n2236__));
  not1  g0440(.din(n2844_lo), .dout(new_new_n2237__));
  buf1  g0441(.din(n2856_lo), .dout(new_new_n2238__));
  buf1  g0442(.din(n2859_lo), .dout(new_new_n2240__));
  buf1  g0443(.din(n2862_lo), .dout(new_new_n2242__));
  buf1  g0444(.din(n2865_lo), .dout(new_new_n2244__));
  not1  g0445(.din(n2865_lo), .dout(new_new_n2245__));
  buf1  g0446(.din(n2868_lo), .dout(new_new_n2246__));
  buf1  g0447(.din(n2871_lo), .dout(new_new_n2248__));
  buf1  g0448(.din(n2874_lo), .dout(new_new_n2250__));
  buf1  g0449(.din(n2877_lo), .dout(new_new_n2252__));
  not1  g0450(.din(n2877_lo), .dout(new_new_n2253__));
  buf1  g0451(.din(n2880_lo), .dout(new_new_n2254__));
  buf1  g0452(.din(n2883_lo), .dout(new_new_n2256__));
  buf1  g0453(.din(n2886_lo), .dout(new_new_n2258__));
  buf1  g0454(.din(n2889_lo), .dout(new_new_n2260__));
  not1  g0455(.din(n2889_lo), .dout(new_new_n2261__));
  buf1  g0456(.din(n2892_lo), .dout(new_new_n2262__));
  buf1  g0457(.din(n2895_lo), .dout(new_new_n2264__));
  buf1  g0458(.din(n2898_lo), .dout(new_new_n2266__));
  not1  g0459(.din(n2901_lo), .dout(new_new_n2269__));
  buf1  g0460(.din(n2904_lo), .dout(new_new_n2270__));
  buf1  g0461(.din(n2907_lo), .dout(new_new_n2272__));
  buf1  g0462(.din(n2916_lo), .dout(new_new_n2274__));
  buf1  g0463(.din(n2919_lo), .dout(new_new_n2276__));
  not1  g0464(.din(n2925_lo), .dout(new_new_n2279__));
  buf1  g0465(.din(n2928_lo), .dout(new_new_n2280__));
  buf1  g0466(.din(n2940_lo), .dout(new_new_n2282__));
  buf1  g0467(.din(n2943_lo), .dout(new_new_n2284__));
  buf1  g0468(.din(n2952_lo), .dout(new_new_n2286__));
  buf1  g0469(.din(n2955_lo), .dout(new_new_n2288__));
  buf1  g0470(.din(n2961_lo), .dout(new_new_n2290__));
  not1  g0471(.din(n2961_lo), .dout(new_new_n2291__));
  buf1  g0472(.din(n2964_lo), .dout(new_new_n2292__));
  buf1  g0473(.din(n2967_lo), .dout(new_new_n2294__));
  buf1  g0474(.din(n2970_lo), .dout(new_new_n2296__));
  not1  g0475(.din(n2970_lo), .dout(new_new_n2297__));
  buf1  g0476(.din(n2976_lo), .dout(new_new_n2298__));
  buf1  g0477(.din(n2979_lo), .dout(new_new_n2300__));
  buf1  g0478(.din(n2982_lo), .dout(new_new_n2302__));
  not1  g0479(.din(n2982_lo), .dout(new_new_n2303__));
  buf1  g0480(.din(n2988_lo), .dout(new_new_n2304__));
  buf1  g0481(.din(n2991_lo), .dout(new_new_n2306__));
  buf1  g0482(.din(n2994_lo), .dout(new_new_n2308__));
  not1  g0483(.din(n2994_lo), .dout(new_new_n2309__));
  buf1  g0484(.din(n2997_lo), .dout(new_new_n2310__));
  buf1  g0485(.din(n3000_lo), .dout(new_new_n2312__));
  buf1  g0486(.din(n3003_lo), .dout(new_new_n2314__));
  buf1  g0487(.din(n3006_lo), .dout(new_new_n2316__));
  not1  g0488(.din(n3006_lo), .dout(new_new_n2317__));
  buf1  g0489(.din(n3012_lo), .dout(new_new_n2318__));
  buf1  g0490(.din(n3015_lo), .dout(new_new_n2320__));
  buf1  g0491(.din(n3018_lo), .dout(new_new_n2322__));
  not1  g0492(.din(n3018_lo), .dout(new_new_n2323__));
  not1  g0493(.din(n3021_lo), .dout(new_new_n2325__));
  buf1  g0494(.din(n3024_lo), .dout(new_new_n2326__));
  buf1  g0495(.din(n3027_lo), .dout(new_new_n2328__));
  buf1  g0496(.din(n3030_lo), .dout(new_new_n2330__));
  not1  g0497(.din(n3030_lo), .dout(new_new_n2331__));
  buf1  g0498(.din(n3033_lo), .dout(new_new_n2332__));
  not1  g0499(.din(n3033_lo), .dout(new_new_n2333__));
  buf1  g0500(.din(n3036_lo), .dout(new_new_n2334__));
  buf1  g0501(.din(n3039_lo), .dout(new_new_n2336__));
  buf1  g0502(.din(n3045_lo), .dout(new_new_n2338__));
  not1  g0503(.din(n3045_lo), .dout(new_new_n2339__));
  buf1  g0504(.din(n3048_lo), .dout(new_new_n2340__));
  buf1  g0505(.din(n3051_lo), .dout(new_new_n2342__));
  buf1  g0506(.din(n3054_lo), .dout(new_new_n2344__));
  not1  g0507(.din(n3057_lo), .dout(new_new_n2347__));
  buf1  g0508(.din(n3060_lo), .dout(new_new_n2348__));
  buf1  g0509(.din(n3063_lo), .dout(new_new_n2350__));
  buf1  g0510(.din(n3069_lo), .dout(new_new_n2352__));
  not1  g0511(.din(n3069_lo), .dout(new_new_n2353__));
  buf1  g0512(.din(n3072_lo), .dout(new_new_n2354__));
  buf1  g0513(.din(n3075_lo), .dout(new_new_n2356__));
  buf1  g0514(.din(n3081_lo), .dout(new_new_n2358__));
  buf1  g0515(.din(n3084_lo), .dout(new_new_n2360__));
  buf1  g0516(.din(n3087_lo), .dout(new_new_n2362__));
  not1  g0517(.din(n3093_lo), .dout(new_new_n2365__));
  buf1  g0518(.din(n3096_lo), .dout(new_new_n2366__));
  buf1  g0519(.din(n3099_lo), .dout(new_new_n2368__));
  buf1  g0520(.din(n3102_lo), .dout(new_new_n2370__));
  not1  g0521(.din(n3102_lo), .dout(new_new_n2371__));
  buf1  g0522(.din(n3105_lo), .dout(new_new_n2372__));
  buf1  g0523(.din(n3108_lo), .dout(new_new_n2374__));
  buf1  g0524(.din(n3111_lo), .dout(new_new_n2376__));
  buf1  g0525(.din(n3114_lo), .dout(new_new_n2378__));
  not1  g0526(.din(n3114_lo), .dout(new_new_n2379__));
  buf1  g0527(.din(n3117_lo), .dout(new_new_n2380__));
  not1  g0528(.din(n3117_lo), .dout(new_new_n2381__));
  buf1  g0529(.din(n3120_lo), .dout(new_new_n2382__));
  buf1  g0530(.din(n3123_lo), .dout(new_new_n2384__));
  buf1  g0531(.din(n3126_lo), .dout(new_new_n2386__));
  not1  g0532(.din(n3126_lo), .dout(new_new_n2387__));
  buf1  g0533(.din(n3129_lo), .dout(new_new_n2388__));
  not1  g0534(.din(n3129_lo), .dout(new_new_n2389__));
  buf1  g0535(.din(n3132_lo), .dout(new_new_n2390__));
  buf1  g0536(.din(n3135_lo), .dout(new_new_n2392__));
  buf1  g0537(.din(n3138_lo), .dout(new_new_n2394__));
  not1  g0538(.din(n3138_lo), .dout(new_new_n2395__));
  buf1  g0539(.din(n3141_lo), .dout(new_new_n2396__));
  buf1  g0540(.din(n3156_lo), .dout(new_new_n2398__));
  not1  g0541(.din(n3156_lo), .dout(new_new_n2399__));
  buf1  g0542(.din(n3168_lo), .dout(new_new_n2400__));
  buf1  g0543(.din(n3171_lo), .dout(new_new_n2402__));
  buf1  g0544(.din(n3174_lo), .dout(new_new_n2404__));
  buf1  g0545(.din(n3177_lo), .dout(new_new_n2406__));
  not1  g0546(.din(n3177_lo), .dout(new_new_n2407__));
  buf1  g0547(.din(n3180_lo), .dout(new_new_n2408__));
  buf1  g0548(.din(n3183_lo), .dout(new_new_n2410__));
  buf1  g0549(.din(n3192_lo), .dout(new_new_n2412__));
  buf1  g0550(.din(n3195_lo), .dout(new_new_n2414__));
  buf1  g0551(.din(n3204_lo), .dout(new_new_n2416__));
  buf1  g0552(.din(n3207_lo), .dout(new_new_n2418__));
  buf1  g0553(.din(n3210_lo), .dout(new_new_n2420__));
  not1  g0554(.din(n3210_lo), .dout(new_new_n2421__));
  buf1  g0555(.din(n3216_lo), .dout(new_new_n2422__));
  buf1  g0556(.din(n3219_lo), .dout(new_new_n2424__));
  buf1  g0557(.din(n3222_lo), .dout(new_new_n2426__));
  not1  g0558(.din(n3222_lo), .dout(new_new_n2427__));
  buf1  g0559(.din(n3228_lo), .dout(new_new_n2428__));
  buf1  g0560(.din(n3231_lo), .dout(new_new_n2430__));
  buf1  g0561(.din(n3240_lo), .dout(new_new_n2432__));
  buf1  g0562(.din(n3243_lo), .dout(new_new_n2434__));
  buf1  g0563(.din(n3252_lo), .dout(new_new_n2436__));
  buf1  g0564(.din(n3255_lo), .dout(new_new_n2438__));
  buf1  g0565(.din(n3258_lo), .dout(new_new_n2440__));
  not1  g0566(.din(n3258_lo), .dout(new_new_n2441__));
  buf1  g0567(.din(n3264_lo), .dout(new_new_n2442__));
  buf1  g0568(.din(n3267_lo), .dout(new_new_n2444__));
  buf1  g0569(.din(n3270_lo), .dout(new_new_n2446__));
  not1  g0570(.din(n3270_lo), .dout(new_new_n2447__));
  buf1  g0571(.din(n3276_lo), .dout(new_new_n2448__));
  buf1  g0572(.din(n3279_lo), .dout(new_new_n2450__));
  buf1  g0573(.din(n3282_lo), .dout(new_new_n2452__));
  not1  g0574(.din(n3282_lo), .dout(new_new_n2453__));
  buf1  g0575(.din(n3288_lo), .dout(new_new_n2454__));
  buf1  g0576(.din(n3291_lo), .dout(new_new_n2456__));
  buf1  g0577(.din(n3294_lo), .dout(new_new_n2458__));
  not1  g0578(.din(n3294_lo), .dout(new_new_n2459__));
  not1  g0579(.din(n3603_o2), .dout(new_new_n2461__));
  not1  g0580(.din(n3604_o2), .dout(new_new_n2463__));
  not1  g0581(.din(n1391_inv), .dout(new_new_n2465__));
  buf1  g0582(.din(n3798_o2), .dout(new_new_n2466__));
  not1  g0583(.din(n3798_o2), .dout(new_new_n2467__));
  buf1  g0584(.din(n3846_o2), .dout(new_new_n2468__));
  not1  g0585(.din(n3846_o2), .dout(new_new_n2469__));
  buf1  g0586(.din(n4019_o2), .dout(new_new_n2470__));
  buf1  g0587(.din(n4017_o2), .dout(new_new_n2472__));
  not1  g0588(.din(n4017_o2), .dout(new_new_n2473__));
  buf1  g0589(.din(n2177_o2), .dout(new_new_n2474__));
  not1  g0590(.din(n2150_o2), .dout(new_new_n2477__));
  not1  g0591(.din(n2154_o2), .dout(new_new_n2479__));
  buf1  g0592(.din(n2184_o2), .dout(new_new_n2480__));
  buf1  g0593(.din(n2515_o2), .dout(new_new_n2482__));
  buf1  g0594(.din(n3837_o2), .dout(new_new_n2484__));
  not1  g0595(.din(n3837_o2), .dout(new_new_n2485__));
  not1  g0596(.din(n2167_o2), .dout(new_new_n2487__));
  not1  g0597(.din(n2118_o2), .dout(new_new_n2489__));
  buf1  g0598(.din(n2186_o2), .dout(new_new_n2490__));
  not1  g0599(.din(n2174_o2), .dout(new_new_n2493__));
  buf1  g0600(.din(n3964_o2), .dout(new_new_n2494__));
  not1  g0601(.din(n3964_o2), .dout(new_new_n2495__));
  buf1  g0602(.din(n4005_o2), .dout(new_new_n2496__));
  not1  g0603(.din(n4005_o2), .dout(new_new_n2497__));
  buf1  g0604(.din(n4006_o2), .dout(new_new_n2498__));
  not1  g0605(.din(n4006_o2), .dout(new_new_n2499__));
  not1  g0606(.din(n1445_inv), .dout(new_new_n2501__));
  buf1  g0607(.din(n2176_o2), .dout(new_new_n2502__));
  buf1  g0608(.din(n2227_o2), .dout(new_new_n2504__));
  buf1  g0609(.din(n2236_o2), .dout(new_new_n2506__));
  buf1  g0610(.din(n2245_o2), .dout(new_new_n2508__));
  buf1  g0611(.din(n2518_o2), .dout(new_new_n2510__));
  not1  g0612(.din(n2518_o2), .dout(new_new_n2511__));
  buf1  g0613(.din(n4023_o2), .dout(new_new_n2512__));
  buf1  g0614(.din(n1466_inv), .dout(new_new_n2514__));
  buf1  g0615(.din(n4038_o2), .dout(new_new_n2516__));
  not1  g0616(.din(n4038_o2), .dout(new_new_n2517__));
  buf1  g0617(.din(n4039_o2), .dout(new_new_n2518__));
  not1  g0618(.din(n4039_o2), .dout(new_new_n2519__));
  buf1  g0619(.din(n1475_inv), .dout(new_new_n2520__));
  not1  g0620(.din(n1475_inv), .dout(new_new_n2521__));
  not1  g0621(.din(n2119_o2), .dout(new_new_n2523__));
  buf1  g0622(.din(n2275_o2), .dout(new_new_n2524__));
  not1  g0623(.din(n2275_o2), .dout(new_new_n2525__));
  buf1  g0624(.din(n2595_o2), .dout(new_new_n2526__));
  not1  g0625(.din(n2595_o2), .dout(new_new_n2527__));
  buf1  g0626(.din(n2594_o2), .dout(new_new_n2528__));
  not1  g0627(.din(n2594_o2), .dout(new_new_n2529__));
  buf1  g0628(.din(lo498_buf_o2), .dout(new_new_n2530__));
  not1  g0629(.din(lo498_buf_o2), .dout(new_new_n2531__));
  buf1  g0630(.din(lo502_buf_o2), .dout(new_new_n2532__));
  not1  g0631(.din(lo502_buf_o2), .dout(new_new_n2533__));
  buf1  g0632(.din(lo550_buf_o2), .dout(new_new_n2534__));
  not1  g0633(.din(lo550_buf_o2), .dout(new_new_n2535__));
  buf1  g0634(.din(n2596_o2), .dout(new_new_n2536__));
  not1  g0635(.din(n2596_o2), .dout(new_new_n2537__));
  buf1  g0636(.din(n2593_o2), .dout(new_new_n2538__));
  not1  g0637(.din(n2668_o2), .dout(new_new_n2541__));
  buf1  g0638(.din(lo542_buf_o2), .dout(new_new_n2542__));
  not1  g0639(.din(lo542_buf_o2), .dout(new_new_n2543__));
  buf1  g0640(.din(n2667_o2), .dout(new_new_n2544__));
  buf1  g0641(.din(n2404_o2), .dout(new_new_n2546__));
  buf1  g0642(.din(n2410_o2), .dout(new_new_n2548__));
  not1  g0643(.din(n2419_o2), .dout(new_new_n2551__));
  buf1  g0644(.din(n2392_o2), .dout(new_new_n2552__));
  not1  g0645(.din(n2369_o2), .dout(new_new_n2555__));
  not1  g0646(.din(n2397_o2), .dout(new_new_n2557__));
  not1  g0647(.din(n2601_o2), .dout(new_new_n2559__));
  not1  g0648(.din(n2658_o2), .dout(new_new_n2561__));
  buf1  g0649(.din(n2574_o2), .dout(new_new_n2562__));
  not1  g0650(.din(n2574_o2), .dout(new_new_n2563__));
  buf1  g0651(.din(n2205_o2), .dout(new_new_n2564__));
  not1  g0652(.din(n2205_o2), .dout(new_new_n2565__));
  buf1  g0653(.din(lo510_buf_o2), .dout(new_new_n2566__));
  not1  g0654(.din(lo510_buf_o2), .dout(new_new_n2567__));
  buf1  g0655(.din(lo514_buf_o2), .dout(new_new_n2568__));
  not1  g0656(.din(lo514_buf_o2), .dout(new_new_n2569__));
  buf1  g0657(.din(lo554_buf_o2), .dout(new_new_n2570__));
  not1  g0658(.din(lo554_buf_o2), .dout(new_new_n2571__));
  buf1  g0659(.din(lo558_buf_o2), .dout(new_new_n2572__));
  not1  g0660(.din(lo558_buf_o2), .dout(new_new_n2573__));
  buf1  g0661(.din(lo578_buf_o2), .dout(new_new_n2574__));
  not1  g0662(.din(lo578_buf_o2), .dout(new_new_n2575__));
  buf1  g0663(.din(n2254_o2), .dout(new_new_n2576__));
  not1  g0664(.din(n2254_o2), .dout(new_new_n2577__));
  not1  g0665(.din(n2421_o2), .dout(new_new_n2579__));
  not1  g0666(.din(n2422_o2), .dout(new_new_n2581__));
  not1  g0667(.din(n2130_o2), .dout(new_new_n2583__));
  not1  g0668(.din(n2127_o2), .dout(new_new_n2585__));
  not1  g0669(.din(n2131_o2), .dout(new_new_n2587__));
  not1  g0670(.din(n2128_o2), .dout(new_new_n2589__));
  buf1  g0671(.din(n2264_o2), .dout(new_new_n2590__));
  not1  g0672(.din(n2264_o2), .dout(new_new_n2591__));
  buf1  g0673(.din(n2467_o2), .dout(new_new_n2592__));
  buf1  g0674(.din(n2471_o2), .dout(new_new_n2594__));
  buf1  g0675(.din(n2488_o2), .dout(new_new_n2596__));
  buf1  g0676(.din(n2478_o2), .dout(new_new_n2598__));
  buf1  g0677(.din(n2486_o2), .dout(new_new_n2600__));
  buf1  g0678(.din(n2485_o2), .dout(new_new_n2602__));
  buf1  g0679(.din(n2498_o2), .dout(new_new_n2604__));
  buf1  g0680(.din(n2495_o2), .dout(new_new_n2606__));
  buf1  g0681(.din(n2496_o2), .dout(new_new_n2608__));
  buf1  g0682(.din(n2458_o2), .dout(new_new_n2610__));
  buf1  g0683(.din(n2643_o2), .dout(new_new_n2612__));
  not1  g0684(.din(n2643_o2), .dout(new_new_n2613__));
  buf1  g0685(.din(n2462_o2), .dout(new_new_n2614__));
  buf1  g0686(.din(n2468_o2), .dout(new_new_n2616__));
  buf1  g0687(.din(n2639_o2), .dout(new_new_n2618__));
  not1  g0688(.din(n2639_o2), .dout(new_new_n2619__));
  buf1  g0689(.din(n2499_o2), .dout(new_new_n2620__));
  buf1  g0690(.din(n2472_o2), .dout(new_new_n2622__));
  buf1  g0691(.din(n2474_o2), .dout(new_new_n2624__));
  buf1  g0692(.din(n2489_o2), .dout(new_new_n2626__));
  buf1  g0693(.din(n2321_o2), .dout(new_new_n2628__));
  not1  g0694(.din(n2321_o2), .dout(new_new_n2629__));
  buf1  g0695(.din(n2322_o2), .dout(new_new_n2630__));
  not1  g0696(.din(n2322_o2), .dout(new_new_n2631__));
  buf1  g0697(.din(n2640_o2), .dout(new_new_n2632__));
  buf1  g0698(.din(n2642_o2), .dout(new_new_n2634__));
  buf1  g0699(.din(n2187_o2), .dout(new_new_n2636__));
  not1  g0700(.din(n2187_o2), .dout(new_new_n2637__));
  buf1  g0701(.din(n2373_o2), .dout(new_new_n2638__));
  not1  g0702(.din(n2373_o2), .dout(new_new_n2639__));
  buf1  g0703(.din(n2603_o2), .dout(new_new_n2640__));
  buf1  g0704(.din(n2388_o2), .dout(new_new_n2642__));
  not1  g0705(.din(n2388_o2), .dout(new_new_n2643__));
  buf1  g0706(.din(n2437_o2), .dout(new_new_n2644__));
  not1  g0707(.din(n2437_o2), .dout(new_new_n2645__));
  buf1  g0708(.din(n2356_o2), .dout(new_new_n2646__));
  not1  g0709(.din(n2356_o2), .dout(new_new_n2647__));
  buf1  g0710(.din(n2452_o2), .dout(new_new_n2648__));
  not1  g0711(.din(n2452_o2), .dout(new_new_n2649__));
  buf1  g0712(.din(n2347_o2), .dout(new_new_n2650__));
  not1  g0713(.din(n2347_o2), .dout(new_new_n2651__));
  buf1  g0714(.din(n2329_o2), .dout(new_new_n2652__));
  not1  g0715(.din(n2329_o2), .dout(new_new_n2653__));
  buf1  g0716(.din(n2669_o2), .dout(new_new_n2654__));
  not1  g0717(.din(n2669_o2), .dout(new_new_n2655__));
  buf1  g0718(.din(n2332_o2), .dout(new_new_n2656__));
  not1  g0719(.din(n2332_o2), .dout(new_new_n2657__));
  buf1  g0720(.din(n2664_o2), .dout(new_new_n2658__));
  not1  g0721(.din(n2664_o2), .dout(new_new_n2659__));
  buf1  g0722(.din(n2665_o2), .dout(new_new_n2660__));
  buf1  g0723(.din(n2653_o2), .dout(new_new_n2662__));
  not1  g0724(.din(n2653_o2), .dout(new_new_n2663__));
  buf1  g0725(.din(n2654_o2), .dout(new_new_n2664__));
  buf1  g0726(.din(n2636_o2), .dout(new_new_n2666__));
  buf1  g0727(.din(n2660_o2), .dout(new_new_n2668__));
  buf1  g0728(.din(n2318_o2), .dout(new_new_n2670__));
  not1  g0729(.din(n2318_o2), .dout(new_new_n2671__));
  buf1  g0730(.din(n2319_o2), .dout(new_new_n2672__));
  not1  g0731(.din(n2319_o2), .dout(new_new_n2673__));
  buf1  g0732(.din(n2586_o2), .dout(new_new_n2674__));
  not1  g0733(.din(n2586_o2), .dout(new_new_n2675__));
  buf1  g0734(.din(n2587_o2), .dout(new_new_n2676__));
  not1  g0735(.din(n2587_o2), .dout(new_new_n2677__));
  buf1  g0736(.din(n2288_o2), .dout(new_new_n2678__));
  not1  g0737(.din(n2288_o2), .dout(new_new_n2679__));
  buf1  g0738(.din(n2344_o2), .dout(new_new_n2680__));
  not1  g0739(.din(n2344_o2), .dout(new_new_n2681__));
  buf1  g0740(.din(n2530_o2), .dout(new_new_n2682__));
  not1  g0741(.din(n2530_o2), .dout(new_new_n2683__));
  buf1  g0742(.din(n2303_o2), .dout(new_new_n2684__));
  not1  g0743(.din(n2303_o2), .dout(new_new_n2685__));
  buf1  g0744(.din(n2566_o2), .dout(new_new_n2686__));
  not1  g0745(.din(n2566_o2), .dout(new_new_n2687__));
  buf1  g0746(.din(n2567_o2), .dout(new_new_n2688__));
  not1  g0747(.din(n2567_o2), .dout(new_new_n2689__));
  buf1  g0748(.din(n2554_o2), .dout(new_new_n2690__));
  not1  g0749(.din(n2554_o2), .dout(new_new_n2691__));
  buf1  g0750(.din(n2194_o2), .dout(new_new_n2692__));
  not1  g0751(.din(n2194_o2), .dout(new_new_n2693__));
  buf1  g0752(.din(lo582_buf_o2), .dout(new_new_n2694__));
  not1  g0753(.din(lo582_buf_o2), .dout(new_new_n2695__));
  buf1  g0754(.din(lo030_buf_o2), .dout(new_new_n2696__));
  not1  g0755(.din(lo030_buf_o2), .dout(new_new_n2697__));
  buf1  g0756(.din(lo174_buf_o2), .dout(new_new_n2698__));
  not1  g0757(.din(lo174_buf_o2), .dout(new_new_n2699__));
  buf1  g0758(.din(lo178_buf_o2), .dout(new_new_n2700__));
  not1  g0759(.din(lo178_buf_o2), .dout(new_new_n2701__));
  buf1  g0760(.din(lo186_buf_o2), .dout(new_new_n2702__));
  not1  g0761(.din(lo186_buf_o2), .dout(new_new_n2703__));
  buf1  g0762(.din(lo266_buf_o2), .dout(new_new_n2704__));
  not1  g0763(.din(lo266_buf_o2), .dout(new_new_n2705__));
  buf1  g0764(.din(lo306_buf_o2), .dout(new_new_n2706__));
  not1  g0765(.din(lo306_buf_o2), .dout(new_new_n2707__));
  buf1  g0766(.din(lo346_buf_o2), .dout(new_new_n2708__));
  not1  g0767(.din(lo346_buf_o2), .dout(new_new_n2709__));
  buf1  g0768(.din(lo386_buf_o2), .dout(new_new_n2710__));
  not1  g0769(.din(lo386_buf_o2), .dout(new_new_n2711__));
  buf1  g0770(.din(lo426_buf_o2), .dout(new_new_n2712__));
  not1  g0771(.din(lo426_buf_o2), .dout(new_new_n2713__));
  buf1  g0772(.din(lo590_buf_o2), .dout(new_new_n2714__));
  not1  g0773(.din(lo590_buf_o2), .dout(new_new_n2715__));
  buf1  g0774(.din(lo594_buf_o2), .dout(new_new_n2716__));
  not1  g0775(.din(lo594_buf_o2), .dout(new_new_n2717__));
  buf1  g0776(.din(lo606_buf_o2), .dout(new_new_n2718__));
  not1  g0777(.din(lo606_buf_o2), .dout(new_new_n2719__));
  buf1  g0778(.din(lo610_buf_o2), .dout(new_new_n2720__));
  not1  g0779(.din(lo610_buf_o2), .dout(new_new_n2721__));
  buf1  g0780(.din(n2238_o2), .dout(new_new_n2722__));
  not1  g0781(.din(n2238_o2), .dout(new_new_n2723__));
  buf1  g0782(.din(n2229_o2), .dout(new_new_n2724__));
  not1  g0783(.din(n2229_o2), .dout(new_new_n2725__));
  buf1  g0784(.din(n2242_o2), .dout(new_new_n2726__));
  not1  g0785(.din(n2242_o2), .dout(new_new_n2727__));
  buf1  g0786(.din(n2233_o2), .dout(new_new_n2728__));
  not1  g0787(.din(n2233_o2), .dout(new_new_n2729__));
  buf1  g0788(.din(n2168_o2), .dout(new_new_n2730__));
  not1  g0789(.din(n2168_o2), .dout(new_new_n2731__));
  buf1  g0790(.din(n2237_o2), .dout(new_new_n2732__));
  not1  g0791(.din(n2237_o2), .dout(new_new_n2733__));
  buf1  g0792(.din(n2228_o2), .dout(new_new_n2734__));
  not1  g0793(.din(n2228_o2), .dout(new_new_n2735__));
  buf1  g0794(.din(n2172_o2), .dout(new_new_n2736__));
  not1  g0795(.din(n2172_o2), .dout(new_new_n2737__));
  buf1  g0796(.din(n2223_o2), .dout(new_new_n2738__));
  not1  g0797(.din(n2223_o2), .dout(new_new_n2739__));
  buf1  g0798(.din(n2222_o2), .dout(new_new_n2740__));
  not1  g0799(.din(n2222_o2), .dout(new_new_n2741__));
  buf1  g0800(.din(n2170_o2), .dout(new_new_n2742__));
  not1  g0801(.din(n2170_o2), .dout(new_new_n2743__));
  buf1  g0802(.din(n2181_o2), .dout(new_new_n2744__));
  not1  g0803(.din(n2181_o2), .dout(new_new_n2745__));
  buf1  g0804(.din(n2510_o2), .dout(new_new_n2746__));
  not1  g0805(.din(n2510_o2), .dout(new_new_n2747__));
  not1  g0806(.din(n2621_o2), .dout(new_new_n2749__));
  buf1  g0807(.din(lo466_buf_o2), .dout(new_new_n2750__));
  not1  g0808(.din(lo466_buf_o2), .dout(new_new_n2751__));
  buf1  g0809(.din(lo478_buf_o2), .dout(new_new_n2752__));
  not1  g0810(.din(lo478_buf_o2), .dout(new_new_n2753__));
  buf1  g0811(.din(n2149_o2), .dout(new_new_n2754__));
  not1  g0812(.din(n2149_o2), .dout(new_new_n2755__));
  buf1  g0813(.din(n2429_o2), .dout(new_new_n2756__));
  not1  g0814(.din(n2429_o2), .dout(new_new_n2757__));
  buf1  g0815(.din(n2444_o2), .dout(new_new_n2758__));
  not1  g0816(.din(n2444_o2), .dout(new_new_n2759__));
  buf1  g0817(.din(n2153_o2), .dout(new_new_n2760__));
  not1  g0818(.din(n2153_o2), .dout(new_new_n2761__));
  buf1  g0819(.din(n2433_o2), .dout(new_new_n2762__));
  not1  g0820(.din(n2433_o2), .dout(new_new_n2763__));
  buf1  g0821(.din(n2448_o2), .dout(new_new_n2764__));
  not1  g0822(.din(n2448_o2), .dout(new_new_n2765__));
  buf1  g0823(.din(n2367_o2), .dout(new_new_n2766__));
  not1  g0824(.din(n2367_o2), .dout(new_new_n2767__));
  buf1  g0825(.din(n2386_o2), .dout(new_new_n2768__));
  not1  g0826(.din(n2386_o2), .dout(new_new_n2769__));
  buf1  g0827(.din(n2539_o2), .dout(new_new_n2770__));
  not1  g0828(.din(n2539_o2), .dout(new_new_n2771__));
  buf1  g0829(.din(n2183_o2), .dout(new_new_n2772__));
  not1  g0830(.din(n2183_o2), .dout(new_new_n2773__));
  buf1  g0831(.din(n2220_o2), .dout(new_new_n2774__));
  not1  g0832(.din(n2220_o2), .dout(new_new_n2775__));
  buf1  g0833(.din(n2514_o2), .dout(new_new_n2776__));
  not1  g0834(.din(n2514_o2), .dout(new_new_n2777__));
  buf1  g0835(.din(n2196_o2), .dout(new_new_n2778__));
  not1  g0836(.din(n2616_o2), .dout(new_new_n2781__));
  not1  g0837(.din(n2612_o2), .dout(new_new_n2783__));
  not1  g0838(.din(n2627_o2), .dout(new_new_n2785__));
  buf1  g0839(.din(n2140_o2), .dout(new_new_n2786__));
  buf1  g0840(.din(n1877_inv), .dout(new_new_n2788__));
  not1  g0841(.din(lo149_buf_o2), .dout(new_new_n2791__));
  buf1  g0842(.din(lo197_buf_o2), .dout(new_new_n2792__));
  buf1  g0843(.din(lo118_buf_o2), .dout(new_new_n2794__));
  not1  g0844(.din(lo118_buf_o2), .dout(new_new_n2795__));
  buf1  g0845(.din(lo158_buf_o2), .dout(new_new_n2796__));
  buf1  g0846(.din(lo166_buf_o2), .dout(new_new_n2798__));
  buf1  g0847(.din(lo242_buf_o2), .dout(new_new_n2800__));
  buf1  g0848(.din(lo286_buf_o2), .dout(new_new_n2802__));
  buf1  g0849(.din(lo506_buf_o2), .dout(new_new_n2804__));
  not1  g0850(.din(lo506_buf_o2), .dout(new_new_n2805__));
  buf1  g0851(.din(n2198_o2), .dout(new_new_n2806__));
  buf1  g0852(.din(n2202_o2), .dout(new_new_n2808__));
  buf1  g0853(.din(n2197_o2), .dout(new_new_n2810__));
  buf1  g0854(.din(n1913_inv), .dout(new_new_n2812__));
  not1  g0855(.din(n1913_inv), .dout(new_new_n2813__));
  buf1  g0856(.din(n2146_o2), .dout(new_new_n2814__));
  not1  g0857(.din(n2146_o2), .dout(new_new_n2815__));
  buf1  g0858(.din(n1919_inv), .dout(new_new_n2816__));
  not1  g0859(.din(n1919_inv), .dout(new_new_n2817__));
  not1  g0860(.din(lo312_buf_o2), .dout(new_new_n2819__));
  buf1  g0861(.din(lo316_buf_o2), .dout(new_new_n2820__));
  not1  g0862(.din(lo352_buf_o2), .dout(new_new_n2823__));
  buf1  g0863(.din(lo356_buf_o2), .dout(new_new_n2824__));
  not1  g0864(.din(lo392_buf_o2), .dout(new_new_n2827__));
  buf1  g0865(.din(lo396_buf_o2), .dout(new_new_n2828__));
  not1  g0866(.din(lo432_buf_o2), .dout(new_new_n2831__));
  buf1  g0867(.din(lo436_buf_o2), .dout(new_new_n2832__));
  buf1  g0868(.din(lo576_buf_o2), .dout(new_new_n2834__));
  not1  g0869(.din(lo576_buf_o2), .dout(new_new_n2835__));
  or1   g0870(.dina(new_new_n2523__), .dinb(new_new_n2489__), .dout(new_new_n2836__));
  or1   g0871(.dina(new_new_n1763__), .dinb(new_new_n1701__), .dout(new_new_n2837__));
  or1   g0872(.dina(new_new_n2837__), .dinb(new_new_n4161__), .dout(new_new_n2838__));
  and1  g0873(.dina(new_new_n4163__), .dinb(new_new_n2056__), .dout(new_new_n2839__));
  or1   g0874(.dina(new_new_n4161__), .dinb(new_new_n1735__), .dout(new_new_n2840__));
  or1   g0875(.dina(new_new_n4166__), .dinb(new_new_n2235__), .dout(new_new_n2841__));
  or1   g0876(.dina(new_new_n4166__), .dinb(new_new_n2407__), .dout(new_new_n2842__));
  or1   g0877(.dina(new_new_n2589__), .dinb(new_new_n2585__), .dout(new_new_n2843__));
  or1   g0878(.dina(new_new_n2587__), .dinb(new_new_n2583__), .dout(new_new_n2844__));
  or1   g0879(.dina(new_new_n4167__), .dinb(new_new_n4168__), .dout(new_new_n2845__));
  and1  g0880(.dina(new_new_n4167__), .dinb(new_new_n2406__), .dout(new_new_n2846__));
  and1  g0881(.dina(new_new_n4168__), .dinb(new_new_n2234__), .dout(new_new_n2847__));
  or1   g0882(.dina(new_new_n2847__), .dinb(new_new_n2846__), .dout(new_new_n2848__));
  and1  g0883(.dina(new_new_n2463__), .dinb(new_new_n2461__), .dout(new_new_n2849__));
  and1  g0884(.dina(new_new_n2479__), .dinb(new_new_n2477__), .dout(new_new_n2850__));
  and1  g0885(.dina(new_new_n2493__), .dinb(new_new_n2487__), .dout(new_new_n2851__));
  or1   g0886(.dina(new_new_n2480__), .dinb(new_new_n2474__), .dout(new_new_n2852__));
  or1   g0887(.dina(new_new_n2466__), .dinb(new_new_n4170__), .dout(new_new_n2853__));
  or1   g0888(.dina(new_new_n2244__), .dinb(new_new_n2217__), .dout(new_new_n2854__));
  or1   g0889(.dina(new_new_n2854__), .dinb(new_new_n4172__), .dout(new_new_n2855__));
  or1   g0890(.dina(new_new_n4173__), .dinb(new_new_n1867__), .dout(new_new_n2856__));
  and1  g0891(.dina(new_new_n1708__), .dinb(new_new_n1692__), .dout(new_new_n2857__));
  or1   g0892(.dina(new_new_n2857__), .dinb(new_new_n4173__), .dout(new_new_n2858__));
  or1   g0893(.dina(new_new_n4174__), .dinb(new_new_n4176__), .dout(new_new_n2859__));
  or1   g0894(.dina(new_new_n4178__), .dinb(new_new_n4180__), .dout(new_new_n2860__));
  and1  g0895(.dina(new_new_n2860__), .dinb(new_new_n2859__), .dout(new_new_n2861__));
  and1  g0896(.dina(new_new_n2473__), .dinb(new_new_n4180__), .dout(new_new_n2862__));
  and1  g0897(.dina(new_new_n4182__), .dinb(new_new_n4176__), .dout(new_new_n2863__));
  or1   g0898(.dina(new_new_n2863__), .dinb(new_new_n2862__), .dout(new_new_n2864__));
  and1  g0899(.dina(new_new_n4170__), .dinb(new_new_n4183__), .dout(new_new_n2865__));
  or1   g0900(.dina(new_new_n2865__), .dinb(new_new_n4184__), .dout(new_new_n2866__));
  or1   g0901(.dina(new_new_n2467__), .dinb(new_new_n4177__), .dout(new_new_n2867__));
  or1   g0902(.dina(new_new_n4186__), .dinb(new_new_n4181__), .dout(new_new_n2868__));
  and1  g0903(.dina(new_new_n2868__), .dinb(new_new_n2867__), .dout(new_new_n2869__));
  or1   g0904(.dina(new_new_n2525__), .dinb(new_new_n2388__), .dout(new_new_n2870__));
  or1   g0905(.dina(new_new_n2524__), .dinb(new_new_n2389__), .dout(new_new_n2871__));
  and1  g0906(.dina(new_new_n2871__), .dinb(new_new_n2870__), .dout(new_new_n2872__));
  or1   g0907(.dina(new_new_n2872__), .dinb(new_new_n2396__), .dout(new_new_n2873__));
  or1   g0908(.dina(new_new_n2685__), .dinb(new_new_n2679__), .dout(new_new_n2874__));
  or1   g0909(.dina(new_new_n2684__), .dinb(new_new_n2678__), .dout(new_new_n2875__));
  and1  g0910(.dina(new_new_n2875__), .dinb(new_new_n1754__), .dout(new_new_n2876__));
  and1  g0911(.dina(new_new_n2876__), .dinb(new_new_n2874__), .dout(new_new_n2877__));
  and1  g0912(.dina(new_new_n2673__), .dinb(new_new_n2671__), .dout(new_new_n2878__));
  or1   g0913(.dina(new_new_n2672__), .dinb(new_new_n2670__), .dout(new_new_n2879__));
  and1  g0914(.dina(new_new_n2631__), .dinb(new_new_n2629__), .dout(new_new_n2880__));
  or1   g0915(.dina(new_new_n2630__), .dinb(new_new_n2628__), .dout(new_new_n2881__));
  or1   g0916(.dina(new_new_n2880__), .dinb(new_new_n2879__), .dout(new_new_n2882__));
  or1   g0917(.dina(new_new_n2881__), .dinb(new_new_n2878__), .dout(new_new_n2883__));
  and1  g0918(.dina(new_new_n2883__), .dinb(new_new_n2882__), .dout(new_new_n2884__));
  and1  g0919(.dina(new_new_n4187__), .dinb(new_new_n4188__), .dout(new_new_n2885__));
  or1   g0920(.dina(new_new_n4189__), .dinb(new_new_n4190__), .dout(new_new_n2886__));
  and1  g0921(.dina(new_new_n4189__), .dinb(new_new_n4190__), .dout(new_new_n2887__));
  or1   g0922(.dina(new_new_n4187__), .dinb(new_new_n4188__), .dout(new_new_n2888__));
  and1  g0923(.dina(new_new_n2888__), .dinb(new_new_n2886__), .dout(new_new_n2889__));
  or1   g0924(.dina(new_new_n2887__), .dinb(new_new_n2885__), .dout(new_new_n2890__));
  and1  g0925(.dina(new_new_n4191__), .dinb(new_new_n4192__), .dout(new_new_n2891__));
  or1   g0926(.dina(new_new_n4193__), .dinb(new_new_n4194__), .dout(new_new_n2892__));
  and1  g0927(.dina(new_new_n4193__), .dinb(new_new_n4194__), .dout(new_new_n2893__));
  or1   g0928(.dina(new_new_n4191__), .dinb(new_new_n4192__), .dout(new_new_n2894__));
  and1  g0929(.dina(new_new_n2894__), .dinb(new_new_n2892__), .dout(new_new_n2895__));
  or1   g0930(.dina(new_new_n2893__), .dinb(new_new_n2891__), .dout(new_new_n2896__));
  or1   g0931(.dina(new_new_n2896__), .dinb(new_new_n2889__), .dout(new_new_n2897__));
  or1   g0932(.dina(new_new_n2895__), .dinb(new_new_n2890__), .dout(new_new_n2898__));
  and1  g0933(.dina(new_new_n2898__), .dinb(new_new_n2897__), .dout(new_new_n2899__));
  and1  g0934(.dina(new_new_n2646__), .dinb(new_new_n2381__), .dout(new_new_n2900__));
  and1  g0935(.dina(new_new_n2555__), .dinb(new_new_n2358__), .dout(new_new_n2901__));
  and1  g0936(.dina(new_new_n2638__), .dinb(new_new_n2291__), .dout(new_new_n2902__));
  or1   g0937(.dina(new_new_n2902__), .dinb(new_new_n2901__), .dout(new_new_n2903__));
  or1   g0938(.dina(new_new_n2903__), .dinb(new_new_n2900__), .dout(new_new_n2904__));
  and1  g0939(.dina(new_new_n2643__), .dinb(new_new_n2332__), .dout(new_new_n2905__));
  and1  g0940(.dina(new_new_n2552__), .dinb(new_new_n2365__), .dout(new_new_n2906__));
  or1   g0941(.dina(new_new_n2906__), .dinb(new_new_n2905__), .dout(new_new_n2907__));
  and1  g0942(.dina(new_new_n2557__), .dinb(new_new_n2372__), .dout(new_new_n2908__));
  and1  g0943(.dina(new_new_n2642__), .dinb(new_new_n2333__), .dout(new_new_n2909__));
  or1   g0944(.dina(new_new_n2909__), .dinb(new_new_n2908__), .dout(new_new_n2910__));
  or1   g0945(.dina(new_new_n2910__), .dinb(new_new_n2907__), .dout(new_new_n2911__));
  and1  g0946(.dina(new_new_n2546__), .dinb(new_new_n2279__), .dout(new_new_n2912__));
  and1  g0947(.dina(new_new_n2639__), .dinb(new_new_n2290__), .dout(new_new_n2913__));
  or1   g0948(.dina(new_new_n2913__), .dinb(new_new_n2912__), .dout(new_new_n2914__));
  and1  g0949(.dina(new_new_n2548__), .dinb(new_new_n2325__), .dout(new_new_n2915__));
  and1  g0950(.dina(new_new_n2647__), .dinb(new_new_n2380__), .dout(new_new_n2916__));
  or1   g0951(.dina(new_new_n2916__), .dinb(new_new_n2915__), .dout(new_new_n2917__));
  or1   g0952(.dina(new_new_n2917__), .dinb(new_new_n2914__), .dout(new_new_n2918__));
  or1   g0953(.dina(new_new_n2918__), .dinb(new_new_n2911__), .dout(new_new_n2919__));
  or1   g0954(.dina(new_new_n2919__), .dinb(new_new_n2904__), .dout(new_new_n2920__));
  and1  g0955(.dina(new_new_n2551__), .dinb(new_new_n2310__), .dout(new_new_n2921__));
  and1  g0956(.dina(new_new_n2581__), .dinb(new_new_n2579__), .dout(new_new_n2922__));
  or1   g0957(.dina(new_new_n2922__), .dinb(new_new_n1747__), .dout(new_new_n2923__));
  or1   g0958(.dina(new_new_n2923__), .dinb(new_new_n2921__), .dout(new_new_n2924__));
  and1  g0959(.dina(new_new_n2644__), .dinb(new_new_n2353__), .dout(new_new_n2925__));
  and1  g0960(.dina(new_new_n2645__), .dinb(new_new_n2352__), .dout(new_new_n2926__));
  or1   g0961(.dina(new_new_n2926__), .dinb(new_new_n2925__), .dout(new_new_n2927__));
  and1  g0962(.dina(new_new_n2649__), .dinb(new_new_n2338__), .dout(new_new_n2928__));
  and1  g0963(.dina(new_new_n2648__), .dinb(new_new_n2339__), .dout(new_new_n2929__));
  or1   g0964(.dina(new_new_n2929__), .dinb(new_new_n2928__), .dout(new_new_n2930__));
  or1   g0965(.dina(new_new_n2930__), .dinb(new_new_n2927__), .dout(new_new_n2931__));
  or1   g0966(.dina(new_new_n2931__), .dinb(new_new_n2924__), .dout(new_new_n2932__));
  or1   g0967(.dina(new_new_n2614__), .dinb(new_new_n2610__), .dout(new_new_n2933__));
  or1   g0968(.dina(new_new_n2616__), .dinb(new_new_n2592__), .dout(new_new_n2934__));
  or1   g0969(.dina(new_new_n2934__), .dinb(new_new_n2933__), .dout(new_new_n2935__));
  or1   g0970(.dina(new_new_n2622__), .dinb(new_new_n2594__), .dout(new_new_n2936__));
  or1   g0971(.dina(new_new_n2624__), .dinb(new_new_n2598__), .dout(new_new_n2937__));
  or1   g0972(.dina(new_new_n2937__), .dinb(new_new_n2936__), .dout(new_new_n2938__));
  or1   g0973(.dina(new_new_n2938__), .dinb(new_new_n2935__), .dout(new_new_n2939__));
  or1   g0974(.dina(new_new_n2602__), .dinb(new_new_n2600__), .dout(new_new_n2940__));
  or1   g0975(.dina(new_new_n2626__), .dinb(new_new_n2596__), .dout(new_new_n2941__));
  or1   g0976(.dina(new_new_n2941__), .dinb(new_new_n2940__), .dout(new_new_n2942__));
  or1   g0977(.dina(new_new_n2608__), .dinb(new_new_n2606__), .dout(new_new_n2943__));
  or1   g0978(.dina(new_new_n2620__), .dinb(new_new_n2604__), .dout(new_new_n2944__));
  or1   g0979(.dina(new_new_n2944__), .dinb(new_new_n2943__), .dout(new_new_n2945__));
  or1   g0980(.dina(new_new_n2945__), .dinb(new_new_n2942__), .dout(new_new_n2946__));
  or1   g0981(.dina(new_new_n2946__), .dinb(new_new_n2939__), .dout(new_new_n2947__));
  or1   g0982(.dina(new_new_n2947__), .dinb(new_new_n2932__), .dout(new_new_n2948__));
  or1   g0983(.dina(new_new_n2948__), .dinb(new_new_n2920__), .dout(new_new_n2949__));
  and1  g0984(.dina(new_new_n4174__), .dinb(new_new_n4183__), .dout(new_new_n2950__));
  or1   g0985(.dina(new_new_n4184__), .dinb(new_new_n2227__), .dout(new_new_n2951__));
  and1  g0986(.dina(new_new_n2950__), .dinb(new_new_n2511__), .dout(new_new_n2952__));
  and1  g0987(.dina(new_new_n2951__), .dinb(new_new_n2510__), .dout(new_new_n2953__));
  or1   g0988(.dina(new_new_n2953__), .dinb(new_new_n2952__), .dout(new_new_n2954__));
  and1  g0989(.dina(new_new_n2954__), .dinb(new_new_n4169__), .dout(new_new_n2955__));
  and1  g0990(.dina(new_new_n4195__), .dinb(new_new_n2252__), .dout(new_new_n2956__));
  or1   g0991(.dina(new_new_n2956__), .dinb(new_new_n2955__), .dout(new_new_n2957__));
  or1   g0992(.dina(new_new_n2690__), .dinb(new_new_n2682__), .dout(new_new_n2958__));
  or1   g0993(.dina(new_new_n2691__), .dinb(new_new_n2683__), .dout(new_new_n2959__));
  and1  g0994(.dina(new_new_n2959__), .dinb(new_new_n4196__), .dout(new_new_n2960__));
  and1  g0995(.dina(new_new_n2960__), .dinb(new_new_n2958__), .dout(new_new_n2961__));
  or1   g0996(.dina(new_new_n4195__), .dinb(new_new_n4177__), .dout(new_new_n2962__));
  and1  g0997(.dina(new_new_n2689__), .dinb(new_new_n2687__), .dout(new_new_n2963__));
  or1   g0998(.dina(new_new_n2688__), .dinb(new_new_n2686__), .dout(new_new_n2964__));
  and1  g0999(.dina(new_new_n4197__), .dinb(new_new_n4198__), .dout(new_new_n2965__));
  or1   g1000(.dina(new_new_n4186__), .dinb(new_new_n4199__), .dout(new_new_n2966__));
  and1  g1001(.dina(new_new_n4185__), .dinb(new_new_n4199__), .dout(new_new_n2967__));
  or1   g1002(.dina(new_new_n4197__), .dinb(new_new_n4198__), .dout(new_new_n2968__));
  and1  g1003(.dina(new_new_n2968__), .dinb(new_new_n2966__), .dout(new_new_n2969__));
  or1   g1004(.dina(new_new_n2967__), .dinb(new_new_n2965__), .dout(new_new_n2970__));
  or1   g1005(.dina(new_new_n2969__), .dinb(new_new_n4200__), .dout(new_new_n2971__));
  or1   g1006(.dina(new_new_n2970__), .dinb(new_new_n4201__), .dout(new_new_n2972__));
  and1  g1007(.dina(new_new_n2972__), .dinb(new_new_n2971__), .dout(new_new_n2973__));
  or1   g1008(.dina(new_new_n2973__), .dinb(new_new_n4181__), .dout(new_new_n2974__));
  and1  g1009(.dina(new_new_n2974__), .dinb(new_new_n2962__), .dout(new_new_n2975__));
  and1  g1010(.dina(new_new_n2677__), .dinb(new_new_n2674__), .dout(new_new_n2976__));
  or1   g1011(.dina(new_new_n2676__), .dinb(new_new_n2675__), .dout(new_new_n2977__));
  or1   g1012(.dina(new_new_n2977__), .dinb(new_new_n4200__), .dout(new_new_n2978__));
  or1   g1013(.dina(new_new_n2976__), .dinb(new_new_n4201__), .dout(new_new_n2979__));
  and1  g1014(.dina(new_new_n2979__), .dinb(new_new_n4196__), .dout(new_new_n2980__));
  and1  g1015(.dina(new_new_n2980__), .dinb(new_new_n2978__), .dout(new_new_n2981__));
  or1   g1016(.dina(new_new_n2559__), .dinb(new_new_n2538__), .dout(new_new_n2982__));
  or1   g1017(.dina(new_new_n2666__), .dinb(new_new_n2640__), .dout(new_new_n2983__));
  and1  g1018(.dina(new_new_n2983__), .dinb(new_new_n2982__), .dout(new_new_n2984__));
  or1   g1019(.dina(new_new_n2632__), .dinb(new_new_n2618__), .dout(new_new_n2985__));
  or1   g1020(.dina(new_new_n2634__), .dinb(new_new_n2612__), .dout(new_new_n2986__));
  or1   g1021(.dina(new_new_n2986__), .dinb(new_new_n4202__), .dout(new_new_n2987__));
  or1   g1022(.dina(new_new_n2987__), .dinb(new_new_n2984__), .dout(new_new_n2988__));
  or1   g1023(.dina(new_new_n4202__), .dinb(new_new_n2613__), .dout(new_new_n2989__));
  and1  g1024(.dina(new_new_n2989__), .dinb(new_new_n2619__), .dout(new_new_n2990__));
  and1  g1025(.dina(new_new_n2990__), .dinb(new_new_n2988__), .dout(new_new_n2991__));
  or1   g1026(.dina(new_new_n2664__), .dinb(new_new_n2662__), .dout(new_new_n2992__));
  or1   g1027(.dina(new_new_n4203__), .dinb(new_new_n4204__), .dout(new_new_n2993__));
  or1   g1028(.dina(new_new_n2660__), .dinb(new_new_n2658__), .dout(new_new_n2994__));
  and1  g1029(.dina(new_new_n2544__), .dinb(new_new_n2541__), .dout(new_new_n2995__));
  or1   g1030(.dina(new_new_n2995__), .dinb(new_new_n2654__), .dout(new_new_n2996__));
  or1   g1031(.dina(new_new_n2996__), .dinb(new_new_n4205__), .dout(new_new_n2997__));
  or1   g1032(.dina(new_new_n2997__), .dinb(new_new_n4206__), .dout(new_new_n2998__));
  or1   g1033(.dina(new_new_n2998__), .dinb(new_new_n2991__), .dout(new_new_n2999__));
  or1   g1034(.dina(new_new_n4204__), .dinb(new_new_n2655__), .dout(new_new_n3000__));
  or1   g1035(.dina(new_new_n3000__), .dinb(new_new_n4205__), .dout(new_new_n3001__));
  and1  g1036(.dina(new_new_n3001__), .dinb(new_new_n2561__), .dout(new_new_n3002__));
  or1   g1037(.dina(new_new_n3002__), .dinb(new_new_n4203__), .dout(new_new_n3003__));
  or1   g1038(.dina(new_new_n4206__), .dinb(new_new_n2659__), .dout(new_new_n3004__));
  and1  g1039(.dina(new_new_n3004__), .dinb(new_new_n2663__), .dout(new_new_n3005__));
  and1  g1040(.dina(new_new_n3005__), .dinb(new_new_n3003__), .dout(new_new_n3006__));
  and1  g1041(.dina(new_new_n3006__), .dinb(new_new_n2999__), .dout(new_new_n3007__));
  or1   g1042(.dina(new_new_n4207__), .dinb(new_new_n4208__), .dout(new_new_n3008__));
  or1   g1043(.dina(new_new_n3008__), .dinb(new_new_n4209__), .dout(new_new_n3009__));
  or1   g1044(.dina(new_new_n4210__), .dinb(new_new_n4172__), .dout(new_new_n3010__));
  or1   g1045(.dina(new_new_n3010__), .dinb(new_new_n4211__), .dout(new_new_n3011__));
  or1   g1046(.dina(new_new_n3011__), .dinb(new_new_n3009__), .dout(new_new_n3012__));
  and1  g1047(.dina(new_new_n2702__), .dinb(new_new_n4213__), .dout(new_new_n3013__));
  or1   g1048(.dina(new_new_n2703__), .dinb(new_new_n4216__), .dout(new_new_n3014__));
  and1  g1049(.dina(new_new_n2754__), .dinb(new_new_n4220__), .dout(new_new_n3015__));
  or1   g1050(.dina(new_new_n2755__), .dinb(new_new_n4227__), .dout(new_new_n3016__));
  and1  g1051(.dina(new_new_n2760__), .dinb(new_new_n4227__), .dout(new_new_n3017__));
  or1   g1052(.dina(new_new_n2761__), .dinb(new_new_n4220__), .dout(new_new_n3018__));
  and1  g1053(.dina(new_new_n2773__), .dinb(new_new_n2744__), .dout(new_new_n3019__));
  or1   g1054(.dina(new_new_n2772__), .dinb(new_new_n2745__), .dout(new_new_n3020__));
  and1  g1055(.dina(new_new_n2777__), .dinb(new_new_n2747__), .dout(new_new_n3021__));
  or1   g1056(.dina(new_new_n2776__), .dinb(new_new_n2746__), .dout(new_new_n3022__));
  and1  g1057(.dina(new_new_n4213__), .dinb(new_new_n1942__), .dout(new_new_n3023__));
  or1   g1058(.dina(new_new_n4216__), .dinb(new_new_n1943__), .dout(new_new_n3024__));
  and1  g1059(.dina(new_new_n4233__), .dinb(new_new_n4235__), .dout(new_new_n3025__));
  or1   g1060(.dina(new_new_n4237__), .dinb(new_new_n4239__), .dout(new_new_n3026__));
  and1  g1061(.dina(new_new_n3020__), .dinb(new_new_n3014__), .dout(new_new_n3027__));
  or1   g1062(.dina(new_new_n4240__), .dinb(new_new_n4241__), .dout(new_new_n3028__));
  and1  g1063(.dina(new_new_n2731__), .dinb(new_new_n4244__), .dout(new_new_n3029__));
  or1   g1064(.dina(new_new_n2730__), .dinb(new_new_n4249__), .dout(new_new_n3030__));
  and1  g1065(.dina(new_new_n2743__), .dinb(new_new_n2737__), .dout(new_new_n3031__));
  or1   g1066(.dina(new_new_n2742__), .dinb(new_new_n2736__), .dout(new_new_n3032__));
  and1  g1067(.dina(new_new_n3031__), .dinb(new_new_n3030__), .dout(new_new_n3033__));
  or1   g1068(.dina(new_new_n3032__), .dinb(new_new_n3029__), .dout(new_new_n3034__));
  and1  g1069(.dina(new_new_n2693__), .dinb(new_new_n2637__), .dout(new_new_n3035__));
  or1   g1070(.dina(new_new_n2692__), .dinb(new_new_n2636__), .dout(new_new_n3036__));
  and1  g1071(.dina(new_new_n3034__), .dinb(new_new_n3024__), .dout(new_new_n3037__));
  or1   g1072(.dina(new_new_n4252__), .dinb(new_new_n4253__), .dout(new_new_n3038__));
  and1  g1073(.dina(new_new_n2740__), .dinb(new_new_n2739__), .dout(new_new_n3039__));
  or1   g1074(.dina(new_new_n2741__), .dinb(new_new_n2738__), .dout(new_new_n3040__));
  and1  g1075(.dina(new_new_n3040__), .dinb(new_new_n4254__), .dout(new_new_n3041__));
  or1   g1076(.dina(new_new_n3039__), .dinb(new_new_n4255__), .dout(new_new_n3042__));
  and1  g1077(.dina(new_new_n2705__), .dinb(new_new_n4249__), .dout(new_new_n3043__));
  or1   g1078(.dina(new_new_n2704__), .dinb(new_new_n4244__), .dout(new_new_n3044__));
  and1  g1079(.dina(new_new_n3043__), .dinb(new_new_n4255__), .dout(new_new_n3045__));
  or1   g1080(.dina(new_new_n3044__), .dinb(new_new_n4254__), .dout(new_new_n3046__));
  and1  g1081(.dina(new_new_n3046__), .dinb(new_new_n3042__), .dout(new_new_n3047__));
  or1   g1082(.dina(new_new_n3045__), .dinb(new_new_n3041__), .dout(new_new_n3048__));
  and1  g1083(.dina(new_new_n2735__), .dinb(new_new_n2725__), .dout(new_new_n3049__));
  or1   g1084(.dina(new_new_n2734__), .dinb(new_new_n2724__), .dout(new_new_n3050__));
  and1  g1085(.dina(new_new_n3050__), .dinb(new_new_n4250__), .dout(new_new_n3051__));
  or1   g1086(.dina(new_new_n3049__), .dinb(new_new_n4245__), .dout(new_new_n3052__));
  and1  g1087(.dina(new_new_n2700__), .dinb(new_new_n4214__), .dout(new_new_n3053__));
  or1   g1088(.dina(new_new_n2701__), .dinb(new_new_n4217__), .dout(new_new_n3054__));
  and1  g1089(.dina(new_new_n2728__), .dinb(new_new_n4245__), .dout(new_new_n3055__));
  or1   g1090(.dina(new_new_n2729__), .dinb(new_new_n4250__), .dout(new_new_n3056__));
  and1  g1091(.dina(new_new_n3056__), .dinb(new_new_n3054__), .dout(new_new_n3057__));
  or1   g1092(.dina(new_new_n3055__), .dinb(new_new_n3053__), .dout(new_new_n3058__));
  and1  g1093(.dina(new_new_n3057__), .dinb(new_new_n3052__), .dout(new_new_n3059__));
  or1   g1094(.dina(new_new_n3058__), .dinb(new_new_n3051__), .dout(new_new_n3060__));
  and1  g1095(.dina(new_new_n2733__), .dinb(new_new_n2723__), .dout(new_new_n3061__));
  or1   g1096(.dina(new_new_n2732__), .dinb(new_new_n2722__), .dout(new_new_n3062__));
  and1  g1097(.dina(new_new_n3062__), .dinb(new_new_n4251__), .dout(new_new_n3063__));
  or1   g1098(.dina(new_new_n3061__), .dinb(new_new_n4246__), .dout(new_new_n3064__));
  and1  g1099(.dina(new_new_n2698__), .dinb(new_new_n4214__), .dout(new_new_n3065__));
  or1   g1100(.dina(new_new_n2699__), .dinb(new_new_n4217__), .dout(new_new_n3066__));
  and1  g1101(.dina(new_new_n2726__), .dinb(new_new_n4246__), .dout(new_new_n3067__));
  or1   g1102(.dina(new_new_n2727__), .dinb(new_new_n4251__), .dout(new_new_n3068__));
  and1  g1103(.dina(new_new_n3068__), .dinb(new_new_n3066__), .dout(new_new_n3069__));
  or1   g1104(.dina(new_new_n3067__), .dinb(new_new_n3065__), .dout(new_new_n3070__));
  and1  g1105(.dina(new_new_n3069__), .dinb(new_new_n3064__), .dout(new_new_n3071__));
  or1   g1106(.dina(new_new_n3070__), .dinb(new_new_n3063__), .dout(new_new_n3072__));
  and1  g1107(.dina(new_new_n4257__), .dinb(new_new_n4258__), .dout(new_new_n3073__));
  or1   g1108(.dina(new_new_n4259__), .dinb(new_new_n4261__), .dout(new_new_n3074__));
  and1  g1109(.dina(new_new_n4259__), .dinb(new_new_n4261__), .dout(new_new_n3075__));
  or1   g1110(.dina(new_new_n4257__), .dinb(new_new_n4258__), .dout(new_new_n3076__));
  and1  g1111(.dina(new_new_n3076__), .dinb(new_new_n3074__), .dout(new_new_n3077__));
  or1   g1112(.dina(new_new_n3075__), .dinb(new_new_n3073__), .dout(new_new_n3078__));
  or1   g1113(.dina(new_new_n4263__), .dinb(new_new_n4265__), .dout(new_new_n3079__));
  and1  g1114(.dina(new_new_n2706__), .dinb(new_new_n4267__), .dout(new_new_n3080__));
  or1   g1115(.dina(new_new_n2707__), .dinb(new_new_n4270__), .dout(new_new_n3081__));
  and1  g1116(.dina(new_new_n2712__), .dinb(new_new_n4270__), .dout(new_new_n3082__));
  or1   g1117(.dina(new_new_n2713__), .dinb(new_new_n4267__), .dout(new_new_n3083__));
  and1  g1118(.dina(new_new_n3083__), .dinb(new_new_n3081__), .dout(new_new_n3084__));
  or1   g1119(.dina(new_new_n3082__), .dinb(new_new_n3080__), .dout(new_new_n3085__));
  and1  g1120(.dina(new_new_n3085__), .dinb(new_new_n4221__), .dout(new_new_n3086__));
  or1   g1121(.dina(new_new_n3084__), .dinb(new_new_n4228__), .dout(new_new_n3087__));
  and1  g1122(.dina(new_new_n2708__), .dinb(new_new_n4268__), .dout(new_new_n3088__));
  or1   g1123(.dina(new_new_n2709__), .dinb(new_new_n4271__), .dout(new_new_n3089__));
  and1  g1124(.dina(new_new_n2710__), .dinb(new_new_n4271__), .dout(new_new_n3090__));
  or1   g1125(.dina(new_new_n2711__), .dinb(new_new_n4268__), .dout(new_new_n3091__));
  and1  g1126(.dina(new_new_n3091__), .dinb(new_new_n3089__), .dout(new_new_n3092__));
  or1   g1127(.dina(new_new_n3090__), .dinb(new_new_n3088__), .dout(new_new_n3093__));
  and1  g1128(.dina(new_new_n3093__), .dinb(new_new_n4228__), .dout(new_new_n3094__));
  or1   g1129(.dina(new_new_n3092__), .dinb(new_new_n4221__), .dout(new_new_n3095__));
  and1  g1130(.dina(new_new_n3095__), .dinb(new_new_n3087__), .dout(new_new_n3096__));
  or1   g1131(.dina(new_new_n3094__), .dinb(new_new_n3086__), .dout(new_new_n3097__));
  and1  g1132(.dina(new_new_n2815__), .dinb(new_new_n2794__), .dout(new_new_n3098__));
  or1   g1133(.dina(new_new_n4272__), .dinb(new_new_n2795__), .dout(new_new_n3099__));
  and1  g1134(.dina(new_new_n4273__), .dinb(new_new_n2805__), .dout(new_new_n3100__));
  or1   g1135(.dina(new_new_n2817__), .dinb(new_new_n2804__), .dout(new_new_n3101__));
  and1  g1136(.dina(new_new_n4274__), .dinb(new_new_n4275__), .dout(new_new_n3102__));
  or1   g1137(.dina(new_new_n3101__), .dinb(new_new_n3099__), .dout(new_new_n3103__));
  or1   g1138(.dina(new_new_n4277__), .dinb(new_new_n4279__), .dout(new_new_n3104__));
  and1  g1139(.dina(new_new_n2529__), .dinb(new_new_n2526__), .dout(new_new_n3105__));
  or1   g1140(.dina(new_new_n2528__), .dinb(new_new_n2527__), .dout(new_new_n3106__));
  or1   g1141(.dina(new_new_n4282__), .dinb(new_new_n4285__), .dout(new_new_n3107__));
  and1  g1142(.dina(new_new_n4288__), .dinb(new_new_n4290__), .dout(new_new_n3108__));
  and1  g1143(.dina(new_new_n4294__), .dinb(new_new_n1714__), .dout(new_new_n3109__));
  and1  g1144(.dina(new_new_n4301__), .dinb(new_new_n4306__), .dout(new_new_n3110__));
  or1   g1145(.dina(new_new_n3110__), .dinb(new_new_n3109__), .dout(new_new_n3111__));
  and1  g1146(.dina(new_new_n1804__), .dinb(new_new_n4294__), .dout(new_new_n3112__));
  and1  g1147(.dina(new_new_n4312__), .dinb(new_new_n4306__), .dout(new_new_n3113__));
  or1   g1148(.dina(new_new_n3113__), .dinb(new_new_n3112__), .dout(new_new_n3114__));
  and1  g1149(.dina(new_new_n1798__), .dinb(new_new_n4293__), .dout(new_new_n3115__));
  and1  g1150(.dina(new_new_n4314__), .dinb(new_new_n4305__), .dout(new_new_n3116__));
  or1   g1151(.dina(new_new_n3116__), .dinb(new_new_n3115__), .dout(new_new_n3117__));
  and1  g1152(.dina(new_new_n4317__), .dinb(new_new_n1822__), .dout(new_new_n3118__));
  and1  g1153(.dina(new_new_n4323__), .dinb(new_new_n4327__), .dout(new_new_n3119__));
  or1   g1154(.dina(new_new_n3119__), .dinb(new_new_n3118__), .dout(new_new_n3120__));
  and1  g1155(.dina(new_new_n1846__), .dinb(new_new_n4317__), .dout(new_new_n3121__));
  and1  g1156(.dina(new_new_n4333__), .dinb(new_new_n4327__), .dout(new_new_n3122__));
  or1   g1157(.dina(new_new_n3122__), .dinb(new_new_n3121__), .dout(new_new_n3123__));
  and1  g1158(.dina(new_new_n1852__), .dinb(new_new_n4318__), .dout(new_new_n3124__));
  and1  g1159(.dina(new_new_n4335__), .dinb(new_new_n4328__), .dout(new_new_n3125__));
  or1   g1160(.dina(new_new_n3125__), .dinb(new_new_n3124__), .dout(new_new_n3126__));
  and1  g1161(.dina(new_new_n4336__), .dinb(new_new_n2537__), .dout(new_new_n3127__));
  and1  g1162(.dina(new_new_n4338__), .dinb(new_new_n4342__), .dout(new_new_n3128__));
  and1  g1163(.dina(new_new_n4336__), .dinb(new_new_n2536__), .dout(new_new_n3129__));
  and1  g1164(.dina(new_new_n4345__), .dinb(new_new_n4263__), .dout(new_new_n3130__));
  or1   g1165(.dina(new_new_n3130__), .dinb(new_new_n3128__), .dout(new_new_n3131__));
  and1  g1166(.dina(new_new_n2758__), .dinb(new_new_n4223__), .dout(new_new_n3132__));
  or1   g1167(.dina(new_new_n2759__), .dinb(new_new_n4230__), .dout(new_new_n3133__));
  and1  g1168(.dina(new_new_n2764__), .dinb(new_new_n4230__), .dout(new_new_n3134__));
  or1   g1169(.dina(new_new_n2765__), .dinb(new_new_n4223__), .dout(new_new_n3135__));
  and1  g1170(.dina(new_new_n3135__), .dinb(new_new_n3133__), .dout(new_new_n3136__));
  or1   g1171(.dina(new_new_n3134__), .dinb(new_new_n3132__), .dout(new_new_n3137__));
  and1  g1172(.dina(new_new_n4348__), .dinb(new_new_n4288__), .dout(new_new_n3138__));
  or1   g1173(.dina(new_new_n4351__), .dinb(new_new_n4282__), .dout(new_new_n3139__));
  and1  g1174(.dina(new_new_n4287__), .dinb(new_new_n4352__), .dout(new_new_n3140__));
  or1   g1175(.dina(new_new_n4281__), .dinb(new_new_n4354__), .dout(new_new_n3141__));
  or1   g1176(.dina(new_new_n3141__), .dinb(new_new_n3138__), .dout(new_new_n3142__));
  and1  g1177(.dina(new_new_n4357__), .dinb(new_new_n4301__), .dout(new_new_n3143__));
  or1   g1178(.dina(new_new_n4360__), .dinb(new_new_n4361__), .dout(new_new_n3144__));
  and1  g1179(.dina(new_new_n4360__), .dinb(new_new_n4361__), .dout(new_new_n3145__));
  or1   g1180(.dina(new_new_n4357__), .dinb(new_new_n4300__), .dout(new_new_n3146__));
  and1  g1181(.dina(new_new_n3146__), .dinb(new_new_n3144__), .dout(new_new_n3147__));
  or1   g1182(.dina(new_new_n3145__), .dinb(new_new_n3143__), .dout(new_new_n3148__));
  and1  g1183(.dina(new_new_n3147__), .dinb(new_new_n4362__), .dout(new_new_n3149__));
  and1  g1184(.dina(new_new_n3148__), .dinb(new_new_n3077__), .dout(new_new_n3150__));
  or1   g1185(.dina(new_new_n3150__), .dinb(new_new_n3149__), .dout(new_new_n3151__));
  or1   g1186(.dina(new_new_n2810__), .dinb(new_new_n2806__), .dout(new_new_n3152__));
  and1  g1187(.dina(new_new_n3152__), .dinb(new_new_n4366__), .dout(new_new_n3153__));
  and1  g1188(.dina(new_new_n4375__), .dinb(new_new_n2798__), .dout(new_new_n3154__));
  and1  g1189(.dina(new_new_n2808__), .dinb(new_new_n4379__), .dout(new_new_n3155__));
  or1   g1190(.dina(new_new_n3155__), .dinb(new_new_n3154__), .dout(new_new_n3156__));
  or1   g1191(.dina(new_new_n3156__), .dinb(new_new_n3153__), .dout(new_new_n3157__));
  and1  g1192(.dina(new_new_n2802__), .dinb(new_new_n4384__), .dout(new_new_n3158__));
  and1  g1193(.dina(new_new_n2796__), .dinb(new_new_n4393__), .dout(new_new_n3159__));
  or1   g1194(.dina(new_new_n3159__), .dinb(new_new_n3158__), .dout(new_new_n3160__));
  and1  g1195(.dina(new_new_n3160__), .dinb(new_new_n4366__), .dout(new_new_n3161__));
  and1  g1196(.dina(new_new_n4375__), .dinb(new_new_n2792__), .dout(new_new_n3162__));
  and1  g1197(.dina(new_new_n2800__), .dinb(new_new_n4393__), .dout(new_new_n3163__));
  and1  g1198(.dina(new_new_n3163__), .dinb(new_new_n4379__), .dout(new_new_n3164__));
  or1   g1199(.dina(new_new_n3164__), .dinb(new_new_n3162__), .dout(new_new_n3165__));
  or1   g1200(.dina(new_new_n3165__), .dinb(new_new_n3161__), .dout(new_new_n3166__));
  and1  g1201(.dina(new_new_n4318__), .dinb(new_new_n1828__), .dout(new_new_n3167__));
  and1  g1202(.dina(new_new_n4405__), .dinb(new_new_n4328__), .dout(new_new_n3168__));
  and1  g1203(.dina(new_new_n4406__), .dinb(new_new_n4407__), .dout(new_new_n3169__));
  and1  g1204(.dina(new_new_n4408__), .dinb(new_new_n4409__), .dout(new_new_n3170__));
  and1  g1205(.dina(new_new_n4410__), .dinb(new_new_n4411__), .dout(new_new_n3171__));
  and1  g1206(.dina(new_new_n4412__), .dinb(new_new_n4413__), .dout(new_new_n3172__));
  or1   g1207(.dina(new_new_n4302__), .dinb(new_new_n4414__), .dout(new_new_n3173__));
  and1  g1208(.dina(new_new_n1774__), .dinb(new_new_n4295__), .dout(new_new_n3174__));
  and1  g1209(.dina(new_new_n4262__), .dinb(new_new_n4307__), .dout(new_new_n3175__));
  or1   g1210(.dina(new_new_n3175__), .dinb(new_new_n3174__), .dout(new_new_n3176__));
  or1   g1211(.dina(new_new_n4415__), .dinb(new_new_n4417__), .dout(new_new_n3177__));
  and1  g1212(.dina(new_new_n4415__), .dinb(new_new_n4417__), .dout(new_new_n3178__));
  or1   g1213(.dina(new_new_n4419__), .dinb(new_new_n4421__), .dout(new_new_n3179__));
  and1  g1214(.dina(new_new_n1780__), .dinb(new_new_n4295__), .dout(new_new_n3180__));
  and1  g1215(.dina(new_new_n4358__), .dinb(new_new_n4307__), .dout(new_new_n3181__));
  or1   g1216(.dina(new_new_n3181__), .dinb(new_new_n3180__), .dout(new_new_n3182__));
  or1   g1217(.dina(new_new_n4422__), .dinb(new_new_n4424__), .dout(new_new_n3183__));
  and1  g1218(.dina(new_new_n4422__), .dinb(new_new_n4424__), .dout(new_new_n3184__));
  and1  g1219(.dina(new_new_n1786__), .dinb(new_new_n4297__), .dout(new_new_n3185__));
  and1  g1220(.dina(new_new_n4427__), .dinb(new_new_n4309__), .dout(new_new_n3186__));
  or1   g1221(.dina(new_new_n3186__), .dinb(new_new_n3185__), .dout(new_new_n3187__));
  and1  g1222(.dina(new_new_n4429__), .dinb(new_new_n4431__), .dout(new_new_n3188__));
  or1   g1223(.dina(new_new_n4429__), .dinb(new_new_n4431__), .dout(new_new_n3189__));
  and1  g1224(.dina(new_new_n1792__), .dinb(new_new_n4297__), .dout(new_new_n3190__));
  and1  g1225(.dina(new_new_n4277__), .dinb(new_new_n4309__), .dout(new_new_n3191__));
  or1   g1226(.dina(new_new_n3191__), .dinb(new_new_n3190__), .dout(new_new_n3192__));
  and1  g1227(.dina(new_new_n4433__), .dinb(new_new_n4342__), .dout(new_new_n3193__));
  or1   g1228(.dina(new_new_n4433__), .dinb(new_new_n4341__), .dout(new_new_n3194__));
  and1  g1229(.dina(new_new_n4434__), .dinb(new_new_n4436__), .dout(new_new_n3195__));
  and1  g1230(.dina(new_new_n4338__), .dinb(new_new_n4436__), .dout(new_new_n3196__));
  and1  g1231(.dina(new_new_n4298__), .dinb(new_new_n1726__), .dout(new_new_n3197__));
  and1  g1232(.dina(new_new_n4439__), .dinb(new_new_n4310__), .dout(new_new_n3198__));
  or1   g1233(.dina(new_new_n3198__), .dinb(new_new_n3197__), .dout(new_new_n3199__));
  and1  g1234(.dina(new_new_n4440__), .dinb(new_new_n4442__), .dout(new_new_n3200__));
  or1   g1235(.dina(new_new_n4440__), .dinb(new_new_n4442__), .dout(new_new_n3201__));
  and1  g1236(.dina(new_new_n4339__), .dinb(new_new_n4443__), .dout(new_new_n3202__));
  or1   g1237(.dina(new_new_n4444__), .dinb(new_new_n4445__), .dout(new_new_n3203__));
  and1  g1238(.dina(new_new_n4446__), .dinb(new_new_n4239__), .dout(new_new_n3204__));
  or1   g1239(.dina(new_new_n4447__), .dinb(new_new_n4237__), .dout(new_new_n3205__));
  and1  g1240(.dina(new_new_n4448__), .dinb(new_new_n4265__), .dout(new_new_n3206__));
  and1  g1241(.dina(new_new_n2395__), .dinb(new_new_n4449__), .dout(new_new_n3207__));
  and1  g1242(.dina(new_new_n4450__), .dinb(new_new_n2387__), .dout(new_new_n3208__));
  and1  g1243(.dina(new_new_n4345__), .dinb(new_new_n4451__), .dout(new_new_n3209__));
  and1  g1244(.dina(new_new_n4346__), .dinb(new_new_n4452__), .dout(new_new_n3210__));
  or1   g1245(.dina(new_new_n2813__), .dinb(new_new_n1951__), .dout(new_new_n3211__));
  and1  g1246(.dina(new_new_n4298__), .dinb(new_new_n1720__), .dout(new_new_n3212__));
  and1  g1247(.dina(new_new_n4454__), .dinb(new_new_n4310__), .dout(new_new_n3213__));
  or1   g1248(.dina(new_new_n3213__), .dinb(new_new_n3212__), .dout(new_new_n3214__));
  or1   g1249(.dina(new_new_n4456__), .dinb(new_new_n4457__), .dout(new_new_n3215__));
  and1  g1250(.dina(new_new_n4320__), .dinb(new_new_n1810__), .dout(new_new_n3216__));
  and1  g1251(.dina(new_new_n4459__), .dinb(new_new_n4330__), .dout(new_new_n3217__));
  or1   g1252(.dina(new_new_n3217__), .dinb(new_new_n3216__), .dout(new_new_n3218__));
  and1  g1253(.dina(new_new_n4320__), .dinb(new_new_n1816__), .dout(new_new_n3219__));
  and1  g1254(.dina(new_new_n2756__), .dinb(new_new_n4224__), .dout(new_new_n3220__));
  or1   g1255(.dina(new_new_n2757__), .dinb(new_new_n4231__), .dout(new_new_n3221__));
  and1  g1256(.dina(new_new_n2762__), .dinb(new_new_n4231__), .dout(new_new_n3222__));
  or1   g1257(.dina(new_new_n2763__), .dinb(new_new_n4224__), .dout(new_new_n3223__));
  and1  g1258(.dina(new_new_n3223__), .dinb(new_new_n3221__), .dout(new_new_n3224__));
  or1   g1259(.dina(new_new_n3222__), .dinb(new_new_n3220__), .dout(new_new_n3225__));
  and1  g1260(.dina(new_new_n4461__), .dinb(new_new_n4330__), .dout(new_new_n3226__));
  or1   g1261(.dina(new_new_n3226__), .dinb(new_new_n3219__), .dout(new_new_n3227__));
  and1  g1262(.dina(new_new_n1858__), .dinb(new_new_n4321__), .dout(new_new_n3228__));
  and1  g1263(.dina(new_new_n3018__), .dinb(new_new_n3016__), .dout(new_new_n3229__));
  or1   g1264(.dina(new_new_n4463__), .dinb(new_new_n4464__), .dout(new_new_n3230__));
  and1  g1265(.dina(new_new_n4466__), .dinb(new_new_n4331__), .dout(new_new_n3231__));
  or1   g1266(.dina(new_new_n3231__), .dinb(new_new_n3228__), .dout(new_new_n3232__));
  and1  g1267(.dina(new_new_n1840__), .dinb(new_new_n4321__), .dout(new_new_n3233__));
  and1  g1268(.dina(new_new_n4348__), .dinb(new_new_n4331__), .dout(new_new_n3234__));
  or1   g1269(.dina(new_new_n3234__), .dinb(new_new_n3233__), .dout(new_new_n3235__));
  and1  g1270(.dina(new_new_n4467__), .dinb(new_new_n4432__), .dout(new_new_n3236__));
  and1  g1271(.dina(new_new_n2569__), .dinb(new_new_n2296__), .dout(new_new_n3237__));
  or1   g1272(.dina(new_new_n3237__), .dinb(new_new_n3236__), .dout(new_new_n3238__));
  and1  g1273(.dina(new_new_n4445__), .dinb(new_new_n2316__), .dout(new_new_n3239__));
  and1  g1274(.dina(new_new_n4285__), .dinb(new_new_n4443__), .dout(new_new_n3240__));
  or1   g1275(.dina(new_new_n3240__), .dinb(new_new_n3239__), .dout(new_new_n3241__));
  or1   g1276(.dina(new_new_n4468__), .dinb(new_new_n4469__), .dout(new_new_n3242__));
  and1  g1277(.dina(new_new_n4352__), .dinb(new_new_n4470__), .dout(new_new_n3243__));
  and1  g1278(.dina(new_new_n4354__), .dinb(new_new_n4471__), .dout(new_new_n3244__));
  or1   g1279(.dina(new_new_n3244__), .dinb(new_new_n3243__), .dout(new_new_n3245__));
  or1   g1280(.dina(new_new_n4283__), .dinb(new_new_n4473__), .dout(new_new_n3246__));
  and1  g1281(.dina(new_new_n4289__), .dinb(new_new_n4471__), .dout(new_new_n3247__));
  and1  g1282(.dina(new_new_n4474__), .dinb(new_new_n4475__), .dout(new_new_n3248__));
  or1   g1283(.dina(new_new_n4474__), .dinb(new_new_n4475__), .dout(new_new_n3249__));
  or1   g1284(.dina(new_new_n4461__), .dinb(new_new_n4283__), .dout(new_new_n3250__));
  and1  g1285(.dina(new_new_n4289__), .dinb(new_new_n4477__), .dout(new_new_n3251__));
  and1  g1286(.dina(new_new_n4478__), .dinb(new_new_n4479__), .dout(new_new_n3252__));
  or1   g1287(.dina(new_new_n4478__), .dinb(new_new_n4479__), .dout(new_new_n3253__));
  or1   g1288(.dina(new_new_n4427__), .dinb(new_new_n4279__), .dout(new_new_n3254__));
  and1  g1289(.dina(new_new_n4339__), .dinb(new_new_n4432__), .dout(new_new_n3255__));
  and1  g1290(.dina(new_new_n4346__), .dinb(new_new_n4264__), .dout(new_new_n3256__));
  or1   g1291(.dina(new_new_n3256__), .dinb(new_new_n3255__), .dout(new_new_n3257__));
  and1  g1292(.dina(new_new_n4480__), .dinb(new_new_n4481__), .dout(new_new_n3258__));
  or1   g1293(.dina(new_new_n4480__), .dinb(new_new_n4481__), .dout(new_new_n3259__));
  and1  g1294(.dina(new_new_n4482__), .dinb(new_new_n4454__), .dout(new_new_n3260__));
  and1  g1295(.dina(new_new_n4483__), .dinb(new_new_n4358__), .dout(new_new_n3261__));
  and1  g1296(.dina(new_new_n2785__), .dinb(new_new_n2749__), .dout(new_new_n3262__));
  or1   g1297(.dina(new_new_n3262__), .dinb(new_new_n3261__), .dout(new_new_n3263__));
  or1   g1298(.dina(new_new_n4482__), .dinb(new_new_n4455__), .dout(new_new_n3264__));
  or1   g1299(.dina(new_new_n4483__), .dinb(new_new_n4359__), .dout(new_new_n3265__));
  and1  g1300(.dina(new_new_n3265__), .dinb(new_new_n3264__), .dout(new_new_n3266__));
  and1  g1301(.dina(new_new_n3266__), .dinb(new_new_n3263__), .dout(new_new_n3267__));
  or1   g1302(.dina(new_new_n3267__), .dinb(new_new_n3260__), .dout(new_new_n3268__));
  and1  g1303(.dina(new_new_n3268__), .dinb(new_new_n3259__), .dout(new_new_n3269__));
  or1   g1304(.dina(new_new_n3269__), .dinb(new_new_n3258__), .dout(new_new_n3270__));
  or1   g1305(.dina(new_new_n3140__), .dinb(new_new_n3139__), .dout(new_new_n3271__));
  and1  g1306(.dina(new_new_n3271__), .dinb(new_new_n4484__), .dout(new_new_n3272__));
  or1   g1307(.dina(new_new_n4485__), .dinb(new_new_n4486__), .dout(new_new_n3273__));
  and1  g1308(.dina(new_new_n3273__), .dinb(new_new_n4487__), .dout(new_new_n3274__));
  and1  g1309(.dina(new_new_n4236__), .dinb(new_new_n4238__), .dout(new_new_n3275__));
  or1   g1310(.dina(new_new_n4233__), .dinb(new_new_n4235__), .dout(new_new_n3276__));
  and1  g1311(.dina(new_new_n3276__), .dinb(new_new_n3026__), .dout(new_new_n3277__));
  or1   g1312(.dina(new_new_n3275__), .dinb(new_new_n4488__), .dout(new_new_n3278__));
  and1  g1313(.dina(new_new_n4477__), .dinb(new_new_n4489__), .dout(new_new_n3279__));
  or1   g1314(.dina(new_new_n4491__), .dinb(new_new_n4492__), .dout(new_new_n3280__));
  and1  g1315(.dina(new_new_n4491__), .dinb(new_new_n4492__), .dout(new_new_n3281__));
  or1   g1316(.dina(new_new_n4476__), .dinb(new_new_n4489__), .dout(new_new_n3282__));
  and1  g1317(.dina(new_new_n3282__), .dinb(new_new_n3280__), .dout(new_new_n3283__));
  or1   g1318(.dina(new_new_n3281__), .dinb(new_new_n3279__), .dout(new_new_n3284__));
  or1   g1319(.dina(new_new_n3284__), .dinb(new_new_n3277__), .dout(new_new_n3285__));
  or1   g1320(.dina(new_new_n3283__), .dinb(new_new_n3278__), .dout(new_new_n3286__));
  and1  g1321(.dina(new_new_n3286__), .dinb(new_new_n3285__), .dout(new_new_n3287__));
  or1   g1322(.dina(new_new_n4493__), .dinb(new_new_n4494__), .dout(new_new_n3288__));
  and1  g1323(.dina(new_new_n4493__), .dinb(new_new_n4494__), .dout(new_new_n3289__));
  and1  g1324(.dina(new_new_n4495__), .dinb(new_new_n4428__), .dout(new_new_n3290__));
  and1  g1325(.dina(new_new_n3035__), .dinb(new_new_n3027__), .dout(new_new_n3291__));
  or1   g1326(.dina(new_new_n3291__), .dinb(new_new_n3290__), .dout(new_new_n3292__));
  and1  g1327(.dina(new_new_n4496__), .dinb(new_new_n4498__), .dout(new_new_n3293__));
  or1   g1328(.dina(new_new_n4496__), .dinb(new_new_n4498__), .dout(new_new_n3294__));
  and1  g1329(.dina(new_new_n4499__), .dinb(new_new_n4500__), .dout(new_new_n3295__));
  or1   g1330(.dina(new_new_n4501__), .dinb(new_new_n4502__), .dout(new_new_n3296__));
  and1  g1331(.dina(new_new_n4501__), .dinb(new_new_n4502__), .dout(new_new_n3297__));
  or1   g1332(.dina(new_new_n4499__), .dinb(new_new_n4500__), .dout(new_new_n3298__));
  and1  g1333(.dina(new_new_n3298__), .dinb(new_new_n3296__), .dout(new_new_n3299__));
  or1   g1334(.dina(new_new_n3297__), .dinb(new_new_n3295__), .dout(new_new_n3300__));
  and1  g1335(.dina(new_new_n4421__), .dinb(new_new_n4503__), .dout(new_new_n3301__));
  or1   g1336(.dina(new_new_n4505__), .dinb(new_new_n4418__), .dout(new_new_n3302__));
  and1  g1337(.dina(new_new_n4505__), .dinb(new_new_n4418__), .dout(new_new_n3303__));
  or1   g1338(.dina(new_new_n4420__), .dinb(new_new_n4503__), .dout(new_new_n3304__));
  and1  g1339(.dina(new_new_n3304__), .dinb(new_new_n3302__), .dout(new_new_n3305__));
  or1   g1340(.dina(new_new_n3303__), .dinb(new_new_n3301__), .dout(new_new_n3306__));
  and1  g1341(.dina(new_new_n3305__), .dinb(new_new_n3300__), .dout(new_new_n3307__));
  and1  g1342(.dina(new_new_n3306__), .dinb(new_new_n3299__), .dout(new_new_n3308__));
  or1   g1343(.dina(new_new_n3308__), .dinb(new_new_n3307__), .dout(new_new_n3309__));
  and1  g1344(.dina(new_new_n4437__), .dinb(new_new_n4506__), .dout(new_new_n3310__));
  or1   g1345(.dina(new_new_n4508__), .dinb(new_new_n4343__), .dout(new_new_n3311__));
  and1  g1346(.dina(new_new_n4508__), .dinb(new_new_n4343__), .dout(new_new_n3312__));
  or1   g1347(.dina(new_new_n4437__), .dinb(new_new_n4506__), .dout(new_new_n3313__));
  and1  g1348(.dina(new_new_n3313__), .dinb(new_new_n3311__), .dout(new_new_n3314__));
  or1   g1349(.dina(new_new_n3312__), .dinb(new_new_n3310__), .dout(new_new_n3315__));
  and1  g1350(.dina(new_new_n4425__), .dinb(new_new_n4509__), .dout(new_new_n3316__));
  or1   g1351(.dina(new_new_n4510__), .dinb(new_new_n4511__), .dout(new_new_n3317__));
  and1  g1352(.dina(new_new_n4510__), .dinb(new_new_n4511__), .dout(new_new_n3318__));
  or1   g1353(.dina(new_new_n4425__), .dinb(new_new_n4509__), .dout(new_new_n3319__));
  and1  g1354(.dina(new_new_n3319__), .dinb(new_new_n3317__), .dout(new_new_n3320__));
  or1   g1355(.dina(new_new_n3318__), .dinb(new_new_n3316__), .dout(new_new_n3321__));
  and1  g1356(.dina(new_new_n3320__), .dinb(new_new_n3314__), .dout(new_new_n3322__));
  and1  g1357(.dina(new_new_n3321__), .dinb(new_new_n3315__), .dout(new_new_n3323__));
  or1   g1358(.dina(new_new_n3323__), .dinb(new_new_n3322__), .dout(new_new_n3324__));
  and1  g1359(.dina(new_new_n4466__), .dinb(new_new_n4512__), .dout(new_new_n3325__));
  or1   g1360(.dina(new_new_n4513__), .dinb(new_new_n4335__), .dout(new_new_n3326__));
  and1  g1361(.dina(new_new_n4513__), .dinb(new_new_n4334__), .dout(new_new_n3327__));
  or1   g1362(.dina(new_new_n4465__), .dinb(new_new_n4512__), .dout(new_new_n3328__));
  and1  g1363(.dina(new_new_n3328__), .dinb(new_new_n3326__), .dout(new_new_n3329__));
  or1   g1364(.dina(new_new_n3327__), .dinb(new_new_n3325__), .dout(new_new_n3330__));
  or1   g1365(.dina(new_new_n3329__), .dinb(new_new_n3096__), .dout(new_new_n3331__));
  or1   g1366(.dina(new_new_n3330__), .dinb(new_new_n4405__), .dout(new_new_n3332__));
  and1  g1367(.dina(new_new_n3332__), .dinb(new_new_n3331__), .dout(new_new_n3333__));
  and1  g1368(.dina(new_new_n4514__), .dinb(new_new_n4515__), .dout(new_new_n3334__));
  or1   g1369(.dina(new_new_n4516__), .dinb(new_new_n4517__), .dout(new_new_n3335__));
  and1  g1370(.dina(new_new_n4516__), .dinb(new_new_n4517__), .dout(new_new_n3336__));
  or1   g1371(.dina(new_new_n4514__), .dinb(new_new_n4515__), .dout(new_new_n3337__));
  and1  g1372(.dina(new_new_n3337__), .dinb(new_new_n3335__), .dout(new_new_n3338__));
  or1   g1373(.dina(new_new_n3336__), .dinb(new_new_n3334__), .dout(new_new_n3339__));
  and1  g1374(.dina(new_new_n4518__), .dinb(new_new_n4519__), .dout(new_new_n3340__));
  or1   g1375(.dina(new_new_n4520__), .dinb(new_new_n4521__), .dout(new_new_n3341__));
  and1  g1376(.dina(new_new_n4520__), .dinb(new_new_n4521__), .dout(new_new_n3342__));
  or1   g1377(.dina(new_new_n4518__), .dinb(new_new_n4519__), .dout(new_new_n3343__));
  and1  g1378(.dina(new_new_n3343__), .dinb(new_new_n3341__), .dout(new_new_n3344__));
  or1   g1379(.dina(new_new_n3342__), .dinb(new_new_n3340__), .dout(new_new_n3345__));
  and1  g1380(.dina(new_new_n4522__), .dinb(new_new_n4523__), .dout(new_new_n3346__));
  or1   g1381(.dina(new_new_n4524__), .dinb(new_new_n4525__), .dout(new_new_n3347__));
  and1  g1382(.dina(new_new_n4524__), .dinb(new_new_n4525__), .dout(new_new_n3348__));
  or1   g1383(.dina(new_new_n4522__), .dinb(new_new_n4523__), .dout(new_new_n3349__));
  and1  g1384(.dina(new_new_n3349__), .dinb(new_new_n3347__), .dout(new_new_n3350__));
  or1   g1385(.dina(new_new_n3348__), .dinb(new_new_n3346__), .dout(new_new_n3351__));
  and1  g1386(.dina(new_new_n4526__), .dinb(new_new_n4527__), .dout(new_new_n3352__));
  or1   g1387(.dina(new_new_n4528__), .dinb(new_new_n4529__), .dout(new_new_n3353__));
  and1  g1388(.dina(new_new_n4528__), .dinb(new_new_n4529__), .dout(new_new_n3354__));
  or1   g1389(.dina(new_new_n4526__), .dinb(new_new_n4527__), .dout(new_new_n3355__));
  and1  g1390(.dina(new_new_n3355__), .dinb(new_new_n3353__), .dout(new_new_n3356__));
  or1   g1391(.dina(new_new_n3354__), .dinb(new_new_n3352__), .dout(new_new_n3357__));
  or1   g1392(.dina(new_new_n3357__), .dinb(new_new_n3350__), .dout(new_new_n3358__));
  or1   g1393(.dina(new_new_n3356__), .dinb(new_new_n3351__), .dout(new_new_n3359__));
  and1  g1394(.dina(new_new_n3359__), .dinb(new_new_n3358__), .dout(new_new_n3360__));
  and1  g1395(.dina(new_new_n4314__), .dinb(new_new_n3037__), .dout(new_new_n3361__));
  and1  g1396(.dina(new_new_n4452__), .dinb(new_new_n4278__), .dout(new_new_n3362__));
  or1   g1397(.dina(new_new_n3362__), .dinb(new_new_n3361__), .dout(new_new_n3363__));
  or1   g1398(.dina(new_new_n4290__), .dinb(new_new_n4439__), .dout(new_new_n3364__));
  or1   g1399(.dina(new_new_n4312__), .dinb(new_new_n4451__), .dout(new_new_n3365__));
  and1  g1400(.dina(new_new_n3365__), .dinb(new_new_n3364__), .dout(new_new_n3366__));
  and1  g1401(.dina(new_new_n4530__), .dinb(new_new_n4531__), .dout(new_new_n3367__));
  or1   g1402(.dina(new_new_n4530__), .dinb(new_new_n4531__), .dout(new_new_n3368__));
  and1  g1403(.dina(new_new_n4532__), .dinb(new_new_n4459__), .dout(new_new_n3369__));
  or1   g1404(.dina(new_new_n4533__), .dinb(new_new_n4473__), .dout(new_new_n3370__));
  and1  g1405(.dina(new_new_n4533__), .dinb(new_new_n4472__), .dout(new_new_n3371__));
  or1   g1406(.dina(new_new_n4532__), .dinb(new_new_n4458__), .dout(new_new_n3372__));
  and1  g1407(.dina(new_new_n3372__), .dinb(new_new_n3370__), .dout(new_new_n3373__));
  or1   g1408(.dina(new_new_n3371__), .dinb(new_new_n3369__), .dout(new_new_n3374__));
  and1  g1409(.dina(new_new_n4333__), .dinb(new_new_n4534__), .dout(new_new_n3375__));
  or1   g1410(.dina(new_new_n4535__), .dinb(new_new_n4323__), .dout(new_new_n3376__));
  and1  g1411(.dina(new_new_n4535__), .dinb(new_new_n4324__), .dout(new_new_n3377__));
  or1   g1412(.dina(new_new_n4332__), .dinb(new_new_n4534__), .dout(new_new_n3378__));
  and1  g1413(.dina(new_new_n3378__), .dinb(new_new_n3376__), .dout(new_new_n3379__));
  or1   g1414(.dina(new_new_n3377__), .dinb(new_new_n3375__), .dout(new_new_n3380__));
  and1  g1415(.dina(new_new_n4536__), .dinb(new_new_n4537__), .dout(new_new_n3381__));
  or1   g1416(.dina(new_new_n4538__), .dinb(new_new_n4539__), .dout(new_new_n3382__));
  and1  g1417(.dina(new_new_n4538__), .dinb(new_new_n4539__), .dout(new_new_n3383__));
  or1   g1418(.dina(new_new_n4536__), .dinb(new_new_n4537__), .dout(new_new_n3384__));
  and1  g1419(.dina(new_new_n3384__), .dinb(new_new_n3382__), .dout(new_new_n3385__));
  or1   g1420(.dina(new_new_n3383__), .dinb(new_new_n3381__), .dout(new_new_n3386__));
  and1  g1421(.dina(new_new_n4540__), .dinb(new_new_n4349__), .dout(new_new_n3387__));
  or1   g1422(.dina(new_new_n4462__), .dinb(new_new_n4351__), .dout(new_new_n3388__));
  and1  g1423(.dina(new_new_n4462__), .dinb(new_new_n4350__), .dout(new_new_n3389__));
  or1   g1424(.dina(new_new_n4540__), .dinb(new_new_n4349__), .dout(new_new_n3390__));
  and1  g1425(.dina(new_new_n3390__), .dinb(new_new_n3388__), .dout(new_new_n3391__));
  or1   g1426(.dina(new_new_n3389__), .dinb(new_new_n3387__), .dout(new_new_n3392__));
  and1  g1427(.dina(new_new_n3391__), .dinb(new_new_n3386__), .dout(new_new_n3393__));
  and1  g1428(.dina(new_new_n3392__), .dinb(new_new_n3385__), .dout(new_new_n3394__));
  or1   g1429(.dina(new_new_n3394__), .dinb(new_new_n3393__), .dout(new_new_n3395__));
  or1   g1430(.dina(new_new_n4384__), .dinb(new_new_n1995__), .dout(new_new_n3396__));
  and1  g1431(.dina(new_new_n3396__), .dinb(new_new_n4378__), .dout(new_new_n3397__));
  and1  g1432(.dina(new_new_n2791__), .dinb(new_new_n4394__), .dout(new_new_n3398__));
  and1  g1433(.dina(new_new_n3398__), .dinb(new_new_n4367__), .dout(new_new_n3399__));
  and1  g1434(.dina(new_new_n4385__), .dinb(new_new_n2039__), .dout(new_new_n3400__));
  or1   g1435(.dina(new_new_n3400__), .dinb(new_new_n3399__), .dout(new_new_n3401__));
  or1   g1436(.dina(new_new_n3401__), .dinb(new_new_n3397__), .dout(new_new_n3402__));
  and1  g1437(.dina(new_new_n4394__), .dinb(new_new_n1890__), .dout(new_new_n3403__));
  and1  g1438(.dina(new_new_n4396__), .dinb(new_new_n1894__), .dout(new_new_n3404__));
  and1  g1439(.dina(new_new_n4396__), .dinb(new_new_n1974__), .dout(new_new_n3405__));
  and1  g1440(.dina(new_new_n4397__), .dinb(new_new_n1978__), .dout(new_new_n3406__));
  and1  g1441(.dina(new_new_n4397__), .dinb(new_new_n1986__), .dout(new_new_n3407__));
  and1  g1442(.dina(new_new_n4385__), .dinb(new_new_n2018__), .dout(new_new_n3408__));
  and1  g1443(.dina(new_new_n4386__), .dinb(new_new_n2022__), .dout(new_new_n3409__));
  and1  g1444(.dina(new_new_n4386__), .dinb(new_new_n2031__), .dout(new_new_n3410__));
  and1  g1445(.dina(new_new_n4367__), .dinb(new_new_n1899__), .dout(new_new_n3411__));
  or1   g1446(.dina(new_new_n4369__), .dinb(new_new_n1982__), .dout(new_new_n3412__));
  and1  g1447(.dina(new_new_n4400__), .dinb(new_new_n1903__), .dout(new_new_n3413__));
  and1  g1448(.dina(new_new_n3413__), .dinb(new_new_n4369__), .dout(new_new_n3414__));
  and1  g1449(.dina(new_new_n4400__), .dinb(new_new_n1990__), .dout(new_new_n3415__));
  or1   g1450(.dina(new_new_n3415__), .dinb(new_new_n4368__), .dout(new_new_n3416__));
  and1  g1451(.dina(new_new_n4388__), .dinb(new_new_n2048__), .dout(new_new_n3417__));
  and1  g1452(.dina(new_new_n4401__), .dinb(new_new_n1918__), .dout(new_new_n3418__));
  or1   g1453(.dina(new_new_n3418__), .dinb(new_new_n3417__), .dout(new_new_n3419__));
  and1  g1454(.dina(new_new_n3419__), .dinb(new_new_n4371__), .dout(new_new_n3420__));
  or1   g1455(.dina(new_new_n4542__), .dinb(new_new_n4544__), .dout(new_new_n3421__));
  or1   g1456(.dina(new_new_n4547__), .dinb(new_new_n4549__), .dout(new_new_n3422__));
  and1  g1457(.dina(new_new_n3422__), .dinb(new_new_n3421__), .dout(new_new_n3423__));
  and1  g1458(.dina(new_new_n4550__), .dinb(new_new_n4552__), .dout(new_new_n3424__));
  and1  g1459(.dina(new_new_n4556__), .dinb(new_new_n2076__), .dout(new_new_n3425__));
  and1  g1460(.dina(new_new_n4567__), .dinb(new_new_n2184__), .dout(new_new_n3426__));
  or1   g1461(.dina(new_new_n3426__), .dinb(new_new_n3425__), .dout(new_new_n3427__));
  and1  g1462(.dina(new_new_n4556__), .dinb(new_new_n2084__), .dout(new_new_n3428__));
  and1  g1463(.dina(new_new_n4567__), .dinb(new_new_n2192__), .dout(new_new_n3429__));
  or1   g1464(.dina(new_new_n3429__), .dinb(new_new_n3428__), .dout(new_new_n3430__));
  and1  g1465(.dina(new_new_n4557__), .dinb(new_new_n2088__), .dout(new_new_n3431__));
  and1  g1466(.dina(new_new_n4568__), .dinb(new_new_n2196__), .dout(new_new_n3432__));
  or1   g1467(.dina(new_new_n3432__), .dinb(new_new_n3431__), .dout(new_new_n3433__));
  and1  g1468(.dina(new_new_n4557__), .dinb(new_new_n2112__), .dout(new_new_n3434__));
  and1  g1469(.dina(new_new_n4568__), .dinb(new_new_n2148__), .dout(new_new_n3435__));
  or1   g1470(.dina(new_new_n3435__), .dinb(new_new_n3434__), .dout(new_new_n3436__));
  and1  g1471(.dina(new_new_n4559__), .dinb(new_new_n2120__), .dout(new_new_n3437__));
  and1  g1472(.dina(new_new_n4570__), .dinb(new_new_n2156__), .dout(new_new_n3438__));
  or1   g1473(.dina(new_new_n3438__), .dinb(new_new_n3437__), .dout(new_new_n3439__));
  and1  g1474(.dina(new_new_n4559__), .dinb(new_new_n2124__), .dout(new_new_n3440__));
  and1  g1475(.dina(new_new_n4570__), .dinb(new_new_n2160__), .dout(new_new_n3441__));
  or1   g1476(.dina(new_new_n3441__), .dinb(new_new_n3440__), .dout(new_new_n3442__));
  and1  g1477(.dina(new_new_n4560__), .dinb(new_new_n2080__), .dout(new_new_n3443__));
  and1  g1478(.dina(new_new_n4571__), .dinb(new_new_n2188__), .dout(new_new_n3444__));
  or1   g1479(.dina(new_new_n3444__), .dinb(new_new_n3443__), .dout(new_new_n3445__));
  and1  g1480(.dina(new_new_n3445__), .dinb(new_new_n4577__), .dout(new_new_n3446__));
  and1  g1481(.dina(new_new_n4560__), .dinb(new_new_n2116__), .dout(new_new_n3447__));
  and1  g1482(.dina(new_new_n4571__), .dinb(new_new_n2152__), .dout(new_new_n3448__));
  or1   g1483(.dina(new_new_n3448__), .dinb(new_new_n3447__), .dout(new_new_n3449__));
  and1  g1484(.dina(new_new_n3449__), .dinb(new_new_n4580__), .dout(new_new_n3450__));
  or1   g1485(.dina(new_new_n3450__), .dinb(new_new_n3446__), .dout(new_new_n3451__));
  and1  g1486(.dina(new_new_n4562__), .dinb(new_new_n2060__), .dout(new_new_n3452__));
  and1  g1487(.dina(new_new_n4574__), .dinb(new_new_n2168__), .dout(new_new_n3453__));
  or1   g1488(.dina(new_new_n3453__), .dinb(new_new_n3452__), .dout(new_new_n3454__));
  and1  g1489(.dina(new_new_n3454__), .dinb(new_new_n4577__), .dout(new_new_n3455__));
  and1  g1490(.dina(new_new_n4562__), .dinb(new_new_n2096__), .dout(new_new_n3456__));
  and1  g1491(.dina(new_new_n4574__), .dinb(new_new_n2132__), .dout(new_new_n3457__));
  or1   g1492(.dina(new_new_n3457__), .dinb(new_new_n3456__), .dout(new_new_n3458__));
  and1  g1493(.dina(new_new_n3458__), .dinb(new_new_n4580__), .dout(new_new_n3459__));
  or1   g1494(.dina(new_new_n3459__), .dinb(new_new_n3455__), .dout(new_new_n3460__));
  and1  g1495(.dina(new_new_n4563__), .dinb(new_new_n2092__), .dout(new_new_n3461__));
  and1  g1496(.dina(new_new_n4573__), .dinb(new_new_n2200__), .dout(new_new_n3462__));
  or1   g1497(.dina(new_new_n3462__), .dinb(new_new_n3461__), .dout(new_new_n3463__));
  and1  g1498(.dina(new_new_n3463__), .dinb(new_new_n4578__), .dout(new_new_n3464__));
  and1  g1499(.dina(new_new_n4563__), .dinb(new_new_n2128__), .dout(new_new_n3465__));
  and1  g1500(.dina(new_new_n4575__), .dinb(new_new_n2164__), .dout(new_new_n3466__));
  or1   g1501(.dina(new_new_n3466__), .dinb(new_new_n3465__), .dout(new_new_n3467__));
  and1  g1502(.dina(new_new_n3467__), .dinb(new_new_n4579__), .dout(new_new_n3468__));
  or1   g1503(.dina(new_new_n3468__), .dinb(new_new_n3464__), .dout(new_new_n3469__));
  and1  g1504(.dina(new_new_n4401__), .dinb(new_new_n1907__), .dout(new_new_n3470__));
  and1  g1505(.dina(new_new_n3470__), .dinb(new_new_n4371__), .dout(new_new_n3471__));
  and1  g1506(.dina(new_new_n4388__), .dinb(new_new_n2035__), .dout(new_new_n3472__));
  or1   g1507(.dina(new_new_n3472__), .dinb(new_new_n3471__), .dout(new_new_n3473__));
  and1  g1508(.dina(new_new_n4389__), .dinb(new_new_n2042__), .dout(new_new_n3474__));
  and1  g1509(.dina(new_new_n4403__), .dinb(new_new_n1912__), .dout(new_new_n3475__));
  or1   g1510(.dina(new_new_n3475__), .dinb(new_new_n3474__), .dout(new_new_n3476__));
  and1  g1511(.dina(new_new_n3476__), .dinb(new_new_n4372__), .dout(new_new_n3477__));
  and1  g1512(.dina(new_new_n4374__), .dinb(new_new_n1954__), .dout(new_new_n3478__));
  and1  g1513(.dina(new_new_n4403__), .dinb(new_new_n1998__), .dout(new_new_n3479__));
  and1  g1514(.dina(new_new_n3479__), .dinb(new_new_n4380__), .dout(new_new_n3480__));
  or1   g1515(.dina(new_new_n3480__), .dinb(new_new_n3478__), .dout(new_new_n3481__));
  or1   g1516(.dina(new_new_n3481__), .dinb(new_new_n3477__), .dout(new_new_n3482__));
  and1  g1517(.dina(new_new_n4376__), .dinb(new_new_n1960__), .dout(new_new_n3483__));
  and1  g1518(.dina(new_new_n4402__), .dinb(new_new_n2004__), .dout(new_new_n3484__));
  and1  g1519(.dina(new_new_n3484__), .dinb(new_new_n4380__), .dout(new_new_n3485__));
  or1   g1520(.dina(new_new_n3485__), .dinb(new_new_n3483__), .dout(new_new_n3486__));
  and1  g1521(.dina(new_new_n4581__), .dinb(new_new_n4582__), .dout(new_new_n3487__));
  or1   g1522(.dina(new_new_n4542__), .dinb(new_new_n4583__), .dout(new_new_n3488__));
  or1   g1523(.dina(new_new_n4547__), .dinb(new_new_n4584__), .dout(new_new_n3489__));
  and1  g1524(.dina(new_new_n3489__), .dinb(new_new_n3488__), .dout(new_new_n3490__));
  or1   g1525(.dina(new_new_n4543__), .dinb(new_new_n4585__), .dout(new_new_n3491__));
  or1   g1526(.dina(new_new_n4546__), .dinb(new_new_n4586__), .dout(new_new_n3492__));
  and1  g1527(.dina(new_new_n3492__), .dinb(new_new_n3491__), .dout(new_new_n3493__));
  or1   g1528(.dina(new_new_n4550__), .dinb(new_new_n4552__), .dout(new_new_n3494__));
  and1  g1529(.dina(new_new_n4548__), .dinb(new_new_n4587__), .dout(new_new_n3495__));
  and1  g1530(.dina(new_new_n4543__), .dinb(new_new_n4588__), .dout(new_new_n3496__));
  or1   g1531(.dina(new_new_n3496__), .dinb(new_new_n4589__), .dout(new_new_n3497__));
  or1   g1532(.dina(new_new_n3497__), .dinb(new_new_n3495__), .dout(new_new_n3498__));
  and1  g1533(.dina(new_new_n3498__), .dinb(new_new_n3494__), .dout(new_new_n3499__));
  or1   g1534(.dina(new_new_n4592__), .dinb(new_new_n2819__), .dout(new_new_n3500__));
  or1   g1535(.dina(new_new_n4595__), .dinb(new_new_n2831__), .dout(new_new_n3501__));
  and1  g1536(.dina(new_new_n3501__), .dinb(new_new_n3500__), .dout(new_new_n3502__));
  or1   g1537(.dina(new_new_n3502__), .dinb(new_new_n4597__), .dout(new_new_n3503__));
  or1   g1538(.dina(new_new_n4592__), .dinb(new_new_n2823__), .dout(new_new_n3504__));
  or1   g1539(.dina(new_new_n4595__), .dinb(new_new_n2827__), .dout(new_new_n3505__));
  and1  g1540(.dina(new_new_n3505__), .dinb(new_new_n3504__), .dout(new_new_n3506__));
  or1   g1541(.dina(new_new_n3506__), .dinb(new_new_n4599__), .dout(new_new_n3507__));
  and1  g1542(.dina(new_new_n4600__), .dinb(new_new_n1878__), .dout(new_new_n3508__));
  and1  g1543(.dina(new_new_n4600__), .dinb(new_new_n1962__), .dout(new_new_n3509__));
  and1  g1544(.dina(new_new_n4602__), .dinb(new_new_n2006__), .dout(new_new_n3510__));
  and1  g1545(.dina(new_new_n2237__), .dinb(new_new_n4602__), .dout(new_new_n3511__));
  and1  g1546(.dina(new_new_n4603__), .dinb(new_new_n4604__), .dout(new_new_n3512__));
  and1  g1547(.dina(new_new_n4596__), .dinb(new_new_n2820__), .dout(new_new_n3513__));
  and1  g1548(.dina(new_new_n4591__), .dinb(new_new_n2832__), .dout(new_new_n3514__));
  or1   g1549(.dina(new_new_n3514__), .dinb(new_new_n3513__), .dout(new_new_n3515__));
  and1  g1550(.dina(new_new_n3515__), .dinb(new_new_n4599__), .dout(new_new_n3516__));
  and1  g1551(.dina(new_new_n4596__), .dinb(new_new_n2824__), .dout(new_new_n3517__));
  and1  g1552(.dina(new_new_n4593__), .dinb(new_new_n2828__), .dout(new_new_n3518__));
  or1   g1553(.dina(new_new_n3518__), .dinb(new_new_n3517__), .dout(new_new_n3519__));
  and1  g1554(.dina(new_new_n3519__), .dinb(new_new_n4597__), .dout(new_new_n3520__));
  or1   g1555(.dina(new_new_n3520__), .dinb(new_new_n3516__), .dout(new_new_n3521__));
  buf1  g1556(.din(new_new_n4163__), .dout(G2531));
  buf1  g1557(.din(new_new_n4164__), .dout(G2532));
  buf1  g1558(.din(G2532), .dout(G2533));
  buf1  g1559(.din(new_new_n4605__), .dout(G2534));
  buf1  g1560(.din(G2534), .dout(G2535));
  buf1  g1561(.din(new_new_n4607__), .dout(G2536));
  buf1  g1562(.din(G2536), .dout(G2537));
  buf1  g1563(.din(new_new_n4606__), .dout(G2538));
  buf1  g1564(.din(new_new_n1887__), .dout(G2539));
  buf1  g1565(.din(new_new_n2177__), .dout(G2540));
  buf1  g1566(.din(new_new_n2015__), .dout(G2541));
  buf1  g1567(.din(new_new_n2069__), .dout(G2542));
  buf1  g1568(.din(new_new_n1971__), .dout(G2543));
  buf1  g1569(.din(new_new_n2141__), .dout(G2544));
  buf1  g1570(.din(new_new_n1929__), .dout(G2545));
  buf1  g1571(.din(new_new_n2105__), .dout(G2546));
  buf1  g1572(.din(new_new_n2836__), .dout(G2547));
  buf1  g1573(.din(new_new_n2838__), .dout(G2548));
  buf1  g1574(.din(new_new_n2208__), .dout(G2549));
  buf1  g1575(.din(new_new_n2839__), .dout(G2550));
  buf1  g1576(.din(new_new_n4165__), .dout(G2551));
  buf1  g1577(.din(new_new_n2841__), .dout(G2552));
  buf1  g1578(.din(new_new_n2842__), .dout(G2553));
  buf1  g1579(.din(new_new_n4608__), .dout(G2554));
  buf1  g1580(.din(G2554), .dout(G2555));
  buf1  g1581(.din(new_new_n4171__), .dout(G2556));
  buf1  g1582(.din(new_new_n2849__), .dout(G2557));
  buf1  g1583(.din(new_new_n2850__), .dout(G2558));
  buf1  g1584(.din(new_new_n2465__), .dout(G2559));
  buf1  g1585(.din(new_new_n2851__), .dout(G2560));
  not1  g1586(.din(new_new_n4182__), .dout(G2561));
  buf1  g1587(.din(new_new_n2501__), .dout(G2562));
  buf1  g1588(.din(new_new_n2853__), .dout(G2563));
  buf1  g1589(.din(new_new_n2856__), .dout(G2564));
  buf1  g1590(.din(new_new_n2858__), .dout(G2565));
  buf1  g1591(.din(new_new_n2472__), .dout(G2566));
  buf1  g1592(.din(new_new_n4178__), .dout(G2567));
  buf1  g1593(.din(new_new_n2490__), .dout(G2568));
  buf1  g1594(.din(new_new_n2502__), .dout(G2569));
  buf1  g1595(.din(new_new_n2504__), .dout(G2570));
  buf1  g1596(.din(new_new_n2506__), .dout(G2571));
  buf1  g1597(.din(new_new_n2508__), .dout(G2572));
  buf1  g1598(.din(new_new_n4609__), .dout(G2573));
  buf1  g1599(.din(G2573), .dout(G2574));
  not1  g1600(.din(new_new_n4610__), .dout(G2575));
  buf1  g1601(.din(G2575), .dout(G2576));
  buf1  g1602(.din(new_new_n2866__), .dout(G2577));
  buf1  g1603(.din(new_new_n4611__), .dout(G2578));
  buf1  g1604(.din(G2578), .dout(G2579));
  buf1  g1605(.din(new_new_n2873__), .dout(G2580));
  not1  g1606(.din(new_new_n4208__), .dout(G2581));
  buf1  g1607(.din(new_new_n4207__), .dout(G2582));
  buf1  g1608(.din(new_new_n4209__), .dout(G2583));
  buf1  g1609(.din(new_new_n4612__), .dout(G2584));
  buf1  g1610(.din(G2584), .dout(G2585));
  buf1  g1611(.din(new_new_n2957__), .dout(G2586));
  not1  g1612(.din(new_new_n4210__), .dout(G2587));
  buf1  g1613(.din(new_new_n4613__), .dout(G2588));
  buf1  g1614(.din(G2588), .dout(G2589));
  not1  g1615(.din(new_new_n4211__), .dout(G2590));
  buf1  g1616(.din(new_new_n3007__), .dout(G2591));
  buf1  g1617(.din(new_new_n4615__), .dout(G2592));
  buf1  g1618(.din(new_new_n4614__), .dout(G2593));
  buf1  g1619(.din(G2593), .dout(G2594));
  buf1  g1620(.din(new_new_n1372__), .dout(n6254));
  buf1  g1621(.din(new_new_n1686__), .dout(n6257));
  buf1  g1622(.din(new_new_n1688__), .dout(n6260));
  buf1  g1623(.din(new_new_n1690__), .dout(n6263));
  buf1  g1624(.din(new_new_n1374__), .dout(n6266));
  buf1  g1625(.din(new_new_n1694__), .dout(n6269));
  buf1  g1626(.din(new_new_n1696__), .dout(n6272));
  buf1  g1627(.din(new_new_n1698__), .dout(n6275));
  buf1  g1628(.din(new_new_n1376__), .dout(n6278));
  buf1  g1629(.din(new_new_n1702__), .dout(n6281));
  buf1  g1630(.din(new_new_n1704__), .dout(n6284));
  buf1  g1631(.din(new_new_n1706__), .dout(n6287));
  buf1  g1632(.din(new_new_n1378__), .dout(n6290));
  buf1  g1633(.din(new_new_n1710__), .dout(n6293));
  buf1  g1634(.din(new_new_n1712__), .dout(n6296));
  buf1  g1635(.din(new_new_n1380__), .dout(n6299));
  buf1  g1636(.din(new_new_n1716__), .dout(n6302));
  buf1  g1637(.din(new_new_n1718__), .dout(n6305));
  buf1  g1638(.din(new_new_n1382__), .dout(n6308));
  buf1  g1639(.din(new_new_n1722__), .dout(n6311));
  buf1  g1640(.din(new_new_n1724__), .dout(n6314));
  buf1  g1641(.din(new_new_n1384__), .dout(n6317));
  buf1  g1642(.din(new_new_n1728__), .dout(n6320));
  buf1  g1643(.din(new_new_n1730__), .dout(n6323));
  buf1  g1644(.din(new_new_n1732__), .dout(n6326));
  buf1  g1645(.din(new_new_n1386__), .dout(n6329));
  buf1  g1646(.din(new_new_n1736__), .dout(n6332));
  buf1  g1647(.din(new_new_n1388__), .dout(n6335));
  buf1  g1648(.din(new_new_n1740__), .dout(n6338));
  buf1  g1649(.din(new_new_n1742__), .dout(n6341));
  buf1  g1650(.din(new_new_n1744__), .dout(n6344));
  buf1  g1651(.din(new_new_n1390__), .dout(n6347));
  buf1  g1652(.din(new_new_n1748__), .dout(n6350));
  buf1  g1653(.din(new_new_n1750__), .dout(n6353));
  buf1  g1654(.din(new_new_n1752__), .dout(n6356));
  buf1  g1655(.din(new_new_n1392__), .dout(n6359));
  buf1  g1656(.din(new_new_n1756__), .dout(n6362));
  buf1  g1657(.din(new_new_n1758__), .dout(n6365));
  buf1  g1658(.din(new_new_n1760__), .dout(n6368));
  buf1  g1659(.din(new_new_n1394__), .dout(n6371));
  buf1  g1660(.din(new_new_n1764__), .dout(n6374));
  buf1  g1661(.din(new_new_n1766__), .dout(n6377));
  buf1  g1662(.din(new_new_n1396__), .dout(n6380));
  buf1  g1663(.din(new_new_n1770__), .dout(n6383));
  buf1  g1664(.din(new_new_n1772__), .dout(n6386));
  buf1  g1665(.din(new_new_n1398__), .dout(n6389));
  buf1  g1666(.din(new_new_n1776__), .dout(n6392));
  buf1  g1667(.din(new_new_n1778__), .dout(n6395));
  buf1  g1668(.din(new_new_n1400__), .dout(n6398));
  buf1  g1669(.din(new_new_n1782__), .dout(n6401));
  buf1  g1670(.din(new_new_n1784__), .dout(n6404));
  buf1  g1671(.din(new_new_n1402__), .dout(n6407));
  buf1  g1672(.din(new_new_n1788__), .dout(n6410));
  buf1  g1673(.din(new_new_n1790__), .dout(n6413));
  buf1  g1674(.din(new_new_n1404__), .dout(n6416));
  buf1  g1675(.din(new_new_n1794__), .dout(n6419));
  buf1  g1676(.din(new_new_n1796__), .dout(n6422));
  buf1  g1677(.din(new_new_n1406__), .dout(n6425));
  buf1  g1678(.din(new_new_n1800__), .dout(n6428));
  buf1  g1679(.din(new_new_n1802__), .dout(n6431));
  buf1  g1680(.din(new_new_n1408__), .dout(n6434));
  buf1  g1681(.din(new_new_n1806__), .dout(n6437));
  buf1  g1682(.din(new_new_n1808__), .dout(n6440));
  buf1  g1683(.din(new_new_n1410__), .dout(n6443));
  buf1  g1684(.din(new_new_n1812__), .dout(n6446));
  buf1  g1685(.din(new_new_n1814__), .dout(n6449));
  buf1  g1686(.din(new_new_n1412__), .dout(n6452));
  buf1  g1687(.din(new_new_n1818__), .dout(n6455));
  buf1  g1688(.din(new_new_n1820__), .dout(n6458));
  buf1  g1689(.din(new_new_n1414__), .dout(n6461));
  buf1  g1690(.din(new_new_n1824__), .dout(n6464));
  buf1  g1691(.din(new_new_n1826__), .dout(n6467));
  buf1  g1692(.din(new_new_n1416__), .dout(n6470));
  buf1  g1693(.din(new_new_n1830__), .dout(n6473));
  buf1  g1694(.din(new_new_n1832__), .dout(n6476));
  buf1  g1695(.din(new_new_n1418__), .dout(n6479));
  buf1  g1696(.din(new_new_n1836__), .dout(n6482));
  buf1  g1697(.din(new_new_n1838__), .dout(n6485));
  buf1  g1698(.din(new_new_n1420__), .dout(n6488));
  buf1  g1699(.din(new_new_n1842__), .dout(n6491));
  buf1  g1700(.din(new_new_n1844__), .dout(n6494));
  buf1  g1701(.din(new_new_n1422__), .dout(n6497));
  buf1  g1702(.din(new_new_n1848__), .dout(n6500));
  buf1  g1703(.din(new_new_n1850__), .dout(n6503));
  buf1  g1704(.din(new_new_n1424__), .dout(n6506));
  buf1  g1705(.din(new_new_n1854__), .dout(n6509));
  buf1  g1706(.din(new_new_n1856__), .dout(n6512));
  buf1  g1707(.din(new_new_n1426__), .dout(n6515));
  buf1  g1708(.din(new_new_n1860__), .dout(n6518));
  buf1  g1709(.din(new_new_n1862__), .dout(n6521));
  buf1  g1710(.din(new_new_n1864__), .dout(n6524));
  buf1  g1711(.din(new_new_n1428__), .dout(n6527));
  buf1  g1712(.din(new_new_n1868__), .dout(n6530));
  buf1  g1713(.din(new_new_n1870__), .dout(n6533));
  buf1  g1714(.din(new_new_n1872__), .dout(n6536));
  buf1  g1715(.din(new_new_n1430__), .dout(n6539));
  buf1  g1716(.din(new_new_n1432__), .dout(n6542));
  buf1  g1717(.din(new_new_n1434__), .dout(n6545));
  buf1  g1718(.din(new_new_n1880__), .dout(n6548));
  buf1  g1719(.din(new_new_n1882__), .dout(n6551));
  buf1  g1720(.din(new_new_n4407__), .dout(n6554));
  buf1  g1721(.din(new_new_n1436__), .dout(n6557));
  buf1  g1722(.din(new_new_n1888__), .dout(n6560));
  buf1  g1723(.din(new_new_n1438__), .dout(n6563));
  buf1  g1724(.din(new_new_n1892__), .dout(n6566));
  buf1  g1725(.din(new_new_n1440__), .dout(n6569));
  buf1  g1726(.din(new_new_n1896__), .dout(n6572));
  buf1  g1727(.din(new_new_n1442__), .dout(n6575));
  buf1  g1728(.din(new_new_n1900__), .dout(n6578));
  buf1  g1729(.din(new_new_n1444__), .dout(n6581));
  buf1  g1730(.din(new_new_n1904__), .dout(n6584));
  buf1  g1731(.din(new_new_n1446__), .dout(n6587));
  buf1  g1732(.din(new_new_n1448__), .dout(n6590));
  buf1  g1733(.din(new_new_n1910__), .dout(n6593));
  buf1  g1734(.din(new_new_n1450__), .dout(n6596));
  buf1  g1735(.din(new_new_n1452__), .dout(n6599));
  buf1  g1736(.din(new_new_n1916__), .dout(n6602));
  buf1  g1737(.din(new_new_n1454__), .dout(n6605));
  buf1  g1738(.din(new_new_n1456__), .dout(n6608));
  buf1  g1739(.din(new_new_n1922__), .dout(n6611));
  buf1  g1740(.din(new_new_n1924__), .dout(n6614));
  buf1  g1741(.din(new_new_n4409__), .dout(n6617));
  buf1  g1742(.din(new_new_n1458__), .dout(n6620));
  buf1  g1743(.din(new_new_n1930__), .dout(n6623));
  buf1  g1744(.din(new_new_n1460__), .dout(n6626));
  buf1  g1745(.din(new_new_n1934__), .dout(n6629));
  buf1  g1746(.din(new_new_n1462__), .dout(n6632));
  buf1  g1747(.din(new_new_n1938__), .dout(n6635));
  buf1  g1748(.din(new_new_n1940__), .dout(n6638));
  buf1  g1749(.din(new_new_n1464__), .dout(n6641));
  buf1  g1750(.din(new_new_n1944__), .dout(n6644));
  buf1  g1751(.din(new_new_n1466__), .dout(n6647));
  buf1  g1752(.din(new_new_n1948__), .dout(n6650));
  buf1  g1753(.din(new_new_n1468__), .dout(n6653));
  buf1  g1754(.din(new_new_n1952__), .dout(n6656));
  buf1  g1755(.din(new_new_n1470__), .dout(n6659));
  buf1  g1756(.din(new_new_n1472__), .dout(n6662));
  buf1  g1757(.din(new_new_n1958__), .dout(n6665));
  buf1  g1758(.din(new_new_n1474__), .dout(n6668));
  buf1  g1759(.din(new_new_n1476__), .dout(n6671));
  buf1  g1760(.din(new_new_n1964__), .dout(n6674));
  buf1  g1761(.din(new_new_n1966__), .dout(n6677));
  buf1  g1762(.din(new_new_n4408__), .dout(n6680));
  buf1  g1763(.din(new_new_n1478__), .dout(n6683));
  buf1  g1764(.din(new_new_n1972__), .dout(n6686));
  buf1  g1765(.din(new_new_n1480__), .dout(n6689));
  buf1  g1766(.din(new_new_n1976__), .dout(n6692));
  buf1  g1767(.din(new_new_n1482__), .dout(n6695));
  buf1  g1768(.din(new_new_n1980__), .dout(n6698));
  buf1  g1769(.din(new_new_n1484__), .dout(n6701));
  buf1  g1770(.din(new_new_n1984__), .dout(n6704));
  buf1  g1771(.din(new_new_n1486__), .dout(n6707));
  buf1  g1772(.din(new_new_n1988__), .dout(n6710));
  buf1  g1773(.din(new_new_n1488__), .dout(n6713));
  buf1  g1774(.din(new_new_n1992__), .dout(n6716));
  buf1  g1775(.din(new_new_n1490__), .dout(n6719));
  buf1  g1776(.din(new_new_n1996__), .dout(n6722));
  buf1  g1777(.din(new_new_n1492__), .dout(n6725));
  buf1  g1778(.din(new_new_n1494__), .dout(n6728));
  buf1  g1779(.din(new_new_n2002__), .dout(n6731));
  buf1  g1780(.din(new_new_n1496__), .dout(n6734));
  buf1  g1781(.din(new_new_n1498__), .dout(n6737));
  buf1  g1782(.din(new_new_n2008__), .dout(n6740));
  buf1  g1783(.din(new_new_n2010__), .dout(n6743));
  buf1  g1784(.din(new_new_n4406__), .dout(n6746));
  buf1  g1785(.din(new_new_n1500__), .dout(n6749));
  buf1  g1786(.din(new_new_n2016__), .dout(n6752));
  buf1  g1787(.din(new_new_n1502__), .dout(n6755));
  buf1  g1788(.din(new_new_n2020__), .dout(n6758));
  buf1  g1789(.din(new_new_n1504__), .dout(n6761));
  buf1  g1790(.din(new_new_n2024__), .dout(n6764));
  buf1  g1791(.din(new_new_n1506__), .dout(n6767));
  buf1  g1792(.din(new_new_n2028__), .dout(n6770));
  buf1  g1793(.din(new_new_n1508__), .dout(n6773));
  buf1  g1794(.din(new_new_n2032__), .dout(n6776));
  buf1  g1795(.din(new_new_n1510__), .dout(n6779));
  buf1  g1796(.din(new_new_n2036__), .dout(n6782));
  buf1  g1797(.din(new_new_n1512__), .dout(n6785));
  buf1  g1798(.din(new_new_n2040__), .dout(n6788));
  buf1  g1799(.din(new_new_n1514__), .dout(n6791));
  buf1  g1800(.din(new_new_n1516__), .dout(n6794));
  buf1  g1801(.din(new_new_n2046__), .dout(n6797));
  buf1  g1802(.din(new_new_n1518__), .dout(n6800));
  buf1  g1803(.din(new_new_n2050__), .dout(n6803));
  buf1  g1804(.din(new_new_n2052__), .dout(n6806));
  buf1  g1805(.din(new_new_n2054__), .dout(n6809));
  buf1  g1806(.din(new_new_n1520__), .dout(n6812));
  buf1  g1807(.din(new_new_n2058__), .dout(n6815));
  buf1  g1808(.din(new_new_n1522__), .dout(n6818));
  buf1  g1809(.din(new_new_n2062__), .dout(n6821));
  buf1  g1810(.din(new_new_n2064__), .dout(n6824));
  buf1  g1811(.din(new_new_n4411__), .dout(n6827));
  buf1  g1812(.din(new_new_n1524__), .dout(n6830));
  buf1  g1813(.din(new_new_n2070__), .dout(n6833));
  buf1  g1814(.din(new_new_n1526__), .dout(n6836));
  buf1  g1815(.din(new_new_n2074__), .dout(n6839));
  buf1  g1816(.din(new_new_n1532__), .dout(n6842));
  buf1  g1817(.din(new_new_n2078__), .dout(n6845));
  buf1  g1818(.din(new_new_n1534__), .dout(n6848));
  buf1  g1819(.din(new_new_n2082__), .dout(n6851));
  buf1  g1820(.din(new_new_n1536__), .dout(n6854));
  buf1  g1821(.din(new_new_n2086__), .dout(n6857));
  buf1  g1822(.din(new_new_n1538__), .dout(n6860));
  buf1  g1823(.din(new_new_n2090__), .dout(n6863));
  buf1  g1824(.din(new_new_n1540__), .dout(n6866));
  buf1  g1825(.din(new_new_n2094__), .dout(n6869));
  buf1  g1826(.din(new_new_n1542__), .dout(n6872));
  buf1  g1827(.din(new_new_n2098__), .dout(n6875));
  buf1  g1828(.din(new_new_n2100__), .dout(n6878));
  buf1  g1829(.din(new_new_n4413__), .dout(n6881));
  buf1  g1830(.din(new_new_n1544__), .dout(n6884));
  buf1  g1831(.din(new_new_n2106__), .dout(n6887));
  buf1  g1832(.din(new_new_n1546__), .dout(n6890));
  buf1  g1833(.din(new_new_n2110__), .dout(n6893));
  buf1  g1834(.din(new_new_n1552__), .dout(n6896));
  buf1  g1835(.din(new_new_n2114__), .dout(n6899));
  buf1  g1836(.din(new_new_n1554__), .dout(n6902));
  buf1  g1837(.din(new_new_n2118__), .dout(n6905));
  buf1  g1838(.din(new_new_n1556__), .dout(n6908));
  buf1  g1839(.din(new_new_n2122__), .dout(n6911));
  buf1  g1840(.din(new_new_n1558__), .dout(n6914));
  buf1  g1841(.din(new_new_n2126__), .dout(n6917));
  buf1  g1842(.din(new_new_n1560__), .dout(n6920));
  buf1  g1843(.din(new_new_n2130__), .dout(n6923));
  buf1  g1844(.din(new_new_n1562__), .dout(n6926));
  buf1  g1845(.din(new_new_n2134__), .dout(n6929));
  buf1  g1846(.din(new_new_n2136__), .dout(n6932));
  buf1  g1847(.din(new_new_n4412__), .dout(n6935));
  buf1  g1848(.din(new_new_n1564__), .dout(n6938));
  buf1  g1849(.din(new_new_n2142__), .dout(n6941));
  buf1  g1850(.din(new_new_n1566__), .dout(n6944));
  buf1  g1851(.din(new_new_n2146__), .dout(n6947));
  buf1  g1852(.din(new_new_n1572__), .dout(n6950));
  buf1  g1853(.din(new_new_n2150__), .dout(n6953));
  buf1  g1854(.din(new_new_n1574__), .dout(n6956));
  buf1  g1855(.din(new_new_n2154__), .dout(n6959));
  buf1  g1856(.din(new_new_n1576__), .dout(n6962));
  buf1  g1857(.din(new_new_n2158__), .dout(n6965));
  buf1  g1858(.din(new_new_n1578__), .dout(n6968));
  buf1  g1859(.din(new_new_n2162__), .dout(n6971));
  buf1  g1860(.din(new_new_n1580__), .dout(n6974));
  buf1  g1861(.din(new_new_n2166__), .dout(n6977));
  buf1  g1862(.din(new_new_n1582__), .dout(n6980));
  buf1  g1863(.din(new_new_n2170__), .dout(n6983));
  buf1  g1864(.din(new_new_n2172__), .dout(n6986));
  buf1  g1865(.din(new_new_n4410__), .dout(n6989));
  buf1  g1866(.din(new_new_n1584__), .dout(n6992));
  buf1  g1867(.din(new_new_n2178__), .dout(n6995));
  buf1  g1868(.din(new_new_n1586__), .dout(n6998));
  buf1  g1869(.din(new_new_n2182__), .dout(n7001));
  buf1  g1870(.din(new_new_n1592__), .dout(n7004));
  buf1  g1871(.din(new_new_n2186__), .dout(n7007));
  buf1  g1872(.din(new_new_n1594__), .dout(n7010));
  buf1  g1873(.din(new_new_n2190__), .dout(n7013));
  buf1  g1874(.din(new_new_n1596__), .dout(n7016));
  buf1  g1875(.din(new_new_n2194__), .dout(n7019));
  buf1  g1876(.din(new_new_n1598__), .dout(n7022));
  buf1  g1877(.din(new_new_n2198__), .dout(n7025));
  buf1  g1878(.din(new_new_n1600__), .dout(n7028));
  buf1  g1879(.din(new_new_n2202__), .dout(n7031));
  buf1  g1880(.din(new_new_n2204__), .dout(n7034));
  buf1  g1881(.din(new_new_n2206__), .dout(n7037));
  buf1  g1882(.din(new_new_n1602__), .dout(n7040));
  buf1  g1883(.din(new_new_n2210__), .dout(n7043));
  buf1  g1884(.din(new_new_n2212__), .dout(n7046));
  buf1  g1885(.din(new_new_n2214__), .dout(n7049));
  buf1  g1886(.din(new_new_n1604__), .dout(n7052));
  buf1  g1887(.din(new_new_n1606__), .dout(n7055));
  buf1  g1888(.din(new_new_n2220__), .dout(n7058));
  buf1  g1889(.din(new_new_n2222__), .dout(n7061));
  buf1  g1890(.din(new_new_n4414__), .dout(n7064));
  buf1  g1891(.din(new_new_n1608__), .dout(n7067));
  buf1  g1892(.din(new_new_n2228__), .dout(n7070));
  buf1  g1893(.din(new_new_n2230__), .dout(n7073));
  buf1  g1894(.din(new_new_n2232__), .dout(n7076));
  buf1  g1895(.din(new_new_n1610__), .dout(n7079));
  buf1  g1896(.din(new_new_n1612__), .dout(n7082));
  buf1  g1897(.din(new_new_n2238__), .dout(n7085));
  buf1  g1898(.din(new_new_n2240__), .dout(n7088));
  buf1  g1899(.din(new_new_n2242__), .dout(n7091));
  buf1  g1900(.din(new_new_n1614__), .dout(n7094));
  buf1  g1901(.din(new_new_n2246__), .dout(n7097));
  buf1  g1902(.din(new_new_n2248__), .dout(n7100));
  buf1  g1903(.din(new_new_n2250__), .dout(n7103));
  buf1  g1904(.din(new_new_n1616__), .dout(n7106));
  buf1  g1905(.din(new_new_n2254__), .dout(n7109));
  buf1  g1906(.din(new_new_n2256__), .dout(n7112));
  buf1  g1907(.din(new_new_n2258__), .dout(n7115));
  buf1  g1908(.din(new_new_n1618__), .dout(n7118));
  buf1  g1909(.din(new_new_n2262__), .dout(n7121));
  buf1  g1910(.din(new_new_n2264__), .dout(n7124));
  buf1  g1911(.din(new_new_n2266__), .dout(n7127));
  buf1  g1912(.din(new_new_n1620__), .dout(n7130));
  buf1  g1913(.din(new_new_n2270__), .dout(n7133));
  buf1  g1914(.din(new_new_n1622__), .dout(n7136));
  buf1  g1915(.din(new_new_n2274__), .dout(n7139));
  buf1  g1916(.din(new_new_n4504__), .dout(n7142));
  buf1  g1917(.din(new_new_n1624__), .dout(n7145));
  buf1  g1918(.din(new_new_n1626__), .dout(n7148));
  buf1  g1919(.din(new_new_n2282__), .dout(n7151));
  buf1  g1920(.din(new_new_n1628__), .dout(n7154));
  buf1  g1921(.din(new_new_n2286__), .dout(n7157));
  buf1  g1922(.din(new_new_n4467__), .dout(n7160));
  buf1  g1923(.din(new_new_n1630__), .dout(n7163));
  buf1  g1924(.din(new_new_n2292__), .dout(n7166));
  buf1  g1925(.din(new_new_n2294__), .dout(n7169));
  buf1  g1926(.din(new_new_n1632__), .dout(n7172));
  buf1  g1927(.din(new_new_n2298__), .dout(n7175));
  buf1  g1928(.din(new_new_n2300__), .dout(n7178));
  buf1  g1929(.din(new_new_n1634__), .dout(n7181));
  buf1  g1930(.din(new_new_n2304__), .dout(n7184));
  buf1  g1931(.din(new_new_n2306__), .dout(n7187));
  buf1  g1932(.din(new_new_n4507__), .dout(n7190));
  buf1  g1933(.din(new_new_n1636__), .dout(n7193));
  buf1  g1934(.din(new_new_n2312__), .dout(n7196));
  buf1  g1935(.din(new_new_n2314__), .dout(n7199));
  buf1  g1936(.din(new_new_n1638__), .dout(n7202));
  buf1  g1937(.din(new_new_n2318__), .dout(n7205));
  buf1  g1938(.din(new_new_n2320__), .dout(n7208));
  buf1  g1939(.din(new_new_n4284__), .dout(n7211));
  buf1  g1940(.din(new_new_n1640__), .dout(n7214));
  buf1  g1941(.din(new_new_n2326__), .dout(n7217));
  buf1  g1942(.din(new_new_n2328__), .dout(n7220));
  buf1  g1943(.din(new_new_n4470__), .dout(n7223));
  buf1  g1944(.din(new_new_n1642__), .dout(n7226));
  buf1  g1945(.din(new_new_n2334__), .dout(n7229));
  buf1  g1946(.din(new_new_n4353__), .dout(n7232));
  buf1  g1947(.din(new_new_n1644__), .dout(n7235));
  buf1  g1948(.din(new_new_n2340__), .dout(n7238));
  buf1  g1949(.din(new_new_n2342__), .dout(n7241));
  buf1  g1950(.din(new_new_n2344__), .dout(n7244));
  buf1  g1951(.din(new_new_n1646__), .dout(n7247));
  buf1  g1952(.din(new_new_n2348__), .dout(n7250));
  buf1  g1953(.din(new_new_n4490__), .dout(n7253));
  buf1  g1954(.din(new_new_n1648__), .dout(n7256));
  buf1  g1955(.din(new_new_n2354__), .dout(n7259));
  buf1  g1956(.din(new_new_n4234__), .dout(n7262));
  buf1  g1957(.din(new_new_n1650__), .dout(n7265));
  buf1  g1958(.din(new_new_n2360__), .dout(n7268));
  buf1  g1959(.din(new_new_n4232__), .dout(n7271));
  buf1  g1960(.din(new_new_n1652__), .dout(n7274));
  buf1  g1961(.din(new_new_n2366__), .dout(n7277));
  buf1  g1962(.din(new_new_n2368__), .dout(n7280));
  buf1  g1963(.din(new_new_n4486__), .dout(n7283));
  buf1  g1964(.din(new_new_n1654__), .dout(n7286));
  buf1  g1965(.din(new_new_n2374__), .dout(n7289));
  buf1  g1966(.din(new_new_n2376__), .dout(n7292));
  buf1  g1967(.din(new_new_n4485__), .dout(n7295));
  buf1  g1968(.din(new_new_n1656__), .dout(n7298));
  buf1  g1969(.din(new_new_n2382__), .dout(n7301));
  buf1  g1970(.din(new_new_n2384__), .dout(n7304));
  buf1  g1971(.din(new_new_n4449__), .dout(n7307));
  buf1  g1972(.din(new_new_n1658__), .dout(n7310));
  buf1  g1973(.din(new_new_n2390__), .dout(n7313));
  buf1  g1974(.din(new_new_n2392__), .dout(n7316));
  buf1  g1975(.din(new_new_n4450__), .dout(n7319));
  buf1  g1976(.din(new_new_n1662__), .dout(n7322));
  buf1  g1977(.din(new_new_n1664__), .dout(n7325));
  buf1  g1978(.din(new_new_n2400__), .dout(n7328));
  buf1  g1979(.din(new_new_n2402__), .dout(n7331));
  buf1  g1980(.din(new_new_n2404__), .dout(n7334));
  buf1  g1981(.din(new_new_n1666__), .dout(n7337));
  buf1  g1982(.din(new_new_n2408__), .dout(n7340));
  buf1  g1983(.din(new_new_n1668__), .dout(n7343));
  buf1  g1984(.din(new_new_n2412__), .dout(n7346));
  buf1  g1985(.din(new_new_n1670__), .dout(n7349));
  buf1  g1986(.din(new_new_n2416__), .dout(n7352));
  buf1  g1987(.din(new_new_n2418__), .dout(n7355));
  buf1  g1988(.din(new_new_n1672__), .dout(n7358));
  buf1  g1989(.din(new_new_n2422__), .dout(n7361));
  buf1  g1990(.din(new_new_n2424__), .dout(n7364));
  buf1  g1991(.din(new_new_n1674__), .dout(n7367));
  buf1  g1992(.din(new_new_n2428__), .dout(n7370));
  buf1  g1993(.din(new_new_n1676__), .dout(n7373));
  buf1  g1994(.din(new_new_n2432__), .dout(n7376));
  buf1  g1995(.din(new_new_n1678__), .dout(n7379));
  buf1  g1996(.din(new_new_n2436__), .dout(n7382));
  buf1  g1997(.din(new_new_n2438__), .dout(n7385));
  buf1  g1998(.din(new_new_n1680__), .dout(n7388));
  buf1  g1999(.din(new_new_n2442__), .dout(n7391));
  buf1  g2000(.din(new_new_n2444__), .dout(n7394));
  buf1  g2001(.din(new_new_n1682__), .dout(n7397));
  buf1  g2002(.din(new_new_n2448__), .dout(n7400));
  buf1  g2003(.din(new_new_n2450__), .dout(n7403));
  buf1  g2004(.din(new_new_n1684__), .dout(n7406));
  buf1  g2005(.din(new_new_n2454__), .dout(n7409));
  buf1  g2006(.din(new_new_n2456__), .dout(n7412));
  buf1  g2007(.din(new_new_n2512__), .dout(n7415));
  buf1  g2008(.din(new_new_n2514__), .dout(n7418));
  buf1  g2009(.din(new_new_n4324__), .dout(n7421));
  buf1  g2010(.din(new_new_n4262__), .dout(n7424));
  buf1  g2011(.din(new_new_n4302__), .dout(n7427));
  buf1  g2012(.din(new_new_n4455__), .dout(n7430));
  buf1  g2013(.din(new_new_n4359__), .dout(n7433));
  buf1  g2014(.din(new_new_n4241__), .dout(n7436));
  buf1  g2015(.din(new_new_n4464__), .dout(n7439));
  buf1  g2016(.din(new_new_n4463__), .dout(n7442));
  buf1  g2017(.din(new_new_n4240__), .dout(n7445));
  buf1  g2018(.din(new_new_n4256__), .dout(n7448));
  buf1  g2019(.din(new_new_n4575__), .dout(n7451));
  buf1  g2020(.din(new_new_n4253__), .dout(n7454));
  buf1  g2021(.din(new_new_n4488__), .dout(n7457));
  buf1  g2022(.din(new_new_n4428__), .dout(n7460));
  buf1  g2023(.din(new_new_n4252__), .dout(n7463));
  buf1  g2024(.din(new_new_n4578__), .dout(n7466));
  buf1  g2025(.din(new_new_n4389__), .dout(n7469));
  buf1  g2026(.din(new_new_n4372__), .dout(n7472));
  buf1  g2027(.din(new_new_n4495__), .dout(n7475));
  buf1  g2028(.din(new_new_n4278__), .dout(n7478));
  buf1  g2029(.din(new_new_n4313__), .dout(n7481));
  buf1  g2030(.din(new_new_n4438__), .dout(n7484));
  buf1  g2031(.din(new_new_n4311__), .dout(n7487));
  buf1  g2032(.din(new_new_n4362__), .dout(n7490));
  buf1  g2033(.din(new_new_n2786__), .dout(n7493));
  buf1  g2034(.din(new_new_n2788__), .dout(n7496));
  buf1  g2035(.din(new_new_n4376__), .dout(n7499));
  buf1  g2036(.din(new_new_n4272__), .dout(n7502));
  buf1  g2037(.din(new_new_n4273__), .dout(n7505));
  not1  g2038(.din(new_new_n4487__), .dout(n7508));
  buf1  g2039(.din(new_new_n4404__), .dout(n7511));
  buf1  g2040(.din(new_new_n4275__), .dout(n7514));
  buf1  g2041(.din(new_new_n4274__), .dout(n7517));
  buf1  g2042(.din(new_new_n4588__), .dout(n7520));
  buf1  g2043(.din(new_new_n4549__), .dout(n7523));
  buf1  g2044(.din(new_new_n4544__), .dout(n7526));
  buf1  g2045(.din(new_new_n4548__), .dout(n7529));
  not1  g2046(.din(new_new_n4457__), .dout(n7532));
  not1  g2047(.din(new_new_n4469__), .dout(n7535));
  buf1  g2048(.din(new_new_n4587__), .dout(n7538));
  buf1  g2049(.din(new_new_n4468__), .dout(n7541));
  buf1  g2050(.din(new_new_n4419__), .dout(n7544));
  buf1  g2051(.din(new_new_n4444__), .dout(n7547));
  buf1  g2052(.din(new_new_n4434__), .dout(n7550));
  buf1  g2053(.din(new_new_n4447__), .dout(n7553));
  buf1  g2054(.din(new_new_n4446__), .dout(n7556));
  buf1  g2055(.din(new_new_n4448__), .dout(n7559));
  buf1  g2056(.din(new_new_n4456__), .dout(n7562));
  not1  g2057(.din(new_new_n4484__), .dout(n7565));
  not1  g2058(.din(new_new_n4497__), .dout(n7568));
  buf1  g2059(.din(new_new_n4589__), .dout(n7571));
  buf1  g2060(.din(new_new_n4584__), .dout(n7574));
  buf1  g2061(.din(new_new_n4586__), .dout(n7577));
  buf1  g2062(.din(new_new_n4583__), .dout(n7580));
  buf1  g2063(.din(new_new_n4585__), .dout(n7583));
  buf1  g2064(.din(new_new_n4593__), .dout(n7586));
  buf1  g2065(.din(new_new_n4551__), .dout(n7589));
  buf1  g2066(.din(new_new_n3167__), .dout(n7592));
  buf1  g2067(.din(new_new_n3168__), .dout(n7595));
  buf1  g2068(.din(new_new_n3169__), .dout(n7598));
  buf1  g2069(.din(new_new_n3170__), .dout(n7601));
  buf1  g2070(.din(new_new_n3171__), .dout(n7604));
  buf1  g2071(.din(new_new_n3172__), .dout(n7607));
  buf1  g2072(.din(new_new_n3173__), .dout(n7610));
  not1  g2073(.din(new_new_n3177__), .dout(n7613));
  buf1  g2074(.din(new_new_n3178__), .dout(n7616));
  not1  g2075(.din(new_new_n3179__), .dout(n7619));
  not1  g2076(.din(new_new_n3183__), .dout(n7622));
  buf1  g2077(.din(new_new_n3184__), .dout(n7625));
  buf1  g2078(.din(new_new_n3188__), .dout(n7628));
  not1  g2079(.din(new_new_n3189__), .dout(n7631));
  buf1  g2080(.din(new_new_n3193__), .dout(n7634));
  not1  g2081(.din(new_new_n3194__), .dout(n7637));
  buf1  g2082(.din(new_new_n3195__), .dout(n7640));
  buf1  g2083(.din(new_new_n3196__), .dout(n7643));
  buf1  g2084(.din(new_new_n3200__), .dout(n7646));
  not1  g2085(.din(new_new_n3201__), .dout(n7649));
  buf1  g2086(.din(new_new_n3202__), .dout(n7652));
  not1  g2087(.din(new_new_n3203__), .dout(n7655));
  buf1  g2088(.din(new_new_n3204__), .dout(n7658));
  not1  g2089(.din(new_new_n3205__), .dout(n7661));
  buf1  g2090(.din(new_new_n3206__), .dout(n7664));
  buf1  g2091(.din(new_new_n3207__), .dout(n7667));
  buf1  g2092(.din(new_new_n3208__), .dout(n7670));
  buf1  g2093(.din(new_new_n3209__), .dout(n7673));
  buf1  g2094(.din(new_new_n3210__), .dout(n7676));
  not1  g2095(.din(new_new_n4582__), .dout(n7679));
  buf1  g2096(.din(new_new_n3214__), .dout(n7682));
  not1  g2097(.din(new_new_n3215__), .dout(n7685));
  buf1  g2098(.din(new_new_n3218__), .dout(n7688));
  buf1  g2099(.din(new_new_n3227__), .dout(n7691));
  buf1  g2100(.din(new_new_n3232__), .dout(n7694));
  buf1  g2101(.din(new_new_n3235__), .dout(n7697));
  buf1  g2102(.din(new_new_n3238__), .dout(n7700));
  buf1  g2103(.din(new_new_n3241__), .dout(n7703));
  not1  g2104(.din(new_new_n3242__), .dout(n7706));
  buf1  g2105(.din(new_new_n3245__), .dout(n7709));
  buf1  g2106(.din(new_new_n3248__), .dout(n7712));
  not1  g2107(.din(new_new_n3249__), .dout(n7715));
  buf1  g2108(.din(new_new_n3252__), .dout(n7718));
  not1  g2109(.din(new_new_n3253__), .dout(n7721));
  not1  g2110(.din(new_new_n3270__), .dout(n7724));
  not1  g2111(.din(new_new_n3272__), .dout(n7727));
  not1  g2112(.din(new_new_n3288__), .dout(n7730));
  buf1  g2113(.din(new_new_n3289__), .dout(n7733));
  not1  g2114(.din(new_new_n3293__), .dout(n7736));
  not1  g2115(.din(new_new_n3294__), .dout(n7739));
  buf1  g2116(.din(new_new_n3309__), .dout(n7742));
  buf1  g2117(.din(new_new_n3324__), .dout(n7745));
  buf1  g2118(.din(new_new_n3333__), .dout(n7748));
  buf1  g2119(.din(new_new_n3360__), .dout(n7751));
  buf1  g2120(.din(new_new_n3367__), .dout(n7754));
  not1  g2121(.din(new_new_n3368__), .dout(n7757));
  buf1  g2122(.din(new_new_n3395__), .dout(n7760));
  not1  g2123(.din(new_new_n4581__), .dout(n7763));
  buf1  g2124(.din(new_new_n4598__), .dout(n7766));
  buf1  g2125(.din(new_new_n1738__), .dout(n7769));
  buf1  g2126(.din(new_new_n1932__), .dout(n7772));
  buf1  g2127(.din(new_new_n1936__), .dout(n7775));
  buf1  g2128(.din(new_new_n1946__), .dout(n7778));
  buf1  g2129(.din(new_new_n2026__), .dout(n7781));
  buf1  g2130(.din(new_new_n2072__), .dout(n7784));
  buf1  g2131(.din(new_new_n2108__), .dout(n7787));
  buf1  g2132(.din(new_new_n2144__), .dout(n7790));
  buf1  g2133(.din(new_new_n2180__), .dout(n7793));
  buf1  g2134(.din(new_new_n2410__), .dout(n7796));
  buf1  g2135(.din(new_new_n2414__), .dout(n7799));
  buf1  g2136(.din(new_new_n2430__), .dout(n7802));
  buf1  g2137(.din(new_new_n2434__), .dout(n7805));
  buf1  g2138(.din(new_new_n3403__), .dout(n7808));
  buf1  g2139(.din(new_new_n3404__), .dout(n7811));
  buf1  g2140(.din(new_new_n3405__), .dout(n7814));
  buf1  g2141(.din(new_new_n3406__), .dout(n7817));
  buf1  g2142(.din(new_new_n3407__), .dout(n7820));
  buf1  g2143(.din(new_new_n3408__), .dout(n7823));
  buf1  g2144(.din(new_new_n3409__), .dout(n7826));
  buf1  g2145(.din(new_new_n3410__), .dout(n7829));
  buf1  g2146(.din(new_new_n3411__), .dout(n7832));
  buf1  g2147(.din(new_new_n3412__), .dout(n7835));
  buf1  g2148(.din(new_new_n3414__), .dout(n7838));
  buf1  g2149(.din(new_new_n3416__), .dout(n7841));
  buf1  g2150(.din(new_new_n3420__), .dout(n7844));
  buf1  g2151(.din(new_new_n3424__), .dout(n7847));
  buf1  g2152(.din(new_new_n4601__), .dout(n7850));
  buf1  g2153(.din(new_new_n2236__), .dout(n7853));
  buf1  g2154(.din(new_new_n3427__), .dout(n7856));
  buf1  g2155(.din(new_new_n3430__), .dout(n7859));
  buf1  g2156(.din(new_new_n3433__), .dout(n7862));
  buf1  g2157(.din(new_new_n3436__), .dout(n7865));
  buf1  g2158(.din(new_new_n3439__), .dout(n7868));
  buf1  g2159(.din(new_new_n3442__), .dout(n7871));
  buf1  g2160(.din(new_new_n3451__), .dout(n7874));
  buf1  g2161(.din(new_new_n3460__), .dout(n7877));
  buf1  g2162(.din(new_new_n3469__), .dout(n7880));
  buf1  g2163(.din(new_new_n3473__), .dout(n7883));
  buf1  g2164(.din(new_new_n3482__), .dout(n7886));
  buf1  g2165(.din(new_new_n3486__), .dout(n7889));
  not1  g2166(.din(new_new_n3487__), .dout(n7892));
  buf1  g2167(.din(new_new_n3490__), .dout(n7895));
  buf1  g2168(.din(new_new_n3493__), .dout(n7898));
  buf1  g2169(.din(new_new_n3499__), .dout(n7901));
  not1  g2170(.din(new_new_n4604__), .dout(n7904));
  not1  g2171(.din(new_new_n4603__), .dout(n7907));
  buf1  g2172(.din(new_new_n1908__), .dout(n7910));
  buf1  g2173(.din(new_new_n1956__), .dout(n7913));
  buf1  g2174(.din(new_new_n1876__), .dout(n7916));
  buf1  g2175(.din(new_new_n1914__), .dout(n7919));
  buf1  g2176(.din(new_new_n1920__), .dout(n7922));
  buf1  g2177(.din(new_new_n2000__), .dout(n7925));
  buf1  g2178(.din(new_new_n2044__), .dout(n7928));
  buf1  g2179(.din(new_new_n2280__), .dout(n7931));
  buf1  g2180(.din(new_new_n3508__), .dout(n7934));
  buf1  g2181(.din(new_new_n3509__), .dout(n7937));
  buf1  g2182(.din(new_new_n3510__), .dout(n7940));
  buf1  g2183(.din(new_new_n3511__), .dout(n7943));
  not1  g2184(.din(new_new_n3512__), .dout(n7946));
  buf1  g2185(.din(new_new_n3521__), .dout(n7949));
  buf1  g2186(.din(new_new_n1528__), .dout(n7952));
  buf1  g2187(.din(new_new_n1530__), .dout(n7955));
  buf1  g2188(.din(new_new_n1548__), .dout(n7958));
  buf1  g2189(.din(new_new_n1550__), .dout(n7961));
  buf1  g2190(.din(new_new_n1568__), .dout(n7964));
  buf1  g2191(.din(new_new_n1570__), .dout(n7967));
  buf1  g2192(.din(new_new_n1588__), .dout(n7970));
  buf1  g2193(.din(new_new_n1590__), .dout(n7973));
  buf1  g2194(.din(new_new_n1660__), .dout(n7976));
  buf1  g2195(.din(new_new_n2245__), .dout(new_new_n4161__));
  buf1  g2196(.din(new_new_n2209__), .dout(new_new_n4162__));
  buf1  g2197(.din(new_new_n4162__), .dout(new_new_n4163__));
  buf1  g2198(.din(new_new_n4162__), .dout(new_new_n4164__));
  buf1  g2199(.din(new_new_n2840__), .dout(new_new_n4165__));
  buf1  g2200(.din(new_new_n4165__), .dout(new_new_n4166__));
  buf1  g2201(.din(new_new_n2844__), .dout(new_new_n4167__));
  buf1  g2202(.din(new_new_n2843__), .dout(new_new_n4168__));
  buf1  g2203(.din(new_new_n2253__), .dout(new_new_n4169__));
  buf1  g2204(.din(new_new_n4169__), .dout(new_new_n4170__));
  buf1  g2205(.din(new_new_n2848__), .dout(new_new_n4171__));
  buf1  g2206(.din(new_new_n4171__), .dout(new_new_n4172__));
  buf1  g2207(.din(new_new_n2855__), .dout(new_new_n4173__));
  buf1  g2208(.din(new_new_n2469__), .dout(new_new_n4174__));
  buf1  g2209(.din(new_new_n2260__), .dout(new_new_n4175__));
  buf1  g2210(.din(new_new_n4175__), .dout(new_new_n4176__));
  buf1  g2211(.din(new_new_n4175__), .dout(new_new_n4177__));
  buf1  g2212(.din(new_new_n2470__), .dout(new_new_n4178__));
  buf1  g2213(.din(new_new_n2261__), .dout(new_new_n4179__));
  buf1  g2214(.din(new_new_n4179__), .dout(new_new_n4180__));
  buf1  g2215(.din(new_new_n4179__), .dout(new_new_n4181__));
  buf1  g2216(.din(new_new_n2852__), .dout(new_new_n4182__));
  buf1  g2217(.din(new_new_n2226__), .dout(new_new_n4183__));
  buf1  g2218(.din(new_new_n2468__), .dout(new_new_n4184__));
  buf1  g2219(.din(new_new_n2591__), .dout(new_new_n4185__));
  buf1  g2220(.din(new_new_n4185__), .dout(new_new_n4186__));
  buf1  g2221(.din(new_new_n2657__), .dout(new_new_n4187__));
  buf1  g2222(.din(new_new_n2652__), .dout(new_new_n4188__));
  buf1  g2223(.din(new_new_n2656__), .dout(new_new_n4189__));
  buf1  g2224(.din(new_new_n2653__), .dout(new_new_n4190__));
  buf1  g2225(.din(new_new_n2680__), .dout(new_new_n4191__));
  buf1  g2226(.din(new_new_n2651__), .dout(new_new_n4192__));
  buf1  g2227(.din(new_new_n2681__), .dout(new_new_n4193__));
  buf1  g2228(.din(new_new_n2650__), .dout(new_new_n4194__));
  buf1  g2229(.din(new_new_n2482__), .dout(new_new_n4195__));
  buf1  g2230(.din(new_new_n1875__), .dout(new_new_n4196__));
  buf1  g2231(.din(new_new_n2590__), .dout(new_new_n4197__));
  buf1  g2232(.din(new_new_n2563__), .dout(new_new_n4198__));
  buf1  g2233(.din(new_new_n2562__), .dout(new_new_n4199__));
  buf1  g2234(.din(new_new_n2963__), .dout(new_new_n4200__));
  buf1  g2235(.din(new_new_n2964__), .dout(new_new_n4201__));
  buf1  g2236(.din(new_new_n2985__), .dout(new_new_n4202__));
  buf1  g2237(.din(new_new_n2992__), .dout(new_new_n4203__));
  buf1  g2238(.din(new_new_n2668__), .dout(new_new_n4204__));
  buf1  g2239(.din(new_new_n2994__), .dout(new_new_n4205__));
  buf1  g2240(.din(new_new_n2993__), .dout(new_new_n4206__));
  buf1  g2241(.din(new_new_n2884__), .dout(new_new_n4207__));
  buf1  g2242(.din(new_new_n2877__), .dout(new_new_n4208__));
  buf1  g2243(.din(new_new_n2899__), .dout(new_new_n4209__));
  buf1  g2244(.din(new_new_n2961__), .dout(new_new_n4210__));
  buf1  g2245(.din(new_new_n2981__), .dout(new_new_n4211__));
  buf1  g2246(.din(new_new_n2516__), .dout(new_new_n4212__));
  buf1  g2247(.din(new_new_n4212__), .dout(new_new_n4213__));
  buf1  g2248(.din(new_new_n4212__), .dout(new_new_n4214__));
  buf1  g2249(.din(new_new_n2517__), .dout(new_new_n4215__));
  buf1  g2250(.din(new_new_n4215__), .dout(new_new_n4216__));
  buf1  g2251(.din(new_new_n4215__), .dout(new_new_n4217__));
  buf1  g2252(.din(new_new_n2494__), .dout(new_new_n4218__));
  buf1  g2253(.din(new_new_n4218__), .dout(new_new_n4219__));
  buf1  g2254(.din(new_new_n4219__), .dout(new_new_n4220__));
  buf1  g2255(.din(new_new_n4219__), .dout(new_new_n4221__));
  buf1  g2256(.din(new_new_n4218__), .dout(new_new_n4222__));
  buf1  g2257(.din(new_new_n4222__), .dout(new_new_n4223__));
  buf1  g2258(.din(new_new_n4222__), .dout(new_new_n4224__));
  buf1  g2259(.din(new_new_n2495__), .dout(new_new_n4225__));
  buf1  g2260(.din(new_new_n4225__), .dout(new_new_n4226__));
  buf1  g2261(.din(new_new_n4226__), .dout(new_new_n4227__));
  buf1  g2262(.din(new_new_n4226__), .dout(new_new_n4228__));
  buf1  g2263(.din(new_new_n4225__), .dout(new_new_n4229__));
  buf1  g2264(.din(new_new_n4229__), .dout(new_new_n4230__));
  buf1  g2265(.din(new_new_n4229__), .dout(new_new_n4231__));
  buf1  g2266(.din(new_new_n2572__), .dout(new_new_n4232__));
  buf1  g2267(.din(new_new_n4232__), .dout(new_new_n4233__));
  buf1  g2268(.din(new_new_n2570__), .dout(new_new_n4234__));
  buf1  g2269(.din(new_new_n4234__), .dout(new_new_n4235__));
  buf1  g2270(.din(new_new_n2573__), .dout(new_new_n4236__));
  buf1  g2271(.din(new_new_n4236__), .dout(new_new_n4237__));
  buf1  g2272(.din(new_new_n2571__), .dout(new_new_n4238__));
  buf1  g2273(.din(new_new_n4238__), .dout(new_new_n4239__));
  buf1  g2274(.din(new_new_n3019__), .dout(new_new_n4240__));
  buf1  g2275(.din(new_new_n3013__), .dout(new_new_n4241__));
  buf1  g2276(.din(new_new_n2499__), .dout(new_new_n4242__));
  buf1  g2277(.din(new_new_n4242__), .dout(new_new_n4243__));
  buf1  g2278(.din(new_new_n4243__), .dout(new_new_n4244__));
  buf1  g2279(.din(new_new_n4243__), .dout(new_new_n4245__));
  buf1  g2280(.din(new_new_n4242__), .dout(new_new_n4246__));
  buf1  g2281(.din(new_new_n2498__), .dout(new_new_n4247__));
  buf1  g2282(.din(new_new_n4247__), .dout(new_new_n4248__));
  buf1  g2283(.din(new_new_n4248__), .dout(new_new_n4249__));
  buf1  g2284(.din(new_new_n4248__), .dout(new_new_n4250__));
  buf1  g2285(.din(new_new_n4247__), .dout(new_new_n4251__));
  buf1  g2286(.din(new_new_n3033__), .dout(new_new_n4252__));
  buf1  g2287(.din(new_new_n3023__), .dout(new_new_n4253__));
  buf1  g2288(.din(new_new_n2497__), .dout(new_new_n4254__));
  buf1  g2289(.din(new_new_n2496__), .dout(new_new_n4255__));
  buf1  g2290(.din(new_new_n3022__), .dout(new_new_n4256__));
  buf1  g2291(.din(new_new_n4256__), .dout(new_new_n4257__));
  buf1  g2292(.din(new_new_n2565__), .dout(new_new_n4258__));
  buf1  g2293(.din(new_new_n3021__), .dout(new_new_n4259__));
  buf1  g2294(.din(new_new_n2564__), .dout(new_new_n4260__));
  buf1  g2295(.din(new_new_n4260__), .dout(new_new_n4261__));
  buf1  g2296(.din(new_new_n4260__), .dout(new_new_n4262__));
  buf1  g2297(.din(new_new_n2379__), .dout(new_new_n4263__));
  buf1  g2298(.din(new_new_n2371__), .dout(new_new_n4264__));
  buf1  g2299(.din(new_new_n4264__), .dout(new_new_n4265__));
  buf1  g2300(.din(new_new_n2485__), .dout(new_new_n4266__));
  buf1  g2301(.din(new_new_n4266__), .dout(new_new_n4267__));
  buf1  g2302(.din(new_new_n4266__), .dout(new_new_n4268__));
  buf1  g2303(.din(new_new_n2484__), .dout(new_new_n4269__));
  buf1  g2304(.din(new_new_n4269__), .dout(new_new_n4270__));
  buf1  g2305(.din(new_new_n4269__), .dout(new_new_n4271__));
  buf1  g2306(.din(new_new_n2814__), .dout(new_new_n4272__));
  buf1  g2307(.din(new_new_n2816__), .dout(new_new_n4273__));
  buf1  g2308(.din(new_new_n3100__), .dout(new_new_n4274__));
  buf1  g2309(.din(new_new_n3098__), .dout(new_new_n4275__));
  buf1  g2310(.din(new_new_n3038__), .dout(new_new_n4276__));
  buf1  g2311(.din(new_new_n4276__), .dout(new_new_n4277__));
  buf1  g2312(.din(new_new_n4276__), .dout(new_new_n4278__));
  buf1  g2313(.din(new_new_n2697__), .dout(new_new_n4279__));
  buf1  g2314(.din(new_new_n3106__), .dout(new_new_n4280__));
  buf1  g2315(.din(new_new_n4280__), .dout(new_new_n4281__));
  buf1  g2316(.din(new_new_n4281__), .dout(new_new_n4282__));
  buf1  g2317(.din(new_new_n4280__), .dout(new_new_n4283__));
  buf1  g2318(.din(new_new_n2322__), .dout(new_new_n4284__));
  buf1  g2319(.din(new_new_n4284__), .dout(new_new_n4285__));
  buf1  g2320(.din(new_new_n3105__), .dout(new_new_n4286__));
  buf1  g2321(.din(new_new_n4286__), .dout(new_new_n4287__));
  buf1  g2322(.din(new_new_n4287__), .dout(new_new_n4288__));
  buf1  g2323(.din(new_new_n4286__), .dout(new_new_n4289__));
  buf1  g2324(.din(new_new_n3071__), .dout(new_new_n4290__));
  buf1  g2325(.din(new_new_n1768__), .dout(new_new_n4291__));
  buf1  g2326(.din(new_new_n4291__), .dout(new_new_n4292__));
  buf1  g2327(.din(new_new_n4292__), .dout(new_new_n4293__));
  buf1  g2328(.din(new_new_n4293__), .dout(new_new_n4294__));
  buf1  g2329(.din(new_new_n4292__), .dout(new_new_n4295__));
  buf1  g2330(.din(new_new_n4291__), .dout(new_new_n4296__));
  buf1  g2331(.din(new_new_n4296__), .dout(new_new_n4297__));
  buf1  g2332(.din(new_new_n4296__), .dout(new_new_n4298__));
  buf1  g2333(.din(new_new_n2576__), .dout(new_new_n4299__));
  buf1  g2334(.din(new_new_n4299__), .dout(new_new_n4300__));
  buf1  g2335(.din(new_new_n4300__), .dout(new_new_n4301__));
  buf1  g2336(.din(new_new_n4299__), .dout(new_new_n4302__));
  buf1  g2337(.din(new_new_n1769__), .dout(new_new_n4303__));
  buf1  g2338(.din(new_new_n4303__), .dout(new_new_n4304__));
  buf1  g2339(.din(new_new_n4304__), .dout(new_new_n4305__));
  buf1  g2340(.din(new_new_n4305__), .dout(new_new_n4306__));
  buf1  g2341(.din(new_new_n4304__), .dout(new_new_n4307__));
  buf1  g2342(.din(new_new_n4303__), .dout(new_new_n4308__));
  buf1  g2343(.din(new_new_n4308__), .dout(new_new_n4309__));
  buf1  g2344(.din(new_new_n4308__), .dout(new_new_n4310__));
  buf1  g2345(.din(new_new_n3072__), .dout(new_new_n4311__));
  buf1  g2346(.din(new_new_n4311__), .dout(new_new_n4312__));
  buf1  g2347(.din(new_new_n3047__), .dout(new_new_n4313__));
  buf1  g2348(.din(new_new_n4313__), .dout(new_new_n4314__));
  buf1  g2349(.din(new_new_n1834__), .dout(new_new_n4315__));
  buf1  g2350(.din(new_new_n4315__), .dout(new_new_n4316__));
  buf1  g2351(.din(new_new_n4316__), .dout(new_new_n4317__));
  buf1  g2352(.din(new_new_n4316__), .dout(new_new_n4318__));
  buf1  g2353(.din(new_new_n4315__), .dout(new_new_n4319__));
  buf1  g2354(.din(new_new_n4319__), .dout(new_new_n4320__));
  buf1  g2355(.din(new_new_n4319__), .dout(new_new_n4321__));
  buf1  g2356(.din(new_new_n2520__), .dout(new_new_n4322__));
  buf1  g2357(.din(new_new_n4322__), .dout(new_new_n4323__));
  buf1  g2358(.din(new_new_n4322__), .dout(new_new_n4324__));
  buf1  g2359(.din(new_new_n1835__), .dout(new_new_n4325__));
  buf1  g2360(.din(new_new_n4325__), .dout(new_new_n4326__));
  buf1  g2361(.din(new_new_n4326__), .dout(new_new_n4327__));
  buf1  g2362(.din(new_new_n4326__), .dout(new_new_n4328__));
  buf1  g2363(.din(new_new_n4325__), .dout(new_new_n4329__));
  buf1  g2364(.din(new_new_n4329__), .dout(new_new_n4330__));
  buf1  g2365(.din(new_new_n4329__), .dout(new_new_n4331__));
  buf1  g2366(.din(new_new_n2766__), .dout(new_new_n4332__));
  buf1  g2367(.din(new_new_n4332__), .dout(new_new_n4333__));
  buf1  g2368(.din(new_new_n2518__), .dout(new_new_n4334__));
  buf1  g2369(.din(new_new_n4334__), .dout(new_new_n4335__));
  buf1  g2370(.din(new_new_n2696__), .dout(new_new_n4336__));
  buf1  g2371(.din(new_new_n3127__), .dout(new_new_n4337__));
  buf1  g2372(.din(new_new_n4337__), .dout(new_new_n4338__));
  buf1  g2373(.din(new_new_n4337__), .dout(new_new_n4339__));
  buf1  g2374(.din(new_new_n2303__), .dout(new_new_n4340__));
  buf1  g2375(.din(new_new_n4340__), .dout(new_new_n4341__));
  buf1  g2376(.din(new_new_n4341__), .dout(new_new_n4342__));
  buf1  g2377(.din(new_new_n4340__), .dout(new_new_n4343__));
  buf1  g2378(.din(new_new_n3129__), .dout(new_new_n4344__));
  buf1  g2379(.din(new_new_n4344__), .dout(new_new_n4345__));
  buf1  g2380(.din(new_new_n4344__), .dout(new_new_n4346__));
  buf1  g2381(.din(new_new_n3137__), .dout(new_new_n4347__));
  buf1  g2382(.din(new_new_n4347__), .dout(new_new_n4348__));
  buf1  g2383(.din(new_new_n4347__), .dout(new_new_n4349__));
  buf1  g2384(.din(new_new_n3136__), .dout(new_new_n4350__));
  buf1  g2385(.din(new_new_n4350__), .dout(new_new_n4351__));
  buf1  g2386(.din(new_new_n2543__), .dout(new_new_n4352__));
  buf1  g2387(.din(new_new_n2542__), .dout(new_new_n4353__));
  buf1  g2388(.din(new_new_n4353__), .dout(new_new_n4354__));
  buf1  g2389(.din(new_new_n2774__), .dout(new_new_n4355__));
  buf1  g2390(.din(new_new_n4355__), .dout(new_new_n4356__));
  buf1  g2391(.din(new_new_n4356__), .dout(new_new_n4357__));
  buf1  g2392(.din(new_new_n4356__), .dout(new_new_n4358__));
  buf1  g2393(.din(new_new_n4355__), .dout(new_new_n4359__));
  buf1  g2394(.din(new_new_n2775__), .dout(new_new_n4360__));
  buf1  g2395(.din(new_new_n2577__), .dout(new_new_n4361__));
  buf1  g2396(.din(new_new_n3078__), .dout(new_new_n4362__));
  buf1  g2397(.din(new_new_n2752__), .dout(new_new_n4363__));
  buf1  g2398(.din(new_new_n4363__), .dout(new_new_n4364__));
  buf1  g2399(.din(new_new_n4364__), .dout(new_new_n4365__));
  buf1  g2400(.din(new_new_n4365__), .dout(new_new_n4366__));
  buf1  g2401(.din(new_new_n4365__), .dout(new_new_n4367__));
  buf1  g2402(.din(new_new_n4364__), .dout(new_new_n4368__));
  buf1  g2403(.din(new_new_n4368__), .dout(new_new_n4369__));
  buf1  g2404(.din(new_new_n4363__), .dout(new_new_n4370__));
  buf1  g2405(.din(new_new_n4370__), .dout(new_new_n4371__));
  buf1  g2406(.din(new_new_n4370__), .dout(new_new_n4372__));
  buf1  g2407(.din(new_new_n2812__), .dout(new_new_n4373__));
  buf1  g2408(.din(new_new_n4373__), .dout(new_new_n4374__));
  buf1  g2409(.din(new_new_n4374__), .dout(new_new_n4375__));
  buf1  g2410(.din(new_new_n4373__), .dout(new_new_n4376__));
  buf1  g2411(.din(new_new_n2753__), .dout(new_new_n4377__));
  buf1  g2412(.din(new_new_n4377__), .dout(new_new_n4378__));
  buf1  g2413(.din(new_new_n4378__), .dout(new_new_n4379__));
  buf1  g2414(.din(new_new_n4377__), .dout(new_new_n4380__));
  buf1  g2415(.din(new_new_n2750__), .dout(new_new_n4381__));
  buf1  g2416(.din(new_new_n4381__), .dout(new_new_n4382__));
  buf1  g2417(.din(new_new_n4382__), .dout(new_new_n4383__));
  buf1  g2418(.din(new_new_n4383__), .dout(new_new_n4384__));
  buf1  g2419(.din(new_new_n4383__), .dout(new_new_n4385__));
  buf1  g2420(.din(new_new_n4382__), .dout(new_new_n4386__));
  buf1  g2421(.din(new_new_n4381__), .dout(new_new_n4387__));
  buf1  g2422(.din(new_new_n4387__), .dout(new_new_n4388__));
  buf1  g2423(.din(new_new_n4387__), .dout(new_new_n4389__));
  buf1  g2424(.din(new_new_n2751__), .dout(new_new_n4390__));
  buf1  g2425(.din(new_new_n4390__), .dout(new_new_n4391__));
  buf1  g2426(.din(new_new_n4391__), .dout(new_new_n4392__));
  buf1  g2427(.din(new_new_n4392__), .dout(new_new_n4393__));
  buf1  g2428(.din(new_new_n4392__), .dout(new_new_n4394__));
  buf1  g2429(.din(new_new_n4391__), .dout(new_new_n4395__));
  buf1  g2430(.din(new_new_n4395__), .dout(new_new_n4396__));
  buf1  g2431(.din(new_new_n4395__), .dout(new_new_n4397__));
  buf1  g2432(.din(new_new_n4390__), .dout(new_new_n4398__));
  buf1  g2433(.din(new_new_n4398__), .dout(new_new_n4399__));
  buf1  g2434(.din(new_new_n4399__), .dout(new_new_n4400__));
  buf1  g2435(.din(new_new_n4399__), .dout(new_new_n4401__));
  buf1  g2436(.din(new_new_n4398__), .dout(new_new_n4402__));
  buf1  g2437(.din(new_new_n4402__), .dout(new_new_n4403__));
  buf1  g2438(.din(new_new_n3097__), .dout(new_new_n4404__));
  buf1  g2439(.din(new_new_n4404__), .dout(new_new_n4405__));
  buf1  g2440(.din(new_new_n2012__), .dout(new_new_n4406__));
  buf1  g2441(.din(new_new_n1884__), .dout(new_new_n4407__));
  buf1  g2442(.din(new_new_n1968__), .dout(new_new_n4408__));
  buf1  g2443(.din(new_new_n1926__), .dout(new_new_n4409__));
  buf1  g2444(.din(new_new_n2174__), .dout(new_new_n4410__));
  buf1  g2445(.din(new_new_n2066__), .dout(new_new_n4411__));
  buf1  g2446(.din(new_new_n2138__), .dout(new_new_n4412__));
  buf1  g2447(.din(new_new_n2102__), .dout(new_new_n4413__));
  buf1  g2448(.din(new_new_n2224__), .dout(new_new_n4414__));
  buf1  g2449(.din(new_new_n3176__), .dout(new_new_n4415__));
  buf1  g2450(.din(new_new_n2531__), .dout(new_new_n4416__));
  buf1  g2451(.din(new_new_n4416__), .dout(new_new_n4417__));
  buf1  g2452(.din(new_new_n4416__), .dout(new_new_n4418__));
  buf1  g2453(.din(new_new_n3111__), .dout(new_new_n4419__));
  buf1  g2454(.din(new_new_n2533__), .dout(new_new_n4420__));
  buf1  g2455(.din(new_new_n4420__), .dout(new_new_n4421__));
  buf1  g2456(.din(new_new_n3182__), .dout(new_new_n4422__));
  buf1  g2457(.din(new_new_n2567__), .dout(new_new_n4423__));
  buf1  g2458(.din(new_new_n4423__), .dout(new_new_n4424__));
  buf1  g2459(.din(new_new_n4423__), .dout(new_new_n4425__));
  buf1  g2460(.din(new_new_n3028__), .dout(new_new_n4426__));
  buf1  g2461(.din(new_new_n4426__), .dout(new_new_n4427__));
  buf1  g2462(.din(new_new_n4426__), .dout(new_new_n4428__));
  buf1  g2463(.din(new_new_n3187__), .dout(new_new_n4429__));
  buf1  g2464(.din(new_new_n2297__), .dout(new_new_n4430__));
  buf1  g2465(.din(new_new_n4430__), .dout(new_new_n4431__));
  buf1  g2466(.din(new_new_n4430__), .dout(new_new_n4432__));
  buf1  g2467(.din(new_new_n3192__), .dout(new_new_n4433__));
  buf1  g2468(.din(new_new_n3117__), .dout(new_new_n4434__));
  buf1  g2469(.din(new_new_n2309__), .dout(new_new_n4435__));
  buf1  g2470(.din(new_new_n4435__), .dout(new_new_n4436__));
  buf1  g2471(.din(new_new_n4435__), .dout(new_new_n4437__));
  buf1  g2472(.din(new_new_n3060__), .dout(new_new_n4438__));
  buf1  g2473(.din(new_new_n4438__), .dout(new_new_n4439__));
  buf1  g2474(.din(new_new_n3199__), .dout(new_new_n4440__));
  buf1  g2475(.din(new_new_n2317__), .dout(new_new_n4441__));
  buf1  g2476(.din(new_new_n4441__), .dout(new_new_n4442__));
  buf1  g2477(.din(new_new_n4441__), .dout(new_new_n4443__));
  buf1  g2478(.din(new_new_n3114__), .dout(new_new_n4444__));
  buf1  g2479(.din(new_new_n2323__), .dout(new_new_n4445__));
  buf1  g2480(.din(new_new_n3123__), .dout(new_new_n4446__));
  buf1  g2481(.din(new_new_n3120__), .dout(new_new_n4447__));
  buf1  g2482(.din(new_new_n3126__), .dout(new_new_n4448__));
  buf1  g2483(.din(new_new_n2386__), .dout(new_new_n4449__));
  buf1  g2484(.din(new_new_n2394__), .dout(new_new_n4450__));
  buf1  g2485(.din(new_new_n3059__), .dout(new_new_n4451__));
  buf1  g2486(.din(new_new_n3048__), .dout(new_new_n4452__));
  buf1  g2487(.din(new_new_n2778__), .dout(new_new_n4453__));
  buf1  g2488(.din(new_new_n4453__), .dout(new_new_n4454__));
  buf1  g2489(.din(new_new_n4453__), .dout(new_new_n4455__));
  buf1  g2490(.din(new_new_n3131__), .dout(new_new_n4456__));
  buf1  g2491(.din(new_new_n3104__), .dout(new_new_n4457__));
  buf1  g2492(.din(new_new_n2768__), .dout(new_new_n4458__));
  buf1  g2493(.din(new_new_n4458__), .dout(new_new_n4459__));
  buf1  g2494(.din(new_new_n3225__), .dout(new_new_n4460__));
  buf1  g2495(.din(new_new_n4460__), .dout(new_new_n4461__));
  buf1  g2496(.din(new_new_n4460__), .dout(new_new_n4462__));
  buf1  g2497(.din(new_new_n3017__), .dout(new_new_n4463__));
  buf1  g2498(.din(new_new_n3015__), .dout(new_new_n4464__));
  buf1  g2499(.din(new_new_n3230__), .dout(new_new_n4465__));
  buf1  g2500(.din(new_new_n4465__), .dout(new_new_n4466__));
  buf1  g2501(.din(new_new_n2568__), .dout(new_new_n4467__));
  buf1  g2502(.din(new_new_n3108__), .dout(new_new_n4468__));
  buf1  g2503(.din(new_new_n3107__), .dout(new_new_n4469__));
  buf1  g2504(.din(new_new_n2330__), .dout(new_new_n4470__));
  buf1  g2505(.din(new_new_n2331__), .dout(new_new_n4471__));
  buf1  g2506(.din(new_new_n2769__), .dout(new_new_n4472__));
  buf1  g2507(.din(new_new_n4472__), .dout(new_new_n4473__));
  buf1  g2508(.din(new_new_n3247__), .dout(new_new_n4474__));
  buf1  g2509(.din(new_new_n3246__), .dout(new_new_n4475__));
  buf1  g2510(.din(new_new_n2535__), .dout(new_new_n4476__));
  buf1  g2511(.din(new_new_n4476__), .dout(new_new_n4477__));
  buf1  g2512(.din(new_new_n3251__), .dout(new_new_n4478__));
  buf1  g2513(.din(new_new_n3250__), .dout(new_new_n4479__));
  buf1  g2514(.din(new_new_n3257__), .dout(new_new_n4480__));
  buf1  g2515(.din(new_new_n3254__), .dout(new_new_n4481__));
  buf1  g2516(.din(new_new_n2783__), .dout(new_new_n4482__));
  buf1  g2517(.din(new_new_n2781__), .dout(new_new_n4483__));
  buf1  g2518(.din(new_new_n3142__), .dout(new_new_n4484__));
  buf1  g2519(.din(new_new_n2378__), .dout(new_new_n4485__));
  buf1  g2520(.din(new_new_n2370__), .dout(new_new_n4486__));
  buf1  g2521(.din(new_new_n3079__), .dout(new_new_n4487__));
  buf1  g2522(.din(new_new_n3025__), .dout(new_new_n4488__));
  buf1  g2523(.din(new_new_n2459__), .dout(new_new_n4489__));
  buf1  g2524(.din(new_new_n2534__), .dout(new_new_n4490__));
  buf1  g2525(.din(new_new_n4490__), .dout(new_new_n4491__));
  buf1  g2526(.din(new_new_n2458__), .dout(new_new_n4492__));
  buf1  g2527(.din(new_new_n3287__), .dout(new_new_n4493__));
  buf1  g2528(.din(new_new_n3274__), .dout(new_new_n4494__));
  buf1  g2529(.din(new_new_n3036__), .dout(new_new_n4495__));
  buf1  g2530(.din(new_new_n3292__), .dout(new_new_n4496__));
  buf1  g2531(.din(new_new_n3151__), .dout(new_new_n4497__));
  buf1  g2532(.din(new_new_n4497__), .dout(new_new_n4498__));
  buf1  g2533(.din(new_new_n2447__), .dout(new_new_n4499__));
  buf1  g2534(.din(new_new_n2440__), .dout(new_new_n4500__));
  buf1  g2535(.din(new_new_n2446__), .dout(new_new_n4501__));
  buf1  g2536(.din(new_new_n2441__), .dout(new_new_n4502__));
  buf1  g2537(.din(new_new_n2530__), .dout(new_new_n4503__));
  buf1  g2538(.din(new_new_n2532__), .dout(new_new_n4504__));
  buf1  g2539(.din(new_new_n4504__), .dout(new_new_n4505__));
  buf1  g2540(.din(new_new_n2302__), .dout(new_new_n4506__));
  buf1  g2541(.din(new_new_n2308__), .dout(new_new_n4507__));
  buf1  g2542(.din(new_new_n4507__), .dout(new_new_n4508__));
  buf1  g2543(.din(new_new_n2453__), .dout(new_new_n4509__));
  buf1  g2544(.din(new_new_n2566__), .dout(new_new_n4510__));
  buf1  g2545(.din(new_new_n2452__), .dout(new_new_n4511__));
  buf1  g2546(.din(new_new_n2519__), .dout(new_new_n4512__));
  buf1  g2547(.din(new_new_n3229__), .dout(new_new_n4513__));
  buf1  g2548(.din(new_new_n2721__), .dout(new_new_n4514__));
  buf1  g2549(.din(new_new_n2718__), .dout(new_new_n4515__));
  buf1  g2550(.din(new_new_n2720__), .dout(new_new_n4516__));
  buf1  g2551(.din(new_new_n2719__), .dout(new_new_n4517__));
  buf1  g2552(.din(new_new_n2717__), .dout(new_new_n4518__));
  buf1  g2553(.din(new_new_n2714__), .dout(new_new_n4519__));
  buf1  g2554(.din(new_new_n2716__), .dout(new_new_n4520__));
  buf1  g2555(.din(new_new_n2715__), .dout(new_new_n4521__));
  buf1  g2556(.din(new_new_n3344__), .dout(new_new_n4522__));
  buf1  g2557(.din(new_new_n3338__), .dout(new_new_n4523__));
  buf1  g2558(.din(new_new_n3345__), .dout(new_new_n4524__));
  buf1  g2559(.din(new_new_n3339__), .dout(new_new_n4525__));
  buf1  g2560(.din(new_new_n2427__), .dout(new_new_n4526__));
  buf1  g2561(.din(new_new_n2420__), .dout(new_new_n4527__));
  buf1  g2562(.din(new_new_n2426__), .dout(new_new_n4528__));
  buf1  g2563(.din(new_new_n2421__), .dout(new_new_n4529__));
  buf1  g2564(.din(new_new_n3366__), .dout(new_new_n4530__));
  buf1  g2565(.din(new_new_n3363__), .dout(new_new_n4531__));
  buf1  g2566(.din(new_new_n2770__), .dout(new_new_n4532__));
  buf1  g2567(.din(new_new_n2771__), .dout(new_new_n4533__));
  buf1  g2568(.din(new_new_n2521__), .dout(new_new_n4534__));
  buf1  g2569(.din(new_new_n2767__), .dout(new_new_n4535__));
  buf1  g2570(.din(new_new_n3379__), .dout(new_new_n4536__));
  buf1  g2571(.din(new_new_n3373__), .dout(new_new_n4537__));
  buf1  g2572(.din(new_new_n3380__), .dout(new_new_n4538__));
  buf1  g2573(.din(new_new_n3374__), .dout(new_new_n4539__));
  buf1  g2574(.din(new_new_n3224__), .dout(new_new_n4540__));
  buf1  g2575(.din(new_new_n3103__), .dout(new_new_n4541__));
  buf1  g2576(.din(new_new_n4541__), .dout(new_new_n4542__));
  buf1  g2577(.din(new_new_n4541__), .dout(new_new_n4543__));
  buf1  g2578(.din(new_new_n2350__), .dout(new_new_n4544__));
  buf1  g2579(.din(new_new_n3102__), .dout(new_new_n4545__));
  buf1  g2580(.din(new_new_n4545__), .dout(new_new_n4546__));
  buf1  g2581(.din(new_new_n4546__), .dout(new_new_n4547__));
  buf1  g2582(.din(new_new_n4545__), .dout(new_new_n4548__));
  buf1  g2583(.din(new_new_n2276__), .dout(new_new_n4549__));
  buf1  g2584(.din(new_new_n3423__), .dout(new_new_n4550__));
  buf1  g2585(.din(new_new_n3166__), .dout(new_new_n4551__));
  buf1  g2586(.din(new_new_n4551__), .dout(new_new_n4552__));
  buf1  g2587(.din(new_new_n2575__), .dout(new_new_n4553__));
  buf1  g2588(.din(new_new_n4553__), .dout(new_new_n4554__));
  buf1  g2589(.din(new_new_n4554__), .dout(new_new_n4555__));
  buf1  g2590(.din(new_new_n4555__), .dout(new_new_n4556__));
  buf1  g2591(.din(new_new_n4555__), .dout(new_new_n4557__));
  buf1  g2592(.din(new_new_n4554__), .dout(new_new_n4558__));
  buf1  g2593(.din(new_new_n4558__), .dout(new_new_n4559__));
  buf1  g2594(.din(new_new_n4558__), .dout(new_new_n4560__));
  buf1  g2595(.din(new_new_n4553__), .dout(new_new_n4561__));
  buf1  g2596(.din(new_new_n4561__), .dout(new_new_n4562__));
  buf1  g2597(.din(new_new_n4561__), .dout(new_new_n4563__));
  buf1  g2598(.din(new_new_n2574__), .dout(new_new_n4564__));
  buf1  g2599(.din(new_new_n4564__), .dout(new_new_n4565__));
  buf1  g2600(.din(new_new_n4565__), .dout(new_new_n4566__));
  buf1  g2601(.din(new_new_n4566__), .dout(new_new_n4567__));
  buf1  g2602(.din(new_new_n4566__), .dout(new_new_n4568__));
  buf1  g2603(.din(new_new_n4565__), .dout(new_new_n4569__));
  buf1  g2604(.din(new_new_n4569__), .dout(new_new_n4570__));
  buf1  g2605(.din(new_new_n4569__), .dout(new_new_n4571__));
  buf1  g2606(.din(new_new_n4564__), .dout(new_new_n4572__));
  buf1  g2607(.din(new_new_n4572__), .dout(new_new_n4573__));
  buf1  g2608(.din(new_new_n4573__), .dout(new_new_n4574__));
  buf1  g2609(.din(new_new_n4572__), .dout(new_new_n4575__));
  buf1  g2610(.din(new_new_n2694__), .dout(new_new_n4576__));
  buf1  g2611(.din(new_new_n4576__), .dout(new_new_n4577__));
  buf1  g2612(.din(new_new_n4576__), .dout(new_new_n4578__));
  buf1  g2613(.din(new_new_n2695__), .dout(new_new_n4579__));
  buf1  g2614(.din(new_new_n4579__), .dout(new_new_n4580__));
  buf1  g2615(.din(new_new_n3402__), .dout(new_new_n4581__));
  buf1  g2616(.din(new_new_n3211__), .dout(new_new_n4582__));
  buf1  g2617(.din(new_new_n2356__), .dout(new_new_n4583__));
  buf1  g2618(.din(new_new_n2284__), .dout(new_new_n4584__));
  buf1  g2619(.din(new_new_n2362__), .dout(new_new_n4585__));
  buf1  g2620(.din(new_new_n2288__), .dout(new_new_n4586__));
  buf1  g2621(.din(new_new_n2336__), .dout(new_new_n4587__));
  buf1  g2622(.din(new_new_n2272__), .dout(new_new_n4588__));
  buf1  g2623(.din(new_new_n3157__), .dout(new_new_n4589__));
  buf1  g2624(.din(new_new_n2834__), .dout(new_new_n4590__));
  buf1  g2625(.din(new_new_n4590__), .dout(new_new_n4591__));
  buf1  g2626(.din(new_new_n4591__), .dout(new_new_n4592__));
  buf1  g2627(.din(new_new_n4590__), .dout(new_new_n4593__));
  buf1  g2628(.din(new_new_n2835__), .dout(new_new_n4594__));
  buf1  g2629(.din(new_new_n4594__), .dout(new_new_n4595__));
  buf1  g2630(.din(new_new_n4594__), .dout(new_new_n4596__));
  buf1  g2631(.din(new_new_n2399__), .dout(new_new_n4597__));
  buf1  g2632(.din(new_new_n2398__), .dout(new_new_n4598__));
  buf1  g2633(.din(new_new_n4598__), .dout(new_new_n4599__));
  buf1  g2634(.din(new_new_n2219__), .dout(new_new_n4600__));
  buf1  g2635(.din(new_new_n2218__), .dout(new_new_n4601__));
  buf1  g2636(.din(new_new_n4601__), .dout(new_new_n4602__));
  buf1  g2637(.din(new_new_n3507__), .dout(new_new_n4603__));
  buf1  g2638(.din(new_new_n3503__), .dout(new_new_n4604__));
  buf1  g2639(.din(new_new_n2269__), .dout(new_new_n4605__));
  buf1  g2640(.din(new_new_n2347__), .dout(new_new_n4606__));
  buf1  g2641(.din(new_new_n4606__), .dout(new_new_n4607__));
  buf1  g2642(.din(new_new_n2845__), .dout(new_new_n4608__));
  buf1  g2643(.din(new_new_n2861__), .dout(new_new_n4609__));
  buf1  g2644(.din(new_new_n2864__), .dout(new_new_n4610__));
  buf1  g2645(.din(new_new_n2869__), .dout(new_new_n4611__));
  buf1  g2646(.din(new_new_n2949__), .dout(new_new_n4612__));
  buf1  g2647(.din(new_new_n2975__), .dout(new_new_n4613__));
  buf1  g2648(.din(new_new_n3012__), .dout(new_new_n4614__));
  zero1 g2649(.dout(new_new_n4615__));
  always @ (posedge clock) begin
    n1416_lo <= n6254;
    n1419_lo <= n6257;
    n1422_lo <= n6260;
    n1425_lo <= n6263;
    n1428_lo <= n6266;
    n1431_lo <= n6269;
    n1434_lo <= n6272;
    n1437_lo <= n6275;
    n1440_lo <= n6278;
    n1443_lo <= n6281;
    n1446_lo <= n6284;
    n1449_lo <= n6287;
    n1452_lo <= n6290;
    n1455_lo <= n6293;
    n1458_lo <= n6296;
    n1464_lo <= n6299;
    n1467_lo <= n6302;
    n1470_lo <= n6305;
    n1476_lo <= n6308;
    n1479_lo <= n6311;
    n1482_lo <= n6314;
    n1488_lo <= n6317;
    n1491_lo <= n6320;
    n1494_lo <= n6323;
    n1497_lo <= n6326;
    n1500_lo <= n6329;
    n1503_lo <= n6332;
    n1512_lo <= n6335;
    n1515_lo <= n6338;
    n1518_lo <= n6341;
    n1521_lo <= n6344;
    n1524_lo <= n6347;
    n1527_lo <= n6350;
    n1530_lo <= n6353;
    n1533_lo <= n6356;
    n1536_lo <= n6359;
    n1539_lo <= n6362;
    n1542_lo <= n6365;
    n1545_lo <= n6368;
    n1548_lo <= n6371;
    n1551_lo <= n6374;
    n1554_lo <= n6377;
    n1560_lo <= n6380;
    n1563_lo <= n6383;
    n1566_lo <= n6386;
    n1572_lo <= n6389;
    n1575_lo <= n6392;
    n1578_lo <= n6395;
    n1584_lo <= n6398;
    n1587_lo <= n6401;
    n1590_lo <= n6404;
    n1596_lo <= n6407;
    n1599_lo <= n6410;
    n1602_lo <= n6413;
    n1608_lo <= n6416;
    n1611_lo <= n6419;
    n1614_lo <= n6422;
    n1620_lo <= n6425;
    n1623_lo <= n6428;
    n1626_lo <= n6431;
    n1632_lo <= n6434;
    n1635_lo <= n6437;
    n1638_lo <= n6440;
    n1644_lo <= n6443;
    n1647_lo <= n6446;
    n1650_lo <= n6449;
    n1656_lo <= n6452;
    n1659_lo <= n6455;
    n1662_lo <= n6458;
    n1668_lo <= n6461;
    n1671_lo <= n6464;
    n1674_lo <= n6467;
    n1680_lo <= n6470;
    n1683_lo <= n6473;
    n1686_lo <= n6476;
    n1692_lo <= n6479;
    n1695_lo <= n6482;
    n1698_lo <= n6485;
    n1704_lo <= n6488;
    n1707_lo <= n6491;
    n1710_lo <= n6494;
    n1716_lo <= n6497;
    n1719_lo <= n6500;
    n1722_lo <= n6503;
    n1728_lo <= n6506;
    n1731_lo <= n6509;
    n1734_lo <= n6512;
    n1740_lo <= n6515;
    n1743_lo <= n6518;
    n1746_lo <= n6521;
    n1749_lo <= n6524;
    n1752_lo <= n6527;
    n1755_lo <= n6530;
    n1758_lo <= n6533;
    n1761_lo <= n6536;
    n1764_lo <= n6539;
    n1776_lo <= n6542;
    n1788_lo <= n6545;
    n1791_lo <= n6548;
    n1794_lo <= n6551;
    n1797_lo <= n6554;
    n1800_lo <= n6557;
    n1803_lo <= n6560;
    n1812_lo <= n6563;
    n1815_lo <= n6566;
    n1824_lo <= n6569;
    n1827_lo <= n6572;
    n1836_lo <= n6575;
    n1839_lo <= n6578;
    n1848_lo <= n6581;
    n1851_lo <= n6584;
    n1860_lo <= n6587;
    n1872_lo <= n6590;
    n1875_lo <= n6593;
    n1884_lo <= n6596;
    n1896_lo <= n6599;
    n1899_lo <= n6602;
    n1908_lo <= n6605;
    n1920_lo <= n6608;
    n1923_lo <= n6611;
    n1926_lo <= n6614;
    n1929_lo <= n6617;
    n1932_lo <= n6620;
    n1935_lo <= n6623;
    n1944_lo <= n6626;
    n1947_lo <= n6629;
    n1956_lo <= n6632;
    n1959_lo <= n6635;
    n1962_lo <= n6638;
    n1968_lo <= n6641;
    n1971_lo <= n6644;
    n1980_lo <= n6647;
    n1983_lo <= n6650;
    n1992_lo <= n6653;
    n1995_lo <= n6656;
    n2004_lo <= n6659;
    n2016_lo <= n6662;
    n2019_lo <= n6665;
    n2028_lo <= n6668;
    n2040_lo <= n6671;
    n2043_lo <= n6674;
    n2046_lo <= n6677;
    n2049_lo <= n6680;
    n2052_lo <= n6683;
    n2055_lo <= n6686;
    n2064_lo <= n6689;
    n2067_lo <= n6692;
    n2076_lo <= n6695;
    n2079_lo <= n6698;
    n2088_lo <= n6701;
    n2091_lo <= n6704;
    n2100_lo <= n6707;
    n2103_lo <= n6710;
    n2112_lo <= n6713;
    n2115_lo <= n6716;
    n2124_lo <= n6719;
    n2127_lo <= n6722;
    n2136_lo <= n6725;
    n2148_lo <= n6728;
    n2151_lo <= n6731;
    n2160_lo <= n6734;
    n2172_lo <= n6737;
    n2175_lo <= n6740;
    n2178_lo <= n6743;
    n2181_lo <= n6746;
    n2184_lo <= n6749;
    n2187_lo <= n6752;
    n2196_lo <= n6755;
    n2199_lo <= n6758;
    n2208_lo <= n6761;
    n2211_lo <= n6764;
    n2220_lo <= n6767;
    n2223_lo <= n6770;
    n2232_lo <= n6773;
    n2235_lo <= n6776;
    n2244_lo <= n6779;
    n2247_lo <= n6782;
    n2256_lo <= n6785;
    n2259_lo <= n6788;
    n2268_lo <= n6791;
    n2280_lo <= n6794;
    n2283_lo <= n6797;
    n2292_lo <= n6800;
    n2295_lo <= n6803;
    n2298_lo <= n6806;
    n2301_lo <= n6809;
    n2304_lo <= n6812;
    n2307_lo <= n6815;
    n2316_lo <= n6818;
    n2319_lo <= n6821;
    n2322_lo <= n6824;
    n2325_lo <= n6827;
    n2328_lo <= n6830;
    n2331_lo <= n6833;
    n2340_lo <= n6836;
    n2343_lo <= n6839;
    n2376_lo <= n6842;
    n2379_lo <= n6845;
    n2388_lo <= n6848;
    n2391_lo <= n6851;
    n2400_lo <= n6854;
    n2403_lo <= n6857;
    n2412_lo <= n6860;
    n2415_lo <= n6863;
    n2424_lo <= n6866;
    n2427_lo <= n6869;
    n2436_lo <= n6872;
    n2439_lo <= n6875;
    n2442_lo <= n6878;
    n2445_lo <= n6881;
    n2448_lo <= n6884;
    n2451_lo <= n6887;
    n2460_lo <= n6890;
    n2463_lo <= n6893;
    n2496_lo <= n6896;
    n2499_lo <= n6899;
    n2508_lo <= n6902;
    n2511_lo <= n6905;
    n2520_lo <= n6908;
    n2523_lo <= n6911;
    n2532_lo <= n6914;
    n2535_lo <= n6917;
    n2544_lo <= n6920;
    n2547_lo <= n6923;
    n2556_lo <= n6926;
    n2559_lo <= n6929;
    n2562_lo <= n6932;
    n2565_lo <= n6935;
    n2568_lo <= n6938;
    n2571_lo <= n6941;
    n2580_lo <= n6944;
    n2583_lo <= n6947;
    n2616_lo <= n6950;
    n2619_lo <= n6953;
    n2628_lo <= n6956;
    n2631_lo <= n6959;
    n2640_lo <= n6962;
    n2643_lo <= n6965;
    n2652_lo <= n6968;
    n2655_lo <= n6971;
    n2664_lo <= n6974;
    n2667_lo <= n6977;
    n2676_lo <= n6980;
    n2679_lo <= n6983;
    n2682_lo <= n6986;
    n2685_lo <= n6989;
    n2688_lo <= n6992;
    n2691_lo <= n6995;
    n2700_lo <= n6998;
    n2703_lo <= n7001;
    n2736_lo <= n7004;
    n2739_lo <= n7007;
    n2748_lo <= n7010;
    n2751_lo <= n7013;
    n2760_lo <= n7016;
    n2763_lo <= n7019;
    n2772_lo <= n7022;
    n2775_lo <= n7025;
    n2784_lo <= n7028;
    n2787_lo <= n7031;
    n2790_lo <= n7034;
    n2793_lo <= n7037;
    n2796_lo <= n7040;
    n2799_lo <= n7043;
    n2802_lo <= n7046;
    n2805_lo <= n7049;
    n2808_lo <= n7052;
    n2820_lo <= n7055;
    n2823_lo <= n7058;
    n2826_lo <= n7061;
    n2829_lo <= n7064;
    n2832_lo <= n7067;
    n2835_lo <= n7070;
    n2838_lo <= n7073;
    n2841_lo <= n7076;
    n2844_lo <= n7079;
    n2856_lo <= n7082;
    n2859_lo <= n7085;
    n2862_lo <= n7088;
    n2865_lo <= n7091;
    n2868_lo <= n7094;
    n2871_lo <= n7097;
    n2874_lo <= n7100;
    n2877_lo <= n7103;
    n2880_lo <= n7106;
    n2883_lo <= n7109;
    n2886_lo <= n7112;
    n2889_lo <= n7115;
    n2892_lo <= n7118;
    n2895_lo <= n7121;
    n2898_lo <= n7124;
    n2901_lo <= n7127;
    n2904_lo <= n7130;
    n2907_lo <= n7133;
    n2916_lo <= n7136;
    n2919_lo <= n7139;
    n2925_lo <= n7142;
    n2928_lo <= n7145;
    n2940_lo <= n7148;
    n2943_lo <= n7151;
    n2952_lo <= n7154;
    n2955_lo <= n7157;
    n2961_lo <= n7160;
    n2964_lo <= n7163;
    n2967_lo <= n7166;
    n2970_lo <= n7169;
    n2976_lo <= n7172;
    n2979_lo <= n7175;
    n2982_lo <= n7178;
    n2988_lo <= n7181;
    n2991_lo <= n7184;
    n2994_lo <= n7187;
    n2997_lo <= n7190;
    n3000_lo <= n7193;
    n3003_lo <= n7196;
    n3006_lo <= n7199;
    n3012_lo <= n7202;
    n3015_lo <= n7205;
    n3018_lo <= n7208;
    n3021_lo <= n7211;
    n3024_lo <= n7214;
    n3027_lo <= n7217;
    n3030_lo <= n7220;
    n3033_lo <= n7223;
    n3036_lo <= n7226;
    n3039_lo <= n7229;
    n3045_lo <= n7232;
    n3048_lo <= n7235;
    n3051_lo <= n7238;
    n3054_lo <= n7241;
    n3057_lo <= n7244;
    n3060_lo <= n7247;
    n3063_lo <= n7250;
    n3069_lo <= n7253;
    n3072_lo <= n7256;
    n3075_lo <= n7259;
    n3081_lo <= n7262;
    n3084_lo <= n7265;
    n3087_lo <= n7268;
    n3093_lo <= n7271;
    n3096_lo <= n7274;
    n3099_lo <= n7277;
    n3102_lo <= n7280;
    n3105_lo <= n7283;
    n3108_lo <= n7286;
    n3111_lo <= n7289;
    n3114_lo <= n7292;
    n3117_lo <= n7295;
    n3120_lo <= n7298;
    n3123_lo <= n7301;
    n3126_lo <= n7304;
    n3129_lo <= n7307;
    n3132_lo <= n7310;
    n3135_lo <= n7313;
    n3138_lo <= n7316;
    n3141_lo <= n7319;
    n3156_lo <= n7322;
    n3168_lo <= n7325;
    n3171_lo <= n7328;
    n3174_lo <= n7331;
    n3177_lo <= n7334;
    n3180_lo <= n7337;
    n3183_lo <= n7340;
    n3192_lo <= n7343;
    n3195_lo <= n7346;
    n3204_lo <= n7349;
    n3207_lo <= n7352;
    n3210_lo <= n7355;
    n3216_lo <= n7358;
    n3219_lo <= n7361;
    n3222_lo <= n7364;
    n3228_lo <= n7367;
    n3231_lo <= n7370;
    n3240_lo <= n7373;
    n3243_lo <= n7376;
    n3252_lo <= n7379;
    n3255_lo <= n7382;
    n3258_lo <= n7385;
    n3264_lo <= n7388;
    n3267_lo <= n7391;
    n3270_lo <= n7394;
    n3276_lo <= n7397;
    n3279_lo <= n7400;
    n3282_lo <= n7403;
    n3288_lo <= n7406;
    n3291_lo <= n7409;
    n3294_lo <= n7412;
    n3603_o2 <= n7415;
    n3604_o2 <= n7418;
    n1391_inv <= n7421;
    n3798_o2 <= n7424;
    n3846_o2 <= n7427;
    n4019_o2 <= n7430;
    n4017_o2 <= n7433;
    n2177_o2 <= n7436;
    n2150_o2 <= n7439;
    n2154_o2 <= n7442;
    n2184_o2 <= n7445;
    n2515_o2 <= n7448;
    n3837_o2 <= n7451;
    n2167_o2 <= n7454;
    n2118_o2 <= n7457;
    n2186_o2 <= n7460;
    n2174_o2 <= n7463;
    n3964_o2 <= n7466;
    n4005_o2 <= n7469;
    n4006_o2 <= n7472;
    n1445_inv <= n7475;
    n2176_o2 <= n7478;
    n2227_o2 <= n7481;
    n2236_o2 <= n7484;
    n2245_o2 <= n7487;
    n2518_o2 <= n7490;
    n4023_o2 <= n7493;
    n1466_inv <= n7496;
    n4038_o2 <= n7499;
    n4039_o2 <= n7502;
    n1475_inv <= n7505;
    n2119_o2 <= n7508;
    n2275_o2 <= n7511;
    n2595_o2 <= n7514;
    n2594_o2 <= n7517;
    lo498_buf_o2 <= n7520;
    lo502_buf_o2 <= n7523;
    lo550_buf_o2 <= n7526;
    n2596_o2 <= n7529;
    n2593_o2 <= n7532;
    n2668_o2 <= n7535;
    lo542_buf_o2 <= n7538;
    n2667_o2 <= n7541;
    n2404_o2 <= n7544;
    n2410_o2 <= n7547;
    n2419_o2 <= n7550;
    n2392_o2 <= n7553;
    n2369_o2 <= n7556;
    n2397_o2 <= n7559;
    n2601_o2 <= n7562;
    n2658_o2 <= n7565;
    n2574_o2 <= n7568;
    n2205_o2 <= n7571;
    lo510_buf_o2 <= n7574;
    lo514_buf_o2 <= n7577;
    lo554_buf_o2 <= n7580;
    lo558_buf_o2 <= n7583;
    lo578_buf_o2 <= n7586;
    n2254_o2 <= n7589;
    n2421_o2 <= n7592;
    n2422_o2 <= n7595;
    n2130_o2 <= n7598;
    n2127_o2 <= n7601;
    n2131_o2 <= n7604;
    n2128_o2 <= n7607;
    n2264_o2 <= n7610;
    n2467_o2 <= n7613;
    n2471_o2 <= n7616;
    n2488_o2 <= n7619;
    n2478_o2 <= n7622;
    n2486_o2 <= n7625;
    n2485_o2 <= n7628;
    n2498_o2 <= n7631;
    n2495_o2 <= n7634;
    n2496_o2 <= n7637;
    n2458_o2 <= n7640;
    n2643_o2 <= n7643;
    n2462_o2 <= n7646;
    n2468_o2 <= n7649;
    n2639_o2 <= n7652;
    n2499_o2 <= n7655;
    n2472_o2 <= n7658;
    n2474_o2 <= n7661;
    n2489_o2 <= n7664;
    n2321_o2 <= n7667;
    n2322_o2 <= n7670;
    n2640_o2 <= n7673;
    n2642_o2 <= n7676;
    n2187_o2 <= n7679;
    n2373_o2 <= n7682;
    n2603_o2 <= n7685;
    n2388_o2 <= n7688;
    n2437_o2 <= n7691;
    n2356_o2 <= n7694;
    n2452_o2 <= n7697;
    n2347_o2 <= n7700;
    n2329_o2 <= n7703;
    n2669_o2 <= n7706;
    n2332_o2 <= n7709;
    n2664_o2 <= n7712;
    n2665_o2 <= n7715;
    n2653_o2 <= n7718;
    n2654_o2 <= n7721;
    n2636_o2 <= n7724;
    n2660_o2 <= n7727;
    n2318_o2 <= n7730;
    n2319_o2 <= n7733;
    n2586_o2 <= n7736;
    n2587_o2 <= n7739;
    n2288_o2 <= n7742;
    n2344_o2 <= n7745;
    n2530_o2 <= n7748;
    n2303_o2 <= n7751;
    n2566_o2 <= n7754;
    n2567_o2 <= n7757;
    n2554_o2 <= n7760;
    n2194_o2 <= n7763;
    lo582_buf_o2 <= n7766;
    lo030_buf_o2 <= n7769;
    lo174_buf_o2 <= n7772;
    lo178_buf_o2 <= n7775;
    lo186_buf_o2 <= n7778;
    lo266_buf_o2 <= n7781;
    lo306_buf_o2 <= n7784;
    lo346_buf_o2 <= n7787;
    lo386_buf_o2 <= n7790;
    lo426_buf_o2 <= n7793;
    lo590_buf_o2 <= n7796;
    lo594_buf_o2 <= n7799;
    lo606_buf_o2 <= n7802;
    lo610_buf_o2 <= n7805;
    n2238_o2 <= n7808;
    n2229_o2 <= n7811;
    n2242_o2 <= n7814;
    n2233_o2 <= n7817;
    n2168_o2 <= n7820;
    n2237_o2 <= n7823;
    n2228_o2 <= n7826;
    n2172_o2 <= n7829;
    n2223_o2 <= n7832;
    n2222_o2 <= n7835;
    n2170_o2 <= n7838;
    n2181_o2 <= n7841;
    n2510_o2 <= n7844;
    n2621_o2 <= n7847;
    lo466_buf_o2 <= n7850;
    lo478_buf_o2 <= n7853;
    n2149_o2 <= n7856;
    n2429_o2 <= n7859;
    n2444_o2 <= n7862;
    n2153_o2 <= n7865;
    n2433_o2 <= n7868;
    n2448_o2 <= n7871;
    n2367_o2 <= n7874;
    n2386_o2 <= n7877;
    n2539_o2 <= n7880;
    n2183_o2 <= n7883;
    n2220_o2 <= n7886;
    n2514_o2 <= n7889;
    n2196_o2 <= n7892;
    n2616_o2 <= n7895;
    n2612_o2 <= n7898;
    n2627_o2 <= n7901;
    n2140_o2 <= n7904;
    n1877_inv <= n7907;
    lo149_buf_o2 <= n7910;
    lo197_buf_o2 <= n7913;
    lo118_buf_o2 <= n7916;
    lo158_buf_o2 <= n7919;
    lo166_buf_o2 <= n7922;
    lo242_buf_o2 <= n7925;
    lo286_buf_o2 <= n7928;
    lo506_buf_o2 <= n7931;
    n2198_o2 <= n7934;
    n2202_o2 <= n7937;
    n2197_o2 <= n7940;
    n1913_inv <= n7943;
    n2146_o2 <= n7946;
    n1919_inv <= n7949;
    lo312_buf_o2 <= n7952;
    lo316_buf_o2 <= n7955;
    lo352_buf_o2 <= n7958;
    lo356_buf_o2 <= n7961;
    lo392_buf_o2 <= n7964;
    lo396_buf_o2 <= n7967;
    lo432_buf_o2 <= n7970;
    lo436_buf_o2 <= n7973;
    lo576_buf_o2 <= n7976;
  end
  initial begin
    n1416_lo <= 1'b0;
    n1419_lo <= 1'b0;
    n1422_lo <= 1'b0;
    n1425_lo <= 1'b0;
    n1428_lo <= 1'b0;
    n1431_lo <= 1'b0;
    n1434_lo <= 1'b0;
    n1437_lo <= 1'b0;
    n1440_lo <= 1'b0;
    n1443_lo <= 1'b0;
    n1446_lo <= 1'b0;
    n1449_lo <= 1'b0;
    n1452_lo <= 1'b0;
    n1455_lo <= 1'b0;
    n1458_lo <= 1'b0;
    n1464_lo <= 1'b0;
    n1467_lo <= 1'b0;
    n1470_lo <= 1'b0;
    n1476_lo <= 1'b0;
    n1479_lo <= 1'b0;
    n1482_lo <= 1'b0;
    n1488_lo <= 1'b0;
    n1491_lo <= 1'b0;
    n1494_lo <= 1'b0;
    n1497_lo <= 1'b0;
    n1500_lo <= 1'b0;
    n1503_lo <= 1'b0;
    n1512_lo <= 1'b0;
    n1515_lo <= 1'b0;
    n1518_lo <= 1'b0;
    n1521_lo <= 1'b0;
    n1524_lo <= 1'b0;
    n1527_lo <= 1'b0;
    n1530_lo <= 1'b0;
    n1533_lo <= 1'b0;
    n1536_lo <= 1'b0;
    n1539_lo <= 1'b0;
    n1542_lo <= 1'b0;
    n1545_lo <= 1'b0;
    n1548_lo <= 1'b0;
    n1551_lo <= 1'b0;
    n1554_lo <= 1'b0;
    n1560_lo <= 1'b0;
    n1563_lo <= 1'b0;
    n1566_lo <= 1'b0;
    n1572_lo <= 1'b0;
    n1575_lo <= 1'b0;
    n1578_lo <= 1'b0;
    n1584_lo <= 1'b0;
    n1587_lo <= 1'b0;
    n1590_lo <= 1'b0;
    n1596_lo <= 1'b0;
    n1599_lo <= 1'b0;
    n1602_lo <= 1'b0;
    n1608_lo <= 1'b0;
    n1611_lo <= 1'b0;
    n1614_lo <= 1'b0;
    n1620_lo <= 1'b0;
    n1623_lo <= 1'b0;
    n1626_lo <= 1'b0;
    n1632_lo <= 1'b0;
    n1635_lo <= 1'b0;
    n1638_lo <= 1'b0;
    n1644_lo <= 1'b0;
    n1647_lo <= 1'b0;
    n1650_lo <= 1'b0;
    n1656_lo <= 1'b0;
    n1659_lo <= 1'b0;
    n1662_lo <= 1'b0;
    n1668_lo <= 1'b0;
    n1671_lo <= 1'b0;
    n1674_lo <= 1'b0;
    n1680_lo <= 1'b0;
    n1683_lo <= 1'b0;
    n1686_lo <= 1'b0;
    n1692_lo <= 1'b0;
    n1695_lo <= 1'b0;
    n1698_lo <= 1'b0;
    n1704_lo <= 1'b0;
    n1707_lo <= 1'b0;
    n1710_lo <= 1'b0;
    n1716_lo <= 1'b0;
    n1719_lo <= 1'b0;
    n1722_lo <= 1'b0;
    n1728_lo <= 1'b0;
    n1731_lo <= 1'b0;
    n1734_lo <= 1'b0;
    n1740_lo <= 1'b0;
    n1743_lo <= 1'b0;
    n1746_lo <= 1'b0;
    n1749_lo <= 1'b0;
    n1752_lo <= 1'b0;
    n1755_lo <= 1'b0;
    n1758_lo <= 1'b0;
    n1761_lo <= 1'b0;
    n1764_lo <= 1'b0;
    n1776_lo <= 1'b0;
    n1788_lo <= 1'b0;
    n1791_lo <= 1'b0;
    n1794_lo <= 1'b0;
    n1797_lo <= 1'b0;
    n1800_lo <= 1'b0;
    n1803_lo <= 1'b0;
    n1812_lo <= 1'b0;
    n1815_lo <= 1'b0;
    n1824_lo <= 1'b0;
    n1827_lo <= 1'b0;
    n1836_lo <= 1'b0;
    n1839_lo <= 1'b0;
    n1848_lo <= 1'b0;
    n1851_lo <= 1'b0;
    n1860_lo <= 1'b0;
    n1872_lo <= 1'b0;
    n1875_lo <= 1'b0;
    n1884_lo <= 1'b0;
    n1896_lo <= 1'b0;
    n1899_lo <= 1'b0;
    n1908_lo <= 1'b0;
    n1920_lo <= 1'b0;
    n1923_lo <= 1'b0;
    n1926_lo <= 1'b0;
    n1929_lo <= 1'b0;
    n1932_lo <= 1'b0;
    n1935_lo <= 1'b0;
    n1944_lo <= 1'b0;
    n1947_lo <= 1'b0;
    n1956_lo <= 1'b0;
    n1959_lo <= 1'b0;
    n1962_lo <= 1'b0;
    n1968_lo <= 1'b0;
    n1971_lo <= 1'b0;
    n1980_lo <= 1'b0;
    n1983_lo <= 1'b0;
    n1992_lo <= 1'b0;
    n1995_lo <= 1'b0;
    n2004_lo <= 1'b0;
    n2016_lo <= 1'b0;
    n2019_lo <= 1'b0;
    n2028_lo <= 1'b0;
    n2040_lo <= 1'b0;
    n2043_lo <= 1'b0;
    n2046_lo <= 1'b0;
    n2049_lo <= 1'b0;
    n2052_lo <= 1'b0;
    n2055_lo <= 1'b0;
    n2064_lo <= 1'b0;
    n2067_lo <= 1'b0;
    n2076_lo <= 1'b0;
    n2079_lo <= 1'b0;
    n2088_lo <= 1'b0;
    n2091_lo <= 1'b0;
    n2100_lo <= 1'b0;
    n2103_lo <= 1'b0;
    n2112_lo <= 1'b0;
    n2115_lo <= 1'b0;
    n2124_lo <= 1'b0;
    n2127_lo <= 1'b0;
    n2136_lo <= 1'b0;
    n2148_lo <= 1'b0;
    n2151_lo <= 1'b0;
    n2160_lo <= 1'b0;
    n2172_lo <= 1'b0;
    n2175_lo <= 1'b0;
    n2178_lo <= 1'b0;
    n2181_lo <= 1'b0;
    n2184_lo <= 1'b0;
    n2187_lo <= 1'b0;
    n2196_lo <= 1'b0;
    n2199_lo <= 1'b0;
    n2208_lo <= 1'b0;
    n2211_lo <= 1'b0;
    n2220_lo <= 1'b0;
    n2223_lo <= 1'b0;
    n2232_lo <= 1'b0;
    n2235_lo <= 1'b0;
    n2244_lo <= 1'b0;
    n2247_lo <= 1'b0;
    n2256_lo <= 1'b0;
    n2259_lo <= 1'b0;
    n2268_lo <= 1'b0;
    n2280_lo <= 1'b0;
    n2283_lo <= 1'b0;
    n2292_lo <= 1'b0;
    n2295_lo <= 1'b0;
    n2298_lo <= 1'b0;
    n2301_lo <= 1'b0;
    n2304_lo <= 1'b0;
    n2307_lo <= 1'b0;
    n2316_lo <= 1'b0;
    n2319_lo <= 1'b0;
    n2322_lo <= 1'b0;
    n2325_lo <= 1'b0;
    n2328_lo <= 1'b0;
    n2331_lo <= 1'b0;
    n2340_lo <= 1'b0;
    n2343_lo <= 1'b0;
    n2376_lo <= 1'b0;
    n2379_lo <= 1'b0;
    n2388_lo <= 1'b0;
    n2391_lo <= 1'b0;
    n2400_lo <= 1'b0;
    n2403_lo <= 1'b0;
    n2412_lo <= 1'b0;
    n2415_lo <= 1'b0;
    n2424_lo <= 1'b0;
    n2427_lo <= 1'b0;
    n2436_lo <= 1'b0;
    n2439_lo <= 1'b0;
    n2442_lo <= 1'b0;
    n2445_lo <= 1'b0;
    n2448_lo <= 1'b0;
    n2451_lo <= 1'b0;
    n2460_lo <= 1'b0;
    n2463_lo <= 1'b0;
    n2496_lo <= 1'b0;
    n2499_lo <= 1'b0;
    n2508_lo <= 1'b0;
    n2511_lo <= 1'b0;
    n2520_lo <= 1'b0;
    n2523_lo <= 1'b0;
    n2532_lo <= 1'b0;
    n2535_lo <= 1'b0;
    n2544_lo <= 1'b0;
    n2547_lo <= 1'b0;
    n2556_lo <= 1'b0;
    n2559_lo <= 1'b0;
    n2562_lo <= 1'b0;
    n2565_lo <= 1'b0;
    n2568_lo <= 1'b0;
    n2571_lo <= 1'b0;
    n2580_lo <= 1'b0;
    n2583_lo <= 1'b0;
    n2616_lo <= 1'b0;
    n2619_lo <= 1'b0;
    n2628_lo <= 1'b0;
    n2631_lo <= 1'b0;
    n2640_lo <= 1'b0;
    n2643_lo <= 1'b0;
    n2652_lo <= 1'b0;
    n2655_lo <= 1'b0;
    n2664_lo <= 1'b0;
    n2667_lo <= 1'b0;
    n2676_lo <= 1'b0;
    n2679_lo <= 1'b0;
    n2682_lo <= 1'b0;
    n2685_lo <= 1'b0;
    n2688_lo <= 1'b0;
    n2691_lo <= 1'b0;
    n2700_lo <= 1'b0;
    n2703_lo <= 1'b0;
    n2736_lo <= 1'b0;
    n2739_lo <= 1'b0;
    n2748_lo <= 1'b0;
    n2751_lo <= 1'b0;
    n2760_lo <= 1'b0;
    n2763_lo <= 1'b0;
    n2772_lo <= 1'b0;
    n2775_lo <= 1'b0;
    n2784_lo <= 1'b0;
    n2787_lo <= 1'b0;
    n2790_lo <= 1'b0;
    n2793_lo <= 1'b0;
    n2796_lo <= 1'b0;
    n2799_lo <= 1'b0;
    n2802_lo <= 1'b0;
    n2805_lo <= 1'b0;
    n2808_lo <= 1'b0;
    n2820_lo <= 1'b0;
    n2823_lo <= 1'b0;
    n2826_lo <= 1'b0;
    n2829_lo <= 1'b0;
    n2832_lo <= 1'b0;
    n2835_lo <= 1'b0;
    n2838_lo <= 1'b0;
    n2841_lo <= 1'b0;
    n2844_lo <= 1'b0;
    n2856_lo <= 1'b0;
    n2859_lo <= 1'b0;
    n2862_lo <= 1'b0;
    n2865_lo <= 1'b0;
    n2868_lo <= 1'b0;
    n2871_lo <= 1'b0;
    n2874_lo <= 1'b0;
    n2877_lo <= 1'b0;
    n2880_lo <= 1'b0;
    n2883_lo <= 1'b0;
    n2886_lo <= 1'b0;
    n2889_lo <= 1'b0;
    n2892_lo <= 1'b0;
    n2895_lo <= 1'b0;
    n2898_lo <= 1'b0;
    n2901_lo <= 1'b0;
    n2904_lo <= 1'b0;
    n2907_lo <= 1'b0;
    n2916_lo <= 1'b0;
    n2919_lo <= 1'b0;
    n2925_lo <= 1'b0;
    n2928_lo <= 1'b0;
    n2940_lo <= 1'b0;
    n2943_lo <= 1'b0;
    n2952_lo <= 1'b0;
    n2955_lo <= 1'b0;
    n2961_lo <= 1'b0;
    n2964_lo <= 1'b0;
    n2967_lo <= 1'b0;
    n2970_lo <= 1'b0;
    n2976_lo <= 1'b0;
    n2979_lo <= 1'b0;
    n2982_lo <= 1'b0;
    n2988_lo <= 1'b0;
    n2991_lo <= 1'b0;
    n2994_lo <= 1'b0;
    n2997_lo <= 1'b0;
    n3000_lo <= 1'b0;
    n3003_lo <= 1'b0;
    n3006_lo <= 1'b0;
    n3012_lo <= 1'b0;
    n3015_lo <= 1'b0;
    n3018_lo <= 1'b0;
    n3021_lo <= 1'b0;
    n3024_lo <= 1'b0;
    n3027_lo <= 1'b0;
    n3030_lo <= 1'b0;
    n3033_lo <= 1'b0;
    n3036_lo <= 1'b0;
    n3039_lo <= 1'b0;
    n3045_lo <= 1'b0;
    n3048_lo <= 1'b0;
    n3051_lo <= 1'b0;
    n3054_lo <= 1'b0;
    n3057_lo <= 1'b0;
    n3060_lo <= 1'b0;
    n3063_lo <= 1'b0;
    n3069_lo <= 1'b0;
    n3072_lo <= 1'b0;
    n3075_lo <= 1'b0;
    n3081_lo <= 1'b0;
    n3084_lo <= 1'b0;
    n3087_lo <= 1'b0;
    n3093_lo <= 1'b0;
    n3096_lo <= 1'b0;
    n3099_lo <= 1'b0;
    n3102_lo <= 1'b0;
    n3105_lo <= 1'b0;
    n3108_lo <= 1'b0;
    n3111_lo <= 1'b0;
    n3114_lo <= 1'b0;
    n3117_lo <= 1'b0;
    n3120_lo <= 1'b0;
    n3123_lo <= 1'b0;
    n3126_lo <= 1'b0;
    n3129_lo <= 1'b0;
    n3132_lo <= 1'b0;
    n3135_lo <= 1'b0;
    n3138_lo <= 1'b0;
    n3141_lo <= 1'b0;
    n3156_lo <= 1'b0;
    n3168_lo <= 1'b0;
    n3171_lo <= 1'b0;
    n3174_lo <= 1'b0;
    n3177_lo <= 1'b0;
    n3180_lo <= 1'b0;
    n3183_lo <= 1'b0;
    n3192_lo <= 1'b0;
    n3195_lo <= 1'b0;
    n3204_lo <= 1'b0;
    n3207_lo <= 1'b0;
    n3210_lo <= 1'b0;
    n3216_lo <= 1'b0;
    n3219_lo <= 1'b0;
    n3222_lo <= 1'b0;
    n3228_lo <= 1'b0;
    n3231_lo <= 1'b0;
    n3240_lo <= 1'b0;
    n3243_lo <= 1'b0;
    n3252_lo <= 1'b0;
    n3255_lo <= 1'b0;
    n3258_lo <= 1'b0;
    n3264_lo <= 1'b0;
    n3267_lo <= 1'b0;
    n3270_lo <= 1'b0;
    n3276_lo <= 1'b0;
    n3279_lo <= 1'b0;
    n3282_lo <= 1'b0;
    n3288_lo <= 1'b0;
    n3291_lo <= 1'b0;
    n3294_lo <= 1'b0;
    n3603_o2 <= 1'b0;
    n3604_o2 <= 1'b0;
    n1391_inv <= 1'b0;
    n3798_o2 <= 1'b0;
    n3846_o2 <= 1'b0;
    n4019_o2 <= 1'b0;
    n4017_o2 <= 1'b0;
    n2177_o2 <= 1'b0;
    n2150_o2 <= 1'b0;
    n2154_o2 <= 1'b0;
    n2184_o2 <= 1'b0;
    n2515_o2 <= 1'b0;
    n3837_o2 <= 1'b0;
    n2167_o2 <= 1'b0;
    n2118_o2 <= 1'b0;
    n2186_o2 <= 1'b0;
    n2174_o2 <= 1'b0;
    n3964_o2 <= 1'b0;
    n4005_o2 <= 1'b0;
    n4006_o2 <= 1'b0;
    n1445_inv <= 1'b0;
    n2176_o2 <= 1'b0;
    n2227_o2 <= 1'b0;
    n2236_o2 <= 1'b0;
    n2245_o2 <= 1'b0;
    n2518_o2 <= 1'b0;
    n4023_o2 <= 1'b0;
    n1466_inv <= 1'b0;
    n4038_o2 <= 1'b0;
    n4039_o2 <= 1'b0;
    n1475_inv <= 1'b0;
    n2119_o2 <= 1'b0;
    n2275_o2 <= 1'b0;
    n2595_o2 <= 1'b0;
    n2594_o2 <= 1'b0;
    lo498_buf_o2 <= 1'b0;
    lo502_buf_o2 <= 1'b0;
    lo550_buf_o2 <= 1'b0;
    n2596_o2 <= 1'b0;
    n2593_o2 <= 1'b0;
    n2668_o2 <= 1'b0;
    lo542_buf_o2 <= 1'b0;
    n2667_o2 <= 1'b0;
    n2404_o2 <= 1'b0;
    n2410_o2 <= 1'b0;
    n2419_o2 <= 1'b0;
    n2392_o2 <= 1'b0;
    n2369_o2 <= 1'b0;
    n2397_o2 <= 1'b0;
    n2601_o2 <= 1'b0;
    n2658_o2 <= 1'b0;
    n2574_o2 <= 1'b0;
    n2205_o2 <= 1'b0;
    lo510_buf_o2 <= 1'b0;
    lo514_buf_o2 <= 1'b0;
    lo554_buf_o2 <= 1'b0;
    lo558_buf_o2 <= 1'b0;
    lo578_buf_o2 <= 1'b0;
    n2254_o2 <= 1'b0;
    n2421_o2 <= 1'b0;
    n2422_o2 <= 1'b0;
    n2130_o2 <= 1'b0;
    n2127_o2 <= 1'b0;
    n2131_o2 <= 1'b0;
    n2128_o2 <= 1'b0;
    n2264_o2 <= 1'b0;
    n2467_o2 <= 1'b0;
    n2471_o2 <= 1'b0;
    n2488_o2 <= 1'b0;
    n2478_o2 <= 1'b0;
    n2486_o2 <= 1'b0;
    n2485_o2 <= 1'b0;
    n2498_o2 <= 1'b0;
    n2495_o2 <= 1'b0;
    n2496_o2 <= 1'b0;
    n2458_o2 <= 1'b0;
    n2643_o2 <= 1'b0;
    n2462_o2 <= 1'b0;
    n2468_o2 <= 1'b0;
    n2639_o2 <= 1'b0;
    n2499_o2 <= 1'b0;
    n2472_o2 <= 1'b0;
    n2474_o2 <= 1'b0;
    n2489_o2 <= 1'b0;
    n2321_o2 <= 1'b0;
    n2322_o2 <= 1'b0;
    n2640_o2 <= 1'b0;
    n2642_o2 <= 1'b0;
    n2187_o2 <= 1'b0;
    n2373_o2 <= 1'b0;
    n2603_o2 <= 1'b0;
    n2388_o2 <= 1'b0;
    n2437_o2 <= 1'b0;
    n2356_o2 <= 1'b0;
    n2452_o2 <= 1'b0;
    n2347_o2 <= 1'b0;
    n2329_o2 <= 1'b0;
    n2669_o2 <= 1'b0;
    n2332_o2 <= 1'b0;
    n2664_o2 <= 1'b0;
    n2665_o2 <= 1'b0;
    n2653_o2 <= 1'b0;
    n2654_o2 <= 1'b0;
    n2636_o2 <= 1'b0;
    n2660_o2 <= 1'b0;
    n2318_o2 <= 1'b0;
    n2319_o2 <= 1'b0;
    n2586_o2 <= 1'b0;
    n2587_o2 <= 1'b0;
    n2288_o2 <= 1'b0;
    n2344_o2 <= 1'b0;
    n2530_o2 <= 1'b0;
    n2303_o2 <= 1'b0;
    n2566_o2 <= 1'b0;
    n2567_o2 <= 1'b0;
    n2554_o2 <= 1'b0;
    n2194_o2 <= 1'b0;
    lo582_buf_o2 <= 1'b0;
    lo030_buf_o2 <= 1'b0;
    lo174_buf_o2 <= 1'b0;
    lo178_buf_o2 <= 1'b0;
    lo186_buf_o2 <= 1'b0;
    lo266_buf_o2 <= 1'b0;
    lo306_buf_o2 <= 1'b0;
    lo346_buf_o2 <= 1'b0;
    lo386_buf_o2 <= 1'b0;
    lo426_buf_o2 <= 1'b0;
    lo590_buf_o2 <= 1'b0;
    lo594_buf_o2 <= 1'b0;
    lo606_buf_o2 <= 1'b0;
    lo610_buf_o2 <= 1'b0;
    n2238_o2 <= 1'b0;
    n2229_o2 <= 1'b0;
    n2242_o2 <= 1'b0;
    n2233_o2 <= 1'b0;
    n2168_o2 <= 1'b0;
    n2237_o2 <= 1'b0;
    n2228_o2 <= 1'b0;
    n2172_o2 <= 1'b0;
    n2223_o2 <= 1'b0;
    n2222_o2 <= 1'b0;
    n2170_o2 <= 1'b0;
    n2181_o2 <= 1'b0;
    n2510_o2 <= 1'b0;
    n2621_o2 <= 1'b0;
    lo466_buf_o2 <= 1'b0;
    lo478_buf_o2 <= 1'b0;
    n2149_o2 <= 1'b0;
    n2429_o2 <= 1'b0;
    n2444_o2 <= 1'b0;
    n2153_o2 <= 1'b0;
    n2433_o2 <= 1'b0;
    n2448_o2 <= 1'b0;
    n2367_o2 <= 1'b0;
    n2386_o2 <= 1'b0;
    n2539_o2 <= 1'b0;
    n2183_o2 <= 1'b0;
    n2220_o2 <= 1'b0;
    n2514_o2 <= 1'b0;
    n2196_o2 <= 1'b0;
    n2616_o2 <= 1'b0;
    n2612_o2 <= 1'b0;
    n2627_o2 <= 1'b0;
    n2140_o2 <= 1'b0;
    n1877_inv <= 1'b0;
    lo149_buf_o2 <= 1'b0;
    lo197_buf_o2 <= 1'b0;
    lo118_buf_o2 <= 1'b0;
    lo158_buf_o2 <= 1'b0;
    lo166_buf_o2 <= 1'b0;
    lo242_buf_o2 <= 1'b0;
    lo286_buf_o2 <= 1'b0;
    lo506_buf_o2 <= 1'b0;
    n2198_o2 <= 1'b0;
    n2202_o2 <= 1'b0;
    n2197_o2 <= 1'b0;
    n1913_inv <= 1'b0;
    n2146_o2 <= 1'b0;
    n1919_inv <= 1'b0;
    lo312_buf_o2 <= 1'b0;
    lo316_buf_o2 <= 1'b0;
    lo352_buf_o2 <= 1'b0;
    lo356_buf_o2 <= 1'b0;
    lo392_buf_o2 <= 1'b0;
    lo396_buf_o2 <= 1'b0;
    lo432_buf_o2 <= 1'b0;
    lo436_buf_o2 <= 1'b0;
    lo576_buf_o2 <= 1'b0;
  end
endmodule


