// Benchmark "mymod" written by ABC on Wed Nov  1 23:37:36 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36,
    G426, G427, G428, G429, G430, G431, G432  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36;
  output G426, G427, G428, G429, G430, G431, G432;
  reg n229_lo, n253_lo, n256_lo, n259_lo, n262_lo, n277_lo, n301_lo,
    n304_lo, n307_lo, n310_lo, n325_lo, n349_lo, n352_lo, n355_lo, n358_lo,
    n373_lo, n397_lo, n400_lo, n403_lo, n406_lo, n421_lo, n445_lo, n448_lo,
    n451_lo, n454_lo, n469_lo, n493_lo, n496_lo, n499_lo, n502_lo, n517_lo,
    n520_lo, n541_lo, n544_lo, n547_lo, n550_lo, n565_lo, n589_lo, n592_lo,
    n595_lo, n598_lo, n613_lo, n625_lo, n628_lo, n631_lo, n634_lo, n852_o2,
    n853_o2, n955_o2, n956_o2, n531_o2, n549_o2, n537_o2, n540_o2, n546_o2,
    n534_o2, n552_o2, n543_o2, n961_o2, n223_inv, n555_o2, n1009_o2,
    n1010_o2, n1011_o2, n1012_o2, lo026_buf_o2, lo074_buf_o2, lo090_buf_o2,
    lo122_buf_o2, n510_o2, n498_o2, n516_o2, n507_o2, lo106_buf_o2,
    n519_o2, n1029_o2, n1041_o2, n1043_o2, n1045_o2, n558_o2, n563_o2,
    lo094_buf_o2, lo102_buf_o2, n522_o2, n298_inv, n486_o2, n304_inv,
    n564_o2, n528_o2, n492_o2, n530_o2, n548_o2, n536_o2, n539_o2,
    lo025_buf_o2, lo073_buf_o2, lo089_buf_o2, lo121_buf_o2, n509_o2,
    n513_o2, n501_o2, n504_o2, n495_o2, n497_o2, n515_o2, n506_o2,
    lo010_buf_o2, lo042_buf_o2, lo058_buf_o2, lo138_buf_o2, lo014_buf_o2,
    lo022_buf_o2, lo030_buf_o2, lo038_buf_o2, lo046_buf_o2, lo054_buf_o2,
    lo126_buf_o2, lo134_buf_o2, lo093_buf_o2, lo101_buf_o2, lo002_buf_o2,
    lo006_buf_o2, lo062_buf_o2, lo070_buf_o2, lo078_buf_o2, lo086_buf_o2,
    lo110_buf_o2, lo118_buf_o2, n476_o2, n482_o2, n478_o2, n479_o2;
  wire new_new_n308__, new_new_n310__, new_new_n312__, new_new_n314__,
    new_new_n315__, new_new_n316__, new_new_n318__, new_new_n320__,
    new_new_n322__, new_new_n323__, new_new_n324__, new_new_n326__,
    new_new_n328__, new_new_n330__, new_new_n331__, new_new_n332__,
    new_new_n334__, new_new_n336__, new_new_n338__, new_new_n340__,
    new_new_n342__, new_new_n344__, new_new_n346__, new_new_n348__,
    new_new_n350__, new_new_n352__, new_new_n354__, new_new_n356__,
    new_new_n358__, new_new_n360__, new_new_n362__, new_new_n364__,
    new_new_n366__, new_new_n368__, new_new_n370__, new_new_n371__,
    new_new_n372__, new_new_n374__, new_new_n376__, new_new_n378__,
    new_new_n380__, new_new_n382__, new_new_n384__, new_new_n386__,
    new_new_n389__, new_new_n390__, new_new_n392__, new_new_n394__,
    new_new_n396__, new_new_n398__, new_new_n400__, new_new_n402__,
    new_new_n404__, new_new_n406__, new_new_n408__, new_new_n409__,
    new_new_n410__, new_new_n412__, new_new_n414__, new_new_n416__,
    new_new_n418__, new_new_n419__, new_new_n420__, new_new_n422__,
    new_new_n424__, new_new_n426__, new_new_n428__, new_new_n429__,
    new_new_n430__, new_new_n432__, new_new_n434__, new_new_n436__,
    new_new_n438__, new_new_n440__, new_new_n442__, new_new_n444__,
    new_new_n446__, new_new_n448__, new_new_n450__, new_new_n451__,
    new_new_n452__, new_new_n454__, new_new_n456__, new_new_n458__,
    new_new_n460__, new_new_n462__, new_new_n464__, new_new_n466__,
    new_new_n468__, new_new_n470__, new_new_n472__, new_new_n474__,
    new_new_n476__, new_new_n478__, new_new_n480__, new_new_n482__,
    new_new_n483__, new_new_n484__, new_new_n485__, new_new_n487__,
    new_new_n489__, new_new_n490__, new_new_n491__, new_new_n493__,
    new_new_n495__, new_new_n496__, new_new_n498__, new_new_n500__,
    new_new_n501__, new_new_n503__, new_new_n505__, new_new_n507__,
    new_new_n509__, new_new_n510__, new_new_n512__, new_new_n514__,
    new_new_n516__, new_new_n519__, new_new_n521__, new_new_n523__,
    new_new_n525__, new_new_n526__, new_new_n529__, new_new_n531__,
    new_new_n533__, new_new_n535__, new_new_n537__, new_new_n538__,
    new_new_n540__, new_new_n542__, new_new_n545__, new_new_n546__,
    new_new_n548__, new_new_n550__, new_new_n552__, new_new_n554__,
    new_new_n555__, new_new_n556__, new_new_n558__, new_new_n560__,
    new_new_n562__, new_new_n564__, new_new_n566__, new_new_n568__,
    new_new_n570__, new_new_n572__, new_new_n574__, new_new_n576__,
    new_new_n578__, new_new_n579__, new_new_n580__, new_new_n581__,
    new_new_n582__, new_new_n583__, new_new_n584__, new_new_n585__,
    new_new_n586__, new_new_n588__, new_new_n590__, new_new_n592__,
    new_new_n593__, new_new_n594__, new_new_n595__, new_new_n596__,
    new_new_n597__, new_new_n598__, new_new_n599__, new_new_n600__,
    new_new_n602__, new_new_n604__, new_new_n607__, new_new_n608__,
    new_new_n611__, new_new_n612__, new_new_n615__, new_new_n616__,
    new_new_n617__, new_new_n618__, new_new_n620__, new_new_n621__,
    new_new_n622__, new_new_n623__, new_new_n624__, new_new_n625__,
    new_new_n626__, new_new_n628__, new_new_n629__, new_new_n630__,
    new_new_n632__, new_new_n633__, new_new_n634__, new_new_n636__,
    new_new_n638__, new_new_n640__, new_new_n642__, new_new_n644__,
    new_new_n645__, new_new_n646__, new_new_n647__, new_new_n648__,
    new_new_n649__, new_new_n650__, new_new_n651__, new_new_n652__,
    new_new_n653__, new_new_n654__, new_new_n655__, new_new_n656__,
    new_new_n657__, new_new_n658__, new_new_n659__, new_new_n660__,
    new_new_n661__, new_new_n662__, new_new_n663__, new_new_n664__,
    new_new_n665__, new_new_n666__, new_new_n667__, new_new_n668__,
    new_new_n669__, new_new_n670__, new_new_n671__, new_new_n672__,
    new_new_n673__, new_new_n674__, new_new_n675__, new_new_n676__,
    new_new_n677__, new_new_n678__, new_new_n679__, new_new_n680__,
    new_new_n681__, new_new_n682__, new_new_n683__, new_new_n684__,
    new_new_n685__, new_new_n686__, new_new_n687__, new_new_n688__,
    new_new_n689__, new_new_n690__, new_new_n691__, new_new_n692__,
    new_new_n693__, new_new_n694__, new_new_n695__, new_new_n696__,
    new_new_n697__, new_new_n698__, new_new_n699__, new_new_n700__,
    new_new_n701__, new_new_n702__, new_new_n703__, new_new_n704__,
    new_new_n705__, new_new_n706__, new_new_n707__, new_new_n708__,
    new_new_n709__, new_new_n710__, new_new_n711__, new_new_n712__,
    new_new_n713__, new_new_n714__, new_new_n715__, new_new_n716__,
    new_new_n717__, new_new_n718__, new_new_n719__, new_new_n720__,
    new_new_n721__, new_new_n722__, new_new_n723__, new_new_n724__,
    new_new_n725__, new_new_n726__, new_new_n727__, new_new_n728__,
    new_new_n729__, new_new_n730__, new_new_n731__, new_new_n732__,
    new_new_n733__, new_new_n734__, new_new_n735__, new_new_n736__,
    new_new_n737__, new_new_n738__, new_new_n739__, new_new_n740__,
    new_new_n741__, new_new_n742__, new_new_n743__, new_new_n744__,
    new_new_n745__, new_new_n746__, new_new_n747__, new_new_n748__,
    new_new_n749__, new_new_n750__, new_new_n751__, new_new_n752__,
    new_new_n753__, new_new_n754__, new_new_n755__, new_new_n756__,
    new_new_n757__, new_new_n758__, new_new_n759__, new_new_n760__,
    new_new_n761__, new_new_n762__, new_new_n763__, new_new_n764__,
    new_new_n765__, new_new_n766__, new_new_n767__, new_new_n768__,
    new_new_n769__, new_new_n770__, new_new_n771__, new_new_n772__,
    new_new_n773__, new_new_n774__, new_new_n775__, new_new_n776__,
    new_new_n777__, new_new_n778__, new_new_n779__, new_new_n919__,
    new_new_n920__, new_new_n921__, new_new_n922__, new_new_n923__,
    new_new_n924__, new_new_n925__, new_new_n926__, new_new_n927__,
    new_new_n928__, new_new_n929__, new_new_n930__, new_new_n931__,
    new_new_n932__, new_new_n933__, new_new_n934__, new_new_n935__,
    new_new_n936__, new_new_n937__, new_new_n938__, new_new_n939__,
    new_new_n940__, new_new_n941__, new_new_n942__, new_new_n943__,
    new_new_n944__, new_new_n945__, new_new_n946__, new_new_n947__,
    new_new_n948__, new_new_n949__, new_new_n950__, new_new_n951__,
    new_new_n952__, new_new_n953__, new_new_n954__, new_new_n955__,
    new_new_n956__, new_new_n957__, new_new_n958__, new_new_n959__,
    new_new_n960__, new_new_n961__, new_new_n962__, new_new_n963__,
    new_new_n964__, new_new_n965__, new_new_n966__, new_new_n967__,
    new_new_n968__, new_new_n969__, new_new_n970__, new_new_n971__,
    new_new_n972__, new_new_n973__, new_new_n974__, new_new_n975__,
    new_new_n976__, new_new_n977__, new_new_n978__, new_new_n979__,
    new_new_n980__, new_new_n981__, new_new_n982__, new_new_n983__,
    new_new_n984__, new_new_n985__, new_new_n986__, new_new_n987__,
    new_new_n988__, new_new_n989__, new_new_n990__, new_new_n991__,
    new_new_n992__, new_new_n993__, new_new_n994__, new_new_n995__,
    new_new_n996__, new_new_n997__, new_new_n998__, n1312, n1315, n1318,
    n1321, n1324, n1327, n1330, n1333, n1336, n1339, n1342, n1345, n1348,
    n1351, n1354, n1357, n1360, n1363, n1366, n1369, n1372, n1375, n1378,
    n1381, n1384, n1387, n1390, n1393, n1396, n1399, n1402, n1405, n1408,
    n1411, n1414, n1417, n1420, n1423, n1426, n1429, n1432, n1435, n1438,
    n1441, n1444, n1447, n1450, n1453, n1456, n1459, n1462, n1465, n1468,
    n1471, n1474, n1477, n1480, n1483, n1486, n1489, n1492, n1495, n1498,
    n1501, n1504, n1507, n1510, n1513, n1516, n1519, n1522, n1525, n1528,
    n1531, n1534, n1537, n1540, n1543, n1546, n1549, n1552, n1555, n1558,
    n1561, n1564, n1567, n1570, n1573, n1576, n1579, n1582, n1585, n1588,
    n1591, n1594, n1597, n1600, n1603, n1606, n1609, n1612, n1615, n1618,
    n1621, n1624, n1627, n1630, n1633, n1636, n1639, n1642, n1645, n1648,
    n1651, n1654, n1657, n1660, n1663, n1666, n1669, n1672, n1675, n1678,
    n1681, n1684, n1687, n1690, n1693, n1696, n1699, n1702, n1705;
  buf1  g000(.din(G1), .dout(new_new_n308__));
  buf1  g001(.din(G2), .dout(new_new_n310__));
  buf1  g002(.din(G3), .dout(new_new_n312__));
  buf1  g003(.din(G4), .dout(new_new_n314__));
  not1  g004(.din(G4), .dout(new_new_n315__));
  buf1  g005(.din(G5), .dout(new_new_n316__));
  buf1  g006(.din(G6), .dout(new_new_n318__));
  buf1  g007(.din(G7), .dout(new_new_n320__));
  buf1  g008(.din(G8), .dout(new_new_n322__));
  not1  g009(.din(G8), .dout(new_new_n323__));
  buf1  g010(.din(G9), .dout(new_new_n324__));
  buf1  g011(.din(G10), .dout(new_new_n326__));
  buf1  g012(.din(G11), .dout(new_new_n328__));
  buf1  g013(.din(G12), .dout(new_new_n330__));
  not1  g014(.din(G12), .dout(new_new_n331__));
  buf1  g015(.din(G13), .dout(new_new_n332__));
  buf1  g016(.din(G14), .dout(new_new_n334__));
  buf1  g017(.din(G15), .dout(new_new_n336__));
  buf1  g018(.din(G16), .dout(new_new_n338__));
  buf1  g019(.din(G17), .dout(new_new_n340__));
  buf1  g020(.din(G18), .dout(new_new_n342__));
  buf1  g021(.din(G19), .dout(new_new_n344__));
  buf1  g022(.din(G20), .dout(new_new_n346__));
  buf1  g023(.din(G21), .dout(new_new_n348__));
  buf1  g024(.din(G22), .dout(new_new_n350__));
  buf1  g025(.din(G23), .dout(new_new_n352__));
  buf1  g026(.din(G24), .dout(new_new_n354__));
  buf1  g027(.din(G25), .dout(new_new_n356__));
  buf1  g028(.din(G26), .dout(new_new_n358__));
  buf1  g029(.din(G27), .dout(new_new_n360__));
  buf1  g030(.din(G28), .dout(new_new_n362__));
  buf1  g031(.din(G29), .dout(new_new_n364__));
  buf1  g032(.din(G30), .dout(new_new_n366__));
  buf1  g033(.din(G31), .dout(new_new_n368__));
  buf1  g034(.din(G32), .dout(new_new_n370__));
  not1  g035(.din(G32), .dout(new_new_n371__));
  buf1  g036(.din(G33), .dout(new_new_n372__));
  buf1  g037(.din(G34), .dout(new_new_n374__));
  buf1  g038(.din(G35), .dout(new_new_n376__));
  buf1  g039(.din(G36), .dout(new_new_n378__));
  buf1  g040(.din(n229_lo), .dout(new_new_n380__));
  buf1  g041(.din(n253_lo), .dout(new_new_n382__));
  buf1  g042(.din(n256_lo), .dout(new_new_n384__));
  buf1  g043(.din(n259_lo), .dout(new_new_n386__));
  not1  g044(.din(n262_lo), .dout(new_new_n389__));
  buf1  g045(.din(n277_lo), .dout(new_new_n390__));
  buf1  g046(.din(n301_lo), .dout(new_new_n392__));
  buf1  g047(.din(n304_lo), .dout(new_new_n394__));
  buf1  g048(.din(n307_lo), .dout(new_new_n396__));
  buf1  g049(.din(n310_lo), .dout(new_new_n398__));
  buf1  g050(.din(n325_lo), .dout(new_new_n400__));
  buf1  g051(.din(n349_lo), .dout(new_new_n402__));
  buf1  g052(.din(n352_lo), .dout(new_new_n404__));
  buf1  g053(.din(n355_lo), .dout(new_new_n406__));
  buf1  g054(.din(n358_lo), .dout(new_new_n408__));
  not1  g055(.din(n358_lo), .dout(new_new_n409__));
  buf1  g056(.din(n373_lo), .dout(new_new_n410__));
  buf1  g057(.din(n397_lo), .dout(new_new_n412__));
  buf1  g058(.din(n400_lo), .dout(new_new_n414__));
  buf1  g059(.din(n403_lo), .dout(new_new_n416__));
  buf1  g060(.din(n406_lo), .dout(new_new_n418__));
  not1  g061(.din(n406_lo), .dout(new_new_n419__));
  buf1  g062(.din(n421_lo), .dout(new_new_n420__));
  buf1  g063(.din(n445_lo), .dout(new_new_n422__));
  buf1  g064(.din(n448_lo), .dout(new_new_n424__));
  buf1  g065(.din(n451_lo), .dout(new_new_n426__));
  buf1  g066(.din(n454_lo), .dout(new_new_n428__));
  not1  g067(.din(n454_lo), .dout(new_new_n429__));
  buf1  g068(.din(n469_lo), .dout(new_new_n430__));
  buf1  g069(.din(n493_lo), .dout(new_new_n432__));
  buf1  g070(.din(n496_lo), .dout(new_new_n434__));
  buf1  g071(.din(n499_lo), .dout(new_new_n436__));
  buf1  g072(.din(n502_lo), .dout(new_new_n438__));
  buf1  g073(.din(n517_lo), .dout(new_new_n440__));
  buf1  g074(.din(n520_lo), .dout(new_new_n442__));
  buf1  g075(.din(n541_lo), .dout(new_new_n444__));
  buf1  g076(.din(n544_lo), .dout(new_new_n446__));
  buf1  g077(.din(n547_lo), .dout(new_new_n448__));
  buf1  g078(.din(n550_lo), .dout(new_new_n450__));
  not1  g079(.din(n550_lo), .dout(new_new_n451__));
  buf1  g080(.din(n565_lo), .dout(new_new_n452__));
  buf1  g081(.din(n589_lo), .dout(new_new_n454__));
  buf1  g082(.din(n592_lo), .dout(new_new_n456__));
  buf1  g083(.din(n595_lo), .dout(new_new_n458__));
  buf1  g084(.din(n598_lo), .dout(new_new_n460__));
  buf1  g085(.din(n613_lo), .dout(new_new_n462__));
  buf1  g086(.din(n625_lo), .dout(new_new_n464__));
  buf1  g087(.din(n628_lo), .dout(new_new_n466__));
  buf1  g088(.din(n631_lo), .dout(new_new_n468__));
  buf1  g089(.din(n634_lo), .dout(new_new_n470__));
  buf1  g090(.din(n852_o2), .dout(new_new_n472__));
  buf1  g091(.din(n853_o2), .dout(new_new_n474__));
  buf1  g092(.din(n955_o2), .dout(new_new_n476__));
  buf1  g093(.din(n956_o2), .dout(new_new_n478__));
  buf1  g094(.din(n531_o2), .dout(new_new_n480__));
  buf1  g095(.din(n549_o2), .dout(new_new_n482__));
  not1  g096(.din(n549_o2), .dout(new_new_n483__));
  buf1  g097(.din(n537_o2), .dout(new_new_n484__));
  not1  g098(.din(n537_o2), .dout(new_new_n485__));
  not1  g099(.din(n540_o2), .dout(new_new_n487__));
  not1  g100(.din(n546_o2), .dout(new_new_n489__));
  buf1  g101(.din(n534_o2), .dout(new_new_n490__));
  not1  g102(.din(n534_o2), .dout(new_new_n491__));
  not1  g103(.din(n552_o2), .dout(new_new_n493__));
  not1  g104(.din(n543_o2), .dout(new_new_n495__));
  buf1  g105(.din(n961_o2), .dout(new_new_n496__));
  buf1  g106(.din(n223_inv), .dout(new_new_n498__));
  buf1  g107(.din(n555_o2), .dout(new_new_n500__));
  not1  g108(.din(n555_o2), .dout(new_new_n501__));
  not1  g109(.din(n1009_o2), .dout(new_new_n503__));
  not1  g110(.din(n1010_o2), .dout(new_new_n505__));
  not1  g111(.din(n1011_o2), .dout(new_new_n507__));
  not1  g112(.din(n1012_o2), .dout(new_new_n509__));
  buf1  g113(.din(lo026_buf_o2), .dout(new_new_n510__));
  buf1  g114(.din(lo074_buf_o2), .dout(new_new_n512__));
  buf1  g115(.din(lo090_buf_o2), .dout(new_new_n514__));
  buf1  g116(.din(lo122_buf_o2), .dout(new_new_n516__));
  not1  g117(.din(n510_o2), .dout(new_new_n519__));
  not1  g118(.din(n498_o2), .dout(new_new_n521__));
  not1  g119(.din(n516_o2), .dout(new_new_n523__));
  not1  g120(.din(n507_o2), .dout(new_new_n525__));
  buf1  g121(.din(lo106_buf_o2), .dout(new_new_n526__));
  not1  g122(.din(n519_o2), .dout(new_new_n529__));
  not1  g123(.din(n1029_o2), .dout(new_new_n531__));
  not1  g124(.din(n1041_o2), .dout(new_new_n533__));
  not1  g125(.din(n1043_o2), .dout(new_new_n535__));
  not1  g126(.din(n1045_o2), .dout(new_new_n537__));
  buf1  g127(.din(n558_o2), .dout(new_new_n538__));
  buf1  g128(.din(n563_o2), .dout(new_new_n540__));
  buf1  g129(.din(lo094_buf_o2), .dout(new_new_n542__));
  not1  g130(.din(lo102_buf_o2), .dout(new_new_n545__));
  buf1  g131(.din(n522_o2), .dout(new_new_n546__));
  buf1  g132(.din(n298_inv), .dout(new_new_n548__));
  buf1  g133(.din(n486_o2), .dout(new_new_n550__));
  buf1  g134(.din(n304_inv), .dout(new_new_n552__));
  buf1  g135(.din(n564_o2), .dout(new_new_n554__));
  not1  g136(.din(n564_o2), .dout(new_new_n555__));
  buf1  g137(.din(n528_o2), .dout(new_new_n556__));
  buf1  g138(.din(n492_o2), .dout(new_new_n558__));
  buf1  g139(.din(n530_o2), .dout(new_new_n560__));
  buf1  g140(.din(n548_o2), .dout(new_new_n562__));
  buf1  g141(.din(n536_o2), .dout(new_new_n564__));
  buf1  g142(.din(n539_o2), .dout(new_new_n566__));
  buf1  g143(.din(lo025_buf_o2), .dout(new_new_n568__));
  buf1  g144(.din(lo073_buf_o2), .dout(new_new_n570__));
  buf1  g145(.din(lo089_buf_o2), .dout(new_new_n572__));
  buf1  g146(.din(lo121_buf_o2), .dout(new_new_n574__));
  buf1  g147(.din(n509_o2), .dout(new_new_n576__));
  buf1  g148(.din(n513_o2), .dout(new_new_n578__));
  not1  g149(.din(n513_o2), .dout(new_new_n579__));
  buf1  g150(.din(n501_o2), .dout(new_new_n580__));
  not1  g151(.din(n501_o2), .dout(new_new_n581__));
  buf1  g152(.din(n504_o2), .dout(new_new_n582__));
  not1  g153(.din(n504_o2), .dout(new_new_n583__));
  buf1  g154(.din(n495_o2), .dout(new_new_n584__));
  not1  g155(.din(n495_o2), .dout(new_new_n585__));
  buf1  g156(.din(n497_o2), .dout(new_new_n586__));
  buf1  g157(.din(n515_o2), .dout(new_new_n588__));
  buf1  g158(.din(n506_o2), .dout(new_new_n590__));
  buf1  g159(.din(lo010_buf_o2), .dout(new_new_n592__));
  not1  g160(.din(lo010_buf_o2), .dout(new_new_n593__));
  buf1  g161(.din(lo042_buf_o2), .dout(new_new_n594__));
  not1  g162(.din(lo042_buf_o2), .dout(new_new_n595__));
  buf1  g163(.din(lo058_buf_o2), .dout(new_new_n596__));
  not1  g164(.din(lo058_buf_o2), .dout(new_new_n597__));
  buf1  g165(.din(lo138_buf_o2), .dout(new_new_n598__));
  not1  g166(.din(lo138_buf_o2), .dout(new_new_n599__));
  buf1  g167(.din(lo014_buf_o2), .dout(new_new_n600__));
  buf1  g168(.din(lo022_buf_o2), .dout(new_new_n602__));
  buf1  g169(.din(lo030_buf_o2), .dout(new_new_n604__));
  not1  g170(.din(lo038_buf_o2), .dout(new_new_n607__));
  buf1  g171(.din(lo046_buf_o2), .dout(new_new_n608__));
  not1  g172(.din(lo054_buf_o2), .dout(new_new_n611__));
  buf1  g173(.din(lo126_buf_o2), .dout(new_new_n612__));
  not1  g174(.din(lo134_buf_o2), .dout(new_new_n615__));
  buf1  g175(.din(lo093_buf_o2), .dout(new_new_n616__));
  not1  g176(.din(lo093_buf_o2), .dout(new_new_n617__));
  buf1  g177(.din(lo101_buf_o2), .dout(new_new_n618__));
  buf1  g178(.din(lo002_buf_o2), .dout(new_new_n620__));
  not1  g179(.din(lo002_buf_o2), .dout(new_new_n621__));
  buf1  g180(.din(lo006_buf_o2), .dout(new_new_n622__));
  not1  g181(.din(lo006_buf_o2), .dout(new_new_n623__));
  buf1  g182(.din(lo062_buf_o2), .dout(new_new_n624__));
  not1  g183(.din(lo062_buf_o2), .dout(new_new_n625__));
  buf1  g184(.din(lo070_buf_o2), .dout(new_new_n626__));
  buf1  g185(.din(lo078_buf_o2), .dout(new_new_n628__));
  not1  g186(.din(lo078_buf_o2), .dout(new_new_n629__));
  buf1  g187(.din(lo086_buf_o2), .dout(new_new_n630__));
  buf1  g188(.din(lo110_buf_o2), .dout(new_new_n632__));
  not1  g189(.din(lo110_buf_o2), .dout(new_new_n633__));
  buf1  g190(.din(lo118_buf_o2), .dout(new_new_n634__));
  buf1  g191(.din(n476_o2), .dout(new_new_n636__));
  buf1  g192(.din(n482_o2), .dout(new_new_n638__));
  buf1  g193(.din(n478_o2), .dout(new_new_n640__));
  buf1  g194(.din(n479_o2), .dout(new_new_n642__));
  or1   g195(.dina(new_new_n472__), .dinb(new_new_n474__), .dout(new_new_n644__));
  or1   g196(.dina(new_new_n476__), .dinb(new_new_n478__), .dout(new_new_n645__));
  or1   g197(.dina(new_new_n538__), .dinb(new_new_n540__), .dout(new_new_n646__));
  or1   g198(.dina(new_new_n389__), .dinb(new_new_n921__), .dout(new_new_n647__));
  and1  g199(.dina(new_new_n480__), .dinb(new_new_n647__), .dout(new_new_n648__));
  and1  g200(.dina(new_new_n460__), .dinb(new_new_n925__), .dout(new_new_n649__));
  or1   g201(.dina(new_new_n495__), .dinb(new_new_n649__), .dout(new_new_n650__));
  and1  g202(.dina(new_new_n450__), .dinb(new_new_n925__), .dout(new_new_n651__));
  or1   g203(.dina(new_new_n451__), .dinb(new_new_n921__), .dout(new_new_n652__));
  and1  g204(.dina(new_new_n500__), .dinb(new_new_n652__), .dout(new_new_n653__));
  or1   g205(.dina(new_new_n501__), .dinb(new_new_n651__), .dout(new_new_n654__));
  and1  g206(.dina(new_new_n930__), .dinb(new_new_n931__), .dout(new_new_n655__));
  and1  g207(.dina(new_new_n438__), .dinb(new_new_n926__), .dout(new_new_n656__));
  or1   g208(.dina(new_new_n493__), .dinb(new_new_n656__), .dout(new_new_n657__));
  and1  g209(.dina(new_new_n470__), .dinb(new_new_n926__), .dout(new_new_n658__));
  or1   g210(.dina(new_new_n487__), .dinb(new_new_n658__), .dout(new_new_n659__));
  and1  g211(.dina(new_new_n932__), .dinb(new_new_n659__), .dout(new_new_n660__));
  and1  g212(.dina(new_new_n655__), .dinb(new_new_n660__), .dout(new_new_n661__));
  and1  g213(.dina(new_new_n408__), .dinb(new_new_n928__), .dout(new_new_n662__));
  or1   g214(.dina(new_new_n409__), .dinb(new_new_n920__), .dout(new_new_n663__));
  and1  g215(.dina(new_new_n482__), .dinb(new_new_n663__), .dout(new_new_n664__));
  or1   g216(.dina(new_new_n483__), .dinb(new_new_n662__), .dout(new_new_n665__));
  and1  g217(.dina(new_new_n428__), .dinb(new_new_n928__), .dout(new_new_n666__));
  or1   g218(.dina(new_new_n429__), .dinb(new_new_n922__), .dout(new_new_n667__));
  and1  g219(.dina(new_new_n490__), .dinb(new_new_n667__), .dout(new_new_n668__));
  or1   g220(.dina(new_new_n491__), .dinb(new_new_n666__), .dout(new_new_n669__));
  and1  g221(.dina(new_new_n933__), .dinb(new_new_n669__), .dout(new_new_n670__));
  or1   g222(.dina(new_new_n934__), .dinb(new_new_n935__), .dout(new_new_n671__));
  and1  g223(.dina(new_new_n398__), .dinb(new_new_n929__), .dout(new_new_n672__));
  or1   g224(.dina(new_new_n489__), .dinb(new_new_n672__), .dout(new_new_n673__));
  and1  g225(.dina(new_new_n418__), .dinb(new_new_n929__), .dout(new_new_n674__));
  or1   g226(.dina(new_new_n419__), .dinb(new_new_n922__), .dout(new_new_n675__));
  and1  g227(.dina(new_new_n484__), .dinb(new_new_n675__), .dout(new_new_n676__));
  or1   g228(.dina(new_new_n485__), .dinb(new_new_n674__), .dout(new_new_n677__));
  and1  g229(.dina(new_new_n936__), .dinb(new_new_n937__), .dout(new_new_n678__));
  and1  g230(.dina(new_new_n670__), .dinb(new_new_n678__), .dout(new_new_n679__));
  and1  g231(.dina(new_new_n661__), .dinb(new_new_n938__), .dout(new_new_n680__));
  or1   g232(.dina(new_new_n648__), .dinb(new_new_n680__), .dout(new_new_n681__));
  or1   g233(.dina(new_new_n932__), .dinb(new_new_n939__), .dout(new_new_n682__));
  or1   g234(.dina(new_new_n671__), .dinb(new_new_n682__), .dout(new_new_n683__));
  and1  g235(.dina(new_new_n936__), .dinb(new_new_n683__), .dout(new_new_n684__));
  or1   g236(.dina(new_new_n935__), .dinb(new_new_n939__), .dout(new_new_n685__));
  or1   g237(.dina(new_new_n931__), .dinb(new_new_n685__), .dout(new_new_n686__));
  and1  g238(.dina(new_new_n933__), .dinb(new_new_n686__), .dout(new_new_n687__));
  and1  g239(.dina(new_new_n940__), .dinb(new_new_n687__), .dout(new_new_n688__));
  or1   g240(.dina(new_new_n930__), .dinb(new_new_n653__), .dout(new_new_n689__));
  and1  g241(.dina(new_new_n937__), .dinb(new_new_n689__), .dout(new_new_n690__));
  or1   g242(.dina(new_new_n934__), .dinb(new_new_n690__), .dout(new_new_n691__));
  and1  g243(.dina(new_new_n940__), .dinb(new_new_n691__), .dout(new_new_n692__));
  or1   g244(.dina(new_new_n509__), .dinb(new_new_n560__), .dout(new_new_n693__));
  or1   g245(.dina(new_new_n503__), .dinb(new_new_n562__), .dout(new_new_n694__));
  or1   g246(.dina(new_new_n505__), .dinb(new_new_n564__), .dout(new_new_n695__));
  or1   g247(.dina(new_new_n507__), .dinb(new_new_n566__), .dout(new_new_n696__));
  and1  g248(.dina(new_new_n510__), .dinb(new_new_n943__), .dout(new_new_n697__));
  or1   g249(.dina(new_new_n519__), .dinb(new_new_n697__), .dout(new_new_n698__));
  and1  g250(.dina(new_new_n512__), .dinb(new_new_n943__), .dout(new_new_n699__));
  or1   g251(.dina(new_new_n521__), .dinb(new_new_n699__), .dout(new_new_n700__));
  and1  g252(.dina(new_new_n514__), .dinb(new_new_n942__), .dout(new_new_n701__));
  or1   g253(.dina(new_new_n523__), .dinb(new_new_n701__), .dout(new_new_n702__));
  and1  g254(.dina(new_new_n516__), .dinb(new_new_n944__), .dout(new_new_n703__));
  or1   g255(.dina(new_new_n525__), .dinb(new_new_n703__), .dout(new_new_n704__));
  and1  g256(.dina(new_new_n526__), .dinb(new_new_n944__), .dout(new_new_n705__));
  or1   g257(.dina(new_new_n529__), .dinb(new_new_n705__), .dout(new_new_n706__));
  or1   g258(.dina(new_new_n531__), .dinb(new_new_n576__), .dout(new_new_n707__));
  or1   g259(.dina(new_new_n533__), .dinb(new_new_n586__), .dout(new_new_n708__));
  or1   g260(.dina(new_new_n535__), .dinb(new_new_n588__), .dout(new_new_n709__));
  or1   g261(.dina(new_new_n537__), .dinb(new_new_n590__), .dout(new_new_n710__));
  and1  g262(.dina(new_new_n542__), .dinb(new_new_n558__), .dout(new_new_n711__));
  or1   g263(.dina(new_new_n545__), .dinb(new_new_n711__), .dout(new_new_n712__));
  or1   g264(.dina(new_new_n945__), .dinb(new_new_n946__), .dout(new_new_n713__));
  or1   g265(.dina(new_new_n947__), .dinb(new_new_n948__), .dout(new_new_n714__));
  or1   g266(.dina(new_new_n949__), .dinb(new_new_n950__), .dout(new_new_n715__));
  and1  g267(.dina(new_new_n714__), .dinb(new_new_n715__), .dout(new_new_n716__));
  and1  g268(.dina(new_new_n713__), .dinb(new_new_n716__), .dout(new_new_n717__));
  or1   g269(.dina(new_new_n951__), .dinb(new_new_n952__), .dout(new_new_n718__));
  or1   g270(.dina(new_new_n953__), .dinb(new_new_n954__), .dout(new_new_n719__));
  and1  g271(.dina(new_new_n718__), .dinb(new_new_n719__), .dout(new_new_n720__));
  or1   g272(.dina(new_new_n955__), .dinb(new_new_n956__), .dout(new_new_n721__));
  or1   g273(.dina(new_new_n957__), .dinb(new_new_n958__), .dout(new_new_n722__));
  and1  g274(.dina(new_new_n721__), .dinb(new_new_n722__), .dout(new_new_n723__));
  or1   g275(.dina(new_new_n959__), .dinb(new_new_n960__), .dout(new_new_n724__));
  or1   g276(.dina(new_new_n961__), .dinb(new_new_n962__), .dout(new_new_n725__));
  and1  g277(.dina(new_new_n724__), .dinb(new_new_n725__), .dout(new_new_n726__));
  and1  g278(.dina(new_new_n723__), .dinb(new_new_n726__), .dout(new_new_n727__));
  and1  g279(.dina(new_new_n720__), .dinb(new_new_n727__), .dout(new_new_n728__));
  or1   g280(.dina(new_new_n963__), .dinb(new_new_n964__), .dout(new_new_n729__));
  or1   g281(.dina(new_new_n965__), .dinb(new_new_n966__), .dout(new_new_n730__));
  or1   g282(.dina(new_new_n967__), .dinb(new_new_n968__), .dout(new_new_n731__));
  and1  g283(.dina(new_new_n730__), .dinb(new_new_n731__), .dout(new_new_n732__));
  and1  g284(.dina(new_new_n729__), .dinb(new_new_n732__), .dout(new_new_n733__));
  or1   g285(.dina(new_new_n969__), .dinb(new_new_n970__), .dout(new_new_n734__));
  or1   g286(.dina(new_new_n971__), .dinb(new_new_n972__), .dout(new_new_n735__));
  and1  g287(.dina(new_new_n734__), .dinb(new_new_n735__), .dout(new_new_n736__));
  or1   g288(.dina(new_new_n585__), .dinb(new_new_n592__), .dout(new_new_n737__));
  or1   g289(.dina(new_new_n583__), .dinb(new_new_n598__), .dout(new_new_n738__));
  and1  g290(.dina(new_new_n737__), .dinb(new_new_n738__), .dout(new_new_n739__));
  or1   g291(.dina(new_new_n581__), .dinb(new_new_n596__), .dout(new_new_n740__));
  or1   g292(.dina(new_new_n579__), .dinb(new_new_n594__), .dout(new_new_n741__));
  and1  g293(.dina(new_new_n740__), .dinb(new_new_n741__), .dout(new_new_n742__));
  and1  g294(.dina(new_new_n739__), .dinb(new_new_n742__), .dout(new_new_n743__));
  and1  g295(.dina(new_new_n736__), .dinb(new_new_n743__), .dout(new_new_n744__));
  and1  g296(.dina(new_new_n617__), .dinb(new_new_n973__), .dout(new_new_n745__));
  and1  g297(.dina(new_new_n633__), .dinb(new_new_n974__), .dout(new_new_n746__));
  and1  g298(.dina(new_new_n621__), .dinb(new_new_n622__), .dout(new_new_n747__));
  or1   g299(.dina(new_new_n746__), .dinb(new_new_n747__), .dout(new_new_n748__));
  or1   g300(.dina(new_new_n745__), .dinb(new_new_n748__), .dout(new_new_n749__));
  and1  g301(.dina(new_new_n625__), .dinb(new_new_n975__), .dout(new_new_n750__));
  and1  g302(.dina(new_new_n629__), .dinb(new_new_n976__), .dout(new_new_n751__));
  or1   g303(.dina(new_new_n750__), .dinb(new_new_n751__), .dout(new_new_n752__));
  or1   g304(.dina(new_new_n636__), .dinb(new_new_n642__), .dout(new_new_n753__));
  or1   g305(.dina(new_new_n638__), .dinb(new_new_n640__), .dout(new_new_n754__));
  or1   g306(.dina(new_new_n753__), .dinb(new_new_n754__), .dout(new_new_n755__));
  or1   g307(.dina(new_new_n752__), .dinb(new_new_n755__), .dout(new_new_n756__));
  and1  g308(.dina(new_new_n977__), .dinb(new_new_n978__), .dout(new_new_n757__));
  and1  g309(.dina(new_new_n979__), .dinb(new_new_n980__), .dout(new_new_n758__));
  or1   g310(.dina(new_new_n981__), .dinb(new_new_n982__), .dout(new_new_n759__));
  or1   g311(.dina(new_new_n593__), .dinb(new_new_n985__), .dout(new_new_n760__));
  or1   g312(.dina(new_new_n595__), .dinb(new_new_n985__), .dout(new_new_n761__));
  or1   g313(.dina(new_new_n597__), .dinb(new_new_n984__), .dout(new_new_n762__));
  or1   g314(.dina(new_new_n599__), .dinb(new_new_n986__), .dout(new_new_n763__));
  and1  g315(.dina(new_new_n600__), .dinb(new_new_n990__), .dout(new_new_n764__));
  and1  g316(.dina(new_new_n604__), .dinb(new_new_n990__), .dout(new_new_n765__));
  or1   g317(.dina(new_new_n607__), .dinb(new_new_n765__), .dout(new_new_n766__));
  and1  g318(.dina(new_new_n608__), .dinb(new_new_n989__), .dout(new_new_n767__));
  or1   g319(.dina(new_new_n611__), .dinb(new_new_n767__), .dout(new_new_n768__));
  and1  g320(.dina(new_new_n612__), .dinb(new_new_n991__), .dout(new_new_n769__));
  or1   g321(.dina(new_new_n615__), .dinb(new_new_n769__), .dout(new_new_n770__));
  and1  g322(.dina(new_new_n620__), .dinb(new_new_n991__), .dout(new_new_n771__));
  or1   g323(.dina(new_new_n623__), .dinb(new_new_n771__), .dout(new_new_n772__));
  and1  g324(.dina(new_new_n624__), .dinb(new_new_n993__), .dout(new_new_n773__));
  and1  g325(.dina(new_new_n628__), .dinb(new_new_n993__), .dout(new_new_n774__));
  and1  g326(.dina(new_new_n632__), .dinb(new_new_n994__), .dout(new_new_n775__));
  and1  g327(.dina(new_new_n315__), .dinb(new_new_n995__), .dout(new_new_n776__));
  and1  g328(.dina(new_new_n323__), .dinb(new_new_n996__), .dout(new_new_n777__));
  and1  g329(.dina(new_new_n331__), .dinb(new_new_n997__), .dout(new_new_n778__));
  and1  g330(.dina(new_new_n371__), .dinb(new_new_n998__), .dout(new_new_n779__));
  buf1  g331(.din(new_new_n644__), .dout(G426));
  buf1  g332(.din(new_new_n645__), .dout(G427));
  buf1  g333(.din(new_new_n646__), .dout(G428));
  not1  g334(.din(new_new_n681__), .dout(G429));
  not1  g335(.din(new_new_n938__), .dout(G430));
  not1  g336(.din(new_new_n688__), .dout(G431));
  not1  g337(.din(new_new_n692__), .dout(G432));
  buf1  g338(.din(new_new_n312__), .dout(n1312));
  buf1  g339(.din(new_new_n316__), .dout(n1315));
  buf1  g340(.din(new_new_n382__), .dout(n1318));
  buf1  g341(.din(new_new_n384__), .dout(n1321));
  buf1  g342(.din(new_new_n955__), .dout(n1324));
  buf1  g343(.din(new_new_n320__), .dout(n1327));
  buf1  g344(.din(new_new_n324__), .dout(n1330));
  buf1  g345(.din(new_new_n392__), .dout(n1333));
  buf1  g346(.din(new_new_n394__), .dout(n1336));
  buf1  g347(.din(new_new_n949__), .dout(n1339));
  buf1  g348(.din(new_new_n328__), .dout(n1342));
  buf1  g349(.din(new_new_n332__), .dout(n1345));
  buf1  g350(.din(new_new_n402__), .dout(n1348));
  buf1  g351(.din(new_new_n404__), .dout(n1351));
  buf1  g352(.din(new_new_n961__), .dout(n1354));
  buf1  g353(.din(new_new_n336__), .dout(n1357));
  buf1  g354(.din(new_new_n340__), .dout(n1360));
  buf1  g355(.din(new_new_n412__), .dout(n1363));
  buf1  g356(.din(new_new_n414__), .dout(n1366));
  buf1  g357(.din(new_new_n959__), .dout(n1369));
  buf1  g358(.din(new_new_n344__), .dout(n1372));
  buf1  g359(.din(new_new_n348__), .dout(n1375));
  buf1  g360(.din(new_new_n422__), .dout(n1378));
  buf1  g361(.din(new_new_n424__), .dout(n1381));
  buf1  g362(.din(new_new_n951__), .dout(n1384));
  buf1  g363(.din(new_new_n352__), .dout(n1387));
  buf1  g364(.din(new_new_n356__), .dout(n1390));
  buf1  g365(.din(new_new_n432__), .dout(n1393));
  buf1  g366(.din(new_new_n434__), .dout(n1396));
  buf1  g367(.din(new_new_n953__), .dout(n1399));
  buf1  g368(.din(new_new_n360__), .dout(n1402));
  buf1  g369(.din(new_new_n440__), .dout(n1405));
  buf1  g370(.din(new_new_n364__), .dout(n1408));
  buf1  g371(.din(new_new_n444__), .dout(n1411));
  buf1  g372(.din(new_new_n446__), .dout(n1414));
  buf1  g373(.din(new_new_n945__), .dout(n1417));
  buf1  g374(.din(new_new_n368__), .dout(n1420));
  buf1  g375(.din(new_new_n372__), .dout(n1423));
  buf1  g376(.din(new_new_n454__), .dout(n1426));
  buf1  g377(.din(new_new_n456__), .dout(n1429));
  buf1  g378(.din(new_new_n947__), .dout(n1432));
  buf1  g379(.din(new_new_n376__), .dout(n1435));
  buf1  g380(.din(new_new_n378__), .dout(n1438));
  buf1  g381(.din(new_new_n464__), .dout(n1441));
  buf1  g382(.din(new_new_n466__), .dout(n1444));
  buf1  g383(.din(new_new_n957__), .dout(n1447));
  buf1  g384(.din(new_new_n496__), .dout(n1450));
  buf1  g385(.din(new_new_n498__), .dout(n1453));
  buf1  g386(.din(new_new_n546__), .dout(n1456));
  buf1  g387(.din(new_new_n548__), .dout(n1459));
  not1  g388(.din(new_new_n956__), .dout(n1462));
  not1  g389(.din(new_new_n962__), .dout(n1465));
  not1  g390(.din(new_new_n960__), .dout(n1468));
  not1  g391(.din(new_new_n958__), .dout(n1471));
  not1  g392(.din(new_new_n950__), .dout(n1474));
  not1  g393(.din(new_new_n952__), .dout(n1477));
  not1  g394(.din(new_new_n954__), .dout(n1480));
  not1  g395(.din(new_new_n948__), .dout(n1483));
  buf1  g396(.din(new_new_n550__), .dout(n1486));
  buf1  g397(.din(new_new_n552__), .dout(n1489));
  not1  g398(.din(new_new_n946__), .dout(n1492));
  buf1  g399(.din(new_new_n578__), .dout(n1495));
  buf1  g400(.din(new_new_n580__), .dout(n1498));
  buf1  g401(.din(new_new_n582__), .dout(n1501));
  buf1  g402(.din(new_new_n584__), .dout(n1504));
  buf1  g403(.din(new_new_n967__), .dout(n1507));
  buf1  g404(.din(new_new_n969__), .dout(n1510));
  buf1  g405(.din(new_new_n971__), .dout(n1513));
  buf1  g406(.din(new_new_n965__), .dout(n1516));
  not1  g407(.din(new_new_n968__), .dout(n1519));
  not1  g408(.din(new_new_n970__), .dout(n1522));
  not1  g409(.din(new_new_n972__), .dout(n1525));
  not1  g410(.din(new_new_n966__), .dout(n1528));
  buf1  g411(.din(new_new_n963__), .dout(n1531));
  not1  g412(.din(new_new_n964__), .dout(n1534));
  buf1  g413(.din(new_new_n602__), .dout(n1537));
  buf1  g414(.din(new_new_n975__), .dout(n1540));
  buf1  g415(.din(new_new_n976__), .dout(n1543));
  buf1  g416(.din(new_new_n974__), .dout(n1546));
  not1  g417(.din(new_new_n977__), .dout(n1549));
  not1  g418(.din(new_new_n978__), .dout(n1552));
  buf1  g419(.din(new_new_n616__), .dout(n1555));
  buf1  g420(.din(new_new_n973__), .dout(n1558));
  not1  g421(.din(new_new_n979__), .dout(n1561));
  not1  g422(.din(new_new_n980__), .dout(n1564));
  buf1  g423(.din(new_new_n981__), .dout(n1567));
  buf1  g424(.din(new_new_n982__), .dout(n1570));
  not1  g425(.din(new_new_n757__), .dout(n1573));
  not1  g426(.din(new_new_n986__), .dout(n1576));
  buf1  g427(.din(new_new_n994__), .dout(n1579));
  not1  g428(.din(new_new_n760__), .dout(n1582));
  not1  g429(.din(new_new_n761__), .dout(n1585));
  not1  g430(.din(new_new_n762__), .dout(n1588));
  not1  g431(.din(new_new_n763__), .dout(n1591));
  buf1  g432(.din(new_new_n390__), .dout(n1594));
  buf1  g433(.din(new_new_n420__), .dout(n1597));
  buf1  g434(.din(new_new_n430__), .dout(n1600));
  buf1  g435(.din(new_new_n452__), .dout(n1603));
  buf1  g436(.din(new_new_n764__), .dout(n1606));
  not1  g437(.din(new_new_n766__), .dout(n1609));
  not1  g438(.din(new_new_n768__), .dout(n1612));
  not1  g439(.din(new_new_n770__), .dout(n1615));
  not1  g440(.din(new_new_n772__), .dout(n1618));
  buf1  g441(.din(new_new_n773__), .dout(n1621));
  buf1  g442(.din(new_new_n774__), .dout(n1624));
  buf1  g443(.din(new_new_n775__), .dout(n1627));
  buf1  g444(.din(new_new_n380__), .dout(n1630));
  buf1  g445(.din(new_new_n400__), .dout(n1633));
  buf1  g446(.din(new_new_n410__), .dout(n1636));
  buf1  g447(.din(new_new_n462__), .dout(n1639));
  buf1  g448(.din(new_new_n314__), .dout(n1642));
  buf1  g449(.din(new_new_n995__), .dout(n1645));
  buf1  g450(.din(new_new_n322__), .dout(n1648));
  buf1  g451(.din(new_new_n996__), .dout(n1651));
  buf1  g452(.din(new_new_n330__), .dout(n1654));
  buf1  g453(.din(new_new_n997__), .dout(n1657));
  buf1  g454(.din(new_new_n370__), .dout(n1660));
  buf1  g455(.din(new_new_n998__), .dout(n1663));
  buf1  g456(.din(new_new_n354__), .dout(n1666));
  buf1  g457(.din(new_new_n358__), .dout(n1669));
  buf1  g458(.din(new_new_n308__), .dout(n1672));
  buf1  g459(.din(new_new_n310__), .dout(n1675));
  buf1  g460(.din(new_new_n338__), .dout(n1678));
  buf1  g461(.din(new_new_n342__), .dout(n1681));
  buf1  g462(.din(new_new_n346__), .dout(n1684));
  buf1  g463(.din(new_new_n350__), .dout(n1687));
  buf1  g464(.din(new_new_n362__), .dout(n1690));
  buf1  g465(.din(new_new_n366__), .dout(n1693));
  buf1  g466(.din(new_new_n776__), .dout(n1696));
  buf1  g467(.din(new_new_n777__), .dout(n1699));
  buf1  g468(.din(new_new_n778__), .dout(n1702));
  buf1  g469(.din(new_new_n779__), .dout(n1705));
  buf1  g470(.din(new_new_n555__), .dout(new_new_n919__));
  buf1  g471(.din(new_new_n919__), .dout(new_new_n920__));
  buf1  g472(.din(new_new_n920__), .dout(new_new_n921__));
  buf1  g473(.din(new_new_n919__), .dout(new_new_n922__));
  buf1  g474(.din(new_new_n554__), .dout(new_new_n923__));
  buf1  g475(.din(new_new_n923__), .dout(new_new_n924__));
  buf1  g476(.din(new_new_n924__), .dout(new_new_n925__));
  buf1  g477(.din(new_new_n924__), .dout(new_new_n926__));
  buf1  g478(.din(new_new_n923__), .dout(new_new_n927__));
  buf1  g479(.din(new_new_n927__), .dout(new_new_n928__));
  buf1  g480(.din(new_new_n927__), .dout(new_new_n929__));
  buf1  g481(.din(new_new_n650__), .dout(new_new_n930__));
  buf1  g482(.din(new_new_n654__), .dout(new_new_n931__));
  buf1  g483(.din(new_new_n657__), .dout(new_new_n932__));
  buf1  g484(.din(new_new_n665__), .dout(new_new_n933__));
  buf1  g485(.din(new_new_n664__), .dout(new_new_n934__));
  buf1  g486(.din(new_new_n668__), .dout(new_new_n935__));
  buf1  g487(.din(new_new_n673__), .dout(new_new_n936__));
  buf1  g488(.din(new_new_n677__), .dout(new_new_n937__));
  buf1  g489(.din(new_new_n679__), .dout(new_new_n938__));
  buf1  g490(.din(new_new_n676__), .dout(new_new_n939__));
  buf1  g491(.din(new_new_n684__), .dout(new_new_n940__));
  buf1  g492(.din(new_new_n556__), .dout(new_new_n941__));
  buf1  g493(.din(new_new_n941__), .dout(new_new_n942__));
  buf1  g494(.din(new_new_n942__), .dout(new_new_n943__));
  buf1  g495(.din(new_new_n941__), .dout(new_new_n944__));
  buf1  g496(.din(new_new_n448__), .dout(new_new_n945__));
  buf1  g497(.din(new_new_n706__), .dout(new_new_n946__));
  buf1  g498(.din(new_new_n458__), .dout(new_new_n947__));
  buf1  g499(.din(new_new_n704__), .dout(new_new_n948__));
  buf1  g500(.din(new_new_n396__), .dout(new_new_n949__));
  buf1  g501(.din(new_new_n698__), .dout(new_new_n950__));
  buf1  g502(.din(new_new_n426__), .dout(new_new_n951__));
  buf1  g503(.din(new_new_n700__), .dout(new_new_n952__));
  buf1  g504(.din(new_new_n436__), .dout(new_new_n953__));
  buf1  g505(.din(new_new_n702__), .dout(new_new_n954__));
  buf1  g506(.din(new_new_n386__), .dout(new_new_n955__));
  buf1  g507(.din(new_new_n693__), .dout(new_new_n956__));
  buf1  g508(.din(new_new_n468__), .dout(new_new_n957__));
  buf1  g509(.din(new_new_n696__), .dout(new_new_n958__));
  buf1  g510(.din(new_new_n416__), .dout(new_new_n959__));
  buf1  g511(.din(new_new_n695__), .dout(new_new_n960__));
  buf1  g512(.din(new_new_n406__), .dout(new_new_n961__));
  buf1  g513(.din(new_new_n694__), .dout(new_new_n962__));
  buf1  g514(.din(new_new_n442__), .dout(new_new_n963__));
  buf1  g515(.din(new_new_n712__), .dout(new_new_n964__));
  buf1  g516(.din(new_new_n574__), .dout(new_new_n965__));
  buf1  g517(.din(new_new_n710__), .dout(new_new_n966__));
  buf1  g518(.din(new_new_n568__), .dout(new_new_n967__));
  buf1  g519(.din(new_new_n707__), .dout(new_new_n968__));
  buf1  g520(.din(new_new_n570__), .dout(new_new_n969__));
  buf1  g521(.din(new_new_n708__), .dout(new_new_n970__));
  buf1  g522(.din(new_new_n572__), .dout(new_new_n971__));
  buf1  g523(.din(new_new_n709__), .dout(new_new_n972__));
  buf1  g524(.din(new_new_n618__), .dout(new_new_n973__));
  buf1  g525(.din(new_new_n634__), .dout(new_new_n974__));
  buf1  g526(.din(new_new_n626__), .dout(new_new_n975__));
  buf1  g527(.din(new_new_n630__), .dout(new_new_n976__));
  buf1  g528(.din(new_new_n717__), .dout(new_new_n977__));
  buf1  g529(.din(new_new_n728__), .dout(new_new_n978__));
  buf1  g530(.din(new_new_n733__), .dout(new_new_n979__));
  buf1  g531(.din(new_new_n744__), .dout(new_new_n980__));
  buf1  g532(.din(new_new_n749__), .dout(new_new_n981__));
  buf1  g533(.din(new_new_n756__), .dout(new_new_n982__));
  buf1  g534(.din(new_new_n758__), .dout(new_new_n983__));
  buf1  g535(.din(new_new_n983__), .dout(new_new_n984__));
  buf1  g536(.din(new_new_n984__), .dout(new_new_n985__));
  buf1  g537(.din(new_new_n983__), .dout(new_new_n986__));
  buf1  g538(.din(new_new_n759__), .dout(new_new_n987__));
  buf1  g539(.din(new_new_n987__), .dout(new_new_n988__));
  buf1  g540(.din(new_new_n988__), .dout(new_new_n989__));
  buf1  g541(.din(new_new_n989__), .dout(new_new_n990__));
  buf1  g542(.din(new_new_n988__), .dout(new_new_n991__));
  buf1  g543(.din(new_new_n987__), .dout(new_new_n992__));
  buf1  g544(.din(new_new_n992__), .dout(new_new_n993__));
  buf1  g545(.din(new_new_n992__), .dout(new_new_n994__));
  buf1  g546(.din(new_new_n318__), .dout(new_new_n995__));
  buf1  g547(.din(new_new_n326__), .dout(new_new_n996__));
  buf1  g548(.din(new_new_n334__), .dout(new_new_n997__));
  buf1  g549(.din(new_new_n374__), .dout(new_new_n998__));
  always @ (posedge clock) begin
    n229_lo <= n1312;
    n253_lo <= n1315;
    n256_lo <= n1318;
    n259_lo <= n1321;
    n262_lo <= n1324;
    n277_lo <= n1327;
    n301_lo <= n1330;
    n304_lo <= n1333;
    n307_lo <= n1336;
    n310_lo <= n1339;
    n325_lo <= n1342;
    n349_lo <= n1345;
    n352_lo <= n1348;
    n355_lo <= n1351;
    n358_lo <= n1354;
    n373_lo <= n1357;
    n397_lo <= n1360;
    n400_lo <= n1363;
    n403_lo <= n1366;
    n406_lo <= n1369;
    n421_lo <= n1372;
    n445_lo <= n1375;
    n448_lo <= n1378;
    n451_lo <= n1381;
    n454_lo <= n1384;
    n469_lo <= n1387;
    n493_lo <= n1390;
    n496_lo <= n1393;
    n499_lo <= n1396;
    n502_lo <= n1399;
    n517_lo <= n1402;
    n520_lo <= n1405;
    n541_lo <= n1408;
    n544_lo <= n1411;
    n547_lo <= n1414;
    n550_lo <= n1417;
    n565_lo <= n1420;
    n589_lo <= n1423;
    n592_lo <= n1426;
    n595_lo <= n1429;
    n598_lo <= n1432;
    n613_lo <= n1435;
    n625_lo <= n1438;
    n628_lo <= n1441;
    n631_lo <= n1444;
    n634_lo <= n1447;
    n852_o2 <= n1450;
    n853_o2 <= n1453;
    n955_o2 <= n1456;
    n956_o2 <= n1459;
    n531_o2 <= n1462;
    n549_o2 <= n1465;
    n537_o2 <= n1468;
    n540_o2 <= n1471;
    n546_o2 <= n1474;
    n534_o2 <= n1477;
    n552_o2 <= n1480;
    n543_o2 <= n1483;
    n961_o2 <= n1486;
    n223_inv <= n1489;
    n555_o2 <= n1492;
    n1009_o2 <= n1495;
    n1010_o2 <= n1498;
    n1011_o2 <= n1501;
    n1012_o2 <= n1504;
    lo026_buf_o2 <= n1507;
    lo074_buf_o2 <= n1510;
    lo090_buf_o2 <= n1513;
    lo122_buf_o2 <= n1516;
    n510_o2 <= n1519;
    n498_o2 <= n1522;
    n516_o2 <= n1525;
    n507_o2 <= n1528;
    lo106_buf_o2 <= n1531;
    n519_o2 <= n1534;
    n1029_o2 <= n1537;
    n1041_o2 <= n1540;
    n1043_o2 <= n1543;
    n1045_o2 <= n1546;
    n558_o2 <= n1549;
    n563_o2 <= n1552;
    lo094_buf_o2 <= n1555;
    lo102_buf_o2 <= n1558;
    n522_o2 <= n1561;
    n298_inv <= n1564;
    n486_o2 <= n1567;
    n304_inv <= n1570;
    n564_o2 <= n1573;
    n528_o2 <= n1576;
    n492_o2 <= n1579;
    n530_o2 <= n1582;
    n548_o2 <= n1585;
    n536_o2 <= n1588;
    n539_o2 <= n1591;
    lo025_buf_o2 <= n1594;
    lo073_buf_o2 <= n1597;
    lo089_buf_o2 <= n1600;
    lo121_buf_o2 <= n1603;
    n509_o2 <= n1606;
    n513_o2 <= n1609;
    n501_o2 <= n1612;
    n504_o2 <= n1615;
    n495_o2 <= n1618;
    n497_o2 <= n1621;
    n515_o2 <= n1624;
    n506_o2 <= n1627;
    lo010_buf_o2 <= n1630;
    lo042_buf_o2 <= n1633;
    lo058_buf_o2 <= n1636;
    lo138_buf_o2 <= n1639;
    lo014_buf_o2 <= n1642;
    lo022_buf_o2 <= n1645;
    lo030_buf_o2 <= n1648;
    lo038_buf_o2 <= n1651;
    lo046_buf_o2 <= n1654;
    lo054_buf_o2 <= n1657;
    lo126_buf_o2 <= n1660;
    lo134_buf_o2 <= n1663;
    lo093_buf_o2 <= n1666;
    lo101_buf_o2 <= n1669;
    lo002_buf_o2 <= n1672;
    lo006_buf_o2 <= n1675;
    lo062_buf_o2 <= n1678;
    lo070_buf_o2 <= n1681;
    lo078_buf_o2 <= n1684;
    lo086_buf_o2 <= n1687;
    lo110_buf_o2 <= n1690;
    lo118_buf_o2 <= n1693;
    n476_o2 <= n1696;
    n482_o2 <= n1699;
    n478_o2 <= n1702;
    n479_o2 <= n1705;
  end
  initial begin
    n229_lo <= 1'b0;
    n253_lo <= 1'b0;
    n256_lo <= 1'b0;
    n259_lo <= 1'b0;
    n262_lo <= 1'b0;
    n277_lo <= 1'b0;
    n301_lo <= 1'b0;
    n304_lo <= 1'b0;
    n307_lo <= 1'b0;
    n310_lo <= 1'b0;
    n325_lo <= 1'b0;
    n349_lo <= 1'b0;
    n352_lo <= 1'b0;
    n355_lo <= 1'b0;
    n358_lo <= 1'b0;
    n373_lo <= 1'b0;
    n397_lo <= 1'b0;
    n400_lo <= 1'b0;
    n403_lo <= 1'b0;
    n406_lo <= 1'b0;
    n421_lo <= 1'b0;
    n445_lo <= 1'b0;
    n448_lo <= 1'b0;
    n451_lo <= 1'b0;
    n454_lo <= 1'b0;
    n469_lo <= 1'b0;
    n493_lo <= 1'b0;
    n496_lo <= 1'b0;
    n499_lo <= 1'b0;
    n502_lo <= 1'b0;
    n517_lo <= 1'b0;
    n520_lo <= 1'b0;
    n541_lo <= 1'b0;
    n544_lo <= 1'b0;
    n547_lo <= 1'b0;
    n550_lo <= 1'b0;
    n565_lo <= 1'b0;
    n589_lo <= 1'b0;
    n592_lo <= 1'b0;
    n595_lo <= 1'b0;
    n598_lo <= 1'b0;
    n613_lo <= 1'b0;
    n625_lo <= 1'b0;
    n628_lo <= 1'b0;
    n631_lo <= 1'b0;
    n634_lo <= 1'b0;
    n852_o2 <= 1'b0;
    n853_o2 <= 1'b0;
    n955_o2 <= 1'b0;
    n956_o2 <= 1'b0;
    n531_o2 <= 1'b0;
    n549_o2 <= 1'b0;
    n537_o2 <= 1'b0;
    n540_o2 <= 1'b0;
    n546_o2 <= 1'b0;
    n534_o2 <= 1'b0;
    n552_o2 <= 1'b0;
    n543_o2 <= 1'b0;
    n961_o2 <= 1'b0;
    n223_inv <= 1'b0;
    n555_o2 <= 1'b0;
    n1009_o2 <= 1'b0;
    n1010_o2 <= 1'b0;
    n1011_o2 <= 1'b0;
    n1012_o2 <= 1'b0;
    lo026_buf_o2 <= 1'b0;
    lo074_buf_o2 <= 1'b0;
    lo090_buf_o2 <= 1'b0;
    lo122_buf_o2 <= 1'b0;
    n510_o2 <= 1'b0;
    n498_o2 <= 1'b0;
    n516_o2 <= 1'b0;
    n507_o2 <= 1'b0;
    lo106_buf_o2 <= 1'b0;
    n519_o2 <= 1'b0;
    n1029_o2 <= 1'b0;
    n1041_o2 <= 1'b0;
    n1043_o2 <= 1'b0;
    n1045_o2 <= 1'b0;
    n558_o2 <= 1'b0;
    n563_o2 <= 1'b0;
    lo094_buf_o2 <= 1'b0;
    lo102_buf_o2 <= 1'b0;
    n522_o2 <= 1'b0;
    n298_inv <= 1'b0;
    n486_o2 <= 1'b0;
    n304_inv <= 1'b0;
    n564_o2 <= 1'b0;
    n528_o2 <= 1'b0;
    n492_o2 <= 1'b0;
    n530_o2 <= 1'b0;
    n548_o2 <= 1'b0;
    n536_o2 <= 1'b0;
    n539_o2 <= 1'b0;
    lo025_buf_o2 <= 1'b0;
    lo073_buf_o2 <= 1'b0;
    lo089_buf_o2 <= 1'b0;
    lo121_buf_o2 <= 1'b0;
    n509_o2 <= 1'b0;
    n513_o2 <= 1'b0;
    n501_o2 <= 1'b0;
    n504_o2 <= 1'b0;
    n495_o2 <= 1'b0;
    n497_o2 <= 1'b0;
    n515_o2 <= 1'b0;
    n506_o2 <= 1'b0;
    lo010_buf_o2 <= 1'b0;
    lo042_buf_o2 <= 1'b0;
    lo058_buf_o2 <= 1'b0;
    lo138_buf_o2 <= 1'b0;
    lo014_buf_o2 <= 1'b0;
    lo022_buf_o2 <= 1'b0;
    lo030_buf_o2 <= 1'b0;
    lo038_buf_o2 <= 1'b0;
    lo046_buf_o2 <= 1'b0;
    lo054_buf_o2 <= 1'b0;
    lo126_buf_o2 <= 1'b0;
    lo134_buf_o2 <= 1'b0;
    lo093_buf_o2 <= 1'b0;
    lo101_buf_o2 <= 1'b0;
    lo002_buf_o2 <= 1'b0;
    lo006_buf_o2 <= 1'b0;
    lo062_buf_o2 <= 1'b0;
    lo070_buf_o2 <= 1'b0;
    lo078_buf_o2 <= 1'b0;
    lo086_buf_o2 <= 1'b0;
    lo110_buf_o2 <= 1'b0;
    lo118_buf_o2 <= 1'b0;
    n476_o2 <= 1'b0;
    n482_o2 <= 1'b0;
    n478_o2 <= 1'b0;
    n479_o2 <= 1'b0;
  end
endmodule


