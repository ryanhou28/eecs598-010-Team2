
module mymod
(
  G1_p,
  G1_n,
  G2_p,
  G2_n,
  G3_p,
  G3_n,
  G4_p,
  G4_n,
  G5_p,
  G5_n,
  G6_p,
  G6_n,
  G7_p,
  G7_n,
  G8_p,
  G8_n,
  G9_p,
  G9_n,
  G10_p,
  G10_n,
  G11_p,
  G11_n,
  G12_p,
  G12_n,
  G13_p,
  G13_n,
  G14_p,
  G14_n,
  G15_p,
  G15_n,
  G16_p,
  G16_n,
  G17_p,
  G17_n,
  G18_p,
  G18_n,
  G19_p,
  G19_n,
  G20_p,
  G20_n,
  G21_p,
  G21_n,
  G22_p,
  G22_n,
  G23_p,
  G23_n,
  G24_p,
  G24_n,
  G25_p,
  G25_n,
  G26_p,
  G26_n,
  G27_p,
  G27_n,
  G28_p,
  G28_n,
  G29_p,
  G29_n,
  G30_p,
  G30_n,
  G31_p,
  G31_n,
  G32_p,
  G32_n,
  G33_p,
  G33_n,
  G34_p,
  G34_n,
  G35_p,
  G35_n,
  G36_p,
  G36_n,
  G37_p,
  G37_n,
  G38_p,
  G38_n,
  G39_p,
  G39_n,
  G40_p,
  G40_n,
  G41_p,
  G41_n,
  G42_p,
  G42_n,
  G43_p,
  G43_n,
  G44_p,
  G44_n,
  G45_p,
  G45_n,
  G46_p,
  G46_n,
  G47_p,
  G47_n,
  G48_p,
  G48_n,
  G49_p,
  G49_n,
  G50_p,
  G50_n,
  G3519_p,
  G3520_p,
  G3521_p,
  G3522_p,
  G3523_p,
  G3524_p,
  G3525_p,
  G3526_p,
  G3527_p,
  G3528_p,
  G3529_p,
  G3530_p,
  G3531_p,
  G3532_p,
  G3533_p,
  G3534_p,
  G3535_p,
  G3536_p,
  G3537_p,
  G3538_n,
  G3539_p,
  G3540_p
);

  input G1_p;input G1_n;input G2_p;input G2_n;input G3_p;input G3_n;input G4_p;input G4_n;input G5_p;input G5_n;input G6_p;input G6_n;input G7_p;input G7_n;input G8_p;input G8_n;input G9_p;input G9_n;input G10_p;input G10_n;input G11_p;input G11_n;input G12_p;input G12_n;input G13_p;input G13_n;input G14_p;input G14_n;input G15_p;input G15_n;input G16_p;input G16_n;input G17_p;input G17_n;input G18_p;input G18_n;input G19_p;input G19_n;input G20_p;input G20_n;input G21_p;input G21_n;input G22_p;input G22_n;input G23_p;input G23_n;input G24_p;input G24_n;input G25_p;input G25_n;input G26_p;input G26_n;input G27_p;input G27_n;input G28_p;input G28_n;input G29_p;input G29_n;input G30_p;input G30_n;input G31_p;input G31_n;input G32_p;input G32_n;input G33_p;input G33_n;input G34_p;input G34_n;input G35_p;input G35_n;input G36_p;input G36_n;input G37_p;input G37_n;input G38_p;input G38_n;input G39_p;input G39_n;input G40_p;input G40_n;input G41_p;input G41_n;input G42_p;input G42_n;input G43_p;input G43_n;input G44_p;input G44_n;input G45_p;input G45_n;input G46_p;input G46_n;input G47_p;input G47_n;input G48_p;input G48_n;input G49_p;input G49_n;input G50_p;input G50_n;
  output G3519_p;output G3520_p;output G3521_p;output G3522_p;output G3523_p;output G3524_p;output G3525_p;output G3526_p;output G3527_p;output G3528_p;output G3529_p;output G3530_p;output G3531_p;output G3532_p;output G3533_p;output G3534_p;output G3535_p;output G3536_p;output G3537_p;output G3538_n;output G3539_p;output G3540_p;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire g51_p;
  wire g51_n;
  wire g52_p;
  wire g52_n;
  wire g53_p;
  wire g53_n;
  wire g54_p;
  wire g54_n;
  wire g55_p;
  wire g55_n;
  wire g56_p;
  wire g56_n;
  wire g57_p;
  wire g57_n;
  wire g58_p;
  wire g58_n;
  wire g59_p;
  wire g59_n;
  wire g60_p;
  wire g60_n;
  wire g61_p;
  wire g61_n;
  wire g62_p;
  wire g62_n;
  wire g63_p;
  wire g63_n;
  wire g64_p;
  wire g64_n;
  wire g65_p;
  wire g65_n;
  wire g66_p;
  wire g66_n;
  wire g67_p;
  wire g67_n;
  wire g68_p;
  wire g68_n;
  wire g69_p;
  wire g69_n;
  wire g70_p;
  wire g70_n;
  wire g71_p;
  wire g71_n;
  wire g72_p;
  wire g72_n;
  wire g73_p;
  wire g73_n;
  wire g74_p;
  wire g74_n;
  wire g75_p;
  wire g75_n;
  wire g76_p;
  wire g76_n;
  wire g77_p;
  wire g77_n;
  wire g78_p;
  wire g78_n;
  wire g79_p;
  wire g79_n;
  wire g80_p;
  wire g80_n;
  wire g81_p;
  wire g81_n;
  wire g82_p;
  wire g82_n;
  wire g83_p;
  wire g83_n;
  wire g84_p;
  wire g84_n;
  wire g85_p;
  wire g85_n;
  wire g86_p;
  wire g86_n;
  wire g87_p;
  wire g87_n;
  wire g88_p;
  wire g88_n;
  wire g89_p;
  wire g89_n;
  wire g90_p;
  wire g90_n;
  wire g91_p;
  wire g91_n;
  wire g92_p;
  wire g92_n;
  wire g93_p;
  wire g93_n;
  wire g94_p;
  wire g94_n;
  wire g95_p;
  wire g95_n;
  wire g96_p;
  wire g96_n;
  wire g97_p;
  wire g97_n;
  wire g98_p;
  wire g98_n;
  wire g99_p;
  wire g99_n;
  wire g100_p;
  wire g100_n;
  wire g101_p;
  wire g101_n;
  wire g102_p;
  wire g102_n;
  wire g103_p;
  wire g103_n;
  wire g104_p;
  wire g104_n;
  wire g105_p;
  wire g105_n;
  wire g106_p;
  wire g106_n;
  wire g107_p;
  wire g107_n;
  wire g108_p;
  wire g108_n;
  wire g109_p;
  wire g109_n;
  wire g110_p;
  wire g110_n;
  wire g111_p;
  wire g111_n;
  wire g112_p;
  wire g112_n;
  wire g113_p;
  wire g113_n;
  wire g114_p;
  wire g114_n;
  wire g115_p;
  wire g115_n;
  wire g116_p;
  wire g116_n;
  wire g117_p;
  wire g117_n;
  wire g118_p;
  wire g118_n;
  wire g119_p;
  wire g119_n;
  wire g120_p;
  wire g120_n;
  wire g121_p;
  wire g121_n;
  wire g122_p;
  wire g122_n;
  wire g123_p;
  wire g123_n;
  wire g124_p;
  wire g124_n;
  wire g125_p;
  wire g125_n;
  wire g126_p;
  wire g126_n;
  wire g127_p;
  wire g127_n;
  wire g128_p;
  wire g128_n;
  wire g129_p;
  wire g129_n;
  wire g130_p;
  wire g130_n;
  wire g131_p;
  wire g131_n;
  wire g132_p;
  wire g132_n;
  wire g133_p;
  wire g133_n;
  wire g134_p;
  wire g134_n;
  wire g135_p;
  wire g135_n;
  wire g136_p;
  wire g136_n;
  wire g137_p;
  wire g137_n;
  wire g138_p;
  wire g138_n;
  wire g139_p;
  wire g139_n;
  wire g140_p;
  wire g140_n;
  wire g141_p;
  wire g141_n;
  wire g142_p;
  wire g142_n;
  wire g143_p;
  wire g143_n;
  wire g144_p;
  wire g144_n;
  wire g145_p;
  wire g145_n;
  wire g146_p;
  wire g146_n;
  wire g147_p;
  wire g147_n;
  wire g148_p;
  wire g148_n;
  wire g149_p;
  wire g149_n;
  wire g150_p;
  wire g150_n;
  wire g151_p;
  wire g151_n;
  wire g152_p;
  wire g152_n;
  wire g153_p;
  wire g153_n;
  wire g154_p;
  wire g154_n;
  wire g155_p;
  wire g155_n;
  wire g156_p;
  wire g156_n;
  wire g157_p;
  wire g157_n;
  wire g158_p;
  wire g158_n;
  wire g159_p;
  wire g159_n;
  wire g160_p;
  wire g160_n;
  wire g161_p;
  wire g161_n;
  wire g162_p;
  wire g162_n;
  wire g163_p;
  wire g163_n;
  wire g164_p;
  wire g164_n;
  wire g165_p;
  wire g165_n;
  wire g166_p;
  wire g166_n;
  wire g167_p;
  wire g167_n;
  wire g168_p;
  wire g168_n;
  wire g169_p;
  wire g169_n;
  wire g170_p;
  wire g170_n;
  wire g171_p;
  wire g171_n;
  wire g172_p;
  wire g172_n;
  wire g173_p;
  wire g173_n;
  wire g174_p;
  wire g174_n;
  wire g175_p;
  wire g175_n;
  wire g176_p;
  wire g176_n;
  wire g177_p;
  wire g177_n;
  wire g178_p;
  wire g178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire g686_p;
  wire g686_n;
  wire g687_p;
  wire g687_n;
  wire g688_p;
  wire g688_n;
  wire g689_p;
  wire g689_n;
  wire g690_p;
  wire g690_n;
  wire g691_p;
  wire g691_n;
  wire g692_p;
  wire g692_n;
  wire g693_p;
  wire g693_n;
  wire g694_p;
  wire g694_n;
  wire g695_p;
  wire g695_n;
  wire g696_p;
  wire g696_n;
  wire g697_p;
  wire g697_n;
  wire g698_p;
  wire g698_n;
  wire g699_p;
  wire g699_n;
  wire g700_p;
  wire g700_n;
  wire g701_p;
  wire g701_n;
  wire g702_p;
  wire g702_n;
  wire g703_p;
  wire g703_n;
  wire g704_p;
  wire g704_n;
  wire g705_p;
  wire g705_n;
  wire g706_p;
  wire g706_n;
  wire g707_p;
  wire g707_n;
  wire g708_p;
  wire g708_n;
  wire g709_p;
  wire g709_n;
  wire g710_p;
  wire g710_n;
  wire g711_p;
  wire g711_n;
  wire g712_p;
  wire g712_n;
  wire g713_p;
  wire g713_n;
  wire g714_p;
  wire g714_n;
  wire g715_p;
  wire g715_n;
  wire g716_p;
  wire g716_n;
  wire g717_p;
  wire g717_n;
  wire g718_p;
  wire g718_n;
  wire g719_p;
  wire g719_n;
  wire g720_p;
  wire g720_n;
  wire g721_p;
  wire g721_n;
  wire g722_p;
  wire g722_n;
  wire g723_p;
  wire g723_n;
  wire g724_p;
  wire g724_n;
  wire g725_p;
  wire g725_n;
  wire g726_p;
  wire g726_n;
  wire g727_p;
  wire g727_n;
  wire g728_p;
  wire g728_n;
  wire g729_p;
  wire g729_n;
  wire g730_p;
  wire g730_n;
  wire g731_p;
  wire g731_n;
  wire g732_p;
  wire g732_n;
  wire g733_p;
  wire g733_n;
  wire g734_p;
  wire g734_n;
  wire g735_p;
  wire g735_n;
  wire g736_p;
  wire g736_n;
  wire g737_p;
  wire g737_n;
  wire g738_p;
  wire g738_n;
  wire g739_p;
  wire g739_n;
  wire g740_p;
  wire g740_n;
  wire g741_p;
  wire g741_n;
  wire g742_p;
  wire g742_n;
  wire g743_p;
  wire g743_n;
  wire g744_p;
  wire g744_n;
  wire g745_p;
  wire g745_n;
  wire g746_p;
  wire g746_n;
  wire g747_p;
  wire g747_n;
  wire g748_p;
  wire g748_n;
  wire g749_p;
  wire g749_n;
  wire g750_p;
  wire g750_n;
  wire g751_p;
  wire g751_n;
  wire g752_p;
  wire g752_n;
  wire g753_p;
  wire g753_n;
  wire g754_p;
  wire g754_n;
  wire g755_p;
  wire g755_n;
  wire g756_p;
  wire g756_n;
  wire g757_p;
  wire g757_n;
  wire g758_p;
  wire g758_n;
  wire g759_p;
  wire g759_n;
  wire g760_p;
  wire g760_n;
  wire g761_p;
  wire g761_n;
  wire g762_p;
  wire g762_n;
  wire g763_p;
  wire g763_n;
  wire g764_p;
  wire g764_n;
  wire g765_p;
  wire g765_n;
  wire g766_p;
  wire g766_n;
  wire g767_p;
  wire g767_n;
  wire g768_p;
  wire g768_n;
  wire g769_p;
  wire g769_n;
  wire g770_p;
  wire g770_n;
  wire g771_p;
  wire g771_n;
  wire g772_p;
  wire g772_n;
  wire g773_p;
  wire g773_n;
  wire g774_p;
  wire g774_n;
  wire g775_p;
  wire g775_n;
  wire g776_p;
  wire g776_n;
  wire g777_p;
  wire g777_n;
  wire g778_p;
  wire g778_n;
  wire g779_p;
  wire g779_n;
  wire g780_p;
  wire g780_n;
  wire g781_p;
  wire g781_n;
  wire g782_p;
  wire g782_n;
  wire g783_p;
  wire g783_n;
  wire g784_p;
  wire g784_n;
  wire g785_p;
  wire g785_n;
  wire g786_p;
  wire g786_n;
  wire g787_p;
  wire g787_n;
  wire g788_p;
  wire g788_n;
  wire g789_p;
  wire g789_n;
  wire g790_p;
  wire g790_n;
  wire g791_p;
  wire g791_n;
  wire g792_p;
  wire g792_n;
  wire g793_p;
  wire g793_n;
  wire g794_p;
  wire g794_n;
  wire g795_p;
  wire g795_n;
  wire g796_p;
  wire g796_n;
  wire g797_p;
  wire g797_n;
  wire g798_p;
  wire g798_n;
  wire g799_p;
  wire g799_n;
  wire g800_p;
  wire g800_n;
  wire g801_p;
  wire g801_n;
  wire g802_p;
  wire g802_n;
  wire g803_p;
  wire g803_n;
  wire g804_p;
  wire g804_n;
  wire g805_p;
  wire g805_n;
  wire g806_p;
  wire g806_n;
  wire g807_p;
  wire g807_n;
  wire g808_p;
  wire g808_n;
  wire g809_p;
  wire g809_n;
  wire g810_p;
  wire g810_n;
  wire g811_p;
  wire g811_n;
  wire g812_p;
  wire g812_n;
  wire g813_p;
  wire g813_n;
  wire g814_p;
  wire g814_n;
  wire g815_p;
  wire g815_n;
  wire g816_p;
  wire g816_n;
  wire g817_p;
  wire g817_n;
  wire g818_p;
  wire g818_n;
  wire g819_p;
  wire g819_n;
  wire g820_p;
  wire g820_n;
  wire g821_p;
  wire g821_n;
  wire g822_p;
  wire g822_n;
  wire g823_p;
  wire g823_n;
  wire g824_p;
  wire g824_n;
  wire g825_p;
  wire g825_n;
  wire g826_p;
  wire g826_n;
  wire g827_p;
  wire g827_n;
  wire g828_p;
  wire g828_n;
  wire g829_p;
  wire g829_n;
  wire g830_p;
  wire g830_n;
  wire g831_p;
  wire g831_n;
  wire g832_p;
  wire g832_n;
  wire g833_p;
  wire g833_n;
  wire g834_p;
  wire g834_n;
  wire g835_p;
  wire g835_n;
  wire g836_p;
  wire g836_n;
  wire g837_p;
  wire g837_n;
  wire g838_p;
  wire g838_n;
  wire g839_p;
  wire g839_n;
  wire g840_p;
  wire g840_n;
  wire g841_p;
  wire g841_n;
  wire g842_p;
  wire g842_n;
  wire g843_p;
  wire g843_n;
  wire g844_p;
  wire g844_n;
  wire g845_p;
  wire g845_n;
  wire g846_p;
  wire g846_n;
  wire g847_p;
  wire g847_n;
  wire g848_p;
  wire g848_n;
  wire g849_p;
  wire g849_n;
  wire g850_p;
  wire g850_n;
  wire g851_p;
  wire g851_n;
  wire g852_p;
  wire g852_n;
  wire g853_p;
  wire g853_n;
  wire g854_p;
  wire g854_n;
  wire g855_p;
  wire g855_n;
  wire g856_p;
  wire g856_n;
  wire g857_p;
  wire g857_n;
  wire g858_p;
  wire g858_n;
  wire g859_p;
  wire g859_n;
  wire g860_p;
  wire g860_n;
  wire g861_p;
  wire g861_n;
  wire g862_p;
  wire g862_n;
  wire g863_p;
  wire g863_n;
  wire g864_p;
  wire g864_n;
  wire g865_p;
  wire g865_n;
  wire g866_p;
  wire g866_n;
  wire g867_p;
  wire g867_n;
  wire g868_p;
  wire g868_n;
  wire g869_p;
  wire g869_n;
  wire g870_p;
  wire g870_n;
  wire g871_p;
  wire g871_n;
  wire g872_p;
  wire g872_n;
  wire g873_p;
  wire g873_n;
  wire g874_p;
  wire g874_n;
  wire g875_p;
  wire g875_n;
  wire g876_p;
  wire g876_n;
  wire g877_p;
  wire g877_n;
  wire g878_p;
  wire g878_n;
  wire g879_p;
  wire g879_n;
  wire g880_p;
  wire g880_n;
  wire g881_p;
  wire g881_n;
  wire g882_p;
  wire g882_n;
  wire g883_p;
  wire g883_n;
  wire g884_p;
  wire g884_n;
  wire g885_p;
  wire g885_n;
  wire g886_p;
  wire g886_n;
  wire g887_p;
  wire g887_n;
  wire g888_p;
  wire g888_n;
  wire g889_p;
  wire g889_n;
  wire g890_p;
  wire g890_n;
  wire g891_p;
  wire g891_n;
  wire g892_p;
  wire g892_n;
  wire g893_p;
  wire g893_n;
  wire g894_p;
  wire g894_n;
  wire g895_p;
  wire g895_n;
  wire g896_p;
  wire g896_n;
  wire g897_p;
  wire g897_n;
  wire g898_p;
  wire g898_n;
  wire g899_p;
  wire g899_n;
  wire g900_p;
  wire g900_n;
  wire g901_p;
  wire g901_n;
  wire g902_p;
  wire g902_n;
  wire g903_p;
  wire g903_n;
  wire g904_p;
  wire g904_n;
  wire G7_n_spl_;
  wire G7_n_spl_0;
  wire G7_n_spl_00;
  wire G7_n_spl_000;
  wire G7_n_spl_0000;
  wire G7_n_spl_001;
  wire G7_n_spl_01;
  wire G7_n_spl_010;
  wire G7_n_spl_011;
  wire G7_n_spl_1;
  wire G7_n_spl_10;
  wire G7_n_spl_100;
  wire G7_n_spl_101;
  wire G7_n_spl_11;
  wire G7_n_spl_110;
  wire G7_n_spl_111;
  wire G8_n_spl_;
  wire G8_n_spl_0;
  wire G8_n_spl_00;
  wire G8_n_spl_000;
  wire G8_n_spl_001;
  wire G8_n_spl_01;
  wire G8_n_spl_010;
  wire G8_n_spl_011;
  wire G8_n_spl_1;
  wire G8_n_spl_10;
  wire G8_n_spl_100;
  wire G8_n_spl_101;
  wire G8_n_spl_11;
  wire G8_n_spl_110;
  wire G7_p_spl_;
  wire G7_p_spl_0;
  wire G7_p_spl_00;
  wire G7_p_spl_000;
  wire G7_p_spl_0000;
  wire G7_p_spl_0001;
  wire G7_p_spl_001;
  wire G7_p_spl_01;
  wire G7_p_spl_010;
  wire G7_p_spl_011;
  wire G7_p_spl_1;
  wire G7_p_spl_10;
  wire G7_p_spl_100;
  wire G7_p_spl_101;
  wire G7_p_spl_11;
  wire G7_p_spl_110;
  wire G7_p_spl_111;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire G8_p_spl_00;
  wire G8_p_spl_000;
  wire G8_p_spl_001;
  wire G8_p_spl_01;
  wire G8_p_spl_010;
  wire G8_p_spl_011;
  wire G8_p_spl_1;
  wire G8_p_spl_10;
  wire G8_p_spl_100;
  wire G8_p_spl_101;
  wire G8_p_spl_11;
  wire G8_p_spl_110;
  wire G8_p_spl_111;
  wire G9_n_spl_;
  wire G9_n_spl_0;
  wire G9_n_spl_00;
  wire G9_n_spl_000;
  wire G9_n_spl_001;
  wire G9_n_spl_01;
  wire G9_n_spl_010;
  wire G9_n_spl_011;
  wire G9_n_spl_1;
  wire G9_n_spl_10;
  wire G9_n_spl_100;
  wire G9_n_spl_101;
  wire G9_n_spl_11;
  wire G9_n_spl_110;
  wire g51_p_spl_;
  wire G9_p_spl_;
  wire G9_p_spl_0;
  wire G9_p_spl_00;
  wire G9_p_spl_000;
  wire G9_p_spl_001;
  wire G9_p_spl_01;
  wire G9_p_spl_010;
  wire G9_p_spl_011;
  wire G9_p_spl_1;
  wire G9_p_spl_10;
  wire G9_p_spl_100;
  wire G9_p_spl_101;
  wire G9_p_spl_11;
  wire G9_p_spl_110;
  wire g51_n_spl_;
  wire G10_n_spl_;
  wire G10_n_spl_0;
  wire G10_n_spl_00;
  wire G10_n_spl_000;
  wire G10_n_spl_001;
  wire G10_n_spl_01;
  wire G10_n_spl_010;
  wire G10_n_spl_011;
  wire G10_n_spl_1;
  wire G10_n_spl_10;
  wire G10_n_spl_100;
  wire G10_n_spl_101;
  wire G10_n_spl_11;
  wire G10_n_spl_110;
  wire g52_p_spl_;
  wire G12_n_spl_;
  wire G12_n_spl_0;
  wire G12_n_spl_00;
  wire G12_n_spl_000;
  wire G12_n_spl_001;
  wire G12_n_spl_01;
  wire G12_n_spl_010;
  wire G12_n_spl_011;
  wire G12_n_spl_1;
  wire G12_n_spl_10;
  wire G12_n_spl_100;
  wire G12_n_spl_101;
  wire G12_n_spl_11;
  wire G13_n_spl_;
  wire G13_n_spl_0;
  wire G13_n_spl_00;
  wire G13_n_spl_000;
  wire G13_n_spl_001;
  wire G13_n_spl_01;
  wire G13_n_spl_010;
  wire G13_n_spl_011;
  wire G13_n_spl_1;
  wire G13_n_spl_10;
  wire G13_n_spl_100;
  wire G13_n_spl_101;
  wire G13_n_spl_11;
  wire G13_n_spl_110;
  wire G12_p_spl_;
  wire G12_p_spl_0;
  wire G12_p_spl_00;
  wire G12_p_spl_000;
  wire G12_p_spl_001;
  wire G12_p_spl_01;
  wire G12_p_spl_010;
  wire G12_p_spl_011;
  wire G12_p_spl_1;
  wire G12_p_spl_10;
  wire G12_p_spl_100;
  wire G12_p_spl_101;
  wire G12_p_spl_11;
  wire G12_p_spl_110;
  wire G13_p_spl_;
  wire G13_p_spl_0;
  wire G13_p_spl_00;
  wire G13_p_spl_000;
  wire G13_p_spl_001;
  wire G13_p_spl_01;
  wire G13_p_spl_010;
  wire G13_p_spl_011;
  wire G13_p_spl_1;
  wire G13_p_spl_10;
  wire G13_p_spl_100;
  wire G13_p_spl_101;
  wire G13_p_spl_11;
  wire G13_p_spl_110;
  wire G13_p_spl_111;
  wire G11_p_spl_;
  wire G11_p_spl_0;
  wire G11_p_spl_00;
  wire G11_p_spl_000;
  wire G11_p_spl_001;
  wire G11_p_spl_01;
  wire G11_p_spl_010;
  wire G11_p_spl_011;
  wire G11_p_spl_1;
  wire G11_p_spl_10;
  wire G11_p_spl_100;
  wire G11_p_spl_101;
  wire G11_p_spl_11;
  wire g54_n_spl_;
  wire G11_n_spl_;
  wire G11_n_spl_0;
  wire G11_n_spl_00;
  wire G11_n_spl_000;
  wire G11_n_spl_001;
  wire G11_n_spl_01;
  wire G11_n_spl_010;
  wire G11_n_spl_011;
  wire G11_n_spl_1;
  wire G11_n_spl_10;
  wire G11_n_spl_100;
  wire G11_n_spl_11;
  wire g54_p_spl_;
  wire G1_n_spl_;
  wire G1_n_spl_0;
  wire G1_n_spl_00;
  wire G1_n_spl_000;
  wire G1_n_spl_001;
  wire G1_n_spl_01;
  wire G1_n_spl_010;
  wire G1_n_spl_1;
  wire G1_n_spl_10;
  wire G1_n_spl_11;
  wire G3_n_spl_;
  wire G3_n_spl_0;
  wire G3_n_spl_00;
  wire G3_n_spl_000;
  wire G3_n_spl_0000;
  wire G3_n_spl_0001;
  wire G3_n_spl_001;
  wire G3_n_spl_0010;
  wire G3_n_spl_01;
  wire G3_n_spl_010;
  wire G3_n_spl_011;
  wire G3_n_spl_1;
  wire G3_n_spl_10;
  wire G3_n_spl_100;
  wire G3_n_spl_101;
  wire G3_n_spl_11;
  wire G3_n_spl_110;
  wire G3_n_spl_111;
  wire G34_n_spl_;
  wire G34_n_spl_0;
  wire G34_n_spl_00;
  wire G34_n_spl_01;
  wire G34_n_spl_1;
  wire G34_n_spl_10;
  wire G32_n_spl_;
  wire G32_n_spl_0;
  wire G32_n_spl_00;
  wire G32_n_spl_01;
  wire G32_n_spl_1;
  wire G36_n_spl_;
  wire G36_n_spl_0;
  wire G36_n_spl_00;
  wire G36_n_spl_01;
  wire G36_n_spl_1;
  wire G10_p_spl_;
  wire G10_p_spl_0;
  wire G10_p_spl_00;
  wire G10_p_spl_000;
  wire G10_p_spl_001;
  wire G10_p_spl_01;
  wire G10_p_spl_010;
  wire G10_p_spl_011;
  wire G10_p_spl_1;
  wire G10_p_spl_10;
  wire G10_p_spl_100;
  wire G10_p_spl_101;
  wire G10_p_spl_11;
  wire G33_n_spl_;
  wire G33_n_spl_0;
  wire G33_n_spl_00;
  wire G33_n_spl_01;
  wire G33_n_spl_1;
  wire G14_p_spl_;
  wire G14_p_spl_0;
  wire G14_p_spl_00;
  wire G14_p_spl_000;
  wire G14_p_spl_001;
  wire G14_p_spl_01;
  wire G14_p_spl_010;
  wire G14_p_spl_011;
  wire G14_p_spl_1;
  wire G14_p_spl_10;
  wire G14_p_spl_100;
  wire G14_p_spl_101;
  wire G14_p_spl_11;
  wire G14_p_spl_110;
  wire G14_p_spl_111;
  wire G37_n_spl_;
  wire G37_n_spl_0;
  wire G37_n_spl_1;
  wire G31_n_spl_;
  wire G31_n_spl_0;
  wire G31_n_spl_00;
  wire G31_n_spl_01;
  wire G31_n_spl_1;
  wire G35_n_spl_;
  wire G35_n_spl_0;
  wire G35_n_spl_00;
  wire G35_n_spl_01;
  wire G35_n_spl_1;
  wire G35_n_spl_10;
  wire G30_n_spl_;
  wire G30_n_spl_0;
  wire G30_n_spl_00;
  wire G30_n_spl_01;
  wire G30_n_spl_1;
  wire G2_p_spl_;
  wire G2_p_spl_0;
  wire G2_p_spl_00;
  wire G2_p_spl_1;
  wire G1_p_spl_;
  wire G1_p_spl_0;
  wire G1_p_spl_00;
  wire G1_p_spl_000;
  wire G1_p_spl_01;
  wire G1_p_spl_1;
  wire G1_p_spl_10;
  wire G1_p_spl_11;
  wire G2_n_spl_;
  wire G2_n_spl_0;
  wire G2_n_spl_00;
  wire G2_n_spl_1;
  wire g73_p_spl_;
  wire g73_p_spl_0;
  wire G3_p_spl_;
  wire G3_p_spl_0;
  wire G3_p_spl_00;
  wire G3_p_spl_000;
  wire G3_p_spl_0000;
  wire G3_p_spl_0001;
  wire G3_p_spl_001;
  wire G3_p_spl_01;
  wire G3_p_spl_010;
  wire G3_p_spl_011;
  wire G3_p_spl_1;
  wire G3_p_spl_10;
  wire G3_p_spl_100;
  wire G3_p_spl_101;
  wire G3_p_spl_11;
  wire G3_p_spl_110;
  wire G3_p_spl_111;
  wire g73_n_spl_;
  wire g73_n_spl_0;
  wire g75_n_spl_;
  wire g75_p_spl_;
  wire g74_n_spl_;
  wire g76_n_spl_;
  wire g78_p_spl_;
  wire g78_n_spl_;
  wire g79_n_spl_;
  wire g79_n_spl_0;
  wire g79_n_spl_1;
  wire G36_p_spl_;
  wire G36_p_spl_0;
  wire G36_p_spl_1;
  wire G37_p_spl_;
  wire G37_p_spl_0;
  wire G34_p_spl_;
  wire G34_p_spl_0;
  wire G34_p_spl_00;
  wire G34_p_spl_1;
  wire G35_p_spl_;
  wire G35_p_spl_0;
  wire G35_p_spl_00;
  wire G35_p_spl_1;
  wire g87_p_spl_;
  wire g90_n_spl_;
  wire g87_n_spl_;
  wire g90_p_spl_;
  wire G32_p_spl_;
  wire G32_p_spl_0;
  wire G32_p_spl_00;
  wire G32_p_spl_1;
  wire G33_p_spl_;
  wire G33_p_spl_0;
  wire G33_p_spl_00;
  wire G33_p_spl_1;
  wire G30_p_spl_;
  wire G30_p_spl_0;
  wire G30_p_spl_00;
  wire G30_p_spl_1;
  wire G31_p_spl_;
  wire G31_p_spl_0;
  wire G31_p_spl_00;
  wire G31_p_spl_1;
  wire g96_n_spl_;
  wire g99_p_spl_;
  wire g96_p_spl_;
  wire g99_n_spl_;
  wire g102_p_spl_;
  wire g102_n_spl_;
  wire g106_n_spl_;
  wire g106_p_spl_;
  wire G14_n_spl_;
  wire G14_n_spl_0;
  wire G14_n_spl_00;
  wire G14_n_spl_000;
  wire G14_n_spl_001;
  wire G14_n_spl_01;
  wire G14_n_spl_010;
  wire G14_n_spl_011;
  wire G14_n_spl_1;
  wire G14_n_spl_10;
  wire G14_n_spl_100;
  wire G14_n_spl_101;
  wire G14_n_spl_11;
  wire G14_n_spl_110;
  wire G14_n_spl_111;
  wire g108_p_spl_;
  wire g111_n_spl_;
  wire g108_n_spl_;
  wire g111_p_spl_;
  wire g117_n_spl_;
  wire g117_p_spl_;
  wire g116_p_spl_;
  wire g119_n_spl_;
  wire g116_n_spl_;
  wire g119_p_spl_;
  wire g122_p_spl_;
  wire g122_n_spl_;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_00;
  wire G4_p_spl_000;
  wire G4_p_spl_0000;
  wire G4_p_spl_00000;
  wire G4_p_spl_00001;
  wire G4_p_spl_0001;
  wire G4_p_spl_00010;
  wire G4_p_spl_00011;
  wire G4_p_spl_001;
  wire G4_p_spl_0010;
  wire G4_p_spl_0011;
  wire G4_p_spl_01;
  wire G4_p_spl_010;
  wire G4_p_spl_0100;
  wire G4_p_spl_0101;
  wire G4_p_spl_011;
  wire G4_p_spl_0110;
  wire G4_p_spl_0111;
  wire G4_p_spl_1;
  wire G4_p_spl_10;
  wire G4_p_spl_100;
  wire G4_p_spl_1000;
  wire G4_p_spl_1001;
  wire G4_p_spl_101;
  wire G4_p_spl_1010;
  wire G4_p_spl_1011;
  wire G4_p_spl_11;
  wire G4_p_spl_110;
  wire G4_p_spl_1100;
  wire G4_p_spl_1101;
  wire G4_p_spl_111;
  wire G4_p_spl_1110;
  wire G4_p_spl_1111;
  wire G4_n_spl_;
  wire G4_n_spl_0;
  wire G4_n_spl_00;
  wire G4_n_spl_000;
  wire G4_n_spl_0000;
  wire G4_n_spl_00000;
  wire G4_n_spl_00001;
  wire G4_n_spl_0001;
  wire G4_n_spl_00010;
  wire G4_n_spl_00011;
  wire G4_n_spl_001;
  wire G4_n_spl_0010;
  wire G4_n_spl_0011;
  wire G4_n_spl_01;
  wire G4_n_spl_010;
  wire G4_n_spl_0100;
  wire G4_n_spl_0101;
  wire G4_n_spl_011;
  wire G4_n_spl_0110;
  wire G4_n_spl_0111;
  wire G4_n_spl_1;
  wire G4_n_spl_10;
  wire G4_n_spl_100;
  wire G4_n_spl_1000;
  wire G4_n_spl_1001;
  wire G4_n_spl_101;
  wire G4_n_spl_1010;
  wire G4_n_spl_1011;
  wire G4_n_spl_11;
  wire G4_n_spl_110;
  wire G4_n_spl_1100;
  wire G4_n_spl_1101;
  wire G4_n_spl_111;
  wire G4_n_spl_1110;
  wire G4_n_spl_1111;
  wire g126_n_spl_;
  wire g126_p_spl_;
  wire g129_p_spl_;
  wire g129_p_spl_0;
  wire g129_p_spl_00;
  wire g129_p_spl_000;
  wire g129_p_spl_001;
  wire g129_p_spl_01;
  wire g129_p_spl_1;
  wire g129_p_spl_10;
  wire g129_p_spl_11;
  wire g130_n_spl_;
  wire g130_n_spl_0;
  wire g130_n_spl_00;
  wire g130_n_spl_01;
  wire g130_n_spl_1;
  wire g130_n_spl_10;
  wire g130_n_spl_11;
  wire g129_n_spl_;
  wire g129_n_spl_0;
  wire g129_n_spl_00;
  wire g129_n_spl_000;
  wire g129_n_spl_001;
  wire g129_n_spl_01;
  wire g129_n_spl_1;
  wire g129_n_spl_10;
  wire g129_n_spl_11;
  wire g130_p_spl_;
  wire g130_p_spl_0;
  wire g130_p_spl_00;
  wire g130_p_spl_01;
  wire g130_p_spl_1;
  wire g130_p_spl_10;
  wire g130_p_spl_11;
  wire g131_p_spl_;
  wire g131_n_spl_;
  wire g133_n_spl_;
  wire g133_n_spl_0;
  wire g133_n_spl_1;
  wire g134_n_spl_;
  wire g134_n_spl_0;
  wire g133_p_spl_;
  wire g133_p_spl_0;
  wire g133_p_spl_1;
  wire g134_p_spl_;
  wire g134_p_spl_0;
  wire g137_n_spl_;
  wire g137_n_spl_0;
  wire g137_n_spl_00;
  wire g137_n_spl_000;
  wire g137_n_spl_01;
  wire g137_n_spl_1;
  wire g137_n_spl_10;
  wire g137_n_spl_11;
  wire g137_p_spl_;
  wire g137_p_spl_0;
  wire g137_p_spl_00;
  wire g137_p_spl_000;
  wire g137_p_spl_01;
  wire g137_p_spl_1;
  wire g137_p_spl_10;
  wire g137_p_spl_11;
  wire g138_p_spl_;
  wire g138_p_spl_0;
  wire g138_p_spl_00;
  wire g138_p_spl_01;
  wire g138_p_spl_1;
  wire g138_p_spl_10;
  wire g138_p_spl_11;
  wire g138_n_spl_;
  wire g138_n_spl_0;
  wire g138_n_spl_00;
  wire g138_n_spl_01;
  wire g138_n_spl_1;
  wire g138_n_spl_10;
  wire g138_n_spl_11;
  wire G39_p_spl_;
  wire G39_p_spl_0;
  wire G39_p_spl_00;
  wire G39_p_spl_000;
  wire G39_p_spl_01;
  wire G39_p_spl_1;
  wire G39_p_spl_10;
  wire G39_p_spl_11;
  wire G39_n_spl_;
  wire G39_n_spl_0;
  wire G39_n_spl_00;
  wire G39_n_spl_000;
  wire G39_n_spl_01;
  wire G39_n_spl_1;
  wire G39_n_spl_10;
  wire G39_n_spl_11;
  wire G5_p_spl_;
  wire G5_p_spl_0;
  wire G5_p_spl_00;
  wire G5_p_spl_01;
  wire G5_p_spl_1;
  wire G5_n_spl_;
  wire G5_n_spl_0;
  wire G5_n_spl_00;
  wire G5_n_spl_01;
  wire G5_n_spl_1;
  wire g146_n_spl_;
  wire g146_p_spl_;
  wire g147_n_spl_;
  wire g147_n_spl_0;
  wire g147_n_spl_00;
  wire g147_n_spl_000;
  wire g147_n_spl_01;
  wire g147_n_spl_1;
  wire g147_n_spl_10;
  wire g147_n_spl_11;
  wire g147_p_spl_;
  wire g147_p_spl_0;
  wire g147_p_spl_00;
  wire g147_p_spl_000;
  wire g147_p_spl_01;
  wire g147_p_spl_1;
  wire g147_p_spl_10;
  wire g147_p_spl_11;
  wire G6_n_spl_;
  wire G6_n_spl_0;
  wire G6_n_spl_00;
  wire G6_n_spl_01;
  wire G6_n_spl_1;
  wire G6_n_spl_10;
  wire G6_p_spl_;
  wire G6_p_spl_0;
  wire G6_p_spl_00;
  wire G6_p_spl_01;
  wire G6_p_spl_1;
  wire G6_p_spl_10;
  wire g149_p_spl_;
  wire g149_p_spl_0;
  wire g149_n_spl_;
  wire g149_n_spl_0;
  wire g148_p_spl_;
  wire g148_p_spl_0;
  wire g150_p_spl_;
  wire g150_p_spl_0;
  wire g150_p_spl_1;
  wire g148_n_spl_;
  wire g148_n_spl_0;
  wire g150_n_spl_;
  wire g150_n_spl_0;
  wire g150_n_spl_1;
  wire g153_p_spl_;
  wire g153_p_spl_0;
  wire g153_p_spl_00;
  wire g153_p_spl_01;
  wire g153_p_spl_1;
  wire g153_p_spl_10;
  wire g153_p_spl_11;
  wire g153_n_spl_;
  wire g153_n_spl_0;
  wire g153_n_spl_00;
  wire g153_n_spl_01;
  wire g153_n_spl_1;
  wire g153_n_spl_10;
  wire g153_n_spl_11;
  wire G41_n_spl_;
  wire G41_n_spl_0;
  wire G41_n_spl_00;
  wire G41_n_spl_01;
  wire G41_n_spl_1;
  wire G41_n_spl_10;
  wire G41_p_spl_;
  wire G41_p_spl_0;
  wire G41_p_spl_00;
  wire G41_p_spl_01;
  wire G41_p_spl_1;
  wire G41_p_spl_10;
  wire g151_n_spl_;
  wire g151_n_spl_0;
  wire g151_p_spl_;
  wire g151_p_spl_0;
  wire G25_n_spl_;
  wire G26_n_spl_;
  wire G26_n_spl_0;
  wire G25_p_spl_;
  wire G26_p_spl_;
  wire G26_p_spl_0;
  wire g161_p_spl_;
  wire g161_p_spl_0;
  wire g161_p_spl_1;
  wire g162_n_spl_;
  wire g162_n_spl_0;
  wire g162_n_spl_00;
  wire g162_n_spl_000;
  wire g162_n_spl_01;
  wire g162_n_spl_1;
  wire g162_n_spl_10;
  wire g162_n_spl_11;
  wire g161_n_spl_;
  wire g161_n_spl_0;
  wire g161_n_spl_1;
  wire g162_p_spl_;
  wire g162_p_spl_0;
  wire g162_p_spl_00;
  wire g162_p_spl_000;
  wire g162_p_spl_01;
  wire g162_p_spl_1;
  wire g162_p_spl_10;
  wire g162_p_spl_11;
  wire g145_p_spl_;
  wire g145_p_spl_0;
  wire g145_n_spl_;
  wire g145_n_spl_0;
  wire G23_n_spl_;
  wire G24_n_spl_;
  wire G24_n_spl_0;
  wire G24_n_spl_1;
  wire G23_p_spl_;
  wire G24_p_spl_;
  wire G24_p_spl_0;
  wire G24_p_spl_1;
  wire g165_n_spl_;
  wire g165_n_spl_0;
  wire g165_n_spl_00;
  wire g165_n_spl_01;
  wire g165_n_spl_1;
  wire g165_n_spl_10;
  wire g165_n_spl_11;
  wire g165_p_spl_;
  wire g165_p_spl_0;
  wire g165_p_spl_00;
  wire g165_p_spl_01;
  wire g165_p_spl_1;
  wire g165_p_spl_10;
  wire g165_p_spl_11;
  wire g167_n_spl_;
  wire g167_n_spl_0;
  wire g167_p_spl_;
  wire g167_p_spl_0;
  wire g169_n_spl_;
  wire g169_p_spl_;
  wire G40_n_spl_;
  wire G40_n_spl_0;
  wire G40_n_spl_00;
  wire G40_n_spl_01;
  wire G40_n_spl_1;
  wire G40_n_spl_10;
  wire G40_p_spl_;
  wire G40_p_spl_0;
  wire G40_p_spl_00;
  wire G40_p_spl_01;
  wire G40_p_spl_1;
  wire G40_p_spl_10;
  wire g186_p_spl_;
  wire g186_p_spl_0;
  wire g186_p_spl_1;
  wire g186_n_spl_;
  wire g186_n_spl_0;
  wire g186_n_spl_1;
  wire g177_p_spl_;
  wire g177_p_spl_0;
  wire g177_n_spl_;
  wire g177_n_spl_0;
  wire g190_n_spl_;
  wire g190_n_spl_0;
  wire g190_p_spl_;
  wire g190_p_spl_0;
  wire g196_n_spl_;
  wire g196_p_spl_;
  wire g212_p_spl_;
  wire g212_p_spl_0;
  wire g212_p_spl_1;
  wire g212_n_spl_;
  wire g212_n_spl_0;
  wire g212_n_spl_1;
  wire g202_p_spl_;
  wire g202_p_spl_0;
  wire g202_n_spl_;
  wire g202_n_spl_0;
  wire g216_n_spl_;
  wire g216_p_spl_;
  wire g223_n_spl_;
  wire g238_p_spl_;
  wire g238_p_spl_0;
  wire g238_p_spl_1;
  wire g238_n_spl_;
  wire g238_n_spl_0;
  wire g238_n_spl_1;
  wire g229_p_spl_;
  wire g229_p_spl_0;
  wire g229_n_spl_;
  wire g229_n_spl_0;
  wire g242_n_spl_;
  wire g242_n_spl_0;
  wire g242_p_spl_;
  wire g242_p_spl_0;
  wire g217_p_spl_;
  wire g217_p_spl_0;
  wire g217_p_spl_1;
  wire g243_p_spl_;
  wire g243_p_spl_0;
  wire g217_n_spl_;
  wire g217_n_spl_0;
  wire g217_n_spl_1;
  wire g243_n_spl_;
  wire g243_n_spl_0;
  wire g191_p_spl_;
  wire g191_p_spl_0;
  wire g244_p_spl_;
  wire g191_n_spl_;
  wire g191_n_spl_0;
  wire g244_n_spl_;
  wire g168_p_spl_;
  wire g168_p_spl_0;
  wire g245_p_spl_;
  wire g168_n_spl_;
  wire g168_n_spl_0;
  wire g245_n_spl_;
  wire g248_n_spl_;
  wire g248_n_spl_0;
  wire g248_n_spl_1;
  wire g248_p_spl_;
  wire g248_p_spl_0;
  wire g248_p_spl_1;
  wire g259_p_spl_;
  wire g259_p_spl_0;
  wire g259_p_spl_00;
  wire g259_p_spl_1;
  wire g259_n_spl_;
  wire g259_n_spl_0;
  wire g259_n_spl_00;
  wire g259_n_spl_1;
  wire g260_n_spl_;
  wire g260_n_spl_0;
  wire g260_n_spl_1;
  wire g260_p_spl_;
  wire g260_p_spl_0;
  wire g260_p_spl_1;
  wire g269_p_spl_;
  wire g269_n_spl_;
  wire g257_p_spl_;
  wire g257_p_spl_0;
  wire g257_n_spl_;
  wire g257_n_spl_0;
  wire g273_n_spl_;
  wire g273_n_spl_0;
  wire g273_p_spl_;
  wire g273_p_spl_0;
  wire g291_p_spl_;
  wire g291_n_spl_;
  wire g282_p_spl_;
  wire g282_p_spl_0;
  wire g282_n_spl_;
  wire g282_n_spl_0;
  wire g295_n_spl_;
  wire g295_n_spl_0;
  wire g295_p_spl_;
  wire g295_p_spl_0;
  wire G21_p_spl_;
  wire G21_p_spl_0;
  wire G21_p_spl_00;
  wire G21_p_spl_01;
  wire G21_p_spl_1;
  wire G21_p_spl_10;
  wire G21_p_spl_11;
  wire G21_n_spl_;
  wire G21_n_spl_0;
  wire G21_n_spl_00;
  wire G21_n_spl_01;
  wire G21_n_spl_1;
  wire G21_n_spl_10;
  wire G21_n_spl_11;
  wire G29_n_spl_;
  wire G29_p_spl_;
  wire g315_p_spl_;
  wire g315_n_spl_;
  wire g306_p_spl_;
  wire g306_p_spl_0;
  wire g306_n_spl_;
  wire g306_n_spl_0;
  wire g319_n_spl_;
  wire g319_p_spl_;
  wire g326_n_spl_;
  wire G22_p_spl_;
  wire G22_p_spl_0;
  wire G22_p_spl_00;
  wire G22_p_spl_01;
  wire G22_p_spl_1;
  wire G22_p_spl_10;
  wire G22_p_spl_11;
  wire G22_n_spl_;
  wire G22_n_spl_0;
  wire G22_n_spl_00;
  wire G22_n_spl_01;
  wire G22_n_spl_1;
  wire G22_n_spl_10;
  wire G22_n_spl_11;
  wire g341_p_spl_;
  wire g341_n_spl_;
  wire g332_p_spl_;
  wire g332_p_spl_0;
  wire g332_n_spl_;
  wire g332_n_spl_0;
  wire g345_n_spl_;
  wire g345_n_spl_0;
  wire g345_p_spl_;
  wire g345_p_spl_0;
  wire g320_p_spl_;
  wire g320_p_spl_0;
  wire g320_p_spl_1;
  wire g346_p_spl_;
  wire g346_p_spl_0;
  wire g320_n_spl_;
  wire g320_n_spl_0;
  wire g320_n_spl_1;
  wire g346_n_spl_;
  wire g346_n_spl_0;
  wire g296_p_spl_;
  wire g296_p_spl_0;
  wire g347_p_spl_;
  wire g296_n_spl_;
  wire g296_n_spl_0;
  wire g347_n_spl_;
  wire g274_p_spl_;
  wire g274_p_spl_0;
  wire g348_p_spl_;
  wire g274_n_spl_;
  wire g274_n_spl_0;
  wire g348_n_spl_;
  wire g246_p_spl_;
  wire g349_p_spl_;
  wire g349_p_spl_0;
  wire g349_p_spl_1;
  wire g356_n_spl_;
  wire g363_n_spl_;
  wire G27_p_spl_;
  wire G27_p_spl_0;
  wire g79_p_spl_;
  wire g79_p_spl_0;
  wire G27_n_spl_;
  wire G48_p_spl_;
  wire g365_p_spl_;
  wire g365_p_spl_0;
  wire g365_p_spl_1;
  wire G48_n_spl_;
  wire g365_n_spl_;
  wire g365_n_spl_0;
  wire g365_n_spl_1;
  wire g366_p_spl_;
  wire g366_p_spl_0;
  wire g366_p_spl_00;
  wire g366_p_spl_000;
  wire g366_p_spl_001;
  wire g366_p_spl_01;
  wire g366_p_spl_010;
  wire g366_p_spl_011;
  wire g366_p_spl_1;
  wire g366_p_spl_10;
  wire g366_p_spl_100;
  wire g366_p_spl_101;
  wire g366_p_spl_11;
  wire g366_n_spl_;
  wire g366_n_spl_0;
  wire g366_n_spl_00;
  wire g366_n_spl_000;
  wire g366_n_spl_001;
  wire g366_n_spl_01;
  wire g366_n_spl_010;
  wire g366_n_spl_011;
  wire g366_n_spl_1;
  wire g366_n_spl_10;
  wire g366_n_spl_100;
  wire g366_n_spl_101;
  wire g366_n_spl_11;
  wire g367_n_spl_;
  wire g367_p_spl_;
  wire g371_n_spl_;
  wire g371_p_spl_;
  wire G47_p_spl_;
  wire G47_p_spl_0;
  wire G47_p_spl_00;
  wire G47_p_spl_01;
  wire G47_p_spl_1;
  wire G47_p_spl_10;
  wire g374_p_spl_;
  wire g374_p_spl_0;
  wire g374_p_spl_1;
  wire G47_n_spl_;
  wire G47_n_spl_0;
  wire G47_n_spl_00;
  wire G47_n_spl_01;
  wire G47_n_spl_1;
  wire G47_n_spl_10;
  wire g374_n_spl_;
  wire g374_n_spl_0;
  wire g374_n_spl_1;
  wire g370_n_spl_;
  wire g370_n_spl_0;
  wire g370_n_spl_1;
  wire g370_p_spl_;
  wire g370_p_spl_0;
  wire g370_p_spl_1;
  wire g76_p_spl_;
  wire g377_n_spl_;
  wire g377_n_spl_0;
  wire g377_n_spl_00;
  wire g377_n_spl_01;
  wire g377_n_spl_1;
  wire g377_n_spl_10;
  wire g377_n_spl_11;
  wire g379_p_spl_;
  wire g379_p_spl_0;
  wire g379_p_spl_00;
  wire g379_p_spl_01;
  wire g379_p_spl_1;
  wire g379_p_spl_10;
  wire g382_p_spl_;
  wire g382_n_spl_;
  wire g377_p_spl_;
  wire g377_p_spl_0;
  wire g377_p_spl_00;
  wire g377_p_spl_01;
  wire g377_p_spl_1;
  wire g377_p_spl_10;
  wire g384_p_spl_;
  wire g384_p_spl_0;
  wire g384_p_spl_00;
  wire g384_p_spl_01;
  wire g384_p_spl_1;
  wire g384_p_spl_10;
  wire g384_n_spl_;
  wire g384_n_spl_0;
  wire g384_n_spl_00;
  wire g384_n_spl_01;
  wire g384_n_spl_1;
  wire g384_n_spl_10;
  wire g387_n_spl_;
  wire g387_n_spl_0;
  wire g387_p_spl_;
  wire g387_p_spl_0;
  wire g385_n_spl_;
  wire g385_n_spl_0;
  wire g385_n_spl_00;
  wire g385_n_spl_000;
  wire g385_n_spl_001;
  wire g385_n_spl_01;
  wire g385_n_spl_1;
  wire g385_n_spl_10;
  wire g385_n_spl_11;
  wire g385_p_spl_;
  wire g385_p_spl_0;
  wire g385_p_spl_00;
  wire g385_p_spl_000;
  wire g385_p_spl_001;
  wire g385_p_spl_01;
  wire g385_p_spl_1;
  wire g385_p_spl_10;
  wire g385_p_spl_11;
  wire g390_p_spl_;
  wire g390_p_spl_0;
  wire g390_p_spl_1;
  wire g390_n_spl_;
  wire g390_n_spl_0;
  wire g390_n_spl_1;
  wire g394_n_spl_;
  wire g394_n_spl_0;
  wire g394_n_spl_00;
  wire g394_n_spl_01;
  wire g394_n_spl_1;
  wire g394_p_spl_;
  wire g394_p_spl_0;
  wire g394_p_spl_00;
  wire g394_p_spl_01;
  wire g394_p_spl_1;
  wire g55_n_spl_;
  wire g393_p_spl_;
  wire g393_p_spl_0;
  wire g393_p_spl_00;
  wire g393_p_spl_000;
  wire g393_p_spl_001;
  wire g393_p_spl_01;
  wire g393_p_spl_010;
  wire g393_p_spl_011;
  wire g393_p_spl_1;
  wire g393_p_spl_10;
  wire g393_p_spl_100;
  wire g393_p_spl_101;
  wire g393_p_spl_11;
  wire g393_p_spl_110;
  wire g393_p_spl_111;
  wire g393_n_spl_;
  wire g393_n_spl_0;
  wire g393_n_spl_00;
  wire g393_n_spl_000;
  wire g393_n_spl_001;
  wire g393_n_spl_01;
  wire g393_n_spl_010;
  wire g393_n_spl_011;
  wire g393_n_spl_1;
  wire g393_n_spl_10;
  wire g393_n_spl_100;
  wire g393_n_spl_101;
  wire g393_n_spl_11;
  wire g393_n_spl_110;
  wire g393_n_spl_111;
  wire g404_n_spl_;
  wire g404_n_spl_0;
  wire g404_p_spl_;
  wire g404_p_spl_0;
  wire g403_n_spl_;
  wire g403_n_spl_0;
  wire g403_n_spl_1;
  wire g405_p_spl_;
  wire g403_p_spl_;
  wire g403_p_spl_0;
  wire g403_p_spl_1;
  wire g405_n_spl_;
  wire G45_p_spl_;
  wire g406_n_spl_;
  wire g406_n_spl_0;
  wire g406_n_spl_00;
  wire g406_n_spl_000;
  wire g406_n_spl_0000;
  wire g406_n_spl_001;
  wire g406_n_spl_01;
  wire g406_n_spl_010;
  wire g406_n_spl_011;
  wire g406_n_spl_1;
  wire g406_n_spl_10;
  wire g406_n_spl_100;
  wire g406_n_spl_101;
  wire g406_n_spl_11;
  wire g406_n_spl_110;
  wire g406_n_spl_111;
  wire G45_n_spl_;
  wire g406_p_spl_;
  wire g406_p_spl_0;
  wire g406_p_spl_00;
  wire g406_p_spl_000;
  wire g406_p_spl_0000;
  wire g406_p_spl_001;
  wire g406_p_spl_01;
  wire g406_p_spl_010;
  wire g406_p_spl_011;
  wire g406_p_spl_1;
  wire g406_p_spl_10;
  wire g406_p_spl_100;
  wire g406_p_spl_101;
  wire g406_p_spl_11;
  wire g406_p_spl_110;
  wire g406_p_spl_111;
  wire g408_p_spl_;
  wire g408_n_spl_;
  wire G44_p_spl_;
  wire G44_p_spl_0;
  wire g409_n_spl_;
  wire g409_n_spl_0;
  wire g409_n_spl_00;
  wire g409_n_spl_000;
  wire g409_n_spl_001;
  wire g409_n_spl_01;
  wire g409_n_spl_010;
  wire g409_n_spl_011;
  wire g409_n_spl_1;
  wire g409_n_spl_10;
  wire g409_n_spl_100;
  wire g409_n_spl_101;
  wire g409_n_spl_11;
  wire g409_n_spl_110;
  wire g409_n_spl_111;
  wire G44_n_spl_;
  wire G44_n_spl_0;
  wire g409_p_spl_;
  wire g409_p_spl_0;
  wire g409_p_spl_00;
  wire g409_p_spl_000;
  wire g409_p_spl_001;
  wire g409_p_spl_01;
  wire g409_p_spl_010;
  wire g409_p_spl_011;
  wire g409_p_spl_1;
  wire g409_p_spl_10;
  wire g409_p_spl_100;
  wire g409_p_spl_101;
  wire g409_p_spl_11;
  wire g409_p_spl_110;
  wire g409_p_spl_111;
  wire G42_p_spl_;
  wire G42_p_spl_0;
  wire G42_p_spl_1;
  wire g412_n_spl_;
  wire g412_n_spl_0;
  wire g412_n_spl_00;
  wire g412_n_spl_000;
  wire g412_n_spl_0000;
  wire g412_n_spl_0001;
  wire g412_n_spl_001;
  wire g412_n_spl_0010;
  wire g412_n_spl_01;
  wire g412_n_spl_010;
  wire g412_n_spl_011;
  wire g412_n_spl_1;
  wire g412_n_spl_10;
  wire g412_n_spl_100;
  wire g412_n_spl_101;
  wire g412_n_spl_11;
  wire g412_n_spl_110;
  wire g412_n_spl_111;
  wire G42_n_spl_;
  wire G42_n_spl_0;
  wire G42_n_spl_1;
  wire g412_p_spl_;
  wire g412_p_spl_0;
  wire g412_p_spl_00;
  wire g412_p_spl_000;
  wire g412_p_spl_0000;
  wire g412_p_spl_0001;
  wire g412_p_spl_001;
  wire g412_p_spl_0010;
  wire g412_p_spl_01;
  wire g412_p_spl_010;
  wire g412_p_spl_011;
  wire g412_p_spl_1;
  wire g412_p_spl_10;
  wire g412_p_spl_100;
  wire g412_p_spl_101;
  wire g412_p_spl_11;
  wire g412_p_spl_110;
  wire g412_p_spl_111;
  wire g414_n_spl_;
  wire g414_n_spl_0;
  wire g414_n_spl_00;
  wire g414_n_spl_000;
  wire g414_n_spl_0000;
  wire g414_n_spl_0001;
  wire g414_n_spl_001;
  wire g414_n_spl_01;
  wire g414_n_spl_010;
  wire g414_n_spl_011;
  wire g414_n_spl_1;
  wire g414_n_spl_10;
  wire g414_n_spl_100;
  wire g414_n_spl_101;
  wire g414_n_spl_11;
  wire g414_n_spl_110;
  wire g414_n_spl_111;
  wire g414_p_spl_;
  wire g414_p_spl_0;
  wire g414_p_spl_00;
  wire g414_p_spl_000;
  wire g414_p_spl_0000;
  wire g414_p_spl_0001;
  wire g414_p_spl_001;
  wire g414_p_spl_01;
  wire g414_p_spl_010;
  wire g414_p_spl_011;
  wire g414_p_spl_1;
  wire g414_p_spl_10;
  wire g414_p_spl_100;
  wire g414_p_spl_101;
  wire g414_p_spl_11;
  wire g414_p_spl_110;
  wire g414_p_spl_111;
  wire G43_p_spl_;
  wire G43_p_spl_0;
  wire G43_p_spl_1;
  wire G43_n_spl_;
  wire G43_n_spl_0;
  wire G43_n_spl_1;
  wire g416_p_spl_;
  wire g416_n_spl_;
  wire g423_n_spl_;
  wire g423_n_spl_0;
  wire g423_n_spl_00;
  wire g423_n_spl_000;
  wire g423_n_spl_001;
  wire g423_n_spl_01;
  wire g423_n_spl_010;
  wire g423_n_spl_011;
  wire g423_n_spl_1;
  wire g423_n_spl_10;
  wire g423_n_spl_11;
  wire g423_p_spl_;
  wire g423_p_spl_0;
  wire g423_p_spl_00;
  wire g423_p_spl_000;
  wire g423_p_spl_001;
  wire g423_p_spl_01;
  wire g423_p_spl_010;
  wire g423_p_spl_011;
  wire g423_p_spl_1;
  wire g423_p_spl_10;
  wire g423_p_spl_11;
  wire g425_n_spl_;
  wire g425_n_spl_0;
  wire g425_n_spl_00;
  wire g425_n_spl_000;
  wire g425_n_spl_001;
  wire g425_n_spl_01;
  wire g425_n_spl_010;
  wire g425_n_spl_011;
  wire g425_n_spl_1;
  wire g425_n_spl_10;
  wire g425_n_spl_100;
  wire g425_n_spl_101;
  wire g425_n_spl_11;
  wire g425_p_spl_;
  wire g425_p_spl_0;
  wire g425_p_spl_00;
  wire g425_p_spl_000;
  wire g425_p_spl_001;
  wire g425_p_spl_01;
  wire g425_p_spl_010;
  wire g425_p_spl_011;
  wire g425_p_spl_1;
  wire g425_p_spl_10;
  wire g425_p_spl_100;
  wire g425_p_spl_101;
  wire g425_p_spl_11;
  wire g432_n_spl_;
  wire g432_p_spl_;
  wire g430_n_spl_;
  wire g430_p_spl_;
  wire g438_n_spl_;
  wire g438_p_spl_;
  wire g440_n_spl_;
  wire g441_n_spl_;
  wire g440_p_spl_;
  wire g441_p_spl_;
  wire g439_p_spl_;
  wire g439_n_spl_;
  wire g453_n_spl_;
  wire g453_p_spl_;
  wire g452_p_spl_;
  wire g452_p_spl_0;
  wire g452_p_spl_1;
  wire g456_p_spl_;
  wire g456_p_spl_0;
  wire g456_p_spl_1;
  wire g452_n_spl_;
  wire g452_n_spl_0;
  wire g452_n_spl_1;
  wire g456_n_spl_;
  wire g456_n_spl_0;
  wire g456_n_spl_1;
  wire G20_p_spl_;
  wire G20_p_spl_0;
  wire G20_p_spl_00;
  wire G20_p_spl_1;
  wire G20_n_spl_;
  wire G20_n_spl_0;
  wire G20_n_spl_00;
  wire G20_n_spl_1;
  wire G18_p_spl_;
  wire G18_p_spl_0;
  wire G18_p_spl_1;
  wire G18_n_spl_;
  wire G18_n_spl_0;
  wire G18_n_spl_1;
  wire G19_p_spl_;
  wire G19_p_spl_0;
  wire G19_p_spl_00;
  wire G19_p_spl_1;
  wire G19_n_spl_;
  wire G19_n_spl_0;
  wire G19_n_spl_00;
  wire G19_n_spl_1;
  wire g480_n_spl_;
  wire g480_p_spl_;
  wire g500_p_spl_;
  wire g500_p_spl_0;
  wire g500_n_spl_;
  wire g500_n_spl_0;
  wire g379_n_spl_;
  wire g379_n_spl_0;
  wire g379_n_spl_00;
  wire g379_n_spl_01;
  wire g379_n_spl_1;
  wire g503_n_spl_;
  wire g503_p_spl_;
  wire g501_p_spl_;
  wire g504_p_spl_;
  wire g501_n_spl_;
  wire g504_n_spl_;
  wire g510_n_spl_;
  wire g510_p_spl_;
  wire g514_n_spl_;
  wire g514_p_spl_;
  wire g513_p_spl_;
  wire g513_p_spl_0;
  wire g513_p_spl_00;
  wire g513_p_spl_1;
  wire g517_p_spl_;
  wire g517_p_spl_0;
  wire g517_p_spl_00;
  wire g517_p_spl_1;
  wire g513_n_spl_;
  wire g513_n_spl_0;
  wire g513_n_spl_00;
  wire g513_n_spl_1;
  wire g517_n_spl_;
  wire g517_n_spl_0;
  wire g517_n_spl_00;
  wire g517_n_spl_1;
  wire g518_p_spl_;
  wire g519_p_spl_;
  wire g518_n_spl_;
  wire g519_n_spl_;
  wire g349_n_spl_;
  wire g520_n_spl_;
  wire g521_p_spl_;
  wire g521_p_spl_0;
  wire g520_p_spl_;
  wire g521_n_spl_;
  wire g521_n_spl_0;
  wire g528_p_spl_;
  wire g528_n_spl_;
  wire g530_n_spl_;
  wire g530_n_spl_0;
  wire g530_p_spl_;
  wire g530_p_spl_0;
  wire g527_n_spl_;
  wire g527_n_spl_0;
  wire g534_n_spl_;
  wire g534_n_spl_0;
  wire g534_n_spl_1;
  wire g527_p_spl_;
  wire g527_p_spl_0;
  wire g534_p_spl_;
  wire g534_p_spl_0;
  wire g534_p_spl_1;
  wire g552_n_spl_;
  wire g552_p_spl_;
  wire g555_p_spl_;
  wire g555_p_spl_0;
  wire g555_n_spl_;
  wire g555_n_spl_0;
  wire g569_n_spl_;
  wire g569_p_spl_;
  wire g579_n_spl_;
  wire g579_p_spl_;
  wire g594_n_spl_;
  wire g594_p_spl_;
  wire g376_p_spl_;
  wire g376_p_spl_0;
  wire g597_n_spl_;
  wire g597_n_spl_0;
  wire g597_n_spl_00;
  wire g597_n_spl_1;
  wire g376_n_spl_;
  wire g597_p_spl_;
  wire g597_p_spl_0;
  wire g597_p_spl_00;
  wire g597_p_spl_1;
  wire g600_n_spl_;
  wire g600_p_spl_;
  wire g601_n_spl_;
  wire g601_p_spl_;
  wire g603_n_spl_;
  wire g603_p_spl_;
  wire g605_p_spl_;
  wire g605_n_spl_;
  wire g598_n_spl_;
  wire g608_n_spl_;
  wire g598_p_spl_;
  wire g608_p_spl_;
  wire g613_n_spl_;
  wire g613_p_spl_;
  wire g617_p_spl_;
  wire g617_n_spl_;
  wire g616_n_spl_;
  wire g616_n_spl_0;
  wire g616_n_spl_1;
  wire g620_n_spl_;
  wire g620_n_spl_0;
  wire g620_n_spl_1;
  wire g616_p_spl_;
  wire g616_p_spl_0;
  wire g616_p_spl_1;
  wire g620_p_spl_;
  wire g620_p_spl_0;
  wire g620_p_spl_1;
  wire g628_n_spl_;
  wire g628_n_spl_0;
  wire g628_p_spl_;
  wire g628_p_spl_0;
  wire g653_n_spl_;
  wire g654_n_spl_;
  wire g653_p_spl_;
  wire g654_p_spl_;
  wire g649_p_spl_;
  wire g649_n_spl_;
  wire g685_p_spl_;
  wire g685_n_spl_;
  wire g706_n_spl_;
  wire g706_p_spl_;
  wire g705_n_spl_;
  wire g705_p_spl_;
  wire g723_p_spl_;
  wire g723_n_spl_;
  wire g726_p_spl_;
  wire g726_n_spl_;
  wire g724_p_spl_;
  wire g724_p_spl_0;
  wire g729_p_spl_;
  wire g724_n_spl_;
  wire g724_n_spl_0;
  wire g729_n_spl_;
  wire g730_n_spl_;
  wire g730_n_spl_0;
  wire g730_p_spl_;
  wire g730_p_spl_0;
  wire g733_p_spl_;
  wire g735_n_spl_;
  wire g733_n_spl_;
  wire g735_p_spl_;
  wire g738_n_spl_;
  wire g738_n_spl_0;
  wire g738_n_spl_1;
  wire g740_n_spl_;
  wire g740_n_spl_0;
  wire g738_p_spl_;
  wire g738_p_spl_0;
  wire g738_p_spl_1;
  wire g740_p_spl_;
  wire g740_p_spl_0;
  wire g732_p_spl_;
  wire g732_p_spl_0;
  wire g732_p_spl_1;
  wire g741_n_spl_;
  wire g741_n_spl_0;
  wire g732_n_spl_;
  wire g732_n_spl_0;
  wire g732_n_spl_1;
  wire g741_p_spl_;
  wire g741_p_spl_0;
  wire G17_p_spl_;
  wire G17_p_spl_0;
  wire G17_n_spl_;
  wire G17_n_spl_0;
  wire G16_n_spl_;
  wire G16_p_spl_;
  wire g779_n_spl_;
  wire g779_p_spl_;
  wire g782_p_spl_;
  wire g782_p_spl_0;
  wire g782_n_spl_;
  wire g782_n_spl_0;
  wire g818_p_spl_;
  wire g818_n_spl_;
  wire g626_p_spl_;
  wire g722_p_spl_;
  wire g626_n_spl_;
  wire g626_n_spl_0;
  wire g722_n_spl_;
  wire g722_n_spl_0;
  wire g778_p_spl_;
  wire g827_p_spl_;
  wire g778_n_spl_;
  wire g778_n_spl_0;
  wire g827_n_spl_;
  wire g827_n_spl_0;
  wire g509_p_spl_;
  wire g866_p_spl_;
  wire g509_n_spl_;
  wire g509_n_spl_0;
  wire g866_n_spl_;
  wire g866_n_spl_0;
  wire g451_p_spl_;
  wire g679_p_spl_;
  wire g451_n_spl_;
  wire g451_n_spl_0;
  wire g679_n_spl_;
  wire g679_n_spl_0;
  wire g869_n_spl_;
  wire g870_n_spl_;
  wire g868_n_spl_;
  wire g868_n_spl_0;
  wire g867_n_spl_;
  wire g874_n_spl_;
  wire g873_n_spl_;
  wire g879_p_spl_;
  wire g881_n_spl_;
  wire g879_n_spl_;
  wire g881_p_spl_;
  wire G50_n_spl_;
  wire g888_n_spl_;
  wire g888_n_spl_0;
  wire g888_n_spl_1;
  wire G50_p_spl_;
  wire g888_p_spl_;
  wire g888_p_spl_0;
  wire g888_p_spl_1;
  wire g886_p_spl_;
  wire g886_p_spl_0;
  wire g886_p_spl_1;
  wire g892_n_spl_;
  wire g886_n_spl_;
  wire g886_n_spl_0;
  wire g886_n_spl_1;
  wire g892_p_spl_;
  wire g884_n_spl_;
  wire g884_p_spl_;

  LA
  g_g51_p
  (
    .dout(g51_p),
    .din1(G7_n_spl_0000),
    .din2(G8_n_spl_000)
  );


  FA
  g_g51_n
  (
    .dout(g51_n),
    .din1(G7_p_spl_0000),
    .din2(G8_p_spl_000)
  );


  LA
  g_g52_p
  (
    .dout(g52_p),
    .din1(G9_n_spl_000),
    .din2(g51_p_spl_)
  );


  FA
  g_g52_n
  (
    .dout(g52_n),
    .din1(G9_p_spl_000),
    .din2(g51_n_spl_)
  );


  LA
  g_g53_p
  (
    .dout(g53_p),
    .din1(G10_n_spl_000),
    .din2(g52_p_spl_)
  );


  LA
  g_g54_p
  (
    .dout(g54_p),
    .din1(G12_n_spl_000),
    .din2(G13_n_spl_000)
  );


  FA
  g_g54_n
  (
    .dout(g54_n),
    .din1(G12_p_spl_000),
    .din2(G13_p_spl_000)
  );


  LA
  g_g55_p
  (
    .dout(g55_p),
    .din1(G11_p_spl_000),
    .din2(g54_n_spl_)
  );


  FA
  g_g55_n
  (
    .dout(g55_n),
    .din1(G11_n_spl_000),
    .din2(g54_p_spl_)
  );


  LA
  g_g56_p
  (
    .dout(g56_p),
    .din1(G1_n_spl_000),
    .din2(G3_n_spl_0000)
  );


  FA
  g_g57_n
  (
    .dout(g57_n),
    .din1(G11_p_spl_000),
    .din2(G34_n_spl_00)
  );


  FA
  g_g58_n
  (
    .dout(g58_n),
    .din1(G9_p_spl_000),
    .din2(G32_n_spl_00)
  );


  LA
  g_g59_p
  (
    .dout(g59_p),
    .din1(g57_n),
    .din2(g58_n)
  );


  FA
  g_g60_n
  (
    .dout(g60_n),
    .din1(G13_p_spl_000),
    .din2(G36_n_spl_00)
  );


  FA
  g_g61_n
  (
    .dout(g61_n),
    .din1(G10_p_spl_000),
    .din2(G33_n_spl_00)
  );


  LA
  g_g62_p
  (
    .dout(g62_p),
    .din1(g60_n),
    .din2(g61_n)
  );


  LA
  g_g63_p
  (
    .dout(g63_p),
    .din1(g59_p),
    .din2(g62_p)
  );


  FA
  g_g64_n
  (
    .dout(g64_n),
    .din1(G14_p_spl_000),
    .din2(G37_n_spl_0)
  );


  FA
  g_g65_n
  (
    .dout(g65_n),
    .din1(G8_p_spl_000),
    .din2(G31_n_spl_00)
  );


  LA
  g_g66_p
  (
    .dout(g66_p),
    .din1(g64_n),
    .din2(g65_n)
  );


  FA
  g_g67_n
  (
    .dout(g67_n),
    .din1(G12_p_spl_000),
    .din2(G35_n_spl_00)
  );


  FA
  g_g68_n
  (
    .dout(g68_n),
    .din1(G7_p_spl_0000),
    .din2(G30_n_spl_00)
  );


  LA
  g_g69_p
  (
    .dout(g69_p),
    .din1(g67_n),
    .din2(g68_n)
  );


  LA
  g_g70_p
  (
    .dout(g70_p),
    .din1(g66_p),
    .din2(g69_p)
  );


  LA
  g_g71_p
  (
    .dout(g71_p),
    .din1(g63_p),
    .din2(g70_p)
  );


  FA
  g_g72_n
  (
    .dout(g72_n),
    .din1(g56_p),
    .din2(g71_p)
  );


  LA
  g_g73_p
  (
    .dout(g73_p),
    .din1(G1_n_spl_000),
    .din2(G2_p_spl_00)
  );


  FA
  g_g73_n
  (
    .dout(g73_n),
    .din1(G1_p_spl_000),
    .din2(G2_n_spl_00)
  );


  LA
  g_g74_p
  (
    .dout(g74_p),
    .din1(G3_n_spl_0000),
    .din2(g73_p_spl_0)
  );


  FA
  g_g74_n
  (
    .dout(g74_n),
    .din1(G3_p_spl_0000),
    .din2(g73_n_spl_0)
  );


  LA
  g_g75_p
  (
    .dout(g75_p),
    .din1(G8_n_spl_000),
    .din2(G9_n_spl_000)
  );


  FA
  g_g75_n
  (
    .dout(g75_n),
    .din1(G8_p_spl_001),
    .din2(G9_p_spl_001)
  );


  LA
  g_g76_p
  (
    .dout(g76_p),
    .din1(G7_n_spl_0000),
    .din2(g75_n_spl_)
  );


  FA
  g_g76_n
  (
    .dout(g76_n),
    .din1(G7_p_spl_0001),
    .din2(g75_p_spl_)
  );


  FA
  g_g77_n
  (
    .dout(g77_n),
    .din1(g74_n_spl_),
    .din2(g76_n_spl_)
  );


  LA
  g_g78_p
  (
    .dout(g78_p),
    .din1(G1_n_spl_001),
    .din2(G2_n_spl_00)
  );


  FA
  g_g78_n
  (
    .dout(g78_n),
    .din1(G1_p_spl_000),
    .din2(G2_p_spl_00)
  );


  LA
  g_g79_p
  (
    .dout(g79_p),
    .din1(G3_n_spl_0001),
    .din2(g78_p_spl_)
  );


  FA
  g_g79_n
  (
    .dout(g79_n),
    .din1(G3_p_spl_0000),
    .din2(g78_n_spl_)
  );


  LA
  g_g80_p
  (
    .dout(g80_p),
    .din1(G35_n_spl_00),
    .din2(G36_n_spl_00)
  );


  FA
  g_g81_n
  (
    .dout(g81_n),
    .din1(G34_n_spl_00),
    .din2(g80_p)
  );


  FA
  g_g82_n
  (
    .dout(g82_n),
    .din1(g79_n_spl_0),
    .din2(g81_n)
  );


  LA
  g_g83_p
  (
    .dout(g83_p),
    .din1(g77_n),
    .din2(g82_n)
  );


  LA
  g_g84_p
  (
    .dout(g84_p),
    .din1(g72_n),
    .din2(g83_p)
  );


  LA
  g_g85_p
  (
    .dout(g85_p),
    .din1(G36_n_spl_01),
    .din2(G37_n_spl_0)
  );


  FA
  g_g85_n
  (
    .dout(g85_n),
    .din1(G36_p_spl_0),
    .din2(G37_p_spl_0)
  );


  LA
  g_g86_p
  (
    .dout(g86_p),
    .din1(G36_p_spl_0),
    .din2(G37_p_spl_0)
  );


  FA
  g_g86_n
  (
    .dout(g86_n),
    .din1(G36_n_spl_01),
    .din2(G37_n_spl_1)
  );


  LA
  g_g87_p
  (
    .dout(g87_p),
    .din1(g85_n),
    .din2(g86_n)
  );


  FA
  g_g87_n
  (
    .dout(g87_n),
    .din1(g85_p),
    .din2(g86_p)
  );


  LA
  g_g88_p
  (
    .dout(g88_p),
    .din1(G34_n_spl_01),
    .din2(G35_n_spl_01)
  );


  FA
  g_g88_n
  (
    .dout(g88_n),
    .din1(G34_p_spl_00),
    .din2(G35_p_spl_00)
  );


  LA
  g_g89_p
  (
    .dout(g89_p),
    .din1(G34_p_spl_00),
    .din2(G35_p_spl_00)
  );


  FA
  g_g89_n
  (
    .dout(g89_n),
    .din1(G34_n_spl_01),
    .din2(G35_n_spl_01)
  );


  LA
  g_g90_p
  (
    .dout(g90_p),
    .din1(g88_n),
    .din2(g89_n)
  );


  FA
  g_g90_n
  (
    .dout(g90_n),
    .din1(g88_p),
    .din2(g89_p)
  );


  LA
  g_g91_p
  (
    .dout(g91_p),
    .din1(g87_p_spl_),
    .din2(g90_n_spl_)
  );


  FA
  g_g91_n
  (
    .dout(g91_n),
    .din1(g87_n_spl_),
    .din2(g90_p_spl_)
  );


  LA
  g_g92_p
  (
    .dout(g92_p),
    .din1(g87_n_spl_),
    .din2(g90_p_spl_)
  );


  FA
  g_g92_n
  (
    .dout(g92_n),
    .din1(g87_p_spl_),
    .din2(g90_n_spl_)
  );


  LA
  g_g93_p
  (
    .dout(g93_p),
    .din1(g91_n),
    .din2(g92_n)
  );


  FA
  g_g93_n
  (
    .dout(g93_n),
    .din1(g91_p),
    .din2(g92_p)
  );


  LA
  g_g94_p
  (
    .dout(g94_p),
    .din1(G32_n_spl_00),
    .din2(G33_n_spl_00)
  );


  FA
  g_g94_n
  (
    .dout(g94_n),
    .din1(G32_p_spl_00),
    .din2(G33_p_spl_00)
  );


  LA
  g_g95_p
  (
    .dout(g95_p),
    .din1(G32_p_spl_00),
    .din2(G33_p_spl_00)
  );


  FA
  g_g95_n
  (
    .dout(g95_n),
    .din1(G32_n_spl_01),
    .din2(G33_n_spl_01)
  );


  LA
  g_g96_p
  (
    .dout(g96_p),
    .din1(g94_n),
    .din2(g95_n)
  );


  FA
  g_g96_n
  (
    .dout(g96_n),
    .din1(g94_p),
    .din2(g95_p)
  );


  LA
  g_g97_p
  (
    .dout(g97_p),
    .din1(G30_n_spl_00),
    .din2(G31_n_spl_00)
  );


  FA
  g_g97_n
  (
    .dout(g97_n),
    .din1(G30_p_spl_00),
    .din2(G31_p_spl_00)
  );


  LA
  g_g98_p
  (
    .dout(g98_p),
    .din1(G30_p_spl_00),
    .din2(G31_p_spl_00)
  );


  FA
  g_g98_n
  (
    .dout(g98_n),
    .din1(G30_n_spl_01),
    .din2(G31_n_spl_01)
  );


  LA
  g_g99_p
  (
    .dout(g99_p),
    .din1(g97_n),
    .din2(g98_n)
  );


  FA
  g_g99_n
  (
    .dout(g99_n),
    .din1(g97_p),
    .din2(g98_p)
  );


  LA
  g_g100_p
  (
    .dout(g100_p),
    .din1(g96_n_spl_),
    .din2(g99_p_spl_)
  );


  FA
  g_g100_n
  (
    .dout(g100_n),
    .din1(g96_p_spl_),
    .din2(g99_n_spl_)
  );


  LA
  g_g101_p
  (
    .dout(g101_p),
    .din1(g96_p_spl_),
    .din2(g99_n_spl_)
  );


  FA
  g_g101_n
  (
    .dout(g101_n),
    .din1(g96_n_spl_),
    .din2(g99_p_spl_)
  );


  LA
  g_g102_p
  (
    .dout(g102_p),
    .din1(g100_n),
    .din2(g101_n)
  );


  FA
  g_g102_n
  (
    .dout(g102_n),
    .din1(g100_p),
    .din2(g101_p)
  );


  FA
  g_g103_n
  (
    .dout(g103_n),
    .din1(g93_p),
    .din2(g102_p_spl_)
  );


  FA
  g_g104_n
  (
    .dout(g104_n),
    .din1(g93_n),
    .din2(g102_n_spl_)
  );


  LA
  g_g105_p
  (
    .dout(g105_p),
    .din1(g103_n),
    .din2(g104_n)
  );


  LA
  g_g106_p
  (
    .dout(g106_p),
    .din1(G11_n_spl_000),
    .din2(G12_n_spl_000)
  );


  FA
  g_g106_n
  (
    .dout(g106_n),
    .din1(G11_p_spl_001),
    .din2(G12_p_spl_001)
  );


  LA
  g_g107_p
  (
    .dout(g107_p),
    .din1(G11_p_spl_001),
    .din2(G12_p_spl_001)
  );


  FA
  g_g107_n
  (
    .dout(g107_n),
    .din1(G11_n_spl_001),
    .din2(G12_n_spl_001)
  );


  LA
  g_g108_p
  (
    .dout(g108_p),
    .din1(g106_n_spl_),
    .din2(g107_n)
  );


  FA
  g_g108_n
  (
    .dout(g108_n),
    .din1(g106_p_spl_),
    .din2(g107_p)
  );


  LA
  g_g109_p
  (
    .dout(g109_p),
    .din1(G13_n_spl_000),
    .din2(G14_n_spl_000)
  );


  FA
  g_g109_n
  (
    .dout(g109_n),
    .din1(G13_p_spl_001),
    .din2(G14_p_spl_000)
  );


  LA
  g_g110_p
  (
    .dout(g110_p),
    .din1(G13_p_spl_001),
    .din2(G14_p_spl_001)
  );


  FA
  g_g110_n
  (
    .dout(g110_n),
    .din1(G13_n_spl_001),
    .din2(G14_n_spl_000)
  );


  LA
  g_g111_p
  (
    .dout(g111_p),
    .din1(g109_n),
    .din2(g110_n)
  );


  FA
  g_g111_n
  (
    .dout(g111_n),
    .din1(g109_p),
    .din2(g110_p)
  );


  LA
  g_g112_p
  (
    .dout(g112_p),
    .din1(g108_p_spl_),
    .din2(g111_n_spl_)
  );


  FA
  g_g112_n
  (
    .dout(g112_n),
    .din1(g108_n_spl_),
    .din2(g111_p_spl_)
  );


  LA
  g_g113_p
  (
    .dout(g113_p),
    .din1(g108_n_spl_),
    .din2(g111_p_spl_)
  );


  FA
  g_g113_n
  (
    .dout(g113_n),
    .din1(g108_p_spl_),
    .din2(g111_n_spl_)
  );


  LA
  g_g114_p
  (
    .dout(g114_p),
    .din1(g112_n),
    .din2(g113_n)
  );


  FA
  g_g114_n
  (
    .dout(g114_n),
    .din1(g112_p),
    .din2(g113_p)
  );


  LA
  g_g115_p
  (
    .dout(g115_p),
    .din1(G7_p_spl_0001),
    .din2(G8_p_spl_001)
  );


  FA
  g_g115_n
  (
    .dout(g115_n),
    .din1(G7_n_spl_000),
    .din2(G8_n_spl_001)
  );


  LA
  g_g116_p
  (
    .dout(g116_p),
    .din1(g51_n_spl_),
    .din2(g115_n)
  );


  FA
  g_g116_n
  (
    .dout(g116_n),
    .din1(g51_p_spl_),
    .din2(g115_p)
  );


  LA
  g_g117_p
  (
    .dout(g117_p),
    .din1(G9_n_spl_001),
    .din2(G10_n_spl_000)
  );


  FA
  g_g117_n
  (
    .dout(g117_n),
    .din1(G9_p_spl_001),
    .din2(G10_p_spl_000)
  );


  LA
  g_g118_p
  (
    .dout(g118_p),
    .din1(G9_p_spl_010),
    .din2(G10_p_spl_001)
  );


  FA
  g_g118_n
  (
    .dout(g118_n),
    .din1(G9_n_spl_001),
    .din2(G10_n_spl_001)
  );


  LA
  g_g119_p
  (
    .dout(g119_p),
    .din1(g117_n_spl_),
    .din2(g118_n)
  );


  FA
  g_g119_n
  (
    .dout(g119_n),
    .din1(g117_p_spl_),
    .din2(g118_p)
  );


  LA
  g_g120_p
  (
    .dout(g120_p),
    .din1(g116_p_spl_),
    .din2(g119_n_spl_)
  );


  FA
  g_g120_n
  (
    .dout(g120_n),
    .din1(g116_n_spl_),
    .din2(g119_p_spl_)
  );


  LA
  g_g121_p
  (
    .dout(g121_p),
    .din1(g116_n_spl_),
    .din2(g119_p_spl_)
  );


  FA
  g_g121_n
  (
    .dout(g121_n),
    .din1(g116_p_spl_),
    .din2(g119_n_spl_)
  );


  LA
  g_g122_p
  (
    .dout(g122_p),
    .din1(g120_n),
    .din2(g121_n)
  );


  FA
  g_g122_n
  (
    .dout(g122_n),
    .din1(g120_p),
    .din2(g121_p)
  );


  LA
  g_g123_p
  (
    .dout(g123_p),
    .din1(g114_n),
    .din2(g122_p_spl_)
  );


  LA
  g_g124_p
  (
    .dout(g124_p),
    .din1(g114_p),
    .din2(g122_n_spl_)
  );


  FA
  g_g125_n
  (
    .dout(g125_n),
    .din1(g123_p),
    .din2(g124_p)
  );


  LA
  g_g126_p
  (
    .dout(g126_p),
    .din1(G1_p_spl_00),
    .din2(G2_p_spl_0)
  );


  FA
  g_g126_n
  (
    .dout(g126_n),
    .din1(G1_n_spl_001),
    .din2(G2_n_spl_0)
  );


  LA
  g_g127_p
  (
    .dout(g127_p),
    .din1(G1_p_spl_01),
    .din2(G3_p_spl_0001)
  );


  FA
  g_g127_n
  (
    .dout(g127_n),
    .din1(G1_n_spl_010),
    .din2(G3_n_spl_0001)
  );


  LA
  g_g128_p
  (
    .dout(g128_p),
    .din1(G4_p_spl_00000),
    .din2(g127_p)
  );


  FA
  g_g128_n
  (
    .dout(g128_n),
    .din1(G4_n_spl_00000),
    .din2(g127_n)
  );


  LA
  g_g129_p
  (
    .dout(g129_p),
    .din1(g126_n_spl_),
    .din2(g128_n)
  );


  FA
  g_g129_n
  (
    .dout(g129_n),
    .din1(g126_p_spl_),
    .din2(g128_p)
  );


  LA
  g_g130_p
  (
    .dout(g130_p),
    .din1(G3_p_spl_0001),
    .din2(g73_p_spl_0)
  );


  FA
  g_g130_n
  (
    .dout(g130_n),
    .din1(G3_n_spl_0010),
    .din2(g73_n_spl_0)
  );


  LA
  g_g131_p
  (
    .dout(g131_p),
    .din1(g129_p_spl_000),
    .din2(g130_n_spl_00)
  );


  FA
  g_g131_n
  (
    .dout(g131_n),
    .din1(g129_n_spl_000),
    .din2(g130_p_spl_00)
  );


  LA
  g_g132_p
  (
    .dout(g132_p),
    .din1(G1_n_spl_010),
    .din2(G4_p_spl_00000)
  );


  FA
  g_g132_n
  (
    .dout(g132_n),
    .din1(G1_p_spl_01),
    .din2(G4_n_spl_00000)
  );


  LA
  g_g133_p
  (
    .dout(g133_p),
    .din1(g131_p_spl_),
    .din2(g132_n)
  );


  FA
  g_g133_n
  (
    .dout(g133_n),
    .din1(g131_n_spl_),
    .din2(g132_p)
  );


  LA
  g_g134_p
  (
    .dout(g134_p),
    .din1(G3_p_spl_001),
    .din2(g129_n_spl_000)
  );


  FA
  g_g134_n
  (
    .dout(g134_n),
    .din1(G3_n_spl_0010),
    .din2(g129_p_spl_000)
  );


  LA
  g_g135_p
  (
    .dout(g135_p),
    .din1(g133_n_spl_0),
    .din2(g134_n_spl_0)
  );


  FA
  g_g135_n
  (
    .dout(g135_n),
    .din1(g133_p_spl_0),
    .din2(g134_p_spl_0)
  );


  LA
  g_g136_p
  (
    .dout(g136_p),
    .din1(G14_p_spl_001),
    .din2(g135_n)
  );


  FA
  g_g136_n
  (
    .dout(g136_n),
    .din1(G14_n_spl_001),
    .din2(g135_p)
  );


  LA
  g_g137_p
  (
    .dout(g137_p),
    .din1(G3_n_spl_001),
    .din2(G4_p_spl_00001)
  );


  FA
  g_g137_n
  (
    .dout(g137_n),
    .din1(G3_p_spl_001),
    .din2(G4_n_spl_00001)
  );


  LA
  g_g138_p
  (
    .dout(g138_p),
    .din1(G3_n_spl_010),
    .din2(g137_n_spl_000)
  );


  FA
  g_g138_n
  (
    .dout(g138_n),
    .din1(G3_p_spl_010),
    .din2(g137_p_spl_000)
  );


  LA
  g_g139_p
  (
    .dout(g139_p),
    .din1(G12_n_spl_001),
    .din2(g138_p_spl_00)
  );


  FA
  g_g139_n
  (
    .dout(g139_n),
    .din1(G12_p_spl_010),
    .din2(g138_n_spl_00)
  );


  LA
  g_g140_p
  (
    .dout(g140_p),
    .din1(G39_p_spl_000),
    .din2(g137_p_spl_000)
  );


  FA
  g_g140_n
  (
    .dout(g140_n),
    .din1(G39_n_spl_000),
    .din2(g137_n_spl_000)
  );


  LA
  g_g141_p
  (
    .dout(g141_p),
    .din1(g139_n),
    .din2(g140_n)
  );


  FA
  g_g141_n
  (
    .dout(g141_n),
    .din1(g139_p),
    .din2(g140_p)
  );


  LA
  g_g142_p
  (
    .dout(g142_p),
    .din1(g129_n_spl_001),
    .din2(g141_n)
  );


  FA
  g_g142_n
  (
    .dout(g142_n),
    .din1(g129_p_spl_001),
    .din2(g141_p)
  );


  LA
  g_g143_p
  (
    .dout(g143_p),
    .din1(G14_n_spl_001),
    .din2(g130_p_spl_00)
  );


  FA
  g_g143_n
  (
    .dout(g143_n),
    .din1(G14_p_spl_010),
    .din2(g130_n_spl_00)
  );


  LA
  g_g144_p
  (
    .dout(g144_p),
    .din1(g142_n),
    .din2(g143_n)
  );


  FA
  g_g144_n
  (
    .dout(g144_n),
    .din1(g142_p),
    .din2(g143_p)
  );


  LA
  g_g145_p
  (
    .dout(g145_p),
    .din1(g136_n),
    .din2(g144_p)
  );


  FA
  g_g145_n
  (
    .dout(g145_n),
    .din1(g136_p),
    .din2(g144_n)
  );


  LA
  g_g146_p
  (
    .dout(g146_p),
    .din1(G4_p_spl_00001),
    .din2(G5_p_spl_00)
  );


  FA
  g_g146_n
  (
    .dout(g146_n),
    .din1(G4_n_spl_00001),
    .din2(G5_n_spl_00)
  );


  LA
  g_g147_p
  (
    .dout(g147_p),
    .din1(g126_p_spl_),
    .din2(g146_n_spl_)
  );


  FA
  g_g147_n
  (
    .dout(g147_n),
    .din1(g126_n_spl_),
    .din2(g146_p_spl_)
  );


  LA
  g_g148_p
  (
    .dout(g148_p),
    .din1(G38_p),
    .din2(g147_n_spl_000)
  );


  FA
  g_g148_n
  (
    .dout(g148_n),
    .din1(G38_n),
    .din2(g147_p_spl_000)
  );


  LA
  g_g149_p
  (
    .dout(g149_p),
    .din1(G1_n_spl_01),
    .din2(G6_n_spl_00)
  );


  FA
  g_g149_n
  (
    .dout(g149_n),
    .din1(G1_p_spl_10),
    .din2(G6_p_spl_00)
  );


  LA
  g_g150_p
  (
    .dout(g150_p),
    .din1(G5_n_spl_00),
    .din2(g149_p_spl_0)
  );


  FA
  g_g150_n
  (
    .dout(g150_n),
    .din1(G5_p_spl_00),
    .din2(g149_n_spl_0)
  );


  LA
  g_g151_p
  (
    .dout(g151_p),
    .din1(g148_p_spl_0),
    .din2(g150_p_spl_0)
  );


  FA
  g_g151_n
  (
    .dout(g151_n),
    .din1(g148_n_spl_0),
    .din2(g150_n_spl_0)
  );


  LA
  g_g152_p
  (
    .dout(g152_p),
    .din1(G37_p_spl_),
    .din2(g150_n_spl_0)
  );


  FA
  g_g152_n
  (
    .dout(g152_n),
    .din1(G37_n_spl_1),
    .din2(g150_p_spl_0)
  );


  LA
  g_g153_p
  (
    .dout(g153_p),
    .din1(G4_n_spl_00010),
    .din2(G49_n)
  );


  FA
  g_g153_n
  (
    .dout(g153_n),
    .din1(G4_p_spl_00010),
    .din2(G49_p)
  );


  LA
  g_g154_p
  (
    .dout(g154_p),
    .din1(G35_p_spl_0),
    .din2(g153_p_spl_00)
  );


  FA
  g_g154_n
  (
    .dout(g154_n),
    .din1(G35_n_spl_10),
    .din2(g153_n_spl_00)
  );


  LA
  g_g155_p
  (
    .dout(g155_p),
    .din1(g152_n),
    .din2(g154_n)
  );


  FA
  g_g155_n
  (
    .dout(g155_n),
    .din1(g152_p),
    .din2(g154_p)
  );


  LA
  g_g156_p
  (
    .dout(g156_p),
    .din1(G4_n_spl_00010),
    .din2(G41_n_spl_00)
  );


  FA
  g_g156_n
  (
    .dout(g156_n),
    .din1(G4_p_spl_00010),
    .din2(G41_p_spl_00)
  );


  LA
  g_g157_p
  (
    .dout(g157_p),
    .din1(G4_p_spl_00011),
    .din2(G36_n_spl_1)
  );


  FA
  g_g157_n
  (
    .dout(g157_n),
    .din1(G4_n_spl_00011),
    .din2(G36_p_spl_1)
  );


  LA
  g_g158_p
  (
    .dout(g158_p),
    .din1(g156_n),
    .din2(g157_n)
  );


  FA
  g_g158_n
  (
    .dout(g158_n),
    .din1(g156_p),
    .din2(g157_p)
  );


  LA
  g_g159_p
  (
    .dout(g159_p),
    .din1(g155_p),
    .din2(g158_n)
  );


  FA
  g_g159_n
  (
    .dout(g159_n),
    .din1(g155_n),
    .din2(g158_p)
  );


  LA
  g_g160_p
  (
    .dout(g160_p),
    .din1(g147_n_spl_000),
    .din2(g159_n)
  );


  FA
  g_g160_n
  (
    .dout(g160_n),
    .din1(g147_p_spl_000),
    .din2(g159_p)
  );


  LA
  g_g161_p
  (
    .dout(g161_p),
    .din1(g151_n_spl_0),
    .din2(g160_n)
  );


  FA
  g_g161_n
  (
    .dout(g161_n),
    .din1(g151_p_spl_0),
    .din2(g160_p)
  );


  LA
  g_g162_p
  (
    .dout(g162_p),
    .din1(G25_n_spl_),
    .din2(G26_n_spl_0)
  );


  FA
  g_g162_n
  (
    .dout(g162_n),
    .din1(G25_p_spl_),
    .din2(G26_p_spl_0)
  );


  LA
  g_g163_p
  (
    .dout(g163_p),
    .din1(g161_p_spl_0),
    .din2(g162_n_spl_000)
  );


  FA
  g_g163_n
  (
    .dout(g163_n),
    .din1(g161_n_spl_0),
    .din2(g162_p_spl_000)
  );


  LA
  g_g164_p
  (
    .dout(g164_p),
    .din1(g145_p_spl_0),
    .din2(g163_n)
  );


  FA
  g_g164_n
  (
    .dout(g164_n),
    .din1(g145_n_spl_0),
    .din2(g163_p)
  );


  LA
  g_g165_p
  (
    .dout(g165_p),
    .din1(G23_n_spl_),
    .din2(G24_n_spl_0)
  );


  FA
  g_g165_n
  (
    .dout(g165_n),
    .din1(G23_p_spl_),
    .din2(G24_p_spl_0)
  );


  LA
  g_g166_p
  (
    .dout(g166_p),
    .din1(g145_n_spl_0),
    .din2(g161_p_spl_0)
  );


  FA
  g_g166_n
  (
    .dout(g166_n),
    .din1(g145_p_spl_0),
    .din2(g161_n_spl_0)
  );


  LA
  g_g167_p
  (
    .dout(g167_p),
    .din1(g165_n_spl_00),
    .din2(g166_p)
  );


  FA
  g_g167_n
  (
    .dout(g167_n),
    .din1(g165_p_spl_00),
    .din2(g166_n)
  );


  LA
  g_g168_p
  (
    .dout(g168_p),
    .din1(g164_n),
    .din2(g167_n_spl_0)
  );


  FA
  g_g168_n
  (
    .dout(g168_n),
    .din1(g164_p),
    .din2(g167_p_spl_0)
  );


  LA
  g_g169_p
  (
    .dout(g169_p),
    .din1(g130_n_spl_01),
    .din2(g134_n_spl_0)
  );


  FA
  g_g169_n
  (
    .dout(g169_n),
    .din1(g130_p_spl_01),
    .din2(g134_p_spl_0)
  );


  LA
  g_g170_p
  (
    .dout(g170_p),
    .din1(G13_n_spl_001),
    .din2(g169_n_spl_)
  );


  FA
  g_g170_n
  (
    .dout(g170_n),
    .din1(G13_p_spl_010),
    .din2(g169_p_spl_)
  );


  LA
  g_g171_p
  (
    .dout(g171_p),
    .din1(G11_n_spl_001),
    .din2(g138_p_spl_00)
  );


  FA
  g_g171_n
  (
    .dout(g171_n),
    .din1(G11_p_spl_010),
    .din2(g138_n_spl_00)
  );


  LA
  g_g172_p
  (
    .dout(g172_p),
    .din1(G14_p_spl_010),
    .din2(g137_p_spl_00)
  );


  FA
  g_g172_n
  (
    .dout(g172_n),
    .din1(G14_n_spl_010),
    .din2(g137_n_spl_00)
  );


  LA
  g_g173_p
  (
    .dout(g173_p),
    .din1(g171_n),
    .din2(g172_n)
  );


  FA
  g_g173_n
  (
    .dout(g173_n),
    .din1(g171_p),
    .din2(g172_p)
  );


  LA
  g_g174_p
  (
    .dout(g174_p),
    .din1(g129_n_spl_001),
    .din2(g173_n)
  );


  FA
  g_g174_n
  (
    .dout(g174_n),
    .din1(g129_p_spl_001),
    .din2(g173_p)
  );


  LA
  g_g175_p
  (
    .dout(g175_p),
    .din1(G13_p_spl_010),
    .din2(g133_p_spl_0)
  );


  FA
  g_g175_n
  (
    .dout(g175_n),
    .din1(G13_n_spl_010),
    .din2(g133_n_spl_0)
  );


  LA
  g_g176_p
  (
    .dout(g176_p),
    .din1(g174_n),
    .din2(g175_n)
  );


  FA
  g_g176_n
  (
    .dout(g176_n),
    .din1(g174_p),
    .din2(g175_p)
  );


  LA
  g_g177_p
  (
    .dout(g177_p),
    .din1(g170_n),
    .din2(g176_p)
  );


  FA
  g_g177_n
  (
    .dout(g177_n),
    .din1(g170_p),
    .din2(g176_n)
  );


  LA
  g_g178_p
  (
    .dout(g178_p),
    .din1(G36_p_spl_1),
    .din2(g150_n_spl_1)
  );


  FA
  g_g178_n
  (
    .dout(g178_n),
    .din1(G36_n_spl_1),
    .din2(g150_p_spl_1)
  );


  LA
  g_g179_p
  (
    .dout(g179_p),
    .din1(G34_p_spl_0),
    .din2(g153_p_spl_00)
  );


  FA
  g_g179_n
  (
    .dout(g179_n),
    .din1(G34_n_spl_10),
    .din2(g153_n_spl_00)
  );


  LA
  g_g180_p
  (
    .dout(g180_p),
    .din1(g178_n),
    .din2(g179_n)
  );


  FA
  g_g180_n
  (
    .dout(g180_n),
    .din1(g178_p),
    .din2(g179_p)
  );


  LA
  g_g181_p
  (
    .dout(g181_p),
    .din1(G4_n_spl_00011),
    .din2(G40_n_spl_00)
  );


  FA
  g_g181_n
  (
    .dout(g181_n),
    .din1(G4_p_spl_00011),
    .din2(G40_p_spl_00)
  );


  LA
  g_g182_p
  (
    .dout(g182_p),
    .din1(G4_p_spl_0010),
    .din2(G35_n_spl_10)
  );


  FA
  g_g182_n
  (
    .dout(g182_n),
    .din1(G4_n_spl_0010),
    .din2(G35_p_spl_1)
  );


  LA
  g_g183_p
  (
    .dout(g183_p),
    .din1(g181_n),
    .din2(g182_n)
  );


  FA
  g_g183_n
  (
    .dout(g183_n),
    .din1(g181_p),
    .din2(g182_p)
  );


  LA
  g_g184_p
  (
    .dout(g184_p),
    .din1(g180_p),
    .din2(g183_n)
  );


  FA
  g_g184_n
  (
    .dout(g184_n),
    .din1(g180_n),
    .din2(g183_p)
  );


  LA
  g_g185_p
  (
    .dout(g185_p),
    .din1(g147_n_spl_00),
    .din2(g184_n)
  );


  FA
  g_g185_n
  (
    .dout(g185_n),
    .din1(g147_p_spl_00),
    .din2(g184_p)
  );


  LA
  g_g186_p
  (
    .dout(g186_p),
    .din1(g151_n_spl_0),
    .din2(g185_n)
  );


  FA
  g_g186_n
  (
    .dout(g186_n),
    .din1(g151_p_spl_0),
    .din2(g185_p)
  );


  LA
  g_g187_p
  (
    .dout(g187_p),
    .din1(g162_n_spl_000),
    .din2(g186_p_spl_0)
  );


  FA
  g_g187_n
  (
    .dout(g187_n),
    .din1(g162_p_spl_000),
    .din2(g186_n_spl_0)
  );


  LA
  g_g188_p
  (
    .dout(g188_p),
    .din1(g177_p_spl_0),
    .din2(g187_n)
  );


  FA
  g_g188_n
  (
    .dout(g188_n),
    .din1(g177_n_spl_0),
    .din2(g187_p)
  );


  LA
  g_g189_p
  (
    .dout(g189_p),
    .din1(g165_n_spl_00),
    .din2(g177_n_spl_0)
  );


  FA
  g_g189_n
  (
    .dout(g189_n),
    .din1(g165_p_spl_00),
    .din2(g177_p_spl_0)
  );


  LA
  g_g190_p
  (
    .dout(g190_p),
    .din1(g186_p_spl_0),
    .din2(g189_p)
  );


  FA
  g_g190_n
  (
    .dout(g190_n),
    .din1(g186_n_spl_0),
    .din2(g189_n)
  );


  LA
  g_g191_p
  (
    .dout(g191_p),
    .din1(g188_n),
    .din2(g190_n_spl_0)
  );


  FA
  g_g191_n
  (
    .dout(g191_n),
    .din1(g188_p),
    .din2(g190_p_spl_0)
  );


  LA
  g_g192_p
  (
    .dout(g192_p),
    .din1(G11_p_spl_010),
    .din2(g133_n_spl_1)
  );


  FA
  g_g192_n
  (
    .dout(g192_n),
    .din1(G11_n_spl_010),
    .din2(g133_p_spl_1)
  );


  LA
  g_g193_p
  (
    .dout(g193_p),
    .din1(G11_n_spl_010),
    .din2(g130_n_spl_01)
  );


  FA
  g_g193_n
  (
    .dout(g193_n),
    .din1(G11_p_spl_011),
    .din2(g130_p_spl_01)
  );


  LA
  g_g194_p
  (
    .dout(g194_p),
    .din1(g192_n),
    .din2(g193_n)
  );


  FA
  g_g194_n
  (
    .dout(g194_n),
    .din1(g192_p),
    .din2(g193_p)
  );


  LA
  g_g195_p
  (
    .dout(g195_p),
    .din1(G12_n_spl_010),
    .din2(g137_p_spl_01)
  );


  FA
  g_g195_n
  (
    .dout(g195_n),
    .din1(G12_p_spl_010),
    .din2(g137_n_spl_01)
  );


  LA
  g_g196_p
  (
    .dout(g196_p),
    .din1(G13_n_spl_010),
    .din2(g106_p_spl_)
  );


  FA
  g_g196_n
  (
    .dout(g196_n),
    .din1(G13_p_spl_011),
    .din2(g106_n_spl_)
  );


  LA
  g_g197_p
  (
    .dout(g197_p),
    .din1(G3_p_spl_010),
    .din2(g196_n_spl_)
  );


  FA
  g_g197_n
  (
    .dout(g197_n),
    .din1(G3_n_spl_010),
    .din2(g196_p_spl_)
  );


  LA
  g_g198_p
  (
    .dout(g198_p),
    .din1(G9_n_spl_010),
    .din2(g138_p_spl_01)
  );


  FA
  g_g198_n
  (
    .dout(g198_n),
    .din1(G9_p_spl_010),
    .din2(g138_n_spl_01)
  );


  LA
  g_g199_p
  (
    .dout(g199_p),
    .din1(g197_n),
    .din2(g198_n)
  );


  FA
  g_g199_n
  (
    .dout(g199_n),
    .din1(g197_p),
    .din2(g198_p)
  );


  LA
  g_g200_p
  (
    .dout(g200_p),
    .din1(g195_n),
    .din2(g199_p)
  );


  FA
  g_g200_n
  (
    .dout(g200_n),
    .din1(g195_p),
    .din2(g199_n)
  );


  LA
  g_g201_p
  (
    .dout(g201_p),
    .din1(g129_n_spl_01),
    .din2(g200_n)
  );


  FA
  g_g201_n
  (
    .dout(g201_n),
    .din1(g129_p_spl_01),
    .din2(g200_p)
  );


  LA
  g_g202_p
  (
    .dout(g202_p),
    .din1(g194_n),
    .din2(g201_n)
  );


  FA
  g_g202_n
  (
    .dout(g202_n),
    .din1(g194_p),
    .din2(g201_p)
  );


  LA
  g_g203_p
  (
    .dout(g203_p),
    .din1(g148_p_spl_0),
    .din2(g149_p_spl_0)
  );


  FA
  g_g203_n
  (
    .dout(g203_n),
    .din1(g148_n_spl_0),
    .din2(g149_n_spl_0)
  );


  LA
  g_g204_p
  (
    .dout(g204_p),
    .din1(G4_p_spl_0010),
    .din2(G33_p_spl_0)
  );


  FA
  g_g204_n
  (
    .dout(g204_n),
    .din1(G4_n_spl_0010),
    .din2(G33_n_spl_01)
  );


  LA
  g_g205_p
  (
    .dout(g205_p),
    .din1(G4_n_spl_0011),
    .din2(G14_p_spl_011)
  );


  FA
  g_g205_n
  (
    .dout(g205_n),
    .din1(G4_p_spl_0011),
    .din2(G14_n_spl_010)
  );


  LA
  g_g206_p
  (
    .dout(g206_p),
    .din1(g204_n),
    .din2(g205_n)
  );


  FA
  g_g206_n
  (
    .dout(g206_n),
    .din1(g204_p),
    .din2(g205_p)
  );


  LA
  g_g207_p
  (
    .dout(g207_p),
    .din1(G34_p_spl_1),
    .din2(g149_n_spl_)
  );


  FA
  g_g207_n
  (
    .dout(g207_n),
    .din1(G34_n_spl_10),
    .din2(g149_p_spl_)
  );


  LA
  g_g208_p
  (
    .dout(g208_p),
    .din1(G32_p_spl_0),
    .din2(g153_p_spl_01)
  );


  FA
  g_g208_n
  (
    .dout(g208_n),
    .din1(G32_n_spl_01),
    .din2(g153_n_spl_01)
  );


  LA
  g_g209_p
  (
    .dout(g209_p),
    .din1(g207_n),
    .din2(g208_n)
  );


  FA
  g_g209_n
  (
    .dout(g209_n),
    .din1(g207_p),
    .din2(g208_p)
  );


  LA
  g_g210_p
  (
    .dout(g210_p),
    .din1(g206_p),
    .din2(g209_p)
  );


  FA
  g_g210_n
  (
    .dout(g210_n),
    .din1(g206_n),
    .din2(g209_n)
  );


  LA
  g_g211_p
  (
    .dout(g211_p),
    .din1(g147_n_spl_01),
    .din2(g210_n)
  );


  FA
  g_g211_n
  (
    .dout(g211_n),
    .din1(g147_p_spl_01),
    .din2(g210_p)
  );


  LA
  g_g212_p
  (
    .dout(g212_p),
    .din1(g203_n),
    .din2(g211_n)
  );


  FA
  g_g212_n
  (
    .dout(g212_n),
    .din1(g203_p),
    .din2(g211_p)
  );


  LA
  g_g213_p
  (
    .dout(g213_p),
    .din1(g162_n_spl_00),
    .din2(g212_p_spl_0)
  );


  FA
  g_g213_n
  (
    .dout(g213_n),
    .din1(g162_p_spl_00),
    .din2(g212_n_spl_0)
  );


  LA
  g_g214_p
  (
    .dout(g214_p),
    .din1(g202_p_spl_0),
    .din2(g213_n)
  );


  FA
  g_g214_n
  (
    .dout(g214_n),
    .din1(g202_n_spl_0),
    .din2(g213_p)
  );


  LA
  g_g215_p
  (
    .dout(g215_p),
    .din1(g165_n_spl_01),
    .din2(g202_n_spl_0)
  );


  FA
  g_g215_n
  (
    .dout(g215_n),
    .din1(g165_p_spl_01),
    .din2(g202_p_spl_0)
  );


  LA
  g_g216_p
  (
    .dout(g216_p),
    .din1(g212_p_spl_0),
    .din2(g215_p)
  );


  FA
  g_g216_n
  (
    .dout(g216_n),
    .din1(g212_n_spl_0),
    .din2(g215_n)
  );


  LA
  g_g217_p
  (
    .dout(g217_p),
    .din1(g214_n),
    .din2(g216_n_spl_)
  );


  FA
  g_g217_n
  (
    .dout(g217_n),
    .din1(g214_p),
    .din2(g216_p_spl_)
  );


  LA
  g_g218_p
  (
    .dout(g218_p),
    .din1(G12_p_spl_011),
    .din2(g133_n_spl_1)
  );


  FA
  g_g218_n
  (
    .dout(g218_n),
    .din1(G12_n_spl_010),
    .din2(g133_p_spl_1)
  );


  LA
  g_g219_p
  (
    .dout(g219_p),
    .din1(G12_n_spl_011),
    .din2(g130_n_spl_10)
  );


  FA
  g_g219_n
  (
    .dout(g219_n),
    .din1(G12_p_spl_011),
    .din2(g130_p_spl_10)
  );


  LA
  g_g220_p
  (
    .dout(g220_p),
    .din1(g218_n),
    .din2(g219_n)
  );


  FA
  g_g220_n
  (
    .dout(g220_n),
    .din1(g218_p),
    .din2(g219_p)
  );


  LA
  g_g221_p
  (
    .dout(g221_p),
    .din1(G13_p_spl_011),
    .din2(g137_p_spl_01)
  );


  FA
  g_g221_n
  (
    .dout(g221_n),
    .din1(G13_n_spl_011),
    .din2(g137_n_spl_01)
  );


  LA
  g_g222_p
  (
    .dout(g222_p),
    .din1(G12_p_spl_100),
    .din2(G13_p_spl_100)
  );


  FA
  g_g222_n
  (
    .dout(g222_n),
    .din1(G12_n_spl_011),
    .din2(G13_n_spl_011)
  );


  LA
  g_g223_p
  (
    .dout(g223_p),
    .din1(g54_n_spl_),
    .din2(g222_n)
  );


  FA
  g_g223_n
  (
    .dout(g223_n),
    .din1(g54_p_spl_),
    .din2(g222_p)
  );


  LA
  g_g224_p
  (
    .dout(g224_p),
    .din1(G3_p_spl_011),
    .din2(g223_p)
  );


  FA
  g_g224_n
  (
    .dout(g224_n),
    .din1(G3_n_spl_011),
    .din2(g223_n_spl_)
  );


  LA
  g_g225_p
  (
    .dout(g225_p),
    .din1(G10_p_spl_001),
    .din2(g138_p_spl_01)
  );


  FA
  g_g225_n
  (
    .dout(g225_n),
    .din1(G10_n_spl_001),
    .din2(g138_n_spl_01)
  );


  LA
  g_g226_p
  (
    .dout(g226_p),
    .din1(g224_n),
    .din2(g225_n)
  );


  FA
  g_g226_n
  (
    .dout(g226_n),
    .din1(g224_p),
    .din2(g225_p)
  );


  LA
  g_g227_p
  (
    .dout(g227_p),
    .din1(g221_n),
    .din2(g226_p)
  );


  FA
  g_g227_n
  (
    .dout(g227_n),
    .din1(g221_p),
    .din2(g226_n)
  );


  LA
  g_g228_p
  (
    .dout(g228_p),
    .din1(g129_n_spl_01),
    .din2(g227_n)
  );


  FA
  g_g228_n
  (
    .dout(g228_n),
    .din1(g129_p_spl_01),
    .din2(g227_p)
  );


  LA
  g_g229_p
  (
    .dout(g229_p),
    .din1(g220_n),
    .din2(g228_n)
  );


  FA
  g_g229_n
  (
    .dout(g229_n),
    .din1(g220_p),
    .din2(g228_p)
  );


  LA
  g_g230_p
  (
    .dout(g230_p),
    .din1(G35_p_spl_1),
    .din2(g150_n_spl_1)
  );


  FA
  g_g230_n
  (
    .dout(g230_n),
    .din1(G35_n_spl_1),
    .din2(g150_p_spl_1)
  );


  LA
  g_g231_p
  (
    .dout(g231_p),
    .din1(G33_p_spl_1),
    .din2(g153_p_spl_01)
  );


  FA
  g_g231_n
  (
    .dout(g231_n),
    .din1(G33_n_spl_1),
    .din2(g153_n_spl_01)
  );


  LA
  g_g232_p
  (
    .dout(g232_p),
    .din1(g230_n),
    .din2(g231_n)
  );


  FA
  g_g232_n
  (
    .dout(g232_n),
    .din1(g230_p),
    .din2(g231_p)
  );


  LA
  g_g233_p
  (
    .dout(g233_p),
    .din1(G4_n_spl_0011),
    .din2(G39_n_spl_000)
  );


  FA
  g_g233_n
  (
    .dout(g233_n),
    .din1(G4_p_spl_0011),
    .din2(G39_p_spl_000)
  );


  LA
  g_g234_p
  (
    .dout(g234_p),
    .din1(G4_p_spl_0100),
    .din2(G34_n_spl_1)
  );


  FA
  g_g234_n
  (
    .dout(g234_n),
    .din1(G4_n_spl_0100),
    .din2(G34_p_spl_1)
  );


  LA
  g_g235_p
  (
    .dout(g235_p),
    .din1(g233_n),
    .din2(g234_n)
  );


  FA
  g_g235_n
  (
    .dout(g235_n),
    .din1(g233_p),
    .din2(g234_p)
  );


  LA
  g_g236_p
  (
    .dout(g236_p),
    .din1(g232_p),
    .din2(g235_n)
  );


  FA
  g_g236_n
  (
    .dout(g236_n),
    .din1(g232_n),
    .din2(g235_p)
  );


  LA
  g_g237_p
  (
    .dout(g237_p),
    .din1(g147_n_spl_01),
    .din2(g236_n)
  );


  FA
  g_g237_n
  (
    .dout(g237_n),
    .din1(g147_p_spl_01),
    .din2(g236_p)
  );


  LA
  g_g238_p
  (
    .dout(g238_p),
    .din1(g151_n_spl_),
    .din2(g237_n)
  );


  FA
  g_g238_n
  (
    .dout(g238_n),
    .din1(g151_p_spl_),
    .din2(g237_p)
  );


  LA
  g_g239_p
  (
    .dout(g239_p),
    .din1(g162_n_spl_01),
    .din2(g238_p_spl_0)
  );


  FA
  g_g239_n
  (
    .dout(g239_n),
    .din1(g162_p_spl_01),
    .din2(g238_n_spl_0)
  );


  LA
  g_g240_p
  (
    .dout(g240_p),
    .din1(g229_p_spl_0),
    .din2(g239_n)
  );


  FA
  g_g240_n
  (
    .dout(g240_n),
    .din1(g229_n_spl_0),
    .din2(g239_p)
  );


  LA
  g_g241_p
  (
    .dout(g241_p),
    .din1(g165_n_spl_01),
    .din2(g229_n_spl_0)
  );


  FA
  g_g241_n
  (
    .dout(g241_n),
    .din1(g165_p_spl_01),
    .din2(g229_p_spl_0)
  );


  LA
  g_g242_p
  (
    .dout(g242_p),
    .din1(g238_p_spl_0),
    .din2(g241_p)
  );


  FA
  g_g242_n
  (
    .dout(g242_n),
    .din1(g238_n_spl_0),
    .din2(g241_n)
  );


  LA
  g_g243_p
  (
    .dout(g243_p),
    .din1(g240_n),
    .din2(g242_n_spl_0)
  );


  FA
  g_g243_n
  (
    .dout(g243_n),
    .din1(g240_p),
    .din2(g242_p_spl_0)
  );


  LA
  g_g244_p
  (
    .dout(g244_p),
    .din1(g217_p_spl_0),
    .din2(g243_p_spl_0)
  );


  FA
  g_g244_n
  (
    .dout(g244_n),
    .din1(g217_n_spl_0),
    .din2(g243_n_spl_0)
  );


  LA
  g_g245_p
  (
    .dout(g245_p),
    .din1(g191_p_spl_0),
    .din2(g244_p_spl_)
  );


  FA
  g_g245_n
  (
    .dout(g245_n),
    .din1(g191_n_spl_0),
    .din2(g244_n_spl_)
  );


  LA
  g_g246_p
  (
    .dout(g246_p),
    .din1(g168_p_spl_0),
    .din2(g245_p_spl_)
  );


  FA
  g_g246_n
  (
    .dout(g246_n),
    .din1(g168_n_spl_0),
    .din2(g245_n_spl_)
  );


  LA
  g_g247_p
  (
    .dout(g247_p),
    .din1(G1_n_spl_10),
    .din2(G3_p_spl_011)
  );


  FA
  g_g247_n
  (
    .dout(g247_n),
    .din1(G1_p_spl_10),
    .din2(G3_n_spl_011)
  );


  LA
  g_g248_p
  (
    .dout(g248_p),
    .din1(g131_p_spl_),
    .din2(g247_n)
  );


  FA
  g_g248_n
  (
    .dout(g248_n),
    .din1(g131_n_spl_),
    .din2(g247_p)
  );


  LA
  g_g249_p
  (
    .dout(g249_p),
    .din1(g134_n_spl_),
    .din2(g248_n_spl_0)
  );


  FA
  g_g249_n
  (
    .dout(g249_n),
    .din1(g134_p_spl_),
    .din2(g248_p_spl_0)
  );


  LA
  g_g250_p
  (
    .dout(g250_p),
    .din1(G10_p_spl_010),
    .din2(g249_n)
  );


  FA
  g_g250_n
  (
    .dout(g250_n),
    .din1(G10_n_spl_010),
    .din2(g249_p)
  );


  LA
  g_g251_p
  (
    .dout(g251_p),
    .din1(G8_n_spl_001),
    .din2(g138_p_spl_10)
  );


  FA
  g_g251_n
  (
    .dout(g251_n),
    .din1(G8_p_spl_010),
    .din2(g138_n_spl_10)
  );


  LA
  g_g252_p
  (
    .dout(g252_p),
    .din1(G11_n_spl_011),
    .din2(g137_p_spl_10)
  );


  FA
  g_g252_n
  (
    .dout(g252_n),
    .din1(G11_p_spl_011),
    .din2(g137_n_spl_10)
  );


  LA
  g_g253_p
  (
    .dout(g253_p),
    .din1(g251_n),
    .din2(g252_n)
  );


  FA
  g_g253_n
  (
    .dout(g253_n),
    .din1(g251_p),
    .din2(g252_p)
  );


  LA
  g_g254_p
  (
    .dout(g254_p),
    .din1(g129_n_spl_10),
    .din2(g253_n)
  );


  FA
  g_g254_n
  (
    .dout(g254_n),
    .din1(g129_p_spl_10),
    .din2(g253_p)
  );


  LA
  g_g255_p
  (
    .dout(g255_p),
    .din1(G10_n_spl_010),
    .din2(g130_p_spl_10)
  );


  FA
  g_g255_n
  (
    .dout(g255_n),
    .din1(G10_p_spl_010),
    .din2(g130_n_spl_10)
  );


  LA
  g_g256_p
  (
    .dout(g256_p),
    .din1(g254_n),
    .din2(g255_n)
  );


  FA
  g_g256_n
  (
    .dout(g256_n),
    .din1(g254_p),
    .din2(g255_p)
  );


  LA
  g_g257_p
  (
    .dout(g257_p),
    .din1(g250_n),
    .din2(g256_p)
  );


  FA
  g_g257_n
  (
    .dout(g257_n),
    .din1(g250_p),
    .din2(g256_n)
  );


  LA
  g_g258_p
  (
    .dout(g258_p),
    .din1(G5_n_spl_01),
    .din2(G6_n_spl_00)
  );


  FA
  g_g258_n
  (
    .dout(g258_n),
    .din1(G5_p_spl_01),
    .din2(G6_p_spl_00)
  );


  LA
  g_g259_p
  (
    .dout(g259_p),
    .din1(G1_n_spl_10),
    .din2(g258_n)
  );


  FA
  g_g259_n
  (
    .dout(g259_n),
    .din1(G1_p_spl_11),
    .din2(g258_p)
  );


  LA
  g_g260_p
  (
    .dout(g260_p),
    .din1(g148_p_spl_),
    .din2(g259_p_spl_00)
  );


  FA
  g_g260_n
  (
    .dout(g260_n),
    .din1(g148_n_spl_),
    .din2(g259_n_spl_00)
  );


  LA
  g_g261_p
  (
    .dout(g261_p),
    .din1(G33_p_spl_1),
    .din2(g259_n_spl_00)
  );


  FA
  g_g261_n
  (
    .dout(g261_n),
    .din1(G33_n_spl_1),
    .din2(g259_p_spl_00)
  );


  LA
  g_g262_p
  (
    .dout(g262_p),
    .din1(G31_p_spl_0),
    .din2(g153_p_spl_10)
  );


  FA
  g_g262_n
  (
    .dout(g262_n),
    .din1(G31_n_spl_01),
    .din2(g153_n_spl_10)
  );


  LA
  g_g263_p
  (
    .dout(g263_p),
    .din1(g261_n),
    .din2(g262_n)
  );


  FA
  g_g263_n
  (
    .dout(g263_n),
    .din1(g261_p),
    .din2(g262_p)
  );


  LA
  g_g264_p
  (
    .dout(g264_p),
    .din1(G4_n_spl_0100),
    .din2(G13_n_spl_100)
  );


  FA
  g_g264_n
  (
    .dout(g264_n),
    .din1(G4_p_spl_0100),
    .din2(G13_p_spl_100)
  );


  LA
  g_g265_p
  (
    .dout(g265_p),
    .din1(G4_p_spl_0101),
    .din2(G32_n_spl_1)
  );


  FA
  g_g265_n
  (
    .dout(g265_n),
    .din1(G4_n_spl_0101),
    .din2(G32_p_spl_1)
  );


  LA
  g_g266_p
  (
    .dout(g266_p),
    .din1(g264_n),
    .din2(g265_n)
  );


  FA
  g_g266_n
  (
    .dout(g266_n),
    .din1(g264_p),
    .din2(g265_p)
  );


  LA
  g_g267_p
  (
    .dout(g267_p),
    .din1(g263_p),
    .din2(g266_n)
  );


  FA
  g_g267_n
  (
    .dout(g267_n),
    .din1(g263_n),
    .din2(g266_p)
  );


  LA
  g_g268_p
  (
    .dout(g268_p),
    .din1(g147_n_spl_10),
    .din2(g267_n)
  );


  FA
  g_g268_n
  (
    .dout(g268_n),
    .din1(g147_p_spl_10),
    .din2(g267_p)
  );


  LA
  g_g269_p
  (
    .dout(g269_p),
    .din1(g260_n_spl_0),
    .din2(g268_n)
  );


  FA
  g_g269_n
  (
    .dout(g269_n),
    .din1(g260_p_spl_0),
    .din2(g268_p)
  );


  LA
  g_g270_p
  (
    .dout(g270_p),
    .din1(g162_n_spl_01),
    .din2(g269_p_spl_)
  );


  FA
  g_g270_n
  (
    .dout(g270_n),
    .din1(g162_p_spl_01),
    .din2(g269_n_spl_)
  );


  LA
  g_g271_p
  (
    .dout(g271_p),
    .din1(g257_p_spl_0),
    .din2(g270_n)
  );


  FA
  g_g271_n
  (
    .dout(g271_n),
    .din1(g257_n_spl_0),
    .din2(g270_p)
  );


  LA
  g_g272_p
  (
    .dout(g272_p),
    .din1(g165_n_spl_10),
    .din2(g257_n_spl_0)
  );


  FA
  g_g272_n
  (
    .dout(g272_n),
    .din1(g165_p_spl_10),
    .din2(g257_p_spl_0)
  );


  LA
  g_g273_p
  (
    .dout(g273_p),
    .din1(g269_p_spl_),
    .din2(g272_p)
  );


  FA
  g_g273_n
  (
    .dout(g273_n),
    .din1(g269_n_spl_),
    .din2(g272_n)
  );


  LA
  g_g274_p
  (
    .dout(g274_p),
    .din1(g271_n),
    .din2(g273_n_spl_0)
  );


  FA
  g_g274_n
  (
    .dout(g274_n),
    .din1(g271_p),
    .din2(g273_p_spl_0)
  );


  LA
  g_g275_p
  (
    .dout(g275_p),
    .din1(G9_n_spl_010),
    .din2(g169_n_spl_)
  );


  FA
  g_g275_n
  (
    .dout(g275_n),
    .din1(G9_p_spl_011),
    .din2(g169_p_spl_)
  );


  LA
  g_g276_p
  (
    .dout(g276_p),
    .din1(G7_p_spl_001),
    .din2(g138_p_spl_10)
  );


  FA
  g_g276_n
  (
    .dout(g276_n),
    .din1(G7_n_spl_001),
    .din2(g138_n_spl_10)
  );


  LA
  g_g277_p
  (
    .dout(g277_p),
    .din1(G10_p_spl_011),
    .din2(g137_p_spl_10)
  );


  FA
  g_g277_n
  (
    .dout(g277_n),
    .din1(G10_n_spl_011),
    .din2(g137_n_spl_10)
  );


  LA
  g_g278_p
  (
    .dout(g278_p),
    .din1(g276_n),
    .din2(g277_n)
  );


  FA
  g_g278_n
  (
    .dout(g278_n),
    .din1(g276_p),
    .din2(g277_p)
  );


  LA
  g_g279_p
  (
    .dout(g279_p),
    .din1(g129_n_spl_10),
    .din2(g278_n)
  );


  FA
  g_g279_n
  (
    .dout(g279_n),
    .din1(g129_p_spl_10),
    .din2(g278_p)
  );


  LA
  g_g280_p
  (
    .dout(g280_p),
    .din1(G9_p_spl_011),
    .din2(g248_p_spl_0)
  );


  FA
  g_g280_n
  (
    .dout(g280_n),
    .din1(G9_n_spl_011),
    .din2(g248_n_spl_0)
  );


  LA
  g_g281_p
  (
    .dout(g281_p),
    .din1(g279_n),
    .din2(g280_n)
  );


  FA
  g_g281_n
  (
    .dout(g281_n),
    .din1(g279_p),
    .din2(g280_p)
  );


  LA
  g_g282_p
  (
    .dout(g282_p),
    .din1(g275_n),
    .din2(g281_p)
  );


  FA
  g_g282_n
  (
    .dout(g282_n),
    .din1(g275_p),
    .din2(g281_n)
  );


  LA
  g_g283_p
  (
    .dout(g283_p),
    .din1(G32_p_spl_1),
    .din2(g259_n_spl_0)
  );


  FA
  g_g283_n
  (
    .dout(g283_n),
    .din1(G32_n_spl_1),
    .din2(g259_p_spl_0)
  );


  LA
  g_g284_p
  (
    .dout(g284_p),
    .din1(G30_p_spl_0),
    .din2(g153_p_spl_10)
  );


  FA
  g_g284_n
  (
    .dout(g284_n),
    .din1(G30_n_spl_01),
    .din2(g153_n_spl_10)
  );


  LA
  g_g285_p
  (
    .dout(g285_p),
    .din1(g283_n),
    .din2(g284_n)
  );


  FA
  g_g285_n
  (
    .dout(g285_n),
    .din1(g283_p),
    .din2(g284_p)
  );


  LA
  g_g286_p
  (
    .dout(g286_p),
    .din1(G4_n_spl_0101),
    .din2(G12_n_spl_100)
  );


  FA
  g_g286_n
  (
    .dout(g286_n),
    .din1(G4_p_spl_0101),
    .din2(G12_p_spl_100)
  );


  LA
  g_g287_p
  (
    .dout(g287_p),
    .din1(G4_p_spl_0110),
    .din2(G31_n_spl_1)
  );


  FA
  g_g287_n
  (
    .dout(g287_n),
    .din1(G4_n_spl_0110),
    .din2(G31_p_spl_1)
  );


  LA
  g_g288_p
  (
    .dout(g288_p),
    .din1(g286_n),
    .din2(g287_n)
  );


  FA
  g_g288_n
  (
    .dout(g288_n),
    .din1(g286_p),
    .din2(g287_p)
  );


  LA
  g_g289_p
  (
    .dout(g289_p),
    .din1(g285_p),
    .din2(g288_n)
  );


  FA
  g_g289_n
  (
    .dout(g289_n),
    .din1(g285_n),
    .din2(g288_p)
  );


  LA
  g_g290_p
  (
    .dout(g290_p),
    .din1(g147_n_spl_10),
    .din2(g289_n)
  );


  FA
  g_g290_n
  (
    .dout(g290_n),
    .din1(g147_p_spl_10),
    .din2(g289_p)
  );


  LA
  g_g291_p
  (
    .dout(g291_p),
    .din1(g260_n_spl_0),
    .din2(g290_n)
  );


  FA
  g_g291_n
  (
    .dout(g291_n),
    .din1(g260_p_spl_0),
    .din2(g290_p)
  );


  LA
  g_g292_p
  (
    .dout(g292_p),
    .din1(g162_n_spl_10),
    .din2(g291_p_spl_)
  );


  FA
  g_g292_n
  (
    .dout(g292_n),
    .din1(g162_p_spl_10),
    .din2(g291_n_spl_)
  );


  LA
  g_g293_p
  (
    .dout(g293_p),
    .din1(g282_p_spl_0),
    .din2(g292_n)
  );


  FA
  g_g293_n
  (
    .dout(g293_n),
    .din1(g282_n_spl_0),
    .din2(g292_p)
  );


  LA
  g_g294_p
  (
    .dout(g294_p),
    .din1(g165_n_spl_10),
    .din2(g282_n_spl_0)
  );


  FA
  g_g294_n
  (
    .dout(g294_n),
    .din1(g165_p_spl_10),
    .din2(g282_p_spl_0)
  );


  LA
  g_g295_p
  (
    .dout(g295_p),
    .din1(g291_p_spl_),
    .din2(g294_p)
  );


  FA
  g_g295_n
  (
    .dout(g295_n),
    .din1(g291_n_spl_),
    .din2(g294_n)
  );


  LA
  g_g296_p
  (
    .dout(g296_p),
    .din1(g293_n),
    .din2(g295_n_spl_0)
  );


  FA
  g_g296_n
  (
    .dout(g296_n),
    .din1(g293_p),
    .din2(g295_p_spl_0)
  );


  LA
  g_g297_p
  (
    .dout(g297_p),
    .din1(G7_p_spl_001),
    .din2(g248_n_spl_1)
  );


  FA
  g_g297_n
  (
    .dout(g297_n),
    .din1(G7_n_spl_001),
    .din2(g248_p_spl_1)
  );


  LA
  g_g298_p
  (
    .dout(g298_p),
    .din1(G7_n_spl_010),
    .din2(g130_n_spl_11)
  );


  FA
  g_g298_n
  (
    .dout(g298_n),
    .din1(G7_p_spl_010),
    .din2(g130_p_spl_11)
  );


  LA
  g_g299_p
  (
    .dout(g299_p),
    .din1(g297_n),
    .din2(g298_n)
  );


  FA
  g_g299_n
  (
    .dout(g299_n),
    .din1(g297_p),
    .din2(g298_p)
  );


  LA
  g_g300_p
  (
    .dout(g300_p),
    .din1(G8_n_spl_010),
    .din2(g137_p_spl_11)
  );


  FA
  g_g300_n
  (
    .dout(g300_n),
    .din1(G8_p_spl_010),
    .din2(g137_n_spl_11)
  );


  LA
  g_g301_p
  (
    .dout(g301_p),
    .din1(G3_p_spl_100),
    .din2(g52_n)
  );


  FA
  g_g301_n
  (
    .dout(g301_n),
    .din1(G3_n_spl_100),
    .din2(g52_p_spl_)
  );


  LA
  g_g302_p
  (
    .dout(g302_p),
    .din1(G21_p_spl_00),
    .din2(g138_p_spl_11)
  );


  FA
  g_g302_n
  (
    .dout(g302_n),
    .din1(G21_n_spl_00),
    .din2(g138_n_spl_11)
  );


  LA
  g_g303_p
  (
    .dout(g303_p),
    .din1(g301_n),
    .din2(g302_n)
  );


  FA
  g_g303_n
  (
    .dout(g303_n),
    .din1(g301_p),
    .din2(g302_p)
  );


  LA
  g_g304_p
  (
    .dout(g304_p),
    .din1(g300_n),
    .din2(g303_p)
  );


  FA
  g_g304_n
  (
    .dout(g304_n),
    .din1(g300_p),
    .din2(g303_n)
  );


  LA
  g_g305_p
  (
    .dout(g305_p),
    .din1(g129_n_spl_11),
    .din2(g304_n)
  );


  FA
  g_g305_n
  (
    .dout(g305_n),
    .din1(g129_p_spl_11),
    .din2(g304_p)
  );


  LA
  g_g306_p
  (
    .dout(g306_p),
    .din1(g299_n),
    .din2(g305_n)
  );


  FA
  g_g306_n
  (
    .dout(g306_n),
    .din1(g299_p),
    .din2(g305_p)
  );


  LA
  g_g307_p
  (
    .dout(g307_p),
    .din1(G30_p_spl_1),
    .din2(g259_n_spl_1)
  );


  FA
  g_g307_n
  (
    .dout(g307_n),
    .din1(G30_n_spl_1),
    .din2(g259_p_spl_1)
  );


  LA
  g_g308_p
  (
    .dout(g308_p),
    .din1(G28_p),
    .din2(g153_p_spl_11)
  );


  FA
  g_g308_n
  (
    .dout(g308_n),
    .din1(G28_n),
    .din2(g153_n_spl_11)
  );


  LA
  g_g309_p
  (
    .dout(g309_p),
    .din1(g307_n),
    .din2(g308_n)
  );


  FA
  g_g309_n
  (
    .dout(g309_n),
    .din1(g307_p),
    .din2(g308_p)
  );


  LA
  g_g310_p
  (
    .dout(g310_p),
    .din1(G4_n_spl_0110),
    .din2(G10_n_spl_011)
  );


  FA
  g_g310_n
  (
    .dout(g310_n),
    .din1(G4_p_spl_0110),
    .din2(G10_p_spl_011)
  );


  LA
  g_g311_p
  (
    .dout(g311_p),
    .din1(G4_p_spl_0111),
    .din2(G29_n_spl_)
  );


  FA
  g_g311_n
  (
    .dout(g311_n),
    .din1(G4_n_spl_0111),
    .din2(G29_p_spl_)
  );


  LA
  g_g312_p
  (
    .dout(g312_p),
    .din1(g310_n),
    .din2(g311_n)
  );


  FA
  g_g312_n
  (
    .dout(g312_n),
    .din1(g310_p),
    .din2(g311_p)
  );


  LA
  g_g313_p
  (
    .dout(g313_p),
    .din1(g309_p),
    .din2(g312_n)
  );


  FA
  g_g313_n
  (
    .dout(g313_n),
    .din1(g309_n),
    .din2(g312_p)
  );


  LA
  g_g314_p
  (
    .dout(g314_p),
    .din1(g147_n_spl_11),
    .din2(g313_n)
  );


  FA
  g_g314_n
  (
    .dout(g314_n),
    .din1(g147_p_spl_11),
    .din2(g313_p)
  );


  LA
  g_g315_p
  (
    .dout(g315_p),
    .din1(g260_n_spl_1),
    .din2(g314_n)
  );


  FA
  g_g315_n
  (
    .dout(g315_n),
    .din1(g260_p_spl_1),
    .din2(g314_p)
  );


  LA
  g_g316_p
  (
    .dout(g316_p),
    .din1(g162_n_spl_10),
    .din2(g315_p_spl_)
  );


  FA
  g_g316_n
  (
    .dout(g316_n),
    .din1(g162_p_spl_10),
    .din2(g315_n_spl_)
  );


  LA
  g_g317_p
  (
    .dout(g317_p),
    .din1(g306_p_spl_0),
    .din2(g316_n)
  );


  FA
  g_g317_n
  (
    .dout(g317_n),
    .din1(g306_n_spl_0),
    .din2(g316_p)
  );


  LA
  g_g318_p
  (
    .dout(g318_p),
    .din1(g165_n_spl_11),
    .din2(g306_n_spl_0)
  );


  FA
  g_g318_n
  (
    .dout(g318_n),
    .din1(g165_p_spl_11),
    .din2(g306_p_spl_0)
  );


  LA
  g_g319_p
  (
    .dout(g319_p),
    .din1(g315_p_spl_),
    .din2(g318_p)
  );


  FA
  g_g319_n
  (
    .dout(g319_n),
    .din1(g315_n_spl_),
    .din2(g318_n)
  );


  LA
  g_g320_p
  (
    .dout(g320_p),
    .din1(g317_n),
    .din2(g319_n_spl_)
  );


  FA
  g_g320_n
  (
    .dout(g320_n),
    .din1(g317_p),
    .din2(g319_p_spl_)
  );


  LA
  g_g321_p
  (
    .dout(g321_p),
    .din1(G8_p_spl_011),
    .din2(g248_n_spl_1)
  );


  FA
  g_g321_n
  (
    .dout(g321_n),
    .din1(G8_n_spl_010),
    .din2(g248_p_spl_1)
  );


  LA
  g_g322_p
  (
    .dout(g322_p),
    .din1(G8_n_spl_011),
    .din2(g130_n_spl_11)
  );


  FA
  g_g322_n
  (
    .dout(g322_n),
    .din1(G8_p_spl_011),
    .din2(g130_p_spl_11)
  );


  LA
  g_g323_p
  (
    .dout(g323_p),
    .din1(g321_n),
    .din2(g322_n)
  );


  FA
  g_g323_n
  (
    .dout(g323_n),
    .din1(g321_p),
    .din2(g322_p)
  );


  LA
  g_g324_p
  (
    .dout(g324_p),
    .din1(G9_n_spl_011),
    .din2(g137_p_spl_11)
  );


  FA
  g_g324_n
  (
    .dout(g324_n),
    .din1(G9_p_spl_100),
    .din2(g137_n_spl_11)
  );


  LA
  g_g325_p
  (
    .dout(g325_p),
    .din1(G8_p_spl_100),
    .din2(G9_p_spl_100)
  );


  FA
  g_g325_n
  (
    .dout(g325_n),
    .din1(G8_n_spl_011),
    .din2(G9_n_spl_100)
  );


  LA
  g_g326_p
  (
    .dout(g326_p),
    .din1(g75_n_spl_),
    .din2(g325_n)
  );


  FA
  g_g326_n
  (
    .dout(g326_n),
    .din1(g75_p_spl_),
    .din2(g325_p)
  );


  LA
  g_g327_p
  (
    .dout(g327_p),
    .din1(G3_p_spl_100),
    .din2(g326_p)
  );


  FA
  g_g327_n
  (
    .dout(g327_n),
    .din1(G3_n_spl_100),
    .din2(g326_n_spl_)
  );


  LA
  g_g328_p
  (
    .dout(g328_p),
    .din1(G22_p_spl_00),
    .din2(g138_p_spl_11)
  );


  FA
  g_g328_n
  (
    .dout(g328_n),
    .din1(G22_n_spl_00),
    .din2(g138_n_spl_11)
  );


  LA
  g_g329_p
  (
    .dout(g329_p),
    .din1(g327_n),
    .din2(g328_n)
  );


  FA
  g_g329_n
  (
    .dout(g329_n),
    .din1(g327_p),
    .din2(g328_p)
  );


  LA
  g_g330_p
  (
    .dout(g330_p),
    .din1(g324_n),
    .din2(g329_p)
  );


  FA
  g_g330_n
  (
    .dout(g330_n),
    .din1(g324_p),
    .din2(g329_n)
  );


  LA
  g_g331_p
  (
    .dout(g331_p),
    .din1(g129_n_spl_11),
    .din2(g330_n)
  );


  FA
  g_g331_n
  (
    .dout(g331_n),
    .din1(g129_p_spl_11),
    .din2(g330_p)
  );


  LA
  g_g332_p
  (
    .dout(g332_p),
    .din1(g323_n),
    .din2(g331_n)
  );


  FA
  g_g332_n
  (
    .dout(g332_n),
    .din1(g323_p),
    .din2(g331_p)
  );


  LA
  g_g333_p
  (
    .dout(g333_p),
    .din1(G31_p_spl_1),
    .din2(g259_n_spl_1)
  );


  FA
  g_g333_n
  (
    .dout(g333_n),
    .din1(G31_n_spl_1),
    .din2(g259_p_spl_1)
  );


  LA
  g_g334_p
  (
    .dout(g334_p),
    .din1(G29_p_spl_),
    .din2(g153_p_spl_11)
  );


  FA
  g_g334_n
  (
    .dout(g334_n),
    .din1(G29_n_spl_),
    .din2(g153_n_spl_11)
  );


  LA
  g_g335_p
  (
    .dout(g335_p),
    .din1(g333_n),
    .din2(g334_n)
  );


  FA
  g_g335_n
  (
    .dout(g335_n),
    .din1(g333_p),
    .din2(g334_p)
  );


  LA
  g_g336_p
  (
    .dout(g336_p),
    .din1(G4_n_spl_0111),
    .din2(G11_n_spl_011)
  );


  FA
  g_g336_n
  (
    .dout(g336_n),
    .din1(G4_p_spl_0111),
    .din2(G11_p_spl_100)
  );


  LA
  g_g337_p
  (
    .dout(g337_p),
    .din1(G4_p_spl_1000),
    .din2(G30_n_spl_1)
  );


  FA
  g_g337_n
  (
    .dout(g337_n),
    .din1(G4_n_spl_1000),
    .din2(G30_p_spl_1)
  );


  LA
  g_g338_p
  (
    .dout(g338_p),
    .din1(g336_n),
    .din2(g337_n)
  );


  FA
  g_g338_n
  (
    .dout(g338_n),
    .din1(g336_p),
    .din2(g337_p)
  );


  LA
  g_g339_p
  (
    .dout(g339_p),
    .din1(g335_p),
    .din2(g338_n)
  );


  FA
  g_g339_n
  (
    .dout(g339_n),
    .din1(g335_n),
    .din2(g338_p)
  );


  LA
  g_g340_p
  (
    .dout(g340_p),
    .din1(g147_n_spl_11),
    .din2(g339_n)
  );


  FA
  g_g340_n
  (
    .dout(g340_n),
    .din1(g147_p_spl_11),
    .din2(g339_p)
  );


  LA
  g_g341_p
  (
    .dout(g341_p),
    .din1(g260_n_spl_1),
    .din2(g340_n)
  );


  FA
  g_g341_n
  (
    .dout(g341_n),
    .din1(g260_p_spl_1),
    .din2(g340_p)
  );


  LA
  g_g342_p
  (
    .dout(g342_p),
    .din1(g162_n_spl_11),
    .din2(g341_p_spl_)
  );


  FA
  g_g342_n
  (
    .dout(g342_n),
    .din1(g162_p_spl_11),
    .din2(g341_n_spl_)
  );


  LA
  g_g343_p
  (
    .dout(g343_p),
    .din1(g332_p_spl_0),
    .din2(g342_n)
  );


  FA
  g_g343_n
  (
    .dout(g343_n),
    .din1(g332_n_spl_0),
    .din2(g342_p)
  );


  LA
  g_g344_p
  (
    .dout(g344_p),
    .din1(g165_n_spl_11),
    .din2(g332_n_spl_0)
  );


  FA
  g_g344_n
  (
    .dout(g344_n),
    .din1(g165_p_spl_11),
    .din2(g332_p_spl_0)
  );


  LA
  g_g345_p
  (
    .dout(g345_p),
    .din1(g341_p_spl_),
    .din2(g344_p)
  );


  FA
  g_g345_n
  (
    .dout(g345_n),
    .din1(g341_n_spl_),
    .din2(g344_n)
  );


  LA
  g_g346_p
  (
    .dout(g346_p),
    .din1(g343_n),
    .din2(g345_n_spl_0)
  );


  FA
  g_g346_n
  (
    .dout(g346_n),
    .din1(g343_p),
    .din2(g345_p_spl_0)
  );


  LA
  g_g347_p
  (
    .dout(g347_p),
    .din1(g320_p_spl_0),
    .din2(g346_p_spl_0)
  );


  FA
  g_g347_n
  (
    .dout(g347_n),
    .din1(g320_n_spl_0),
    .din2(g346_n_spl_0)
  );


  LA
  g_g348_p
  (
    .dout(g348_p),
    .din1(g296_p_spl_0),
    .din2(g347_p_spl_)
  );


  FA
  g_g348_n
  (
    .dout(g348_n),
    .din1(g296_n_spl_0),
    .din2(g347_n_spl_)
  );


  LA
  g_g349_p
  (
    .dout(g349_p),
    .din1(g274_p_spl_0),
    .din2(g348_p_spl_)
  );


  FA
  g_g349_n
  (
    .dout(g349_n),
    .din1(g274_n_spl_0),
    .din2(g348_n_spl_)
  );


  LA
  g_g350_p
  (
    .dout(g350_p),
    .din1(g246_p_spl_),
    .din2(g349_p_spl_0)
  );


  LA
  g_g351_p
  (
    .dout(g351_p),
    .din1(g190_p_spl_0),
    .din2(g244_p_spl_)
  );


  FA
  g_g351_n
  (
    .dout(g351_n),
    .din1(g190_n_spl_0),
    .din2(g244_n_spl_)
  );


  LA
  g_g352_p
  (
    .dout(g352_p),
    .din1(g217_p_spl_0),
    .din2(g242_p_spl_0)
  );


  FA
  g_g352_n
  (
    .dout(g352_n),
    .din1(g217_n_spl_0),
    .din2(g242_n_spl_0)
  );


  LA
  g_g353_p
  (
    .dout(g353_p),
    .din1(g351_n),
    .din2(g352_n)
  );


  FA
  g_g353_n
  (
    .dout(g353_n),
    .din1(g351_p),
    .din2(g352_p)
  );


  LA
  g_g354_p
  (
    .dout(g354_p),
    .din1(g167_p_spl_0),
    .din2(g245_p_spl_)
  );


  FA
  g_g354_n
  (
    .dout(g354_n),
    .din1(g167_n_spl_0),
    .din2(g245_n_spl_)
  );


  LA
  g_g355_p
  (
    .dout(g355_p),
    .din1(g216_n_spl_),
    .din2(g354_n)
  );


  FA
  g_g355_n
  (
    .dout(g355_n),
    .din1(g216_p_spl_),
    .din2(g354_p)
  );


  LA
  g_g356_p
  (
    .dout(g356_p),
    .din1(g353_p),
    .din2(g355_p)
  );


  FA
  g_g356_n
  (
    .dout(g356_n),
    .din1(g353_n),
    .din2(g355_n)
  );


  LA
  g_g357_p
  (
    .dout(g357_p),
    .din1(g349_p_spl_0),
    .din2(g356_n_spl_)
  );


  LA
  g_g358_p
  (
    .dout(g358_p),
    .din1(g295_p_spl_0),
    .din2(g347_p_spl_)
  );


  FA
  g_g358_n
  (
    .dout(g358_n),
    .din1(g295_n_spl_0),
    .din2(g347_n_spl_)
  );


  LA
  g_g359_p
  (
    .dout(g359_p),
    .din1(g320_p_spl_0),
    .din2(g345_p_spl_0)
  );


  FA
  g_g359_n
  (
    .dout(g359_n),
    .din1(g320_n_spl_0),
    .din2(g345_n_spl_0)
  );


  LA
  g_g360_p
  (
    .dout(g360_p),
    .din1(g358_n),
    .din2(g359_n)
  );


  FA
  g_g360_n
  (
    .dout(g360_n),
    .din1(g358_p),
    .din2(g359_p)
  );


  LA
  g_g361_p
  (
    .dout(g361_p),
    .din1(g273_p_spl_0),
    .din2(g348_p_spl_)
  );


  FA
  g_g361_n
  (
    .dout(g361_n),
    .din1(g273_n_spl_0),
    .din2(g348_n_spl_)
  );


  LA
  g_g362_p
  (
    .dout(g362_p),
    .din1(g319_n_spl_),
    .din2(g361_n)
  );


  FA
  g_g362_n
  (
    .dout(g362_n),
    .din1(g319_p_spl_),
    .din2(g361_p)
  );


  LA
  g_g363_p
  (
    .dout(g363_p),
    .din1(g360_p),
    .din2(g362_p)
  );


  FA
  g_g363_n
  (
    .dout(g363_n),
    .din1(g360_n),
    .din2(g362_n)
  );


  FA
  g_g364_n
  (
    .dout(g364_n),
    .din1(g357_p),
    .din2(g363_n_spl_)
  );


  LA
  g_g365_p
  (
    .dout(g365_p),
    .din1(G27_p_spl_0),
    .din2(g79_p_spl_0)
  );


  FA
  g_g365_n
  (
    .dout(g365_n),
    .din1(G27_n_spl_),
    .din2(g79_n_spl_0)
  );


  LA
  g_g366_p
  (
    .dout(g366_p),
    .din1(G48_p_spl_),
    .din2(g365_p_spl_0)
  );


  FA
  g_g366_n
  (
    .dout(g366_n),
    .din1(G48_n_spl_),
    .din2(g365_n_spl_0)
  );


  LA
  g_g367_p
  (
    .dout(g367_p),
    .din1(g177_n_spl_),
    .din2(g366_p_spl_000)
  );


  FA
  g_g367_n
  (
    .dout(g367_n),
    .din1(g177_p_spl_),
    .din2(g366_n_spl_000)
  );


  LA
  g_g368_p
  (
    .dout(g368_p),
    .din1(g191_n_spl_0),
    .din2(g367_n_spl_)
  );


  FA
  g_g368_n
  (
    .dout(g368_n),
    .din1(g191_p_spl_0),
    .din2(g367_p_spl_)
  );


  LA
  g_g369_p
  (
    .dout(g369_p),
    .din1(g191_p_spl_),
    .din2(g367_p_spl_)
  );


  FA
  g_g369_n
  (
    .dout(g369_n),
    .din1(g191_n_spl_),
    .din2(g367_n_spl_)
  );


  LA
  g_g370_p
  (
    .dout(g370_p),
    .din1(g368_n),
    .din2(g369_n)
  );


  FA
  g_g370_n
  (
    .dout(g370_n),
    .din1(g368_p),
    .din2(g369_p)
  );


  LA
  g_g371_p
  (
    .dout(g371_p),
    .din1(g145_n_spl_),
    .din2(g366_p_spl_000)
  );


  FA
  g_g371_n
  (
    .dout(g371_n),
    .din1(g145_p_spl_),
    .din2(g366_n_spl_000)
  );


  LA
  g_g372_p
  (
    .dout(g372_p),
    .din1(g168_n_spl_0),
    .din2(g371_n_spl_)
  );


  FA
  g_g372_n
  (
    .dout(g372_n),
    .din1(g168_p_spl_0),
    .din2(g371_p_spl_)
  );


  LA
  g_g373_p
  (
    .dout(g373_p),
    .din1(g168_p_spl_),
    .din2(g371_p_spl_)
  );


  FA
  g_g373_n
  (
    .dout(g373_n),
    .din1(g168_n_spl_),
    .din2(g371_n_spl_)
  );


  LA
  g_g374_p
  (
    .dout(g374_p),
    .din1(g372_n),
    .din2(g373_n)
  );


  FA
  g_g374_n
  (
    .dout(g374_n),
    .din1(g372_p),
    .din2(g373_p)
  );


  LA
  g_g375_p
  (
    .dout(g375_p),
    .din1(G47_p_spl_00),
    .din2(g374_p_spl_0)
  );


  FA
  g_g375_n
  (
    .dout(g375_n),
    .din1(G47_n_spl_00),
    .din2(g374_n_spl_0)
  );


  LA
  g_g376_p
  (
    .dout(g376_p),
    .din1(g370_n_spl_0),
    .din2(g375_p)
  );


  FA
  g_g376_n
  (
    .dout(g376_n),
    .din1(g370_p_spl_0),
    .din2(g375_n)
  );


  LA
  g_g377_p
  (
    .dout(g377_p),
    .din1(G5_p_spl_01),
    .din2(g79_p_spl_0)
  );


  FA
  g_g377_n
  (
    .dout(g377_n),
    .din1(G5_n_spl_01),
    .din2(g79_n_spl_1)
  );


  LA
  g_g378_p
  (
    .dout(g378_p),
    .din1(g76_p_spl_),
    .din2(g377_n_spl_00)
  );


  LA
  g_g379_p
  (
    .dout(g379_p),
    .din1(g356_n_spl_),
    .din2(g366_n_spl_001)
  );


  FA
  g_g379_n
  (
    .dout(g379_n),
    .din1(g356_p),
    .din2(g366_p_spl_001)
  );


  LA
  g_g380_p
  (
    .dout(g380_p),
    .din1(G1_n_spl_11),
    .din2(g379_p_spl_00)
  );


  FA
  g_g381_n
  (
    .dout(g381_n),
    .din1(g378_p),
    .din2(g380_p)
  );


  LA
  g_g382_p
  (
    .dout(g382_p),
    .din1(G2_n_spl_1),
    .din2(G3_n_spl_101)
  );


  FA
  g_g382_n
  (
    .dout(g382_n),
    .din1(G2_p_spl_1),
    .din2(G3_p_spl_101)
  );


  LA
  g_g383_p
  (
    .dout(g383_p),
    .din1(G6_p_spl_01),
    .din2(g382_p_spl_)
  );


  FA
  g_g383_n
  (
    .dout(g383_n),
    .din1(G6_n_spl_01),
    .din2(g382_n_spl_)
  );


  LA
  g_g384_p
  (
    .dout(g384_p),
    .din1(G1_n_spl_11),
    .din2(g383_n)
  );


  FA
  g_g384_n
  (
    .dout(g384_n),
    .din1(G1_p_spl_11),
    .din2(g383_p)
  );


  LA
  g_g385_p
  (
    .dout(g385_p),
    .din1(g377_p_spl_00),
    .din2(g384_p_spl_00)
  );


  FA
  g_g385_n
  (
    .dout(g385_n),
    .din1(g377_n_spl_00),
    .din2(g384_n_spl_00)
  );


  LA
  g_g386_p
  (
    .dout(g386_p),
    .din1(G47_n_spl_00),
    .din2(g374_p_spl_0)
  );


  FA
  g_g386_n
  (
    .dout(g386_n),
    .din1(G47_p_spl_00),
    .din2(g374_n_spl_0)
  );


  LA
  g_g387_p
  (
    .dout(g387_p),
    .din1(G47_p_spl_01),
    .din2(g374_n_spl_1)
  );


  FA
  g_g387_n
  (
    .dout(g387_n),
    .din1(G47_n_spl_01),
    .din2(g374_p_spl_1)
  );


  LA
  g_g388_p
  (
    .dout(g388_p),
    .din1(g386_n),
    .din2(g387_n_spl_0)
  );


  FA
  g_g388_n
  (
    .dout(g388_n),
    .din1(g386_p),
    .din2(g387_p_spl_0)
  );


  LA
  g_g389_p
  (
    .dout(g389_p),
    .din1(g385_n_spl_000),
    .din2(g388_p)
  );


  FA
  g_g389_n
  (
    .dout(g389_n),
    .din1(g385_p_spl_000),
    .din2(g388_n)
  );


  LA
  g_g390_p
  (
    .dout(g390_p),
    .din1(G4_p_spl_1000),
    .din2(g382_p_spl_)
  );


  FA
  g_g390_n
  (
    .dout(g390_n),
    .din1(G4_n_spl_1000),
    .din2(g382_n_spl_)
  );


  LA
  g_g391_p
  (
    .dout(g391_p),
    .din1(g374_p_spl_1),
    .din2(g390_p_spl_0)
  );


  FA
  g_g391_n
  (
    .dout(g391_n),
    .din1(g374_n_spl_1),
    .din2(g390_n_spl_0)
  );


  LA
  g_g392_p
  (
    .dout(g392_p),
    .din1(G3_p_spl_101),
    .din2(G23_n_spl_)
  );


  FA
  g_g392_n
  (
    .dout(g392_n),
    .din1(G3_n_spl_101),
    .din2(G23_p_spl_)
  );


  LA
  g_g393_p
  (
    .dout(g393_p),
    .din1(g73_p_spl_),
    .din2(g392_n)
  );


  FA
  g_g393_n
  (
    .dout(g393_n),
    .din1(g73_n_spl_),
    .din2(g392_p)
  );


  LA
  g_g394_p
  (
    .dout(g394_p),
    .din1(G4_n_spl_1001),
    .din2(g79_p_spl_)
  );


  FA
  g_g394_n
  (
    .dout(g394_n),
    .din1(G4_p_spl_1001),
    .din2(g79_n_spl_1)
  );


  LA
  g_g395_p
  (
    .dout(g395_p),
    .din1(G14_p_spl_011),
    .din2(g394_n_spl_00)
  );


  FA
  g_g395_n
  (
    .dout(g395_n),
    .din1(G14_n_spl_011),
    .din2(g394_p_spl_00)
  );


  LA
  g_g396_p
  (
    .dout(g396_p),
    .din1(G6_n_spl_01),
    .din2(g122_n_spl_)
  );


  FA
  g_g396_n
  (
    .dout(g396_n),
    .din1(G6_p_spl_01),
    .din2(g122_p_spl_)
  );


  LA
  g_g397_p
  (
    .dout(g397_p),
    .din1(G6_p_spl_10),
    .din2(g76_n_spl_)
  );


  FA
  g_g397_n
  (
    .dout(g397_n),
    .din1(G6_n_spl_10),
    .din2(g76_p_spl_)
  );


  LA
  g_g398_p
  (
    .dout(g398_p),
    .din1(g55_p),
    .din2(g397_n)
  );


  FA
  g_g398_n
  (
    .dout(g398_n),
    .din1(g55_n_spl_),
    .din2(g397_p)
  );


  LA
  g_g399_p
  (
    .dout(g399_p),
    .din1(g396_n),
    .din2(g398_p)
  );


  FA
  g_g399_n
  (
    .dout(g399_n),
    .din1(g396_p),
    .din2(g398_n)
  );


  LA
  g_g400_p
  (
    .dout(g400_p),
    .din1(g394_p_spl_00),
    .din2(g399_p)
  );


  FA
  g_g400_n
  (
    .dout(g400_n),
    .din1(g394_n_spl_00),
    .din2(g399_n)
  );


  LA
  g_g401_p
  (
    .dout(g401_p),
    .din1(g395_n),
    .din2(g400_n)
  );


  FA
  g_g401_n
  (
    .dout(g401_n),
    .din1(g395_p),
    .din2(g400_p)
  );


  LA
  g_g402_p
  (
    .dout(g402_p),
    .din1(g393_p_spl_000),
    .din2(g401_n)
  );


  FA
  g_g402_n
  (
    .dout(g402_n),
    .din1(g393_n_spl_000),
    .din2(g401_p)
  );


  LA
  g_g403_p
  (
    .dout(g403_p),
    .din1(G3_p_spl_110),
    .din2(G25_p_spl_)
  );


  FA
  g_g403_n
  (
    .dout(g403_n),
    .din1(G3_n_spl_110),
    .din2(G25_n_spl_)
  );


  LA
  g_g404_p
  (
    .dout(g404_p),
    .din1(G3_p_spl_110),
    .din2(G24_p_spl_0)
  );


  FA
  g_g404_n
  (
    .dout(g404_n),
    .din1(G3_n_spl_110),
    .din2(G24_n_spl_0)
  );


  LA
  g_g405_p
  (
    .dout(g405_p),
    .din1(G26_p_spl_0),
    .din2(g404_n_spl_0)
  );


  FA
  g_g405_n
  (
    .dout(g405_n),
    .din1(G26_n_spl_0),
    .din2(g404_p_spl_0)
  );


  LA
  g_g406_p
  (
    .dout(g406_p),
    .din1(g403_n_spl_0),
    .din2(g405_p_spl_)
  );


  FA
  g_g406_n
  (
    .dout(g406_n),
    .din1(g403_p_spl_0),
    .din2(g405_n_spl_)
  );


  LA
  g_g407_p
  (
    .dout(g407_p),
    .din1(G45_p_spl_),
    .din2(g406_n_spl_0000)
  );


  FA
  g_g407_n
  (
    .dout(g407_n),
    .din1(G45_n_spl_),
    .din2(g406_p_spl_0000)
  );


  LA
  g_g408_p
  (
    .dout(g408_p),
    .din1(G26_n_spl_),
    .din2(g404_n_spl_0)
  );


  FA
  g_g408_n
  (
    .dout(g408_n),
    .din1(G26_p_spl_),
    .din2(g404_p_spl_0)
  );


  LA
  g_g409_p
  (
    .dout(g409_p),
    .din1(g403_n_spl_0),
    .din2(g408_p_spl_)
  );


  FA
  g_g409_n
  (
    .dout(g409_n),
    .din1(g403_p_spl_0),
    .din2(g408_n_spl_)
  );


  LA
  g_g410_p
  (
    .dout(g410_p),
    .din1(G44_p_spl_0),
    .din2(g409_n_spl_000)
  );


  FA
  g_g410_n
  (
    .dout(g410_n),
    .din1(G44_n_spl_0),
    .din2(g409_p_spl_000)
  );


  LA
  g_g411_p
  (
    .dout(g411_p),
    .din1(g407_n),
    .din2(g410_n)
  );


  FA
  g_g411_n
  (
    .dout(g411_n),
    .din1(g407_p),
    .din2(g410_p)
  );


  LA
  g_g412_p
  (
    .dout(g412_p),
    .din1(g403_p_spl_1),
    .din2(g408_p_spl_)
  );


  FA
  g_g412_n
  (
    .dout(g412_n),
    .din1(g403_n_spl_1),
    .din2(g408_n_spl_)
  );


  LA
  g_g413_p
  (
    .dout(g413_p),
    .din1(G42_p_spl_0),
    .din2(g412_n_spl_0000)
  );


  FA
  g_g413_n
  (
    .dout(g413_n),
    .din1(G42_n_spl_0),
    .din2(g412_p_spl_0000)
  );


  LA
  g_g414_p
  (
    .dout(g414_p),
    .din1(g403_p_spl_1),
    .din2(g405_p_spl_)
  );


  FA
  g_g414_n
  (
    .dout(g414_n),
    .din1(g403_n_spl_1),
    .din2(g405_n_spl_)
  );


  LA
  g_g415_p
  (
    .dout(g415_p),
    .din1(G39_p_spl_00),
    .din2(g414_n_spl_0000)
  );


  FA
  g_g415_n
  (
    .dout(g415_n),
    .din1(G39_n_spl_00),
    .din2(g414_p_spl_0000)
  );


  LA
  g_g416_p
  (
    .dout(g416_p),
    .din1(g413_n),
    .din2(g415_n)
  );


  FA
  g_g416_n
  (
    .dout(g416_n),
    .din1(g413_p),
    .din2(g415_p)
  );


  LA
  g_g417_p
  (
    .dout(g417_p),
    .din1(G46_p),
    .din2(g412_n_spl_0000)
  );


  FA
  g_g417_n
  (
    .dout(g417_n),
    .din1(G46_n),
    .din2(g412_p_spl_0000)
  );


  LA
  g_g418_p
  (
    .dout(g418_p),
    .din1(G43_p_spl_0),
    .din2(g414_n_spl_0000)
  );


  FA
  g_g418_n
  (
    .dout(g418_n),
    .din1(G43_n_spl_0),
    .din2(g414_p_spl_0000)
  );


  LA
  g_g419_p
  (
    .dout(g419_p),
    .din1(g417_n),
    .din2(g418_n)
  );


  FA
  g_g419_n
  (
    .dout(g419_n),
    .din1(g417_p),
    .din2(g418_p)
  );


  LA
  g_g420_p
  (
    .dout(g420_p),
    .din1(g416_p_spl_),
    .din2(g419_p)
  );


  FA
  g_g420_n
  (
    .dout(g420_n),
    .din1(g416_n_spl_),
    .din2(g419_n)
  );


  LA
  g_g421_p
  (
    .dout(g421_p),
    .din1(g411_p),
    .din2(g420_p)
  );


  FA
  g_g421_n
  (
    .dout(g421_n),
    .din1(g411_n),
    .din2(g420_n)
  );


  LA
  g_g422_p
  (
    .dout(g422_p),
    .din1(G3_p_spl_111),
    .din2(g162_n_spl_11)
  );


  FA
  g_g422_n
  (
    .dout(g422_n),
    .din1(G3_n_spl_111),
    .din2(g162_p_spl_11)
  );


  LA
  g_g423_p
  (
    .dout(g423_p),
    .din1(g404_n_spl_),
    .din2(g422_n)
  );


  FA
  g_g423_n
  (
    .dout(g423_n),
    .din1(g404_p_spl_),
    .din2(g422_p)
  );


  LA
  g_g424_p
  (
    .dout(g424_p),
    .din1(G40_p_spl_00),
    .din2(g423_n_spl_000)
  );


  FA
  g_g424_n
  (
    .dout(g424_n),
    .din1(G40_n_spl_00),
    .din2(g423_p_spl_000)
  );


  LA
  g_g425_p
  (
    .dout(g425_p),
    .din1(G3_p_spl_111),
    .din2(g406_p_spl_0000)
  );


  FA
  g_g425_n
  (
    .dout(g425_n),
    .din1(G3_n_spl_111),
    .din2(g406_n_spl_0000)
  );


  LA
  g_g426_p
  (
    .dout(g426_p),
    .din1(G41_p_spl_00),
    .din2(g425_n_spl_000)
  );


  FA
  g_g426_n
  (
    .dout(g426_n),
    .din1(G41_n_spl_00),
    .din2(g425_p_spl_000)
  );


  LA
  g_g427_p
  (
    .dout(g427_p),
    .din1(G4_p_spl_1001),
    .din2(g426_n)
  );


  FA
  g_g427_n
  (
    .dout(g427_n),
    .din1(G4_n_spl_1001),
    .din2(g426_p)
  );


  LA
  g_g428_p
  (
    .dout(g428_p),
    .din1(g424_n),
    .din2(g427_p)
  );


  FA
  g_g428_n
  (
    .dout(g428_n),
    .din1(g424_p),
    .din2(g427_n)
  );


  LA
  g_g429_p
  (
    .dout(g429_p),
    .din1(g421_p),
    .din2(g428_p)
  );


  FA
  g_g429_n
  (
    .dout(g429_n),
    .din1(g421_n),
    .din2(g428_n)
  );


  LA
  g_g430_p
  (
    .dout(g430_p),
    .din1(G11_n_spl_100),
    .din2(g425_n_spl_000)
  );


  FA
  g_g430_n
  (
    .dout(g430_n),
    .din1(G11_p_spl_100),
    .din2(g425_p_spl_000)
  );


  LA
  g_g431_p
  (
    .dout(g431_p),
    .din1(G10_n_spl_100),
    .din2(g412_n_spl_0001)
  );


  FA
  g_g431_n
  (
    .dout(g431_n),
    .din1(G10_p_spl_100),
    .din2(g412_p_spl_0001)
  );


  LA
  g_g432_p
  (
    .dout(g432_p),
    .din1(G13_n_spl_100),
    .din2(g414_n_spl_0001)
  );


  FA
  g_g432_n
  (
    .dout(g432_n),
    .din1(G13_p_spl_101),
    .din2(g414_p_spl_0001)
  );


  LA
  g_g433_p
  (
    .dout(g433_p),
    .din1(g431_n),
    .din2(g432_n_spl_)
  );


  FA
  g_g433_n
  (
    .dout(g433_n),
    .din1(g431_p),
    .din2(g432_p_spl_)
  );


  LA
  g_g434_p
  (
    .dout(g434_p),
    .din1(g430_n_spl_),
    .din2(g433_p)
  );


  FA
  g_g434_n
  (
    .dout(g434_n),
    .din1(g430_p_spl_),
    .din2(g433_n)
  );


  LA
  g_g435_p
  (
    .dout(g435_p),
    .din1(G7_n_spl_010),
    .din2(g406_n_spl_000)
  );


  FA
  g_g435_n
  (
    .dout(g435_n),
    .din1(G7_p_spl_010),
    .din2(g406_p_spl_000)
  );


  LA
  g_g436_p
  (
    .dout(g436_p),
    .din1(G8_n_spl_100),
    .din2(g409_n_spl_000)
  );


  FA
  g_g436_n
  (
    .dout(g436_n),
    .din1(G8_p_spl_100),
    .din2(g409_p_spl_000)
  );


  LA
  g_g437_p
  (
    .dout(g437_p),
    .din1(g435_n),
    .din2(g436_n)
  );


  FA
  g_g437_n
  (
    .dout(g437_n),
    .din1(g435_p),
    .din2(g436_p)
  );


  LA
  g_g438_p
  (
    .dout(g438_p),
    .din1(G9_n_spl_100),
    .din2(g414_n_spl_0001)
  );


  FA
  g_g438_n
  (
    .dout(g438_n),
    .din1(G9_p_spl_101),
    .din2(g414_p_spl_0001)
  );


  LA
  g_g439_p
  (
    .dout(g439_p),
    .din1(G4_n_spl_1010),
    .din2(g438_n_spl_)
  );


  FA
  g_g439_n
  (
    .dout(g439_n),
    .din1(G4_p_spl_1010),
    .din2(g438_p_spl_)
  );


  LA
  g_g440_p
  (
    .dout(g440_p),
    .din1(G12_n_spl_100),
    .din2(g423_n_spl_000)
  );


  FA
  g_g440_n
  (
    .dout(g440_n),
    .din1(G12_p_spl_101),
    .din2(g423_p_spl_000)
  );


  LA
  g_g441_p
  (
    .dout(g441_p),
    .din1(G22_p_spl_00),
    .din2(g412_n_spl_0001)
  );


  FA
  g_g441_n
  (
    .dout(g441_n),
    .din1(G22_n_spl_00),
    .din2(g412_p_spl_0001)
  );


  LA
  g_g442_p
  (
    .dout(g442_p),
    .din1(g440_n_spl_),
    .din2(g441_n_spl_)
  );


  FA
  g_g442_n
  (
    .dout(g442_n),
    .din1(g440_p_spl_),
    .din2(g441_p_spl_)
  );


  LA
  g_g443_p
  (
    .dout(g443_p),
    .din1(g439_p_spl_),
    .din2(g442_p)
  );


  FA
  g_g443_n
  (
    .dout(g443_n),
    .din1(g439_n_spl_),
    .din2(g442_n)
  );


  LA
  g_g444_p
  (
    .dout(g444_p),
    .din1(g437_p),
    .din2(g443_p)
  );


  FA
  g_g444_n
  (
    .dout(g444_n),
    .din1(g437_n),
    .din2(g443_n)
  );


  LA
  g_g445_p
  (
    .dout(g445_p),
    .din1(g434_p),
    .din2(g444_p)
  );


  FA
  g_g445_n
  (
    .dout(g445_n),
    .din1(g434_n),
    .din2(g444_n)
  );


  LA
  g_g446_p
  (
    .dout(g446_p),
    .din1(g429_n),
    .din2(g445_n)
  );


  FA
  g_g446_n
  (
    .dout(g446_n),
    .din1(g429_p),
    .din2(g445_p)
  );


  LA
  g_g447_p
  (
    .dout(g447_p),
    .din1(g393_n_spl_000),
    .din2(g446_p)
  );


  FA
  g_g447_n
  (
    .dout(g447_n),
    .din1(g393_p_spl_000),
    .din2(g446_n)
  );


  LA
  g_g448_p
  (
    .dout(g448_p),
    .din1(g402_n),
    .din2(g447_n)
  );


  FA
  g_g448_n
  (
    .dout(g448_n),
    .din1(g402_p),
    .din2(g447_p)
  );


  LA
  g_g449_p
  (
    .dout(g449_p),
    .din1(g391_n),
    .din2(g448_n)
  );


  FA
  g_g449_n
  (
    .dout(g449_n),
    .din1(g391_p),
    .din2(g448_p)
  );


  LA
  g_g450_p
  (
    .dout(g450_p),
    .din1(g385_p_spl_000),
    .din2(g449_p)
  );


  FA
  g_g450_n
  (
    .dout(g450_n),
    .din1(g385_n_spl_000),
    .din2(g449_n)
  );


  LA
  g_g451_p
  (
    .dout(g451_p),
    .din1(g389_n),
    .din2(g450_n)
  );


  FA
  g_g451_n
  (
    .dout(g451_n),
    .din1(g389_p),
    .din2(g450_p)
  );


  LA
  g_g452_p
  (
    .dout(g452_p),
    .din1(G2_n_spl_1),
    .din2(G4_p_spl_1010)
  );


  FA
  g_g452_n
  (
    .dout(g452_n),
    .din1(G2_p_spl_1),
    .din2(G4_n_spl_1010)
  );


  LA
  g_g453_p
  (
    .dout(g453_p),
    .din1(g257_n_spl_),
    .din2(g366_p_spl_001)
  );


  FA
  g_g453_n
  (
    .dout(g453_n),
    .din1(g257_p_spl_),
    .din2(g366_n_spl_001)
  );


  LA
  g_g454_p
  (
    .dout(g454_p),
    .din1(g274_n_spl_0),
    .din2(g453_n_spl_)
  );


  FA
  g_g454_n
  (
    .dout(g454_n),
    .din1(g274_p_spl_0),
    .din2(g453_p_spl_)
  );


  LA
  g_g455_p
  (
    .dout(g455_p),
    .din1(g274_p_spl_),
    .din2(g453_p_spl_)
  );


  FA
  g_g455_n
  (
    .dout(g455_n),
    .din1(g274_n_spl_),
    .din2(g453_n_spl_)
  );


  LA
  g_g456_p
  (
    .dout(g456_p),
    .din1(g454_n),
    .din2(g455_n)
  );


  FA
  g_g456_n
  (
    .dout(g456_n),
    .din1(g454_p),
    .din2(g455_p)
  );


  LA
  g_g457_p
  (
    .dout(g457_p),
    .din1(g452_p_spl_0),
    .din2(g456_p_spl_0)
  );


  FA
  g_g457_n
  (
    .dout(g457_n),
    .din1(g452_n_spl_0),
    .din2(g456_n_spl_0)
  );


  LA
  g_g458_p
  (
    .dout(g458_p),
    .din1(G10_n_spl_100),
    .din2(g393_p_spl_001)
  );


  FA
  g_g458_n
  (
    .dout(g458_n),
    .din1(G10_p_spl_100),
    .din2(g393_n_spl_001)
  );


  LA
  g_g459_p
  (
    .dout(g459_p),
    .din1(g385_p_spl_001),
    .din2(g458_n)
  );


  FA
  g_g459_n
  (
    .dout(g459_n),
    .din1(g385_n_spl_001),
    .din2(g458_p)
  );


  LA
  g_g460_p
  (
    .dout(g460_p),
    .din1(G8_n_spl_100),
    .din2(g423_n_spl_001)
  );


  FA
  g_g460_n
  (
    .dout(g460_n),
    .din1(G8_p_spl_101),
    .din2(g423_p_spl_001)
  );


  LA
  g_g461_p
  (
    .dout(g461_p),
    .din1(g441_n_spl_),
    .din2(g460_n)
  );


  FA
  g_g461_n
  (
    .dout(g461_n),
    .din1(g441_p_spl_),
    .din2(g460_p)
  );


  LA
  g_g462_p
  (
    .dout(g462_p),
    .din1(G20_p_spl_00),
    .din2(g409_n_spl_001)
  );


  FA
  g_g462_n
  (
    .dout(g462_n),
    .din1(G20_n_spl_00),
    .din2(g409_p_spl_001)
  );


  LA
  g_g463_p
  (
    .dout(g463_p),
    .din1(G21_p_spl_00),
    .din2(g414_n_spl_001)
  );


  FA
  g_g463_n
  (
    .dout(g463_n),
    .din1(G21_n_spl_00),
    .din2(g414_p_spl_001)
  );


  LA
  g_g464_p
  (
    .dout(g464_p),
    .din1(g462_n),
    .din2(g463_n)
  );


  FA
  g_g464_n
  (
    .dout(g464_n),
    .din1(g462_p),
    .din2(g463_p)
  );


  LA
  g_g465_p
  (
    .dout(g465_p),
    .din1(g439_p_spl_),
    .din2(g464_p)
  );


  FA
  g_g465_n
  (
    .dout(g465_n),
    .din1(g439_n_spl_),
    .din2(g464_n)
  );


  LA
  g_g466_p
  (
    .dout(g466_p),
    .din1(g461_p),
    .din2(g465_p)
  );


  FA
  g_g466_n
  (
    .dout(g466_n),
    .din1(g461_n),
    .din2(g465_n)
  );


  LA
  g_g467_p
  (
    .dout(g467_p),
    .din1(G18_p_spl_0),
    .din2(g412_n_spl_0010)
  );


  FA
  g_g467_n
  (
    .dout(g467_n),
    .din1(G18_n_spl_0),
    .din2(g412_p_spl_0010)
  );


  LA
  g_g468_p
  (
    .dout(g468_p),
    .din1(G7_n_spl_011),
    .din2(g425_n_spl_001)
  );


  FA
  g_g468_n
  (
    .dout(g468_n),
    .din1(G7_p_spl_011),
    .din2(g425_p_spl_001)
  );


  LA
  g_g469_p
  (
    .dout(g469_p),
    .din1(G19_p_spl_00),
    .din2(g406_n_spl_001)
  );


  FA
  g_g469_n
  (
    .dout(g469_n),
    .din1(G19_n_spl_00),
    .din2(g406_p_spl_001)
  );


  LA
  g_g470_p
  (
    .dout(g470_p),
    .din1(g468_n),
    .din2(g469_n)
  );


  FA
  g_g470_n
  (
    .dout(g470_n),
    .din1(g468_p),
    .din2(g469_p)
  );


  LA
  g_g471_p
  (
    .dout(g471_p),
    .din1(g467_n),
    .din2(g470_p)
  );


  FA
  g_g471_n
  (
    .dout(g471_n),
    .din1(g467_p),
    .din2(g470_n)
  );


  LA
  g_g472_p
  (
    .dout(g472_p),
    .din1(g466_p),
    .din2(g471_p)
  );


  FA
  g_g472_n
  (
    .dout(g472_n),
    .din1(g466_n),
    .din2(g471_n)
  );


  LA
  g_g473_p
  (
    .dout(g473_p),
    .din1(G13_n_spl_101),
    .din2(g425_n_spl_001)
  );


  FA
  g_g473_n
  (
    .dout(g473_n),
    .din1(G13_p_spl_101),
    .din2(g425_p_spl_001)
  );


  LA
  g_g474_p
  (
    .dout(g474_p),
    .din1(g416_p_spl_),
    .din2(g440_n_spl_)
  );


  FA
  g_g474_n
  (
    .dout(g474_n),
    .din1(g416_n_spl_),
    .din2(g440_p_spl_)
  );


  LA
  g_g475_p
  (
    .dout(g475_p),
    .din1(g473_n),
    .din2(g474_p)
  );


  FA
  g_g475_n
  (
    .dout(g475_n),
    .din1(g473_p),
    .din2(g474_n)
  );


  LA
  g_g476_p
  (
    .dout(g476_p),
    .din1(G40_p_spl_01),
    .din2(g409_n_spl_001)
  );


  FA
  g_g476_n
  (
    .dout(g476_n),
    .din1(G40_n_spl_01),
    .din2(g409_p_spl_001)
  );


  LA
  g_g477_p
  (
    .dout(g477_p),
    .din1(G14_n_spl_011),
    .din2(g412_n_spl_0010)
  );


  FA
  g_g477_n
  (
    .dout(g477_n),
    .din1(G14_p_spl_100),
    .din2(g412_p_spl_0010)
  );


  LA
  g_g478_p
  (
    .dout(g478_p),
    .din1(g476_n),
    .din2(g477_n)
  );


  FA
  g_g478_n
  (
    .dout(g478_n),
    .din1(g476_p),
    .din2(g477_p)
  );


  LA
  g_g479_p
  (
    .dout(g479_p),
    .din1(G41_p_spl_01),
    .din2(g406_n_spl_001)
  );


  FA
  g_g479_n
  (
    .dout(g479_n),
    .din1(G41_n_spl_01),
    .din2(g406_p_spl_001)
  );


  LA
  g_g480_p
  (
    .dout(g480_p),
    .din1(G11_n_spl_100),
    .din2(g414_n_spl_001)
  );


  FA
  g_g480_n
  (
    .dout(g480_n),
    .din1(G11_p_spl_101),
    .din2(g414_p_spl_001)
  );


  LA
  g_g481_p
  (
    .dout(g481_p),
    .din1(g479_n),
    .din2(g480_n_spl_)
  );


  FA
  g_g481_n
  (
    .dout(g481_n),
    .din1(g479_p),
    .din2(g480_p_spl_)
  );


  LA
  g_g482_p
  (
    .dout(g482_p),
    .din1(g478_p),
    .din2(g481_p)
  );


  FA
  g_g482_n
  (
    .dout(g482_n),
    .din1(g478_n),
    .din2(g481_n)
  );


  LA
  g_g483_p
  (
    .dout(g483_p),
    .din1(G4_p_spl_1011),
    .din2(g482_p)
  );


  FA
  g_g483_n
  (
    .dout(g483_n),
    .din1(G4_n_spl_1011),
    .din2(g482_n)
  );


  LA
  g_g484_p
  (
    .dout(g484_p),
    .din1(g475_p),
    .din2(g483_p)
  );


  FA
  g_g484_n
  (
    .dout(g484_n),
    .din1(g475_n),
    .din2(g483_n)
  );


  LA
  g_g485_p
  (
    .dout(g485_p),
    .din1(g472_n),
    .din2(g484_n)
  );


  FA
  g_g485_n
  (
    .dout(g485_n),
    .din1(g472_p),
    .din2(g484_p)
  );


  LA
  g_g486_p
  (
    .dout(g486_p),
    .din1(g393_n_spl_001),
    .din2(g485_n)
  );


  FA
  g_g486_n
  (
    .dout(g486_n),
    .din1(g393_p_spl_001),
    .din2(g485_p)
  );


  LA
  g_g487_p
  (
    .dout(g487_p),
    .din1(g459_p),
    .din2(g486_n)
  );


  FA
  g_g487_n
  (
    .dout(g487_n),
    .din1(g459_n),
    .din2(g486_p)
  );


  LA
  g_g488_p
  (
    .dout(g488_p),
    .din1(g457_n),
    .din2(g487_p)
  );


  FA
  g_g488_n
  (
    .dout(g488_n),
    .din1(g457_p),
    .din2(g487_n)
  );


  LA
  g_g489_p
  (
    .dout(g489_p),
    .din1(g212_n_spl_1),
    .din2(g238_n_spl_1)
  );


  FA
  g_g489_n
  (
    .dout(g489_n),
    .din1(g212_p_spl_1),
    .din2(g238_p_spl_1)
  );


  LA
  g_g490_p
  (
    .dout(g490_p),
    .din1(g161_n_spl_1),
    .din2(g186_n_spl_1)
  );


  FA
  g_g490_n
  (
    .dout(g490_n),
    .din1(g161_p_spl_1),
    .din2(g186_p_spl_1)
  );


  LA
  g_g491_p
  (
    .dout(g491_p),
    .din1(g489_p),
    .din2(g490_p)
  );


  FA
  g_g491_n
  (
    .dout(g491_n),
    .din1(g489_n),
    .din2(g490_n)
  );


  LA
  g_g492_p
  (
    .dout(g492_p),
    .din1(G24_p_spl_1),
    .din2(g491_n)
  );


  FA
  g_g492_n
  (
    .dout(g492_n),
    .din1(G24_n_spl_1),
    .din2(g491_p)
  );


  LA
  g_g493_p
  (
    .dout(g493_p),
    .din1(g212_p_spl_1),
    .din2(g238_p_spl_1)
  );


  FA
  g_g493_n
  (
    .dout(g493_n),
    .din1(g212_n_spl_1),
    .din2(g238_n_spl_1)
  );


  LA
  g_g494_p
  (
    .dout(g494_p),
    .din1(g161_p_spl_1),
    .din2(g186_p_spl_1)
  );


  FA
  g_g494_n
  (
    .dout(g494_n),
    .din1(g161_n_spl_1),
    .din2(g186_n_spl_1)
  );


  LA
  g_g495_p
  (
    .dout(g495_p),
    .din1(g493_p),
    .din2(g494_p)
  );


  FA
  g_g495_n
  (
    .dout(g495_n),
    .din1(g493_n),
    .din2(g494_n)
  );


  LA
  g_g496_p
  (
    .dout(g496_p),
    .din1(G24_n_spl_1),
    .din2(g495_n)
  );


  FA
  g_g496_n
  (
    .dout(g496_n),
    .din1(G24_p_spl_1),
    .din2(g495_p)
  );


  LA
  g_g497_p
  (
    .dout(g497_p),
    .din1(g492_n),
    .din2(g496_n)
  );


  FA
  g_g497_n
  (
    .dout(g497_n),
    .din1(g492_p),
    .din2(g496_p)
  );


  LA
  g_g498_p
  (
    .dout(g498_p),
    .din1(g366_n_spl_010),
    .din2(g497_n)
  );


  FA
  g_g498_n
  (
    .dout(g498_n),
    .din1(g366_p_spl_010),
    .din2(g497_p)
  );


  LA
  g_g499_p
  (
    .dout(g499_p),
    .din1(g246_n),
    .din2(g366_p_spl_010)
  );


  FA
  g_g499_n
  (
    .dout(g499_n),
    .din1(g246_p_spl_),
    .din2(g366_n_spl_010)
  );


  LA
  g_g500_p
  (
    .dout(g500_p),
    .din1(g498_n),
    .din2(g499_n)
  );


  FA
  g_g500_n
  (
    .dout(g500_n),
    .din1(g498_p),
    .din2(g499_p)
  );


  LA
  g_g501_p
  (
    .dout(g501_p),
    .din1(G47_p_spl_01),
    .din2(g500_p_spl_0)
  );


  FA
  g_g501_n
  (
    .dout(g501_n),
    .din1(G47_n_spl_01),
    .din2(g500_n_spl_0)
  );


  LA
  g_g502_p
  (
    .dout(g502_p),
    .din1(g379_p_spl_00),
    .din2(g456_n_spl_0)
  );


  FA
  g_g502_n
  (
    .dout(g502_n),
    .din1(g379_n_spl_00),
    .din2(g456_p_spl_0)
  );


  LA
  g_g503_p
  (
    .dout(g503_p),
    .din1(g379_n_spl_00),
    .din2(g456_p_spl_1)
  );


  FA
  g_g503_n
  (
    .dout(g503_n),
    .din1(g379_p_spl_01),
    .din2(g456_n_spl_1)
  );


  LA
  g_g504_p
  (
    .dout(g504_p),
    .din1(g502_n),
    .din2(g503_n_spl_)
  );


  FA
  g_g504_n
  (
    .dout(g504_n),
    .din1(g502_p),
    .din2(g503_p_spl_)
  );


  LA
  g_g505_p
  (
    .dout(g505_p),
    .din1(g501_p_spl_),
    .din2(g504_p_spl_)
  );


  FA
  g_g505_n
  (
    .dout(g505_n),
    .din1(g501_n_spl_),
    .din2(g504_n_spl_)
  );


  LA
  g_g506_p
  (
    .dout(g506_p),
    .din1(g501_n_spl_),
    .din2(g504_n_spl_)
  );


  FA
  g_g506_n
  (
    .dout(g506_n),
    .din1(g501_p_spl_),
    .din2(g504_p_spl_)
  );


  LA
  g_g507_p
  (
    .dout(g507_p),
    .din1(g505_n),
    .din2(g506_n)
  );


  FA
  g_g507_n
  (
    .dout(g507_n),
    .din1(g505_p),
    .din2(g506_p)
  );


  LA
  g_g508_p
  (
    .dout(g508_p),
    .din1(g385_n_spl_001),
    .din2(g507_n)
  );


  FA
  g_g508_n
  (
    .dout(g508_n),
    .din1(g385_p_spl_001),
    .din2(g507_p)
  );


  LA
  g_g509_p
  (
    .dout(g509_p),
    .din1(g488_n),
    .din2(g508_n)
  );


  FA
  g_g509_n
  (
    .dout(g509_n),
    .din1(g488_p),
    .din2(g508_p)
  );


  LA
  g_g510_p
  (
    .dout(g510_p),
    .din1(g282_n_spl_),
    .din2(g366_p_spl_011)
  );


  FA
  g_g510_n
  (
    .dout(g510_n),
    .din1(g282_p_spl_),
    .din2(g366_n_spl_011)
  );


  LA
  g_g511_p
  (
    .dout(g511_p),
    .din1(g296_n_spl_0),
    .din2(g510_n_spl_)
  );


  FA
  g_g511_n
  (
    .dout(g511_n),
    .din1(g296_p_spl_0),
    .din2(g510_p_spl_)
  );


  LA
  g_g512_p
  (
    .dout(g512_p),
    .din1(g296_p_spl_),
    .din2(g510_p_spl_)
  );


  FA
  g_g512_n
  (
    .dout(g512_n),
    .din1(g296_n_spl_),
    .din2(g510_n_spl_)
  );


  LA
  g_g513_p
  (
    .dout(g513_p),
    .din1(g511_n),
    .din2(g512_n)
  );


  FA
  g_g513_n
  (
    .dout(g513_n),
    .din1(g511_p),
    .din2(g512_p)
  );


  LA
  g_g514_p
  (
    .dout(g514_p),
    .din1(g332_n_spl_),
    .din2(g365_p_spl_0)
  );


  FA
  g_g514_n
  (
    .dout(g514_n),
    .din1(g332_p_spl_),
    .din2(g365_n_spl_0)
  );


  LA
  g_g515_p
  (
    .dout(g515_p),
    .din1(g346_n_spl_0),
    .din2(g514_n_spl_)
  );


  FA
  g_g515_n
  (
    .dout(g515_n),
    .din1(g346_p_spl_0),
    .din2(g514_p_spl_)
  );


  LA
  g_g516_p
  (
    .dout(g516_p),
    .din1(g346_p_spl_),
    .din2(g514_p_spl_)
  );


  FA
  g_g516_n
  (
    .dout(g516_n),
    .din1(g346_n_spl_),
    .din2(g514_n_spl_)
  );


  LA
  g_g517_p
  (
    .dout(g517_p),
    .din1(g515_n),
    .din2(g516_n)
  );


  FA
  g_g517_n
  (
    .dout(g517_n),
    .din1(g515_p),
    .din2(g516_p)
  );


  LA
  g_g518_p
  (
    .dout(g518_p),
    .din1(g513_p_spl_00),
    .din2(g517_p_spl_00)
  );


  FA
  g_g518_n
  (
    .dout(g518_n),
    .din1(g513_n_spl_00),
    .din2(g517_n_spl_00)
  );


  LA
  g_g519_p
  (
    .dout(g519_p),
    .din1(g456_p_spl_1),
    .din2(g500_n_spl_0)
  );


  FA
  g_g519_n
  (
    .dout(g519_n),
    .din1(g456_n_spl_1),
    .din2(g500_p_spl_0)
  );


  LA
  g_g520_p
  (
    .dout(g520_p),
    .din1(g518_p_spl_),
    .din2(g519_p_spl_)
  );


  FA
  g_g520_n
  (
    .dout(g520_n),
    .din1(g518_n_spl_),
    .din2(g519_n_spl_)
  );


  LA
  g_g521_p
  (
    .dout(g521_p),
    .din1(g349_n_spl_),
    .din2(g500_n_spl_)
  );


  FA
  g_g521_n
  (
    .dout(g521_n),
    .din1(g349_p_spl_1),
    .din2(g500_p_spl_)
  );


  LA
  g_g522_p
  (
    .dout(g522_p),
    .din1(g520_n_spl_),
    .din2(g521_p_spl_0)
  );


  FA
  g_g522_n
  (
    .dout(g522_n),
    .din1(g520_p_spl_),
    .din2(g521_n_spl_0)
  );


  LA
  g_g523_p
  (
    .dout(g523_p),
    .din1(g520_p_spl_),
    .din2(g521_n_spl_0)
  );


  FA
  g_g523_n
  (
    .dout(g523_n),
    .din1(g520_n_spl_),
    .din2(g521_p_spl_0)
  );


  LA
  g_g524_p
  (
    .dout(g524_p),
    .din1(g522_n),
    .din2(g523_n)
  );


  FA
  g_g524_n
  (
    .dout(g524_n),
    .din1(g522_p),
    .din2(g523_p)
  );


  LA
  g_g525_p
  (
    .dout(g525_p),
    .din1(G47_p_spl_10),
    .din2(g524_n)
  );


  FA
  g_g525_n
  (
    .dout(g525_n),
    .din1(G47_n_spl_10),
    .din2(g524_p)
  );


  LA
  g_g526_p
  (
    .dout(g526_p),
    .din1(g349_n_spl_),
    .din2(g379_n_spl_01)
  );


  FA
  g_g526_n
  (
    .dout(g526_n),
    .din1(g349_p_spl_1),
    .din2(g379_p_spl_01)
  );


  LA
  g_g527_p
  (
    .dout(g527_p),
    .din1(g363_p),
    .din2(g526_n)
  );


  FA
  g_g527_n
  (
    .dout(g527_n),
    .din1(g363_n_spl_),
    .din2(g526_p)
  );


  LA
  g_g528_p
  (
    .dout(g528_p),
    .din1(g295_p_spl_),
    .din2(g366_n_spl_011)
  );


  FA
  g_g528_n
  (
    .dout(g528_n),
    .din1(g295_n_spl_),
    .din2(g366_p_spl_011)
  );


  LA
  g_g529_p
  (
    .dout(g529_p),
    .din1(g517_p_spl_00),
    .din2(g528_p_spl_)
  );


  FA
  g_g529_n
  (
    .dout(g529_n),
    .din1(g517_n_spl_00),
    .din2(g528_n_spl_)
  );


  LA
  g_g530_p
  (
    .dout(g530_p),
    .din1(g273_p_spl_),
    .din2(g366_n_spl_100)
  );


  FA
  g_g530_n
  (
    .dout(g530_n),
    .din1(g273_n_spl_),
    .din2(g366_p_spl_100)
  );


  LA
  g_g531_p
  (
    .dout(g531_p),
    .din1(g518_p_spl_),
    .din2(g530_n_spl_0)
  );


  FA
  g_g531_n
  (
    .dout(g531_n),
    .din1(g518_n_spl_),
    .din2(g530_p_spl_0)
  );


  LA
  g_g532_p
  (
    .dout(g532_p),
    .din1(g345_p_spl_),
    .din2(g365_n_spl_1)
  );


  FA
  g_g532_n
  (
    .dout(g532_n),
    .din1(g345_n_spl_),
    .din2(g365_p_spl_1)
  );


  LA
  g_g533_p
  (
    .dout(g533_p),
    .din1(g531_n),
    .din2(g532_n)
  );


  FA
  g_g533_n
  (
    .dout(g533_n),
    .din1(g531_p),
    .din2(g532_p)
  );


  LA
  g_g534_p
  (
    .dout(g534_p),
    .din1(g529_n),
    .din2(g533_p)
  );


  FA
  g_g534_n
  (
    .dout(g534_n),
    .din1(g529_p),
    .din2(g533_n)
  );


  LA
  g_g535_p
  (
    .dout(g535_p),
    .din1(g527_n_spl_0),
    .din2(g534_n_spl_0)
  );


  FA
  g_g535_n
  (
    .dout(g535_n),
    .din1(g527_p_spl_0),
    .din2(g534_p_spl_0)
  );


  LA
  g_g536_p
  (
    .dout(g536_p),
    .din1(g527_p_spl_0),
    .din2(g534_p_spl_0)
  );


  FA
  g_g536_n
  (
    .dout(g536_n),
    .din1(g527_n_spl_0),
    .din2(g534_n_spl_0)
  );


  LA
  g_g537_p
  (
    .dout(g537_p),
    .din1(g535_n),
    .din2(g536_n)
  );


  FA
  g_g537_n
  (
    .dout(g537_n),
    .din1(g535_p),
    .din2(g536_p)
  );


  LA
  g_g538_p
  (
    .dout(g538_p),
    .din1(g525_p),
    .din2(g537_n)
  );


  LA
  g_g539_p
  (
    .dout(g539_p),
    .din1(g525_n),
    .din2(g537_p)
  );


  FA
  g_g540_n
  (
    .dout(g540_n),
    .din1(g538_p),
    .din2(g539_p)
  );


  LA
  g_g541_p
  (
    .dout(g541_p),
    .din1(g74_n_spl_),
    .din2(g78_n_spl_)
  );


  LA
  g_g542_p
  (
    .dout(g542_p),
    .din1(g540_n),
    .din2(g541_p)
  );


  LA
  g_g543_p
  (
    .dout(g543_p),
    .din1(G10_n_spl_101),
    .din2(g326_n_spl_)
  );


  FA
  g_g544_n
  (
    .dout(g544_n),
    .din1(G7_p_spl_011),
    .din2(g543_p)
  );


  FA
  g_g545_n
  (
    .dout(g545_n),
    .din1(G7_n_spl_011),
    .din2(G9_n_spl_101)
  );


  LA
  g_g546_p
  (
    .dout(g546_p),
    .din1(g78_p_spl_),
    .din2(g545_n)
  );


  LA
  g_g547_p
  (
    .dout(g547_p),
    .din1(g544_n),
    .din2(g546_p)
  );


  LA
  g_g548_p
  (
    .dout(g548_p),
    .din1(G14_n_spl_100),
    .din2(g74_p)
  );


  LA
  g_g549_p
  (
    .dout(g549_p),
    .din1(g223_n_spl_),
    .din2(g548_p)
  );


  FA
  g_g550_n
  (
    .dout(g550_n),
    .din1(g547_p),
    .din2(g549_p)
  );


  FA
  g_g551_n
  (
    .dout(g551_n),
    .din1(g542_p),
    .din2(g550_n)
  );


  LA
  g_g552_p
  (
    .dout(g552_p),
    .din1(g202_n_spl_),
    .din2(g366_p_spl_100)
  );


  FA
  g_g552_n
  (
    .dout(g552_n),
    .din1(g202_p_spl_),
    .din2(g366_n_spl_100)
  );


  LA
  g_g553_p
  (
    .dout(g553_p),
    .din1(g217_n_spl_1),
    .din2(g552_n_spl_)
  );


  FA
  g_g553_n
  (
    .dout(g553_n),
    .din1(g217_p_spl_1),
    .din2(g552_p_spl_)
  );


  LA
  g_g554_p
  (
    .dout(g554_p),
    .din1(g217_p_spl_1),
    .din2(g552_p_spl_)
  );


  FA
  g_g554_n
  (
    .dout(g554_n),
    .din1(g217_n_spl_1),
    .din2(g552_n_spl_)
  );


  LA
  g_g555_p
  (
    .dout(g555_p),
    .din1(g553_n),
    .din2(g554_n)
  );


  FA
  g_g555_n
  (
    .dout(g555_n),
    .din1(g553_p),
    .din2(g554_p)
  );


  LA
  g_g556_p
  (
    .dout(g556_p),
    .din1(g390_p_spl_0),
    .din2(g555_p_spl_0)
  );


  FA
  g_g556_n
  (
    .dout(g556_n),
    .din1(g390_n_spl_0),
    .din2(g555_n_spl_0)
  );


  LA
  g_g557_p
  (
    .dout(g557_p),
    .din1(G11_p_spl_101),
    .din2(g394_n_spl_01)
  );


  FA
  g_g557_n
  (
    .dout(g557_n),
    .din1(G11_n_spl_10),
    .din2(g394_p_spl_01)
  );


  LA
  g_g558_p
  (
    .dout(g558_p),
    .din1(g393_p_spl_010),
    .din2(g557_n)
  );


  FA
  g_g558_n
  (
    .dout(g558_n),
    .din1(g393_n_spl_010),
    .din2(g557_p)
  );


  LA
  g_g559_p
  (
    .dout(g559_p),
    .din1(g385_p_spl_01),
    .din2(g558_n)
  );


  FA
  g_g559_n
  (
    .dout(g559_n),
    .din1(g385_n_spl_01),
    .din2(g558_p)
  );


  LA
  g_g560_p
  (
    .dout(g560_p),
    .din1(G41_p_spl_01),
    .din2(g409_n_spl_010)
  );


  FA
  g_g560_n
  (
    .dout(g560_n),
    .din1(G41_n_spl_01),
    .din2(g409_p_spl_010)
  );


  LA
  g_g561_p
  (
    .dout(g561_p),
    .din1(G42_p_spl_0),
    .din2(g406_n_spl_010)
  );


  FA
  g_g561_n
  (
    .dout(g561_n),
    .din1(G42_n_spl_0),
    .din2(g406_p_spl_010)
  );


  LA
  g_g562_p
  (
    .dout(g562_p),
    .din1(G4_p_spl_1011),
    .din2(g561_n)
  );


  FA
  g_g562_n
  (
    .dout(g562_n),
    .din1(G4_n_spl_1011),
    .din2(g561_p)
  );


  LA
  g_g563_p
  (
    .dout(g563_p),
    .din1(g560_n),
    .din2(g562_p)
  );


  FA
  g_g563_n
  (
    .dout(g563_n),
    .din1(g560_p),
    .din2(g562_n)
  );


  LA
  g_g564_p
  (
    .dout(g564_p),
    .din1(G13_n_spl_101),
    .din2(g423_n_spl_001)
  );


  FA
  g_g564_n
  (
    .dout(g564_n),
    .din1(G13_p_spl_110),
    .din2(g423_p_spl_001)
  );


  LA
  g_g565_p
  (
    .dout(g565_p),
    .din1(G14_n_spl_100),
    .din2(g425_n_spl_010)
  );


  FA
  g_g565_n
  (
    .dout(g565_n),
    .din1(G14_p_spl_100),
    .din2(g425_p_spl_010)
  );


  LA
  g_g566_p
  (
    .dout(g566_p),
    .din1(g564_n),
    .din2(g565_n)
  );


  FA
  g_g566_n
  (
    .dout(g566_n),
    .din1(g564_p),
    .din2(g565_p)
  );


  LA
  g_g567_p
  (
    .dout(g567_p),
    .din1(G39_n_spl_01),
    .din2(G43_n_spl_0)
  );


  FA
  g_g567_n
  (
    .dout(g567_n),
    .din1(G39_p_spl_01),
    .din2(G43_p_spl_0)
  );


  LA
  g_g568_p
  (
    .dout(g568_p),
    .din1(g412_n_spl_001),
    .din2(g567_n)
  );


  FA
  g_g568_n
  (
    .dout(g568_n),
    .din1(g412_p_spl_001),
    .din2(g567_p)
  );


  LA
  g_g569_p
  (
    .dout(g569_p),
    .din1(G12_p_spl_101),
    .din2(G40_n_spl_01)
  );


  FA
  g_g569_n
  (
    .dout(g569_n),
    .din1(G12_n_spl_101),
    .din2(G40_p_spl_01)
  );


  LA
  g_g570_p
  (
    .dout(g570_p),
    .din1(g414_n_spl_010),
    .din2(g569_n_spl_)
  );


  FA
  g_g570_n
  (
    .dout(g570_n),
    .din1(g414_p_spl_010),
    .din2(g569_p_spl_)
  );


  LA
  g_g571_p
  (
    .dout(g571_p),
    .din1(g568_n),
    .din2(g570_n)
  );


  FA
  g_g571_n
  (
    .dout(g571_n),
    .din1(g568_p),
    .din2(g570_p)
  );


  LA
  g_g572_p
  (
    .dout(g572_p),
    .din1(g566_p),
    .din2(g571_p)
  );


  FA
  g_g572_n
  (
    .dout(g572_n),
    .din1(g566_n),
    .din2(g571_n)
  );


  LA
  g_g573_p
  (
    .dout(g573_p),
    .din1(g563_p),
    .din2(g572_p)
  );


  FA
  g_g573_n
  (
    .dout(g573_n),
    .din1(g563_n),
    .din2(g572_n)
  );


  LA
  g_g574_p
  (
    .dout(g574_p),
    .din1(G8_n_spl_101),
    .din2(g425_n_spl_010)
  );


  FA
  g_g574_n
  (
    .dout(g574_n),
    .din1(G8_p_spl_101),
    .din2(g425_p_spl_010)
  );


  LA
  g_g575_p
  (
    .dout(g575_p),
    .din1(G7_n_spl_100),
    .din2(g412_n_spl_010)
  );


  FA
  g_g575_n
  (
    .dout(g575_n),
    .din1(G7_p_spl_100),
    .din2(g412_p_spl_010)
  );


  LA
  g_g576_p
  (
    .dout(g576_p),
    .din1(G10_n_spl_101),
    .din2(g414_n_spl_010)
  );


  FA
  g_g576_n
  (
    .dout(g576_n),
    .din1(G10_p_spl_101),
    .din2(g414_p_spl_010)
  );


  LA
  g_g577_p
  (
    .dout(g577_p),
    .din1(g575_n),
    .din2(g576_n)
  );


  FA
  g_g577_n
  (
    .dout(g577_n),
    .din1(g575_p),
    .din2(g576_p)
  );


  LA
  g_g578_p
  (
    .dout(g578_p),
    .din1(g574_n),
    .din2(g577_p)
  );


  FA
  g_g578_n
  (
    .dout(g578_n),
    .din1(g574_p),
    .din2(g577_n)
  );


  LA
  g_g579_p
  (
    .dout(g579_p),
    .din1(G9_n_spl_101),
    .din2(g423_n_spl_010)
  );


  FA
  g_g579_n
  (
    .dout(g579_n),
    .din1(G9_p_spl_101),
    .din2(g423_p_spl_010)
  );


  LA
  g_g580_p
  (
    .dout(g580_p),
    .din1(G20_p_spl_00),
    .din2(g406_n_spl_010)
  );


  FA
  g_g580_n
  (
    .dout(g580_n),
    .din1(G20_n_spl_00),
    .din2(g406_p_spl_010)
  );


  LA
  g_g581_p
  (
    .dout(g581_p),
    .din1(G21_p_spl_01),
    .din2(g409_n_spl_010)
  );


  FA
  g_g581_n
  (
    .dout(g581_n),
    .din1(G21_n_spl_01),
    .din2(g409_p_spl_010)
  );


  LA
  g_g582_p
  (
    .dout(g582_p),
    .din1(g580_n),
    .din2(g581_n)
  );


  FA
  g_g582_n
  (
    .dout(g582_n),
    .din1(g580_p),
    .din2(g581_p)
  );


  LA
  g_g583_p
  (
    .dout(g583_p),
    .din1(g579_n_spl_),
    .din2(g582_p)
  );


  FA
  g_g583_n
  (
    .dout(g583_n),
    .din1(g579_p_spl_),
    .din2(g582_n)
  );


  LA
  g_g584_p
  (
    .dout(g584_p),
    .din1(G19_p_spl_00),
    .din2(g412_n_spl_010)
  );


  FA
  g_g584_n
  (
    .dout(g584_n),
    .din1(G19_n_spl_00),
    .din2(g412_p_spl_010)
  );


  LA
  g_g585_p
  (
    .dout(g585_p),
    .din1(G22_p_spl_01),
    .din2(g414_n_spl_011)
  );


  FA
  g_g585_n
  (
    .dout(g585_n),
    .din1(G22_n_spl_01),
    .din2(g414_p_spl_011)
  );


  LA
  g_g586_p
  (
    .dout(g586_p),
    .din1(g584_n),
    .din2(g585_n)
  );


  FA
  g_g586_n
  (
    .dout(g586_n),
    .din1(g584_p),
    .din2(g585_p)
  );


  LA
  g_g587_p
  (
    .dout(g587_p),
    .din1(G4_n_spl_1100),
    .din2(g586_p)
  );


  FA
  g_g587_n
  (
    .dout(g587_n),
    .din1(G4_p_spl_1100),
    .din2(g586_n)
  );


  LA
  g_g588_p
  (
    .dout(g588_p),
    .din1(g583_p),
    .din2(g587_p)
  );


  FA
  g_g588_n
  (
    .dout(g588_n),
    .din1(g583_n),
    .din2(g587_n)
  );


  LA
  g_g589_p
  (
    .dout(g589_p),
    .din1(g578_p),
    .din2(g588_p)
  );


  FA
  g_g589_n
  (
    .dout(g589_n),
    .din1(g578_n),
    .din2(g588_n)
  );


  LA
  g_g590_p
  (
    .dout(g590_p),
    .din1(g573_n),
    .din2(g589_n)
  );


  FA
  g_g590_n
  (
    .dout(g590_n),
    .din1(g573_p),
    .din2(g589_p)
  );


  LA
  g_g591_p
  (
    .dout(g591_p),
    .din1(g393_n_spl_010),
    .din2(g590_n)
  );


  FA
  g_g591_n
  (
    .dout(g591_n),
    .din1(g393_p_spl_010),
    .din2(g590_p)
  );


  LA
  g_g592_p
  (
    .dout(g592_p),
    .din1(g559_p),
    .din2(g591_n)
  );


  FA
  g_g592_n
  (
    .dout(g592_n),
    .din1(g559_n),
    .din2(g591_p)
  );


  LA
  g_g593_p
  (
    .dout(g593_p),
    .din1(g556_n),
    .din2(g592_p)
  );


  FA
  g_g593_n
  (
    .dout(g593_n),
    .din1(g556_p),
    .din2(g592_n)
  );


  LA
  g_g594_p
  (
    .dout(g594_p),
    .din1(g229_n_spl_),
    .din2(g366_p_spl_101)
  );


  FA
  g_g594_n
  (
    .dout(g594_n),
    .din1(g229_p_spl_),
    .din2(g366_n_spl_101)
  );


  LA
  g_g595_p
  (
    .dout(g595_p),
    .din1(g243_n_spl_0),
    .din2(g594_n_spl_)
  );


  FA
  g_g595_n
  (
    .dout(g595_n),
    .din1(g243_p_spl_0),
    .din2(g594_p_spl_)
  );


  LA
  g_g596_p
  (
    .dout(g596_p),
    .din1(g243_p_spl_),
    .din2(g594_p_spl_)
  );


  FA
  g_g596_n
  (
    .dout(g596_n),
    .din1(g243_n_spl_),
    .din2(g594_n_spl_)
  );


  LA
  g_g597_p
  (
    .dout(g597_p),
    .din1(g595_n),
    .din2(g596_n)
  );


  FA
  g_g597_n
  (
    .dout(g597_n),
    .din1(g595_p),
    .din2(g596_p)
  );


  LA
  g_g598_p
  (
    .dout(g598_p),
    .din1(g376_p_spl_0),
    .din2(g597_n_spl_00)
  );


  FA
  g_g598_n
  (
    .dout(g598_n),
    .din1(g376_n_spl_),
    .din2(g597_p_spl_00)
  );


  LA
  g_g599_p
  (
    .dout(g599_p),
    .din1(g242_p_spl_),
    .din2(g366_n_spl_101)
  );


  FA
  g_g599_n
  (
    .dout(g599_n),
    .din1(g242_n_spl_),
    .din2(g366_p_spl_101)
  );


  LA
  g_g600_p
  (
    .dout(g600_p),
    .din1(g167_p_spl_),
    .din2(g366_n_spl_11)
  );


  FA
  g_g600_n
  (
    .dout(g600_n),
    .din1(g167_n_spl_),
    .din2(g366_p_spl_11)
  );


  LA
  g_g601_p
  (
    .dout(g601_p),
    .din1(g370_n_spl_0),
    .din2(g600_n_spl_)
  );


  FA
  g_g601_n
  (
    .dout(g601_n),
    .din1(g370_p_spl_0),
    .din2(g600_p_spl_)
  );


  LA
  g_g602_p
  (
    .dout(g602_p),
    .din1(g190_p_spl_),
    .din2(g366_n_spl_11)
  );


  FA
  g_g602_n
  (
    .dout(g602_n),
    .din1(g190_n_spl_),
    .din2(g366_p_spl_11)
  );


  LA
  g_g603_p
  (
    .dout(g603_p),
    .din1(g601_n_spl_),
    .din2(g602_n)
  );


  FA
  g_g603_n
  (
    .dout(g603_n),
    .din1(g601_p_spl_),
    .din2(g602_p)
  );


  LA
  g_g604_p
  (
    .dout(g604_p),
    .din1(g597_n_spl_00),
    .din2(g603_n_spl_)
  );


  FA
  g_g604_n
  (
    .dout(g604_n),
    .din1(g597_p_spl_00),
    .din2(g603_p_spl_)
  );


  LA
  g_g605_p
  (
    .dout(g605_p),
    .din1(g599_n),
    .din2(g604_n)
  );


  FA
  g_g605_n
  (
    .dout(g605_n),
    .din1(g599_p),
    .din2(g604_p)
  );


  LA
  g_g606_p
  (
    .dout(g606_p),
    .din1(g555_n_spl_0),
    .din2(g605_p_spl_)
  );


  FA
  g_g606_n
  (
    .dout(g606_n),
    .din1(g555_p_spl_0),
    .din2(g605_n_spl_)
  );


  LA
  g_g607_p
  (
    .dout(g607_p),
    .din1(g555_p_spl_),
    .din2(g605_n_spl_)
  );


  FA
  g_g607_n
  (
    .dout(g607_n),
    .din1(g555_n_spl_),
    .din2(g605_p_spl_)
  );


  LA
  g_g608_p
  (
    .dout(g608_p),
    .din1(g606_n),
    .din2(g607_n)
  );


  FA
  g_g608_n
  (
    .dout(g608_n),
    .din1(g606_p),
    .din2(g607_p)
  );


  LA
  g_g609_p
  (
    .dout(g609_p),
    .din1(g598_n_spl_),
    .din2(g608_n_spl_)
  );


  FA
  g_g609_n
  (
    .dout(g609_n),
    .din1(g598_p_spl_),
    .din2(g608_p_spl_)
  );


  LA
  g_g610_p
  (
    .dout(g610_p),
    .din1(g598_p_spl_),
    .din2(g608_p_spl_)
  );


  FA
  g_g610_n
  (
    .dout(g610_n),
    .din1(g598_n_spl_),
    .din2(g608_n_spl_)
  );


  LA
  g_g611_p
  (
    .dout(g611_p),
    .din1(g609_n),
    .din2(g610_n)
  );


  FA
  g_g611_n
  (
    .dout(g611_n),
    .din1(g609_p),
    .din2(g610_p)
  );


  LA
  g_g612_p
  (
    .dout(g612_p),
    .din1(g370_p_spl_1),
    .din2(g600_p_spl_)
  );


  FA
  g_g612_n
  (
    .dout(g612_n),
    .din1(g370_n_spl_1),
    .din2(g600_n_spl_)
  );


  LA
  g_g613_p
  (
    .dout(g613_p),
    .din1(g601_n_spl_),
    .din2(g612_n)
  );


  FA
  g_g613_n
  (
    .dout(g613_n),
    .din1(g601_p_spl_),
    .din2(g612_p)
  );


  LA
  g_g614_p
  (
    .dout(g614_p),
    .din1(g387_n_spl_0),
    .din2(g613_n_spl_)
  );


  FA
  g_g614_n
  (
    .dout(g614_n),
    .din1(g387_p_spl_0),
    .din2(g613_p_spl_)
  );


  LA
  g_g615_p
  (
    .dout(g615_p),
    .din1(g387_p_spl_),
    .din2(g613_p_spl_)
  );


  FA
  g_g615_n
  (
    .dout(g615_n),
    .din1(g387_n_spl_),
    .din2(g613_n_spl_)
  );


  LA
  g_g616_p
  (
    .dout(g616_p),
    .din1(g614_n),
    .din2(g615_n)
  );


  FA
  g_g616_n
  (
    .dout(g616_n),
    .din1(g614_p),
    .din2(g615_p)
  );


  LA
  g_g617_p
  (
    .dout(g617_p),
    .din1(g376_n_spl_),
    .din2(g603_n_spl_)
  );


  FA
  g_g617_n
  (
    .dout(g617_n),
    .din1(g376_p_spl_0),
    .din2(g603_p_spl_)
  );


  LA
  g_g618_p
  (
    .dout(g618_p),
    .din1(g597_p_spl_0),
    .din2(g617_p_spl_)
  );


  FA
  g_g618_n
  (
    .dout(g618_n),
    .din1(g597_n_spl_0),
    .din2(g617_n_spl_)
  );


  LA
  g_g619_p
  (
    .dout(g619_p),
    .din1(g597_n_spl_1),
    .din2(g617_n_spl_)
  );


  FA
  g_g619_n
  (
    .dout(g619_n),
    .din1(g597_p_spl_1),
    .din2(g617_p_spl_)
  );


  LA
  g_g620_p
  (
    .dout(g620_p),
    .din1(g618_n),
    .din2(g619_n)
  );


  FA
  g_g620_n
  (
    .dout(g620_n),
    .din1(g618_p),
    .din2(g619_p)
  );


  LA
  g_g621_p
  (
    .dout(g621_p),
    .din1(g616_n_spl_0),
    .din2(g620_n_spl_0)
  );


  FA
  g_g621_n
  (
    .dout(g621_n),
    .din1(g616_p_spl_0),
    .din2(g620_p_spl_0)
  );


  LA
  g_g622_p
  (
    .dout(g622_p),
    .din1(g379_p_spl_10),
    .din2(g621_n)
  );


  FA
  g_g622_n
  (
    .dout(g622_n),
    .din1(g379_n_spl_01),
    .din2(g621_p)
  );


  LA
  g_g623_p
  (
    .dout(g623_p),
    .din1(g377_n_spl_01),
    .din2(g622_n)
  );


  FA
  g_g623_n
  (
    .dout(g623_n),
    .din1(g377_p_spl_00),
    .din2(g622_p)
  );


  LA
  g_g624_p
  (
    .dout(g624_p),
    .din1(g384_p_spl_00),
    .din2(g623_n)
  );


  FA
  g_g624_n
  (
    .dout(g624_n),
    .din1(g384_n_spl_00),
    .din2(g623_p)
  );


  LA
  g_g625_p
  (
    .dout(g625_p),
    .din1(g611_n),
    .din2(g624_n)
  );


  FA
  g_g625_n
  (
    .dout(g625_n),
    .din1(g611_p),
    .din2(g624_p)
  );


  LA
  g_g626_p
  (
    .dout(g626_p),
    .din1(g593_n),
    .din2(g625_n)
  );


  FA
  g_g626_n
  (
    .dout(g626_n),
    .din1(g593_p),
    .din2(g625_p)
  );


  LA
  g_g627_p
  (
    .dout(g627_p),
    .din1(g379_p_spl_10),
    .din2(g616_p_spl_0)
  );


  FA
  g_g627_n
  (
    .dout(g627_n),
    .din1(g379_n_spl_1),
    .din2(g616_n_spl_0)
  );


  LA
  g_g628_p
  (
    .dout(g628_p),
    .din1(g379_n_spl_1),
    .din2(g616_n_spl_1)
  );


  FA
  g_g628_n
  (
    .dout(g628_n),
    .din1(g379_p_spl_1),
    .din2(g616_p_spl_1)
  );


  LA
  g_g629_p
  (
    .dout(g629_p),
    .din1(g627_n),
    .din2(g628_n_spl_0)
  );


  FA
  g_g629_n
  (
    .dout(g629_n),
    .din1(g627_p),
    .din2(g628_p_spl_0)
  );


  LA
  g_g630_p
  (
    .dout(g630_p),
    .din1(g377_n_spl_01),
    .din2(g629_p)
  );


  FA
  g_g630_n
  (
    .dout(g630_n),
    .din1(g377_p_spl_01),
    .din2(g629_n)
  );


  LA
  g_g631_p
  (
    .dout(g631_p),
    .din1(g384_n_spl_01),
    .din2(g616_n_spl_1)
  );


  FA
  g_g631_n
  (
    .dout(g631_n),
    .din1(g384_p_spl_01),
    .din2(g616_p_spl_1)
  );


  LA
  g_g632_p
  (
    .dout(g632_p),
    .din1(G39_p_spl_01),
    .din2(g423_n_spl_010)
  );


  FA
  g_g632_n
  (
    .dout(g632_n),
    .din1(G39_n_spl_01),
    .din2(g423_p_spl_010)
  );


  LA
  g_g633_p
  (
    .dout(g633_p),
    .din1(G40_p_spl_10),
    .din2(g425_n_spl_011)
  );


  FA
  g_g633_n
  (
    .dout(g633_n),
    .din1(G40_n_spl_10),
    .din2(g425_p_spl_011)
  );


  LA
  g_g634_p
  (
    .dout(g634_p),
    .din1(g632_n),
    .din2(g633_n)
  );


  FA
  g_g634_n
  (
    .dout(g634_n),
    .din1(g632_p),
    .din2(g633_p)
  );


  LA
  g_g635_p
  (
    .dout(g635_p),
    .din1(G43_p_spl_1),
    .din2(g409_n_spl_011)
  );


  FA
  g_g635_n
  (
    .dout(g635_n),
    .din1(G43_n_spl_1),
    .din2(g409_p_spl_011)
  );


  LA
  g_g636_p
  (
    .dout(g636_p),
    .din1(G44_p_spl_0),
    .din2(g406_n_spl_011)
  );


  FA
  g_g636_n
  (
    .dout(g636_n),
    .din1(G44_n_spl_0),
    .din2(g406_p_spl_011)
  );


  LA
  g_g637_p
  (
    .dout(g637_p),
    .din1(G4_p_spl_1100),
    .din2(g636_n)
  );


  FA
  g_g637_n
  (
    .dout(g637_n),
    .din1(G4_n_spl_1100),
    .din2(g636_p)
  );


  LA
  g_g638_p
  (
    .dout(g638_p),
    .din1(g635_n),
    .din2(g637_p)
  );


  FA
  g_g638_n
  (
    .dout(g638_n),
    .din1(g635_p),
    .din2(g637_n)
  );


  LA
  g_g639_p
  (
    .dout(g639_p),
    .din1(g634_p),
    .din2(g638_p)
  );


  FA
  g_g639_n
  (
    .dout(g639_n),
    .din1(g634_n),
    .din2(g638_n)
  );


  LA
  g_g640_p
  (
    .dout(g640_p),
    .din1(G41_n_spl_10),
    .din2(G45_n_spl_)
  );


  FA
  g_g640_n
  (
    .dout(g640_n),
    .din1(G41_p_spl_10),
    .din2(G45_p_spl_)
  );


  LA
  g_g641_p
  (
    .dout(g641_p),
    .din1(g412_n_spl_011),
    .din2(g640_n)
  );


  FA
  g_g641_n
  (
    .dout(g641_n),
    .din1(g412_p_spl_011),
    .din2(g640_p)
  );


  LA
  g_g642_p
  (
    .dout(g642_p),
    .din1(G14_p_spl_101),
    .din2(G42_n_spl_1)
  );


  FA
  g_g642_n
  (
    .dout(g642_n),
    .din1(G14_n_spl_101),
    .din2(G42_p_spl_1)
  );


  LA
  g_g643_p
  (
    .dout(g643_p),
    .din1(g414_n_spl_011),
    .din2(g642_n)
  );


  FA
  g_g643_n
  (
    .dout(g643_n),
    .din1(g414_p_spl_011),
    .din2(g642_p)
  );


  LA
  g_g644_p
  (
    .dout(g644_p),
    .din1(g641_n),
    .din2(g643_n)
  );


  FA
  g_g644_n
  (
    .dout(g644_n),
    .din1(g641_p),
    .din2(g643_p)
  );


  LA
  g_g645_p
  (
    .dout(g645_p),
    .din1(g639_p),
    .din2(g644_p)
  );


  FA
  g_g645_n
  (
    .dout(g645_n),
    .din1(g639_n),
    .din2(g644_n)
  );


  LA
  g_g646_p
  (
    .dout(g646_p),
    .din1(G12_n_spl_101),
    .din2(g414_n_spl_100)
  );


  FA
  g_g646_n
  (
    .dout(g646_n),
    .din1(G12_p_spl_110),
    .din2(g414_p_spl_100)
  );


  LA
  g_g647_p
  (
    .dout(g647_p),
    .din1(G10_n_spl_110),
    .din2(g425_n_spl_011)
  );


  FA
  g_g647_n
  (
    .dout(g647_n),
    .din1(G10_p_spl_101),
    .din2(g425_p_spl_011)
  );


  LA
  g_g648_p
  (
    .dout(g648_p),
    .din1(g646_n),
    .din2(g647_n)
  );


  FA
  g_g648_n
  (
    .dout(g648_n),
    .din1(g646_p),
    .din2(g647_p)
  );


  LA
  g_g649_p
  (
    .dout(g649_p),
    .din1(G4_n_spl_1101),
    .din2(g648_p)
  );


  FA
  g_g649_n
  (
    .dout(g649_n),
    .din1(G4_p_spl_1101),
    .din2(g648_n)
  );


  LA
  g_g650_p
  (
    .dout(g650_p),
    .din1(G22_p_spl_01),
    .din2(g406_n_spl_011)
  );


  FA
  g_g650_n
  (
    .dout(g650_n),
    .din1(G22_n_spl_01),
    .din2(g406_p_spl_011)
  );


  LA
  g_g651_p
  (
    .dout(g651_p),
    .din1(G7_n_spl_100),
    .din2(g409_n_spl_011)
  );


  FA
  g_g651_n
  (
    .dout(g651_n),
    .din1(G7_p_spl_100),
    .din2(g409_p_spl_011)
  );


  LA
  g_g652_p
  (
    .dout(g652_p),
    .din1(g650_n),
    .din2(g651_n)
  );


  FA
  g_g652_n
  (
    .dout(g652_n),
    .din1(g650_p),
    .din2(g651_p)
  );


  LA
  g_g653_p
  (
    .dout(g653_p),
    .din1(G8_n_spl_101),
    .din2(g414_n_spl_100)
  );


  FA
  g_g653_n
  (
    .dout(g653_n),
    .din1(G8_p_spl_110),
    .din2(g414_p_spl_100)
  );


  LA
  g_g654_p
  (
    .dout(g654_p),
    .din1(G11_n_spl_11),
    .din2(g423_n_spl_011)
  );


  FA
  g_g654_n
  (
    .dout(g654_n),
    .din1(G11_p_spl_11),
    .din2(g423_p_spl_011)
  );


  LA
  g_g655_p
  (
    .dout(g655_p),
    .din1(g653_n_spl_),
    .din2(g654_n_spl_)
  );


  FA
  g_g655_n
  (
    .dout(g655_n),
    .din1(g653_p_spl_),
    .din2(g654_p_spl_)
  );


  LA
  g_g656_p
  (
    .dout(g656_p),
    .din1(G9_p_spl_110),
    .din2(G21_n_spl_01)
  );


  FA
  g_g656_n
  (
    .dout(g656_n),
    .din1(G9_n_spl_110),
    .din2(G21_p_spl_01)
  );


  LA
  g_g657_p
  (
    .dout(g657_p),
    .din1(g412_n_spl_011),
    .din2(g656_n)
  );


  FA
  g_g657_n
  (
    .dout(g657_n),
    .din1(g412_p_spl_011),
    .din2(g656_p)
  );


  LA
  g_g658_p
  (
    .dout(g658_p),
    .din1(g655_p),
    .din2(g657_n)
  );


  FA
  g_g658_n
  (
    .dout(g658_n),
    .din1(g655_n),
    .din2(g657_p)
  );


  LA
  g_g659_p
  (
    .dout(g659_p),
    .din1(g652_p),
    .din2(g658_p)
  );


  FA
  g_g659_n
  (
    .dout(g659_n),
    .din1(g652_n),
    .din2(g658_n)
  );


  LA
  g_g660_p
  (
    .dout(g660_p),
    .din1(g649_p_spl_),
    .din2(g659_p)
  );


  FA
  g_g660_n
  (
    .dout(g660_n),
    .din1(g649_n_spl_),
    .din2(g659_n)
  );


  LA
  g_g661_p
  (
    .dout(g661_p),
    .din1(g645_n),
    .din2(g660_n)
  );


  FA
  g_g661_n
  (
    .dout(g661_n),
    .din1(g645_p),
    .din2(g660_p)
  );


  LA
  g_g662_p
  (
    .dout(g662_p),
    .din1(g393_n_spl_011),
    .din2(g661_n)
  );


  FA
  g_g662_n
  (
    .dout(g662_n),
    .din1(g393_p_spl_011),
    .din2(g661_p)
  );


  LA
  g_g663_p
  (
    .dout(g663_p),
    .din1(G6_n_spl_10),
    .din2(g102_p_spl_)
  );


  FA
  g_g663_n
  (
    .dout(g663_n),
    .din1(G6_p_spl_10),
    .din2(g102_n_spl_)
  );


  LA
  g_g664_p
  (
    .dout(g664_p),
    .din1(G7_n_spl_101),
    .din2(G8_p_spl_110)
  );


  FA
  g_g664_n
  (
    .dout(g664_n),
    .din1(G7_p_spl_101),
    .din2(G8_n_spl_110)
  );


  LA
  g_g665_p
  (
    .dout(g665_p),
    .din1(g117_n_spl_),
    .din2(g664_p)
  );


  FA
  g_g665_n
  (
    .dout(g665_n),
    .din1(g117_p_spl_),
    .din2(g664_n)
  );


  LA
  g_g666_p
  (
    .dout(g666_p),
    .din1(G6_p_spl_1),
    .din2(g665_p)
  );


  FA
  g_g666_n
  (
    .dout(g666_n),
    .din1(G6_n_spl_1),
    .din2(g665_n)
  );


  LA
  g_g667_p
  (
    .dout(g667_p),
    .din1(g663_n),
    .din2(g666_n)
  );


  FA
  g_g667_n
  (
    .dout(g667_n),
    .din1(g663_p),
    .din2(g666_p)
  );


  LA
  g_g668_p
  (
    .dout(g668_p),
    .din1(g196_p_spl_),
    .din2(g667_n)
  );


  FA
  g_g668_n
  (
    .dout(g668_n),
    .din1(g196_n_spl_),
    .din2(g667_p)
  );


  LA
  g_g669_p
  (
    .dout(g669_p),
    .din1(G14_n_spl_101),
    .din2(g668_p)
  );


  FA
  g_g669_n
  (
    .dout(g669_n),
    .din1(G14_p_spl_101),
    .din2(g668_n)
  );


  LA
  g_g670_p
  (
    .dout(g670_p),
    .din1(g394_p_spl_01),
    .din2(g669_p)
  );


  FA
  g_g670_n
  (
    .dout(g670_n),
    .din1(g394_n_spl_01),
    .din2(g669_n)
  );


  LA
  g_g671_p
  (
    .dout(g671_p),
    .din1(G13_p_spl_110),
    .din2(g394_n_spl_1)
  );


  FA
  g_g671_n
  (
    .dout(g671_n),
    .din1(G13_n_spl_110),
    .din2(g394_p_spl_1)
  );


  LA
  g_g672_p
  (
    .dout(g672_p),
    .din1(g670_n),
    .din2(g671_n)
  );


  FA
  g_g672_n
  (
    .dout(g672_n),
    .din1(g670_p),
    .din2(g671_p)
  );


  LA
  g_g673_p
  (
    .dout(g673_p),
    .din1(g393_p_spl_011),
    .din2(g672_p)
  );


  FA
  g_g673_n
  (
    .dout(g673_n),
    .din1(g393_n_spl_011),
    .din2(g672_n)
  );


  LA
  g_g674_p
  (
    .dout(g674_p),
    .din1(g370_p_spl_1),
    .din2(g390_p_spl_1)
  );


  FA
  g_g674_n
  (
    .dout(g674_n),
    .din1(g370_n_spl_1),
    .din2(g390_n_spl_1)
  );


  LA
  g_g675_p
  (
    .dout(g675_p),
    .din1(g385_p_spl_01),
    .din2(g674_n)
  );


  FA
  g_g675_n
  (
    .dout(g675_n),
    .din1(g385_n_spl_01),
    .din2(g674_p)
  );


  LA
  g_g676_p
  (
    .dout(g676_p),
    .din1(g673_n),
    .din2(g675_p)
  );


  FA
  g_g676_n
  (
    .dout(g676_n),
    .din1(g673_p),
    .din2(g675_n)
  );


  LA
  g_g677_p
  (
    .dout(g677_p),
    .din1(g662_n),
    .din2(g676_p)
  );


  FA
  g_g677_n
  (
    .dout(g677_n),
    .din1(g662_p),
    .din2(g676_n)
  );


  LA
  g_g678_p
  (
    .dout(g678_p),
    .din1(g631_n),
    .din2(g677_n)
  );


  FA
  g_g678_n
  (
    .dout(g678_n),
    .din1(g631_p),
    .din2(g677_p)
  );


  LA
  g_g679_p
  (
    .dout(g679_p),
    .din1(g630_n),
    .din2(g678_p)
  );


  FA
  g_g679_n
  (
    .dout(g679_n),
    .din1(g630_p),
    .din2(g678_n)
  );


  LA
  g_g680_p
  (
    .dout(g680_p),
    .din1(g620_p_spl_0),
    .din2(g628_n_spl_0)
  );


  FA
  g_g680_n
  (
    .dout(g680_n),
    .din1(g620_n_spl_0),
    .din2(g628_p_spl_0)
  );


  LA
  g_g681_p
  (
    .dout(g681_p),
    .din1(g620_n_spl_1),
    .din2(g628_p_spl_)
  );


  FA
  g_g681_n
  (
    .dout(g681_n),
    .din1(g620_p_spl_1),
    .din2(g628_n_spl_)
  );


  LA
  g_g682_p
  (
    .dout(g682_p),
    .din1(g680_n),
    .din2(g681_n)
  );


  FA
  g_g682_n
  (
    .dout(g682_n),
    .din1(g680_p),
    .din2(g681_p)
  );


  LA
  g_g683_p
  (
    .dout(g683_p),
    .din1(g377_n_spl_10),
    .din2(g682_n)
  );


  FA
  g_g683_n
  (
    .dout(g683_n),
    .din1(g377_p_spl_01),
    .din2(g682_p)
  );


  LA
  g_g684_p
  (
    .dout(g684_p),
    .din1(g384_n_spl_01),
    .din2(g620_n_spl_1)
  );


  FA
  g_g684_n
  (
    .dout(g684_n),
    .din1(g384_p_spl_01),
    .din2(g620_p_spl_1)
  );


  LA
  g_g685_p
  (
    .dout(g685_p),
    .din1(G4_p_spl_1101),
    .din2(g432_n_spl_)
  );


  FA
  g_g685_n
  (
    .dout(g685_n),
    .din1(G4_n_spl_1101),
    .din2(g432_p_spl_)
  );


  LA
  g_g686_p
  (
    .dout(g686_p),
    .din1(G43_p_spl_1),
    .din2(g406_n_spl_100)
  );


  FA
  g_g686_n
  (
    .dout(g686_n),
    .din1(G43_n_spl_1),
    .din2(g406_p_spl_100)
  );


  LA
  g_g687_p
  (
    .dout(g687_p),
    .din1(g685_p_spl_),
    .din2(g686_n)
  );


  FA
  g_g687_n
  (
    .dout(g687_n),
    .din1(g685_n_spl_),
    .din2(g686_p)
  );


  LA
  g_g688_p
  (
    .dout(g688_p),
    .din1(G14_n_spl_110),
    .din2(g423_n_spl_011)
  );


  FA
  g_g688_n
  (
    .dout(g688_n),
    .din1(G14_p_spl_110),
    .din2(g423_p_spl_011)
  );


  LA
  g_g689_p
  (
    .dout(g689_p),
    .din1(G41_p_spl_10),
    .din2(g414_n_spl_101)
  );


  FA
  g_g689_n
  (
    .dout(g689_n),
    .din1(G41_n_spl_10),
    .din2(g414_p_spl_101)
  );


  LA
  g_g690_p
  (
    .dout(g690_p),
    .din1(G42_p_spl_1),
    .din2(g409_n_spl_100)
  );


  FA
  g_g690_n
  (
    .dout(g690_n),
    .din1(G42_n_spl_1),
    .din2(g409_p_spl_100)
  );


  LA
  g_g691_p
  (
    .dout(g691_p),
    .din1(g689_n),
    .din2(g690_n)
  );


  FA
  g_g691_n
  (
    .dout(g691_n),
    .din1(g689_p),
    .din2(g690_p)
  );


  LA
  g_g692_p
  (
    .dout(g692_p),
    .din1(g688_n),
    .din2(g691_p)
  );


  FA
  g_g692_n
  (
    .dout(g692_n),
    .din1(g688_p),
    .din2(g691_n)
  );


  LA
  g_g693_p
  (
    .dout(g693_p),
    .din1(g687_p),
    .din2(g692_p)
  );


  FA
  g_g693_n
  (
    .dout(g693_n),
    .din1(g687_n),
    .din2(g692_n)
  );


  LA
  g_g694_p
  (
    .dout(g694_p),
    .din1(G39_p_spl_10),
    .din2(g425_n_spl_100)
  );


  FA
  g_g694_n
  (
    .dout(g694_n),
    .din1(G39_n_spl_10),
    .din2(g425_p_spl_100)
  );


  LA
  g_g695_p
  (
    .dout(g695_p),
    .din1(G40_n_spl_10),
    .din2(G44_n_spl_)
  );


  FA
  g_g695_n
  (
    .dout(g695_n),
    .din1(G40_p_spl_10),
    .din2(G44_p_spl_)
  );


  LA
  g_g696_p
  (
    .dout(g696_p),
    .din1(g412_n_spl_100),
    .din2(g695_n)
  );


  FA
  g_g696_n
  (
    .dout(g696_n),
    .din1(g412_p_spl_100),
    .din2(g695_p)
  );


  LA
  g_g697_p
  (
    .dout(g697_p),
    .din1(g694_n),
    .din2(g696_n)
  );


  FA
  g_g697_n
  (
    .dout(g697_n),
    .din1(g694_p),
    .din2(g696_p)
  );


  LA
  g_g698_p
  (
    .dout(g698_p),
    .din1(g693_p),
    .din2(g697_p)
  );


  FA
  g_g698_n
  (
    .dout(g698_n),
    .din1(g693_n),
    .din2(g697_n)
  );


  LA
  g_g699_p
  (
    .dout(g699_p),
    .din1(G21_p_spl_10),
    .din2(g406_n_spl_100)
  );


  FA
  g_g699_n
  (
    .dout(g699_n),
    .din1(G21_n_spl_10),
    .din2(g406_p_spl_100)
  );


  LA
  g_g700_p
  (
    .dout(g700_p),
    .din1(G22_p_spl_10),
    .din2(g409_n_spl_100)
  );


  FA
  g_g700_n
  (
    .dout(g700_n),
    .din1(G22_n_spl_10),
    .din2(g409_p_spl_100)
  );


  LA
  g_g701_p
  (
    .dout(g701_p),
    .din1(g699_n),
    .din2(g700_n)
  );


  FA
  g_g701_n
  (
    .dout(g701_n),
    .din1(g699_p),
    .din2(g700_p)
  );


  LA
  g_g702_p
  (
    .dout(g702_p),
    .din1(G9_n_spl_110),
    .din2(g425_n_spl_100)
  );


  FA
  g_g702_n
  (
    .dout(g702_n),
    .din1(G9_p_spl_110),
    .din2(g425_p_spl_100)
  );


  LA
  g_g703_p
  (
    .dout(g703_p),
    .din1(G4_n_spl_1110),
    .din2(g702_n)
  );


  FA
  g_g703_n
  (
    .dout(g703_n),
    .din1(G4_p_spl_1110),
    .din2(g702_p)
  );


  LA
  g_g704_p
  (
    .dout(g704_p),
    .din1(g701_p),
    .din2(g703_p)
  );


  FA
  g_g704_n
  (
    .dout(g704_n),
    .din1(g701_n),
    .din2(g703_n)
  );


  LA
  g_g705_p
  (
    .dout(g705_p),
    .din1(G10_n_spl_110),
    .din2(g423_n_spl_10)
  );


  FA
  g_g705_n
  (
    .dout(g705_n),
    .din1(G10_p_spl_11),
    .din2(g423_p_spl_10)
  );


  LA
  g_g706_p
  (
    .dout(g706_p),
    .din1(G8_p_spl_111),
    .din2(G20_n_spl_0)
  );


  FA
  g_g706_n
  (
    .dout(g706_n),
    .din1(G8_n_spl_110),
    .din2(G20_p_spl_0)
  );


  LA
  g_g707_p
  (
    .dout(g707_p),
    .din1(g412_n_spl_100),
    .din2(g706_n_spl_)
  );


  FA
  g_g707_n
  (
    .dout(g707_n),
    .din1(g412_p_spl_100),
    .din2(g706_p_spl_)
  );


  LA
  g_g708_p
  (
    .dout(g708_p),
    .din1(g705_n_spl_),
    .din2(g707_n)
  );


  FA
  g_g708_n
  (
    .dout(g708_n),
    .din1(g705_p_spl_),
    .din2(g707_p)
  );


  LA
  g_g709_p
  (
    .dout(g709_p),
    .din1(G7_n_spl_101),
    .din2(g414_n_spl_101)
  );


  FA
  g_g709_n
  (
    .dout(g709_n),
    .din1(G7_p_spl_101),
    .din2(g414_p_spl_101)
  );


  LA
  g_g710_p
  (
    .dout(g710_p),
    .din1(g480_n_spl_),
    .din2(g709_n)
  );


  FA
  g_g710_n
  (
    .dout(g710_n),
    .din1(g480_p_spl_),
    .din2(g709_p)
  );


  LA
  g_g711_p
  (
    .dout(g711_p),
    .din1(g708_p),
    .din2(g710_p)
  );


  FA
  g_g711_n
  (
    .dout(g711_n),
    .din1(g708_n),
    .din2(g710_n)
  );


  LA
  g_g712_p
  (
    .dout(g712_p),
    .din1(g704_p),
    .din2(g711_p)
  );


  FA
  g_g712_n
  (
    .dout(g712_n),
    .din1(g704_n),
    .din2(g711_n)
  );


  LA
  g_g713_p
  (
    .dout(g713_p),
    .din1(g698_n),
    .din2(g712_n)
  );


  FA
  g_g713_n
  (
    .dout(g713_n),
    .din1(g698_p),
    .din2(g712_p)
  );


  LA
  g_g714_p
  (
    .dout(g714_p),
    .din1(g393_n_spl_100),
    .din2(g713_n)
  );


  FA
  g_g714_n
  (
    .dout(g714_n),
    .din1(g393_p_spl_100),
    .din2(g713_p)
  );


  LA
  g_g715_p
  (
    .dout(g715_p),
    .din1(g390_p_spl_1),
    .din2(g597_p_spl_1)
  );


  FA
  g_g715_n
  (
    .dout(g715_n),
    .din1(g390_n_spl_1),
    .din2(g597_n_spl_1)
  );


  LA
  g_g716_p
  (
    .dout(g716_p),
    .din1(G12_p_spl_110),
    .din2(g394_n_spl_1)
  );


  FA
  g_g716_n
  (
    .dout(g716_n),
    .din1(G12_n_spl_11),
    .din2(g394_p_spl_1)
  );


  LA
  g_g717_p
  (
    .dout(g717_p),
    .din1(g393_p_spl_100),
    .din2(g716_n)
  );


  FA
  g_g717_n
  (
    .dout(g717_n),
    .din1(g393_n_spl_100),
    .din2(g716_p)
  );


  LA
  g_g718_p
  (
    .dout(g718_p),
    .din1(g385_p_spl_10),
    .din2(g717_n)
  );


  FA
  g_g718_n
  (
    .dout(g718_n),
    .din1(g385_n_spl_10),
    .din2(g717_p)
  );


  LA
  g_g719_p
  (
    .dout(g719_p),
    .din1(g715_n),
    .din2(g718_p)
  );


  FA
  g_g719_n
  (
    .dout(g719_n),
    .din1(g715_p),
    .din2(g718_n)
  );


  LA
  g_g720_p
  (
    .dout(g720_p),
    .din1(g714_n),
    .din2(g719_p)
  );


  FA
  g_g720_n
  (
    .dout(g720_n),
    .din1(g714_p),
    .din2(g719_n)
  );


  LA
  g_g721_p
  (
    .dout(g721_p),
    .din1(g684_n),
    .din2(g720_n)
  );


  FA
  g_g721_n
  (
    .dout(g721_n),
    .din1(g684_p),
    .din2(g720_p)
  );


  LA
  g_g722_p
  (
    .dout(g722_p),
    .din1(g683_n),
    .din2(g721_p)
  );


  FA
  g_g722_n
  (
    .dout(g722_n),
    .din1(g683_p),
    .din2(g721_n)
  );


  LA
  g_g723_p
  (
    .dout(g723_p),
    .din1(G47_p_spl_10),
    .din2(g519_p_spl_)
  );


  FA
  g_g723_n
  (
    .dout(g723_n),
    .din1(G47_n_spl_10),
    .din2(g519_n_spl_)
  );


  LA
  g_g724_p
  (
    .dout(g724_p),
    .din1(g513_p_spl_00),
    .din2(g723_p_spl_)
  );


  FA
  g_g724_n
  (
    .dout(g724_n),
    .din1(g513_n_spl_00),
    .din2(g723_n_spl_)
  );


  LA
  g_g725_p
  (
    .dout(g725_p),
    .din1(g513_p_spl_0),
    .din2(g530_n_spl_0)
  );


  FA
  g_g725_n
  (
    .dout(g725_n),
    .din1(g513_n_spl_0),
    .din2(g530_p_spl_0)
  );


  LA
  g_g726_p
  (
    .dout(g726_p),
    .din1(g528_n_spl_),
    .din2(g725_n)
  );


  FA
  g_g726_n
  (
    .dout(g726_n),
    .din1(g528_p_spl_),
    .din2(g725_p)
  );


  LA
  g_g727_p
  (
    .dout(g727_p),
    .din1(g517_p_spl_0),
    .din2(g726_p_spl_)
  );


  FA
  g_g727_n
  (
    .dout(g727_n),
    .din1(g517_n_spl_0),
    .din2(g726_n_spl_)
  );


  LA
  g_g728_p
  (
    .dout(g728_p),
    .din1(g517_n_spl_1),
    .din2(g726_n_spl_)
  );


  FA
  g_g728_n
  (
    .dout(g728_n),
    .din1(g517_p_spl_1),
    .din2(g726_p_spl_)
  );


  LA
  g_g729_p
  (
    .dout(g729_p),
    .din1(g727_n),
    .din2(g728_n)
  );


  FA
  g_g729_n
  (
    .dout(g729_n),
    .din1(g727_p),
    .din2(g728_p)
  );


  LA
  g_g730_p
  (
    .dout(g730_p),
    .din1(g724_p_spl_0),
    .din2(g729_p_spl_)
  );


  FA
  g_g730_n
  (
    .dout(g730_n),
    .din1(g724_n_spl_0),
    .din2(g729_n_spl_)
  );


  LA
  g_g731_p
  (
    .dout(g731_p),
    .din1(g724_n_spl_0),
    .din2(g729_n_spl_)
  );


  FA
  g_g731_n
  (
    .dout(g731_n),
    .din1(g724_p_spl_0),
    .din2(g729_p_spl_)
  );


  LA
  g_g732_p
  (
    .dout(g732_p),
    .din1(g730_n_spl_0),
    .din2(g731_n)
  );


  FA
  g_g732_n
  (
    .dout(g732_n),
    .din1(g730_p_spl_0),
    .din2(g731_p)
  );


  LA
  g_g733_p
  (
    .dout(g733_p),
    .din1(g503_n_spl_),
    .din2(g530_n_spl_)
  );


  FA
  g_g733_n
  (
    .dout(g733_n),
    .din1(g503_p_spl_),
    .din2(g530_p_spl_)
  );


  LA
  g_g734_p
  (
    .dout(g734_p),
    .din1(g513_n_spl_1),
    .din2(g723_n_spl_)
  );


  FA
  g_g734_n
  (
    .dout(g734_n),
    .din1(g513_p_spl_1),
    .din2(g723_p_spl_)
  );


  LA
  g_g735_p
  (
    .dout(g735_p),
    .din1(g724_n_spl_),
    .din2(g734_n)
  );


  FA
  g_g735_n
  (
    .dout(g735_n),
    .din1(g724_p_spl_),
    .din2(g734_p)
  );


  LA
  g_g736_p
  (
    .dout(g736_p),
    .din1(g733_p_spl_),
    .din2(g735_n_spl_)
  );


  FA
  g_g736_n
  (
    .dout(g736_n),
    .din1(g733_n_spl_),
    .din2(g735_p_spl_)
  );


  LA
  g_g737_p
  (
    .dout(g737_p),
    .din1(g733_n_spl_),
    .din2(g735_p_spl_)
  );


  FA
  g_g737_n
  (
    .dout(g737_n),
    .din1(g733_p_spl_),
    .din2(g735_n_spl_)
  );


  LA
  g_g738_p
  (
    .dout(g738_p),
    .din1(g736_n),
    .din2(g737_n)
  );


  FA
  g_g738_n
  (
    .dout(g738_n),
    .din1(g736_p),
    .din2(g737_p)
  );


  LA
  g_g739_p
  (
    .dout(g739_p),
    .din1(G47_p_spl_1),
    .din2(g527_n_spl_)
  );


  FA
  g_g739_n
  (
    .dout(g739_n),
    .din1(G47_n_spl_1),
    .din2(g527_p_spl_)
  );


  LA
  g_g740_p
  (
    .dout(g740_p),
    .din1(g521_p_spl_),
    .din2(g739_p)
  );


  FA
  g_g740_n
  (
    .dout(g740_n),
    .din1(g521_n_spl_),
    .din2(g739_n)
  );


  LA
  g_g741_p
  (
    .dout(g741_p),
    .din1(g738_n_spl_0),
    .din2(g740_n_spl_0)
  );


  FA
  g_g741_n
  (
    .dout(g741_n),
    .din1(g738_p_spl_0),
    .din2(g740_p_spl_0)
  );


  LA
  g_g742_p
  (
    .dout(g742_p),
    .din1(g732_p_spl_0),
    .din2(g741_n_spl_0)
  );


  FA
  g_g742_n
  (
    .dout(g742_n),
    .din1(g732_n_spl_0),
    .din2(g741_p_spl_0)
  );


  LA
  g_g743_p
  (
    .dout(g743_p),
    .din1(g732_n_spl_0),
    .din2(g741_p_spl_0)
  );


  FA
  g_g743_n
  (
    .dout(g743_n),
    .din1(g732_p_spl_0),
    .din2(g741_n_spl_0)
  );


  LA
  g_g744_p
  (
    .dout(g744_p),
    .din1(g742_n),
    .din2(g743_n)
  );


  FA
  g_g744_n
  (
    .dout(g744_n),
    .din1(g742_p),
    .din2(g743_p)
  );


  LA
  g_g745_p
  (
    .dout(g745_p),
    .din1(g377_n_spl_10),
    .din2(g744_n)
  );


  FA
  g_g745_n
  (
    .dout(g745_n),
    .din1(g377_p_spl_10),
    .din2(g744_p)
  );


  LA
  g_g746_p
  (
    .dout(g746_p),
    .din1(g452_p_spl_0),
    .din2(g517_p_spl_1)
  );


  FA
  g_g746_n
  (
    .dout(g746_n),
    .din1(g452_n_spl_0),
    .din2(g517_n_spl_1)
  );


  LA
  g_g747_p
  (
    .dout(g747_p),
    .din1(G8_n_spl_11),
    .din2(g393_p_spl_101)
  );


  FA
  g_g747_n
  (
    .dout(g747_n),
    .din1(G8_p_spl_111),
    .din2(g393_n_spl_101)
  );


  LA
  g_g748_p
  (
    .dout(g748_p),
    .din1(g385_p_spl_10),
    .din2(g747_n)
  );


  FA
  g_g748_n
  (
    .dout(g748_n),
    .din1(g385_n_spl_10),
    .din2(g747_p)
  );


  LA
  g_g749_p
  (
    .dout(g749_p),
    .din1(g430_n_spl_),
    .din2(g438_n_spl_)
  );


  FA
  g_g749_n
  (
    .dout(g749_n),
    .din1(g430_p_spl_),
    .din2(g438_p_spl_)
  );


  LA
  g_g750_p
  (
    .dout(g750_p),
    .din1(G39_p_spl_10),
    .din2(g406_n_spl_101)
  );


  FA
  g_g750_n
  (
    .dout(g750_n),
    .din1(G39_n_spl_10),
    .din2(g406_p_spl_101)
  );


  LA
  g_g751_p
  (
    .dout(g751_p),
    .din1(G14_n_spl_110),
    .din2(g409_n_spl_101)
  );


  FA
  g_g751_n
  (
    .dout(g751_n),
    .din1(G14_p_spl_110),
    .din2(g409_p_spl_101)
  );


  LA
  g_g752_p
  (
    .dout(g752_p),
    .din1(g750_n),
    .din2(g751_n)
  );


  FA
  g_g752_n
  (
    .dout(g752_n),
    .din1(g750_p),
    .din2(g751_p)
  );


  LA
  g_g753_p
  (
    .dout(g753_p),
    .din1(g705_n_spl_),
    .din2(g752_p)
  );


  FA
  g_g753_n
  (
    .dout(g753_n),
    .din1(g705_p_spl_),
    .din2(g752_n)
  );


  LA
  g_g754_p
  (
    .dout(g754_p),
    .din1(g412_n_spl_101),
    .din2(g569_n_spl_)
  );


  FA
  g_g754_n
  (
    .dout(g754_n),
    .din1(g412_p_spl_101),
    .din2(g569_p_spl_)
  );


  LA
  g_g755_p
  (
    .dout(g755_p),
    .din1(g685_p_spl_),
    .din2(g754_n)
  );


  FA
  g_g755_n
  (
    .dout(g755_n),
    .din1(g685_n_spl_),
    .din2(g754_p)
  );


  LA
  g_g756_p
  (
    .dout(g756_p),
    .din1(g753_p),
    .din2(g755_p)
  );


  FA
  g_g756_n
  (
    .dout(g756_n),
    .din1(g753_n),
    .din2(g755_n)
  );


  LA
  g_g757_p
  (
    .dout(g757_p),
    .din1(g749_p),
    .din2(g756_p)
  );


  FA
  g_g757_n
  (
    .dout(g757_n),
    .din1(g749_n),
    .din2(g756_n)
  );


  LA
  g_g758_p
  (
    .dout(g758_p),
    .din1(G21_p_spl_10),
    .din2(g425_n_spl_101)
  );


  FA
  g_g758_n
  (
    .dout(g758_n),
    .din1(G21_n_spl_10),
    .din2(g425_p_spl_101)
  );


  LA
  g_g759_p
  (
    .dout(g759_p),
    .din1(G17_p_spl_0),
    .din2(g406_n_spl_101)
  );


  FA
  g_g759_n
  (
    .dout(g759_n),
    .din1(G17_n_spl_0),
    .din2(g406_p_spl_101)
  );


  LA
  g_g760_p
  (
    .dout(g760_p),
    .din1(g758_n),
    .din2(g759_n)
  );


  FA
  g_g760_n
  (
    .dout(g760_n),
    .din1(g758_p),
    .din2(g759_p)
  );


  LA
  g_g761_p
  (
    .dout(g761_p),
    .din1(G22_p_spl_10),
    .din2(g423_n_spl_10)
  );


  FA
  g_g761_n
  (
    .dout(g761_n),
    .din1(G22_n_spl_10),
    .din2(g423_p_spl_10)
  );


  LA
  g_g762_p
  (
    .dout(g762_p),
    .din1(G4_n_spl_1110),
    .din2(g761_n)
  );


  FA
  g_g762_n
  (
    .dout(g762_n),
    .din1(G4_p_spl_1110),
    .din2(g761_p)
  );


  LA
  g_g763_p
  (
    .dout(g763_p),
    .din1(G18_p_spl_0),
    .din2(g409_n_spl_101)
  );


  FA
  g_g763_n
  (
    .dout(g763_n),
    .din1(G18_n_spl_0),
    .din2(g409_p_spl_101)
  );


  LA
  g_g764_p
  (
    .dout(g764_p),
    .din1(G16_n_spl_),
    .din2(G20_n_spl_1)
  );


  FA
  g_g764_n
  (
    .dout(g764_n),
    .din1(G16_p_spl_),
    .din2(G20_p_spl_1)
  );


  LA
  g_g765_p
  (
    .dout(g765_p),
    .din1(g412_n_spl_101),
    .din2(g764_n)
  );


  FA
  g_g765_n
  (
    .dout(g765_n),
    .din1(g412_p_spl_101),
    .din2(g764_p)
  );


  LA
  g_g766_p
  (
    .dout(g766_p),
    .din1(G7_p_spl_110),
    .din2(G19_n_spl_0)
  );


  FA
  g_g766_n
  (
    .dout(g766_n),
    .din1(G7_n_spl_110),
    .din2(G19_p_spl_0)
  );


  LA
  g_g767_p
  (
    .dout(g767_p),
    .din1(g414_n_spl_110),
    .din2(g766_n)
  );


  FA
  g_g767_n
  (
    .dout(g767_n),
    .din1(g414_p_spl_110),
    .din2(g766_p)
  );


  LA
  g_g768_p
  (
    .dout(g768_p),
    .din1(g765_n),
    .din2(g767_n)
  );


  FA
  g_g768_n
  (
    .dout(g768_n),
    .din1(g765_p),
    .din2(g767_p)
  );


  LA
  g_g769_p
  (
    .dout(g769_p),
    .din1(g763_n),
    .din2(g768_p)
  );


  FA
  g_g769_n
  (
    .dout(g769_n),
    .din1(g763_p),
    .din2(g768_n)
  );


  LA
  g_g770_p
  (
    .dout(g770_p),
    .din1(g762_p),
    .din2(g769_p)
  );


  FA
  g_g770_n
  (
    .dout(g770_n),
    .din1(g762_n),
    .din2(g769_n)
  );


  LA
  g_g771_p
  (
    .dout(g771_p),
    .din1(g760_p),
    .din2(g770_p)
  );


  FA
  g_g771_n
  (
    .dout(g771_n),
    .din1(g760_n),
    .din2(g770_n)
  );


  LA
  g_g772_p
  (
    .dout(g772_p),
    .din1(g757_n),
    .din2(g771_n)
  );


  FA
  g_g772_n
  (
    .dout(g772_n),
    .din1(g757_p),
    .din2(g771_p)
  );


  LA
  g_g773_p
  (
    .dout(g773_p),
    .din1(g393_n_spl_101),
    .din2(g772_n)
  );


  FA
  g_g773_n
  (
    .dout(g773_n),
    .din1(g393_p_spl_101),
    .din2(g772_p)
  );


  LA
  g_g774_p
  (
    .dout(g774_p),
    .din1(g748_p),
    .din2(g773_n)
  );


  FA
  g_g774_n
  (
    .dout(g774_n),
    .din1(g748_n),
    .din2(g773_p)
  );


  LA
  g_g775_p
  (
    .dout(g775_p),
    .din1(g746_n),
    .din2(g774_p)
  );


  FA
  g_g775_n
  (
    .dout(g775_n),
    .din1(g746_p),
    .din2(g774_n)
  );


  LA
  g_g776_p
  (
    .dout(g776_p),
    .din1(g384_n_spl_10),
    .din2(g732_n_spl_1)
  );


  FA
  g_g776_n
  (
    .dout(g776_n),
    .din1(g384_p_spl_10),
    .din2(g732_p_spl_1)
  );


  LA
  g_g777_p
  (
    .dout(g777_p),
    .din1(g775_n),
    .din2(g776_n)
  );


  FA
  g_g777_n
  (
    .dout(g777_n),
    .din1(g775_p),
    .din2(g776_p)
  );


  LA
  g_g778_p
  (
    .dout(g778_p),
    .din1(g745_n),
    .din2(g777_p)
  );


  FA
  g_g778_n
  (
    .dout(g778_n),
    .din1(g745_p),
    .din2(g777_n)
  );


  LA
  g_g779_p
  (
    .dout(g779_p),
    .din1(g306_n_spl_),
    .din2(g365_p_spl_1)
  );


  FA
  g_g779_n
  (
    .dout(g779_n),
    .din1(g306_p_spl_),
    .din2(g365_n_spl_1)
  );


  LA
  g_g780_p
  (
    .dout(g780_p),
    .din1(g320_n_spl_1),
    .din2(g779_n_spl_)
  );


  FA
  g_g780_n
  (
    .dout(g780_n),
    .din1(g320_p_spl_1),
    .din2(g779_p_spl_)
  );


  LA
  g_g781_p
  (
    .dout(g781_p),
    .din1(g320_p_spl_1),
    .din2(g779_p_spl_)
  );


  FA
  g_g781_n
  (
    .dout(g781_n),
    .din1(g320_n_spl_1),
    .din2(g779_n_spl_)
  );


  LA
  g_g782_p
  (
    .dout(g782_p),
    .din1(g780_n),
    .din2(g781_n)
  );


  FA
  g_g782_n
  (
    .dout(g782_n),
    .din1(g780_p),
    .din2(g781_p)
  );


  LA
  g_g783_p
  (
    .dout(g783_p),
    .din1(g452_p_spl_1),
    .din2(g782_p_spl_0)
  );


  FA
  g_g783_n
  (
    .dout(g783_n),
    .din1(g452_n_spl_1),
    .din2(g782_n_spl_0)
  );


  LA
  g_g784_p
  (
    .dout(g784_p),
    .din1(G11_p_spl_11),
    .din2(G39_n_spl_11)
  );


  FA
  g_g784_n
  (
    .dout(g784_n),
    .din1(G11_n_spl_11),
    .din2(G39_p_spl_11)
  );


  LA
  g_g785_p
  (
    .dout(g785_p),
    .din1(g412_n_spl_110),
    .din2(g784_n)
  );


  FA
  g_g785_n
  (
    .dout(g785_n),
    .din1(g412_p_spl_110),
    .din2(g784_p)
  );


  LA
  g_g786_p
  (
    .dout(g786_p),
    .din1(G5_p_spl_1),
    .din2(g579_n_spl_)
  );


  FA
  g_g786_n
  (
    .dout(g786_n),
    .din1(G5_n_spl_1),
    .din2(g579_p_spl_)
  );


  LA
  g_g787_p
  (
    .dout(g787_p),
    .din1(g649_p_spl_),
    .din2(g786_p)
  );


  FA
  g_g787_n
  (
    .dout(g787_n),
    .din1(g649_n_spl_),
    .din2(g786_n)
  );


  LA
  g_g788_p
  (
    .dout(g788_p),
    .din1(G14_n_spl_111),
    .din2(g406_n_spl_110)
  );


  FA
  g_g788_n
  (
    .dout(g788_n),
    .din1(G14_p_spl_111),
    .din2(g406_p_spl_110)
  );


  LA
  g_g789_p
  (
    .dout(g789_p),
    .din1(G13_n_spl_110),
    .din2(g409_n_spl_110)
  );


  FA
  g_g789_n
  (
    .dout(g789_n),
    .din1(G13_p_spl_111),
    .din2(g409_p_spl_110)
  );


  LA
  g_g790_p
  (
    .dout(g790_p),
    .din1(g788_n),
    .din2(g789_n)
  );


  FA
  g_g790_n
  (
    .dout(g790_n),
    .din1(g788_p),
    .din2(g789_p)
  );


  LA
  g_g791_p
  (
    .dout(g791_p),
    .din1(g653_n_spl_),
    .din2(g790_p)
  );


  FA
  g_g791_n
  (
    .dout(g791_n),
    .din1(g653_p_spl_),
    .din2(g790_n)
  );


  LA
  g_g792_p
  (
    .dout(g792_p),
    .din1(g787_p),
    .din2(g791_p)
  );


  FA
  g_g792_n
  (
    .dout(g792_n),
    .din1(g787_n),
    .din2(g791_n)
  );


  LA
  g_g793_p
  (
    .dout(g793_p),
    .din1(g785_n),
    .din2(g792_p)
  );


  FA
  g_g793_n
  (
    .dout(g793_n),
    .din1(g785_p),
    .din2(g792_n)
  );


  LA
  g_g794_p
  (
    .dout(g794_p),
    .din1(G5_n_spl_1),
    .din2(G7_n_spl_110)
  );


  FA
  g_g794_n
  (
    .dout(g794_n),
    .din1(G5_p_spl_1),
    .din2(G7_p_spl_110)
  );


  LA
  g_g795_p
  (
    .dout(g795_p),
    .din1(G17_p_spl_0),
    .din2(g409_n_spl_110)
  );


  FA
  g_g795_n
  (
    .dout(g795_n),
    .din1(G17_n_spl_0),
    .din2(g409_p_spl_110)
  );


  LA
  g_g796_p
  (
    .dout(g796_p),
    .din1(G15_n),
    .din2(G19_n_spl_1)
  );


  FA
  g_g796_n
  (
    .dout(g796_n),
    .din1(G15_p),
    .din2(G19_p_spl_1)
  );


  LA
  g_g797_p
  (
    .dout(g797_p),
    .din1(g412_n_spl_110),
    .din2(g796_n)
  );


  FA
  g_g797_n
  (
    .dout(g797_n),
    .din1(g412_p_spl_110),
    .din2(g796_p)
  );


  LA
  g_g798_p
  (
    .dout(g798_p),
    .din1(G18_n_spl_1),
    .din2(G22_n_spl_11)
  );


  FA
  g_g798_n
  (
    .dout(g798_n),
    .din1(G18_p_spl_1),
    .din2(G22_p_spl_11)
  );


  LA
  g_g799_p
  (
    .dout(g799_p),
    .din1(g414_n_spl_110),
    .din2(g798_n)
  );


  FA
  g_g799_n
  (
    .dout(g799_n),
    .din1(g414_p_spl_110),
    .din2(g798_p)
  );


  LA
  g_g800_p
  (
    .dout(g800_p),
    .din1(g797_n),
    .din2(g799_n)
  );


  FA
  g_g800_n
  (
    .dout(g800_n),
    .din1(g797_p),
    .din2(g799_p)
  );


  LA
  g_g801_p
  (
    .dout(g801_p),
    .din1(g795_n),
    .din2(g800_p)
  );


  FA
  g_g801_n
  (
    .dout(g801_n),
    .din1(g795_p),
    .din2(g800_n)
  );


  LA
  g_g802_p
  (
    .dout(g802_p),
    .din1(G21_p_spl_11),
    .din2(g423_n_spl_11)
  );


  FA
  g_g802_n
  (
    .dout(g802_n),
    .din1(G21_n_spl_11),
    .din2(g423_p_spl_11)
  );


  LA
  g_g803_p
  (
    .dout(g803_p),
    .din1(g146_p_spl_),
    .din2(g802_n)
  );


  FA
  g_g803_n
  (
    .dout(g803_n),
    .din1(g146_n_spl_),
    .din2(g802_p)
  );


  LA
  g_g804_p
  (
    .dout(g804_p),
    .din1(G20_p_spl_1),
    .din2(g425_n_spl_101)
  );


  FA
  g_g804_n
  (
    .dout(g804_n),
    .din1(G20_n_spl_1),
    .din2(g425_p_spl_101)
  );


  LA
  g_g805_p
  (
    .dout(g805_p),
    .din1(G16_p_spl_),
    .din2(g406_n_spl_110)
  );


  FA
  g_g805_n
  (
    .dout(g805_n),
    .din1(G16_n_spl_),
    .din2(g406_p_spl_110)
  );


  LA
  g_g806_p
  (
    .dout(g806_p),
    .din1(g804_n),
    .din2(g805_n)
  );


  FA
  g_g806_n
  (
    .dout(g806_n),
    .din1(g804_p),
    .din2(g805_p)
  );


  LA
  g_g807_p
  (
    .dout(g807_p),
    .din1(g803_p),
    .din2(g806_p)
  );


  FA
  g_g807_n
  (
    .dout(g807_n),
    .din1(g803_n),
    .din2(g806_n)
  );


  LA
  g_g808_p
  (
    .dout(g808_p),
    .din1(g801_p),
    .din2(g807_p)
  );


  FA
  g_g808_n
  (
    .dout(g808_n),
    .din1(g801_n),
    .din2(g807_n)
  );


  LA
  g_g809_p
  (
    .dout(g809_p),
    .din1(g794_n),
    .din2(g808_n)
  );


  FA
  g_g809_n
  (
    .dout(g809_n),
    .din1(g794_p),
    .din2(g808_p)
  );


  LA
  g_g810_p
  (
    .dout(g810_p),
    .din1(g793_n),
    .din2(g809_p)
  );


  FA
  g_g810_n
  (
    .dout(g810_n),
    .din1(g793_p),
    .din2(g809_n)
  );


  LA
  g_g811_p
  (
    .dout(g811_p),
    .din1(g393_n_spl_110),
    .din2(g810_n)
  );


  FA
  g_g811_n
  (
    .dout(g811_n),
    .din1(g393_p_spl_110),
    .din2(g810_p)
  );


  LA
  g_g812_p
  (
    .dout(g812_p),
    .din1(G7_n_spl_111),
    .din2(g393_p_spl_110)
  );


  FA
  g_g812_n
  (
    .dout(g812_n),
    .din1(G7_p_spl_111),
    .din2(g393_n_spl_110)
  );


  LA
  g_g813_p
  (
    .dout(g813_p),
    .din1(g385_p_spl_11),
    .din2(g812_n)
  );


  FA
  g_g813_n
  (
    .dout(g813_n),
    .din1(g385_n_spl_11),
    .din2(g812_p)
  );


  LA
  g_g814_p
  (
    .dout(g814_p),
    .din1(g811_n),
    .din2(g813_p)
  );


  FA
  g_g814_n
  (
    .dout(g814_n),
    .din1(g811_p),
    .din2(g813_n)
  );


  LA
  g_g815_p
  (
    .dout(g815_p),
    .din1(g783_n),
    .din2(g814_p)
  );


  FA
  g_g815_n
  (
    .dout(g815_n),
    .din1(g783_p),
    .din2(g814_n)
  );


  LA
  g_g816_p
  (
    .dout(g816_p),
    .din1(g534_p_spl_1),
    .din2(g782_n_spl_0)
  );


  FA
  g_g816_n
  (
    .dout(g816_n),
    .din1(g534_n_spl_1),
    .din2(g782_p_spl_0)
  );


  LA
  g_g817_p
  (
    .dout(g817_p),
    .din1(g534_n_spl_1),
    .din2(g782_p_spl_)
  );


  FA
  g_g817_n
  (
    .dout(g817_n),
    .din1(g534_p_spl_1),
    .din2(g782_n_spl_)
  );


  LA
  g_g818_p
  (
    .dout(g818_p),
    .din1(g816_n),
    .din2(g817_n)
  );


  FA
  g_g818_n
  (
    .dout(g818_n),
    .din1(g816_p),
    .din2(g817_p)
  );


  LA
  g_g819_p
  (
    .dout(g819_p),
    .din1(g730_n_spl_0),
    .din2(g818_p_spl_)
  );


  FA
  g_g819_n
  (
    .dout(g819_n),
    .din1(g730_p_spl_0),
    .din2(g818_n_spl_)
  );


  LA
  g_g820_p
  (
    .dout(g820_p),
    .din1(g730_p_spl_),
    .din2(g818_n_spl_)
  );


  FA
  g_g820_n
  (
    .dout(g820_n),
    .din1(g730_n_spl_),
    .din2(g818_p_spl_)
  );


  LA
  g_g821_p
  (
    .dout(g821_p),
    .din1(g819_n),
    .din2(g820_n)
  );


  FA
  g_g821_n
  (
    .dout(g821_n),
    .din1(g819_p),
    .din2(g820_p)
  );


  LA
  g_g822_p
  (
    .dout(g822_p),
    .din1(g732_n_spl_1),
    .din2(g738_n_spl_0)
  );


  FA
  g_g822_n
  (
    .dout(g822_n),
    .din1(g732_p_spl_1),
    .din2(g738_p_spl_0)
  );


  LA
  g_g823_p
  (
    .dout(g823_p),
    .din1(g740_p_spl_0),
    .din2(g822_n)
  );


  FA
  g_g823_n
  (
    .dout(g823_n),
    .din1(g740_n_spl_0),
    .din2(g822_p)
  );


  LA
  g_g824_p
  (
    .dout(g824_p),
    .din1(g377_n_spl_11),
    .din2(g823_n)
  );


  FA
  g_g824_n
  (
    .dout(g824_n),
    .din1(g377_p_spl_10),
    .din2(g823_p)
  );


  LA
  g_g825_p
  (
    .dout(g825_p),
    .din1(g384_p_spl_10),
    .din2(g824_n)
  );


  FA
  g_g825_n
  (
    .dout(g825_n),
    .din1(g384_n_spl_10),
    .din2(g824_p)
  );


  LA
  g_g826_p
  (
    .dout(g826_p),
    .din1(g821_n),
    .din2(g825_n)
  );


  FA
  g_g826_n
  (
    .dout(g826_n),
    .din1(g821_p),
    .din2(g825_p)
  );


  LA
  g_g827_p
  (
    .dout(g827_p),
    .din1(g815_n),
    .din2(g826_n)
  );


  FA
  g_g827_n
  (
    .dout(g827_n),
    .din1(g815_p),
    .din2(g826_p)
  );


  LA
  g_g828_p
  (
    .dout(g828_p),
    .din1(g452_p_spl_1),
    .din2(g513_p_spl_1)
  );


  FA
  g_g828_n
  (
    .dout(g828_n),
    .din1(g452_n_spl_1),
    .din2(g513_n_spl_1)
  );


  LA
  g_g829_p
  (
    .dout(g829_p),
    .din1(G9_n_spl_11),
    .din2(g393_p_spl_111)
  );


  FA
  g_g829_n
  (
    .dout(g829_n),
    .din1(G9_p_spl_11),
    .din2(g393_n_spl_111)
  );


  LA
  g_g830_p
  (
    .dout(g830_p),
    .din1(g385_p_spl_11),
    .din2(g829_n)
  );


  FA
  g_g830_n
  (
    .dout(g830_n),
    .din1(g385_n_spl_11),
    .din2(g829_p)
  );


  LA
  g_g831_p
  (
    .dout(g831_p),
    .din1(G13_p_spl_111),
    .din2(G41_n_spl_1)
  );


  FA
  g_g831_n
  (
    .dout(g831_n),
    .din1(G13_n_spl_11),
    .din2(G41_p_spl_1)
  );


  LA
  g_g832_p
  (
    .dout(g832_p),
    .din1(g412_n_spl_111),
    .din2(g831_n)
  );


  FA
  g_g832_n
  (
    .dout(g832_n),
    .din1(g412_p_spl_111),
    .din2(g831_p)
  );


  LA
  g_g833_p
  (
    .dout(g833_p),
    .din1(G10_p_spl_11),
    .din2(G14_p_spl_111)
  );


  FA
  g_g833_n
  (
    .dout(g833_n),
    .din1(G10_n_spl_11),
    .din2(G14_n_spl_111)
  );


  LA
  g_g834_p
  (
    .dout(g834_p),
    .din1(g414_n_spl_111),
    .din2(g833_n)
  );


  FA
  g_g834_n
  (
    .dout(g834_n),
    .din1(g414_p_spl_111),
    .din2(g833_p)
  );


  LA
  g_g835_p
  (
    .dout(g835_p),
    .din1(g832_n),
    .din2(g834_n)
  );


  FA
  g_g835_n
  (
    .dout(g835_n),
    .din1(g832_p),
    .din2(g834_p)
  );


  LA
  g_g836_p
  (
    .dout(g836_p),
    .din1(g654_n_spl_),
    .din2(g835_p)
  );


  FA
  g_g836_n
  (
    .dout(g836_n),
    .din1(g654_p_spl_),
    .din2(g835_n)
  );


  LA
  g_g837_p
  (
    .dout(g837_p),
    .din1(G39_p_spl_11),
    .din2(g409_n_spl_111)
  );


  FA
  g_g837_n
  (
    .dout(g837_n),
    .din1(G39_n_spl_11),
    .din2(g409_p_spl_111)
  );


  LA
  g_g838_p
  (
    .dout(g838_p),
    .din1(G4_p_spl_1111),
    .din2(g837_n)
  );


  FA
  g_g838_n
  (
    .dout(g838_n),
    .din1(G4_n_spl_1111),
    .din2(g837_p)
  );


  LA
  g_g839_p
  (
    .dout(g839_p),
    .din1(G40_p_spl_1),
    .din2(g406_n_spl_111)
  );


  FA
  g_g839_n
  (
    .dout(g839_n),
    .din1(G40_n_spl_1),
    .din2(g406_p_spl_111)
  );


  LA
  g_g840_p
  (
    .dout(g840_p),
    .din1(G12_n_spl_11),
    .din2(g425_n_spl_11)
  );


  FA
  g_g840_n
  (
    .dout(g840_n),
    .din1(G12_p_spl_11),
    .din2(g425_p_spl_11)
  );


  LA
  g_g841_p
  (
    .dout(g841_p),
    .din1(g839_n),
    .din2(g840_n)
  );


  FA
  g_g841_n
  (
    .dout(g841_n),
    .din1(g839_p),
    .din2(g840_p)
  );


  LA
  g_g842_p
  (
    .dout(g842_p),
    .din1(g838_p),
    .din2(g841_p)
  );


  FA
  g_g842_n
  (
    .dout(g842_n),
    .din1(g838_n),
    .din2(g841_n)
  );


  LA
  g_g843_p
  (
    .dout(g843_p),
    .din1(g836_p),
    .din2(g842_p)
  );


  FA
  g_g843_n
  (
    .dout(g843_n),
    .din1(g836_n),
    .din2(g842_n)
  );


  LA
  g_g844_p
  (
    .dout(g844_p),
    .din1(G22_p_spl_11),
    .din2(g425_n_spl_11)
  );


  FA
  g_g844_n
  (
    .dout(g844_n),
    .din1(G22_n_spl_11),
    .din2(g425_p_spl_11)
  );


  LA
  g_g845_p
  (
    .dout(g845_p),
    .din1(G17_n_spl_),
    .din2(G21_n_spl_11)
  );


  FA
  g_g845_n
  (
    .dout(g845_n),
    .din1(G17_p_spl_),
    .din2(G21_p_spl_11)
  );


  LA
  g_g846_p
  (
    .dout(g846_p),
    .din1(g412_n_spl_111),
    .din2(g845_n)
  );


  FA
  g_g846_n
  (
    .dout(g846_n),
    .din1(g412_p_spl_111),
    .din2(g845_p)
  );


  LA
  g_g847_p
  (
    .dout(g847_p),
    .din1(g414_n_spl_111),
    .din2(g706_n_spl_)
  );


  FA
  g_g847_n
  (
    .dout(g847_n),
    .din1(g414_p_spl_111),
    .din2(g706_p_spl_)
  );


  LA
  g_g848_p
  (
    .dout(g848_p),
    .din1(g846_n),
    .din2(g847_n)
  );


  FA
  g_g848_n
  (
    .dout(g848_n),
    .din1(g846_p),
    .din2(g847_p)
  );


  LA
  g_g849_p
  (
    .dout(g849_p),
    .din1(g844_n),
    .din2(g848_p)
  );


  FA
  g_g849_n
  (
    .dout(g849_n),
    .din1(g844_p),
    .din2(g848_n)
  );


  LA
  g_g850_p
  (
    .dout(g850_p),
    .din1(G7_n_spl_111),
    .din2(g423_n_spl_11)
  );


  FA
  g_g850_n
  (
    .dout(g850_n),
    .din1(G7_p_spl_111),
    .din2(g423_p_spl_11)
  );


  LA
  g_g851_p
  (
    .dout(g851_p),
    .din1(G4_n_spl_1111),
    .din2(g850_n)
  );


  FA
  g_g851_n
  (
    .dout(g851_n),
    .din1(G4_p_spl_1111),
    .din2(g850_p)
  );


  LA
  g_g852_p
  (
    .dout(g852_p),
    .din1(G19_p_spl_1),
    .din2(g409_n_spl_111)
  );


  FA
  g_g852_n
  (
    .dout(g852_n),
    .din1(G19_n_spl_1),
    .din2(g409_p_spl_111)
  );


  LA
  g_g853_p
  (
    .dout(g853_p),
    .din1(G18_p_spl_1),
    .din2(g406_n_spl_111)
  );


  FA
  g_g853_n
  (
    .dout(g853_n),
    .din1(G18_n_spl_1),
    .din2(g406_p_spl_111)
  );


  LA
  g_g854_p
  (
    .dout(g854_p),
    .din1(g852_n),
    .din2(g853_n)
  );


  FA
  g_g854_n
  (
    .dout(g854_n),
    .din1(g852_p),
    .din2(g853_p)
  );


  LA
  g_g855_p
  (
    .dout(g855_p),
    .din1(g851_p),
    .din2(g854_p)
  );


  FA
  g_g855_n
  (
    .dout(g855_n),
    .din1(g851_n),
    .din2(g854_n)
  );


  LA
  g_g856_p
  (
    .dout(g856_p),
    .din1(g849_p),
    .din2(g855_p)
  );


  FA
  g_g856_n
  (
    .dout(g856_n),
    .din1(g849_n),
    .din2(g855_n)
  );


  LA
  g_g857_p
  (
    .dout(g857_p),
    .din1(g843_n),
    .din2(g856_n)
  );


  FA
  g_g857_n
  (
    .dout(g857_n),
    .din1(g843_p),
    .din2(g856_p)
  );


  LA
  g_g858_p
  (
    .dout(g858_p),
    .din1(g393_n_spl_111),
    .din2(g857_n)
  );


  FA
  g_g858_n
  (
    .dout(g858_n),
    .din1(g393_p_spl_111),
    .din2(g857_p)
  );


  LA
  g_g859_p
  (
    .dout(g859_p),
    .din1(g830_p),
    .din2(g858_n)
  );


  FA
  g_g859_n
  (
    .dout(g859_n),
    .din1(g830_n),
    .din2(g858_p)
  );


  LA
  g_g860_p
  (
    .dout(g860_p),
    .din1(g828_n),
    .din2(g859_p)
  );


  FA
  g_g860_n
  (
    .dout(g860_n),
    .din1(g828_p),
    .din2(g859_n)
  );


  LA
  g_g861_p
  (
    .dout(g861_p),
    .din1(g738_p_spl_1),
    .din2(g740_p_spl_)
  );


  FA
  g_g861_n
  (
    .dout(g861_n),
    .din1(g738_n_spl_1),
    .din2(g740_n_spl_)
  );


  LA
  g_g862_p
  (
    .dout(g862_p),
    .din1(g384_n_spl_1),
    .din2(g738_n_spl_1)
  );


  FA
  g_g862_n
  (
    .dout(g862_n),
    .din1(g384_p_spl_1),
    .din2(g738_p_spl_1)
  );


  LA
  g_g863_p
  (
    .dout(g863_p),
    .din1(g377_n_spl_11),
    .din2(g741_n_spl_)
  );


  FA
  g_g863_n
  (
    .dout(g863_n),
    .din1(g377_p_spl_1),
    .din2(g741_p_spl_)
  );


  LA
  g_g864_p
  (
    .dout(g864_p),
    .din1(g862_n),
    .din2(g863_n)
  );


  FA
  g_g864_n
  (
    .dout(g864_n),
    .din1(g862_p),
    .din2(g863_p)
  );


  LA
  g_g865_p
  (
    .dout(g865_p),
    .din1(g861_n),
    .din2(g864_n)
  );


  FA
  g_g865_n
  (
    .dout(g865_n),
    .din1(g861_p),
    .din2(g864_p)
  );


  LA
  g_g866_p
  (
    .dout(g866_p),
    .din1(g860_n),
    .din2(g865_n)
  );


  FA
  g_g866_n
  (
    .dout(g866_n),
    .din1(g860_p),
    .din2(g865_p)
  );


  LA
  g_g867_p
  (
    .dout(g867_p),
    .din1(g626_p_spl_),
    .din2(g722_p_spl_)
  );


  FA
  g_g867_n
  (
    .dout(g867_n),
    .din1(g626_n_spl_0),
    .din2(g722_n_spl_0)
  );


  LA
  g_g868_p
  (
    .dout(g868_p),
    .din1(g778_p_spl_),
    .din2(g827_p_spl_)
  );


  FA
  g_g868_n
  (
    .dout(g868_n),
    .din1(g778_n_spl_0),
    .din2(g827_n_spl_0)
  );


  LA
  g_g869_p
  (
    .dout(g869_p),
    .din1(g509_p_spl_),
    .din2(g866_p_spl_)
  );


  FA
  g_g869_n
  (
    .dout(g869_n),
    .din1(g509_n_spl_0),
    .din2(g866_n_spl_0)
  );


  LA
  g_g870_p
  (
    .dout(g870_p),
    .din1(g451_p_spl_),
    .din2(g679_p_spl_)
  );


  FA
  g_g870_n
  (
    .dout(g870_n),
    .din1(g451_n_spl_0),
    .din2(g679_n_spl_0)
  );


  FA
  g_g871_n
  (
    .dout(g871_n),
    .din1(g869_n_spl_),
    .din2(g870_n_spl_)
  );


  FA
  g_g872_n
  (
    .dout(g872_n),
    .din1(g868_n_spl_0),
    .din2(g871_n)
  );


  FA
  g_g873_n
  (
    .dout(g873_n),
    .din1(g867_n_spl_),
    .din2(g872_n)
  );


  LA
  g_g874_p
  (
    .dout(g874_p),
    .din1(G27_p_spl_0),
    .din2(G48_p_spl_)
  );


  FA
  g_g874_n
  (
    .dout(g874_n),
    .din1(G27_n_spl_),
    .din2(G48_n_spl_)
  );


  FA
  g_g875_n
  (
    .dout(g875_n),
    .din1(g868_n_spl_0),
    .din2(g874_n_spl_)
  );


  LA
  g_g876_p
  (
    .dout(g876_p),
    .din1(G27_p_spl_),
    .din2(g875_n)
  );


  LA
  g_g877_p
  (
    .dout(g877_p),
    .din1(g873_n_spl_),
    .din2(g876_p)
  );


  LA
  g_g878_p
  (
    .dout(g878_p),
    .din1(g451_n_spl_0),
    .din2(g679_n_spl_0)
  );


  FA
  g_g878_n
  (
    .dout(g878_n),
    .din1(g451_p_spl_),
    .din2(g679_p_spl_)
  );


  LA
  g_g879_p
  (
    .dout(g879_p),
    .din1(g870_n_spl_),
    .din2(g878_n)
  );


  FA
  g_g879_n
  (
    .dout(g879_n),
    .din1(g870_p),
    .din2(g878_p)
  );


  LA
  g_g880_p
  (
    .dout(g880_p),
    .din1(g626_n_spl_0),
    .din2(g722_n_spl_0)
  );


  FA
  g_g880_n
  (
    .dout(g880_n),
    .din1(g626_p_spl_),
    .din2(g722_p_spl_)
  );


  LA
  g_g881_p
  (
    .dout(g881_p),
    .din1(g867_n_spl_),
    .din2(g880_n)
  );


  FA
  g_g881_n
  (
    .dout(g881_n),
    .din1(g867_p),
    .din2(g880_p)
  );


  LA
  g_g882_p
  (
    .dout(g882_p),
    .din1(g879_p_spl_),
    .din2(g881_n_spl_)
  );


  FA
  g_g882_n
  (
    .dout(g882_n),
    .din1(g879_n_spl_),
    .din2(g881_p_spl_)
  );


  LA
  g_g883_p
  (
    .dout(g883_p),
    .din1(g879_n_spl_),
    .din2(g881_p_spl_)
  );


  FA
  g_g883_n
  (
    .dout(g883_n),
    .din1(g879_p_spl_),
    .din2(g881_n_spl_)
  );


  LA
  g_g884_p
  (
    .dout(g884_p),
    .din1(g882_n),
    .din2(g883_n)
  );


  FA
  g_g884_n
  (
    .dout(g884_n),
    .din1(g882_p),
    .din2(g883_p)
  );


  LA
  g_g885_p
  (
    .dout(g885_p),
    .din1(g509_n_spl_0),
    .din2(g866_n_spl_0)
  );


  FA
  g_g885_n
  (
    .dout(g885_n),
    .din1(g509_p_spl_),
    .din2(g866_p_spl_)
  );


  LA
  g_g886_p
  (
    .dout(g886_p),
    .din1(g869_n_spl_),
    .din2(g885_n)
  );


  FA
  g_g886_n
  (
    .dout(g886_n),
    .din1(g869_p),
    .din2(g885_p)
  );


  LA
  g_g887_p
  (
    .dout(g887_p),
    .din1(g778_n_spl_0),
    .din2(g827_n_spl_0)
  );


  FA
  g_g887_n
  (
    .dout(g887_n),
    .din1(g778_p_spl_),
    .din2(g827_p_spl_)
  );


  LA
  g_g888_p
  (
    .dout(g888_p),
    .din1(g868_n_spl_),
    .din2(g887_n)
  );


  FA
  g_g888_n
  (
    .dout(g888_n),
    .din1(g868_p),
    .din2(g887_p)
  );


  LA
  g_g889_p
  (
    .dout(g889_p),
    .din1(G50_n_spl_),
    .din2(g888_n_spl_0)
  );


  FA
  g_g889_n
  (
    .dout(g889_n),
    .din1(G50_p_spl_),
    .din2(g888_p_spl_0)
  );


  LA
  g_g890_p
  (
    .dout(g890_p),
    .din1(G50_p_spl_),
    .din2(g888_p_spl_0)
  );


  FA
  g_g890_n
  (
    .dout(g890_n),
    .din1(G50_n_spl_),
    .din2(g888_n_spl_0)
  );


  LA
  g_g891_p
  (
    .dout(g891_p),
    .din1(g874_n_spl_),
    .din2(g890_n)
  );


  FA
  g_g891_n
  (
    .dout(g891_n),
    .din1(g874_p),
    .din2(g890_p)
  );


  LA
  g_g892_p
  (
    .dout(g892_p),
    .din1(g889_n),
    .din2(g891_p)
  );


  FA
  g_g892_n
  (
    .dout(g892_n),
    .din1(g889_p),
    .din2(g891_n)
  );


  LA
  g_g893_p
  (
    .dout(g893_p),
    .din1(g886_p_spl_0),
    .din2(g892_n_spl_)
  );


  FA
  g_g893_n
  (
    .dout(g893_n),
    .din1(g886_n_spl_0),
    .din2(g892_p_spl_)
  );


  LA
  g_g894_p
  (
    .dout(g894_p),
    .din1(g886_n_spl_0),
    .din2(g892_p_spl_)
  );


  FA
  g_g894_n
  (
    .dout(g894_n),
    .din1(g886_p_spl_0),
    .din2(g892_n_spl_)
  );


  LA
  g_g895_p
  (
    .dout(g895_p),
    .din1(g893_n),
    .din2(g894_n)
  );


  FA
  g_g895_n
  (
    .dout(g895_n),
    .din1(g893_p),
    .din2(g894_p)
  );


  LA
  g_g896_p
  (
    .dout(g896_p),
    .din1(g884_n_spl_),
    .din2(g895_p)
  );


  LA
  g_g897_p
  (
    .dout(g897_p),
    .din1(g884_p_spl_),
    .din2(g895_n)
  );


  FA
  g_g898_n
  (
    .dout(g898_n),
    .din1(g896_p),
    .din2(g897_p)
  );


  LA
  g_g899_p
  (
    .dout(g899_p),
    .din1(g886_n_spl_1),
    .din2(g888_n_spl_1)
  );


  FA
  g_g899_n
  (
    .dout(g899_n),
    .din1(g886_p_spl_1),
    .din2(g888_p_spl_1)
  );


  LA
  g_g900_p
  (
    .dout(g900_p),
    .din1(g886_p_spl_1),
    .din2(g888_p_spl_1)
  );


  FA
  g_g900_n
  (
    .dout(g900_n),
    .din1(g886_n_spl_1),
    .din2(g888_n_spl_1)
  );


  LA
  g_g901_p
  (
    .dout(g901_p),
    .din1(g899_n),
    .din2(g900_n)
  );


  FA
  g_g901_n
  (
    .dout(g901_n),
    .din1(g899_p),
    .din2(g900_p)
  );


  FA
  g_g902_n
  (
    .dout(g902_n),
    .din1(g884_p_spl_),
    .din2(g901_p)
  );


  FA
  g_g903_n
  (
    .dout(g903_n),
    .din1(g884_n_spl_),
    .din2(g901_n)
  );


  LA
  g_g904_p
  (
    .dout(g904_p),
    .din1(g902_n),
    .din2(g903_n)
  );


  buf

  (
    G3519_p,
    g53_p
  );


  buf

  (
    G3520_p,
    g55_n_spl_
  );


  buf

  (
    G3521_p,
    g84_p
  );


  buf

  (
    G3522_p,
    g105_p
  );


  buf

  (
    G3523_p,
    g125_n
  );


  buf

  (
    G3524_p,
    g350_p
  );


  buf

  (
    G3525_p,
    g364_n
  );


  buf

  (
    G3526_p,
    g376_p_spl_
  );


  buf

  (
    G3527_p,
    g381_n
  );


  buf

  (
    G3528_p,
    g451_n_spl_
  );


  buf

  (
    G3529_p,
    g509_n_spl_
  );


  buf

  (
    G3530_p,
    g551_n
  );


  buf

  (
    G3531_p,
    g626_n_spl_
  );


  buf

  (
    G3532_p,
    g679_n_spl_
  );


  buf

  (
    G3533_p,
    g722_n_spl_
  );


  buf

  (
    G3534_p,
    g778_n_spl_
  );


  buf

  (
    G3535_p,
    g827_n_spl_
  );


  buf

  (
    G3536_p,
    g866_n_spl_
  );


  buf

  (
    G3537_p,
    g873_n_spl_
  );


  buf

  (
    G3538_n,
    g877_p
  );


  buf

  (
    G3539_p,
    g898_n
  );


  buf

  (
    G3540_p,
    g904_p
  );


  buf

  (
    G7_n_spl_,
    G7_n
  );


  buf

  (
    G7_n_spl_0,
    G7_n_spl_
  );


  buf

  (
    G7_n_spl_00,
    G7_n_spl_0
  );


  buf

  (
    G7_n_spl_000,
    G7_n_spl_00
  );


  buf

  (
    G7_n_spl_0000,
    G7_n_spl_000
  );


  buf

  (
    G7_n_spl_001,
    G7_n_spl_00
  );


  buf

  (
    G7_n_spl_01,
    G7_n_spl_0
  );


  buf

  (
    G7_n_spl_010,
    G7_n_spl_01
  );


  buf

  (
    G7_n_spl_011,
    G7_n_spl_01
  );


  buf

  (
    G7_n_spl_1,
    G7_n_spl_
  );


  buf

  (
    G7_n_spl_10,
    G7_n_spl_1
  );


  buf

  (
    G7_n_spl_100,
    G7_n_spl_10
  );


  buf

  (
    G7_n_spl_101,
    G7_n_spl_10
  );


  buf

  (
    G7_n_spl_11,
    G7_n_spl_1
  );


  buf

  (
    G7_n_spl_110,
    G7_n_spl_11
  );


  buf

  (
    G7_n_spl_111,
    G7_n_spl_11
  );


  buf

  (
    G8_n_spl_,
    G8_n
  );


  buf

  (
    G8_n_spl_0,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_00,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_000,
    G8_n_spl_00
  );


  buf

  (
    G8_n_spl_001,
    G8_n_spl_00
  );


  buf

  (
    G8_n_spl_01,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_010,
    G8_n_spl_01
  );


  buf

  (
    G8_n_spl_011,
    G8_n_spl_01
  );


  buf

  (
    G8_n_spl_1,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_10,
    G8_n_spl_1
  );


  buf

  (
    G8_n_spl_100,
    G8_n_spl_10
  );


  buf

  (
    G8_n_spl_101,
    G8_n_spl_10
  );


  buf

  (
    G8_n_spl_11,
    G8_n_spl_1
  );


  buf

  (
    G8_n_spl_110,
    G8_n_spl_11
  );


  buf

  (
    G7_p_spl_,
    G7_p
  );


  buf

  (
    G7_p_spl_0,
    G7_p_spl_
  );


  buf

  (
    G7_p_spl_00,
    G7_p_spl_0
  );


  buf

  (
    G7_p_spl_000,
    G7_p_spl_00
  );


  buf

  (
    G7_p_spl_0000,
    G7_p_spl_000
  );


  buf

  (
    G7_p_spl_0001,
    G7_p_spl_000
  );


  buf

  (
    G7_p_spl_001,
    G7_p_spl_00
  );


  buf

  (
    G7_p_spl_01,
    G7_p_spl_0
  );


  buf

  (
    G7_p_spl_010,
    G7_p_spl_01
  );


  buf

  (
    G7_p_spl_011,
    G7_p_spl_01
  );


  buf

  (
    G7_p_spl_1,
    G7_p_spl_
  );


  buf

  (
    G7_p_spl_10,
    G7_p_spl_1
  );


  buf

  (
    G7_p_spl_100,
    G7_p_spl_10
  );


  buf

  (
    G7_p_spl_101,
    G7_p_spl_10
  );


  buf

  (
    G7_p_spl_11,
    G7_p_spl_1
  );


  buf

  (
    G7_p_spl_110,
    G7_p_spl_11
  );


  buf

  (
    G7_p_spl_111,
    G7_p_spl_11
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_00,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_000,
    G8_p_spl_00
  );


  buf

  (
    G8_p_spl_001,
    G8_p_spl_00
  );


  buf

  (
    G8_p_spl_01,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_010,
    G8_p_spl_01
  );


  buf

  (
    G8_p_spl_011,
    G8_p_spl_01
  );


  buf

  (
    G8_p_spl_1,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_10,
    G8_p_spl_1
  );


  buf

  (
    G8_p_spl_100,
    G8_p_spl_10
  );


  buf

  (
    G8_p_spl_101,
    G8_p_spl_10
  );


  buf

  (
    G8_p_spl_11,
    G8_p_spl_1
  );


  buf

  (
    G8_p_spl_110,
    G8_p_spl_11
  );


  buf

  (
    G8_p_spl_111,
    G8_p_spl_11
  );


  buf

  (
    G9_n_spl_,
    G9_n
  );


  buf

  (
    G9_n_spl_0,
    G9_n_spl_
  );


  buf

  (
    G9_n_spl_00,
    G9_n_spl_0
  );


  buf

  (
    G9_n_spl_000,
    G9_n_spl_00
  );


  buf

  (
    G9_n_spl_001,
    G9_n_spl_00
  );


  buf

  (
    G9_n_spl_01,
    G9_n_spl_0
  );


  buf

  (
    G9_n_spl_010,
    G9_n_spl_01
  );


  buf

  (
    G9_n_spl_011,
    G9_n_spl_01
  );


  buf

  (
    G9_n_spl_1,
    G9_n_spl_
  );


  buf

  (
    G9_n_spl_10,
    G9_n_spl_1
  );


  buf

  (
    G9_n_spl_100,
    G9_n_spl_10
  );


  buf

  (
    G9_n_spl_101,
    G9_n_spl_10
  );


  buf

  (
    G9_n_spl_11,
    G9_n_spl_1
  );


  buf

  (
    G9_n_spl_110,
    G9_n_spl_11
  );


  buf

  (
    g51_p_spl_,
    g51_p
  );


  buf

  (
    G9_p_spl_,
    G9_p
  );


  buf

  (
    G9_p_spl_0,
    G9_p_spl_
  );


  buf

  (
    G9_p_spl_00,
    G9_p_spl_0
  );


  buf

  (
    G9_p_spl_000,
    G9_p_spl_00
  );


  buf

  (
    G9_p_spl_001,
    G9_p_spl_00
  );


  buf

  (
    G9_p_spl_01,
    G9_p_spl_0
  );


  buf

  (
    G9_p_spl_010,
    G9_p_spl_01
  );


  buf

  (
    G9_p_spl_011,
    G9_p_spl_01
  );


  buf

  (
    G9_p_spl_1,
    G9_p_spl_
  );


  buf

  (
    G9_p_spl_10,
    G9_p_spl_1
  );


  buf

  (
    G9_p_spl_100,
    G9_p_spl_10
  );


  buf

  (
    G9_p_spl_101,
    G9_p_spl_10
  );


  buf

  (
    G9_p_spl_11,
    G9_p_spl_1
  );


  buf

  (
    G9_p_spl_110,
    G9_p_spl_11
  );


  buf

  (
    g51_n_spl_,
    g51_n
  );


  buf

  (
    G10_n_spl_,
    G10_n
  );


  buf

  (
    G10_n_spl_0,
    G10_n_spl_
  );


  buf

  (
    G10_n_spl_00,
    G10_n_spl_0
  );


  buf

  (
    G10_n_spl_000,
    G10_n_spl_00
  );


  buf

  (
    G10_n_spl_001,
    G10_n_spl_00
  );


  buf

  (
    G10_n_spl_01,
    G10_n_spl_0
  );


  buf

  (
    G10_n_spl_010,
    G10_n_spl_01
  );


  buf

  (
    G10_n_spl_011,
    G10_n_spl_01
  );


  buf

  (
    G10_n_spl_1,
    G10_n_spl_
  );


  buf

  (
    G10_n_spl_10,
    G10_n_spl_1
  );


  buf

  (
    G10_n_spl_100,
    G10_n_spl_10
  );


  buf

  (
    G10_n_spl_101,
    G10_n_spl_10
  );


  buf

  (
    G10_n_spl_11,
    G10_n_spl_1
  );


  buf

  (
    G10_n_spl_110,
    G10_n_spl_11
  );


  buf

  (
    g52_p_spl_,
    g52_p
  );


  buf

  (
    G12_n_spl_,
    G12_n
  );


  buf

  (
    G12_n_spl_0,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_00,
    G12_n_spl_0
  );


  buf

  (
    G12_n_spl_000,
    G12_n_spl_00
  );


  buf

  (
    G12_n_spl_001,
    G12_n_spl_00
  );


  buf

  (
    G12_n_spl_01,
    G12_n_spl_0
  );


  buf

  (
    G12_n_spl_010,
    G12_n_spl_01
  );


  buf

  (
    G12_n_spl_011,
    G12_n_spl_01
  );


  buf

  (
    G12_n_spl_1,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_10,
    G12_n_spl_1
  );


  buf

  (
    G12_n_spl_100,
    G12_n_spl_10
  );


  buf

  (
    G12_n_spl_101,
    G12_n_spl_10
  );


  buf

  (
    G12_n_spl_11,
    G12_n_spl_1
  );


  buf

  (
    G13_n_spl_,
    G13_n
  );


  buf

  (
    G13_n_spl_0,
    G13_n_spl_
  );


  buf

  (
    G13_n_spl_00,
    G13_n_spl_0
  );


  buf

  (
    G13_n_spl_000,
    G13_n_spl_00
  );


  buf

  (
    G13_n_spl_001,
    G13_n_spl_00
  );


  buf

  (
    G13_n_spl_01,
    G13_n_spl_0
  );


  buf

  (
    G13_n_spl_010,
    G13_n_spl_01
  );


  buf

  (
    G13_n_spl_011,
    G13_n_spl_01
  );


  buf

  (
    G13_n_spl_1,
    G13_n_spl_
  );


  buf

  (
    G13_n_spl_10,
    G13_n_spl_1
  );


  buf

  (
    G13_n_spl_100,
    G13_n_spl_10
  );


  buf

  (
    G13_n_spl_101,
    G13_n_spl_10
  );


  buf

  (
    G13_n_spl_11,
    G13_n_spl_1
  );


  buf

  (
    G13_n_spl_110,
    G13_n_spl_11
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G12_p_spl_0,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_00,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_000,
    G12_p_spl_00
  );


  buf

  (
    G12_p_spl_001,
    G12_p_spl_00
  );


  buf

  (
    G12_p_spl_01,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_010,
    G12_p_spl_01
  );


  buf

  (
    G12_p_spl_011,
    G12_p_spl_01
  );


  buf

  (
    G12_p_spl_1,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_10,
    G12_p_spl_1
  );


  buf

  (
    G12_p_spl_100,
    G12_p_spl_10
  );


  buf

  (
    G12_p_spl_101,
    G12_p_spl_10
  );


  buf

  (
    G12_p_spl_11,
    G12_p_spl_1
  );


  buf

  (
    G12_p_spl_110,
    G12_p_spl_11
  );


  buf

  (
    G13_p_spl_,
    G13_p
  );


  buf

  (
    G13_p_spl_0,
    G13_p_spl_
  );


  buf

  (
    G13_p_spl_00,
    G13_p_spl_0
  );


  buf

  (
    G13_p_spl_000,
    G13_p_spl_00
  );


  buf

  (
    G13_p_spl_001,
    G13_p_spl_00
  );


  buf

  (
    G13_p_spl_01,
    G13_p_spl_0
  );


  buf

  (
    G13_p_spl_010,
    G13_p_spl_01
  );


  buf

  (
    G13_p_spl_011,
    G13_p_spl_01
  );


  buf

  (
    G13_p_spl_1,
    G13_p_spl_
  );


  buf

  (
    G13_p_spl_10,
    G13_p_spl_1
  );


  buf

  (
    G13_p_spl_100,
    G13_p_spl_10
  );


  buf

  (
    G13_p_spl_101,
    G13_p_spl_10
  );


  buf

  (
    G13_p_spl_11,
    G13_p_spl_1
  );


  buf

  (
    G13_p_spl_110,
    G13_p_spl_11
  );


  buf

  (
    G13_p_spl_111,
    G13_p_spl_11
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    G11_p_spl_0,
    G11_p_spl_
  );


  buf

  (
    G11_p_spl_00,
    G11_p_spl_0
  );


  buf

  (
    G11_p_spl_000,
    G11_p_spl_00
  );


  buf

  (
    G11_p_spl_001,
    G11_p_spl_00
  );


  buf

  (
    G11_p_spl_01,
    G11_p_spl_0
  );


  buf

  (
    G11_p_spl_010,
    G11_p_spl_01
  );


  buf

  (
    G11_p_spl_011,
    G11_p_spl_01
  );


  buf

  (
    G11_p_spl_1,
    G11_p_spl_
  );


  buf

  (
    G11_p_spl_10,
    G11_p_spl_1
  );


  buf

  (
    G11_p_spl_100,
    G11_p_spl_10
  );


  buf

  (
    G11_p_spl_101,
    G11_p_spl_10
  );


  buf

  (
    G11_p_spl_11,
    G11_p_spl_1
  );


  buf

  (
    g54_n_spl_,
    g54_n
  );


  buf

  (
    G11_n_spl_,
    G11_n
  );


  buf

  (
    G11_n_spl_0,
    G11_n_spl_
  );


  buf

  (
    G11_n_spl_00,
    G11_n_spl_0
  );


  buf

  (
    G11_n_spl_000,
    G11_n_spl_00
  );


  buf

  (
    G11_n_spl_001,
    G11_n_spl_00
  );


  buf

  (
    G11_n_spl_01,
    G11_n_spl_0
  );


  buf

  (
    G11_n_spl_010,
    G11_n_spl_01
  );


  buf

  (
    G11_n_spl_011,
    G11_n_spl_01
  );


  buf

  (
    G11_n_spl_1,
    G11_n_spl_
  );


  buf

  (
    G11_n_spl_10,
    G11_n_spl_1
  );


  buf

  (
    G11_n_spl_100,
    G11_n_spl_10
  );


  buf

  (
    G11_n_spl_11,
    G11_n_spl_1
  );


  buf

  (
    g54_p_spl_,
    g54_p
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G1_n_spl_0,
    G1_n_spl_
  );


  buf

  (
    G1_n_spl_00,
    G1_n_spl_0
  );


  buf

  (
    G1_n_spl_000,
    G1_n_spl_00
  );


  buf

  (
    G1_n_spl_001,
    G1_n_spl_00
  );


  buf

  (
    G1_n_spl_01,
    G1_n_spl_0
  );


  buf

  (
    G1_n_spl_010,
    G1_n_spl_01
  );


  buf

  (
    G1_n_spl_1,
    G1_n_spl_
  );


  buf

  (
    G1_n_spl_10,
    G1_n_spl_1
  );


  buf

  (
    G1_n_spl_11,
    G1_n_spl_1
  );


  buf

  (
    G3_n_spl_,
    G3_n
  );


  buf

  (
    G3_n_spl_0,
    G3_n_spl_
  );


  buf

  (
    G3_n_spl_00,
    G3_n_spl_0
  );


  buf

  (
    G3_n_spl_000,
    G3_n_spl_00
  );


  buf

  (
    G3_n_spl_0000,
    G3_n_spl_000
  );


  buf

  (
    G3_n_spl_0001,
    G3_n_spl_000
  );


  buf

  (
    G3_n_spl_001,
    G3_n_spl_00
  );


  buf

  (
    G3_n_spl_0010,
    G3_n_spl_001
  );


  buf

  (
    G3_n_spl_01,
    G3_n_spl_0
  );


  buf

  (
    G3_n_spl_010,
    G3_n_spl_01
  );


  buf

  (
    G3_n_spl_011,
    G3_n_spl_01
  );


  buf

  (
    G3_n_spl_1,
    G3_n_spl_
  );


  buf

  (
    G3_n_spl_10,
    G3_n_spl_1
  );


  buf

  (
    G3_n_spl_100,
    G3_n_spl_10
  );


  buf

  (
    G3_n_spl_101,
    G3_n_spl_10
  );


  buf

  (
    G3_n_spl_11,
    G3_n_spl_1
  );


  buf

  (
    G3_n_spl_110,
    G3_n_spl_11
  );


  buf

  (
    G3_n_spl_111,
    G3_n_spl_11
  );


  buf

  (
    G34_n_spl_,
    G34_n
  );


  buf

  (
    G34_n_spl_0,
    G34_n_spl_
  );


  buf

  (
    G34_n_spl_00,
    G34_n_spl_0
  );


  buf

  (
    G34_n_spl_01,
    G34_n_spl_0
  );


  buf

  (
    G34_n_spl_1,
    G34_n_spl_
  );


  buf

  (
    G34_n_spl_10,
    G34_n_spl_1
  );


  buf

  (
    G32_n_spl_,
    G32_n
  );


  buf

  (
    G32_n_spl_0,
    G32_n_spl_
  );


  buf

  (
    G32_n_spl_00,
    G32_n_spl_0
  );


  buf

  (
    G32_n_spl_01,
    G32_n_spl_0
  );


  buf

  (
    G32_n_spl_1,
    G32_n_spl_
  );


  buf

  (
    G36_n_spl_,
    G36_n
  );


  buf

  (
    G36_n_spl_0,
    G36_n_spl_
  );


  buf

  (
    G36_n_spl_00,
    G36_n_spl_0
  );


  buf

  (
    G36_n_spl_01,
    G36_n_spl_0
  );


  buf

  (
    G36_n_spl_1,
    G36_n_spl_
  );


  buf

  (
    G10_p_spl_,
    G10_p
  );


  buf

  (
    G10_p_spl_0,
    G10_p_spl_
  );


  buf

  (
    G10_p_spl_00,
    G10_p_spl_0
  );


  buf

  (
    G10_p_spl_000,
    G10_p_spl_00
  );


  buf

  (
    G10_p_spl_001,
    G10_p_spl_00
  );


  buf

  (
    G10_p_spl_01,
    G10_p_spl_0
  );


  buf

  (
    G10_p_spl_010,
    G10_p_spl_01
  );


  buf

  (
    G10_p_spl_011,
    G10_p_spl_01
  );


  buf

  (
    G10_p_spl_1,
    G10_p_spl_
  );


  buf

  (
    G10_p_spl_10,
    G10_p_spl_1
  );


  buf

  (
    G10_p_spl_100,
    G10_p_spl_10
  );


  buf

  (
    G10_p_spl_101,
    G10_p_spl_10
  );


  buf

  (
    G10_p_spl_11,
    G10_p_spl_1
  );


  buf

  (
    G33_n_spl_,
    G33_n
  );


  buf

  (
    G33_n_spl_0,
    G33_n_spl_
  );


  buf

  (
    G33_n_spl_00,
    G33_n_spl_0
  );


  buf

  (
    G33_n_spl_01,
    G33_n_spl_0
  );


  buf

  (
    G33_n_spl_1,
    G33_n_spl_
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G14_p_spl_0,
    G14_p_spl_
  );


  buf

  (
    G14_p_spl_00,
    G14_p_spl_0
  );


  buf

  (
    G14_p_spl_000,
    G14_p_spl_00
  );


  buf

  (
    G14_p_spl_001,
    G14_p_spl_00
  );


  buf

  (
    G14_p_spl_01,
    G14_p_spl_0
  );


  buf

  (
    G14_p_spl_010,
    G14_p_spl_01
  );


  buf

  (
    G14_p_spl_011,
    G14_p_spl_01
  );


  buf

  (
    G14_p_spl_1,
    G14_p_spl_
  );


  buf

  (
    G14_p_spl_10,
    G14_p_spl_1
  );


  buf

  (
    G14_p_spl_100,
    G14_p_spl_10
  );


  buf

  (
    G14_p_spl_101,
    G14_p_spl_10
  );


  buf

  (
    G14_p_spl_11,
    G14_p_spl_1
  );


  buf

  (
    G14_p_spl_110,
    G14_p_spl_11
  );


  buf

  (
    G14_p_spl_111,
    G14_p_spl_11
  );


  buf

  (
    G37_n_spl_,
    G37_n
  );


  buf

  (
    G37_n_spl_0,
    G37_n_spl_
  );


  buf

  (
    G37_n_spl_1,
    G37_n_spl_
  );


  buf

  (
    G31_n_spl_,
    G31_n
  );


  buf

  (
    G31_n_spl_0,
    G31_n_spl_
  );


  buf

  (
    G31_n_spl_00,
    G31_n_spl_0
  );


  buf

  (
    G31_n_spl_01,
    G31_n_spl_0
  );


  buf

  (
    G31_n_spl_1,
    G31_n_spl_
  );


  buf

  (
    G35_n_spl_,
    G35_n
  );


  buf

  (
    G35_n_spl_0,
    G35_n_spl_
  );


  buf

  (
    G35_n_spl_00,
    G35_n_spl_0
  );


  buf

  (
    G35_n_spl_01,
    G35_n_spl_0
  );


  buf

  (
    G35_n_spl_1,
    G35_n_spl_
  );


  buf

  (
    G35_n_spl_10,
    G35_n_spl_1
  );


  buf

  (
    G30_n_spl_,
    G30_n
  );


  buf

  (
    G30_n_spl_0,
    G30_n_spl_
  );


  buf

  (
    G30_n_spl_00,
    G30_n_spl_0
  );


  buf

  (
    G30_n_spl_01,
    G30_n_spl_0
  );


  buf

  (
    G30_n_spl_1,
    G30_n_spl_
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G2_p_spl_0,
    G2_p_spl_
  );


  buf

  (
    G2_p_spl_00,
    G2_p_spl_0
  );


  buf

  (
    G2_p_spl_1,
    G2_p_spl_
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G1_p_spl_0,
    G1_p_spl_
  );


  buf

  (
    G1_p_spl_00,
    G1_p_spl_0
  );


  buf

  (
    G1_p_spl_000,
    G1_p_spl_00
  );


  buf

  (
    G1_p_spl_01,
    G1_p_spl_0
  );


  buf

  (
    G1_p_spl_1,
    G1_p_spl_
  );


  buf

  (
    G1_p_spl_10,
    G1_p_spl_1
  );


  buf

  (
    G1_p_spl_11,
    G1_p_spl_1
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G2_n_spl_0,
    G2_n_spl_
  );


  buf

  (
    G2_n_spl_00,
    G2_n_spl_0
  );


  buf

  (
    G2_n_spl_1,
    G2_n_spl_
  );


  buf

  (
    g73_p_spl_,
    g73_p
  );


  buf

  (
    g73_p_spl_0,
    g73_p_spl_
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G3_p_spl_0,
    G3_p_spl_
  );


  buf

  (
    G3_p_spl_00,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_000,
    G3_p_spl_00
  );


  buf

  (
    G3_p_spl_0000,
    G3_p_spl_000
  );


  buf

  (
    G3_p_spl_0001,
    G3_p_spl_000
  );


  buf

  (
    G3_p_spl_001,
    G3_p_spl_00
  );


  buf

  (
    G3_p_spl_01,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_010,
    G3_p_spl_01
  );


  buf

  (
    G3_p_spl_011,
    G3_p_spl_01
  );


  buf

  (
    G3_p_spl_1,
    G3_p_spl_
  );


  buf

  (
    G3_p_spl_10,
    G3_p_spl_1
  );


  buf

  (
    G3_p_spl_100,
    G3_p_spl_10
  );


  buf

  (
    G3_p_spl_101,
    G3_p_spl_10
  );


  buf

  (
    G3_p_spl_11,
    G3_p_spl_1
  );


  buf

  (
    G3_p_spl_110,
    G3_p_spl_11
  );


  buf

  (
    G3_p_spl_111,
    G3_p_spl_11
  );


  buf

  (
    g73_n_spl_,
    g73_n
  );


  buf

  (
    g73_n_spl_0,
    g73_n_spl_
  );


  buf

  (
    g75_n_spl_,
    g75_n
  );


  buf

  (
    g75_p_spl_,
    g75_p
  );


  buf

  (
    g74_n_spl_,
    g74_n
  );


  buf

  (
    g76_n_spl_,
    g76_n
  );


  buf

  (
    g78_p_spl_,
    g78_p
  );


  buf

  (
    g78_n_spl_,
    g78_n
  );


  buf

  (
    g79_n_spl_,
    g79_n
  );


  buf

  (
    g79_n_spl_0,
    g79_n_spl_
  );


  buf

  (
    g79_n_spl_1,
    g79_n_spl_
  );


  buf

  (
    G36_p_spl_,
    G36_p
  );


  buf

  (
    G36_p_spl_0,
    G36_p_spl_
  );


  buf

  (
    G36_p_spl_1,
    G36_p_spl_
  );


  buf

  (
    G37_p_spl_,
    G37_p
  );


  buf

  (
    G37_p_spl_0,
    G37_p_spl_
  );


  buf

  (
    G34_p_spl_,
    G34_p
  );


  buf

  (
    G34_p_spl_0,
    G34_p_spl_
  );


  buf

  (
    G34_p_spl_00,
    G34_p_spl_0
  );


  buf

  (
    G34_p_spl_1,
    G34_p_spl_
  );


  buf

  (
    G35_p_spl_,
    G35_p
  );


  buf

  (
    G35_p_spl_0,
    G35_p_spl_
  );


  buf

  (
    G35_p_spl_00,
    G35_p_spl_0
  );


  buf

  (
    G35_p_spl_1,
    G35_p_spl_
  );


  buf

  (
    g87_p_spl_,
    g87_p
  );


  buf

  (
    g90_n_spl_,
    g90_n
  );


  buf

  (
    g87_n_spl_,
    g87_n
  );


  buf

  (
    g90_p_spl_,
    g90_p
  );


  buf

  (
    G32_p_spl_,
    G32_p
  );


  buf

  (
    G32_p_spl_0,
    G32_p_spl_
  );


  buf

  (
    G32_p_spl_00,
    G32_p_spl_0
  );


  buf

  (
    G32_p_spl_1,
    G32_p_spl_
  );


  buf

  (
    G33_p_spl_,
    G33_p
  );


  buf

  (
    G33_p_spl_0,
    G33_p_spl_
  );


  buf

  (
    G33_p_spl_00,
    G33_p_spl_0
  );


  buf

  (
    G33_p_spl_1,
    G33_p_spl_
  );


  buf

  (
    G30_p_spl_,
    G30_p
  );


  buf

  (
    G30_p_spl_0,
    G30_p_spl_
  );


  buf

  (
    G30_p_spl_00,
    G30_p_spl_0
  );


  buf

  (
    G30_p_spl_1,
    G30_p_spl_
  );


  buf

  (
    G31_p_spl_,
    G31_p
  );


  buf

  (
    G31_p_spl_0,
    G31_p_spl_
  );


  buf

  (
    G31_p_spl_00,
    G31_p_spl_0
  );


  buf

  (
    G31_p_spl_1,
    G31_p_spl_
  );


  buf

  (
    g96_n_spl_,
    g96_n
  );


  buf

  (
    g99_p_spl_,
    g99_p
  );


  buf

  (
    g96_p_spl_,
    g96_p
  );


  buf

  (
    g99_n_spl_,
    g99_n
  );


  buf

  (
    g102_p_spl_,
    g102_p
  );


  buf

  (
    g102_n_spl_,
    g102_n
  );


  buf

  (
    g106_n_spl_,
    g106_n
  );


  buf

  (
    g106_p_spl_,
    g106_p
  );


  buf

  (
    G14_n_spl_,
    G14_n
  );


  buf

  (
    G14_n_spl_0,
    G14_n_spl_
  );


  buf

  (
    G14_n_spl_00,
    G14_n_spl_0
  );


  buf

  (
    G14_n_spl_000,
    G14_n_spl_00
  );


  buf

  (
    G14_n_spl_001,
    G14_n_spl_00
  );


  buf

  (
    G14_n_spl_01,
    G14_n_spl_0
  );


  buf

  (
    G14_n_spl_010,
    G14_n_spl_01
  );


  buf

  (
    G14_n_spl_011,
    G14_n_spl_01
  );


  buf

  (
    G14_n_spl_1,
    G14_n_spl_
  );


  buf

  (
    G14_n_spl_10,
    G14_n_spl_1
  );


  buf

  (
    G14_n_spl_100,
    G14_n_spl_10
  );


  buf

  (
    G14_n_spl_101,
    G14_n_spl_10
  );


  buf

  (
    G14_n_spl_11,
    G14_n_spl_1
  );


  buf

  (
    G14_n_spl_110,
    G14_n_spl_11
  );


  buf

  (
    G14_n_spl_111,
    G14_n_spl_11
  );


  buf

  (
    g108_p_spl_,
    g108_p
  );


  buf

  (
    g111_n_spl_,
    g111_n
  );


  buf

  (
    g108_n_spl_,
    g108_n
  );


  buf

  (
    g111_p_spl_,
    g111_p
  );


  buf

  (
    g117_n_spl_,
    g117_n
  );


  buf

  (
    g117_p_spl_,
    g117_p
  );


  buf

  (
    g116_p_spl_,
    g116_p
  );


  buf

  (
    g119_n_spl_,
    g119_n
  );


  buf

  (
    g116_n_spl_,
    g116_n
  );


  buf

  (
    g119_p_spl_,
    g119_p
  );


  buf

  (
    g122_p_spl_,
    g122_p
  );


  buf

  (
    g122_n_spl_,
    g122_n
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_00,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_000,
    G4_p_spl_00
  );


  buf

  (
    G4_p_spl_0000,
    G4_p_spl_000
  );


  buf

  (
    G4_p_spl_00000,
    G4_p_spl_0000
  );


  buf

  (
    G4_p_spl_00001,
    G4_p_spl_0000
  );


  buf

  (
    G4_p_spl_0001,
    G4_p_spl_000
  );


  buf

  (
    G4_p_spl_00010,
    G4_p_spl_0001
  );


  buf

  (
    G4_p_spl_00011,
    G4_p_spl_0001
  );


  buf

  (
    G4_p_spl_001,
    G4_p_spl_00
  );


  buf

  (
    G4_p_spl_0010,
    G4_p_spl_001
  );


  buf

  (
    G4_p_spl_0011,
    G4_p_spl_001
  );


  buf

  (
    G4_p_spl_01,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_010,
    G4_p_spl_01
  );


  buf

  (
    G4_p_spl_0100,
    G4_p_spl_010
  );


  buf

  (
    G4_p_spl_0101,
    G4_p_spl_010
  );


  buf

  (
    G4_p_spl_011,
    G4_p_spl_01
  );


  buf

  (
    G4_p_spl_0110,
    G4_p_spl_011
  );


  buf

  (
    G4_p_spl_0111,
    G4_p_spl_011
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_10,
    G4_p_spl_1
  );


  buf

  (
    G4_p_spl_100,
    G4_p_spl_10
  );


  buf

  (
    G4_p_spl_1000,
    G4_p_spl_100
  );


  buf

  (
    G4_p_spl_1001,
    G4_p_spl_100
  );


  buf

  (
    G4_p_spl_101,
    G4_p_spl_10
  );


  buf

  (
    G4_p_spl_1010,
    G4_p_spl_101
  );


  buf

  (
    G4_p_spl_1011,
    G4_p_spl_101
  );


  buf

  (
    G4_p_spl_11,
    G4_p_spl_1
  );


  buf

  (
    G4_p_spl_110,
    G4_p_spl_11
  );


  buf

  (
    G4_p_spl_1100,
    G4_p_spl_110
  );


  buf

  (
    G4_p_spl_1101,
    G4_p_spl_110
  );


  buf

  (
    G4_p_spl_111,
    G4_p_spl_11
  );


  buf

  (
    G4_p_spl_1110,
    G4_p_spl_111
  );


  buf

  (
    G4_p_spl_1111,
    G4_p_spl_111
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    G4_n_spl_0,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_00,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_000,
    G4_n_spl_00
  );


  buf

  (
    G4_n_spl_0000,
    G4_n_spl_000
  );


  buf

  (
    G4_n_spl_00000,
    G4_n_spl_0000
  );


  buf

  (
    G4_n_spl_00001,
    G4_n_spl_0000
  );


  buf

  (
    G4_n_spl_0001,
    G4_n_spl_000
  );


  buf

  (
    G4_n_spl_00010,
    G4_n_spl_0001
  );


  buf

  (
    G4_n_spl_00011,
    G4_n_spl_0001
  );


  buf

  (
    G4_n_spl_001,
    G4_n_spl_00
  );


  buf

  (
    G4_n_spl_0010,
    G4_n_spl_001
  );


  buf

  (
    G4_n_spl_0011,
    G4_n_spl_001
  );


  buf

  (
    G4_n_spl_01,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_010,
    G4_n_spl_01
  );


  buf

  (
    G4_n_spl_0100,
    G4_n_spl_010
  );


  buf

  (
    G4_n_spl_0101,
    G4_n_spl_010
  );


  buf

  (
    G4_n_spl_011,
    G4_n_spl_01
  );


  buf

  (
    G4_n_spl_0110,
    G4_n_spl_011
  );


  buf

  (
    G4_n_spl_0111,
    G4_n_spl_011
  );


  buf

  (
    G4_n_spl_1,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_10,
    G4_n_spl_1
  );


  buf

  (
    G4_n_spl_100,
    G4_n_spl_10
  );


  buf

  (
    G4_n_spl_1000,
    G4_n_spl_100
  );


  buf

  (
    G4_n_spl_1001,
    G4_n_spl_100
  );


  buf

  (
    G4_n_spl_101,
    G4_n_spl_10
  );


  buf

  (
    G4_n_spl_1010,
    G4_n_spl_101
  );


  buf

  (
    G4_n_spl_1011,
    G4_n_spl_101
  );


  buf

  (
    G4_n_spl_11,
    G4_n_spl_1
  );


  buf

  (
    G4_n_spl_110,
    G4_n_spl_11
  );


  buf

  (
    G4_n_spl_1100,
    G4_n_spl_110
  );


  buf

  (
    G4_n_spl_1101,
    G4_n_spl_110
  );


  buf

  (
    G4_n_spl_111,
    G4_n_spl_11
  );


  buf

  (
    G4_n_spl_1110,
    G4_n_spl_111
  );


  buf

  (
    G4_n_spl_1111,
    G4_n_spl_111
  );


  buf

  (
    g126_n_spl_,
    g126_n
  );


  buf

  (
    g126_p_spl_,
    g126_p
  );


  buf

  (
    g129_p_spl_,
    g129_p
  );


  buf

  (
    g129_p_spl_0,
    g129_p_spl_
  );


  buf

  (
    g129_p_spl_00,
    g129_p_spl_0
  );


  buf

  (
    g129_p_spl_000,
    g129_p_spl_00
  );


  buf

  (
    g129_p_spl_001,
    g129_p_spl_00
  );


  buf

  (
    g129_p_spl_01,
    g129_p_spl_0
  );


  buf

  (
    g129_p_spl_1,
    g129_p_spl_
  );


  buf

  (
    g129_p_spl_10,
    g129_p_spl_1
  );


  buf

  (
    g129_p_spl_11,
    g129_p_spl_1
  );


  buf

  (
    g130_n_spl_,
    g130_n
  );


  buf

  (
    g130_n_spl_0,
    g130_n_spl_
  );


  buf

  (
    g130_n_spl_00,
    g130_n_spl_0
  );


  buf

  (
    g130_n_spl_01,
    g130_n_spl_0
  );


  buf

  (
    g130_n_spl_1,
    g130_n_spl_
  );


  buf

  (
    g130_n_spl_10,
    g130_n_spl_1
  );


  buf

  (
    g130_n_spl_11,
    g130_n_spl_1
  );


  buf

  (
    g129_n_spl_,
    g129_n
  );


  buf

  (
    g129_n_spl_0,
    g129_n_spl_
  );


  buf

  (
    g129_n_spl_00,
    g129_n_spl_0
  );


  buf

  (
    g129_n_spl_000,
    g129_n_spl_00
  );


  buf

  (
    g129_n_spl_001,
    g129_n_spl_00
  );


  buf

  (
    g129_n_spl_01,
    g129_n_spl_0
  );


  buf

  (
    g129_n_spl_1,
    g129_n_spl_
  );


  buf

  (
    g129_n_spl_10,
    g129_n_spl_1
  );


  buf

  (
    g129_n_spl_11,
    g129_n_spl_1
  );


  buf

  (
    g130_p_spl_,
    g130_p
  );


  buf

  (
    g130_p_spl_0,
    g130_p_spl_
  );


  buf

  (
    g130_p_spl_00,
    g130_p_spl_0
  );


  buf

  (
    g130_p_spl_01,
    g130_p_spl_0
  );


  buf

  (
    g130_p_spl_1,
    g130_p_spl_
  );


  buf

  (
    g130_p_spl_10,
    g130_p_spl_1
  );


  buf

  (
    g130_p_spl_11,
    g130_p_spl_1
  );


  buf

  (
    g131_p_spl_,
    g131_p
  );


  buf

  (
    g131_n_spl_,
    g131_n
  );


  buf

  (
    g133_n_spl_,
    g133_n
  );


  buf

  (
    g133_n_spl_0,
    g133_n_spl_
  );


  buf

  (
    g133_n_spl_1,
    g133_n_spl_
  );


  buf

  (
    g134_n_spl_,
    g134_n
  );


  buf

  (
    g134_n_spl_0,
    g134_n_spl_
  );


  buf

  (
    g133_p_spl_,
    g133_p
  );


  buf

  (
    g133_p_spl_0,
    g133_p_spl_
  );


  buf

  (
    g133_p_spl_1,
    g133_p_spl_
  );


  buf

  (
    g134_p_spl_,
    g134_p
  );


  buf

  (
    g134_p_spl_0,
    g134_p_spl_
  );


  buf

  (
    g137_n_spl_,
    g137_n
  );


  buf

  (
    g137_n_spl_0,
    g137_n_spl_
  );


  buf

  (
    g137_n_spl_00,
    g137_n_spl_0
  );


  buf

  (
    g137_n_spl_000,
    g137_n_spl_00
  );


  buf

  (
    g137_n_spl_01,
    g137_n_spl_0
  );


  buf

  (
    g137_n_spl_1,
    g137_n_spl_
  );


  buf

  (
    g137_n_spl_10,
    g137_n_spl_1
  );


  buf

  (
    g137_n_spl_11,
    g137_n_spl_1
  );


  buf

  (
    g137_p_spl_,
    g137_p
  );


  buf

  (
    g137_p_spl_0,
    g137_p_spl_
  );


  buf

  (
    g137_p_spl_00,
    g137_p_spl_0
  );


  buf

  (
    g137_p_spl_000,
    g137_p_spl_00
  );


  buf

  (
    g137_p_spl_01,
    g137_p_spl_0
  );


  buf

  (
    g137_p_spl_1,
    g137_p_spl_
  );


  buf

  (
    g137_p_spl_10,
    g137_p_spl_1
  );


  buf

  (
    g137_p_spl_11,
    g137_p_spl_1
  );


  buf

  (
    g138_p_spl_,
    g138_p
  );


  buf

  (
    g138_p_spl_0,
    g138_p_spl_
  );


  buf

  (
    g138_p_spl_00,
    g138_p_spl_0
  );


  buf

  (
    g138_p_spl_01,
    g138_p_spl_0
  );


  buf

  (
    g138_p_spl_1,
    g138_p_spl_
  );


  buf

  (
    g138_p_spl_10,
    g138_p_spl_1
  );


  buf

  (
    g138_p_spl_11,
    g138_p_spl_1
  );


  buf

  (
    g138_n_spl_,
    g138_n
  );


  buf

  (
    g138_n_spl_0,
    g138_n_spl_
  );


  buf

  (
    g138_n_spl_00,
    g138_n_spl_0
  );


  buf

  (
    g138_n_spl_01,
    g138_n_spl_0
  );


  buf

  (
    g138_n_spl_1,
    g138_n_spl_
  );


  buf

  (
    g138_n_spl_10,
    g138_n_spl_1
  );


  buf

  (
    g138_n_spl_11,
    g138_n_spl_1
  );


  buf

  (
    G39_p_spl_,
    G39_p
  );


  buf

  (
    G39_p_spl_0,
    G39_p_spl_
  );


  buf

  (
    G39_p_spl_00,
    G39_p_spl_0
  );


  buf

  (
    G39_p_spl_000,
    G39_p_spl_00
  );


  buf

  (
    G39_p_spl_01,
    G39_p_spl_0
  );


  buf

  (
    G39_p_spl_1,
    G39_p_spl_
  );


  buf

  (
    G39_p_spl_10,
    G39_p_spl_1
  );


  buf

  (
    G39_p_spl_11,
    G39_p_spl_1
  );


  buf

  (
    G39_n_spl_,
    G39_n
  );


  buf

  (
    G39_n_spl_0,
    G39_n_spl_
  );


  buf

  (
    G39_n_spl_00,
    G39_n_spl_0
  );


  buf

  (
    G39_n_spl_000,
    G39_n_spl_00
  );


  buf

  (
    G39_n_spl_01,
    G39_n_spl_0
  );


  buf

  (
    G39_n_spl_1,
    G39_n_spl_
  );


  buf

  (
    G39_n_spl_10,
    G39_n_spl_1
  );


  buf

  (
    G39_n_spl_11,
    G39_n_spl_1
  );


  buf

  (
    G5_p_spl_,
    G5_p
  );


  buf

  (
    G5_p_spl_0,
    G5_p_spl_
  );


  buf

  (
    G5_p_spl_00,
    G5_p_spl_0
  );


  buf

  (
    G5_p_spl_01,
    G5_p_spl_0
  );


  buf

  (
    G5_p_spl_1,
    G5_p_spl_
  );


  buf

  (
    G5_n_spl_,
    G5_n
  );


  buf

  (
    G5_n_spl_0,
    G5_n_spl_
  );


  buf

  (
    G5_n_spl_00,
    G5_n_spl_0
  );


  buf

  (
    G5_n_spl_01,
    G5_n_spl_0
  );


  buf

  (
    G5_n_spl_1,
    G5_n_spl_
  );


  buf

  (
    g146_n_spl_,
    g146_n
  );


  buf

  (
    g146_p_spl_,
    g146_p
  );


  buf

  (
    g147_n_spl_,
    g147_n
  );


  buf

  (
    g147_n_spl_0,
    g147_n_spl_
  );


  buf

  (
    g147_n_spl_00,
    g147_n_spl_0
  );


  buf

  (
    g147_n_spl_000,
    g147_n_spl_00
  );


  buf

  (
    g147_n_spl_01,
    g147_n_spl_0
  );


  buf

  (
    g147_n_spl_1,
    g147_n_spl_
  );


  buf

  (
    g147_n_spl_10,
    g147_n_spl_1
  );


  buf

  (
    g147_n_spl_11,
    g147_n_spl_1
  );


  buf

  (
    g147_p_spl_,
    g147_p
  );


  buf

  (
    g147_p_spl_0,
    g147_p_spl_
  );


  buf

  (
    g147_p_spl_00,
    g147_p_spl_0
  );


  buf

  (
    g147_p_spl_000,
    g147_p_spl_00
  );


  buf

  (
    g147_p_spl_01,
    g147_p_spl_0
  );


  buf

  (
    g147_p_spl_1,
    g147_p_spl_
  );


  buf

  (
    g147_p_spl_10,
    g147_p_spl_1
  );


  buf

  (
    g147_p_spl_11,
    g147_p_spl_1
  );


  buf

  (
    G6_n_spl_,
    G6_n
  );


  buf

  (
    G6_n_spl_0,
    G6_n_spl_
  );


  buf

  (
    G6_n_spl_00,
    G6_n_spl_0
  );


  buf

  (
    G6_n_spl_01,
    G6_n_spl_0
  );


  buf

  (
    G6_n_spl_1,
    G6_n_spl_
  );


  buf

  (
    G6_n_spl_10,
    G6_n_spl_1
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G6_p_spl_0,
    G6_p_spl_
  );


  buf

  (
    G6_p_spl_00,
    G6_p_spl_0
  );


  buf

  (
    G6_p_spl_01,
    G6_p_spl_0
  );


  buf

  (
    G6_p_spl_1,
    G6_p_spl_
  );


  buf

  (
    G6_p_spl_10,
    G6_p_spl_1
  );


  buf

  (
    g149_p_spl_,
    g149_p
  );


  buf

  (
    g149_p_spl_0,
    g149_p_spl_
  );


  buf

  (
    g149_n_spl_,
    g149_n
  );


  buf

  (
    g149_n_spl_0,
    g149_n_spl_
  );


  buf

  (
    g148_p_spl_,
    g148_p
  );


  buf

  (
    g148_p_spl_0,
    g148_p_spl_
  );


  buf

  (
    g150_p_spl_,
    g150_p
  );


  buf

  (
    g150_p_spl_0,
    g150_p_spl_
  );


  buf

  (
    g150_p_spl_1,
    g150_p_spl_
  );


  buf

  (
    g148_n_spl_,
    g148_n
  );


  buf

  (
    g148_n_spl_0,
    g148_n_spl_
  );


  buf

  (
    g150_n_spl_,
    g150_n
  );


  buf

  (
    g150_n_spl_0,
    g150_n_spl_
  );


  buf

  (
    g150_n_spl_1,
    g150_n_spl_
  );


  buf

  (
    g153_p_spl_,
    g153_p
  );


  buf

  (
    g153_p_spl_0,
    g153_p_spl_
  );


  buf

  (
    g153_p_spl_00,
    g153_p_spl_0
  );


  buf

  (
    g153_p_spl_01,
    g153_p_spl_0
  );


  buf

  (
    g153_p_spl_1,
    g153_p_spl_
  );


  buf

  (
    g153_p_spl_10,
    g153_p_spl_1
  );


  buf

  (
    g153_p_spl_11,
    g153_p_spl_1
  );


  buf

  (
    g153_n_spl_,
    g153_n
  );


  buf

  (
    g153_n_spl_0,
    g153_n_spl_
  );


  buf

  (
    g153_n_spl_00,
    g153_n_spl_0
  );


  buf

  (
    g153_n_spl_01,
    g153_n_spl_0
  );


  buf

  (
    g153_n_spl_1,
    g153_n_spl_
  );


  buf

  (
    g153_n_spl_10,
    g153_n_spl_1
  );


  buf

  (
    g153_n_spl_11,
    g153_n_spl_1
  );


  buf

  (
    G41_n_spl_,
    G41_n
  );


  buf

  (
    G41_n_spl_0,
    G41_n_spl_
  );


  buf

  (
    G41_n_spl_00,
    G41_n_spl_0
  );


  buf

  (
    G41_n_spl_01,
    G41_n_spl_0
  );


  buf

  (
    G41_n_spl_1,
    G41_n_spl_
  );


  buf

  (
    G41_n_spl_10,
    G41_n_spl_1
  );


  buf

  (
    G41_p_spl_,
    G41_p
  );


  buf

  (
    G41_p_spl_0,
    G41_p_spl_
  );


  buf

  (
    G41_p_spl_00,
    G41_p_spl_0
  );


  buf

  (
    G41_p_spl_01,
    G41_p_spl_0
  );


  buf

  (
    G41_p_spl_1,
    G41_p_spl_
  );


  buf

  (
    G41_p_spl_10,
    G41_p_spl_1
  );


  buf

  (
    g151_n_spl_,
    g151_n
  );


  buf

  (
    g151_n_spl_0,
    g151_n_spl_
  );


  buf

  (
    g151_p_spl_,
    g151_p
  );


  buf

  (
    g151_p_spl_0,
    g151_p_spl_
  );


  buf

  (
    G25_n_spl_,
    G25_n
  );


  buf

  (
    G26_n_spl_,
    G26_n
  );


  buf

  (
    G26_n_spl_0,
    G26_n_spl_
  );


  buf

  (
    G25_p_spl_,
    G25_p
  );


  buf

  (
    G26_p_spl_,
    G26_p
  );


  buf

  (
    G26_p_spl_0,
    G26_p_spl_
  );


  buf

  (
    g161_p_spl_,
    g161_p
  );


  buf

  (
    g161_p_spl_0,
    g161_p_spl_
  );


  buf

  (
    g161_p_spl_1,
    g161_p_spl_
  );


  buf

  (
    g162_n_spl_,
    g162_n
  );


  buf

  (
    g162_n_spl_0,
    g162_n_spl_
  );


  buf

  (
    g162_n_spl_00,
    g162_n_spl_0
  );


  buf

  (
    g162_n_spl_000,
    g162_n_spl_00
  );


  buf

  (
    g162_n_spl_01,
    g162_n_spl_0
  );


  buf

  (
    g162_n_spl_1,
    g162_n_spl_
  );


  buf

  (
    g162_n_spl_10,
    g162_n_spl_1
  );


  buf

  (
    g162_n_spl_11,
    g162_n_spl_1
  );


  buf

  (
    g161_n_spl_,
    g161_n
  );


  buf

  (
    g161_n_spl_0,
    g161_n_spl_
  );


  buf

  (
    g161_n_spl_1,
    g161_n_spl_
  );


  buf

  (
    g162_p_spl_,
    g162_p
  );


  buf

  (
    g162_p_spl_0,
    g162_p_spl_
  );


  buf

  (
    g162_p_spl_00,
    g162_p_spl_0
  );


  buf

  (
    g162_p_spl_000,
    g162_p_spl_00
  );


  buf

  (
    g162_p_spl_01,
    g162_p_spl_0
  );


  buf

  (
    g162_p_spl_1,
    g162_p_spl_
  );


  buf

  (
    g162_p_spl_10,
    g162_p_spl_1
  );


  buf

  (
    g162_p_spl_11,
    g162_p_spl_1
  );


  buf

  (
    g145_p_spl_,
    g145_p
  );


  buf

  (
    g145_p_spl_0,
    g145_p_spl_
  );


  buf

  (
    g145_n_spl_,
    g145_n
  );


  buf

  (
    g145_n_spl_0,
    g145_n_spl_
  );


  buf

  (
    G23_n_spl_,
    G23_n
  );


  buf

  (
    G24_n_spl_,
    G24_n
  );


  buf

  (
    G24_n_spl_0,
    G24_n_spl_
  );


  buf

  (
    G24_n_spl_1,
    G24_n_spl_
  );


  buf

  (
    G23_p_spl_,
    G23_p
  );


  buf

  (
    G24_p_spl_,
    G24_p
  );


  buf

  (
    G24_p_spl_0,
    G24_p_spl_
  );


  buf

  (
    G24_p_spl_1,
    G24_p_spl_
  );


  buf

  (
    g165_n_spl_,
    g165_n
  );


  buf

  (
    g165_n_spl_0,
    g165_n_spl_
  );


  buf

  (
    g165_n_spl_00,
    g165_n_spl_0
  );


  buf

  (
    g165_n_spl_01,
    g165_n_spl_0
  );


  buf

  (
    g165_n_spl_1,
    g165_n_spl_
  );


  buf

  (
    g165_n_spl_10,
    g165_n_spl_1
  );


  buf

  (
    g165_n_spl_11,
    g165_n_spl_1
  );


  buf

  (
    g165_p_spl_,
    g165_p
  );


  buf

  (
    g165_p_spl_0,
    g165_p_spl_
  );


  buf

  (
    g165_p_spl_00,
    g165_p_spl_0
  );


  buf

  (
    g165_p_spl_01,
    g165_p_spl_0
  );


  buf

  (
    g165_p_spl_1,
    g165_p_spl_
  );


  buf

  (
    g165_p_spl_10,
    g165_p_spl_1
  );


  buf

  (
    g165_p_spl_11,
    g165_p_spl_1
  );


  buf

  (
    g167_n_spl_,
    g167_n
  );


  buf

  (
    g167_n_spl_0,
    g167_n_spl_
  );


  buf

  (
    g167_p_spl_,
    g167_p
  );


  buf

  (
    g167_p_spl_0,
    g167_p_spl_
  );


  buf

  (
    g169_n_spl_,
    g169_n
  );


  buf

  (
    g169_p_spl_,
    g169_p
  );


  buf

  (
    G40_n_spl_,
    G40_n
  );


  buf

  (
    G40_n_spl_0,
    G40_n_spl_
  );


  buf

  (
    G40_n_spl_00,
    G40_n_spl_0
  );


  buf

  (
    G40_n_spl_01,
    G40_n_spl_0
  );


  buf

  (
    G40_n_spl_1,
    G40_n_spl_
  );


  buf

  (
    G40_n_spl_10,
    G40_n_spl_1
  );


  buf

  (
    G40_p_spl_,
    G40_p
  );


  buf

  (
    G40_p_spl_0,
    G40_p_spl_
  );


  buf

  (
    G40_p_spl_00,
    G40_p_spl_0
  );


  buf

  (
    G40_p_spl_01,
    G40_p_spl_0
  );


  buf

  (
    G40_p_spl_1,
    G40_p_spl_
  );


  buf

  (
    G40_p_spl_10,
    G40_p_spl_1
  );


  buf

  (
    g186_p_spl_,
    g186_p
  );


  buf

  (
    g186_p_spl_0,
    g186_p_spl_
  );


  buf

  (
    g186_p_spl_1,
    g186_p_spl_
  );


  buf

  (
    g186_n_spl_,
    g186_n
  );


  buf

  (
    g186_n_spl_0,
    g186_n_spl_
  );


  buf

  (
    g186_n_spl_1,
    g186_n_spl_
  );


  buf

  (
    g177_p_spl_,
    g177_p
  );


  buf

  (
    g177_p_spl_0,
    g177_p_spl_
  );


  buf

  (
    g177_n_spl_,
    g177_n
  );


  buf

  (
    g177_n_spl_0,
    g177_n_spl_
  );


  buf

  (
    g190_n_spl_,
    g190_n
  );


  buf

  (
    g190_n_spl_0,
    g190_n_spl_
  );


  buf

  (
    g190_p_spl_,
    g190_p
  );


  buf

  (
    g190_p_spl_0,
    g190_p_spl_
  );


  buf

  (
    g196_n_spl_,
    g196_n
  );


  buf

  (
    g196_p_spl_,
    g196_p
  );


  buf

  (
    g212_p_spl_,
    g212_p
  );


  buf

  (
    g212_p_spl_0,
    g212_p_spl_
  );


  buf

  (
    g212_p_spl_1,
    g212_p_spl_
  );


  buf

  (
    g212_n_spl_,
    g212_n
  );


  buf

  (
    g212_n_spl_0,
    g212_n_spl_
  );


  buf

  (
    g212_n_spl_1,
    g212_n_spl_
  );


  buf

  (
    g202_p_spl_,
    g202_p
  );


  buf

  (
    g202_p_spl_0,
    g202_p_spl_
  );


  buf

  (
    g202_n_spl_,
    g202_n
  );


  buf

  (
    g202_n_spl_0,
    g202_n_spl_
  );


  buf

  (
    g216_n_spl_,
    g216_n
  );


  buf

  (
    g216_p_spl_,
    g216_p
  );


  buf

  (
    g223_n_spl_,
    g223_n
  );


  buf

  (
    g238_p_spl_,
    g238_p
  );


  buf

  (
    g238_p_spl_0,
    g238_p_spl_
  );


  buf

  (
    g238_p_spl_1,
    g238_p_spl_
  );


  buf

  (
    g238_n_spl_,
    g238_n
  );


  buf

  (
    g238_n_spl_0,
    g238_n_spl_
  );


  buf

  (
    g238_n_spl_1,
    g238_n_spl_
  );


  buf

  (
    g229_p_spl_,
    g229_p
  );


  buf

  (
    g229_p_spl_0,
    g229_p_spl_
  );


  buf

  (
    g229_n_spl_,
    g229_n
  );


  buf

  (
    g229_n_spl_0,
    g229_n_spl_
  );


  buf

  (
    g242_n_spl_,
    g242_n
  );


  buf

  (
    g242_n_spl_0,
    g242_n_spl_
  );


  buf

  (
    g242_p_spl_,
    g242_p
  );


  buf

  (
    g242_p_spl_0,
    g242_p_spl_
  );


  buf

  (
    g217_p_spl_,
    g217_p
  );


  buf

  (
    g217_p_spl_0,
    g217_p_spl_
  );


  buf

  (
    g217_p_spl_1,
    g217_p_spl_
  );


  buf

  (
    g243_p_spl_,
    g243_p
  );


  buf

  (
    g243_p_spl_0,
    g243_p_spl_
  );


  buf

  (
    g217_n_spl_,
    g217_n
  );


  buf

  (
    g217_n_spl_0,
    g217_n_spl_
  );


  buf

  (
    g217_n_spl_1,
    g217_n_spl_
  );


  buf

  (
    g243_n_spl_,
    g243_n
  );


  buf

  (
    g243_n_spl_0,
    g243_n_spl_
  );


  buf

  (
    g191_p_spl_,
    g191_p
  );


  buf

  (
    g191_p_spl_0,
    g191_p_spl_
  );


  buf

  (
    g244_p_spl_,
    g244_p
  );


  buf

  (
    g191_n_spl_,
    g191_n
  );


  buf

  (
    g191_n_spl_0,
    g191_n_spl_
  );


  buf

  (
    g244_n_spl_,
    g244_n
  );


  buf

  (
    g168_p_spl_,
    g168_p
  );


  buf

  (
    g168_p_spl_0,
    g168_p_spl_
  );


  buf

  (
    g245_p_spl_,
    g245_p
  );


  buf

  (
    g168_n_spl_,
    g168_n
  );


  buf

  (
    g168_n_spl_0,
    g168_n_spl_
  );


  buf

  (
    g245_n_spl_,
    g245_n
  );


  buf

  (
    g248_n_spl_,
    g248_n
  );


  buf

  (
    g248_n_spl_0,
    g248_n_spl_
  );


  buf

  (
    g248_n_spl_1,
    g248_n_spl_
  );


  buf

  (
    g248_p_spl_,
    g248_p
  );


  buf

  (
    g248_p_spl_0,
    g248_p_spl_
  );


  buf

  (
    g248_p_spl_1,
    g248_p_spl_
  );


  buf

  (
    g259_p_spl_,
    g259_p
  );


  buf

  (
    g259_p_spl_0,
    g259_p_spl_
  );


  buf

  (
    g259_p_spl_00,
    g259_p_spl_0
  );


  buf

  (
    g259_p_spl_1,
    g259_p_spl_
  );


  buf

  (
    g259_n_spl_,
    g259_n
  );


  buf

  (
    g259_n_spl_0,
    g259_n_spl_
  );


  buf

  (
    g259_n_spl_00,
    g259_n_spl_0
  );


  buf

  (
    g259_n_spl_1,
    g259_n_spl_
  );


  buf

  (
    g260_n_spl_,
    g260_n
  );


  buf

  (
    g260_n_spl_0,
    g260_n_spl_
  );


  buf

  (
    g260_n_spl_1,
    g260_n_spl_
  );


  buf

  (
    g260_p_spl_,
    g260_p
  );


  buf

  (
    g260_p_spl_0,
    g260_p_spl_
  );


  buf

  (
    g260_p_spl_1,
    g260_p_spl_
  );


  buf

  (
    g269_p_spl_,
    g269_p
  );


  buf

  (
    g269_n_spl_,
    g269_n
  );


  buf

  (
    g257_p_spl_,
    g257_p
  );


  buf

  (
    g257_p_spl_0,
    g257_p_spl_
  );


  buf

  (
    g257_n_spl_,
    g257_n
  );


  buf

  (
    g257_n_spl_0,
    g257_n_spl_
  );


  buf

  (
    g273_n_spl_,
    g273_n
  );


  buf

  (
    g273_n_spl_0,
    g273_n_spl_
  );


  buf

  (
    g273_p_spl_,
    g273_p
  );


  buf

  (
    g273_p_spl_0,
    g273_p_spl_
  );


  buf

  (
    g291_p_spl_,
    g291_p
  );


  buf

  (
    g291_n_spl_,
    g291_n
  );


  buf

  (
    g282_p_spl_,
    g282_p
  );


  buf

  (
    g282_p_spl_0,
    g282_p_spl_
  );


  buf

  (
    g282_n_spl_,
    g282_n
  );


  buf

  (
    g282_n_spl_0,
    g282_n_spl_
  );


  buf

  (
    g295_n_spl_,
    g295_n
  );


  buf

  (
    g295_n_spl_0,
    g295_n_spl_
  );


  buf

  (
    g295_p_spl_,
    g295_p
  );


  buf

  (
    g295_p_spl_0,
    g295_p_spl_
  );


  buf

  (
    G21_p_spl_,
    G21_p
  );


  buf

  (
    G21_p_spl_0,
    G21_p_spl_
  );


  buf

  (
    G21_p_spl_00,
    G21_p_spl_0
  );


  buf

  (
    G21_p_spl_01,
    G21_p_spl_0
  );


  buf

  (
    G21_p_spl_1,
    G21_p_spl_
  );


  buf

  (
    G21_p_spl_10,
    G21_p_spl_1
  );


  buf

  (
    G21_p_spl_11,
    G21_p_spl_1
  );


  buf

  (
    G21_n_spl_,
    G21_n
  );


  buf

  (
    G21_n_spl_0,
    G21_n_spl_
  );


  buf

  (
    G21_n_spl_00,
    G21_n_spl_0
  );


  buf

  (
    G21_n_spl_01,
    G21_n_spl_0
  );


  buf

  (
    G21_n_spl_1,
    G21_n_spl_
  );


  buf

  (
    G21_n_spl_10,
    G21_n_spl_1
  );


  buf

  (
    G21_n_spl_11,
    G21_n_spl_1
  );


  buf

  (
    G29_n_spl_,
    G29_n
  );


  buf

  (
    G29_p_spl_,
    G29_p
  );


  buf

  (
    g315_p_spl_,
    g315_p
  );


  buf

  (
    g315_n_spl_,
    g315_n
  );


  buf

  (
    g306_p_spl_,
    g306_p
  );


  buf

  (
    g306_p_spl_0,
    g306_p_spl_
  );


  buf

  (
    g306_n_spl_,
    g306_n
  );


  buf

  (
    g306_n_spl_0,
    g306_n_spl_
  );


  buf

  (
    g319_n_spl_,
    g319_n
  );


  buf

  (
    g319_p_spl_,
    g319_p
  );


  buf

  (
    g326_n_spl_,
    g326_n
  );


  buf

  (
    G22_p_spl_,
    G22_p
  );


  buf

  (
    G22_p_spl_0,
    G22_p_spl_
  );


  buf

  (
    G22_p_spl_00,
    G22_p_spl_0
  );


  buf

  (
    G22_p_spl_01,
    G22_p_spl_0
  );


  buf

  (
    G22_p_spl_1,
    G22_p_spl_
  );


  buf

  (
    G22_p_spl_10,
    G22_p_spl_1
  );


  buf

  (
    G22_p_spl_11,
    G22_p_spl_1
  );


  buf

  (
    G22_n_spl_,
    G22_n
  );


  buf

  (
    G22_n_spl_0,
    G22_n_spl_
  );


  buf

  (
    G22_n_spl_00,
    G22_n_spl_0
  );


  buf

  (
    G22_n_spl_01,
    G22_n_spl_0
  );


  buf

  (
    G22_n_spl_1,
    G22_n_spl_
  );


  buf

  (
    G22_n_spl_10,
    G22_n_spl_1
  );


  buf

  (
    G22_n_spl_11,
    G22_n_spl_1
  );


  buf

  (
    g341_p_spl_,
    g341_p
  );


  buf

  (
    g341_n_spl_,
    g341_n
  );


  buf

  (
    g332_p_spl_,
    g332_p
  );


  buf

  (
    g332_p_spl_0,
    g332_p_spl_
  );


  buf

  (
    g332_n_spl_,
    g332_n
  );


  buf

  (
    g332_n_spl_0,
    g332_n_spl_
  );


  buf

  (
    g345_n_spl_,
    g345_n
  );


  buf

  (
    g345_n_spl_0,
    g345_n_spl_
  );


  buf

  (
    g345_p_spl_,
    g345_p
  );


  buf

  (
    g345_p_spl_0,
    g345_p_spl_
  );


  buf

  (
    g320_p_spl_,
    g320_p
  );


  buf

  (
    g320_p_spl_0,
    g320_p_spl_
  );


  buf

  (
    g320_p_spl_1,
    g320_p_spl_
  );


  buf

  (
    g346_p_spl_,
    g346_p
  );


  buf

  (
    g346_p_spl_0,
    g346_p_spl_
  );


  buf

  (
    g320_n_spl_,
    g320_n
  );


  buf

  (
    g320_n_spl_0,
    g320_n_spl_
  );


  buf

  (
    g320_n_spl_1,
    g320_n_spl_
  );


  buf

  (
    g346_n_spl_,
    g346_n
  );


  buf

  (
    g346_n_spl_0,
    g346_n_spl_
  );


  buf

  (
    g296_p_spl_,
    g296_p
  );


  buf

  (
    g296_p_spl_0,
    g296_p_spl_
  );


  buf

  (
    g347_p_spl_,
    g347_p
  );


  buf

  (
    g296_n_spl_,
    g296_n
  );


  buf

  (
    g296_n_spl_0,
    g296_n_spl_
  );


  buf

  (
    g347_n_spl_,
    g347_n
  );


  buf

  (
    g274_p_spl_,
    g274_p
  );


  buf

  (
    g274_p_spl_0,
    g274_p_spl_
  );


  buf

  (
    g348_p_spl_,
    g348_p
  );


  buf

  (
    g274_n_spl_,
    g274_n
  );


  buf

  (
    g274_n_spl_0,
    g274_n_spl_
  );


  buf

  (
    g348_n_spl_,
    g348_n
  );


  buf

  (
    g246_p_spl_,
    g246_p
  );


  buf

  (
    g349_p_spl_,
    g349_p
  );


  buf

  (
    g349_p_spl_0,
    g349_p_spl_
  );


  buf

  (
    g349_p_spl_1,
    g349_p_spl_
  );


  buf

  (
    g356_n_spl_,
    g356_n
  );


  buf

  (
    g363_n_spl_,
    g363_n
  );


  buf

  (
    G27_p_spl_,
    G27_p
  );


  buf

  (
    G27_p_spl_0,
    G27_p_spl_
  );


  buf

  (
    g79_p_spl_,
    g79_p
  );


  buf

  (
    g79_p_spl_0,
    g79_p_spl_
  );


  buf

  (
    G27_n_spl_,
    G27_n
  );


  buf

  (
    G48_p_spl_,
    G48_p
  );


  buf

  (
    g365_p_spl_,
    g365_p
  );


  buf

  (
    g365_p_spl_0,
    g365_p_spl_
  );


  buf

  (
    g365_p_spl_1,
    g365_p_spl_
  );


  buf

  (
    G48_n_spl_,
    G48_n
  );


  buf

  (
    g365_n_spl_,
    g365_n
  );


  buf

  (
    g365_n_spl_0,
    g365_n_spl_
  );


  buf

  (
    g365_n_spl_1,
    g365_n_spl_
  );


  buf

  (
    g366_p_spl_,
    g366_p
  );


  buf

  (
    g366_p_spl_0,
    g366_p_spl_
  );


  buf

  (
    g366_p_spl_00,
    g366_p_spl_0
  );


  buf

  (
    g366_p_spl_000,
    g366_p_spl_00
  );


  buf

  (
    g366_p_spl_001,
    g366_p_spl_00
  );


  buf

  (
    g366_p_spl_01,
    g366_p_spl_0
  );


  buf

  (
    g366_p_spl_010,
    g366_p_spl_01
  );


  buf

  (
    g366_p_spl_011,
    g366_p_spl_01
  );


  buf

  (
    g366_p_spl_1,
    g366_p_spl_
  );


  buf

  (
    g366_p_spl_10,
    g366_p_spl_1
  );


  buf

  (
    g366_p_spl_100,
    g366_p_spl_10
  );


  buf

  (
    g366_p_spl_101,
    g366_p_spl_10
  );


  buf

  (
    g366_p_spl_11,
    g366_p_spl_1
  );


  buf

  (
    g366_n_spl_,
    g366_n
  );


  buf

  (
    g366_n_spl_0,
    g366_n_spl_
  );


  buf

  (
    g366_n_spl_00,
    g366_n_spl_0
  );


  buf

  (
    g366_n_spl_000,
    g366_n_spl_00
  );


  buf

  (
    g366_n_spl_001,
    g366_n_spl_00
  );


  buf

  (
    g366_n_spl_01,
    g366_n_spl_0
  );


  buf

  (
    g366_n_spl_010,
    g366_n_spl_01
  );


  buf

  (
    g366_n_spl_011,
    g366_n_spl_01
  );


  buf

  (
    g366_n_spl_1,
    g366_n_spl_
  );


  buf

  (
    g366_n_spl_10,
    g366_n_spl_1
  );


  buf

  (
    g366_n_spl_100,
    g366_n_spl_10
  );


  buf

  (
    g366_n_spl_101,
    g366_n_spl_10
  );


  buf

  (
    g366_n_spl_11,
    g366_n_spl_1
  );


  buf

  (
    g367_n_spl_,
    g367_n
  );


  buf

  (
    g367_p_spl_,
    g367_p
  );


  buf

  (
    g371_n_spl_,
    g371_n
  );


  buf

  (
    g371_p_spl_,
    g371_p
  );


  buf

  (
    G47_p_spl_,
    G47_p
  );


  buf

  (
    G47_p_spl_0,
    G47_p_spl_
  );


  buf

  (
    G47_p_spl_00,
    G47_p_spl_0
  );


  buf

  (
    G47_p_spl_01,
    G47_p_spl_0
  );


  buf

  (
    G47_p_spl_1,
    G47_p_spl_
  );


  buf

  (
    G47_p_spl_10,
    G47_p_spl_1
  );


  buf

  (
    g374_p_spl_,
    g374_p
  );


  buf

  (
    g374_p_spl_0,
    g374_p_spl_
  );


  buf

  (
    g374_p_spl_1,
    g374_p_spl_
  );


  buf

  (
    G47_n_spl_,
    G47_n
  );


  buf

  (
    G47_n_spl_0,
    G47_n_spl_
  );


  buf

  (
    G47_n_spl_00,
    G47_n_spl_0
  );


  buf

  (
    G47_n_spl_01,
    G47_n_spl_0
  );


  buf

  (
    G47_n_spl_1,
    G47_n_spl_
  );


  buf

  (
    G47_n_spl_10,
    G47_n_spl_1
  );


  buf

  (
    g374_n_spl_,
    g374_n
  );


  buf

  (
    g374_n_spl_0,
    g374_n_spl_
  );


  buf

  (
    g374_n_spl_1,
    g374_n_spl_
  );


  buf

  (
    g370_n_spl_,
    g370_n
  );


  buf

  (
    g370_n_spl_0,
    g370_n_spl_
  );


  buf

  (
    g370_n_spl_1,
    g370_n_spl_
  );


  buf

  (
    g370_p_spl_,
    g370_p
  );


  buf

  (
    g370_p_spl_0,
    g370_p_spl_
  );


  buf

  (
    g370_p_spl_1,
    g370_p_spl_
  );


  buf

  (
    g76_p_spl_,
    g76_p
  );


  buf

  (
    g377_n_spl_,
    g377_n
  );


  buf

  (
    g377_n_spl_0,
    g377_n_spl_
  );


  buf

  (
    g377_n_spl_00,
    g377_n_spl_0
  );


  buf

  (
    g377_n_spl_01,
    g377_n_spl_0
  );


  buf

  (
    g377_n_spl_1,
    g377_n_spl_
  );


  buf

  (
    g377_n_spl_10,
    g377_n_spl_1
  );


  buf

  (
    g377_n_spl_11,
    g377_n_spl_1
  );


  buf

  (
    g379_p_spl_,
    g379_p
  );


  buf

  (
    g379_p_spl_0,
    g379_p_spl_
  );


  buf

  (
    g379_p_spl_00,
    g379_p_spl_0
  );


  buf

  (
    g379_p_spl_01,
    g379_p_spl_0
  );


  buf

  (
    g379_p_spl_1,
    g379_p_spl_
  );


  buf

  (
    g379_p_spl_10,
    g379_p_spl_1
  );


  buf

  (
    g382_p_spl_,
    g382_p
  );


  buf

  (
    g382_n_spl_,
    g382_n
  );


  buf

  (
    g377_p_spl_,
    g377_p
  );


  buf

  (
    g377_p_spl_0,
    g377_p_spl_
  );


  buf

  (
    g377_p_spl_00,
    g377_p_spl_0
  );


  buf

  (
    g377_p_spl_01,
    g377_p_spl_0
  );


  buf

  (
    g377_p_spl_1,
    g377_p_spl_
  );


  buf

  (
    g377_p_spl_10,
    g377_p_spl_1
  );


  buf

  (
    g384_p_spl_,
    g384_p
  );


  buf

  (
    g384_p_spl_0,
    g384_p_spl_
  );


  buf

  (
    g384_p_spl_00,
    g384_p_spl_0
  );


  buf

  (
    g384_p_spl_01,
    g384_p_spl_0
  );


  buf

  (
    g384_p_spl_1,
    g384_p_spl_
  );


  buf

  (
    g384_p_spl_10,
    g384_p_spl_1
  );


  buf

  (
    g384_n_spl_,
    g384_n
  );


  buf

  (
    g384_n_spl_0,
    g384_n_spl_
  );


  buf

  (
    g384_n_spl_00,
    g384_n_spl_0
  );


  buf

  (
    g384_n_spl_01,
    g384_n_spl_0
  );


  buf

  (
    g384_n_spl_1,
    g384_n_spl_
  );


  buf

  (
    g384_n_spl_10,
    g384_n_spl_1
  );


  buf

  (
    g387_n_spl_,
    g387_n
  );


  buf

  (
    g387_n_spl_0,
    g387_n_spl_
  );


  buf

  (
    g387_p_spl_,
    g387_p
  );


  buf

  (
    g387_p_spl_0,
    g387_p_spl_
  );


  buf

  (
    g385_n_spl_,
    g385_n
  );


  buf

  (
    g385_n_spl_0,
    g385_n_spl_
  );


  buf

  (
    g385_n_spl_00,
    g385_n_spl_0
  );


  buf

  (
    g385_n_spl_000,
    g385_n_spl_00
  );


  buf

  (
    g385_n_spl_001,
    g385_n_spl_00
  );


  buf

  (
    g385_n_spl_01,
    g385_n_spl_0
  );


  buf

  (
    g385_n_spl_1,
    g385_n_spl_
  );


  buf

  (
    g385_n_spl_10,
    g385_n_spl_1
  );


  buf

  (
    g385_n_spl_11,
    g385_n_spl_1
  );


  buf

  (
    g385_p_spl_,
    g385_p
  );


  buf

  (
    g385_p_spl_0,
    g385_p_spl_
  );


  buf

  (
    g385_p_spl_00,
    g385_p_spl_0
  );


  buf

  (
    g385_p_spl_000,
    g385_p_spl_00
  );


  buf

  (
    g385_p_spl_001,
    g385_p_spl_00
  );


  buf

  (
    g385_p_spl_01,
    g385_p_spl_0
  );


  buf

  (
    g385_p_spl_1,
    g385_p_spl_
  );


  buf

  (
    g385_p_spl_10,
    g385_p_spl_1
  );


  buf

  (
    g385_p_spl_11,
    g385_p_spl_1
  );


  buf

  (
    g390_p_spl_,
    g390_p
  );


  buf

  (
    g390_p_spl_0,
    g390_p_spl_
  );


  buf

  (
    g390_p_spl_1,
    g390_p_spl_
  );


  buf

  (
    g390_n_spl_,
    g390_n
  );


  buf

  (
    g390_n_spl_0,
    g390_n_spl_
  );


  buf

  (
    g390_n_spl_1,
    g390_n_spl_
  );


  buf

  (
    g394_n_spl_,
    g394_n
  );


  buf

  (
    g394_n_spl_0,
    g394_n_spl_
  );


  buf

  (
    g394_n_spl_00,
    g394_n_spl_0
  );


  buf

  (
    g394_n_spl_01,
    g394_n_spl_0
  );


  buf

  (
    g394_n_spl_1,
    g394_n_spl_
  );


  buf

  (
    g394_p_spl_,
    g394_p
  );


  buf

  (
    g394_p_spl_0,
    g394_p_spl_
  );


  buf

  (
    g394_p_spl_00,
    g394_p_spl_0
  );


  buf

  (
    g394_p_spl_01,
    g394_p_spl_0
  );


  buf

  (
    g394_p_spl_1,
    g394_p_spl_
  );


  buf

  (
    g55_n_spl_,
    g55_n
  );


  buf

  (
    g393_p_spl_,
    g393_p
  );


  buf

  (
    g393_p_spl_0,
    g393_p_spl_
  );


  buf

  (
    g393_p_spl_00,
    g393_p_spl_0
  );


  buf

  (
    g393_p_spl_000,
    g393_p_spl_00
  );


  buf

  (
    g393_p_spl_001,
    g393_p_spl_00
  );


  buf

  (
    g393_p_spl_01,
    g393_p_spl_0
  );


  buf

  (
    g393_p_spl_010,
    g393_p_spl_01
  );


  buf

  (
    g393_p_spl_011,
    g393_p_spl_01
  );


  buf

  (
    g393_p_spl_1,
    g393_p_spl_
  );


  buf

  (
    g393_p_spl_10,
    g393_p_spl_1
  );


  buf

  (
    g393_p_spl_100,
    g393_p_spl_10
  );


  buf

  (
    g393_p_spl_101,
    g393_p_spl_10
  );


  buf

  (
    g393_p_spl_11,
    g393_p_spl_1
  );


  buf

  (
    g393_p_spl_110,
    g393_p_spl_11
  );


  buf

  (
    g393_p_spl_111,
    g393_p_spl_11
  );


  buf

  (
    g393_n_spl_,
    g393_n
  );


  buf

  (
    g393_n_spl_0,
    g393_n_spl_
  );


  buf

  (
    g393_n_spl_00,
    g393_n_spl_0
  );


  buf

  (
    g393_n_spl_000,
    g393_n_spl_00
  );


  buf

  (
    g393_n_spl_001,
    g393_n_spl_00
  );


  buf

  (
    g393_n_spl_01,
    g393_n_spl_0
  );


  buf

  (
    g393_n_spl_010,
    g393_n_spl_01
  );


  buf

  (
    g393_n_spl_011,
    g393_n_spl_01
  );


  buf

  (
    g393_n_spl_1,
    g393_n_spl_
  );


  buf

  (
    g393_n_spl_10,
    g393_n_spl_1
  );


  buf

  (
    g393_n_spl_100,
    g393_n_spl_10
  );


  buf

  (
    g393_n_spl_101,
    g393_n_spl_10
  );


  buf

  (
    g393_n_spl_11,
    g393_n_spl_1
  );


  buf

  (
    g393_n_spl_110,
    g393_n_spl_11
  );


  buf

  (
    g393_n_spl_111,
    g393_n_spl_11
  );


  buf

  (
    g404_n_spl_,
    g404_n
  );


  buf

  (
    g404_n_spl_0,
    g404_n_spl_
  );


  buf

  (
    g404_p_spl_,
    g404_p
  );


  buf

  (
    g404_p_spl_0,
    g404_p_spl_
  );


  buf

  (
    g403_n_spl_,
    g403_n
  );


  buf

  (
    g403_n_spl_0,
    g403_n_spl_
  );


  buf

  (
    g403_n_spl_1,
    g403_n_spl_
  );


  buf

  (
    g405_p_spl_,
    g405_p
  );


  buf

  (
    g403_p_spl_,
    g403_p
  );


  buf

  (
    g403_p_spl_0,
    g403_p_spl_
  );


  buf

  (
    g403_p_spl_1,
    g403_p_spl_
  );


  buf

  (
    g405_n_spl_,
    g405_n
  );


  buf

  (
    G45_p_spl_,
    G45_p
  );


  buf

  (
    g406_n_spl_,
    g406_n
  );


  buf

  (
    g406_n_spl_0,
    g406_n_spl_
  );


  buf

  (
    g406_n_spl_00,
    g406_n_spl_0
  );


  buf

  (
    g406_n_spl_000,
    g406_n_spl_00
  );


  buf

  (
    g406_n_spl_0000,
    g406_n_spl_000
  );


  buf

  (
    g406_n_spl_001,
    g406_n_spl_00
  );


  buf

  (
    g406_n_spl_01,
    g406_n_spl_0
  );


  buf

  (
    g406_n_spl_010,
    g406_n_spl_01
  );


  buf

  (
    g406_n_spl_011,
    g406_n_spl_01
  );


  buf

  (
    g406_n_spl_1,
    g406_n_spl_
  );


  buf

  (
    g406_n_spl_10,
    g406_n_spl_1
  );


  buf

  (
    g406_n_spl_100,
    g406_n_spl_10
  );


  buf

  (
    g406_n_spl_101,
    g406_n_spl_10
  );


  buf

  (
    g406_n_spl_11,
    g406_n_spl_1
  );


  buf

  (
    g406_n_spl_110,
    g406_n_spl_11
  );


  buf

  (
    g406_n_spl_111,
    g406_n_spl_11
  );


  buf

  (
    G45_n_spl_,
    G45_n
  );


  buf

  (
    g406_p_spl_,
    g406_p
  );


  buf

  (
    g406_p_spl_0,
    g406_p_spl_
  );


  buf

  (
    g406_p_spl_00,
    g406_p_spl_0
  );


  buf

  (
    g406_p_spl_000,
    g406_p_spl_00
  );


  buf

  (
    g406_p_spl_0000,
    g406_p_spl_000
  );


  buf

  (
    g406_p_spl_001,
    g406_p_spl_00
  );


  buf

  (
    g406_p_spl_01,
    g406_p_spl_0
  );


  buf

  (
    g406_p_spl_010,
    g406_p_spl_01
  );


  buf

  (
    g406_p_spl_011,
    g406_p_spl_01
  );


  buf

  (
    g406_p_spl_1,
    g406_p_spl_
  );


  buf

  (
    g406_p_spl_10,
    g406_p_spl_1
  );


  buf

  (
    g406_p_spl_100,
    g406_p_spl_10
  );


  buf

  (
    g406_p_spl_101,
    g406_p_spl_10
  );


  buf

  (
    g406_p_spl_11,
    g406_p_spl_1
  );


  buf

  (
    g406_p_spl_110,
    g406_p_spl_11
  );


  buf

  (
    g406_p_spl_111,
    g406_p_spl_11
  );


  buf

  (
    g408_p_spl_,
    g408_p
  );


  buf

  (
    g408_n_spl_,
    g408_n
  );


  buf

  (
    G44_p_spl_,
    G44_p
  );


  buf

  (
    G44_p_spl_0,
    G44_p_spl_
  );


  buf

  (
    g409_n_spl_,
    g409_n
  );


  buf

  (
    g409_n_spl_0,
    g409_n_spl_
  );


  buf

  (
    g409_n_spl_00,
    g409_n_spl_0
  );


  buf

  (
    g409_n_spl_000,
    g409_n_spl_00
  );


  buf

  (
    g409_n_spl_001,
    g409_n_spl_00
  );


  buf

  (
    g409_n_spl_01,
    g409_n_spl_0
  );


  buf

  (
    g409_n_spl_010,
    g409_n_spl_01
  );


  buf

  (
    g409_n_spl_011,
    g409_n_spl_01
  );


  buf

  (
    g409_n_spl_1,
    g409_n_spl_
  );


  buf

  (
    g409_n_spl_10,
    g409_n_spl_1
  );


  buf

  (
    g409_n_spl_100,
    g409_n_spl_10
  );


  buf

  (
    g409_n_spl_101,
    g409_n_spl_10
  );


  buf

  (
    g409_n_spl_11,
    g409_n_spl_1
  );


  buf

  (
    g409_n_spl_110,
    g409_n_spl_11
  );


  buf

  (
    g409_n_spl_111,
    g409_n_spl_11
  );


  buf

  (
    G44_n_spl_,
    G44_n
  );


  buf

  (
    G44_n_spl_0,
    G44_n_spl_
  );


  buf

  (
    g409_p_spl_,
    g409_p
  );


  buf

  (
    g409_p_spl_0,
    g409_p_spl_
  );


  buf

  (
    g409_p_spl_00,
    g409_p_spl_0
  );


  buf

  (
    g409_p_spl_000,
    g409_p_spl_00
  );


  buf

  (
    g409_p_spl_001,
    g409_p_spl_00
  );


  buf

  (
    g409_p_spl_01,
    g409_p_spl_0
  );


  buf

  (
    g409_p_spl_010,
    g409_p_spl_01
  );


  buf

  (
    g409_p_spl_011,
    g409_p_spl_01
  );


  buf

  (
    g409_p_spl_1,
    g409_p_spl_
  );


  buf

  (
    g409_p_spl_10,
    g409_p_spl_1
  );


  buf

  (
    g409_p_spl_100,
    g409_p_spl_10
  );


  buf

  (
    g409_p_spl_101,
    g409_p_spl_10
  );


  buf

  (
    g409_p_spl_11,
    g409_p_spl_1
  );


  buf

  (
    g409_p_spl_110,
    g409_p_spl_11
  );


  buf

  (
    g409_p_spl_111,
    g409_p_spl_11
  );


  buf

  (
    G42_p_spl_,
    G42_p
  );


  buf

  (
    G42_p_spl_0,
    G42_p_spl_
  );


  buf

  (
    G42_p_spl_1,
    G42_p_spl_
  );


  buf

  (
    g412_n_spl_,
    g412_n
  );


  buf

  (
    g412_n_spl_0,
    g412_n_spl_
  );


  buf

  (
    g412_n_spl_00,
    g412_n_spl_0
  );


  buf

  (
    g412_n_spl_000,
    g412_n_spl_00
  );


  buf

  (
    g412_n_spl_0000,
    g412_n_spl_000
  );


  buf

  (
    g412_n_spl_0001,
    g412_n_spl_000
  );


  buf

  (
    g412_n_spl_001,
    g412_n_spl_00
  );


  buf

  (
    g412_n_spl_0010,
    g412_n_spl_001
  );


  buf

  (
    g412_n_spl_01,
    g412_n_spl_0
  );


  buf

  (
    g412_n_spl_010,
    g412_n_spl_01
  );


  buf

  (
    g412_n_spl_011,
    g412_n_spl_01
  );


  buf

  (
    g412_n_spl_1,
    g412_n_spl_
  );


  buf

  (
    g412_n_spl_10,
    g412_n_spl_1
  );


  buf

  (
    g412_n_spl_100,
    g412_n_spl_10
  );


  buf

  (
    g412_n_spl_101,
    g412_n_spl_10
  );


  buf

  (
    g412_n_spl_11,
    g412_n_spl_1
  );


  buf

  (
    g412_n_spl_110,
    g412_n_spl_11
  );


  buf

  (
    g412_n_spl_111,
    g412_n_spl_11
  );


  buf

  (
    G42_n_spl_,
    G42_n
  );


  buf

  (
    G42_n_spl_0,
    G42_n_spl_
  );


  buf

  (
    G42_n_spl_1,
    G42_n_spl_
  );


  buf

  (
    g412_p_spl_,
    g412_p
  );


  buf

  (
    g412_p_spl_0,
    g412_p_spl_
  );


  buf

  (
    g412_p_spl_00,
    g412_p_spl_0
  );


  buf

  (
    g412_p_spl_000,
    g412_p_spl_00
  );


  buf

  (
    g412_p_spl_0000,
    g412_p_spl_000
  );


  buf

  (
    g412_p_spl_0001,
    g412_p_spl_000
  );


  buf

  (
    g412_p_spl_001,
    g412_p_spl_00
  );


  buf

  (
    g412_p_spl_0010,
    g412_p_spl_001
  );


  buf

  (
    g412_p_spl_01,
    g412_p_spl_0
  );


  buf

  (
    g412_p_spl_010,
    g412_p_spl_01
  );


  buf

  (
    g412_p_spl_011,
    g412_p_spl_01
  );


  buf

  (
    g412_p_spl_1,
    g412_p_spl_
  );


  buf

  (
    g412_p_spl_10,
    g412_p_spl_1
  );


  buf

  (
    g412_p_spl_100,
    g412_p_spl_10
  );


  buf

  (
    g412_p_spl_101,
    g412_p_spl_10
  );


  buf

  (
    g412_p_spl_11,
    g412_p_spl_1
  );


  buf

  (
    g412_p_spl_110,
    g412_p_spl_11
  );


  buf

  (
    g412_p_spl_111,
    g412_p_spl_11
  );


  buf

  (
    g414_n_spl_,
    g414_n
  );


  buf

  (
    g414_n_spl_0,
    g414_n_spl_
  );


  buf

  (
    g414_n_spl_00,
    g414_n_spl_0
  );


  buf

  (
    g414_n_spl_000,
    g414_n_spl_00
  );


  buf

  (
    g414_n_spl_0000,
    g414_n_spl_000
  );


  buf

  (
    g414_n_spl_0001,
    g414_n_spl_000
  );


  buf

  (
    g414_n_spl_001,
    g414_n_spl_00
  );


  buf

  (
    g414_n_spl_01,
    g414_n_spl_0
  );


  buf

  (
    g414_n_spl_010,
    g414_n_spl_01
  );


  buf

  (
    g414_n_spl_011,
    g414_n_spl_01
  );


  buf

  (
    g414_n_spl_1,
    g414_n_spl_
  );


  buf

  (
    g414_n_spl_10,
    g414_n_spl_1
  );


  buf

  (
    g414_n_spl_100,
    g414_n_spl_10
  );


  buf

  (
    g414_n_spl_101,
    g414_n_spl_10
  );


  buf

  (
    g414_n_spl_11,
    g414_n_spl_1
  );


  buf

  (
    g414_n_spl_110,
    g414_n_spl_11
  );


  buf

  (
    g414_n_spl_111,
    g414_n_spl_11
  );


  buf

  (
    g414_p_spl_,
    g414_p
  );


  buf

  (
    g414_p_spl_0,
    g414_p_spl_
  );


  buf

  (
    g414_p_spl_00,
    g414_p_spl_0
  );


  buf

  (
    g414_p_spl_000,
    g414_p_spl_00
  );


  buf

  (
    g414_p_spl_0000,
    g414_p_spl_000
  );


  buf

  (
    g414_p_spl_0001,
    g414_p_spl_000
  );


  buf

  (
    g414_p_spl_001,
    g414_p_spl_00
  );


  buf

  (
    g414_p_spl_01,
    g414_p_spl_0
  );


  buf

  (
    g414_p_spl_010,
    g414_p_spl_01
  );


  buf

  (
    g414_p_spl_011,
    g414_p_spl_01
  );


  buf

  (
    g414_p_spl_1,
    g414_p_spl_
  );


  buf

  (
    g414_p_spl_10,
    g414_p_spl_1
  );


  buf

  (
    g414_p_spl_100,
    g414_p_spl_10
  );


  buf

  (
    g414_p_spl_101,
    g414_p_spl_10
  );


  buf

  (
    g414_p_spl_11,
    g414_p_spl_1
  );


  buf

  (
    g414_p_spl_110,
    g414_p_spl_11
  );


  buf

  (
    g414_p_spl_111,
    g414_p_spl_11
  );


  buf

  (
    G43_p_spl_,
    G43_p
  );


  buf

  (
    G43_p_spl_0,
    G43_p_spl_
  );


  buf

  (
    G43_p_spl_1,
    G43_p_spl_
  );


  buf

  (
    G43_n_spl_,
    G43_n
  );


  buf

  (
    G43_n_spl_0,
    G43_n_spl_
  );


  buf

  (
    G43_n_spl_1,
    G43_n_spl_
  );


  buf

  (
    g416_p_spl_,
    g416_p
  );


  buf

  (
    g416_n_spl_,
    g416_n
  );


  buf

  (
    g423_n_spl_,
    g423_n
  );


  buf

  (
    g423_n_spl_0,
    g423_n_spl_
  );


  buf

  (
    g423_n_spl_00,
    g423_n_spl_0
  );


  buf

  (
    g423_n_spl_000,
    g423_n_spl_00
  );


  buf

  (
    g423_n_spl_001,
    g423_n_spl_00
  );


  buf

  (
    g423_n_spl_01,
    g423_n_spl_0
  );


  buf

  (
    g423_n_spl_010,
    g423_n_spl_01
  );


  buf

  (
    g423_n_spl_011,
    g423_n_spl_01
  );


  buf

  (
    g423_n_spl_1,
    g423_n_spl_
  );


  buf

  (
    g423_n_spl_10,
    g423_n_spl_1
  );


  buf

  (
    g423_n_spl_11,
    g423_n_spl_1
  );


  buf

  (
    g423_p_spl_,
    g423_p
  );


  buf

  (
    g423_p_spl_0,
    g423_p_spl_
  );


  buf

  (
    g423_p_spl_00,
    g423_p_spl_0
  );


  buf

  (
    g423_p_spl_000,
    g423_p_spl_00
  );


  buf

  (
    g423_p_spl_001,
    g423_p_spl_00
  );


  buf

  (
    g423_p_spl_01,
    g423_p_spl_0
  );


  buf

  (
    g423_p_spl_010,
    g423_p_spl_01
  );


  buf

  (
    g423_p_spl_011,
    g423_p_spl_01
  );


  buf

  (
    g423_p_spl_1,
    g423_p_spl_
  );


  buf

  (
    g423_p_spl_10,
    g423_p_spl_1
  );


  buf

  (
    g423_p_spl_11,
    g423_p_spl_1
  );


  buf

  (
    g425_n_spl_,
    g425_n
  );


  buf

  (
    g425_n_spl_0,
    g425_n_spl_
  );


  buf

  (
    g425_n_spl_00,
    g425_n_spl_0
  );


  buf

  (
    g425_n_spl_000,
    g425_n_spl_00
  );


  buf

  (
    g425_n_spl_001,
    g425_n_spl_00
  );


  buf

  (
    g425_n_spl_01,
    g425_n_spl_0
  );


  buf

  (
    g425_n_spl_010,
    g425_n_spl_01
  );


  buf

  (
    g425_n_spl_011,
    g425_n_spl_01
  );


  buf

  (
    g425_n_spl_1,
    g425_n_spl_
  );


  buf

  (
    g425_n_spl_10,
    g425_n_spl_1
  );


  buf

  (
    g425_n_spl_100,
    g425_n_spl_10
  );


  buf

  (
    g425_n_spl_101,
    g425_n_spl_10
  );


  buf

  (
    g425_n_spl_11,
    g425_n_spl_1
  );


  buf

  (
    g425_p_spl_,
    g425_p
  );


  buf

  (
    g425_p_spl_0,
    g425_p_spl_
  );


  buf

  (
    g425_p_spl_00,
    g425_p_spl_0
  );


  buf

  (
    g425_p_spl_000,
    g425_p_spl_00
  );


  buf

  (
    g425_p_spl_001,
    g425_p_spl_00
  );


  buf

  (
    g425_p_spl_01,
    g425_p_spl_0
  );


  buf

  (
    g425_p_spl_010,
    g425_p_spl_01
  );


  buf

  (
    g425_p_spl_011,
    g425_p_spl_01
  );


  buf

  (
    g425_p_spl_1,
    g425_p_spl_
  );


  buf

  (
    g425_p_spl_10,
    g425_p_spl_1
  );


  buf

  (
    g425_p_spl_100,
    g425_p_spl_10
  );


  buf

  (
    g425_p_spl_101,
    g425_p_spl_10
  );


  buf

  (
    g425_p_spl_11,
    g425_p_spl_1
  );


  buf

  (
    g432_n_spl_,
    g432_n
  );


  buf

  (
    g432_p_spl_,
    g432_p
  );


  buf

  (
    g430_n_spl_,
    g430_n
  );


  buf

  (
    g430_p_spl_,
    g430_p
  );


  buf

  (
    g438_n_spl_,
    g438_n
  );


  buf

  (
    g438_p_spl_,
    g438_p
  );


  buf

  (
    g440_n_spl_,
    g440_n
  );


  buf

  (
    g441_n_spl_,
    g441_n
  );


  buf

  (
    g440_p_spl_,
    g440_p
  );


  buf

  (
    g441_p_spl_,
    g441_p
  );


  buf

  (
    g439_p_spl_,
    g439_p
  );


  buf

  (
    g439_n_spl_,
    g439_n
  );


  buf

  (
    g453_n_spl_,
    g453_n
  );


  buf

  (
    g453_p_spl_,
    g453_p
  );


  buf

  (
    g452_p_spl_,
    g452_p
  );


  buf

  (
    g452_p_spl_0,
    g452_p_spl_
  );


  buf

  (
    g452_p_spl_1,
    g452_p_spl_
  );


  buf

  (
    g456_p_spl_,
    g456_p
  );


  buf

  (
    g456_p_spl_0,
    g456_p_spl_
  );


  buf

  (
    g456_p_spl_1,
    g456_p_spl_
  );


  buf

  (
    g452_n_spl_,
    g452_n
  );


  buf

  (
    g452_n_spl_0,
    g452_n_spl_
  );


  buf

  (
    g452_n_spl_1,
    g452_n_spl_
  );


  buf

  (
    g456_n_spl_,
    g456_n
  );


  buf

  (
    g456_n_spl_0,
    g456_n_spl_
  );


  buf

  (
    g456_n_spl_1,
    g456_n_spl_
  );


  buf

  (
    G20_p_spl_,
    G20_p
  );


  buf

  (
    G20_p_spl_0,
    G20_p_spl_
  );


  buf

  (
    G20_p_spl_00,
    G20_p_spl_0
  );


  buf

  (
    G20_p_spl_1,
    G20_p_spl_
  );


  buf

  (
    G20_n_spl_,
    G20_n
  );


  buf

  (
    G20_n_spl_0,
    G20_n_spl_
  );


  buf

  (
    G20_n_spl_00,
    G20_n_spl_0
  );


  buf

  (
    G20_n_spl_1,
    G20_n_spl_
  );


  buf

  (
    G18_p_spl_,
    G18_p
  );


  buf

  (
    G18_p_spl_0,
    G18_p_spl_
  );


  buf

  (
    G18_p_spl_1,
    G18_p_spl_
  );


  buf

  (
    G18_n_spl_,
    G18_n
  );


  buf

  (
    G18_n_spl_0,
    G18_n_spl_
  );


  buf

  (
    G18_n_spl_1,
    G18_n_spl_
  );


  buf

  (
    G19_p_spl_,
    G19_p
  );


  buf

  (
    G19_p_spl_0,
    G19_p_spl_
  );


  buf

  (
    G19_p_spl_00,
    G19_p_spl_0
  );


  buf

  (
    G19_p_spl_1,
    G19_p_spl_
  );


  buf

  (
    G19_n_spl_,
    G19_n
  );


  buf

  (
    G19_n_spl_0,
    G19_n_spl_
  );


  buf

  (
    G19_n_spl_00,
    G19_n_spl_0
  );


  buf

  (
    G19_n_spl_1,
    G19_n_spl_
  );


  buf

  (
    g480_n_spl_,
    g480_n
  );


  buf

  (
    g480_p_spl_,
    g480_p
  );


  buf

  (
    g500_p_spl_,
    g500_p
  );


  buf

  (
    g500_p_spl_0,
    g500_p_spl_
  );


  buf

  (
    g500_n_spl_,
    g500_n
  );


  buf

  (
    g500_n_spl_0,
    g500_n_spl_
  );


  buf

  (
    g379_n_spl_,
    g379_n
  );


  buf

  (
    g379_n_spl_0,
    g379_n_spl_
  );


  buf

  (
    g379_n_spl_00,
    g379_n_spl_0
  );


  buf

  (
    g379_n_spl_01,
    g379_n_spl_0
  );


  buf

  (
    g379_n_spl_1,
    g379_n_spl_
  );


  buf

  (
    g503_n_spl_,
    g503_n
  );


  buf

  (
    g503_p_spl_,
    g503_p
  );


  buf

  (
    g501_p_spl_,
    g501_p
  );


  buf

  (
    g504_p_spl_,
    g504_p
  );


  buf

  (
    g501_n_spl_,
    g501_n
  );


  buf

  (
    g504_n_spl_,
    g504_n
  );


  buf

  (
    g510_n_spl_,
    g510_n
  );


  buf

  (
    g510_p_spl_,
    g510_p
  );


  buf

  (
    g514_n_spl_,
    g514_n
  );


  buf

  (
    g514_p_spl_,
    g514_p
  );


  buf

  (
    g513_p_spl_,
    g513_p
  );


  buf

  (
    g513_p_spl_0,
    g513_p_spl_
  );


  buf

  (
    g513_p_spl_00,
    g513_p_spl_0
  );


  buf

  (
    g513_p_spl_1,
    g513_p_spl_
  );


  buf

  (
    g517_p_spl_,
    g517_p
  );


  buf

  (
    g517_p_spl_0,
    g517_p_spl_
  );


  buf

  (
    g517_p_spl_00,
    g517_p_spl_0
  );


  buf

  (
    g517_p_spl_1,
    g517_p_spl_
  );


  buf

  (
    g513_n_spl_,
    g513_n
  );


  buf

  (
    g513_n_spl_0,
    g513_n_spl_
  );


  buf

  (
    g513_n_spl_00,
    g513_n_spl_0
  );


  buf

  (
    g513_n_spl_1,
    g513_n_spl_
  );


  buf

  (
    g517_n_spl_,
    g517_n
  );


  buf

  (
    g517_n_spl_0,
    g517_n_spl_
  );


  buf

  (
    g517_n_spl_00,
    g517_n_spl_0
  );


  buf

  (
    g517_n_spl_1,
    g517_n_spl_
  );


  buf

  (
    g518_p_spl_,
    g518_p
  );


  buf

  (
    g519_p_spl_,
    g519_p
  );


  buf

  (
    g518_n_spl_,
    g518_n
  );


  buf

  (
    g519_n_spl_,
    g519_n
  );


  buf

  (
    g349_n_spl_,
    g349_n
  );


  buf

  (
    g520_n_spl_,
    g520_n
  );


  buf

  (
    g521_p_spl_,
    g521_p
  );


  buf

  (
    g521_p_spl_0,
    g521_p_spl_
  );


  buf

  (
    g520_p_spl_,
    g520_p
  );


  buf

  (
    g521_n_spl_,
    g521_n
  );


  buf

  (
    g521_n_spl_0,
    g521_n_spl_
  );


  buf

  (
    g528_p_spl_,
    g528_p
  );


  buf

  (
    g528_n_spl_,
    g528_n
  );


  buf

  (
    g530_n_spl_,
    g530_n
  );


  buf

  (
    g530_n_spl_0,
    g530_n_spl_
  );


  buf

  (
    g530_p_spl_,
    g530_p
  );


  buf

  (
    g530_p_spl_0,
    g530_p_spl_
  );


  buf

  (
    g527_n_spl_,
    g527_n
  );


  buf

  (
    g527_n_spl_0,
    g527_n_spl_
  );


  buf

  (
    g534_n_spl_,
    g534_n
  );


  buf

  (
    g534_n_spl_0,
    g534_n_spl_
  );


  buf

  (
    g534_n_spl_1,
    g534_n_spl_
  );


  buf

  (
    g527_p_spl_,
    g527_p
  );


  buf

  (
    g527_p_spl_0,
    g527_p_spl_
  );


  buf

  (
    g534_p_spl_,
    g534_p
  );


  buf

  (
    g534_p_spl_0,
    g534_p_spl_
  );


  buf

  (
    g534_p_spl_1,
    g534_p_spl_
  );


  buf

  (
    g552_n_spl_,
    g552_n
  );


  buf

  (
    g552_p_spl_,
    g552_p
  );


  buf

  (
    g555_p_spl_,
    g555_p
  );


  buf

  (
    g555_p_spl_0,
    g555_p_spl_
  );


  buf

  (
    g555_n_spl_,
    g555_n
  );


  buf

  (
    g555_n_spl_0,
    g555_n_spl_
  );


  buf

  (
    g569_n_spl_,
    g569_n
  );


  buf

  (
    g569_p_spl_,
    g569_p
  );


  buf

  (
    g579_n_spl_,
    g579_n
  );


  buf

  (
    g579_p_spl_,
    g579_p
  );


  buf

  (
    g594_n_spl_,
    g594_n
  );


  buf

  (
    g594_p_spl_,
    g594_p
  );


  buf

  (
    g376_p_spl_,
    g376_p
  );


  buf

  (
    g376_p_spl_0,
    g376_p_spl_
  );


  buf

  (
    g597_n_spl_,
    g597_n
  );


  buf

  (
    g597_n_spl_0,
    g597_n_spl_
  );


  buf

  (
    g597_n_spl_00,
    g597_n_spl_0
  );


  buf

  (
    g597_n_spl_1,
    g597_n_spl_
  );


  buf

  (
    g376_n_spl_,
    g376_n
  );


  buf

  (
    g597_p_spl_,
    g597_p
  );


  buf

  (
    g597_p_spl_0,
    g597_p_spl_
  );


  buf

  (
    g597_p_spl_00,
    g597_p_spl_0
  );


  buf

  (
    g597_p_spl_1,
    g597_p_spl_
  );


  buf

  (
    g600_n_spl_,
    g600_n
  );


  buf

  (
    g600_p_spl_,
    g600_p
  );


  buf

  (
    g601_n_spl_,
    g601_n
  );


  buf

  (
    g601_p_spl_,
    g601_p
  );


  buf

  (
    g603_n_spl_,
    g603_n
  );


  buf

  (
    g603_p_spl_,
    g603_p
  );


  buf

  (
    g605_p_spl_,
    g605_p
  );


  buf

  (
    g605_n_spl_,
    g605_n
  );


  buf

  (
    g598_n_spl_,
    g598_n
  );


  buf

  (
    g608_n_spl_,
    g608_n
  );


  buf

  (
    g598_p_spl_,
    g598_p
  );


  buf

  (
    g608_p_spl_,
    g608_p
  );


  buf

  (
    g613_n_spl_,
    g613_n
  );


  buf

  (
    g613_p_spl_,
    g613_p
  );


  buf

  (
    g617_p_spl_,
    g617_p
  );


  buf

  (
    g617_n_spl_,
    g617_n
  );


  buf

  (
    g616_n_spl_,
    g616_n
  );


  buf

  (
    g616_n_spl_0,
    g616_n_spl_
  );


  buf

  (
    g616_n_spl_1,
    g616_n_spl_
  );


  buf

  (
    g620_n_spl_,
    g620_n
  );


  buf

  (
    g620_n_spl_0,
    g620_n_spl_
  );


  buf

  (
    g620_n_spl_1,
    g620_n_spl_
  );


  buf

  (
    g616_p_spl_,
    g616_p
  );


  buf

  (
    g616_p_spl_0,
    g616_p_spl_
  );


  buf

  (
    g616_p_spl_1,
    g616_p_spl_
  );


  buf

  (
    g620_p_spl_,
    g620_p
  );


  buf

  (
    g620_p_spl_0,
    g620_p_spl_
  );


  buf

  (
    g620_p_spl_1,
    g620_p_spl_
  );


  buf

  (
    g628_n_spl_,
    g628_n
  );


  buf

  (
    g628_n_spl_0,
    g628_n_spl_
  );


  buf

  (
    g628_p_spl_,
    g628_p
  );


  buf

  (
    g628_p_spl_0,
    g628_p_spl_
  );


  buf

  (
    g653_n_spl_,
    g653_n
  );


  buf

  (
    g654_n_spl_,
    g654_n
  );


  buf

  (
    g653_p_spl_,
    g653_p
  );


  buf

  (
    g654_p_spl_,
    g654_p
  );


  buf

  (
    g649_p_spl_,
    g649_p
  );


  buf

  (
    g649_n_spl_,
    g649_n
  );


  buf

  (
    g685_p_spl_,
    g685_p
  );


  buf

  (
    g685_n_spl_,
    g685_n
  );


  buf

  (
    g706_n_spl_,
    g706_n
  );


  buf

  (
    g706_p_spl_,
    g706_p
  );


  buf

  (
    g705_n_spl_,
    g705_n
  );


  buf

  (
    g705_p_spl_,
    g705_p
  );


  buf

  (
    g723_p_spl_,
    g723_p
  );


  buf

  (
    g723_n_spl_,
    g723_n
  );


  buf

  (
    g726_p_spl_,
    g726_p
  );


  buf

  (
    g726_n_spl_,
    g726_n
  );


  buf

  (
    g724_p_spl_,
    g724_p
  );


  buf

  (
    g724_p_spl_0,
    g724_p_spl_
  );


  buf

  (
    g729_p_spl_,
    g729_p
  );


  buf

  (
    g724_n_spl_,
    g724_n
  );


  buf

  (
    g724_n_spl_0,
    g724_n_spl_
  );


  buf

  (
    g729_n_spl_,
    g729_n
  );


  buf

  (
    g730_n_spl_,
    g730_n
  );


  buf

  (
    g730_n_spl_0,
    g730_n_spl_
  );


  buf

  (
    g730_p_spl_,
    g730_p
  );


  buf

  (
    g730_p_spl_0,
    g730_p_spl_
  );


  buf

  (
    g733_p_spl_,
    g733_p
  );


  buf

  (
    g735_n_spl_,
    g735_n
  );


  buf

  (
    g733_n_spl_,
    g733_n
  );


  buf

  (
    g735_p_spl_,
    g735_p
  );


  buf

  (
    g738_n_spl_,
    g738_n
  );


  buf

  (
    g738_n_spl_0,
    g738_n_spl_
  );


  buf

  (
    g738_n_spl_1,
    g738_n_spl_
  );


  buf

  (
    g740_n_spl_,
    g740_n
  );


  buf

  (
    g740_n_spl_0,
    g740_n_spl_
  );


  buf

  (
    g738_p_spl_,
    g738_p
  );


  buf

  (
    g738_p_spl_0,
    g738_p_spl_
  );


  buf

  (
    g738_p_spl_1,
    g738_p_spl_
  );


  buf

  (
    g740_p_spl_,
    g740_p
  );


  buf

  (
    g740_p_spl_0,
    g740_p_spl_
  );


  buf

  (
    g732_p_spl_,
    g732_p
  );


  buf

  (
    g732_p_spl_0,
    g732_p_spl_
  );


  buf

  (
    g732_p_spl_1,
    g732_p_spl_
  );


  buf

  (
    g741_n_spl_,
    g741_n
  );


  buf

  (
    g741_n_spl_0,
    g741_n_spl_
  );


  buf

  (
    g732_n_spl_,
    g732_n
  );


  buf

  (
    g732_n_spl_0,
    g732_n_spl_
  );


  buf

  (
    g732_n_spl_1,
    g732_n_spl_
  );


  buf

  (
    g741_p_spl_,
    g741_p
  );


  buf

  (
    g741_p_spl_0,
    g741_p_spl_
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


  buf

  (
    G17_p_spl_0,
    G17_p_spl_
  );


  buf

  (
    G17_n_spl_,
    G17_n
  );


  buf

  (
    G17_n_spl_0,
    G17_n_spl_
  );


  buf

  (
    G16_n_spl_,
    G16_n
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    g779_n_spl_,
    g779_n
  );


  buf

  (
    g779_p_spl_,
    g779_p
  );


  buf

  (
    g782_p_spl_,
    g782_p
  );


  buf

  (
    g782_p_spl_0,
    g782_p_spl_
  );


  buf

  (
    g782_n_spl_,
    g782_n
  );


  buf

  (
    g782_n_spl_0,
    g782_n_spl_
  );


  buf

  (
    g818_p_spl_,
    g818_p
  );


  buf

  (
    g818_n_spl_,
    g818_n
  );


  buf

  (
    g626_p_spl_,
    g626_p
  );


  buf

  (
    g722_p_spl_,
    g722_p
  );


  buf

  (
    g626_n_spl_,
    g626_n
  );


  buf

  (
    g626_n_spl_0,
    g626_n_spl_
  );


  buf

  (
    g722_n_spl_,
    g722_n
  );


  buf

  (
    g722_n_spl_0,
    g722_n_spl_
  );


  buf

  (
    g778_p_spl_,
    g778_p
  );


  buf

  (
    g827_p_spl_,
    g827_p
  );


  buf

  (
    g778_n_spl_,
    g778_n
  );


  buf

  (
    g778_n_spl_0,
    g778_n_spl_
  );


  buf

  (
    g827_n_spl_,
    g827_n
  );


  buf

  (
    g827_n_spl_0,
    g827_n_spl_
  );


  buf

  (
    g509_p_spl_,
    g509_p
  );


  buf

  (
    g866_p_spl_,
    g866_p
  );


  buf

  (
    g509_n_spl_,
    g509_n
  );


  buf

  (
    g509_n_spl_0,
    g509_n_spl_
  );


  buf

  (
    g866_n_spl_,
    g866_n
  );


  buf

  (
    g866_n_spl_0,
    g866_n_spl_
  );


  buf

  (
    g451_p_spl_,
    g451_p
  );


  buf

  (
    g679_p_spl_,
    g679_p
  );


  buf

  (
    g451_n_spl_,
    g451_n
  );


  buf

  (
    g451_n_spl_0,
    g451_n_spl_
  );


  buf

  (
    g679_n_spl_,
    g679_n
  );


  buf

  (
    g679_n_spl_0,
    g679_n_spl_
  );


  buf

  (
    g869_n_spl_,
    g869_n
  );


  buf

  (
    g870_n_spl_,
    g870_n
  );


  buf

  (
    g868_n_spl_,
    g868_n
  );


  buf

  (
    g868_n_spl_0,
    g868_n_spl_
  );


  buf

  (
    g867_n_spl_,
    g867_n
  );


  buf

  (
    g874_n_spl_,
    g874_n
  );


  buf

  (
    g873_n_spl_,
    g873_n
  );


  buf

  (
    g879_p_spl_,
    g879_p
  );


  buf

  (
    g881_n_spl_,
    g881_n
  );


  buf

  (
    g879_n_spl_,
    g879_n
  );


  buf

  (
    g881_p_spl_,
    g881_p
  );


  buf

  (
    G50_n_spl_,
    G50_n
  );


  buf

  (
    g888_n_spl_,
    g888_n
  );


  buf

  (
    g888_n_spl_0,
    g888_n_spl_
  );


  buf

  (
    g888_n_spl_1,
    g888_n_spl_
  );


  buf

  (
    G50_p_spl_,
    G50_p
  );


  buf

  (
    g888_p_spl_,
    g888_p
  );


  buf

  (
    g888_p_spl_0,
    g888_p_spl_
  );


  buf

  (
    g888_p_spl_1,
    g888_p_spl_
  );


  buf

  (
    g886_p_spl_,
    g886_p
  );


  buf

  (
    g886_p_spl_0,
    g886_p_spl_
  );


  buf

  (
    g886_p_spl_1,
    g886_p_spl_
  );


  buf

  (
    g892_n_spl_,
    g892_n
  );


  buf

  (
    g886_n_spl_,
    g886_n
  );


  buf

  (
    g886_n_spl_0,
    g886_n_spl_
  );


  buf

  (
    g886_n_spl_1,
    g886_n_spl_
  );


  buf

  (
    g892_p_spl_,
    g892_p
  );


  buf

  (
    g884_n_spl_,
    g884_n
  );


  buf

  (
    g884_p_spl_,
    g884_p
  );


endmodule
