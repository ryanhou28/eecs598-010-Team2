// Benchmark "mymod" written by ABC on Sun Oct 29 19:31:50 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58,
    G59, G60,
    G855, G856, G857, G858, G859, G860, G861, G862, G863, G864, G865, G866,
    G867, G868, G869, G870, G871, G872, G873, G874, G875, G876, G877, G878,
    G879, G880  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G58, G59, G60;
  output G855, G856, G857, G858, G859, G860, G861, G862, G863, G864, G865,
    G866, G867, G868, G869, G870, G871, G872, G873, G874, G875, G876, G877,
    G878, G879, G880;
  reg n480_lo, n492_lo, n495_lo, n498_lo, n501_lo, n504_lo, n516_lo,
    n528_lo, n531_lo, n540_lo, n543_lo, n546_lo, n549_lo, n552_lo, n564_lo,
    n579_lo, n600_lo, n603_lo, n606_lo, n609_lo, n612_lo, n615_lo, n618_lo,
    n621_lo, n627_lo, n630_lo, n633_lo, n639_lo, n642_lo, n645_lo, n648_lo,
    n660_lo, n663_lo, n672_lo, n675_lo, n678_lo, n681_lo, n684_lo, n687_lo,
    n690_lo, n693_lo, n696_lo, n699_lo, n702_lo, n705_lo, n708_lo, n711_lo,
    n714_lo, n717_lo, n720_lo, n723_lo, n726_lo, n729_lo, n732_lo, n735_lo,
    n738_lo, n741_lo, n744_lo, n747_lo, n750_lo, n756_lo, n759_lo, n762_lo,
    n768_lo, n771_lo, n774_lo, n780_lo, n783_lo, n786_lo, n792_lo, n795_lo,
    n804_lo, n807_lo, n816_lo, n819_lo, n828_lo, n831_lo, n843_lo, n846_lo,
    n849_lo, n852_lo, n855_lo, n858_lo, n861_lo, n864_lo, n867_lo, n870_lo,
    n879_lo, n891_lo, n903_lo, n915_lo, n918_lo, n927_lo, n951_lo, n954_lo,
    n957_lo, n960_lo, n963_lo, n966_lo, n972_lo, n975_lo, n978_lo, n984_lo,
    n987_lo, n990_lo, n996_lo, n999_lo, n1002_lo, n1008_lo, n1011_lo,
    n1014_lo, n1020_lo, n1023_lo, n1026_lo, n1032_lo, n1035_lo, n1038_lo,
    n1044_lo, n1047_lo, n1050_lo, n1053_lo, n1056_lo, n1059_lo, n1062_lo,
    n1065_lo, n1068_lo, n1071_lo, n1074_lo, n1077_lo, n1080_lo, n1083_lo,
    n1086_lo, n1089_lo, n1092_lo, n1095_lo, n1098_lo, n1101_lo, n1104_lo,
    n1107_lo, n1110_lo, n1113_lo, n1116_lo, n1119_lo, n1122_lo, n1125_lo,
    n1128_lo, n1131_lo, n1134_lo, n1137_lo, n1140_lo, n1143_lo, n1146_lo,
    n1149_lo, n1152_lo, n1155_lo, n1158_lo, n1167_lo, n1170_lo, n1173_lo,
    n1176_lo, n1179_lo, n1529_o2, n1616_o2, n1655_o2, n1656_o2, n1657_o2,
    n1730_o2, n1731_o2, n1732_o2, n1729_o2, n1805_o2, n1808_o2, n1807_o2,
    n1809_o2, n1663_o2, n1664_o2, n1704_o2, n1705_o2, n1706_o2, n1707_o2,
    n1708_o2, n1709_o2, G280_o2, G655_o2, G663_o2, G672_o2, G538_o2,
    n1780_o2, n1781_o2, n1797_o2, n1798_o2, n1799_o2, n1800_o2, G578_o2,
    n1828_o2, n801_lo_buf_o2, G693_o2, G702_o2, G712_o2, G685_o2, G658_o2,
    G667_o2, G677_o2, G650_o2, G798_o2, n1017_lo_buf_o2, n1029_lo_buf_o2,
    n1041_lo_buf_o2, G558_o2, G562_o2, G566_o2, n1835_o2, n1836_o2,
    n1837_o2, n765_lo_buf_o2, n777_lo_buf_o2, n789_lo_buf_o2, G617_o2,
    G626_o2, G636_o2, n489_lo_buf_o2, n513_lo_buf_o2, n561_lo_buf_o2,
    n597_lo_buf_o2, n657_lo_buf_o2, G276_o2, n1005_lo_buf_o2,
    n1161_lo_buf_o2, G620_o2, G629_o2, G639_o2, G554_o2, G690_o2, G698_o2,
    G707_o2, G319_o2, G389_o2, n753_lo_buf_o2, G647_o2, G769_o2, G785_o2,
    G808_o2, G445_o2, G448_o2, G477_o2, G480_o2, G436_o2, G786_o2, G787_o2,
    G826_o2, G827_o2, G825_o2, G610_o2, n537_lo_buf_o2, n669_lo_buf_o2,
    n969_lo_buf_o2, n981_lo_buf_o2, n993_lo_buf_o2, G309_o2, G461_o2,
    G487_o2, G460_o2, G468_o2, G287_o2, G613_o2, n585_lo_buf_o2,
    n813_lo_buf_o2, n825_lo_buf_o2, n837_lo_buf_o2, n897_lo_buf_o2,
    n909_lo_buf_o2, n933_lo_buf_o2, G451_o2, G682_o2, G756_o2, G542_o2,
    G546_o2, G550_o2, G310_o2, n798_lo_buf_o2, n882_lo_buf_o2, G427_o2,
    G497_o2, G499_o2, G501_o2, G498_o2, G500_o2, G502_o2, G369_o2,
    n939_lo_buf_o2, n486_lo_buf_o2, n510_lo_buf_o2, n558_lo_buf_o2,
    n594_lo_buf_o2, n654_lo_buf_o2, n477_lo_buf_o2, n525_lo_buf_o2,
    n573_lo_buf_o2;
  wire new_new_n683__, new_new_n685__, new_new_n687__, new_new_n689__,
    new_new_n691__, new_new_n693__, new_new_n695__, new_new_n697__,
    new_new_n699__, new_new_n701__, new_new_n703__, new_new_n705__,
    new_new_n707__, new_new_n709__, new_new_n711__, new_new_n713__,
    new_new_n715__, new_new_n717__, new_new_n719__, new_new_n721__,
    new_new_n723__, new_new_n725__, new_new_n727__, new_new_n729__,
    new_new_n731__, new_new_n733__, new_new_n735__, new_new_n737__,
    new_new_n739__, new_new_n741__, new_new_n743__, new_new_n745__,
    new_new_n747__, new_new_n749__, new_new_n751__, new_new_n753__,
    new_new_n755__, new_new_n757__, new_new_n759__, new_new_n761__,
    new_new_n763__, new_new_n765__, new_new_n767__, new_new_n769__,
    new_new_n771__, new_new_n773__, new_new_n775__, new_new_n777__,
    new_new_n779__, new_new_n781__, new_new_n783__, new_new_n785__,
    new_new_n787__, new_new_n789__, new_new_n791__, new_new_n793__,
    new_new_n795__, new_new_n797__, new_new_n799__, new_new_n801__,
    new_new_n803__, new_new_n804__, new_new_n806__, new_new_n807__,
    new_new_n809__, new_new_n811__, new_new_n812__, new_new_n813__,
    new_new_n814__, new_new_n815__, new_new_n816__, new_new_n817__,
    new_new_n818__, new_new_n819__, new_new_n820__, new_new_n822__,
    new_new_n823__, new_new_n825__, new_new_n827__, new_new_n830__,
    new_new_n832__, new_new_n833__, new_new_n834__, new_new_n835__,
    new_new_n836__, new_new_n837__, new_new_n839__, new_new_n841__,
    new_new_n842__, new_new_n844__, new_new_n845__, new_new_n847__,
    new_new_n850__, new_new_n851__, new_new_n853__, new_new_n856__,
    new_new_n857__, new_new_n859__, new_new_n861__, new_new_n864__,
    new_new_n865__, new_new_n866__, new_new_n867__, new_new_n868__,
    new_new_n869__, new_new_n870__, new_new_n871__, new_new_n873__,
    new_new_n875__, new_new_n878__, new_new_n879__, new_new_n881__,
    new_new_n883__, new_new_n886__, new_new_n887__, new_new_n889__,
    new_new_n891__, new_new_n893__, new_new_n895__, new_new_n897__,
    new_new_n899__, new_new_n901__, new_new_n903__, new_new_n905__,
    new_new_n907__, new_new_n909__, new_new_n911__, new_new_n913__,
    new_new_n915__, new_new_n917__, new_new_n919__, new_new_n921__,
    new_new_n924__, new_new_n925__, new_new_n927__, new_new_n928__,
    new_new_n930__, new_new_n931__, new_new_n933__, new_new_n934__,
    new_new_n936__, new_new_n937__, new_new_n939__, new_new_n940__,
    new_new_n942__, new_new_n943__, new_new_n946__, new_new_n947__,
    new_new_n950__, new_new_n951__, new_new_n954__, new_new_n955__,
    new_new_n957__, new_new_n959__, new_new_n961__, new_new_n963__,
    new_new_n964__, new_new_n965__, new_new_n967__, new_new_n969__,
    new_new_n971__, new_new_n972__, new_new_n973__, new_new_n975__,
    new_new_n976__, new_new_n977__, new_new_n979__, new_new_n981__,
    new_new_n983__, new_new_n986__, new_new_n987__, new_new_n989__,
    new_new_n991__, new_new_n993__, new_new_n994__, new_new_n996__,
    new_new_n997__, new_new_n999__, new_new_n1002__, new_new_n1003__,
    new_new_n1005__, new_new_n1008__, new_new_n1009__, new_new_n1011__,
    new_new_n1014__, new_new_n1015__, new_new_n1017__, new_new_n1018__,
    new_new_n1020__, new_new_n1021__, new_new_n1023__, new_new_n1024__,
    new_new_n1026__, new_new_n1027__, new_new_n1029__, new_new_n1030__,
    new_new_n1032__, new_new_n1033__, new_new_n1035__, new_new_n1036__,
    new_new_n1038__, new_new_n1039__, new_new_n1041__, new_new_n1043__,
    new_new_n1045__, new_new_n1046__, new_new_n1047__, new_new_n1049__,
    new_new_n1051__, new_new_n1054__, new_new_n1055__, new_new_n1057__,
    new_new_n1059__, new_new_n1062__, new_new_n1063__, new_new_n1065__,
    new_new_n1067__, new_new_n1070__, new_new_n1071__, new_new_n1073__,
    new_new_n1075__, new_new_n1078__, new_new_n1079__, new_new_n1081__,
    new_new_n1083__, new_new_n1086__, new_new_n1087__, new_new_n1089__,
    new_new_n1091__, new_new_n1094__, new_new_n1095__, new_new_n1097__,
    new_new_n1099__, new_new_n1102__, new_new_n1103__, new_new_n1105__,
    new_new_n1107__, new_new_n1110__, new_new_n1111__, new_new_n1113__,
    new_new_n1114__, new_new_n1115__, new_new_n1117__, new_new_n1119__,
    new_new_n1122__, new_new_n1123__, new_new_n1126__, new_new_n1128__,
    new_new_n1130__, new_new_n1132__, new_new_n1134__, new_new_n1136__,
    new_new_n1138__, new_new_n1140__, new_new_n1142__, new_new_n1144__,
    new_new_n1146__, new_new_n1148__, new_new_n1150__, new_new_n1151__,
    new_new_n1152__, new_new_n1153__, new_new_n1155__, new_new_n1156__,
    new_new_n1157__, new_new_n1159__, new_new_n1160__, new_new_n1161__,
    new_new_n1162__, new_new_n1163__, new_new_n1165__, new_new_n1168__,
    new_new_n1170__, new_new_n1172__, new_new_n1174__, new_new_n1176__,
    new_new_n1177__, new_new_n1179__, new_new_n1182__, new_new_n1183__,
    new_new_n1184__, new_new_n1185__, new_new_n1186__, new_new_n1187__,
    new_new_n1188__, new_new_n1190__, new_new_n1191__, new_new_n1193__,
    new_new_n1194__, new_new_n1196__, new_new_n1198__, new_new_n1200__,
    new_new_n1202__, new_new_n1204__, new_new_n1206__, new_new_n1208__,
    new_new_n1210__, new_new_n1212__, new_new_n1213__, new_new_n1214__,
    new_new_n1215__, new_new_n1216__, new_new_n1217__, new_new_n1218__,
    new_new_n1219__, new_new_n1221__, new_new_n1223__, new_new_n1225__,
    new_new_n1227__, new_new_n1230__, new_new_n1231__, new_new_n1232__,
    new_new_n1233__, new_new_n1234__, new_new_n1235__, new_new_n1236__,
    new_new_n1237__, new_new_n1238__, new_new_n1239__, new_new_n1240__,
    new_new_n1241__, new_new_n1242__, new_new_n1243__, new_new_n1245__,
    new_new_n1246__, new_new_n1247__, new_new_n1249__, new_new_n1251__,
    new_new_n1253__, new_new_n1255__, new_new_n1256__, new_new_n1257__,
    new_new_n1258__, new_new_n1259__, new_new_n1260__, new_new_n1261__,
    new_new_n1262__, new_new_n1263__, new_new_n1264__, new_new_n1265__,
    new_new_n1267__, new_new_n1269__, new_new_n1270__, new_new_n1271__,
    new_new_n1272__, new_new_n1273__, new_new_n1276__, new_new_n1277__,
    new_new_n1278__, new_new_n1280__, new_new_n1282__, new_new_n1284__,
    new_new_n1286__, new_new_n1287__, new_new_n1288__, new_new_n1289__,
    new_new_n1290__, new_new_n1291__, new_new_n1292__, new_new_n1293__,
    new_new_n1294__, new_new_n1296__, new_new_n1298__, new_new_n1300__,
    new_new_n1302__, new_new_n1304__, new_new_n1306__, new_new_n1307__,
    new_new_n1308__, new_new_n1309__, new_new_n1311__, new_new_n1313__,
    new_new_n1314__, new_new_n1315__, new_new_n1316__, new_new_n1317__,
    new_new_n1318__, new_new_n1319__, new_new_n1320__, new_new_n1321__,
    new_new_n1322__, new_new_n1323__, new_new_n1324__, new_new_n1325__,
    new_new_n1326__, new_new_n1327__, new_new_n1330__, new_new_n1331__,
    new_new_n1332__, new_new_n1333__, new_new_n1334__, new_new_n1335__,
    new_new_n1337__, new_new_n1339__, new_new_n1342__, new_new_n1344__,
    new_new_n1346__, new_new_n1347__, new_new_n1348__, new_new_n1349__,
    new_new_n1350__, new_new_n1351__, new_new_n1352__, new_new_n1353__,
    new_new_n1354__, new_new_n1355__, new_new_n1356__, new_new_n1357__,
    new_new_n1358__, new_new_n1359__, new_new_n1361__, new_new_n1362__,
    new_new_n1364__, new_new_n1366__, new_new_n1368__, new_new_n1370__,
    new_new_n1372__, new_new_n1374__, new_new_n1376__, new_new_n1378__,
    new_new_n1379__, new_new_n1381__, new_new_n1382__, new_new_n1383__,
    new_new_n1385__, new_new_n1386__, new_new_n1387__, new_new_n1388__,
    new_new_n1389__, new_new_n1390__, new_new_n1391__, new_new_n1392__,
    new_new_n1393__, new_new_n1394__, new_new_n1395__, new_new_n1396__,
    new_new_n1397__, new_new_n1398__, new_new_n1399__, new_new_n1400__,
    new_new_n1401__, new_new_n1402__, new_new_n1403__, new_new_n1404__,
    new_new_n1405__, new_new_n1406__, new_new_n1407__, new_new_n1408__,
    new_new_n1409__, new_new_n1410__, new_new_n1411__, new_new_n1412__,
    new_new_n1413__, new_new_n1414__, new_new_n1415__, new_new_n1416__,
    new_new_n1417__, new_new_n1418__, new_new_n1419__, new_new_n1420__,
    new_new_n1421__, new_new_n1422__, new_new_n1423__, new_new_n1424__,
    new_new_n1425__, new_new_n1426__, new_new_n1427__, new_new_n1428__,
    new_new_n1429__, new_new_n1430__, new_new_n1431__, new_new_n1432__,
    new_new_n1433__, new_new_n1434__, new_new_n1435__, new_new_n1436__,
    new_new_n1437__, new_new_n1438__, new_new_n1439__, new_new_n1440__,
    new_new_n1441__, new_new_n1442__, new_new_n1443__, new_new_n1444__,
    new_new_n1445__, new_new_n1446__, new_new_n1447__, new_new_n1448__,
    new_new_n1449__, new_new_n1450__, new_new_n1451__, new_new_n1452__,
    new_new_n1453__, new_new_n1454__, new_new_n1455__, new_new_n1456__,
    new_new_n1457__, new_new_n1458__, new_new_n1459__, new_new_n1460__,
    new_new_n1461__, new_new_n1462__, new_new_n1463__, new_new_n1464__,
    new_new_n1465__, new_new_n1466__, new_new_n1467__, new_new_n1468__,
    new_new_n1469__, new_new_n1470__, new_new_n1471__, new_new_n1472__,
    new_new_n1473__, new_new_n1474__, new_new_n1475__, new_new_n1476__,
    new_new_n1477__, new_new_n1478__, new_new_n1479__, new_new_n1480__,
    new_new_n1481__, new_new_n1482__, new_new_n1483__, new_new_n1484__,
    new_new_n1485__, new_new_n1486__, new_new_n1487__, new_new_n1488__,
    new_new_n1489__, new_new_n1490__, new_new_n1491__, new_new_n1492__,
    new_new_n1493__, new_new_n1494__, new_new_n1495__, new_new_n1496__,
    new_new_n1497__, new_new_n1498__, new_new_n1499__, new_new_n1500__,
    new_new_n1501__, new_new_n1502__, new_new_n1503__, new_new_n1504__,
    new_new_n1505__, new_new_n1506__, new_new_n1507__, new_new_n1508__,
    new_new_n1509__, new_new_n1510__, new_new_n1511__, new_new_n1512__,
    new_new_n1513__, new_new_n1514__, new_new_n1515__, new_new_n1516__,
    new_new_n1517__, new_new_n1518__, new_new_n1519__, new_new_n1520__,
    new_new_n1521__, new_new_n1522__, new_new_n1523__, new_new_n1524__,
    new_new_n1525__, new_new_n1526__, new_new_n1527__, new_new_n1528__,
    new_new_n1529__, new_new_n1530__, new_new_n1531__, new_new_n1532__,
    new_new_n1533__, new_new_n1534__, new_new_n1535__, new_new_n1536__,
    new_new_n1537__, new_new_n1538__, new_new_n1539__, new_new_n1540__,
    new_new_n1541__, new_new_n1542__, new_new_n1543__, new_new_n1544__,
    new_new_n1545__, new_new_n1546__, new_new_n1547__, new_new_n1548__,
    new_new_n1549__, new_new_n1550__, new_new_n1551__, new_new_n1552__,
    new_new_n1553__, new_new_n1554__, new_new_n1555__, new_new_n1556__,
    new_new_n1557__, new_new_n1558__, new_new_n1559__, new_new_n1560__,
    new_new_n1561__, new_new_n1562__, new_new_n1563__, new_new_n1564__,
    new_new_n1565__, new_new_n1566__, new_new_n1567__, new_new_n1568__,
    new_new_n1569__, new_new_n1570__, new_new_n1571__, new_new_n1572__,
    new_new_n1573__, new_new_n1574__, new_new_n1575__, new_new_n1576__,
    new_new_n1577__, new_new_n1578__, new_new_n1579__, new_new_n1580__,
    new_new_n1581__, new_new_n1582__, new_new_n1583__, new_new_n1584__,
    new_new_n1585__, new_new_n1586__, new_new_n1587__, new_new_n1588__,
    new_new_n1589__, new_new_n1590__, new_new_n1591__, new_new_n1592__,
    new_new_n1593__, new_new_n1594__, new_new_n1595__, new_new_n1596__,
    new_new_n1597__, new_new_n1598__, new_new_n1599__, new_new_n1600__,
    new_new_n1601__, new_new_n1602__, new_new_n1603__, new_new_n1604__,
    new_new_n1605__, new_new_n1606__, new_new_n1607__, new_new_n1608__,
    new_new_n1609__, new_new_n1610__, new_new_n1611__, new_new_n1612__,
    new_new_n1613__, new_new_n1614__, new_new_n1615__, new_new_n1616__,
    new_new_n1617__, new_new_n1618__, new_new_n1619__, new_new_n1620__,
    new_new_n1621__, new_new_n1622__, new_new_n1623__, new_new_n1624__,
    new_new_n1625__, new_new_n1626__, new_new_n1627__, new_new_n1628__,
    new_new_n1629__, new_new_n1630__, new_new_n1631__, new_new_n1632__,
    new_new_n1633__, new_new_n1634__, new_new_n1635__, new_new_n1636__,
    new_new_n1637__, new_new_n1638__, new_new_n1639__, new_new_n1640__,
    new_new_n1641__, new_new_n1642__, new_new_n1643__, new_new_n1644__,
    new_new_n1645__, new_new_n1646__, new_new_n1647__, new_new_n1648__,
    new_new_n1649__, new_new_n1650__, new_new_n1651__, new_new_n1652__,
    new_new_n1653__, new_new_n1654__, new_new_n1655__, new_new_n1656__,
    new_new_n1657__, new_new_n1658__, new_new_n1659__, new_new_n1660__,
    new_new_n1661__, new_new_n1662__, new_new_n1663__, new_new_n1664__,
    new_new_n1665__, new_new_n1666__, new_new_n1667__, new_new_n1668__,
    new_new_n1669__, new_new_n1670__, new_new_n1671__, new_new_n1672__,
    new_new_n1673__, new_new_n1674__, new_new_n1675__, new_new_n1676__,
    new_new_n1677__, new_new_n1678__, new_new_n1679__, new_new_n1680__,
    new_new_n1681__, new_new_n1682__, new_new_n1683__, new_new_n1684__,
    new_new_n1685__, new_new_n1686__, new_new_n1687__, new_new_n1688__,
    new_new_n1689__, new_new_n1690__, new_new_n1691__, new_new_n1692__,
    new_new_n1693__, new_new_n1694__, new_new_n1695__, new_new_n1696__,
    new_new_n1697__, new_new_n1698__, new_new_n1699__, new_new_n1700__,
    new_new_n1701__, new_new_n1702__, new_new_n1703__, new_new_n1704__,
    new_new_n1705__, new_new_n1706__, new_new_n1707__, new_new_n1708__,
    new_new_n1709__, new_new_n1710__, new_new_n1711__, new_new_n1712__,
    new_new_n1713__, new_new_n1714__, new_new_n1715__, new_new_n1716__,
    new_new_n1717__, new_new_n1718__, new_new_n1719__, new_new_n1720__,
    new_new_n1721__, new_new_n1722__, new_new_n1723__, new_new_n1724__,
    new_new_n1725__, new_new_n1726__, new_new_n1727__, new_new_n1728__,
    new_new_n1729__, new_new_n1730__, new_new_n1731__, new_new_n1732__,
    new_new_n1733__, new_new_n1734__, new_new_n1735__, new_new_n1736__,
    new_new_n1737__, new_new_n1738__, new_new_n1739__, new_new_n1740__,
    new_new_n1741__, new_new_n1742__, new_new_n1743__, new_new_n1744__,
    new_new_n1745__, new_new_n1746__, new_new_n1747__, new_new_n1748__,
    new_new_n1749__, new_new_n1750__, new_new_n1751__, new_new_n1752__,
    new_new_n1753__, new_new_n1754__, new_new_n1755__, new_new_n1756__,
    new_new_n1757__, new_new_n1758__, new_new_n1759__, new_new_n1760__,
    new_new_n1761__, new_new_n1762__, new_new_n1763__, new_new_n1764__,
    new_new_n1765__, new_new_n1766__, new_new_n1767__, new_new_n1768__,
    new_new_n1769__, new_new_n1770__, new_new_n1771__, new_new_n1772__,
    new_new_n1773__, new_new_n1774__, new_new_n1775__, new_new_n1776__,
    new_new_n1777__, new_new_n1778__, new_new_n1779__, new_new_n1780__,
    new_new_n1781__, new_new_n1782__, new_new_n1783__, new_new_n1784__,
    new_new_n1785__, new_new_n1786__, new_new_n1787__, new_new_n1788__,
    new_new_n1789__, new_new_n1790__, new_new_n1791__, new_new_n1792__,
    new_new_n1793__, new_new_n1794__, new_new_n1795__, new_new_n1796__,
    new_new_n1797__, new_new_n1798__, new_new_n1799__, new_new_n1800__,
    new_new_n1801__, new_new_n1802__, new_new_n1803__, new_new_n1804__,
    new_new_n1805__, new_new_n1806__, new_new_n1807__, new_new_n1808__,
    new_new_n1809__, new_new_n1810__, new_new_n1811__, new_new_n1812__,
    new_new_n1813__, new_new_n1814__, new_new_n1815__, new_new_n1816__,
    new_new_n2141__, new_new_n2142__, new_new_n2143__, new_new_n2144__,
    new_new_n2145__, new_new_n2146__, new_new_n2147__, new_new_n2148__,
    new_new_n2149__, new_new_n2150__, new_new_n2151__, new_new_n2152__,
    new_new_n2153__, new_new_n2154__, new_new_n2155__, new_new_n2156__,
    new_new_n2157__, new_new_n2158__, new_new_n2159__, new_new_n2160__,
    new_new_n2161__, new_new_n2162__, new_new_n2163__, new_new_n2164__,
    new_new_n2165__, new_new_n2166__, new_new_n2167__, new_new_n2168__,
    new_new_n2169__, new_new_n2170__, new_new_n2171__, new_new_n2172__,
    new_new_n2173__, new_new_n2174__, new_new_n2175__, new_new_n2176__,
    new_new_n2177__, new_new_n2178__, new_new_n2179__, new_new_n2180__,
    new_new_n2181__, new_new_n2182__, new_new_n2183__, new_new_n2184__,
    new_new_n2185__, new_new_n2186__, new_new_n2187__, new_new_n2188__,
    new_new_n2189__, new_new_n2190__, new_new_n2191__, new_new_n2192__,
    new_new_n2193__, new_new_n2194__, new_new_n2195__, new_new_n2196__,
    new_new_n2197__, new_new_n2198__, new_new_n2199__, new_new_n2200__,
    new_new_n2201__, new_new_n2202__, new_new_n2203__, new_new_n2204__,
    new_new_n2205__, new_new_n2206__, new_new_n2207__, new_new_n2208__,
    new_new_n2209__, new_new_n2210__, new_new_n2211__, new_new_n2212__,
    new_new_n2213__, new_new_n2214__, new_new_n2215__, new_new_n2216__,
    new_new_n2217__, new_new_n2218__, new_new_n2219__, new_new_n2220__,
    new_new_n2221__, new_new_n2222__, new_new_n2223__, new_new_n2224__,
    new_new_n2225__, new_new_n2226__, new_new_n2227__, new_new_n2228__,
    new_new_n2229__, new_new_n2230__, new_new_n2231__, new_new_n2232__,
    new_new_n2233__, new_new_n2234__, new_new_n2235__, new_new_n2236__,
    new_new_n2237__, new_new_n2238__, new_new_n2239__, new_new_n2240__,
    new_new_n2241__, new_new_n2242__, new_new_n2243__, new_new_n2244__,
    new_new_n2245__, new_new_n2246__, new_new_n2247__, new_new_n2248__,
    new_new_n2249__, new_new_n2250__, new_new_n2251__, new_new_n2252__,
    new_new_n2253__, new_new_n2254__, new_new_n2255__, new_new_n2256__,
    new_new_n2257__, new_new_n2258__, new_new_n2259__, new_new_n2260__,
    new_new_n2261__, new_new_n2262__, new_new_n2263__, new_new_n2264__,
    new_new_n2265__, new_new_n2266__, new_new_n2267__, new_new_n2268__,
    new_new_n2269__, new_new_n2270__, new_new_n2271__, new_new_n2272__,
    new_new_n2273__, new_new_n2274__, new_new_n2275__, new_new_n2276__,
    new_new_n2277__, new_new_n2278__, new_new_n2279__, new_new_n2280__,
    new_new_n2281__, new_new_n2282__, new_new_n2283__, new_new_n2284__,
    new_new_n2285__, new_new_n2286__, new_new_n2287__, new_new_n2288__,
    new_new_n2289__, new_new_n2290__, new_new_n2291__, new_new_n2292__,
    new_new_n2293__, new_new_n2294__, new_new_n2295__, new_new_n2296__,
    new_new_n2297__, new_new_n2298__, new_new_n2299__, new_new_n2300__,
    new_new_n2301__, new_new_n2302__, new_new_n2303__, new_new_n2304__,
    new_new_n2305__, new_new_n2306__, new_new_n2307__, new_new_n2308__,
    new_new_n2309__, new_new_n2310__, new_new_n2311__, new_new_n2312__,
    new_new_n2313__, new_new_n2314__, new_new_n2315__, new_new_n2316__,
    new_new_n2317__, new_new_n2318__, new_new_n2319__, new_new_n2320__,
    new_new_n2321__, new_new_n2322__, new_new_n2323__, new_new_n2324__,
    new_new_n2325__, new_new_n2326__, new_new_n2327__, new_new_n2328__,
    new_new_n2329__, new_new_n2330__, new_new_n2331__, new_new_n2332__,
    new_new_n2333__, new_new_n2334__, new_new_n2335__, new_new_n2336__,
    new_new_n2337__, new_new_n2338__, new_new_n2339__, new_new_n2340__,
    new_new_n2341__, new_new_n2342__, new_new_n2343__, new_new_n2344__,
    new_new_n2345__, new_new_n2346__, new_new_n2347__, new_new_n2348__,
    new_new_n2349__, new_new_n2350__, new_new_n2351__, new_new_n2352__,
    new_new_n2353__, new_new_n2354__, new_new_n2355__, new_new_n2356__,
    new_new_n2357__, new_new_n2358__, new_new_n2359__, new_new_n2360__,
    new_new_n2361__, new_new_n2362__, new_new_n2363__, new_new_n2364__,
    new_new_n2365__, new_new_n2366__, new_new_n2367__, new_new_n2368__,
    new_new_n2369__, new_new_n2370__, new_new_n2371__, new_new_n2372__,
    new_new_n2373__, new_new_n2374__, new_new_n2375__, new_new_n2376__,
    new_new_n2377__, new_new_n2378__, new_new_n2379__, new_new_n2380__,
    new_new_n2381__, new_new_n2382__, new_new_n2383__, new_new_n2384__,
    new_new_n2385__, new_new_n2386__, new_new_n2387__, new_new_n2388__,
    new_new_n2389__, new_new_n2390__, new_new_n2391__, new_new_n2392__,
    new_new_n2393__, new_new_n2394__, new_new_n2395__, new_new_n2396__,
    new_new_n2397__, new_new_n2398__, new_new_n2399__, new_new_n2400__,
    new_new_n2401__, new_new_n2402__, new_new_n2403__, new_new_n2404__,
    new_new_n2405__, new_new_n2406__, new_new_n2407__, new_new_n2408__,
    new_new_n2409__, new_new_n2410__, new_new_n2411__, new_new_n2412__,
    new_new_n2413__, new_new_n2414__, new_new_n2415__, new_new_n2416__,
    new_new_n2417__, new_new_n2418__, new_new_n2419__, new_new_n2420__,
    new_new_n2421__, new_new_n2422__, new_new_n2423__, new_new_n2424__,
    new_new_n2425__, new_new_n2426__, new_new_n2427__, new_new_n2428__,
    new_new_n2429__, new_new_n2430__, new_new_n2431__, new_new_n2432__,
    new_new_n2433__, new_new_n2434__, new_new_n2435__, new_new_n2436__,
    new_new_n2437__, new_new_n2438__, new_new_n2439__, new_new_n2440__,
    new_new_n2441__, new_new_n2442__, new_new_n2443__, new_new_n2444__,
    n3413, n3416, n3419, n3422, n3425, n3428, n3431, n3434, n3437, n3440,
    n3443, n3446, n3449, n3452, n3455, n3458, n3461, n3464, n3467, n3470,
    n3473, n3476, n3479, n3482, n3485, n3488, n3491, n3494, n3497, n3500,
    n3503, n3506, n3509, n3512, n3515, n3518, n3521, n3524, n3527, n3530,
    n3533, n3536, n3539, n3542, n3545, n3548, n3551, n3554, n3557, n3560,
    n3563, n3566, n3569, n3572, n3575, n3578, n3581, n3584, n3587, n3590,
    n3593, n3596, n3599, n3602, n3605, n3608, n3611, n3614, n3617, n3620,
    n3623, n3626, n3629, n3632, n3635, n3638, n3641, n3644, n3647, n3650,
    n3653, n3656, n3659, n3662, n3665, n3668, n3671, n3674, n3677, n3680,
    n3683, n3686, n3689, n3692, n3695, n3698, n3701, n3704, n3707, n3710,
    n3713, n3716, n3719, n3722, n3725, n3728, n3731, n3734, n3737, n3740,
    n3743, n3746, n3749, n3752, n3755, n3758, n3761, n3764, n3767, n3770,
    n3773, n3776, n3779, n3782, n3785, n3788, n3791, n3794, n3797, n3800,
    n3803, n3806, n3809, n3812, n3815, n3818, n3821, n3824, n3827, n3830,
    n3833, n3836, n3839, n3842, n3845, n3848, n3851, n3854, n3857, n3860,
    n3863, n3866, n3869, n3872, n3875, n3878, n3881, n3884, n3887, n3890,
    n3893, n3896, n3899, n3902, n3905, n3908, n3911, n3914, n3917, n3920,
    n3923, n3926, n3929, n3932, n3935, n3938, n3941, n3944, n3947, n3950,
    n3953, n3956, n3959, n3962, n3965, n3968, n3971, n3974, n3977, n3980,
    n3983, n3986, n3989, n3992, n3995, n3998, n4001, n4004, n4007, n4010,
    n4013, n4016, n4019, n4022, n4025, n4028, n4031, n4034, n4037, n4040,
    n4043, n4046, n4049, n4052, n4055, n4058, n4061, n4064, n4067, n4070,
    n4073, n4076, n4079, n4082, n4085, n4088, n4091, n4094, n4097, n4100,
    n4103, n4106, n4109, n4112, n4115, n4118, n4121, n4124, n4127, n4130,
    n4133, n4136, n4139, n4142, n4145, n4148, n4151, n4154, n4157, n4160,
    n4163, n4166, n4169, n4172, n4175, n4178, n4181, n4184, n4187, n4190,
    n4193, n4196, n4199, n4202, n4205, n4208, n4211, n4214, n4217, n4220,
    n4223, n4226, n4229, n4232, n4235, n4238, n4241, n4244, n4247, n4250,
    n4253, n4256, n4259, n4262, n4265, n4268, n4271, n4274, n4277, n4280,
    n4283, n4286, n4289, n4292, n4295, n4298, n4301, n4304;
  buf1  g0000(.din(G1), .dout(new_new_n683__));
  buf1  g0001(.din(G2), .dout(new_new_n685__));
  buf1  g0002(.din(G3), .dout(new_new_n687__));
  buf1  g0003(.din(G4), .dout(new_new_n689__));
  buf1  g0004(.din(G5), .dout(new_new_n691__));
  buf1  g0005(.din(G6), .dout(new_new_n693__));
  buf1  g0006(.din(G7), .dout(new_new_n695__));
  buf1  g0007(.din(G8), .dout(new_new_n697__));
  buf1  g0008(.din(G9), .dout(new_new_n699__));
  buf1  g0009(.din(G10), .dout(new_new_n701__));
  buf1  g0010(.din(G11), .dout(new_new_n703__));
  buf1  g0011(.din(G12), .dout(new_new_n705__));
  buf1  g0012(.din(G13), .dout(new_new_n707__));
  buf1  g0013(.din(G14), .dout(new_new_n709__));
  buf1  g0014(.din(G15), .dout(new_new_n711__));
  buf1  g0015(.din(G16), .dout(new_new_n713__));
  buf1  g0016(.din(G17), .dout(new_new_n715__));
  buf1  g0017(.din(G18), .dout(new_new_n717__));
  buf1  g0018(.din(G19), .dout(new_new_n719__));
  buf1  g0019(.din(G20), .dout(new_new_n721__));
  buf1  g0020(.din(G21), .dout(new_new_n723__));
  buf1  g0021(.din(G22), .dout(new_new_n725__));
  buf1  g0022(.din(G23), .dout(new_new_n727__));
  buf1  g0023(.din(G24), .dout(new_new_n729__));
  buf1  g0024(.din(G25), .dout(new_new_n731__));
  buf1  g0025(.din(G26), .dout(new_new_n733__));
  buf1  g0026(.din(G27), .dout(new_new_n735__));
  buf1  g0027(.din(G28), .dout(new_new_n737__));
  buf1  g0028(.din(G29), .dout(new_new_n739__));
  buf1  g0029(.din(G30), .dout(new_new_n741__));
  buf1  g0030(.din(G31), .dout(new_new_n743__));
  buf1  g0031(.din(G32), .dout(new_new_n745__));
  buf1  g0032(.din(G33), .dout(new_new_n747__));
  buf1  g0033(.din(G34), .dout(new_new_n749__));
  buf1  g0034(.din(G35), .dout(new_new_n751__));
  buf1  g0035(.din(G36), .dout(new_new_n753__));
  buf1  g0036(.din(G37), .dout(new_new_n755__));
  buf1  g0037(.din(G38), .dout(new_new_n757__));
  buf1  g0038(.din(G39), .dout(new_new_n759__));
  buf1  g0039(.din(G40), .dout(new_new_n761__));
  buf1  g0040(.din(G41), .dout(new_new_n763__));
  buf1  g0041(.din(G42), .dout(new_new_n765__));
  buf1  g0042(.din(G43), .dout(new_new_n767__));
  buf1  g0043(.din(G44), .dout(new_new_n769__));
  buf1  g0044(.din(G45), .dout(new_new_n771__));
  buf1  g0045(.din(G46), .dout(new_new_n773__));
  buf1  g0046(.din(G47), .dout(new_new_n775__));
  buf1  g0047(.din(G48), .dout(new_new_n777__));
  buf1  g0048(.din(G49), .dout(new_new_n779__));
  buf1  g0049(.din(G50), .dout(new_new_n781__));
  buf1  g0050(.din(G51), .dout(new_new_n783__));
  buf1  g0051(.din(G52), .dout(new_new_n785__));
  buf1  g0052(.din(G53), .dout(new_new_n787__));
  buf1  g0053(.din(G54), .dout(new_new_n789__));
  buf1  g0054(.din(G55), .dout(new_new_n791__));
  buf1  g0055(.din(G56), .dout(new_new_n793__));
  buf1  g0056(.din(G57), .dout(new_new_n795__));
  buf1  g0057(.din(G58), .dout(new_new_n797__));
  buf1  g0058(.din(G59), .dout(new_new_n799__));
  buf1  g0059(.din(G60), .dout(new_new_n801__));
  buf1  g0060(.din(n480_lo), .dout(new_new_n803__));
  not1  g0061(.din(n480_lo), .dout(new_new_n804__));
  not1  g0062(.din(n492_lo), .dout(new_new_n806__));
  buf1  g0063(.din(n495_lo), .dout(new_new_n807__));
  buf1  g0064(.din(n498_lo), .dout(new_new_n809__));
  buf1  g0065(.din(n501_lo), .dout(new_new_n811__));
  not1  g0066(.din(n501_lo), .dout(new_new_n812__));
  buf1  g0067(.din(n504_lo), .dout(new_new_n813__));
  not1  g0068(.din(n504_lo), .dout(new_new_n814__));
  buf1  g0069(.din(n516_lo), .dout(new_new_n815__));
  not1  g0070(.din(n516_lo), .dout(new_new_n816__));
  buf1  g0071(.din(n528_lo), .dout(new_new_n817__));
  not1  g0072(.din(n528_lo), .dout(new_new_n818__));
  buf1  g0073(.din(n531_lo), .dout(new_new_n819__));
  not1  g0074(.din(n531_lo), .dout(new_new_n820__));
  not1  g0075(.din(n540_lo), .dout(new_new_n822__));
  buf1  g0076(.din(n543_lo), .dout(new_new_n823__));
  buf1  g0077(.din(n546_lo), .dout(new_new_n825__));
  buf1  g0078(.din(n549_lo), .dout(new_new_n827__));
  not1  g0079(.din(n552_lo), .dout(new_new_n830__));
  not1  g0080(.din(n564_lo), .dout(new_new_n832__));
  buf1  g0081(.din(n579_lo), .dout(new_new_n833__));
  not1  g0082(.din(n579_lo), .dout(new_new_n834__));
  buf1  g0083(.din(n600_lo), .dout(new_new_n835__));
  not1  g0084(.din(n600_lo), .dout(new_new_n836__));
  buf1  g0085(.din(n603_lo), .dout(new_new_n837__));
  buf1  g0086(.din(n606_lo), .dout(new_new_n839__));
  buf1  g0087(.din(n609_lo), .dout(new_new_n841__));
  not1  g0088(.din(n609_lo), .dout(new_new_n842__));
  not1  g0089(.din(n612_lo), .dout(new_new_n844__));
  buf1  g0090(.din(n615_lo), .dout(new_new_n845__));
  buf1  g0091(.din(n618_lo), .dout(new_new_n847__));
  not1  g0092(.din(n621_lo), .dout(new_new_n850__));
  buf1  g0093(.din(n627_lo), .dout(new_new_n851__));
  buf1  g0094(.din(n630_lo), .dout(new_new_n853__));
  not1  g0095(.din(n633_lo), .dout(new_new_n856__));
  buf1  g0096(.din(n639_lo), .dout(new_new_n857__));
  buf1  g0097(.din(n642_lo), .dout(new_new_n859__));
  buf1  g0098(.din(n645_lo), .dout(new_new_n861__));
  not1  g0099(.din(n648_lo), .dout(new_new_n864__));
  buf1  g0100(.din(n660_lo), .dout(new_new_n865__));
  not1  g0101(.din(n660_lo), .dout(new_new_n866__));
  buf1  g0102(.din(n663_lo), .dout(new_new_n867__));
  not1  g0103(.din(n663_lo), .dout(new_new_n868__));
  buf1  g0104(.din(n672_lo), .dout(new_new_n869__));
  not1  g0105(.din(n672_lo), .dout(new_new_n870__));
  buf1  g0106(.din(n675_lo), .dout(new_new_n871__));
  buf1  g0107(.din(n678_lo), .dout(new_new_n873__));
  buf1  g0108(.din(n681_lo), .dout(new_new_n875__));
  not1  g0109(.din(n684_lo), .dout(new_new_n878__));
  buf1  g0110(.din(n687_lo), .dout(new_new_n879__));
  buf1  g0111(.din(n690_lo), .dout(new_new_n881__));
  buf1  g0112(.din(n693_lo), .dout(new_new_n883__));
  not1  g0113(.din(n696_lo), .dout(new_new_n886__));
  buf1  g0114(.din(n699_lo), .dout(new_new_n887__));
  buf1  g0115(.din(n702_lo), .dout(new_new_n889__));
  buf1  g0116(.din(n705_lo), .dout(new_new_n891__));
  buf1  g0117(.din(n708_lo), .dout(new_new_n893__));
  buf1  g0118(.din(n711_lo), .dout(new_new_n895__));
  buf1  g0119(.din(n714_lo), .dout(new_new_n897__));
  buf1  g0120(.din(n717_lo), .dout(new_new_n899__));
  buf1  g0121(.din(n720_lo), .dout(new_new_n901__));
  buf1  g0122(.din(n723_lo), .dout(new_new_n903__));
  buf1  g0123(.din(n726_lo), .dout(new_new_n905__));
  buf1  g0124(.din(n729_lo), .dout(new_new_n907__));
  buf1  g0125(.din(n732_lo), .dout(new_new_n909__));
  buf1  g0126(.din(n735_lo), .dout(new_new_n911__));
  buf1  g0127(.din(n738_lo), .dout(new_new_n913__));
  buf1  g0128(.din(n741_lo), .dout(new_new_n915__));
  buf1  g0129(.din(n744_lo), .dout(new_new_n917__));
  buf1  g0130(.din(n747_lo), .dout(new_new_n919__));
  buf1  g0131(.din(n750_lo), .dout(new_new_n921__));
  not1  g0132(.din(n756_lo), .dout(new_new_n924__));
  buf1  g0133(.din(n759_lo), .dout(new_new_n925__));
  buf1  g0134(.din(n762_lo), .dout(new_new_n927__));
  not1  g0135(.din(n762_lo), .dout(new_new_n928__));
  not1  g0136(.din(n768_lo), .dout(new_new_n930__));
  buf1  g0137(.din(n771_lo), .dout(new_new_n931__));
  buf1  g0138(.din(n774_lo), .dout(new_new_n933__));
  not1  g0139(.din(n774_lo), .dout(new_new_n934__));
  not1  g0140(.din(n780_lo), .dout(new_new_n936__));
  buf1  g0141(.din(n783_lo), .dout(new_new_n937__));
  buf1  g0142(.din(n786_lo), .dout(new_new_n939__));
  not1  g0143(.din(n786_lo), .dout(new_new_n940__));
  not1  g0144(.din(n792_lo), .dout(new_new_n942__));
  buf1  g0145(.din(n795_lo), .dout(new_new_n943__));
  not1  g0146(.din(n804_lo), .dout(new_new_n946__));
  buf1  g0147(.din(n807_lo), .dout(new_new_n947__));
  not1  g0148(.din(n816_lo), .dout(new_new_n950__));
  buf1  g0149(.din(n819_lo), .dout(new_new_n951__));
  not1  g0150(.din(n828_lo), .dout(new_new_n954__));
  buf1  g0151(.din(n831_lo), .dout(new_new_n955__));
  buf1  g0152(.din(n843_lo), .dout(new_new_n957__));
  buf1  g0153(.din(n846_lo), .dout(new_new_n959__));
  buf1  g0154(.din(n849_lo), .dout(new_new_n961__));
  buf1  g0155(.din(n852_lo), .dout(new_new_n963__));
  not1  g0156(.din(n852_lo), .dout(new_new_n964__));
  buf1  g0157(.din(n855_lo), .dout(new_new_n965__));
  buf1  g0158(.din(n858_lo), .dout(new_new_n967__));
  buf1  g0159(.din(n861_lo), .dout(new_new_n969__));
  buf1  g0160(.din(n864_lo), .dout(new_new_n971__));
  not1  g0161(.din(n864_lo), .dout(new_new_n972__));
  buf1  g0162(.din(n867_lo), .dout(new_new_n973__));
  buf1  g0163(.din(n870_lo), .dout(new_new_n975__));
  not1  g0164(.din(n870_lo), .dout(new_new_n976__));
  buf1  g0165(.din(n879_lo), .dout(new_new_n977__));
  buf1  g0166(.din(n891_lo), .dout(new_new_n979__));
  buf1  g0167(.din(n903_lo), .dout(new_new_n981__));
  buf1  g0168(.din(n915_lo), .dout(new_new_n983__));
  not1  g0169(.din(n918_lo), .dout(new_new_n986__));
  buf1  g0170(.din(n927_lo), .dout(new_new_n987__));
  buf1  g0171(.din(n951_lo), .dout(new_new_n989__));
  buf1  g0172(.din(n954_lo), .dout(new_new_n991__));
  buf1  g0173(.din(n957_lo), .dout(new_new_n993__));
  not1  g0174(.din(n957_lo), .dout(new_new_n994__));
  not1  g0175(.din(n960_lo), .dout(new_new_n996__));
  buf1  g0176(.din(n963_lo), .dout(new_new_n997__));
  buf1  g0177(.din(n966_lo), .dout(new_new_n999__));
  not1  g0178(.din(n972_lo), .dout(new_new_n1002__));
  buf1  g0179(.din(n975_lo), .dout(new_new_n1003__));
  buf1  g0180(.din(n978_lo), .dout(new_new_n1005__));
  not1  g0181(.din(n984_lo), .dout(new_new_n1008__));
  buf1  g0182(.din(n987_lo), .dout(new_new_n1009__));
  buf1  g0183(.din(n990_lo), .dout(new_new_n1011__));
  not1  g0184(.din(n996_lo), .dout(new_new_n1014__));
  buf1  g0185(.din(n999_lo), .dout(new_new_n1015__));
  buf1  g0186(.din(n1002_lo), .dout(new_new_n1017__));
  not1  g0187(.din(n1002_lo), .dout(new_new_n1018__));
  not1  g0188(.din(n1008_lo), .dout(new_new_n1020__));
  buf1  g0189(.din(n1011_lo), .dout(new_new_n1021__));
  buf1  g0190(.din(n1014_lo), .dout(new_new_n1023__));
  not1  g0191(.din(n1014_lo), .dout(new_new_n1024__));
  not1  g0192(.din(n1020_lo), .dout(new_new_n1026__));
  buf1  g0193(.din(n1023_lo), .dout(new_new_n1027__));
  buf1  g0194(.din(n1026_lo), .dout(new_new_n1029__));
  not1  g0195(.din(n1026_lo), .dout(new_new_n1030__));
  not1  g0196(.din(n1032_lo), .dout(new_new_n1032__));
  buf1  g0197(.din(n1035_lo), .dout(new_new_n1033__));
  buf1  g0198(.din(n1038_lo), .dout(new_new_n1035__));
  not1  g0199(.din(n1038_lo), .dout(new_new_n1036__));
  not1  g0200(.din(n1044_lo), .dout(new_new_n1038__));
  buf1  g0201(.din(n1047_lo), .dout(new_new_n1039__));
  buf1  g0202(.din(n1050_lo), .dout(new_new_n1041__));
  buf1  g0203(.din(n1053_lo), .dout(new_new_n1043__));
  buf1  g0204(.din(n1056_lo), .dout(new_new_n1045__));
  not1  g0205(.din(n1056_lo), .dout(new_new_n1046__));
  buf1  g0206(.din(n1059_lo), .dout(new_new_n1047__));
  buf1  g0207(.din(n1062_lo), .dout(new_new_n1049__));
  buf1  g0208(.din(n1065_lo), .dout(new_new_n1051__));
  not1  g0209(.din(n1068_lo), .dout(new_new_n1054__));
  buf1  g0210(.din(n1071_lo), .dout(new_new_n1055__));
  buf1  g0211(.din(n1074_lo), .dout(new_new_n1057__));
  buf1  g0212(.din(n1077_lo), .dout(new_new_n1059__));
  not1  g0213(.din(n1080_lo), .dout(new_new_n1062__));
  buf1  g0214(.din(n1083_lo), .dout(new_new_n1063__));
  buf1  g0215(.din(n1086_lo), .dout(new_new_n1065__));
  buf1  g0216(.din(n1089_lo), .dout(new_new_n1067__));
  not1  g0217(.din(n1092_lo), .dout(new_new_n1070__));
  buf1  g0218(.din(n1095_lo), .dout(new_new_n1071__));
  buf1  g0219(.din(n1098_lo), .dout(new_new_n1073__));
  buf1  g0220(.din(n1101_lo), .dout(new_new_n1075__));
  not1  g0221(.din(n1104_lo), .dout(new_new_n1078__));
  buf1  g0222(.din(n1107_lo), .dout(new_new_n1079__));
  buf1  g0223(.din(n1110_lo), .dout(new_new_n1081__));
  buf1  g0224(.din(n1113_lo), .dout(new_new_n1083__));
  not1  g0225(.din(n1116_lo), .dout(new_new_n1086__));
  buf1  g0226(.din(n1119_lo), .dout(new_new_n1087__));
  buf1  g0227(.din(n1122_lo), .dout(new_new_n1089__));
  buf1  g0228(.din(n1125_lo), .dout(new_new_n1091__));
  not1  g0229(.din(n1128_lo), .dout(new_new_n1094__));
  buf1  g0230(.din(n1131_lo), .dout(new_new_n1095__));
  buf1  g0231(.din(n1134_lo), .dout(new_new_n1097__));
  buf1  g0232(.din(n1137_lo), .dout(new_new_n1099__));
  not1  g0233(.din(n1140_lo), .dout(new_new_n1102__));
  buf1  g0234(.din(n1143_lo), .dout(new_new_n1103__));
  buf1  g0235(.din(n1146_lo), .dout(new_new_n1105__));
  buf1  g0236(.din(n1149_lo), .dout(new_new_n1107__));
  not1  g0237(.din(n1152_lo), .dout(new_new_n1110__));
  buf1  g0238(.din(n1155_lo), .dout(new_new_n1111__));
  buf1  g0239(.din(n1158_lo), .dout(new_new_n1113__));
  not1  g0240(.din(n1158_lo), .dout(new_new_n1114__));
  buf1  g0241(.din(n1167_lo), .dout(new_new_n1115__));
  buf1  g0242(.din(n1170_lo), .dout(new_new_n1117__));
  buf1  g0243(.din(n1173_lo), .dout(new_new_n1119__));
  not1  g0244(.din(n1176_lo), .dout(new_new_n1122__));
  buf1  g0245(.din(n1179_lo), .dout(new_new_n1123__));
  not1  g0246(.din(n1529_o2), .dout(new_new_n1126__));
  not1  g0247(.din(n1616_o2), .dout(new_new_n1128__));
  not1  g0248(.din(n1655_o2), .dout(new_new_n1130__));
  not1  g0249(.din(n1656_o2), .dout(new_new_n1132__));
  not1  g0250(.din(n1657_o2), .dout(new_new_n1134__));
  not1  g0251(.din(n1730_o2), .dout(new_new_n1136__));
  not1  g0252(.din(n1731_o2), .dout(new_new_n1138__));
  not1  g0253(.din(n1732_o2), .dout(new_new_n1140__));
  not1  g0254(.din(n1729_o2), .dout(new_new_n1142__));
  not1  g0255(.din(n1805_o2), .dout(new_new_n1144__));
  not1  g0256(.din(n1808_o2), .dout(new_new_n1146__));
  not1  g0257(.din(n1807_o2), .dout(new_new_n1148__));
  not1  g0258(.din(n1809_o2), .dout(new_new_n1150__));
  buf1  g0259(.din(n1663_o2), .dout(new_new_n1151__));
  not1  g0260(.din(n1663_o2), .dout(new_new_n1152__));
  buf1  g0261(.din(n1664_o2), .dout(new_new_n1153__));
  buf1  g0262(.din(n1704_o2), .dout(new_new_n1155__));
  not1  g0263(.din(n1704_o2), .dout(new_new_n1156__));
  buf1  g0264(.din(n1705_o2), .dout(new_new_n1157__));
  buf1  g0265(.din(n1706_o2), .dout(new_new_n1159__));
  not1  g0266(.din(n1706_o2), .dout(new_new_n1160__));
  buf1  g0267(.din(n1707_o2), .dout(new_new_n1161__));
  not1  g0268(.din(n1707_o2), .dout(new_new_n1162__));
  buf1  g0269(.din(n1708_o2), .dout(new_new_n1163__));
  buf1  g0270(.din(n1709_o2), .dout(new_new_n1165__));
  not1  g0271(.din(G280_o2), .dout(new_new_n1168__));
  not1  g0272(.din(G655_o2), .dout(new_new_n1170__));
  not1  g0273(.din(G663_o2), .dout(new_new_n1172__));
  not1  g0274(.din(G672_o2), .dout(new_new_n1174__));
  not1  g0275(.din(G538_o2), .dout(new_new_n1176__));
  buf1  g0276(.din(n1780_o2), .dout(new_new_n1177__));
  buf1  g0277(.din(n1781_o2), .dout(new_new_n1179__));
  not1  g0278(.din(n1797_o2), .dout(new_new_n1182__));
  buf1  g0279(.din(n1798_o2), .dout(new_new_n1183__));
  not1  g0280(.din(n1798_o2), .dout(new_new_n1184__));
  buf1  g0281(.din(n1799_o2), .dout(new_new_n1185__));
  not1  g0282(.din(n1799_o2), .dout(new_new_n1186__));
  buf1  g0283(.din(n1800_o2), .dout(new_new_n1187__));
  not1  g0284(.din(n1800_o2), .dout(new_new_n1188__));
  not1  g0285(.din(G578_o2), .dout(new_new_n1190__));
  buf1  g0286(.din(n1828_o2), .dout(new_new_n1191__));
  buf1  g0287(.din(n801_lo_buf_o2), .dout(new_new_n1193__));
  not1  g0288(.din(n801_lo_buf_o2), .dout(new_new_n1194__));
  not1  g0289(.din(G693_o2), .dout(new_new_n1196__));
  not1  g0290(.din(G702_o2), .dout(new_new_n1198__));
  not1  g0291(.din(G712_o2), .dout(new_new_n1200__));
  not1  g0292(.din(G685_o2), .dout(new_new_n1202__));
  not1  g0293(.din(G658_o2), .dout(new_new_n1204__));
  not1  g0294(.din(G667_o2), .dout(new_new_n1206__));
  not1  g0295(.din(G677_o2), .dout(new_new_n1208__));
  not1  g0296(.din(G650_o2), .dout(new_new_n1210__));
  not1  g0297(.din(G798_o2), .dout(new_new_n1212__));
  buf1  g0298(.din(n1017_lo_buf_o2), .dout(new_new_n1213__));
  not1  g0299(.din(n1017_lo_buf_o2), .dout(new_new_n1214__));
  buf1  g0300(.din(n1029_lo_buf_o2), .dout(new_new_n1215__));
  not1  g0301(.din(n1029_lo_buf_o2), .dout(new_new_n1216__));
  buf1  g0302(.din(n1041_lo_buf_o2), .dout(new_new_n1217__));
  not1  g0303(.din(n1041_lo_buf_o2), .dout(new_new_n1218__));
  buf1  g0304(.din(G558_o2), .dout(new_new_n1219__));
  buf1  g0305(.din(G562_o2), .dout(new_new_n1221__));
  buf1  g0306(.din(G566_o2), .dout(new_new_n1223__));
  buf1  g0307(.din(n1835_o2), .dout(new_new_n1225__));
  buf1  g0308(.din(n1836_o2), .dout(new_new_n1227__));
  not1  g0309(.din(n1837_o2), .dout(new_new_n1230__));
  buf1  g0310(.din(n765_lo_buf_o2), .dout(new_new_n1231__));
  not1  g0311(.din(n765_lo_buf_o2), .dout(new_new_n1232__));
  buf1  g0312(.din(n777_lo_buf_o2), .dout(new_new_n1233__));
  not1  g0313(.din(n777_lo_buf_o2), .dout(new_new_n1234__));
  buf1  g0314(.din(n789_lo_buf_o2), .dout(new_new_n1235__));
  not1  g0315(.din(n789_lo_buf_o2), .dout(new_new_n1236__));
  buf1  g0316(.din(G617_o2), .dout(new_new_n1237__));
  not1  g0317(.din(G617_o2), .dout(new_new_n1238__));
  buf1  g0318(.din(G626_o2), .dout(new_new_n1239__));
  not1  g0319(.din(G626_o2), .dout(new_new_n1240__));
  buf1  g0320(.din(G636_o2), .dout(new_new_n1241__));
  not1  g0321(.din(G636_o2), .dout(new_new_n1242__));
  buf1  g0322(.din(n489_lo_buf_o2), .dout(new_new_n1243__));
  buf1  g0323(.din(n513_lo_buf_o2), .dout(new_new_n1245__));
  not1  g0324(.din(n513_lo_buf_o2), .dout(new_new_n1246__));
  buf1  g0325(.din(n561_lo_buf_o2), .dout(new_new_n1247__));
  buf1  g0326(.din(n597_lo_buf_o2), .dout(new_new_n1249__));
  buf1  g0327(.din(n657_lo_buf_o2), .dout(new_new_n1251__));
  buf1  g0328(.din(G276_o2), .dout(new_new_n1253__));
  buf1  g0329(.din(n1005_lo_buf_o2), .dout(new_new_n1255__));
  not1  g0330(.din(n1005_lo_buf_o2), .dout(new_new_n1256__));
  buf1  g0331(.din(n1161_lo_buf_o2), .dout(new_new_n1257__));
  not1  g0332(.din(n1161_lo_buf_o2), .dout(new_new_n1258__));
  buf1  g0333(.din(G620_o2), .dout(new_new_n1259__));
  not1  g0334(.din(G620_o2), .dout(new_new_n1260__));
  buf1  g0335(.din(G629_o2), .dout(new_new_n1261__));
  not1  g0336(.din(G629_o2), .dout(new_new_n1262__));
  buf1  g0337(.din(G639_o2), .dout(new_new_n1263__));
  not1  g0338(.din(G639_o2), .dout(new_new_n1264__));
  buf1  g0339(.din(G554_o2), .dout(new_new_n1265__));
  buf1  g0340(.din(G690_o2), .dout(new_new_n1267__));
  buf1  g0341(.din(G698_o2), .dout(new_new_n1269__));
  not1  g0342(.din(G698_o2), .dout(new_new_n1270__));
  buf1  g0343(.din(G707_o2), .dout(new_new_n1271__));
  not1  g0344(.din(G707_o2), .dout(new_new_n1272__));
  buf1  g0345(.din(G319_o2), .dout(new_new_n1273__));
  not1  g0346(.din(G389_o2), .dout(new_new_n1276__));
  buf1  g0347(.din(n753_lo_buf_o2), .dout(new_new_n1277__));
  not1  g0348(.din(n753_lo_buf_o2), .dout(new_new_n1278__));
  not1  g0349(.din(G647_o2), .dout(new_new_n1280__));
  not1  g0350(.din(G769_o2), .dout(new_new_n1282__));
  not1  g0351(.din(G785_o2), .dout(new_new_n1284__));
  not1  g0352(.din(G808_o2), .dout(new_new_n1286__));
  buf1  g0353(.din(G445_o2), .dout(new_new_n1287__));
  not1  g0354(.din(G445_o2), .dout(new_new_n1288__));
  buf1  g0355(.din(G448_o2), .dout(new_new_n1289__));
  not1  g0356(.din(G448_o2), .dout(new_new_n1290__));
  buf1  g0357(.din(G477_o2), .dout(new_new_n1291__));
  not1  g0358(.din(G477_o2), .dout(new_new_n1292__));
  buf1  g0359(.din(G480_o2), .dout(new_new_n1293__));
  not1  g0360(.din(G480_o2), .dout(new_new_n1294__));
  not1  g0361(.din(G436_o2), .dout(new_new_n1296__));
  not1  g0362(.din(G786_o2), .dout(new_new_n1298__));
  not1  g0363(.din(G787_o2), .dout(new_new_n1300__));
  not1  g0364(.din(G826_o2), .dout(new_new_n1302__));
  not1  g0365(.din(G827_o2), .dout(new_new_n1304__));
  not1  g0366(.din(G825_o2), .dout(new_new_n1306__));
  buf1  g0367(.din(G610_o2), .dout(new_new_n1307__));
  not1  g0368(.din(G610_o2), .dout(new_new_n1308__));
  buf1  g0369(.din(n537_lo_buf_o2), .dout(new_new_n1309__));
  buf1  g0370(.din(n669_lo_buf_o2), .dout(new_new_n1311__));
  buf1  g0371(.din(n969_lo_buf_o2), .dout(new_new_n1313__));
  not1  g0372(.din(n969_lo_buf_o2), .dout(new_new_n1314__));
  buf1  g0373(.din(n981_lo_buf_o2), .dout(new_new_n1315__));
  not1  g0374(.din(n981_lo_buf_o2), .dout(new_new_n1316__));
  buf1  g0375(.din(n993_lo_buf_o2), .dout(new_new_n1317__));
  not1  g0376(.din(n993_lo_buf_o2), .dout(new_new_n1318__));
  buf1  g0377(.din(G309_o2), .dout(new_new_n1319__));
  not1  g0378(.din(G309_o2), .dout(new_new_n1320__));
  buf1  g0379(.din(G461_o2), .dout(new_new_n1321__));
  not1  g0380(.din(G461_o2), .dout(new_new_n1322__));
  buf1  g0381(.din(G487_o2), .dout(new_new_n1323__));
  not1  g0382(.din(G487_o2), .dout(new_new_n1324__));
  buf1  g0383(.din(G460_o2), .dout(new_new_n1325__));
  not1  g0384(.din(G460_o2), .dout(new_new_n1326__));
  buf1  g0385(.din(G468_o2), .dout(new_new_n1327__));
  not1  g0386(.din(G287_o2), .dout(new_new_n1330__));
  buf1  g0387(.din(G613_o2), .dout(new_new_n1331__));
  not1  g0388(.din(G613_o2), .dout(new_new_n1332__));
  buf1  g0389(.din(n585_lo_buf_o2), .dout(new_new_n1333__));
  not1  g0390(.din(n585_lo_buf_o2), .dout(new_new_n1334__));
  buf1  g0391(.din(n813_lo_buf_o2), .dout(new_new_n1335__));
  buf1  g0392(.din(n825_lo_buf_o2), .dout(new_new_n1337__));
  buf1  g0393(.din(n837_lo_buf_o2), .dout(new_new_n1339__));
  not1  g0394(.din(n897_lo_buf_o2), .dout(new_new_n1342__));
  not1  g0395(.din(n909_lo_buf_o2), .dout(new_new_n1344__));
  not1  g0396(.din(n933_lo_buf_o2), .dout(new_new_n1346__));
  buf1  g0397(.din(G451_o2), .dout(new_new_n1347__));
  not1  g0398(.din(G451_o2), .dout(new_new_n1348__));
  buf1  g0399(.din(G682_o2), .dout(new_new_n1349__));
  not1  g0400(.din(G682_o2), .dout(new_new_n1350__));
  buf1  g0401(.din(G756_o2), .dout(new_new_n1351__));
  not1  g0402(.din(G756_o2), .dout(new_new_n1352__));
  buf1  g0403(.din(G542_o2), .dout(new_new_n1353__));
  not1  g0404(.din(G542_o2), .dout(new_new_n1354__));
  buf1  g0405(.din(G546_o2), .dout(new_new_n1355__));
  not1  g0406(.din(G546_o2), .dout(new_new_n1356__));
  buf1  g0407(.din(G550_o2), .dout(new_new_n1357__));
  not1  g0408(.din(G550_o2), .dout(new_new_n1358__));
  buf1  g0409(.din(G310_o2), .dout(new_new_n1359__));
  buf1  g0410(.din(n798_lo_buf_o2), .dout(new_new_n1361__));
  not1  g0411(.din(n798_lo_buf_o2), .dout(new_new_n1362__));
  not1  g0412(.din(n882_lo_buf_o2), .dout(new_new_n1364__));
  not1  g0413(.din(G427_o2), .dout(new_new_n1366__));
  not1  g0414(.din(G497_o2), .dout(new_new_n1368__));
  not1  g0415(.din(G499_o2), .dout(new_new_n1370__));
  not1  g0416(.din(G501_o2), .dout(new_new_n1372__));
  not1  g0417(.din(G498_o2), .dout(new_new_n1374__));
  not1  g0418(.din(G500_o2), .dout(new_new_n1376__));
  not1  g0419(.din(G502_o2), .dout(new_new_n1378__));
  buf1  g0420(.din(G369_o2), .dout(new_new_n1379__));
  buf1  g0421(.din(n939_lo_buf_o2), .dout(new_new_n1381__));
  not1  g0422(.din(n939_lo_buf_o2), .dout(new_new_n1382__));
  buf1  g0423(.din(n486_lo_buf_o2), .dout(new_new_n1383__));
  buf1  g0424(.din(n510_lo_buf_o2), .dout(new_new_n1385__));
  not1  g0425(.din(n510_lo_buf_o2), .dout(new_new_n1386__));
  buf1  g0426(.din(n558_lo_buf_o2), .dout(new_new_n1387__));
  not1  g0427(.din(n558_lo_buf_o2), .dout(new_new_n1388__));
  buf1  g0428(.din(n594_lo_buf_o2), .dout(new_new_n1389__));
  not1  g0429(.din(n594_lo_buf_o2), .dout(new_new_n1390__));
  buf1  g0430(.din(n654_lo_buf_o2), .dout(new_new_n1391__));
  not1  g0431(.din(n654_lo_buf_o2), .dout(new_new_n1392__));
  buf1  g0432(.din(n477_lo_buf_o2), .dout(new_new_n1393__));
  not1  g0433(.din(n477_lo_buf_o2), .dout(new_new_n1394__));
  buf1  g0434(.din(n525_lo_buf_o2), .dout(new_new_n1395__));
  not1  g0435(.din(n525_lo_buf_o2), .dout(new_new_n1396__));
  buf1  g0436(.din(n573_lo_buf_o2), .dout(new_new_n1397__));
  not1  g0437(.din(n573_lo_buf_o2), .dout(new_new_n1398__));
  or1   g0438(.dina(new_new_n866__), .dinb(new_new_n2142__), .dout(new_new_n1399__));
  or1   g0439(.dina(new_new_n1399__), .dinb(new_new_n2144__), .dout(new_new_n1400__));
  or1   g0440(.dina(new_new_n2145__), .dinb(new_new_n2142__), .dout(new_new_n1401__));
  or1   g0441(.dina(new_new_n2146__), .dinb(new_new_n2147__), .dout(new_new_n1402__));
  or1   g0442(.dina(new_new_n2146__), .dinb(new_new_n2144__), .dout(new_new_n1403__));
  or1   g0443(.dina(new_new_n886__), .dinb(new_new_n878__), .dout(new_new_n1404__));
  or1   g0444(.dina(new_new_n806__), .dinb(new_new_n2148__), .dout(new_new_n1405__));
  or1   g0445(.dina(new_new_n1405__), .dinb(new_new_n2149__), .dout(new_new_n1406__));
  or1   g0446(.dina(new_new_n1406__), .dinb(new_new_n2150__), .dout(new_new_n1407__));
  and1  g0447(.dina(new_new_n817__), .dinb(new_new_n803__), .dout(new_new_n1408__));
  or1   g0448(.dina(new_new_n818__), .dinb(new_new_n2148__), .dout(new_new_n1409__));
  and1  g0449(.dina(new_new_n1408__), .dinb(new_new_n813__), .dout(new_new_n1410__));
  or1   g0450(.dina(new_new_n1409__), .dinb(new_new_n2149__), .dout(new_new_n1411__));
  and1  g0451(.dina(new_new_n1410__), .dinb(new_new_n815__), .dout(new_new_n1412__));
  or1   g0452(.dina(new_new_n1411__), .dinb(new_new_n2150__), .dout(new_new_n1413__));
  and1  g0453(.dina(new_new_n1412__), .dinb(new_new_n2152__), .dout(new_new_n1414__));
  and1  g0454(.dina(new_new_n865__), .dinb(new_new_n835__), .dout(new_new_n1415__));
  and1  g0455(.dina(new_new_n1415__), .dinb(new_new_n869__), .dout(new_new_n1416__));
  or1   g0456(.dina(new_new_n2153__), .dinb(new_new_n2145__), .dout(new_new_n1417__));
  or1   g0457(.dina(new_new_n2154__), .dinb(new_new_n2147__), .dout(new_new_n1418__));
  or1   g0458(.dina(new_new_n2154__), .dinb(new_new_n2143__), .dout(new_new_n1419__));
  or1   g0459(.dina(new_new_n901__), .dinb(new_new_n893__), .dout(new_new_n1420__));
  and1  g0460(.dina(new_new_n2155__), .dinb(new_new_n917__), .dout(new_new_n1421__));
  or1   g0461(.dina(new_new_n1413__), .dinb(new_new_n2152__), .dout(new_new_n1422__));
  or1   g0462(.dina(new_new_n2156__), .dinb(new_new_n2141__), .dout(new_new_n1423__));
  or1   g0463(.dina(new_new_n1423__), .dinb(new_new_n2157__), .dout(new_new_n1424__));
  or1   g0464(.dina(new_new_n2156__), .dinb(new_new_n2153__), .dout(new_new_n1425__));
  or1   g0465(.dina(new_new_n1425__), .dinb(new_new_n864__), .dout(new_new_n1426__));
  or1   g0466(.dina(new_new_n1426__), .dinb(new_new_n2157__), .dout(new_new_n1427__));
  and1  g0467(.dina(new_new_n2155__), .dinb(new_new_n909__), .dout(new_new_n1428__));
  and1  g0468(.dina(new_new_n2158__), .dinb(new_new_n2160__), .dout(new_new_n1429__));
  or1   g0469(.dina(new_new_n2162__), .dinb(new_new_n2164__), .dout(new_new_n1430__));
  and1  g0470(.dina(new_new_n2162__), .dinb(new_new_n2164__), .dout(new_new_n1431__));
  or1   g0471(.dina(new_new_n2158__), .dinb(new_new_n2160__), .dout(new_new_n1432__));
  and1  g0472(.dina(new_new_n1432__), .dinb(new_new_n1430__), .dout(new_new_n1433__));
  or1   g0473(.dina(new_new_n1431__), .dinb(new_new_n1429__), .dout(new_new_n1434__));
  and1  g0474(.dina(new_new_n2166__), .dinb(new_new_n2167__), .dout(new_new_n1435__));
  or1   g0475(.dina(new_new_n2168__), .dinb(new_new_n2169__), .dout(new_new_n1436__));
  and1  g0476(.dina(new_new_n2168__), .dinb(new_new_n2169__), .dout(new_new_n1437__));
  or1   g0477(.dina(new_new_n2166__), .dinb(new_new_n2167__), .dout(new_new_n1438__));
  and1  g0478(.dina(new_new_n1438__), .dinb(new_new_n1436__), .dout(new_new_n1439__));
  or1   g0479(.dina(new_new_n1437__), .dinb(new_new_n1435__), .dout(new_new_n1440__));
  and1  g0480(.dina(new_new_n1440__), .dinb(new_new_n1434__), .dout(new_new_n1441__));
  and1  g0481(.dina(new_new_n1439__), .dinb(new_new_n1433__), .dout(new_new_n1442__));
  or1   g0482(.dina(new_new_n1442__), .dinb(new_new_n1441__), .dout(new_new_n1443__));
  and1  g0483(.dina(new_new_n2170__), .dinb(new_new_n2161__), .dout(new_new_n1444__));
  or1   g0484(.dina(new_new_n2171__), .dinb(new_new_n2165__), .dout(new_new_n1445__));
  and1  g0485(.dina(new_new_n2171__), .dinb(new_new_n2165__), .dout(new_new_n1446__));
  or1   g0486(.dina(new_new_n2170__), .dinb(new_new_n2161__), .dout(new_new_n1447__));
  and1  g0487(.dina(new_new_n1447__), .dinb(new_new_n1445__), .dout(new_new_n1448__));
  or1   g0488(.dina(new_new_n1446__), .dinb(new_new_n1444__), .dout(new_new_n1449__));
  and1  g0489(.dina(new_new_n2172__), .dinb(new_new_n2173__), .dout(new_new_n1450__));
  or1   g0490(.dina(new_new_n2174__), .dinb(new_new_n2175__), .dout(new_new_n1451__));
  and1  g0491(.dina(new_new_n2174__), .dinb(new_new_n2175__), .dout(new_new_n1452__));
  or1   g0492(.dina(new_new_n2172__), .dinb(new_new_n2173__), .dout(new_new_n1453__));
  and1  g0493(.dina(new_new_n1453__), .dinb(new_new_n1451__), .dout(new_new_n1454__));
  or1   g0494(.dina(new_new_n1452__), .dinb(new_new_n1450__), .dout(new_new_n1455__));
  and1  g0495(.dina(new_new_n1455__), .dinb(new_new_n1449__), .dout(new_new_n1456__));
  and1  g0496(.dina(new_new_n1454__), .dinb(new_new_n1448__), .dout(new_new_n1457__));
  or1   g0497(.dina(new_new_n1457__), .dinb(new_new_n1456__), .dout(new_new_n1458__));
  or1   g0498(.dina(new_new_n2178__), .dinb(new_new_n954__), .dout(new_new_n1459__));
  or1   g0499(.dina(new_new_n1282__), .dinb(new_new_n2185__), .dout(new_new_n1460__));
  and1  g0500(.dina(new_new_n1460__), .dinb(new_new_n1459__), .dout(new_new_n1461__));
  or1   g0501(.dina(new_new_n1200__), .dinb(new_new_n2192__), .dout(new_new_n1462__));
  or1   g0502(.dina(new_new_n1140__), .dinb(new_new_n2199__), .dout(new_new_n1463__));
  and1  g0503(.dina(new_new_n1463__), .dinb(new_new_n1462__), .dout(new_new_n1464__));
  or1   g0504(.dina(new_new_n1122__), .dinb(new_new_n2205__), .dout(new_new_n1465__));
  or1   g0505(.dina(new_new_n1134__), .dinb(new_new_n2208__), .dout(new_new_n1466__));
  and1  g0506(.dina(new_new_n1466__), .dinb(new_new_n1465__), .dout(new_new_n1467__));
  or1   g0507(.dina(new_new_n2215__), .dinb(new_new_n1038__), .dout(new_new_n1468__));
  and1  g0508(.dina(new_new_n1464__), .dinb(new_new_n1461__), .dout(new_new_n1469__));
  and1  g0509(.dina(new_new_n1469__), .dinb(new_new_n1467__), .dout(new_new_n1470__));
  and1  g0510(.dina(new_new_n1470__), .dinb(new_new_n1468__), .dout(new_new_n1471__));
  or1   g0511(.dina(new_new_n2178__), .dinb(new_new_n942__), .dout(new_new_n1472__));
  or1   g0512(.dina(new_new_n1284__), .dinb(new_new_n2185__), .dout(new_new_n1473__));
  and1  g0513(.dina(new_new_n1473__), .dinb(new_new_n1472__), .dout(new_new_n1474__));
  or1   g0514(.dina(new_new_n1202__), .dinb(new_new_n2192__), .dout(new_new_n1475__));
  or1   g0515(.dina(new_new_n1144__), .dinb(new_new_n2199__), .dout(new_new_n1476__));
  and1  g0516(.dina(new_new_n1476__), .dinb(new_new_n1475__), .dout(new_new_n1477__));
  or1   g0517(.dina(new_new_n1142__), .dinb(new_new_n2208__), .dout(new_new_n1478__));
  or1   g0518(.dina(new_new_n2215__), .dinb(new_new_n1020__), .dout(new_new_n1479__));
  and1  g0519(.dina(new_new_n1479__), .dinb(new_new_n1478__), .dout(new_new_n1480__));
  and1  g0520(.dina(new_new_n1477__), .dinb(new_new_n1474__), .dout(new_new_n1481__));
  and1  g0521(.dina(new_new_n1481__), .dinb(new_new_n1480__), .dout(new_new_n1482__));
  or1   g0522(.dina(new_new_n2179__), .dinb(new_new_n946__), .dout(new_new_n1483__));
  or1   g0523(.dina(new_new_n1298__), .dinb(new_new_n2186__), .dout(new_new_n1484__));
  and1  g0524(.dina(new_new_n1484__), .dinb(new_new_n1483__), .dout(new_new_n1485__));
  or1   g0525(.dina(new_new_n1196__), .dinb(new_new_n2193__), .dout(new_new_n1486__));
  or1   g0526(.dina(new_new_n1136__), .dinb(new_new_n2200__), .dout(new_new_n1487__));
  and1  g0527(.dina(new_new_n1487__), .dinb(new_new_n1486__), .dout(new_new_n1488__));
  or1   g0528(.dina(new_new_n1102__), .dinb(new_new_n2205__), .dout(new_new_n1489__));
  or1   g0529(.dina(new_new_n1130__), .dinb(new_new_n2209__), .dout(new_new_n1490__));
  and1  g0530(.dina(new_new_n1490__), .dinb(new_new_n1489__), .dout(new_new_n1491__));
  or1   g0531(.dina(new_new_n2216__), .dinb(new_new_n1026__), .dout(new_new_n1492__));
  and1  g0532(.dina(new_new_n1488__), .dinb(new_new_n1485__), .dout(new_new_n1493__));
  and1  g0533(.dina(new_new_n1493__), .dinb(new_new_n1491__), .dout(new_new_n1494__));
  and1  g0534(.dina(new_new_n1494__), .dinb(new_new_n1492__), .dout(new_new_n1495__));
  or1   g0535(.dina(new_new_n2179__), .dinb(new_new_n950__), .dout(new_new_n1496__));
  or1   g0536(.dina(new_new_n1300__), .dinb(new_new_n2186__), .dout(new_new_n1497__));
  and1  g0537(.dina(new_new_n1497__), .dinb(new_new_n1496__), .dout(new_new_n1498__));
  or1   g0538(.dina(new_new_n1198__), .dinb(new_new_n2193__), .dout(new_new_n1499__));
  or1   g0539(.dina(new_new_n1138__), .dinb(new_new_n2200__), .dout(new_new_n1500__));
  and1  g0540(.dina(new_new_n1500__), .dinb(new_new_n1499__), .dout(new_new_n1501__));
  or1   g0541(.dina(new_new_n1110__), .dinb(new_new_n2204__), .dout(new_new_n1502__));
  or1   g0542(.dina(new_new_n1132__), .dinb(new_new_n2209__), .dout(new_new_n1503__));
  and1  g0543(.dina(new_new_n1503__), .dinb(new_new_n1502__), .dout(new_new_n1504__));
  or1   g0544(.dina(new_new_n2216__), .dinb(new_new_n1032__), .dout(new_new_n1505__));
  and1  g0545(.dina(new_new_n1501__), .dinb(new_new_n1498__), .dout(new_new_n1506__));
  and1  g0546(.dina(new_new_n1506__), .dinb(new_new_n1504__), .dout(new_new_n1507__));
  and1  g0547(.dina(new_new_n1507__), .dinb(new_new_n1505__), .dout(new_new_n1508__));
  or1   g0548(.dina(new_new_n1212__), .dinb(new_new_n1190__), .dout(new_new_n1509__));
  and1  g0549(.dina(new_new_n1509__), .dinb(new_new_n2220__), .dout(new_new_n1510__));
  or1   g0550(.dina(new_new_n2181__), .dinb(new_new_n936__), .dout(new_new_n1511__));
  or1   g0551(.dina(new_new_n1286__), .dinb(new_new_n2188__), .dout(new_new_n1512__));
  and1  g0552(.dina(new_new_n1512__), .dinb(new_new_n1511__), .dout(new_new_n1513__));
  or1   g0553(.dina(new_new_n1208__), .dinb(new_new_n2195__), .dout(new_new_n1514__));
  or1   g0554(.dina(new_new_n1174__), .dinb(new_new_n2202__), .dout(new_new_n1515__));
  and1  g0555(.dina(new_new_n1515__), .dinb(new_new_n1514__), .dout(new_new_n1516__));
  or1   g0556(.dina(new_new_n1150__), .dinb(new_new_n2211__), .dout(new_new_n1517__));
  or1   g0557(.dina(new_new_n2218__), .dinb(new_new_n1014__), .dout(new_new_n1518__));
  and1  g0558(.dina(new_new_n1518__), .dinb(new_new_n1517__), .dout(new_new_n1519__));
  and1  g0559(.dina(new_new_n1516__), .dinb(new_new_n1513__), .dout(new_new_n1520__));
  and1  g0560(.dina(new_new_n1520__), .dinb(new_new_n1519__), .dout(new_new_n1521__));
  or1   g0561(.dina(new_new_n1128__), .dinb(new_new_n2181__), .dout(new_new_n1522__));
  or1   g0562(.dina(new_new_n1306__), .dinb(new_new_n2188__), .dout(new_new_n1523__));
  and1  g0563(.dina(new_new_n1523__), .dinb(new_new_n1522__), .dout(new_new_n1524__));
  or1   g0564(.dina(new_new_n1210__), .dinb(new_new_n2195__), .dout(new_new_n1525__));
  or1   g0565(.dina(new_new_n2220__), .dinb(new_new_n2202__), .dout(new_new_n1526__));
  and1  g0566(.dina(new_new_n1526__), .dinb(new_new_n1525__), .dout(new_new_n1527__));
  or1   g0567(.dina(new_new_n1176__), .dinb(new_new_n2211__), .dout(new_new_n1528__));
  or1   g0568(.dina(new_new_n2218__), .dinb(new_new_n996__), .dout(new_new_n1529__));
  and1  g0569(.dina(new_new_n1529__), .dinb(new_new_n1528__), .dout(new_new_n1530__));
  and1  g0570(.dina(new_new_n1527__), .dinb(new_new_n1524__), .dout(new_new_n1531__));
  and1  g0571(.dina(new_new_n1531__), .dinb(new_new_n1530__), .dout(new_new_n1532__));
  or1   g0572(.dina(new_new_n2182__), .dinb(new_new_n924__), .dout(new_new_n1533__));
  or1   g0573(.dina(new_new_n1302__), .dinb(new_new_n2189__), .dout(new_new_n1534__));
  and1  g0574(.dina(new_new_n1534__), .dinb(new_new_n1533__), .dout(new_new_n1535__));
  or1   g0575(.dina(new_new_n1204__), .dinb(new_new_n2196__), .dout(new_new_n1536__));
  or1   g0576(.dina(new_new_n1170__), .dinb(new_new_n2203__), .dout(new_new_n1537__));
  and1  g0577(.dina(new_new_n1537__), .dinb(new_new_n1536__), .dout(new_new_n1538__));
  or1   g0578(.dina(new_new_n1148__), .dinb(new_new_n2212__), .dout(new_new_n1539__));
  or1   g0579(.dina(new_new_n2219__), .dinb(new_new_n1002__), .dout(new_new_n1540__));
  and1  g0580(.dina(new_new_n1540__), .dinb(new_new_n1539__), .dout(new_new_n1541__));
  and1  g0581(.dina(new_new_n1538__), .dinb(new_new_n1535__), .dout(new_new_n1542__));
  and1  g0582(.dina(new_new_n1542__), .dinb(new_new_n1541__), .dout(new_new_n1543__));
  or1   g0583(.dina(new_new_n2182__), .dinb(new_new_n930__), .dout(new_new_n1544__));
  or1   g0584(.dina(new_new_n1304__), .dinb(new_new_n2189__), .dout(new_new_n1545__));
  and1  g0585(.dina(new_new_n1545__), .dinb(new_new_n1544__), .dout(new_new_n1546__));
  or1   g0586(.dina(new_new_n1206__), .dinb(new_new_n2196__), .dout(new_new_n1547__));
  or1   g0587(.dina(new_new_n1172__), .dinb(new_new_n2203__), .dout(new_new_n1548__));
  and1  g0588(.dina(new_new_n1548__), .dinb(new_new_n1547__), .dout(new_new_n1549__));
  or1   g0589(.dina(new_new_n1146__), .dinb(new_new_n2212__), .dout(new_new_n1550__));
  or1   g0590(.dina(new_new_n2219__), .dinb(new_new_n1008__), .dout(new_new_n1551__));
  and1  g0591(.dina(new_new_n1551__), .dinb(new_new_n1550__), .dout(new_new_n1552__));
  and1  g0592(.dina(new_new_n1549__), .dinb(new_new_n1546__), .dout(new_new_n1553__));
  and1  g0593(.dina(new_new_n1553__), .dinb(new_new_n1552__), .dout(new_new_n1554__));
  or1   g0594(.dina(new_new_n1156__), .dinb(new_new_n1152__), .dout(new_new_n1555__));
  or1   g0595(.dina(new_new_n1555__), .dinb(new_new_n812__), .dout(new_new_n1556__));
  or1   g0596(.dina(new_new_n1556__), .dinb(new_new_n1182__), .dout(new_new_n1557__));
  and1  g0597(.dina(new_new_n2222__), .dinb(new_new_n2225__), .dout(new_new_n1558__));
  or1   g0598(.dina(new_new_n2227__), .dinb(new_new_n2229__), .dout(new_new_n1559__));
  and1  g0599(.dina(new_new_n2232__), .dinb(new_new_n2235__), .dout(new_new_n1560__));
  or1   g0600(.dina(new_new_n2237__), .dinb(new_new_n2239__), .dout(new_new_n1561__));
  and1  g0601(.dina(new_new_n2242__), .dinb(new_new_n2245__), .dout(new_new_n1562__));
  or1   g0602(.dina(new_new_n2247__), .dinb(new_new_n2249__), .dout(new_new_n1563__));
  and1  g0603(.dina(new_new_n1324__), .dinb(new_new_n1320__), .dout(new_new_n1564__));
  or1   g0604(.dina(new_new_n1323__), .dinb(new_new_n1319__), .dout(new_new_n1565__));
  and1  g0605(.dina(new_new_n1326__), .dinb(new_new_n1322__), .dout(new_new_n1566__));
  or1   g0606(.dina(new_new_n1325__), .dinb(new_new_n1321__), .dout(new_new_n1567__));
  and1  g0607(.dina(new_new_n1566__), .dinb(new_new_n1564__), .dout(new_new_n1568__));
  or1   g0608(.dina(new_new_n1567__), .dinb(new_new_n1565__), .dout(new_new_n1569__));
  and1  g0609(.dina(new_new_n2251__), .dinb(new_new_n2253__), .dout(new_new_n1570__));
  or1   g0610(.dina(new_new_n2256__), .dinb(new_new_n2259__), .dout(new_new_n1571__));
  and1  g0611(.dina(new_new_n1259__), .dinb(new_new_n1238__), .dout(new_new_n1572__));
  or1   g0612(.dina(new_new_n1260__), .dinb(new_new_n1237__), .dout(new_new_n1573__));
  and1  g0613(.dina(new_new_n2262__), .dinb(new_new_n1240__), .dout(new_new_n1574__));
  or1   g0614(.dina(new_new_n2264__), .dinb(new_new_n1239__), .dout(new_new_n1575__));
  and1  g0615(.dina(new_new_n2266__), .dinb(new_new_n1242__), .dout(new_new_n1576__));
  or1   g0616(.dina(new_new_n2268__), .dinb(new_new_n1241__), .dout(new_new_n1577__));
  and1  g0617(.dina(new_new_n2269__), .dinb(new_new_n1308__), .dout(new_new_n1578__));
  or1   g0618(.dina(new_new_n2270__), .dinb(new_new_n1307__), .dout(new_new_n1579__));
  and1  g0619(.dina(new_new_n2227__), .dinb(new_new_n2229__), .dout(new_new_n1580__));
  or1   g0620(.dina(new_new_n2222__), .dinb(new_new_n2225__), .dout(new_new_n1581__));
  and1  g0621(.dina(new_new_n2272__), .dinb(new_new_n2273__), .dout(new_new_n1582__));
  or1   g0622(.dina(new_new_n2275__), .dinb(new_new_n2277__), .dout(new_new_n1583__));
  and1  g0623(.dina(new_new_n2237__), .dinb(new_new_n2239__), .dout(new_new_n1584__));
  or1   g0624(.dina(new_new_n2232__), .dinb(new_new_n2235__), .dout(new_new_n1585__));
  and1  g0625(.dina(new_new_n2279__), .dinb(new_new_n2282__), .dout(new_new_n1586__));
  or1   g0626(.dina(new_new_n2284__), .dinb(new_new_n2287__), .dout(new_new_n1587__));
  and1  g0627(.dina(new_new_n2247__), .dinb(new_new_n2249__), .dout(new_new_n1588__));
  or1   g0628(.dina(new_new_n2242__), .dinb(new_new_n2245__), .dout(new_new_n1589__));
  and1  g0629(.dina(new_new_n2290__), .dinb(new_new_n2293__), .dout(new_new_n1590__));
  or1   g0630(.dina(new_new_n2296__), .dinb(new_new_n2300__), .dout(new_new_n1591__));
  and1  g0631(.dina(new_new_n2256__), .dinb(new_new_n2259__), .dout(new_new_n1592__));
  or1   g0632(.dina(new_new_n2251__), .dinb(new_new_n2253__), .dout(new_new_n1593__));
  and1  g0633(.dina(new_new_n1593__), .dinb(new_new_n2302__), .dout(new_new_n1594__));
  or1   g0634(.dina(new_new_n2303__), .dinb(new_new_n1570__), .dout(new_new_n1595__));
  and1  g0635(.dina(new_new_n2272__), .dinb(new_new_n2287__), .dout(new_new_n1596__));
  or1   g0636(.dina(new_new_n2275__), .dinb(new_new_n2282__), .dout(new_new_n1597__));
  and1  g0637(.dina(new_new_n2279__), .dinb(new_new_n2271__), .dout(new_new_n1598__));
  or1   g0638(.dina(new_new_n2284__), .dinb(new_new_n2274__), .dout(new_new_n1599__));
  and1  g0639(.dina(new_new_n2304__), .dinb(new_new_n2300__), .dout(new_new_n1600__));
  or1   g0640(.dina(new_new_n2305__), .dinb(new_new_n2293__), .dout(new_new_n1601__));
  and1  g0641(.dina(new_new_n2306__), .dinb(new_new_n2269__), .dout(new_new_n1602__));
  or1   g0642(.dina(new_new_n2307__), .dinb(new_new_n2270__), .dout(new_new_n1603__));
  and1  g0643(.dina(new_new_n1603__), .dinb(new_new_n1350__), .dout(new_new_n1604__));
  or1   g0644(.dina(new_new_n1602__), .dinb(new_new_n2308__), .dout(new_new_n1605__));
  and1  g0645(.dina(new_new_n2304__), .dinb(new_new_n2290__), .dout(new_new_n1606__));
  or1   g0646(.dina(new_new_n2305__), .dinb(new_new_n2296__), .dout(new_new_n1607__));
  and1  g0647(.dina(new_new_n1606__), .dinb(new_new_n2310__), .dout(new_new_n1608__));
  or1   g0648(.dina(new_new_n1607__), .dinb(new_new_n2313__), .dout(new_new_n1609__));
  and1  g0649(.dina(new_new_n1597__), .dinb(new_new_n2273__), .dout(new_new_n1610__));
  or1   g0650(.dina(new_new_n1596__), .dinb(new_new_n2277__), .dout(new_new_n1611__));
  and1  g0651(.dina(new_new_n1610__), .dinb(new_new_n1601__), .dout(new_new_n1612__));
  or1   g0652(.dina(new_new_n1611__), .dinb(new_new_n1600__), .dout(new_new_n1613__));
  and1  g0653(.dina(new_new_n1612__), .dinb(new_new_n1609__), .dout(new_new_n1614__));
  or1   g0654(.dina(new_new_n1613__), .dinb(new_new_n1608__), .dout(new_new_n1615__));
  or1   g0655(.dina(new_new_n2315__), .dinb(new_new_n1366__), .dout(new_new_n1616__));
  and1  g0656(.dina(new_new_n1374__), .dinb(new_new_n1368__), .dout(new_new_n1617__));
  and1  g0657(.dina(new_new_n1617__), .dinb(new_new_n2317__), .dout(new_new_n1618__));
  and1  g0658(.dina(new_new_n1376__), .dinb(new_new_n1370__), .dout(new_new_n1619__));
  and1  g0659(.dina(new_new_n1619__), .dinb(new_new_n2317__), .dout(new_new_n1620__));
  and1  g0660(.dina(new_new_n1378__), .dinb(new_new_n1372__), .dout(new_new_n1621__));
  and1  g0661(.dina(new_new_n1621__), .dinb(new_new_n2318__), .dout(new_new_n1622__));
  or1   g0662(.dina(new_new_n2320__), .dinb(new_new_n2321__), .dout(new_new_n1623__));
  or1   g0663(.dina(new_new_n2323__), .dinb(new_new_n2324__), .dout(new_new_n1624__));
  or1   g0664(.dina(new_new_n2326__), .dinb(new_new_n2327__), .dout(new_new_n1625__));
  and1  g0665(.dina(new_new_n2328__), .dinb(new_new_n2330__), .dout(new_new_n1626__));
  or1   g0666(.dina(new_new_n1396__), .dinb(new_new_n2331__), .dout(new_new_n1627__));
  and1  g0667(.dina(new_new_n1626__), .dinb(new_new_n2333__), .dout(new_new_n1628__));
  or1   g0668(.dina(new_new_n1627__), .dinb(new_new_n1398__), .dout(new_new_n1629__));
  and1  g0669(.dina(new_new_n2320__), .dinb(new_new_n2321__), .dout(new_new_n1630__));
  and1  g0670(.dina(new_new_n2323__), .dinb(new_new_n2324__), .dout(new_new_n1631__));
  and1  g0671(.dina(new_new_n2326__), .dinb(new_new_n2327__), .dout(new_new_n1632__));
  or1   g0672(.dina(new_new_n2334__), .dinb(new_new_n1327__), .dout(new_new_n1633__));
  or1   g0673(.dina(new_new_n1362__), .dinb(new_new_n2336__), .dout(new_new_n1634__));
  and1  g0674(.dina(new_new_n1634__), .dinb(new_new_n1633__), .dout(new_new_n1635__));
  and1  g0675(.dina(new_new_n1635__), .dinb(new_new_n2318__), .dout(new_new_n1636__));
  or1   g0676(.dina(new_new_n2338__), .dinb(new_new_n1382__), .dout(new_new_n1637__));
  or1   g0677(.dina(new_new_n2339__), .dinb(new_new_n2341__), .dout(new_new_n1638__));
  or1   g0678(.dina(new_new_n1577__), .dinb(new_new_n2343__), .dout(new_new_n1639__));
  and1  g0679(.dina(new_new_n1639__), .dinb(new_new_n1638__), .dout(new_new_n1640__));
  or1   g0680(.dina(new_new_n2344__), .dinb(new_new_n2306__), .dout(new_new_n1641__));
  or1   g0681(.dina(new_new_n1579__), .dinb(new_new_n2307__), .dout(new_new_n1642__));
  and1  g0682(.dina(new_new_n1642__), .dinb(new_new_n1641__), .dout(new_new_n1643__));
  or1   g0683(.dina(new_new_n2310__), .dinb(new_new_n2345__), .dout(new_new_n1644__));
  or1   g0684(.dina(new_new_n2313__), .dinb(new_new_n1591__), .dout(new_new_n1645__));
  and1  g0685(.dina(new_new_n1645__), .dinb(new_new_n1644__), .dout(new_new_n1646__));
  and1  g0686(.dina(new_new_n2347__), .dinb(new_new_n2349__), .dout(new_new_n1647__));
  or1   g0687(.dina(new_new_n2350__), .dinb(new_new_n2351__), .dout(new_new_n1648__));
  and1  g0688(.dina(new_new_n2350__), .dinb(new_new_n2351__), .dout(new_new_n1649__));
  or1   g0689(.dina(new_new_n2347__), .dinb(new_new_n2349__), .dout(new_new_n1650__));
  and1  g0690(.dina(new_new_n1650__), .dinb(new_new_n1648__), .dout(new_new_n1651__));
  or1   g0691(.dina(new_new_n1649__), .dinb(new_new_n1647__), .dout(new_new_n1652__));
  and1  g0692(.dina(new_new_n2353__), .dinb(new_new_n2355__), .dout(new_new_n1653__));
  or1   g0693(.dina(new_new_n2356__), .dinb(new_new_n2357__), .dout(new_new_n1654__));
  and1  g0694(.dina(new_new_n2356__), .dinb(new_new_n2357__), .dout(new_new_n1655__));
  or1   g0695(.dina(new_new_n2353__), .dinb(new_new_n2355__), .dout(new_new_n1656__));
  and1  g0696(.dina(new_new_n1656__), .dinb(new_new_n1654__), .dout(new_new_n1657__));
  or1   g0697(.dina(new_new_n1655__), .dinb(new_new_n1653__), .dout(new_new_n1658__));
  or1   g0698(.dina(new_new_n1657__), .dinb(new_new_n1651__), .dout(new_new_n1659__));
  or1   g0699(.dina(new_new_n1658__), .dinb(new_new_n1652__), .dout(new_new_n1660__));
  and1  g0700(.dina(new_new_n1660__), .dinb(new_new_n1659__), .dout(new_new_n1661__));
  and1  g0701(.dina(new_new_n2359__), .dinb(new_new_n2361__), .dout(new_new_n1662__));
  or1   g0702(.dina(new_new_n2362__), .dinb(new_new_n2363__), .dout(new_new_n1663__));
  and1  g0703(.dina(new_new_n2362__), .dinb(new_new_n2363__), .dout(new_new_n1664__));
  or1   g0704(.dina(new_new_n2359__), .dinb(new_new_n2361__), .dout(new_new_n1665__));
  and1  g0705(.dina(new_new_n1665__), .dinb(new_new_n1663__), .dout(new_new_n1666__));
  or1   g0706(.dina(new_new_n1664__), .dinb(new_new_n1662__), .dout(new_new_n1667__));
  and1  g0707(.dina(new_new_n2364__), .dinb(new_new_n2366__), .dout(new_new_n1668__));
  or1   g0708(.dina(new_new_n2367__), .dinb(new_new_n2368__), .dout(new_new_n1669__));
  and1  g0709(.dina(new_new_n2367__), .dinb(new_new_n2368__), .dout(new_new_n1670__));
  or1   g0710(.dina(new_new_n2364__), .dinb(new_new_n2366__), .dout(new_new_n1671__));
  and1  g0711(.dina(new_new_n1671__), .dinb(new_new_n1669__), .dout(new_new_n1672__));
  or1   g0712(.dina(new_new_n1670__), .dinb(new_new_n1668__), .dout(new_new_n1673__));
  or1   g0713(.dina(new_new_n1672__), .dinb(new_new_n1666__), .dout(new_new_n1674__));
  or1   g0714(.dina(new_new_n1673__), .dinb(new_new_n1667__), .dout(new_new_n1675__));
  and1  g0715(.dina(new_new_n1675__), .dinb(new_new_n1674__), .dout(new_new_n1676__));
  and1  g0716(.dina(new_new_n2224__), .dinb(new_new_n2258__), .dout(new_new_n1677__));
  or1   g0717(.dina(new_new_n2230__), .dinb(new_new_n2254__), .dout(new_new_n1678__));
  and1  g0718(.dina(new_new_n2230__), .dinb(new_new_n2254__), .dout(new_new_n1679__));
  or1   g0719(.dina(new_new_n2226__), .dinb(new_new_n2260__), .dout(new_new_n1680__));
  and1  g0720(.dina(new_new_n1680__), .dinb(new_new_n1678__), .dout(new_new_n1681__));
  or1   g0721(.dina(new_new_n1679__), .dinb(new_new_n1677__), .dout(new_new_n1682__));
  and1  g0722(.dina(new_new_n2244__), .dinb(new_new_n2234__), .dout(new_new_n1683__));
  or1   g0723(.dina(new_new_n2250__), .dinb(new_new_n2240__), .dout(new_new_n1684__));
  and1  g0724(.dina(new_new_n2250__), .dinb(new_new_n2240__), .dout(new_new_n1685__));
  or1   g0725(.dina(new_new_n2246__), .dinb(new_new_n2236__), .dout(new_new_n1686__));
  and1  g0726(.dina(new_new_n1686__), .dinb(new_new_n1684__), .dout(new_new_n1687__));
  or1   g0727(.dina(new_new_n1685__), .dinb(new_new_n1683__), .dout(new_new_n1688__));
  or1   g0728(.dina(new_new_n1687__), .dinb(new_new_n1681__), .dout(new_new_n1689__));
  or1   g0729(.dina(new_new_n1688__), .dinb(new_new_n1682__), .dout(new_new_n1690__));
  and1  g0730(.dina(new_new_n1690__), .dinb(new_new_n1689__), .dout(new_new_n1691__));
  and1  g0731(.dina(new_new_n2370__), .dinb(new_new_n2372__), .dout(new_new_n1692__));
  or1   g0732(.dina(new_new_n2373__), .dinb(new_new_n2374__), .dout(new_new_n1693__));
  and1  g0733(.dina(new_new_n2373__), .dinb(new_new_n2374__), .dout(new_new_n1694__));
  or1   g0734(.dina(new_new_n2370__), .dinb(new_new_n2372__), .dout(new_new_n1695__));
  and1  g0735(.dina(new_new_n1695__), .dinb(new_new_n1693__), .dout(new_new_n1696__));
  or1   g0736(.dina(new_new_n1694__), .dinb(new_new_n1692__), .dout(new_new_n1697__));
  and1  g0737(.dina(new_new_n2376__), .dinb(new_new_n2378__), .dout(new_new_n1698__));
  or1   g0738(.dina(new_new_n2379__), .dinb(new_new_n2380__), .dout(new_new_n1699__));
  and1  g0739(.dina(new_new_n2379__), .dinb(new_new_n2380__), .dout(new_new_n1700__));
  or1   g0740(.dina(new_new_n2376__), .dinb(new_new_n2378__), .dout(new_new_n1701__));
  and1  g0741(.dina(new_new_n1701__), .dinb(new_new_n1699__), .dout(new_new_n1702__));
  or1   g0742(.dina(new_new_n1700__), .dinb(new_new_n1698__), .dout(new_new_n1703__));
  or1   g0743(.dina(new_new_n1702__), .dinb(new_new_n1696__), .dout(new_new_n1704__));
  or1   g0744(.dina(new_new_n1703__), .dinb(new_new_n1697__), .dout(new_new_n1705__));
  and1  g0745(.dina(new_new_n1705__), .dinb(new_new_n1704__), .dout(new_new_n1706__));
  or1   g0746(.dina(new_new_n1162__), .dinb(new_new_n1160__), .dout(new_new_n1707__));
  or1   g0747(.dina(new_new_n1707__), .dinb(new_new_n842__), .dout(new_new_n1708__));
  or1   g0748(.dina(new_new_n1708__), .dinb(new_new_n850__), .dout(new_new_n1709__));
  or1   g0749(.dina(new_new_n1709__), .dinb(new_new_n2381__), .dout(new_new_n1710__));
  or1   g0750(.dina(new_new_n1710__), .dinb(new_new_n856__), .dout(new_new_n1711__));
  and1  g0751(.dina(new_new_n2383__), .dinb(new_new_n2262__), .dout(new_new_n1712__));
  or1   g0752(.dina(new_new_n2384__), .dinb(new_new_n2264__), .dout(new_new_n1713__));
  and1  g0753(.dina(new_new_n2266__), .dinb(new_new_n2261__), .dout(new_new_n1714__));
  or1   g0754(.dina(new_new_n2268__), .dinb(new_new_n2263__), .dout(new_new_n1715__));
  and1  g0755(.dina(new_new_n1714__), .dinb(new_new_n2341__), .dout(new_new_n1716__));
  or1   g0756(.dina(new_new_n1715__), .dinb(new_new_n2343__), .dout(new_new_n1717__));
  and1  g0757(.dina(new_new_n1713__), .dinb(new_new_n1270__), .dout(new_new_n1718__));
  or1   g0758(.dina(new_new_n1712__), .dinb(new_new_n2385__), .dout(new_new_n1719__));
  and1  g0759(.dina(new_new_n1718__), .dinb(new_new_n1717__), .dout(new_new_n1720__));
  or1   g0760(.dina(new_new_n1719__), .dinb(new_new_n1716__), .dout(new_new_n1721__));
  or1   g0761(.dina(new_new_n1721__), .dinb(new_new_n2386__), .dout(new_new_n1722__));
  or1   g0762(.dina(new_new_n1720__), .dinb(new_new_n1573__), .dout(new_new_n1723__));
  and1  g0763(.dina(new_new_n1723__), .dinb(new_new_n1722__), .dout(new_new_n1724__));
  and1  g0764(.dina(new_new_n2265__), .dinb(new_new_n2340__), .dout(new_new_n1725__));
  or1   g0765(.dina(new_new_n2267__), .dinb(new_new_n2342__), .dout(new_new_n1726__));
  and1  g0766(.dina(new_new_n1726__), .dinb(new_new_n2384__), .dout(new_new_n1727__));
  or1   g0767(.dina(new_new_n1725__), .dinb(new_new_n2383__), .dout(new_new_n1728__));
  or1   g0768(.dina(new_new_n1728__), .dinb(new_new_n2387__), .dout(new_new_n1729__));
  or1   g0769(.dina(new_new_n1727__), .dinb(new_new_n1575__), .dout(new_new_n1730__));
  and1  g0770(.dina(new_new_n1730__), .dinb(new_new_n1729__), .dout(new_new_n1731__));
  and1  g0771(.dina(new_new_n2280__), .dinb(new_new_n2299__), .dout(new_new_n1732__));
  or1   g0772(.dina(new_new_n2285__), .dinb(new_new_n2294__), .dout(new_new_n1733__));
  and1  g0773(.dina(new_new_n2291__), .dinb(new_new_n2280__), .dout(new_new_n1734__));
  or1   g0774(.dina(new_new_n2297__), .dinb(new_new_n2285__), .dout(new_new_n1735__));
  and1  g0775(.dina(new_new_n1734__), .dinb(new_new_n2311__), .dout(new_new_n1736__));
  or1   g0776(.dina(new_new_n1735__), .dinb(new_new_n2314__), .dout(new_new_n1737__));
  and1  g0777(.dina(new_new_n1733__), .dinb(new_new_n2281__), .dout(new_new_n1738__));
  or1   g0778(.dina(new_new_n1732__), .dinb(new_new_n2288__), .dout(new_new_n1739__));
  and1  g0779(.dina(new_new_n1738__), .dinb(new_new_n1737__), .dout(new_new_n1740__));
  or1   g0780(.dina(new_new_n1739__), .dinb(new_new_n1736__), .dout(new_new_n1741__));
  or1   g0781(.dina(new_new_n1741__), .dinb(new_new_n2388__), .dout(new_new_n1742__));
  or1   g0782(.dina(new_new_n1740__), .dinb(new_new_n1583__), .dout(new_new_n1743__));
  and1  g0783(.dina(new_new_n1743__), .dinb(new_new_n1742__), .dout(new_new_n1744__));
  and1  g0784(.dina(new_new_n2311__), .dinb(new_new_n2291__), .dout(new_new_n1745__));
  or1   g0785(.dina(new_new_n2314__), .dinb(new_new_n2297__), .dout(new_new_n1746__));
  and1  g0786(.dina(new_new_n1746__), .dinb(new_new_n2294__), .dout(new_new_n1747__));
  or1   g0787(.dina(new_new_n1745__), .dinb(new_new_n2301__), .dout(new_new_n1748__));
  or1   g0788(.dina(new_new_n1748__), .dinb(new_new_n2389__), .dout(new_new_n1749__));
  or1   g0789(.dina(new_new_n1747__), .dinb(new_new_n1587__), .dout(new_new_n1750__));
  and1  g0790(.dina(new_new_n1750__), .dinb(new_new_n1749__), .dout(new_new_n1751__));
  or1   g0791(.dina(new_new_n2390__), .dinb(new_new_n2391__), .dout(new_new_n1752__));
  or1   g0792(.dina(new_new_n1614__), .dinb(new_new_n1595__), .dout(new_new_n1753__));
  and1  g0793(.dina(new_new_n1753__), .dinb(new_new_n1752__), .dout(new_new_n1754__));
  or1   g0794(.dina(new_new_n2393__), .dinb(new_new_n2394__), .dout(new_new_n1755__));
  and1  g0795(.dina(new_new_n2395__), .dinb(new_new_n975__), .dout(new_new_n1756__));
  or1   g0796(.dina(new_new_n2396__), .dinb(new_new_n2397__), .dout(new_new_n1757__));
  or1   g0797(.dina(new_new_n1757__), .dinb(new_new_n1330__), .dout(new_new_n1758__));
  or1   g0798(.dina(new_new_n1758__), .dinb(new_new_n1359__), .dout(new_new_n1759__));
  and1  g0799(.dina(new_new_n1347__), .dinb(new_new_n2398__), .dout(new_new_n1760__));
  or1   g0800(.dina(new_new_n2396__), .dinb(new_new_n1273__), .dout(new_new_n1761__));
  or1   g0801(.dina(new_new_n1761__), .dinb(new_new_n1334__), .dout(new_new_n1762__));
  or1   g0802(.dina(new_new_n2400__), .dinb(new_new_n2334__), .dout(new_new_n1763__));
  and1  g0803(.dina(new_new_n2402__), .dinb(new_new_n2404__), .dout(new_new_n1764__));
  and1  g0804(.dina(new_new_n1764__), .dinb(new_new_n2407__), .dout(new_new_n1765__));
  or1   g0805(.dina(new_new_n1765__), .dinb(new_new_n2331__), .dout(new_new_n1766__));
  or1   g0806(.dina(new_new_n2409__), .dinb(new_new_n820__), .dout(new_new_n1767__));
  or1   g0807(.dina(new_new_n1767__), .dinb(new_new_n868__), .dout(new_new_n1768__));
  and1  g0808(.dina(new_new_n2393__), .dinb(new_new_n2394__), .dout(new_new_n1769__));
  or1   g0809(.dina(new_new_n2410__), .dinb(new_new_n2407__), .dout(new_new_n1770__));
  or1   g0810(.dina(new_new_n2411__), .dinb(new_new_n1386__), .dout(new_new_n1771__));
  and1  g0811(.dina(new_new_n1771__), .dinb(new_new_n1770__), .dout(new_new_n1772__));
  and1  g0812(.dina(new_new_n1772__), .dinb(new_new_n2412__), .dout(new_new_n1773__));
  and1  g0813(.dina(new_new_n1773__), .dinb(new_new_n1381__), .dout(new_new_n1774__));
  and1  g0814(.dina(new_new_n1774__), .dinb(new_new_n2404__), .dout(new_new_n1775__));
  and1  g0815(.dina(new_new_n2330__), .dinb(new_new_n2413__), .dout(new_new_n1776__));
  and1  g0816(.dina(new_new_n1776__), .dinb(new_new_n2333__), .dout(new_new_n1777__));
  and1  g0817(.dina(new_new_n1777__), .dinb(new_new_n2408__), .dout(new_new_n1778__));
  or1   g0818(.dina(new_new_n2409__), .dinb(new_new_n2338__), .dout(new_new_n1779__));
  or1   g0819(.dina(new_new_n1779__), .dinb(new_new_n2411__), .dout(new_new_n1780__));
  and1  g0820(.dina(new_new_n1780__), .dinb(new_new_n1778__), .dout(new_new_n1781__));
  or1   g0821(.dina(new_new_n1781__), .dinb(new_new_n1775__), .dout(new_new_n1782__));
  or1   g0822(.dina(new_new_n2415__), .dinb(new_new_n2417__), .dout(new_new_n1783__));
  or1   g0823(.dina(new_new_n2418__), .dinb(new_new_n2415__), .dout(new_new_n1784__));
  or1   g0824(.dina(new_new_n2419__), .dinb(new_new_n2421__), .dout(new_new_n1785__));
  or1   g0825(.dina(new_new_n2419__), .dinb(new_new_n2422__), .dout(new_new_n1786__));
  or1   g0826(.dina(new_new_n1786__), .dinb(new_new_n1114__), .dout(new_new_n1787__));
  and1  g0827(.dina(new_new_n1783__), .dinb(new_new_n2424__), .dout(new_new_n1788__));
  and1  g0828(.dina(new_new_n1788__), .dinb(new_new_n1785__), .dout(new_new_n1789__));
  and1  g0829(.dina(new_new_n1789__), .dinb(new_new_n1787__), .dout(new_new_n1790__));
  or1   g0830(.dina(new_new_n1230__), .dinb(new_new_n2426__), .dout(new_new_n1791__));
  or1   g0831(.dina(new_new_n2336__), .dinb(new_new_n928__), .dout(new_new_n1792__));
  and1  g0832(.dina(new_new_n1792__), .dinb(new_new_n1791__), .dout(new_new_n1793__));
  or1   g0833(.dina(new_new_n2400__), .dinb(new_new_n1342__), .dout(new_new_n1794__));
  and1  g0834(.dina(new_new_n1794__), .dinb(new_new_n2428__), .dout(new_new_n1795__));
  and1  g0835(.dina(new_new_n1795__), .dinb(new_new_n1793__), .dout(new_new_n1796__));
  or1   g0836(.dina(new_new_n2397__), .dinb(new_new_n2426__), .dout(new_new_n1797__));
  or1   g0837(.dina(new_new_n2337__), .dinb(new_new_n934__), .dout(new_new_n1798__));
  and1  g0838(.dina(new_new_n1798__), .dinb(new_new_n1797__), .dout(new_new_n1799__));
  or1   g0839(.dina(new_new_n2401__), .dinb(new_new_n1344__), .dout(new_new_n1800__));
  and1  g0840(.dina(new_new_n1800__), .dinb(new_new_n2428__), .dout(new_new_n1801__));
  and1  g0841(.dina(new_new_n1801__), .dinb(new_new_n1799__), .dout(new_new_n1802__));
  or1   g0842(.dina(new_new_n986__), .dinb(new_new_n2425__), .dout(new_new_n1803__));
  or1   g0843(.dina(new_new_n2337__), .dinb(new_new_n940__), .dout(new_new_n1804__));
  and1  g0844(.dina(new_new_n1804__), .dinb(new_new_n1803__), .dout(new_new_n1805__));
  or1   g0845(.dina(new_new_n2401__), .dinb(new_new_n1346__), .dout(new_new_n1806__));
  and1  g0846(.dina(new_new_n1806__), .dinb(new_new_n2429__), .dout(new_new_n1807__));
  and1  g0847(.dina(new_new_n1807__), .dinb(new_new_n1805__), .dout(new_new_n1808__));
  or1   g0848(.dina(new_new_n2430__), .dinb(new_new_n1629__), .dout(new_new_n1809__));
  or1   g0849(.dina(new_new_n1809__), .dinb(new_new_n834__), .dout(new_new_n1810__));
  and1  g0850(.dina(new_new_n2432__), .dinb(new_new_n2434__), .dout(new_new_n1811__));
  and1  g0851(.dina(new_new_n2432__), .dinb(new_new_n2435__), .dout(new_new_n1812__));
  and1  g0852(.dina(new_new_n2433__), .dinb(new_new_n2436__), .dout(new_new_n1813__));
  and1  g0853(.dina(new_new_n2438__), .dinb(new_new_n2440__), .dout(new_new_n1814__));
  and1  g0854(.dina(new_new_n2438__), .dinb(new_new_n2441__), .dout(new_new_n1815__));
  and1  g0855(.dina(new_new_n2439__), .dinb(new_new_n2442__), .dout(new_new_n1816__));
  buf1  g0856(.din(new_new_n1400__), .dout(G855));
  buf1  g0857(.din(new_new_n1402__), .dout(G856));
  buf1  g0858(.din(new_new_n2151__), .dout(G857));
  buf1  g0859(.din(new_new_n1404__), .dout(G858));
  buf1  g0860(.din(new_new_n1407__), .dout(G859));
  buf1  g0861(.din(new_new_n1414__), .dout(G860));
  buf1  g0862(.din(new_new_n1416__), .dout(G861));
  not1  g0863(.din(new_new_n1418__), .dout(G862));
  not1  g0864(.din(new_new_n1419__), .dout(G863));
  not1  g0865(.din(new_new_n1421__), .dout(G864));
  not1  g0866(.din(new_new_n1422__), .dout(G865));
  buf1  g0867(.din(new_new_n1126__), .dout(G866));
  buf1  g0868(.din(new_new_n1424__), .dout(G867));
  buf1  g0869(.din(new_new_n1427__), .dout(G868));
  not1  g0870(.din(new_new_n1428__), .dout(G869));
  buf1  g0871(.din(new_new_n1443__), .dout(G870));
  buf1  g0872(.din(new_new_n1458__), .dout(G871));
  buf1  g0873(.din(new_new_n1471__), .dout(G872));
  buf1  g0874(.din(new_new_n1482__), .dout(G873));
  buf1  g0875(.din(new_new_n1495__), .dout(G874));
  buf1  g0876(.din(new_new_n1508__), .dout(G875));
  buf1  g0877(.din(new_new_n1510__), .dout(G876));
  buf1  g0878(.din(new_new_n1521__), .dout(G877));
  buf1  g0879(.din(new_new_n1532__), .dout(G878));
  buf1  g0880(.din(new_new_n1543__), .dout(G879));
  buf1  g0881(.din(new_new_n1554__), .dout(G880));
  buf1  g0882(.din(new_new_n1151__), .dout(n3413));
  buf1  g0883(.din(new_new_n1155__), .dout(n3416));
  buf1  g0884(.din(new_new_n687__), .dout(n3419));
  buf1  g0885(.din(new_new_n807__), .dout(n3422));
  buf1  g0886(.din(new_new_n809__), .dout(n3425));
  buf1  g0887(.din(new_new_n811__), .dout(n3428));
  buf1  g0888(.din(new_new_n1157__), .dout(n3431));
  buf1  g0889(.din(new_new_n1153__), .dout(n3434));
  buf1  g0890(.din(new_new_n693__), .dout(n3437));
  buf1  g0891(.din(new_new_n1177__), .dout(n3440));
  buf1  g0892(.din(new_new_n695__), .dout(n3443));
  buf1  g0893(.din(new_new_n823__), .dout(n3446));
  buf1  g0894(.din(new_new_n825__), .dout(n3449));
  buf1  g0895(.din(new_new_n827__), .dout(n3452));
  buf1  g0896(.din(new_new_n1159__), .dout(n3455));
  buf1  g0897(.din(new_new_n701__), .dout(n3458));
  buf1  g0898(.din(new_new_n1161__), .dout(n3461));
  buf1  g0899(.din(new_new_n705__), .dout(n3464));
  buf1  g0900(.din(new_new_n837__), .dout(n3467));
  buf1  g0901(.din(new_new_n839__), .dout(n3470));
  buf1  g0902(.din(new_new_n841__), .dout(n3473));
  buf1  g0903(.din(new_new_n707__), .dout(n3476));
  buf1  g0904(.din(new_new_n845__), .dout(n3479));
  buf1  g0905(.din(new_new_n847__), .dout(n3482));
  buf1  g0906(.din(new_new_n709__), .dout(n3485));
  buf1  g0907(.din(new_new_n851__), .dout(n3488));
  buf1  g0908(.din(new_new_n853__), .dout(n3491));
  buf1  g0909(.din(new_new_n711__), .dout(n3494));
  buf1  g0910(.din(new_new_n857__), .dout(n3497));
  buf1  g0911(.din(new_new_n859__), .dout(n3500));
  buf1  g0912(.din(new_new_n861__), .dout(n3503));
  buf1  g0913(.din(new_new_n1163__), .dout(n3506));
  buf1  g0914(.din(new_new_n715__), .dout(n3509));
  buf1  g0915(.din(new_new_n1179__), .dout(n3512));
  buf1  g0916(.din(new_new_n717__), .dout(n3515));
  buf1  g0917(.din(new_new_n871__), .dout(n3518));
  buf1  g0918(.din(new_new_n873__), .dout(n3521));
  buf1  g0919(.din(new_new_n875__), .dout(n3524));
  buf1  g0920(.din(new_new_n719__), .dout(n3527));
  buf1  g0921(.din(new_new_n879__), .dout(n3530));
  buf1  g0922(.din(new_new_n881__), .dout(n3533));
  buf1  g0923(.din(new_new_n883__), .dout(n3536));
  buf1  g0924(.din(new_new_n721__), .dout(n3539));
  buf1  g0925(.din(new_new_n887__), .dout(n3542));
  buf1  g0926(.din(new_new_n889__), .dout(n3545));
  buf1  g0927(.din(new_new_n891__), .dout(n3548));
  buf1  g0928(.din(new_new_n723__), .dout(n3551));
  buf1  g0929(.din(new_new_n895__), .dout(n3554));
  buf1  g0930(.din(new_new_n897__), .dout(n3557));
  buf1  g0931(.din(new_new_n899__), .dout(n3560));
  buf1  g0932(.din(new_new_n725__), .dout(n3563));
  buf1  g0933(.din(new_new_n903__), .dout(n3566));
  buf1  g0934(.din(new_new_n905__), .dout(n3569));
  buf1  g0935(.din(new_new_n907__), .dout(n3572));
  buf1  g0936(.din(new_new_n727__), .dout(n3575));
  buf1  g0937(.din(new_new_n911__), .dout(n3578));
  buf1  g0938(.din(new_new_n913__), .dout(n3581));
  buf1  g0939(.din(new_new_n915__), .dout(n3584));
  buf1  g0940(.din(new_new_n729__), .dout(n3587));
  buf1  g0941(.din(new_new_n919__), .dout(n3590));
  buf1  g0942(.din(new_new_n2346__), .dout(n3593));
  buf1  g0943(.din(new_new_n731__), .dout(n3596));
  buf1  g0944(.din(new_new_n925__), .dout(n3599));
  buf1  g0945(.din(new_new_n2348__), .dout(n3602));
  buf1  g0946(.din(new_new_n733__), .dout(n3605));
  buf1  g0947(.din(new_new_n931__), .dout(n3608));
  buf1  g0948(.din(new_new_n2354__), .dout(n3611));
  buf1  g0949(.din(new_new_n735__), .dout(n3614));
  buf1  g0950(.din(new_new_n937__), .dout(n3617));
  buf1  g0951(.din(new_new_n2352__), .dout(n3620));
  buf1  g0952(.din(new_new_n737__), .dout(n3623));
  buf1  g0953(.din(new_new_n2358__), .dout(n3626));
  buf1  g0954(.din(new_new_n739__), .dout(n3629));
  buf1  g0955(.din(new_new_n2360__), .dout(n3632));
  buf1  g0956(.din(new_new_n741__), .dout(n3635));
  buf1  g0957(.din(new_new_n2365__), .dout(n3638));
  buf1  g0958(.din(new_new_n743__), .dout(n3641));
  buf1  g0959(.din(new_new_n745__), .dout(n3644));
  buf1  g0960(.din(new_new_n957__), .dout(n3647));
  buf1  g0961(.din(new_new_n959__), .dout(n3650));
  buf1  g0962(.din(new_new_n961__), .dout(n3653));
  buf1  g0963(.din(new_new_n747__), .dout(n3656));
  buf1  g0964(.din(new_new_n965__), .dout(n3659));
  buf1  g0965(.din(new_new_n967__), .dout(n3662));
  buf1  g0966(.din(new_new_n969__), .dout(n3665));
  buf1  g0967(.din(new_new_n749__), .dout(n3668));
  buf1  g0968(.din(new_new_n973__), .dout(n3671));
  buf1  g0969(.din(new_new_n751__), .dout(n3674));
  buf1  g0970(.din(new_new_n753__), .dout(n3677));
  buf1  g0971(.din(new_new_n755__), .dout(n3680));
  buf1  g0972(.din(new_new_n757__), .dout(n3683));
  buf1  g0973(.din(new_new_n983__), .dout(n3686));
  buf1  g0974(.din(new_new_n759__), .dout(n3689));
  buf1  g0975(.din(new_new_n763__), .dout(n3692));
  buf1  g0976(.din(new_new_n989__), .dout(n3695));
  buf1  g0977(.din(new_new_n991__), .dout(n3698));
  buf1  g0978(.din(new_new_n2260__), .dout(n3701));
  buf1  g0979(.din(new_new_n765__), .dout(n3704));
  buf1  g0980(.din(new_new_n997__), .dout(n3707));
  buf1  g0981(.din(new_new_n2226__), .dout(n3710));
  buf1  g0982(.din(new_new_n767__), .dout(n3713));
  buf1  g0983(.din(new_new_n1003__), .dout(n3716));
  buf1  g0984(.din(new_new_n2236__), .dout(n3719));
  buf1  g0985(.din(new_new_n769__), .dout(n3722));
  buf1  g0986(.din(new_new_n1009__), .dout(n3725));
  buf1  g0987(.din(new_new_n2246__), .dout(n3728));
  buf1  g0988(.din(new_new_n771__), .dout(n3731));
  buf1  g0989(.din(new_new_n1015__), .dout(n3734));
  buf1  g0990(.din(new_new_n2369__), .dout(n3737));
  buf1  g0991(.din(new_new_n773__), .dout(n3740));
  buf1  g0992(.din(new_new_n1021__), .dout(n3743));
  buf1  g0993(.din(new_new_n2371__), .dout(n3746));
  buf1  g0994(.din(new_new_n775__), .dout(n3749));
  buf1  g0995(.din(new_new_n1027__), .dout(n3752));
  buf1  g0996(.din(new_new_n2377__), .dout(n3755));
  buf1  g0997(.din(new_new_n777__), .dout(n3758));
  buf1  g0998(.din(new_new_n1033__), .dout(n3761));
  buf1  g0999(.din(new_new_n2375__), .dout(n3764));
  buf1  g1000(.din(new_new_n779__), .dout(n3767));
  buf1  g1001(.din(new_new_n1039__), .dout(n3770));
  buf1  g1002(.din(new_new_n1041__), .dout(n3773));
  buf1  g1003(.din(new_new_n1043__), .dout(n3776));
  buf1  g1004(.din(new_new_n781__), .dout(n3779));
  buf1  g1005(.din(new_new_n1047__), .dout(n3782));
  buf1  g1006(.din(new_new_n1049__), .dout(n3785));
  buf1  g1007(.din(new_new_n1051__), .dout(n3788));
  buf1  g1008(.din(new_new_n783__), .dout(n3791));
  buf1  g1009(.din(new_new_n1055__), .dout(n3794));
  buf1  g1010(.din(new_new_n1057__), .dout(n3797));
  buf1  g1011(.din(new_new_n1059__), .dout(n3800));
  buf1  g1012(.din(new_new_n785__), .dout(n3803));
  buf1  g1013(.din(new_new_n1063__), .dout(n3806));
  buf1  g1014(.din(new_new_n1065__), .dout(n3809));
  buf1  g1015(.din(new_new_n1067__), .dout(n3812));
  buf1  g1016(.din(new_new_n787__), .dout(n3815));
  buf1  g1017(.din(new_new_n1071__), .dout(n3818));
  buf1  g1018(.din(new_new_n1073__), .dout(n3821));
  buf1  g1019(.din(new_new_n1075__), .dout(n3824));
  buf1  g1020(.din(new_new_n789__), .dout(n3827));
  buf1  g1021(.din(new_new_n1079__), .dout(n3830));
  buf1  g1022(.din(new_new_n1081__), .dout(n3833));
  buf1  g1023(.din(new_new_n1083__), .dout(n3836));
  buf1  g1024(.din(new_new_n791__), .dout(n3839));
  buf1  g1025(.din(new_new_n1087__), .dout(n3842));
  buf1  g1026(.din(new_new_n1089__), .dout(n3845));
  buf1  g1027(.din(new_new_n1091__), .dout(n3848));
  buf1  g1028(.din(new_new_n793__), .dout(n3851));
  buf1  g1029(.din(new_new_n1095__), .dout(n3854));
  buf1  g1030(.din(new_new_n1097__), .dout(n3857));
  buf1  g1031(.din(new_new_n1099__), .dout(n3860));
  buf1  g1032(.din(new_new_n795__), .dout(n3863));
  buf1  g1033(.din(new_new_n1103__), .dout(n3866));
  buf1  g1034(.din(new_new_n1105__), .dout(n3869));
  buf1  g1035(.din(new_new_n1107__), .dout(n3872));
  buf1  g1036(.din(new_new_n797__), .dout(n3875));
  buf1  g1037(.din(new_new_n1111__), .dout(n3878));
  buf1  g1038(.din(new_new_n799__), .dout(n3881));
  buf1  g1039(.din(new_new_n1115__), .dout(n3884));
  buf1  g1040(.din(new_new_n1117__), .dout(n3887));
  buf1  g1041(.din(new_new_n1119__), .dout(n3890));
  buf1  g1042(.din(new_new_n801__), .dout(n3893));
  buf1  g1043(.din(new_new_n1165__), .dout(n3896));
  buf1  g1044(.din(new_new_n1191__), .dout(n3899));
  buf1  g1045(.din(new_new_n1219__), .dout(n3902));
  buf1  g1046(.din(new_new_n1221__), .dout(n3905));
  buf1  g1047(.din(new_new_n1223__), .dout(n3908));
  buf1  g1048(.din(new_new_n1267__), .dout(n3911));
  buf1  g1049(.din(new_new_n2385__), .dout(n3914));
  buf1  g1050(.din(new_new_n2382__), .dout(n3917));
  buf1  g1051(.din(new_new_n1265__), .dout(n3920));
  buf1  g1052(.din(new_new_n2308__), .dout(n3923));
  buf1  g1053(.din(new_new_n2231__), .dout(n3926));
  buf1  g1054(.din(new_new_n2221__), .dout(n3929));
  buf1  g1055(.din(new_new_n2241__), .dout(n3932));
  buf1  g1056(.din(new_new_n1225__), .dout(n3935));
  buf1  g1057(.din(new_new_n1227__), .dout(n3938));
  buf1  g1058(.din(new_new_n2395__), .dout(n3941));
  buf1  g1059(.din(new_new_n1245__), .dout(n3944));
  buf1  g1060(.din(new_new_n1247__), .dout(n3947));
  buf1  g1061(.din(new_new_n1249__), .dout(n3950));
  buf1  g1062(.din(new_new_n1251__), .dout(n3953));
  buf1  g1063(.din(new_new_n1253__), .dout(n3956));
  not1  g1064(.din(new_new_n2381__), .dout(n3959));
  buf1  g1065(.din(new_new_n2276__), .dout(n3962));
  buf1  g1066(.din(new_new_n2288__), .dout(n3965));
  buf1  g1067(.din(new_new_n2301__), .dout(n3968));
  buf1  g1068(.din(new_new_n2255__), .dout(n3971));
  buf1  g1069(.din(new_new_n1309__), .dout(n3974));
  buf1  g1070(.din(new_new_n1311__), .dout(n3977));
  buf1  g1071(.din(new_new_n1333__), .dout(n3980));
  buf1  g1072(.din(new_new_n1335__), .dout(n3983));
  buf1  g1073(.din(new_new_n1337__), .dout(n3986));
  buf1  g1074(.din(new_new_n1339__), .dout(n3989));
  buf1  g1075(.din(new_new_n2302__), .dout(n3992));
  buf1  g1076(.din(new_new_n2315__), .dout(n3995));
  buf1  g1077(.din(new_new_n1361__), .dout(n3998));
  buf1  g1078(.din(new_new_n2386__), .dout(n4001));
  buf1  g1079(.din(new_new_n2387__), .dout(n4004));
  buf1  g1080(.din(new_new_n2339__), .dout(n4007));
  buf1  g1081(.din(new_new_n2344__), .dout(n4010));
  buf1  g1082(.din(new_new_n2388__), .dout(n4013));
  buf1  g1083(.din(new_new_n2389__), .dout(n4016));
  buf1  g1084(.din(new_new_n2345__), .dout(n4019));
  buf1  g1085(.din(new_new_n2391__), .dout(n4022));
  buf1  g1086(.din(new_new_n2390__), .dout(n4025));
  buf1  g1087(.din(new_new_n1023__), .dout(n4028));
  buf1  g1088(.din(new_new_n1029__), .dout(n4031));
  buf1  g1089(.din(new_new_n1035__), .dout(n4034));
  not1  g1090(.din(new_new_n2319__), .dout(n4037));
  not1  g1091(.din(new_new_n2322__), .dout(n4040));
  not1  g1092(.din(new_new_n2325__), .dout(n4043));
  buf1  g1093(.din(new_new_n2329__), .dout(n4046));
  buf1  g1094(.din(new_new_n2328__), .dout(n4049));
  buf1  g1095(.din(new_new_n2332__), .dout(n4052));
  buf1  g1096(.din(new_new_n927__), .dout(n4055));
  buf1  g1097(.din(new_new_n933__), .dout(n4058));
  buf1  g1098(.din(new_new_n939__), .dout(n4061));
  not1  g1099(.din(new_new_n2424__), .dout(n4064));
  not1  g1100(.din(new_new_n2417__), .dout(n4067));
  not1  g1101(.din(new_new_n2421__), .dout(n4070));
  buf1  g1102(.din(new_new_n2413__), .dout(n4073));
  buf1  g1103(.din(new_new_n2408__), .dout(n4076));
  buf1  g1104(.din(new_new_n2410__), .dout(n4079));
  buf1  g1105(.din(new_new_n2412__), .dout(n4082));
  buf1  g1106(.din(new_new_n1391__), .dout(n4085));
  buf1  g1107(.din(new_new_n2405__), .dout(n4088));
  buf1  g1108(.din(new_new_n1017__), .dout(n4091));
  buf1  g1109(.din(new_new_n1113__), .dout(n4094));
  not1  g1110(.din(new_new_n2414__), .dout(n4097));
  not1  g1111(.din(new_new_n2418__), .dout(n4100));
  not1  g1112(.din(new_new_n2422__), .dout(n4103));
  not1  g1113(.din(new_new_n2392__), .dout(n4106));
  not1  g1114(.din(new_new_n2423__), .dout(n4109));
  not1  g1115(.din(new_new_n2416__), .dout(n4112));
  not1  g1116(.din(new_new_n2420__), .dout(n4115));
  not1  g1117(.din(new_new_n2402__), .dout(n4118));
  buf1  g1118(.din(n4088), .dout(n4121));
  buf1  g1119(.din(new_new_n2398__), .dout(n4124));
  buf1  g1120(.din(new_new_n2303__), .dout(n4127));
  buf1  g1121(.din(new_new_n1640__), .dout(n4130));
  buf1  g1122(.din(new_new_n1643__), .dout(n4133));
  buf1  g1123(.din(new_new_n1646__), .dout(n4136));
  buf1  g1124(.din(new_new_n1661__), .dout(n4139));
  buf1  g1125(.din(new_new_n1676__), .dout(n4142));
  buf1  g1126(.din(new_new_n1691__), .dout(n4145));
  buf1  g1127(.din(new_new_n1706__), .dout(n4148));
  not1  g1128(.din(new_new_n1711__), .dout(n4151));
  buf1  g1129(.din(new_new_n1724__), .dout(n4154));
  buf1  g1130(.din(new_new_n1731__), .dout(n4157));
  buf1  g1131(.din(new_new_n1744__), .dout(n4160));
  buf1  g1132(.din(new_new_n1751__), .dout(n4163));
  buf1  g1133(.din(new_new_n1754__), .dout(n4166));
  not1  g1134(.din(new_new_n2443__), .dout(n4169));
  buf1  g1135(.din(new_new_n819__), .dout(n4172));
  buf1  g1136(.din(new_new_n867__), .dout(n4175));
  buf1  g1137(.din(new_new_n999__), .dout(n4178));
  buf1  g1138(.din(new_new_n1005__), .dout(n4181));
  buf1  g1139(.din(new_new_n1011__), .dout(n4184));
  buf1  g1140(.din(new_new_n1756__), .dout(n4187));
  not1  g1141(.din(new_new_n2429__), .dout(n4190));
  buf1  g1142(.din(new_new_n1760__), .dout(n4193));
  not1  g1143(.din(new_new_n1763__), .dout(n4196));
  not1  g1144(.din(new_new_n2433__), .dout(n4199));
  not1  g1145(.din(new_new_n2430__), .dout(n4202));
  not1  g1146(.din(new_new_n1769__), .dout(n4205));
  buf1  g1147(.din(new_new_n833__), .dout(n4208));
  buf1  g1148(.din(new_new_n2440__), .dout(n4211));
  buf1  g1149(.din(new_new_n2441__), .dout(n4214));
  buf1  g1150(.din(new_new_n2442__), .dout(n4217));
  buf1  g1151(.din(new_new_n2434__), .dout(n4220));
  buf1  g1152(.din(new_new_n2435__), .dout(n4223));
  buf1  g1153(.din(new_new_n2436__), .dout(n4226));
  buf1  g1154(.din(new_new_n2439__), .dout(n4229));
  buf1  g1155(.din(n4169), .dout(n4232));
  not1  g1156(.din(new_new_n1790__), .dout(n4235));
  not1  g1157(.din(new_new_n1796__), .dout(n4238));
  not1  g1158(.din(new_new_n1802__), .dout(n4241));
  not1  g1159(.din(new_new_n1808__), .dout(n4244));
  buf1  g1160(.din(new_new_n2444__), .dout(n4247));
  buf1  g1161(.din(new_new_n943__), .dout(n4250));
  buf1  g1162(.din(new_new_n977__), .dout(n4253));
  not1  g1163(.din(new_new_n1810__), .dout(n4256));
  buf1  g1164(.din(new_new_n1811__), .dout(n4259));
  buf1  g1165(.din(new_new_n1812__), .dout(n4262));
  buf1  g1166(.din(new_new_n1813__), .dout(n4265));
  buf1  g1167(.din(new_new_n1814__), .dout(n4268));
  buf1  g1168(.din(new_new_n1815__), .dout(n4271));
  buf1  g1169(.din(new_new_n1816__), .dout(n4274));
  buf1  g1170(.din(n4247), .dout(n4277));
  buf1  g1171(.din(new_new_n761__), .dout(n4280));
  buf1  g1172(.din(new_new_n685__), .dout(n4283));
  buf1  g1173(.din(new_new_n689__), .dout(n4286));
  buf1  g1174(.din(new_new_n697__), .dout(n4289));
  buf1  g1175(.din(new_new_n703__), .dout(n4292));
  buf1  g1176(.din(new_new_n713__), .dout(n4295));
  buf1  g1177(.din(new_new_n683__), .dout(n4298));
  buf1  g1178(.din(new_new_n691__), .dout(n4301));
  buf1  g1179(.din(new_new_n699__), .dout(n4304));
  buf1  g1180(.din(new_new_n822__), .dout(new_new_n2141__));
  buf1  g1181(.din(new_new_n2141__), .dout(new_new_n2142__));
  buf1  g1182(.din(new_new_n832__), .dout(new_new_n2143__));
  buf1  g1183(.din(new_new_n2143__), .dout(new_new_n2144__));
  buf1  g1184(.din(new_new_n830__), .dout(new_new_n2145__));
  buf1  g1185(.din(new_new_n1401__), .dout(new_new_n2146__));
  buf1  g1186(.din(new_new_n870__), .dout(new_new_n2147__));
  buf1  g1187(.din(new_new_n804__), .dout(new_new_n2148__));
  buf1  g1188(.din(new_new_n814__), .dout(new_new_n2149__));
  buf1  g1189(.din(new_new_n816__), .dout(new_new_n2150__));
  buf1  g1190(.din(new_new_n1403__), .dout(new_new_n2151__));
  buf1  g1191(.din(new_new_n2151__), .dout(new_new_n2152__));
  buf1  g1192(.din(new_new_n836__), .dout(new_new_n2153__));
  buf1  g1193(.din(new_new_n1417__), .dout(new_new_n2154__));
  buf1  g1194(.din(new_new_n1420__), .dout(new_new_n2155__));
  buf1  g1195(.din(new_new_n844__), .dout(new_new_n2156__));
  buf1  g1196(.din(new_new_n1168__), .dout(new_new_n2157__));
  buf1  g1197(.din(new_new_n1287__), .dout(new_new_n2158__));
  buf1  g1198(.din(new_new_n963__), .dout(new_new_n2159__));
  buf1  g1199(.din(new_new_n2159__), .dout(new_new_n2160__));
  buf1  g1200(.din(new_new_n2159__), .dout(new_new_n2161__));
  buf1  g1201(.din(new_new_n1288__), .dout(new_new_n2162__));
  buf1  g1202(.din(new_new_n964__), .dout(new_new_n2163__));
  buf1  g1203(.din(new_new_n2163__), .dout(new_new_n2164__));
  buf1  g1204(.din(new_new_n2163__), .dout(new_new_n2165__));
  buf1  g1205(.din(new_new_n1289__), .dout(new_new_n2166__));
  buf1  g1206(.din(new_new_n971__), .dout(new_new_n2167__));
  buf1  g1207(.din(new_new_n1290__), .dout(new_new_n2168__));
  buf1  g1208(.din(new_new_n972__), .dout(new_new_n2169__));
  buf1  g1209(.din(new_new_n1291__), .dout(new_new_n2170__));
  buf1  g1210(.din(new_new_n1292__), .dout(new_new_n2171__));
  buf1  g1211(.din(new_new_n1293__), .dout(new_new_n2172__));
  buf1  g1212(.din(new_new_n1045__), .dout(new_new_n2173__));
  buf1  g1213(.din(new_new_n1294__), .dout(new_new_n2174__));
  buf1  g1214(.din(new_new_n1046__), .dout(new_new_n2175__));
  buf1  g1215(.din(new_new_n1054__), .dout(new_new_n2176__));
  buf1  g1216(.din(new_new_n2176__), .dout(new_new_n2177__));
  buf1  g1217(.din(new_new_n2177__), .dout(new_new_n2178__));
  buf1  g1218(.din(new_new_n2177__), .dout(new_new_n2179__));
  buf1  g1219(.din(new_new_n2176__), .dout(new_new_n2180__));
  buf1  g1220(.din(new_new_n2180__), .dout(new_new_n2181__));
  buf1  g1221(.din(new_new_n2180__), .dout(new_new_n2182__));
  buf1  g1222(.din(new_new_n1062__), .dout(new_new_n2183__));
  buf1  g1223(.din(new_new_n2183__), .dout(new_new_n2184__));
  buf1  g1224(.din(new_new_n2184__), .dout(new_new_n2185__));
  buf1  g1225(.din(new_new_n2184__), .dout(new_new_n2186__));
  buf1  g1226(.din(new_new_n2183__), .dout(new_new_n2187__));
  buf1  g1227(.din(new_new_n2187__), .dout(new_new_n2188__));
  buf1  g1228(.din(new_new_n2187__), .dout(new_new_n2189__));
  buf1  g1229(.din(new_new_n1070__), .dout(new_new_n2190__));
  buf1  g1230(.din(new_new_n2190__), .dout(new_new_n2191__));
  buf1  g1231(.din(new_new_n2191__), .dout(new_new_n2192__));
  buf1  g1232(.din(new_new_n2191__), .dout(new_new_n2193__));
  buf1  g1233(.din(new_new_n2190__), .dout(new_new_n2194__));
  buf1  g1234(.din(new_new_n2194__), .dout(new_new_n2195__));
  buf1  g1235(.din(new_new_n2194__), .dout(new_new_n2196__));
  buf1  g1236(.din(new_new_n1078__), .dout(new_new_n2197__));
  buf1  g1237(.din(new_new_n2197__), .dout(new_new_n2198__));
  buf1  g1238(.din(new_new_n2198__), .dout(new_new_n2199__));
  buf1  g1239(.din(new_new_n2198__), .dout(new_new_n2200__));
  buf1  g1240(.din(new_new_n2197__), .dout(new_new_n2201__));
  buf1  g1241(.din(new_new_n2201__), .dout(new_new_n2202__));
  buf1  g1242(.din(new_new_n2201__), .dout(new_new_n2203__));
  buf1  g1243(.din(new_new_n1094__), .dout(new_new_n2204__));
  buf1  g1244(.din(new_new_n2204__), .dout(new_new_n2205__));
  buf1  g1245(.din(new_new_n1086__), .dout(new_new_n2206__));
  buf1  g1246(.din(new_new_n2206__), .dout(new_new_n2207__));
  buf1  g1247(.din(new_new_n2207__), .dout(new_new_n2208__));
  buf1  g1248(.din(new_new_n2207__), .dout(new_new_n2209__));
  buf1  g1249(.din(new_new_n2206__), .dout(new_new_n2210__));
  buf1  g1250(.din(new_new_n2210__), .dout(new_new_n2211__));
  buf1  g1251(.din(new_new_n2210__), .dout(new_new_n2212__));
  buf1  g1252(.din(new_new_n1296__), .dout(new_new_n2213__));
  buf1  g1253(.din(new_new_n2213__), .dout(new_new_n2214__));
  buf1  g1254(.din(new_new_n2214__), .dout(new_new_n2215__));
  buf1  g1255(.din(new_new_n2214__), .dout(new_new_n2216__));
  buf1  g1256(.din(new_new_n2213__), .dout(new_new_n2217__));
  buf1  g1257(.din(new_new_n2217__), .dout(new_new_n2218__));
  buf1  g1258(.din(new_new_n2217__), .dout(new_new_n2219__));
  buf1  g1259(.din(new_new_n1280__), .dout(new_new_n2220__));
  buf1  g1260(.din(new_new_n1353__), .dout(new_new_n2221__));
  buf1  g1261(.din(new_new_n2221__), .dout(new_new_n2222__));
  buf1  g1262(.din(new_new_n1313__), .dout(new_new_n2223__));
  buf1  g1263(.din(new_new_n2223__), .dout(new_new_n2224__));
  buf1  g1264(.din(new_new_n2224__), .dout(new_new_n2225__));
  buf1  g1265(.din(new_new_n2223__), .dout(new_new_n2226__));
  buf1  g1266(.din(new_new_n1354__), .dout(new_new_n2227__));
  buf1  g1267(.din(new_new_n1314__), .dout(new_new_n2228__));
  buf1  g1268(.din(new_new_n2228__), .dout(new_new_n2229__));
  buf1  g1269(.din(new_new_n2228__), .dout(new_new_n2230__));
  buf1  g1270(.din(new_new_n1355__), .dout(new_new_n2231__));
  buf1  g1271(.din(new_new_n2231__), .dout(new_new_n2232__));
  buf1  g1272(.din(new_new_n1315__), .dout(new_new_n2233__));
  buf1  g1273(.din(new_new_n2233__), .dout(new_new_n2234__));
  buf1  g1274(.din(new_new_n2234__), .dout(new_new_n2235__));
  buf1  g1275(.din(new_new_n2233__), .dout(new_new_n2236__));
  buf1  g1276(.din(new_new_n1356__), .dout(new_new_n2237__));
  buf1  g1277(.din(new_new_n1316__), .dout(new_new_n2238__));
  buf1  g1278(.din(new_new_n2238__), .dout(new_new_n2239__));
  buf1  g1279(.din(new_new_n2238__), .dout(new_new_n2240__));
  buf1  g1280(.din(new_new_n1357__), .dout(new_new_n2241__));
  buf1  g1281(.din(new_new_n2241__), .dout(new_new_n2242__));
  buf1  g1282(.din(new_new_n1317__), .dout(new_new_n2243__));
  buf1  g1283(.din(new_new_n2243__), .dout(new_new_n2244__));
  buf1  g1284(.din(new_new_n2244__), .dout(new_new_n2245__));
  buf1  g1285(.din(new_new_n2243__), .dout(new_new_n2246__));
  buf1  g1286(.din(new_new_n1358__), .dout(new_new_n2247__));
  buf1  g1287(.din(new_new_n1318__), .dout(new_new_n2248__));
  buf1  g1288(.din(new_new_n2248__), .dout(new_new_n2249__));
  buf1  g1289(.din(new_new_n2248__), .dout(new_new_n2250__));
  buf1  g1290(.din(new_new_n1568__), .dout(new_new_n2251__));
  buf1  g1291(.din(new_new_n994__), .dout(new_new_n2252__));
  buf1  g1292(.din(new_new_n2252__), .dout(new_new_n2253__));
  buf1  g1293(.din(new_new_n2252__), .dout(new_new_n2254__));
  buf1  g1294(.din(new_new_n1569__), .dout(new_new_n2255__));
  buf1  g1295(.din(new_new_n2255__), .dout(new_new_n2256__));
  buf1  g1296(.din(new_new_n993__), .dout(new_new_n2257__));
  buf1  g1297(.din(new_new_n2257__), .dout(new_new_n2258__));
  buf1  g1298(.din(new_new_n2258__), .dout(new_new_n2259__));
  buf1  g1299(.din(new_new_n2257__), .dout(new_new_n2260__));
  buf1  g1300(.din(new_new_n1261__), .dout(new_new_n2261__));
  buf1  g1301(.din(new_new_n2261__), .dout(new_new_n2262__));
  buf1  g1302(.din(new_new_n1262__), .dout(new_new_n2263__));
  buf1  g1303(.din(new_new_n2263__), .dout(new_new_n2264__));
  buf1  g1304(.din(new_new_n1263__), .dout(new_new_n2265__));
  buf1  g1305(.din(new_new_n2265__), .dout(new_new_n2266__));
  buf1  g1306(.din(new_new_n1264__), .dout(new_new_n2267__));
  buf1  g1307(.din(new_new_n2267__), .dout(new_new_n2268__));
  buf1  g1308(.din(new_new_n1331__), .dout(new_new_n2269__));
  buf1  g1309(.din(new_new_n1332__), .dout(new_new_n2270__));
  buf1  g1310(.din(new_new_n1581__), .dout(new_new_n2271__));
  buf1  g1311(.din(new_new_n2271__), .dout(new_new_n2272__));
  buf1  g1312(.din(new_new_n1559__), .dout(new_new_n2273__));
  buf1  g1313(.din(new_new_n1580__), .dout(new_new_n2274__));
  buf1  g1314(.din(new_new_n2274__), .dout(new_new_n2275__));
  buf1  g1315(.din(new_new_n1558__), .dout(new_new_n2276__));
  buf1  g1316(.din(new_new_n2276__), .dout(new_new_n2277__));
  buf1  g1317(.din(new_new_n1585__), .dout(new_new_n2278__));
  buf1  g1318(.din(new_new_n2278__), .dout(new_new_n2279__));
  buf1  g1319(.din(new_new_n2278__), .dout(new_new_n2280__));
  buf1  g1320(.din(new_new_n1561__), .dout(new_new_n2281__));
  buf1  g1321(.din(new_new_n2281__), .dout(new_new_n2282__));
  buf1  g1322(.din(new_new_n1584__), .dout(new_new_n2283__));
  buf1  g1323(.din(new_new_n2283__), .dout(new_new_n2284__));
  buf1  g1324(.din(new_new_n2283__), .dout(new_new_n2285__));
  buf1  g1325(.din(new_new_n1560__), .dout(new_new_n2286__));
  buf1  g1326(.din(new_new_n2286__), .dout(new_new_n2287__));
  buf1  g1327(.din(new_new_n2286__), .dout(new_new_n2288__));
  buf1  g1328(.din(new_new_n1589__), .dout(new_new_n2289__));
  buf1  g1329(.din(new_new_n2289__), .dout(new_new_n2290__));
  buf1  g1330(.din(new_new_n2289__), .dout(new_new_n2291__));
  buf1  g1331(.din(new_new_n1563__), .dout(new_new_n2292__));
  buf1  g1332(.din(new_new_n2292__), .dout(new_new_n2293__));
  buf1  g1333(.din(new_new_n2292__), .dout(new_new_n2294__));
  buf1  g1334(.din(new_new_n1588__), .dout(new_new_n2295__));
  buf1  g1335(.din(new_new_n2295__), .dout(new_new_n2296__));
  buf1  g1336(.din(new_new_n2295__), .dout(new_new_n2297__));
  buf1  g1337(.din(new_new_n1562__), .dout(new_new_n2298__));
  buf1  g1338(.din(new_new_n2298__), .dout(new_new_n2299__));
  buf1  g1339(.din(new_new_n2299__), .dout(new_new_n2300__));
  buf1  g1340(.din(new_new_n2298__), .dout(new_new_n2301__));
  buf1  g1341(.din(new_new_n1571__), .dout(new_new_n2302__));
  buf1  g1342(.din(new_new_n1592__), .dout(new_new_n2303__));
  buf1  g1343(.din(new_new_n1598__), .dout(new_new_n2304__));
  buf1  g1344(.din(new_new_n1599__), .dout(new_new_n2305__));
  buf1  g1345(.din(new_new_n1351__), .dout(new_new_n2306__));
  buf1  g1346(.din(new_new_n1352__), .dout(new_new_n2307__));
  buf1  g1347(.din(new_new_n1349__), .dout(new_new_n2308__));
  buf1  g1348(.din(new_new_n1605__), .dout(new_new_n2309__));
  buf1  g1349(.din(new_new_n2309__), .dout(new_new_n2310__));
  buf1  g1350(.din(new_new_n2309__), .dout(new_new_n2311__));
  buf1  g1351(.din(new_new_n1604__), .dout(new_new_n2312__));
  buf1  g1352(.din(new_new_n2312__), .dout(new_new_n2313__));
  buf1  g1353(.din(new_new_n2312__), .dout(new_new_n2314__));
  buf1  g1354(.din(new_new_n1379__), .dout(new_new_n2315__));
  buf1  g1355(.din(new_new_n1616__), .dout(new_new_n2316__));
  buf1  g1356(.din(new_new_n2316__), .dout(new_new_n2317__));
  buf1  g1357(.din(new_new_n2316__), .dout(new_new_n2318__));
  buf1  g1358(.din(new_new_n1618__), .dout(new_new_n2319__));
  buf1  g1359(.din(new_new_n2319__), .dout(new_new_n2320__));
  buf1  g1360(.din(new_new_n1024__), .dout(new_new_n2321__));
  buf1  g1361(.din(new_new_n1620__), .dout(new_new_n2322__));
  buf1  g1362(.din(new_new_n2322__), .dout(new_new_n2323__));
  buf1  g1363(.din(new_new_n1030__), .dout(new_new_n2324__));
  buf1  g1364(.din(new_new_n1622__), .dout(new_new_n2325__));
  buf1  g1365(.din(new_new_n2325__), .dout(new_new_n2326__));
  buf1  g1366(.din(new_new_n1036__), .dout(new_new_n2327__));
  buf1  g1367(.din(new_new_n1395__), .dout(new_new_n2328__));
  buf1  g1368(.din(new_new_n1393__), .dout(new_new_n2329__));
  buf1  g1369(.din(new_new_n2329__), .dout(new_new_n2330__));
  buf1  g1370(.din(new_new_n1394__), .dout(new_new_n2331__));
  buf1  g1371(.din(new_new_n1397__), .dout(new_new_n2332__));
  buf1  g1372(.din(new_new_n2332__), .dout(new_new_n2333__));
  buf1  g1373(.din(new_new_n1364__), .dout(new_new_n2334__));
  buf1  g1374(.din(new_new_n1348__), .dout(new_new_n2335__));
  buf1  g1375(.din(new_new_n2335__), .dout(new_new_n2336__));
  buf1  g1376(.din(new_new_n2335__), .dout(new_new_n2337__));
  buf1  g1377(.din(new_new_n1390__), .dout(new_new_n2338__));
  buf1  g1378(.din(new_new_n1576__), .dout(new_new_n2339__));
  buf1  g1379(.din(new_new_n1257__), .dout(new_new_n2340__));
  buf1  g1380(.din(new_new_n2340__), .dout(new_new_n2341__));
  buf1  g1381(.din(new_new_n1258__), .dout(new_new_n2342__));
  buf1  g1382(.din(new_new_n2342__), .dout(new_new_n2343__));
  buf1  g1383(.din(new_new_n1578__), .dout(new_new_n2344__));
  buf1  g1384(.din(new_new_n1590__), .dout(new_new_n2345__));
  buf1  g1385(.din(new_new_n1277__), .dout(new_new_n2346__));
  buf1  g1386(.din(new_new_n2346__), .dout(new_new_n2347__));
  buf1  g1387(.din(new_new_n1231__), .dout(new_new_n2348__));
  buf1  g1388(.din(new_new_n2348__), .dout(new_new_n2349__));
  buf1  g1389(.din(new_new_n1278__), .dout(new_new_n2350__));
  buf1  g1390(.din(new_new_n1232__), .dout(new_new_n2351__));
  buf1  g1391(.din(new_new_n1235__), .dout(new_new_n2352__));
  buf1  g1392(.din(new_new_n2352__), .dout(new_new_n2353__));
  buf1  g1393(.din(new_new_n1233__), .dout(new_new_n2354__));
  buf1  g1394(.din(new_new_n2354__), .dout(new_new_n2355__));
  buf1  g1395(.din(new_new_n1236__), .dout(new_new_n2356__));
  buf1  g1396(.din(new_new_n1234__), .dout(new_new_n2357__));
  buf1  g1397(.din(new_new_n1193__), .dout(new_new_n2358__));
  buf1  g1398(.din(new_new_n2358__), .dout(new_new_n2359__));
  buf1  g1399(.din(new_new_n1183__), .dout(new_new_n2360__));
  buf1  g1400(.din(new_new_n2360__), .dout(new_new_n2361__));
  buf1  g1401(.din(new_new_n1194__), .dout(new_new_n2362__));
  buf1  g1402(.din(new_new_n1184__), .dout(new_new_n2363__));
  buf1  g1403(.din(new_new_n1187__), .dout(new_new_n2364__));
  buf1  g1404(.din(new_new_n1185__), .dout(new_new_n2365__));
  buf1  g1405(.din(new_new_n2365__), .dout(new_new_n2366__));
  buf1  g1406(.din(new_new_n1188__), .dout(new_new_n2367__));
  buf1  g1407(.din(new_new_n1186__), .dout(new_new_n2368__));
  buf1  g1408(.din(new_new_n1255__), .dout(new_new_n2369__));
  buf1  g1409(.din(new_new_n2369__), .dout(new_new_n2370__));
  buf1  g1410(.din(new_new_n1213__), .dout(new_new_n2371__));
  buf1  g1411(.din(new_new_n2371__), .dout(new_new_n2372__));
  buf1  g1412(.din(new_new_n1256__), .dout(new_new_n2373__));
  buf1  g1413(.din(new_new_n1214__), .dout(new_new_n2374__));
  buf1  g1414(.din(new_new_n1217__), .dout(new_new_n2375__));
  buf1  g1415(.din(new_new_n2375__), .dout(new_new_n2376__));
  buf1  g1416(.din(new_new_n1215__), .dout(new_new_n2377__));
  buf1  g1417(.din(new_new_n2377__), .dout(new_new_n2378__));
  buf1  g1418(.din(new_new_n1218__), .dout(new_new_n2379__));
  buf1  g1419(.din(new_new_n1216__), .dout(new_new_n2380__));
  buf1  g1420(.din(new_new_n1557__), .dout(new_new_n2381__));
  buf1  g1421(.din(new_new_n1271__), .dout(new_new_n2382__));
  buf1  g1422(.din(new_new_n2382__), .dout(new_new_n2383__));
  buf1  g1423(.din(new_new_n1272__), .dout(new_new_n2384__));
  buf1  g1424(.din(new_new_n1269__), .dout(new_new_n2385__));
  buf1  g1425(.din(new_new_n1572__), .dout(new_new_n2386__));
  buf1  g1426(.din(new_new_n1574__), .dout(new_new_n2387__));
  buf1  g1427(.din(new_new_n1582__), .dout(new_new_n2388__));
  buf1  g1428(.din(new_new_n1586__), .dout(new_new_n2389__));
  buf1  g1429(.din(new_new_n1615__), .dout(new_new_n2390__));
  buf1  g1430(.din(new_new_n1594__), .dout(new_new_n2391__));
  buf1  g1431(.din(new_new_n1636__), .dout(new_new_n2392__));
  buf1  g1432(.din(new_new_n2392__), .dout(new_new_n2393__));
  buf1  g1433(.din(new_new_n1018__), .dout(new_new_n2394__));
  buf1  g1434(.din(new_new_n1243__), .dout(new_new_n2395__));
  buf1  g1435(.din(new_new_n1276__), .dout(new_new_n2396__));
  buf1  g1436(.din(new_new_n1246__), .dout(new_new_n2397__));
  buf1  g1437(.din(new_new_n921__), .dout(new_new_n2398__));
  buf1  g1438(.din(new_new_n1762__), .dout(new_new_n2399__));
  buf1  g1439(.din(new_new_n2399__), .dout(new_new_n2400__));
  buf1  g1440(.din(new_new_n2399__), .dout(new_new_n2401__));
  buf1  g1441(.din(new_new_n1637__), .dout(new_new_n2402__));
  buf1  g1442(.din(new_new_n1628__), .dout(new_new_n2403__));
  buf1  g1443(.din(new_new_n2403__), .dout(new_new_n2404__));
  buf1  g1444(.din(new_new_n2403__), .dout(new_new_n2405__));
  buf1  g1445(.din(new_new_n1385__), .dout(new_new_n2406__));
  buf1  g1446(.din(new_new_n2406__), .dout(new_new_n2407__));
  buf1  g1447(.din(new_new_n2406__), .dout(new_new_n2408__));
  buf1  g1448(.din(new_new_n1392__), .dout(new_new_n2409__));
  buf1  g1449(.din(new_new_n1387__), .dout(new_new_n2410__));
  buf1  g1450(.din(new_new_n1388__), .dout(new_new_n2411__));
  buf1  g1451(.din(new_new_n1389__), .dout(new_new_n2412__));
  buf1  g1452(.din(new_new_n1383__), .dout(new_new_n2413__));
  buf1  g1453(.din(new_new_n1630__), .dout(new_new_n2414__));
  buf1  g1454(.din(new_new_n2414__), .dout(new_new_n2415__));
  buf1  g1455(.din(new_new_n1624__), .dout(new_new_n2416__));
  buf1  g1456(.din(new_new_n2416__), .dout(new_new_n2417__));
  buf1  g1457(.din(new_new_n1631__), .dout(new_new_n2418__));
  buf1  g1458(.din(new_new_n1784__), .dout(new_new_n2419__));
  buf1  g1459(.din(new_new_n1625__), .dout(new_new_n2420__));
  buf1  g1460(.din(new_new_n2420__), .dout(new_new_n2421__));
  buf1  g1461(.din(new_new_n1632__), .dout(new_new_n2422__));
  buf1  g1462(.din(new_new_n1623__), .dout(new_new_n2423__));
  buf1  g1463(.din(new_new_n2423__), .dout(new_new_n2424__));
  buf1  g1464(.din(new_new_n976__), .dout(new_new_n2425__));
  buf1  g1465(.din(new_new_n2425__), .dout(new_new_n2426__));
  buf1  g1466(.din(new_new_n1759__), .dout(new_new_n2427__));
  buf1  g1467(.din(new_new_n2427__), .dout(new_new_n2428__));
  buf1  g1468(.din(new_new_n2427__), .dout(new_new_n2429__));
  buf1  g1469(.din(new_new_n1768__), .dout(new_new_n2430__));
  buf1  g1470(.din(new_new_n1766__), .dout(new_new_n2431__));
  buf1  g1471(.din(new_new_n2431__), .dout(new_new_n2432__));
  buf1  g1472(.din(new_new_n2431__), .dout(new_new_n2433__));
  buf1  g1473(.din(new_new_n979__), .dout(new_new_n2434__));
  buf1  g1474(.din(new_new_n981__), .dout(new_new_n2435__));
  buf1  g1475(.din(new_new_n987__), .dout(new_new_n2436__));
  buf1  g1476(.din(new_new_n1782__), .dout(new_new_n2437__));
  buf1  g1477(.din(new_new_n2437__), .dout(new_new_n2438__));
  buf1  g1478(.din(new_new_n2437__), .dout(new_new_n2439__));
  buf1  g1479(.din(new_new_n947__), .dout(new_new_n2440__));
  buf1  g1480(.din(new_new_n951__), .dout(new_new_n2441__));
  buf1  g1481(.din(new_new_n955__), .dout(new_new_n2442__));
  buf1  g1482(.din(new_new_n1755__), .dout(new_new_n2443__));
  buf1  g1483(.din(new_new_n1123__), .dout(new_new_n2444__));
  always @ (posedge clock) begin
    n480_lo <= n3413;
    n492_lo <= n3416;
    n495_lo <= n3419;
    n498_lo <= n3422;
    n501_lo <= n3425;
    n504_lo <= n3428;
    n516_lo <= n3431;
    n528_lo <= n3434;
    n531_lo <= n3437;
    n540_lo <= n3440;
    n543_lo <= n3443;
    n546_lo <= n3446;
    n549_lo <= n3449;
    n552_lo <= n3452;
    n564_lo <= n3455;
    n579_lo <= n3458;
    n600_lo <= n3461;
    n603_lo <= n3464;
    n606_lo <= n3467;
    n609_lo <= n3470;
    n612_lo <= n3473;
    n615_lo <= n3476;
    n618_lo <= n3479;
    n621_lo <= n3482;
    n627_lo <= n3485;
    n630_lo <= n3488;
    n633_lo <= n3491;
    n639_lo <= n3494;
    n642_lo <= n3497;
    n645_lo <= n3500;
    n648_lo <= n3503;
    n660_lo <= n3506;
    n663_lo <= n3509;
    n672_lo <= n3512;
    n675_lo <= n3515;
    n678_lo <= n3518;
    n681_lo <= n3521;
    n684_lo <= n3524;
    n687_lo <= n3527;
    n690_lo <= n3530;
    n693_lo <= n3533;
    n696_lo <= n3536;
    n699_lo <= n3539;
    n702_lo <= n3542;
    n705_lo <= n3545;
    n708_lo <= n3548;
    n711_lo <= n3551;
    n714_lo <= n3554;
    n717_lo <= n3557;
    n720_lo <= n3560;
    n723_lo <= n3563;
    n726_lo <= n3566;
    n729_lo <= n3569;
    n732_lo <= n3572;
    n735_lo <= n3575;
    n738_lo <= n3578;
    n741_lo <= n3581;
    n744_lo <= n3584;
    n747_lo <= n3587;
    n750_lo <= n3590;
    n756_lo <= n3593;
    n759_lo <= n3596;
    n762_lo <= n3599;
    n768_lo <= n3602;
    n771_lo <= n3605;
    n774_lo <= n3608;
    n780_lo <= n3611;
    n783_lo <= n3614;
    n786_lo <= n3617;
    n792_lo <= n3620;
    n795_lo <= n3623;
    n804_lo <= n3626;
    n807_lo <= n3629;
    n816_lo <= n3632;
    n819_lo <= n3635;
    n828_lo <= n3638;
    n831_lo <= n3641;
    n843_lo <= n3644;
    n846_lo <= n3647;
    n849_lo <= n3650;
    n852_lo <= n3653;
    n855_lo <= n3656;
    n858_lo <= n3659;
    n861_lo <= n3662;
    n864_lo <= n3665;
    n867_lo <= n3668;
    n870_lo <= n3671;
    n879_lo <= n3674;
    n891_lo <= n3677;
    n903_lo <= n3680;
    n915_lo <= n3683;
    n918_lo <= n3686;
    n927_lo <= n3689;
    n951_lo <= n3692;
    n954_lo <= n3695;
    n957_lo <= n3698;
    n960_lo <= n3701;
    n963_lo <= n3704;
    n966_lo <= n3707;
    n972_lo <= n3710;
    n975_lo <= n3713;
    n978_lo <= n3716;
    n984_lo <= n3719;
    n987_lo <= n3722;
    n990_lo <= n3725;
    n996_lo <= n3728;
    n999_lo <= n3731;
    n1002_lo <= n3734;
    n1008_lo <= n3737;
    n1011_lo <= n3740;
    n1014_lo <= n3743;
    n1020_lo <= n3746;
    n1023_lo <= n3749;
    n1026_lo <= n3752;
    n1032_lo <= n3755;
    n1035_lo <= n3758;
    n1038_lo <= n3761;
    n1044_lo <= n3764;
    n1047_lo <= n3767;
    n1050_lo <= n3770;
    n1053_lo <= n3773;
    n1056_lo <= n3776;
    n1059_lo <= n3779;
    n1062_lo <= n3782;
    n1065_lo <= n3785;
    n1068_lo <= n3788;
    n1071_lo <= n3791;
    n1074_lo <= n3794;
    n1077_lo <= n3797;
    n1080_lo <= n3800;
    n1083_lo <= n3803;
    n1086_lo <= n3806;
    n1089_lo <= n3809;
    n1092_lo <= n3812;
    n1095_lo <= n3815;
    n1098_lo <= n3818;
    n1101_lo <= n3821;
    n1104_lo <= n3824;
    n1107_lo <= n3827;
    n1110_lo <= n3830;
    n1113_lo <= n3833;
    n1116_lo <= n3836;
    n1119_lo <= n3839;
    n1122_lo <= n3842;
    n1125_lo <= n3845;
    n1128_lo <= n3848;
    n1131_lo <= n3851;
    n1134_lo <= n3854;
    n1137_lo <= n3857;
    n1140_lo <= n3860;
    n1143_lo <= n3863;
    n1146_lo <= n3866;
    n1149_lo <= n3869;
    n1152_lo <= n3872;
    n1155_lo <= n3875;
    n1158_lo <= n3878;
    n1167_lo <= n3881;
    n1170_lo <= n3884;
    n1173_lo <= n3887;
    n1176_lo <= n3890;
    n1179_lo <= n3893;
    n1529_o2 <= n3896;
    n1616_o2 <= n3899;
    n1655_o2 <= n3902;
    n1656_o2 <= n3905;
    n1657_o2 <= n3908;
    n1730_o2 <= n3911;
    n1731_o2 <= n3914;
    n1732_o2 <= n3917;
    n1729_o2 <= n3920;
    n1805_o2 <= n3923;
    n1808_o2 <= n3926;
    n1807_o2 <= n3929;
    n1809_o2 <= n3932;
    n1663_o2 <= n3935;
    n1664_o2 <= n3938;
    n1704_o2 <= n3941;
    n1705_o2 <= n3944;
    n1706_o2 <= n3947;
    n1707_o2 <= n3950;
    n1708_o2 <= n3953;
    n1709_o2 <= n3956;
    G280_o2 <= n3959;
    G655_o2 <= n3962;
    G663_o2 <= n3965;
    G672_o2 <= n3968;
    G538_o2 <= n3971;
    n1780_o2 <= n3974;
    n1781_o2 <= n3977;
    n1797_o2 <= n3980;
    n1798_o2 <= n3983;
    n1799_o2 <= n3986;
    n1800_o2 <= n3989;
    G578_o2 <= n3992;
    n1828_o2 <= n3995;
    n801_lo_buf_o2 <= n3998;
    G693_o2 <= n4001;
    G702_o2 <= n4004;
    G712_o2 <= n4007;
    G685_o2 <= n4010;
    G658_o2 <= n4013;
    G667_o2 <= n4016;
    G677_o2 <= n4019;
    G650_o2 <= n4022;
    G798_o2 <= n4025;
    n1017_lo_buf_o2 <= n4028;
    n1029_lo_buf_o2 <= n4031;
    n1041_lo_buf_o2 <= n4034;
    G558_o2 <= n4037;
    G562_o2 <= n4040;
    G566_o2 <= n4043;
    n1835_o2 <= n4046;
    n1836_o2 <= n4049;
    n1837_o2 <= n4052;
    n765_lo_buf_o2 <= n4055;
    n777_lo_buf_o2 <= n4058;
    n789_lo_buf_o2 <= n4061;
    G617_o2 <= n4064;
    G626_o2 <= n4067;
    G636_o2 <= n4070;
    n489_lo_buf_o2 <= n4073;
    n513_lo_buf_o2 <= n4076;
    n561_lo_buf_o2 <= n4079;
    n597_lo_buf_o2 <= n4082;
    n657_lo_buf_o2 <= n4085;
    G276_o2 <= n4088;
    n1005_lo_buf_o2 <= n4091;
    n1161_lo_buf_o2 <= n4094;
    G620_o2 <= n4097;
    G629_o2 <= n4100;
    G639_o2 <= n4103;
    G554_o2 <= n4106;
    G690_o2 <= n4109;
    G698_o2 <= n4112;
    G707_o2 <= n4115;
    G319_o2 <= n4118;
    G389_o2 <= n4121;
    n753_lo_buf_o2 <= n4124;
    G647_o2 <= n4127;
    G769_o2 <= n4130;
    G785_o2 <= n4133;
    G808_o2 <= n4136;
    G445_o2 <= n4139;
    G448_o2 <= n4142;
    G477_o2 <= n4145;
    G480_o2 <= n4148;
    G436_o2 <= n4151;
    G786_o2 <= n4154;
    G787_o2 <= n4157;
    G826_o2 <= n4160;
    G827_o2 <= n4163;
    G825_o2 <= n4166;
    G610_o2 <= n4169;
    n537_lo_buf_o2 <= n4172;
    n669_lo_buf_o2 <= n4175;
    n969_lo_buf_o2 <= n4178;
    n981_lo_buf_o2 <= n4181;
    n993_lo_buf_o2 <= n4184;
    G309_o2 <= n4187;
    G461_o2 <= n4190;
    G487_o2 <= n4193;
    G460_o2 <= n4196;
    G468_o2 <= n4199;
    G287_o2 <= n4202;
    G613_o2 <= n4205;
    n585_lo_buf_o2 <= n4208;
    n813_lo_buf_o2 <= n4211;
    n825_lo_buf_o2 <= n4214;
    n837_lo_buf_o2 <= n4217;
    n897_lo_buf_o2 <= n4220;
    n909_lo_buf_o2 <= n4223;
    n933_lo_buf_o2 <= n4226;
    G451_o2 <= n4229;
    G682_o2 <= n4232;
    G756_o2 <= n4235;
    G542_o2 <= n4238;
    G546_o2 <= n4241;
    G550_o2 <= n4244;
    G310_o2 <= n4247;
    n798_lo_buf_o2 <= n4250;
    n882_lo_buf_o2 <= n4253;
    G427_o2 <= n4256;
    G497_o2 <= n4259;
    G499_o2 <= n4262;
    G501_o2 <= n4265;
    G498_o2 <= n4268;
    G500_o2 <= n4271;
    G502_o2 <= n4274;
    G369_o2 <= n4277;
    n939_lo_buf_o2 <= n4280;
    n486_lo_buf_o2 <= n4283;
    n510_lo_buf_o2 <= n4286;
    n558_lo_buf_o2 <= n4289;
    n594_lo_buf_o2 <= n4292;
    n654_lo_buf_o2 <= n4295;
    n477_lo_buf_o2 <= n4298;
    n525_lo_buf_o2 <= n4301;
    n573_lo_buf_o2 <= n4304;
  end
  initial begin
    n480_lo <= 1'b0;
    n492_lo <= 1'b0;
    n495_lo <= 1'b0;
    n498_lo <= 1'b0;
    n501_lo <= 1'b0;
    n504_lo <= 1'b0;
    n516_lo <= 1'b0;
    n528_lo <= 1'b0;
    n531_lo <= 1'b0;
    n540_lo <= 1'b0;
    n543_lo <= 1'b0;
    n546_lo <= 1'b0;
    n549_lo <= 1'b0;
    n552_lo <= 1'b0;
    n564_lo <= 1'b0;
    n579_lo <= 1'b0;
    n600_lo <= 1'b0;
    n603_lo <= 1'b0;
    n606_lo <= 1'b0;
    n609_lo <= 1'b0;
    n612_lo <= 1'b0;
    n615_lo <= 1'b0;
    n618_lo <= 1'b0;
    n621_lo <= 1'b0;
    n627_lo <= 1'b0;
    n630_lo <= 1'b0;
    n633_lo <= 1'b0;
    n639_lo <= 1'b0;
    n642_lo <= 1'b0;
    n645_lo <= 1'b0;
    n648_lo <= 1'b0;
    n660_lo <= 1'b0;
    n663_lo <= 1'b0;
    n672_lo <= 1'b0;
    n675_lo <= 1'b0;
    n678_lo <= 1'b0;
    n681_lo <= 1'b0;
    n684_lo <= 1'b0;
    n687_lo <= 1'b0;
    n690_lo <= 1'b0;
    n693_lo <= 1'b0;
    n696_lo <= 1'b0;
    n699_lo <= 1'b0;
    n702_lo <= 1'b0;
    n705_lo <= 1'b0;
    n708_lo <= 1'b0;
    n711_lo <= 1'b0;
    n714_lo <= 1'b0;
    n717_lo <= 1'b0;
    n720_lo <= 1'b0;
    n723_lo <= 1'b0;
    n726_lo <= 1'b0;
    n729_lo <= 1'b0;
    n732_lo <= 1'b0;
    n735_lo <= 1'b0;
    n738_lo <= 1'b0;
    n741_lo <= 1'b0;
    n744_lo <= 1'b0;
    n747_lo <= 1'b0;
    n750_lo <= 1'b0;
    n756_lo <= 1'b0;
    n759_lo <= 1'b0;
    n762_lo <= 1'b0;
    n768_lo <= 1'b0;
    n771_lo <= 1'b0;
    n774_lo <= 1'b0;
    n780_lo <= 1'b0;
    n783_lo <= 1'b0;
    n786_lo <= 1'b0;
    n792_lo <= 1'b0;
    n795_lo <= 1'b0;
    n804_lo <= 1'b0;
    n807_lo <= 1'b0;
    n816_lo <= 1'b0;
    n819_lo <= 1'b0;
    n828_lo <= 1'b0;
    n831_lo <= 1'b0;
    n843_lo <= 1'b0;
    n846_lo <= 1'b0;
    n849_lo <= 1'b0;
    n852_lo <= 1'b0;
    n855_lo <= 1'b0;
    n858_lo <= 1'b0;
    n861_lo <= 1'b0;
    n864_lo <= 1'b0;
    n867_lo <= 1'b0;
    n870_lo <= 1'b0;
    n879_lo <= 1'b0;
    n891_lo <= 1'b0;
    n903_lo <= 1'b0;
    n915_lo <= 1'b0;
    n918_lo <= 1'b0;
    n927_lo <= 1'b0;
    n951_lo <= 1'b0;
    n954_lo <= 1'b0;
    n957_lo <= 1'b0;
    n960_lo <= 1'b0;
    n963_lo <= 1'b0;
    n966_lo <= 1'b0;
    n972_lo <= 1'b0;
    n975_lo <= 1'b0;
    n978_lo <= 1'b0;
    n984_lo <= 1'b0;
    n987_lo <= 1'b0;
    n990_lo <= 1'b0;
    n996_lo <= 1'b0;
    n999_lo <= 1'b0;
    n1002_lo <= 1'b0;
    n1008_lo <= 1'b0;
    n1011_lo <= 1'b0;
    n1014_lo <= 1'b0;
    n1020_lo <= 1'b0;
    n1023_lo <= 1'b0;
    n1026_lo <= 1'b0;
    n1032_lo <= 1'b0;
    n1035_lo <= 1'b0;
    n1038_lo <= 1'b0;
    n1044_lo <= 1'b0;
    n1047_lo <= 1'b0;
    n1050_lo <= 1'b0;
    n1053_lo <= 1'b0;
    n1056_lo <= 1'b0;
    n1059_lo <= 1'b0;
    n1062_lo <= 1'b0;
    n1065_lo <= 1'b0;
    n1068_lo <= 1'b0;
    n1071_lo <= 1'b0;
    n1074_lo <= 1'b0;
    n1077_lo <= 1'b0;
    n1080_lo <= 1'b0;
    n1083_lo <= 1'b0;
    n1086_lo <= 1'b0;
    n1089_lo <= 1'b0;
    n1092_lo <= 1'b0;
    n1095_lo <= 1'b0;
    n1098_lo <= 1'b0;
    n1101_lo <= 1'b0;
    n1104_lo <= 1'b0;
    n1107_lo <= 1'b0;
    n1110_lo <= 1'b0;
    n1113_lo <= 1'b0;
    n1116_lo <= 1'b0;
    n1119_lo <= 1'b0;
    n1122_lo <= 1'b0;
    n1125_lo <= 1'b0;
    n1128_lo <= 1'b0;
    n1131_lo <= 1'b0;
    n1134_lo <= 1'b0;
    n1137_lo <= 1'b0;
    n1140_lo <= 1'b0;
    n1143_lo <= 1'b0;
    n1146_lo <= 1'b0;
    n1149_lo <= 1'b0;
    n1152_lo <= 1'b0;
    n1155_lo <= 1'b0;
    n1158_lo <= 1'b0;
    n1167_lo <= 1'b0;
    n1170_lo <= 1'b0;
    n1173_lo <= 1'b0;
    n1176_lo <= 1'b0;
    n1179_lo <= 1'b0;
    n1529_o2 <= 1'b0;
    n1616_o2 <= 1'b0;
    n1655_o2 <= 1'b0;
    n1656_o2 <= 1'b0;
    n1657_o2 <= 1'b0;
    n1730_o2 <= 1'b0;
    n1731_o2 <= 1'b0;
    n1732_o2 <= 1'b0;
    n1729_o2 <= 1'b0;
    n1805_o2 <= 1'b0;
    n1808_o2 <= 1'b0;
    n1807_o2 <= 1'b0;
    n1809_o2 <= 1'b0;
    n1663_o2 <= 1'b0;
    n1664_o2 <= 1'b0;
    n1704_o2 <= 1'b0;
    n1705_o2 <= 1'b0;
    n1706_o2 <= 1'b0;
    n1707_o2 <= 1'b0;
    n1708_o2 <= 1'b0;
    n1709_o2 <= 1'b0;
    G280_o2 <= 1'b0;
    G655_o2 <= 1'b0;
    G663_o2 <= 1'b0;
    G672_o2 <= 1'b0;
    G538_o2 <= 1'b0;
    n1780_o2 <= 1'b0;
    n1781_o2 <= 1'b0;
    n1797_o2 <= 1'b0;
    n1798_o2 <= 1'b0;
    n1799_o2 <= 1'b0;
    n1800_o2 <= 1'b0;
    G578_o2 <= 1'b0;
    n1828_o2 <= 1'b0;
    n801_lo_buf_o2 <= 1'b0;
    G693_o2 <= 1'b0;
    G702_o2 <= 1'b0;
    G712_o2 <= 1'b0;
    G685_o2 <= 1'b0;
    G658_o2 <= 1'b0;
    G667_o2 <= 1'b0;
    G677_o2 <= 1'b0;
    G650_o2 <= 1'b0;
    G798_o2 <= 1'b0;
    n1017_lo_buf_o2 <= 1'b0;
    n1029_lo_buf_o2 <= 1'b0;
    n1041_lo_buf_o2 <= 1'b0;
    G558_o2 <= 1'b0;
    G562_o2 <= 1'b0;
    G566_o2 <= 1'b0;
    n1835_o2 <= 1'b0;
    n1836_o2 <= 1'b0;
    n1837_o2 <= 1'b0;
    n765_lo_buf_o2 <= 1'b0;
    n777_lo_buf_o2 <= 1'b0;
    n789_lo_buf_o2 <= 1'b0;
    G617_o2 <= 1'b0;
    G626_o2 <= 1'b0;
    G636_o2 <= 1'b0;
    n489_lo_buf_o2 <= 1'b0;
    n513_lo_buf_o2 <= 1'b0;
    n561_lo_buf_o2 <= 1'b0;
    n597_lo_buf_o2 <= 1'b0;
    n657_lo_buf_o2 <= 1'b0;
    G276_o2 <= 1'b0;
    n1005_lo_buf_o2 <= 1'b0;
    n1161_lo_buf_o2 <= 1'b0;
    G620_o2 <= 1'b0;
    G629_o2 <= 1'b0;
    G639_o2 <= 1'b0;
    G554_o2 <= 1'b0;
    G690_o2 <= 1'b0;
    G698_o2 <= 1'b0;
    G707_o2 <= 1'b0;
    G319_o2 <= 1'b0;
    G389_o2 <= 1'b0;
    n753_lo_buf_o2 <= 1'b0;
    G647_o2 <= 1'b0;
    G769_o2 <= 1'b0;
    G785_o2 <= 1'b0;
    G808_o2 <= 1'b0;
    G445_o2 <= 1'b0;
    G448_o2 <= 1'b0;
    G477_o2 <= 1'b0;
    G480_o2 <= 1'b0;
    G436_o2 <= 1'b0;
    G786_o2 <= 1'b0;
    G787_o2 <= 1'b0;
    G826_o2 <= 1'b0;
    G827_o2 <= 1'b0;
    G825_o2 <= 1'b0;
    G610_o2 <= 1'b0;
    n537_lo_buf_o2 <= 1'b0;
    n669_lo_buf_o2 <= 1'b0;
    n969_lo_buf_o2 <= 1'b0;
    n981_lo_buf_o2 <= 1'b0;
    n993_lo_buf_o2 <= 1'b0;
    G309_o2 <= 1'b0;
    G461_o2 <= 1'b0;
    G487_o2 <= 1'b0;
    G460_o2 <= 1'b0;
    G468_o2 <= 1'b0;
    G287_o2 <= 1'b0;
    G613_o2 <= 1'b0;
    n585_lo_buf_o2 <= 1'b0;
    n813_lo_buf_o2 <= 1'b0;
    n825_lo_buf_o2 <= 1'b0;
    n837_lo_buf_o2 <= 1'b0;
    n897_lo_buf_o2 <= 1'b0;
    n909_lo_buf_o2 <= 1'b0;
    n933_lo_buf_o2 <= 1'b0;
    G451_o2 <= 1'b0;
    G682_o2 <= 1'b0;
    G756_o2 <= 1'b0;
    G542_o2 <= 1'b0;
    G546_o2 <= 1'b0;
    G550_o2 <= 1'b0;
    G310_o2 <= 1'b0;
    n798_lo_buf_o2 <= 1'b0;
    n882_lo_buf_o2 <= 1'b0;
    G427_o2 <= 1'b0;
    G497_o2 <= 1'b0;
    G499_o2 <= 1'b0;
    G501_o2 <= 1'b0;
    G498_o2 <= 1'b0;
    G500_o2 <= 1'b0;
    G502_o2 <= 1'b0;
    G369_o2 <= 1'b0;
    n939_lo_buf_o2 <= 1'b0;
    n486_lo_buf_o2 <= 1'b0;
    n510_lo_buf_o2 <= 1'b0;
    n558_lo_buf_o2 <= 1'b0;
    n594_lo_buf_o2 <= 1'b0;
    n654_lo_buf_o2 <= 1'b0;
    n477_lo_buf_o2 <= 1'b0;
    n525_lo_buf_o2 <= 1'b0;
    n573_lo_buf_o2 <= 1'b0;
  end
endmodule


