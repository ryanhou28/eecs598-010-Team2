// Benchmark "mymod" written by ABC on Sun Oct 29 19:31:53 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33,
    G1884, G1885, G1886, G1887, G1888, G1889, G1890, G1891, G1892, G1893,
    G1894, G1895, G1896, G1897, G1898, G1899, G1900, G1901, G1902, G1903,
    G1904, G1905, G1906, G1907, G1908  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33;
  output G1884, G1885, G1886, G1887, G1888, G1889, G1890, G1891, G1892, G1893,
    G1894, G1895, G1896, G1897, G1898, G1899, G1900, G1901, G1902, G1903,
    G1904, G1905, G1906, G1907, G1908;
  reg n949_lo, n961_lo, n973_lo, n976_lo, n985_lo, n997_lo, n1009_lo,
    n1021_lo, n1024_lo, n1033_lo, n1036_lo, n1045_lo, n1057_lo, n1069_lo,
    n1081_lo, n1093_lo, n1105_lo, n1117_lo, n1129_lo, n1132_lo, n1141_lo,
    n1144_lo, n1156_lo, n1159_lo, n1165_lo, n1168_lo, n1180_lo, n1189_lo,
    n1192_lo, n1201_lo, n1204_lo, n1216_lo, n1228_lo, n1231_lo, n1237_lo,
    n1240_lo, n1243_lo, n1249_lo, n1252_lo, n1255_lo, n1261_lo, n1264_lo,
    n1267_lo, n1273_lo, n1276_lo, n1279_lo, n1282_lo, n1285_lo, n1288_lo,
    n1291_lo, n1294_lo, n1297_lo, n1300_lo, n1303_lo, n1309_lo, n1312_lo,
    n1315_lo, n1318_lo, n1321_lo, n1324_lo, n1333_lo, n1874_o2, n2180_o2,
    n2372_o2, n2190_o2, n2191_o2, n2212_o2, n2213_o2, n2214_o2, n2215_o2,
    n2275_o2, n2276_o2, n2290_o2, n2291_o2, n2681_o2, n2680_o2, n2683_o2,
    n2684_o2, n2686_o2, n2319_o2, n2320_o2, n304_inv, G554_o2, G557_o2,
    G185_o2, G188_o2, G191_o2, G194_o2, G1182_o2, G1222_o2, G1247_o2,
    G1371_o2, G1383_o2, G1386_o2, n2416_o2, n2428_o2, n2438_o2, n2439_o2,
    n2440_o2, n2444_o2, n2497_o2, n2498_o2, n2503_o2, n2505_o2, n2529_o2,
    n2562_o2, n2570_o2, n2571_o2, n2574_o2, n2575_o2, G546_o2, G550_o2,
    n2633_o2, n2639_o2, n2642_o2, n2645_o2, n2679_o2, n2662_o2, n2724_o2,
    G382_o2, G199_o2, G202_o2, G225_o2, G248_o2, G260_o2, n2716_o2,
    n2737_o2, n1174_lo_buf_o2, n1198_lo_buf_o2, G371_o2, G1059_o2,
    n2586_o2, n2587_o2, n460_inv, n2648_o2, n2649_o2, n2650_o2, n2651_o2,
    n2652_o2, G365_o2, G1496_o2, G1502_o2, n2700_o2, n2701_o2, n2733_o2,
    n2734_o2, n2744_o2, n2747_o2, n2754_o2, n2755_o2, n511_inv, G1609_o2,
    G1625_o2, G738_o2, G755_o2, G1511_o2, G1522_o2, G1538_o2, G1549_o2,
    G1563_o2, G1584_o2, G1576_o2, G1598_o2, G1395_o2, G1410_o2, G1420_o2,
    G1434_o2, n562_inv, n1162_lo_buf_o2, n1102_lo_buf_o2, G359_o2,
    n982_lo_buf_o2, n1030_lo_buf_o2, n1042_lo_buf_o2, n583_inv, G606_o2,
    G1118_o2, G1069_o2, G1145_o2, G1209_o2, G1189_o2, G1699_o2, G1702_o2,
    G1705_o2, G1708_o2, G1684_o2, G1687_o2, G1690_o2, G1693_o2, G1696_o2,
    G1642_o2, G1645_o2, G1648_o2, G1651_o2, G1654_o2, G1657_o2, G1660_o2,
    n1222_lo_buf_o2, n1330_lo_buf_o2, n658_inv, n661_inv, n1306_lo_buf_o2,
    n1150_lo_buf_o2, G175_o2, G241_o2, G356_o2, G989_o2, G984_o2, n685_inv,
    n688_inv, n958_lo_buf_o2, n1114_lo_buf_o2, G182_o2, G1215_o2, G971_o2,
    G938_o2, G1198_o2, G1203_o2, G1218_o2, G785_o2, G1168_o2, G1130_o2,
    G1185_o2, G1250_o2, G1225_o2, G1791_o2, G1788_o2, G981_o2, n745_inv,
    n748_inv, G1062_o2, n970_lo_buf_o2, n1006_lo_buf_o2, n1078_lo_buf_o2,
    n1126_lo_buf_o2, n766_inv, G165_o2, n1234_lo_buf_o2, n1246_lo_buf_o2,
    n1258_lo_buf_o2, n1270_lo_buf_o2, G368_o2, G428_o2, G212_o2, G841_o2,
    G788_o2, n1186_lo_buf_o2, G391_o2, G387_o2, G645_o2, G1140_o2,
    G1178_o2, G1370_o2, n820_inv, G1357_o2, G816_o2, G1369_o2, G901_o2,
    G1056_o2, G1107_o2, G1087_o2, G1135_o2, n1018_lo_buf_o2,
    n1090_lo_buf_o2, n853_inv, G131_o2, n859_inv, n862_inv, G338_o2,
    n1171_lo_buf_o2, n1195_lo_buf_o2, G419_o2, G425_o2, G497_o2, G416_o2,
    G491_o2, G500_o2, G353_o2, G641_o2, G1117_o2, G1096_o2, G1143_o2,
    G1112_o2, n1138_lo_buf_o2, n1210_lo_buf_o2, G687_o2, G541_o2, G802_o2,
    G813_o2, G810_o2, G987_o2, G898_o2, n946_lo_buf_o2, n1054_lo_buf_o2,
    G728_o2, G856_o2, n949_1_inv, G942_o2, G1099_o2, G1154_o2, G1131_o2,
    G1169_o2, G134_o2, n970_inv, G470_o2, G344_o2, G362_o2, G482_o2,
    G660_o2, G672_o2, n1096_lo_buf_o2, G479_o2, G669_o2, n994_lo_buf_o2,
    n1066_lo_buf_o2, n1006_inv, G147_o2, G473_o2, G488_o2, G589_o2,
    G663_o2, G684_o2, G605_o2, G774_o2, G782_o2;
  wire new_n709_, new_n711_, new_n713_, new_n715_, new_n717_, new_n719_,
    new_n721_, new_n723_, new_n725_, new_n727_, new_n729_, new_n731_,
    new_n733_, new_n735_, new_n737_, new_n739_, new_n741_, new_n743_,
    new_n745_, new_n747_, new_n749_, new_n751_, new_n753_, new_n755_,
    new_n757_, new_n759_, new_n761_, new_n763_, new_n765_, new_n767_,
    new_n769_, new_n771_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n907_, new_n909_, new_n911_,
    new_n913_, new_n915_, new_n917_, new_n919_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n935_, new_n937_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n965_, new_n966_, new_n967_, new_n969_, new_n971_,
    new_n973_, new_n974_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1025_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1033_,
    new_n1035_, new_n1037_, new_n1039_, new_n1041_, new_n1043_, new_n1045_,
    new_n1047_, new_n1049_, new_n1051_, new_n1052_, new_n1053_, new_n1055_,
    new_n1058_, new_n1059_, new_n1061_, new_n1063_, new_n1065_, new_n1067_,
    new_n1068_, new_n1069_, new_n1071_, new_n1073_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1111_, new_n1112_, new_n1113_,
    new_n1115_, new_n1117_, new_n1119_, new_n1121_, new_n1123_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1168_, new_n1169_, new_n1171_, new_n1173_, new_n1175_, new_n1177_,
    new_n1178_, new_n1179_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1185_, new_n1187_, new_n1189_, new_n1191_, new_n1193_, new_n1195_,
    new_n1197_, new_n1199_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1231_, new_n1233_, new_n1234_, new_n1235_, new_n1237_,
    new_n1239_, new_n1241_, new_n1243_, new_n1245_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1259_, new_n1260_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1301_, new_n1303_, new_n1304_, new_n1305_, new_n1306_,
    new_n1307_, new_n1309_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1361_, new_n1363_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1389_, new_n1390_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_,
    new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_,
    new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_,
    new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_,
    new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_,
    new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_,
    new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_,
    new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_,
    new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_,
    new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_,
    new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_,
    new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_,
    new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_,
    new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_,
    new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_,
    new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_,
    new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_,
    new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_,
    new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_,
    new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_,
    new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_,
    new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_,
    new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_,
    new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_,
    new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_,
    new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_,
    new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_,
    new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_,
    new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_,
    new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_,
    new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_,
    new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_,
    new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_,
    new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_,
    new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_,
    new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_,
    new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_,
    new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_,
    new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_,
    new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_,
    new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_,
    new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_,
    new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_,
    new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_,
    new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_,
    new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_,
    new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_,
    new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_,
    new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_,
    new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_,
    new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_,
    new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_,
    new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_,
    new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_,
    new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_,
    new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_,
    new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_,
    new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_,
    new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_,
    new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_,
    new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_,
    new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_,
    new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_,
    new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_,
    new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_,
    new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_,
    new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_,
    new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_,
    new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_,
    new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_,
    new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_,
    new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_,
    new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_,
    new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_,
    new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_,
    new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_,
    new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_,
    new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_,
    new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_,
    new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_,
    new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_,
    new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_,
    new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_,
    new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_,
    new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_,
    new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_,
    new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_,
    new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_,
    new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_,
    new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_,
    new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_,
    new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_,
    new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_,
    new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_,
    new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_,
    new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_,
    new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_,
    new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_,
    new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_,
    new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_,
    new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_,
    new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_,
    new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_,
    new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_,
    new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_,
    new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_,
    new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_,
    new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_,
    new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_,
    new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_,
    new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_,
    new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_,
    new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_,
    new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_,
    new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_,
    new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_,
    new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_,
    new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_,
    new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_,
    new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_,
    new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_,
    new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_,
    new_n2183_, new_n2184_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_,
    new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_,
    new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_,
    new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_,
    new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_,
    new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_,
    new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_,
    new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_,
    new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_,
    new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_,
    new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_,
    new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_,
    new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_,
    new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_,
    new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_,
    new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_,
    new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_,
    new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_,
    new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_,
    new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_,
    new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_,
    new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_,
    new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_,
    new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_,
    new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_,
    new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_,
    new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_,
    new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_,
    new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_,
    new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_,
    new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_,
    new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_,
    new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_,
    new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_,
    new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_,
    new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_,
    new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_,
    new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_,
    new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_,
    new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_,
    new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_,
    new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_,
    new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_,
    new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_,
    new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_,
    new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_,
    new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_,
    new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_, new_n2982_,
    new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_, new_n2988_,
    new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_,
    new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_, new_n3000_,
    new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_,
    new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_, new_n3012_,
    new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_,
    new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_,
    new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_,
    new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_,
    new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_,
    new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_,
    new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_,
    new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_,
    new_n3061_, new_n3062_, new_n3063_, new_n3064_, n949_li, n961_li,
    n973_li, n976_li, n985_li, n997_li, n1009_li, n1021_li, n1024_li,
    n1033_li, n1036_li, n1045_li, n1057_li, n1069_li, n1081_li, n1093_li,
    n1105_li, n1117_li, n1129_li, n1132_li, n1141_li, n1144_li, n1156_li,
    n1159_li, n1165_li, n1168_li, n1180_li, n1189_li, n1192_li, n1201_li,
    n1204_li, n1216_li, n1228_li, n1231_li, n1237_li, n1240_li, n1243_li,
    n1249_li, n1252_li, n1255_li, n1261_li, n1264_li, n1267_li, n1273_li,
    n1276_li, n1279_li, n1282_li, n1285_li, n1288_li, n1291_li, n1294_li,
    n1297_li, n1300_li, n1303_li, n1309_li, n1312_li, n1315_li, n1318_li,
    n1321_li, n1324_li, n1333_li, n1874_i2, n2180_i2, n2372_i2, n2190_i2,
    n2191_i2, n2212_i2, n2213_i2, n2214_i2, n2215_i2, n2275_i2, n2276_i2,
    n2290_i2, n2291_i2, n2681_i2, n2680_i2, n2683_i2, n2684_i2, n2686_i2,
    n2319_i2, n2320_i2, n2321_i2, G554_i2, G557_i2, G185_i2, G188_i2,
    G191_i2, G194_i2, G1182_i2, G1222_i2, G1247_i2, G1371_i2, G1383_i2,
    G1386_i2, n2416_i2, n2428_i2, n2438_i2, n2439_i2, n2440_i2, n2444_i2,
    n2497_i2, n2498_i2, n2503_i2, n2505_i2, n2529_i2, n2562_i2, n2570_i2,
    n2571_i2, n2574_i2, n2575_i2, G546_i2, G550_i2, n2633_i2, n2639_i2,
    n2642_i2, n2645_i2, n2679_i2, n2662_i2, n2724_i2, G382_i2, G199_i2,
    G202_i2, G225_i2, G248_i2, G260_i2, n2716_i2, n2737_i2,
    n1174_lo_buf_i2, n1198_lo_buf_i2, G371_i2, G1059_i2, n2586_i2,
    n2587_i2, G1019_i2, n2648_i2, n2649_i2, n2650_i2, n2651_i2, n2652_i2,
    G365_i2, G1496_i2, G1502_i2, n2700_i2, n2701_i2, n2733_i2, n2734_i2,
    n2744_i2, n2747_i2, n2754_i2, n2755_i2, n2756_i2, G1609_i2, G1625_i2,
    G738_i2, G755_i2, G1511_i2, G1522_i2, G1538_i2, G1549_i2, G1563_i2,
    G1584_i2, G1576_i2, G1598_i2, G1395_i2, G1410_i2, G1420_i2, G1434_i2,
    G1240_i2, n1162_lo_buf_i2, n1102_lo_buf_i2, G359_i2, n982_lo_buf_i2,
    n1030_lo_buf_i2, n1042_lo_buf_i2, G161_i2, G606_i2, G1118_i2, G1069_i2,
    G1145_i2, G1209_i2, G1189_i2, G1699_i2, G1702_i2, G1705_i2, G1708_i2,
    G1684_i2, G1687_i2, G1690_i2, G1693_i2, G1696_i2, G1642_i2, G1645_i2,
    G1648_i2, G1651_i2, G1654_i2, G1657_i2, G1660_i2, n1222_lo_buf_i2,
    n1330_lo_buf_i2, G123_i2, G142_i2, n1306_lo_buf_i2, n1150_lo_buf_i2,
    G175_i2, G241_i2, G356_i2, G989_i2, G984_i2, G1009_i2, G1012_i2,
    n958_lo_buf_i2, n1114_lo_buf_i2, G182_i2, G1215_i2, G971_i2, G938_i2,
    G1198_i2, G1203_i2, G1218_i2, G785_i2, G1168_i2, G1130_i2, G1185_i2,
    G1250_i2, G1225_i2, G1791_i2, G1788_i2, G981_i2, G1031_i2, G1015_i2,
    G1062_i2, n970_lo_buf_i2, n1006_lo_buf_i2, n1078_lo_buf_i2,
    n1126_lo_buf_i2, G116_i2, G165_i2, n1234_lo_buf_i2, n1246_lo_buf_i2,
    n1258_lo_buf_i2, n1270_lo_buf_i2, G368_i2, G428_i2, G212_i2, G841_i2,
    G788_i2, n1186_lo_buf_i2, G391_i2, G387_i2, G645_i2, G1140_i2,
    G1178_i2, G1370_i2, G1205_i2, G1357_i2, G816_i2, G1369_i2, G901_i2,
    G1056_i2, G1107_i2, G1087_i2, G1135_i2, n1018_lo_buf_i2,
    n1090_lo_buf_i2, G119_i2, G131_i2, G154_i2, G169_i2, G338_i2,
    n1171_lo_buf_i2, n1195_lo_buf_i2, G419_i2, G425_i2, G497_i2, G416_i2,
    G491_i2, G500_i2, G353_i2, G641_i2, G1117_i2, G1096_i2, G1143_i2,
    G1112_i2, n1138_lo_buf_i2, n1210_lo_buf_i2, G687_i2, G541_i2, G802_i2,
    G813_i2, G810_i2, G987_i2, G898_i2, n946_lo_buf_i2, n1054_lo_buf_i2,
    G728_i2, G856_i2, G831_i2, G942_i2, G1099_i2, G1154_i2, G1131_i2,
    G1169_i2, G134_i2, G157_i2, G470_i2, G344_i2, G362_i2, G482_i2,
    G660_i2, G672_i2, n1096_lo_buf_i2, G479_i2, G669_i2, n994_lo_buf_i2,
    n1066_lo_buf_i2, G112_i2, G147_i2, G473_i2, G488_i2, G589_i2, G663_i2,
    G684_i2, G605_i2, G774_i2, G782_i2;
  assign new_n709_ = G1;
  assign new_n711_ = G2;
  assign new_n713_ = G3;
  assign new_n715_ = G4;
  assign new_n717_ = G5;
  assign new_n719_ = G6;
  assign new_n721_ = G7;
  assign new_n723_ = G8;
  assign new_n725_ = G9;
  assign new_n727_ = G10;
  assign new_n729_ = G11;
  assign new_n731_ = G12;
  assign new_n733_ = G13;
  assign new_n735_ = G14;
  assign new_n737_ = G15;
  assign new_n739_ = G16;
  assign new_n741_ = G17;
  assign new_n743_ = G18;
  assign new_n745_ = G19;
  assign new_n747_ = G20;
  assign new_n749_ = G21;
  assign new_n751_ = G22;
  assign new_n753_ = G23;
  assign new_n755_ = G24;
  assign new_n757_ = G25;
  assign new_n759_ = G26;
  assign new_n761_ = G27;
  assign new_n763_ = G28;
  assign new_n765_ = G29;
  assign new_n767_ = G30;
  assign new_n769_ = G31;
  assign new_n771_ = G32;
  assign new_n773_ = G33;
  assign new_n775_ = n949_lo;
  assign new_n776_ = ~n949_lo;
  assign new_n777_ = n961_lo;
  assign new_n778_ = ~n961_lo;
  assign new_n779_ = n973_lo;
  assign new_n780_ = ~n973_lo;
  assign new_n781_ = n976_lo;
  assign new_n782_ = ~n976_lo;
  assign new_n783_ = n985_lo;
  assign new_n784_ = ~n985_lo;
  assign new_n785_ = n997_lo;
  assign new_n786_ = ~n997_lo;
  assign new_n787_ = n1009_lo;
  assign new_n788_ = ~n1009_lo;
  assign new_n789_ = n1021_lo;
  assign new_n790_ = ~n1021_lo;
  assign new_n791_ = n1024_lo;
  assign new_n792_ = ~n1024_lo;
  assign new_n793_ = n1033_lo;
  assign new_n794_ = ~n1033_lo;
  assign new_n795_ = n1036_lo;
  assign new_n796_ = ~n1036_lo;
  assign new_n797_ = n1045_lo;
  assign new_n798_ = ~n1045_lo;
  assign new_n799_ = n1057_lo;
  assign new_n800_ = ~n1057_lo;
  assign new_n801_ = n1069_lo;
  assign new_n802_ = ~n1069_lo;
  assign new_n803_ = n1081_lo;
  assign new_n804_ = ~n1081_lo;
  assign new_n805_ = n1093_lo;
  assign new_n806_ = ~n1093_lo;
  assign new_n807_ = n1105_lo;
  assign new_n808_ = ~n1105_lo;
  assign new_n809_ = n1117_lo;
  assign new_n810_ = ~n1117_lo;
  assign new_n811_ = n1129_lo;
  assign new_n812_ = ~n1129_lo;
  assign new_n813_ = n1132_lo;
  assign new_n815_ = n1141_lo;
  assign new_n816_ = ~n1141_lo;
  assign new_n817_ = n1144_lo;
  assign new_n818_ = ~n1144_lo;
  assign new_n819_ = n1156_lo;
  assign new_n821_ = n1159_lo;
  assign new_n822_ = ~n1159_lo;
  assign new_n823_ = n1165_lo;
  assign new_n824_ = ~n1165_lo;
  assign new_n825_ = n1168_lo;
  assign new_n827_ = n1180_lo;
  assign new_n829_ = n1189_lo;
  assign new_n830_ = ~n1189_lo;
  assign new_n831_ = n1192_lo;
  assign new_n833_ = n1201_lo;
  assign new_n834_ = ~n1201_lo;
  assign new_n835_ = n1204_lo;
  assign new_n837_ = n1216_lo;
  assign new_n838_ = ~n1216_lo;
  assign new_n839_ = n1228_lo;
  assign new_n841_ = n1231_lo;
  assign new_n843_ = n1237_lo;
  assign new_n844_ = ~n1237_lo;
  assign new_n845_ = n1240_lo;
  assign new_n847_ = n1243_lo;
  assign new_n849_ = n1249_lo;
  assign new_n850_ = ~n1249_lo;
  assign new_n851_ = n1252_lo;
  assign new_n853_ = n1255_lo;
  assign new_n855_ = n1261_lo;
  assign new_n856_ = ~n1261_lo;
  assign new_n857_ = n1264_lo;
  assign new_n859_ = n1267_lo;
  assign new_n861_ = n1273_lo;
  assign new_n862_ = ~n1273_lo;
  assign new_n863_ = n1276_lo;
  assign new_n865_ = n1279_lo;
  assign new_n867_ = n1282_lo;
  assign new_n868_ = ~n1282_lo;
  assign new_n869_ = n1285_lo;
  assign new_n870_ = ~n1285_lo;
  assign new_n871_ = n1288_lo;
  assign new_n873_ = n1291_lo;
  assign new_n875_ = n1294_lo;
  assign new_n876_ = ~n1294_lo;
  assign new_n877_ = n1297_lo;
  assign new_n878_ = ~n1297_lo;
  assign new_n879_ = n1300_lo;
  assign new_n881_ = n1303_lo;
  assign new_n883_ = n1309_lo;
  assign new_n884_ = ~n1309_lo;
  assign new_n885_ = n1312_lo;
  assign new_n887_ = n1315_lo;
  assign new_n889_ = n1318_lo;
  assign new_n890_ = ~n1318_lo;
  assign new_n891_ = n1321_lo;
  assign new_n892_ = ~n1321_lo;
  assign new_n893_ = n1324_lo;
  assign new_n894_ = ~n1324_lo;
  assign new_n895_ = n1333_lo;
  assign new_n896_ = ~n1333_lo;
  assign new_n897_ = n1874_o2;
  assign new_n898_ = ~n1874_o2;
  assign new_n899_ = n2180_o2;
  assign new_n900_ = ~n2180_o2;
  assign new_n901_ = n2372_o2;
  assign new_n902_ = ~n2372_o2;
  assign new_n903_ = n2190_o2;
  assign new_n905_ = n2191_o2;
  assign new_n907_ = n2212_o2;
  assign new_n909_ = n2213_o2;
  assign new_n911_ = n2214_o2;
  assign new_n913_ = n2215_o2;
  assign new_n915_ = n2275_o2;
  assign new_n917_ = n2276_o2;
  assign new_n919_ = n2290_o2;
  assign new_n921_ = n2291_o2;
  assign new_n923_ = n2681_o2;
  assign new_n924_ = ~n2681_o2;
  assign new_n925_ = n2680_o2;
  assign new_n926_ = ~n2680_o2;
  assign new_n927_ = n2683_o2;
  assign new_n928_ = ~n2683_o2;
  assign new_n929_ = n2684_o2;
  assign new_n930_ = ~n2684_o2;
  assign new_n931_ = n2686_o2;
  assign new_n932_ = ~n2686_o2;
  assign new_n933_ = n2319_o2;
  assign new_n935_ = n2320_o2;
  assign new_n937_ = n304_inv;
  assign new_n939_ = G554_o2;
  assign new_n940_ = ~G554_o2;
  assign new_n941_ = G557_o2;
  assign new_n942_ = ~G557_o2;
  assign new_n943_ = G185_o2;
  assign new_n944_ = ~G185_o2;
  assign new_n945_ = G188_o2;
  assign new_n946_ = ~G188_o2;
  assign new_n947_ = G191_o2;
  assign new_n948_ = ~G191_o2;
  assign new_n949_ = G194_o2;
  assign new_n950_ = ~G194_o2;
  assign new_n951_ = G1182_o2;
  assign new_n952_ = ~G1182_o2;
  assign new_n953_ = G1222_o2;
  assign new_n954_ = ~G1222_o2;
  assign new_n955_ = G1247_o2;
  assign new_n956_ = ~G1247_o2;
  assign new_n957_ = G1371_o2;
  assign new_n958_ = ~G1371_o2;
  assign new_n959_ = G1383_o2;
  assign new_n960_ = ~G1383_o2;
  assign new_n961_ = G1386_o2;
  assign new_n962_ = ~G1386_o2;
  assign new_n963_ = n2416_o2;
  assign new_n965_ = n2428_o2;
  assign new_n966_ = ~n2428_o2;
  assign new_n967_ = n2438_o2;
  assign new_n969_ = n2439_o2;
  assign new_n971_ = n2440_o2;
  assign new_n973_ = n2444_o2;
  assign new_n974_ = ~n2444_o2;
  assign new_n976_ = ~n2497_o2;
  assign new_n977_ = n2498_o2;
  assign new_n978_ = ~n2498_o2;
  assign new_n979_ = n2503_o2;
  assign new_n980_ = ~n2503_o2;
  assign new_n981_ = n2505_o2;
  assign new_n982_ = ~n2505_o2;
  assign new_n983_ = n2529_o2;
  assign new_n984_ = ~n2529_o2;
  assign new_n985_ = n2562_o2;
  assign new_n986_ = ~n2562_o2;
  assign new_n987_ = n2570_o2;
  assign new_n988_ = ~n2570_o2;
  assign new_n989_ = n2571_o2;
  assign new_n990_ = ~n2571_o2;
  assign new_n991_ = n2574_o2;
  assign new_n992_ = ~n2574_o2;
  assign new_n993_ = n2575_o2;
  assign new_n994_ = ~n2575_o2;
  assign new_n995_ = G546_o2;
  assign new_n996_ = ~G546_o2;
  assign new_n997_ = G550_o2;
  assign new_n998_ = ~G550_o2;
  assign new_n999_ = n2633_o2;
  assign new_n1000_ = ~n2633_o2;
  assign new_n1001_ = n2639_o2;
  assign new_n1002_ = ~n2639_o2;
  assign new_n1003_ = n2642_o2;
  assign new_n1004_ = ~n2642_o2;
  assign new_n1005_ = n2645_o2;
  assign new_n1006_ = ~n2645_o2;
  assign new_n1007_ = n2679_o2;
  assign new_n1009_ = n2662_o2;
  assign new_n1010_ = ~n2662_o2;
  assign new_n1011_ = n2724_o2;
  assign new_n1012_ = ~n2724_o2;
  assign new_n1014_ = ~G382_o2;
  assign new_n1015_ = G199_o2;
  assign new_n1016_ = ~G199_o2;
  assign new_n1017_ = G202_o2;
  assign new_n1018_ = ~G202_o2;
  assign new_n1020_ = ~G225_o2;
  assign new_n1021_ = G248_o2;
  assign new_n1022_ = ~G248_o2;
  assign new_n1023_ = G260_o2;
  assign new_n1024_ = ~G260_o2;
  assign new_n1025_ = n2716_o2;
  assign new_n1028_ = ~n2737_o2;
  assign new_n1029_ = n1174_lo_buf_o2;
  assign new_n1030_ = ~n1174_lo_buf_o2;
  assign new_n1031_ = n1198_lo_buf_o2;
  assign new_n1033_ = G371_o2;
  assign new_n1035_ = G1059_o2;
  assign new_n1037_ = n2586_o2;
  assign new_n1039_ = n2587_o2;
  assign new_n1041_ = n460_inv;
  assign new_n1043_ = n2648_o2;
  assign new_n1045_ = n2649_o2;
  assign new_n1047_ = n2650_o2;
  assign new_n1049_ = n2651_o2;
  assign new_n1051_ = n2652_o2;
  assign new_n1052_ = ~n2652_o2;
  assign new_n1053_ = G365_o2;
  assign new_n1055_ = G1496_o2;
  assign new_n1058_ = ~G1502_o2;
  assign new_n1059_ = n2700_o2;
  assign new_n1061_ = n2701_o2;
  assign new_n1063_ = n2733_o2;
  assign new_n1065_ = n2734_o2;
  assign new_n1067_ = n2744_o2;
  assign new_n1068_ = ~n2744_o2;
  assign new_n1069_ = n2747_o2;
  assign new_n1071_ = n2754_o2;
  assign new_n1073_ = n2755_o2;
  assign new_n1075_ = n511_inv;
  assign new_n1076_ = ~n511_inv;
  assign new_n1077_ = G1609_o2;
  assign new_n1078_ = ~G1609_o2;
  assign new_n1079_ = G1625_o2;
  assign new_n1080_ = ~G1625_o2;
  assign new_n1081_ = G738_o2;
  assign new_n1082_ = ~G738_o2;
  assign new_n1083_ = G755_o2;
  assign new_n1084_ = ~G755_o2;
  assign new_n1085_ = G1511_o2;
  assign new_n1086_ = ~G1511_o2;
  assign new_n1087_ = G1522_o2;
  assign new_n1088_ = ~G1522_o2;
  assign new_n1089_ = G1538_o2;
  assign new_n1090_ = ~G1538_o2;
  assign new_n1091_ = G1549_o2;
  assign new_n1092_ = ~G1549_o2;
  assign new_n1093_ = G1563_o2;
  assign new_n1094_ = ~G1563_o2;
  assign new_n1095_ = G1584_o2;
  assign new_n1096_ = ~G1584_o2;
  assign new_n1097_ = G1576_o2;
  assign new_n1098_ = ~G1576_o2;
  assign new_n1099_ = G1598_o2;
  assign new_n1100_ = ~G1598_o2;
  assign new_n1101_ = G1395_o2;
  assign new_n1102_ = ~G1395_o2;
  assign new_n1103_ = G1410_o2;
  assign new_n1104_ = ~G1410_o2;
  assign new_n1105_ = G1420_o2;
  assign new_n1106_ = ~G1420_o2;
  assign new_n1107_ = G1434_o2;
  assign new_n1108_ = ~G1434_o2;
  assign new_n1109_ = n562_inv;
  assign new_n1111_ = n1162_lo_buf_o2;
  assign new_n1112_ = ~n1162_lo_buf_o2;
  assign new_n1113_ = n1102_lo_buf_o2;
  assign new_n1115_ = G359_o2;
  assign new_n1117_ = n982_lo_buf_o2;
  assign new_n1119_ = n1030_lo_buf_o2;
  assign new_n1121_ = n1042_lo_buf_o2;
  assign new_n1123_ = n583_inv;
  assign new_n1125_ = G606_o2;
  assign new_n1126_ = ~G606_o2;
  assign new_n1127_ = G1118_o2;
  assign new_n1128_ = ~G1118_o2;
  assign new_n1129_ = G1069_o2;
  assign new_n1130_ = ~G1069_o2;
  assign new_n1131_ = G1145_o2;
  assign new_n1132_ = ~G1145_o2;
  assign new_n1133_ = G1209_o2;
  assign new_n1134_ = ~G1209_o2;
  assign new_n1135_ = G1189_o2;
  assign new_n1136_ = ~G1189_o2;
  assign new_n1137_ = G1699_o2;
  assign new_n1138_ = ~G1699_o2;
  assign new_n1139_ = G1702_o2;
  assign new_n1140_ = ~G1702_o2;
  assign new_n1141_ = G1705_o2;
  assign new_n1142_ = ~G1705_o2;
  assign new_n1143_ = G1708_o2;
  assign new_n1144_ = ~G1708_o2;
  assign new_n1145_ = G1684_o2;
  assign new_n1146_ = ~G1684_o2;
  assign new_n1147_ = G1687_o2;
  assign new_n1148_ = ~G1687_o2;
  assign new_n1149_ = G1690_o2;
  assign new_n1150_ = ~G1690_o2;
  assign new_n1151_ = G1693_o2;
  assign new_n1152_ = ~G1693_o2;
  assign new_n1153_ = G1696_o2;
  assign new_n1154_ = ~G1696_o2;
  assign new_n1155_ = G1642_o2;
  assign new_n1156_ = ~G1642_o2;
  assign new_n1157_ = G1645_o2;
  assign new_n1158_ = ~G1645_o2;
  assign new_n1159_ = G1648_o2;
  assign new_n1160_ = ~G1648_o2;
  assign new_n1161_ = G1651_o2;
  assign new_n1162_ = ~G1651_o2;
  assign new_n1163_ = G1654_o2;
  assign new_n1164_ = ~G1654_o2;
  assign new_n1165_ = G1657_o2;
  assign new_n1166_ = ~G1657_o2;
  assign new_n1167_ = G1660_o2;
  assign new_n1168_ = ~G1660_o2;
  assign new_n1169_ = n1222_lo_buf_o2;
  assign new_n1171_ = n1330_lo_buf_o2;
  assign new_n1173_ = n658_inv;
  assign new_n1175_ = n661_inv;
  assign new_n1177_ = n1306_lo_buf_o2;
  assign new_n1178_ = ~n1306_lo_buf_o2;
  assign new_n1179_ = n1150_lo_buf_o2;
  assign new_n1181_ = G175_o2;
  assign new_n1182_ = ~G175_o2;
  assign new_n1183_ = G241_o2;
  assign new_n1184_ = ~G241_o2;
  assign new_n1185_ = G356_o2;
  assign new_n1187_ = G989_o2;
  assign new_n1189_ = G984_o2;
  assign new_n1191_ = n685_inv;
  assign new_n1193_ = n688_inv;
  assign new_n1195_ = n958_lo_buf_o2;
  assign new_n1197_ = n1114_lo_buf_o2;
  assign new_n1199_ = G182_o2;
  assign new_n1201_ = G1215_o2;
  assign new_n1202_ = ~G1215_o2;
  assign new_n1203_ = G971_o2;
  assign new_n1204_ = ~G971_o2;
  assign new_n1205_ = G938_o2;
  assign new_n1206_ = ~G938_o2;
  assign new_n1207_ = G1198_o2;
  assign new_n1208_ = ~G1198_o2;
  assign new_n1209_ = G1203_o2;
  assign new_n1210_ = ~G1203_o2;
  assign new_n1211_ = G1218_o2;
  assign new_n1212_ = ~G1218_o2;
  assign new_n1213_ = G785_o2;
  assign new_n1214_ = ~G785_o2;
  assign new_n1215_ = G1168_o2;
  assign new_n1216_ = ~G1168_o2;
  assign new_n1217_ = G1130_o2;
  assign new_n1218_ = ~G1130_o2;
  assign new_n1219_ = G1185_o2;
  assign new_n1220_ = ~G1185_o2;
  assign new_n1221_ = G1250_o2;
  assign new_n1222_ = ~G1250_o2;
  assign new_n1223_ = G1225_o2;
  assign new_n1224_ = ~G1225_o2;
  assign new_n1225_ = G1791_o2;
  assign new_n1226_ = ~G1791_o2;
  assign new_n1227_ = G1788_o2;
  assign new_n1228_ = ~G1788_o2;
  assign new_n1229_ = G981_o2;
  assign new_n1231_ = n745_inv;
  assign new_n1233_ = n748_inv;
  assign new_n1234_ = ~n748_inv;
  assign new_n1235_ = G1062_o2;
  assign new_n1237_ = n970_lo_buf_o2;
  assign new_n1239_ = n1006_lo_buf_o2;
  assign new_n1241_ = n1078_lo_buf_o2;
  assign new_n1243_ = n1126_lo_buf_o2;
  assign new_n1245_ = n766_inv;
  assign new_n1247_ = G165_o2;
  assign new_n1248_ = ~G165_o2;
  assign new_n1249_ = n1234_lo_buf_o2;
  assign new_n1250_ = ~n1234_lo_buf_o2;
  assign new_n1251_ = n1246_lo_buf_o2;
  assign new_n1252_ = ~n1246_lo_buf_o2;
  assign new_n1253_ = n1258_lo_buf_o2;
  assign new_n1254_ = ~n1258_lo_buf_o2;
  assign new_n1255_ = n1270_lo_buf_o2;
  assign new_n1256_ = ~n1270_lo_buf_o2;
  assign new_n1257_ = G368_o2;
  assign new_n1259_ = G428_o2;
  assign new_n1260_ = ~G428_o2;
  assign new_n1261_ = G212_o2;
  assign new_n1262_ = ~G212_o2;
  assign new_n1263_ = G841_o2;
  assign new_n1264_ = ~G841_o2;
  assign new_n1265_ = G788_o2;
  assign new_n1266_ = ~G788_o2;
  assign new_n1267_ = n1186_lo_buf_o2;
  assign new_n1269_ = G391_o2;
  assign new_n1270_ = ~G391_o2;
  assign new_n1271_ = G387_o2;
  assign new_n1272_ = ~G387_o2;
  assign new_n1273_ = G645_o2;
  assign new_n1274_ = ~G645_o2;
  assign new_n1275_ = G1140_o2;
  assign new_n1276_ = ~G1140_o2;
  assign new_n1277_ = G1178_o2;
  assign new_n1278_ = ~G1178_o2;
  assign new_n1279_ = G1370_o2;
  assign new_n1280_ = ~G1370_o2;
  assign new_n1281_ = n820_inv;
  assign new_n1282_ = ~n820_inv;
  assign new_n1283_ = G1357_o2;
  assign new_n1284_ = ~G1357_o2;
  assign new_n1285_ = G816_o2;
  assign new_n1286_ = ~G816_o2;
  assign new_n1287_ = G1369_o2;
  assign new_n1288_ = ~G1369_o2;
  assign new_n1289_ = G901_o2;
  assign new_n1290_ = ~G901_o2;
  assign new_n1291_ = G1056_o2;
  assign new_n1292_ = ~G1056_o2;
  assign new_n1293_ = G1107_o2;
  assign new_n1294_ = ~G1107_o2;
  assign new_n1295_ = G1087_o2;
  assign new_n1296_ = ~G1087_o2;
  assign new_n1297_ = G1135_o2;
  assign new_n1298_ = ~G1135_o2;
  assign new_n1299_ = n1018_lo_buf_o2;
  assign new_n1301_ = n1090_lo_buf_o2;
  assign new_n1303_ = n853_inv;
  assign new_n1304_ = ~n853_inv;
  assign new_n1305_ = G131_o2;
  assign new_n1306_ = ~G131_o2;
  assign new_n1307_ = n859_inv;
  assign new_n1309_ = n862_inv;
  assign new_n1311_ = G338_o2;
  assign new_n1312_ = ~G338_o2;
  assign new_n1313_ = n1171_lo_buf_o2;
  assign new_n1314_ = ~n1171_lo_buf_o2;
  assign new_n1315_ = n1195_lo_buf_o2;
  assign new_n1316_ = ~n1195_lo_buf_o2;
  assign new_n1317_ = G419_o2;
  assign new_n1318_ = ~G419_o2;
  assign new_n1319_ = G425_o2;
  assign new_n1320_ = ~G425_o2;
  assign new_n1321_ = G497_o2;
  assign new_n1322_ = ~G497_o2;
  assign new_n1323_ = G416_o2;
  assign new_n1324_ = ~G416_o2;
  assign new_n1325_ = G491_o2;
  assign new_n1326_ = ~G491_o2;
  assign new_n1327_ = G500_o2;
  assign new_n1328_ = ~G500_o2;
  assign new_n1329_ = G353_o2;
  assign new_n1330_ = ~G353_o2;
  assign new_n1331_ = G641_o2;
  assign new_n1332_ = ~G641_o2;
  assign new_n1333_ = G1117_o2;
  assign new_n1334_ = ~G1117_o2;
  assign new_n1335_ = G1096_o2;
  assign new_n1336_ = ~G1096_o2;
  assign new_n1337_ = G1143_o2;
  assign new_n1338_ = ~G1143_o2;
  assign new_n1339_ = G1112_o2;
  assign new_n1340_ = ~G1112_o2;
  assign new_n1341_ = n1138_lo_buf_o2;
  assign new_n1342_ = ~n1138_lo_buf_o2;
  assign new_n1343_ = n1210_lo_buf_o2;
  assign new_n1344_ = ~n1210_lo_buf_o2;
  assign new_n1345_ = G687_o2;
  assign new_n1346_ = ~G687_o2;
  assign new_n1347_ = G541_o2;
  assign new_n1348_ = ~G541_o2;
  assign new_n1349_ = G802_o2;
  assign new_n1350_ = ~G802_o2;
  assign new_n1351_ = G813_o2;
  assign new_n1352_ = ~G813_o2;
  assign new_n1353_ = G810_o2;
  assign new_n1354_ = ~G810_o2;
  assign new_n1355_ = G987_o2;
  assign new_n1356_ = ~G987_o2;
  assign new_n1357_ = G898_o2;
  assign new_n1358_ = ~G898_o2;
  assign new_n1359_ = n946_lo_buf_o2;
  assign new_n1361_ = n1054_lo_buf_o2;
  assign new_n1363_ = G728_o2;
  assign new_n1364_ = ~G728_o2;
  assign new_n1365_ = G856_o2;
  assign new_n1366_ = ~G856_o2;
  assign new_n1367_ = n949_1_inv;
  assign new_n1368_ = ~n949_1_inv;
  assign new_n1369_ = G942_o2;
  assign new_n1370_ = ~G942_o2;
  assign new_n1371_ = G1099_o2;
  assign new_n1372_ = ~G1099_o2;
  assign new_n1373_ = G1154_o2;
  assign new_n1374_ = ~G1154_o2;
  assign new_n1375_ = G1131_o2;
  assign new_n1376_ = ~G1131_o2;
  assign new_n1377_ = G1169_o2;
  assign new_n1378_ = ~G1169_o2;
  assign new_n1379_ = G134_o2;
  assign new_n1380_ = ~G134_o2;
  assign new_n1381_ = n970_inv;
  assign new_n1383_ = G470_o2;
  assign new_n1384_ = ~G470_o2;
  assign new_n1385_ = G344_o2;
  assign new_n1386_ = ~G344_o2;
  assign new_n1387_ = G362_o2;
  assign new_n1389_ = G482_o2;
  assign new_n1390_ = ~G482_o2;
  assign new_n1391_ = G660_o2;
  assign new_n1392_ = ~G660_o2;
  assign new_n1393_ = G672_o2;
  assign new_n1394_ = ~G672_o2;
  assign new_n1395_ = n1096_lo_buf_o2;
  assign new_n1396_ = ~n1096_lo_buf_o2;
  assign new_n1397_ = G479_o2;
  assign new_n1398_ = ~G479_o2;
  assign new_n1399_ = G669_o2;
  assign new_n1400_ = ~G669_o2;
  assign new_n1401_ = n994_lo_buf_o2;
  assign new_n1402_ = ~n994_lo_buf_o2;
  assign new_n1403_ = n1066_lo_buf_o2;
  assign new_n1404_ = ~n1066_lo_buf_o2;
  assign new_n1405_ = n1006_inv;
  assign new_n1406_ = ~n1006_inv;
  assign new_n1407_ = G147_o2;
  assign new_n1408_ = ~G147_o2;
  assign new_n1409_ = G473_o2;
  assign new_n1410_ = ~G473_o2;
  assign new_n1411_ = G488_o2;
  assign new_n1412_ = ~G488_o2;
  assign new_n1413_ = G589_o2;
  assign new_n1414_ = ~G589_o2;
  assign new_n1415_ = G663_o2;
  assign new_n1416_ = ~G663_o2;
  assign new_n1417_ = G684_o2;
  assign new_n1418_ = ~G684_o2;
  assign new_n1419_ = G605_o2;
  assign new_n1420_ = ~G605_o2;
  assign new_n1421_ = G774_o2;
  assign new_n1422_ = ~G774_o2;
  assign new_n1423_ = G782_o2;
  assign new_n1424_ = ~G782_o2;
  assign new_n1425_ = new_n2535_ & new_n2536_;
  assign new_n1426_ = new_n2537_ | new_n2538_;
  assign new_n1427_ = new_n2540_ & new_n2543_;
  assign new_n1428_ = new_n2547_ | new_n2550_;
  assign new_n1429_ = new_n1427_ & new_n2555_;
  assign new_n1430_ = new_n1428_ | new_n2562_;
  assign new_n1431_ = new_n1429_ & new_n2566_;
  assign new_n1432_ = new_n1430_ | new_n2573_;
  assign new_n1433_ = new_n1431_ & new_n775_;
  assign new_n1434_ = new_n1432_ & new_n776_;
  assign new_n1435_ = new_n1434_ | new_n1433_;
  assign new_n1436_ = new_n2540_ & new_n2580_;
  assign new_n1437_ = new_n2547_ | new_n2583_;
  assign new_n1438_ = new_n2584_ & new_n2587_;
  assign new_n1439_ = new_n2591_ | new_n2594_;
  assign new_n1440_ = new_n1438_ & new_n2566_;
  assign new_n1441_ = new_n1439_ | new_n2573_;
  assign new_n1442_ = new_n1440_ & new_n777_;
  assign new_n1443_ = new_n1441_ & new_n778_;
  assign new_n1444_ = new_n1443_ | new_n1442_;
  assign new_n1445_ = new_n2584_ & new_n2599_;
  assign new_n1446_ = new_n2591_ | new_n2602_;
  assign new_n1447_ = new_n1445_ & new_n2567_;
  assign new_n1448_ = new_n1446_ | new_n2574_;
  assign new_n1449_ = new_n1447_ & new_n779_;
  assign new_n1450_ = new_n1448_ & new_n780_;
  assign new_n1451_ = new_n1450_ | new_n1449_;
  assign new_n1452_ = new_n2539_ & new_n2605_;
  assign new_n1453_ = new_n2546_ | new_n2608_;
  assign new_n1454_ = new_n1452_ & new_n2555_;
  assign new_n1455_ = new_n1453_ | new_n2562_;
  assign new_n1456_ = new_n1454_ & new_n2567_;
  assign new_n1457_ = new_n1455_ | new_n2574_;
  assign new_n1458_ = new_n1456_ & new_n783_;
  assign new_n1459_ = new_n1457_ & new_n784_;
  assign new_n1460_ = new_n1459_ | new_n1458_;
  assign new_n1461_ = new_n2535_ & new_n2610_;
  assign new_n1462_ = new_n2537_ | new_n2612_;
  assign new_n1463_ = new_n1461_ & new_n2614_;
  assign new_n1464_ = new_n1462_ | new_n2617_;
  assign new_n1465_ = new_n1463_ & new_n2599_;
  assign new_n1466_ = new_n1464_ | new_n2602_;
  assign new_n1467_ = new_n1465_ & new_n2621_;
  assign new_n1468_ = new_n1466_ | new_n2628_;
  assign new_n1469_ = new_n1467_ & new_n799_;
  assign new_n1470_ = new_n1468_ & new_n800_;
  assign new_n1471_ = new_n1470_ | new_n1469_;
  assign new_n1472_ = new_n2633_ & new_n2610_;
  assign new_n1473_ = new_n2634_ | new_n2612_;
  assign new_n1474_ = new_n2635_ & new_n2543_;
  assign new_n1475_ = new_n2636_ | new_n2550_;
  assign new_n1476_ = new_n1474_ & new_n2637_;
  assign new_n1477_ = new_n1475_ | new_n2638_;
  assign new_n1478_ = new_n1476_ & new_n2621_;
  assign new_n1479_ = new_n1477_ | new_n2628_;
  assign new_n1480_ = new_n1478_ & new_n809_;
  assign new_n1481_ = new_n1479_ & new_n810_;
  assign new_n1482_ = new_n1481_ | new_n1480_;
  assign new_n1483_ = new_n2635_ & new_n2614_;
  assign new_n1484_ = new_n2636_ | new_n2617_;
  assign new_n1485_ = new_n1483_ & new_n2587_;
  assign new_n1486_ = new_n1484_ | new_n2594_;
  assign new_n1487_ = new_n1485_ & new_n2622_;
  assign new_n1488_ = new_n1486_ | new_n2629_;
  assign new_n1489_ = new_n1487_ & new_n811_;
  assign new_n1490_ = new_n1488_ & new_n812_;
  assign new_n1491_ = new_n1490_ | new_n1489_;
  assign new_n1492_ = new_n2536_ & new_n2640_;
  assign new_n1493_ = new_n2538_ | new_n2642_;
  assign new_n1494_ = new_n1492_ & new_n2544_;
  assign new_n1495_ = new_n1493_ | new_n2549_;
  assign new_n1496_ = new_n1494_ & new_n2588_;
  assign new_n1497_ = new_n1495_ | new_n2595_;
  assign new_n1498_ = new_n1496_ & new_n2569_;
  assign new_n1499_ = new_n1497_ | new_n2576_;
  assign new_n1500_ = new_n1498_ & new_n785_;
  assign new_n1501_ = new_n1499_ & new_n786_;
  assign new_n1502_ = new_n1501_ | new_n1500_;
  assign new_n1503_ = new_n2609_ & new_n2640_;
  assign new_n1504_ = new_n2611_ | new_n2642_;
  assign new_n1505_ = new_n2644_ & new_n2544_;
  assign new_n1506_ = new_n2647_ | new_n2551_;
  assign new_n1507_ = new_n1505_ & new_n2598_;
  assign new_n1508_ = new_n1506_ | new_n2603_;
  assign new_n1509_ = new_n1507_ & new_n2569_;
  assign new_n1510_ = new_n1508_ | new_n2576_;
  assign new_n1511_ = new_n1509_ & new_n787_;
  assign new_n1512_ = new_n1510_ & new_n788_;
  assign new_n1513_ = new_n1512_ | new_n1511_;
  assign new_n1514_ = new_n2644_ & new_n2615_;
  assign new_n1515_ = new_n2647_ | new_n2618_;
  assign new_n1516_ = new_n1514_ & new_n2556_;
  assign new_n1517_ = new_n1515_ | new_n2563_;
  assign new_n1518_ = new_n1516_ & new_n2570_;
  assign new_n1519_ = new_n1517_ | new_n2577_;
  assign new_n1520_ = new_n1518_ & new_n789_;
  assign new_n1521_ = new_n1519_ & new_n790_;
  assign new_n1522_ = new_n1521_ | new_n1520_;
  assign new_n1523_ = new_n2645_ & new_n2580_;
  assign new_n1524_ = new_n2648_ | new_n2583_;
  assign new_n1525_ = new_n2649_ & new_n2637_;
  assign new_n1526_ = new_n1524_ | new_n2638_;
  assign new_n1527_ = new_n1525_ & new_n2570_;
  assign new_n1528_ = new_n1526_ | new_n2577_;
  assign new_n1529_ = new_n1527_ & new_n793_;
  assign new_n1530_ = new_n1528_ & new_n794_;
  assign new_n1531_ = new_n1530_ | new_n1529_;
  assign new_n1532_ = new_n2645_ & new_n2605_;
  assign new_n1533_ = new_n2648_ | new_n2608_;
  assign new_n1534_ = new_n1532_ & new_n2588_;
  assign new_n1535_ = new_n1533_ | new_n2595_;
  assign new_n1536_ = new_n1534_ & new_n2622_;
  assign new_n1537_ = new_n1535_ | new_n2629_;
  assign new_n1538_ = new_n1536_ & new_n797_;
  assign new_n1539_ = new_n1537_ & new_n798_;
  assign new_n1540_ = new_n1539_ | new_n1538_;
  assign new_n1541_ = new_n2633_ & new_n2651_;
  assign new_n1542_ = new_n2634_ | new_n1078_;
  assign new_n1543_ = new_n2653_ & new_n2545_;
  assign new_n1544_ = new_n2656_ | new_n2551_;
  assign new_n1545_ = new_n2657_ & new_n2590_;
  assign new_n1546_ = new_n2658_ | new_n2596_;
  assign new_n1547_ = new_n1545_ & new_n2624_;
  assign new_n1548_ = new_n1546_ | new_n2631_;
  assign new_n1549_ = new_n1547_ & new_n801_;
  assign new_n1550_ = new_n1548_ & new_n802_;
  assign new_n1551_ = new_n1550_ | new_n1549_;
  assign new_n1552_ = new_n2657_ & new_n2600_;
  assign new_n1553_ = new_n2658_ | new_n2603_;
  assign new_n1554_ = new_n1552_ & new_n2624_;
  assign new_n1555_ = new_n1553_ | new_n2631_;
  assign new_n1556_ = new_n1554_ & new_n803_;
  assign new_n1557_ = new_n1555_ & new_n804_;
  assign new_n1558_ = new_n1557_ | new_n1556_;
  assign new_n1559_ = new_n2653_ & new_n2615_;
  assign new_n1560_ = new_n2656_ | new_n2618_;
  assign new_n1561_ = new_n1559_ & new_n2556_;
  assign new_n1562_ = new_n1560_ | new_n2563_;
  assign new_n1563_ = new_n1561_ & new_n2625_;
  assign new_n1564_ = new_n1562_ | new_n2632_;
  assign new_n1565_ = new_n1563_ & new_n805_;
  assign new_n1566_ = new_n1564_ & new_n806_;
  assign new_n1567_ = new_n1566_ | new_n1565_;
  assign new_n1568_ = new_n2654_ & new_n2606_;
  assign new_n1569_ = new_n2655_ | new_n2607_;
  assign new_n1570_ = new_n1568_ & new_n2590_;
  assign new_n1571_ = new_n1569_ | new_n2596_;
  assign new_n1572_ = new_n1570_ & new_n2625_;
  assign new_n1573_ = new_n1571_ | new_n2632_;
  assign new_n1574_ = new_n1572_ & new_n807_;
  assign new_n1575_ = new_n1573_ & new_n808_;
  assign new_n1576_ = new_n1575_ | new_n1574_;
  assign new_n1577_ = new_n955_ | new_n941_;
  assign new_n1578_ = new_n956_ | new_n942_;
  assign new_n1579_ = new_n1578_ & new_n1577_;
  assign new_n1580_ = new_n952_ | new_n949_;
  assign new_n1581_ = new_n951_ | new_n950_;
  assign new_n1582_ = new_n1581_ & new_n1580_;
  assign new_n1583_ = new_n954_ | new_n947_;
  assign new_n1584_ = new_n953_ | new_n948_;
  assign new_n1585_ = new_n1584_ & new_n1583_;
  assign new_n1586_ = new_n957_ | new_n945_;
  assign new_n1587_ = new_n958_ | new_n946_;
  assign new_n1588_ = new_n1587_ & new_n1586_;
  assign new_n1589_ = new_n962_ | new_n943_;
  assign new_n1590_ = new_n961_ | new_n944_;
  assign new_n1591_ = new_n1590_ & new_n1589_;
  assign new_n1592_ = new_n959_ | new_n939_;
  assign new_n1593_ = new_n960_ | new_n940_;
  assign new_n1594_ = new_n1593_ & new_n1592_;
  assign new_n1595_ = new_n1582_ & new_n1579_;
  assign new_n1596_ = new_n1595_ & new_n1585_;
  assign new_n1597_ = new_n1596_ & new_n1588_;
  assign new_n1598_ = new_n1597_ & new_n996_;
  assign new_n1599_ = new_n1598_ & new_n1591_;
  assign new_n1600_ = new_n1599_ & new_n1594_;
  assign new_n1601_ = new_n1600_ & new_n998_;
  assign new_n1602_ = new_n1601_ | new_n1023_;
  assign new_n1603_ = new_n2659_ | new_n2661_;
  assign new_n1604_ = new_n1603_ | new_n2661_;
  assign new_n1605_ = new_n1024_ & new_n1020_;
  assign new_n1606_ = new_n1605_ & new_n1014_;
  assign new_n1607_ = new_n2649_ & new_n2557_;
  assign new_n1608_ = new_n1607_ & new_n2664_;
  assign new_n1609_ = new_n2654_ & new_n2581_;
  assign new_n1610_ = new_n1609_ & new_n2557_;
  assign new_n1611_ = new_n1610_ & new_n2664_;
  assign new_n1612_ = new_n2641_ & new_n2651_;
  assign new_n1613_ = new_n2670_ & new_n2545_;
  assign new_n1614_ = new_n1613_ & new_n2559_;
  assign new_n1615_ = new_n1614_ & new_n2665_;
  assign new_n1616_ = new_n2670_ & new_n2581_;
  assign new_n1617_ = new_n2671_ & new_n2589_;
  assign new_n1618_ = new_n1617_ & new_n2665_;
  assign new_n1619_ = new_n2671_ & new_n2600_;
  assign new_n1620_ = new_n1619_ & new_n2667_;
  assign new_n1621_ = new_n2669_ & new_n2606_;
  assign new_n1622_ = new_n1621_ & new_n2559_;
  assign new_n1623_ = new_n1622_ & new_n2667_;
  assign new_n1624_ = new_n1058_ & new_n997_;
  assign new_n1625_ = new_n1624_ & new_n2650_;
  assign new_n1626_ = new_n1625_ & new_n2582_;
  assign new_n1627_ = new_n1626_ & new_n2560_;
  assign new_n1628_ = new_n1627_ & new_n2668_;
  assign new_n1629_ = new_n1055_ & new_n995_;
  assign new_n1630_ = new_n1629_ & new_n2641_;
  assign new_n1631_ = new_n1630_ & new_n2582_;
  assign new_n1632_ = new_n1631_ & new_n2560_;
  assign new_n1633_ = new_n1632_ & new_n2668_;
  assign new_n1634_ = new_n1611_ | new_n1608_;
  assign new_n1635_ = new_n1634_ | new_n1615_;
  assign new_n1636_ = new_n1635_ | new_n1618_;
  assign new_n1637_ = new_n1636_ | new_n1620_;
  assign new_n1638_ = new_n1637_ | new_n1623_;
  assign new_n1639_ = new_n1638_ | new_n1628_;
  assign new_n1640_ = new_n1639_ | new_n1633_;
  assign new_n1641_ = new_n1228_ & new_n1226_;
  assign new_n1642_ = new_n1227_ | new_n1225_;
  assign new_n1643_ = new_n2674_ | new_n1640_;
  assign new_n1644_ = new_n2659_ | new_n892_;
  assign new_n1645_ = new_n1644_ | new_n1643_;
  assign new_n1646_ = new_n1645_ & new_n1604_;
  assign new_n1647_ = new_n1213_ & new_n1131_;
  assign new_n1648_ = new_n1214_ | new_n1132_;
  assign new_n1649_ = new_n1220_ & new_n1126_;
  assign new_n1650_ = new_n1219_ | new_n1125_;
  assign new_n1651_ = new_n1650_ & new_n1648_;
  assign new_n1652_ = new_n1649_ | new_n1647_;
  assign new_n1653_ = new_n2678_ & new_n2679_;
  assign new_n1654_ = new_n2680_ | new_n2681_;
  assign new_n1655_ = new_n2680_ & new_n2681_;
  assign new_n1656_ = new_n2678_ | new_n2679_;
  assign new_n1657_ = new_n1656_ & new_n1654_;
  assign new_n1658_ = new_n1655_ | new_n1653_;
  assign new_n1659_ = new_n925_ & new_n815_;
  assign new_n1660_ = new_n926_ | new_n816_;
  assign new_n1661_ = new_n1659_ & new_n2684_;
  assign new_n1662_ = new_n1660_ | new_n2689_;
  assign new_n1663_ = new_n1661_ & new_n2674_;
  assign new_n1664_ = new_n1662_ | new_n2694_;
  assign new_n1665_ = new_n1664_ & new_n1658_;
  assign new_n1666_ = new_n1663_ & new_n1657_;
  assign new_n1667_ = new_n1666_ | new_n1665_;
  assign new_n1668_ = new_n2699_ | new_n2660_;
  assign new_n1669_ = new_n2703_ & new_n1667_;
  assign new_n1670_ = new_n1206_ & new_n1204_;
  assign new_n1671_ = new_n1205_ | new_n1203_;
  assign new_n1672_ = new_n1215_ & new_n1133_;
  assign new_n1673_ = new_n1216_ | new_n1134_;
  assign new_n1674_ = new_n1222_ & new_n1128_;
  assign new_n1675_ = new_n1221_ | new_n1127_;
  assign new_n1676_ = new_n1675_ & new_n1673_;
  assign new_n1677_ = new_n1674_ | new_n1672_;
  assign new_n1678_ = new_n2706_ & new_n2707_;
  assign new_n1679_ = new_n2708_ | new_n2709_;
  assign new_n1680_ = new_n2708_ & new_n2709_;
  assign new_n1681_ = new_n2706_ | new_n2707_;
  assign new_n1682_ = new_n1681_ & new_n1679_;
  assign new_n1683_ = new_n1680_ | new_n1678_;
  assign new_n1684_ = new_n2684_ & new_n843_;
  assign new_n1685_ = new_n2689_ | new_n844_;
  assign new_n1686_ = new_n1684_ & new_n2675_;
  assign new_n1687_ = new_n1685_ | new_n2694_;
  assign new_n1688_ = new_n1687_ & new_n1683_;
  assign new_n1689_ = new_n1686_ & new_n1682_;
  assign new_n1690_ = new_n1689_ | new_n1688_;
  assign new_n1691_ = new_n1690_ & new_n2703_;
  assign new_n1692_ = new_n2685_ & new_n855_;
  assign new_n1693_ = new_n2690_ | new_n856_;
  assign new_n1694_ = new_n1692_ & new_n2675_;
  assign new_n1695_ = new_n1693_ | new_n2695_;
  assign new_n1696_ = new_n1695_ & new_n930_;
  assign new_n1697_ = new_n1694_ & new_n929_;
  assign new_n1698_ = new_n1697_ | new_n1696_;
  assign new_n1699_ = new_n1698_ & new_n2704_;
  assign new_n1700_ = new_n2685_ & new_n861_;
  assign new_n1701_ = new_n2690_ | new_n862_;
  assign new_n1702_ = new_n1700_ & new_n2677_;
  assign new_n1703_ = new_n1701_ | new_n2695_;
  assign new_n1704_ = new_n1703_ & new_n928_;
  assign new_n1705_ = new_n1702_ & new_n927_;
  assign new_n1706_ = new_n1705_ | new_n1704_;
  assign new_n1707_ = new_n1706_ & new_n2704_;
  assign new_n1708_ = new_n923_ & new_n823_;
  assign new_n1709_ = new_n924_ | new_n824_;
  assign new_n1710_ = new_n1708_ & new_n2686_;
  assign new_n1711_ = new_n1709_ | new_n2691_;
  assign new_n1712_ = new_n1710_ & new_n2677_;
  assign new_n1713_ = new_n1711_ | new_n2696_;
  assign new_n1714_ = new_n1713_ & new_n931_;
  assign new_n1715_ = new_n1712_ & new_n932_;
  assign new_n1716_ = new_n1715_ | new_n1714_;
  assign new_n1717_ = new_n1716_ & new_n2705_;
  assign new_n1718_ = new_n1158_ & new_n1156_;
  assign new_n1719_ = new_n1157_ | new_n1155_;
  assign new_n1720_ = new_n1718_ & new_n1160_;
  assign new_n1721_ = new_n1719_ | new_n1159_;
  assign new_n1722_ = new_n1720_ & new_n1162_;
  assign new_n1723_ = new_n1721_ | new_n1161_;
  assign new_n1724_ = new_n1722_ & new_n1146_;
  assign new_n1725_ = new_n1723_ | new_n1145_;
  assign new_n1726_ = new_n1724_ & new_n1148_;
  assign new_n1727_ = new_n1725_ | new_n1147_;
  assign new_n1728_ = new_n1726_ & new_n1150_;
  assign new_n1729_ = new_n1727_ | new_n1149_;
  assign new_n1730_ = new_n1728_ & new_n1152_;
  assign new_n1731_ = new_n1729_ | new_n1151_;
  assign new_n1732_ = new_n1731_ & new_n2711_;
  assign new_n1733_ = new_n1730_ | new_n2699_;
  assign new_n1734_ = new_n1207_ & new_n1202_;
  assign new_n1735_ = new_n1208_ | new_n1201_;
  assign new_n1736_ = new_n2713_ & new_n1016_;
  assign new_n1737_ = new_n2714_ | new_n1015_;
  assign new_n1738_ = new_n1737_ & new_n1734_;
  assign new_n1739_ = new_n1736_ | new_n1735_;
  assign new_n1740_ = new_n2715_ & new_n2716_;
  assign new_n1741_ = new_n2717_ | new_n2718_;
  assign new_n1742_ = new_n2717_ & new_n2718_;
  assign new_n1743_ = new_n2715_ | new_n2716_;
  assign new_n1744_ = new_n1743_ & new_n1741_;
  assign new_n1745_ = new_n1742_ | new_n1740_;
  assign new_n1746_ = new_n869_ & new_n829_;
  assign new_n1747_ = new_n870_ | new_n830_;
  assign new_n1748_ = new_n1747_ & new_n2711_;
  assign new_n1749_ = new_n1746_ | new_n2698_;
  assign new_n1750_ = new_n1749_ & new_n1745_;
  assign new_n1751_ = new_n1748_ & new_n1744_;
  assign new_n1752_ = new_n1751_ | new_n1750_;
  assign new_n1753_ = new_n1164_ & new_n1154_;
  assign new_n1754_ = new_n1163_ | new_n1153_;
  assign new_n1755_ = new_n1753_ & new_n1138_;
  assign new_n1756_ = new_n1754_ | new_n1137_;
  assign new_n1757_ = new_n1755_ & new_n1140_;
  assign new_n1758_ = new_n1756_ | new_n1139_;
  assign new_n1759_ = new_n1757_ & new_n1142_;
  assign new_n1760_ = new_n1758_ | new_n1141_;
  assign new_n1761_ = new_n1759_ & new_n1144_;
  assign new_n1762_ = new_n1760_ | new_n1143_;
  assign new_n1763_ = new_n1761_ & new_n1166_;
  assign new_n1764_ = new_n1762_ | new_n1165_;
  assign new_n1765_ = new_n1763_ & new_n1168_;
  assign new_n1766_ = new_n1764_ | new_n1167_;
  assign new_n1767_ = new_n1766_ & new_n2712_;
  assign new_n1768_ = new_n1765_ | new_n2700_;
  assign new_n1769_ = new_n2713_ & new_n1018_;
  assign new_n1770_ = new_n2714_ | new_n1017_;
  assign new_n1771_ = new_n1211_ & new_n1210_;
  assign new_n1772_ = new_n1212_ | new_n1209_;
  assign new_n1773_ = new_n1771_ & new_n1770_;
  assign new_n1774_ = new_n1772_ | new_n1769_;
  assign new_n1775_ = new_n2719_ & new_n2720_;
  assign new_n1776_ = new_n2721_ | new_n2722_;
  assign new_n1777_ = new_n2721_ & new_n2722_;
  assign new_n1778_ = new_n2719_ | new_n2720_;
  assign new_n1779_ = new_n1778_ & new_n1776_;
  assign new_n1780_ = new_n1777_ | new_n1775_;
  assign new_n1781_ = new_n877_ & new_n833_;
  assign new_n1782_ = new_n878_ | new_n834_;
  assign new_n1783_ = new_n1782_ & new_n2712_;
  assign new_n1784_ = new_n1781_ | new_n2700_;
  assign new_n1785_ = new_n1784_ & new_n1780_;
  assign new_n1786_ = new_n1783_ & new_n1779_;
  assign new_n1787_ = new_n1786_ | new_n1785_;
  assign new_n1788_ = new_n1218_ & new_n1135_;
  assign new_n1789_ = new_n1217_ | new_n1136_;
  assign new_n1790_ = new_n1224_ & new_n1129_;
  assign new_n1791_ = new_n1223_ | new_n1130_;
  assign new_n1792_ = new_n1791_ & new_n1789_;
  assign new_n1793_ = new_n1790_ | new_n1788_;
  assign new_n1794_ = new_n2686_ & new_n849_;
  assign new_n1795_ = new_n2691_ | new_n850_;
  assign new_n1796_ = new_n1794_ & new_n2676_;
  assign new_n1797_ = new_n1795_ | new_n2696_;
  assign new_n1798_ = new_n2723_ & new_n2724_;
  assign new_n1799_ = new_n2725_ | new_n2726_;
  assign new_n1800_ = new_n2725_ & new_n2726_;
  assign new_n1801_ = new_n2723_ | new_n2724_;
  assign new_n1802_ = new_n1801_ & new_n1799_;
  assign new_n1803_ = new_n1800_ | new_n1798_;
  assign new_n1804_ = new_n2727_ & new_n2728_;
  assign new_n1805_ = new_n2729_ | new_n2730_;
  assign new_n1806_ = new_n2729_ & new_n2730_;
  assign new_n1807_ = new_n2727_ | new_n2728_;
  assign new_n1808_ = new_n1807_ & new_n1805_;
  assign new_n1809_ = new_n1806_ | new_n1804_;
  assign new_n1810_ = new_n1808_ & new_n1803_;
  assign new_n1811_ = new_n1809_ & new_n1802_;
  assign new_n1812_ = new_n1811_ | new_n1810_;
  assign new_n1813_ = new_n1812_ & new_n2705_;
  assign new_n1814_ = new_n2732_ & new_n2733_;
  assign new_n1815_ = new_n2734_ | new_n1012_;
  assign new_n1816_ = new_n2736_ & new_n2737_;
  assign new_n1817_ = new_n2738_ | new_n1112_;
  assign new_n1818_ = new_n2739_ & new_n2742_;
  assign new_n1819_ = new_n1276_ | new_n2747_;
  assign new_n1820_ = new_n2750_ & new_n2742_;
  assign new_n1821_ = new_n1278_ | new_n2747_;
  assign new_n1822_ = new_n1282_ & new_n2743_;
  assign new_n1823_ = new_n2751_ | new_n2748_;
  assign new_n1824_ = new_n1284_ & new_n2743_;
  assign new_n1825_ = new_n1283_ | new_n2748_;
  assign new_n1826_ = new_n1288_ & new_n2744_;
  assign new_n1827_ = new_n1287_ | new_n2749_;
  assign new_n1828_ = new_n1279_ & new_n2744_;
  assign new_n1829_ = new_n1280_ | new_n2749_;
  assign new_n1830_ = new_n2732_ & new_n983_;
  assign new_n1831_ = new_n2734_ | new_n984_;
  assign new_n1832_ = new_n2736_ & new_n1029_;
  assign new_n1833_ = new_n2738_ | new_n1030_;
  assign new_n1834_ = new_n1199_ | new_n976_;
  assign new_n1835_ = new_n2752_ & new_n1182_;
  assign new_n1836_ = new_n1342_ | new_n1181_;
  assign new_n1837_ = new_n1835_ & new_n2754_;
  assign new_n1838_ = new_n1836_ | new_n2757_;
  assign new_n1839_ = new_n2759_ & new_n2754_;
  assign new_n1840_ = new_n1316_ | new_n2757_;
  assign new_n1841_ = new_n2760_ | new_n2761_;
  assign new_n1842_ = new_n1826_ | new_n1815_;
  assign new_n1843_ = new_n1842_ & new_n1841_;
  assign new_n1844_ = new_n1829_ | new_n2763_;
  assign new_n1845_ = new_n2764_ | new_n1250_;
  assign new_n1846_ = new_n1845_ & new_n1844_;
  assign new_n1847_ = new_n2766_ & new_n2767_;
  assign new_n1848_ = new_n2769_ & new_n2770_;
  assign new_n1849_ = new_n2771_ & new_n868_;
  assign new_n1850_ = new_n1849_ & new_n2773_;
  assign new_n1851_ = new_n1850_ & new_n2775_;
  assign new_n1852_ = new_n2773_ & new_n890_;
  assign new_n1853_ = new_n1852_ & new_n2775_;
  assign new_n1854_ = new_n2777_ | new_n1851_;
  assign new_n1855_ = new_n2771_ & new_n876_;
  assign new_n1856_ = new_n1855_ & new_n2772_;
  assign new_n1857_ = new_n1856_ & new_n2776_;
  assign new_n1858_ = new_n1857_ | new_n2777_;
  assign new_n1859_ = new_n2766_ | new_n1831_;
  assign new_n1860_ = new_n2769_ | new_n1833_;
  assign new_n1861_ = new_n2778_ | new_n2779_;
  assign new_n1862_ = new_n1822_ | new_n1817_;
  assign new_n1863_ = new_n1862_ & new_n1861_;
  assign new_n1864_ = new_n2780_ | new_n2782_;
  assign new_n1865_ = new_n1824_ | new_n1252_;
  assign new_n1866_ = new_n1865_ & new_n1864_;
  assign new_n1867_ = new_n1866_ & new_n1863_;
  assign new_n1868_ = new_n1819_ | new_n2784_;
  assign new_n1869_ = new_n2785_ | new_n1256_;
  assign new_n1870_ = new_n1869_ & new_n1868_;
  assign new_n1871_ = new_n1821_ | new_n2787_;
  assign new_n1872_ = new_n2788_ | new_n1254_;
  assign new_n1873_ = new_n1872_ & new_n1871_;
  assign new_n1874_ = new_n1873_ & new_n1870_;
  assign new_n1875_ = new_n1340_ & new_n1337_;
  assign new_n1876_ = new_n1339_ | new_n1338_;
  assign new_n1877_ = new_n2789_ & new_n2790_;
  assign new_n1878_ = new_n2791_ | new_n2793_;
  assign new_n1879_ = new_n2791_ & new_n2793_;
  assign new_n1880_ = new_n2789_ | new_n2790_;
  assign new_n1881_ = new_n1880_ & new_n1878_;
  assign new_n1882_ = new_n1879_ | new_n1877_;
  assign new_n1883_ = new_n988_ & new_n985_;
  assign new_n1884_ = new_n987_ & new_n986_;
  assign new_n1885_ = new_n1884_ | new_n1883_;
  assign new_n1886_ = new_n1005_ & new_n1000_;
  assign new_n1887_ = new_n1006_ & new_n999_;
  assign new_n1888_ = new_n1887_ | new_n1886_;
  assign new_n1889_ = new_n1003_ & new_n1002_;
  assign new_n1890_ = new_n1004_ & new_n1001_;
  assign new_n1891_ = new_n1890_ | new_n1889_;
  assign new_n1892_ = new_n2795_ & new_n2797_;
  assign new_n1893_ = new_n1892_ & new_n2800_;
  assign new_n1894_ = new_n1893_ & new_n2806_;
  assign new_n1895_ = new_n1894_ & new_n2811_;
  assign new_n1896_ = new_n2814_ & new_n2816_;
  assign new_n1897_ = new_n1896_ & new_n2800_;
  assign new_n1898_ = new_n1897_ & new_n2806_;
  assign new_n1899_ = new_n2817_ & new_n2819_;
  assign new_n1900_ = new_n2817_ & new_n2811_;
  assign new_n1901_ = new_n2795_ & new_n2814_;
  assign new_n1902_ = new_n1901_ & new_n2801_;
  assign new_n1903_ = new_n1902_ & new_n2807_;
  assign new_n1904_ = new_n2820_ & new_n2819_;
  assign new_n1905_ = new_n2820_ & new_n2812_;
  assign new_n1906_ = new_n2821_ & new_n2822_;
  assign new_n1907_ = new_n2823_ | new_n2824_;
  assign new_n1908_ = new_n2823_ & new_n2824_;
  assign new_n1909_ = new_n2821_ | new_n2822_;
  assign new_n1910_ = new_n1909_ & new_n1907_;
  assign new_n1911_ = new_n1908_ | new_n1906_;
  assign new_n1912_ = new_n1911_ & new_n2826_;
  assign new_n1913_ = new_n1910_ & new_n2829_;
  assign new_n1914_ = new_n1913_ | new_n1912_;
  assign new_n1915_ = new_n2831_ & new_n2832_;
  assign new_n1916_ = new_n2833_ | new_n2834_;
  assign new_n1917_ = new_n2833_ & new_n2834_;
  assign new_n1918_ = new_n2831_ | new_n2832_;
  assign new_n1919_ = new_n1918_ & new_n1916_;
  assign new_n1920_ = new_n1917_ | new_n1915_;
  assign new_n1921_ = new_n1920_ & new_n2836_;
  assign new_n1922_ = new_n1919_ & new_n2838_;
  assign new_n1923_ = new_n1922_ | new_n1921_;
  assign new_n1924_ = new_n1421_ & new_n1383_;
  assign new_n1925_ = new_n1422_ | new_n1384_;
  assign new_n1926_ = new_n1414_ & new_n1392_;
  assign new_n1927_ = new_n1413_ | new_n1391_;
  assign new_n1928_ = new_n1927_ & new_n1925_;
  assign new_n1929_ = new_n1926_ | new_n1924_;
  assign new_n1930_ = new_n1929_ & new_n2840_;
  assign new_n1931_ = new_n1928_ & new_n2841_;
  assign new_n1932_ = new_n1931_ | new_n1930_;
  assign new_n1933_ = new_n1423_ & new_n1389_;
  assign new_n1934_ = new_n1424_ | new_n1390_;
  assign new_n1935_ = new_n1420_ & new_n1394_;
  assign new_n1936_ = new_n1419_ | new_n1393_;
  assign new_n1937_ = new_n1936_ & new_n1934_;
  assign new_n1938_ = new_n1935_ | new_n1933_;
  assign new_n1939_ = new_n1938_ & new_n2826_;
  assign new_n1940_ = new_n1937_ & new_n2829_;
  assign new_n1941_ = new_n1940_ | new_n1939_;
  assign new_n1942_ = new_n991_ & new_n989_;
  assign new_n1943_ = new_n992_ & new_n990_;
  assign new_n1944_ = new_n1943_ | new_n1942_;
  assign new_n1945_ = new_n2842_ | new_n2843_;
  assign new_n1946_ = new_n1009_ & new_n979_;
  assign new_n1947_ = new_n1010_ & new_n980_;
  assign new_n1948_ = new_n1947_ | new_n1946_;
  assign new_n1949_ = new_n2844_ | new_n2845_;
  assign new_n1950_ = new_n2844_ & new_n2845_;
  assign new_n1951_ = new_n2842_ & new_n2843_;
  assign new_n1952_ = new_n1265_ & new_n1264_;
  assign new_n1953_ = new_n1266_ | new_n1263_;
  assign new_n1954_ = new_n2846_ & new_n2847_;
  assign new_n1955_ = new_n2848_ | new_n2849_;
  assign new_n1956_ = new_n2848_ & new_n2849_;
  assign new_n1957_ = new_n2846_ | new_n2847_;
  assign new_n1958_ = new_n1957_ & new_n1955_;
  assign new_n1959_ = new_n1956_ | new_n1954_;
  assign new_n1960_ = new_n1958_ & new_n993_;
  assign new_n1961_ = new_n1959_ & new_n994_;
  assign new_n1962_ = new_n1961_ | new_n1960_;
  assign new_n1963_ = new_n982_ & new_n973_;
  assign new_n1964_ = new_n981_ & new_n974_;
  assign new_n1965_ = new_n1964_ | new_n1963_;
  assign new_n1966_ = new_n2850_ & new_n2851_;
  assign new_n1967_ = new_n2850_ | new_n2851_;
  assign new_n1968_ = new_n2854_ | new_n2857_;
  assign new_n1969_ = new_n1968_ | new_n2860_;
  assign new_n1970_ = new_n1969_ | new_n2860_;
  assign new_n1971_ = new_n1970_ | new_n2861_;
  assign new_n1972_ = new_n1971_ | new_n2861_;
  assign new_n1973_ = new_n1972_ | new_n2854_;
  assign new_n1974_ = new_n1973_ | new_n2855_;
  assign new_n1975_ = new_n2867_ | new_n2871_;
  assign new_n1976_ = new_n1975_ | new_n2871_;
  assign new_n1977_ = new_n1976_ | new_n2872_;
  assign new_n1978_ = new_n1977_ | new_n2872_;
  assign new_n1979_ = new_n2876_ & new_n2878_;
  assign new_n1980_ = new_n2879_ | new_n2880_;
  assign new_n1981_ = new_n2879_ & new_n2880_;
  assign new_n1982_ = new_n2876_ | new_n2878_;
  assign new_n1983_ = new_n1982_ & new_n1980_;
  assign new_n1984_ = new_n1981_ | new_n1979_;
  assign new_n1985_ = new_n1984_ & new_n2840_;
  assign new_n1986_ = new_n1983_ & new_n2841_;
  assign new_n1987_ = new_n1986_ | new_n1985_;
  assign new_n1988_ = new_n2881_ & new_n2882_;
  assign new_n1989_ = new_n2883_ | new_n2884_;
  assign new_n1990_ = new_n2883_ & new_n2884_;
  assign new_n1991_ = new_n2881_ | new_n2882_;
  assign new_n1992_ = new_n1991_ & new_n1989_;
  assign new_n1993_ = new_n1990_ | new_n1988_;
  assign new_n1994_ = new_n1993_ & new_n2886_;
  assign new_n1995_ = new_n1992_ & new_n1404_;
  assign new_n1996_ = new_n1995_ | new_n1994_;
  assign new_n1997_ = new_n2888_ & new_n2890_;
  assign new_n1998_ = new_n2888_ | new_n2890_;
  assign new_n1999_ = new_n2892_ | new_n2894_;
  assign new_n2000_ = new_n2897_ | new_n2894_;
  assign new_n2001_ = new_n2899_ & new_n2900_;
  assign new_n2002_ = new_n2901_ | new_n2902_;
  assign new_n2003_ = new_n2901_ & new_n2902_;
  assign new_n2004_ = new_n2899_ | new_n2900_;
  assign new_n2005_ = new_n2004_ & new_n2002_;
  assign new_n2006_ = new_n2003_ | new_n2001_;
  assign new_n2007_ = new_n2903_ & new_n2904_;
  assign new_n2008_ = new_n2905_ | new_n2906_;
  assign new_n2009_ = new_n2905_ & new_n2906_;
  assign new_n2010_ = new_n2903_ | new_n2904_;
  assign new_n2011_ = new_n2010_ & new_n2008_;
  assign new_n2012_ = new_n2009_ | new_n2007_;
  assign new_n2013_ = new_n2907_ & new_n2908_;
  assign new_n2014_ = new_n2909_ | new_n2910_;
  assign new_n2015_ = new_n2909_ & new_n2910_;
  assign new_n2016_ = new_n2907_ | new_n2908_;
  assign new_n2017_ = new_n2016_ & new_n2014_;
  assign new_n2018_ = new_n2015_ | new_n2013_;
  assign new_n2019_ = new_n2911_ & new_n2912_;
  assign new_n2020_ = new_n2897_ | new_n822_;
  assign new_n2021_ = new_n2019_ & new_n2755_;
  assign new_n2022_ = new_n2020_ | new_n2758_;
  assign new_n2023_ = new_n2022_ & new_n2018_;
  assign new_n2024_ = new_n2021_ & new_n2017_;
  assign new_n2025_ = new_n2024_ | new_n2023_;
  assign new_n2026_ = new_n2913_ & new_n2914_;
  assign new_n2027_ = new_n2915_ | new_n2916_;
  assign new_n2028_ = new_n2915_ & new_n2916_;
  assign new_n2029_ = new_n2913_ | new_n2914_;
  assign new_n2030_ = new_n2029_ & new_n2027_;
  assign new_n2031_ = new_n2028_ | new_n2026_;
  assign new_n2032_ = new_n2917_ & new_n2918_;
  assign new_n2033_ = new_n2919_ | new_n2920_;
  assign new_n2034_ = new_n2919_ & new_n2920_;
  assign new_n2035_ = new_n2917_ | new_n2918_;
  assign new_n2036_ = new_n2035_ & new_n2033_;
  assign new_n2037_ = new_n2034_ | new_n2032_;
  assign new_n2038_ = new_n2921_ & new_n2922_;
  assign new_n2039_ = new_n2923_ | new_n2924_;
  assign new_n2040_ = new_n2923_ & new_n2924_;
  assign new_n2041_ = new_n2921_ | new_n2922_;
  assign new_n2042_ = new_n2041_ & new_n2039_;
  assign new_n2043_ = new_n2040_ | new_n2038_;
  assign new_n2044_ = new_n2925_ & new_n2926_;
  assign new_n2045_ = new_n2927_ | new_n2928_;
  assign new_n2046_ = new_n2927_ & new_n2928_;
  assign new_n2047_ = new_n2925_ | new_n2926_;
  assign new_n2048_ = new_n2047_ & new_n2045_;
  assign new_n2049_ = new_n2046_ | new_n2044_;
  assign new_n2050_ = new_n2929_ & new_n2930_;
  assign new_n2051_ = new_n2931_ | new_n2932_;
  assign new_n2052_ = new_n2931_ & new_n2932_;
  assign new_n2053_ = new_n2929_ | new_n2930_;
  assign new_n2054_ = new_n2053_ & new_n2051_;
  assign new_n2055_ = new_n2052_ | new_n2050_;
  assign new_n2056_ = new_n2054_ & new_n2043_;
  assign new_n2057_ = new_n2055_ & new_n2042_;
  assign new_n2058_ = new_n2057_ | new_n2056_;
  assign new_n2059_ = new_n2933_ & new_n2934_;
  assign new_n2060_ = new_n2935_ | new_n2936_;
  assign new_n2061_ = new_n2935_ & new_n2936_;
  assign new_n2062_ = new_n2933_ | new_n2934_;
  assign new_n2063_ = new_n2062_ & new_n2060_;
  assign new_n2064_ = new_n2061_ | new_n2059_;
  assign new_n2065_ = new_n2937_ & new_n2939_;
  assign new_n2066_ = new_n2940_ | new_n2941_;
  assign new_n2067_ = new_n2940_ & new_n2941_;
  assign new_n2068_ = new_n2937_ | new_n2939_;
  assign new_n2069_ = new_n2068_ & new_n2066_;
  assign new_n2070_ = new_n2067_ | new_n2065_;
  assign new_n2071_ = new_n1377_ & new_n1292_;
  assign new_n2072_ = new_n1378_ | new_n1291_;
  assign new_n2073_ = new_n1371_ & new_n1298_;
  assign new_n2074_ = new_n1372_ | new_n1297_;
  assign new_n2075_ = new_n2074_ & new_n2072_;
  assign new_n2076_ = new_n2073_ | new_n2071_;
  assign new_n2077_ = new_n2942_ & new_n2944_;
  assign new_n2078_ = new_n2946_ | new_n2947_;
  assign new_n2079_ = new_n2946_ & new_n2947_;
  assign new_n2080_ = new_n2942_ | new_n2944_;
  assign new_n2081_ = new_n2080_ & new_n2078_;
  assign new_n2082_ = new_n2079_ | new_n2077_;
  assign new_n2083_ = new_n2082_ & new_n2070_;
  assign new_n2084_ = new_n2081_ & new_n2069_;
  assign new_n2085_ = new_n2084_ | new_n2083_;
  assign new_n2086_ = new_n1363_ & new_n1290_;
  assign new_n2087_ = new_n1364_ | new_n1289_;
  assign new_n2088_ = new_n1369_ & new_n1274_;
  assign new_n2089_ = new_n1370_ | new_n1273_;
  assign new_n2090_ = new_n2089_ & new_n2087_;
  assign new_n2091_ = new_n2088_ | new_n2086_;
  assign new_n2092_ = new_n1348_ & new_n1285_;
  assign new_n2093_ = new_n1347_ | new_n1286_;
  assign new_n2094_ = new_n1366_ & new_n1259_;
  assign new_n2095_ = new_n1365_ | new_n1260_;
  assign new_n2096_ = new_n2095_ & new_n2093_;
  assign new_n2097_ = new_n2094_ | new_n2092_;
  assign new_n2098_ = new_n2948_ & new_n2949_;
  assign new_n2099_ = new_n2950_ | new_n2951_;
  assign new_n2100_ = new_n2950_ & new_n2951_;
  assign new_n2101_ = new_n2948_ | new_n2949_;
  assign new_n2102_ = new_n2101_ & new_n2099_;
  assign new_n2103_ = new_n2100_ | new_n2098_;
  assign new_n2104_ = new_n2911_ & new_n2952_;
  assign new_n2105_ = new_n2898_ | new_n1314_;
  assign new_n2106_ = new_n2104_ & new_n2755_;
  assign new_n2107_ = new_n2105_ | new_n2758_;
  assign new_n2108_ = new_n2953_ & new_n2954_;
  assign new_n2109_ = new_n2955_ | new_n2891_;
  assign new_n2110_ = new_n2955_ & new_n2891_;
  assign new_n2111_ = new_n2953_ | new_n2954_;
  assign new_n2112_ = new_n2111_ & new_n2109_;
  assign new_n2113_ = new_n2110_ | new_n2108_;
  assign new_n2114_ = new_n2112_ | new_n2102_;
  assign new_n2115_ = new_n2113_ | new_n2103_;
  assign new_n2116_ = new_n2115_ & new_n2114_;
  assign new_n2117_ = new_n2957_ & new_n2959_;
  assign new_n2118_ = new_n2960_ | new_n2961_;
  assign new_n2119_ = new_n2960_ & new_n2961_;
  assign new_n2120_ = new_n2957_ | new_n2959_;
  assign new_n2121_ = new_n2120_ & new_n2118_;
  assign new_n2122_ = new_n2119_ | new_n2117_;
  assign new_n2123_ = new_n1374_ & new_n1295_;
  assign new_n2124_ = new_n1373_ | new_n1296_;
  assign new_n2125_ = new_n1376_ & new_n1293_;
  assign new_n2126_ = new_n1375_ | new_n1294_;
  assign new_n2127_ = new_n2126_ & new_n2124_;
  assign new_n2128_ = new_n2125_ | new_n2123_;
  assign new_n2129_ = new_n2962_ & new_n2963_;
  assign new_n2130_ = new_n2964_ | new_n2966_;
  assign new_n2131_ = new_n2964_ & new_n2966_;
  assign new_n2132_ = new_n2962_ | new_n2963_;
  assign new_n2133_ = new_n2132_ & new_n2130_;
  assign new_n2134_ = new_n2131_ | new_n2129_;
  assign new_n2135_ = new_n2133_ | new_n2122_;
  assign new_n2136_ = new_n2134_ | new_n2121_;
  assign new_n2137_ = new_n2136_ & new_n2135_;
  assign new_n2138_ = new_n2827_ & new_n2968_;
  assign new_n2139_ = new_n2830_ & new_n2970_;
  assign new_n2140_ = new_n2139_ | new_n2138_;
  assign new_n2141_ = new_n1336_ & new_n1334_;
  assign new_n2142_ = new_n1335_ | new_n1333_;
  assign new_n2143_ = new_n2971_ & new_n2973_;
  assign new_n2144_ = new_n2974_ | new_n2975_;
  assign new_n2145_ = new_n2974_ & new_n2975_;
  assign new_n2146_ = new_n2971_ | new_n2973_;
  assign new_n2147_ = new_n2146_ & new_n2144_;
  assign new_n2148_ = new_n2145_ | new_n2143_;
  assign new_n2149_ = new_n2147_ & new_n1882_;
  assign new_n2150_ = new_n2148_ & new_n2976_;
  assign new_n2151_ = new_n2150_ | new_n2149_;
  assign new_n2152_ = new_n1396_ | new_n2978_;
  assign new_n2153_ = new_n2981_ | new_n2984_;
  assign new_n2154_ = new_n2153_ & new_n2152_;
  assign new_n2155_ = new_n2986_ & new_n2987_;
  assign new_n2156_ = new_n2990_ & new_n2978_;
  assign new_n2157_ = new_n2990_ | new_n2977_;
  assign new_n2158_ = new_n2994_ | new_n2996_;
  assign new_n2159_ = new_n2994_ & new_n2996_;
  assign new_n2160_ = new_n838_ & new_n2997_;
  assign new_n2161_ = new_n2999_ | new_n818_;
  assign new_n2162_ = new_n2160_ & new_n2986_;
  assign new_n2163_ = new_n2161_ | new_n3001_;
  assign new_n2164_ = new_n2163_ & new_n3002_;
  assign new_n2165_ = new_n2162_ & new_n3003_;
  assign new_n2166_ = new_n2165_ | new_n2164_;
  assign new_n2167_ = new_n2830_ & new_n3002_;
  assign new_n2168_ = new_n2827_ & new_n3003_;
  assign new_n2169_ = new_n2168_ | new_n2167_;
  assign new_n2170_ = new_n1306_ & new_n3005_;
  assign new_n2171_ = new_n1305_ & new_n3007_;
  assign new_n2172_ = new_n2171_ | new_n2170_;
  assign new_n2173_ = new_n3008_ & new_n2970_;
  assign new_n2174_ = new_n3009_ | new_n2968_;
  assign new_n2175_ = new_n3009_ & new_n2967_;
  assign new_n2176_ = new_n3008_ | new_n2969_;
  assign new_n2177_ = new_n2176_ & new_n2174_;
  assign new_n2178_ = new_n2175_ | new_n2173_;
  assign new_n2179_ = new_n2178_ & new_n2836_;
  assign new_n2180_ = new_n2177_ & new_n2838_;
  assign new_n2181_ = new_n2180_ | new_n2179_;
  assign new_n2182_ = new_n3005_ & new_n782_;
  assign new_n2183_ = new_n3007_ & new_n3012_;
  assign new_n2184_ = new_n2183_ | new_n2182_;
  assign G1884 = new_n1435_;
  assign G1885 = new_n1444_;
  assign G1886 = new_n1451_;
  assign G1887 = new_n1460_;
  assign G1888 = new_n1471_;
  assign G1889 = new_n1482_;
  assign G1890 = new_n1491_;
  assign G1891 = new_n1502_;
  assign G1892 = new_n1513_;
  assign G1893 = new_n1522_;
  assign G1894 = new_n1531_;
  assign G1895 = new_n1540_;
  assign G1896 = new_n1551_;
  assign G1897 = new_n1558_;
  assign G1898 = new_n1567_;
  assign G1899 = new_n1576_;
  assign G1900 = new_n1646_;
  assign G1901 = new_n1669_;
  assign G1902 = new_n1691_;
  assign G1903 = new_n1699_;
  assign G1904 = new_n1707_;
  assign G1905 = new_n1717_;
  assign G1906 = new_n1752_;
  assign G1907 = new_n1787_;
  assign G1908 = new_n1813_;
  assign n949_li = new_n919_;
  assign n961_li = new_n903_;
  assign n973_li = new_n907_;
  assign n976_li = new_n715_;
  assign n985_li = new_n967_;
  assign n997_li = new_n933_;
  assign n1009_li = new_n909_;
  assign n1021_li = new_n915_;
  assign n1024_li = new_n723_;
  assign n1033_li = new_n969_;
  assign n1036_li = new_n725_;
  assign n1045_li = new_n971_;
  assign n1057_li = new_n921_;
  assign n1069_li = new_n935_;
  assign n1081_li = new_n911_;
  assign n1093_li = new_n917_;
  assign n1105_li = new_n963_;
  assign n1117_li = new_n905_;
  assign n1129_li = new_n913_;
  assign n1132_li = new_n741_;
  assign n1141_li = new_n2733_;
  assign n1144_li = new_n743_;
  assign n1156_li = new_n745_;
  assign n1159_li = new_n819_;
  assign n1165_li = new_n2737_;
  assign n1168_li = new_n747_;
  assign n1180_li = new_n749_;
  assign n1189_li = new_n1007_;
  assign n1192_li = new_n751_;
  assign n1201_li = new_n1031_;
  assign n1204_li = new_n753_;
  assign n1216_li = new_n755_;
  assign n1228_li = new_n757_;
  assign n1231_li = new_n839_;
  assign n1237_li = new_n2763_;
  assign n1240_li = new_n759_;
  assign n1243_li = new_n845_;
  assign n1249_li = new_n2782_;
  assign n1252_li = new_n761_;
  assign n1255_li = new_n851_;
  assign n1261_li = new_n2787_;
  assign n1264_li = new_n763_;
  assign n1267_li = new_n857_;
  assign n1273_li = new_n2784_;
  assign n1276_li = new_n765_;
  assign n1279_li = new_n863_;
  assign n1282_li = new_n865_;
  assign n1285_li = new_n3015_;
  assign n1288_li = new_n767_;
  assign n1291_li = new_n871_;
  assign n1294_li = new_n873_;
  assign n1297_li = new_n3016_;
  assign n1300_li = new_n769_;
  assign n1303_li = new_n879_;
  assign n1309_li = new_n1177_;
  assign n1312_li = new_n771_;
  assign n1315_li = new_n885_;
  assign n1318_li = new_n887_;
  assign n1321_li = new_n3017_;
  assign n1324_li = new_n773_;
  assign n1333_li = new_n3019_;
  assign n1874_i2 = new_n937_;
  assign n2180_i2 = new_n1033_;
  assign n2372_i2 = new_n1109_;
  assign n2190_i2 = new_n1037_;
  assign n2191_i2 = new_n1039_;
  assign n2212_i2 = new_n1043_;
  assign n2213_i2 = new_n1045_;
  assign n2214_i2 = new_n1047_;
  assign n2215_i2 = new_n1049_;
  assign n2275_i2 = new_n1059_;
  assign n2276_i2 = new_n1061_;
  assign n2290_i2 = new_n1063_;
  assign n2291_i2 = new_n1065_;
  assign n2681_i2 = new_n2735_;
  assign n2680_i2 = new_n2731_;
  assign n2683_i2 = new_n2739_;
  assign n2684_i2 = new_n2750_;
  assign n2686_i2 = new_n2751_;
  assign n2319_i2 = new_n1071_;
  assign n2320_i2 = new_n1073_;
  assign n2321_i2 = new_n2958_;
  assign G554_i2 = new_n2761_;
  assign G557_i2 = new_n2779_;
  assign G185_i2 = new_n2762_;
  assign G188_i2 = new_n2781_;
  assign G191_i2 = new_n2786_;
  assign G194_i2 = new_n2783_;
  assign G1182_i2 = new_n2785_;
  assign G1222_i2 = new_n2788_;
  assign G1247_i2 = new_n2778_;
  assign G1371_i2 = new_n2780_;
  assign G1383_i2 = new_n2760_;
  assign G1386_i2 = new_n2764_;
  assign n2416_i2 = new_n1113_;
  assign n2428_i2 = new_n1115_;
  assign n2438_i2 = new_n1117_;
  assign n2439_i2 = new_n1119_;
  assign n2440_i2 = new_n1121_;
  assign n2444_i2 = new_n1123_;
  assign n2497_i2 = new_n2892_;
  assign n2498_i2 = new_n1171_;
  assign n2503_i2 = new_n1173_;
  assign n2505_i2 = new_n1175_;
  assign n2529_i2 = new_n1179_;
  assign n2562_i2 = new_n1185_;
  assign n2570_i2 = new_n1187_;
  assign n2571_i2 = new_n1189_;
  assign n2574_i2 = new_n1191_;
  assign n2575_i2 = new_n1193_;
  assign G546_i2 = new_n2767_;
  assign G550_i2 = new_n2770_;
  assign n2633_i2 = new_n1229_;
  assign n2639_i2 = new_n1231_;
  assign n2642_i2 = new_n2945_;
  assign n2645_i2 = new_n1235_;
  assign n2679_i2 = new_n1267_;
  assign n2662_i2 = new_n1257_;
  assign n2724_i2 = new_n2752_;
  assign G382_i2 = ~new_n2776_;
  assign G199_i2 = n1285_li;
  assign G202_i2 = n1297_li;
  assign G225_i2 = n1321_li;
  assign G248_i2 = n1333_li;
  assign G260_i2 = new_n3018_;
  assign n2716_i2 = new_n2972_;
  assign n2737_i2 = new_n2792_;
  assign n1174_lo_buf_i2 = new_n2952_;
  assign n1198_lo_buf_i2 = new_n2759_;
  assign G371_i2 = new_n2956_;
  assign G1059_i2 = n2642_i2;
  assign n2586_i2 = new_n1195_;
  assign n2587_i2 = new_n1197_;
  assign G1019_i2 = new_n2965_;
  assign n2648_i2 = new_n1237_;
  assign n2649_i2 = new_n1239_;
  assign n2650_i2 = new_n1241_;
  assign n2651_i2 = new_n1243_;
  assign n2652_i2 = new_n1245_;
  assign G365_i2 = new_n2938_;
  assign G1496_i2 = new_n2765_;
  assign G1502_i2 = ~new_n2768_;
  assign n2700_i2 = new_n1299_;
  assign n2701_i2 = new_n1301_;
  assign n2733_i2 = new_n1359_;
  assign n2734_i2 = new_n1361_;
  assign n2744_i2 = new_n1381_;
  assign n2747_i2 = new_n1387_;
  assign n2754_i2 = new_n2837_;
  assign n2755_i2 = new_n2886_;
  assign n2756_i2 = new_n2839_;
  assign G1609_i2 = new_n2797_;
  assign G1625_i2 = new_n2816_;
  assign G738_i2 = ~new_n2818_;
  assign G755_i2 = ~new_n2812_;
  assign G1511_i2 = ~new_n2815_;
  assign G1522_i2 = G1511_i2;
  assign G1538_i2 = ~new_n2796_;
  assign G1549_i2 = G1538_i2;
  assign G1563_i2 = new_n2801_;
  assign G1584_i2 = new_n2803_;
  assign G1576_i2 = G1584_i2;
  assign G1598_i2 = new_n2802_;
  assign G1395_i2 = ~new_n2807_;
  assign G1410_i2 = ~new_n2809_;
  assign G1420_i2 = G1410_i2;
  assign G1434_i2 = ~new_n2808_;
  assign G1240_i2 = new_n2976_;
  assign n1162_lo_buf_i2 = new_n2912_;
  assign n1102_lo_buf_i2 = new_n2981_;
  assign G359_i2 = new_n2887_;
  assign n982_lo_buf_i2 = new_n3012_;
  assign n1030_lo_buf_i2 = new_n3006_;
  assign n1042_lo_buf_i2 = new_n2984_;
  assign G161_i2 = new_n2980_;
  assign G606_i2 = new_n3020_;
  assign G1118_i2 = new_n3021_;
  assign G1069_i2 = new_n3022_;
  assign G1145_i2 = new_n3023_;
  assign G1209_i2 = new_n3024_;
  assign G1189_i2 = new_n3025_;
  assign G1699_i2 = new_n2863_;
  assign G1702_i2 = G1699_i2;
  assign G1705_i2 = new_n2864_;
  assign G1708_i2 = G1705_i2;
  assign G1684_i2 = new_n2874_;
  assign G1687_i2 = G1684_i2;
  assign G1690_i2 = new_n2875_;
  assign G1693_i2 = G1690_i2;
  assign G1696_i2 = new_n2857_;
  assign G1642_i2 = new_n2867_;
  assign G1645_i2 = new_n2866_;
  assign G1648_i2 = new_n2868_;
  assign G1651_i2 = G1648_i2;
  assign G1654_i2 = new_n2855_;
  assign G1657_i2 = new_n2856_;
  assign G1660_i2 = G1657_i2;
  assign n1222_lo_buf_i2 = new_n2999_;
  assign n1330_lo_buf_i2 = new_n3001_;
  assign G123_i2 = new_n3013_;
  assign G142_i2 = new_n2985_;
  assign n1306_lo_buf_i2 = new_n2895_;
  assign n1150_lo_buf_i2 = new_n2997_;
  assign G175_i2 = new_n2998_;
  assign G241_i2 = new_n3000_;
  assign G356_i2 = G142_i2;
  assign G989_i2 = new_n2991_;
  assign G984_i2 = new_n2995_;
  assign G1009_i2 = new_n2993_;
  assign G1012_i2 = new_n3027_;
  assign n958_lo_buf_i2 = new_n3031_;
  assign n1114_lo_buf_i2 = new_n3035_;
  assign G182_i2 = new_n2898_;
  assign G1215_i2 = ~new_n1945_;
  assign G971_i2 = ~new_n1949_;
  assign G938_i2 = new_n1950_;
  assign G1198_i2 = ~new_n1951_;
  assign G1203_i2 = new_n1966_;
  assign G1218_i2 = new_n1967_;
  assign G785_i2 = G606_i2;
  assign G1168_i2 = G1118_i2;
  assign G1130_i2 = G1069_i2;
  assign G1185_i2 = G1145_i2;
  assign G1250_i2 = G1209_i2;
  assign G1225_i2 = G1189_i2;
  assign G1791_i2 = new_n1974_;
  assign G1788_i2 = new_n1978_;
  assign G981_i2 = new_n3038_;
  assign G1031_i2 = G989_i2;
  assign G1015_i2 = new_n3040_;
  assign G1062_i2 = G1012_i2;
  assign n970_lo_buf_i2 = new_n3042_;
  assign n1006_lo_buf_i2 = new_n3045_;
  assign n1078_lo_buf_i2 = new_n3048_;
  assign n1126_lo_buf_i2 = new_n3052_;
  assign G116_i2 = n958_lo_buf_i2;
  assign G165_i2 = n1114_lo_buf_i2;
  assign n1234_lo_buf_i2 = new_n841_;
  assign n1246_lo_buf_i2 = new_n847_;
  assign n1258_lo_buf_i2 = new_n853_;
  assign n1270_lo_buf_i2 = new_n859_;
  assign G368_i2 = new_n2982_;
  assign G428_i2 = G123_i2;
  assign G212_i2 = n1306_lo_buf_i2;
  assign G841_i2 = new_n1997_;
  assign G788_i2 = new_n1998_;
  assign n1186_lo_buf_i2 = new_n2987_;
  assign G391_i2 = new_n1999_;
  assign G387_i2 = new_n2000_;
  assign G645_i2 = new_n3055_;
  assign G1140_i2 = new_n2025_;
  assign G1178_i2 = new_n2058_;
  assign G1370_i2 = new_n2085_;
  assign G1205_i2 = new_n2116_;
  assign G1357_i2 = new_n2137_;
  assign G816_i2 = new_n3056_;
  assign G1369_i2 = new_n2151_;
  assign G901_i2 = new_n3058_;
  assign G1056_i2 = G981_i2;
  assign G1107_i2 = new_n2992_;
  assign G1087_i2 = G1015_i2;
  assign G1135_i2 = new_n3028_;
  assign n1018_lo_buf_i2 = new_n3060_;
  assign n1090_lo_buf_i2 = new_n3062_;
  assign G119_i2 = n970_lo_buf_i2;
  assign G131_i2 = n1006_lo_buf_i2;
  assign G154_i2 = n1078_lo_buf_i2;
  assign G169_i2 = n1126_lo_buf_i2;
  assign G338_i2 = new_n3030_;
  assign n1171_lo_buf_i2 = new_n825_;
  assign n1195_lo_buf_i2 = new_n831_;
  assign G419_i2 = new_n2877_;
  assign G425_i2 = new_n1307_;
  assign G497_i2 = n2754_i2;
  assign G416_i2 = G359_i2;
  assign G491_i2 = new_n3014_;
  assign G500_i2 = n1030_lo_buf_i2;
  assign G353_i2 = new_n2155_;
  assign G641_i2 = G645_i2;
  assign G1117_i2 = new_n2156_;
  assign G1096_i2 = ~new_n2157_;
  assign G1143_i2 = new_n2158_;
  assign G1112_i2 = new_n2159_;
  assign n1138_lo_buf_i2 = new_n813_;
  assign n1210_lo_buf_i2 = new_n835_;
  assign G687_i2 = G368_i2;
  assign G541_i2 = G491_i2;
  assign G802_i2 = new_n2166_;
  assign G813_i2 = new_n2169_;
  assign G810_i2 = new_n2172_;
  assign G987_i2 = new_n2181_;
  assign G898_i2 = G901_i2;
  assign n946_lo_buf_i2 = new_n3063_;
  assign n1054_lo_buf_i2 = new_n3064_;
  assign G728_i2 = new_n3054_;
  assign G856_i2 = G816_i2;
  assign G831_i2 = new_n2184_;
  assign G942_i2 = new_n3057_;
  assign G1099_i2 = new_n3037_;
  assign G1154_i2 = G1107_i2;
  assign G1131_i2 = new_n3039_;
  assign G1169_i2 = G1135_i2;
  assign G134_i2 = n1018_lo_buf_i2;
  assign G157_i2 = n1090_lo_buf_i2;
  assign G470_i2 = new_n3043_;
  assign G344_i2 = new_n3046_;
  assign G362_i2 = new_n3049_;
  assign G482_i2 = new_n3051_;
  assign G660_i2 = new_n3032_;
  assign G672_i2 = new_n3034_;
  assign n1096_lo_buf_i2 = new_n735_;
  assign G479_i2 = new_n3053_;
  assign G669_i2 = new_n3036_;
  assign n994_lo_buf_i2 = new_n717_;
  assign n1066_lo_buf_i2 = new_n729_;
  assign G112_i2 = n946_lo_buf_i2;
  assign G147_i2 = n1054_lo_buf_i2;
  assign G473_i2 = new_n3059_;
  assign G488_i2 = new_n3061_;
  assign G589_i2 = G470_i2;
  assign G663_i2 = G344_i2;
  assign G684_i2 = G362_i2;
  assign G605_i2 = G479_i2;
  assign G774_i2 = G660_i2;
  assign G782_i2 = G669_i2;
  assign new_n2535_ = new_n1090_;
  assign new_n2536_ = new_n1086_;
  assign new_n2537_ = new_n1089_;
  assign new_n2538_ = new_n1085_;
  assign new_n2539_ = new_n1425_;
  assign new_n2540_ = new_n2539_;
  assign new_n2541_ = new_n1095_;
  assign new_n2542_ = new_n2541_;
  assign new_n2543_ = new_n2542_;
  assign new_n2544_ = new_n2542_;
  assign new_n2545_ = new_n2541_;
  assign new_n2546_ = new_n1426_;
  assign new_n2547_ = new_n2546_;
  assign new_n2548_ = new_n1096_;
  assign new_n2549_ = new_n2548_;
  assign new_n2550_ = new_n2549_;
  assign new_n2551_ = new_n2548_;
  assign new_n2552_ = new_n1102_;
  assign new_n2553_ = new_n2552_;
  assign new_n2554_ = new_n2553_;
  assign new_n2555_ = new_n2554_;
  assign new_n2556_ = new_n2554_;
  assign new_n2557_ = new_n2553_;
  assign new_n2558_ = new_n2552_;
  assign new_n2559_ = new_n2558_;
  assign new_n2560_ = new_n2558_;
  assign new_n2561_ = new_n1101_;
  assign new_n2562_ = new_n2561_;
  assign new_n2563_ = new_n2561_;
  assign new_n2564_ = new_n1082_;
  assign new_n2565_ = new_n2564_;
  assign new_n2566_ = new_n2565_;
  assign new_n2567_ = new_n2565_;
  assign new_n2568_ = new_n2564_;
  assign new_n2569_ = new_n2568_;
  assign new_n2570_ = new_n2568_;
  assign new_n2571_ = new_n1081_;
  assign new_n2572_ = new_n2571_;
  assign new_n2573_ = new_n2572_;
  assign new_n2574_ = new_n2572_;
  assign new_n2575_ = new_n2571_;
  assign new_n2576_ = new_n2575_;
  assign new_n2577_ = new_n2575_;
  assign new_n2578_ = new_n1093_;
  assign new_n2579_ = new_n2578_;
  assign new_n2580_ = new_n2579_;
  assign new_n2581_ = new_n2579_;
  assign new_n2582_ = new_n2578_;
  assign new_n2583_ = new_n1094_;
  assign new_n2584_ = new_n1436_;
  assign new_n2585_ = new_n1106_;
  assign new_n2586_ = new_n2585_;
  assign new_n2587_ = new_n2586_;
  assign new_n2588_ = new_n2586_;
  assign new_n2589_ = new_n2585_;
  assign new_n2590_ = new_n2589_;
  assign new_n2591_ = new_n1437_;
  assign new_n2592_ = new_n1105_;
  assign new_n2593_ = new_n2592_;
  assign new_n2594_ = new_n2593_;
  assign new_n2595_ = new_n2593_;
  assign new_n2596_ = new_n2592_;
  assign new_n2597_ = new_n1104_;
  assign new_n2598_ = new_n2597_;
  assign new_n2599_ = new_n2598_;
  assign new_n2600_ = new_n2597_;
  assign new_n2601_ = new_n1103_;
  assign new_n2602_ = new_n2601_;
  assign new_n2603_ = new_n2601_;
  assign new_n2604_ = new_n1097_;
  assign new_n2605_ = new_n2604_;
  assign new_n2606_ = new_n2604_;
  assign new_n2607_ = new_n1098_;
  assign new_n2608_ = new_n2607_;
  assign new_n2609_ = new_n1088_;
  assign new_n2610_ = new_n2609_;
  assign new_n2611_ = new_n1087_;
  assign new_n2612_ = new_n2611_;
  assign new_n2613_ = new_n1099_;
  assign new_n2614_ = new_n2613_;
  assign new_n2615_ = new_n2613_;
  assign new_n2616_ = new_n1100_;
  assign new_n2617_ = new_n2616_;
  assign new_n2618_ = new_n2616_;
  assign new_n2619_ = new_n1084_;
  assign new_n2620_ = new_n2619_;
  assign new_n2621_ = new_n2620_;
  assign new_n2622_ = new_n2620_;
  assign new_n2623_ = new_n2619_;
  assign new_n2624_ = new_n2623_;
  assign new_n2625_ = new_n2623_;
  assign new_n2626_ = new_n1083_;
  assign new_n2627_ = new_n2626_;
  assign new_n2628_ = new_n2627_;
  assign new_n2629_ = new_n2627_;
  assign new_n2630_ = new_n2626_;
  assign new_n2631_ = new_n2630_;
  assign new_n2632_ = new_n2630_;
  assign new_n2633_ = new_n1092_;
  assign new_n2634_ = new_n1091_;
  assign new_n2635_ = new_n1472_;
  assign new_n2636_ = new_n1473_;
  assign new_n2637_ = new_n1108_;
  assign new_n2638_ = new_n1107_;
  assign new_n2639_ = new_n1079_;
  assign new_n2640_ = new_n2639_;
  assign new_n2641_ = new_n2639_;
  assign new_n2642_ = new_n1080_;
  assign new_n2643_ = new_n1503_;
  assign new_n2644_ = new_n2643_;
  assign new_n2645_ = new_n2643_;
  assign new_n2646_ = new_n1504_;
  assign new_n2647_ = new_n2646_;
  assign new_n2648_ = new_n2646_;
  assign new_n2649_ = new_n1523_;
  assign new_n2650_ = new_n1077_;
  assign new_n2651_ = new_n2650_;
  assign new_n2652_ = new_n1541_;
  assign new_n2653_ = new_n2652_;
  assign new_n2654_ = new_n2652_;
  assign new_n2655_ = new_n1542_;
  assign new_n2656_ = new_n2655_;
  assign new_n2657_ = new_n1543_;
  assign new_n2658_ = new_n1544_;
  assign new_n2659_ = new_n1602_;
  assign new_n2660_ = new_n891_;
  assign new_n2661_ = new_n2660_;
  assign new_n2662_ = new_n1606_;
  assign new_n2663_ = new_n2662_;
  assign new_n2664_ = new_n2663_;
  assign new_n2665_ = new_n2663_;
  assign new_n2666_ = new_n2662_;
  assign new_n2667_ = new_n2666_;
  assign new_n2668_ = new_n2666_;
  assign new_n2669_ = new_n1612_;
  assign new_n2670_ = new_n2669_;
  assign new_n2671_ = new_n1616_;
  assign new_n2672_ = new_n1642_;
  assign new_n2673_ = new_n2672_;
  assign new_n2674_ = new_n2673_;
  assign new_n2675_ = new_n2673_;
  assign new_n2676_ = new_n2672_;
  assign new_n2677_ = new_n2676_;
  assign new_n2678_ = new_n1652_;
  assign new_n2679_ = new_n902_;
  assign new_n2680_ = new_n1651_;
  assign new_n2681_ = new_n901_;
  assign new_n2682_ = new_n884_;
  assign new_n2683_ = new_n2682_;
  assign new_n2684_ = new_n2683_;
  assign new_n2685_ = new_n2683_;
  assign new_n2686_ = new_n2682_;
  assign new_n2687_ = new_n883_;
  assign new_n2688_ = new_n2687_;
  assign new_n2689_ = new_n2688_;
  assign new_n2690_ = new_n2688_;
  assign new_n2691_ = new_n2687_;
  assign new_n2692_ = new_n1641_;
  assign new_n2693_ = new_n2692_;
  assign new_n2694_ = new_n2693_;
  assign new_n2695_ = new_n2693_;
  assign new_n2696_ = new_n2692_;
  assign new_n2697_ = new_n895_;
  assign new_n2698_ = new_n2697_;
  assign new_n2699_ = new_n2698_;
  assign new_n2700_ = new_n2697_;
  assign new_n2701_ = new_n1668_;
  assign new_n2702_ = new_n2701_;
  assign new_n2703_ = new_n2702_;
  assign new_n2704_ = new_n2702_;
  assign new_n2705_ = new_n2701_;
  assign new_n2706_ = new_n1676_;
  assign new_n2707_ = new_n1670_;
  assign new_n2708_ = new_n1677_;
  assign new_n2709_ = new_n1671_;
  assign new_n2710_ = new_n896_;
  assign new_n2711_ = new_n2710_;
  assign new_n2712_ = new_n2710_;
  assign new_n2713_ = new_n1022_;
  assign new_n2714_ = new_n1021_;
  assign new_n2715_ = new_n1739_;
  assign new_n2716_ = new_n1732_;
  assign new_n2717_ = new_n1738_;
  assign new_n2718_ = new_n1733_;
  assign new_n2719_ = new_n1774_;
  assign new_n2720_ = new_n1767_;
  assign new_n2721_ = new_n1773_;
  assign new_n2722_ = new_n1768_;
  assign new_n2723_ = new_n1797_;
  assign new_n2724_ = new_n1793_;
  assign new_n2725_ = new_n1796_;
  assign new_n2726_ = new_n1792_;
  assign new_n2727_ = new_n899_;
  assign new_n2728_ = new_n897_;
  assign new_n2729_ = new_n900_;
  assign new_n2730_ = new_n898_;
  assign new_n2731_ = new_n1269_;
  assign new_n2732_ = new_n2731_;
  assign new_n2733_ = new_n1011_;
  assign new_n2734_ = new_n1270_;
  assign new_n2735_ = new_n1271_;
  assign new_n2736_ = new_n2735_;
  assign new_n2737_ = new_n1111_;
  assign new_n2738_ = new_n1272_;
  assign new_n2739_ = new_n1275_;
  assign new_n2740_ = new_n1262_;
  assign new_n2741_ = new_n2740_;
  assign new_n2742_ = new_n2741_;
  assign new_n2743_ = new_n2741_;
  assign new_n2744_ = new_n2740_;
  assign new_n2745_ = new_n1261_;
  assign new_n2746_ = new_n2745_;
  assign new_n2747_ = new_n2746_;
  assign new_n2748_ = new_n2746_;
  assign new_n2749_ = new_n2745_;
  assign new_n2750_ = new_n1277_;
  assign new_n2751_ = new_n1281_;
  assign new_n2752_ = new_n1341_;
  assign new_n2753_ = new_n1184_;
  assign new_n2754_ = new_n2753_;
  assign new_n2755_ = new_n2753_;
  assign new_n2756_ = new_n1183_;
  assign new_n2757_ = new_n2756_;
  assign new_n2758_ = new_n2756_;
  assign new_n2759_ = new_n1315_;
  assign new_n2760_ = new_n1827_;
  assign new_n2761_ = new_n1814_;
  assign new_n2762_ = new_n1249_;
  assign new_n2763_ = new_n2762_;
  assign new_n2764_ = new_n1828_;
  assign new_n2765_ = new_n1843_;
  assign new_n2766_ = new_n2765_;
  assign new_n2767_ = new_n1830_;
  assign new_n2768_ = new_n1846_;
  assign new_n2769_ = new_n2768_;
  assign new_n2770_ = new_n1832_;
  assign new_n2771_ = new_n1178_;
  assign new_n2772_ = new_n978_;
  assign new_n2773_ = new_n2772_;
  assign new_n2774_ = new_n1834_;
  assign new_n2775_ = new_n2774_;
  assign new_n2776_ = new_n2774_;
  assign new_n2777_ = new_n1853_;
  assign new_n2778_ = new_n1823_;
  assign new_n2779_ = new_n1816_;
  assign new_n2780_ = new_n1825_;
  assign new_n2781_ = new_n1251_;
  assign new_n2782_ = new_n2781_;
  assign new_n2783_ = new_n1255_;
  assign new_n2784_ = new_n2783_;
  assign new_n2785_ = new_n1818_;
  assign new_n2786_ = new_n1253_;
  assign new_n2787_ = new_n2786_;
  assign new_n2788_ = new_n1820_;
  assign new_n2789_ = new_n1876_;
  assign new_n2790_ = new_n1368_;
  assign new_n2791_ = new_n1875_;
  assign new_n2792_ = new_n1367_;
  assign new_n2793_ = new_n2792_;
  assign new_n2794_ = new_n1860_;
  assign new_n2795_ = new_n2794_;
  assign new_n2796_ = new_n2794_;
  assign new_n2797_ = new_n1847_;
  assign new_n2798_ = new_n1867_;
  assign new_n2799_ = new_n2798_;
  assign new_n2800_ = new_n2799_;
  assign new_n2801_ = new_n2799_;
  assign new_n2802_ = new_n2798_;
  assign new_n2803_ = new_n2802_;
  assign new_n2804_ = new_n1874_;
  assign new_n2805_ = new_n2804_;
  assign new_n2806_ = new_n2805_;
  assign new_n2807_ = new_n2805_;
  assign new_n2808_ = new_n2804_;
  assign new_n2809_ = new_n2808_;
  assign new_n2810_ = new_n1858_;
  assign new_n2811_ = new_n2810_;
  assign new_n2812_ = new_n2810_;
  assign new_n2813_ = new_n1859_;
  assign new_n2814_ = new_n2813_;
  assign new_n2815_ = new_n2813_;
  assign new_n2816_ = new_n1848_;
  assign new_n2817_ = new_n1898_;
  assign new_n2818_ = new_n1854_;
  assign new_n2819_ = new_n2818_;
  assign new_n2820_ = new_n1903_;
  assign new_n2821_ = new_n1399_;
  assign new_n2822_ = new_n1397_;
  assign new_n2823_ = new_n1400_;
  assign new_n2824_ = new_n1398_;
  assign new_n2825_ = new_n1407_;
  assign new_n2826_ = new_n2825_;
  assign new_n2827_ = new_n2825_;
  assign new_n2828_ = new_n1408_;
  assign new_n2829_ = new_n2828_;
  assign new_n2830_ = new_n2828_;
  assign new_n2831_ = new_n1415_;
  assign new_n2832_ = new_n1409_;
  assign new_n2833_ = new_n1416_;
  assign new_n2834_ = new_n1410_;
  assign new_n2835_ = new_n1401_;
  assign new_n2836_ = new_n2835_;
  assign new_n2837_ = new_n2835_;
  assign new_n2838_ = new_n1402_;
  assign new_n2839_ = new_n1405_;
  assign new_n2840_ = new_n2839_;
  assign new_n2841_ = new_n1406_;
  assign new_n2842_ = new_n1944_;
  assign new_n2843_ = new_n1028_;
  assign new_n2844_ = new_n1948_;
  assign new_n2845_ = new_n1053_;
  assign new_n2846_ = new_n1953_;
  assign new_n2847_ = new_n965_;
  assign new_n2848_ = new_n1952_;
  assign new_n2849_ = new_n966_;
  assign new_n2850_ = new_n1965_;
  assign new_n2851_ = new_n1962_;
  assign new_n2852_ = new_n1905_;
  assign new_n2853_ = new_n2852_;
  assign new_n2854_ = new_n2853_;
  assign new_n2855_ = new_n2853_;
  assign new_n2856_ = new_n2852_;
  assign new_n2857_ = new_n1900_;
  assign new_n2858_ = new_n1895_;
  assign new_n2859_ = new_n2858_;
  assign new_n2860_ = new_n2859_;
  assign new_n2861_ = new_n2859_;
  assign new_n2862_ = new_n2858_;
  assign new_n2863_ = new_n2862_;
  assign new_n2864_ = new_n2862_;
  assign new_n2865_ = new_n1904_;
  assign new_n2866_ = new_n2865_;
  assign new_n2867_ = new_n2866_;
  assign new_n2868_ = new_n2865_;
  assign new_n2869_ = new_n1899_;
  assign new_n2870_ = new_n2869_;
  assign new_n2871_ = new_n2870_;
  assign new_n2872_ = new_n2870_;
  assign new_n2873_ = new_n2869_;
  assign new_n2874_ = new_n2873_;
  assign new_n2875_ = new_n2873_;
  assign new_n2876_ = new_n1311_;
  assign new_n2877_ = new_n1303_;
  assign new_n2878_ = new_n2877_;
  assign new_n2879_ = new_n1312_;
  assign new_n2880_ = new_n1304_;
  assign new_n2881_ = new_n1417_;
  assign new_n2882_ = new_n1411_;
  assign new_n2883_ = new_n1418_;
  assign new_n2884_ = new_n1412_;
  assign new_n2885_ = new_n1403_;
  assign new_n2886_ = new_n2885_;
  assign new_n2887_ = new_n2885_;
  assign new_n2888_ = new_n1069_;
  assign new_n2889_ = new_n1067_;
  assign new_n2890_ = new_n2889_;
  assign new_n2891_ = new_n2889_;
  assign new_n2892_ = new_n1169_;
  assign new_n2893_ = new_n881_;
  assign new_n2894_ = new_n2893_;
  assign new_n2895_ = new_n2893_;
  assign new_n2896_ = new_n1343_;
  assign new_n2897_ = new_n2896_;
  assign new_n2898_ = new_n2896_;
  assign new_n2899_ = new_n1353_;
  assign new_n2900_ = new_n1318_;
  assign new_n2901_ = new_n1354_;
  assign new_n2902_ = new_n1317_;
  assign new_n2903_ = new_n1351_;
  assign new_n2904_ = new_n1320_;
  assign new_n2905_ = new_n1352_;
  assign new_n2906_ = new_n1319_;
  assign new_n2907_ = new_n2011_;
  assign new_n2908_ = new_n2006_;
  assign new_n2909_ = new_n2012_;
  assign new_n2910_ = new_n2005_;
  assign new_n2911_ = new_n1344_;
  assign new_n2912_ = new_n821_;
  assign new_n2913_ = new_n1358_;
  assign new_n2914_ = new_n1331_;
  assign new_n2915_ = new_n1357_;
  assign new_n2916_ = new_n1332_;
  assign new_n2917_ = new_n1349_;
  assign new_n2918_ = new_n1324_;
  assign new_n2919_ = new_n1350_;
  assign new_n2920_ = new_n1323_;
  assign new_n2921_ = new_n2036_;
  assign new_n2922_ = new_n2031_;
  assign new_n2923_ = new_n2037_;
  assign new_n2924_ = new_n2030_;
  assign new_n2925_ = new_n1327_;
  assign new_n2926_ = new_n1322_;
  assign new_n2927_ = new_n1328_;
  assign new_n2928_ = new_n1321_;
  assign new_n2929_ = new_n2049_;
  assign new_n2930_ = new_n1052_;
  assign new_n2931_ = new_n2048_;
  assign new_n2932_ = new_n1051_;
  assign new_n2933_ = new_n1345_;
  assign new_n2934_ = new_n1325_;
  assign new_n2935_ = new_n1346_;
  assign new_n2936_ = new_n1326_;
  assign new_n2937_ = new_n2064_;
  assign new_n2938_ = new_n1839_;
  assign new_n2939_ = new_n2938_;
  assign new_n2940_ = new_n2063_;
  assign new_n2941_ = new_n1840_;
  assign new_n2942_ = new_n2076_;
  assign new_n2943_ = new_n1233_;
  assign new_n2944_ = new_n2943_;
  assign new_n2945_ = new_n2943_;
  assign new_n2946_ = new_n2075_;
  assign new_n2947_ = new_n1234_;
  assign new_n2948_ = new_n2097_;
  assign new_n2949_ = new_n2090_;
  assign new_n2950_ = new_n2096_;
  assign new_n2951_ = new_n2091_;
  assign new_n2952_ = new_n1313_;
  assign new_n2953_ = new_n2106_;
  assign new_n2954_ = new_n1068_;
  assign new_n2955_ = new_n2107_;
  assign new_n2956_ = new_n1837_;
  assign new_n2957_ = new_n2956_;
  assign new_n2958_ = new_n1075_;
  assign new_n2959_ = new_n2958_;
  assign new_n2960_ = new_n1838_;
  assign new_n2961_ = new_n1076_;
  assign new_n2962_ = new_n2128_;
  assign new_n2963_ = new_n1356_;
  assign new_n2964_ = new_n2127_;
  assign new_n2965_ = new_n1355_;
  assign new_n2966_ = new_n2965_;
  assign new_n2967_ = new_n1380_;
  assign new_n2968_ = new_n2967_;
  assign new_n2969_ = new_n1379_;
  assign new_n2970_ = new_n2969_;
  assign new_n2971_ = new_n2142_;
  assign new_n2972_ = new_n1329_;
  assign new_n2973_ = new_n2972_;
  assign new_n2974_ = new_n2141_;
  assign new_n2975_ = new_n1330_;
  assign new_n2976_ = new_n1881_;
  assign new_n2977_ = new_n796_;
  assign new_n2978_ = new_n2977_;
  assign new_n2979_ = new_n1395_;
  assign new_n2980_ = new_n2979_;
  assign new_n2981_ = new_n2980_;
  assign new_n2982_ = new_n2979_;
  assign new_n2983_ = new_n795_;
  assign new_n2984_ = new_n2983_;
  assign new_n2985_ = new_n2983_;
  assign new_n2986_ = new_n894_;
  assign new_n2987_ = new_n827_;
  assign new_n2988_ = new_n1914_;
  assign new_n2989_ = new_n2988_;
  assign new_n2990_ = new_n2989_;
  assign new_n2991_ = new_n2989_;
  assign new_n2992_ = new_n2988_;
  assign new_n2993_ = new_n1932_;
  assign new_n2994_ = new_n2993_;
  assign new_n2995_ = new_n1923_;
  assign new_n2996_ = new_n2995_;
  assign new_n2997_ = new_n817_;
  assign new_n2998_ = new_n837_;
  assign new_n2999_ = new_n2998_;
  assign new_n3000_ = new_n893_;
  assign new_n3001_ = new_n3000_;
  assign new_n3002_ = new_n1247_;
  assign new_n3003_ = new_n1248_;
  assign new_n3004_ = new_n791_;
  assign new_n3005_ = new_n3004_;
  assign new_n3006_ = new_n3004_;
  assign new_n3007_ = new_n792_;
  assign new_n3008_ = new_n1385_;
  assign new_n3009_ = new_n1386_;
  assign new_n3010_ = new_n781_;
  assign new_n3011_ = new_n3010_;
  assign new_n3012_ = new_n3011_;
  assign new_n3013_ = new_n3011_;
  assign new_n3014_ = new_n3010_;
  assign new_n3015_ = new_n867_;
  assign new_n3016_ = new_n875_;
  assign new_n3017_ = new_n889_;
  assign new_n3018_ = new_n977_;
  assign new_n3019_ = new_n3018_;
  assign new_n3020_ = new_n1025_;
  assign new_n3021_ = new_n1035_;
  assign new_n3022_ = new_n1041_;
  assign new_n3023_ = new_n1885_;
  assign new_n3024_ = new_n1888_;
  assign new_n3025_ = new_n1891_;
  assign new_n3026_ = new_n1941_;
  assign new_n3027_ = new_n3026_;
  assign new_n3028_ = new_n3026_;
  assign new_n3029_ = new_n711_;
  assign new_n3030_ = new_n3029_;
  assign new_n3031_ = new_n3030_;
  assign new_n3032_ = new_n3029_;
  assign new_n3033_ = new_n737_;
  assign new_n3034_ = new_n3033_;
  assign new_n3035_ = new_n3034_;
  assign new_n3036_ = new_n3033_;
  assign new_n3037_ = new_n1987_;
  assign new_n3038_ = new_n3037_;
  assign new_n3039_ = new_n1996_;
  assign new_n3040_ = new_n3039_;
  assign new_n3041_ = new_n713_;
  assign new_n3042_ = new_n3041_;
  assign new_n3043_ = new_n3041_;
  assign new_n3044_ = new_n719_;
  assign new_n3045_ = new_n3044_;
  assign new_n3046_ = new_n3044_;
  assign new_n3047_ = new_n731_;
  assign new_n3048_ = new_n3047_;
  assign new_n3049_ = new_n3047_;
  assign new_n3050_ = new_n739_;
  assign new_n3051_ = new_n3050_;
  assign new_n3052_ = new_n3051_;
  assign new_n3053_ = new_n3050_;
  assign new_n3054_ = new_n1309_;
  assign new_n3055_ = new_n3054_;
  assign new_n3056_ = new_n2140_;
  assign new_n3057_ = new_n2154_;
  assign new_n3058_ = new_n3057_;
  assign new_n3059_ = new_n721_;
  assign new_n3060_ = new_n3059_;
  assign new_n3061_ = new_n733_;
  assign new_n3062_ = new_n3061_;
  assign new_n3063_ = new_n709_;
  assign new_n3064_ = new_n727_;
  always @ (posedge clock) begin
    n949_lo <= n949_li;
    n961_lo <= n961_li;
    n973_lo <= n973_li;
    n976_lo <= n976_li;
    n985_lo <= n985_li;
    n997_lo <= n997_li;
    n1009_lo <= n1009_li;
    n1021_lo <= n1021_li;
    n1024_lo <= n1024_li;
    n1033_lo <= n1033_li;
    n1036_lo <= n1036_li;
    n1045_lo <= n1045_li;
    n1057_lo <= n1057_li;
    n1069_lo <= n1069_li;
    n1081_lo <= n1081_li;
    n1093_lo <= n1093_li;
    n1105_lo <= n1105_li;
    n1117_lo <= n1117_li;
    n1129_lo <= n1129_li;
    n1132_lo <= n1132_li;
    n1141_lo <= n1141_li;
    n1144_lo <= n1144_li;
    n1156_lo <= n1156_li;
    n1159_lo <= n1159_li;
    n1165_lo <= n1165_li;
    n1168_lo <= n1168_li;
    n1180_lo <= n1180_li;
    n1189_lo <= n1189_li;
    n1192_lo <= n1192_li;
    n1201_lo <= n1201_li;
    n1204_lo <= n1204_li;
    n1216_lo <= n1216_li;
    n1228_lo <= n1228_li;
    n1231_lo <= n1231_li;
    n1237_lo <= n1237_li;
    n1240_lo <= n1240_li;
    n1243_lo <= n1243_li;
    n1249_lo <= n1249_li;
    n1252_lo <= n1252_li;
    n1255_lo <= n1255_li;
    n1261_lo <= n1261_li;
    n1264_lo <= n1264_li;
    n1267_lo <= n1267_li;
    n1273_lo <= n1273_li;
    n1276_lo <= n1276_li;
    n1279_lo <= n1279_li;
    n1282_lo <= n1282_li;
    n1285_lo <= n1285_li;
    n1288_lo <= n1288_li;
    n1291_lo <= n1291_li;
    n1294_lo <= n1294_li;
    n1297_lo <= n1297_li;
    n1300_lo <= n1300_li;
    n1303_lo <= n1303_li;
    n1309_lo <= n1309_li;
    n1312_lo <= n1312_li;
    n1315_lo <= n1315_li;
    n1318_lo <= n1318_li;
    n1321_lo <= n1321_li;
    n1324_lo <= n1324_li;
    n1333_lo <= n1333_li;
    n1874_o2 <= n1874_i2;
    n2180_o2 <= n2180_i2;
    n2372_o2 <= n2372_i2;
    n2190_o2 <= n2190_i2;
    n2191_o2 <= n2191_i2;
    n2212_o2 <= n2212_i2;
    n2213_o2 <= n2213_i2;
    n2214_o2 <= n2214_i2;
    n2215_o2 <= n2215_i2;
    n2275_o2 <= n2275_i2;
    n2276_o2 <= n2276_i2;
    n2290_o2 <= n2290_i2;
    n2291_o2 <= n2291_i2;
    n2681_o2 <= n2681_i2;
    n2680_o2 <= n2680_i2;
    n2683_o2 <= n2683_i2;
    n2684_o2 <= n2684_i2;
    n2686_o2 <= n2686_i2;
    n2319_o2 <= n2319_i2;
    n2320_o2 <= n2320_i2;
    n304_inv <= n2321_i2;
    G554_o2 <= G554_i2;
    G557_o2 <= G557_i2;
    G185_o2 <= G185_i2;
    G188_o2 <= G188_i2;
    G191_o2 <= G191_i2;
    G194_o2 <= G194_i2;
    G1182_o2 <= G1182_i2;
    G1222_o2 <= G1222_i2;
    G1247_o2 <= G1247_i2;
    G1371_o2 <= G1371_i2;
    G1383_o2 <= G1383_i2;
    G1386_o2 <= G1386_i2;
    n2416_o2 <= n2416_i2;
    n2428_o2 <= n2428_i2;
    n2438_o2 <= n2438_i2;
    n2439_o2 <= n2439_i2;
    n2440_o2 <= n2440_i2;
    n2444_o2 <= n2444_i2;
    n2497_o2 <= n2497_i2;
    n2498_o2 <= n2498_i2;
    n2503_o2 <= n2503_i2;
    n2505_o2 <= n2505_i2;
    n2529_o2 <= n2529_i2;
    n2562_o2 <= n2562_i2;
    n2570_o2 <= n2570_i2;
    n2571_o2 <= n2571_i2;
    n2574_o2 <= n2574_i2;
    n2575_o2 <= n2575_i2;
    G546_o2 <= G546_i2;
    G550_o2 <= G550_i2;
    n2633_o2 <= n2633_i2;
    n2639_o2 <= n2639_i2;
    n2642_o2 <= n2642_i2;
    n2645_o2 <= n2645_i2;
    n2679_o2 <= n2679_i2;
    n2662_o2 <= n2662_i2;
    n2724_o2 <= n2724_i2;
    G382_o2 <= G382_i2;
    G199_o2 <= G199_i2;
    G202_o2 <= G202_i2;
    G225_o2 <= G225_i2;
    G248_o2 <= G248_i2;
    G260_o2 <= G260_i2;
    n2716_o2 <= n2716_i2;
    n2737_o2 <= n2737_i2;
    n1174_lo_buf_o2 <= n1174_lo_buf_i2;
    n1198_lo_buf_o2 <= n1198_lo_buf_i2;
    G371_o2 <= G371_i2;
    G1059_o2 <= G1059_i2;
    n2586_o2 <= n2586_i2;
    n2587_o2 <= n2587_i2;
    n460_inv <= G1019_i2;
    n2648_o2 <= n2648_i2;
    n2649_o2 <= n2649_i2;
    n2650_o2 <= n2650_i2;
    n2651_o2 <= n2651_i2;
    n2652_o2 <= n2652_i2;
    G365_o2 <= G365_i2;
    G1496_o2 <= G1496_i2;
    G1502_o2 <= G1502_i2;
    n2700_o2 <= n2700_i2;
    n2701_o2 <= n2701_i2;
    n2733_o2 <= n2733_i2;
    n2734_o2 <= n2734_i2;
    n2744_o2 <= n2744_i2;
    n2747_o2 <= n2747_i2;
    n2754_o2 <= n2754_i2;
    n2755_o2 <= n2755_i2;
    n511_inv <= n2756_i2;
    G1609_o2 <= G1609_i2;
    G1625_o2 <= G1625_i2;
    G738_o2 <= G738_i2;
    G755_o2 <= G755_i2;
    G1511_o2 <= G1511_i2;
    G1522_o2 <= G1522_i2;
    G1538_o2 <= G1538_i2;
    G1549_o2 <= G1549_i2;
    G1563_o2 <= G1563_i2;
    G1584_o2 <= G1584_i2;
    G1576_o2 <= G1576_i2;
    G1598_o2 <= G1598_i2;
    G1395_o2 <= G1395_i2;
    G1410_o2 <= G1410_i2;
    G1420_o2 <= G1420_i2;
    G1434_o2 <= G1434_i2;
    n562_inv <= G1240_i2;
    n1162_lo_buf_o2 <= n1162_lo_buf_i2;
    n1102_lo_buf_o2 <= n1102_lo_buf_i2;
    G359_o2 <= G359_i2;
    n982_lo_buf_o2 <= n982_lo_buf_i2;
    n1030_lo_buf_o2 <= n1030_lo_buf_i2;
    n1042_lo_buf_o2 <= n1042_lo_buf_i2;
    n583_inv <= G161_i2;
    G606_o2 <= G606_i2;
    G1118_o2 <= G1118_i2;
    G1069_o2 <= G1069_i2;
    G1145_o2 <= G1145_i2;
    G1209_o2 <= G1209_i2;
    G1189_o2 <= G1189_i2;
    G1699_o2 <= G1699_i2;
    G1702_o2 <= G1702_i2;
    G1705_o2 <= G1705_i2;
    G1708_o2 <= G1708_i2;
    G1684_o2 <= G1684_i2;
    G1687_o2 <= G1687_i2;
    G1690_o2 <= G1690_i2;
    G1693_o2 <= G1693_i2;
    G1696_o2 <= G1696_i2;
    G1642_o2 <= G1642_i2;
    G1645_o2 <= G1645_i2;
    G1648_o2 <= G1648_i2;
    G1651_o2 <= G1651_i2;
    G1654_o2 <= G1654_i2;
    G1657_o2 <= G1657_i2;
    G1660_o2 <= G1660_i2;
    n1222_lo_buf_o2 <= n1222_lo_buf_i2;
    n1330_lo_buf_o2 <= n1330_lo_buf_i2;
    n658_inv <= G123_i2;
    n661_inv <= G142_i2;
    n1306_lo_buf_o2 <= n1306_lo_buf_i2;
    n1150_lo_buf_o2 <= n1150_lo_buf_i2;
    G175_o2 <= G175_i2;
    G241_o2 <= G241_i2;
    G356_o2 <= G356_i2;
    G989_o2 <= G989_i2;
    G984_o2 <= G984_i2;
    n685_inv <= G1009_i2;
    n688_inv <= G1012_i2;
    n958_lo_buf_o2 <= n958_lo_buf_i2;
    n1114_lo_buf_o2 <= n1114_lo_buf_i2;
    G182_o2 <= G182_i2;
    G1215_o2 <= G1215_i2;
    G971_o2 <= G971_i2;
    G938_o2 <= G938_i2;
    G1198_o2 <= G1198_i2;
    G1203_o2 <= G1203_i2;
    G1218_o2 <= G1218_i2;
    G785_o2 <= G785_i2;
    G1168_o2 <= G1168_i2;
    G1130_o2 <= G1130_i2;
    G1185_o2 <= G1185_i2;
    G1250_o2 <= G1250_i2;
    G1225_o2 <= G1225_i2;
    G1791_o2 <= G1791_i2;
    G1788_o2 <= G1788_i2;
    G981_o2 <= G981_i2;
    n745_inv <= G1031_i2;
    n748_inv <= G1015_i2;
    G1062_o2 <= G1062_i2;
    n970_lo_buf_o2 <= n970_lo_buf_i2;
    n1006_lo_buf_o2 <= n1006_lo_buf_i2;
    n1078_lo_buf_o2 <= n1078_lo_buf_i2;
    n1126_lo_buf_o2 <= n1126_lo_buf_i2;
    n766_inv <= G116_i2;
    G165_o2 <= G165_i2;
    n1234_lo_buf_o2 <= n1234_lo_buf_i2;
    n1246_lo_buf_o2 <= n1246_lo_buf_i2;
    n1258_lo_buf_o2 <= n1258_lo_buf_i2;
    n1270_lo_buf_o2 <= n1270_lo_buf_i2;
    G368_o2 <= G368_i2;
    G428_o2 <= G428_i2;
    G212_o2 <= G212_i2;
    G841_o2 <= G841_i2;
    G788_o2 <= G788_i2;
    n1186_lo_buf_o2 <= n1186_lo_buf_i2;
    G391_o2 <= G391_i2;
    G387_o2 <= G387_i2;
    G645_o2 <= G645_i2;
    G1140_o2 <= G1140_i2;
    G1178_o2 <= G1178_i2;
    G1370_o2 <= G1370_i2;
    n820_inv <= G1205_i2;
    G1357_o2 <= G1357_i2;
    G816_o2 <= G816_i2;
    G1369_o2 <= G1369_i2;
    G901_o2 <= G901_i2;
    G1056_o2 <= G1056_i2;
    G1107_o2 <= G1107_i2;
    G1087_o2 <= G1087_i2;
    G1135_o2 <= G1135_i2;
    n1018_lo_buf_o2 <= n1018_lo_buf_i2;
    n1090_lo_buf_o2 <= n1090_lo_buf_i2;
    n853_inv <= G119_i2;
    G131_o2 <= G131_i2;
    n859_inv <= G154_i2;
    n862_inv <= G169_i2;
    G338_o2 <= G338_i2;
    n1171_lo_buf_o2 <= n1171_lo_buf_i2;
    n1195_lo_buf_o2 <= n1195_lo_buf_i2;
    G419_o2 <= G419_i2;
    G425_o2 <= G425_i2;
    G497_o2 <= G497_i2;
    G416_o2 <= G416_i2;
    G491_o2 <= G491_i2;
    G500_o2 <= G500_i2;
    G353_o2 <= G353_i2;
    G641_o2 <= G641_i2;
    G1117_o2 <= G1117_i2;
    G1096_o2 <= G1096_i2;
    G1143_o2 <= G1143_i2;
    G1112_o2 <= G1112_i2;
    n1138_lo_buf_o2 <= n1138_lo_buf_i2;
    n1210_lo_buf_o2 <= n1210_lo_buf_i2;
    G687_o2 <= G687_i2;
    G541_o2 <= G541_i2;
    G802_o2 <= G802_i2;
    G813_o2 <= G813_i2;
    G810_o2 <= G810_i2;
    G987_o2 <= G987_i2;
    G898_o2 <= G898_i2;
    n946_lo_buf_o2 <= n946_lo_buf_i2;
    n1054_lo_buf_o2 <= n1054_lo_buf_i2;
    G728_o2 <= G728_i2;
    G856_o2 <= G856_i2;
    n949_1_inv <= G831_i2;
    G942_o2 <= G942_i2;
    G1099_o2 <= G1099_i2;
    G1154_o2 <= G1154_i2;
    G1131_o2 <= G1131_i2;
    G1169_o2 <= G1169_i2;
    G134_o2 <= G134_i2;
    n970_inv <= G157_i2;
    G470_o2 <= G470_i2;
    G344_o2 <= G344_i2;
    G362_o2 <= G362_i2;
    G482_o2 <= G482_i2;
    G660_o2 <= G660_i2;
    G672_o2 <= G672_i2;
    n1096_lo_buf_o2 <= n1096_lo_buf_i2;
    G479_o2 <= G479_i2;
    G669_o2 <= G669_i2;
    n994_lo_buf_o2 <= n994_lo_buf_i2;
    n1066_lo_buf_o2 <= n1066_lo_buf_i2;
    n1006_inv <= G112_i2;
    G147_o2 <= G147_i2;
    G473_o2 <= G473_i2;
    G488_o2 <= G488_i2;
    G589_o2 <= G589_i2;
    G663_o2 <= G663_i2;
    G684_o2 <= G684_i2;
    G605_o2 <= G605_i2;
    G774_o2 <= G774_i2;
    G782_o2 <= G782_i2;
  end
  initial begin
    n949_lo <= 1'b0;
    n961_lo <= 1'b0;
    n973_lo <= 1'b0;
    n976_lo <= 1'b0;
    n985_lo <= 1'b0;
    n997_lo <= 1'b0;
    n1009_lo <= 1'b0;
    n1021_lo <= 1'b0;
    n1024_lo <= 1'b0;
    n1033_lo <= 1'b0;
    n1036_lo <= 1'b0;
    n1045_lo <= 1'b0;
    n1057_lo <= 1'b0;
    n1069_lo <= 1'b0;
    n1081_lo <= 1'b0;
    n1093_lo <= 1'b0;
    n1105_lo <= 1'b0;
    n1117_lo <= 1'b0;
    n1129_lo <= 1'b0;
    n1132_lo <= 1'b0;
    n1141_lo <= 1'b0;
    n1144_lo <= 1'b0;
    n1156_lo <= 1'b0;
    n1159_lo <= 1'b0;
    n1165_lo <= 1'b0;
    n1168_lo <= 1'b0;
    n1180_lo <= 1'b0;
    n1189_lo <= 1'b0;
    n1192_lo <= 1'b0;
    n1201_lo <= 1'b0;
    n1204_lo <= 1'b0;
    n1216_lo <= 1'b0;
    n1228_lo <= 1'b0;
    n1231_lo <= 1'b0;
    n1237_lo <= 1'b0;
    n1240_lo <= 1'b0;
    n1243_lo <= 1'b0;
    n1249_lo <= 1'b0;
    n1252_lo <= 1'b0;
    n1255_lo <= 1'b0;
    n1261_lo <= 1'b0;
    n1264_lo <= 1'b0;
    n1267_lo <= 1'b0;
    n1273_lo <= 1'b0;
    n1276_lo <= 1'b0;
    n1279_lo <= 1'b0;
    n1282_lo <= 1'b0;
    n1285_lo <= 1'b0;
    n1288_lo <= 1'b0;
    n1291_lo <= 1'b0;
    n1294_lo <= 1'b0;
    n1297_lo <= 1'b0;
    n1300_lo <= 1'b0;
    n1303_lo <= 1'b0;
    n1309_lo <= 1'b0;
    n1312_lo <= 1'b0;
    n1315_lo <= 1'b0;
    n1318_lo <= 1'b0;
    n1321_lo <= 1'b0;
    n1324_lo <= 1'b0;
    n1333_lo <= 1'b0;
    n1874_o2 <= 1'b0;
    n2180_o2 <= 1'b0;
    n2372_o2 <= 1'b0;
    n2190_o2 <= 1'b0;
    n2191_o2 <= 1'b0;
    n2212_o2 <= 1'b0;
    n2213_o2 <= 1'b0;
    n2214_o2 <= 1'b0;
    n2215_o2 <= 1'b0;
    n2275_o2 <= 1'b0;
    n2276_o2 <= 1'b0;
    n2290_o2 <= 1'b0;
    n2291_o2 <= 1'b0;
    n2681_o2 <= 1'b0;
    n2680_o2 <= 1'b0;
    n2683_o2 <= 1'b0;
    n2684_o2 <= 1'b0;
    n2686_o2 <= 1'b0;
    n2319_o2 <= 1'b0;
    n2320_o2 <= 1'b0;
    n304_inv <= 1'b0;
    G554_o2 <= 1'b0;
    G557_o2 <= 1'b0;
    G185_o2 <= 1'b0;
    G188_o2 <= 1'b0;
    G191_o2 <= 1'b0;
    G194_o2 <= 1'b0;
    G1182_o2 <= 1'b0;
    G1222_o2 <= 1'b0;
    G1247_o2 <= 1'b0;
    G1371_o2 <= 1'b0;
    G1383_o2 <= 1'b0;
    G1386_o2 <= 1'b0;
    n2416_o2 <= 1'b0;
    n2428_o2 <= 1'b0;
    n2438_o2 <= 1'b0;
    n2439_o2 <= 1'b0;
    n2440_o2 <= 1'b0;
    n2444_o2 <= 1'b0;
    n2497_o2 <= 1'b0;
    n2498_o2 <= 1'b0;
    n2503_o2 <= 1'b0;
    n2505_o2 <= 1'b0;
    n2529_o2 <= 1'b0;
    n2562_o2 <= 1'b0;
    n2570_o2 <= 1'b0;
    n2571_o2 <= 1'b0;
    n2574_o2 <= 1'b0;
    n2575_o2 <= 1'b0;
    G546_o2 <= 1'b0;
    G550_o2 <= 1'b0;
    n2633_o2 <= 1'b0;
    n2639_o2 <= 1'b0;
    n2642_o2 <= 1'b0;
    n2645_o2 <= 1'b0;
    n2679_o2 <= 1'b0;
    n2662_o2 <= 1'b0;
    n2724_o2 <= 1'b0;
    G382_o2 <= 1'b0;
    G199_o2 <= 1'b0;
    G202_o2 <= 1'b0;
    G225_o2 <= 1'b0;
    G248_o2 <= 1'b0;
    G260_o2 <= 1'b0;
    n2716_o2 <= 1'b0;
    n2737_o2 <= 1'b0;
    n1174_lo_buf_o2 <= 1'b0;
    n1198_lo_buf_o2 <= 1'b0;
    G371_o2 <= 1'b0;
    G1059_o2 <= 1'b0;
    n2586_o2 <= 1'b0;
    n2587_o2 <= 1'b0;
    n460_inv <= 1'b0;
    n2648_o2 <= 1'b0;
    n2649_o2 <= 1'b0;
    n2650_o2 <= 1'b0;
    n2651_o2 <= 1'b0;
    n2652_o2 <= 1'b0;
    G365_o2 <= 1'b0;
    G1496_o2 <= 1'b0;
    G1502_o2 <= 1'b0;
    n2700_o2 <= 1'b0;
    n2701_o2 <= 1'b0;
    n2733_o2 <= 1'b0;
    n2734_o2 <= 1'b0;
    n2744_o2 <= 1'b0;
    n2747_o2 <= 1'b0;
    n2754_o2 <= 1'b0;
    n2755_o2 <= 1'b0;
    n511_inv <= 1'b0;
    G1609_o2 <= 1'b0;
    G1625_o2 <= 1'b0;
    G738_o2 <= 1'b0;
    G755_o2 <= 1'b0;
    G1511_o2 <= 1'b0;
    G1522_o2 <= 1'b0;
    G1538_o2 <= 1'b0;
    G1549_o2 <= 1'b0;
    G1563_o2 <= 1'b0;
    G1584_o2 <= 1'b0;
    G1576_o2 <= 1'b0;
    G1598_o2 <= 1'b0;
    G1395_o2 <= 1'b0;
    G1410_o2 <= 1'b0;
    G1420_o2 <= 1'b0;
    G1434_o2 <= 1'b0;
    n562_inv <= 1'b0;
    n1162_lo_buf_o2 <= 1'b0;
    n1102_lo_buf_o2 <= 1'b0;
    G359_o2 <= 1'b0;
    n982_lo_buf_o2 <= 1'b0;
    n1030_lo_buf_o2 <= 1'b0;
    n1042_lo_buf_o2 <= 1'b0;
    n583_inv <= 1'b0;
    G606_o2 <= 1'b0;
    G1118_o2 <= 1'b0;
    G1069_o2 <= 1'b0;
    G1145_o2 <= 1'b0;
    G1209_o2 <= 1'b0;
    G1189_o2 <= 1'b0;
    G1699_o2 <= 1'b0;
    G1702_o2 <= 1'b0;
    G1705_o2 <= 1'b0;
    G1708_o2 <= 1'b0;
    G1684_o2 <= 1'b0;
    G1687_o2 <= 1'b0;
    G1690_o2 <= 1'b0;
    G1693_o2 <= 1'b0;
    G1696_o2 <= 1'b0;
    G1642_o2 <= 1'b0;
    G1645_o2 <= 1'b0;
    G1648_o2 <= 1'b0;
    G1651_o2 <= 1'b0;
    G1654_o2 <= 1'b0;
    G1657_o2 <= 1'b0;
    G1660_o2 <= 1'b0;
    n1222_lo_buf_o2 <= 1'b0;
    n1330_lo_buf_o2 <= 1'b0;
    n658_inv <= 1'b0;
    n661_inv <= 1'b0;
    n1306_lo_buf_o2 <= 1'b0;
    n1150_lo_buf_o2 <= 1'b0;
    G175_o2 <= 1'b0;
    G241_o2 <= 1'b0;
    G356_o2 <= 1'b0;
    G989_o2 <= 1'b0;
    G984_o2 <= 1'b0;
    n685_inv <= 1'b0;
    n688_inv <= 1'b0;
    n958_lo_buf_o2 <= 1'b0;
    n1114_lo_buf_o2 <= 1'b0;
    G182_o2 <= 1'b0;
    G1215_o2 <= 1'b0;
    G971_o2 <= 1'b0;
    G938_o2 <= 1'b0;
    G1198_o2 <= 1'b0;
    G1203_o2 <= 1'b0;
    G1218_o2 <= 1'b0;
    G785_o2 <= 1'b0;
    G1168_o2 <= 1'b0;
    G1130_o2 <= 1'b0;
    G1185_o2 <= 1'b0;
    G1250_o2 <= 1'b0;
    G1225_o2 <= 1'b0;
    G1791_o2 <= 1'b0;
    G1788_o2 <= 1'b0;
    G981_o2 <= 1'b0;
    n745_inv <= 1'b0;
    n748_inv <= 1'b0;
    G1062_o2 <= 1'b0;
    n970_lo_buf_o2 <= 1'b0;
    n1006_lo_buf_o2 <= 1'b0;
    n1078_lo_buf_o2 <= 1'b0;
    n1126_lo_buf_o2 <= 1'b0;
    n766_inv <= 1'b0;
    G165_o2 <= 1'b0;
    n1234_lo_buf_o2 <= 1'b0;
    n1246_lo_buf_o2 <= 1'b0;
    n1258_lo_buf_o2 <= 1'b0;
    n1270_lo_buf_o2 <= 1'b0;
    G368_o2 <= 1'b0;
    G428_o2 <= 1'b0;
    G212_o2 <= 1'b0;
    G841_o2 <= 1'b0;
    G788_o2 <= 1'b0;
    n1186_lo_buf_o2 <= 1'b0;
    G391_o2 <= 1'b0;
    G387_o2 <= 1'b0;
    G645_o2 <= 1'b0;
    G1140_o2 <= 1'b0;
    G1178_o2 <= 1'b0;
    G1370_o2 <= 1'b0;
    n820_inv <= 1'b0;
    G1357_o2 <= 1'b0;
    G816_o2 <= 1'b0;
    G1369_o2 <= 1'b0;
    G901_o2 <= 1'b0;
    G1056_o2 <= 1'b0;
    G1107_o2 <= 1'b0;
    G1087_o2 <= 1'b0;
    G1135_o2 <= 1'b0;
    n1018_lo_buf_o2 <= 1'b0;
    n1090_lo_buf_o2 <= 1'b0;
    n853_inv <= 1'b0;
    G131_o2 <= 1'b0;
    n859_inv <= 1'b0;
    n862_inv <= 1'b0;
    G338_o2 <= 1'b0;
    n1171_lo_buf_o2 <= 1'b0;
    n1195_lo_buf_o2 <= 1'b0;
    G419_o2 <= 1'b0;
    G425_o2 <= 1'b0;
    G497_o2 <= 1'b0;
    G416_o2 <= 1'b0;
    G491_o2 <= 1'b0;
    G500_o2 <= 1'b0;
    G353_o2 <= 1'b0;
    G641_o2 <= 1'b0;
    G1117_o2 <= 1'b0;
    G1096_o2 <= 1'b0;
    G1143_o2 <= 1'b0;
    G1112_o2 <= 1'b0;
    n1138_lo_buf_o2 <= 1'b0;
    n1210_lo_buf_o2 <= 1'b0;
    G687_o2 <= 1'b0;
    G541_o2 <= 1'b0;
    G802_o2 <= 1'b0;
    G813_o2 <= 1'b0;
    G810_o2 <= 1'b0;
    G987_o2 <= 1'b0;
    G898_o2 <= 1'b0;
    n946_lo_buf_o2 <= 1'b0;
    n1054_lo_buf_o2 <= 1'b0;
    G728_o2 <= 1'b0;
    G856_o2 <= 1'b0;
    n949_1_inv <= 1'b0;
    G942_o2 <= 1'b0;
    G1099_o2 <= 1'b0;
    G1154_o2 <= 1'b0;
    G1131_o2 <= 1'b0;
    G1169_o2 <= 1'b0;
    G134_o2 <= 1'b0;
    n970_inv <= 1'b0;
    G470_o2 <= 1'b0;
    G344_o2 <= 1'b0;
    G362_o2 <= 1'b0;
    G482_o2 <= 1'b0;
    G660_o2 <= 1'b0;
    G672_o2 <= 1'b0;
    n1096_lo_buf_o2 <= 1'b0;
    G479_o2 <= 1'b0;
    G669_o2 <= 1'b0;
    n994_lo_buf_o2 <= 1'b0;
    n1066_lo_buf_o2 <= 1'b0;
    n1006_inv <= 1'b0;
    G147_o2 <= 1'b0;
    G473_o2 <= 1'b0;
    G488_o2 <= 1'b0;
    G589_o2 <= 1'b0;
    G663_o2 <= 1'b0;
    G684_o2 <= 1'b0;
    G605_o2 <= 1'b0;
    G774_o2 <= 1'b0;
    G782_o2 <= 1'b0;
  end
endmodule


