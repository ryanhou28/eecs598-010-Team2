// Benchmark "c5315" written by ABC on Sun Oct 29 16:27:00 2023

module c5315_clk (  clk,
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58,
    G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70, G71, G72,
    G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86,
    G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G109, G110, G111, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G124,
    G125, G126, G127, G128, G129, G130, G131, G132, G133, G134, G135, G136,
    G137, G138, G139, G140, G141, G142, G143, G144, G145, G146, G147, G148,
    G149, G150, G151, G152, G153, G154, G155, G156, G157, G158, G159, G160,
    G161, G162, G163, G164, G165, G166, G167, G168, G169, G170, G171, G172,
    G173, G174, G175, G176, G177, G178,
    G5193, G5194, G5195, G5196, G5197, G5198, G5199, G5200, G5201, G5202,
    G5203, G5204, G5205, G5206, G5207, G5208, G5209, G5210, G5211, G5212,
    G5213, G5214, G5215, G5216, G5217, G5218, G5219, G5220, G5221, G5222,
    G5223, G5224, G5225, G5226, G5227, G5228, G5229, G5230, G5231, G5232,
    G5233, G5234, G5235, G5236, G5237, G5238, G5239, G5240, G5241, G5242,
    G5243, G5244, G5245, G5246, G5247, G5248, G5249, G5250, G5251, G5252,
    G5253, G5254, G5255, G5256, G5257, G5258, G5259, G5260, G5261, G5262,
    G5263, G5264, G5265, G5266, G5267, G5268, G5269, G5270, G5271, G5272,
    G5273, G5274, G5275, G5276, G5277, G5278, G5279, G5280, G5281, G5282,
    G5283, G5284, G5285, G5286, G5287, G5288, G5289, G5290, G5291, G5292,
    G5293, G5294, G5295, G5296, G5297, G5298, G5299, G5300, G5301, G5302,
    G5303, G5304, G5305, G5306, G5307, G5308, G5309, G5310, G5311, G5312,
    G5313, G5314, G5315  );
  
  input clk, G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70,
    G71, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98,
    G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G110,
    G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G133, G134,
    G135, G136, G137, G138, G139, G140, G141, G142, G143, G144, G145, G146,
    G147, G148, G149, G150, G151, G152, G153, G154, G155, G156, G157, G158,
    G159, G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G170,
    G171, G172, G173, G174, G175, G176, G177, G178;
  output G5193, G5194, G5195, G5196, G5197, G5198, G5199, G5200, G5201, G5202,
    G5203, G5204, G5205, G5206, G5207, G5208, G5209, G5210, G5211, G5212,
    G5213, G5214, G5215, G5216, G5217, G5218, G5219, G5220, G5221, G5222,
    G5223, G5224, G5225, G5226, G5227, G5228, G5229, G5230, G5231, G5232,
    G5233, G5234, G5235, G5236, G5237, G5238, G5239, G5240, G5241, G5242,
    G5243, G5244, G5245, G5246, G5247, G5248, G5249, G5250, G5251, G5252,
    G5253, G5254, G5255, G5256, G5257, G5258, G5259, G5260, G5261, G5262,
    G5263, G5264, G5265, G5266, G5267, G5268, G5269, G5270, G5271, G5272,
    G5273, G5274, G5275, G5276, G5277, G5278, G5279, G5280, G5281, G5282,
    G5283, G5284, G5285, G5286, G5287, G5288, G5289, G5290, G5291, G5292,
    G5293, G5294, G5295, G5296, G5297, G5298, G5299, G5300, G5301, G5302,
    G5303, G5304, G5305, G5306, G5307, G5308, G5309, G5310, G5311, G5312,
    G5313, G5314, G5315;
  reg n2610_lo, n2613_lo, n2616_lo, n2619_lo, n2622_lo, n2625_lo, n2628_lo,
    n2631_lo, n2634_lo, n2637_lo, n2640_lo, n2643_lo, n2646_lo, n2649_lo,
    n2652_lo, n2655_lo, n2658_lo, n2661_lo, n2664_lo, n2667_lo, n2670_lo,
    n2673_lo, n2676_lo, n2679_lo, n2682_lo, n2685_lo, n2688_lo, n2691_lo,
    n2694_lo, n2697_lo, n2700_lo, n2703_lo, n2706_lo, n2709_lo, n2712_lo,
    n2715_lo, n2718_lo, n2721_lo, n2724_lo, n2727_lo, n2730_lo, n2733_lo,
    n2736_lo, n2739_lo, n2742_lo, n2745_lo, n2748_lo, n2751_lo, n2754_lo,
    n2757_lo, n2760_lo, n2763_lo, n2766_lo, n2769_lo, n2772_lo, n2775_lo,
    n2778_lo, n2781_lo, n2784_lo, n2787_lo, n2790_lo, n2793_lo, n2796_lo,
    n2799_lo, n2802_lo, n2805_lo, n2808_lo, n2811_lo, n2814_lo, n2817_lo,
    n2820_lo, n2823_lo, n2826_lo, n2829_lo, n2832_lo, n2835_lo, n2838_lo,
    n2841_lo, n2844_lo, n2847_lo, n2850_lo, n2853_lo, n2856_lo, n2859_lo,
    n2862_lo, n2865_lo, n2868_lo, n2871_lo, n2874_lo, n2877_lo, n2880_lo,
    n2883_lo, n2886_lo, n2889_lo, n2892_lo, n2895_lo, n2898_lo, n2901_lo,
    n2904_lo, n2907_lo, n2910_lo, n2913_lo, n2916_lo, n2919_lo, n2922_lo,
    n2925_lo, n2928_lo, n2931_lo, n2934_lo, n2937_lo, n2940_lo, n2943_lo,
    n2946_lo, n2949_lo, n2952_lo, n2955_lo, n2958_lo, n2961_lo, n2964_lo,
    n2967_lo, n2970_lo, n2973_lo, n2976_lo, n2979_lo, n2982_lo, n2985_lo,
    n2988_lo, n2991_lo, n2994_lo, n2997_lo, n3000_lo, n3003_lo, n3006_lo,
    n3009_lo, n3012_lo, n3015_lo, n3018_lo, n3021_lo, n3024_lo, n3027_lo,
    n3030_lo, n3033_lo, n3036_lo, n3039_lo, n3042_lo, n3045_lo, n3048_lo,
    n3051_lo, n3054_lo, n3057_lo, n3060_lo, n3063_lo, n3066_lo, n3069_lo,
    n3072_lo, n3075_lo, n3078_lo, n3081_lo, n3084_lo, n3087_lo, n3090_lo,
    n3093_lo, n3096_lo, n3099_lo, n3102_lo, n3105_lo, n3108_lo, n3111_lo,
    n3114_lo, n3117_lo, n3120_lo, n3123_lo, n3126_lo, n3129_lo, n3132_lo,
    n3135_lo, n3138_lo, n3141_lo, n3144_lo, n3147_lo, n3150_lo, n3153_lo,
    n3156_lo, n3159_lo, n3162_lo, n3165_lo, n3168_lo, n3171_lo, n3174_lo,
    n3177_lo, n3180_lo, n3183_lo, n3186_lo, n3189_lo, n3192_lo, n3195_lo,
    n3198_lo, n3201_lo, n3204_lo, n3207_lo, n3210_lo, n3213_lo, n3216_lo,
    n3219_lo, n3222_lo, n3225_lo, n3228_lo, n3231_lo, n3234_lo, n3237_lo,
    n3240_lo, n3243_lo, n3246_lo, n3249_lo, n3252_lo, n3255_lo, n3258_lo,
    n3261_lo, n3264_lo, n3267_lo, n3270_lo, n3273_lo, n3276_lo, n3279_lo,
    n3282_lo, n3285_lo, n3288_lo, n3291_lo, n3294_lo, n3297_lo, n3300_lo,
    n3303_lo, n3306_lo, n3309_lo, n3312_lo, n3315_lo, n3318_lo, n3321_lo,
    n3324_lo, n3327_lo, n3330_lo, n3333_lo, n3336_lo, n3339_lo, n3342_lo,
    n3345_lo, n3348_lo, n3351_lo, n3354_lo, n3357_lo, n3360_lo, n3363_lo,
    n3366_lo, n3369_lo, n3372_lo, n3375_lo, n3378_lo, n3381_lo, n3384_lo,
    n3387_lo, n3390_lo, n3393_lo, n3396_lo, n3399_lo, n3402_lo, n3405_lo,
    n3408_lo, n3411_lo, n3414_lo, n3417_lo, n3420_lo, n3423_lo, n3426_lo,
    n3429_lo, n3432_lo, n3435_lo, n3438_lo, n3441_lo, n3444_lo, n3447_lo,
    n3450_lo, n3453_lo, n3456_lo, n3459_lo, n3462_lo, n3465_lo, n3468_lo,
    n3471_lo, n3474_lo, n3477_lo, n3480_lo, n3483_lo, n3486_lo, n3489_lo,
    n3492_lo, n3495_lo, n3498_lo, n3501_lo, n3504_lo, n3507_lo, n3510_lo,
    n3513_lo, n3516_lo, n3519_lo, n3522_lo, n3525_lo, n3528_lo, n3531_lo,
    n3534_lo, n3537_lo, n3540_lo, n3543_lo, n3546_lo, n3549_lo, n3552_lo,
    n3555_lo, n3558_lo, n3561_lo, n3564_lo, n3567_lo, n3570_lo, n3573_lo,
    n3576_lo, n3579_lo, n3582_lo, n3585_lo, n3588_lo, n3591_lo, n3594_lo,
    n3597_lo, n3600_lo, n3603_lo, n3606_lo, n3609_lo, n3612_lo, n3615_lo,
    n3618_lo, n3621_lo, n3624_lo, n3627_lo, n3630_lo, n3633_lo, n3636_lo,
    n3639_lo, n3642_lo, n3645_lo, n3648_lo, n3651_lo, n3654_lo, n3657_lo,
    n3660_lo, n3663_lo, n3666_lo, n3669_lo, n3672_lo, n3675_lo, n3678_lo,
    n3681_lo, n3684_lo, n3687_lo, n3690_lo, n3693_lo, n3696_lo, n3699_lo,
    n3702_lo, n3705_lo, n3708_lo, n3711_lo, n3714_lo, n3717_lo, n3720_lo,
    n3723_lo, n3726_lo, n3729_lo, n3732_lo, n3735_lo, n3738_lo, n3741_lo,
    n3744_lo, n3747_lo, n3750_lo, n3753_lo, n3756_lo, n3759_lo, n3762_lo,
    n3765_lo, n3768_lo, n3771_lo, n3774_lo, n3777_lo, n3780_lo, n3783_lo,
    n3786_lo, n3789_lo, n3792_lo, n3795_lo, n3798_lo, n3801_lo, n3804_lo,
    n3807_lo, n3810_lo, n3813_lo, n3816_lo, n3819_lo, n3822_lo, n3825_lo,
    n3828_lo, n3831_lo, n3834_lo, n3837_lo, n3840_lo, n3843_lo, n3846_lo,
    n3849_lo, n3852_lo, n3855_lo, n3858_lo, n3861_lo, n3864_lo, n3867_lo,
    n3870_lo, n3873_lo, n3876_lo, n3879_lo, n3882_lo, n3885_lo, n3888_lo,
    n3891_lo, n3894_lo, n3897_lo, n3900_lo, n3903_lo, n3906_lo, n3909_lo,
    n3912_lo, n3915_lo, n3918_lo, n3921_lo, n3924_lo, n3927_lo, n3930_lo,
    n3933_lo, n3936_lo, n3939_lo, n3942_lo, n3945_lo, n3948_lo, n3951_lo,
    n3954_lo, n3957_lo, n3960_lo, n3963_lo, n3966_lo, n3969_lo, n3972_lo,
    n3975_lo, n3978_lo, n3981_lo, n3984_lo, n3987_lo, n3990_lo, n3993_lo,
    n3996_lo, n3999_lo, n4002_lo, n4005_lo, n4008_lo, n4011_lo, n4014_lo,
    n4017_lo, n4020_lo, n4023_lo, n4026_lo, n4029_lo, n4032_lo, n4035_lo,
    n4038_lo, n4041_lo, n4044_lo, n4047_lo, n4050_lo, n4053_lo, n4056_lo,
    n4059_lo, n4062_lo, n4065_lo, n4068_lo, n4071_lo, n4074_lo, n4077_lo,
    n4080_lo, n4083_lo, n4086_lo, n4089_lo, n4092_lo, n4095_lo, n4098_lo,
    n4101_lo, n4104_lo, n4107_lo, n4110_lo, n4113_lo, n4116_lo, n4119_lo,
    n4122_lo, n4125_lo, n4128_lo, n4131_lo, n4134_lo, n4137_lo, n4140_lo,
    n4143_lo, n4146_lo, n4149_lo, n4152_lo, n4155_lo, n4158_lo, n4161_lo,
    n4164_lo, n4167_lo, n4170_lo, n4173_lo, n4176_lo, n4179_lo, n4182_lo,
    n4185_lo, n4188_lo, n4191_lo, n4194_lo, n4197_lo, n4200_lo, n4203_lo,
    n4206_lo, n4209_lo, n4212_lo, n4215_lo, n4218_lo, n4221_lo, n4224_lo,
    n4227_lo, n4230_lo, n4233_lo, n4236_lo, n4239_lo, n4242_lo, n4245_lo,
    n4248_lo, n4251_lo, n4254_lo, n4257_lo, n4260_lo, n4263_lo, n4266_lo,
    n4269_lo, n4272_lo, n4275_lo, n4278_lo, n4281_lo, n4284_lo, n4287_lo,
    n4290_lo, n4293_lo, n4296_lo, n4299_lo, n4302_lo, n4305_lo, n4308_lo,
    n4311_lo, n4314_lo, n4317_lo, n4320_lo, n4323_lo, n4326_lo, n4329_lo,
    n4332_lo, n4335_lo, n4338_lo, n4341_lo, n4344_lo, n4347_lo, n4350_lo,
    n4353_lo, n4356_lo, n4359_lo, n4362_lo, n4365_lo, n4368_lo, n4371_lo,
    n4374_lo, n4377_lo, n4380_lo, n4383_lo, n4386_lo, n4389_lo, n4392_lo,
    n4395_lo, n4398_lo, n4401_lo, n4404_lo, n4407_lo, n4410_lo, n4413_lo,
    n4416_lo, n4419_lo, n4422_lo, n4425_lo, n4428_lo, n4431_lo, n4434_lo,
    n4437_lo, n4440_lo, n4443_lo, n4446_lo, n4449_lo, n4452_lo, n4455_lo,
    n4458_lo, n4461_lo, n4464_lo, n4467_lo, n4470_lo, n4473_lo, n4476_lo,
    n4479_lo, n4482_lo, n4485_lo, n4488_lo, n4491_lo, n4494_lo, n4497_lo,
    n4500_lo, n4503_lo, n4506_lo, n4509_lo, n4512_lo, n4515_lo, n4518_lo,
    n4521_lo, n4524_lo, n4527_lo, n4530_lo, n4533_lo, n4536_lo, n4539_lo,
    n4542_lo, n4545_lo, n4548_lo, n4551_lo, n4554_lo, n4557_lo, n4560_lo,
    n4563_lo, n4566_lo, n4569_lo, n4572_lo, n4575_lo, n4578_lo, n4581_lo,
    n4584_lo, n4587_lo, n4590_lo, n4593_lo, n4596_lo, n4599_lo, n4602_lo,
    n4605_lo, n4608_lo, n4611_lo, n4614_lo, n4617_lo, n4620_lo, n4623_lo,
    n4626_lo, n4629_lo, n4632_lo, n4635_lo, n4638_lo, n4641_lo, n4644_lo,
    n4647_lo, n4650_lo, n4653_lo, n4656_lo, n4659_lo, n4662_lo, n4665_lo,
    n4668_lo, n4671_lo, n4674_lo, n4677_lo, n4680_lo, n4683_lo, n4686_lo,
    n4689_lo, n4692_lo, n4695_lo, n4698_lo, n4701_lo, n4704_lo, n4707_lo,
    n4710_lo, n4713_lo, n4716_lo, n4719_lo, n4722_lo, n4725_lo, n4728_lo,
    n4731_lo, n4734_lo, n4737_lo, n4740_lo, n4743_lo;
  wire new_G632_, new_G633_, new_G634_, new_G647_, new_G659_, new_G671_,
    new_G684_, new_G685_, new_G686_, new_G687_, new_G688_, new_G689_,
    new_G690_, new_G694_, new_G706_, new_G718_, new_G730_, new_G742_,
    new_G746_, new_G749_, new_G752_, new_G756_, new_G768_, new_G780_,
    new_G792_, new_G804_, new_G813_, new_G825_, new_G836_, new_G848_,
    new_G860_, new_G872_, new_G884_, new_G896_, new_G908_, new_G911_,
    new_G914_, new_G917_, new_G920_, new_G923_, new_G926_, new_G929_,
    new_G932_, new_G935_, new_G938_, new_G941_, new_G944_, new_G947_,
    new_G950_, new_G953_, new_G956_, new_G963_, new_G970_, new_G976_,
    new_G980_, new_G983_, new_G993_, new_G996_, new_G999_, new_G1002_,
    new_G1005_, new_G1008_, new_G1011_, new_G1014_, new_G1017_, new_G1020_,
    new_G1023_, new_G1026_, new_G1029_, new_G1032_, new_G1035_, new_G1038_,
    new_G1041_, new_G1044_, new_G1047_, new_G1050_, new_G1053_, new_G1060_,
    new_G1067_, new_G1070_, new_G1075_, new_G1081_, new_G1084_, new_G1087_,
    new_G1090_, new_G1093_, new_G1096_, new_G1099_, new_G1102_, new_G1105_,
    new_G1108_, new_G1111_, new_G1114_, new_G1117_, new_G1120_, new_G1123_,
    new_G1126_, new_G1129_, new_G1132_, new_G1135_, new_G1138_, new_G1141_,
    new_G1144_, new_G1147_, new_G1150_, new_G1162_, new_G1172_, new_G1184_,
    new_G1196_, new_G1208_, new_G1214_, new_G1218_, new_G1230_, new_G1242_,
    new_G1245_, new_G1248_, new_G1256_, new_G1264_, new_G1272_, new_G1280_,
    new_G1287_, new_G1294_, new_G1301_, new_G1308_, new_G1311_, new_G1314_,
    new_G1317_, new_G1320_, new_G1323_, new_G1326_, new_G1329_, new_G1332_,
    new_G1335_, new_G1338_, new_G1341_, new_G1344_, new_G1347_, new_G1350_,
    new_G1353_, new_G1356_, new_G1359_, new_G1362_, new_G1365_, new_G1368_,
    new_G1371_, new_G1374_, new_G1377_, new_G1380_, new_G1383_, new_G1386_,
    new_G1389_, new_G1392_, new_G1395_, new_G1398_, new_G1401_, new_G1404_,
    new_G1407_, new_G1410_, new_G1413_, new_G1416_, new_G1419_, new_G1422_,
    new_G1425_, new_G1428_, new_G1431_, new_G1434_, new_G1437_, new_G1440_,
    new_G1443_, new_G1446_, new_G1449_, new_G1452_, new_G1455_, new_G1458_,
    new_G1459_, new_G1460_, new_G1461_, new_G1462_, new_G1463_, new_G1464_,
    new_G1465_, new_G1466_, new_G1467_, new_G1468_, new_G1469_, new_G1470_,
    new_G1471_, new_G1472_, new_G1473_, new_G1474_, new_G1475_, new_G1476_,
    new_G1477_, new_G1478_, new_G1479_, new_G1480_, new_G1481_, new_G1482_,
    new_G1483_, new_G1484_, new_G1485_, new_G1486_, new_G1487_, new_G1488_,
    new_G1489_, new_G1490_, new_G1491_, new_G1492_, new_G1493_, new_G1494_,
    new_G1495_, new_G1496_, new_G1497_, new_G1498_, new_G1499_, new_G1500_,
    new_G1501_, new_G1502_, new_G1503_, new_G1504_, new_G1505_, new_G1506_,
    new_G1507_, new_G1508_, new_G1509_, new_G1510_, new_G1511_, new_G1512_,
    new_G1513_, new_G1514_, new_G1515_, new_G1516_, new_G1517_, new_G1518_,
    new_G1519_, new_G1520_, new_G1526_, new_G1537_, new_G1548_, new_G1554_,
    new_G1565_, new_G1576_, new_G1577_, new_G1582_, new_G1583_, new_G1584_,
    new_G1585_, new_G1586_, new_G1587_, new_G1588_, new_G1589_, new_G1590_,
    new_G1591_, new_G1592_, new_G1593_, new_G1594_, new_G1595_, new_G1601_,
    new_G1612_, new_G1623_, new_G1629_, new_G1640_, new_G1651_, new_G1652_,
    new_G1663_, new_G1674_, new_G1685_, new_G1696_, new_G1697_, new_G1698_,
    new_G1699_, new_G1700_, new_G1701_, new_G1702_, new_G1703_, new_G1704_,
    new_G1705_, new_G1706_, new_G1707_, new_G1708_, new_G1709_, new_G1710_,
    new_G1711_, new_G1712_, new_G1713_, new_G1714_, new_G1715_, new_G1716_,
    new_G1717_, new_G1718_, new_G1719_, new_G1720_, new_G1721_, new_G1722_,
    new_G1723_, new_G1724_, new_G1725_, new_G1726_, new_G1727_, new_G1728_,
    new_G1734_, new_G1740_, new_G1741_, new_G1742_, new_G1743_, new_G1744_,
    new_G1745_, new_G1746_, new_G1747_, new_G1748_, new_G1749_, new_G1750_,
    new_G1755_, new_G1764_, new_G1774_, new_G1775_, new_G1776_, new_G1777_,
    new_G1778_, new_G1779_, new_G1780_, new_G1781_, new_G1782_, new_G1783_,
    new_G1784_, new_G1785_, new_G1786_, new_G1787_, new_G1788_, new_G1789_,
    new_G1790_, new_G1791_, new_G1792_, new_G1793_, new_G1794_, new_G1795_,
    new_G1796_, new_G1797_, new_G1798_, new_G1799_, new_G1800_, new_G1801_,
    new_G1802_, new_G1803_, new_G1804_, new_G1805_, new_G1806_, new_G1807_,
    new_G1808_, new_G1809_, new_G1810_, new_G1811_, new_G1812_, new_G1813_,
    new_G1814_, new_G1815_, new_G1821_, new_G1827_, new_G1828_, new_G1829_,
    new_G1830_, new_G1831_, new_G1832_, new_G1833_, new_G1834_, new_G1835_,
    new_G1836_, new_G1837_, new_G1842_, new_G1843_, new_G1844_, new_G1845_,
    new_G1846_, new_G1847_, new_G1848_, new_G1849_, new_G1850_, new_G1851_,
    new_G1852_, new_G1853_, new_G1854_, new_G1855_, new_G1856_, new_G1857_,
    new_G1858_, new_G1859_, new_G1860_, new_G1861_, new_G1862_, new_G1863_,
    new_G1864_, new_G1865_, new_G1866_, new_G1867_, new_G1868_, new_G1869_,
    new_G1870_, new_G1871_, new_G1872_, new_G1873_, new_G1876_, new_G1879_,
    new_G1880_, new_G1883_, new_G1886_, new_G1887_, new_G1888_, new_G1889_,
    new_G1890_, new_G1891_, new_G1892_, new_G1893_, new_G1894_, new_G1895_,
    new_G1896_, new_G1897_, new_G1898_, new_G1899_, new_G1900_, new_G1901_,
    new_G1902_, new_G1903_, new_G1904_, new_G1905_, new_G1906_, new_G1907_,
    new_G1908_, new_G1911_, new_G1914_, new_G1925_, new_G1936_, new_G1941_,
    new_G1944_, new_G1945_, new_G1946_, new_G1947_, new_G1948_, new_G1959_,
    new_G1970_, new_G1981_, new_G1992_, new_G2003_, new_G2014_, new_G2015_,
    new_G2016_, new_G2017_, new_G2018_, new_G2019_, new_G2020_, new_G2031_,
    new_G2042_, new_G2053_, new_G2064_, new_G2067_, new_G2068_, new_G2069_,
    new_G2070_, new_G2071_, new_G2072_, new_G2073_, new_G2076_, new_G2077_,
    new_G2078_, new_G2079_, new_G2080_, new_G2081_, new_G2082_, new_G2083_,
    new_G2084_, new_G2085_, new_G2086_, new_G2087_, new_G2088_, new_G2089_,
    new_G2090_, new_G2091_, new_G2092_, new_G2093_, new_G2094_, new_G2095_,
    new_G2096_, new_G2097_, new_G2098_, new_G2099_, new_G2100_, new_G2101_,
    new_G2102_, new_G2103_, new_G2104_, new_G2105_, new_G2108_, new_G2109_,
    new_G2110_, new_G2111_, new_G2112_, new_G2113_, new_G2114_, new_G2115_,
    new_G2116_, new_G2117_, new_G2118_, new_G2119_, new_G2120_, new_G2121_,
    new_G2122_, new_G2123_, new_G2124_, new_G2125_, new_G2126_, new_G2127_,
    new_G2128_, new_G2129_, new_G2130_, new_G2131_, new_G2132_, new_G2133_,
    new_G2134_, new_G2135_, new_G2136_, new_G2137_, new_G2138_, new_G2139_,
    new_G2140_, new_G2141_, new_G2142_, new_G2143_, new_G2144_, new_G2145_,
    new_G2146_, new_G2147_, new_G2148_, new_G2149_, new_G2150_, new_G2151_,
    new_G2152_, new_G2153_, new_G2154_, new_G2155_, new_G2156_, new_G2157_,
    new_G2158_, new_G2159_, new_G2160_, new_G2161_, new_G2162_, new_G2163_,
    new_G2164_, new_G2165_, new_G2166_, new_G2167_, new_G2168_, new_G2169_,
    new_G2170_, new_G2171_, new_G2172_, new_G2173_, new_G2174_, new_G2175_,
    new_G2176_, new_G2177_, new_G2178_, new_G2179_, new_G2180_, new_G2181_,
    new_G2182_, new_G2183_, new_G2184_, new_G2185_, new_G2186_, new_G2187_,
    new_G2188_, new_G2189_, new_G2190_, new_G2191_, new_G2192_, new_G2193_,
    new_G2194_, new_G2195_, new_G2196_, new_G2197_, new_G2198_, new_G2199_,
    new_G2200_, new_G2201_, new_G2202_, new_G2203_, new_G2204_, new_G2205_,
    new_G2206_, new_G2207_, new_G2208_, new_G2209_, new_G2210_, new_G2211_,
    new_G2212_, new_G2213_, new_G2214_, new_G2215_, new_G2216_, new_G2217_,
    new_G2218_, new_G2219_, new_G2220_, new_G2221_, new_G2222_, new_G2223_,
    new_G2224_, new_G2225_, new_G2226_, new_G2227_, new_G2228_, new_G2229_,
    new_G2230_, new_G2231_, new_G2240_, new_G2241_, new_G2242_, new_G2243_,
    new_G2244_, new_G2245_, new_G2248_, new_G2249_, new_G2250_, new_G2251_,
    new_G2252_, new_G2253_, new_G2254_, new_G2255_, new_G2256_, new_G2257_,
    new_G2258_, new_G2259_, new_G2260_, new_G2261_, new_G2262_, new_G2263_,
    new_G2264_, new_G2265_, new_G2266_, new_G2267_, new_G2268_, new_G2269_,
    new_G2270_, new_G2271_, new_G2277_, new_G2278_, new_G2279_, new_G2280_,
    new_G2281_, new_G2282_, new_G2283_, new_G2284_, new_G2285_, new_G2286_,
    new_G2287_, new_G2288_, new_G2289_, new_G2290_, new_G2291_, new_G2292_,
    new_G2293_, new_G2294_, new_G2295_, new_G2296_, new_G2297_, new_G2298_,
    new_G2299_, new_G2300_, new_G2301_, new_G2302_, new_G2303_, new_G2304_,
    new_G2305_, new_G2306_, new_G2307_, new_G2308_, new_G2309_, new_G2310_,
    new_G2314_, new_G2318_, new_G2319_, new_G2320_, new_G2321_, new_G2322_,
    new_G2323_, new_G2324_, new_G2325_, new_G2326_, new_G2327_, new_G2328_,
    new_G2332_, new_G2336_, new_G2339_, new_G2340_, new_G2341_, new_G2342_,
    new_G2343_, new_G2344_, new_G2345_, new_G2346_, new_G2347_, new_G2348_,
    new_G2349_, new_G2352_, new_G2355_, new_G2358_, new_G2361_, new_G2362_,
    new_G2363_, new_G2366_, new_G2367_, new_G2368_, new_G2369_, new_G2370_,
    new_G2371_, new_G2372_, new_G2373_, new_G2374_, new_G2375_, new_G2376_,
    new_G2377_, new_G2378_, new_G2379_, new_G2386_, new_G2392_, new_G2398_,
    new_G2404_, new_G2410_, new_G2418_, new_G2424_, new_G2430_, new_G2436_,
    new_G2437_, new_G2438_, new_G2441_, new_G2442_, new_G2443_, new_G2444_,
    new_G2445_, new_G2446_, new_G2447_, new_G2448_, new_G2454_, new_G2460_,
    new_G2466_, new_G2472_, new_G2480_, new_G2486_, new_G2492_, new_G2499_,
    new_G2500_, new_G2501_, new_G2502_, new_G2503_, new_G2504_, new_G2505_,
    new_G2506_, new_G2507_, new_G2508_, new_G2511_, new_G2512_, new_G2513_,
    new_G2514_, new_G2515_, new_G2516_, new_G2517_, new_G2520_, new_G2523_,
    new_G2526_, new_G2527_, new_G2528_, new_G2529_, new_G2530_, new_G2531_,
    new_G2532_, new_G2533_, new_G2534_, new_G2535_, new_G2536_, new_G2537_,
    new_G2538_, new_G2539_, new_G2540_, new_G2543_, new_G2547_, new_G2550_,
    new_G2553_, new_G2556_, new_G2559_, new_G2562_, new_G2565_, new_G2568_,
    new_G2571_, new_G2574_, new_G2577_, new_G2580_, new_G2583_, new_G2586_,
    new_G2589_, new_G2590_, new_G2591_, new_G2592_, new_G2593_, new_G2596_,
    new_G2599_, new_G2600_, new_G2601_, new_G2602_, new_G2603_, new_G2606_,
    new_G2609_, new_G2612_, new_G2615_, new_G2618_, new_G2621_, new_G2624_,
    new_G2625_, new_G2626_, new_G2629_, new_G2632_, new_G2635_, new_G2638_,
    new_G2641_, new_G2644_, new_G2647_, new_G2650_, new_G2653_, new_G2656_,
    new_G2659_, new_G2662_, new_G2663_, new_G2666_, new_G2667_, new_G2668_,
    new_G2669_, new_G2670_, new_G2671_, new_G2672_, new_G2673_, new_G2674_,
    new_G2675_, new_G2679_, new_G2685_, new_G2692_, new_G2693_, new_G2696_,
    new_G2700_, new_G2705_, new_G2711_, new_G2715_, new_G2720_, new_G2726_,
    new_G2727_, new_G2731_, new_G2737_, new_G2744_, new_G2752_, new_G2759_,
    new_G2770_, new_G2774_, new_G2780_, new_G2787_, new_G2788_, new_G2792_,
    new_G2797_, new_G2804_, new_G2810_, new_G2817_, new_G2828_, new_G2832_,
    new_G2837_, new_G2843_, new_G2844_, new_G2850_, new_G2857_, new_G2865_,
    new_G2872_, new_G2875_, new_G2876_, new_G2877_, new_G2878_, new_G2879_,
    new_G2883_, new_G2887_, new_G2888_, new_G2891_, new_G2894_, new_G2897_,
    new_G2900_, new_G2903_, new_G2906_, new_G2909_, new_G2912_, new_G2915_,
    new_G2918_, new_G2921_, new_G2924_, new_G2927_, new_G2930_, new_G2933_,
    new_G2936_, new_G2939_, new_G2942_, new_G2945_, new_G2948_, new_G2951_,
    new_G2954_, new_G2957_, new_G2960_, new_G2963_, new_G2966_, new_G2969_,
    new_G2972_, new_G2975_, new_G2978_, new_G2981_, new_G2984_, new_G2987_,
    new_G2990_, new_G2993_, new_G2996_, new_G2999_, new_G3002_, new_G3005_,
    new_G3008_, new_G3011_, new_G3014_, new_G3017_, new_G3020_, new_G3023_,
    new_G3026_, new_G3029_, new_G3032_, new_G3035_, new_G3038_, new_G3039_,
    new_G3040_, new_G3041_, new_G3042_, new_G3043_, new_G3044_, new_G3045_,
    new_G3046_, new_G3047_, new_G3048_, new_G3049_, new_G3050_, new_G3051_,
    new_G3052_, new_G3053_, new_G3054_, new_G3055_, new_G3056_, new_G3057_,
    new_G3058_, new_G3059_, new_G3060_, new_G3063_, new_G3064_, new_G3065_,
    new_G3066_, new_G3067_, new_G3068_, new_G3069_, new_G3070_, new_G3071_,
    new_G3072_, new_G3073_, new_G3074_, new_G3075_, new_G3076_, new_G3077_,
    new_G3078_, new_G3079_, new_G3080_, new_G3081_, new_G3082_, new_G3083_,
    new_G3084_, new_G3085_, new_G3086_, new_G3087_, new_G3088_, new_G3089_,
    new_G3090_, new_G3091_, new_G3092_, new_G3093_, new_G3094_, new_G3097_,
    new_G3098_, new_G3099_, new_G3100_, new_G3101_, new_G3102_, new_G3103_,
    new_G3104_, new_G3105_, new_G3106_, new_G3107_, new_G3108_, new_G3109_,
    new_G3110_, new_G3111_, new_G3112_, new_G3113_, new_G3114_, new_G3115_,
    new_G3116_, new_G3117_, new_G3118_, new_G3119_, new_G3120_, new_G3121_,
    new_G3122_, new_G3123_, new_G3124_, new_G3125_, new_G3126_, new_G3127_,
    new_G3128_, new_G3129_, new_G3130_, new_G3131_, new_G3132_, new_G3133_,
    new_G3134_, new_G3135_, new_G3136_, new_G3137_, new_G3138_, new_G3139_,
    new_G3140_, new_G3141_, new_G3142_, new_G3143_, new_G3144_, new_G3145_,
    new_G3146_, new_G3147_, new_G3148_, new_G3149_, new_G3150_, new_G3151_,
    new_G3152_, new_G3153_, new_G3154_, new_G3155_, new_G3156_, new_G3157_,
    new_G3158_, new_G3159_, new_G3160_, new_G3161_, new_G3162_, new_G3163_,
    new_G3164_, new_G3165_, new_G3166_, new_G3167_, new_G3168_, new_G3169_,
    new_G3170_, new_G3171_, new_G3172_, new_G3173_, new_G3174_, new_G3175_,
    new_G3176_, new_G3177_, new_G3178_, new_G3179_, new_G3180_, new_G3181_,
    new_G3182_, new_G3183_, new_G3184_, new_G3185_, new_G3186_, new_G3187_,
    new_G3188_, new_G3189_, new_G3190_, new_G3191_, new_G3192_, new_G3195_,
    new_G3196_, new_G3197_, new_G3198_, new_G3199_, new_G3202_, new_G3203_,
    new_G3204_, new_G3205_, new_G3206_, new_G3207_, new_G3208_, new_G3211_,
    new_G3214_, new_G3215_, new_G3218_, new_G3219_, new_G3222_, new_G3225_,
    new_G3228_, new_G3231_, new_G3234_, new_G3237_, new_G3240_, new_G3241_,
    new_G3244_, new_G3247_, new_G3250_, new_G3253_, new_G3256_, new_G3259_,
    new_G3262_, new_G3265_, new_G3266_, new_G3267_, new_G3268_, new_G3269_,
    new_G3270_, new_G3271_, new_G3272_, new_G3273_, new_G3274_, new_G3275_,
    new_G3276_, new_G3277_, new_G3280_, new_G3281_, new_G3282_, new_G3283_,
    new_G3284_, new_G3285_, new_G3286_, new_G3287_, new_G3288_, new_G3289_,
    new_G3290_, new_G3291_, new_G3292_, new_G3293_, new_G3294_, new_G3295_,
    new_G3296_, new_G3297_, new_G3298_, new_G3299_, new_G3300_, new_G3301_,
    new_G3302_, new_G3303_, new_G3313_, new_G3314_, new_G3315_, new_G3316_,
    new_G3317_, new_G3331_, new_G3332_, new_G3333_, new_G3334_, new_G3335_,
    new_G3336_, new_G3337_, new_G3338_, new_G3339_, new_G3340_, new_G3341_,
    new_G3342_, new_G3343_, new_G3344_, new_G3348_, new_G3351_, new_G3355_,
    new_G3358_, new_G3359_, new_G3360_, new_G3363_, new_G3364_, new_G3365_,
    new_G3366_, new_G3367_, new_G3368_, new_G3369_, new_G3370_, new_G3371_,
    new_G3374_, new_G3377_, new_G3380_, new_G3383_, new_G3386_, new_G3393_,
    new_G3404_, new_G3415_, new_G3421_, new_G3428_, new_G3438_, new_G3449_,
    new_G3459_, new_G3466_, new_G3467_, new_G3474_, new_G3485_, new_G3495_,
    new_G3503_, new_G3517_, new_G3533_, new_G3546_, new_G3552_, new_G3559_,
    new_G3570_, new_G3576_, new_G3583_, new_G3594_, new_G3604_, new_G3605_,
    new_G3606_, new_G3607_, new_G3608_, new_G3609_, new_G3610_, new_G3611_,
    new_G3621_, new_G3629_, new_G3645_, new_G3658_, new_G3664_, new_G3665_,
    new_G3666_, new_G3670_, new_G3674_, new_G3677_, new_G3681_, new_G3685_,
    new_G3688_, new_G3689_, new_G3690_, new_G3691_, new_G3692_, new_G3693_,
    new_G3694_, new_G3695_, new_G3696_, new_G3697_, new_G3700_, new_G3703_,
    new_G3706_, new_G3709_, new_G3710_, new_G3713_, new_G3714_, new_G3715_,
    new_G3716_, new_G3717_, new_G3718_, new_G3719_, new_G3720_, new_G3723_,
    new_G3726_, new_G3729_, new_G3732_, new_G3735_, new_G3738_, new_G3739_,
    new_G3742_, new_G3745_, new_G3748_, new_G3751_, new_G3752_, new_G3753_,
    new_G3754_, new_G3755_, new_G3756_, new_G3757_, new_G3758_, new_G3759_,
    new_G3760_, new_G3761_, new_G3762_, new_G3763_, new_G3764_, new_G3765_,
    new_G3768_, new_G3769_, new_G3770_, new_G3771_, new_G3772_, new_G3773_,
    new_G3774_, new_G3775_, new_G3776_, new_G3779_, new_G3780_, new_G3781_,
    new_G3782_, new_G3783_, new_G3784_, new_G3785_, new_G3786_, new_G3787_,
    new_G3788_, new_G3789_, new_G3790_, new_G3791_, new_G3792_, new_G3793_,
    new_G3796_, new_G3797_, new_G3798_, new_G3799_, new_G3800_, new_G3801_,
    new_G3802_, new_G3805_, new_G3806_, new_G3807_, new_G3808_, new_G3809_,
    new_G3810_, new_G3811_, new_G3812_, new_G3813_, new_G3814_, new_G3815_,
    new_G3816_, new_G3817_, new_G3818_, new_G3819_, new_G3820_, new_G3821_,
    new_G3822_, new_G3823_, new_G3824_, new_G3825_, new_G3828_, new_G3829_,
    new_G3830_, new_G3831_, new_G3832_, new_G3833_, new_G3834_, new_G3837_,
    new_G3838_, new_G3839_, new_G3840_, new_G3841_, new_G3842_, new_G3843_,
    new_G3844_, new_G3845_, new_G3846_, new_G3847_, new_G3848_, new_G3849_,
    new_G3852_, new_G3855_, new_G3856_, new_G3857_, new_G3858_, new_G3859_,
    new_G3862_, new_G3863_, new_G3864_, new_G3865_, new_G3866_, new_G3867_,
    new_G3868_, new_G3869_, new_G3870_, new_G3871_, new_G3872_, new_G3873_,
    new_G3874_, new_G3875_, new_G3876_, new_G3877_, new_G3878_, new_G3879_,
    new_G3882_, new_G3885_, new_G3888_, new_G3891_, new_G3894_, new_G3897_,
    new_G3900_, new_G3903_, new_G3904_, new_G3905_, new_G3906_, new_G3909_,
    new_G3912_, new_G3915_, new_G3918_, new_G3921_, new_G3924_, new_G3927_,
    new_G3930_, new_G3933_, new_G3936_, new_G3939_, new_G3942_, new_G3945_,
    new_G3948_, new_G3951_, new_G3954_, new_G3957_, new_G3960_, new_G3963_,
    new_G3966_, new_G3969_, new_G3972_, new_G3975_, new_G3978_, new_G3981_,
    new_G3984_, new_G3987_, new_G3990_, new_G3993_, new_G3996_, new_G3999_,
    new_G4002_, new_G4005_, new_G4008_, new_G4011_, new_G4014_, new_G4017_,
    new_G4020_, new_G4023_, new_G4026_, new_G4029_, new_G4032_, new_G4035_,
    new_G4038_, new_G4039_, new_G4040_, new_G4041_, new_G4042_, new_G4043_,
    new_G4044_, new_G4045_, new_G4046_, new_G4047_, new_G4048_, new_G4051_,
    new_G4054_, new_G4058_, new_G4061_, new_G4064_, new_G4065_, new_G4068_,
    new_G4072_, new_G4075_, new_G4076_, new_G4077_, new_G4080_, new_G4081_,
    new_G4082_, new_G4083_, new_G4084_, new_G4085_, new_G4086_, new_G4087_,
    new_G4088_, new_G4089_, new_G4092_, new_G4095_, new_G4098_, new_G4101_,
    new_G4104_, new_G4107_, new_G4110_, new_G4113_, new_G4116_, new_G4119_,
    new_G4122_, new_G4125_, new_G4128_, new_G4131_, new_G4134_, new_G4137_,
    new_G4140_, new_G4143_, new_G4146_, new_G4149_, new_G4152_, new_G4155_,
    new_G4158_, new_G4161_, new_G4164_, new_G4167_, new_G4170_, new_G4173_,
    new_G4174_, new_G4175_, new_G4176_, new_G4177_, new_G4180_, new_G4183_,
    new_G4184_, new_G4185_, new_G4186_, new_G4187_, new_G4188_, new_G4189_,
    new_G4190_, new_G4191_, new_G4192_, new_G4193_, new_G4194_, new_G4195_,
    new_G4196_, new_G4197_, new_G4198_, new_G4199_, new_G4200_, new_G4201_,
    new_G4202_, new_G4203_, new_G4204_, new_G4205_, new_G4206_, new_G4207_,
    new_G4208_, new_G4209_, new_G4210_, new_G4211_, new_G4212_, new_G4213_,
    new_G4214_, new_G4215_, new_G4216_, new_G4217_, new_G4218_, new_G4219_,
    new_G4220_, new_G4221_, new_G4222_, new_G4223_, new_G4224_, new_G4225_,
    new_G4226_, new_G4227_, new_G4230_, new_G4231_, new_G4232_, new_G4233_,
    new_G4234_, new_G4235_, new_G4236_, new_G4237_, new_G4238_, new_G4239_,
    new_G4240_, new_G4241_, new_G4242_, new_G4243_, new_G4244_, new_G4245_,
    new_G4246_, new_G4247_, new_G4248_, new_G4249_, new_G4250_, new_G4251_,
    new_G4252_, new_G4253_, new_G4254_, new_G4257_, new_G4260_, new_G4261_,
    new_G4262_, new_G4263_, new_G4264_, new_G4265_, new_G4266_, new_G4267_,
    new_G4268_, new_G4269_, new_G4270_, new_G4271_, new_G4272_, new_G4273_,
    new_G4274_, new_G4275_, new_G4276_, new_G4282_, new_G4283_, new_G4284_,
    new_G4285_, new_G4286_, new_G4287_, new_G4288_, new_G4289_, new_G4290_,
    new_G4293_, new_G4294_, new_G4295_, new_G4296_, new_G4297_, new_G4298_,
    new_G4299_, new_G4300_, new_G4301_, new_G4302_, new_G4303_, new_G4309_,
    new_G4310_, new_G4311_, new_G4312_, new_G4313_, new_G4314_, new_G4315_,
    new_G4316_, new_G4319_, new_G4320_, new_G4321_, new_G4322_, new_G4323_,
    new_G4329_, new_G4330_, new_G4331_, new_G4332_, new_G4333_, new_G4334_,
    new_G4335_, new_G4336_, new_G4339_, new_G4340_, new_G4343_, new_G4344_,
    new_G4345_, new_G4346_, new_G4349_, new_G4350_, new_G4351_, new_G4352_,
    new_G4355_, new_G4356_, new_G4359_, new_G4360_, new_G4363_, new_G4364_,
    new_G4367_, new_G4368_, new_G4369_, new_G4370_, new_G4371_, new_G4374_,
    new_G4375_, new_G4376_, new_G4377_, new_G4378_, new_G4381_, new_G4382_,
    new_G4383_, new_G4384_, new_G4385_, new_G4386_, new_G4387_, new_G4388_,
    new_G4389_, new_G4390_, new_G4391_, new_G4392_, new_G4393_, new_G4394_,
    new_G4395_, new_G4396_, new_G4397_, new_G4398_, new_G4399_, new_G4400_,
    new_G4403_, new_G4404_, new_G4405_, new_G4406_, new_G4407_, new_G4408_,
    new_G4409_, new_G4413_, new_G4414_, new_G4415_, new_G4416_, new_G4417_,
    new_G4420_, new_G4423_, new_G4424_, new_G4425_, new_G4426_, new_G4427_,
    new_G4428_, new_G4429_, new_G4430_, new_G4431_, new_G4432_, new_G4437_,
    new_G4440_, new_G4443_, new_G4446_, new_G4449_, new_G4450_, new_G4453_,
    new_G4454_, new_G4455_, new_G4456_, new_G4457_, new_G4458_, new_G4463_,
    new_G4466_, new_G4469_, new_G4472_, new_G4473_, new_G4476_, new_G4477_,
    new_G4478_, new_G4479_, new_G4480_, new_G4483_, new_G4484_, new_G4487_,
    new_G4488_, new_G4489_, new_G4490_, new_G4491_, new_G4492_, new_G4493_,
    new_G4494_, new_G4497_, new_G4498_, new_G4501_, new_G4504_, new_G4507_,
    new_G4508_, new_G4509_, new_G4510_, new_G4511_, new_G4512_, new_G4513_,
    new_G4514_, new_G4515_, new_G4516_, new_G4517_, new_G4518_, new_G4519_,
    new_G4520_, new_G4521_, new_G4522_, new_G4523_, new_G4524_, new_G4525_,
    new_G4526_, new_G4527_, new_G4528_, new_G4529_, new_G4530_, new_G4531_,
    new_G4532_, new_G4533_, new_G4534_, new_G4535_, new_G4536_, new_G4537_,
    new_G4538_, new_G4539_, new_G4540_, new_G4541_, new_G4542_, new_G4543_,
    new_G4544_, new_G4545_, new_G4546_, new_G4547_, new_G4548_, new_G4549_,
    new_G4550_, new_G4551_, new_G4552_, new_G4553_, new_G4554_, new_G4560_,
    new_G4561_, new_G4562_, new_G4568_, new_G4569_, new_G4570_, new_G4571_,
    new_G4572_, new_G4573_, new_G4576_, new_G4579_, new_G4580_, new_G4581_,
    new_G4582_, new_G4583_, new_G4586_, new_G4589_, new_G4592_, new_G4593_,
    new_G4594_, new_G4597_, new_G4600_, new_G4603_, new_G4606_, new_G4613_,
    new_G4616_, new_G4619_, new_G4622_, new_G4623_, new_G4624_, new_G4630_,
    new_G4636_, new_G4642_, new_G4648_, new_G4654_, new_G4655_, new_G4658_,
    new_G4664_, new_G4670_, new_G4671_, new_G4672_, new_G4673_, new_G4674_,
    new_G4675_, new_G4676_, new_G4677_, new_G4678_, new_G4679_, new_G4680_,
    new_G4681_, new_G4684_, new_G4687_, new_G4690_, new_G4691_, new_G4692_,
    new_G4693_, new_G4694_, new_G4697_, new_G4700_, new_G4701_, new_G4702_,
    new_G4703_, new_G4704_, new_G4705_, new_G4706_, new_G4709_, new_G4710_,
    new_G4711_, new_G4712_, new_G4713_, new_G4714_, new_G4715_, new_G4716_,
    new_G4717_, new_G4718_, new_G4719_, new_G4720_, new_G4721_, new_G4722_,
    new_G4723_, new_G4724_, new_G4725_, new_G4726_, new_G4727_, new_G4728_,
    new_G4729_, new_G4730_, new_G4731_, new_G4732_, new_G4733_, new_G4734_,
    new_G4735_, new_G4736_, new_G4737_, new_G4738_, new_G4739_, new_G4740_,
    new_G4741_, new_G4742_, new_G4743_, new_G4744_, new_G4745_, new_G4746_,
    new_G4747_, new_G4748_, new_G4749_, new_G4750_, new_G4751_, new_G4752_,
    new_G4753_, new_G4754_, new_G4755_, new_G4756_, new_G4757_, new_G4758_,
    new_G4761_, new_G4762_, new_G4763_, new_G4764_, new_G4765_, new_G4766_,
    new_G4767_, new_G4768_, new_G4769_, new_G4770_, new_G4771_, new_G4772_,
    new_G4773_, new_G4774_, new_G4775_, new_G4776_, new_G4777_, new_G4778_,
    new_G4779_, new_G4780_, new_G4786_, new_G4792_, new_G4798_, new_G4804_,
    new_G4810_, new_G4816_, new_G4822_, new_G4828_, new_G4831_, new_G4834_,
    new_G4835_, new_G4836_, new_G4837_, new_G4838_, new_G4841_, new_G4844_,
    new_G4847_, new_G4848_, new_G4849_, new_G4850_, new_G4851_, new_G4852_,
    new_G4853_, new_G4854_, new_G4855_, new_G4856_, new_G4857_, new_G4858_,
    new_G4859_, new_G4860_, new_G4861_, new_G4862_, new_G4863_, new_G4864_,
    new_G4865_, new_G4866_, new_G4867_, new_G4868_, new_G4869_, new_G4870_,
    new_G4871_, new_G4872_, new_G4873_, new_G4874_, new_G4875_, new_G4876_,
    new_G4877_, new_G4878_, new_G4879_, new_G4880_, new_G4881_, new_G4882_,
    new_G4883_, new_G4884_, new_G4885_, new_G4886_, new_G4887_, new_G4888_,
    new_G4889_, new_G4890_, new_G4891_, new_G4892_, new_G4895_, new_G4898_,
    new_G4899_, new_G4900_, new_G4901_, new_G4902_, new_G4903_, new_G4904_,
    new_G4907_, new_G4908_, new_G4909_, new_G4910_, new_G4911_, new_G4912_,
    new_G4913_, new_G4914_, new_G4915_, new_G4916_, new_G4917_, new_G4918_,
    new_G4919_, new_G4920_, new_G4923_, new_G4926_, new_G4927_, new_G4928_,
    new_G4929_, new_G4930_, new_G4933_, new_G4936_, new_G4939_, new_G4940_,
    new_G4941_, new_G4942_, new_G4943_, new_G4944_, new_G4945_, new_G4946_,
    new_G4947_, new_G4948_, new_G4951_, new_G4954_, new_G4955_, new_G4956_,
    new_G4957_, new_G4958_, new_G4959_, new_G4960_, new_G4963_, new_G4964_,
    new_G4965_, new_G4966_, new_G4967_, new_G4968_, new_G4971_, new_G4974_,
    new_G4975_, new_G4976_, new_G4977_, new_G4978_, new_G4981_, new_G4984_,
    new_G4987_, new_G4988_, new_G4989_, new_G4990_, new_G4991_, new_G4992_,
    new_G4993_, new_G4994_, new_G4995_, new_G4996_, new_G4999_, new_G5002_,
    new_G5003_, new_G5004_, new_G5005_, new_G5006_, new_G5007_, new_G5008_,
    new_G5011_, new_G5012_, new_G5013_, new_G5014_, new_G5015_, new_G5016_,
    new_G5019_, new_G5022_, new_G5023_, new_G5024_, new_G5025_, new_G5026_,
    new_G5029_, new_G5032_, new_G5035_, new_G5036_, new_G5037_, new_G5038_,
    new_G5039_, new_G5040_, new_G5041_, new_G5042_, new_G5043_, new_G5044_,
    new_G5045_, new_G5046_, new_G5047_, new_G5048_, new_G5051_, new_G5054_,
    new_G5055_, new_G5056_, new_G5059_, new_G5060_, new_G5061_, new_G5062_,
    new_G5063_, new_G5064_, new_G5067_, new_G5070_, new_G5073_, new_G5076_,
    new_G5077_, new_G5078_, new_G5079_, new_G5080_, new_G5083_, new_G5084_,
    new_G5085_, new_G5086_, new_G5087_, new_G5088_, new_G5089_, new_G5090_,
    new_G5091_, new_G5092_, new_G5093_, new_G5094_, new_G5095_, new_G5096_,
    new_G5097_, new_G5098_, new_G5101_, new_G5104_, new_G5107_, new_G5108_,
    new_G5111_, new_G5114_, new_G5115_, new_G5116_, new_G5117_, new_G5118_,
    new_G5119_, new_G5120_, new_G5121_, new_G5122_, new_G5123_, new_G5124_,
    new_G5125_, new_G5126_, new_G5127_, new_G5128_, new_G5129_, new_G5130_,
    new_G5131_, new_G5132_, new_G5133_, new_G5134_, new_G5135_, new_G5138_,
    new_G5141_, new_G5142_, new_G5143_, new_G5144_, new_G5145_, new_G5146_,
    new_G5147_, new_G5150_, new_G5153_, new_G5154_, new_G5155_, new_G5156_,
    new_G5157_, new_G5158_, new_G5159_, new_G5162_, new_G5165_, new_G5166_,
    new_G5167_, new_G5168_, new_G5169_, new_G5172_, new_G5175_, new_G5178_,
    new_G5181_, new_G5182_, new_G5183_, new_G5184_, new_G5185_, new_G5186_,
    new_G5187_, new_G5188_, new_G5189_, new_G5190_, new_G5191_, new_G5192_,
    n2610_li, n2613_li, n2616_li, n2619_li, n2622_li, n2625_li, n2628_li,
    n2631_li, n2634_li, n2637_li, n2640_li, n2643_li, n2646_li, n2649_li,
    n2652_li, n2655_li, n2658_li, n2661_li, n2664_li, n2667_li, n2670_li,
    n2673_li, n2676_li, n2679_li, n2682_li, n2685_li, n2688_li, n2691_li,
    n2694_li, n2697_li, n2700_li, n2703_li, n2706_li, n2709_li, n2712_li,
    n2715_li, n2718_li, n2721_li, n2724_li, n2727_li, n2730_li, n2733_li,
    n2736_li, n2739_li, n2742_li, n2745_li, n2748_li, n2751_li, n2754_li,
    n2757_li, n2760_li, n2763_li, n2766_li, n2769_li, n2772_li, n2775_li,
    n2778_li, n2781_li, n2784_li, n2787_li, n2790_li, n2793_li, n2796_li,
    n2799_li, n2802_li, n2805_li, n2808_li, n2811_li, n2814_li, n2817_li,
    n2820_li, n2823_li, n2826_li, n2829_li, n2832_li, n2835_li, n2838_li,
    n2841_li, n2844_li, n2847_li, n2850_li, n2853_li, n2856_li, n2859_li,
    n2862_li, n2865_li, n2868_li, n2871_li, n2874_li, n2877_li, n2880_li,
    n2883_li, n2886_li, n2889_li, n2892_li, n2895_li, n2898_li, n2901_li,
    n2904_li, n2907_li, n2910_li, n2913_li, n2916_li, n2919_li, n2922_li,
    n2925_li, n2928_li, n2931_li, n2934_li, n2937_li, n2940_li, n2943_li,
    n2946_li, n2949_li, n2952_li, n2955_li, n2958_li, n2961_li, n2964_li,
    n2967_li, n2970_li, n2973_li, n2976_li, n2979_li, n2982_li, n2985_li,
    n2988_li, n2991_li, n2994_li, n2997_li, n3000_li, n3003_li, n3006_li,
    n3009_li, n3012_li, n3015_li, n3018_li, n3021_li, n3024_li, n3027_li,
    n3030_li, n3033_li, n3036_li, n3039_li, n3042_li, n3045_li, n3048_li,
    n3051_li, n3054_li, n3057_li, n3060_li, n3063_li, n3066_li, n3069_li,
    n3072_li, n3075_li, n3078_li, n3081_li, n3084_li, n3087_li, n3090_li,
    n3093_li, n3096_li, n3099_li, n3102_li, n3105_li, n3108_li, n3111_li,
    n3114_li, n3117_li, n3120_li, n3123_li, n3126_li, n3129_li, n3132_li,
    n3135_li, n3138_li, n3141_li, n3144_li, n3147_li, n3150_li, n3153_li,
    n3156_li, n3159_li, n3162_li, n3165_li, n3168_li, n3171_li, n3174_li,
    n3177_li, n3180_li, n3183_li, n3186_li, n3189_li, n3192_li, n3195_li,
    n3198_li, n3201_li, n3204_li, n3207_li, n3210_li, n3213_li, n3216_li,
    n3219_li, n3222_li, n3225_li, n3228_li, n3231_li, n3234_li, n3237_li,
    n3240_li, n3243_li, n3246_li, n3249_li, n3252_li, n3255_li, n3258_li,
    n3261_li, n3264_li, n3267_li, n3270_li, n3273_li, n3276_li, n3279_li,
    n3282_li, n3285_li, n3288_li, n3291_li, n3294_li, n3297_li, n3300_li,
    n3303_li, n3306_li, n3309_li, n3312_li, n3315_li, n3318_li, n3321_li,
    n3324_li, n3327_li, n3330_li, n3333_li, n3336_li, n3339_li, n3342_li,
    n3345_li, n3348_li, n3351_li, n3354_li, n3357_li, n3360_li, n3363_li,
    n3366_li, n3369_li, n3372_li, n3375_li, n3378_li, n3381_li, n3384_li,
    n3387_li, n3390_li, n3393_li, n3396_li, n3399_li, n3402_li, n3405_li,
    n3408_li, n3411_li, n3414_li, n3417_li, n3420_li, n3423_li, n3426_li,
    n3429_li, n3432_li, n3435_li, n3438_li, n3441_li, n3444_li, n3447_li,
    n3450_li, n3453_li, n3456_li, n3459_li, n3462_li, n3465_li, n3468_li,
    n3471_li, n3474_li, n3477_li, n3480_li, n3483_li, n3486_li, n3489_li,
    n3492_li, n3495_li, n3498_li, n3501_li, n3504_li, n3507_li, n3510_li,
    n3513_li, n3516_li, n3519_li, n3522_li, n3525_li, n3528_li, n3531_li,
    n3534_li, n3537_li, n3540_li, n3543_li, n3546_li, n3549_li, n3552_li,
    n3555_li, n3558_li, n3561_li, n3564_li, n3567_li, n3570_li, n3573_li,
    n3576_li, n3579_li, n3582_li, n3585_li, n3588_li, n3591_li, n3594_li,
    n3597_li, n3600_li, n3603_li, n3606_li, n3609_li, n3612_li, n3615_li,
    n3618_li, n3621_li, n3624_li, n3627_li, n3630_li, n3633_li, n3636_li,
    n3639_li, n3642_li, n3645_li, n3648_li, n3651_li, n3654_li, n3657_li,
    n3660_li, n3663_li, n3666_li, n3669_li, n3672_li, n3675_li, n3678_li,
    n3681_li, n3684_li, n3687_li, n3690_li, n3693_li, n3696_li, n3699_li,
    n3702_li, n3705_li, n3708_li, n3711_li, n3714_li, n3717_li, n3720_li,
    n3723_li, n3726_li, n3729_li, n3732_li, n3735_li, n3738_li, n3741_li,
    n3744_li, n3747_li, n3750_li, n3753_li, n3756_li, n3759_li, n3762_li,
    n3765_li, n3768_li, n3771_li, n3774_li, n3777_li, n3780_li, n3783_li,
    n3786_li, n3789_li, n3792_li, n3795_li, n3798_li, n3801_li, n3804_li,
    n3807_li, n3810_li, n3813_li, n3816_li, n3819_li, n3822_li, n3825_li,
    n3828_li, n3831_li, n3834_li, n3837_li, n3840_li, n3843_li, n3846_li,
    n3849_li, n3852_li, n3855_li, n3858_li, n3861_li, n3864_li, n3867_li,
    n3870_li, n3873_li, n3876_li, n3879_li, n3882_li, n3885_li, n3888_li,
    n3891_li, n3894_li, n3897_li, n3900_li, n3903_li, n3906_li, n3909_li,
    n3912_li, n3915_li, n3918_li, n3921_li, n3924_li, n3927_li, n3930_li,
    n3933_li, n3936_li, n3939_li, n3942_li, n3945_li, n3948_li, n3951_li,
    n3954_li, n3957_li, n3960_li, n3963_li, n3966_li, n3969_li, n3972_li,
    n3975_li, n3978_li, n3981_li, n3984_li, n3987_li, n3990_li, n3993_li,
    n3996_li, n3999_li, n4002_li, n4005_li, n4008_li, n4011_li, n4014_li,
    n4017_li, n4020_li, n4023_li, n4026_li, n4029_li, n4032_li, n4035_li,
    n4038_li, n4041_li, n4044_li, n4047_li, n4050_li, n4053_li, n4056_li,
    n4059_li, n4062_li, n4065_li, n4068_li, n4071_li, n4074_li, n4077_li,
    n4080_li, n4083_li, n4086_li, n4089_li, n4092_li, n4095_li, n4098_li,
    n4101_li, n4104_li, n4107_li, n4110_li, n4113_li, n4116_li, n4119_li,
    n4122_li, n4125_li, n4128_li, n4131_li, n4134_li, n4137_li, n4140_li,
    n4143_li, n4146_li, n4149_li, n4152_li, n4155_li, n4158_li, n4161_li,
    n4164_li, n4167_li, n4170_li, n4173_li, n4176_li, n4179_li, n4182_li,
    n4185_li, n4188_li, n4191_li, n4194_li, n4197_li, n4200_li, n4203_li,
    n4206_li, n4209_li, n4212_li, n4215_li, n4218_li, n4221_li, n4224_li,
    n4227_li, n4230_li, n4233_li, n4236_li, n4239_li, n4242_li, n4245_li,
    n4248_li, n4251_li, n4254_li, n4257_li, n4260_li, n4263_li, n4266_li,
    n4269_li, n4272_li, n4275_li, n4278_li, n4281_li, n4284_li, n4287_li,
    n4290_li, n4293_li, n4296_li, n4299_li, n4302_li, n4305_li, n4308_li,
    n4311_li, n4314_li, n4317_li, n4320_li, n4323_li, n4326_li, n4329_li,
    n4332_li, n4335_li, n4338_li, n4341_li, n4344_li, n4347_li, n4350_li,
    n4353_li, n4356_li, n4359_li, n4362_li, n4365_li, n4368_li, n4371_li,
    n4374_li, n4377_li, n4380_li, n4383_li, n4386_li, n4389_li, n4392_li,
    n4395_li, n4398_li, n4401_li, n4404_li, n4407_li, n4410_li, n4413_li,
    n4416_li, n4419_li, n4422_li, n4425_li, n4428_li, n4431_li, n4434_li,
    n4437_li, n4440_li, n4443_li, n4446_li, n4449_li, n4452_li, n4455_li,
    n4458_li, n4461_li, n4464_li, n4467_li, n4470_li, n4473_li, n4476_li,
    n4479_li, n4482_li, n4485_li, n4488_li, n4491_li, n4494_li, n4497_li,
    n4500_li, n4503_li, n4506_li, n4509_li, n4512_li, n4515_li, n4518_li,
    n4521_li, n4524_li, n4527_li, n4530_li, n4533_li, n4536_li, n4539_li,
    n4542_li, n4545_li, n4548_li, n4551_li, n4554_li, n4557_li, n4560_li,
    n4563_li, n4566_li, n4569_li, n4572_li, n4575_li, n4578_li, n4581_li,
    n4584_li, n4587_li, n4590_li, n4593_li, n4596_li, n4599_li, n4602_li,
    n4605_li, n4608_li, n4611_li, n4614_li, n4617_li, n4620_li, n4623_li,
    n4626_li, n4629_li, n4632_li, n4635_li, n4638_li, n4641_li, n4644_li,
    n4647_li, n4650_li, n4653_li, n4656_li, n4659_li, n4662_li, n4665_li,
    n4668_li, n4671_li, n4674_li, n4677_li, n4680_li, n4683_li, n4686_li,
    n4689_li, n4692_li, n4695_li, n4698_li, n4701_li, n4704_li, n4707_li,
    n4710_li, n4713_li, n4716_li, n4719_li, n4722_li, n4725_li, n4728_li,
    n4731_li, n4734_li, n4737_li, n4740_li, n4743_li;
  assign new_G632_ = n3351_lo & n4743_lo;
  assign new_G633_ = ~n4575_lo;
  assign new_G634_ = ~n4599_lo;
  assign new_G647_ = ~n4611_lo;
  assign new_G659_ = ~n4623_lo;
  assign new_G671_ = ~n4635_lo;
  assign new_G684_ = ~n4215_lo | ~n2619_lo;
  assign new_G685_ = ~n4587_lo;
  assign new_G686_ = ~new_G632_;
  assign new_G687_ = new_G633_ & n2739_lo;
  assign new_G688_ = n4239_lo & n4455_lo;
  assign new_G689_ = n4443_lo & n4239_lo & n4467_lo & n4455_lo;
  assign new_G690_ = ~n4491_lo;
  assign new_G694_ = ~n4503_lo;
  assign new_G706_ = ~n4515_lo;
  assign new_G718_ = ~n4503_lo;
  assign new_G730_ = ~n4515_lo;
  assign new_G742_ = ~n3375_lo;
  assign new_G746_ = ~n3375_lo;
  assign new_G749_ = ~n3399_lo;
  assign new_G752_ = ~n4551_lo;
  assign new_G756_ = ~n4527_lo;
  assign new_G768_ = ~n4539_lo;
  assign new_G780_ = ~n4527_lo;
  assign new_G792_ = ~n4539_lo;
  assign new_G804_ = ~n3831_lo;
  assign new_G813_ = ~n3819_lo;
  assign new_G825_ = ~n3819_lo;
  assign new_G836_ = ~n3807_lo;
  assign new_G848_ = ~n3807_lo;
  assign new_G860_ = ~n4683_lo;
  assign new_G872_ = ~n4671_lo;
  assign new_G884_ = ~n4695_lo;
  assign new_G896_ = ~n4707_lo;
  assign new_G908_ = ~n3687_lo;
  assign new_G911_ = ~n3687_lo;
  assign new_G914_ = ~n3711_lo;
  assign new_G917_ = ~n3711_lo;
  assign new_G920_ = ~n3735_lo;
  assign new_G923_ = ~n3735_lo;
  assign new_G926_ = ~n3759_lo;
  assign new_G929_ = ~n3759_lo;
  assign new_G932_ = ~n3843_lo;
  assign new_G935_ = ~n3843_lo;
  assign new_G938_ = ~n3867_lo;
  assign new_G941_ = ~n3867_lo;
  assign new_G944_ = ~n3891_lo;
  assign new_G947_ = ~n3891_lo;
  assign new_G950_ = ~n3915_lo;
  assign new_G953_ = ~n3915_lo;
  assign new_G956_ = ~n4095_lo;
  assign new_G963_ = ~n4095_lo;
  assign new_G970_ = ~n3663_lo;
  assign new_G976_ = n2739_lo & n2751_lo;
  assign new_G980_ = ~n2619_lo;
  assign new_G983_ = ~n4563_lo;
  assign new_G993_ = ~n3963_lo;
  assign new_G996_ = ~n3987_lo;
  assign new_G999_ = ~n4011_lo;
  assign new_G1002_ = ~n4011_lo;
  assign new_G1005_ = ~n4035_lo;
  assign new_G1008_ = ~n4035_lo;
  assign new_G1011_ = ~n4059_lo;
  assign new_G1014_ = ~n4059_lo;
  assign new_G1017_ = ~n4119_lo;
  assign new_G1020_ = ~n4119_lo;
  assign new_G1023_ = ~n4143_lo;
  assign new_G1026_ = ~n4143_lo;
  assign new_G1029_ = ~n3843_lo;
  assign new_G1032_ = ~n3843_lo;
  assign new_G1035_ = ~n3867_lo;
  assign new_G1038_ = ~n3867_lo;
  assign new_G1041_ = ~n3891_lo;
  assign new_G1044_ = ~n3891_lo;
  assign new_G1047_ = ~n3915_lo;
  assign new_G1050_ = ~n3915_lo;
  assign new_G1053_ = ~n4083_lo;
  assign new_G1060_ = ~n4083_lo;
  assign new_G1067_ = ~n4431_lo;
  assign new_G1070_ = n2751_lo & n2739_lo;
  assign new_G1075_ = ~n4563_lo;
  assign new_G1081_ = ~n4059_lo;
  assign new_G1084_ = ~n4059_lo;
  assign new_G1087_ = ~n4119_lo;
  assign new_G1090_ = ~n4119_lo;
  assign new_G1093_ = ~n4143_lo;
  assign new_G1096_ = ~n4143_lo;
  assign new_G1099_ = ~n3963_lo;
  assign new_G1102_ = ~n3987_lo;
  assign new_G1105_ = ~n4011_lo;
  assign new_G1108_ = ~n4011_lo;
  assign new_G1111_ = ~n4035_lo;
  assign new_G1114_ = ~n4035_lo;
  assign new_G1117_ = ~n4167_lo;
  assign new_G1120_ = ~n4167_lo;
  assign new_G1123_ = ~n3687_lo;
  assign new_G1126_ = ~n3687_lo;
  assign new_G1129_ = ~n3711_lo;
  assign new_G1132_ = ~n3711_lo;
  assign new_G1135_ = ~n3735_lo;
  assign new_G1138_ = ~n3735_lo;
  assign new_G1141_ = ~n3759_lo;
  assign new_G1144_ = ~n3759_lo;
  assign new_G1147_ = ~n4059_lo;
  assign new_G1150_ = ~n3783_lo;
  assign new_G1162_ = ~n3783_lo;
  assign new_G1172_ = ~n3831_lo;
  assign new_G1184_ = ~n4683_lo;
  assign new_G1196_ = ~n4671_lo;
  assign new_G1208_ = ~n4731_lo;
  assign new_G1214_ = ~n4719_lo;
  assign new_G1218_ = ~n4695_lo;
  assign new_G1230_ = ~n4707_lo;
  assign new_G1242_ = ~n4647_lo;
  assign new_G1245_ = ~n4659_lo;
  assign new_G1248_ = ~n4719_lo;
  assign new_G1256_ = ~n4731_lo;
  assign new_G1264_ = ~n4719_lo;
  assign new_G1272_ = ~n4731_lo;
  assign new_G1280_ = ~n4719_lo;
  assign new_G1287_ = ~n4731_lo;
  assign new_G1294_ = ~n4719_lo;
  assign new_G1301_ = ~n4731_lo;
  assign new_G1308_ = ~n3975_lo;
  assign new_G1311_ = ~n4311_lo;
  assign new_G1314_ = ~n4323_lo;
  assign new_G1317_ = ~n4335_lo;
  assign new_G1320_ = ~n4287_lo;
  assign new_G1323_ = ~n4299_lo;
  assign new_G1326_ = ~n4251_lo;
  assign new_G1329_ = ~n4263_lo;
  assign new_G1332_ = ~n4275_lo;
  assign new_G1335_ = ~n4227_lo;
  assign new_G1338_ = ~n2631_lo;
  assign new_G1341_ = ~n4311_lo;
  assign new_G1344_ = ~n4323_lo;
  assign new_G1347_ = ~n4335_lo;
  assign new_G1350_ = ~n4299_lo;
  assign new_G1353_ = ~n4251_lo;
  assign new_G1356_ = ~n4263_lo;
  assign new_G1359_ = ~n4275_lo;
  assign new_G1362_ = ~n4287_lo;
  assign new_G1365_ = ~n4227_lo;
  assign new_G1368_ = ~n4347_lo;
  assign new_G1371_ = ~n4359_lo;
  assign new_G1374_ = ~n4371_lo;
  assign new_G1377_ = ~n4383_lo;
  assign new_G1380_ = ~n4395_lo;
  assign new_G1383_ = ~n4407_lo;
  assign new_G1386_ = ~n2859_lo;
  assign new_G1389_ = ~n4347_lo;
  assign new_G1392_ = ~n4371_lo;
  assign new_G1395_ = ~n4383_lo;
  assign new_G1398_ = ~n4395_lo;
  assign new_G1401_ = ~n4407_lo;
  assign new_G1404_ = ~n4359_lo;
  assign new_G1407_ = ~n4167_lo;
  assign new_G1410_ = ~n4191_lo;
  assign new_G1413_ = ~n4119_lo;
  assign new_G1416_ = ~n4143_lo;
  assign new_G1419_ = ~n4011_lo;
  assign new_G1422_ = ~n4035_lo;
  assign new_G1425_ = ~n3963_lo;
  assign new_G1428_ = ~n3987_lo;
  assign new_G1431_ = ~n3915_lo;
  assign new_G1434_ = ~n3939_lo;
  assign new_G1437_ = ~n3867_lo;
  assign new_G1440_ = ~n3891_lo;
  assign new_G1443_ = ~n3759_lo;
  assign new_G1446_ = ~n3843_lo;
  assign new_G1449_ = ~n3711_lo;
  assign new_G1452_ = ~n3735_lo;
  assign new_G1455_ = ~n3687_lo;
  assign new_G1458_ = new_G671_ & n4383_lo;
  assign new_G1459_ = new_G634_ | n4383_lo;
  assign new_G1460_ = n3519_lo & new_G694_ & new_G706_;
  assign new_G1461_ = n3531_lo & new_G694_ & new_G706_;
  assign new_G1462_ = n3507_lo & new_G694_ & new_G706_;
  assign new_G1463_ = n3495_lo & new_G694_ & new_G706_;
  assign new_G1464_ = n3483_lo & new_G694_ & new_G706_;
  assign new_G1465_ = n3579_lo & new_G718_ & new_G730_;
  assign new_G1466_ = n3471_lo & new_G718_ & new_G730_;
  assign new_G1467_ = n3447_lo & new_G718_ & new_G730_;
  assign new_G1468_ = n3423_lo & new_G718_ & new_G730_;
  assign new_G1469_ = n3519_lo & new_G756_ & new_G768_;
  assign new_G1470_ = n3531_lo & new_G756_ & new_G768_;
  assign new_G1471_ = n3507_lo & new_G756_ & new_G768_;
  assign new_G1472_ = n3495_lo & new_G756_ & new_G768_;
  assign new_G1473_ = n3483_lo & new_G756_ & new_G768_;
  assign new_G1474_ = n3579_lo & new_G780_ & new_G792_;
  assign new_G1475_ = n3471_lo & new_G780_ & new_G792_;
  assign new_G1476_ = n3447_lo & new_G780_ & new_G792_;
  assign new_G1477_ = n3423_lo & new_G780_ & new_G792_;
  assign new_G1478_ = n3099_lo & new_G1218_ & new_G1230_;
  assign new_G1479_ = n2871_lo & new_G860_ & new_G872_;
  assign new_G1480_ = n3099_lo & new_G1184_ & new_G1196_;
  assign new_G1481_ = n2823_lo & new_G1184_ & new_G1196_;
  assign new_G1482_ = n3087_lo & new_G1184_ & new_G1196_;
  assign new_G1483_ = n2787_lo & new_G1184_ & new_G1196_;
  assign new_G1484_ = n2775_lo & new_G1184_ & new_G1196_;
  assign new_G1485_ = n2679_lo & new_G860_ & new_G872_;
  assign new_G1486_ = n2667_lo & new_G860_ & new_G872_;
  assign new_G1487_ = n2907_lo & new_G860_ & new_G872_;
  assign new_G1488_ = n2883_lo & new_G860_ & new_G872_;
  assign new_G1489_ = n2823_lo & new_G1218_ & new_G1230_;
  assign new_G1490_ = n3087_lo & new_G1218_ & new_G1230_;
  assign new_G1491_ = n2787_lo & new_G1218_ & new_G1230_;
  assign new_G1492_ = n2775_lo & new_G1218_ & new_G1230_;
  assign new_G1493_ = n2679_lo & new_G884_ & new_G896_;
  assign new_G1494_ = n2667_lo & new_G884_ & new_G896_;
  assign new_G1495_ = n2907_lo & new_G884_ & new_G896_;
  assign new_G1496_ = n2883_lo & new_G884_ & new_G896_;
  assign new_G1497_ = n3255_lo & new_G1245_ & n4647_lo;
  assign new_G1498_ = new_G1264_ & new_G1272_;
  assign new_G1499_ = n2871_lo & new_G884_ & new_G896_;
  assign new_G1500_ = new_G1248_ & new_G1256_;
  assign new_G1501_ = ~new_G1311_;
  assign new_G1502_ = ~new_G1314_;
  assign new_G1503_ = ~new_G1317_;
  assign new_G1504_ = ~new_G1320_;
  assign new_G1505_ = ~new_G1323_;
  assign new_G1506_ = ~new_G1326_;
  assign new_G1507_ = ~new_G1329_;
  assign new_G1508_ = ~new_G1332_;
  assign new_G1509_ = ~new_G1335_;
  assign new_G1510_ = ~new_G1338_;
  assign new_G1511_ = ~new_G1341_;
  assign new_G1512_ = ~new_G1344_;
  assign new_G1513_ = ~new_G1347_;
  assign new_G1514_ = ~new_G1350_;
  assign new_G1515_ = ~new_G1353_;
  assign new_G1516_ = ~new_G1356_;
  assign new_G1517_ = ~new_G1359_;
  assign new_G1518_ = ~new_G1362_;
  assign new_G1519_ = ~new_G1365_;
  assign new_G1520_ = ~new_G742_;
  assign new_G1526_ = ~new_G694_;
  assign new_G1537_ = ~new_G706_;
  assign new_G1548_ = ~new_G742_;
  assign new_G1554_ = ~new_G718_;
  assign new_G1565_ = ~new_G730_;
  assign new_G1576_ = n3555_lo & new_G718_ & new_G730_;
  assign new_G1577_ = ~new_G980_;
  assign new_G1582_ = ~new_G1368_;
  assign new_G1583_ = ~new_G1371_;
  assign new_G1584_ = ~new_G1374_;
  assign new_G1585_ = ~new_G1377_;
  assign new_G1586_ = ~new_G1380_;
  assign new_G1587_ = ~new_G1383_;
  assign new_G1588_ = ~new_G1386_;
  assign new_G1589_ = ~new_G1389_;
  assign new_G1590_ = ~new_G1392_;
  assign new_G1591_ = ~new_G1395_;
  assign new_G1592_ = ~new_G1398_;
  assign new_G1593_ = ~new_G1401_;
  assign new_G1594_ = ~new_G1404_;
  assign new_G1595_ = ~new_G746_;
  assign new_G1601_ = ~new_G756_;
  assign new_G1612_ = ~new_G768_;
  assign new_G1623_ = ~new_G746_;
  assign new_G1629_ = ~new_G780_;
  assign new_G1640_ = ~new_G792_;
  assign new_G1651_ = n3555_lo & new_G780_ & new_G792_;
  assign new_G1652_ = ~new_G860_;
  assign new_G1663_ = ~new_G872_;
  assign new_G1674_ = ~new_G884_;
  assign new_G1685_ = ~new_G896_;
  assign new_G1696_ = ~new_G908_;
  assign new_G1697_ = ~new_G911_;
  assign new_G1698_ = ~new_G914_;
  assign new_G1699_ = ~new_G917_;
  assign new_G1700_ = ~new_G920_;
  assign new_G1701_ = ~new_G923_;
  assign new_G1702_ = ~new_G926_;
  assign new_G1703_ = ~new_G929_;
  assign new_G1704_ = new_G671_ & n4323_lo & new_G911_;
  assign new_G1705_ = new_G671_ & n4335_lo & new_G917_;
  assign new_G1706_ = new_G671_ & n4287_lo & new_G923_;
  assign new_G1707_ = new_G671_ & n4299_lo & new_G929_;
  assign new_G1708_ = new_G634_ & new_G908_;
  assign new_G1709_ = new_G634_ & new_G914_;
  assign new_G1710_ = new_G634_ & new_G920_;
  assign new_G1711_ = new_G634_ & new_G926_;
  assign new_G1712_ = ~new_G932_;
  assign new_G1713_ = ~new_G935_;
  assign new_G1714_ = ~new_G938_;
  assign new_G1715_ = ~new_G941_;
  assign new_G1716_ = ~new_G944_;
  assign new_G1717_ = ~new_G947_;
  assign new_G1718_ = ~new_G950_;
  assign new_G1719_ = ~new_G953_;
  assign new_G1720_ = new_G671_ & n4251_lo & new_G935_;
  assign new_G1721_ = new_G671_ & n4263_lo & new_G941_;
  assign new_G1722_ = new_G671_ & n4275_lo & new_G947_;
  assign new_G1723_ = new_G671_ & n4227_lo & new_G953_;
  assign new_G1724_ = new_G634_ & new_G932_;
  assign new_G1725_ = new_G634_ & new_G938_;
  assign new_G1726_ = new_G634_ & new_G944_;
  assign new_G1727_ = new_G634_ & new_G950_;
  assign new_G1728_ = ~new_G956_;
  assign new_G1734_ = ~new_G963_;
  assign new_G1740_ = n3951_lo & new_G956_;
  assign new_G1741_ = n3927_lo & new_G956_;
  assign new_G1742_ = n3903_lo & new_G956_;
  assign new_G1743_ = n3879_lo & new_G956_;
  assign new_G1744_ = n3855_lo & new_G956_;
  assign new_G1745_ = n3771_lo & new_G963_;
  assign new_G1746_ = n3747_lo & new_G963_;
  assign new_G1747_ = n3723_lo & new_G963_;
  assign new_G1748_ = n3699_lo & new_G963_;
  assign new_G1749_ = n3675_lo & new_G963_;
  assign new_G1750_ = ~new_G749_;
  assign new_G1755_ = ~new_G983_;
  assign new_G1764_ = ~new_G976_;
  assign new_G1774_ = ~new_G993_;
  assign new_G1775_ = ~new_G996_;
  assign new_G1776_ = ~new_G999_;
  assign new_G1777_ = ~new_G1002_;
  assign new_G1778_ = ~new_G1005_;
  assign new_G1779_ = ~new_G1008_;
  assign new_G1780_ = new_G836_ & new_G996_;
  assign new_G1781_ = new_G836_ & n4347_lo & new_G1002_;
  assign new_G1782_ = new_G836_ & n4359_lo & new_G1008_;
  assign new_G1783_ = new_G1150_ & new_G993_;
  assign new_G1784_ = new_G1150_ & new_G999_;
  assign new_G1785_ = new_G1150_ & new_G1005_;
  assign new_G1786_ = ~new_G1011_;
  assign new_G1787_ = ~new_G1014_;
  assign new_G1788_ = ~new_G1017_;
  assign new_G1789_ = ~new_G1020_;
  assign new_G1790_ = ~new_G1023_;
  assign new_G1791_ = ~new_G1026_;
  assign new_G1792_ = new_G671_ & n4371_lo & new_G1014_;
  assign new_G1793_ = ~new_G1458_;
  assign new_G1794_ = new_G671_ & n4395_lo & new_G1020_;
  assign new_G1795_ = new_G671_ & n4407_lo & new_G1026_;
  assign new_G1796_ = new_G634_ & new_G1011_;
  assign new_G1797_ = new_G634_ & new_G1017_;
  assign new_G1798_ = new_G634_ & new_G1023_;
  assign new_G1799_ = ~new_G1029_;
  assign new_G1800_ = ~new_G1032_;
  assign new_G1801_ = ~new_G1035_;
  assign new_G1802_ = ~new_G1038_;
  assign new_G1803_ = ~new_G1041_;
  assign new_G1804_ = ~new_G1044_;
  assign new_G1805_ = ~new_G1047_;
  assign new_G1806_ = ~new_G1050_;
  assign new_G1807_ = new_G836_ & n4251_lo & new_G1032_;
  assign new_G1808_ = new_G836_ & n4263_lo & new_G1038_;
  assign new_G1809_ = new_G836_ & n4275_lo & new_G1044_;
  assign new_G1810_ = new_G836_ & n4227_lo & new_G1050_;
  assign new_G1811_ = new_G1150_ & new_G1029_;
  assign new_G1812_ = new_G1150_ & new_G1035_;
  assign new_G1813_ = new_G1150_ & new_G1041_;
  assign new_G1814_ = new_G1150_ & new_G1047_;
  assign new_G1815_ = ~new_G1053_;
  assign new_G1821_ = ~new_G1060_;
  assign new_G1827_ = n4203_lo & new_G1053_;
  assign new_G1828_ = n4179_lo & new_G1053_;
  assign new_G1829_ = n4155_lo & new_G1053_;
  assign new_G1830_ = n4131_lo & new_G1053_;
  assign new_G1831_ = n4107_lo & new_G1053_;
  assign new_G1832_ = n4071_lo & new_G1060_;
  assign new_G1833_ = n4047_lo & new_G1060_;
  assign new_G1834_ = n4023_lo & new_G1060_;
  assign new_G1835_ = n3999_lo & new_G1060_;
  assign new_G1836_ = n3975_lo & new_G1060_;
  assign new_G1837_ = ~new_G1075_;
  assign new_G1842_ = n2991_lo & new_G1075_;
  assign new_G1843_ = n3003_lo & new_G1075_;
  assign new_G1844_ = n3027_lo & new_G1075_;
  assign new_G1845_ = n3027_lo & new_G1075_;
  assign new_G1846_ = ~new_G1081_;
  assign new_G1847_ = ~new_G1084_;
  assign new_G1848_ = ~new_G1087_;
  assign new_G1849_ = ~new_G1090_;
  assign new_G1850_ = ~new_G1093_;
  assign new_G1851_ = ~new_G1096_;
  assign new_G1852_ = new_G848_ & n4371_lo & new_G1084_;
  assign new_G1853_ = new_G848_ & n4383_lo;
  assign new_G1854_ = new_G848_ & n4395_lo & new_G1090_;
  assign new_G1855_ = new_G848_ & n4407_lo & new_G1096_;
  assign new_G1856_ = new_G1162_ & new_G1081_;
  assign new_G1857_ = new_G1162_ | n4383_lo;
  assign new_G1858_ = new_G1162_ & new_G1087_;
  assign new_G1859_ = new_G1162_ & new_G1093_;
  assign new_G1860_ = ~new_G1099_;
  assign new_G1861_ = ~new_G1102_;
  assign new_G1862_ = ~new_G1105_;
  assign new_G1863_ = ~new_G1108_;
  assign new_G1864_ = ~new_G1111_;
  assign new_G1865_ = ~new_G1114_;
  assign new_G1866_ = new_G848_ & new_G1102_;
  assign new_G1867_ = new_G848_ & n4347_lo & new_G1108_;
  assign new_G1868_ = new_G848_ & n4359_lo & new_G1114_;
  assign new_G1869_ = new_G1162_ & new_G1099_;
  assign new_G1870_ = new_G1162_ & new_G1105_;
  assign new_G1871_ = new_G1162_ & new_G1111_;
  assign new_G1872_ = ~new_G1117_;
  assign new_G1873_ = ~new_G970_;
  assign new_G1876_ = ~new_G970_;
  assign new_G1879_ = ~new_G1120_;
  assign new_G1880_ = ~new_G970_;
  assign new_G1883_ = ~new_G970_;
  assign new_G1886_ = new_G848_ & new_G1117_;
  assign new_G1887_ = new_G848_ & new_G1120_;
  assign new_G1888_ = ~new_G1123_;
  assign new_G1889_ = ~new_G1126_;
  assign new_G1890_ = ~new_G1129_;
  assign new_G1891_ = ~new_G1132_;
  assign new_G1892_ = ~new_G1135_;
  assign new_G1893_ = ~new_G1138_;
  assign new_G1894_ = ~new_G1141_;
  assign new_G1895_ = ~new_G1144_;
  assign new_G1896_ = new_G836_ & n4323_lo & new_G1126_;
  assign new_G1897_ = new_G836_ & n4335_lo & new_G1132_;
  assign new_G1898_ = new_G836_ & n4287_lo & new_G1138_;
  assign new_G1899_ = new_G836_ & n4299_lo & new_G1144_;
  assign new_G1900_ = new_G1150_ & new_G1123_;
  assign new_G1901_ = new_G1150_ & new_G1129_;
  assign new_G1902_ = new_G1150_ & new_G1135_;
  assign new_G1903_ = new_G1150_ & new_G1141_;
  assign new_G1904_ = ~new_G1407_;
  assign new_G1905_ = ~new_G1410_;
  assign new_G1906_ = ~new_G1413_;
  assign new_G1907_ = ~new_G1416_;
  assign new_G1908_ = ~new_G1147_;
  assign new_G1911_ = ~new_G1147_;
  assign new_G1914_ = ~new_G1184_;
  assign new_G1925_ = ~new_G1196_;
  assign new_G1936_ = ~new_G1208_;
  assign new_G1941_ = ~new_G1214_;
  assign new_G1944_ = n3063_lo & new_G1208_;
  assign new_G1945_ = n3051_lo & new_G1208_;
  assign new_G1946_ = n3063_lo & new_G1208_;
  assign new_G1947_ = n3051_lo & new_G1208_;
  assign new_G1948_ = ~new_G1218_;
  assign new_G1959_ = ~new_G1230_;
  assign new_G1970_ = ~new_G1248_;
  assign new_G1981_ = ~new_G1256_;
  assign new_G1992_ = ~new_G1264_;
  assign new_G2003_ = ~new_G1272_;
  assign new_G2014_ = ~new_G1431_;
  assign new_G2015_ = ~new_G1434_;
  assign new_G2016_ = ~new_G1437_;
  assign new_G2017_ = ~new_G1440_;
  assign new_G2018_ = ~new_G1443_;
  assign new_G2019_ = ~new_G1446_;
  assign new_G2020_ = ~new_G1280_;
  assign new_G2031_ = ~new_G1287_;
  assign new_G2042_ = ~new_G1294_;
  assign new_G2053_ = ~new_G1301_;
  assign new_G2064_ = ~new_G1308_;
  assign new_G2067_ = ~new_G1419_;
  assign new_G2068_ = ~new_G1422_;
  assign new_G2069_ = ~new_G1425_;
  assign new_G2070_ = ~new_G1428_;
  assign new_G2071_ = ~new_G1449_;
  assign new_G2072_ = ~new_G1452_;
  assign new_G2073_ = ~new_G970_;
  assign new_G2076_ = ~new_G1455_;
  assign new_G2077_ = n4323_lo & new_G659_ & new_G1697_;
  assign new_G2078_ = n4335_lo & new_G659_ & new_G1699_;
  assign new_G2079_ = n4287_lo & new_G659_ & new_G1701_;
  assign new_G2080_ = n4299_lo & new_G659_ & new_G1703_;
  assign new_G2081_ = new_G647_ & new_G1696_;
  assign new_G2082_ = new_G647_ & new_G1698_;
  assign new_G2083_ = new_G647_ & new_G1700_;
  assign new_G2084_ = new_G647_ & new_G1702_;
  assign new_G2085_ = n4251_lo & new_G659_ & new_G1713_;
  assign new_G2086_ = n4263_lo & new_G659_ & new_G1715_;
  assign new_G2087_ = n4275_lo & new_G659_ & new_G1717_;
  assign new_G2088_ = n4227_lo & new_G659_ & new_G1719_;
  assign new_G2089_ = new_G647_ & new_G1712_;
  assign new_G2090_ = new_G647_ & new_G1714_;
  assign new_G2091_ = new_G647_ & new_G1716_;
  assign new_G2092_ = new_G647_ & new_G1718_;
  assign new_G2093_ = new_G813_ & new_G1775_;
  assign new_G2094_ = n4347_lo & new_G813_ & new_G1777_;
  assign new_G2095_ = n4359_lo & new_G813_ & new_G1779_;
  assign new_G2096_ = new_G1172_ & new_G1774_;
  assign new_G2097_ = new_G1172_ & new_G1776_;
  assign new_G2098_ = new_G1172_ & new_G1778_;
  assign new_G2099_ = n4371_lo & new_G659_ & new_G1787_;
  assign new_G2100_ = n4395_lo & new_G659_ & new_G1789_;
  assign new_G2101_ = n4407_lo & new_G659_ & new_G1791_;
  assign new_G2102_ = new_G647_ & new_G1786_;
  assign new_G2103_ = new_G647_ & new_G1788_;
  assign new_G2104_ = new_G647_ & new_G1790_;
  assign new_G2105_ = new_G1793_ & new_G1459_;
  assign new_G2108_ = n4251_lo & new_G813_ & new_G1800_;
  assign new_G2109_ = n4263_lo & new_G813_ & new_G1802_;
  assign new_G2110_ = n4275_lo & new_G813_ & new_G1804_;
  assign new_G2111_ = n4227_lo & new_G813_ & new_G1806_;
  assign new_G2112_ = new_G1172_ & new_G1799_;
  assign new_G2113_ = new_G1172_ & new_G1801_;
  assign new_G2114_ = new_G1172_ & new_G1803_;
  assign new_G2115_ = new_G1172_ & new_G1805_;
  assign new_G2116_ = n4371_lo & new_G825_ & new_G1847_;
  assign new_G2117_ = ~new_G1853_;
  assign new_G2118_ = n4395_lo & new_G825_ & new_G1849_;
  assign new_G2119_ = n4407_lo & new_G825_ & new_G1851_;
  assign new_G2120_ = new_G804_ & new_G1846_;
  assign new_G2121_ = new_G804_ & new_G1848_;
  assign new_G2122_ = new_G804_ & new_G1850_;
  assign new_G2123_ = new_G825_ & new_G1861_;
  assign new_G2124_ = n4347_lo & new_G825_ & new_G1863_;
  assign new_G2125_ = n4359_lo & new_G825_ & new_G1865_;
  assign new_G2126_ = new_G804_ & new_G1860_;
  assign new_G2127_ = new_G804_ & new_G1862_;
  assign new_G2128_ = new_G804_ & new_G1864_;
  assign new_G2129_ = new_G825_ & new_G1872_;
  assign new_G2130_ = new_G825_ & new_G1879_;
  assign new_G2131_ = n4323_lo & new_G813_ & new_G1889_;
  assign new_G2132_ = n4335_lo & new_G813_ & new_G1891_;
  assign new_G2133_ = n4287_lo & new_G813_ & new_G1893_;
  assign new_G2134_ = n4299_lo & new_G813_ & new_G1895_;
  assign new_G2135_ = new_G1172_ & new_G1888_;
  assign new_G2136_ = new_G1172_ & new_G1890_;
  assign new_G2137_ = new_G1172_ & new_G1892_;
  assign new_G2138_ = new_G1172_ & new_G1894_;
  assign new_G2139_ = ~new_G1410_ | ~new_G1904_;
  assign new_G2140_ = ~new_G1407_ | ~new_G1905_;
  assign new_G2141_ = ~new_G1416_ | ~new_G1906_;
  assign new_G2142_ = ~new_G1413_ | ~new_G1907_;
  assign new_G2143_ = ~new_G1434_ | ~new_G2014_;
  assign new_G2144_ = ~new_G1431_ | ~new_G2015_;
  assign new_G2145_ = ~new_G1440_ | ~new_G2016_;
  assign new_G2146_ = ~new_G1437_ | ~new_G2017_;
  assign new_G2147_ = ~new_G1446_ | ~new_G2018_;
  assign new_G2148_ = ~new_G1443_ | ~new_G2019_;
  assign new_G2149_ = ~new_G1422_ | ~new_G2067_;
  assign new_G2150_ = ~new_G1419_ | ~new_G2068_;
  assign new_G2151_ = ~new_G1428_ | ~new_G2069_;
  assign new_G2152_ = ~new_G1425_ | ~new_G2070_;
  assign new_G2153_ = ~new_G1452_ | ~new_G2071_;
  assign new_G2154_ = ~new_G1449_ | ~new_G2072_;
  assign new_G2155_ = new_G1755_ & new_G1764_;
  assign new_G2156_ = new_G983_ & new_G1764_;
  assign new_G2157_ = n3639_lo & new_G1526_ & new_G706_;
  assign new_G2158_ = n3651_lo & new_G1526_ & new_G706_;
  assign new_G2159_ = n3627_lo & new_G1526_ & new_G706_;
  assign new_G2160_ = n3615_lo & new_G1526_ & new_G706_;
  assign new_G2161_ = n3603_lo & new_G1526_ & new_G706_;
  assign new_G2162_ = n3567_lo & new_G1554_ & new_G730_;
  assign new_G2163_ = n3591_lo & new_G1554_ & new_G730_;
  assign new_G2164_ = n3459_lo & new_G1554_ & new_G730_;
  assign new_G2165_ = n3435_lo & new_G1554_ & new_G730_;
  assign new_G2166_ = new_G1755_ & new_G1764_;
  assign new_G2167_ = new_G983_ & new_G1764_;
  assign new_G2168_ = n3639_lo & new_G1601_ & new_G768_;
  assign new_G2169_ = n3651_lo & new_G1601_ & new_G768_;
  assign new_G2170_ = n3627_lo & new_G1601_ & new_G768_;
  assign new_G2171_ = n3615_lo & new_G1601_ & new_G768_;
  assign new_G2172_ = n3603_lo & new_G1601_ & new_G768_;
  assign new_G2173_ = n3567_lo & new_G1629_ & new_G792_;
  assign new_G2174_ = n3591_lo & new_G1629_ & new_G792_;
  assign new_G2175_ = n3459_lo & new_G1629_ & new_G792_;
  assign new_G2176_ = n3435_lo & new_G1629_ & new_G792_;
  assign new_G2177_ = new_G1755_ & new_G1764_;
  assign new_G2178_ = new_G983_ & new_G1764_;
  assign new_G2179_ = n3111_lo & new_G1948_ & new_G1230_;
  assign new_G2180_ = new_G1755_ & new_G1764_;
  assign new_G2181_ = new_G983_ & new_G1764_;
  assign new_G2182_ = n2643_lo & new_G1652_ & new_G872_;
  assign new_G2183_ = n3111_lo & new_G1914_ & new_G1196_;
  assign new_G2184_ = n2811_lo & new_G1914_ & new_G1196_;
  assign new_G2185_ = n3075_lo & new_G1914_ & new_G1196_;
  assign new_G2186_ = n3039_lo & new_G1914_ & new_G1196_;
  assign new_G2187_ = n2799_lo & new_G1914_ & new_G1196_;
  assign new_G2188_ = n2931_lo & new_G1652_ & new_G872_;
  assign new_G2189_ = n2919_lo & new_G1652_ & new_G872_;
  assign new_G2190_ = n2895_lo & new_G1652_ & new_G872_;
  assign new_G2191_ = n2655_lo & new_G1652_ & new_G872_;
  assign new_G2192_ = n2811_lo & new_G1948_ & new_G1230_;
  assign new_G2193_ = n3075_lo & new_G1948_ & new_G1230_;
  assign new_G2194_ = n3039_lo & new_G1948_ & new_G1230_;
  assign new_G2195_ = n2799_lo & new_G1948_ & new_G1230_;
  assign new_G2196_ = n2931_lo & new_G1674_ & new_G896_;
  assign new_G2197_ = n2919_lo & new_G1674_ & new_G896_;
  assign new_G2198_ = n2895_lo & new_G1674_ & new_G896_;
  assign new_G2199_ = n2655_lo & new_G1674_ & new_G896_;
  assign new_G2200_ = n3219_lo & new_G1992_ & new_G1272_;
  assign new_G2201_ = n2643_lo & new_G1674_ & new_G896_;
  assign new_G2202_ = n3195_lo & new_G1970_ & new_G1256_;
  assign new_G2203_ = n3543_lo & new_G1554_ & new_G730_;
  assign new_G2204_ = n3543_lo & new_G1629_ & new_G792_;
  assign new_G2205_ = new_G1704_ | new_G2077_;
  assign new_G2206_ = new_G1705_ | new_G2078_;
  assign new_G2207_ = new_G1706_ | new_G2079_;
  assign new_G2208_ = new_G1707_ | new_G2080_;
  assign new_G2209_ = n4323_lo | new_G1708_ | new_G2081_;
  assign new_G2210_ = n4335_lo | new_G1709_ | new_G2082_;
  assign new_G2211_ = n4287_lo | new_G1710_ | new_G2083_;
  assign new_G2212_ = n4299_lo | new_G1711_ | new_G2084_;
  assign new_G2213_ = new_G1720_ | new_G2085_;
  assign new_G2214_ = new_G1721_ | new_G2086_;
  assign new_G2215_ = new_G1722_ | new_G2087_;
  assign new_G2216_ = new_G1723_ | new_G2088_;
  assign new_G2217_ = n4251_lo | new_G1724_ | new_G2089_;
  assign new_G2218_ = n4263_lo | new_G1725_ | new_G2090_;
  assign new_G2219_ = n4275_lo | new_G1726_ | new_G2091_;
  assign new_G2220_ = n4227_lo | new_G1727_ | new_G2092_;
  assign new_G2221_ = n3939_lo & new_G1728_;
  assign new_G2222_ = n3915_lo & new_G1728_;
  assign new_G2223_ = n3891_lo & new_G1728_;
  assign new_G2224_ = n3867_lo & new_G1728_;
  assign new_G2225_ = n3843_lo & new_G1728_;
  assign new_G2226_ = n3759_lo & new_G1734_;
  assign new_G2227_ = n3735_lo & new_G1734_;
  assign new_G2228_ = n3711_lo & new_G1734_;
  assign new_G2229_ = n3687_lo & new_G1734_;
  assign new_G2230_ = n3663_lo & new_G1734_;
  assign new_G2231_ = ~new_G1764_;
  assign new_G2240_ = new_G1780_ | new_G2093_;
  assign new_G2241_ = new_G1781_ | new_G2094_;
  assign new_G2242_ = new_G1782_ | new_G2095_;
  assign new_G2243_ = n4347_lo | new_G1784_ | new_G2097_;
  assign new_G2244_ = n4359_lo | new_G1785_ | new_G2098_;
  assign new_G2245_ = new_G1783_ | new_G2096_;
  assign new_G2248_ = new_G1792_ | new_G2099_;
  assign new_G2249_ = new_G1794_ | new_G2100_;
  assign new_G2250_ = new_G1795_ | new_G2101_;
  assign new_G2251_ = n4371_lo | new_G1796_ | new_G2102_;
  assign new_G2252_ = n4395_lo | new_G1797_ | new_G2103_;
  assign new_G2253_ = n4407_lo | new_G1798_ | new_G2104_;
  assign new_G2254_ = new_G1807_ | new_G2108_;
  assign new_G2255_ = new_G1808_ | new_G2109_;
  assign new_G2256_ = new_G1809_ | new_G2110_;
  assign new_G2257_ = new_G1810_ | new_G2111_;
  assign new_G2258_ = n4251_lo | new_G1811_ | new_G2112_;
  assign new_G2259_ = n4263_lo | new_G1812_ | new_G2113_;
  assign new_G2260_ = n4275_lo | new_G1813_ | new_G2114_;
  assign new_G2261_ = n4227_lo | new_G1814_ | new_G2115_;
  assign new_G2262_ = n4191_lo & new_G1815_;
  assign new_G2263_ = n4167_lo & new_G1815_;
  assign new_G2264_ = n4143_lo & new_G1815_;
  assign new_G2265_ = n4119_lo & new_G1815_;
  assign new_G2266_ = n4059_lo & new_G1821_;
  assign new_G2267_ = n4035_lo & new_G1821_;
  assign new_G2268_ = n4011_lo & new_G1821_;
  assign new_G2269_ = n3987_lo & new_G1821_;
  assign new_G2270_ = n3963_lo & new_G1821_;
  assign new_G2271_ = new_G1815_ | new_G1831_;
  assign new_G2277_ = n2991_lo & new_G1837_;
  assign new_G2278_ = n3015_lo & new_G1837_;
  assign new_G2279_ = n2763_lo & new_G1837_;
  assign new_G2280_ = n2763_lo & new_G1837_;
  assign new_G2281_ = new_G1852_ | new_G2116_;
  assign new_G2282_ = new_G1854_ | new_G2118_;
  assign new_G2283_ = new_G1855_ | new_G2119_;
  assign new_G2284_ = n4371_lo | new_G1856_ | new_G2120_;
  assign new_G2285_ = n4395_lo | new_G1858_ | new_G2121_;
  assign new_G2286_ = n4407_lo | new_G1859_ | new_G2122_;
  assign new_G2287_ = new_G1866_ | new_G2123_;
  assign new_G2288_ = new_G1867_ | new_G2124_;
  assign new_G2289_ = new_G1868_ | new_G2125_;
  assign new_G2290_ = n4347_lo | new_G1870_ | new_G2127_;
  assign new_G2291_ = n4359_lo | new_G1871_ | new_G2128_;
  assign new_G2292_ = ~new_G1873_;
  assign new_G2293_ = ~new_G1876_;
  assign new_G2294_ = ~new_G1880_;
  assign new_G2295_ = ~new_G1883_;
  assign new_G2296_ = new_G1886_ | new_G2129_;
  assign new_G2297_ = new_G848_ & n4311_lo & new_G1876_;
  assign new_G2298_ = new_G1887_ | new_G2130_;
  assign new_G2299_ = new_G848_ & n4311_lo & new_G1883_;
  assign new_G2300_ = new_G1162_ & new_G1873_;
  assign new_G2301_ = new_G1162_ & new_G1880_;
  assign new_G2302_ = new_G1896_ | new_G2131_;
  assign new_G2303_ = new_G1897_ | new_G2132_;
  assign new_G2304_ = new_G1898_ | new_G2133_;
  assign new_G2305_ = new_G1899_ | new_G2134_;
  assign new_G2306_ = n4323_lo | new_G1900_ | new_G2135_;
  assign new_G2307_ = n4335_lo | new_G1901_ | new_G2136_;
  assign new_G2308_ = n4287_lo | new_G1902_ | new_G2137_;
  assign new_G2309_ = n4299_lo | new_G1903_ | new_G2138_;
  assign new_G2310_ = ~new_G2139_ | ~new_G2140_;
  assign new_G2314_ = ~new_G2141_ | ~new_G2142_;
  assign new_G2318_ = ~new_G1908_;
  assign new_G2319_ = ~new_G1911_;
  assign new_G2320_ = n3183_lo & new_G1970_ & new_G1256_;
  assign new_G2321_ = n3267_lo & new_G1970_ & new_G1256_;
  assign new_G2322_ = n3279_lo & new_G1970_ & new_G1256_;
  assign new_G2323_ = n3291_lo & new_G1970_ & new_G1256_;
  assign new_G2324_ = n3327_lo & new_G1992_ & new_G1272_;
  assign new_G2325_ = n3303_lo & new_G1992_ & new_G1272_;
  assign new_G2326_ = n3207_lo & new_G1992_ & new_G1272_;
  assign new_G2327_ = n3315_lo & new_G1992_ & new_G1272_;
  assign new_G2328_ = ~new_G2143_ | ~new_G2144_;
  assign new_G2332_ = ~new_G2145_ | ~new_G2146_;
  assign new_G2336_ = ~new_G2147_ | ~new_G2148_;
  assign new_G2339_ = n3243_lo & new_G2020_ & new_G1287_;
  assign new_G2340_ = n3135_lo & new_G2020_ & new_G1287_;
  assign new_G2341_ = n2847_lo & new_G2020_ & new_G1287_;
  assign new_G2342_ = n3147_lo & new_G2020_ & new_G1287_;
  assign new_G2343_ = n3159_lo & new_G2020_ & new_G1287_;
  assign new_G2344_ = n2835_lo & new_G2042_ & new_G1301_;
  assign new_G2345_ = n3123_lo & new_G2042_ & new_G1301_;
  assign new_G2346_ = n3171_lo & new_G2042_ & new_G1301_;
  assign new_G2347_ = n3231_lo & new_G2042_ & new_G1301_;
  assign new_G2348_ = n3255_lo & new_G2042_ & new_G1301_;
  assign new_G2349_ = ~new_G2151_ | ~new_G2152_;
  assign new_G2352_ = ~new_G2149_ | ~new_G2150_;
  assign new_G2355_ = new_G2117_ & new_G1857_;
  assign new_G2358_ = new_G1869_ | new_G2126_;
  assign new_G2361_ = ~new_G2073_;
  assign new_G2362_ = ~new_G2073_ | ~new_G2076_;
  assign new_G2363_ = ~new_G2153_ | ~new_G2154_;
  assign new_G2366_ = ~new_G2105_;
  assign new_G2367_ = new_G2278_ | new_G1843_;
  assign new_G2368_ = new_G2279_ | new_G1844_;
  assign new_G2369_ = new_G2280_ | new_G1845_;
  assign new_G2370_ = new_G2277_ | new_G1842_;
  assign new_G2371_ = ~new_G2205_;
  assign new_G2372_ = ~new_G2206_;
  assign new_G2373_ = ~new_G2207_;
  assign new_G2374_ = ~new_G2208_;
  assign new_G2375_ = ~new_G2213_;
  assign new_G2376_ = ~new_G2214_;
  assign new_G2377_ = ~new_G2215_;
  assign new_G2378_ = ~new_G2216_;
  assign new_G2379_ = new_G2222_ | new_G1741_;
  assign new_G2386_ = new_G2223_ | new_G1742_;
  assign new_G2392_ = new_G2224_ | new_G1743_;
  assign new_G2398_ = new_G2225_ | new_G1744_;
  assign new_G2404_ = new_G2226_ | new_G1745_;
  assign new_G2410_ = new_G2227_ | new_G1746_;
  assign new_G2418_ = new_G2228_ | new_G1747_;
  assign new_G2424_ = new_G2229_ | new_G1748_;
  assign new_G2430_ = new_G2230_ | new_G1749_;
  assign new_G2436_ = ~new_G2241_;
  assign new_G2437_ = ~new_G2242_;
  assign new_G2438_ = ~new_G2240_;
  assign new_G2441_ = ~new_G2248_;
  assign new_G2442_ = ~new_G2249_;
  assign new_G2443_ = ~new_G2250_;
  assign new_G2444_ = ~new_G2254_;
  assign new_G2445_ = ~new_G2255_;
  assign new_G2446_ = ~new_G2256_;
  assign new_G2447_ = ~new_G2257_;
  assign new_G2448_ = new_G2263_ | new_G1828_;
  assign new_G2454_ = new_G2264_ | new_G1829_;
  assign new_G2460_ = new_G2265_ | new_G1830_;
  assign new_G2466_ = new_G2266_ | new_G1832_;
  assign new_G2472_ = new_G2267_ | new_G1833_;
  assign new_G2480_ = new_G2268_ | new_G1834_;
  assign new_G2486_ = new_G2269_ | new_G1835_;
  assign new_G2492_ = new_G2270_ | new_G1836_;
  assign new_G2499_ = ~new_G2281_;
  assign new_G2500_ = ~new_G2282_;
  assign new_G2501_ = ~new_G2283_;
  assign new_G2502_ = ~new_G2288_;
  assign new_G2503_ = ~new_G2289_;
  assign new_G2504_ = n4311_lo & new_G825_ & new_G2293_;
  assign new_G2505_ = n4311_lo & new_G825_ & new_G2295_;
  assign new_G2506_ = new_G804_ & new_G2292_;
  assign new_G2507_ = new_G804_ & new_G2294_;
  assign new_G2508_ = ~new_G2296_;
  assign new_G2511_ = ~new_G2298_;
  assign new_G2512_ = ~new_G2302_;
  assign new_G2513_ = ~new_G2303_;
  assign new_G2514_ = ~new_G2304_;
  assign new_G2515_ = ~new_G2305_;
  assign new_G2516_ = new_G2105_ & new_G1992_ & new_G2003_;
  assign new_G2517_ = new_G2262_ | new_G1827_;
  assign new_G2520_ = new_G2221_ | new_G1740_;
  assign new_G2523_ = ~new_G2287_;
  assign new_G2526_ = ~new_G1455_ | ~new_G2361_;
  assign new_G2527_ = ~new_G2245_;
  assign new_G2528_ = new_G2367_ & new_G1070_;
  assign new_G2529_ = n2703_lo & new_G1755_ & new_G2231_;
  assign new_G2530_ = n2715_lo & new_G983_ & new_G2231_;
  assign new_G2531_ = n2727_lo & new_G1755_ & new_G2231_;
  assign new_G2532_ = n2967_lo & new_G983_ & new_G2231_;
  assign new_G2533_ = new_G2368_ & new_G1070_;
  assign new_G2534_ = n2943_lo & new_G1755_ & new_G2231_;
  assign new_G2535_ = n2691_lo & new_G983_ & new_G2231_;
  assign new_G2536_ = n2979_lo & new_G1755_ & new_G2231_;
  assign new_G2537_ = n2955_lo & new_G983_ & new_G2231_;
  assign new_G2538_ = new_G2369_ & new_G1070_;
  assign new_G2539_ = new_G2370_ & new_G1070_;
  assign new_G2540_ = new_G2271_ & n4383_lo;
  assign new_G2543_ = n4383_lo & new_G2271_;
  assign new_G2547_ = new_G2371_ & new_G2209_;
  assign new_G2550_ = new_G2372_ & new_G2210_;
  assign new_G2553_ = new_G2373_ & new_G2211_;
  assign new_G2556_ = new_G2374_ & new_G2212_;
  assign new_G2559_ = new_G2375_ & new_G2217_;
  assign new_G2562_ = new_G2376_ & new_G2218_;
  assign new_G2565_ = new_G2377_ & new_G2219_;
  assign new_G2568_ = new_G2378_ & new_G2220_;
  assign new_G2571_ = new_G2436_ & new_G2243_;
  assign new_G2574_ = new_G2437_ & new_G2244_;
  assign new_G2577_ = ~new_G2245_;
  assign new_G2580_ = new_G2441_ & new_G2251_;
  assign new_G2583_ = new_G2442_ & new_G2252_;
  assign new_G2586_ = new_G2443_ & new_G2253_;
  assign new_G2589_ = new_G2297_ | new_G2504_;
  assign new_G2590_ = new_G2299_ | new_G2505_;
  assign new_G2591_ = n4311_lo | new_G2300_ | new_G2506_;
  assign new_G2592_ = n4311_lo | new_G2301_ | new_G2507_;
  assign new_G2593_ = ~new_G2310_;
  assign new_G2596_ = ~new_G2314_;
  assign new_G2599_ = new_G2314_ & new_G2310_ & new_G1908_;
  assign new_G2600_ = new_G2511_ & new_G1992_ & new_G2003_;
  assign new_G2601_ = new_G2447_ & new_G2261_;
  assign new_G2602_ = ~new_G2355_;
  assign new_G2603_ = ~new_G2328_;
  assign new_G2606_ = ~new_G2332_;
  assign new_G2609_ = ~new_G2336_;
  assign new_G2612_ = ~new_G2336_;
  assign new_G2615_ = ~new_G2271_;
  assign new_G2618_ = ~new_G2271_;
  assign new_G2621_ = ~new_G2271_;
  assign new_G2624_ = ~new_G2349_;
  assign new_G2625_ = ~new_G2352_;
  assign new_G2626_ = new_G2445_ & new_G2259_;
  assign new_G2629_ = new_G2446_ & new_G2260_;
  assign new_G2632_ = new_G2515_ & new_G2309_;
  assign new_G2635_ = new_G2444_ & new_G2258_;
  assign new_G2638_ = new_G2513_ & new_G2307_;
  assign new_G2641_ = new_G2514_ & new_G2308_;
  assign new_G2644_ = new_G2512_ & new_G2306_;
  assign new_G2647_ = new_G2500_ & new_G2285_;
  assign new_G2650_ = new_G2501_ & new_G2286_;
  assign new_G2653_ = new_G2499_ & new_G2284_;
  assign new_G2656_ = new_G2502_ & new_G2290_;
  assign new_G2659_ = new_G2503_ & new_G2291_;
  assign new_G2662_ = ~new_G2358_;
  assign new_G2663_ = ~new_G2526_ | ~new_G2362_;
  assign new_G2666_ = ~new_G2363_;
  assign new_G2667_ = n4311_lo & new_G2430_;
  assign new_G2668_ = ~new_G2438_;
  assign new_G2669_ = ~new_G2508_;
  assign new_G2670_ = new_G2430_ & n4311_lo;
  assign new_G2671_ = new_G2156_ | new_G2155_ | new_G2529_ | new_G2530_;
  assign new_G2672_ = new_G2167_ | new_G2166_ | new_G2531_ | new_G2532_;
  assign new_G2673_ = new_G2178_ | new_G2177_ | new_G2534_ | new_G2535_;
  assign new_G2674_ = new_G2181_ | new_G2180_ | new_G2536_ | new_G2537_;
  assign new_G2675_ = new_G2424_ & n4323_lo;
  assign new_G2679_ = new_G2418_ & n4335_lo;
  assign new_G2685_ = n4287_lo & new_G2410_;
  assign new_G2692_ = new_G2404_ & n4299_lo;
  assign new_G2693_ = new_G2398_ & n4251_lo;
  assign new_G2696_ = new_G2392_ & n4263_lo;
  assign new_G2700_ = new_G2386_ & n4275_lo;
  assign new_G2705_ = new_G2379_ & n4227_lo;
  assign new_G2711_ = n4323_lo & new_G2424_;
  assign new_G2715_ = n4335_lo & new_G2418_;
  assign new_G2720_ = n4287_lo & new_G2410_;
  assign new_G2726_ = n4299_lo & new_G2404_;
  assign new_G2727_ = n4251_lo & new_G2398_;
  assign new_G2731_ = n4263_lo & new_G2392_;
  assign new_G2737_ = n4275_lo & new_G2386_;
  assign new_G2744_ = n4227_lo & new_G2379_;
  assign new_G2752_ = ~new_G2492_;
  assign new_G2759_ = ~new_G2486_;
  assign new_G2770_ = ~new_G2486_;
  assign new_G2774_ = new_G2480_ & n4347_lo;
  assign new_G2780_ = n4359_lo & new_G2472_;
  assign new_G2787_ = new_G2466_ & n4371_lo;
  assign new_G2788_ = new_G2460_ & n4395_lo;
  assign new_G2792_ = new_G2454_ & n4407_lo;
  assign new_G2797_ = ~new_G2448_;
  assign new_G2804_ = ~new_G2448_;
  assign new_G2810_ = ~new_G2492_;
  assign new_G2817_ = ~new_G2486_;
  assign new_G2828_ = ~new_G2486_;
  assign new_G2832_ = n4347_lo & new_G2480_;
  assign new_G2837_ = n4359_lo & new_G2472_;
  assign new_G2843_ = n4371_lo & new_G2466_;
  assign new_G2844_ = n4395_lo & new_G2460_;
  assign new_G2850_ = n4407_lo & new_G2454_;
  assign new_G2857_ = ~new_G2448_;
  assign new_G2865_ = ~new_G2448_;
  assign new_G2872_ = ~new_G2492_;
  assign new_G2875_ = ~new_G2589_;
  assign new_G2876_ = ~new_G2590_;
  assign new_G2877_ = ~new_G2517_;
  assign new_G2878_ = ~new_G2520_;
  assign new_G2879_ = ~new_G2601_;
  assign new_G2883_ = ~new_G2508_;
  assign new_G2887_ = new_G2438_ & new_G2042_ & new_G2053_;
  assign new_G2888_ = ~new_G2430_;
  assign new_G2891_ = ~new_G2424_;
  assign new_G2894_ = ~new_G2418_;
  assign new_G2897_ = ~new_G2410_;
  assign new_G2900_ = ~new_G2404_;
  assign new_G2903_ = ~new_G2398_;
  assign new_G2906_ = ~new_G2392_;
  assign new_G2909_ = ~new_G2386_;
  assign new_G2912_ = ~new_G2379_;
  assign new_G2915_ = ~n4287_lo & ~new_G2410_;
  assign new_G2918_ = ~new_G2430_;
  assign new_G2921_ = ~new_G2424_;
  assign new_G2924_ = ~new_G2418_;
  assign new_G2927_ = ~new_G2404_;
  assign new_G2930_ = ~new_G2398_;
  assign new_G2933_ = ~new_G2392_;
  assign new_G2936_ = ~new_G2386_;
  assign new_G2939_ = ~new_G2410_;
  assign new_G2942_ = ~new_G2379_;
  assign new_G2945_ = ~n4287_lo & ~new_G2410_;
  assign new_G2948_ = ~n4227_lo & ~new_G2379_;
  assign new_G2951_ = ~new_G2480_;
  assign new_G2954_ = ~new_G2472_;
  assign new_G2957_ = ~new_G2466_;
  assign new_G2960_ = ~new_G2460_;
  assign new_G2963_ = ~new_G2454_;
  assign new_G2966_ = ~n4359_lo & ~new_G2472_;
  assign new_G2969_ = ~new_G2480_;
  assign new_G2972_ = ~new_G2466_;
  assign new_G2975_ = ~new_G2460_;
  assign new_G2978_ = ~new_G2454_;
  assign new_G2981_ = ~new_G2472_;
  assign new_G2984_ = ~n4359_lo & ~new_G2472_;
  assign new_G2987_ = ~new_G2454_;
  assign new_G2990_ = ~new_G2460_;
  assign new_G2993_ = ~new_G2448_;
  assign new_G2996_ = ~new_G2466_;
  assign new_G2999_ = ~new_G2480_;
  assign new_G3002_ = ~new_G2472_;
  assign new_G3005_ = ~new_G2492_;
  assign new_G3008_ = ~new_G2486_;
  assign new_G3011_ = ~new_G2410_;
  assign new_G3014_ = ~new_G2404_;
  assign new_G3017_ = ~new_G2424_;
  assign new_G3020_ = ~new_G2418_;
  assign new_G3023_ = ~new_G2430_;
  assign new_G3026_ = ~new_G2386_;
  assign new_G3029_ = ~new_G2379_;
  assign new_G3032_ = ~new_G2398_;
  assign new_G3035_ = ~new_G2392_;
  assign new_G3038_ = ~new_G2352_ | ~new_G2624_;
  assign new_G3039_ = ~new_G2349_ | ~new_G2625_;
  assign new_G3040_ = ~new_G2523_;
  assign new_G3041_ = ~new_G2523_ | ~new_G2662_;
  assign new_G3042_ = ~new_G2574_;
  assign new_G3043_ = ~new_G2571_;
  assign new_G3044_ = ~new_G2586_;
  assign new_G3045_ = ~new_G2583_;
  assign new_G3046_ = ~new_G2580_;
  assign new_G3047_ = ~new_G2556_;
  assign new_G3048_ = ~new_G2553_;
  assign new_G3049_ = ~new_G2550_;
  assign new_G3050_ = ~new_G2547_;
  assign new_G3051_ = ~new_G2568_;
  assign new_G3052_ = ~new_G2565_;
  assign new_G3053_ = ~new_G2562_;
  assign new_G3054_ = ~new_G2559_;
  assign new_G3055_ = new_G2577_ & new_G1245_ & new_G1242_;
  assign new_G3056_ = ~new_G2615_;
  assign new_G3057_ = ~new_G2615_ | ~new_G1585_;
  assign new_G3058_ = ~new_G2618_ | ~new_G1591_;
  assign new_G3059_ = ~new_G2618_;
  assign new_G3060_ = new_G2875_ & new_G2591_;
  assign new_G3063_ = new_G2876_ & new_G2592_;
  assign new_G3064_ = ~new_G2621_;
  assign new_G3065_ = new_G2593_ & new_G2314_ & new_G2318_;
  assign new_G3066_ = new_G2310_ & new_G2596_ & new_G2319_;
  assign new_G3067_ = new_G2596_ & new_G2593_ & new_G1911_;
  assign new_G3068_ = new_G2568_ & new_G1970_ & new_G1981_;
  assign new_G3069_ = new_G2565_ & new_G1970_ & new_G1981_;
  assign new_G3070_ = new_G2562_ & new_G1970_ & new_G1981_;
  assign new_G3071_ = new_G2559_ & new_G1970_ & new_G1981_;
  assign new_G3072_ = new_G2586_ & new_G1992_ & new_G2003_;
  assign new_G3073_ = new_G2583_ & new_G1992_ & new_G2003_;
  assign new_G3074_ = ~new_G2626_;
  assign new_G3075_ = ~new_G2629_;
  assign new_G3076_ = ~new_G2632_;
  assign new_G3077_ = ~new_G2635_;
  assign new_G3078_ = ~new_G2647_;
  assign new_G3079_ = ~new_G2650_;
  assign new_G3080_ = ~new_G2653_;
  assign new_G3081_ = ~new_G2653_ | ~new_G2602_;
  assign new_G3082_ = ~new_G2609_;
  assign new_G3083_ = ~new_G2612_;
  assign new_G3084_ = new_G2332_ & new_G2328_ & new_G2609_;
  assign new_G3085_ = new_G2606_ & new_G2603_ & new_G2612_;
  assign new_G3086_ = new_G2556_ & new_G2020_ & new_G2031_;
  assign new_G3087_ = new_G2553_ & new_G2020_ & new_G2031_;
  assign new_G3088_ = new_G2550_ & new_G2020_ & new_G2031_;
  assign new_G3089_ = new_G2547_ & new_G2020_ & new_G2031_;
  assign new_G3090_ = new_G2580_ & new_G2042_ & new_G2053_;
  assign new_G3091_ = new_G2574_ & new_G2042_ & new_G2053_;
  assign new_G3092_ = new_G2571_ & new_G2042_ & new_G2053_;
  assign new_G3093_ = new_G2577_ & new_G2042_ & new_G2053_;
  assign new_G3094_ = ~new_G3038_ | ~new_G3039_;
  assign new_G3097_ = ~new_G2638_;
  assign new_G3098_ = ~new_G2641_;
  assign new_G3099_ = ~new_G2644_;
  assign new_G3100_ = ~new_G2656_;
  assign new_G3101_ = ~new_G2659_;
  assign new_G3102_ = ~new_G2358_ | ~new_G3040_;
  assign new_G3103_ = ~new_G2663_;
  assign new_G3104_ = ~new_G2663_ | ~new_G2666_;
  assign new_G3105_ = new_G2527_ & new_G3042_ & new_G3043_ & new_G2668_;
  assign new_G3106_ = new_G3046_ & new_G3044_ & new_G3045_ & new_G2366_;
  assign new_G3107_ = new_G3050_ & new_G3047_ & new_G3048_ & new_G3049_;
  assign new_G3108_ = new_G3054_ & new_G3051_ & new_G3052_ & new_G3053_;
  assign new_G3109_ = new_G2752_ & new_G2770_;
  assign new_G3110_ = new_G2759_ & new_G2752_ & new_G2774_;
  assign new_G3111_ = new_G2810_ & new_G2828_;
  assign new_G3112_ = new_G2817_ & new_G2810_ & new_G2832_;
  assign new_G3113_ = ~new_G2888_;
  assign new_G3114_ = ~new_G2888_ | ~new_G1501_;
  assign new_G3115_ = ~new_G2891_;
  assign new_G3116_ = ~new_G2891_ | ~new_G1502_;
  assign new_G3117_ = ~new_G2894_;
  assign new_G3118_ = ~new_G2894_ | ~new_G1503_;
  assign new_G3119_ = ~new_G2897_;
  assign new_G3120_ = ~new_G2897_ | ~new_G1504_;
  assign new_G3121_ = ~new_G2900_;
  assign new_G3122_ = ~new_G2900_ | ~new_G1505_;
  assign new_G3123_ = ~new_G2903_;
  assign new_G3124_ = ~new_G2903_ | ~new_G1506_;
  assign new_G3125_ = ~new_G2906_;
  assign new_G3126_ = ~new_G2906_ | ~new_G1507_;
  assign new_G3127_ = ~new_G2909_;
  assign new_G3128_ = ~new_G2909_ | ~new_G1508_;
  assign new_G3129_ = ~new_G2912_;
  assign new_G3130_ = ~new_G2912_ | ~new_G1509_;
  assign new_G3131_ = ~new_G2915_;
  assign new_G3132_ = ~new_G2918_ | ~new_G1511_;
  assign new_G3133_ = ~new_G2918_;
  assign new_G3134_ = ~new_G2921_ | ~new_G1512_;
  assign new_G3135_ = ~new_G2921_;
  assign new_G3136_ = ~new_G2924_ | ~new_G1513_;
  assign new_G3137_ = ~new_G2924_;
  assign new_G3138_ = ~new_G2927_ | ~new_G1514_;
  assign new_G3139_ = ~new_G2927_;
  assign new_G3140_ = ~new_G2930_ | ~new_G1515_;
  assign new_G3141_ = ~new_G2930_;
  assign new_G3142_ = ~new_G2933_ | ~new_G1516_;
  assign new_G3143_ = ~new_G2933_;
  assign new_G3144_ = ~new_G2936_ | ~new_G1517_;
  assign new_G3145_ = ~new_G2936_;
  assign new_G3146_ = ~new_G2939_ | ~new_G1518_;
  assign new_G3147_ = ~new_G2939_;
  assign new_G3148_ = ~new_G2942_ | ~new_G1519_;
  assign new_G3149_ = ~new_G2942_;
  assign new_G3150_ = ~new_G2951_;
  assign new_G3151_ = ~new_G2951_ | ~new_G1582_;
  assign new_G3152_ = ~new_G2954_;
  assign new_G3153_ = ~new_G2954_ | ~new_G1583_;
  assign new_G3154_ = ~new_G2957_;
  assign new_G3155_ = ~new_G2957_ | ~new_G1584_;
  assign new_G3156_ = ~new_G1377_ | ~new_G3056_;
  assign new_G3157_ = ~new_G2960_;
  assign new_G3158_ = ~new_G2960_ | ~new_G1586_;
  assign new_G3159_ = ~new_G2963_;
  assign new_G3160_ = ~new_G2963_ | ~new_G1587_;
  assign new_G3161_ = new_G2759_ & new_G2774_;
  assign new_G3162_ = new_G2759_ & new_G2774_;
  assign new_G3163_ = n2859_lo & new_G2797_;
  assign new_G3164_ = ~new_G2966_;
  assign new_G3165_ = ~new_G2969_ | ~new_G1589_;
  assign new_G3166_ = ~new_G2969_;
  assign new_G3167_ = ~new_G2972_ | ~new_G1590_;
  assign new_G3168_ = ~new_G2972_;
  assign new_G3169_ = ~new_G1395_ | ~new_G3059_;
  assign new_G3170_ = ~new_G2975_ | ~new_G1592_;
  assign new_G3171_ = ~new_G2975_;
  assign new_G3172_ = ~new_G2978_ | ~new_G1593_;
  assign new_G3173_ = ~new_G2978_;
  assign new_G3174_ = ~new_G2981_ | ~new_G1594_;
  assign new_G3175_ = ~new_G2981_;
  assign new_G3176_ = new_G2817_ & new_G2832_;
  assign new_G3177_ = new_G2817_ & new_G2832_;
  assign new_G3178_ = ~new_G2987_;
  assign new_G3179_ = ~new_G2990_;
  assign new_G3180_ = ~new_G2993_ | ~new_G2877_;
  assign new_G3181_ = ~new_G2993_;
  assign new_G3182_ = ~new_G2996_;
  assign new_G3183_ = ~new_G2996_ | ~new_G3064_;
  assign new_G3184_ = ~new_G3011_;
  assign new_G3185_ = ~new_G3014_;
  assign new_G3186_ = ~new_G3017_;
  assign new_G3187_ = ~new_G3020_;
  assign new_G3188_ = ~new_G3023_ | ~new_G2878_;
  assign new_G3189_ = ~new_G3023_;
  assign new_G3190_ = ~new_G3065_ & ~new_G2599_;
  assign new_G3191_ = ~new_G3066_ & ~new_G3067_;
  assign new_G3192_ = ~new_G2879_;
  assign new_G3195_ = ~new_G2629_ | ~new_G3074_;
  assign new_G3196_ = ~new_G2626_ | ~new_G3075_;
  assign new_G3197_ = ~new_G2635_ | ~new_G3076_;
  assign new_G3198_ = ~new_G2632_ | ~new_G3077_;
  assign new_G3199_ = ~new_G2883_;
  assign new_G3202_ = ~new_G2650_ | ~new_G3078_;
  assign new_G3203_ = ~new_G2647_ | ~new_G3079_;
  assign new_G3204_ = ~new_G2355_ | ~new_G3080_;
  assign new_G3205_ = new_G2603_ & new_G2332_ & new_G3082_;
  assign new_G3206_ = new_G2328_ & new_G2606_ & new_G3083_;
  assign new_G3207_ = new_G3063_ & new_G2020_ & new_G2031_;
  assign new_G3208_ = ~new_G2872_;
  assign new_G3211_ = ~new_G2685_;
  assign new_G3214_ = ~new_G2945_;
  assign new_G3215_ = ~new_G2720_;
  assign new_G3218_ = ~new_G2948_;
  assign new_G3219_ = ~new_G2744_;
  assign new_G3222_ = ~new_G2797_;
  assign new_G3225_ = ~new_G2752_;
  assign new_G3228_ = ~new_G2752_;
  assign new_G3231_ = ~new_G2759_;
  assign new_G3234_ = ~new_G2759_;
  assign new_G3237_ = ~new_G2780_;
  assign new_G3240_ = ~new_G2984_;
  assign new_G3241_ = ~new_G2810_;
  assign new_G3244_ = ~new_G2817_;
  assign new_G3247_ = ~new_G2837_;
  assign new_G3250_ = ~new_G2810_;
  assign new_G3253_ = ~new_G2817_;
  assign new_G3256_ = ~new_G2865_;
  assign new_G3259_ = ~new_G2857_;
  assign new_G3262_ = ~new_G2865_;
  assign new_G3265_ = ~new_G2999_;
  assign new_G3266_ = ~new_G3002_;
  assign new_G3267_ = ~new_G3005_;
  assign new_G3268_ = ~new_G3008_;
  assign new_G3269_ = ~new_G3026_;
  assign new_G3270_ = ~new_G3029_;
  assign new_G3271_ = ~new_G3032_;
  assign new_G3272_ = ~new_G3035_;
  assign new_G3273_ = ~new_G2641_ | ~new_G3097_;
  assign new_G3274_ = ~new_G2638_ | ~new_G3098_;
  assign new_G3275_ = ~new_G2659_ | ~new_G3100_;
  assign new_G3276_ = ~new_G2656_ | ~new_G3101_;
  assign new_G3277_ = ~new_G3041_ | ~new_G3102_;
  assign new_G3280_ = ~new_G2363_ | ~new_G3103_;
  assign new_G3281_ = ~new_G3060_;
  assign new_G3282_ = ~new_G1311_ | ~new_G3113_;
  assign new_G3283_ = ~new_G1314_ | ~new_G3115_;
  assign new_G3284_ = ~new_G1317_ | ~new_G3117_;
  assign new_G3285_ = ~new_G1320_ | ~new_G3119_;
  assign new_G3286_ = ~new_G1323_ | ~new_G3121_;
  assign new_G3287_ = ~new_G1326_ | ~new_G3123_;
  assign new_G3288_ = ~new_G1329_ | ~new_G3125_;
  assign new_G3289_ = ~new_G1332_ | ~new_G3127_;
  assign new_G3290_ = ~new_G1335_ | ~new_G3129_;
  assign new_G3291_ = ~new_G1341_ | ~new_G3133_;
  assign new_G3292_ = ~new_G1344_ | ~new_G3135_;
  assign new_G3293_ = ~new_G1347_ | ~new_G3137_;
  assign new_G3294_ = ~new_G1350_ | ~new_G3139_;
  assign new_G3295_ = ~new_G1353_ | ~new_G3141_;
  assign new_G3296_ = ~new_G1356_ | ~new_G3143_;
  assign new_G3297_ = ~new_G1359_ | ~new_G3145_;
  assign new_G3298_ = ~new_G1362_ | ~new_G3147_;
  assign new_G3299_ = ~new_G1365_ | ~new_G3149_;
  assign new_G3300_ = ~new_G1368_ | ~new_G3150_;
  assign new_G3301_ = ~new_G1371_ | ~new_G3152_;
  assign new_G3302_ = ~new_G1374_ | ~new_G3154_;
  assign new_G3303_ = ~new_G3156_ | ~new_G3057_;
  assign new_G3313_ = ~new_G1380_ | ~new_G3157_;
  assign new_G3314_ = ~new_G1383_ | ~new_G3159_;
  assign new_G3315_ = ~new_G1389_ | ~new_G3166_;
  assign new_G3316_ = ~new_G1392_ | ~new_G3168_;
  assign new_G3317_ = ~new_G3058_ | ~new_G3169_;
  assign new_G3331_ = ~new_G1398_ | ~new_G3171_;
  assign new_G3332_ = ~new_G1401_ | ~new_G3173_;
  assign new_G3333_ = ~new_G1404_ | ~new_G3175_;
  assign new_G3334_ = ~new_G2990_ | ~new_G3178_;
  assign new_G3335_ = ~new_G2987_ | ~new_G3179_;
  assign new_G3336_ = ~new_G2517_ | ~new_G3181_;
  assign new_G3337_ = ~new_G2621_ | ~new_G3182_;
  assign new_G3338_ = ~new_G3014_ | ~new_G3184_;
  assign new_G3339_ = ~new_G3011_ | ~new_G3185_;
  assign new_G3340_ = ~new_G3020_ | ~new_G3186_;
  assign new_G3341_ = ~new_G3017_ | ~new_G3187_;
  assign new_G3342_ = ~new_G2520_ | ~new_G3189_;
  assign new_G3343_ = ~new_G3094_;
  assign new_G3344_ = ~new_G3195_ | ~new_G3196_;
  assign new_G3348_ = ~new_G3197_ | ~new_G3198_;
  assign new_G3351_ = ~new_G3202_ | ~new_G3203_;
  assign new_G3355_ = ~new_G3204_ | ~new_G3081_;
  assign new_G3358_ = ~new_G3205_ & ~new_G3084_;
  assign new_G3359_ = ~new_G3206_ & ~new_G3085_;
  assign new_G3360_ = new_G2804_ | new_G3163_;
  assign new_G3363_ = ~new_G3002_ | ~new_G3265_;
  assign new_G3364_ = ~new_G2999_ | ~new_G3266_;
  assign new_G3365_ = ~new_G3008_ | ~new_G3267_;
  assign new_G3366_ = ~new_G3005_ | ~new_G3268_;
  assign new_G3367_ = ~new_G3029_ | ~new_G3269_;
  assign new_G3368_ = ~new_G3026_ | ~new_G3270_;
  assign new_G3369_ = ~new_G3035_ | ~new_G3271_;
  assign new_G3370_ = ~new_G3032_ | ~new_G3272_;
  assign new_G3371_ = ~new_G3191_ | ~new_G3190_;
  assign new_G3374_ = ~new_G3060_;
  assign new_G3377_ = ~new_G3273_ | ~new_G3274_;
  assign new_G3380_ = ~new_G3275_ | ~new_G3276_;
  assign new_G3383_ = ~new_G3280_ | ~new_G3104_;
  assign new_G3386_ = ~new_G3282_ | ~new_G3114_;
  assign new_G3393_ = ~new_G3283_ | ~new_G3116_;
  assign new_G3404_ = ~new_G3284_ | ~new_G3118_;
  assign new_G3415_ = ~new_G3285_ | ~new_G3120_;
  assign new_G3421_ = ~new_G3286_ | ~new_G3122_;
  assign new_G3428_ = ~new_G3287_ | ~new_G3124_;
  assign new_G3438_ = ~new_G3288_ | ~new_G3126_;
  assign new_G3449_ = ~new_G3289_ | ~new_G3128_;
  assign new_G3459_ = ~new_G3290_ | ~new_G3130_;
  assign new_G3466_ = ~new_G3211_;
  assign new_G3467_ = ~new_G3132_ | ~new_G3291_;
  assign new_G3474_ = ~new_G3134_ | ~new_G3292_;
  assign new_G3485_ = ~new_G3136_ | ~new_G3293_;
  assign new_G3495_ = ~new_G3138_ | ~new_G3294_;
  assign new_G3503_ = ~new_G3140_ | ~new_G3295_;
  assign new_G3517_ = ~new_G3142_ | ~new_G3296_;
  assign new_G3533_ = ~new_G3144_ | ~new_G3297_;
  assign new_G3546_ = ~new_G3146_ | ~new_G3298_;
  assign new_G3552_ = ~new_G3148_ | ~new_G3299_;
  assign new_G3559_ = ~new_G3300_ | ~new_G3151_;
  assign new_G3570_ = ~new_G3301_ | ~new_G3153_;
  assign new_G3576_ = ~new_G3302_ | ~new_G3155_;
  assign new_G3583_ = ~new_G3313_ | ~new_G3158_;
  assign new_G3594_ = ~new_G3314_ | ~new_G3160_;
  assign new_G3604_ = ~new_G3222_ | ~new_G1588_;
  assign new_G3605_ = ~new_G3222_;
  assign new_G3606_ = ~new_G3225_;
  assign new_G3607_ = ~new_G3228_;
  assign new_G3608_ = ~new_G3231_;
  assign new_G3609_ = ~new_G3234_;
  assign new_G3610_ = ~new_G3237_;
  assign new_G3611_ = ~new_G3165_ | ~new_G3315_;
  assign new_G3621_ = ~new_G3167_ | ~new_G3316_;
  assign new_G3629_ = ~new_G3170_ | ~new_G3331_;
  assign new_G3645_ = ~new_G3172_ | ~new_G3332_;
  assign new_G3658_ = ~new_G3174_ | ~new_G3333_;
  assign new_G3664_ = ~new_G3244_;
  assign new_G3665_ = ~new_G3253_;
  assign new_G3666_ = ~new_G3334_ | ~new_G3335_;
  assign new_G3670_ = ~new_G3180_ | ~new_G3336_;
  assign new_G3674_ = ~new_G3337_ | ~new_G3183_;
  assign new_G3677_ = ~new_G3338_ | ~new_G3339_;
  assign new_G3681_ = ~new_G3340_ | ~new_G3341_;
  assign new_G3685_ = ~new_G3188_ | ~new_G3342_;
  assign new_G3688_ = new_G3208_ & new_G2872_;
  assign new_G3689_ = ~new_G3215_;
  assign new_G3690_ = ~new_G3219_;
  assign new_G3691_ = ~new_G3241_;
  assign new_G3692_ = ~new_G3247_;
  assign new_G3693_ = ~new_G3250_;
  assign new_G3694_ = ~new_G3256_;
  assign new_G3695_ = ~new_G3259_;
  assign new_G3696_ = ~new_G3262_;
  assign new_G3697_ = ~new_G3365_ | ~new_G3366_;
  assign new_G3700_ = ~new_G3363_ | ~new_G3364_;
  assign new_G3703_ = ~new_G3369_ | ~new_G3370_;
  assign new_G3706_ = ~new_G3367_ | ~new_G3368_;
  assign new_G3709_ = ~new_G3277_;
  assign new_G3710_ = ~new_G3359_ | ~new_G3358_;
  assign new_G3713_ = new_G3303_ & new_G2788_;
  assign new_G3714_ = ~new_G1386_ | ~new_G3605_;
  assign new_G3715_ = ~new_G3360_;
  assign new_G3716_ = new_G3317_ & new_G2844_;
  assign new_G3717_ = new_G3317_ & new_G2844_;
  assign new_G3718_ = ~new_G3371_;
  assign new_G3719_ = ~new_G3371_ | ~new_G3343_;
  assign new_G3720_ = ~new_G3344_;
  assign new_G3723_ = ~new_G3351_;
  assign new_G3726_ = ~new_G3348_;
  assign new_G3729_ = ~new_G3348_;
  assign new_G3732_ = ~new_G3355_;
  assign new_G3735_ = ~new_G3355_;
  assign new_G3738_ = ~new_G3383_;
  assign new_G3739_ = new_G3208_ | new_G3688_;
  assign new_G3742_ = ~new_G3303_;
  assign new_G3745_ = ~new_G3317_;
  assign new_G3748_ = ~new_G3317_;
  assign new_G3751_ = ~new_G3374_;
  assign new_G3752_ = ~new_G3374_ | ~new_G3099_;
  assign new_G3753_ = ~new_G3377_;
  assign new_G3754_ = ~new_G3380_;
  assign new_G3755_ = ~new_G3380_ | ~new_G3709_;
  assign new_G3756_ = new_G3467_ & new_G2711_;
  assign new_G3757_ = new_G3474_ & new_G3467_ & new_G2715_;
  assign new_G3758_ = new_G3474_ & new_G3485_ & new_G3467_ & new_G2720_;
  assign new_G3759_ = new_G2759_ & new_G3559_ & new_G2752_ & new_G2780_;
  assign new_G3760_ = new_G3386_ & new_G2675_;
  assign new_G3761_ = new_G3393_ & new_G3386_ & new_G2679_;
  assign new_G3762_ = new_G3393_ & new_G3404_ & new_G3386_ & new_G2685_;
  assign new_G3763_ = new_G2817_ & new_G3611_ & new_G2810_ & new_G2837_;
  assign new_G3764_ = ~new_G3415_;
  assign new_G3765_ = new_G3386_ & new_G3393_ & new_G3415_ & new_G3404_;
  assign new_G3768_ = new_G3393_ & new_G2679_;
  assign new_G3769_ = new_G3404_ & new_G2685_ & new_G3393_;
  assign new_G3770_ = new_G3415_ & new_G3404_ & new_G3393_;
  assign new_G3771_ = new_G3393_ & new_G2679_;
  assign new_G3772_ = new_G2685_ & new_G3404_ & new_G3393_;
  assign new_G3773_ = new_G3404_ & new_G2685_;
  assign new_G3774_ = new_G3415_ & new_G3404_;
  assign new_G3775_ = new_G3404_ & new_G2685_;
  assign new_G3776_ = new_G3421_ & new_G3428_ & new_G3459_ & new_G3438_ & new_G3449_;
  assign new_G3779_ = new_G3421_ & new_G2693_;
  assign new_G3780_ = new_G3428_ & new_G3421_ & new_G2696_;
  assign new_G3781_ = new_G3428_ & new_G3438_ & new_G3421_ & new_G2700_;
  assign new_G3782_ = new_G2705_ & new_G3449_ & new_G3438_ & new_G3421_ & new_G3428_;
  assign new_G3783_ = new_G3428_ & new_G2696_;
  assign new_G3784_ = new_G3438_ & new_G2700_ & new_G3428_;
  assign new_G3785_ = new_G3428_ & new_G3449_ & new_G3438_ & new_G2705_;
  assign new_G3786_ = new_G3449_ & n2631_lo & new_G3459_ & new_G3438_ & new_G3428_;
  assign new_G3787_ = new_G2700_ & new_G3438_;
  assign new_G3788_ = new_G3449_ & new_G3438_ & new_G2705_;
  assign new_G3789_ = new_G3449_ & n2631_lo & new_G3459_ & new_G3438_;
  assign new_G3790_ = new_G3449_ & new_G2705_;
  assign new_G3791_ = n2631_lo & new_G3459_ & new_G3449_;
  assign new_G3792_ = n2631_lo & new_G3459_;
  assign new_G3793_ = new_G3467_ & new_G3546_ & new_G3485_ & new_G3474_;
  assign new_G3796_ = new_G3474_ & new_G2715_;
  assign new_G3797_ = new_G3485_ & new_G2720_ & new_G3474_;
  assign new_G3798_ = new_G3546_ & new_G3485_ & new_G3474_;
  assign new_G3799_ = new_G3474_ & new_G2715_;
  assign new_G3800_ = new_G3485_ & new_G2720_ & new_G3474_;
  assign new_G3801_ = new_G3485_ & new_G2720_;
  assign new_G3802_ = new_G3503_ & new_G3552_ & new_G3533_ & new_G3517_ & new_G3495_;
  assign new_G3805_ = new_G3495_ & new_G2727_;
  assign new_G3806_ = new_G3503_ & new_G3495_ & new_G2731_;
  assign new_G3807_ = new_G3503_ & new_G3517_ & new_G3495_ & new_G2737_;
  assign new_G3808_ = new_G2744_ & new_G3533_ & new_G3517_ & new_G3495_ & new_G3503_;
  assign new_G3809_ = new_G3503_ & new_G2731_;
  assign new_G3810_ = new_G3517_ & new_G2737_ & new_G3503_;
  assign new_G3811_ = new_G3503_ & new_G3533_ & new_G3517_ & new_G2744_;
  assign new_G3812_ = new_G3533_ & new_G3552_ & new_G3517_ & new_G3503_;
  assign new_G3813_ = new_G3503_ & new_G2731_;
  assign new_G3814_ = new_G3517_ & new_G2737_ & new_G3503_;
  assign new_G3815_ = new_G3503_ & new_G3533_ & new_G3517_ & new_G2744_;
  assign new_G3816_ = new_G3517_ & new_G2737_;
  assign new_G3817_ = new_G3533_ & new_G3517_ & new_G2744_;
  assign new_G3818_ = new_G3552_ & new_G3517_ & new_G3533_;
  assign new_G3819_ = new_G3517_ & new_G2737_;
  assign new_G3820_ = new_G3533_ & new_G3517_ & new_G2744_;
  assign new_G3821_ = new_G3533_ & new_G2744_;
  assign new_G3822_ = new_G3546_ & new_G3485_;
  assign new_G3823_ = new_G3552_ & new_G3533_;
  assign new_G3824_ = ~new_G3570_;
  assign new_G3825_ = new_G2752_ & new_G2759_ & new_G3570_ & new_G3559_;
  assign new_G3828_ = new_G3559_ & new_G2780_ & new_G2759_;
  assign new_G3829_ = new_G3570_ & new_G3559_ & new_G2759_;
  assign new_G3830_ = new_G2780_ & new_G3559_ & new_G2759_;
  assign new_G3831_ = new_G3559_ & new_G2780_;
  assign new_G3832_ = new_G3570_ & new_G3559_;
  assign new_G3833_ = new_G3559_ & new_G2780_;
  assign new_G3834_ = new_G3576_ & new_G3303_ & new_G2797_ & new_G3583_ & new_G3594_;
  assign new_G3837_ = new_G3576_ & new_G2540_;
  assign new_G3838_ = new_G3303_ & new_G3576_ & new_G2788_;
  assign new_G3839_ = new_G3303_ & new_G3583_ & new_G3576_ & new_G2792_;
  assign new_G3840_ = new_G2804_ & new_G3594_ & new_G3583_ & new_G3576_ & new_G3303_;
  assign new_G3841_ = new_G3583_ & new_G2792_ & new_G3303_;
  assign new_G3842_ = new_G3303_ & new_G3594_ & new_G3583_ & new_G2804_;
  assign new_G3843_ = new_G3594_ & n2859_lo & new_G2797_ & new_G3583_ & new_G3303_;
  assign new_G3844_ = new_G2792_ & new_G3583_;
  assign new_G3845_ = new_G3594_ & new_G3583_ & new_G2804_;
  assign new_G3846_ = new_G3594_ & n2859_lo & new_G2797_ & new_G3583_;
  assign new_G3847_ = new_G3594_ & new_G2804_;
  assign new_G3848_ = n2859_lo & new_G2797_ & new_G3594_;
  assign new_G3849_ = ~new_G3604_ | ~new_G3714_;
  assign new_G3852_ = new_G2810_ & new_G3658_ & new_G3611_ & new_G2817_;
  assign new_G3855_ = new_G3611_ & new_G2837_ & new_G2817_;
  assign new_G3856_ = new_G3658_ & new_G3611_ & new_G2817_;
  assign new_G3857_ = new_G3611_ & new_G2837_ & new_G2817_;
  assign new_G3858_ = new_G3611_ & new_G2837_;
  assign new_G3859_ = new_G3317_ & new_G2865_ & new_G3645_ & new_G3629_ & new_G3621_;
  assign new_G3862_ = new_G3621_ & new_G2543_;
  assign new_G3863_ = new_G3317_ & new_G3621_ & new_G2844_;
  assign new_G3864_ = new_G3317_ & new_G3629_ & new_G3621_ & new_G2850_;
  assign new_G3865_ = new_G2857_ & new_G3645_ & new_G3629_ & new_G3621_ & new_G3317_;
  assign new_G3866_ = new_G3629_ & new_G2850_ & new_G3317_;
  assign new_G3867_ = new_G3317_ & new_G3645_ & new_G3629_ & new_G2857_;
  assign new_G3868_ = new_G3645_ & new_G2865_ & new_G3629_ & new_G3317_;
  assign new_G3869_ = new_G3629_ & new_G2850_ & new_G3317_;
  assign new_G3870_ = new_G3317_ & new_G3645_ & new_G3629_ & new_G2857_;
  assign new_G3871_ = new_G3629_ & new_G2850_;
  assign new_G3872_ = new_G3645_ & new_G3629_ & new_G2857_;
  assign new_G3873_ = new_G2865_ & new_G3629_ & new_G3645_;
  assign new_G3874_ = new_G3629_ & new_G2850_;
  assign new_G3875_ = new_G3645_ & new_G3629_ & new_G2857_;
  assign new_G3876_ = new_G3645_ & new_G2857_;
  assign new_G3877_ = new_G3658_ & new_G3611_;
  assign new_G3878_ = new_G2865_ & new_G3645_;
  assign new_G3879_ = ~new_G3666_;
  assign new_G3882_ = ~new_G3670_;
  assign new_G3885_ = ~new_G3677_;
  assign new_G3888_ = ~new_G3681_;
  assign new_G3891_ = ~new_G3674_;
  assign new_G3894_ = ~new_G3674_;
  assign new_G3897_ = ~new_G3685_;
  assign new_G3900_ = ~new_G3685_;
  assign new_G3903_ = ~new_G3094_ | ~new_G3718_;
  assign new_G3904_ = ~new_G3710_;
  assign new_G3905_ = ~new_G3710_ | ~new_G3738_;
  assign new_G3906_ = ~new_G3459_;
  assign new_G3909_ = ~new_G3386_;
  assign new_G3912_ = ~new_G3386_;
  assign new_G3915_ = ~new_G3393_;
  assign new_G3918_ = ~new_G3393_;
  assign new_G3921_ = ~new_G3404_;
  assign new_G3924_ = ~new_G3404_;
  assign new_G3927_ = ~new_G3421_;
  assign new_G3930_ = ~new_G3428_;
  assign new_G3933_ = ~new_G3438_;
  assign new_G3936_ = ~new_G3449_;
  assign new_G3939_ = ~new_G3546_;
  assign new_G3942_ = ~new_G3485_;
  assign new_G3945_ = ~new_G3467_;
  assign new_G3948_ = ~new_G3474_;
  assign new_G3951_ = ~new_G3546_;
  assign new_G3954_ = ~new_G3485_;
  assign new_G3957_ = ~new_G3467_;
  assign new_G3960_ = ~new_G3474_;
  assign new_G3963_ = ~new_G3552_;
  assign new_G3966_ = ~new_G3533_;
  assign new_G3969_ = ~new_G3495_;
  assign new_G3972_ = ~new_G3517_;
  assign new_G3975_ = ~new_G3503_;
  assign new_G3978_ = ~new_G3503_;
  assign new_G3981_ = ~new_G3552_;
  assign new_G3984_ = ~new_G3533_;
  assign new_G3987_ = ~new_G3495_;
  assign new_G3990_ = ~new_G3517_;
  assign new_G3993_ = ~new_G3559_;
  assign new_G3996_ = ~new_G3559_;
  assign new_G3999_ = ~new_G3576_;
  assign new_G4002_ = ~new_G3583_;
  assign new_G4005_ = ~new_G3594_;
  assign new_G4008_ = ~new_G3658_;
  assign new_G4011_ = ~new_G3611_;
  assign new_G4014_ = ~new_G3658_;
  assign new_G4017_ = ~new_G3611_;
  assign new_G4020_ = ~new_G3645_;
  assign new_G4023_ = ~new_G3621_;
  assign new_G4026_ = ~new_G3629_;
  assign new_G4029_ = ~new_G3645_;
  assign new_G4032_ = ~new_G3621_;
  assign new_G4035_ = ~new_G3629_;
  assign new_G4038_ = ~new_G3697_;
  assign new_G4039_ = ~new_G3700_;
  assign new_G4040_ = ~new_G3703_;
  assign new_G4041_ = ~new_G3706_;
  assign new_G4042_ = ~new_G2644_ | ~new_G3751_;
  assign new_G4043_ = ~new_G3277_ | ~new_G3754_;
  assign new_G4044_ = new_G3758_ | new_G3757_ | new_G2667_ | new_G3756_;
  assign new_G4045_ = new_G3759_ | new_G3110_ | new_G2492_ | new_G3109_;
  assign new_G4046_ = new_G3762_ | new_G3761_ | new_G2670_ | new_G3760_;
  assign new_G4047_ = new_G3763_ | new_G3112_ | new_G2492_ | new_G3111_;
  assign new_G4048_ = new_G3781_ | new_G3780_ | new_G2692_ | new_G3779_ | new_G3782_;
  assign new_G4051_ = new_G2715_ | new_G3801_;
  assign new_G4054_ = new_G3807_ | new_G3806_ | new_G2726_ | new_G3805_ | new_G3808_;
  assign new_G4058_ = new_G2737_ | new_G3821_;
  assign new_G4061_ = new_G3839_ | new_G3838_ | new_G2787_ | new_G3837_ | new_G3840_;
  assign new_G4064_ = ~new_G3742_;
  assign new_G4065_ = new_G2832_ | new_G3858_;
  assign new_G4068_ = new_G3864_ | new_G3863_ | new_G2843_ | new_G3862_ | new_G3865_;
  assign new_G4072_ = new_G2850_ | new_G3876_;
  assign new_G4075_ = ~new_G3745_;
  assign new_G4076_ = ~new_G3748_;
  assign new_G4077_ = ~new_G3903_ | ~new_G3719_;
  assign new_G4080_ = ~new_G3726_;
  assign new_G4081_ = ~new_G3729_;
  assign new_G4082_ = ~new_G3732_;
  assign new_G4083_ = ~new_G3735_;
  assign new_G4084_ = new_G3344_ & new_G2879_ & new_G3726_;
  assign new_G4085_ = new_G3720_ & new_G3192_ & new_G3729_;
  assign new_G4086_ = new_G3351_ & new_G2883_ & new_G3732_;
  assign new_G4087_ = new_G3723_ & new_G3199_ & new_G3735_;
  assign new_G4088_ = ~new_G3383_ | ~new_G3904_;
  assign new_G4089_ = ~new_G3739_ | ~n3339_lo;
  assign new_G4092_ = new_G3770_ | new_G3769_ | new_G2675_ | new_G3768_;
  assign new_G4095_ = ~new_G3772_ & ~new_G2675_ & ~new_G3771_;
  assign new_G4098_ = new_G3774_ | new_G2679_ | new_G3773_;
  assign new_G4101_ = ~new_G2679_ & ~new_G3775_;
  assign new_G4104_ = new_G3785_ | new_G3784_ | new_G2693_ | new_G3783_ | new_G3786_;
  assign new_G4107_ = new_G3789_ | new_G3788_ | new_G2696_ | new_G3787_;
  assign new_G4110_ = new_G3791_ | new_G2700_ | new_G3790_;
  assign new_G4113_ = new_G2705_ | new_G3792_;
  assign new_G4116_ = new_G3798_ | new_G3797_ | new_G2711_ | new_G3796_;
  assign new_G4119_ = ~new_G3800_ & ~new_G2711_ & ~new_G3799_;
  assign new_G4122_ = new_G3818_ | new_G3817_ | new_G2731_ | new_G3816_;
  assign new_G4125_ = new_G3811_ | new_G3810_ | new_G2727_ | new_G3809_ | new_G3812_;
  assign new_G4128_ = ~new_G3820_ & ~new_G2731_ & ~new_G3819_;
  assign new_G4131_ = ~new_G3815_ & ~new_G3814_ & ~new_G2727_ & ~new_G3813_;
  assign new_G4134_ = new_G3829_ | new_G3828_ | new_G2770_ | new_G3161_;
  assign new_G4137_ = ~new_G3830_ & ~new_G2770_ & ~new_G3162_;
  assign new_G4140_ = new_G3832_ | new_G2774_ | new_G3831_;
  assign new_G4143_ = ~new_G2774_ & ~new_G3833_;
  assign new_G4146_ = new_G3842_ | new_G3841_ | new_G2540_ | new_G3713_ | new_G3843_;
  assign new_G4149_ = new_G3846_ | new_G3845_ | new_G2788_ | new_G3844_;
  assign new_G4152_ = new_G3848_ | new_G2792_ | new_G3847_;
  assign new_G4155_ = new_G3856_ | new_G3855_ | new_G2828_ | new_G3176_;
  assign new_G4158_ = ~new_G3857_ & ~new_G2828_ & ~new_G3177_;
  assign new_G4161_ = new_G3873_ | new_G3872_ | new_G2844_ | new_G3871_;
  assign new_G4164_ = new_G3867_ | new_G3866_ | new_G2543_ | new_G3716_ | new_G3868_;
  assign new_G4167_ = ~new_G3875_ & ~new_G2844_ & ~new_G3874_;
  assign new_G4170_ = ~new_G3870_ & ~new_G3869_ & ~new_G2543_ & ~new_G3717_;
  assign new_G4173_ = ~new_G3700_ | ~new_G4038_;
  assign new_G4174_ = ~new_G3697_ | ~new_G4039_;
  assign new_G4175_ = ~new_G3706_ | ~new_G4040_;
  assign new_G4176_ = ~new_G3703_ | ~new_G4041_;
  assign new_G4177_ = ~new_G4042_ | ~new_G3752_;
  assign new_G4180_ = ~new_G3755_ | ~new_G4043_;
  assign new_G4183_ = ~new_G3849_;
  assign new_G4184_ = ~new_G3906_ | ~new_G1510_;
  assign new_G4185_ = ~new_G3906_;
  assign new_G4186_ = ~new_G3909_;
  assign new_G4187_ = ~new_G3912_;
  assign new_G4188_ = ~new_G3915_;
  assign new_G4189_ = ~new_G3918_;
  assign new_G4190_ = ~new_G3921_ | ~new_G3131_;
  assign new_G4191_ = ~new_G3921_;
  assign new_G4192_ = ~new_G3924_ | ~new_G3466_;
  assign new_G4193_ = ~new_G3924_;
  assign new_G4194_ = new_G3776_ & n2631_lo;
  assign new_G4195_ = ~new_G3927_;
  assign new_G4196_ = ~new_G3930_;
  assign new_G4197_ = ~new_G3933_;
  assign new_G4198_ = ~new_G3936_;
  assign new_G4199_ = ~new_G3802_;
  assign new_G4200_ = ~new_G3948_;
  assign new_G4201_ = ~new_G3960_;
  assign new_G4202_ = ~new_G3975_;
  assign new_G4203_ = ~new_G3978_;
  assign new_G4204_ = ~new_G3993_ | ~new_G3164_;
  assign new_G4205_ = ~new_G3993_;
  assign new_G4206_ = ~new_G3996_ | ~new_G3610_;
  assign new_G4207_ = ~new_G3996_;
  assign new_G4208_ = new_G3834_ & n2859_lo;
  assign new_G4209_ = ~new_G3999_;
  assign new_G4210_ = ~new_G4002_;
  assign new_G4211_ = ~new_G4005_ | ~new_G3715_;
  assign new_G4212_ = ~new_G4005_;
  assign new_G4213_ = ~new_G3859_;
  assign new_G4214_ = ~new_G3891_;
  assign new_G4215_ = ~new_G3894_;
  assign new_G4216_ = ~new_G3897_;
  assign new_G4217_ = ~new_G3900_;
  assign new_G4218_ = new_G3670_ & new_G3666_ & new_G3891_;
  assign new_G4219_ = new_G3882_ & new_G3879_ & new_G3894_;
  assign new_G4220_ = new_G3681_ & new_G3677_ & new_G3897_;
  assign new_G4221_ = new_G3888_ & new_G3885_ & new_G3900_;
  assign new_G4222_ = new_G3849_ & new_G1264_ & new_G2003_;
  assign new_G4223_ = new_G3192_ & new_G3344_ & new_G4080_;
  assign new_G4224_ = new_G2879_ & new_G3720_ & new_G4081_;
  assign new_G4225_ = new_G3199_ & new_G3351_ & new_G4082_;
  assign new_G4226_ = new_G2883_ & new_G3723_ & new_G4083_;
  assign new_G4227_ = ~new_G4088_ | ~new_G3905_;
  assign new_G4230_ = ~new_G3939_;
  assign new_G4231_ = ~new_G3942_;
  assign new_G4232_ = ~new_G3945_;
  assign new_G4233_ = ~new_G3951_;
  assign new_G4234_ = ~new_G3954_;
  assign new_G4235_ = ~new_G3957_;
  assign new_G4236_ = ~new_G3963_;
  assign new_G4237_ = ~new_G3966_;
  assign new_G4238_ = ~new_G3969_;
  assign new_G4239_ = ~new_G3972_;
  assign new_G4240_ = ~new_G3990_;
  assign new_G4241_ = ~new_G3981_;
  assign new_G4242_ = ~new_G3984_;
  assign new_G4243_ = ~new_G3987_;
  assign new_G4244_ = ~new_G4008_;
  assign new_G4245_ = ~new_G4011_;
  assign new_G4246_ = ~new_G4014_;
  assign new_G4247_ = ~new_G4017_;
  assign new_G4248_ = ~new_G4020_;
  assign new_G4249_ = ~new_G4023_;
  assign new_G4250_ = ~new_G4026_;
  assign new_G4251_ = ~new_G4035_;
  assign new_G4252_ = ~new_G4029_;
  assign new_G4253_ = ~new_G4032_;
  assign new_G4254_ = ~new_G4173_ | ~new_G4174_;
  assign new_G4257_ = ~new_G4175_ | ~new_G4176_;
  assign new_G4260_ = new_G3793_ & new_G4054_;
  assign new_G4261_ = new_G4061_ & new_G3825_;
  assign new_G4262_ = new_G4048_ & new_G3765_;
  assign new_G4263_ = new_G3852_ & new_G4068_;
  assign new_G4264_ = ~new_G4077_;
  assign new_G4265_ = ~new_G1338_ | ~new_G4185_;
  assign new_G4266_ = ~new_G4092_;
  assign new_G4267_ = ~new_G4092_ | ~new_G4186_;
  assign new_G4268_ = ~new_G4095_;
  assign new_G4269_ = ~new_G4095_ | ~new_G4187_;
  assign new_G4270_ = ~new_G4098_;
  assign new_G4271_ = ~new_G4098_ | ~new_G4188_;
  assign new_G4272_ = ~new_G4101_;
  assign new_G4273_ = ~new_G4101_ | ~new_G4189_;
  assign new_G4274_ = ~new_G2915_ | ~new_G4191_;
  assign new_G4275_ = ~new_G3211_ | ~new_G4193_;
  assign new_G4276_ = new_G4048_ | new_G4194_;
  assign new_G4282_ = ~new_G4104_;
  assign new_G4283_ = ~new_G4104_ | ~new_G4195_;
  assign new_G4284_ = ~new_G4107_;
  assign new_G4285_ = ~new_G4107_ | ~new_G4196_;
  assign new_G4286_ = ~new_G4110_;
  assign new_G4287_ = ~new_G4110_ | ~new_G4197_;
  assign new_G4288_ = ~new_G4113_;
  assign new_G4289_ = ~new_G4113_ | ~new_G4198_;
  assign new_G4290_ = ~new_G4054_;
  assign new_G4293_ = ~new_G4134_;
  assign new_G4294_ = ~new_G4134_ | ~new_G3606_;
  assign new_G4295_ = ~new_G4137_;
  assign new_G4296_ = ~new_G4137_ | ~new_G3607_;
  assign new_G4297_ = ~new_G4140_;
  assign new_G4298_ = ~new_G4140_ | ~new_G3608_;
  assign new_G4299_ = ~new_G4143_;
  assign new_G4300_ = ~new_G4143_ | ~new_G3609_;
  assign new_G4301_ = ~new_G2966_ | ~new_G4205_;
  assign new_G4302_ = ~new_G3237_ | ~new_G4207_;
  assign new_G4303_ = new_G4061_ | new_G4208_;
  assign new_G4309_ = ~new_G4146_;
  assign new_G4310_ = ~new_G4146_ | ~new_G4209_;
  assign new_G4311_ = ~new_G4149_;
  assign new_G4312_ = ~new_G4149_ | ~new_G4064_;
  assign new_G4313_ = ~new_G4152_;
  assign new_G4314_ = ~new_G4152_ | ~new_G4210_;
  assign new_G4315_ = ~new_G3360_ | ~new_G4212_;
  assign new_G4316_ = ~new_G4068_;
  assign new_G4319_ = new_G3879_ & new_G3670_ & new_G4214_;
  assign new_G4320_ = new_G3666_ & new_G3882_ & new_G4215_;
  assign new_G4321_ = new_G3885_ & new_G3681_ & new_G4216_;
  assign new_G4322_ = new_G3677_ & new_G3888_ & new_G4217_;
  assign new_G4323_ = new_G2324_ | new_G2600_ | new_G4222_;
  assign new_G4329_ = ~new_G4223_ & ~new_G4084_;
  assign new_G4330_ = ~new_G4224_ & ~new_G4085_;
  assign new_G4331_ = ~new_G4225_ & ~new_G4086_;
  assign new_G4332_ = ~new_G4226_ & ~new_G4087_;
  assign new_G4333_ = ~new_G4180_;
  assign new_G4334_ = new_G3739_ & new_G4089_;
  assign new_G4335_ = new_G4089_ & n3339_lo;
  assign new_G4336_ = new_G4051_ | new_G3822_;
  assign new_G4339_ = ~new_G4116_;
  assign new_G4340_ = ~new_G4051_;
  assign new_G4343_ = ~new_G4119_;
  assign new_G4344_ = ~new_G4122_;
  assign new_G4345_ = ~new_G4122_ | ~new_G3218_;
  assign new_G4346_ = new_G4058_ | new_G3823_;
  assign new_G4349_ = ~new_G4125_;
  assign new_G4350_ = ~new_G4128_;
  assign new_G4351_ = ~new_G4128_ | ~new_G3690_;
  assign new_G4352_ = ~new_G4058_;
  assign new_G4355_ = ~new_G4131_;
  assign new_G4356_ = new_G4065_ | new_G3877_;
  assign new_G4359_ = ~new_G4155_;
  assign new_G4360_ = ~new_G4065_;
  assign new_G4363_ = ~new_G4158_;
  assign new_G4364_ = new_G4072_ | new_G3878_;
  assign new_G4367_ = ~new_G4161_;
  assign new_G4368_ = ~new_G4164_;
  assign new_G4369_ = ~new_G4167_;
  assign new_G4370_ = ~new_G4167_ | ~new_G3695_;
  assign new_G4371_ = ~new_G4072_;
  assign new_G4374_ = ~new_G4170_;
  assign new_G4375_ = ~new_G4177_;
  assign new_G4376_ = ~new_G4177_ | ~new_G3753_;
  assign new_G4377_ = ~new_G4227_;
  assign new_G4378_ = ~new_G4184_ | ~new_G4265_;
  assign new_G4381_ = ~new_G3909_ | ~new_G4266_;
  assign new_G4382_ = ~new_G3912_ | ~new_G4268_;
  assign new_G4383_ = ~new_G3915_ | ~new_G4270_;
  assign new_G4384_ = ~new_G3918_ | ~new_G4272_;
  assign new_G4385_ = ~new_G4190_ | ~new_G4274_;
  assign new_G4386_ = ~new_G4192_ | ~new_G4275_;
  assign new_G4387_ = ~new_G3927_ | ~new_G4282_;
  assign new_G4388_ = ~new_G3930_ | ~new_G4284_;
  assign new_G4389_ = ~new_G3933_ | ~new_G4286_;
  assign new_G4390_ = ~new_G3936_ | ~new_G4288_;
  assign new_G4391_ = ~new_G3225_ | ~new_G4293_;
  assign new_G4392_ = ~new_G3228_ | ~new_G4295_;
  assign new_G4393_ = ~new_G3231_ | ~new_G4297_;
  assign new_G4394_ = ~new_G3234_ | ~new_G4299_;
  assign new_G4395_ = ~new_G4204_ | ~new_G4301_;
  assign new_G4396_ = ~new_G4206_ | ~new_G4302_;
  assign new_G4397_ = ~new_G3999_ | ~new_G4309_;
  assign new_G4398_ = ~new_G3742_ | ~new_G4311_;
  assign new_G4399_ = ~new_G4002_ | ~new_G4313_;
  assign new_G4400_ = ~new_G4211_ | ~new_G4315_;
  assign new_G4403_ = ~new_G4319_ & ~new_G4218_;
  assign new_G4404_ = ~new_G4320_ & ~new_G4219_;
  assign new_G4405_ = ~new_G4321_ & ~new_G4220_;
  assign new_G4406_ = ~new_G4322_ & ~new_G4221_;
  assign new_G4407_ = ~new_G4254_;
  assign new_G4408_ = ~new_G4257_;
  assign new_G4409_ = new_G4334_ | new_G4335_;
  assign new_G4413_ = ~new_G2948_ | ~new_G4344_;
  assign new_G4414_ = ~new_G3219_ | ~new_G4350_;
  assign new_G4415_ = ~new_G3259_ | ~new_G4369_;
  assign new_G4416_ = ~new_G3377_ | ~new_G4375_;
  assign new_G4417_ = ~new_G4330_ | ~new_G4329_;
  assign new_G4420_ = ~new_G4332_ | ~new_G4331_;
  assign new_G4423_ = new_G4323_ & new_G1554_ & new_G1565_;
  assign new_G4424_ = new_G4323_ & new_G1629_ & new_G1640_;
  assign new_G4425_ = new_G4323_ & new_G1652_ & new_G1663_;
  assign new_G4426_ = new_G4323_ & new_G1674_ & new_G1685_;
  assign new_G4427_ = ~new_G4381_ | ~new_G4267_;
  assign new_G4428_ = ~new_G4382_ | ~new_G4269_;
  assign new_G4429_ = ~new_G4383_ | ~new_G4271_;
  assign new_G4430_ = ~new_G4384_ | ~new_G4273_;
  assign new_G4431_ = ~new_G4385_;
  assign new_G4432_ = ~new_G4276_;
  assign new_G4437_ = ~new_G4387_ | ~new_G4283_;
  assign new_G4440_ = ~new_G4388_ | ~new_G4285_;
  assign new_G4443_ = ~new_G4389_ | ~new_G4287_;
  assign new_G4446_ = ~new_G4390_ | ~new_G4289_;
  assign new_G4449_ = new_G4276_ & new_G3764_;
  assign new_G4450_ = new_G4290_ & new_G4199_;
  assign new_G4453_ = ~new_G4391_ | ~new_G4294_;
  assign new_G4454_ = ~new_G4392_ | ~new_G4296_;
  assign new_G4455_ = ~new_G4393_ | ~new_G4298_;
  assign new_G4456_ = ~new_G4394_ | ~new_G4300_;
  assign new_G4457_ = ~new_G4395_;
  assign new_G4458_ = ~new_G4303_;
  assign new_G4463_ = ~new_G4397_ | ~new_G4310_;
  assign new_G4466_ = ~new_G4398_ | ~new_G4312_;
  assign new_G4469_ = ~new_G4399_ | ~new_G4314_;
  assign new_G4472_ = new_G4303_ & new_G3824_;
  assign new_G4473_ = new_G4316_ & new_G4213_;
  assign new_G4476_ = ~new_G4336_;
  assign new_G4477_ = ~new_G4336_ | ~new_G3214_;
  assign new_G4478_ = ~new_G4340_;
  assign new_G4479_ = ~new_G4340_ | ~new_G3689_;
  assign new_G4480_ = ~new_G4345_ | ~new_G4413_;
  assign new_G4483_ = ~new_G4346_;
  assign new_G4484_ = ~new_G4351_ | ~new_G4414_;
  assign new_G4487_ = ~new_G4352_;
  assign new_G4488_ = ~new_G4356_;
  assign new_G4489_ = ~new_G4356_ | ~new_G3240_;
  assign new_G4490_ = ~new_G4360_;
  assign new_G4491_ = ~new_G4360_ | ~new_G3692_;
  assign new_G4492_ = ~new_G4364_;
  assign new_G4493_ = ~new_G4364_ | ~new_G4367_;
  assign new_G4494_ = ~new_G4370_ | ~new_G4415_;
  assign new_G4497_ = ~new_G4371_;
  assign new_G4498_ = ~new_G4404_ | ~new_G4403_;
  assign new_G4501_ = ~new_G4406_ | ~new_G4405_;
  assign new_G4504_ = ~new_G4416_ | ~new_G4376_;
  assign new_G4507_ = ~new_G4378_;
  assign new_G4508_ = ~new_G4400_;
  assign new_G4509_ = new_G4409_ & n4659_lo & new_G1242_;
  assign new_G4510_ = ~new_G4428_;
  assign new_G4511_ = ~new_G4430_;
  assign new_G4512_ = new_G4276_ & new_G4427_;
  assign new_G4513_ = new_G4276_ & new_G4429_;
  assign new_G4514_ = new_G4276_ & new_G4431_;
  assign new_G4515_ = ~new_G4454_;
  assign new_G4516_ = ~new_G4456_;
  assign new_G4517_ = new_G4303_ & new_G4453_;
  assign new_G4518_ = new_G4303_ & new_G4455_;
  assign new_G4519_ = new_G4303_ & new_G4457_;
  assign new_G4520_ = new_G4378_ & new_G1248_ & new_G1981_;
  assign new_G4521_ = new_G4400_ & new_G1264_ & new_G2003_;
  assign new_G4522_ = ~new_G4417_;
  assign new_G4523_ = ~new_G4420_;
  assign new_G4524_ = ~new_G4420_ | ~new_G4333_;
  assign new_G4525_ = ~new_G2945_ | ~new_G4476_;
  assign new_G4526_ = ~new_G3215_ | ~new_G4478_;
  assign new_G4527_ = ~new_G2984_ | ~new_G4488_;
  assign new_G4528_ = ~new_G3247_ | ~new_G4490_;
  assign new_G4529_ = ~new_G4161_ | ~new_G4492_;
  assign new_G4530_ = ~new_G4446_;
  assign new_G4531_ = ~new_G4443_;
  assign new_G4532_ = ~new_G4440_;
  assign new_G4533_ = ~new_G4437_;
  assign new_G4534_ = ~new_G4469_;
  assign new_G4535_ = ~new_G4466_;
  assign new_G4536_ = ~new_G4463_;
  assign new_G4537_ = new_G4510_ & new_G4432_;
  assign new_G4538_ = new_G4511_ & new_G4432_;
  assign new_G4539_ = new_G4386_ & new_G4432_;
  assign new_G4540_ = new_G3415_ & new_G4432_;
  assign new_G4541_ = ~new_G4450_;
  assign new_G4542_ = new_G4515_ & new_G4458_;
  assign new_G4543_ = new_G4516_ & new_G4458_;
  assign new_G4544_ = new_G4396_ & new_G4458_;
  assign new_G4545_ = new_G3570_ & new_G4458_;
  assign new_G4546_ = ~new_G4473_;
  assign new_G4547_ = ~new_G4498_;
  assign new_G4548_ = ~new_G4498_ | ~new_G4407_;
  assign new_G4549_ = ~new_G4501_;
  assign new_G4550_ = ~new_G4501_ | ~new_G4408_;
  assign new_G4551_ = new_G4446_ & new_G1248_ & new_G1981_;
  assign new_G4552_ = new_G4443_ & new_G1248_ & new_G1981_;
  assign new_G4553_ = new_G4440_ & new_G1248_ & new_G1981_;
  assign new_G4554_ = new_G2320_ | new_G3068_ | new_G4520_;
  assign new_G4560_ = new_G4469_ & new_G1264_ & new_G2003_;
  assign new_G4561_ = new_G4466_ & new_G1264_ & new_G2003_;
  assign new_G4562_ = new_G2325_ | new_G3072_ | new_G4521_;
  assign new_G4568_ = ~new_G4504_ | ~new_G4522_;
  assign new_G4569_ = ~new_G4504_;
  assign new_G4570_ = ~new_G4180_ | ~new_G4523_;
  assign new_G4571_ = new_G4437_ & new_G1280_ & new_G2031_;
  assign new_G4572_ = new_G4463_ & new_G1294_ & new_G2053_;
  assign new_G4573_ = ~new_G4477_ | ~new_G4525_;
  assign new_G4576_ = ~new_G4479_ | ~new_G4526_;
  assign new_G4579_ = ~new_G4480_;
  assign new_G4580_ = ~new_G4480_ | ~new_G4483_;
  assign new_G4581_ = ~new_G4484_;
  assign new_G4582_ = ~new_G4484_ | ~new_G4487_;
  assign new_G4583_ = ~new_G4489_ | ~new_G4527_;
  assign new_G4586_ = ~new_G4491_ | ~new_G4528_;
  assign new_G4589_ = ~new_G4493_ | ~new_G4529_;
  assign new_G4592_ = ~new_G4494_;
  assign new_G4593_ = ~new_G4494_ | ~new_G4497_;
  assign new_G4594_ = new_G4537_ | new_G4512_;
  assign new_G4597_ = new_G4538_ | new_G4513_;
  assign new_G4600_ = new_G4539_ | new_G4514_;
  assign new_G4603_ = new_G4540_ | new_G4449_;
  assign new_G4606_ = new_G4542_ | new_G4517_;
  assign new_G4613_ = new_G4543_ | new_G4518_;
  assign new_G4616_ = new_G4544_ | new_G4519_;
  assign new_G4619_ = new_G4545_ | new_G4472_;
  assign new_G4622_ = ~new_G4254_ | ~new_G4547_;
  assign new_G4623_ = ~new_G4257_ | ~new_G4549_;
  assign new_G4624_ = new_G2321_ | new_G3069_ | new_G4551_;
  assign new_G4630_ = new_G2322_ | new_G3070_ | new_G4552_;
  assign new_G4636_ = new_G2323_ | new_G3071_ | new_G4553_;
  assign new_G4642_ = new_G2326_ | new_G3073_ | new_G4560_;
  assign new_G4648_ = new_G2327_ | new_G2516_ | new_G4561_;
  assign new_G4654_ = ~new_G4417_ | ~new_G4569_;
  assign new_G4655_ = ~new_G4570_ | ~new_G4524_;
  assign new_G4658_ = new_G2339_ | new_G3086_ | new_G4571_;
  assign new_G4664_ = new_G2344_ | new_G3090_ | new_G4572_;
  assign new_G4670_ = ~new_G4346_ | ~new_G4579_;
  assign new_G4671_ = ~new_G4352_ | ~new_G4581_;
  assign new_G4672_ = ~new_G4371_ | ~new_G4592_;
  assign new_G4673_ = new_G4554_ & new_G718_ & new_G1565_;
  assign new_G4674_ = new_G4562_ & new_G1554_ & new_G1565_;
  assign new_G4675_ = new_G4554_ & new_G780_ & new_G1640_;
  assign new_G4676_ = new_G4562_ & new_G1629_ & new_G1640_;
  assign new_G4677_ = new_G4554_ & new_G860_ & new_G1663_;
  assign new_G4678_ = new_G4562_ & new_G1652_ & new_G1663_;
  assign new_G4679_ = new_G4562_ & new_G1674_ & new_G1685_;
  assign new_G4680_ = new_G4554_ & new_G884_ & new_G1685_;
  assign new_G4681_ = ~new_G4622_ | ~new_G4548_;
  assign new_G4684_ = ~new_G4623_ | ~new_G4550_;
  assign new_G4687_ = ~new_G4568_ | ~new_G4654_;
  assign new_G4690_ = ~new_G4573_;
  assign new_G4691_ = ~new_G4573_ | ~new_G4339_;
  assign new_G4692_ = ~new_G4576_;
  assign new_G4693_ = ~new_G4576_ | ~new_G4343_;
  assign new_G4694_ = ~new_G4670_ | ~new_G4580_;
  assign new_G4697_ = ~new_G4671_ | ~new_G4582_;
  assign new_G4700_ = ~new_G4583_;
  assign new_G4701_ = ~new_G4583_ | ~new_G4359_;
  assign new_G4702_ = ~new_G4586_;
  assign new_G4703_ = ~new_G4586_ | ~new_G4363_;
  assign new_G4704_ = ~new_G4589_;
  assign new_G4705_ = ~new_G4589_ | ~new_G4368_;
  assign new_G4706_ = ~new_G4672_ | ~new_G4593_;
  assign new_G4709_ = ~new_G4603_;
  assign new_G4710_ = ~new_G4600_;
  assign new_G4711_ = ~new_G4597_;
  assign new_G4712_ = ~new_G4594_;
  assign new_G4713_ = ~new_G4619_;
  assign new_G4714_ = ~new_G4616_;
  assign new_G4715_ = ~new_G4613_;
  assign new_G4716_ = ~new_G4606_;
  assign new_G4717_ = new_G4664_ & new_G1526_ & new_G1537_;
  assign new_G4718_ = new_G4658_ & new_G694_ & new_G1537_;
  assign new_G4719_ = new_G1465_ | new_G2162_ | new_G4423_ | new_G4673_;
  assign new_G4720_ = new_G4624_ & new_G718_ & new_G1565_;
  assign new_G4721_ = new_G4642_ & new_G1554_ & new_G1565_;
  assign new_G4722_ = new_G4630_ & new_G718_ & new_G1565_;
  assign new_G4723_ = new_G4648_ & new_G1554_ & new_G1565_;
  assign new_G4724_ = new_G4636_ & new_G718_ & new_G1565_;
  assign new_G4725_ = new_G4664_ & new_G1601_ & new_G1612_;
  assign new_G4726_ = new_G4658_ & new_G756_ & new_G1612_;
  assign new_G4727_ = new_G1474_ | new_G2173_ | new_G4424_ | new_G4675_;
  assign new_G4728_ = new_G4624_ & new_G780_ & new_G1640_;
  assign new_G4729_ = new_G4642_ & new_G1629_ & new_G1640_;
  assign new_G4730_ = new_G4630_ & new_G780_ & new_G1640_;
  assign new_G4731_ = new_G4648_ & new_G1629_ & new_G1640_;
  assign new_G4732_ = new_G4636_ & new_G780_ & new_G1640_;
  assign new_G4733_ = new_G4664_ & new_G1914_ & new_G1925_;
  assign new_G4734_ = new_G4658_ & new_G1184_ & new_G1925_;
  assign new_G4735_ = new_G4648_ & new_G1652_ & new_G1663_;
  assign new_G4736_ = new_G4636_ & new_G860_ & new_G1663_;
  assign new_G4737_ = new_G4642_ & new_G1652_ & new_G1663_;
  assign new_G4738_ = new_G4630_ & new_G860_ & new_G1663_;
  assign new_G4739_ = new_G4624_ & new_G860_ & new_G1663_;
  assign new_G4740_ = new_G4664_ & new_G1948_ & new_G1959_;
  assign new_G4741_ = new_G4658_ & new_G1218_ & new_G1959_;
  assign new_G4742_ = new_G4648_ & new_G1674_ & new_G1685_;
  assign new_G4743_ = new_G4636_ & new_G884_ & new_G1685_;
  assign new_G4744_ = new_G4642_ & new_G1674_ & new_G1685_;
  assign new_G4745_ = new_G4630_ & new_G884_ & new_G1685_;
  assign new_G4746_ = new_G4624_ & new_G884_ & new_G1685_;
  assign new_G4747_ = new_G4606_ & n4659_lo & n4647_lo;
  assign new_G4748_ = ~new_G4655_;
  assign new_G4749_ = new_G4655_ & new_G1941_;
  assign new_G4750_ = new_G4603_ & new_G1280_ & new_G2031_;
  assign new_G4751_ = new_G4600_ & new_G1280_ & new_G2031_;
  assign new_G4752_ = new_G4597_ & new_G1280_ & new_G2031_;
  assign new_G4753_ = new_G4594_ & new_G1280_ & new_G2031_;
  assign new_G4754_ = new_G4619_ & new_G1294_ & new_G2053_;
  assign new_G4755_ = new_G4616_ & new_G1294_ & new_G2053_;
  assign new_G4756_ = new_G4613_ & new_G1294_ & new_G2053_;
  assign new_G4757_ = new_G4606_ & new_G1294_ & new_G2053_;
  assign new_G4758_ = ~new_G4409_ | ~new_G4606_;
  assign new_G4761_ = ~new_G4116_ | ~new_G4690_;
  assign new_G4762_ = ~new_G4119_ | ~new_G4692_;
  assign new_G4763_ = ~new_G4155_ | ~new_G4700_;
  assign new_G4764_ = ~new_G4158_ | ~new_G4702_;
  assign new_G4765_ = ~new_G4164_ | ~new_G4704_;
  assign new_G4766_ = new_G1460_ | new_G2157_ | new_G4717_ | new_G4718_;
  assign new_G4767_ = new_G1466_ | new_G2163_ | new_G4674_ | new_G4720_;
  assign new_G4768_ = new_G1467_ | new_G2164_ | new_G4721_ | new_G4722_;
  assign new_G4769_ = new_G1468_ | new_G2165_ | new_G4723_ | new_G4724_;
  assign new_G4770_ = new_G1469_ | new_G2168_ | new_G4725_ | new_G4726_;
  assign new_G4771_ = new_G1475_ | new_G2174_ | new_G4676_ | new_G4728_;
  assign new_G4772_ = new_G1476_ | new_G2175_ | new_G4729_ | new_G4730_;
  assign new_G4773_ = new_G1477_ | new_G2176_ | new_G4731_ | new_G4732_;
  assign new_G4774_ = new_G4747_ | new_G1497_ | new_G3055_ | new_G4509_;
  assign new_G4775_ = new_G4748_ & new_G1992_ & new_G2003_;
  assign new_G4776_ = ~new_G4681_;
  assign new_G4777_ = ~new_G4684_;
  assign new_G4778_ = ~new_G4687_;
  assign new_G4779_ = new_G4687_ & new_G1941_;
  assign new_G4780_ = new_G2340_ | new_G3087_ | new_G4750_;
  assign new_G4786_ = new_G2341_ | new_G3088_ | new_G4751_;
  assign new_G4792_ = new_G2342_ | new_G3089_ | new_G4752_;
  assign new_G4798_ = new_G2343_ | new_G3207_ | new_G4753_;
  assign new_G4804_ = new_G2345_ | new_G3091_ | new_G4754_;
  assign new_G4810_ = new_G2346_ | new_G3092_ | new_G4755_;
  assign new_G4816_ = new_G2347_ | new_G2887_ | new_G4756_;
  assign new_G4822_ = new_G2348_ | new_G3093_ | new_G4757_;
  assign new_G4828_ = ~new_G4761_ | ~new_G4691_;
  assign new_G4831_ = ~new_G4762_ | ~new_G4693_;
  assign new_G4834_ = ~new_G4694_;
  assign new_G4835_ = ~new_G4694_ | ~new_G4349_;
  assign new_G4836_ = ~new_G4697_;
  assign new_G4837_ = ~new_G4697_ | ~new_G4355_;
  assign new_G4838_ = ~new_G4763_ | ~new_G4701_;
  assign new_G4841_ = ~new_G4764_ | ~new_G4703_;
  assign new_G4844_ = ~new_G4765_ | ~new_G4705_;
  assign new_G4847_ = ~new_G4706_;
  assign new_G4848_ = ~new_G4706_ | ~new_G4374_;
  assign new_G4849_ = new_G4409_ & new_G4758_;
  assign new_G4850_ = new_G4758_ & new_G4606_;
  assign new_G4851_ = new_G4264_ & n4479_lo & new_G4776_ & new_G4777_ & new_G4377_;
  assign new_G4852_ = new_G4778_ & new_G1970_ & new_G1981_;
  assign new_G4853_ = ~new_G4125_ | ~new_G4834_;
  assign new_G4854_ = ~new_G4131_ | ~new_G4836_;
  assign new_G4855_ = ~new_G4170_ | ~new_G4847_;
  assign new_G4856_ = new_G4804_ & new_G1526_ & new_G1537_;
  assign new_G4857_ = new_G4780_ & new_G694_ & new_G1537_;
  assign new_G4858_ = new_G4810_ & new_G1526_ & new_G1537_;
  assign new_G4859_ = new_G4786_ & new_G694_ & new_G1537_;
  assign new_G4860_ = new_G4816_ & new_G1526_ & new_G1537_;
  assign new_G4861_ = new_G4792_ & new_G694_ & new_G1537_;
  assign new_G4862_ = new_G4822_ & new_G1526_ & new_G1537_;
  assign new_G4863_ = new_G4798_ & new_G694_ & new_G1537_;
  assign new_G4864_ = new_G4804_ & new_G1601_ & new_G1612_;
  assign new_G4865_ = new_G4780_ & new_G756_ & new_G1612_;
  assign new_G4866_ = new_G4810_ & new_G1601_ & new_G1612_;
  assign new_G4867_ = new_G4786_ & new_G756_ & new_G1612_;
  assign new_G4868_ = new_G4816_ & new_G1601_ & new_G1612_;
  assign new_G4869_ = new_G4792_ & new_G756_ & new_G1612_;
  assign new_G4870_ = new_G4822_ & new_G1601_ & new_G1612_;
  assign new_G4871_ = new_G4798_ & new_G756_ & new_G1612_;
  assign new_G4872_ = new_G4822_ & new_G1948_ & new_G1959_;
  assign new_G4873_ = new_G4798_ & new_G1218_ & new_G1959_;
  assign new_G4874_ = new_G4822_ & new_G1914_ & new_G1925_;
  assign new_G4875_ = new_G4798_ & new_G1184_ & new_G1925_;
  assign new_G4876_ = new_G4816_ & new_G1914_ & new_G1925_;
  assign new_G4877_ = new_G4792_ & new_G1184_ & new_G1925_;
  assign new_G4878_ = new_G4810_ & new_G1914_ & new_G1925_;
  assign new_G4879_ = new_G4786_ & new_G1184_ & new_G1925_;
  assign new_G4880_ = new_G4804_ & new_G1914_ & new_G1925_;
  assign new_G4881_ = new_G4780_ & new_G1184_ & new_G1925_;
  assign new_G4882_ = new_G4816_ & new_G1948_ & new_G1959_;
  assign new_G4883_ = new_G4792_ & new_G1218_ & new_G1959_;
  assign new_G4884_ = new_G4810_ & new_G1948_ & new_G1959_;
  assign new_G4885_ = new_G4786_ & new_G1218_ & new_G1959_;
  assign new_G4886_ = new_G4804_ & new_G1948_ & new_G1959_;
  assign new_G4887_ = new_G4780_ & new_G1218_ & new_G1959_;
  assign new_G4888_ = ~new_G4828_;
  assign new_G4889_ = ~new_G4828_ | ~new_G4230_;
  assign new_G4890_ = ~new_G4831_;
  assign new_G4891_ = ~new_G4831_ | ~new_G4233_;
  assign new_G4892_ = ~new_G4853_ | ~new_G4835_;
  assign new_G4895_ = ~new_G4854_ | ~new_G4837_;
  assign new_G4898_ = ~new_G4838_;
  assign new_G4899_ = ~new_G4838_ | ~new_G4244_;
  assign new_G4900_ = ~new_G4841_;
  assign new_G4901_ = ~new_G4841_ | ~new_G4246_;
  assign new_G4902_ = ~new_G4844_;
  assign new_G4903_ = ~new_G4844_ | ~new_G3694_;
  assign new_G4904_ = ~new_G4855_ | ~new_G4848_;
  assign new_G4907_ = new_G1461_ | new_G2158_ | new_G4856_ | new_G4857_;
  assign new_G4908_ = new_G1462_ | new_G2159_ | new_G4858_ | new_G4859_;
  assign new_G4909_ = new_G1463_ | new_G2160_ | new_G4860_ | new_G4861_;
  assign new_G4910_ = new_G1464_ | new_G2161_ | new_G4862_ | new_G4863_;
  assign new_G4911_ = new_G1470_ | new_G2169_ | new_G4864_ | new_G4865_;
  assign new_G4912_ = new_G1471_ | new_G2170_ | new_G4866_ | new_G4867_;
  assign new_G4913_ = new_G1472_ | new_G2171_ | new_G4868_ | new_G4869_;
  assign new_G4914_ = new_G1473_ | new_G2172_ | new_G4870_ | new_G4871_;
  assign new_G4915_ = ~new_G3939_ | ~new_G4888_;
  assign new_G4916_ = ~new_G3951_ | ~new_G4890_;
  assign new_G4917_ = ~new_G4008_ | ~new_G4898_;
  assign new_G4918_ = ~new_G4014_ | ~new_G4900_;
  assign new_G4919_ = ~new_G3256_ | ~new_G4902_;
  assign new_G4920_ = ~new_G4915_ | ~new_G4889_;
  assign new_G4923_ = ~new_G4916_ | ~new_G4891_;
  assign new_G4926_ = ~new_G4892_;
  assign new_G4927_ = ~new_G4892_ | ~new_G4236_;
  assign new_G4928_ = ~new_G4895_;
  assign new_G4929_ = ~new_G4895_ | ~new_G4241_;
  assign new_G4930_ = ~new_G4917_ | ~new_G4899_;
  assign new_G4933_ = ~new_G4918_ | ~new_G4901_;
  assign new_G4936_ = ~new_G4919_ | ~new_G4903_;
  assign new_G4939_ = ~new_G4904_;
  assign new_G4940_ = ~new_G4904_ | ~new_G3696_;
  assign new_G4941_ = ~new_G3963_ | ~new_G4926_;
  assign new_G4942_ = ~new_G3981_ | ~new_G4928_;
  assign new_G4943_ = ~new_G3262_ | ~new_G4939_;
  assign new_G4944_ = ~new_G4920_;
  assign new_G4945_ = ~new_G4920_ | ~new_G4231_;
  assign new_G4946_ = ~new_G4923_;
  assign new_G4947_ = ~new_G4923_ | ~new_G4234_;
  assign new_G4948_ = ~new_G4941_ | ~new_G4927_;
  assign new_G4951_ = ~new_G4942_ | ~new_G4929_;
  assign new_G4954_ = ~new_G4930_;
  assign new_G4955_ = ~new_G4930_ | ~new_G4245_;
  assign new_G4956_ = ~new_G4933_;
  assign new_G4957_ = ~new_G4933_ | ~new_G4247_;
  assign new_G4958_ = ~new_G4936_;
  assign new_G4959_ = ~new_G4936_ | ~new_G4248_;
  assign new_G4960_ = ~new_G4943_ | ~new_G4940_;
  assign new_G4963_ = ~new_G3942_ | ~new_G4944_;
  assign new_G4964_ = ~new_G3954_ | ~new_G4946_;
  assign new_G4965_ = ~new_G4011_ | ~new_G4954_;
  assign new_G4966_ = ~new_G4017_ | ~new_G4956_;
  assign new_G4967_ = ~new_G4020_ | ~new_G4958_;
  assign new_G4968_ = ~new_G4963_ | ~new_G4945_;
  assign new_G4971_ = ~new_G4964_ | ~new_G4947_;
  assign new_G4974_ = ~new_G4948_;
  assign new_G4975_ = ~new_G4948_ | ~new_G4237_;
  assign new_G4976_ = ~new_G4951_;
  assign new_G4977_ = ~new_G4951_ | ~new_G4242_;
  assign new_G4978_ = ~new_G4965_ | ~new_G4955_;
  assign new_G4981_ = ~new_G4966_ | ~new_G4957_;
  assign new_G4984_ = ~new_G4967_ | ~new_G4959_;
  assign new_G4987_ = ~new_G4960_;
  assign new_G4988_ = ~new_G4960_ | ~new_G4252_;
  assign new_G4989_ = ~new_G3966_ | ~new_G4974_;
  assign new_G4990_ = ~new_G3984_ | ~new_G4976_;
  assign new_G4991_ = ~new_G4029_ | ~new_G4987_;
  assign new_G4992_ = ~new_G4968_;
  assign new_G4993_ = ~new_G4968_ | ~new_G4232_;
  assign new_G4994_ = ~new_G4971_;
  assign new_G4995_ = ~new_G4971_ | ~new_G4235_;
  assign new_G4996_ = ~new_G4989_ | ~new_G4975_;
  assign new_G4999_ = ~new_G4990_ | ~new_G4977_;
  assign new_G5002_ = ~new_G4978_;
  assign new_G5003_ = ~new_G4978_ | ~new_G3691_;
  assign new_G5004_ = ~new_G4981_;
  assign new_G5005_ = ~new_G4981_ | ~new_G3693_;
  assign new_G5006_ = ~new_G4984_;
  assign new_G5007_ = ~new_G4984_ | ~new_G4249_;
  assign new_G5008_ = ~new_G4991_ | ~new_G4988_;
  assign new_G5011_ = ~new_G3945_ | ~new_G4992_;
  assign new_G5012_ = ~new_G3957_ | ~new_G4994_;
  assign new_G5013_ = ~new_G3241_ | ~new_G5002_;
  assign new_G5014_ = ~new_G3250_ | ~new_G5004_;
  assign new_G5015_ = ~new_G4023_ | ~new_G5006_;
  assign new_G5016_ = ~new_G5011_ | ~new_G4993_;
  assign new_G5019_ = ~new_G5012_ | ~new_G4995_;
  assign new_G5022_ = ~new_G4996_;
  assign new_G5023_ = ~new_G4996_ | ~new_G4238_;
  assign new_G5024_ = ~new_G4999_;
  assign new_G5025_ = ~new_G4999_ | ~new_G4243_;
  assign new_G5026_ = ~new_G5013_ | ~new_G5003_;
  assign new_G5029_ = ~new_G5014_ | ~new_G5005_;
  assign new_G5032_ = ~new_G5015_ | ~new_G5007_;
  assign new_G5035_ = ~new_G5008_;
  assign new_G5036_ = ~new_G5008_ | ~new_G4253_;
  assign new_G5037_ = ~new_G3969_ | ~new_G5022_;
  assign new_G5038_ = ~new_G3987_ | ~new_G5024_;
  assign new_G5039_ = ~new_G4032_ | ~new_G5035_;
  assign new_G5040_ = ~new_G5016_;
  assign new_G5041_ = ~new_G5016_ | ~new_G4200_;
  assign new_G5042_ = ~new_G5019_;
  assign new_G5043_ = ~new_G5019_ | ~new_G4201_;
  assign new_G5044_ = ~new_G5026_;
  assign new_G5045_ = ~new_G5026_ | ~new_G3664_;
  assign new_G5046_ = ~new_G5029_;
  assign new_G5047_ = ~new_G5029_ | ~new_G3665_;
  assign new_G5048_ = ~new_G5037_ | ~new_G5023_;
  assign new_G5051_ = ~new_G5038_ | ~new_G5025_;
  assign new_G5054_ = ~new_G5032_;
  assign new_G5055_ = ~new_G5032_ | ~new_G4250_;
  assign new_G5056_ = ~new_G5039_ | ~new_G5036_;
  assign new_G5059_ = ~new_G3948_ | ~new_G5040_;
  assign new_G5060_ = ~new_G3960_ | ~new_G5042_;
  assign new_G5061_ = ~new_G3244_ | ~new_G5044_;
  assign new_G5062_ = ~new_G3253_ | ~new_G5046_;
  assign new_G5063_ = ~new_G4026_ | ~new_G5054_;
  assign new_G5064_ = ~new_G5059_ | ~new_G5041_;
  assign new_G5067_ = ~new_G5060_ | ~new_G5043_;
  assign new_G5070_ = ~new_G5061_ | ~new_G5045_;
  assign new_G5073_ = ~new_G5062_ | ~new_G5047_;
  assign new_G5076_ = ~new_G5048_;
  assign new_G5077_ = ~new_G5048_ | ~new_G4239_;
  assign new_G5078_ = ~new_G5051_;
  assign new_G5079_ = ~new_G5051_ | ~new_G4240_;
  assign new_G5080_ = ~new_G5063_ | ~new_G5055_;
  assign new_G5083_ = ~new_G5056_;
  assign new_G5084_ = ~new_G5056_ | ~new_G4251_;
  assign new_G5085_ = ~new_G3972_ | ~new_G5076_;
  assign new_G5086_ = ~new_G3990_ | ~new_G5078_;
  assign new_G5087_ = ~new_G4035_ | ~new_G5083_;
  assign new_G5088_ = new_G5067_ & new_G4290_ & new_G690_;
  assign new_G5089_ = new_G5064_ & new_G4054_ & new_G690_;
  assign new_G5090_ = new_G5067_ & new_G4450_ & n4491_lo;
  assign new_G5091_ = new_G5064_ & new_G4541_ & n4491_lo;
  assign new_G5092_ = ~new_G5080_;
  assign new_G5093_ = ~new_G5080_ | ~new_G4075_;
  assign new_G5094_ = new_G5073_ & new_G4316_ & new_G752_;
  assign new_G5095_ = new_G5070_ & new_G4068_ & new_G752_;
  assign new_G5096_ = new_G5073_ & new_G4473_ & n4551_lo;
  assign new_G5097_ = new_G5070_ & new_G4546_ & n4551_lo;
  assign new_G5098_ = ~new_G5085_ | ~new_G5077_;
  assign new_G5101_ = ~new_G5086_ | ~new_G5079_;
  assign new_G5104_ = ~new_G5087_ | ~new_G5084_;
  assign new_G5107_ = ~new_G3745_ | ~new_G5092_;
  assign new_G5108_ = new_G5091_ | new_G5090_ | new_G5088_ | new_G5089_;
  assign new_G5111_ = new_G5097_ | new_G5096_ | new_G5094_ | new_G5095_;
  assign new_G5114_ = ~new_G5098_;
  assign new_G5115_ = ~new_G5098_ | ~new_G4202_;
  assign new_G5116_ = ~new_G5101_;
  assign new_G5117_ = ~new_G5101_ | ~new_G4203_;
  assign new_G5118_ = ~new_G5107_ | ~new_G5093_;
  assign new_G5119_ = ~new_G5104_;
  assign new_G5120_ = ~new_G5104_ | ~new_G4076_;
  assign new_G5121_ = ~new_G3975_ | ~new_G5114_;
  assign new_G5122_ = ~new_G3978_ | ~new_G5116_;
  assign new_G5123_ = ~new_G5108_;
  assign new_G5124_ = ~new_G3748_ | ~new_G5119_;
  assign new_G5125_ = n4551_lo & new_G5118_;
  assign new_G5126_ = ~new_G5111_;
  assign new_G5127_ = ~new_G5121_ | ~new_G5115_;
  assign new_G5128_ = ~new_G5122_ | ~new_G5117_;
  assign new_G5129_ = ~new_G5124_ | ~new_G5120_;
  assign new_G5130_ = ~new_G5128_;
  assign new_G5131_ = n4491_lo & new_G5127_;
  assign new_G5132_ = ~new_G5129_;
  assign new_G5133_ = new_G5130_ & new_G690_;
  assign new_G5134_ = new_G5132_ & new_G752_;
  assign new_G5135_ = new_G5133_ | new_G5131_;
  assign new_G5138_ = new_G5134_ | new_G5125_;
  assign new_G5141_ = ~new_G5135_ | ~new_G5123_;
  assign new_G5142_ = ~new_G5135_;
  assign new_G5143_ = ~new_G5138_ | ~new_G5126_;
  assign new_G5144_ = ~new_G5138_;
  assign new_G5145_ = ~new_G5108_ | ~new_G5142_;
  assign new_G5146_ = ~new_G5111_ | ~new_G5144_;
  assign new_G5147_ = ~new_G5141_ | ~new_G5145_;
  assign new_G5150_ = ~new_G5143_ | ~new_G5146_;
  assign new_G5153_ = new_G5150_ & new_G1264_ & new_G2003_;
  assign new_G5154_ = new_G5147_ & new_G1248_ & new_G1981_;
  assign new_G5155_ = ~new_G5147_;
  assign new_G5156_ = ~new_G5150_;
  assign new_G5157_ = new_G5155_ & new_G1214_;
  assign new_G5158_ = new_G5156_ & new_G1214_;
  assign new_G5159_ = new_G4779_ | new_G5157_;
  assign new_G5162_ = new_G4749_ | new_G5158_;
  assign new_G5165_ = new_G5159_ & new_G1936_;
  assign new_G5166_ = new_G5162_ & new_G1936_;
  assign new_G5167_ = new_G5159_ & new_G1936_;
  assign new_G5168_ = new_G5162_ & new_G1936_;
  assign new_G5169_ = new_G5165_ | new_G1944_;
  assign new_G5172_ = new_G5166_ | new_G1945_;
  assign new_G5175_ = new_G5167_ | new_G1946_;
  assign new_G5178_ = new_G5168_ | new_G1947_;
  assign new_G5181_ = new_G5178_ & new_G1652_ & new_G1663_;
  assign new_G5182_ = new_G5175_ & new_G860_ & new_G1663_;
  assign new_G5183_ = new_G5178_ & new_G1674_ & new_G1685_;
  assign new_G5184_ = new_G5175_ & new_G884_ & new_G1685_;
  assign new_G5185_ = new_G5172_ & new_G1554_ & new_G1565_;
  assign new_G5186_ = new_G5169_ & new_G718_ & new_G1565_;
  assign new_G5187_ = new_G5172_ & new_G1629_ & new_G1640_;
  assign new_G5188_ = new_G5169_ & new_G780_ & new_G1640_;
  assign new_G5189_ = new_G1576_ | new_G2203_ | new_G5185_ | new_G5186_;
  assign new_G5190_ = new_G1651_ | new_G2204_ | new_G5187_ | new_G5188_;
  assign new_G5191_ = new_G5189_ & new_G1548_;
  assign new_G5192_ = new_G5190_ & new_G1623_;
  assign G5193 = ~n3399_lo;
  assign G5194 = ~n3963_lo;
  assign G5195 = ~n4587_lo;
  assign G5196 = ~n4419_lo;
  assign G5197 = ~n4131_lo;
  assign G5198 = ~n4179_lo;
  assign G5199 = n4443_lo & n4479_lo;
  assign G5200 = ~n4431_lo;
  assign G5201 = G5196;
  assign G5202 = G5196;
  assign G5203 = ~n4107_lo;
  assign G5204 = ~n4155_lo;
  assign G5205 = n3399_lo & n3411_lo;
  assign G5206 = ~n3795_lo;
  assign G5207 = ~n4443_lo;
  assign G5208 = ~n4479_lo;
  assign G5209 = ~n4467_lo;
  assign G5210 = ~new_G684_;
  assign G5211 = n3363_lo & new_G685_;
  assign G5212 = ~new_G687_;
  assign G5213 = ~new_G688_;
  assign G5214 = ~new_G742_;
  assign G5215 = ~new_G749_;
  assign G5216 = ~new_G980_;
  assign G5217 = ~new_G1067_;
  assign G5218 = ~new_G1308_;
  assign G5219 = G5217;
  assign G5220 = ~new_G976_ | ~n3387_lo;
  assign G5221 = ~new_G976_;
  assign G5222 = ~new_G1577_;
  assign G5223 = G5222;
  assign G5224 = G5222;
  assign G5225 = G5222;
  assign G5226 = ~new_G2064_;
  assign G5227 = G5226;
  assign G5228 = ~new_G2528_;
  assign G5229 = ~new_G2533_;
  assign G5230 = ~new_G2538_;
  assign G5231 = ~new_G2539_;
  assign G5232 = new_G2671_ & new_G1750_;
  assign G5233 = new_G2672_ & new_G1750_;
  assign G5234 = new_G2673_ & new_G1750_;
  assign G5235 = new_G2674_ & new_G1750_;
  assign G5236 = new_G3105_ & new_G3106_ & new_G2669_;
  assign G5237 = new_G3107_ & new_G3108_ & new_G3281_;
  assign G5238 = new_G3793_ & new_G3802_;
  assign G5239 = new_G3825_ & new_G3834_;
  assign G5240 = new_G3852_ & new_G3859_;
  assign G5241 = new_G3765_ & new_G3776_;
  assign G5242 = ~new_G4077_;
  assign G5243 = ~new_G4227_;
  assign G5244 = new_G4044_ | new_G4260_;
  assign G5245 = new_G4045_ | new_G4261_;
  assign G5246 = new_G4046_ | new_G4262_;
  assign G5247 = new_G4047_ | new_G4263_;
  assign G5248 = ~new_G4323_;
  assign G5249 = ~new_G4562_;
  assign G5250 = ~new_G4554_;
  assign G5251 = ~new_G4606_;
  assign G5252 = new_G1479_ | new_G2182_ | new_G4425_ | new_G4677_;
  assign G5253 = ~new_G4664_;
  assign G5254 = ~new_G4648_;
  assign G5255 = ~new_G4642_;
  assign G5256 = new_G1499_ | new_G2201_ | new_G4426_ | new_G4680_;
  assign G5257 = ~new_G4658_;
  assign G5258 = ~new_G4636_;
  assign G5259 = ~new_G4630_;
  assign G5260 = ~new_G4624_;
  assign G5261 = ~new_G4681_;
  assign G5262 = ~new_G4684_;
  assign G5263 = new_G4712_ & new_G4711_ & new_G4710_ & new_G4532_ & new_G4507_ & new_G4530_ & new_G4531_ & new_G4533_ & new_G4709_;
  assign G5264 = new_G4716_ & new_G4715_ & new_G4714_ & new_G4535_ & new_G4183_ & new_G4508_ & new_G4534_ & new_G4536_ & new_G4713_;
  assign G5265 = new_G4719_ & new_G1548_;
  assign G5266 = new_G4727_ & new_G1623_;
  assign G5267 = new_G1484_ | new_G2187_ | new_G4733_ | new_G4734_;
  assign G5268 = new_G1485_ | new_G2188_ | new_G4735_ | new_G4736_;
  assign G5269 = new_G1486_ | new_G2189_ | new_G4737_ | new_G4738_;
  assign G5270 = new_G1487_ | new_G2190_ | new_G4678_ | new_G4739_;
  assign G5271 = new_G1492_ | new_G2195_ | new_G4740_ | new_G4741_;
  assign G5272 = new_G1493_ | new_G2196_ | new_G4742_ | new_G4743_;
  assign G5273 = new_G1494_ | new_G2197_ | new_G4744_ | new_G4745_;
  assign G5274 = new_G1495_ | new_G2198_ | new_G4679_ | new_G4746_;
  assign G5275 = new_G4766_ & new_G1520_;
  assign G5276 = new_G4767_ & new_G1548_;
  assign G5277 = new_G4768_ & new_G1548_;
  assign G5278 = new_G4769_ & new_G1548_;
  assign G5279 = new_G4770_ & new_G1595_;
  assign G5280 = new_G4771_ & new_G1623_;
  assign G5281 = new_G4772_ & new_G1623_;
  assign G5282 = new_G4773_ & new_G1623_;
  assign G5283 = new_G686_ & new_G4774_;
  assign G5284 = new_G4849_ | new_G4850_;
  assign G5285 = ~new_G4822_;
  assign G5286 = ~new_G4816_;
  assign G5287 = ~new_G4810_;
  assign G5288 = ~new_G4804_;
  assign G5289 = new_G689_ & new_G4851_ & n3795_lo;
  assign G5290 = ~new_G4798_;
  assign G5291 = ~new_G4792_;
  assign G5292 = ~new_G4786_;
  assign G5293 = ~new_G4780_;
  assign G5294 = new_G1478_ | new_G2179_ | new_G4872_ | new_G4873_;
  assign G5295 = new_G1480_ | new_G2183_ | new_G4874_ | new_G4875_;
  assign G5296 = new_G1481_ | new_G2184_ | new_G4876_ | new_G4877_;
  assign G5297 = new_G1482_ | new_G2185_ | new_G4878_ | new_G4879_;
  assign G5298 = new_G1483_ | new_G2186_ | new_G4880_ | new_G4881_;
  assign G5299 = new_G1489_ | new_G2192_ | new_G4882_ | new_G4883_;
  assign G5300 = new_G1490_ | new_G2193_ | new_G4884_ | new_G4885_;
  assign G5301 = new_G1491_ | new_G2194_ | new_G4886_ | new_G4887_;
  assign G5302 = new_G4907_ & new_G1520_;
  assign G5303 = new_G4908_ & new_G1520_;
  assign G5304 = new_G4909_ & new_G1520_;
  assign G5305 = new_G4910_ & new_G1520_;
  assign G5306 = new_G4911_ & new_G1595_;
  assign G5307 = new_G4912_ & new_G1595_;
  assign G5308 = new_G4913_ & new_G1595_;
  assign G5309 = new_G4914_ & new_G1595_;
  assign G5310 = new_G1498_ | new_G2200_ | new_G4775_ | new_G5153_;
  assign G5311 = new_G1500_ | new_G2202_ | new_G4852_ | new_G5154_;
  assign G5312 = new_G1488_ | new_G2191_ | new_G5181_ | new_G5182_;
  assign G5313 = new_G1496_ | new_G2199_ | new_G5183_ | new_G5184_;
  assign G5314 = ~new_G5191_;
  assign G5315 = ~new_G5192_;
  assign n2610_li = G1;
  assign n2613_li = n2610_lo;
  assign n2616_li = n2613_lo;
  assign n2619_li = n2616_lo;
  assign n2622_li = G2;
  assign n2625_li = n2622_lo;
  assign n2628_li = n2625_lo;
  assign n2631_li = n2628_lo;
  assign n2634_li = G3;
  assign n2637_li = n2634_lo;
  assign n2640_li = n2637_lo;
  assign n2643_li = n2640_lo;
  assign n2646_li = G4;
  assign n2649_li = n2646_lo;
  assign n2652_li = n2649_lo;
  assign n2655_li = n2652_lo;
  assign n2658_li = G5;
  assign n2661_li = n2658_lo;
  assign n2664_li = n2661_lo;
  assign n2667_li = n2664_lo;
  assign n2670_li = G6;
  assign n2673_li = n2670_lo;
  assign n2676_li = n2673_lo;
  assign n2679_li = n2676_lo;
  assign n2682_li = G7;
  assign n2685_li = n2682_lo;
  assign n2688_li = n2685_lo;
  assign n2691_li = n2688_lo;
  assign n2694_li = G8;
  assign n2697_li = n2694_lo;
  assign n2700_li = n2697_lo;
  assign n2703_li = n2700_lo;
  assign n2706_li = G9;
  assign n2709_li = n2706_lo;
  assign n2712_li = n2709_lo;
  assign n2715_li = n2712_lo;
  assign n2718_li = G10;
  assign n2721_li = n2718_lo;
  assign n2724_li = n2721_lo;
  assign n2727_li = n2724_lo;
  assign n2730_li = G11;
  assign n2733_li = n2730_lo;
  assign n2736_li = n2733_lo;
  assign n2739_li = n2736_lo;
  assign n2742_li = G12;
  assign n2745_li = n2742_lo;
  assign n2748_li = n2745_lo;
  assign n2751_li = n2748_lo;
  assign n2754_li = G13;
  assign n2757_li = n2754_lo;
  assign n2760_li = n2757_lo;
  assign n2763_li = n2760_lo;
  assign n2766_li = G14;
  assign n2769_li = n2766_lo;
  assign n2772_li = n2769_lo;
  assign n2775_li = n2772_lo;
  assign n2778_li = G15;
  assign n2781_li = n2778_lo;
  assign n2784_li = n2781_lo;
  assign n2787_li = n2784_lo;
  assign n2790_li = G16;
  assign n2793_li = n2790_lo;
  assign n2796_li = n2793_lo;
  assign n2799_li = n2796_lo;
  assign n2802_li = G17;
  assign n2805_li = n2802_lo;
  assign n2808_li = n2805_lo;
  assign n2811_li = n2808_lo;
  assign n2814_li = G18;
  assign n2817_li = n2814_lo;
  assign n2820_li = n2817_lo;
  assign n2823_li = n2820_lo;
  assign n2826_li = G19;
  assign n2829_li = n2826_lo;
  assign n2832_li = n2829_lo;
  assign n2835_li = n2832_lo;
  assign n2838_li = G20;
  assign n2841_li = n2838_lo;
  assign n2844_li = n2841_lo;
  assign n2847_li = n2844_lo;
  assign n2850_li = G21;
  assign n2853_li = n2850_lo;
  assign n2856_li = n2853_lo;
  assign n2859_li = n2856_lo;
  assign n2862_li = G22;
  assign n2865_li = n2862_lo;
  assign n2868_li = n2865_lo;
  assign n2871_li = n2868_lo;
  assign n2874_li = G23;
  assign n2877_li = n2874_lo;
  assign n2880_li = n2877_lo;
  assign n2883_li = n2880_lo;
  assign n2886_li = G24;
  assign n2889_li = n2886_lo;
  assign n2892_li = n2889_lo;
  assign n2895_li = n2892_lo;
  assign n2898_li = G25;
  assign n2901_li = n2898_lo;
  assign n2904_li = n2901_lo;
  assign n2907_li = n2904_lo;
  assign n2910_li = G26;
  assign n2913_li = n2910_lo;
  assign n2916_li = n2913_lo;
  assign n2919_li = n2916_lo;
  assign n2922_li = G27;
  assign n2925_li = n2922_lo;
  assign n2928_li = n2925_lo;
  assign n2931_li = n2928_lo;
  assign n2934_li = G28;
  assign n2937_li = n2934_lo;
  assign n2940_li = n2937_lo;
  assign n2943_li = n2940_lo;
  assign n2946_li = G29;
  assign n2949_li = n2946_lo;
  assign n2952_li = n2949_lo;
  assign n2955_li = n2952_lo;
  assign n2958_li = G30;
  assign n2961_li = n2958_lo;
  assign n2964_li = n2961_lo;
  assign n2967_li = n2964_lo;
  assign n2970_li = G31;
  assign n2973_li = n2970_lo;
  assign n2976_li = n2973_lo;
  assign n2979_li = n2976_lo;
  assign n2982_li = G32;
  assign n2985_li = n2982_lo;
  assign n2988_li = n2985_lo;
  assign n2991_li = n2988_lo;
  assign n2994_li = G33;
  assign n2997_li = n2994_lo;
  assign n3000_li = n2997_lo;
  assign n3003_li = n3000_lo;
  assign n3006_li = G34;
  assign n3009_li = n3006_lo;
  assign n3012_li = n3009_lo;
  assign n3015_li = n3012_lo;
  assign n3018_li = G35;
  assign n3021_li = n3018_lo;
  assign n3024_li = n3021_lo;
  assign n3027_li = n3024_lo;
  assign n3030_li = G36;
  assign n3033_li = n3030_lo;
  assign n3036_li = n3033_lo;
  assign n3039_li = n3036_lo;
  assign n3042_li = G37;
  assign n3045_li = n3042_lo;
  assign n3048_li = n3045_lo;
  assign n3051_li = n3048_lo;
  assign n3054_li = G38;
  assign n3057_li = n3054_lo;
  assign n3060_li = n3057_lo;
  assign n3063_li = n3060_lo;
  assign n3066_li = G39;
  assign n3069_li = n3066_lo;
  assign n3072_li = n3069_lo;
  assign n3075_li = n3072_lo;
  assign n3078_li = G40;
  assign n3081_li = n3078_lo;
  assign n3084_li = n3081_lo;
  assign n3087_li = n3084_lo;
  assign n3090_li = G41;
  assign n3093_li = n3090_lo;
  assign n3096_li = n3093_lo;
  assign n3099_li = n3096_lo;
  assign n3102_li = G42;
  assign n3105_li = n3102_lo;
  assign n3108_li = n3105_lo;
  assign n3111_li = n3108_lo;
  assign n3114_li = G43;
  assign n3117_li = n3114_lo;
  assign n3120_li = n3117_lo;
  assign n3123_li = n3120_lo;
  assign n3126_li = G44;
  assign n3129_li = n3126_lo;
  assign n3132_li = n3129_lo;
  assign n3135_li = n3132_lo;
  assign n3138_li = G45;
  assign n3141_li = n3138_lo;
  assign n3144_li = n3141_lo;
  assign n3147_li = n3144_lo;
  assign n3150_li = G46;
  assign n3153_li = n3150_lo;
  assign n3156_li = n3153_lo;
  assign n3159_li = n3156_lo;
  assign n3162_li = G47;
  assign n3165_li = n3162_lo;
  assign n3168_li = n3165_lo;
  assign n3171_li = n3168_lo;
  assign n3174_li = G48;
  assign n3177_li = n3174_lo;
  assign n3180_li = n3177_lo;
  assign n3183_li = n3180_lo;
  assign n3186_li = G49;
  assign n3189_li = n3186_lo;
  assign n3192_li = n3189_lo;
  assign n3195_li = n3192_lo;
  assign n3198_li = G50;
  assign n3201_li = n3198_lo;
  assign n3204_li = n3201_lo;
  assign n3207_li = n3204_lo;
  assign n3210_li = G51;
  assign n3213_li = n3210_lo;
  assign n3216_li = n3213_lo;
  assign n3219_li = n3216_lo;
  assign n3222_li = G52;
  assign n3225_li = n3222_lo;
  assign n3228_li = n3225_lo;
  assign n3231_li = n3228_lo;
  assign n3234_li = G53;
  assign n3237_li = n3234_lo;
  assign n3240_li = n3237_lo;
  assign n3243_li = n3240_lo;
  assign n3246_li = G54;
  assign n3249_li = n3246_lo;
  assign n3252_li = n3249_lo;
  assign n3255_li = n3252_lo;
  assign n3258_li = G55;
  assign n3261_li = n3258_lo;
  assign n3264_li = n3261_lo;
  assign n3267_li = n3264_lo;
  assign n3270_li = G56;
  assign n3273_li = n3270_lo;
  assign n3276_li = n3273_lo;
  assign n3279_li = n3276_lo;
  assign n3282_li = G57;
  assign n3285_li = n3282_lo;
  assign n3288_li = n3285_lo;
  assign n3291_li = n3288_lo;
  assign n3294_li = G58;
  assign n3297_li = n3294_lo;
  assign n3300_li = n3297_lo;
  assign n3303_li = n3300_lo;
  assign n3306_li = G59;
  assign n3309_li = n3306_lo;
  assign n3312_li = n3309_lo;
  assign n3315_li = n3312_lo;
  assign n3318_li = G60;
  assign n3321_li = n3318_lo;
  assign n3324_li = n3321_lo;
  assign n3327_li = n3324_lo;
  assign n3330_li = G61;
  assign n3333_li = n3330_lo;
  assign n3336_li = n3333_lo;
  assign n3339_li = n3336_lo;
  assign n3342_li = G62;
  assign n3345_li = n3342_lo;
  assign n3348_li = n3345_lo;
  assign n3351_li = n3348_lo;
  assign n3354_li = G63;
  assign n3357_li = n3354_lo;
  assign n3360_li = n3357_lo;
  assign n3363_li = n3360_lo;
  assign n3366_li = G64;
  assign n3369_li = n3366_lo;
  assign n3372_li = n3369_lo;
  assign n3375_li = n3372_lo;
  assign n3378_li = G65;
  assign n3381_li = n3378_lo;
  assign n3384_li = n3381_lo;
  assign n3387_li = n3384_lo;
  assign n3390_li = G66;
  assign n3393_li = n3390_lo;
  assign n3396_li = n3393_lo;
  assign n3399_li = n3396_lo;
  assign n3402_li = G67;
  assign n3405_li = n3402_lo;
  assign n3408_li = n3405_lo;
  assign n3411_li = n3408_lo;
  assign n3414_li = G68;
  assign n3417_li = n3414_lo;
  assign n3420_li = n3417_lo;
  assign n3423_li = n3420_lo;
  assign n3426_li = G69;
  assign n3429_li = n3426_lo;
  assign n3432_li = n3429_lo;
  assign n3435_li = n3432_lo;
  assign n3438_li = G70;
  assign n3441_li = n3438_lo;
  assign n3444_li = n3441_lo;
  assign n3447_li = n3444_lo;
  assign n3450_li = G71;
  assign n3453_li = n3450_lo;
  assign n3456_li = n3453_lo;
  assign n3459_li = n3456_lo;
  assign n3462_li = G72;
  assign n3465_li = n3462_lo;
  assign n3468_li = n3465_lo;
  assign n3471_li = n3468_lo;
  assign n3474_li = G73;
  assign n3477_li = n3474_lo;
  assign n3480_li = n3477_lo;
  assign n3483_li = n3480_lo;
  assign n3486_li = G74;
  assign n3489_li = n3486_lo;
  assign n3492_li = n3489_lo;
  assign n3495_li = n3492_lo;
  assign n3498_li = G75;
  assign n3501_li = n3498_lo;
  assign n3504_li = n3501_lo;
  assign n3507_li = n3504_lo;
  assign n3510_li = G76;
  assign n3513_li = n3510_lo;
  assign n3516_li = n3513_lo;
  assign n3519_li = n3516_lo;
  assign n3522_li = G77;
  assign n3525_li = n3522_lo;
  assign n3528_li = n3525_lo;
  assign n3531_li = n3528_lo;
  assign n3534_li = G78;
  assign n3537_li = n3534_lo;
  assign n3540_li = n3537_lo;
  assign n3543_li = n3540_lo;
  assign n3546_li = G79;
  assign n3549_li = n3546_lo;
  assign n3552_li = n3549_lo;
  assign n3555_li = n3552_lo;
  assign n3558_li = G80;
  assign n3561_li = n3558_lo;
  assign n3564_li = n3561_lo;
  assign n3567_li = n3564_lo;
  assign n3570_li = G81;
  assign n3573_li = n3570_lo;
  assign n3576_li = n3573_lo;
  assign n3579_li = n3576_lo;
  assign n3582_li = G82;
  assign n3585_li = n3582_lo;
  assign n3588_li = n3585_lo;
  assign n3591_li = n3588_lo;
  assign n3594_li = G83;
  assign n3597_li = n3594_lo;
  assign n3600_li = n3597_lo;
  assign n3603_li = n3600_lo;
  assign n3606_li = G84;
  assign n3609_li = n3606_lo;
  assign n3612_li = n3609_lo;
  assign n3615_li = n3612_lo;
  assign n3618_li = G85;
  assign n3621_li = n3618_lo;
  assign n3624_li = n3621_lo;
  assign n3627_li = n3624_lo;
  assign n3630_li = G86;
  assign n3633_li = n3630_lo;
  assign n3636_li = n3633_lo;
  assign n3639_li = n3636_lo;
  assign n3642_li = G87;
  assign n3645_li = n3642_lo;
  assign n3648_li = n3645_lo;
  assign n3651_li = n3648_lo;
  assign n3654_li = G88;
  assign n3657_li = n3654_lo;
  assign n3660_li = n3657_lo;
  assign n3663_li = n3660_lo;
  assign n3666_li = G89;
  assign n3669_li = n3666_lo;
  assign n3672_li = n3669_lo;
  assign n3675_li = n3672_lo;
  assign n3678_li = G90;
  assign n3681_li = n3678_lo;
  assign n3684_li = n3681_lo;
  assign n3687_li = n3684_lo;
  assign n3690_li = G91;
  assign n3693_li = n3690_lo;
  assign n3696_li = n3693_lo;
  assign n3699_li = n3696_lo;
  assign n3702_li = G92;
  assign n3705_li = n3702_lo;
  assign n3708_li = n3705_lo;
  assign n3711_li = n3708_lo;
  assign n3714_li = G93;
  assign n3717_li = n3714_lo;
  assign n3720_li = n3717_lo;
  assign n3723_li = n3720_lo;
  assign n3726_li = G94;
  assign n3729_li = n3726_lo;
  assign n3732_li = n3729_lo;
  assign n3735_li = n3732_lo;
  assign n3738_li = G95;
  assign n3741_li = n3738_lo;
  assign n3744_li = n3741_lo;
  assign n3747_li = n3744_lo;
  assign n3750_li = G96;
  assign n3753_li = n3750_lo;
  assign n3756_li = n3753_lo;
  assign n3759_li = n3756_lo;
  assign n3762_li = G97;
  assign n3765_li = n3762_lo;
  assign n3768_li = n3765_lo;
  assign n3771_li = n3768_lo;
  assign n3774_li = G98;
  assign n3777_li = n3774_lo;
  assign n3780_li = n3777_lo;
  assign n3783_li = n3780_lo;
  assign n3786_li = G99;
  assign n3789_li = n3786_lo;
  assign n3792_li = n3789_lo;
  assign n3795_li = n3792_lo;
  assign n3798_li = G100;
  assign n3801_li = n3798_lo;
  assign n3804_li = n3801_lo;
  assign n3807_li = n3804_lo;
  assign n3810_li = G101;
  assign n3813_li = n3810_lo;
  assign n3816_li = n3813_lo;
  assign n3819_li = n3816_lo;
  assign n3822_li = G102;
  assign n3825_li = n3822_lo;
  assign n3828_li = n3825_lo;
  assign n3831_li = n3828_lo;
  assign n3834_li = G103;
  assign n3837_li = n3834_lo;
  assign n3840_li = n3837_lo;
  assign n3843_li = n3840_lo;
  assign n3846_li = G104;
  assign n3849_li = n3846_lo;
  assign n3852_li = n3849_lo;
  assign n3855_li = n3852_lo;
  assign n3858_li = G105;
  assign n3861_li = n3858_lo;
  assign n3864_li = n3861_lo;
  assign n3867_li = n3864_lo;
  assign n3870_li = G106;
  assign n3873_li = n3870_lo;
  assign n3876_li = n3873_lo;
  assign n3879_li = n3876_lo;
  assign n3882_li = G107;
  assign n3885_li = n3882_lo;
  assign n3888_li = n3885_lo;
  assign n3891_li = n3888_lo;
  assign n3894_li = G108;
  assign n3897_li = n3894_lo;
  assign n3900_li = n3897_lo;
  assign n3903_li = n3900_lo;
  assign n3906_li = G109;
  assign n3909_li = n3906_lo;
  assign n3912_li = n3909_lo;
  assign n3915_li = n3912_lo;
  assign n3918_li = G110;
  assign n3921_li = n3918_lo;
  assign n3924_li = n3921_lo;
  assign n3927_li = n3924_lo;
  assign n3930_li = G111;
  assign n3933_li = n3930_lo;
  assign n3936_li = n3933_lo;
  assign n3939_li = n3936_lo;
  assign n3942_li = G112;
  assign n3945_li = n3942_lo;
  assign n3948_li = n3945_lo;
  assign n3951_li = n3948_lo;
  assign n3954_li = G113;
  assign n3957_li = n3954_lo;
  assign n3960_li = n3957_lo;
  assign n3963_li = n3960_lo;
  assign n3966_li = G114;
  assign n3969_li = n3966_lo;
  assign n3972_li = n3969_lo;
  assign n3975_li = n3972_lo;
  assign n3978_li = G115;
  assign n3981_li = n3978_lo;
  assign n3984_li = n3981_lo;
  assign n3987_li = n3984_lo;
  assign n3990_li = G116;
  assign n3993_li = n3990_lo;
  assign n3996_li = n3993_lo;
  assign n3999_li = n3996_lo;
  assign n4002_li = G117;
  assign n4005_li = n4002_lo;
  assign n4008_li = n4005_lo;
  assign n4011_li = n4008_lo;
  assign n4014_li = G118;
  assign n4017_li = n4014_lo;
  assign n4020_li = n4017_lo;
  assign n4023_li = n4020_lo;
  assign n4026_li = G119;
  assign n4029_li = n4026_lo;
  assign n4032_li = n4029_lo;
  assign n4035_li = n4032_lo;
  assign n4038_li = G120;
  assign n4041_li = n4038_lo;
  assign n4044_li = n4041_lo;
  assign n4047_li = n4044_lo;
  assign n4050_li = G121;
  assign n4053_li = n4050_lo;
  assign n4056_li = n4053_lo;
  assign n4059_li = n4056_lo;
  assign n4062_li = G122;
  assign n4065_li = n4062_lo;
  assign n4068_li = n4065_lo;
  assign n4071_li = n4068_lo;
  assign n4074_li = G123;
  assign n4077_li = n4074_lo;
  assign n4080_li = n4077_lo;
  assign n4083_li = n4080_lo;
  assign n4086_li = G124;
  assign n4089_li = n4086_lo;
  assign n4092_li = n4089_lo;
  assign n4095_li = n4092_lo;
  assign n4098_li = G125;
  assign n4101_li = n4098_lo;
  assign n4104_li = n4101_lo;
  assign n4107_li = n4104_lo;
  assign n4110_li = G126;
  assign n4113_li = n4110_lo;
  assign n4116_li = n4113_lo;
  assign n4119_li = n4116_lo;
  assign n4122_li = G127;
  assign n4125_li = n4122_lo;
  assign n4128_li = n4125_lo;
  assign n4131_li = n4128_lo;
  assign n4134_li = G128;
  assign n4137_li = n4134_lo;
  assign n4140_li = n4137_lo;
  assign n4143_li = n4140_lo;
  assign n4146_li = G129;
  assign n4149_li = n4146_lo;
  assign n4152_li = n4149_lo;
  assign n4155_li = n4152_lo;
  assign n4158_li = G130;
  assign n4161_li = n4158_lo;
  assign n4164_li = n4161_lo;
  assign n4167_li = n4164_lo;
  assign n4170_li = G131;
  assign n4173_li = n4170_lo;
  assign n4176_li = n4173_lo;
  assign n4179_li = n4176_lo;
  assign n4182_li = G132;
  assign n4185_li = n4182_lo;
  assign n4188_li = n4185_lo;
  assign n4191_li = n4188_lo;
  assign n4194_li = G133;
  assign n4197_li = n4194_lo;
  assign n4200_li = n4197_lo;
  assign n4203_li = n4200_lo;
  assign n4206_li = G134;
  assign n4209_li = n4206_lo;
  assign n4212_li = n4209_lo;
  assign n4215_li = n4212_lo;
  assign n4218_li = G135;
  assign n4221_li = n4218_lo;
  assign n4224_li = n4221_lo;
  assign n4227_li = n4224_lo;
  assign n4230_li = G136;
  assign n4233_li = n4230_lo;
  assign n4236_li = n4233_lo;
  assign n4239_li = n4236_lo;
  assign n4242_li = G137;
  assign n4245_li = n4242_lo;
  assign n4248_li = n4245_lo;
  assign n4251_li = n4248_lo;
  assign n4254_li = G138;
  assign n4257_li = n4254_lo;
  assign n4260_li = n4257_lo;
  assign n4263_li = n4260_lo;
  assign n4266_li = G139;
  assign n4269_li = n4266_lo;
  assign n4272_li = n4269_lo;
  assign n4275_li = n4272_lo;
  assign n4278_li = G140;
  assign n4281_li = n4278_lo;
  assign n4284_li = n4281_lo;
  assign n4287_li = n4284_lo;
  assign n4290_li = G141;
  assign n4293_li = n4290_lo;
  assign n4296_li = n4293_lo;
  assign n4299_li = n4296_lo;
  assign n4302_li = G142;
  assign n4305_li = n4302_lo;
  assign n4308_li = n4305_lo;
  assign n4311_li = n4308_lo;
  assign n4314_li = G143;
  assign n4317_li = n4314_lo;
  assign n4320_li = n4317_lo;
  assign n4323_li = n4320_lo;
  assign n4326_li = G144;
  assign n4329_li = n4326_lo;
  assign n4332_li = n4329_lo;
  assign n4335_li = n4332_lo;
  assign n4338_li = G145;
  assign n4341_li = n4338_lo;
  assign n4344_li = n4341_lo;
  assign n4347_li = n4344_lo;
  assign n4350_li = G146;
  assign n4353_li = n4350_lo;
  assign n4356_li = n4353_lo;
  assign n4359_li = n4356_lo;
  assign n4362_li = G147;
  assign n4365_li = n4362_lo;
  assign n4368_li = n4365_lo;
  assign n4371_li = n4368_lo;
  assign n4374_li = G148;
  assign n4377_li = n4374_lo;
  assign n4380_li = n4377_lo;
  assign n4383_li = n4380_lo;
  assign n4386_li = G149;
  assign n4389_li = n4386_lo;
  assign n4392_li = n4389_lo;
  assign n4395_li = n4392_lo;
  assign n4398_li = G150;
  assign n4401_li = n4398_lo;
  assign n4404_li = n4401_lo;
  assign n4407_li = n4404_lo;
  assign n4410_li = G151;
  assign n4413_li = n4410_lo;
  assign n4416_li = n4413_lo;
  assign n4419_li = n4416_lo;
  assign n4422_li = G152;
  assign n4425_li = n4422_lo;
  assign n4428_li = n4425_lo;
  assign n4431_li = n4428_lo;
  assign n4434_li = G153;
  assign n4437_li = n4434_lo;
  assign n4440_li = n4437_lo;
  assign n4443_li = n4440_lo;
  assign n4446_li = G154;
  assign n4449_li = n4446_lo;
  assign n4452_li = n4449_lo;
  assign n4455_li = n4452_lo;
  assign n4458_li = G155;
  assign n4461_li = n4458_lo;
  assign n4464_li = n4461_lo;
  assign n4467_li = n4464_lo;
  assign n4470_li = G156;
  assign n4473_li = n4470_lo;
  assign n4476_li = n4473_lo;
  assign n4479_li = n4476_lo;
  assign n4482_li = G157;
  assign n4485_li = n4482_lo;
  assign n4488_li = n4485_lo;
  assign n4491_li = n4488_lo;
  assign n4494_li = G158;
  assign n4497_li = n4494_lo;
  assign n4500_li = n4497_lo;
  assign n4503_li = n4500_lo;
  assign n4506_li = G159;
  assign n4509_li = n4506_lo;
  assign n4512_li = n4509_lo;
  assign n4515_li = n4512_lo;
  assign n4518_li = G160;
  assign n4521_li = n4518_lo;
  assign n4524_li = n4521_lo;
  assign n4527_li = n4524_lo;
  assign n4530_li = G161;
  assign n4533_li = n4530_lo;
  assign n4536_li = n4533_lo;
  assign n4539_li = n4536_lo;
  assign n4542_li = G162;
  assign n4545_li = n4542_lo;
  assign n4548_li = n4545_lo;
  assign n4551_li = n4548_lo;
  assign n4554_li = G163;
  assign n4557_li = n4554_lo;
  assign n4560_li = n4557_lo;
  assign n4563_li = n4560_lo;
  assign n4566_li = G164;
  assign n4569_li = n4566_lo;
  assign n4572_li = n4569_lo;
  assign n4575_li = n4572_lo;
  assign n4578_li = G165;
  assign n4581_li = n4578_lo;
  assign n4584_li = n4581_lo;
  assign n4587_li = n4584_lo;
  assign n4590_li = G166;
  assign n4593_li = n4590_lo;
  assign n4596_li = n4593_lo;
  assign n4599_li = n4596_lo;
  assign n4602_li = G167;
  assign n4605_li = n4602_lo;
  assign n4608_li = n4605_lo;
  assign n4611_li = n4608_lo;
  assign n4614_li = G168;
  assign n4617_li = n4614_lo;
  assign n4620_li = n4617_lo;
  assign n4623_li = n4620_lo;
  assign n4626_li = G169;
  assign n4629_li = n4626_lo;
  assign n4632_li = n4629_lo;
  assign n4635_li = n4632_lo;
  assign n4638_li = G170;
  assign n4641_li = n4638_lo;
  assign n4644_li = n4641_lo;
  assign n4647_li = n4644_lo;
  assign n4650_li = G171;
  assign n4653_li = n4650_lo;
  assign n4656_li = n4653_lo;
  assign n4659_li = n4656_lo;
  assign n4662_li = G172;
  assign n4665_li = n4662_lo;
  assign n4668_li = n4665_lo;
  assign n4671_li = n4668_lo;
  assign n4674_li = G173;
  assign n4677_li = n4674_lo;
  assign n4680_li = n4677_lo;
  assign n4683_li = n4680_lo;
  assign n4686_li = G174;
  assign n4689_li = n4686_lo;
  assign n4692_li = n4689_lo;
  assign n4695_li = n4692_lo;
  assign n4698_li = G175;
  assign n4701_li = n4698_lo;
  assign n4704_li = n4701_lo;
  assign n4707_li = n4704_lo;
  assign n4710_li = G176;
  assign n4713_li = n4710_lo;
  assign n4716_li = n4713_lo;
  assign n4719_li = n4716_lo;
  assign n4722_li = G177;
  assign n4725_li = n4722_lo;
  assign n4728_li = n4725_lo;
  assign n4731_li = n4728_lo;
  assign n4734_li = G178;
  assign n4737_li = n4734_lo;
  assign n4740_li = n4737_lo;
  assign n4743_li = n4740_lo;
  always @ (posedge clk) begin
    n2610_lo <= n2610_li;
    n2613_lo <= n2613_li;
    n2616_lo <= n2616_li;
    n2619_lo <= n2619_li;
    n2622_lo <= n2622_li;
    n2625_lo <= n2625_li;
    n2628_lo <= n2628_li;
    n2631_lo <= n2631_li;
    n2634_lo <= n2634_li;
    n2637_lo <= n2637_li;
    n2640_lo <= n2640_li;
    n2643_lo <= n2643_li;
    n2646_lo <= n2646_li;
    n2649_lo <= n2649_li;
    n2652_lo <= n2652_li;
    n2655_lo <= n2655_li;
    n2658_lo <= n2658_li;
    n2661_lo <= n2661_li;
    n2664_lo <= n2664_li;
    n2667_lo <= n2667_li;
    n2670_lo <= n2670_li;
    n2673_lo <= n2673_li;
    n2676_lo <= n2676_li;
    n2679_lo <= n2679_li;
    n2682_lo <= n2682_li;
    n2685_lo <= n2685_li;
    n2688_lo <= n2688_li;
    n2691_lo <= n2691_li;
    n2694_lo <= n2694_li;
    n2697_lo <= n2697_li;
    n2700_lo <= n2700_li;
    n2703_lo <= n2703_li;
    n2706_lo <= n2706_li;
    n2709_lo <= n2709_li;
    n2712_lo <= n2712_li;
    n2715_lo <= n2715_li;
    n2718_lo <= n2718_li;
    n2721_lo <= n2721_li;
    n2724_lo <= n2724_li;
    n2727_lo <= n2727_li;
    n2730_lo <= n2730_li;
    n2733_lo <= n2733_li;
    n2736_lo <= n2736_li;
    n2739_lo <= n2739_li;
    n2742_lo <= n2742_li;
    n2745_lo <= n2745_li;
    n2748_lo <= n2748_li;
    n2751_lo <= n2751_li;
    n2754_lo <= n2754_li;
    n2757_lo <= n2757_li;
    n2760_lo <= n2760_li;
    n2763_lo <= n2763_li;
    n2766_lo <= n2766_li;
    n2769_lo <= n2769_li;
    n2772_lo <= n2772_li;
    n2775_lo <= n2775_li;
    n2778_lo <= n2778_li;
    n2781_lo <= n2781_li;
    n2784_lo <= n2784_li;
    n2787_lo <= n2787_li;
    n2790_lo <= n2790_li;
    n2793_lo <= n2793_li;
    n2796_lo <= n2796_li;
    n2799_lo <= n2799_li;
    n2802_lo <= n2802_li;
    n2805_lo <= n2805_li;
    n2808_lo <= n2808_li;
    n2811_lo <= n2811_li;
    n2814_lo <= n2814_li;
    n2817_lo <= n2817_li;
    n2820_lo <= n2820_li;
    n2823_lo <= n2823_li;
    n2826_lo <= n2826_li;
    n2829_lo <= n2829_li;
    n2832_lo <= n2832_li;
    n2835_lo <= n2835_li;
    n2838_lo <= n2838_li;
    n2841_lo <= n2841_li;
    n2844_lo <= n2844_li;
    n2847_lo <= n2847_li;
    n2850_lo <= n2850_li;
    n2853_lo <= n2853_li;
    n2856_lo <= n2856_li;
    n2859_lo <= n2859_li;
    n2862_lo <= n2862_li;
    n2865_lo <= n2865_li;
    n2868_lo <= n2868_li;
    n2871_lo <= n2871_li;
    n2874_lo <= n2874_li;
    n2877_lo <= n2877_li;
    n2880_lo <= n2880_li;
    n2883_lo <= n2883_li;
    n2886_lo <= n2886_li;
    n2889_lo <= n2889_li;
    n2892_lo <= n2892_li;
    n2895_lo <= n2895_li;
    n2898_lo <= n2898_li;
    n2901_lo <= n2901_li;
    n2904_lo <= n2904_li;
    n2907_lo <= n2907_li;
    n2910_lo <= n2910_li;
    n2913_lo <= n2913_li;
    n2916_lo <= n2916_li;
    n2919_lo <= n2919_li;
    n2922_lo <= n2922_li;
    n2925_lo <= n2925_li;
    n2928_lo <= n2928_li;
    n2931_lo <= n2931_li;
    n2934_lo <= n2934_li;
    n2937_lo <= n2937_li;
    n2940_lo <= n2940_li;
    n2943_lo <= n2943_li;
    n2946_lo <= n2946_li;
    n2949_lo <= n2949_li;
    n2952_lo <= n2952_li;
    n2955_lo <= n2955_li;
    n2958_lo <= n2958_li;
    n2961_lo <= n2961_li;
    n2964_lo <= n2964_li;
    n2967_lo <= n2967_li;
    n2970_lo <= n2970_li;
    n2973_lo <= n2973_li;
    n2976_lo <= n2976_li;
    n2979_lo <= n2979_li;
    n2982_lo <= n2982_li;
    n2985_lo <= n2985_li;
    n2988_lo <= n2988_li;
    n2991_lo <= n2991_li;
    n2994_lo <= n2994_li;
    n2997_lo <= n2997_li;
    n3000_lo <= n3000_li;
    n3003_lo <= n3003_li;
    n3006_lo <= n3006_li;
    n3009_lo <= n3009_li;
    n3012_lo <= n3012_li;
    n3015_lo <= n3015_li;
    n3018_lo <= n3018_li;
    n3021_lo <= n3021_li;
    n3024_lo <= n3024_li;
    n3027_lo <= n3027_li;
    n3030_lo <= n3030_li;
    n3033_lo <= n3033_li;
    n3036_lo <= n3036_li;
    n3039_lo <= n3039_li;
    n3042_lo <= n3042_li;
    n3045_lo <= n3045_li;
    n3048_lo <= n3048_li;
    n3051_lo <= n3051_li;
    n3054_lo <= n3054_li;
    n3057_lo <= n3057_li;
    n3060_lo <= n3060_li;
    n3063_lo <= n3063_li;
    n3066_lo <= n3066_li;
    n3069_lo <= n3069_li;
    n3072_lo <= n3072_li;
    n3075_lo <= n3075_li;
    n3078_lo <= n3078_li;
    n3081_lo <= n3081_li;
    n3084_lo <= n3084_li;
    n3087_lo <= n3087_li;
    n3090_lo <= n3090_li;
    n3093_lo <= n3093_li;
    n3096_lo <= n3096_li;
    n3099_lo <= n3099_li;
    n3102_lo <= n3102_li;
    n3105_lo <= n3105_li;
    n3108_lo <= n3108_li;
    n3111_lo <= n3111_li;
    n3114_lo <= n3114_li;
    n3117_lo <= n3117_li;
    n3120_lo <= n3120_li;
    n3123_lo <= n3123_li;
    n3126_lo <= n3126_li;
    n3129_lo <= n3129_li;
    n3132_lo <= n3132_li;
    n3135_lo <= n3135_li;
    n3138_lo <= n3138_li;
    n3141_lo <= n3141_li;
    n3144_lo <= n3144_li;
    n3147_lo <= n3147_li;
    n3150_lo <= n3150_li;
    n3153_lo <= n3153_li;
    n3156_lo <= n3156_li;
    n3159_lo <= n3159_li;
    n3162_lo <= n3162_li;
    n3165_lo <= n3165_li;
    n3168_lo <= n3168_li;
    n3171_lo <= n3171_li;
    n3174_lo <= n3174_li;
    n3177_lo <= n3177_li;
    n3180_lo <= n3180_li;
    n3183_lo <= n3183_li;
    n3186_lo <= n3186_li;
    n3189_lo <= n3189_li;
    n3192_lo <= n3192_li;
    n3195_lo <= n3195_li;
    n3198_lo <= n3198_li;
    n3201_lo <= n3201_li;
    n3204_lo <= n3204_li;
    n3207_lo <= n3207_li;
    n3210_lo <= n3210_li;
    n3213_lo <= n3213_li;
    n3216_lo <= n3216_li;
    n3219_lo <= n3219_li;
    n3222_lo <= n3222_li;
    n3225_lo <= n3225_li;
    n3228_lo <= n3228_li;
    n3231_lo <= n3231_li;
    n3234_lo <= n3234_li;
    n3237_lo <= n3237_li;
    n3240_lo <= n3240_li;
    n3243_lo <= n3243_li;
    n3246_lo <= n3246_li;
    n3249_lo <= n3249_li;
    n3252_lo <= n3252_li;
    n3255_lo <= n3255_li;
    n3258_lo <= n3258_li;
    n3261_lo <= n3261_li;
    n3264_lo <= n3264_li;
    n3267_lo <= n3267_li;
    n3270_lo <= n3270_li;
    n3273_lo <= n3273_li;
    n3276_lo <= n3276_li;
    n3279_lo <= n3279_li;
    n3282_lo <= n3282_li;
    n3285_lo <= n3285_li;
    n3288_lo <= n3288_li;
    n3291_lo <= n3291_li;
    n3294_lo <= n3294_li;
    n3297_lo <= n3297_li;
    n3300_lo <= n3300_li;
    n3303_lo <= n3303_li;
    n3306_lo <= n3306_li;
    n3309_lo <= n3309_li;
    n3312_lo <= n3312_li;
    n3315_lo <= n3315_li;
    n3318_lo <= n3318_li;
    n3321_lo <= n3321_li;
    n3324_lo <= n3324_li;
    n3327_lo <= n3327_li;
    n3330_lo <= n3330_li;
    n3333_lo <= n3333_li;
    n3336_lo <= n3336_li;
    n3339_lo <= n3339_li;
    n3342_lo <= n3342_li;
    n3345_lo <= n3345_li;
    n3348_lo <= n3348_li;
    n3351_lo <= n3351_li;
    n3354_lo <= n3354_li;
    n3357_lo <= n3357_li;
    n3360_lo <= n3360_li;
    n3363_lo <= n3363_li;
    n3366_lo <= n3366_li;
    n3369_lo <= n3369_li;
    n3372_lo <= n3372_li;
    n3375_lo <= n3375_li;
    n3378_lo <= n3378_li;
    n3381_lo <= n3381_li;
    n3384_lo <= n3384_li;
    n3387_lo <= n3387_li;
    n3390_lo <= n3390_li;
    n3393_lo <= n3393_li;
    n3396_lo <= n3396_li;
    n3399_lo <= n3399_li;
    n3402_lo <= n3402_li;
    n3405_lo <= n3405_li;
    n3408_lo <= n3408_li;
    n3411_lo <= n3411_li;
    n3414_lo <= n3414_li;
    n3417_lo <= n3417_li;
    n3420_lo <= n3420_li;
    n3423_lo <= n3423_li;
    n3426_lo <= n3426_li;
    n3429_lo <= n3429_li;
    n3432_lo <= n3432_li;
    n3435_lo <= n3435_li;
    n3438_lo <= n3438_li;
    n3441_lo <= n3441_li;
    n3444_lo <= n3444_li;
    n3447_lo <= n3447_li;
    n3450_lo <= n3450_li;
    n3453_lo <= n3453_li;
    n3456_lo <= n3456_li;
    n3459_lo <= n3459_li;
    n3462_lo <= n3462_li;
    n3465_lo <= n3465_li;
    n3468_lo <= n3468_li;
    n3471_lo <= n3471_li;
    n3474_lo <= n3474_li;
    n3477_lo <= n3477_li;
    n3480_lo <= n3480_li;
    n3483_lo <= n3483_li;
    n3486_lo <= n3486_li;
    n3489_lo <= n3489_li;
    n3492_lo <= n3492_li;
    n3495_lo <= n3495_li;
    n3498_lo <= n3498_li;
    n3501_lo <= n3501_li;
    n3504_lo <= n3504_li;
    n3507_lo <= n3507_li;
    n3510_lo <= n3510_li;
    n3513_lo <= n3513_li;
    n3516_lo <= n3516_li;
    n3519_lo <= n3519_li;
    n3522_lo <= n3522_li;
    n3525_lo <= n3525_li;
    n3528_lo <= n3528_li;
    n3531_lo <= n3531_li;
    n3534_lo <= n3534_li;
    n3537_lo <= n3537_li;
    n3540_lo <= n3540_li;
    n3543_lo <= n3543_li;
    n3546_lo <= n3546_li;
    n3549_lo <= n3549_li;
    n3552_lo <= n3552_li;
    n3555_lo <= n3555_li;
    n3558_lo <= n3558_li;
    n3561_lo <= n3561_li;
    n3564_lo <= n3564_li;
    n3567_lo <= n3567_li;
    n3570_lo <= n3570_li;
    n3573_lo <= n3573_li;
    n3576_lo <= n3576_li;
    n3579_lo <= n3579_li;
    n3582_lo <= n3582_li;
    n3585_lo <= n3585_li;
    n3588_lo <= n3588_li;
    n3591_lo <= n3591_li;
    n3594_lo <= n3594_li;
    n3597_lo <= n3597_li;
    n3600_lo <= n3600_li;
    n3603_lo <= n3603_li;
    n3606_lo <= n3606_li;
    n3609_lo <= n3609_li;
    n3612_lo <= n3612_li;
    n3615_lo <= n3615_li;
    n3618_lo <= n3618_li;
    n3621_lo <= n3621_li;
    n3624_lo <= n3624_li;
    n3627_lo <= n3627_li;
    n3630_lo <= n3630_li;
    n3633_lo <= n3633_li;
    n3636_lo <= n3636_li;
    n3639_lo <= n3639_li;
    n3642_lo <= n3642_li;
    n3645_lo <= n3645_li;
    n3648_lo <= n3648_li;
    n3651_lo <= n3651_li;
    n3654_lo <= n3654_li;
    n3657_lo <= n3657_li;
    n3660_lo <= n3660_li;
    n3663_lo <= n3663_li;
    n3666_lo <= n3666_li;
    n3669_lo <= n3669_li;
    n3672_lo <= n3672_li;
    n3675_lo <= n3675_li;
    n3678_lo <= n3678_li;
    n3681_lo <= n3681_li;
    n3684_lo <= n3684_li;
    n3687_lo <= n3687_li;
    n3690_lo <= n3690_li;
    n3693_lo <= n3693_li;
    n3696_lo <= n3696_li;
    n3699_lo <= n3699_li;
    n3702_lo <= n3702_li;
    n3705_lo <= n3705_li;
    n3708_lo <= n3708_li;
    n3711_lo <= n3711_li;
    n3714_lo <= n3714_li;
    n3717_lo <= n3717_li;
    n3720_lo <= n3720_li;
    n3723_lo <= n3723_li;
    n3726_lo <= n3726_li;
    n3729_lo <= n3729_li;
    n3732_lo <= n3732_li;
    n3735_lo <= n3735_li;
    n3738_lo <= n3738_li;
    n3741_lo <= n3741_li;
    n3744_lo <= n3744_li;
    n3747_lo <= n3747_li;
    n3750_lo <= n3750_li;
    n3753_lo <= n3753_li;
    n3756_lo <= n3756_li;
    n3759_lo <= n3759_li;
    n3762_lo <= n3762_li;
    n3765_lo <= n3765_li;
    n3768_lo <= n3768_li;
    n3771_lo <= n3771_li;
    n3774_lo <= n3774_li;
    n3777_lo <= n3777_li;
    n3780_lo <= n3780_li;
    n3783_lo <= n3783_li;
    n3786_lo <= n3786_li;
    n3789_lo <= n3789_li;
    n3792_lo <= n3792_li;
    n3795_lo <= n3795_li;
    n3798_lo <= n3798_li;
    n3801_lo <= n3801_li;
    n3804_lo <= n3804_li;
    n3807_lo <= n3807_li;
    n3810_lo <= n3810_li;
    n3813_lo <= n3813_li;
    n3816_lo <= n3816_li;
    n3819_lo <= n3819_li;
    n3822_lo <= n3822_li;
    n3825_lo <= n3825_li;
    n3828_lo <= n3828_li;
    n3831_lo <= n3831_li;
    n3834_lo <= n3834_li;
    n3837_lo <= n3837_li;
    n3840_lo <= n3840_li;
    n3843_lo <= n3843_li;
    n3846_lo <= n3846_li;
    n3849_lo <= n3849_li;
    n3852_lo <= n3852_li;
    n3855_lo <= n3855_li;
    n3858_lo <= n3858_li;
    n3861_lo <= n3861_li;
    n3864_lo <= n3864_li;
    n3867_lo <= n3867_li;
    n3870_lo <= n3870_li;
    n3873_lo <= n3873_li;
    n3876_lo <= n3876_li;
    n3879_lo <= n3879_li;
    n3882_lo <= n3882_li;
    n3885_lo <= n3885_li;
    n3888_lo <= n3888_li;
    n3891_lo <= n3891_li;
    n3894_lo <= n3894_li;
    n3897_lo <= n3897_li;
    n3900_lo <= n3900_li;
    n3903_lo <= n3903_li;
    n3906_lo <= n3906_li;
    n3909_lo <= n3909_li;
    n3912_lo <= n3912_li;
    n3915_lo <= n3915_li;
    n3918_lo <= n3918_li;
    n3921_lo <= n3921_li;
    n3924_lo <= n3924_li;
    n3927_lo <= n3927_li;
    n3930_lo <= n3930_li;
    n3933_lo <= n3933_li;
    n3936_lo <= n3936_li;
    n3939_lo <= n3939_li;
    n3942_lo <= n3942_li;
    n3945_lo <= n3945_li;
    n3948_lo <= n3948_li;
    n3951_lo <= n3951_li;
    n3954_lo <= n3954_li;
    n3957_lo <= n3957_li;
    n3960_lo <= n3960_li;
    n3963_lo <= n3963_li;
    n3966_lo <= n3966_li;
    n3969_lo <= n3969_li;
    n3972_lo <= n3972_li;
    n3975_lo <= n3975_li;
    n3978_lo <= n3978_li;
    n3981_lo <= n3981_li;
    n3984_lo <= n3984_li;
    n3987_lo <= n3987_li;
    n3990_lo <= n3990_li;
    n3993_lo <= n3993_li;
    n3996_lo <= n3996_li;
    n3999_lo <= n3999_li;
    n4002_lo <= n4002_li;
    n4005_lo <= n4005_li;
    n4008_lo <= n4008_li;
    n4011_lo <= n4011_li;
    n4014_lo <= n4014_li;
    n4017_lo <= n4017_li;
    n4020_lo <= n4020_li;
    n4023_lo <= n4023_li;
    n4026_lo <= n4026_li;
    n4029_lo <= n4029_li;
    n4032_lo <= n4032_li;
    n4035_lo <= n4035_li;
    n4038_lo <= n4038_li;
    n4041_lo <= n4041_li;
    n4044_lo <= n4044_li;
    n4047_lo <= n4047_li;
    n4050_lo <= n4050_li;
    n4053_lo <= n4053_li;
    n4056_lo <= n4056_li;
    n4059_lo <= n4059_li;
    n4062_lo <= n4062_li;
    n4065_lo <= n4065_li;
    n4068_lo <= n4068_li;
    n4071_lo <= n4071_li;
    n4074_lo <= n4074_li;
    n4077_lo <= n4077_li;
    n4080_lo <= n4080_li;
    n4083_lo <= n4083_li;
    n4086_lo <= n4086_li;
    n4089_lo <= n4089_li;
    n4092_lo <= n4092_li;
    n4095_lo <= n4095_li;
    n4098_lo <= n4098_li;
    n4101_lo <= n4101_li;
    n4104_lo <= n4104_li;
    n4107_lo <= n4107_li;
    n4110_lo <= n4110_li;
    n4113_lo <= n4113_li;
    n4116_lo <= n4116_li;
    n4119_lo <= n4119_li;
    n4122_lo <= n4122_li;
    n4125_lo <= n4125_li;
    n4128_lo <= n4128_li;
    n4131_lo <= n4131_li;
    n4134_lo <= n4134_li;
    n4137_lo <= n4137_li;
    n4140_lo <= n4140_li;
    n4143_lo <= n4143_li;
    n4146_lo <= n4146_li;
    n4149_lo <= n4149_li;
    n4152_lo <= n4152_li;
    n4155_lo <= n4155_li;
    n4158_lo <= n4158_li;
    n4161_lo <= n4161_li;
    n4164_lo <= n4164_li;
    n4167_lo <= n4167_li;
    n4170_lo <= n4170_li;
    n4173_lo <= n4173_li;
    n4176_lo <= n4176_li;
    n4179_lo <= n4179_li;
    n4182_lo <= n4182_li;
    n4185_lo <= n4185_li;
    n4188_lo <= n4188_li;
    n4191_lo <= n4191_li;
    n4194_lo <= n4194_li;
    n4197_lo <= n4197_li;
    n4200_lo <= n4200_li;
    n4203_lo <= n4203_li;
    n4206_lo <= n4206_li;
    n4209_lo <= n4209_li;
    n4212_lo <= n4212_li;
    n4215_lo <= n4215_li;
    n4218_lo <= n4218_li;
    n4221_lo <= n4221_li;
    n4224_lo <= n4224_li;
    n4227_lo <= n4227_li;
    n4230_lo <= n4230_li;
    n4233_lo <= n4233_li;
    n4236_lo <= n4236_li;
    n4239_lo <= n4239_li;
    n4242_lo <= n4242_li;
    n4245_lo <= n4245_li;
    n4248_lo <= n4248_li;
    n4251_lo <= n4251_li;
    n4254_lo <= n4254_li;
    n4257_lo <= n4257_li;
    n4260_lo <= n4260_li;
    n4263_lo <= n4263_li;
    n4266_lo <= n4266_li;
    n4269_lo <= n4269_li;
    n4272_lo <= n4272_li;
    n4275_lo <= n4275_li;
    n4278_lo <= n4278_li;
    n4281_lo <= n4281_li;
    n4284_lo <= n4284_li;
    n4287_lo <= n4287_li;
    n4290_lo <= n4290_li;
    n4293_lo <= n4293_li;
    n4296_lo <= n4296_li;
    n4299_lo <= n4299_li;
    n4302_lo <= n4302_li;
    n4305_lo <= n4305_li;
    n4308_lo <= n4308_li;
    n4311_lo <= n4311_li;
    n4314_lo <= n4314_li;
    n4317_lo <= n4317_li;
    n4320_lo <= n4320_li;
    n4323_lo <= n4323_li;
    n4326_lo <= n4326_li;
    n4329_lo <= n4329_li;
    n4332_lo <= n4332_li;
    n4335_lo <= n4335_li;
    n4338_lo <= n4338_li;
    n4341_lo <= n4341_li;
    n4344_lo <= n4344_li;
    n4347_lo <= n4347_li;
    n4350_lo <= n4350_li;
    n4353_lo <= n4353_li;
    n4356_lo <= n4356_li;
    n4359_lo <= n4359_li;
    n4362_lo <= n4362_li;
    n4365_lo <= n4365_li;
    n4368_lo <= n4368_li;
    n4371_lo <= n4371_li;
    n4374_lo <= n4374_li;
    n4377_lo <= n4377_li;
    n4380_lo <= n4380_li;
    n4383_lo <= n4383_li;
    n4386_lo <= n4386_li;
    n4389_lo <= n4389_li;
    n4392_lo <= n4392_li;
    n4395_lo <= n4395_li;
    n4398_lo <= n4398_li;
    n4401_lo <= n4401_li;
    n4404_lo <= n4404_li;
    n4407_lo <= n4407_li;
    n4410_lo <= n4410_li;
    n4413_lo <= n4413_li;
    n4416_lo <= n4416_li;
    n4419_lo <= n4419_li;
    n4422_lo <= n4422_li;
    n4425_lo <= n4425_li;
    n4428_lo <= n4428_li;
    n4431_lo <= n4431_li;
    n4434_lo <= n4434_li;
    n4437_lo <= n4437_li;
    n4440_lo <= n4440_li;
    n4443_lo <= n4443_li;
    n4446_lo <= n4446_li;
    n4449_lo <= n4449_li;
    n4452_lo <= n4452_li;
    n4455_lo <= n4455_li;
    n4458_lo <= n4458_li;
    n4461_lo <= n4461_li;
    n4464_lo <= n4464_li;
    n4467_lo <= n4467_li;
    n4470_lo <= n4470_li;
    n4473_lo <= n4473_li;
    n4476_lo <= n4476_li;
    n4479_lo <= n4479_li;
    n4482_lo <= n4482_li;
    n4485_lo <= n4485_li;
    n4488_lo <= n4488_li;
    n4491_lo <= n4491_li;
    n4494_lo <= n4494_li;
    n4497_lo <= n4497_li;
    n4500_lo <= n4500_li;
    n4503_lo <= n4503_li;
    n4506_lo <= n4506_li;
    n4509_lo <= n4509_li;
    n4512_lo <= n4512_li;
    n4515_lo <= n4515_li;
    n4518_lo <= n4518_li;
    n4521_lo <= n4521_li;
    n4524_lo <= n4524_li;
    n4527_lo <= n4527_li;
    n4530_lo <= n4530_li;
    n4533_lo <= n4533_li;
    n4536_lo <= n4536_li;
    n4539_lo <= n4539_li;
    n4542_lo <= n4542_li;
    n4545_lo <= n4545_li;
    n4548_lo <= n4548_li;
    n4551_lo <= n4551_li;
    n4554_lo <= n4554_li;
    n4557_lo <= n4557_li;
    n4560_lo <= n4560_li;
    n4563_lo <= n4563_li;
    n4566_lo <= n4566_li;
    n4569_lo <= n4569_li;
    n4572_lo <= n4572_li;
    n4575_lo <= n4575_li;
    n4578_lo <= n4578_li;
    n4581_lo <= n4581_li;
    n4584_lo <= n4584_li;
    n4587_lo <= n4587_li;
    n4590_lo <= n4590_li;
    n4593_lo <= n4593_li;
    n4596_lo <= n4596_li;
    n4599_lo <= n4599_li;
    n4602_lo <= n4602_li;
    n4605_lo <= n4605_li;
    n4608_lo <= n4608_li;
    n4611_lo <= n4611_li;
    n4614_lo <= n4614_li;
    n4617_lo <= n4617_li;
    n4620_lo <= n4620_li;
    n4623_lo <= n4623_li;
    n4626_lo <= n4626_li;
    n4629_lo <= n4629_li;
    n4632_lo <= n4632_li;
    n4635_lo <= n4635_li;
    n4638_lo <= n4638_li;
    n4641_lo <= n4641_li;
    n4644_lo <= n4644_li;
    n4647_lo <= n4647_li;
    n4650_lo <= n4650_li;
    n4653_lo <= n4653_li;
    n4656_lo <= n4656_li;
    n4659_lo <= n4659_li;
    n4662_lo <= n4662_li;
    n4665_lo <= n4665_li;
    n4668_lo <= n4668_li;
    n4671_lo <= n4671_li;
    n4674_lo <= n4674_li;
    n4677_lo <= n4677_li;
    n4680_lo <= n4680_li;
    n4683_lo <= n4683_li;
    n4686_lo <= n4686_li;
    n4689_lo <= n4689_li;
    n4692_lo <= n4692_li;
    n4695_lo <= n4695_li;
    n4698_lo <= n4698_li;
    n4701_lo <= n4701_li;
    n4704_lo <= n4704_li;
    n4707_lo <= n4707_li;
    n4710_lo <= n4710_li;
    n4713_lo <= n4713_li;
    n4716_lo <= n4716_li;
    n4719_lo <= n4719_li;
    n4722_lo <= n4722_li;
    n4725_lo <= n4725_li;
    n4728_lo <= n4728_li;
    n4731_lo <= n4731_li;
    n4734_lo <= n4734_li;
    n4737_lo <= n4737_li;
    n4740_lo <= n4740_li;
    n4743_lo <= n4743_li;
  end
  initial begin
    n2610_lo <= 1'b0;
    n2613_lo <= 1'b0;
    n2616_lo <= 1'b0;
    n2619_lo <= 1'b0;
    n2622_lo <= 1'b0;
    n2625_lo <= 1'b0;
    n2628_lo <= 1'b0;
    n2631_lo <= 1'b0;
    n2634_lo <= 1'b0;
    n2637_lo <= 1'b0;
    n2640_lo <= 1'b0;
    n2643_lo <= 1'b0;
    n2646_lo <= 1'b0;
    n2649_lo <= 1'b0;
    n2652_lo <= 1'b0;
    n2655_lo <= 1'b0;
    n2658_lo <= 1'b0;
    n2661_lo <= 1'b0;
    n2664_lo <= 1'b0;
    n2667_lo <= 1'b0;
    n2670_lo <= 1'b0;
    n2673_lo <= 1'b0;
    n2676_lo <= 1'b0;
    n2679_lo <= 1'b0;
    n2682_lo <= 1'b0;
    n2685_lo <= 1'b0;
    n2688_lo <= 1'b0;
    n2691_lo <= 1'b0;
    n2694_lo <= 1'b0;
    n2697_lo <= 1'b0;
    n2700_lo <= 1'b0;
    n2703_lo <= 1'b0;
    n2706_lo <= 1'b0;
    n2709_lo <= 1'b0;
    n2712_lo <= 1'b0;
    n2715_lo <= 1'b0;
    n2718_lo <= 1'b0;
    n2721_lo <= 1'b0;
    n2724_lo <= 1'b0;
    n2727_lo <= 1'b0;
    n2730_lo <= 1'b0;
    n2733_lo <= 1'b0;
    n2736_lo <= 1'b0;
    n2739_lo <= 1'b0;
    n2742_lo <= 1'b0;
    n2745_lo <= 1'b0;
    n2748_lo <= 1'b0;
    n2751_lo <= 1'b0;
    n2754_lo <= 1'b0;
    n2757_lo <= 1'b0;
    n2760_lo <= 1'b0;
    n2763_lo <= 1'b0;
    n2766_lo <= 1'b0;
    n2769_lo <= 1'b0;
    n2772_lo <= 1'b0;
    n2775_lo <= 1'b0;
    n2778_lo <= 1'b0;
    n2781_lo <= 1'b0;
    n2784_lo <= 1'b0;
    n2787_lo <= 1'b0;
    n2790_lo <= 1'b0;
    n2793_lo <= 1'b0;
    n2796_lo <= 1'b0;
    n2799_lo <= 1'b0;
    n2802_lo <= 1'b0;
    n2805_lo <= 1'b0;
    n2808_lo <= 1'b0;
    n2811_lo <= 1'b0;
    n2814_lo <= 1'b0;
    n2817_lo <= 1'b0;
    n2820_lo <= 1'b0;
    n2823_lo <= 1'b0;
    n2826_lo <= 1'b0;
    n2829_lo <= 1'b0;
    n2832_lo <= 1'b0;
    n2835_lo <= 1'b0;
    n2838_lo <= 1'b0;
    n2841_lo <= 1'b0;
    n2844_lo <= 1'b0;
    n2847_lo <= 1'b0;
    n2850_lo <= 1'b0;
    n2853_lo <= 1'b0;
    n2856_lo <= 1'b0;
    n2859_lo <= 1'b0;
    n2862_lo <= 1'b0;
    n2865_lo <= 1'b0;
    n2868_lo <= 1'b0;
    n2871_lo <= 1'b0;
    n2874_lo <= 1'b0;
    n2877_lo <= 1'b0;
    n2880_lo <= 1'b0;
    n2883_lo <= 1'b0;
    n2886_lo <= 1'b0;
    n2889_lo <= 1'b0;
    n2892_lo <= 1'b0;
    n2895_lo <= 1'b0;
    n2898_lo <= 1'b0;
    n2901_lo <= 1'b0;
    n2904_lo <= 1'b0;
    n2907_lo <= 1'b0;
    n2910_lo <= 1'b0;
    n2913_lo <= 1'b0;
    n2916_lo <= 1'b0;
    n2919_lo <= 1'b0;
    n2922_lo <= 1'b0;
    n2925_lo <= 1'b0;
    n2928_lo <= 1'b0;
    n2931_lo <= 1'b0;
    n2934_lo <= 1'b0;
    n2937_lo <= 1'b0;
    n2940_lo <= 1'b0;
    n2943_lo <= 1'b0;
    n2946_lo <= 1'b0;
    n2949_lo <= 1'b0;
    n2952_lo <= 1'b0;
    n2955_lo <= 1'b0;
    n2958_lo <= 1'b0;
    n2961_lo <= 1'b0;
    n2964_lo <= 1'b0;
    n2967_lo <= 1'b0;
    n2970_lo <= 1'b0;
    n2973_lo <= 1'b0;
    n2976_lo <= 1'b0;
    n2979_lo <= 1'b0;
    n2982_lo <= 1'b0;
    n2985_lo <= 1'b0;
    n2988_lo <= 1'b0;
    n2991_lo <= 1'b0;
    n2994_lo <= 1'b0;
    n2997_lo <= 1'b0;
    n3000_lo <= 1'b0;
    n3003_lo <= 1'b0;
    n3006_lo <= 1'b0;
    n3009_lo <= 1'b0;
    n3012_lo <= 1'b0;
    n3015_lo <= 1'b0;
    n3018_lo <= 1'b0;
    n3021_lo <= 1'b0;
    n3024_lo <= 1'b0;
    n3027_lo <= 1'b0;
    n3030_lo <= 1'b0;
    n3033_lo <= 1'b0;
    n3036_lo <= 1'b0;
    n3039_lo <= 1'b0;
    n3042_lo <= 1'b0;
    n3045_lo <= 1'b0;
    n3048_lo <= 1'b0;
    n3051_lo <= 1'b0;
    n3054_lo <= 1'b0;
    n3057_lo <= 1'b0;
    n3060_lo <= 1'b0;
    n3063_lo <= 1'b0;
    n3066_lo <= 1'b0;
    n3069_lo <= 1'b0;
    n3072_lo <= 1'b0;
    n3075_lo <= 1'b0;
    n3078_lo <= 1'b0;
    n3081_lo <= 1'b0;
    n3084_lo <= 1'b0;
    n3087_lo <= 1'b0;
    n3090_lo <= 1'b0;
    n3093_lo <= 1'b0;
    n3096_lo <= 1'b0;
    n3099_lo <= 1'b0;
    n3102_lo <= 1'b0;
    n3105_lo <= 1'b0;
    n3108_lo <= 1'b0;
    n3111_lo <= 1'b0;
    n3114_lo <= 1'b0;
    n3117_lo <= 1'b0;
    n3120_lo <= 1'b0;
    n3123_lo <= 1'b0;
    n3126_lo <= 1'b0;
    n3129_lo <= 1'b0;
    n3132_lo <= 1'b0;
    n3135_lo <= 1'b0;
    n3138_lo <= 1'b0;
    n3141_lo <= 1'b0;
    n3144_lo <= 1'b0;
    n3147_lo <= 1'b0;
    n3150_lo <= 1'b0;
    n3153_lo <= 1'b0;
    n3156_lo <= 1'b0;
    n3159_lo <= 1'b0;
    n3162_lo <= 1'b0;
    n3165_lo <= 1'b0;
    n3168_lo <= 1'b0;
    n3171_lo <= 1'b0;
    n3174_lo <= 1'b0;
    n3177_lo <= 1'b0;
    n3180_lo <= 1'b0;
    n3183_lo <= 1'b0;
    n3186_lo <= 1'b0;
    n3189_lo <= 1'b0;
    n3192_lo <= 1'b0;
    n3195_lo <= 1'b0;
    n3198_lo <= 1'b0;
    n3201_lo <= 1'b0;
    n3204_lo <= 1'b0;
    n3207_lo <= 1'b0;
    n3210_lo <= 1'b0;
    n3213_lo <= 1'b0;
    n3216_lo <= 1'b0;
    n3219_lo <= 1'b0;
    n3222_lo <= 1'b0;
    n3225_lo <= 1'b0;
    n3228_lo <= 1'b0;
    n3231_lo <= 1'b0;
    n3234_lo <= 1'b0;
    n3237_lo <= 1'b0;
    n3240_lo <= 1'b0;
    n3243_lo <= 1'b0;
    n3246_lo <= 1'b0;
    n3249_lo <= 1'b0;
    n3252_lo <= 1'b0;
    n3255_lo <= 1'b0;
    n3258_lo <= 1'b0;
    n3261_lo <= 1'b0;
    n3264_lo <= 1'b0;
    n3267_lo <= 1'b0;
    n3270_lo <= 1'b0;
    n3273_lo <= 1'b0;
    n3276_lo <= 1'b0;
    n3279_lo <= 1'b0;
    n3282_lo <= 1'b0;
    n3285_lo <= 1'b0;
    n3288_lo <= 1'b0;
    n3291_lo <= 1'b0;
    n3294_lo <= 1'b0;
    n3297_lo <= 1'b0;
    n3300_lo <= 1'b0;
    n3303_lo <= 1'b0;
    n3306_lo <= 1'b0;
    n3309_lo <= 1'b0;
    n3312_lo <= 1'b0;
    n3315_lo <= 1'b0;
    n3318_lo <= 1'b0;
    n3321_lo <= 1'b0;
    n3324_lo <= 1'b0;
    n3327_lo <= 1'b0;
    n3330_lo <= 1'b0;
    n3333_lo <= 1'b0;
    n3336_lo <= 1'b0;
    n3339_lo <= 1'b0;
    n3342_lo <= 1'b0;
    n3345_lo <= 1'b0;
    n3348_lo <= 1'b0;
    n3351_lo <= 1'b0;
    n3354_lo <= 1'b0;
    n3357_lo <= 1'b0;
    n3360_lo <= 1'b0;
    n3363_lo <= 1'b0;
    n3366_lo <= 1'b0;
    n3369_lo <= 1'b0;
    n3372_lo <= 1'b0;
    n3375_lo <= 1'b0;
    n3378_lo <= 1'b0;
    n3381_lo <= 1'b0;
    n3384_lo <= 1'b0;
    n3387_lo <= 1'b0;
    n3390_lo <= 1'b0;
    n3393_lo <= 1'b0;
    n3396_lo <= 1'b0;
    n3399_lo <= 1'b0;
    n3402_lo <= 1'b0;
    n3405_lo <= 1'b0;
    n3408_lo <= 1'b0;
    n3411_lo <= 1'b0;
    n3414_lo <= 1'b0;
    n3417_lo <= 1'b0;
    n3420_lo <= 1'b0;
    n3423_lo <= 1'b0;
    n3426_lo <= 1'b0;
    n3429_lo <= 1'b0;
    n3432_lo <= 1'b0;
    n3435_lo <= 1'b0;
    n3438_lo <= 1'b0;
    n3441_lo <= 1'b0;
    n3444_lo <= 1'b0;
    n3447_lo <= 1'b0;
    n3450_lo <= 1'b0;
    n3453_lo <= 1'b0;
    n3456_lo <= 1'b0;
    n3459_lo <= 1'b0;
    n3462_lo <= 1'b0;
    n3465_lo <= 1'b0;
    n3468_lo <= 1'b0;
    n3471_lo <= 1'b0;
    n3474_lo <= 1'b0;
    n3477_lo <= 1'b0;
    n3480_lo <= 1'b0;
    n3483_lo <= 1'b0;
    n3486_lo <= 1'b0;
    n3489_lo <= 1'b0;
    n3492_lo <= 1'b0;
    n3495_lo <= 1'b0;
    n3498_lo <= 1'b0;
    n3501_lo <= 1'b0;
    n3504_lo <= 1'b0;
    n3507_lo <= 1'b0;
    n3510_lo <= 1'b0;
    n3513_lo <= 1'b0;
    n3516_lo <= 1'b0;
    n3519_lo <= 1'b0;
    n3522_lo <= 1'b0;
    n3525_lo <= 1'b0;
    n3528_lo <= 1'b0;
    n3531_lo <= 1'b0;
    n3534_lo <= 1'b0;
    n3537_lo <= 1'b0;
    n3540_lo <= 1'b0;
    n3543_lo <= 1'b0;
    n3546_lo <= 1'b0;
    n3549_lo <= 1'b0;
    n3552_lo <= 1'b0;
    n3555_lo <= 1'b0;
    n3558_lo <= 1'b0;
    n3561_lo <= 1'b0;
    n3564_lo <= 1'b0;
    n3567_lo <= 1'b0;
    n3570_lo <= 1'b0;
    n3573_lo <= 1'b0;
    n3576_lo <= 1'b0;
    n3579_lo <= 1'b0;
    n3582_lo <= 1'b0;
    n3585_lo <= 1'b0;
    n3588_lo <= 1'b0;
    n3591_lo <= 1'b0;
    n3594_lo <= 1'b0;
    n3597_lo <= 1'b0;
    n3600_lo <= 1'b0;
    n3603_lo <= 1'b0;
    n3606_lo <= 1'b0;
    n3609_lo <= 1'b0;
    n3612_lo <= 1'b0;
    n3615_lo <= 1'b0;
    n3618_lo <= 1'b0;
    n3621_lo <= 1'b0;
    n3624_lo <= 1'b0;
    n3627_lo <= 1'b0;
    n3630_lo <= 1'b0;
    n3633_lo <= 1'b0;
    n3636_lo <= 1'b0;
    n3639_lo <= 1'b0;
    n3642_lo <= 1'b0;
    n3645_lo <= 1'b0;
    n3648_lo <= 1'b0;
    n3651_lo <= 1'b0;
    n3654_lo <= 1'b0;
    n3657_lo <= 1'b0;
    n3660_lo <= 1'b0;
    n3663_lo <= 1'b0;
    n3666_lo <= 1'b0;
    n3669_lo <= 1'b0;
    n3672_lo <= 1'b0;
    n3675_lo <= 1'b0;
    n3678_lo <= 1'b0;
    n3681_lo <= 1'b0;
    n3684_lo <= 1'b0;
    n3687_lo <= 1'b0;
    n3690_lo <= 1'b0;
    n3693_lo <= 1'b0;
    n3696_lo <= 1'b0;
    n3699_lo <= 1'b0;
    n3702_lo <= 1'b0;
    n3705_lo <= 1'b0;
    n3708_lo <= 1'b0;
    n3711_lo <= 1'b0;
    n3714_lo <= 1'b0;
    n3717_lo <= 1'b0;
    n3720_lo <= 1'b0;
    n3723_lo <= 1'b0;
    n3726_lo <= 1'b0;
    n3729_lo <= 1'b0;
    n3732_lo <= 1'b0;
    n3735_lo <= 1'b0;
    n3738_lo <= 1'b0;
    n3741_lo <= 1'b0;
    n3744_lo <= 1'b0;
    n3747_lo <= 1'b0;
    n3750_lo <= 1'b0;
    n3753_lo <= 1'b0;
    n3756_lo <= 1'b0;
    n3759_lo <= 1'b0;
    n3762_lo <= 1'b0;
    n3765_lo <= 1'b0;
    n3768_lo <= 1'b0;
    n3771_lo <= 1'b0;
    n3774_lo <= 1'b0;
    n3777_lo <= 1'b0;
    n3780_lo <= 1'b0;
    n3783_lo <= 1'b0;
    n3786_lo <= 1'b0;
    n3789_lo <= 1'b0;
    n3792_lo <= 1'b0;
    n3795_lo <= 1'b0;
    n3798_lo <= 1'b0;
    n3801_lo <= 1'b0;
    n3804_lo <= 1'b0;
    n3807_lo <= 1'b0;
    n3810_lo <= 1'b0;
    n3813_lo <= 1'b0;
    n3816_lo <= 1'b0;
    n3819_lo <= 1'b0;
    n3822_lo <= 1'b0;
    n3825_lo <= 1'b0;
    n3828_lo <= 1'b0;
    n3831_lo <= 1'b0;
    n3834_lo <= 1'b0;
    n3837_lo <= 1'b0;
    n3840_lo <= 1'b0;
    n3843_lo <= 1'b0;
    n3846_lo <= 1'b0;
    n3849_lo <= 1'b0;
    n3852_lo <= 1'b0;
    n3855_lo <= 1'b0;
    n3858_lo <= 1'b0;
    n3861_lo <= 1'b0;
    n3864_lo <= 1'b0;
    n3867_lo <= 1'b0;
    n3870_lo <= 1'b0;
    n3873_lo <= 1'b0;
    n3876_lo <= 1'b0;
    n3879_lo <= 1'b0;
    n3882_lo <= 1'b0;
    n3885_lo <= 1'b0;
    n3888_lo <= 1'b0;
    n3891_lo <= 1'b0;
    n3894_lo <= 1'b0;
    n3897_lo <= 1'b0;
    n3900_lo <= 1'b0;
    n3903_lo <= 1'b0;
    n3906_lo <= 1'b0;
    n3909_lo <= 1'b0;
    n3912_lo <= 1'b0;
    n3915_lo <= 1'b0;
    n3918_lo <= 1'b0;
    n3921_lo <= 1'b0;
    n3924_lo <= 1'b0;
    n3927_lo <= 1'b0;
    n3930_lo <= 1'b0;
    n3933_lo <= 1'b0;
    n3936_lo <= 1'b0;
    n3939_lo <= 1'b0;
    n3942_lo <= 1'b0;
    n3945_lo <= 1'b0;
    n3948_lo <= 1'b0;
    n3951_lo <= 1'b0;
    n3954_lo <= 1'b0;
    n3957_lo <= 1'b0;
    n3960_lo <= 1'b0;
    n3963_lo <= 1'b0;
    n3966_lo <= 1'b0;
    n3969_lo <= 1'b0;
    n3972_lo <= 1'b0;
    n3975_lo <= 1'b0;
    n3978_lo <= 1'b0;
    n3981_lo <= 1'b0;
    n3984_lo <= 1'b0;
    n3987_lo <= 1'b0;
    n3990_lo <= 1'b0;
    n3993_lo <= 1'b0;
    n3996_lo <= 1'b0;
    n3999_lo <= 1'b0;
    n4002_lo <= 1'b0;
    n4005_lo <= 1'b0;
    n4008_lo <= 1'b0;
    n4011_lo <= 1'b0;
    n4014_lo <= 1'b0;
    n4017_lo <= 1'b0;
    n4020_lo <= 1'b0;
    n4023_lo <= 1'b0;
    n4026_lo <= 1'b0;
    n4029_lo <= 1'b0;
    n4032_lo <= 1'b0;
    n4035_lo <= 1'b0;
    n4038_lo <= 1'b0;
    n4041_lo <= 1'b0;
    n4044_lo <= 1'b0;
    n4047_lo <= 1'b0;
    n4050_lo <= 1'b0;
    n4053_lo <= 1'b0;
    n4056_lo <= 1'b0;
    n4059_lo <= 1'b0;
    n4062_lo <= 1'b0;
    n4065_lo <= 1'b0;
    n4068_lo <= 1'b0;
    n4071_lo <= 1'b0;
    n4074_lo <= 1'b0;
    n4077_lo <= 1'b0;
    n4080_lo <= 1'b0;
    n4083_lo <= 1'b0;
    n4086_lo <= 1'b0;
    n4089_lo <= 1'b0;
    n4092_lo <= 1'b0;
    n4095_lo <= 1'b0;
    n4098_lo <= 1'b0;
    n4101_lo <= 1'b0;
    n4104_lo <= 1'b0;
    n4107_lo <= 1'b0;
    n4110_lo <= 1'b0;
    n4113_lo <= 1'b0;
    n4116_lo <= 1'b0;
    n4119_lo <= 1'b0;
    n4122_lo <= 1'b0;
    n4125_lo <= 1'b0;
    n4128_lo <= 1'b0;
    n4131_lo <= 1'b0;
    n4134_lo <= 1'b0;
    n4137_lo <= 1'b0;
    n4140_lo <= 1'b0;
    n4143_lo <= 1'b0;
    n4146_lo <= 1'b0;
    n4149_lo <= 1'b0;
    n4152_lo <= 1'b0;
    n4155_lo <= 1'b0;
    n4158_lo <= 1'b0;
    n4161_lo <= 1'b0;
    n4164_lo <= 1'b0;
    n4167_lo <= 1'b0;
    n4170_lo <= 1'b0;
    n4173_lo <= 1'b0;
    n4176_lo <= 1'b0;
    n4179_lo <= 1'b0;
    n4182_lo <= 1'b0;
    n4185_lo <= 1'b0;
    n4188_lo <= 1'b0;
    n4191_lo <= 1'b0;
    n4194_lo <= 1'b0;
    n4197_lo <= 1'b0;
    n4200_lo <= 1'b0;
    n4203_lo <= 1'b0;
    n4206_lo <= 1'b0;
    n4209_lo <= 1'b0;
    n4212_lo <= 1'b0;
    n4215_lo <= 1'b0;
    n4218_lo <= 1'b0;
    n4221_lo <= 1'b0;
    n4224_lo <= 1'b0;
    n4227_lo <= 1'b0;
    n4230_lo <= 1'b0;
    n4233_lo <= 1'b0;
    n4236_lo <= 1'b0;
    n4239_lo <= 1'b0;
    n4242_lo <= 1'b0;
    n4245_lo <= 1'b0;
    n4248_lo <= 1'b0;
    n4251_lo <= 1'b0;
    n4254_lo <= 1'b0;
    n4257_lo <= 1'b0;
    n4260_lo <= 1'b0;
    n4263_lo <= 1'b0;
    n4266_lo <= 1'b0;
    n4269_lo <= 1'b0;
    n4272_lo <= 1'b0;
    n4275_lo <= 1'b0;
    n4278_lo <= 1'b0;
    n4281_lo <= 1'b0;
    n4284_lo <= 1'b0;
    n4287_lo <= 1'b0;
    n4290_lo <= 1'b0;
    n4293_lo <= 1'b0;
    n4296_lo <= 1'b0;
    n4299_lo <= 1'b0;
    n4302_lo <= 1'b0;
    n4305_lo <= 1'b0;
    n4308_lo <= 1'b0;
    n4311_lo <= 1'b0;
    n4314_lo <= 1'b0;
    n4317_lo <= 1'b0;
    n4320_lo <= 1'b0;
    n4323_lo <= 1'b0;
    n4326_lo <= 1'b0;
    n4329_lo <= 1'b0;
    n4332_lo <= 1'b0;
    n4335_lo <= 1'b0;
    n4338_lo <= 1'b0;
    n4341_lo <= 1'b0;
    n4344_lo <= 1'b0;
    n4347_lo <= 1'b0;
    n4350_lo <= 1'b0;
    n4353_lo <= 1'b0;
    n4356_lo <= 1'b0;
    n4359_lo <= 1'b0;
    n4362_lo <= 1'b0;
    n4365_lo <= 1'b0;
    n4368_lo <= 1'b0;
    n4371_lo <= 1'b0;
    n4374_lo <= 1'b0;
    n4377_lo <= 1'b0;
    n4380_lo <= 1'b0;
    n4383_lo <= 1'b0;
    n4386_lo <= 1'b0;
    n4389_lo <= 1'b0;
    n4392_lo <= 1'b0;
    n4395_lo <= 1'b0;
    n4398_lo <= 1'b0;
    n4401_lo <= 1'b0;
    n4404_lo <= 1'b0;
    n4407_lo <= 1'b0;
    n4410_lo <= 1'b0;
    n4413_lo <= 1'b0;
    n4416_lo <= 1'b0;
    n4419_lo <= 1'b0;
    n4422_lo <= 1'b0;
    n4425_lo <= 1'b0;
    n4428_lo <= 1'b0;
    n4431_lo <= 1'b0;
    n4434_lo <= 1'b0;
    n4437_lo <= 1'b0;
    n4440_lo <= 1'b0;
    n4443_lo <= 1'b0;
    n4446_lo <= 1'b0;
    n4449_lo <= 1'b0;
    n4452_lo <= 1'b0;
    n4455_lo <= 1'b0;
    n4458_lo <= 1'b0;
    n4461_lo <= 1'b0;
    n4464_lo <= 1'b0;
    n4467_lo <= 1'b0;
    n4470_lo <= 1'b0;
    n4473_lo <= 1'b0;
    n4476_lo <= 1'b0;
    n4479_lo <= 1'b0;
    n4482_lo <= 1'b0;
    n4485_lo <= 1'b0;
    n4488_lo <= 1'b0;
    n4491_lo <= 1'b0;
    n4494_lo <= 1'b0;
    n4497_lo <= 1'b0;
    n4500_lo <= 1'b0;
    n4503_lo <= 1'b0;
    n4506_lo <= 1'b0;
    n4509_lo <= 1'b0;
    n4512_lo <= 1'b0;
    n4515_lo <= 1'b0;
    n4518_lo <= 1'b0;
    n4521_lo <= 1'b0;
    n4524_lo <= 1'b0;
    n4527_lo <= 1'b0;
    n4530_lo <= 1'b0;
    n4533_lo <= 1'b0;
    n4536_lo <= 1'b0;
    n4539_lo <= 1'b0;
    n4542_lo <= 1'b0;
    n4545_lo <= 1'b0;
    n4548_lo <= 1'b0;
    n4551_lo <= 1'b0;
    n4554_lo <= 1'b0;
    n4557_lo <= 1'b0;
    n4560_lo <= 1'b0;
    n4563_lo <= 1'b0;
    n4566_lo <= 1'b0;
    n4569_lo <= 1'b0;
    n4572_lo <= 1'b0;
    n4575_lo <= 1'b0;
    n4578_lo <= 1'b0;
    n4581_lo <= 1'b0;
    n4584_lo <= 1'b0;
    n4587_lo <= 1'b0;
    n4590_lo <= 1'b0;
    n4593_lo <= 1'b0;
    n4596_lo <= 1'b0;
    n4599_lo <= 1'b0;
    n4602_lo <= 1'b0;
    n4605_lo <= 1'b0;
    n4608_lo <= 1'b0;
    n4611_lo <= 1'b0;
    n4614_lo <= 1'b0;
    n4617_lo <= 1'b0;
    n4620_lo <= 1'b0;
    n4623_lo <= 1'b0;
    n4626_lo <= 1'b0;
    n4629_lo <= 1'b0;
    n4632_lo <= 1'b0;
    n4635_lo <= 1'b0;
    n4638_lo <= 1'b0;
    n4641_lo <= 1'b0;
    n4644_lo <= 1'b0;
    n4647_lo <= 1'b0;
    n4650_lo <= 1'b0;
    n4653_lo <= 1'b0;
    n4656_lo <= 1'b0;
    n4659_lo <= 1'b0;
    n4662_lo <= 1'b0;
    n4665_lo <= 1'b0;
    n4668_lo <= 1'b0;
    n4671_lo <= 1'b0;
    n4674_lo <= 1'b0;
    n4677_lo <= 1'b0;
    n4680_lo <= 1'b0;
    n4683_lo <= 1'b0;
    n4686_lo <= 1'b0;
    n4689_lo <= 1'b0;
    n4692_lo <= 1'b0;
    n4695_lo <= 1'b0;
    n4698_lo <= 1'b0;
    n4701_lo <= 1'b0;
    n4704_lo <= 1'b0;
    n4707_lo <= 1'b0;
    n4710_lo <= 1'b0;
    n4713_lo <= 1'b0;
    n4716_lo <= 1'b0;
    n4719_lo <= 1'b0;
    n4722_lo <= 1'b0;
    n4725_lo <= 1'b0;
    n4728_lo <= 1'b0;
    n4731_lo <= 1'b0;
    n4734_lo <= 1'b0;
    n4737_lo <= 1'b0;
    n4740_lo <= 1'b0;
    n4743_lo <= 1'b0;
  end
endmodule


