
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  G1324,
  G1325,
  G1326,
  G1327,
  G1328,
  G1329,
  G1330,
  G1331,
  G1332,
  G1333,
  G1334,
  G1335,
  G1336,
  G1337,
  G1338,
  G1339,
  G1340,
  G1341,
  G1342,
  G1343,
  G1344,
  G1345,
  G1346,
  G1347,
  G1348,
  G1349,
  G1350,
  G1351,
  G1352,
  G1353,
  G1354,
  G1355
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;
  output G1324;output G1325;output G1326;output G1327;output G1328;output G1329;output G1330;output G1331;output G1332;output G1333;output G1334;output G1335;output G1336;output G1337;output G1338;output G1339;output G1340;output G1341;output G1342;output G1343;output G1344;output G1345;output G1346;output G1347;output G1348;output G1349;output G1350;output G1351;output G1352;output G1353;output G1354;output G1355;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire g42_p;
  wire g42_n;
  wire g43_p;
  wire g43_n;
  wire g44_p;
  wire g44_n;
  wire g45_p;
  wire g45_n;
  wire g46_p;
  wire g46_n;
  wire g47_p;
  wire g47_n;
  wire g48_p;
  wire g48_n;
  wire g49_p;
  wire g49_n;
  wire g50_p;
  wire g50_n;
  wire g51_p;
  wire g51_n;
  wire g52_p;
  wire g52_n;
  wire g53_p;
  wire g53_n;
  wire g54_p;
  wire g54_n;
  wire g55_p;
  wire g55_n;
  wire g56_p;
  wire g56_n;
  wire g57_p;
  wire g57_n;
  wire g58_p;
  wire g58_n;
  wire g59_p;
  wire g59_n;
  wire g60_p;
  wire g60_n;
  wire g61_p;
  wire g61_n;
  wire g62_p;
  wire g62_n;
  wire g63_p;
  wire g63_n;
  wire g64_p;
  wire g64_n;
  wire g65_p;
  wire g65_n;
  wire g66_p;
  wire g66_n;
  wire g67_p;
  wire g67_n;
  wire g68_p;
  wire g68_n;
  wire g69_p;
  wire g69_n;
  wire g70_p;
  wire g70_n;
  wire g71_p;
  wire g71_n;
  wire g72_p;
  wire g72_n;
  wire g73_p;
  wire g73_n;
  wire g74_p;
  wire g74_n;
  wire g75_p;
  wire g75_n;
  wire g76_p;
  wire g76_n;
  wire g77_p;
  wire g77_n;
  wire g78_p;
  wire g78_n;
  wire g79_p;
  wire g79_n;
  wire g80_p;
  wire g80_n;
  wire g81_p;
  wire g81_n;
  wire g82_p;
  wire g82_n;
  wire g83_p;
  wire g83_n;
  wire g84_p;
  wire g84_n;
  wire g85_p;
  wire g85_n;
  wire g86_p;
  wire g86_n;
  wire g87_p;
  wire g87_n;
  wire g88_p;
  wire g88_n;
  wire g89_p;
  wire g89_n;
  wire g90_p;
  wire g90_n;
  wire g91_p;
  wire g91_n;
  wire g92_p;
  wire g92_n;
  wire g93_p;
  wire g93_n;
  wire g94_p;
  wire g94_n;
  wire g95_p;
  wire g95_n;
  wire g96_p;
  wire g96_n;
  wire g97_p;
  wire g97_n;
  wire g98_p;
  wire g98_n;
  wire g99_p;
  wire g99_n;
  wire g100_p;
  wire g100_n;
  wire g101_p;
  wire g101_n;
  wire g102_p;
  wire g102_n;
  wire g103_p;
  wire g103_n;
  wire g104_p;
  wire g104_n;
  wire g105_p;
  wire g105_n;
  wire g106_p;
  wire g106_n;
  wire g107_p;
  wire g107_n;
  wire g108_p;
  wire g108_n;
  wire g109_p;
  wire g109_n;
  wire g110_p;
  wire g110_n;
  wire g111_p;
  wire g111_n;
  wire g112_p;
  wire g112_n;
  wire g113_p;
  wire g113_n;
  wire g114_p;
  wire g114_n;
  wire g115_p;
  wire g115_n;
  wire g116_p;
  wire g116_n;
  wire g117_p;
  wire g117_n;
  wire g118_p;
  wire g118_n;
  wire g119_p;
  wire g119_n;
  wire g120_p;
  wire g120_n;
  wire g121_p;
  wire g121_n;
  wire g122_p;
  wire g122_n;
  wire g123_p;
  wire g123_n;
  wire g124_p;
  wire g124_n;
  wire g125_p;
  wire g125_n;
  wire g126_p;
  wire g126_n;
  wire g127_p;
  wire g127_n;
  wire g128_p;
  wire g128_n;
  wire g129_p;
  wire g129_n;
  wire g130_p;
  wire g130_n;
  wire g131_p;
  wire g131_n;
  wire g132_p;
  wire g132_n;
  wire g133_p;
  wire g133_n;
  wire g134_p;
  wire g134_n;
  wire g135_p;
  wire g135_n;
  wire g136_p;
  wire g136_n;
  wire g137_p;
  wire g137_n;
  wire g138_p;
  wire g138_n;
  wire g139_p;
  wire g139_n;
  wire g140_p;
  wire g140_n;
  wire g141_p;
  wire g141_n;
  wire g142_p;
  wire g142_n;
  wire g143_p;
  wire g143_n;
  wire g144_p;
  wire g144_n;
  wire g145_p;
  wire g145_n;
  wire g146_p;
  wire g146_n;
  wire g147_p;
  wire g147_n;
  wire g148_p;
  wire g148_n;
  wire g149_p;
  wire g149_n;
  wire g150_p;
  wire g150_n;
  wire g151_p;
  wire g151_n;
  wire g152_p;
  wire g152_n;
  wire g153_p;
  wire g153_n;
  wire g154_p;
  wire g154_n;
  wire g155_p;
  wire g155_n;
  wire g156_p;
  wire g156_n;
  wire g157_p;
  wire g157_n;
  wire g158_p;
  wire g158_n;
  wire g159_p;
  wire g159_n;
  wire g160_p;
  wire g160_n;
  wire g161_p;
  wire g161_n;
  wire g162_p;
  wire g162_n;
  wire g163_p;
  wire g163_n;
  wire g164_p;
  wire g164_n;
  wire g165_p;
  wire g165_n;
  wire g166_p;
  wire g166_n;
  wire g167_p;
  wire g167_n;
  wire g168_p;
  wire g168_n;
  wire g169_p;
  wire g169_n;
  wire g170_p;
  wire g170_n;
  wire g171_p;
  wire g171_n;
  wire g172_p;
  wire g172_n;
  wire g173_p;
  wire g173_n;
  wire g174_p;
  wire g174_n;
  wire g175_p;
  wire g175_n;
  wire g176_p;
  wire g176_n;
  wire g177_p;
  wire g177_n;
  wire g178_p;
  wire g178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire G9_n_spl_;
  wire G9_n_spl_0;
  wire G9_n_spl_00;
  wire G9_n_spl_1;
  wire G13_n_spl_;
  wire G13_n_spl_0;
  wire G13_n_spl_00;
  wire G13_n_spl_1;
  wire G9_p_spl_;
  wire G9_p_spl_0;
  wire G9_p_spl_00;
  wire G9_p_spl_1;
  wire G13_p_spl_;
  wire G13_p_spl_0;
  wire G13_p_spl_00;
  wire G13_p_spl_1;
  wire G1_p_spl_;
  wire G1_p_spl_0;
  wire G1_p_spl_00;
  wire G1_p_spl_1;
  wire G5_n_spl_;
  wire G5_n_spl_0;
  wire G5_n_spl_00;
  wire G5_n_spl_1;
  wire G1_n_spl_;
  wire G1_n_spl_0;
  wire G1_n_spl_00;
  wire G1_n_spl_1;
  wire G5_p_spl_;
  wire G5_p_spl_0;
  wire G5_p_spl_00;
  wire G5_p_spl_1;
  wire g44_n_spl_;
  wire g47_n_spl_;
  wire g44_p_spl_;
  wire g47_p_spl_;
  wire G41_p_spl_;
  wire G41_p_spl_0;
  wire G41_p_spl_00;
  wire G41_p_spl_01;
  wire G41_p_spl_1;
  wire G41_p_spl_10;
  wire G41_p_spl_11;
  wire G41_n_spl_;
  wire G41_n_spl_0;
  wire G41_n_spl_00;
  wire G41_n_spl_01;
  wire G41_n_spl_1;
  wire G41_n_spl_10;
  wire G41_n_spl_11;
  wire g50_n_spl_;
  wire g51_p_spl_;
  wire g50_p_spl_;
  wire g51_n_spl_;
  wire G19_n_spl_;
  wire G19_n_spl_0;
  wire G19_n_spl_00;
  wire G19_n_spl_1;
  wire G20_n_spl_;
  wire G20_n_spl_0;
  wire G20_n_spl_00;
  wire G20_n_spl_1;
  wire G19_p_spl_;
  wire G19_p_spl_0;
  wire G19_p_spl_00;
  wire G19_p_spl_1;
  wire G20_p_spl_;
  wire G20_p_spl_0;
  wire G20_p_spl_00;
  wire G20_p_spl_1;
  wire G17_p_spl_;
  wire G17_p_spl_0;
  wire G17_p_spl_00;
  wire G17_p_spl_1;
  wire G18_n_spl_;
  wire G18_n_spl_0;
  wire G18_n_spl_00;
  wire G18_n_spl_1;
  wire G17_n_spl_;
  wire G17_n_spl_0;
  wire G17_n_spl_00;
  wire G17_n_spl_1;
  wire G18_p_spl_;
  wire G18_p_spl_0;
  wire G18_p_spl_00;
  wire G18_p_spl_1;
  wire g57_n_spl_;
  wire g60_n_spl_;
  wire g57_p_spl_;
  wire g60_p_spl_;
  wire G23_n_spl_;
  wire G23_n_spl_0;
  wire G23_n_spl_00;
  wire G23_n_spl_1;
  wire G24_n_spl_;
  wire G24_n_spl_0;
  wire G24_n_spl_00;
  wire G24_n_spl_1;
  wire G23_p_spl_;
  wire G23_p_spl_0;
  wire G23_p_spl_00;
  wire G23_p_spl_1;
  wire G24_p_spl_;
  wire G24_p_spl_0;
  wire G24_p_spl_00;
  wire G24_p_spl_1;
  wire G21_p_spl_;
  wire G21_p_spl_0;
  wire G21_p_spl_00;
  wire G21_p_spl_1;
  wire G22_n_spl_;
  wire G22_n_spl_0;
  wire G22_n_spl_00;
  wire G22_n_spl_1;
  wire G21_n_spl_;
  wire G21_n_spl_0;
  wire G21_n_spl_00;
  wire G21_n_spl_1;
  wire G22_p_spl_;
  wire G22_p_spl_0;
  wire G22_p_spl_00;
  wire G22_p_spl_1;
  wire g66_n_spl_;
  wire g69_n_spl_;
  wire g66_p_spl_;
  wire g69_p_spl_;
  wire g63_n_spl_;
  wire g63_n_spl_0;
  wire g63_n_spl_1;
  wire g72_n_spl_;
  wire g72_n_spl_0;
  wire g72_n_spl_1;
  wire g63_p_spl_;
  wire g63_p_spl_0;
  wire g63_p_spl_1;
  wire g72_p_spl_;
  wire g72_p_spl_0;
  wire g72_p_spl_1;
  wire g54_n_spl_;
  wire g75_p_spl_;
  wire g54_p_spl_;
  wire g75_n_spl_;
  wire G25_n_spl_;
  wire G25_n_spl_0;
  wire G25_n_spl_00;
  wire G25_n_spl_1;
  wire G29_n_spl_;
  wire G29_n_spl_0;
  wire G29_n_spl_00;
  wire G29_n_spl_1;
  wire G25_p_spl_;
  wire G25_p_spl_0;
  wire G25_p_spl_00;
  wire G25_p_spl_1;
  wire G29_p_spl_;
  wire G29_p_spl_0;
  wire G29_p_spl_00;
  wire G29_p_spl_1;
  wire g81_n_spl_;
  wire g84_n_spl_;
  wire g81_p_spl_;
  wire g84_p_spl_;
  wire g87_n_spl_;
  wire g88_p_spl_;
  wire g87_p_spl_;
  wire g88_n_spl_;
  wire G7_n_spl_;
  wire G7_n_spl_0;
  wire G7_n_spl_00;
  wire G7_n_spl_1;
  wire G8_n_spl_;
  wire G8_n_spl_0;
  wire G8_n_spl_00;
  wire G8_n_spl_1;
  wire G7_p_spl_;
  wire G7_p_spl_0;
  wire G7_p_spl_00;
  wire G7_p_spl_1;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire G8_p_spl_00;
  wire G8_p_spl_1;
  wire G6_n_spl_;
  wire G6_n_spl_0;
  wire G6_n_spl_00;
  wire G6_n_spl_1;
  wire G6_p_spl_;
  wire G6_p_spl_0;
  wire G6_p_spl_00;
  wire G6_p_spl_1;
  wire g94_n_spl_;
  wire g97_n_spl_;
  wire g94_p_spl_;
  wire g97_p_spl_;
  wire G3_n_spl_;
  wire G3_n_spl_0;
  wire G3_n_spl_00;
  wire G3_n_spl_1;
  wire G4_n_spl_;
  wire G4_n_spl_0;
  wire G4_n_spl_00;
  wire G4_n_spl_1;
  wire G3_p_spl_;
  wire G3_p_spl_0;
  wire G3_p_spl_00;
  wire G3_p_spl_1;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_00;
  wire G4_p_spl_1;
  wire G2_n_spl_;
  wire G2_n_spl_0;
  wire G2_n_spl_00;
  wire G2_n_spl_1;
  wire G2_p_spl_;
  wire G2_p_spl_0;
  wire G2_p_spl_00;
  wire G2_p_spl_1;
  wire g103_n_spl_;
  wire g106_n_spl_;
  wire g103_p_spl_;
  wire g106_p_spl_;
  wire g100_n_spl_;
  wire g100_n_spl_0;
  wire g100_n_spl_1;
  wire g109_n_spl_;
  wire g109_n_spl_0;
  wire g109_n_spl_1;
  wire g100_p_spl_;
  wire g100_p_spl_0;
  wire g100_p_spl_1;
  wire g109_p_spl_;
  wire g109_p_spl_0;
  wire g109_p_spl_1;
  wire g91_n_spl_;
  wire g112_p_spl_;
  wire g91_p_spl_;
  wire g112_n_spl_;
  wire G26_n_spl_;
  wire G26_n_spl_0;
  wire G26_n_spl_00;
  wire G26_n_spl_1;
  wire G30_n_spl_;
  wire G30_n_spl_0;
  wire G30_n_spl_00;
  wire G30_n_spl_1;
  wire G26_p_spl_;
  wire G26_p_spl_0;
  wire G26_p_spl_00;
  wire G26_p_spl_1;
  wire G30_p_spl_;
  wire G30_p_spl_0;
  wire G30_p_spl_00;
  wire G30_p_spl_1;
  wire g118_n_spl_;
  wire g121_n_spl_;
  wire g118_p_spl_;
  wire g121_p_spl_;
  wire g124_n_spl_;
  wire g125_p_spl_;
  wire g124_p_spl_;
  wire g125_n_spl_;
  wire G15_n_spl_;
  wire G15_n_spl_0;
  wire G15_n_spl_00;
  wire G15_n_spl_1;
  wire G16_n_spl_;
  wire G16_n_spl_0;
  wire G16_n_spl_00;
  wire G16_n_spl_1;
  wire G15_p_spl_;
  wire G15_p_spl_0;
  wire G15_p_spl_00;
  wire G15_p_spl_1;
  wire G16_p_spl_;
  wire G16_p_spl_0;
  wire G16_p_spl_00;
  wire G16_p_spl_1;
  wire G14_n_spl_;
  wire G14_n_spl_0;
  wire G14_n_spl_00;
  wire G14_n_spl_1;
  wire G14_p_spl_;
  wire G14_p_spl_0;
  wire G14_p_spl_00;
  wire G14_p_spl_1;
  wire g131_n_spl_;
  wire g134_n_spl_;
  wire g131_p_spl_;
  wire g134_p_spl_;
  wire G11_n_spl_;
  wire G11_n_spl_0;
  wire G11_n_spl_00;
  wire G11_n_spl_1;
  wire G12_n_spl_;
  wire G12_n_spl_0;
  wire G12_n_spl_00;
  wire G12_n_spl_1;
  wire G11_p_spl_;
  wire G11_p_spl_0;
  wire G11_p_spl_00;
  wire G11_p_spl_1;
  wire G12_p_spl_;
  wire G12_p_spl_0;
  wire G12_p_spl_00;
  wire G12_p_spl_1;
  wire G10_n_spl_;
  wire G10_n_spl_0;
  wire G10_n_spl_00;
  wire G10_n_spl_1;
  wire G10_p_spl_;
  wire G10_p_spl_0;
  wire G10_p_spl_00;
  wire G10_p_spl_1;
  wire g140_n_spl_;
  wire g143_n_spl_;
  wire g140_p_spl_;
  wire g143_p_spl_;
  wire g137_n_spl_;
  wire g137_n_spl_0;
  wire g137_n_spl_1;
  wire g146_n_spl_;
  wire g146_n_spl_0;
  wire g146_n_spl_1;
  wire g137_p_spl_;
  wire g137_p_spl_0;
  wire g137_p_spl_1;
  wire g146_p_spl_;
  wire g146_p_spl_0;
  wire g146_p_spl_1;
  wire g128_n_spl_;
  wire g149_p_spl_;
  wire g128_p_spl_;
  wire g149_n_spl_;
  wire g115_n_spl_;
  wire g115_n_spl_0;
  wire g115_n_spl_00;
  wire g115_n_spl_01;
  wire g115_n_spl_1;
  wire g115_n_spl_10;
  wire g152_p_spl_;
  wire g152_p_spl_0;
  wire g152_p_spl_00;
  wire g152_p_spl_01;
  wire g152_p_spl_1;
  wire g152_p_spl_10;
  wire g115_p_spl_;
  wire g115_p_spl_0;
  wire g115_p_spl_00;
  wire g115_p_spl_01;
  wire g115_p_spl_1;
  wire g115_p_spl_10;
  wire g152_n_spl_;
  wire g152_n_spl_0;
  wire g152_n_spl_00;
  wire g152_n_spl_01;
  wire g152_n_spl_1;
  wire g152_n_spl_10;
  wire G28_n_spl_;
  wire G28_n_spl_0;
  wire G28_n_spl_00;
  wire G28_n_spl_1;
  wire G32_n_spl_;
  wire G32_n_spl_0;
  wire G32_n_spl_00;
  wire G32_n_spl_1;
  wire G28_p_spl_;
  wire G28_p_spl_0;
  wire G28_p_spl_00;
  wire G28_p_spl_1;
  wire G32_p_spl_;
  wire G32_p_spl_0;
  wire G32_p_spl_00;
  wire G32_p_spl_1;
  wire g156_n_spl_;
  wire g159_n_spl_;
  wire g156_p_spl_;
  wire g159_p_spl_;
  wire g162_n_spl_;
  wire g163_p_spl_;
  wire g162_p_spl_;
  wire g163_n_spl_;
  wire g166_n_spl_;
  wire g169_p_spl_;
  wire g166_p_spl_;
  wire g169_n_spl_;
  wire G27_n_spl_;
  wire G27_n_spl_0;
  wire G27_n_spl_00;
  wire G27_n_spl_1;
  wire G31_n_spl_;
  wire G31_n_spl_0;
  wire G31_n_spl_00;
  wire G31_n_spl_1;
  wire G27_p_spl_;
  wire G27_p_spl_0;
  wire G27_p_spl_00;
  wire G27_p_spl_1;
  wire G31_p_spl_;
  wire G31_p_spl_0;
  wire G31_p_spl_00;
  wire G31_p_spl_1;
  wire g175_n_spl_;
  wire g178_n_spl_;
  wire g175_p_spl_;
  wire g178_p_spl_;
  wire g181_n_spl_;
  wire g182_p_spl_;
  wire g181_p_spl_;
  wire g182_n_spl_;
  wire g185_n_spl_;
  wire g188_p_spl_;
  wire g185_p_spl_;
  wire g188_n_spl_;
  wire g172_p_spl_;
  wire g172_p_spl_0;
  wire g172_p_spl_00;
  wire g172_p_spl_01;
  wire g172_p_spl_1;
  wire g172_p_spl_10;
  wire g172_p_spl_11;
  wire g191_n_spl_;
  wire g191_n_spl_0;
  wire g191_n_spl_00;
  wire g191_n_spl_01;
  wire g191_n_spl_1;
  wire g191_n_spl_10;
  wire g191_n_spl_11;
  wire g172_n_spl_;
  wire g172_n_spl_0;
  wire g172_n_spl_00;
  wire g172_n_spl_01;
  wire g172_n_spl_1;
  wire g172_n_spl_10;
  wire g172_n_spl_11;
  wire g191_p_spl_;
  wire g191_p_spl_0;
  wire g191_p_spl_00;
  wire g191_p_spl_01;
  wire g191_p_spl_1;
  wire g191_p_spl_10;
  wire g191_p_spl_11;
  wire g195_n_spl_;
  wire g198_n_spl_;
  wire g195_p_spl_;
  wire g198_p_spl_;
  wire g201_n_spl_;
  wire g202_p_spl_;
  wire g201_p_spl_;
  wire g202_n_spl_;
  wire g208_n_spl_;
  wire g211_n_spl_;
  wire g208_p_spl_;
  wire g211_p_spl_;
  wire g214_n_spl_;
  wire g214_n_spl_0;
  wire g214_n_spl_1;
  wire g214_p_spl_;
  wire g214_p_spl_0;
  wire g214_p_spl_1;
  wire g205_n_spl_;
  wire g217_p_spl_;
  wire g205_p_spl_;
  wire g217_n_spl_;
  wire g223_n_spl_;
  wire g226_n_spl_;
  wire g223_p_spl_;
  wire g226_p_spl_;
  wire g229_n_spl_;
  wire g230_p_spl_;
  wire g229_p_spl_;
  wire g230_n_spl_;
  wire g236_n_spl_;
  wire g239_n_spl_;
  wire g236_p_spl_;
  wire g239_p_spl_;
  wire g242_n_spl_;
  wire g242_n_spl_0;
  wire g242_n_spl_1;
  wire g242_p_spl_;
  wire g242_p_spl_0;
  wire g242_p_spl_1;
  wire g233_n_spl_;
  wire g245_p_spl_;
  wire g233_p_spl_;
  wire g245_n_spl_;
  wire g251_n_spl_;
  wire g254_n_spl_;
  wire g251_p_spl_;
  wire g254_p_spl_;
  wire g257_n_spl_;
  wire g258_p_spl_;
  wire g257_p_spl_;
  wire g258_n_spl_;
  wire g261_n_spl_;
  wire g264_p_spl_;
  wire g261_p_spl_;
  wire g264_n_spl_;
  wire g78_n_spl_;
  wire g78_n_spl_0;
  wire g78_n_spl_00;
  wire g78_n_spl_01;
  wire g78_n_spl_1;
  wire g78_n_spl_10;
  wire g267_p_spl_;
  wire g267_p_spl_0;
  wire g267_p_spl_00;
  wire g267_p_spl_01;
  wire g267_p_spl_1;
  wire g267_p_spl_10;
  wire g78_p_spl_;
  wire g78_p_spl_0;
  wire g78_p_spl_00;
  wire g78_p_spl_01;
  wire g78_p_spl_1;
  wire g78_p_spl_10;
  wire g267_n_spl_;
  wire g267_n_spl_0;
  wire g267_n_spl_00;
  wire g267_n_spl_01;
  wire g267_n_spl_1;
  wire g267_n_spl_10;
  wire g248_p_spl_;
  wire g248_p_spl_0;
  wire g248_p_spl_00;
  wire g248_p_spl_01;
  wire g248_p_spl_1;
  wire g248_p_spl_10;
  wire g248_p_spl_11;
  wire g268_p_spl_;
  wire g248_n_spl_;
  wire g248_n_spl_0;
  wire g248_n_spl_00;
  wire g248_n_spl_01;
  wire g248_n_spl_1;
  wire g248_n_spl_10;
  wire g248_n_spl_11;
  wire g268_n_spl_;
  wire g270_p_spl_;
  wire g270_n_spl_;
  wire g269_n_spl_;
  wire g271_n_spl_;
  wire g269_p_spl_;
  wire g271_p_spl_;
  wire g220_p_spl_;
  wire g220_p_spl_0;
  wire g220_p_spl_00;
  wire g220_p_spl_01;
  wire g220_p_spl_1;
  wire g220_p_spl_10;
  wire g220_p_spl_11;
  wire g220_n_spl_;
  wire g220_n_spl_0;
  wire g220_n_spl_00;
  wire g220_n_spl_01;
  wire g220_n_spl_1;
  wire g220_n_spl_10;
  wire g220_n_spl_11;
  wire g274_n_spl_;
  wire g274_n_spl_0;
  wire g274_p_spl_;
  wire g274_p_spl_0;
  wire g192_p_spl_;
  wire g279_n_spl_;
  wire g192_n_spl_;
  wire g279_p_spl_;
  wire g153_p_spl_;
  wire g280_p_spl_;
  wire g153_n_spl_;
  wire g280_n_spl_;
  wire g281_p_spl_;
  wire g281_p_spl_0;
  wire g281_p_spl_1;
  wire g281_n_spl_;
  wire g281_n_spl_0;
  wire g281_n_spl_1;
  wire g298_p_spl_;
  wire g299_p_spl_;
  wire g298_n_spl_;
  wire g299_n_spl_;
  wire g300_p_spl_;
  wire g300_p_spl_0;
  wire g300_p_spl_1;
  wire g300_n_spl_;
  wire g300_n_spl_0;
  wire g300_n_spl_1;
  wire g317_p_spl_;
  wire g317_n_spl_;
  wire g318_p_spl_;
  wire g318_p_spl_0;
  wire g318_p_spl_1;
  wire g318_n_spl_;
  wire g318_n_spl_0;
  wire g318_n_spl_1;
  wire g335_p_spl_;
  wire g335_n_spl_;
  wire g336_p_spl_;
  wire g336_p_spl_0;
  wire g336_p_spl_1;
  wire g336_n_spl_;
  wire g336_n_spl_0;
  wire g336_n_spl_1;
  wire g359_n_spl_;
  wire g359_n_spl_0;
  wire g359_p_spl_;
  wire g359_p_spl_0;
  wire g361_p_spl_;
  wire g361_p_spl_0;
  wire g361_p_spl_1;
  wire g361_n_spl_;
  wire g361_n_spl_0;
  wire g361_n_spl_1;
  wire g378_p_spl_;
  wire g378_n_spl_;
  wire g379_p_spl_;
  wire g379_p_spl_0;
  wire g379_p_spl_1;
  wire g379_n_spl_;
  wire g379_n_spl_0;
  wire g379_n_spl_1;
  wire g397_p_spl_;
  wire g397_p_spl_0;
  wire g397_p_spl_1;
  wire g397_n_spl_;
  wire g397_n_spl_0;
  wire g397_n_spl_1;
  wire g414_p_spl_;
  wire g414_p_spl_0;
  wire g414_p_spl_1;
  wire g414_n_spl_;
  wire g414_n_spl_0;
  wire g414_n_spl_1;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    G37_p,
    G37
  );


  not

  (
    G37_n,
    G37
  );


  buf

  (
    G38_p,
    G38
  );


  not

  (
    G38_n,
    G38
  );


  buf

  (
    G39_p,
    G39
  );


  not

  (
    G39_n,
    G39
  );


  buf

  (
    G40_p,
    G40
  );


  not

  (
    G40_n,
    G40
  );


  buf

  (
    G41_p,
    G41
  );


  not

  (
    G41_n,
    G41
  );


  and

  (
    g42_p,
    G9_n_spl_00,
    G13_n_spl_00
  );


  or

  (
    g42_n,
    G9_p_spl_00,
    G13_p_spl_00
  );


  and

  (
    g43_p,
    G9_p_spl_00,
    G13_p_spl_00
  );


  or

  (
    g43_n,
    G9_n_spl_00,
    G13_n_spl_00
  );


  and

  (
    g44_p,
    g42_n,
    g43_n
  );


  or

  (
    g44_n,
    g42_p,
    g43_p
  );


  and

  (
    g45_p,
    G1_p_spl_00,
    G5_n_spl_00
  );


  or

  (
    g45_n,
    G1_n_spl_00,
    G5_p_spl_00
  );


  and

  (
    g46_p,
    G1_n_spl_00,
    G5_p_spl_00
  );


  or

  (
    g46_n,
    G1_p_spl_00,
    G5_n_spl_00
  );


  and

  (
    g47_p,
    g45_n,
    g46_n
  );


  or

  (
    g47_n,
    g45_p,
    g46_p
  );


  and

  (
    g48_p,
    g44_n_spl_,
    g47_n_spl_
  );


  or

  (
    g48_n,
    g44_p_spl_,
    g47_p_spl_
  );


  and

  (
    g49_p,
    g44_p_spl_,
    g47_p_spl_
  );


  or

  (
    g49_n,
    g44_n_spl_,
    g47_n_spl_
  );


  and

  (
    g50_p,
    g48_n,
    g49_n
  );


  or

  (
    g50_n,
    g48_p,
    g49_p
  );


  and

  (
    g51_p,
    G33_p,
    G41_p_spl_00
  );


  or

  (
    g51_n,
    G33_n,
    G41_n_spl_00
  );


  and

  (
    g52_p,
    g50_n_spl_,
    g51_p_spl_
  );


  or

  (
    g52_n,
    g50_p_spl_,
    g51_n_spl_
  );


  and

  (
    g53_p,
    g50_p_spl_,
    g51_n_spl_
  );


  or

  (
    g53_n,
    g50_n_spl_,
    g51_p_spl_
  );


  and

  (
    g54_p,
    g52_n,
    g53_n
  );


  or

  (
    g54_n,
    g52_p,
    g53_p
  );


  and

  (
    g55_p,
    G19_n_spl_00,
    G20_n_spl_00
  );


  or

  (
    g55_n,
    G19_p_spl_00,
    G20_p_spl_00
  );


  and

  (
    g56_p,
    G19_p_spl_00,
    G20_p_spl_00
  );


  or

  (
    g56_n,
    G19_n_spl_00,
    G20_n_spl_00
  );


  and

  (
    g57_p,
    g55_n,
    g56_n
  );


  or

  (
    g57_n,
    g55_p,
    g56_p
  );


  and

  (
    g58_p,
    G17_p_spl_00,
    G18_n_spl_00
  );


  or

  (
    g58_n,
    G17_n_spl_00,
    G18_p_spl_00
  );


  and

  (
    g59_p,
    G17_n_spl_00,
    G18_p_spl_00
  );


  or

  (
    g59_n,
    G17_p_spl_00,
    G18_n_spl_00
  );


  and

  (
    g60_p,
    g58_n,
    g59_n
  );


  or

  (
    g60_n,
    g58_p,
    g59_p
  );


  and

  (
    g61_p,
    g57_n_spl_,
    g60_n_spl_
  );


  or

  (
    g61_n,
    g57_p_spl_,
    g60_p_spl_
  );


  and

  (
    g62_p,
    g57_p_spl_,
    g60_p_spl_
  );


  or

  (
    g62_n,
    g57_n_spl_,
    g60_n_spl_
  );


  and

  (
    g63_p,
    g61_n,
    g62_n
  );


  or

  (
    g63_n,
    g61_p,
    g62_p
  );


  and

  (
    g64_p,
    G23_n_spl_00,
    G24_n_spl_00
  );


  or

  (
    g64_n,
    G23_p_spl_00,
    G24_p_spl_00
  );


  and

  (
    g65_p,
    G23_p_spl_00,
    G24_p_spl_00
  );


  or

  (
    g65_n,
    G23_n_spl_00,
    G24_n_spl_00
  );


  and

  (
    g66_p,
    g64_n,
    g65_n
  );


  or

  (
    g66_n,
    g64_p,
    g65_p
  );


  and

  (
    g67_p,
    G21_p_spl_00,
    G22_n_spl_00
  );


  or

  (
    g67_n,
    G21_n_spl_00,
    G22_p_spl_00
  );


  and

  (
    g68_p,
    G21_n_spl_00,
    G22_p_spl_00
  );


  or

  (
    g68_n,
    G21_p_spl_00,
    G22_n_spl_00
  );


  and

  (
    g69_p,
    g67_n,
    g68_n
  );


  or

  (
    g69_n,
    g67_p,
    g68_p
  );


  and

  (
    g70_p,
    g66_n_spl_,
    g69_n_spl_
  );


  or

  (
    g70_n,
    g66_p_spl_,
    g69_p_spl_
  );


  and

  (
    g71_p,
    g66_p_spl_,
    g69_p_spl_
  );


  or

  (
    g71_n,
    g66_n_spl_,
    g69_n_spl_
  );


  and

  (
    g72_p,
    g70_n,
    g71_n
  );


  or

  (
    g72_n,
    g70_p,
    g71_p
  );


  and

  (
    g73_p,
    g63_n_spl_0,
    g72_n_spl_0
  );


  or

  (
    g73_n,
    g63_p_spl_0,
    g72_p_spl_0
  );


  and

  (
    g74_p,
    g63_p_spl_0,
    g72_p_spl_0
  );


  or

  (
    g74_n,
    g63_n_spl_0,
    g72_n_spl_0
  );


  and

  (
    g75_p,
    g73_n,
    g74_n
  );


  or

  (
    g75_n,
    g73_p,
    g74_p
  );


  and

  (
    g76_p,
    g54_n_spl_,
    g75_p_spl_
  );


  or

  (
    g76_n,
    g54_p_spl_,
    g75_n_spl_
  );


  and

  (
    g77_p,
    g54_p_spl_,
    g75_n_spl_
  );


  or

  (
    g77_n,
    g54_n_spl_,
    g75_p_spl_
  );


  and

  (
    g78_p,
    g76_n,
    g77_n
  );


  or

  (
    g78_n,
    g76_p,
    g77_p
  );


  and

  (
    g79_p,
    G25_n_spl_00,
    G29_n_spl_00
  );


  or

  (
    g79_n,
    G25_p_spl_00,
    G29_p_spl_00
  );


  and

  (
    g80_p,
    G25_p_spl_00,
    G29_p_spl_00
  );


  or

  (
    g80_n,
    G25_n_spl_00,
    G29_n_spl_00
  );


  and

  (
    g81_p,
    g79_n,
    g80_n
  );


  or

  (
    g81_n,
    g79_p,
    g80_p
  );


  and

  (
    g82_p,
    G17_p_spl_0,
    G21_n_spl_0
  );


  or

  (
    g82_n,
    G17_n_spl_0,
    G21_p_spl_0
  );


  and

  (
    g83_p,
    G17_n_spl_1,
    G21_p_spl_1
  );


  or

  (
    g83_n,
    G17_p_spl_1,
    G21_n_spl_1
  );


  and

  (
    g84_p,
    g82_n,
    g83_n
  );


  or

  (
    g84_n,
    g82_p,
    g83_p
  );


  and

  (
    g85_p,
    g81_n_spl_,
    g84_n_spl_
  );


  or

  (
    g85_n,
    g81_p_spl_,
    g84_p_spl_
  );


  and

  (
    g86_p,
    g81_p_spl_,
    g84_p_spl_
  );


  or

  (
    g86_n,
    g81_n_spl_,
    g84_n_spl_
  );


  and

  (
    g87_p,
    g85_n,
    g86_n
  );


  or

  (
    g87_n,
    g85_p,
    g86_p
  );


  and

  (
    g88_p,
    G37_p,
    G41_p_spl_00
  );


  or

  (
    g88_n,
    G37_n,
    G41_n_spl_00
  );


  and

  (
    g89_p,
    g87_n_spl_,
    g88_p_spl_
  );


  or

  (
    g89_n,
    g87_p_spl_,
    g88_n_spl_
  );


  and

  (
    g90_p,
    g87_p_spl_,
    g88_n_spl_
  );


  or

  (
    g90_n,
    g87_n_spl_,
    g88_p_spl_
  );


  and

  (
    g91_p,
    g89_n,
    g90_n
  );


  or

  (
    g91_n,
    g89_p,
    g90_p
  );


  and

  (
    g92_p,
    G7_n_spl_00,
    G8_n_spl_00
  );


  or

  (
    g92_n,
    G7_p_spl_00,
    G8_p_spl_00
  );


  and

  (
    g93_p,
    G7_p_spl_00,
    G8_p_spl_00
  );


  or

  (
    g93_n,
    G7_n_spl_00,
    G8_n_spl_00
  );


  and

  (
    g94_p,
    g92_n,
    g93_n
  );


  or

  (
    g94_n,
    g92_p,
    g93_p
  );


  and

  (
    g95_p,
    G5_p_spl_0,
    G6_n_spl_00
  );


  or

  (
    g95_n,
    G5_n_spl_0,
    G6_p_spl_00
  );


  and

  (
    g96_p,
    G5_n_spl_1,
    G6_p_spl_00
  );


  or

  (
    g96_n,
    G5_p_spl_1,
    G6_n_spl_00
  );


  and

  (
    g97_p,
    g95_n,
    g96_n
  );


  or

  (
    g97_n,
    g95_p,
    g96_p
  );


  and

  (
    g98_p,
    g94_n_spl_,
    g97_n_spl_
  );


  or

  (
    g98_n,
    g94_p_spl_,
    g97_p_spl_
  );


  and

  (
    g99_p,
    g94_p_spl_,
    g97_p_spl_
  );


  or

  (
    g99_n,
    g94_n_spl_,
    g97_n_spl_
  );


  and

  (
    g100_p,
    g98_n,
    g99_n
  );


  or

  (
    g100_n,
    g98_p,
    g99_p
  );


  and

  (
    g101_p,
    G3_n_spl_00,
    G4_n_spl_00
  );


  or

  (
    g101_n,
    G3_p_spl_00,
    G4_p_spl_00
  );


  and

  (
    g102_p,
    G3_p_spl_00,
    G4_p_spl_00
  );


  or

  (
    g102_n,
    G3_n_spl_00,
    G4_n_spl_00
  );


  and

  (
    g103_p,
    g101_n,
    g102_n
  );


  or

  (
    g103_n,
    g101_p,
    g102_p
  );


  and

  (
    g104_p,
    G1_p_spl_0,
    G2_n_spl_00
  );


  or

  (
    g104_n,
    G1_n_spl_0,
    G2_p_spl_00
  );


  and

  (
    g105_p,
    G1_n_spl_1,
    G2_p_spl_00
  );


  or

  (
    g105_n,
    G1_p_spl_1,
    G2_n_spl_00
  );


  and

  (
    g106_p,
    g104_n,
    g105_n
  );


  or

  (
    g106_n,
    g104_p,
    g105_p
  );


  and

  (
    g107_p,
    g103_n_spl_,
    g106_n_spl_
  );


  or

  (
    g107_n,
    g103_p_spl_,
    g106_p_spl_
  );


  and

  (
    g108_p,
    g103_p_spl_,
    g106_p_spl_
  );


  or

  (
    g108_n,
    g103_n_spl_,
    g106_n_spl_
  );


  and

  (
    g109_p,
    g107_n,
    g108_n
  );


  or

  (
    g109_n,
    g107_p,
    g108_p
  );


  and

  (
    g110_p,
    g100_n_spl_0,
    g109_n_spl_0
  );


  or

  (
    g110_n,
    g100_p_spl_0,
    g109_p_spl_0
  );


  and

  (
    g111_p,
    g100_p_spl_0,
    g109_p_spl_0
  );


  or

  (
    g111_n,
    g100_n_spl_0,
    g109_n_spl_0
  );


  and

  (
    g112_p,
    g110_n,
    g111_n
  );


  or

  (
    g112_n,
    g110_p,
    g111_p
  );


  and

  (
    g113_p,
    g91_n_spl_,
    g112_p_spl_
  );


  or

  (
    g113_n,
    g91_p_spl_,
    g112_n_spl_
  );


  and

  (
    g114_p,
    g91_p_spl_,
    g112_n_spl_
  );


  or

  (
    g114_n,
    g91_n_spl_,
    g112_p_spl_
  );


  and

  (
    g115_p,
    g113_n,
    g114_n
  );


  or

  (
    g115_n,
    g113_p,
    g114_p
  );


  and

  (
    g116_p,
    G26_n_spl_00,
    G30_n_spl_00
  );


  or

  (
    g116_n,
    G26_p_spl_00,
    G30_p_spl_00
  );


  and

  (
    g117_p,
    G26_p_spl_00,
    G30_p_spl_00
  );


  or

  (
    g117_n,
    G26_n_spl_00,
    G30_n_spl_00
  );


  and

  (
    g118_p,
    g116_n,
    g117_n
  );


  or

  (
    g118_n,
    g116_p,
    g117_p
  );


  and

  (
    g119_p,
    G18_p_spl_0,
    G22_n_spl_0
  );


  or

  (
    g119_n,
    G18_n_spl_0,
    G22_p_spl_0
  );


  and

  (
    g120_p,
    G18_n_spl_1,
    G22_p_spl_1
  );


  or

  (
    g120_n,
    G18_p_spl_1,
    G22_n_spl_1
  );


  and

  (
    g121_p,
    g119_n,
    g120_n
  );


  or

  (
    g121_n,
    g119_p,
    g120_p
  );


  and

  (
    g122_p,
    g118_n_spl_,
    g121_n_spl_
  );


  or

  (
    g122_n,
    g118_p_spl_,
    g121_p_spl_
  );


  and

  (
    g123_p,
    g118_p_spl_,
    g121_p_spl_
  );


  or

  (
    g123_n,
    g118_n_spl_,
    g121_n_spl_
  );


  and

  (
    g124_p,
    g122_n,
    g123_n
  );


  or

  (
    g124_n,
    g122_p,
    g123_p
  );


  and

  (
    g125_p,
    G38_p,
    G41_p_spl_01
  );


  or

  (
    g125_n,
    G38_n,
    G41_n_spl_01
  );


  and

  (
    g126_p,
    g124_n_spl_,
    g125_p_spl_
  );


  or

  (
    g126_n,
    g124_p_spl_,
    g125_n_spl_
  );


  and

  (
    g127_p,
    g124_p_spl_,
    g125_n_spl_
  );


  or

  (
    g127_n,
    g124_n_spl_,
    g125_p_spl_
  );


  and

  (
    g128_p,
    g126_n,
    g127_n
  );


  or

  (
    g128_n,
    g126_p,
    g127_p
  );


  and

  (
    g129_p,
    G15_n_spl_00,
    G16_n_spl_00
  );


  or

  (
    g129_n,
    G15_p_spl_00,
    G16_p_spl_00
  );


  and

  (
    g130_p,
    G15_p_spl_00,
    G16_p_spl_00
  );


  or

  (
    g130_n,
    G15_n_spl_00,
    G16_n_spl_00
  );


  and

  (
    g131_p,
    g129_n,
    g130_n
  );


  or

  (
    g131_n,
    g129_p,
    g130_p
  );


  and

  (
    g132_p,
    G13_p_spl_0,
    G14_n_spl_00
  );


  or

  (
    g132_n,
    G13_n_spl_0,
    G14_p_spl_00
  );


  and

  (
    g133_p,
    G13_n_spl_1,
    G14_p_spl_00
  );


  or

  (
    g133_n,
    G13_p_spl_1,
    G14_n_spl_00
  );


  and

  (
    g134_p,
    g132_n,
    g133_n
  );


  or

  (
    g134_n,
    g132_p,
    g133_p
  );


  and

  (
    g135_p,
    g131_n_spl_,
    g134_n_spl_
  );


  or

  (
    g135_n,
    g131_p_spl_,
    g134_p_spl_
  );


  and

  (
    g136_p,
    g131_p_spl_,
    g134_p_spl_
  );


  or

  (
    g136_n,
    g131_n_spl_,
    g134_n_spl_
  );


  and

  (
    g137_p,
    g135_n,
    g136_n
  );


  or

  (
    g137_n,
    g135_p,
    g136_p
  );


  and

  (
    g138_p,
    G11_n_spl_00,
    G12_n_spl_00
  );


  or

  (
    g138_n,
    G11_p_spl_00,
    G12_p_spl_00
  );


  and

  (
    g139_p,
    G11_p_spl_00,
    G12_p_spl_00
  );


  or

  (
    g139_n,
    G11_n_spl_00,
    G12_n_spl_00
  );


  and

  (
    g140_p,
    g138_n,
    g139_n
  );


  or

  (
    g140_n,
    g138_p,
    g139_p
  );


  and

  (
    g141_p,
    G9_p_spl_0,
    G10_n_spl_00
  );


  or

  (
    g141_n,
    G9_n_spl_0,
    G10_p_spl_00
  );


  and

  (
    g142_p,
    G9_n_spl_1,
    G10_p_spl_00
  );


  or

  (
    g142_n,
    G9_p_spl_1,
    G10_n_spl_00
  );


  and

  (
    g143_p,
    g141_n,
    g142_n
  );


  or

  (
    g143_n,
    g141_p,
    g142_p
  );


  and

  (
    g144_p,
    g140_n_spl_,
    g143_n_spl_
  );


  or

  (
    g144_n,
    g140_p_spl_,
    g143_p_spl_
  );


  and

  (
    g145_p,
    g140_p_spl_,
    g143_p_spl_
  );


  or

  (
    g145_n,
    g140_n_spl_,
    g143_n_spl_
  );


  and

  (
    g146_p,
    g144_n,
    g145_n
  );


  or

  (
    g146_n,
    g144_p,
    g145_p
  );


  and

  (
    g147_p,
    g137_n_spl_0,
    g146_n_spl_0
  );


  or

  (
    g147_n,
    g137_p_spl_0,
    g146_p_spl_0
  );


  and

  (
    g148_p,
    g137_p_spl_0,
    g146_p_spl_0
  );


  or

  (
    g148_n,
    g137_n_spl_0,
    g146_n_spl_0
  );


  and

  (
    g149_p,
    g147_n,
    g148_n
  );


  or

  (
    g149_n,
    g147_p,
    g148_p
  );


  and

  (
    g150_p,
    g128_n_spl_,
    g149_p_spl_
  );


  or

  (
    g150_n,
    g128_p_spl_,
    g149_n_spl_
  );


  and

  (
    g151_p,
    g128_p_spl_,
    g149_n_spl_
  );


  or

  (
    g151_n,
    g128_n_spl_,
    g149_p_spl_
  );


  and

  (
    g152_p,
    g150_n,
    g151_n
  );


  or

  (
    g152_n,
    g150_p,
    g151_p
  );


  and

  (
    g153_p,
    g115_n_spl_00,
    g152_p_spl_00
  );


  or

  (
    g153_n,
    g115_p_spl_00,
    g152_n_spl_00
  );


  and

  (
    g154_p,
    G28_n_spl_00,
    G32_n_spl_00
  );


  or

  (
    g154_n,
    G28_p_spl_00,
    G32_p_spl_00
  );


  and

  (
    g155_p,
    G28_p_spl_00,
    G32_p_spl_00
  );


  or

  (
    g155_n,
    G28_n_spl_00,
    G32_n_spl_00
  );


  and

  (
    g156_p,
    g154_n,
    g155_n
  );


  or

  (
    g156_n,
    g154_p,
    g155_p
  );


  and

  (
    g157_p,
    G20_p_spl_0,
    G24_n_spl_0
  );


  or

  (
    g157_n,
    G20_n_spl_0,
    G24_p_spl_0
  );


  and

  (
    g158_p,
    G20_n_spl_1,
    G24_p_spl_1
  );


  or

  (
    g158_n,
    G20_p_spl_1,
    G24_n_spl_1
  );


  and

  (
    g159_p,
    g157_n,
    g158_n
  );


  or

  (
    g159_n,
    g157_p,
    g158_p
  );


  and

  (
    g160_p,
    g156_n_spl_,
    g159_n_spl_
  );


  or

  (
    g160_n,
    g156_p_spl_,
    g159_p_spl_
  );


  and

  (
    g161_p,
    g156_p_spl_,
    g159_p_spl_
  );


  or

  (
    g161_n,
    g156_n_spl_,
    g159_n_spl_
  );


  and

  (
    g162_p,
    g160_n,
    g161_n
  );


  or

  (
    g162_n,
    g160_p,
    g161_p
  );


  and

  (
    g163_p,
    G40_p,
    G41_p_spl_01
  );


  or

  (
    g163_n,
    G40_n,
    G41_n_spl_01
  );


  and

  (
    g164_p,
    g162_n_spl_,
    g163_p_spl_
  );


  or

  (
    g164_n,
    g162_p_spl_,
    g163_n_spl_
  );


  and

  (
    g165_p,
    g162_p_spl_,
    g163_n_spl_
  );


  or

  (
    g165_n,
    g162_n_spl_,
    g163_p_spl_
  );


  and

  (
    g166_p,
    g164_n,
    g165_n
  );


  or

  (
    g166_n,
    g164_p,
    g165_p
  );


  and

  (
    g167_p,
    g100_n_spl_1,
    g137_n_spl_1
  );


  or

  (
    g167_n,
    g100_p_spl_1,
    g137_p_spl_1
  );


  and

  (
    g168_p,
    g100_p_spl_1,
    g137_p_spl_1
  );


  or

  (
    g168_n,
    g100_n_spl_1,
    g137_n_spl_1
  );


  and

  (
    g169_p,
    g167_n,
    g168_n
  );


  or

  (
    g169_n,
    g167_p,
    g168_p
  );


  and

  (
    g170_p,
    g166_n_spl_,
    g169_p_spl_
  );


  or

  (
    g170_n,
    g166_p_spl_,
    g169_n_spl_
  );


  and

  (
    g171_p,
    g166_p_spl_,
    g169_n_spl_
  );


  or

  (
    g171_n,
    g166_n_spl_,
    g169_p_spl_
  );


  and

  (
    g172_p,
    g170_n,
    g171_n
  );


  or

  (
    g172_n,
    g170_p,
    g171_p
  );


  and

  (
    g173_p,
    G27_n_spl_00,
    G31_n_spl_00
  );


  or

  (
    g173_n,
    G27_p_spl_00,
    G31_p_spl_00
  );


  and

  (
    g174_p,
    G27_p_spl_00,
    G31_p_spl_00
  );


  or

  (
    g174_n,
    G27_n_spl_00,
    G31_n_spl_00
  );


  and

  (
    g175_p,
    g173_n,
    g174_n
  );


  or

  (
    g175_n,
    g173_p,
    g174_p
  );


  and

  (
    g176_p,
    G19_p_spl_0,
    G23_n_spl_0
  );


  or

  (
    g176_n,
    G19_n_spl_0,
    G23_p_spl_0
  );


  and

  (
    g177_p,
    G19_n_spl_1,
    G23_p_spl_1
  );


  or

  (
    g177_n,
    G19_p_spl_1,
    G23_n_spl_1
  );


  and

  (
    g178_p,
    g176_n,
    g177_n
  );


  or

  (
    g178_n,
    g176_p,
    g177_p
  );


  and

  (
    g179_p,
    g175_n_spl_,
    g178_n_spl_
  );


  or

  (
    g179_n,
    g175_p_spl_,
    g178_p_spl_
  );


  and

  (
    g180_p,
    g175_p_spl_,
    g178_p_spl_
  );


  or

  (
    g180_n,
    g175_n_spl_,
    g178_n_spl_
  );


  and

  (
    g181_p,
    g179_n,
    g180_n
  );


  or

  (
    g181_n,
    g179_p,
    g180_p
  );


  and

  (
    g182_p,
    G39_p,
    G41_p_spl_10
  );


  or

  (
    g182_n,
    G39_n,
    G41_n_spl_10
  );


  and

  (
    g183_p,
    g181_n_spl_,
    g182_p_spl_
  );


  or

  (
    g183_n,
    g181_p_spl_,
    g182_n_spl_
  );


  and

  (
    g184_p,
    g181_p_spl_,
    g182_n_spl_
  );


  or

  (
    g184_n,
    g181_n_spl_,
    g182_p_spl_
  );


  and

  (
    g185_p,
    g183_n,
    g184_n
  );


  or

  (
    g185_n,
    g183_p,
    g184_p
  );


  and

  (
    g186_p,
    g109_n_spl_1,
    g146_n_spl_1
  );


  or

  (
    g186_n,
    g109_p_spl_1,
    g146_p_spl_1
  );


  and

  (
    g187_p,
    g109_p_spl_1,
    g146_p_spl_1
  );


  or

  (
    g187_n,
    g109_n_spl_1,
    g146_n_spl_1
  );


  and

  (
    g188_p,
    g186_n,
    g187_n
  );


  or

  (
    g188_n,
    g186_p,
    g187_p
  );


  and

  (
    g189_p,
    g185_n_spl_,
    g188_p_spl_
  );


  or

  (
    g189_n,
    g185_p_spl_,
    g188_n_spl_
  );


  and

  (
    g190_p,
    g185_p_spl_,
    g188_n_spl_
  );


  or

  (
    g190_n,
    g185_n_spl_,
    g188_p_spl_
  );


  and

  (
    g191_p,
    g189_n,
    g190_n
  );


  or

  (
    g191_n,
    g189_p,
    g190_p
  );


  and

  (
    g192_p,
    g172_p_spl_00,
    g191_n_spl_00
  );


  or

  (
    g192_n,
    g172_n_spl_00,
    g191_p_spl_00
  );


  and

  (
    g193_p,
    G12_n_spl_0,
    G16_n_spl_0
  );


  or

  (
    g193_n,
    G12_p_spl_0,
    G16_p_spl_0
  );


  and

  (
    g194_p,
    G12_p_spl_1,
    G16_p_spl_1
  );


  or

  (
    g194_n,
    G12_n_spl_1,
    G16_n_spl_1
  );


  and

  (
    g195_p,
    g193_n,
    g194_n
  );


  or

  (
    g195_n,
    g193_p,
    g194_p
  );


  and

  (
    g196_p,
    G4_p_spl_0,
    G8_n_spl_0
  );


  or

  (
    g196_n,
    G4_n_spl_0,
    G8_p_spl_0
  );


  and

  (
    g197_p,
    G4_n_spl_1,
    G8_p_spl_1
  );


  or

  (
    g197_n,
    G4_p_spl_1,
    G8_n_spl_1
  );


  and

  (
    g198_p,
    g196_n,
    g197_n
  );


  or

  (
    g198_n,
    g196_p,
    g197_p
  );


  and

  (
    g199_p,
    g195_n_spl_,
    g198_n_spl_
  );


  or

  (
    g199_n,
    g195_p_spl_,
    g198_p_spl_
  );


  and

  (
    g200_p,
    g195_p_spl_,
    g198_p_spl_
  );


  or

  (
    g200_n,
    g195_n_spl_,
    g198_n_spl_
  );


  and

  (
    g201_p,
    g199_n,
    g200_n
  );


  or

  (
    g201_n,
    g199_p,
    g200_p
  );


  and

  (
    g202_p,
    G36_p,
    G41_p_spl_10
  );


  or

  (
    g202_n,
    G36_n,
    G41_n_spl_10
  );


  and

  (
    g203_p,
    g201_n_spl_,
    g202_p_spl_
  );


  or

  (
    g203_n,
    g201_p_spl_,
    g202_n_spl_
  );


  and

  (
    g204_p,
    g201_p_spl_,
    g202_n_spl_
  );


  or

  (
    g204_n,
    g201_n_spl_,
    g202_p_spl_
  );


  and

  (
    g205_p,
    g203_n,
    g204_n
  );


  or

  (
    g205_n,
    g203_p,
    g204_p
  );


  and

  (
    g206_p,
    G31_n_spl_0,
    G32_n_spl_0
  );


  or

  (
    g206_n,
    G31_p_spl_0,
    G32_p_spl_0
  );


  and

  (
    g207_p,
    G31_p_spl_1,
    G32_p_spl_1
  );


  or

  (
    g207_n,
    G31_n_spl_1,
    G32_n_spl_1
  );


  and

  (
    g208_p,
    g206_n,
    g207_n
  );


  or

  (
    g208_n,
    g206_p,
    g207_p
  );


  and

  (
    g209_p,
    G29_p_spl_0,
    G30_n_spl_0
  );


  or

  (
    g209_n,
    G29_n_spl_0,
    G30_p_spl_0
  );


  and

  (
    g210_p,
    G29_n_spl_1,
    G30_p_spl_1
  );


  or

  (
    g210_n,
    G29_p_spl_1,
    G30_n_spl_1
  );


  and

  (
    g211_p,
    g209_n,
    g210_n
  );


  or

  (
    g211_n,
    g209_p,
    g210_p
  );


  and

  (
    g212_p,
    g208_n_spl_,
    g211_n_spl_
  );


  or

  (
    g212_n,
    g208_p_spl_,
    g211_p_spl_
  );


  and

  (
    g213_p,
    g208_p_spl_,
    g211_p_spl_
  );


  or

  (
    g213_n,
    g208_n_spl_,
    g211_n_spl_
  );


  and

  (
    g214_p,
    g212_n,
    g213_n
  );


  or

  (
    g214_n,
    g212_p,
    g213_p
  );


  and

  (
    g215_p,
    g72_n_spl_1,
    g214_n_spl_0
  );


  or

  (
    g215_n,
    g72_p_spl_1,
    g214_p_spl_0
  );


  and

  (
    g216_p,
    g72_p_spl_1,
    g214_p_spl_0
  );


  or

  (
    g216_n,
    g72_n_spl_1,
    g214_n_spl_0
  );


  and

  (
    g217_p,
    g215_n,
    g216_n
  );


  or

  (
    g217_n,
    g215_p,
    g216_p
  );


  and

  (
    g218_p,
    g205_n_spl_,
    g217_p_spl_
  );


  or

  (
    g218_n,
    g205_p_spl_,
    g217_n_spl_
  );


  and

  (
    g219_p,
    g205_p_spl_,
    g217_n_spl_
  );


  or

  (
    g219_n,
    g205_n_spl_,
    g217_p_spl_
  );


  and

  (
    g220_p,
    g218_n,
    g219_n
  );


  or

  (
    g220_n,
    g218_p,
    g219_p
  );


  and

  (
    g221_p,
    G11_n_spl_0,
    G15_n_spl_0
  );


  or

  (
    g221_n,
    G11_p_spl_0,
    G15_p_spl_0
  );


  and

  (
    g222_p,
    G11_p_spl_1,
    G15_p_spl_1
  );


  or

  (
    g222_n,
    G11_n_spl_1,
    G15_n_spl_1
  );


  and

  (
    g223_p,
    g221_n,
    g222_n
  );


  or

  (
    g223_n,
    g221_p,
    g222_p
  );


  and

  (
    g224_p,
    G3_p_spl_0,
    G7_n_spl_0
  );


  or

  (
    g224_n,
    G3_n_spl_0,
    G7_p_spl_0
  );


  and

  (
    g225_p,
    G3_n_spl_1,
    G7_p_spl_1
  );


  or

  (
    g225_n,
    G3_p_spl_1,
    G7_n_spl_1
  );


  and

  (
    g226_p,
    g224_n,
    g225_n
  );


  or

  (
    g226_n,
    g224_p,
    g225_p
  );


  and

  (
    g227_p,
    g223_n_spl_,
    g226_n_spl_
  );


  or

  (
    g227_n,
    g223_p_spl_,
    g226_p_spl_
  );


  and

  (
    g228_p,
    g223_p_spl_,
    g226_p_spl_
  );


  or

  (
    g228_n,
    g223_n_spl_,
    g226_n_spl_
  );


  and

  (
    g229_p,
    g227_n,
    g228_n
  );


  or

  (
    g229_n,
    g227_p,
    g228_p
  );


  and

  (
    g230_p,
    G35_p,
    G41_p_spl_11
  );


  or

  (
    g230_n,
    G35_n,
    G41_n_spl_11
  );


  and

  (
    g231_p,
    g229_n_spl_,
    g230_p_spl_
  );


  or

  (
    g231_n,
    g229_p_spl_,
    g230_n_spl_
  );


  and

  (
    g232_p,
    g229_p_spl_,
    g230_n_spl_
  );


  or

  (
    g232_n,
    g229_n_spl_,
    g230_p_spl_
  );


  and

  (
    g233_p,
    g231_n,
    g232_n
  );


  or

  (
    g233_n,
    g231_p,
    g232_p
  );


  and

  (
    g234_p,
    G27_n_spl_0,
    G28_n_spl_0
  );


  or

  (
    g234_n,
    G27_p_spl_0,
    G28_p_spl_0
  );


  and

  (
    g235_p,
    G27_p_spl_1,
    G28_p_spl_1
  );


  or

  (
    g235_n,
    G27_n_spl_1,
    G28_n_spl_1
  );


  and

  (
    g236_p,
    g234_n,
    g235_n
  );


  or

  (
    g236_n,
    g234_p,
    g235_p
  );


  and

  (
    g237_p,
    G25_p_spl_0,
    G26_n_spl_0
  );


  or

  (
    g237_n,
    G25_n_spl_0,
    G26_p_spl_0
  );


  and

  (
    g238_p,
    G25_n_spl_1,
    G26_p_spl_1
  );


  or

  (
    g238_n,
    G25_p_spl_1,
    G26_n_spl_1
  );


  and

  (
    g239_p,
    g237_n,
    g238_n
  );


  or

  (
    g239_n,
    g237_p,
    g238_p
  );


  and

  (
    g240_p,
    g236_n_spl_,
    g239_n_spl_
  );


  or

  (
    g240_n,
    g236_p_spl_,
    g239_p_spl_
  );


  and

  (
    g241_p,
    g236_p_spl_,
    g239_p_spl_
  );


  or

  (
    g241_n,
    g236_n_spl_,
    g239_n_spl_
  );


  and

  (
    g242_p,
    g240_n,
    g241_n
  );


  or

  (
    g242_n,
    g240_p,
    g241_p
  );


  and

  (
    g243_p,
    g63_n_spl_1,
    g242_n_spl_0
  );


  or

  (
    g243_n,
    g63_p_spl_1,
    g242_p_spl_0
  );


  and

  (
    g244_p,
    g63_p_spl_1,
    g242_p_spl_0
  );


  or

  (
    g244_n,
    g63_n_spl_1,
    g242_n_spl_0
  );


  and

  (
    g245_p,
    g243_n,
    g244_n
  );


  or

  (
    g245_n,
    g243_p,
    g244_p
  );


  and

  (
    g246_p,
    g233_n_spl_,
    g245_p_spl_
  );


  or

  (
    g246_n,
    g233_p_spl_,
    g245_n_spl_
  );


  and

  (
    g247_p,
    g233_p_spl_,
    g245_n_spl_
  );


  or

  (
    g247_n,
    g233_n_spl_,
    g245_p_spl_
  );


  and

  (
    g248_p,
    g246_n,
    g247_n
  );


  or

  (
    g248_n,
    g246_p,
    g247_p
  );


  and

  (
    g249_p,
    G10_n_spl_0,
    G14_n_spl_0
  );


  or

  (
    g249_n,
    G10_p_spl_0,
    G14_p_spl_0
  );


  and

  (
    g250_p,
    G10_p_spl_1,
    G14_p_spl_1
  );


  or

  (
    g250_n,
    G10_n_spl_1,
    G14_n_spl_1
  );


  and

  (
    g251_p,
    g249_n,
    g250_n
  );


  or

  (
    g251_n,
    g249_p,
    g250_p
  );


  and

  (
    g252_p,
    G2_p_spl_0,
    G6_n_spl_0
  );


  or

  (
    g252_n,
    G2_n_spl_0,
    G6_p_spl_0
  );


  and

  (
    g253_p,
    G2_n_spl_1,
    G6_p_spl_1
  );


  or

  (
    g253_n,
    G2_p_spl_1,
    G6_n_spl_1
  );


  and

  (
    g254_p,
    g252_n,
    g253_n
  );


  or

  (
    g254_n,
    g252_p,
    g253_p
  );


  and

  (
    g255_p,
    g251_n_spl_,
    g254_n_spl_
  );


  or

  (
    g255_n,
    g251_p_spl_,
    g254_p_spl_
  );


  and

  (
    g256_p,
    g251_p_spl_,
    g254_p_spl_
  );


  or

  (
    g256_n,
    g251_n_spl_,
    g254_n_spl_
  );


  and

  (
    g257_p,
    g255_n,
    g256_n
  );


  or

  (
    g257_n,
    g255_p,
    g256_p
  );


  and

  (
    g258_p,
    G34_p,
    G41_p_spl_11
  );


  or

  (
    g258_n,
    G34_n,
    G41_n_spl_11
  );


  and

  (
    g259_p,
    g257_n_spl_,
    g258_p_spl_
  );


  or

  (
    g259_n,
    g257_p_spl_,
    g258_n_spl_
  );


  and

  (
    g260_p,
    g257_p_spl_,
    g258_n_spl_
  );


  or

  (
    g260_n,
    g257_n_spl_,
    g258_p_spl_
  );


  and

  (
    g261_p,
    g259_n,
    g260_n
  );


  or

  (
    g261_n,
    g259_p,
    g260_p
  );


  and

  (
    g262_p,
    g214_n_spl_1,
    g242_n_spl_1
  );


  or

  (
    g262_n,
    g214_p_spl_1,
    g242_p_spl_1
  );


  and

  (
    g263_p,
    g214_p_spl_1,
    g242_p_spl_1
  );


  or

  (
    g263_n,
    g214_n_spl_1,
    g242_n_spl_1
  );


  and

  (
    g264_p,
    g262_n,
    g263_n
  );


  or

  (
    g264_n,
    g262_p,
    g263_p
  );


  and

  (
    g265_p,
    g261_n_spl_,
    g264_p_spl_
  );


  or

  (
    g265_n,
    g261_p_spl_,
    g264_n_spl_
  );


  and

  (
    g266_p,
    g261_p_spl_,
    g264_n_spl_
  );


  or

  (
    g266_n,
    g261_n_spl_,
    g264_p_spl_
  );


  and

  (
    g267_p,
    g265_n,
    g266_n
  );


  or

  (
    g267_n,
    g265_p,
    g266_p
  );


  and

  (
    g268_p,
    g78_n_spl_00,
    g267_p_spl_00
  );


  or

  (
    g268_n,
    g78_p_spl_00,
    g267_n_spl_00
  );


  and

  (
    g269_p,
    g248_p_spl_00,
    g268_p_spl_
  );


  or

  (
    g269_n,
    g248_n_spl_00,
    g268_n_spl_
  );


  and

  (
    g270_p,
    g78_p_spl_00,
    g267_n_spl_00
  );


  or

  (
    g270_n,
    g78_n_spl_00,
    g267_p_spl_00
  );


  and

  (
    g271_p,
    g248_p_spl_00,
    g270_p_spl_
  );


  or

  (
    g271_n,
    g248_n_spl_00,
    g270_n_spl_
  );


  and

  (
    g272_p,
    g269_n_spl_,
    g271_n_spl_
  );


  or

  (
    g272_n,
    g269_p_spl_,
    g271_p_spl_
  );


  and

  (
    g273_p,
    g220_p_spl_00,
    g272_n
  );


  or

  (
    g273_n,
    g220_n_spl_00,
    g272_p
  );


  and

  (
    g274_p,
    g220_p_spl_00,
    g248_n_spl_01
  );


  or

  (
    g274_n,
    g220_n_spl_00,
    g248_p_spl_01
  );


  and

  (
    g275_p,
    g220_n_spl_01,
    g248_p_spl_01
  );


  or

  (
    g275_n,
    g220_p_spl_01,
    g248_n_spl_01
  );


  and

  (
    g276_p,
    g274_n_spl_0,
    g275_n
  );


  or

  (
    g276_n,
    g274_p_spl_0,
    g275_p
  );


  and

  (
    g277_p,
    g267_p_spl_01,
    g276_n
  );


  or

  (
    g277_n,
    g267_n_spl_01,
    g276_p
  );


  and

  (
    g278_p,
    g78_p_spl_01,
    g277_p
  );


  or

  (
    g278_n,
    g78_n_spl_01,
    g277_n
  );


  and

  (
    g279_p,
    g273_n,
    g278_n
  );


  or

  (
    g279_n,
    g273_p,
    g278_p
  );


  and

  (
    g280_p,
    g192_p_spl_,
    g279_n_spl_
  );


  or

  (
    g280_n,
    g192_n_spl_,
    g279_p_spl_
  );


  and

  (
    g281_p,
    g153_p_spl_,
    g280_p_spl_
  );


  or

  (
    g281_n,
    g153_n_spl_,
    g280_n_spl_
  );


  and

  (
    g282_p,
    g78_n_spl_01,
    g281_p_spl_0
  );


  or

  (
    g282_n,
    g78_p_spl_01,
    g281_n_spl_0
  );


  and

  (
    g283_p,
    G1_p_spl_1,
    g282_n
  );


  and

  (
    g284_p,
    G1_n_spl_1,
    g282_p
  );


  or

  (
    g285_n,
    g283_p,
    g284_p
  );


  and

  (
    g286_p,
    g267_n_spl_01,
    g281_p_spl_0
  );


  or

  (
    g286_n,
    g267_p_spl_01,
    g281_n_spl_0
  );


  and

  (
    g287_p,
    G2_p_spl_1,
    g286_n
  );


  and

  (
    g288_p,
    G2_n_spl_1,
    g286_p
  );


  or

  (
    g289_n,
    g287_p,
    g288_p
  );


  and

  (
    g290_p,
    g248_n_spl_10,
    g281_p_spl_1
  );


  or

  (
    g290_n,
    g248_p_spl_10,
    g281_n_spl_1
  );


  and

  (
    g291_p,
    G3_p_spl_1,
    g290_n
  );


  and

  (
    g292_p,
    G3_n_spl_1,
    g290_p
  );


  or

  (
    g293_n,
    g291_p,
    g292_p
  );


  and

  (
    g294_p,
    g220_n_spl_01,
    g281_p_spl_1
  );


  or

  (
    g294_n,
    g220_p_spl_01,
    g281_n_spl_1
  );


  and

  (
    g295_p,
    G4_p_spl_1,
    g294_n
  );


  and

  (
    g296_p,
    G4_n_spl_1,
    g294_p
  );


  or

  (
    g297_n,
    g295_p,
    g296_p
  );


  and

  (
    g298_p,
    g153_p_spl_,
    g191_p_spl_00
  );


  or

  (
    g298_n,
    g153_n_spl_,
    g191_n_spl_00
  );


  and

  (
    g299_p,
    g172_n_spl_00,
    g279_n_spl_
  );


  or

  (
    g299_n,
    g172_p_spl_00,
    g279_p_spl_
  );


  and

  (
    g300_p,
    g298_p_spl_,
    g299_p_spl_
  );


  or

  (
    g300_n,
    g298_n_spl_,
    g299_n_spl_
  );


  and

  (
    g301_p,
    g78_n_spl_10,
    g300_p_spl_0
  );


  or

  (
    g301_n,
    g78_p_spl_10,
    g300_n_spl_0
  );


  and

  (
    g302_p,
    G5_p_spl_1,
    g301_n
  );


  and

  (
    g303_p,
    G5_n_spl_1,
    g301_p
  );


  or

  (
    g304_n,
    g302_p,
    g303_p
  );


  and

  (
    g305_p,
    g267_n_spl_10,
    g300_p_spl_0
  );


  or

  (
    g305_n,
    g267_p_spl_10,
    g300_n_spl_0
  );


  and

  (
    g306_p,
    G6_p_spl_1,
    g305_n
  );


  and

  (
    g307_p,
    G6_n_spl_1,
    g305_p
  );


  or

  (
    g308_n,
    g306_p,
    g307_p
  );


  and

  (
    g309_p,
    g248_n_spl_10,
    g300_p_spl_1
  );


  or

  (
    g309_n,
    g248_p_spl_10,
    g300_n_spl_1
  );


  and

  (
    g310_p,
    G7_p_spl_1,
    g309_n
  );


  and

  (
    g311_p,
    G7_n_spl_1,
    g309_p
  );


  or

  (
    g312_n,
    g310_p,
    g311_p
  );


  and

  (
    g313_p,
    g220_n_spl_10,
    g300_p_spl_1
  );


  or

  (
    g313_n,
    g220_p_spl_10,
    g300_n_spl_1
  );


  and

  (
    g314_p,
    G8_p_spl_1,
    g313_n
  );


  and

  (
    g315_p,
    G8_n_spl_1,
    g313_p
  );


  or

  (
    g316_n,
    g314_p,
    g315_p
  );


  and

  (
    g317_p,
    g115_p_spl_00,
    g152_n_spl_00
  );


  or

  (
    g317_n,
    g115_n_spl_00,
    g152_p_spl_00
  );


  and

  (
    g318_p,
    g280_p_spl_,
    g317_p_spl_
  );


  or

  (
    g318_n,
    g280_n_spl_,
    g317_n_spl_
  );


  and

  (
    g319_p,
    g78_n_spl_10,
    g318_p_spl_0
  );


  or

  (
    g319_n,
    g78_p_spl_10,
    g318_n_spl_0
  );


  and

  (
    g320_p,
    G9_p_spl_1,
    g319_n
  );


  and

  (
    g321_p,
    G9_n_spl_1,
    g319_p
  );


  or

  (
    g322_n,
    g320_p,
    g321_p
  );


  and

  (
    g323_p,
    g267_n_spl_10,
    g318_p_spl_0
  );


  or

  (
    g323_n,
    g267_p_spl_10,
    g318_n_spl_0
  );


  and

  (
    g324_p,
    G10_p_spl_1,
    g323_n
  );


  and

  (
    g325_p,
    G10_n_spl_1,
    g323_p
  );


  or

  (
    g326_n,
    g324_p,
    g325_p
  );


  and

  (
    g327_p,
    g248_n_spl_11,
    g318_p_spl_1
  );


  or

  (
    g327_n,
    g248_p_spl_11,
    g318_n_spl_1
  );


  and

  (
    g328_p,
    G11_p_spl_1,
    g327_n
  );


  and

  (
    g329_p,
    G11_n_spl_1,
    g327_p
  );


  or

  (
    g330_n,
    g328_p,
    g329_p
  );


  and

  (
    g331_p,
    g220_n_spl_10,
    g318_p_spl_1
  );


  or

  (
    g331_n,
    g220_p_spl_10,
    g318_n_spl_1
  );


  and

  (
    g332_p,
    G12_p_spl_1,
    g331_n
  );


  and

  (
    g333_p,
    G12_n_spl_1,
    g331_p
  );


  or

  (
    g334_n,
    g332_p,
    g333_p
  );


  and

  (
    g335_p,
    g191_p_spl_01,
    g317_p_spl_
  );


  or

  (
    g335_n,
    g191_n_spl_01,
    g317_n_spl_
  );


  and

  (
    g336_p,
    g299_p_spl_,
    g335_p_spl_
  );


  or

  (
    g336_n,
    g299_n_spl_,
    g335_n_spl_
  );


  and

  (
    g337_p,
    g78_n_spl_1,
    g336_p_spl_0
  );


  or

  (
    g337_n,
    g78_p_spl_1,
    g336_n_spl_0
  );


  and

  (
    g338_p,
    G13_p_spl_1,
    g337_n
  );


  and

  (
    g339_p,
    G13_n_spl_1,
    g337_p
  );


  or

  (
    g340_n,
    g338_p,
    g339_p
  );


  and

  (
    g341_p,
    g267_n_spl_1,
    g336_p_spl_0
  );


  or

  (
    g341_n,
    g267_p_spl_1,
    g336_n_spl_0
  );


  and

  (
    g342_p,
    G14_p_spl_1,
    g341_n
  );


  and

  (
    g343_p,
    G14_n_spl_1,
    g341_p
  );


  or

  (
    g344_n,
    g342_p,
    g343_p
  );


  and

  (
    g345_p,
    g248_n_spl_11,
    g336_p_spl_1
  );


  or

  (
    g345_n,
    g248_p_spl_11,
    g336_n_spl_1
  );


  and

  (
    g346_p,
    G15_p_spl_1,
    g345_n
  );


  and

  (
    g347_p,
    G15_n_spl_1,
    g345_p
  );


  or

  (
    g348_n,
    g346_p,
    g347_p
  );


  and

  (
    g349_p,
    g220_n_spl_11,
    g336_p_spl_1
  );


  or

  (
    g349_n,
    g220_p_spl_11,
    g336_n_spl_1
  );


  and

  (
    g350_p,
    G16_p_spl_1,
    g349_n
  );


  and

  (
    g351_p,
    G16_n_spl_1,
    g349_p
  );


  or

  (
    g352_n,
    g350_p,
    g351_p
  );


  and

  (
    g353_p,
    g298_n_spl_,
    g335_n_spl_
  );


  or

  (
    g353_n,
    g298_p_spl_,
    g335_p_spl_
  );


  and

  (
    g354_p,
    g172_p_spl_01,
    g353_n
  );


  or

  (
    g354_n,
    g172_n_spl_01,
    g353_p
  );


  and

  (
    g355_p,
    g172_n_spl_01,
    g191_p_spl_01
  );


  or

  (
    g355_n,
    g172_p_spl_01,
    g191_n_spl_01
  );


  and

  (
    g356_p,
    g192_n_spl_,
    g355_n
  );


  or

  (
    g356_n,
    g192_p_spl_,
    g355_p
  );


  and

  (
    g357_p,
    g152_p_spl_01,
    g356_n
  );


  or

  (
    g357_n,
    g152_n_spl_01,
    g356_p
  );


  and

  (
    g358_p,
    g115_p_spl_01,
    g357_p
  );


  or

  (
    g358_n,
    g115_n_spl_01,
    g357_n
  );


  and

  (
    g359_p,
    g354_n,
    g358_n
  );


  or

  (
    g359_n,
    g354_p,
    g358_p
  );


  and

  (
    g360_p,
    g268_p_spl_,
    g359_n_spl_0
  );


  or

  (
    g360_n,
    g268_n_spl_,
    g359_p_spl_0
  );


  and

  (
    g361_p,
    g274_p_spl_0,
    g360_p
  );


  or

  (
    g361_n,
    g274_n_spl_0,
    g360_n
  );


  and

  (
    g362_p,
    g115_n_spl_01,
    g361_p_spl_0
  );


  or

  (
    g362_n,
    g115_p_spl_01,
    g361_n_spl_0
  );


  and

  (
    g363_p,
    G17_p_spl_1,
    g362_n
  );


  and

  (
    g364_p,
    G17_n_spl_1,
    g362_p
  );


  or

  (
    g365_n,
    g363_p,
    g364_p
  );


  and

  (
    g366_p,
    g152_n_spl_01,
    g361_p_spl_0
  );


  or

  (
    g366_n,
    g152_p_spl_01,
    g361_n_spl_0
  );


  and

  (
    g367_p,
    G18_p_spl_1,
    g366_n
  );


  and

  (
    g368_p,
    G18_n_spl_1,
    g366_p
  );


  or

  (
    g369_n,
    g367_p,
    g368_p
  );


  and

  (
    g370_p,
    g191_n_spl_10,
    g361_p_spl_1
  );


  or

  (
    g370_n,
    g191_p_spl_10,
    g361_n_spl_1
  );


  and

  (
    g371_p,
    G19_p_spl_1,
    g370_n
  );


  and

  (
    g372_p,
    G19_n_spl_1,
    g370_p
  );


  or

  (
    g373_n,
    g371_p,
    g372_p
  );


  and

  (
    g374_p,
    g172_n_spl_10,
    g361_p_spl_1
  );


  or

  (
    g374_n,
    g172_p_spl_10,
    g361_n_spl_1
  );


  and

  (
    g375_p,
    G20_p_spl_1,
    g374_n
  );


  and

  (
    g376_p,
    G20_n_spl_1,
    g374_p
  );


  or

  (
    g377_n,
    g375_p,
    g376_p
  );


  and

  (
    g378_p,
    g220_n_spl_11,
    g359_n_spl_0
  );


  or

  (
    g378_n,
    g220_p_spl_11,
    g359_p_spl_0
  );


  and

  (
    g379_p,
    g269_p_spl_,
    g378_p_spl_
  );


  or

  (
    g379_n,
    g269_n_spl_,
    g378_n_spl_
  );


  and

  (
    g380_p,
    g115_n_spl_10,
    g379_p_spl_0
  );


  or

  (
    g380_n,
    g115_p_spl_10,
    g379_n_spl_0
  );


  and

  (
    g381_p,
    G21_p_spl_1,
    g380_n
  );


  and

  (
    g382_p,
    G21_n_spl_1,
    g380_p
  );


  or

  (
    g383_n,
    g381_p,
    g382_p
  );


  and

  (
    g384_p,
    g152_n_spl_10,
    g379_p_spl_0
  );


  or

  (
    g384_n,
    g152_p_spl_10,
    g379_n_spl_0
  );


  and

  (
    g385_p,
    G22_p_spl_1,
    g384_n
  );


  and

  (
    g386_p,
    G22_n_spl_1,
    g384_p
  );


  or

  (
    g387_n,
    g385_p,
    g386_p
  );


  and

  (
    g388_p,
    g191_n_spl_10,
    g379_p_spl_1
  );


  or

  (
    g388_n,
    g191_p_spl_10,
    g379_n_spl_1
  );


  and

  (
    g389_p,
    G23_p_spl_1,
    g388_n
  );


  and

  (
    g390_p,
    G23_n_spl_1,
    g388_p
  );


  or

  (
    g391_n,
    g389_p,
    g390_p
  );


  and

  (
    g392_p,
    g172_n_spl_10,
    g379_p_spl_1
  );


  or

  (
    g392_n,
    g172_p_spl_10,
    g379_n_spl_1
  );


  and

  (
    g393_p,
    G24_p_spl_1,
    g392_n
  );


  and

  (
    g394_p,
    G24_n_spl_1,
    g392_p
  );


  or

  (
    g395_n,
    g393_p,
    g394_p
  );


  and

  (
    g396_p,
    g270_p_spl_,
    g359_n_spl_
  );


  or

  (
    g396_n,
    g270_n_spl_,
    g359_p_spl_
  );


  and

  (
    g397_p,
    g274_p_spl_,
    g396_p
  );


  or

  (
    g397_n,
    g274_n_spl_,
    g396_n
  );


  and

  (
    g398_p,
    g115_n_spl_10,
    g397_p_spl_0
  );


  or

  (
    g398_n,
    g115_p_spl_10,
    g397_n_spl_0
  );


  and

  (
    g399_p,
    G25_p_spl_1,
    g398_n
  );


  and

  (
    g400_p,
    G25_n_spl_1,
    g398_p
  );


  or

  (
    g401_n,
    g399_p,
    g400_p
  );


  and

  (
    g402_p,
    g152_n_spl_10,
    g397_p_spl_0
  );


  or

  (
    g402_n,
    g152_p_spl_10,
    g397_n_spl_0
  );


  and

  (
    g403_p,
    G26_p_spl_1,
    g402_n
  );


  and

  (
    g404_p,
    G26_n_spl_1,
    g402_p
  );


  or

  (
    g405_n,
    g403_p,
    g404_p
  );


  and

  (
    g406_p,
    g191_n_spl_11,
    g397_p_spl_1
  );


  or

  (
    g406_n,
    g191_p_spl_11,
    g397_n_spl_1
  );


  and

  (
    g407_p,
    G27_p_spl_1,
    g406_n
  );


  and

  (
    g408_p,
    G27_n_spl_1,
    g406_p
  );


  or

  (
    g409_n,
    g407_p,
    g408_p
  );


  and

  (
    g410_p,
    g172_n_spl_11,
    g397_p_spl_1
  );


  or

  (
    g410_n,
    g172_p_spl_11,
    g397_n_spl_1
  );


  and

  (
    g411_p,
    G28_p_spl_1,
    g410_n
  );


  and

  (
    g412_p,
    G28_n_spl_1,
    g410_p
  );


  or

  (
    g413_n,
    g411_p,
    g412_p
  );


  and

  (
    g414_p,
    g271_p_spl_,
    g378_p_spl_
  );


  or

  (
    g414_n,
    g271_n_spl_,
    g378_n_spl_
  );


  and

  (
    g415_p,
    g115_n_spl_1,
    g414_p_spl_0
  );


  or

  (
    g415_n,
    g115_p_spl_1,
    g414_n_spl_0
  );


  and

  (
    g416_p,
    G29_p_spl_1,
    g415_n
  );


  and

  (
    g417_p,
    G29_n_spl_1,
    g415_p
  );


  or

  (
    g418_n,
    g416_p,
    g417_p
  );


  and

  (
    g419_p,
    g152_n_spl_1,
    g414_p_spl_0
  );


  or

  (
    g419_n,
    g152_p_spl_1,
    g414_n_spl_0
  );


  and

  (
    g420_p,
    G30_p_spl_1,
    g419_n
  );


  and

  (
    g421_p,
    G30_n_spl_1,
    g419_p
  );


  or

  (
    g422_n,
    g420_p,
    g421_p
  );


  and

  (
    g423_p,
    g191_n_spl_11,
    g414_p_spl_1
  );


  or

  (
    g423_n,
    g191_p_spl_11,
    g414_n_spl_1
  );


  and

  (
    g424_p,
    G31_p_spl_1,
    g423_n
  );


  and

  (
    g425_p,
    G31_n_spl_1,
    g423_p
  );


  or

  (
    g426_n,
    g424_p,
    g425_p
  );


  and

  (
    g427_p,
    g172_n_spl_11,
    g414_p_spl_1
  );


  or

  (
    g427_n,
    g172_p_spl_11,
    g414_n_spl_1
  );


  and

  (
    g428_p,
    G32_p_spl_1,
    g427_n
  );


  and

  (
    g429_p,
    G32_n_spl_1,
    g427_p
  );


  or

  (
    g430_n,
    g428_p,
    g429_p
  );


  not

  (
    G1324,
    g285_n
  );


  not

  (
    G1325,
    g289_n
  );


  not

  (
    G1326,
    g293_n
  );


  not

  (
    G1327,
    g297_n
  );


  not

  (
    G1328,
    g304_n
  );


  not

  (
    G1329,
    g308_n
  );


  not

  (
    G1330,
    g312_n
  );


  not

  (
    G1331,
    g316_n
  );


  not

  (
    G1332,
    g322_n
  );


  not

  (
    G1333,
    g326_n
  );


  not

  (
    G1334,
    g330_n
  );


  not

  (
    G1335,
    g334_n
  );


  not

  (
    G1336,
    g340_n
  );


  not

  (
    G1337,
    g344_n
  );


  not

  (
    G1338,
    g348_n
  );


  not

  (
    G1339,
    g352_n
  );


  not

  (
    G1340,
    g365_n
  );


  not

  (
    G1341,
    g369_n
  );


  not

  (
    G1342,
    g373_n
  );


  not

  (
    G1343,
    g377_n
  );


  not

  (
    G1344,
    g383_n
  );


  not

  (
    G1345,
    g387_n
  );


  not

  (
    G1346,
    g391_n
  );


  not

  (
    G1347,
    g395_n
  );


  not

  (
    G1348,
    g401_n
  );


  not

  (
    G1349,
    g405_n
  );


  not

  (
    G1350,
    g409_n
  );


  not

  (
    G1351,
    g413_n
  );


  not

  (
    G1352,
    g418_n
  );


  not

  (
    G1353,
    g422_n
  );


  not

  (
    G1354,
    g426_n
  );


  not

  (
    G1355,
    g430_n
  );


  buf

  (
    G9_n_spl_,
    G9_n
  );


  buf

  (
    G9_n_spl_0,
    G9_n_spl_
  );


  buf

  (
    G9_n_spl_00,
    G9_n_spl_0
  );


  buf

  (
    G9_n_spl_1,
    G9_n_spl_
  );


  buf

  (
    G13_n_spl_,
    G13_n
  );


  buf

  (
    G13_n_spl_0,
    G13_n_spl_
  );


  buf

  (
    G13_n_spl_00,
    G13_n_spl_0
  );


  buf

  (
    G13_n_spl_1,
    G13_n_spl_
  );


  buf

  (
    G9_p_spl_,
    G9_p
  );


  buf

  (
    G9_p_spl_0,
    G9_p_spl_
  );


  buf

  (
    G9_p_spl_00,
    G9_p_spl_0
  );


  buf

  (
    G9_p_spl_1,
    G9_p_spl_
  );


  buf

  (
    G13_p_spl_,
    G13_p
  );


  buf

  (
    G13_p_spl_0,
    G13_p_spl_
  );


  buf

  (
    G13_p_spl_00,
    G13_p_spl_0
  );


  buf

  (
    G13_p_spl_1,
    G13_p_spl_
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G1_p_spl_0,
    G1_p_spl_
  );


  buf

  (
    G1_p_spl_00,
    G1_p_spl_0
  );


  buf

  (
    G1_p_spl_1,
    G1_p_spl_
  );


  buf

  (
    G5_n_spl_,
    G5_n
  );


  buf

  (
    G5_n_spl_0,
    G5_n_spl_
  );


  buf

  (
    G5_n_spl_00,
    G5_n_spl_0
  );


  buf

  (
    G5_n_spl_1,
    G5_n_spl_
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G1_n_spl_0,
    G1_n_spl_
  );


  buf

  (
    G1_n_spl_00,
    G1_n_spl_0
  );


  buf

  (
    G1_n_spl_1,
    G1_n_spl_
  );


  buf

  (
    G5_p_spl_,
    G5_p
  );


  buf

  (
    G5_p_spl_0,
    G5_p_spl_
  );


  buf

  (
    G5_p_spl_00,
    G5_p_spl_0
  );


  buf

  (
    G5_p_spl_1,
    G5_p_spl_
  );


  buf

  (
    g44_n_spl_,
    g44_n
  );


  buf

  (
    g47_n_spl_,
    g47_n
  );


  buf

  (
    g44_p_spl_,
    g44_p
  );


  buf

  (
    g47_p_spl_,
    g47_p
  );


  buf

  (
    G41_p_spl_,
    G41_p
  );


  buf

  (
    G41_p_spl_0,
    G41_p_spl_
  );


  buf

  (
    G41_p_spl_00,
    G41_p_spl_0
  );


  buf

  (
    G41_p_spl_01,
    G41_p_spl_0
  );


  buf

  (
    G41_p_spl_1,
    G41_p_spl_
  );


  buf

  (
    G41_p_spl_10,
    G41_p_spl_1
  );


  buf

  (
    G41_p_spl_11,
    G41_p_spl_1
  );


  buf

  (
    G41_n_spl_,
    G41_n
  );


  buf

  (
    G41_n_spl_0,
    G41_n_spl_
  );


  buf

  (
    G41_n_spl_00,
    G41_n_spl_0
  );


  buf

  (
    G41_n_spl_01,
    G41_n_spl_0
  );


  buf

  (
    G41_n_spl_1,
    G41_n_spl_
  );


  buf

  (
    G41_n_spl_10,
    G41_n_spl_1
  );


  buf

  (
    G41_n_spl_11,
    G41_n_spl_1
  );


  buf

  (
    g50_n_spl_,
    g50_n
  );


  buf

  (
    g51_p_spl_,
    g51_p
  );


  buf

  (
    g50_p_spl_,
    g50_p
  );


  buf

  (
    g51_n_spl_,
    g51_n
  );


  buf

  (
    G19_n_spl_,
    G19_n
  );


  buf

  (
    G19_n_spl_0,
    G19_n_spl_
  );


  buf

  (
    G19_n_spl_00,
    G19_n_spl_0
  );


  buf

  (
    G19_n_spl_1,
    G19_n_spl_
  );


  buf

  (
    G20_n_spl_,
    G20_n
  );


  buf

  (
    G20_n_spl_0,
    G20_n_spl_
  );


  buf

  (
    G20_n_spl_00,
    G20_n_spl_0
  );


  buf

  (
    G20_n_spl_1,
    G20_n_spl_
  );


  buf

  (
    G19_p_spl_,
    G19_p
  );


  buf

  (
    G19_p_spl_0,
    G19_p_spl_
  );


  buf

  (
    G19_p_spl_00,
    G19_p_spl_0
  );


  buf

  (
    G19_p_spl_1,
    G19_p_spl_
  );


  buf

  (
    G20_p_spl_,
    G20_p
  );


  buf

  (
    G20_p_spl_0,
    G20_p_spl_
  );


  buf

  (
    G20_p_spl_00,
    G20_p_spl_0
  );


  buf

  (
    G20_p_spl_1,
    G20_p_spl_
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


  buf

  (
    G17_p_spl_0,
    G17_p_spl_
  );


  buf

  (
    G17_p_spl_00,
    G17_p_spl_0
  );


  buf

  (
    G17_p_spl_1,
    G17_p_spl_
  );


  buf

  (
    G18_n_spl_,
    G18_n
  );


  buf

  (
    G18_n_spl_0,
    G18_n_spl_
  );


  buf

  (
    G18_n_spl_00,
    G18_n_spl_0
  );


  buf

  (
    G18_n_spl_1,
    G18_n_spl_
  );


  buf

  (
    G17_n_spl_,
    G17_n
  );


  buf

  (
    G17_n_spl_0,
    G17_n_spl_
  );


  buf

  (
    G17_n_spl_00,
    G17_n_spl_0
  );


  buf

  (
    G17_n_spl_1,
    G17_n_spl_
  );


  buf

  (
    G18_p_spl_,
    G18_p
  );


  buf

  (
    G18_p_spl_0,
    G18_p_spl_
  );


  buf

  (
    G18_p_spl_00,
    G18_p_spl_0
  );


  buf

  (
    G18_p_spl_1,
    G18_p_spl_
  );


  buf

  (
    g57_n_spl_,
    g57_n
  );


  buf

  (
    g60_n_spl_,
    g60_n
  );


  buf

  (
    g57_p_spl_,
    g57_p
  );


  buf

  (
    g60_p_spl_,
    g60_p
  );


  buf

  (
    G23_n_spl_,
    G23_n
  );


  buf

  (
    G23_n_spl_0,
    G23_n_spl_
  );


  buf

  (
    G23_n_spl_00,
    G23_n_spl_0
  );


  buf

  (
    G23_n_spl_1,
    G23_n_spl_
  );


  buf

  (
    G24_n_spl_,
    G24_n
  );


  buf

  (
    G24_n_spl_0,
    G24_n_spl_
  );


  buf

  (
    G24_n_spl_00,
    G24_n_spl_0
  );


  buf

  (
    G24_n_spl_1,
    G24_n_spl_
  );


  buf

  (
    G23_p_spl_,
    G23_p
  );


  buf

  (
    G23_p_spl_0,
    G23_p_spl_
  );


  buf

  (
    G23_p_spl_00,
    G23_p_spl_0
  );


  buf

  (
    G23_p_spl_1,
    G23_p_spl_
  );


  buf

  (
    G24_p_spl_,
    G24_p
  );


  buf

  (
    G24_p_spl_0,
    G24_p_spl_
  );


  buf

  (
    G24_p_spl_00,
    G24_p_spl_0
  );


  buf

  (
    G24_p_spl_1,
    G24_p_spl_
  );


  buf

  (
    G21_p_spl_,
    G21_p
  );


  buf

  (
    G21_p_spl_0,
    G21_p_spl_
  );


  buf

  (
    G21_p_spl_00,
    G21_p_spl_0
  );


  buf

  (
    G21_p_spl_1,
    G21_p_spl_
  );


  buf

  (
    G22_n_spl_,
    G22_n
  );


  buf

  (
    G22_n_spl_0,
    G22_n_spl_
  );


  buf

  (
    G22_n_spl_00,
    G22_n_spl_0
  );


  buf

  (
    G22_n_spl_1,
    G22_n_spl_
  );


  buf

  (
    G21_n_spl_,
    G21_n
  );


  buf

  (
    G21_n_spl_0,
    G21_n_spl_
  );


  buf

  (
    G21_n_spl_00,
    G21_n_spl_0
  );


  buf

  (
    G21_n_spl_1,
    G21_n_spl_
  );


  buf

  (
    G22_p_spl_,
    G22_p
  );


  buf

  (
    G22_p_spl_0,
    G22_p_spl_
  );


  buf

  (
    G22_p_spl_00,
    G22_p_spl_0
  );


  buf

  (
    G22_p_spl_1,
    G22_p_spl_
  );


  buf

  (
    g66_n_spl_,
    g66_n
  );


  buf

  (
    g69_n_spl_,
    g69_n
  );


  buf

  (
    g66_p_spl_,
    g66_p
  );


  buf

  (
    g69_p_spl_,
    g69_p
  );


  buf

  (
    g63_n_spl_,
    g63_n
  );


  buf

  (
    g63_n_spl_0,
    g63_n_spl_
  );


  buf

  (
    g63_n_spl_1,
    g63_n_spl_
  );


  buf

  (
    g72_n_spl_,
    g72_n
  );


  buf

  (
    g72_n_spl_0,
    g72_n_spl_
  );


  buf

  (
    g72_n_spl_1,
    g72_n_spl_
  );


  buf

  (
    g63_p_spl_,
    g63_p
  );


  buf

  (
    g63_p_spl_0,
    g63_p_spl_
  );


  buf

  (
    g63_p_spl_1,
    g63_p_spl_
  );


  buf

  (
    g72_p_spl_,
    g72_p
  );


  buf

  (
    g72_p_spl_0,
    g72_p_spl_
  );


  buf

  (
    g72_p_spl_1,
    g72_p_spl_
  );


  buf

  (
    g54_n_spl_,
    g54_n
  );


  buf

  (
    g75_p_spl_,
    g75_p
  );


  buf

  (
    g54_p_spl_,
    g54_p
  );


  buf

  (
    g75_n_spl_,
    g75_n
  );


  buf

  (
    G25_n_spl_,
    G25_n
  );


  buf

  (
    G25_n_spl_0,
    G25_n_spl_
  );


  buf

  (
    G25_n_spl_00,
    G25_n_spl_0
  );


  buf

  (
    G25_n_spl_1,
    G25_n_spl_
  );


  buf

  (
    G29_n_spl_,
    G29_n
  );


  buf

  (
    G29_n_spl_0,
    G29_n_spl_
  );


  buf

  (
    G29_n_spl_00,
    G29_n_spl_0
  );


  buf

  (
    G29_n_spl_1,
    G29_n_spl_
  );


  buf

  (
    G25_p_spl_,
    G25_p
  );


  buf

  (
    G25_p_spl_0,
    G25_p_spl_
  );


  buf

  (
    G25_p_spl_00,
    G25_p_spl_0
  );


  buf

  (
    G25_p_spl_1,
    G25_p_spl_
  );


  buf

  (
    G29_p_spl_,
    G29_p
  );


  buf

  (
    G29_p_spl_0,
    G29_p_spl_
  );


  buf

  (
    G29_p_spl_00,
    G29_p_spl_0
  );


  buf

  (
    G29_p_spl_1,
    G29_p_spl_
  );


  buf

  (
    g81_n_spl_,
    g81_n
  );


  buf

  (
    g84_n_spl_,
    g84_n
  );


  buf

  (
    g81_p_spl_,
    g81_p
  );


  buf

  (
    g84_p_spl_,
    g84_p
  );


  buf

  (
    g87_n_spl_,
    g87_n
  );


  buf

  (
    g88_p_spl_,
    g88_p
  );


  buf

  (
    g87_p_spl_,
    g87_p
  );


  buf

  (
    g88_n_spl_,
    g88_n
  );


  buf

  (
    G7_n_spl_,
    G7_n
  );


  buf

  (
    G7_n_spl_0,
    G7_n_spl_
  );


  buf

  (
    G7_n_spl_00,
    G7_n_spl_0
  );


  buf

  (
    G7_n_spl_1,
    G7_n_spl_
  );


  buf

  (
    G8_n_spl_,
    G8_n
  );


  buf

  (
    G8_n_spl_0,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_00,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_1,
    G8_n_spl_
  );


  buf

  (
    G7_p_spl_,
    G7_p
  );


  buf

  (
    G7_p_spl_0,
    G7_p_spl_
  );


  buf

  (
    G7_p_spl_00,
    G7_p_spl_0
  );


  buf

  (
    G7_p_spl_1,
    G7_p_spl_
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_00,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_1,
    G8_p_spl_
  );


  buf

  (
    G6_n_spl_,
    G6_n
  );


  buf

  (
    G6_n_spl_0,
    G6_n_spl_
  );


  buf

  (
    G6_n_spl_00,
    G6_n_spl_0
  );


  buf

  (
    G6_n_spl_1,
    G6_n_spl_
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G6_p_spl_0,
    G6_p_spl_
  );


  buf

  (
    G6_p_spl_00,
    G6_p_spl_0
  );


  buf

  (
    G6_p_spl_1,
    G6_p_spl_
  );


  buf

  (
    g94_n_spl_,
    g94_n
  );


  buf

  (
    g97_n_spl_,
    g97_n
  );


  buf

  (
    g94_p_spl_,
    g94_p
  );


  buf

  (
    g97_p_spl_,
    g97_p
  );


  buf

  (
    G3_n_spl_,
    G3_n
  );


  buf

  (
    G3_n_spl_0,
    G3_n_spl_
  );


  buf

  (
    G3_n_spl_00,
    G3_n_spl_0
  );


  buf

  (
    G3_n_spl_1,
    G3_n_spl_
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    G4_n_spl_0,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_00,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_1,
    G4_n_spl_
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G3_p_spl_0,
    G3_p_spl_
  );


  buf

  (
    G3_p_spl_00,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_1,
    G3_p_spl_
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_00,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G2_n_spl_0,
    G2_n_spl_
  );


  buf

  (
    G2_n_spl_00,
    G2_n_spl_0
  );


  buf

  (
    G2_n_spl_1,
    G2_n_spl_
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G2_p_spl_0,
    G2_p_spl_
  );


  buf

  (
    G2_p_spl_00,
    G2_p_spl_0
  );


  buf

  (
    G2_p_spl_1,
    G2_p_spl_
  );


  buf

  (
    g103_n_spl_,
    g103_n
  );


  buf

  (
    g106_n_spl_,
    g106_n
  );


  buf

  (
    g103_p_spl_,
    g103_p
  );


  buf

  (
    g106_p_spl_,
    g106_p
  );


  buf

  (
    g100_n_spl_,
    g100_n
  );


  buf

  (
    g100_n_spl_0,
    g100_n_spl_
  );


  buf

  (
    g100_n_spl_1,
    g100_n_spl_
  );


  buf

  (
    g109_n_spl_,
    g109_n
  );


  buf

  (
    g109_n_spl_0,
    g109_n_spl_
  );


  buf

  (
    g109_n_spl_1,
    g109_n_spl_
  );


  buf

  (
    g100_p_spl_,
    g100_p
  );


  buf

  (
    g100_p_spl_0,
    g100_p_spl_
  );


  buf

  (
    g100_p_spl_1,
    g100_p_spl_
  );


  buf

  (
    g109_p_spl_,
    g109_p
  );


  buf

  (
    g109_p_spl_0,
    g109_p_spl_
  );


  buf

  (
    g109_p_spl_1,
    g109_p_spl_
  );


  buf

  (
    g91_n_spl_,
    g91_n
  );


  buf

  (
    g112_p_spl_,
    g112_p
  );


  buf

  (
    g91_p_spl_,
    g91_p
  );


  buf

  (
    g112_n_spl_,
    g112_n
  );


  buf

  (
    G26_n_spl_,
    G26_n
  );


  buf

  (
    G26_n_spl_0,
    G26_n_spl_
  );


  buf

  (
    G26_n_spl_00,
    G26_n_spl_0
  );


  buf

  (
    G26_n_spl_1,
    G26_n_spl_
  );


  buf

  (
    G30_n_spl_,
    G30_n
  );


  buf

  (
    G30_n_spl_0,
    G30_n_spl_
  );


  buf

  (
    G30_n_spl_00,
    G30_n_spl_0
  );


  buf

  (
    G30_n_spl_1,
    G30_n_spl_
  );


  buf

  (
    G26_p_spl_,
    G26_p
  );


  buf

  (
    G26_p_spl_0,
    G26_p_spl_
  );


  buf

  (
    G26_p_spl_00,
    G26_p_spl_0
  );


  buf

  (
    G26_p_spl_1,
    G26_p_spl_
  );


  buf

  (
    G30_p_spl_,
    G30_p
  );


  buf

  (
    G30_p_spl_0,
    G30_p_spl_
  );


  buf

  (
    G30_p_spl_00,
    G30_p_spl_0
  );


  buf

  (
    G30_p_spl_1,
    G30_p_spl_
  );


  buf

  (
    g118_n_spl_,
    g118_n
  );


  buf

  (
    g121_n_spl_,
    g121_n
  );


  buf

  (
    g118_p_spl_,
    g118_p
  );


  buf

  (
    g121_p_spl_,
    g121_p
  );


  buf

  (
    g124_n_spl_,
    g124_n
  );


  buf

  (
    g125_p_spl_,
    g125_p
  );


  buf

  (
    g124_p_spl_,
    g124_p
  );


  buf

  (
    g125_n_spl_,
    g125_n
  );


  buf

  (
    G15_n_spl_,
    G15_n
  );


  buf

  (
    G15_n_spl_0,
    G15_n_spl_
  );


  buf

  (
    G15_n_spl_00,
    G15_n_spl_0
  );


  buf

  (
    G15_n_spl_1,
    G15_n_spl_
  );


  buf

  (
    G16_n_spl_,
    G16_n
  );


  buf

  (
    G16_n_spl_0,
    G16_n_spl_
  );


  buf

  (
    G16_n_spl_00,
    G16_n_spl_0
  );


  buf

  (
    G16_n_spl_1,
    G16_n_spl_
  );


  buf

  (
    G15_p_spl_,
    G15_p
  );


  buf

  (
    G15_p_spl_0,
    G15_p_spl_
  );


  buf

  (
    G15_p_spl_00,
    G15_p_spl_0
  );


  buf

  (
    G15_p_spl_1,
    G15_p_spl_
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    G16_p_spl_0,
    G16_p_spl_
  );


  buf

  (
    G16_p_spl_00,
    G16_p_spl_0
  );


  buf

  (
    G16_p_spl_1,
    G16_p_spl_
  );


  buf

  (
    G14_n_spl_,
    G14_n
  );


  buf

  (
    G14_n_spl_0,
    G14_n_spl_
  );


  buf

  (
    G14_n_spl_00,
    G14_n_spl_0
  );


  buf

  (
    G14_n_spl_1,
    G14_n_spl_
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G14_p_spl_0,
    G14_p_spl_
  );


  buf

  (
    G14_p_spl_00,
    G14_p_spl_0
  );


  buf

  (
    G14_p_spl_1,
    G14_p_spl_
  );


  buf

  (
    g131_n_spl_,
    g131_n
  );


  buf

  (
    g134_n_spl_,
    g134_n
  );


  buf

  (
    g131_p_spl_,
    g131_p
  );


  buf

  (
    g134_p_spl_,
    g134_p
  );


  buf

  (
    G11_n_spl_,
    G11_n
  );


  buf

  (
    G11_n_spl_0,
    G11_n_spl_
  );


  buf

  (
    G11_n_spl_00,
    G11_n_spl_0
  );


  buf

  (
    G11_n_spl_1,
    G11_n_spl_
  );


  buf

  (
    G12_n_spl_,
    G12_n
  );


  buf

  (
    G12_n_spl_0,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_00,
    G12_n_spl_0
  );


  buf

  (
    G12_n_spl_1,
    G12_n_spl_
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    G11_p_spl_0,
    G11_p_spl_
  );


  buf

  (
    G11_p_spl_00,
    G11_p_spl_0
  );


  buf

  (
    G11_p_spl_1,
    G11_p_spl_
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G12_p_spl_0,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_00,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_1,
    G12_p_spl_
  );


  buf

  (
    G10_n_spl_,
    G10_n
  );


  buf

  (
    G10_n_spl_0,
    G10_n_spl_
  );


  buf

  (
    G10_n_spl_00,
    G10_n_spl_0
  );


  buf

  (
    G10_n_spl_1,
    G10_n_spl_
  );


  buf

  (
    G10_p_spl_,
    G10_p
  );


  buf

  (
    G10_p_spl_0,
    G10_p_spl_
  );


  buf

  (
    G10_p_spl_00,
    G10_p_spl_0
  );


  buf

  (
    G10_p_spl_1,
    G10_p_spl_
  );


  buf

  (
    g140_n_spl_,
    g140_n
  );


  buf

  (
    g143_n_spl_,
    g143_n
  );


  buf

  (
    g140_p_spl_,
    g140_p
  );


  buf

  (
    g143_p_spl_,
    g143_p
  );


  buf

  (
    g137_n_spl_,
    g137_n
  );


  buf

  (
    g137_n_spl_0,
    g137_n_spl_
  );


  buf

  (
    g137_n_spl_1,
    g137_n_spl_
  );


  buf

  (
    g146_n_spl_,
    g146_n
  );


  buf

  (
    g146_n_spl_0,
    g146_n_spl_
  );


  buf

  (
    g146_n_spl_1,
    g146_n_spl_
  );


  buf

  (
    g137_p_spl_,
    g137_p
  );


  buf

  (
    g137_p_spl_0,
    g137_p_spl_
  );


  buf

  (
    g137_p_spl_1,
    g137_p_spl_
  );


  buf

  (
    g146_p_spl_,
    g146_p
  );


  buf

  (
    g146_p_spl_0,
    g146_p_spl_
  );


  buf

  (
    g146_p_spl_1,
    g146_p_spl_
  );


  buf

  (
    g128_n_spl_,
    g128_n
  );


  buf

  (
    g149_p_spl_,
    g149_p
  );


  buf

  (
    g128_p_spl_,
    g128_p
  );


  buf

  (
    g149_n_spl_,
    g149_n
  );


  buf

  (
    g115_n_spl_,
    g115_n
  );


  buf

  (
    g115_n_spl_0,
    g115_n_spl_
  );


  buf

  (
    g115_n_spl_00,
    g115_n_spl_0
  );


  buf

  (
    g115_n_spl_01,
    g115_n_spl_0
  );


  buf

  (
    g115_n_spl_1,
    g115_n_spl_
  );


  buf

  (
    g115_n_spl_10,
    g115_n_spl_1
  );


  buf

  (
    g152_p_spl_,
    g152_p
  );


  buf

  (
    g152_p_spl_0,
    g152_p_spl_
  );


  buf

  (
    g152_p_spl_00,
    g152_p_spl_0
  );


  buf

  (
    g152_p_spl_01,
    g152_p_spl_0
  );


  buf

  (
    g152_p_spl_1,
    g152_p_spl_
  );


  buf

  (
    g152_p_spl_10,
    g152_p_spl_1
  );


  buf

  (
    g115_p_spl_,
    g115_p
  );


  buf

  (
    g115_p_spl_0,
    g115_p_spl_
  );


  buf

  (
    g115_p_spl_00,
    g115_p_spl_0
  );


  buf

  (
    g115_p_spl_01,
    g115_p_spl_0
  );


  buf

  (
    g115_p_spl_1,
    g115_p_spl_
  );


  buf

  (
    g115_p_spl_10,
    g115_p_spl_1
  );


  buf

  (
    g152_n_spl_,
    g152_n
  );


  buf

  (
    g152_n_spl_0,
    g152_n_spl_
  );


  buf

  (
    g152_n_spl_00,
    g152_n_spl_0
  );


  buf

  (
    g152_n_spl_01,
    g152_n_spl_0
  );


  buf

  (
    g152_n_spl_1,
    g152_n_spl_
  );


  buf

  (
    g152_n_spl_10,
    g152_n_spl_1
  );


  buf

  (
    G28_n_spl_,
    G28_n
  );


  buf

  (
    G28_n_spl_0,
    G28_n_spl_
  );


  buf

  (
    G28_n_spl_00,
    G28_n_spl_0
  );


  buf

  (
    G28_n_spl_1,
    G28_n_spl_
  );


  buf

  (
    G32_n_spl_,
    G32_n
  );


  buf

  (
    G32_n_spl_0,
    G32_n_spl_
  );


  buf

  (
    G32_n_spl_00,
    G32_n_spl_0
  );


  buf

  (
    G32_n_spl_1,
    G32_n_spl_
  );


  buf

  (
    G28_p_spl_,
    G28_p
  );


  buf

  (
    G28_p_spl_0,
    G28_p_spl_
  );


  buf

  (
    G28_p_spl_00,
    G28_p_spl_0
  );


  buf

  (
    G28_p_spl_1,
    G28_p_spl_
  );


  buf

  (
    G32_p_spl_,
    G32_p
  );


  buf

  (
    G32_p_spl_0,
    G32_p_spl_
  );


  buf

  (
    G32_p_spl_00,
    G32_p_spl_0
  );


  buf

  (
    G32_p_spl_1,
    G32_p_spl_
  );


  buf

  (
    g156_n_spl_,
    g156_n
  );


  buf

  (
    g159_n_spl_,
    g159_n
  );


  buf

  (
    g156_p_spl_,
    g156_p
  );


  buf

  (
    g159_p_spl_,
    g159_p
  );


  buf

  (
    g162_n_spl_,
    g162_n
  );


  buf

  (
    g163_p_spl_,
    g163_p
  );


  buf

  (
    g162_p_spl_,
    g162_p
  );


  buf

  (
    g163_n_spl_,
    g163_n
  );


  buf

  (
    g166_n_spl_,
    g166_n
  );


  buf

  (
    g169_p_spl_,
    g169_p
  );


  buf

  (
    g166_p_spl_,
    g166_p
  );


  buf

  (
    g169_n_spl_,
    g169_n
  );


  buf

  (
    G27_n_spl_,
    G27_n
  );


  buf

  (
    G27_n_spl_0,
    G27_n_spl_
  );


  buf

  (
    G27_n_spl_00,
    G27_n_spl_0
  );


  buf

  (
    G27_n_spl_1,
    G27_n_spl_
  );


  buf

  (
    G31_n_spl_,
    G31_n
  );


  buf

  (
    G31_n_spl_0,
    G31_n_spl_
  );


  buf

  (
    G31_n_spl_00,
    G31_n_spl_0
  );


  buf

  (
    G31_n_spl_1,
    G31_n_spl_
  );


  buf

  (
    G27_p_spl_,
    G27_p
  );


  buf

  (
    G27_p_spl_0,
    G27_p_spl_
  );


  buf

  (
    G27_p_spl_00,
    G27_p_spl_0
  );


  buf

  (
    G27_p_spl_1,
    G27_p_spl_
  );


  buf

  (
    G31_p_spl_,
    G31_p
  );


  buf

  (
    G31_p_spl_0,
    G31_p_spl_
  );


  buf

  (
    G31_p_spl_00,
    G31_p_spl_0
  );


  buf

  (
    G31_p_spl_1,
    G31_p_spl_
  );


  buf

  (
    g175_n_spl_,
    g175_n
  );


  buf

  (
    g178_n_spl_,
    g178_n
  );


  buf

  (
    g175_p_spl_,
    g175_p
  );


  buf

  (
    g178_p_spl_,
    g178_p
  );


  buf

  (
    g181_n_spl_,
    g181_n
  );


  buf

  (
    g182_p_spl_,
    g182_p
  );


  buf

  (
    g181_p_spl_,
    g181_p
  );


  buf

  (
    g182_n_spl_,
    g182_n
  );


  buf

  (
    g185_n_spl_,
    g185_n
  );


  buf

  (
    g188_p_spl_,
    g188_p
  );


  buf

  (
    g185_p_spl_,
    g185_p
  );


  buf

  (
    g188_n_spl_,
    g188_n
  );


  buf

  (
    g172_p_spl_,
    g172_p
  );


  buf

  (
    g172_p_spl_0,
    g172_p_spl_
  );


  buf

  (
    g172_p_spl_00,
    g172_p_spl_0
  );


  buf

  (
    g172_p_spl_01,
    g172_p_spl_0
  );


  buf

  (
    g172_p_spl_1,
    g172_p_spl_
  );


  buf

  (
    g172_p_spl_10,
    g172_p_spl_1
  );


  buf

  (
    g172_p_spl_11,
    g172_p_spl_1
  );


  buf

  (
    g191_n_spl_,
    g191_n
  );


  buf

  (
    g191_n_spl_0,
    g191_n_spl_
  );


  buf

  (
    g191_n_spl_00,
    g191_n_spl_0
  );


  buf

  (
    g191_n_spl_01,
    g191_n_spl_0
  );


  buf

  (
    g191_n_spl_1,
    g191_n_spl_
  );


  buf

  (
    g191_n_spl_10,
    g191_n_spl_1
  );


  buf

  (
    g191_n_spl_11,
    g191_n_spl_1
  );


  buf

  (
    g172_n_spl_,
    g172_n
  );


  buf

  (
    g172_n_spl_0,
    g172_n_spl_
  );


  buf

  (
    g172_n_spl_00,
    g172_n_spl_0
  );


  buf

  (
    g172_n_spl_01,
    g172_n_spl_0
  );


  buf

  (
    g172_n_spl_1,
    g172_n_spl_
  );


  buf

  (
    g172_n_spl_10,
    g172_n_spl_1
  );


  buf

  (
    g172_n_spl_11,
    g172_n_spl_1
  );


  buf

  (
    g191_p_spl_,
    g191_p
  );


  buf

  (
    g191_p_spl_0,
    g191_p_spl_
  );


  buf

  (
    g191_p_spl_00,
    g191_p_spl_0
  );


  buf

  (
    g191_p_spl_01,
    g191_p_spl_0
  );


  buf

  (
    g191_p_spl_1,
    g191_p_spl_
  );


  buf

  (
    g191_p_spl_10,
    g191_p_spl_1
  );


  buf

  (
    g191_p_spl_11,
    g191_p_spl_1
  );


  buf

  (
    g195_n_spl_,
    g195_n
  );


  buf

  (
    g198_n_spl_,
    g198_n
  );


  buf

  (
    g195_p_spl_,
    g195_p
  );


  buf

  (
    g198_p_spl_,
    g198_p
  );


  buf

  (
    g201_n_spl_,
    g201_n
  );


  buf

  (
    g202_p_spl_,
    g202_p
  );


  buf

  (
    g201_p_spl_,
    g201_p
  );


  buf

  (
    g202_n_spl_,
    g202_n
  );


  buf

  (
    g208_n_spl_,
    g208_n
  );


  buf

  (
    g211_n_spl_,
    g211_n
  );


  buf

  (
    g208_p_spl_,
    g208_p
  );


  buf

  (
    g211_p_spl_,
    g211_p
  );


  buf

  (
    g214_n_spl_,
    g214_n
  );


  buf

  (
    g214_n_spl_0,
    g214_n_spl_
  );


  buf

  (
    g214_n_spl_1,
    g214_n_spl_
  );


  buf

  (
    g214_p_spl_,
    g214_p
  );


  buf

  (
    g214_p_spl_0,
    g214_p_spl_
  );


  buf

  (
    g214_p_spl_1,
    g214_p_spl_
  );


  buf

  (
    g205_n_spl_,
    g205_n
  );


  buf

  (
    g217_p_spl_,
    g217_p
  );


  buf

  (
    g205_p_spl_,
    g205_p
  );


  buf

  (
    g217_n_spl_,
    g217_n
  );


  buf

  (
    g223_n_spl_,
    g223_n
  );


  buf

  (
    g226_n_spl_,
    g226_n
  );


  buf

  (
    g223_p_spl_,
    g223_p
  );


  buf

  (
    g226_p_spl_,
    g226_p
  );


  buf

  (
    g229_n_spl_,
    g229_n
  );


  buf

  (
    g230_p_spl_,
    g230_p
  );


  buf

  (
    g229_p_spl_,
    g229_p
  );


  buf

  (
    g230_n_spl_,
    g230_n
  );


  buf

  (
    g236_n_spl_,
    g236_n
  );


  buf

  (
    g239_n_spl_,
    g239_n
  );


  buf

  (
    g236_p_spl_,
    g236_p
  );


  buf

  (
    g239_p_spl_,
    g239_p
  );


  buf

  (
    g242_n_spl_,
    g242_n
  );


  buf

  (
    g242_n_spl_0,
    g242_n_spl_
  );


  buf

  (
    g242_n_spl_1,
    g242_n_spl_
  );


  buf

  (
    g242_p_spl_,
    g242_p
  );


  buf

  (
    g242_p_spl_0,
    g242_p_spl_
  );


  buf

  (
    g242_p_spl_1,
    g242_p_spl_
  );


  buf

  (
    g233_n_spl_,
    g233_n
  );


  buf

  (
    g245_p_spl_,
    g245_p
  );


  buf

  (
    g233_p_spl_,
    g233_p
  );


  buf

  (
    g245_n_spl_,
    g245_n
  );


  buf

  (
    g251_n_spl_,
    g251_n
  );


  buf

  (
    g254_n_spl_,
    g254_n
  );


  buf

  (
    g251_p_spl_,
    g251_p
  );


  buf

  (
    g254_p_spl_,
    g254_p
  );


  buf

  (
    g257_n_spl_,
    g257_n
  );


  buf

  (
    g258_p_spl_,
    g258_p
  );


  buf

  (
    g257_p_spl_,
    g257_p
  );


  buf

  (
    g258_n_spl_,
    g258_n
  );


  buf

  (
    g261_n_spl_,
    g261_n
  );


  buf

  (
    g264_p_spl_,
    g264_p
  );


  buf

  (
    g261_p_spl_,
    g261_p
  );


  buf

  (
    g264_n_spl_,
    g264_n
  );


  buf

  (
    g78_n_spl_,
    g78_n
  );


  buf

  (
    g78_n_spl_0,
    g78_n_spl_
  );


  buf

  (
    g78_n_spl_00,
    g78_n_spl_0
  );


  buf

  (
    g78_n_spl_01,
    g78_n_spl_0
  );


  buf

  (
    g78_n_spl_1,
    g78_n_spl_
  );


  buf

  (
    g78_n_spl_10,
    g78_n_spl_1
  );


  buf

  (
    g267_p_spl_,
    g267_p
  );


  buf

  (
    g267_p_spl_0,
    g267_p_spl_
  );


  buf

  (
    g267_p_spl_00,
    g267_p_spl_0
  );


  buf

  (
    g267_p_spl_01,
    g267_p_spl_0
  );


  buf

  (
    g267_p_spl_1,
    g267_p_spl_
  );


  buf

  (
    g267_p_spl_10,
    g267_p_spl_1
  );


  buf

  (
    g78_p_spl_,
    g78_p
  );


  buf

  (
    g78_p_spl_0,
    g78_p_spl_
  );


  buf

  (
    g78_p_spl_00,
    g78_p_spl_0
  );


  buf

  (
    g78_p_spl_01,
    g78_p_spl_0
  );


  buf

  (
    g78_p_spl_1,
    g78_p_spl_
  );


  buf

  (
    g78_p_spl_10,
    g78_p_spl_1
  );


  buf

  (
    g267_n_spl_,
    g267_n
  );


  buf

  (
    g267_n_spl_0,
    g267_n_spl_
  );


  buf

  (
    g267_n_spl_00,
    g267_n_spl_0
  );


  buf

  (
    g267_n_spl_01,
    g267_n_spl_0
  );


  buf

  (
    g267_n_spl_1,
    g267_n_spl_
  );


  buf

  (
    g267_n_spl_10,
    g267_n_spl_1
  );


  buf

  (
    g248_p_spl_,
    g248_p
  );


  buf

  (
    g248_p_spl_0,
    g248_p_spl_
  );


  buf

  (
    g248_p_spl_00,
    g248_p_spl_0
  );


  buf

  (
    g248_p_spl_01,
    g248_p_spl_0
  );


  buf

  (
    g248_p_spl_1,
    g248_p_spl_
  );


  buf

  (
    g248_p_spl_10,
    g248_p_spl_1
  );


  buf

  (
    g248_p_spl_11,
    g248_p_spl_1
  );


  buf

  (
    g268_p_spl_,
    g268_p
  );


  buf

  (
    g248_n_spl_,
    g248_n
  );


  buf

  (
    g248_n_spl_0,
    g248_n_spl_
  );


  buf

  (
    g248_n_spl_00,
    g248_n_spl_0
  );


  buf

  (
    g248_n_spl_01,
    g248_n_spl_0
  );


  buf

  (
    g248_n_spl_1,
    g248_n_spl_
  );


  buf

  (
    g248_n_spl_10,
    g248_n_spl_1
  );


  buf

  (
    g248_n_spl_11,
    g248_n_spl_1
  );


  buf

  (
    g268_n_spl_,
    g268_n
  );


  buf

  (
    g270_p_spl_,
    g270_p
  );


  buf

  (
    g270_n_spl_,
    g270_n
  );


  buf

  (
    g269_n_spl_,
    g269_n
  );


  buf

  (
    g271_n_spl_,
    g271_n
  );


  buf

  (
    g269_p_spl_,
    g269_p
  );


  buf

  (
    g271_p_spl_,
    g271_p
  );


  buf

  (
    g220_p_spl_,
    g220_p
  );


  buf

  (
    g220_p_spl_0,
    g220_p_spl_
  );


  buf

  (
    g220_p_spl_00,
    g220_p_spl_0
  );


  buf

  (
    g220_p_spl_01,
    g220_p_spl_0
  );


  buf

  (
    g220_p_spl_1,
    g220_p_spl_
  );


  buf

  (
    g220_p_spl_10,
    g220_p_spl_1
  );


  buf

  (
    g220_p_spl_11,
    g220_p_spl_1
  );


  buf

  (
    g220_n_spl_,
    g220_n
  );


  buf

  (
    g220_n_spl_0,
    g220_n_spl_
  );


  buf

  (
    g220_n_spl_00,
    g220_n_spl_0
  );


  buf

  (
    g220_n_spl_01,
    g220_n_spl_0
  );


  buf

  (
    g220_n_spl_1,
    g220_n_spl_
  );


  buf

  (
    g220_n_spl_10,
    g220_n_spl_1
  );


  buf

  (
    g220_n_spl_11,
    g220_n_spl_1
  );


  buf

  (
    g274_n_spl_,
    g274_n
  );


  buf

  (
    g274_n_spl_0,
    g274_n_spl_
  );


  buf

  (
    g274_p_spl_,
    g274_p
  );


  buf

  (
    g274_p_spl_0,
    g274_p_spl_
  );


  buf

  (
    g192_p_spl_,
    g192_p
  );


  buf

  (
    g279_n_spl_,
    g279_n
  );


  buf

  (
    g192_n_spl_,
    g192_n
  );


  buf

  (
    g279_p_spl_,
    g279_p
  );


  buf

  (
    g153_p_spl_,
    g153_p
  );


  buf

  (
    g280_p_spl_,
    g280_p
  );


  buf

  (
    g153_n_spl_,
    g153_n
  );


  buf

  (
    g280_n_spl_,
    g280_n
  );


  buf

  (
    g281_p_spl_,
    g281_p
  );


  buf

  (
    g281_p_spl_0,
    g281_p_spl_
  );


  buf

  (
    g281_p_spl_1,
    g281_p_spl_
  );


  buf

  (
    g281_n_spl_,
    g281_n
  );


  buf

  (
    g281_n_spl_0,
    g281_n_spl_
  );


  buf

  (
    g281_n_spl_1,
    g281_n_spl_
  );


  buf

  (
    g298_p_spl_,
    g298_p
  );


  buf

  (
    g299_p_spl_,
    g299_p
  );


  buf

  (
    g298_n_spl_,
    g298_n
  );


  buf

  (
    g299_n_spl_,
    g299_n
  );


  buf

  (
    g300_p_spl_,
    g300_p
  );


  buf

  (
    g300_p_spl_0,
    g300_p_spl_
  );


  buf

  (
    g300_p_spl_1,
    g300_p_spl_
  );


  buf

  (
    g300_n_spl_,
    g300_n
  );


  buf

  (
    g300_n_spl_0,
    g300_n_spl_
  );


  buf

  (
    g300_n_spl_1,
    g300_n_spl_
  );


  buf

  (
    g317_p_spl_,
    g317_p
  );


  buf

  (
    g317_n_spl_,
    g317_n
  );


  buf

  (
    g318_p_spl_,
    g318_p
  );


  buf

  (
    g318_p_spl_0,
    g318_p_spl_
  );


  buf

  (
    g318_p_spl_1,
    g318_p_spl_
  );


  buf

  (
    g318_n_spl_,
    g318_n
  );


  buf

  (
    g318_n_spl_0,
    g318_n_spl_
  );


  buf

  (
    g318_n_spl_1,
    g318_n_spl_
  );


  buf

  (
    g335_p_spl_,
    g335_p
  );


  buf

  (
    g335_n_spl_,
    g335_n
  );


  buf

  (
    g336_p_spl_,
    g336_p
  );


  buf

  (
    g336_p_spl_0,
    g336_p_spl_
  );


  buf

  (
    g336_p_spl_1,
    g336_p_spl_
  );


  buf

  (
    g336_n_spl_,
    g336_n
  );


  buf

  (
    g336_n_spl_0,
    g336_n_spl_
  );


  buf

  (
    g336_n_spl_1,
    g336_n_spl_
  );


  buf

  (
    g359_n_spl_,
    g359_n
  );


  buf

  (
    g359_n_spl_0,
    g359_n_spl_
  );


  buf

  (
    g359_p_spl_,
    g359_p
  );


  buf

  (
    g359_p_spl_0,
    g359_p_spl_
  );


  buf

  (
    g361_p_spl_,
    g361_p
  );


  buf

  (
    g361_p_spl_0,
    g361_p_spl_
  );


  buf

  (
    g361_p_spl_1,
    g361_p_spl_
  );


  buf

  (
    g361_n_spl_,
    g361_n
  );


  buf

  (
    g361_n_spl_0,
    g361_n_spl_
  );


  buf

  (
    g361_n_spl_1,
    g361_n_spl_
  );


  buf

  (
    g378_p_spl_,
    g378_p
  );


  buf

  (
    g378_n_spl_,
    g378_n
  );


  buf

  (
    g379_p_spl_,
    g379_p
  );


  buf

  (
    g379_p_spl_0,
    g379_p_spl_
  );


  buf

  (
    g379_p_spl_1,
    g379_p_spl_
  );


  buf

  (
    g379_n_spl_,
    g379_n
  );


  buf

  (
    g379_n_spl_0,
    g379_n_spl_
  );


  buf

  (
    g379_n_spl_1,
    g379_n_spl_
  );


  buf

  (
    g397_p_spl_,
    g397_p
  );


  buf

  (
    g397_p_spl_0,
    g397_p_spl_
  );


  buf

  (
    g397_p_spl_1,
    g397_p_spl_
  );


  buf

  (
    g397_n_spl_,
    g397_n
  );


  buf

  (
    g397_n_spl_0,
    g397_n_spl_
  );


  buf

  (
    g397_n_spl_1,
    g397_n_spl_
  );


  buf

  (
    g414_p_spl_,
    g414_p
  );


  buf

  (
    g414_p_spl_0,
    g414_p_spl_
  );


  buf

  (
    g414_p_spl_1,
    g414_p_spl_
  );


  buf

  (
    g414_n_spl_,
    g414_n
  );


  buf

  (
    g414_n_spl_0,
    g414_n_spl_
  );


  buf

  (
    g414_n_spl_1,
    g414_n_spl_
  );


endmodule
