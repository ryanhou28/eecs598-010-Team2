
module mymod
(
  G1_p,
  G1_n,
  G2_p,
  G2_n,
  G3_p,
  G3_n,
  G4_p,
  G4_n,
  G5_p,
  G5_n,
  G6_p,
  G6_n,
  G7_p,
  G7_n,
  G8_p,
  G8_n,
  G9_p,
  G9_n,
  G10_p,
  G10_n,
  G11_p,
  G11_n,
  G12_p,
  G12_n,
  G13_p,
  G13_n,
  G14_p,
  G14_n,
  G15_p,
  G15_n,
  G16_p,
  G16_n,
  G17_p,
  G17_n,
  G18_p,
  G18_n,
  G19_p,
  G19_n,
  G20_p,
  G20_n,
  G21_p,
  G21_n,
  G22_p,
  G22_n,
  G23_p,
  G23_n,
  G24_p,
  G24_n,
  G25_p,
  G25_n,
  G26_p,
  G26_n,
  G27_p,
  G27_n,
  G28_p,
  G28_n,
  G29_p,
  G29_n,
  G30_p,
  G30_n,
  G31_p,
  G31_n,
  G32_p,
  G32_n,
  G33_p,
  G33_n,
  G34_p,
  G34_n,
  G35_p,
  G35_n,
  G36_p,
  G36_n,
  G37_p,
  G37_n,
  G38_p,
  G38_n,
  G39_p,
  G39_n,
  G40_p,
  G40_n,
  G41_p,
  G41_n,
  G42_p,
  G42_n,
  G43_p,
  G43_n,
  G44_p,
  G44_n,
  G45_p,
  G45_n,
  G46_p,
  G46_n,
  G47_p,
  G47_n,
  G48_p,
  G48_n,
  G49_p,
  G49_n,
  G50_p,
  G50_n,
  G51_p,
  G51_n,
  G52_p,
  G52_n,
  G53_p,
  G53_n,
  G54_p,
  G54_n,
  G55_p,
  G55_n,
  G56_p,
  G56_n,
  G57_p,
  G57_n,
  G58_p,
  G58_n,
  G59_p,
  G59_n,
  G60_p,
  G60_n,
  G61_p,
  G61_n,
  G62_p,
  G62_n,
  G63_p,
  G63_n,
  G64_p,
  G64_n,
  G65_p,
  G65_n,
  G66_p,
  G66_n,
  G67_p,
  G67_n,
  G68_p,
  G68_n,
  G69_p,
  G69_n,
  G70_p,
  G70_n,
  G71_p,
  G71_n,
  G72_p,
  G72_n,
  G73_p,
  G73_n,
  G74_p,
  G74_n,
  G75_p,
  G75_n,
  G76_p,
  G76_n,
  G77_p,
  G77_n,
  G78_p,
  G78_n,
  G79_p,
  G79_n,
  G80_p,
  G80_n,
  G81_p,
  G81_n,
  G82_p,
  G82_n,
  G83_p,
  G83_n,
  G84_p,
  G84_n,
  G85_p,
  G85_n,
  G86_p,
  G86_n,
  G87_p,
  G87_n,
  G88_p,
  G88_n,
  G89_p,
  G89_n,
  G90_p,
  G90_n,
  G91_p,
  G91_n,
  G92_p,
  G92_n,
  G93_p,
  G93_n,
  G94_p,
  G94_n,
  G95_p,
  G95_n,
  G96_p,
  G96_n,
  G97_p,
  G97_n,
  G98_p,
  G98_n,
  G99_p,
  G99_n,
  G100_p,
  G100_n,
  G101_p,
  G101_n,
  G102_p,
  G102_n,
  G103_p,
  G103_n,
  G104_p,
  G104_n,
  G105_p,
  G105_n,
  G106_p,
  G106_n,
  G107_p,
  G107_n,
  G108_p,
  G108_n,
  G109_p,
  G109_n,
  G110_p,
  G110_n,
  G111_p,
  G111_n,
  G112_p,
  G112_n,
  G113_p,
  G113_n,
  G114_p,
  G114_n,
  G115_p,
  G115_n,
  G116_p,
  G116_n,
  G117_p,
  G117_n,
  G118_p,
  G118_n,
  G119_p,
  G119_n,
  G120_p,
  G120_n,
  G121_p,
  G121_n,
  G122_p,
  G122_n,
  G123_p,
  G123_n,
  G124_p,
  G124_n,
  G125_p,
  G125_n,
  G126_p,
  G126_n,
  G127_p,
  G127_n,
  G128_p,
  G128_n,
  G129_p,
  G129_n,
  G130_p,
  G130_n,
  G131_p,
  G131_n,
  G132_p,
  G132_n,
  G133_p,
  G133_n,
  G134_p,
  G134_n,
  G135_p,
  G135_n,
  G136_p,
  G136_n,
  G137_p,
  G137_n,
  G138_p,
  G138_n,
  G139_p,
  G139_n,
  G140_p,
  G140_n,
  G141_p,
  G141_n,
  G142_p,
  G142_n,
  G143_p,
  G143_n,
  G144_p,
  G144_n,
  G145_p,
  G145_n,
  G146_p,
  G146_n,
  G147_p,
  G147_n,
  G148_p,
  G148_n,
  G149_p,
  G149_n,
  G150_p,
  G150_n,
  G151_p,
  G151_n,
  G152_p,
  G152_n,
  G153_p,
  G153_n,
  G154_p,
  G154_n,
  G155_p,
  G155_n,
  G156_p,
  G156_n,
  G157_p,
  G157_n,
  G158_p,
  G158_n,
  G159_p,
  G159_n,
  G160_p,
  G160_n,
  G161_p,
  G161_n,
  G162_p,
  G162_n,
  G163_p,
  G163_n,
  G164_p,
  G164_n,
  G165_p,
  G165_n,
  G166_p,
  G166_n,
  G167_p,
  G167_n,
  G168_p,
  G168_n,
  G169_p,
  G169_n,
  G170_p,
  G170_n,
  G171_p,
  G171_n,
  G172_p,
  G172_n,
  G173_p,
  G173_n,
  G174_p,
  G174_n,
  G175_p,
  G175_n,
  G176_p,
  G176_n,
  G177_p,
  G177_n,
  G178_p,
  G178_n,
  G5193_p,
  G5194_p,
  G5195_p,
  G5196_p,
  G5197_p,
  G5198_p,
  G5199_n,
  G5200_p,
  G5201_p,
  G5202_p,
  G5203_p,
  G5204_p,
  G5205_p,
  G5206_p,
  G5207_p,
  G5208_p,
  G5209_p,
  G5210_p,
  G5211_p,
  G5212_p,
  G5213_p,
  G5214_p,
  G5215_p,
  G5216_p,
  G5217_p,
  G5218_p,
  G5219_p,
  G5220_p,
  G5221_p,
  G5222_p,
  G5223_p,
  G5224_p,
  G5225_p,
  G5226_p,
  G5227_p,
  G5228_p,
  G5229_p,
  G5230_p,
  G5231_p,
  G5232_p,
  G5233_p,
  G5234_p,
  G5235_p,
  G5236_n,
  G5237_n,
  G5238_n,
  G5239_p,
  G5240_p,
  G5241_n,
  G5242_n,
  G5243_n,
  G5244_n,
  G5245_p,
  G5246_n,
  G5247_p,
  G5248_n,
  G5249_n,
  G5250_n,
  G5251_p,
  G5252_p,
  G5253_n,
  G5254_n,
  G5255_n,
  G5256_p,
  G5257_n,
  G5258_n,
  G5259_n,
  G5260_n,
  G5261_n,
  G5262_n,
  G5263_n,
  G5264_n,
  G5265_p,
  G5266_p,
  G5267_p,
  G5268_p,
  G5269_p,
  G5270_p,
  G5271_p,
  G5272_p,
  G5273_p,
  G5274_p,
  G5275_p,
  G5276_p,
  G5277_p,
  G5278_p,
  G5279_p,
  G5280_p,
  G5281_p,
  G5282_p,
  G5283_p,
  G5284_p,
  G5285_n,
  G5286_n,
  G5287_n,
  G5288_n,
  G5289_n,
  G5290_n,
  G5291_n,
  G5292_n,
  G5293_n,
  G5294_p,
  G5295_p,
  G5296_p,
  G5297_p,
  G5298_p,
  G5299_p,
  G5300_p,
  G5301_p,
  G5302_p,
  G5303_p,
  G5304_p,
  G5305_p,
  G5306_p,
  G5307_p,
  G5308_p,
  G5309_p,
  G5310_p,
  G5311_p,
  G5312_n,
  G5313_n,
  G5314_p,
  G5315_p
);

  input G1_p;input G1_n;input G2_p;input G2_n;input G3_p;input G3_n;input G4_p;input G4_n;input G5_p;input G5_n;input G6_p;input G6_n;input G7_p;input G7_n;input G8_p;input G8_n;input G9_p;input G9_n;input G10_p;input G10_n;input G11_p;input G11_n;input G12_p;input G12_n;input G13_p;input G13_n;input G14_p;input G14_n;input G15_p;input G15_n;input G16_p;input G16_n;input G17_p;input G17_n;input G18_p;input G18_n;input G19_p;input G19_n;input G20_p;input G20_n;input G21_p;input G21_n;input G22_p;input G22_n;input G23_p;input G23_n;input G24_p;input G24_n;input G25_p;input G25_n;input G26_p;input G26_n;input G27_p;input G27_n;input G28_p;input G28_n;input G29_p;input G29_n;input G30_p;input G30_n;input G31_p;input G31_n;input G32_p;input G32_n;input G33_p;input G33_n;input G34_p;input G34_n;input G35_p;input G35_n;input G36_p;input G36_n;input G37_p;input G37_n;input G38_p;input G38_n;input G39_p;input G39_n;input G40_p;input G40_n;input G41_p;input G41_n;input G42_p;input G42_n;input G43_p;input G43_n;input G44_p;input G44_n;input G45_p;input G45_n;input G46_p;input G46_n;input G47_p;input G47_n;input G48_p;input G48_n;input G49_p;input G49_n;input G50_p;input G50_n;input G51_p;input G51_n;input G52_p;input G52_n;input G53_p;input G53_n;input G54_p;input G54_n;input G55_p;input G55_n;input G56_p;input G56_n;input G57_p;input G57_n;input G58_p;input G58_n;input G59_p;input G59_n;input G60_p;input G60_n;input G61_p;input G61_n;input G62_p;input G62_n;input G63_p;input G63_n;input G64_p;input G64_n;input G65_p;input G65_n;input G66_p;input G66_n;input G67_p;input G67_n;input G68_p;input G68_n;input G69_p;input G69_n;input G70_p;input G70_n;input G71_p;input G71_n;input G72_p;input G72_n;input G73_p;input G73_n;input G74_p;input G74_n;input G75_p;input G75_n;input G76_p;input G76_n;input G77_p;input G77_n;input G78_p;input G78_n;input G79_p;input G79_n;input G80_p;input G80_n;input G81_p;input G81_n;input G82_p;input G82_n;input G83_p;input G83_n;input G84_p;input G84_n;input G85_p;input G85_n;input G86_p;input G86_n;input G87_p;input G87_n;input G88_p;input G88_n;input G89_p;input G89_n;input G90_p;input G90_n;input G91_p;input G91_n;input G92_p;input G92_n;input G93_p;input G93_n;input G94_p;input G94_n;input G95_p;input G95_n;input G96_p;input G96_n;input G97_p;input G97_n;input G98_p;input G98_n;input G99_p;input G99_n;input G100_p;input G100_n;input G101_p;input G101_n;input G102_p;input G102_n;input G103_p;input G103_n;input G104_p;input G104_n;input G105_p;input G105_n;input G106_p;input G106_n;input G107_p;input G107_n;input G108_p;input G108_n;input G109_p;input G109_n;input G110_p;input G110_n;input G111_p;input G111_n;input G112_p;input G112_n;input G113_p;input G113_n;input G114_p;input G114_n;input G115_p;input G115_n;input G116_p;input G116_n;input G117_p;input G117_n;input G118_p;input G118_n;input G119_p;input G119_n;input G120_p;input G120_n;input G121_p;input G121_n;input G122_p;input G122_n;input G123_p;input G123_n;input G124_p;input G124_n;input G125_p;input G125_n;input G126_p;input G126_n;input G127_p;input G127_n;input G128_p;input G128_n;input G129_p;input G129_n;input G130_p;input G130_n;input G131_p;input G131_n;input G132_p;input G132_n;input G133_p;input G133_n;input G134_p;input G134_n;input G135_p;input G135_n;input G136_p;input G136_n;input G137_p;input G137_n;input G138_p;input G138_n;input G139_p;input G139_n;input G140_p;input G140_n;input G141_p;input G141_n;input G142_p;input G142_n;input G143_p;input G143_n;input G144_p;input G144_n;input G145_p;input G145_n;input G146_p;input G146_n;input G147_p;input G147_n;input G148_p;input G148_n;input G149_p;input G149_n;input G150_p;input G150_n;input G151_p;input G151_n;input G152_p;input G152_n;input G153_p;input G153_n;input G154_p;input G154_n;input G155_p;input G155_n;input G156_p;input G156_n;input G157_p;input G157_n;input G158_p;input G158_n;input G159_p;input G159_n;input G160_p;input G160_n;input G161_p;input G161_n;input G162_p;input G162_n;input G163_p;input G163_n;input G164_p;input G164_n;input G165_p;input G165_n;input G166_p;input G166_n;input G167_p;input G167_n;input G168_p;input G168_n;input G169_p;input G169_n;input G170_p;input G170_n;input G171_p;input G171_n;input G172_p;input G172_n;input G173_p;input G173_n;input G174_p;input G174_n;input G175_p;input G175_n;input G176_p;input G176_n;input G177_p;input G177_n;input G178_p;input G178_n;
  output G5193_p;output G5194_p;output G5195_p;output G5196_p;output G5197_p;output G5198_p;output G5199_n;output G5200_p;output G5201_p;output G5202_p;output G5203_p;output G5204_p;output G5205_p;output G5206_p;output G5207_p;output G5208_p;output G5209_p;output G5210_p;output G5211_p;output G5212_p;output G5213_p;output G5214_p;output G5215_p;output G5216_p;output G5217_p;output G5218_p;output G5219_p;output G5220_p;output G5221_p;output G5222_p;output G5223_p;output G5224_p;output G5225_p;output G5226_p;output G5227_p;output G5228_p;output G5229_p;output G5230_p;output G5231_p;output G5232_p;output G5233_p;output G5234_p;output G5235_p;output G5236_n;output G5237_n;output G5238_n;output G5239_p;output G5240_p;output G5241_n;output G5242_n;output G5243_n;output G5244_n;output G5245_p;output G5246_n;output G5247_p;output G5248_n;output G5249_n;output G5250_n;output G5251_p;output G5252_p;output G5253_n;output G5254_n;output G5255_n;output G5256_p;output G5257_n;output G5258_n;output G5259_n;output G5260_n;output G5261_n;output G5262_n;output G5263_n;output G5264_n;output G5265_p;output G5266_p;output G5267_p;output G5268_p;output G5269_p;output G5270_p;output G5271_p;output G5272_p;output G5273_p;output G5274_p;output G5275_p;output G5276_p;output G5277_p;output G5278_p;output G5279_p;output G5280_p;output G5281_p;output G5282_p;output G5283_p;output G5284_p;output G5285_n;output G5286_n;output G5287_n;output G5288_n;output G5289_n;output G5290_n;output G5291_n;output G5292_n;output G5293_n;output G5294_p;output G5295_p;output G5296_p;output G5297_p;output G5298_p;output G5299_p;output G5300_p;output G5301_p;output G5302_p;output G5303_p;output G5304_p;output G5305_p;output G5306_p;output G5307_p;output G5308_p;output G5309_p;output G5310_p;output G5311_p;output G5312_n;output G5313_n;output G5314_p;output G5315_p;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire G51_p;
  wire G51_n;
  wire G52_p;
  wire G52_n;
  wire G53_p;
  wire G53_n;
  wire G54_p;
  wire G54_n;
  wire G55_p;
  wire G55_n;
  wire G56_p;
  wire G56_n;
  wire G57_p;
  wire G57_n;
  wire G58_p;
  wire G58_n;
  wire G59_p;
  wire G59_n;
  wire G60_p;
  wire G60_n;
  wire G61_p;
  wire G61_n;
  wire G62_p;
  wire G62_n;
  wire G63_p;
  wire G63_n;
  wire G64_p;
  wire G64_n;
  wire G65_p;
  wire G65_n;
  wire G66_p;
  wire G66_n;
  wire G67_p;
  wire G67_n;
  wire G68_p;
  wire G68_n;
  wire G69_p;
  wire G69_n;
  wire G70_p;
  wire G70_n;
  wire G71_p;
  wire G71_n;
  wire G72_p;
  wire G72_n;
  wire G73_p;
  wire G73_n;
  wire G74_p;
  wire G74_n;
  wire G75_p;
  wire G75_n;
  wire G76_p;
  wire G76_n;
  wire G77_p;
  wire G77_n;
  wire G78_p;
  wire G78_n;
  wire G79_p;
  wire G79_n;
  wire G80_p;
  wire G80_n;
  wire G81_p;
  wire G81_n;
  wire G82_p;
  wire G82_n;
  wire G83_p;
  wire G83_n;
  wire G84_p;
  wire G84_n;
  wire G85_p;
  wire G85_n;
  wire G86_p;
  wire G86_n;
  wire G87_p;
  wire G87_n;
  wire G88_p;
  wire G88_n;
  wire G89_p;
  wire G89_n;
  wire G90_p;
  wire G90_n;
  wire G91_p;
  wire G91_n;
  wire G92_p;
  wire G92_n;
  wire G93_p;
  wire G93_n;
  wire G94_p;
  wire G94_n;
  wire G95_p;
  wire G95_n;
  wire G96_p;
  wire G96_n;
  wire G97_p;
  wire G97_n;
  wire G98_p;
  wire G98_n;
  wire G99_p;
  wire G99_n;
  wire G100_p;
  wire G100_n;
  wire G101_p;
  wire G101_n;
  wire G102_p;
  wire G102_n;
  wire G103_p;
  wire G103_n;
  wire G104_p;
  wire G104_n;
  wire G105_p;
  wire G105_n;
  wire G106_p;
  wire G106_n;
  wire G107_p;
  wire G107_n;
  wire G108_p;
  wire G108_n;
  wire G109_p;
  wire G109_n;
  wire G110_p;
  wire G110_n;
  wire G111_p;
  wire G111_n;
  wire G112_p;
  wire G112_n;
  wire G113_p;
  wire G113_n;
  wire G114_p;
  wire G114_n;
  wire G115_p;
  wire G115_n;
  wire G116_p;
  wire G116_n;
  wire G117_p;
  wire G117_n;
  wire G118_p;
  wire G118_n;
  wire G119_p;
  wire G119_n;
  wire G120_p;
  wire G120_n;
  wire G121_p;
  wire G121_n;
  wire G122_p;
  wire G122_n;
  wire G123_p;
  wire G123_n;
  wire G124_p;
  wire G124_n;
  wire G125_p;
  wire G125_n;
  wire G126_p;
  wire G126_n;
  wire G127_p;
  wire G127_n;
  wire G128_p;
  wire G128_n;
  wire G129_p;
  wire G129_n;
  wire G130_p;
  wire G130_n;
  wire G131_p;
  wire G131_n;
  wire G132_p;
  wire G132_n;
  wire G133_p;
  wire G133_n;
  wire G134_p;
  wire G134_n;
  wire G135_p;
  wire G135_n;
  wire G136_p;
  wire G136_n;
  wire G137_p;
  wire G137_n;
  wire G138_p;
  wire G138_n;
  wire G139_p;
  wire G139_n;
  wire G140_p;
  wire G140_n;
  wire G141_p;
  wire G141_n;
  wire G142_p;
  wire G142_n;
  wire G143_p;
  wire G143_n;
  wire G144_p;
  wire G144_n;
  wire G145_p;
  wire G145_n;
  wire G146_p;
  wire G146_n;
  wire G147_p;
  wire G147_n;
  wire G148_p;
  wire G148_n;
  wire G149_p;
  wire G149_n;
  wire G150_p;
  wire G150_n;
  wire G151_p;
  wire G151_n;
  wire G152_p;
  wire G152_n;
  wire G153_p;
  wire G153_n;
  wire G154_p;
  wire G154_n;
  wire G155_p;
  wire G155_n;
  wire G156_p;
  wire G156_n;
  wire G157_p;
  wire G157_n;
  wire G158_p;
  wire G158_n;
  wire G159_p;
  wire G159_n;
  wire G160_p;
  wire G160_n;
  wire G161_p;
  wire G161_n;
  wire G162_p;
  wire G162_n;
  wire G163_p;
  wire G163_n;
  wire G164_p;
  wire G164_n;
  wire G165_p;
  wire G165_n;
  wire G166_p;
  wire G166_n;
  wire G167_p;
  wire G167_n;
  wire G168_p;
  wire G168_n;
  wire G169_p;
  wire G169_n;
  wire G170_p;
  wire G170_n;
  wire G171_p;
  wire G171_n;
  wire G172_p;
  wire G172_n;
  wire G173_p;
  wire G173_n;
  wire G174_p;
  wire G174_n;
  wire G175_p;
  wire G175_n;
  wire G176_p;
  wire G176_n;
  wire G177_p;
  wire G177_n;
  wire G178_p;
  wire G178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire g686_p;
  wire g686_n;
  wire g687_p;
  wire g687_n;
  wire g688_p;
  wire g688_n;
  wire g689_p;
  wire g689_n;
  wire g690_p;
  wire g690_n;
  wire g691_p;
  wire g691_n;
  wire g692_p;
  wire g692_n;
  wire g693_p;
  wire g693_n;
  wire g694_p;
  wire g694_n;
  wire g695_p;
  wire g695_n;
  wire g696_p;
  wire g696_n;
  wire g697_p;
  wire g697_n;
  wire g698_p;
  wire g698_n;
  wire g699_p;
  wire g699_n;
  wire g700_p;
  wire g700_n;
  wire g701_p;
  wire g701_n;
  wire g702_p;
  wire g702_n;
  wire g703_p;
  wire g703_n;
  wire g704_p;
  wire g704_n;
  wire g705_p;
  wire g705_n;
  wire g706_p;
  wire g706_n;
  wire g707_p;
  wire g707_n;
  wire g708_p;
  wire g708_n;
  wire g709_p;
  wire g709_n;
  wire g710_p;
  wire g710_n;
  wire g711_p;
  wire g711_n;
  wire g712_p;
  wire g712_n;
  wire g713_p;
  wire g713_n;
  wire g714_p;
  wire g714_n;
  wire g715_p;
  wire g715_n;
  wire g716_p;
  wire g716_n;
  wire g717_p;
  wire g717_n;
  wire g718_p;
  wire g718_n;
  wire g719_p;
  wire g719_n;
  wire g720_p;
  wire g720_n;
  wire g721_p;
  wire g721_n;
  wire g722_p;
  wire g722_n;
  wire g723_p;
  wire g723_n;
  wire g724_p;
  wire g724_n;
  wire g725_p;
  wire g725_n;
  wire g726_p;
  wire g726_n;
  wire g727_p;
  wire g727_n;
  wire g728_p;
  wire g728_n;
  wire g729_p;
  wire g729_n;
  wire g730_p;
  wire g730_n;
  wire g731_p;
  wire g731_n;
  wire g732_p;
  wire g732_n;
  wire g733_p;
  wire g733_n;
  wire g734_p;
  wire g734_n;
  wire g735_p;
  wire g735_n;
  wire g736_p;
  wire g736_n;
  wire g737_p;
  wire g737_n;
  wire g738_p;
  wire g738_n;
  wire g739_p;
  wire g739_n;
  wire g740_p;
  wire g740_n;
  wire g741_p;
  wire g741_n;
  wire g742_p;
  wire g742_n;
  wire g743_p;
  wire g743_n;
  wire g744_p;
  wire g744_n;
  wire g745_p;
  wire g745_n;
  wire g746_p;
  wire g746_n;
  wire g747_p;
  wire g747_n;
  wire g748_p;
  wire g748_n;
  wire g749_p;
  wire g749_n;
  wire g750_p;
  wire g750_n;
  wire g751_p;
  wire g751_n;
  wire g752_p;
  wire g752_n;
  wire g753_p;
  wire g753_n;
  wire g754_p;
  wire g754_n;
  wire g755_p;
  wire g755_n;
  wire g756_p;
  wire g756_n;
  wire g757_p;
  wire g757_n;
  wire g758_p;
  wire g758_n;
  wire g759_p;
  wire g759_n;
  wire g760_p;
  wire g760_n;
  wire g761_p;
  wire g761_n;
  wire g762_p;
  wire g762_n;
  wire g763_p;
  wire g763_n;
  wire g764_p;
  wire g764_n;
  wire g765_p;
  wire g765_n;
  wire g766_p;
  wire g766_n;
  wire g767_p;
  wire g767_n;
  wire g768_p;
  wire g768_n;
  wire g769_p;
  wire g769_n;
  wire g770_p;
  wire g770_n;
  wire g771_p;
  wire g771_n;
  wire g772_p;
  wire g772_n;
  wire g773_p;
  wire g773_n;
  wire g774_p;
  wire g774_n;
  wire g775_p;
  wire g775_n;
  wire g776_p;
  wire g776_n;
  wire g777_p;
  wire g777_n;
  wire g778_p;
  wire g778_n;
  wire g779_p;
  wire g779_n;
  wire g780_p;
  wire g780_n;
  wire g781_p;
  wire g781_n;
  wire g782_p;
  wire g782_n;
  wire g783_p;
  wire g783_n;
  wire g784_p;
  wire g784_n;
  wire g785_p;
  wire g785_n;
  wire g786_p;
  wire g786_n;
  wire g787_p;
  wire g787_n;
  wire g788_p;
  wire g788_n;
  wire g789_p;
  wire g789_n;
  wire g790_p;
  wire g790_n;
  wire g791_p;
  wire g791_n;
  wire g792_p;
  wire g792_n;
  wire g793_p;
  wire g793_n;
  wire g794_p;
  wire g794_n;
  wire g795_p;
  wire g795_n;
  wire g796_p;
  wire g796_n;
  wire g797_p;
  wire g797_n;
  wire g798_p;
  wire g798_n;
  wire g799_p;
  wire g799_n;
  wire g800_p;
  wire g800_n;
  wire g801_p;
  wire g801_n;
  wire g802_p;
  wire g802_n;
  wire g803_p;
  wire g803_n;
  wire g804_p;
  wire g804_n;
  wire g805_p;
  wire g805_n;
  wire g806_p;
  wire g806_n;
  wire g807_p;
  wire g807_n;
  wire g808_p;
  wire g808_n;
  wire g809_p;
  wire g809_n;
  wire g810_p;
  wire g810_n;
  wire g811_p;
  wire g811_n;
  wire g812_p;
  wire g812_n;
  wire g813_p;
  wire g813_n;
  wire g814_p;
  wire g814_n;
  wire g815_p;
  wire g815_n;
  wire g816_p;
  wire g816_n;
  wire g817_p;
  wire g817_n;
  wire g818_p;
  wire g818_n;
  wire g819_p;
  wire g819_n;
  wire g820_p;
  wire g820_n;
  wire g821_p;
  wire g821_n;
  wire g822_p;
  wire g822_n;
  wire g823_p;
  wire g823_n;
  wire g824_p;
  wire g824_n;
  wire g825_p;
  wire g825_n;
  wire g826_p;
  wire g826_n;
  wire g827_p;
  wire g827_n;
  wire g828_p;
  wire g828_n;
  wire g829_p;
  wire g829_n;
  wire g830_p;
  wire g830_n;
  wire g831_p;
  wire g831_n;
  wire g832_p;
  wire g832_n;
  wire g833_p;
  wire g833_n;
  wire g834_p;
  wire g834_n;
  wire g835_p;
  wire g835_n;
  wire g836_p;
  wire g836_n;
  wire g837_p;
  wire g837_n;
  wire g838_p;
  wire g838_n;
  wire g839_p;
  wire g839_n;
  wire g840_p;
  wire g840_n;
  wire g841_p;
  wire g841_n;
  wire g842_p;
  wire g842_n;
  wire g843_p;
  wire g843_n;
  wire g844_p;
  wire g844_n;
  wire g845_p;
  wire g845_n;
  wire g846_p;
  wire g846_n;
  wire g847_p;
  wire g847_n;
  wire g848_p;
  wire g848_n;
  wire g849_p;
  wire g849_n;
  wire g850_p;
  wire g850_n;
  wire g851_p;
  wire g851_n;
  wire g852_p;
  wire g852_n;
  wire g853_p;
  wire g853_n;
  wire g854_p;
  wire g854_n;
  wire g855_p;
  wire g855_n;
  wire g856_p;
  wire g856_n;
  wire g857_p;
  wire g857_n;
  wire g858_p;
  wire g858_n;
  wire g859_p;
  wire g859_n;
  wire g860_p;
  wire g860_n;
  wire g861_p;
  wire g861_n;
  wire g862_p;
  wire g862_n;
  wire g863_p;
  wire g863_n;
  wire g864_p;
  wire g864_n;
  wire g865_p;
  wire g865_n;
  wire g866_p;
  wire g866_n;
  wire g867_p;
  wire g867_n;
  wire g868_p;
  wire g868_n;
  wire g869_p;
  wire g869_n;
  wire g870_p;
  wire g870_n;
  wire g871_p;
  wire g871_n;
  wire g872_p;
  wire g872_n;
  wire g873_p;
  wire g873_n;
  wire g874_p;
  wire g874_n;
  wire g875_p;
  wire g875_n;
  wire g876_p;
  wire g876_n;
  wire g877_p;
  wire g877_n;
  wire g878_p;
  wire g878_n;
  wire g879_p;
  wire g879_n;
  wire g880_p;
  wire g880_n;
  wire g881_p;
  wire g881_n;
  wire g882_p;
  wire g882_n;
  wire g883_p;
  wire g883_n;
  wire g884_p;
  wire g884_n;
  wire g885_p;
  wire g885_n;
  wire g886_p;
  wire g886_n;
  wire g887_p;
  wire g887_n;
  wire g888_p;
  wire g888_n;
  wire g889_p;
  wire g889_n;
  wire g890_p;
  wire g890_n;
  wire g891_p;
  wire g891_n;
  wire g892_p;
  wire g892_n;
  wire g893_p;
  wire g893_n;
  wire g894_p;
  wire g894_n;
  wire g895_p;
  wire g895_n;
  wire g896_p;
  wire g896_n;
  wire g897_p;
  wire g897_n;
  wire g898_p;
  wire g898_n;
  wire g899_p;
  wire g899_n;
  wire g900_p;
  wire g900_n;
  wire g901_p;
  wire g901_n;
  wire g902_p;
  wire g902_n;
  wire g903_p;
  wire g903_n;
  wire g904_p;
  wire g904_n;
  wire g905_p;
  wire g905_n;
  wire g906_p;
  wire g906_n;
  wire g907_p;
  wire g907_n;
  wire g908_p;
  wire g908_n;
  wire g909_p;
  wire g909_n;
  wire g910_p;
  wire g910_n;
  wire g911_p;
  wire g911_n;
  wire g912_p;
  wire g912_n;
  wire g913_p;
  wire g913_n;
  wire g914_p;
  wire g914_n;
  wire g915_p;
  wire g915_n;
  wire g916_p;
  wire g916_n;
  wire g917_p;
  wire g917_n;
  wire g918_p;
  wire g918_n;
  wire g919_p;
  wire g919_n;
  wire g920_p;
  wire g920_n;
  wire g921_p;
  wire g921_n;
  wire g922_p;
  wire g922_n;
  wire g923_p;
  wire g923_n;
  wire g924_p;
  wire g924_n;
  wire g925_p;
  wire g925_n;
  wire g926_p;
  wire g926_n;
  wire g927_p;
  wire g927_n;
  wire g928_p;
  wire g928_n;
  wire g929_p;
  wire g929_n;
  wire g930_p;
  wire g930_n;
  wire g931_p;
  wire g931_n;
  wire g932_p;
  wire g932_n;
  wire g933_p;
  wire g933_n;
  wire g934_p;
  wire g934_n;
  wire g935_p;
  wire g935_n;
  wire g936_p;
  wire g936_n;
  wire g937_p;
  wire g937_n;
  wire g938_p;
  wire g938_n;
  wire g939_p;
  wire g939_n;
  wire g940_p;
  wire g940_n;
  wire g941_p;
  wire g941_n;
  wire g942_p;
  wire g942_n;
  wire g943_p;
  wire g943_n;
  wire g944_p;
  wire g944_n;
  wire g945_p;
  wire g945_n;
  wire g946_p;
  wire g946_n;
  wire g947_p;
  wire g947_n;
  wire g948_p;
  wire g948_n;
  wire g949_p;
  wire g949_n;
  wire g950_p;
  wire g950_n;
  wire g951_p;
  wire g951_n;
  wire g952_p;
  wire g952_n;
  wire g953_p;
  wire g953_n;
  wire g954_p;
  wire g954_n;
  wire g955_p;
  wire g955_n;
  wire g956_p;
  wire g956_n;
  wire g957_p;
  wire g957_n;
  wire g958_p;
  wire g958_n;
  wire g959_p;
  wire g959_n;
  wire g960_p;
  wire g960_n;
  wire g961_p;
  wire g961_n;
  wire g962_p;
  wire g962_n;
  wire g963_p;
  wire g963_n;
  wire g964_p;
  wire g964_n;
  wire g965_p;
  wire g965_n;
  wire g966_p;
  wire g966_n;
  wire g967_p;
  wire g967_n;
  wire g968_p;
  wire g968_n;
  wire g969_p;
  wire g969_n;
  wire g970_p;
  wire g970_n;
  wire g971_p;
  wire g971_n;
  wire g972_p;
  wire g972_n;
  wire g973_p;
  wire g973_n;
  wire g974_p;
  wire g974_n;
  wire g975_p;
  wire g975_n;
  wire g976_p;
  wire g976_n;
  wire g977_p;
  wire g977_n;
  wire g978_p;
  wire g978_n;
  wire g979_p;
  wire g979_n;
  wire g980_p;
  wire g980_n;
  wire g981_p;
  wire g981_n;
  wire g982_p;
  wire g982_n;
  wire g983_p;
  wire g983_n;
  wire g984_p;
  wire g984_n;
  wire g985_p;
  wire g985_n;
  wire g986_p;
  wire g986_n;
  wire g987_p;
  wire g987_n;
  wire g988_p;
  wire g988_n;
  wire g989_p;
  wire g989_n;
  wire g990_p;
  wire g990_n;
  wire g991_p;
  wire g991_n;
  wire g992_p;
  wire g992_n;
  wire g993_p;
  wire g993_n;
  wire g994_p;
  wire g994_n;
  wire g995_p;
  wire g995_n;
  wire g996_p;
  wire g996_n;
  wire g997_p;
  wire g997_n;
  wire g998_p;
  wire g998_n;
  wire g999_p;
  wire g999_n;
  wire g1000_p;
  wire g1000_n;
  wire g1001_p;
  wire g1001_n;
  wire g1002_p;
  wire g1002_n;
  wire g1003_p;
  wire g1003_n;
  wire g1004_p;
  wire g1004_n;
  wire g1005_p;
  wire g1005_n;
  wire g1006_p;
  wire g1006_n;
  wire g1007_p;
  wire g1007_n;
  wire g1008_p;
  wire g1008_n;
  wire g1009_p;
  wire g1009_n;
  wire g1010_p;
  wire g1010_n;
  wire g1011_p;
  wire g1011_n;
  wire g1012_p;
  wire g1012_n;
  wire g1013_p;
  wire g1013_n;
  wire g1014_p;
  wire g1014_n;
  wire g1015_p;
  wire g1015_n;
  wire g1016_p;
  wire g1016_n;
  wire g1017_p;
  wire g1017_n;
  wire g1018_p;
  wire g1018_n;
  wire g1019_p;
  wire g1019_n;
  wire g1020_p;
  wire g1020_n;
  wire g1021_p;
  wire g1021_n;
  wire g1022_p;
  wire g1022_n;
  wire g1023_p;
  wire g1023_n;
  wire g1024_p;
  wire g1024_n;
  wire g1025_p;
  wire g1025_n;
  wire g1026_p;
  wire g1026_n;
  wire g1027_p;
  wire g1027_n;
  wire g1028_p;
  wire g1028_n;
  wire g1029_p;
  wire g1029_n;
  wire g1030_p;
  wire g1030_n;
  wire g1031_p;
  wire g1031_n;
  wire g1032_p;
  wire g1032_n;
  wire g1033_p;
  wire g1033_n;
  wire g1034_p;
  wire g1034_n;
  wire g1035_p;
  wire g1035_n;
  wire g1036_p;
  wire g1036_n;
  wire g1037_p;
  wire g1037_n;
  wire g1038_p;
  wire g1038_n;
  wire g1039_p;
  wire g1039_n;
  wire g1040_p;
  wire g1040_n;
  wire g1041_p;
  wire g1041_n;
  wire g1042_p;
  wire g1042_n;
  wire g1043_p;
  wire g1043_n;
  wire g1044_p;
  wire g1044_n;
  wire g1045_p;
  wire g1045_n;
  wire g1046_p;
  wire g1046_n;
  wire g1047_p;
  wire g1047_n;
  wire g1048_p;
  wire g1048_n;
  wire g1049_p;
  wire g1049_n;
  wire g1050_p;
  wire g1050_n;
  wire g1051_p;
  wire g1051_n;
  wire g1052_p;
  wire g1052_n;
  wire g1053_p;
  wire g1053_n;
  wire g1054_p;
  wire g1054_n;
  wire g1055_p;
  wire g1055_n;
  wire g1056_p;
  wire g1056_n;
  wire g1057_p;
  wire g1057_n;
  wire g1058_p;
  wire g1058_n;
  wire g1059_p;
  wire g1059_n;
  wire g1060_p;
  wire g1060_n;
  wire g1061_p;
  wire g1061_n;
  wire g1062_p;
  wire g1062_n;
  wire g1063_p;
  wire g1063_n;
  wire g1064_p;
  wire g1064_n;
  wire g1065_p;
  wire g1065_n;
  wire g1066_p;
  wire g1066_n;
  wire g1067_p;
  wire g1067_n;
  wire g1068_p;
  wire g1068_n;
  wire g1069_p;
  wire g1069_n;
  wire g1070_p;
  wire g1070_n;
  wire g1071_p;
  wire g1071_n;
  wire g1072_p;
  wire g1072_n;
  wire g1073_p;
  wire g1073_n;
  wire g1074_p;
  wire g1074_n;
  wire g1075_p;
  wire g1075_n;
  wire g1076_p;
  wire g1076_n;
  wire g1077_p;
  wire g1077_n;
  wire g1078_p;
  wire g1078_n;
  wire g1079_p;
  wire g1079_n;
  wire g1080_p;
  wire g1080_n;
  wire g1081_p;
  wire g1081_n;
  wire g1082_p;
  wire g1082_n;
  wire g1083_p;
  wire g1083_n;
  wire g1084_p;
  wire g1084_n;
  wire g1085_p;
  wire g1085_n;
  wire g1086_p;
  wire g1086_n;
  wire g1087_p;
  wire g1087_n;
  wire g1088_p;
  wire g1088_n;
  wire g1089_p;
  wire g1089_n;
  wire g1090_p;
  wire g1090_n;
  wire g1091_p;
  wire g1091_n;
  wire g1092_p;
  wire g1092_n;
  wire g1093_p;
  wire g1093_n;
  wire g1094_p;
  wire g1094_n;
  wire g1095_p;
  wire g1095_n;
  wire g1096_p;
  wire g1096_n;
  wire g1097_p;
  wire g1097_n;
  wire g1098_p;
  wire g1098_n;
  wire g1099_p;
  wire g1099_n;
  wire g1100_p;
  wire g1100_n;
  wire g1101_p;
  wire g1101_n;
  wire g1102_p;
  wire g1102_n;
  wire g1103_p;
  wire g1103_n;
  wire g1104_p;
  wire g1104_n;
  wire g1105_p;
  wire g1105_n;
  wire g1106_p;
  wire g1106_n;
  wire g1107_p;
  wire g1107_n;
  wire g1108_p;
  wire g1108_n;
  wire g1109_p;
  wire g1109_n;
  wire g1110_p;
  wire g1110_n;
  wire g1111_p;
  wire g1111_n;
  wire g1112_p;
  wire g1112_n;
  wire g1113_p;
  wire g1113_n;
  wire g1114_p;
  wire g1114_n;
  wire g1115_p;
  wire g1115_n;
  wire g1116_p;
  wire g1116_n;
  wire g1117_p;
  wire g1117_n;
  wire g1118_p;
  wire g1118_n;
  wire g1119_p;
  wire g1119_n;
  wire g1120_p;
  wire g1120_n;
  wire g1121_p;
  wire g1121_n;
  wire g1122_p;
  wire g1122_n;
  wire g1123_p;
  wire g1123_n;
  wire g1124_p;
  wire g1124_n;
  wire g1125_p;
  wire g1125_n;
  wire g1126_p;
  wire g1126_n;
  wire g1127_p;
  wire g1127_n;
  wire g1128_p;
  wire g1128_n;
  wire g1129_p;
  wire g1129_n;
  wire g1130_p;
  wire g1130_n;
  wire g1131_p;
  wire g1131_n;
  wire g1132_p;
  wire g1132_n;
  wire g1133_p;
  wire g1133_n;
  wire g1134_p;
  wire g1134_n;
  wire g1135_p;
  wire g1135_n;
  wire g1136_p;
  wire g1136_n;
  wire g1137_p;
  wire g1137_n;
  wire g1138_p;
  wire g1138_n;
  wire g1139_p;
  wire g1139_n;
  wire g1140_p;
  wire g1140_n;
  wire g1141_p;
  wire g1141_n;
  wire g1142_p;
  wire g1142_n;
  wire g1143_p;
  wire g1143_n;
  wire g1144_p;
  wire g1144_n;
  wire g1145_p;
  wire g1145_n;
  wire g1146_p;
  wire g1146_n;
  wire g1147_p;
  wire g1147_n;
  wire g1148_p;
  wire g1148_n;
  wire g1149_p;
  wire g1149_n;
  wire g1150_p;
  wire g1150_n;
  wire g1151_p;
  wire g1151_n;
  wire g1152_p;
  wire g1152_n;
  wire g1153_p;
  wire g1153_n;
  wire g1154_p;
  wire g1154_n;
  wire g1155_p;
  wire g1155_n;
  wire g1156_p;
  wire g1156_n;
  wire g1157_p;
  wire g1157_n;
  wire g1158_p;
  wire g1158_n;
  wire g1159_p;
  wire g1159_n;
  wire g1160_p;
  wire g1160_n;
  wire g1161_p;
  wire g1161_n;
  wire g1162_p;
  wire g1162_n;
  wire g1163_p;
  wire g1163_n;
  wire g1164_p;
  wire g1164_n;
  wire g1165_p;
  wire g1165_n;
  wire g1166_p;
  wire g1166_n;
  wire g1167_p;
  wire g1167_n;
  wire g1168_p;
  wire g1168_n;
  wire g1169_p;
  wire g1169_n;
  wire g1170_p;
  wire g1170_n;
  wire g1171_p;
  wire g1171_n;
  wire g1172_p;
  wire g1172_n;
  wire g1173_p;
  wire g1173_n;
  wire g1174_p;
  wire g1174_n;
  wire g1175_p;
  wire g1175_n;
  wire g1176_p;
  wire g1176_n;
  wire g1177_p;
  wire g1177_n;
  wire g1178_p;
  wire g1178_n;
  wire g1179_p;
  wire g1179_n;
  wire g1180_p;
  wire g1180_n;
  wire g1181_p;
  wire g1181_n;
  wire g1182_p;
  wire g1182_n;
  wire g1183_p;
  wire g1183_n;
  wire g1184_p;
  wire g1184_n;
  wire g1185_p;
  wire g1185_n;
  wire g1186_p;
  wire g1186_n;
  wire g1187_p;
  wire g1187_n;
  wire g1188_p;
  wire g1188_n;
  wire g1189_p;
  wire g1189_n;
  wire g1190_p;
  wire g1190_n;
  wire g1191_p;
  wire g1191_n;
  wire g1192_p;
  wire g1192_n;
  wire g1193_p;
  wire g1193_n;
  wire g1194_p;
  wire g1194_n;
  wire g1195_p;
  wire g1195_n;
  wire g1196_p;
  wire g1196_n;
  wire g1197_p;
  wire g1197_n;
  wire g1198_p;
  wire g1198_n;
  wire g1199_p;
  wire g1199_n;
  wire g1200_p;
  wire g1200_n;
  wire g1201_p;
  wire g1201_n;
  wire g1202_p;
  wire g1202_n;
  wire g1203_p;
  wire g1203_n;
  wire g1204_p;
  wire g1204_n;
  wire g1205_p;
  wire g1205_n;
  wire g1206_p;
  wire g1206_n;
  wire g1207_p;
  wire g1207_n;
  wire g1208_p;
  wire g1208_n;
  wire g1209_p;
  wire g1209_n;
  wire g1210_p;
  wire g1210_n;
  wire g1211_p;
  wire g1211_n;
  wire g1212_p;
  wire g1212_n;
  wire g1213_p;
  wire g1213_n;
  wire g1214_p;
  wire g1214_n;
  wire g1215_p;
  wire g1215_n;
  wire g1216_p;
  wire g1216_n;
  wire g1217_p;
  wire g1217_n;
  wire g1218_p;
  wire g1218_n;
  wire g1219_p;
  wire g1219_n;
  wire g1220_p;
  wire g1220_n;
  wire g1221_p;
  wire g1221_n;
  wire g1222_p;
  wire g1222_n;
  wire g1223_p;
  wire g1223_n;
  wire g1224_p;
  wire g1224_n;
  wire g1225_p;
  wire g1225_n;
  wire g1226_p;
  wire g1226_n;
  wire g1227_p;
  wire g1227_n;
  wire g1228_p;
  wire g1228_n;
  wire g1229_p;
  wire g1229_n;
  wire g1230_p;
  wire g1230_n;
  wire g1231_p;
  wire g1231_n;
  wire g1232_p;
  wire g1232_n;
  wire g1233_p;
  wire g1233_n;
  wire g1234_p;
  wire g1234_n;
  wire g1235_p;
  wire g1235_n;
  wire g1236_p;
  wire g1236_n;
  wire g1237_p;
  wire g1237_n;
  wire g1238_p;
  wire g1238_n;
  wire g1239_p;
  wire g1239_n;
  wire g1240_p;
  wire g1240_n;
  wire g1241_p;
  wire g1241_n;
  wire g1242_p;
  wire g1242_n;
  wire g1243_p;
  wire g1243_n;
  wire g1244_p;
  wire g1244_n;
  wire g1245_p;
  wire g1245_n;
  wire g1246_p;
  wire g1246_n;
  wire g1247_p;
  wire g1247_n;
  wire g1248_p;
  wire g1248_n;
  wire g1249_p;
  wire g1249_n;
  wire g1250_p;
  wire g1250_n;
  wire g1251_p;
  wire g1251_n;
  wire g1252_p;
  wire g1252_n;
  wire g1253_p;
  wire g1253_n;
  wire g1254_p;
  wire g1254_n;
  wire g1255_p;
  wire g1255_n;
  wire g1256_p;
  wire g1256_n;
  wire g1257_p;
  wire g1257_n;
  wire g1258_p;
  wire g1258_n;
  wire g1259_p;
  wire g1259_n;
  wire g1260_p;
  wire g1260_n;
  wire g1261_p;
  wire g1261_n;
  wire g1262_p;
  wire g1262_n;
  wire g1263_p;
  wire g1263_n;
  wire g1264_p;
  wire g1264_n;
  wire g1265_p;
  wire g1265_n;
  wire g1266_p;
  wire g1266_n;
  wire g1267_p;
  wire g1267_n;
  wire g1268_p;
  wire g1268_n;
  wire g1269_p;
  wire g1269_n;
  wire g1270_p;
  wire g1270_n;
  wire g1271_p;
  wire g1271_n;
  wire g1272_p;
  wire g1272_n;
  wire g1273_p;
  wire g1273_n;
  wire g1274_p;
  wire g1274_n;
  wire g1275_p;
  wire g1275_n;
  wire g1276_p;
  wire g1276_n;
  wire g1277_p;
  wire g1277_n;
  wire g1278_p;
  wire g1278_n;
  wire g1279_p;
  wire g1279_n;
  wire g1280_p;
  wire g1280_n;
  wire g1281_p;
  wire g1281_n;
  wire g1282_p;
  wire g1282_n;
  wire g1283_p;
  wire g1283_n;
  wire g1284_p;
  wire g1284_n;
  wire g1285_p;
  wire g1285_n;
  wire g1286_p;
  wire g1286_n;
  wire g1287_p;
  wire g1287_n;
  wire g1288_p;
  wire g1288_n;
  wire g1289_p;
  wire g1289_n;
  wire g1290_p;
  wire g1290_n;
  wire g1291_p;
  wire g1291_n;
  wire g1292_p;
  wire g1292_n;
  wire g1293_p;
  wire g1293_n;
  wire g1294_p;
  wire g1294_n;
  wire g1295_p;
  wire g1295_n;
  wire g1296_p;
  wire g1296_n;
  wire g1297_p;
  wire g1297_n;
  wire g1298_p;
  wire g1298_n;
  wire g1299_p;
  wire g1299_n;
  wire g1300_p;
  wire g1300_n;
  wire g1301_p;
  wire g1301_n;
  wire g1302_p;
  wire g1302_n;
  wire g1303_p;
  wire g1303_n;
  wire g1304_p;
  wire g1304_n;
  wire g1305_p;
  wire g1305_n;
  wire g1306_p;
  wire g1306_n;
  wire g1307_p;
  wire g1307_n;
  wire g1308_p;
  wire g1308_n;
  wire g1309_p;
  wire g1309_n;
  wire g1310_p;
  wire g1310_n;
  wire g1311_p;
  wire g1311_n;
  wire g1312_p;
  wire g1312_n;
  wire g1313_p;
  wire g1313_n;
  wire g1314_p;
  wire g1314_n;
  wire g1315_p;
  wire g1315_n;
  wire g1316_p;
  wire g1316_n;
  wire g1317_p;
  wire g1317_n;
  wire g1318_p;
  wire g1318_n;
  wire g1319_p;
  wire g1319_n;
  wire g1320_p;
  wire g1320_n;
  wire g1321_p;
  wire g1321_n;
  wire g1322_p;
  wire g1322_n;
  wire g1323_p;
  wire g1323_n;
  wire g1324_p;
  wire g1324_n;
  wire g1325_p;
  wire g1325_n;
  wire g1326_p;
  wire g1326_n;
  wire g1327_p;
  wire g1327_n;
  wire g1328_p;
  wire g1328_n;
  wire g1329_p;
  wire g1329_n;
  wire g1330_p;
  wire g1330_n;
  wire g1331_p;
  wire g1331_n;
  wire g1332_p;
  wire g1332_n;
  wire g1333_p;
  wire g1333_n;
  wire g1334_p;
  wire g1334_n;
  wire g1335_p;
  wire g1335_n;
  wire g1336_p;
  wire g1336_n;
  wire g1337_p;
  wire g1337_n;
  wire g1338_p;
  wire g1338_n;
  wire g1339_p;
  wire g1339_n;
  wire g1340_p;
  wire g1340_n;
  wire g1341_p;
  wire g1341_n;
  wire g1342_p;
  wire g1342_n;
  wire g1343_p;
  wire g1343_n;
  wire g1344_p;
  wire g1344_n;
  wire g1345_p;
  wire g1345_n;
  wire g1346_p;
  wire g1346_n;
  wire g1347_p;
  wire g1347_n;
  wire g1348_p;
  wire g1348_n;
  wire g1349_p;
  wire g1349_n;
  wire g1350_p;
  wire g1350_n;
  wire g1351_p;
  wire g1351_n;
  wire g1352_p;
  wire g1352_n;
  wire g1353_p;
  wire g1353_n;
  wire g1354_p;
  wire g1354_n;
  wire g1355_p;
  wire g1355_n;
  wire g1356_p;
  wire g1356_n;
  wire g1357_p;
  wire g1357_n;
  wire g1358_p;
  wire g1358_n;
  wire g1359_p;
  wire g1359_n;
  wire g1360_p;
  wire g1360_n;
  wire g1361_p;
  wire g1361_n;
  wire g1362_p;
  wire g1362_n;
  wire g1363_p;
  wire g1363_n;
  wire g1364_p;
  wire g1364_n;
  wire g1365_p;
  wire g1365_n;
  wire g1366_p;
  wire g1366_n;
  wire g1367_p;
  wire g1367_n;
  wire g1368_p;
  wire g1368_n;
  wire g1369_p;
  wire g1369_n;
  wire g1370_p;
  wire g1370_n;
  wire g1371_p;
  wire g1371_n;
  wire g1372_p;
  wire g1372_n;
  wire g1373_p;
  wire g1373_n;
  wire g1374_p;
  wire g1374_n;
  wire g1375_p;
  wire g1375_n;
  wire g1376_p;
  wire g1376_n;
  wire g1377_p;
  wire g1377_n;
  wire g1378_p;
  wire g1378_n;
  wire g1379_p;
  wire g1379_n;
  wire g1380_p;
  wire g1380_n;
  wire g1381_p;
  wire g1381_n;
  wire g1382_p;
  wire g1382_n;
  wire g1383_p;
  wire g1383_n;
  wire g1384_p;
  wire g1384_n;
  wire g1385_p;
  wire g1385_n;
  wire g1386_p;
  wire g1386_n;
  wire g1387_p;
  wire g1387_n;
  wire g1388_p;
  wire g1388_n;
  wire g1389_p;
  wire g1389_n;
  wire g1390_p;
  wire g1390_n;
  wire g1391_p;
  wire g1391_n;
  wire g1392_p;
  wire g1392_n;
  wire g1393_p;
  wire g1393_n;
  wire g1394_p;
  wire g1394_n;
  wire g1395_p;
  wire g1395_n;
  wire g1396_p;
  wire g1396_n;
  wire g1397_p;
  wire g1397_n;
  wire g1398_p;
  wire g1398_n;
  wire g1399_p;
  wire g1399_n;
  wire g1400_p;
  wire g1400_n;
  wire g1401_p;
  wire g1401_n;
  wire g1402_p;
  wire g1402_n;
  wire g1403_p;
  wire g1403_n;
  wire g1404_p;
  wire g1404_n;
  wire g1405_p;
  wire g1405_n;
  wire g1406_p;
  wire g1406_n;
  wire g1407_p;
  wire g1407_n;
  wire g1408_p;
  wire g1408_n;
  wire g1409_p;
  wire g1409_n;
  wire g1410_p;
  wire g1410_n;
  wire g1411_p;
  wire g1411_n;
  wire g1412_p;
  wire g1412_n;
  wire g1413_p;
  wire g1413_n;
  wire g1414_p;
  wire g1414_n;
  wire g1415_p;
  wire g1415_n;
  wire g1416_p;
  wire g1416_n;
  wire g1417_p;
  wire g1417_n;
  wire g1418_p;
  wire g1418_n;
  wire g1419_p;
  wire g1419_n;
  wire g1420_p;
  wire g1420_n;
  wire g1421_p;
  wire g1421_n;
  wire g1422_p;
  wire g1422_n;
  wire g1423_p;
  wire g1423_n;
  wire g1424_p;
  wire g1424_n;
  wire g1425_p;
  wire g1425_n;
  wire g1426_p;
  wire g1426_n;
  wire g1427_p;
  wire g1427_n;
  wire g1428_p;
  wire g1428_n;
  wire g1429_p;
  wire g1429_n;
  wire g1430_p;
  wire g1430_n;
  wire g1431_p;
  wire g1431_n;
  wire g1432_p;
  wire g1432_n;
  wire g1433_p;
  wire g1433_n;
  wire g1434_p;
  wire g1434_n;
  wire g1435_p;
  wire g1435_n;
  wire g1436_p;
  wire g1436_n;
  wire g1437_p;
  wire g1437_n;
  wire g1438_p;
  wire g1438_n;
  wire g1439_p;
  wire g1439_n;
  wire g1440_p;
  wire g1440_n;
  wire g1441_p;
  wire g1441_n;
  wire g1442_p;
  wire g1442_n;
  wire g1443_p;
  wire g1443_n;
  wire g1444_p;
  wire g1444_n;
  wire g1445_p;
  wire g1445_n;
  wire g1446_p;
  wire g1446_n;
  wire g1447_p;
  wire g1447_n;
  wire g1448_p;
  wire g1448_n;
  wire g1449_p;
  wire g1449_n;
  wire g1450_p;
  wire g1450_n;
  wire g1451_p;
  wire g1451_n;
  wire g1452_p;
  wire g1452_n;
  wire g1453_p;
  wire g1453_n;
  wire g1454_p;
  wire g1454_n;
  wire g1455_p;
  wire g1455_n;
  wire g1456_p;
  wire g1456_n;
  wire g1457_p;
  wire g1457_n;
  wire g1458_p;
  wire g1458_n;
  wire g1459_p;
  wire g1459_n;
  wire g1460_p;
  wire g1460_n;
  wire g1461_p;
  wire g1461_n;
  wire g1462_p;
  wire g1462_n;
  wire g1463_p;
  wire g1463_n;
  wire g1464_p;
  wire g1464_n;
  wire g1465_p;
  wire g1465_n;
  wire g1466_p;
  wire g1466_n;
  wire g1467_p;
  wire g1467_n;
  wire g1468_p;
  wire g1468_n;
  wire g1469_p;
  wire g1469_n;
  wire g1470_p;
  wire g1470_n;
  wire g1471_p;
  wire g1471_n;
  wire g1472_p;
  wire g1472_n;
  wire g1473_p;
  wire g1473_n;
  wire g1474_p;
  wire g1474_n;
  wire g1475_p;
  wire g1475_n;
  wire g1476_p;
  wire g1476_n;
  wire g1477_p;
  wire g1477_n;
  wire g1478_p;
  wire g1478_n;
  wire g1479_p;
  wire g1479_n;
  wire g1480_p;
  wire g1480_n;
  wire g1481_p;
  wire g1481_n;
  wire g1482_p;
  wire g1482_n;
  wire g1483_p;
  wire g1483_n;
  wire g1484_p;
  wire g1484_n;
  wire g1485_p;
  wire g1485_n;
  wire g1486_p;
  wire g1486_n;
  wire g1487_p;
  wire g1487_n;
  wire g1488_p;
  wire g1488_n;
  wire g1489_p;
  wire g1489_n;
  wire g1490_p;
  wire g1490_n;
  wire g1491_p;
  wire g1491_n;
  wire g1492_p;
  wire g1492_n;
  wire g1493_p;
  wire g1493_n;
  wire g1494_p;
  wire g1494_n;
  wire g1495_p;
  wire g1495_n;
  wire g1496_p;
  wire g1496_n;
  wire g1497_p;
  wire g1497_n;
  wire g1498_p;
  wire g1498_n;
  wire g1499_p;
  wire g1499_n;
  wire g1500_p;
  wire g1500_n;
  wire g1501_p;
  wire g1501_n;
  wire g1502_p;
  wire g1502_n;
  wire g1503_p;
  wire g1503_n;
  wire g1504_p;
  wire g1504_n;
  wire g1505_p;
  wire g1505_n;
  wire g1506_p;
  wire g1506_n;
  wire g1507_p;
  wire g1507_n;
  wire g1508_p;
  wire g1508_n;
  wire g1509_p;
  wire g1509_n;
  wire g1510_p;
  wire g1510_n;
  wire g1511_p;
  wire g1511_n;
  wire g1512_p;
  wire g1512_n;
  wire g1513_p;
  wire g1513_n;
  wire g1514_p;
  wire g1514_n;
  wire g1515_p;
  wire g1515_n;
  wire g1516_p;
  wire g1516_n;
  wire g1517_p;
  wire g1517_n;
  wire g1518_p;
  wire g1518_n;
  wire g1519_p;
  wire g1519_n;
  wire g1520_p;
  wire g1520_n;
  wire g1521_p;
  wire g1521_n;
  wire g1522_p;
  wire g1522_n;
  wire g1523_p;
  wire g1523_n;
  wire g1524_p;
  wire g1524_n;
  wire g1525_p;
  wire g1525_n;
  wire g1526_p;
  wire g1526_n;
  wire g1527_p;
  wire g1527_n;
  wire g1528_p;
  wire g1528_n;
  wire g1529_p;
  wire g1529_n;
  wire g1530_p;
  wire g1530_n;
  wire g1531_p;
  wire g1531_n;
  wire g1532_p;
  wire g1532_n;
  wire g1533_p;
  wire g1533_n;
  wire g1534_p;
  wire g1534_n;
  wire g1535_p;
  wire g1535_n;
  wire g1536_p;
  wire g1536_n;
  wire g1537_p;
  wire g1537_n;
  wire g1538_p;
  wire g1538_n;
  wire g1539_p;
  wire g1539_n;
  wire g1540_p;
  wire g1540_n;
  wire g1541_p;
  wire g1541_n;
  wire g1542_p;
  wire g1542_n;
  wire g1543_p;
  wire g1543_n;
  wire g1544_p;
  wire g1544_n;
  wire g1545_p;
  wire g1545_n;
  wire G153_n_spl_;
  wire G156_n_spl_;
  wire G66_p_spl_;
  wire G66_p_spl_0;
  wire G66_p_spl_00;
  wire G66_p_spl_01;
  wire G66_p_spl_1;
  wire G1_p_spl_;
  wire G165_n_spl_;
  wire G11_n_spl_;
  wire g185_n_spl_;
  wire g185_n_spl_0;
  wire g185_n_spl_00;
  wire g185_n_spl_000;
  wire g185_n_spl_01;
  wire g185_n_spl_1;
  wire g185_n_spl_10;
  wire g185_n_spl_11;
  wire G163_n_spl_;
  wire G163_n_spl_0;
  wire G163_n_spl_00;
  wire G163_n_spl_01;
  wire G163_n_spl_1;
  wire G163_p_spl_;
  wire G163_p_spl_0;
  wire G163_p_spl_00;
  wire G163_p_spl_01;
  wire G163_p_spl_1;
  wire G128_p_spl_;
  wire G128_p_spl_0;
  wire G128_p_spl_00;
  wire G128_p_spl_000;
  wire G128_p_spl_01;
  wire G128_p_spl_1;
  wire G128_p_spl_10;
  wire G128_p_spl_11;
  wire G168_p_spl_;
  wire G168_p_spl_0;
  wire G168_p_spl_00;
  wire G168_p_spl_000;
  wire G168_p_spl_001;
  wire G168_p_spl_01;
  wire G168_p_spl_010;
  wire G168_p_spl_1;
  wire G168_p_spl_10;
  wire G168_p_spl_11;
  wire G128_n_spl_;
  wire G128_n_spl_0;
  wire G128_n_spl_00;
  wire G128_n_spl_000;
  wire G128_n_spl_01;
  wire G128_n_spl_1;
  wire G128_n_spl_10;
  wire G128_n_spl_11;
  wire G169_p_spl_;
  wire G169_p_spl_0;
  wire G169_p_spl_00;
  wire G169_p_spl_000;
  wire G169_p_spl_001;
  wire G169_p_spl_01;
  wire G169_p_spl_010;
  wire G169_p_spl_011;
  wire G169_p_spl_1;
  wire G169_p_spl_10;
  wire G169_p_spl_11;
  wire G150_p_spl_;
  wire G150_p_spl_0;
  wire G150_p_spl_00;
  wire G150_p_spl_1;
  wire G167_n_spl_;
  wire G167_n_spl_0;
  wire G167_n_spl_00;
  wire G167_n_spl_000;
  wire G167_n_spl_001;
  wire G167_n_spl_01;
  wire G167_n_spl_010;
  wire G167_n_spl_1;
  wire G167_n_spl_10;
  wire G167_n_spl_11;
  wire G166_n_spl_;
  wire G166_n_spl_0;
  wire G166_n_spl_00;
  wire G166_n_spl_000;
  wire G166_n_spl_001;
  wire G166_n_spl_01;
  wire G166_n_spl_010;
  wire G166_n_spl_011;
  wire G166_n_spl_1;
  wire G166_n_spl_10;
  wire G166_n_spl_11;
  wire G150_n_spl_;
  wire G150_n_spl_0;
  wire G150_n_spl_00;
  wire G150_n_spl_1;
  wire G126_p_spl_;
  wire G126_p_spl_0;
  wire G126_p_spl_00;
  wire G126_p_spl_000;
  wire G126_p_spl_01;
  wire G126_p_spl_1;
  wire G126_p_spl_10;
  wire G126_p_spl_11;
  wire G126_n_spl_;
  wire G126_n_spl_0;
  wire G126_n_spl_00;
  wire G126_n_spl_000;
  wire G126_n_spl_01;
  wire G126_n_spl_1;
  wire G126_n_spl_10;
  wire G126_n_spl_11;
  wire G149_p_spl_;
  wire G149_p_spl_0;
  wire G149_p_spl_00;
  wire G149_p_spl_1;
  wire G149_n_spl_;
  wire G149_n_spl_0;
  wire G149_n_spl_00;
  wire G149_n_spl_1;
  wire g224_n_spl_;
  wire g233_n_spl_;
  wire G102_p_spl_;
  wire G102_p_spl_0;
  wire G102_p_spl_00;
  wire G102_p_spl_000;
  wire G102_p_spl_001;
  wire G102_p_spl_01;
  wire G102_p_spl_010;
  wire G102_p_spl_011;
  wire G102_p_spl_1;
  wire G102_p_spl_10;
  wire G102_p_spl_100;
  wire G102_p_spl_101;
  wire G102_p_spl_11;
  wire G102_p_spl_110;
  wire G113_p_spl_;
  wire G113_p_spl_0;
  wire G113_p_spl_00;
  wire G113_p_spl_1;
  wire G102_n_spl_;
  wire G102_n_spl_0;
  wire G102_n_spl_00;
  wire G102_n_spl_000;
  wire G102_n_spl_001;
  wire G102_n_spl_01;
  wire G102_n_spl_010;
  wire G102_n_spl_011;
  wire G102_n_spl_1;
  wire G102_n_spl_10;
  wire G102_n_spl_100;
  wire G102_n_spl_101;
  wire G102_n_spl_11;
  wire G102_n_spl_110;
  wire G113_n_spl_;
  wire G113_n_spl_0;
  wire G113_n_spl_00;
  wire G113_n_spl_01;
  wire G113_n_spl_1;
  wire G98_p_spl_;
  wire G98_p_spl_0;
  wire G98_p_spl_00;
  wire G98_p_spl_000;
  wire G98_p_spl_001;
  wire G98_p_spl_01;
  wire G98_p_spl_010;
  wire G98_p_spl_011;
  wire G98_p_spl_1;
  wire G98_p_spl_10;
  wire G98_p_spl_100;
  wire G98_p_spl_101;
  wire G98_p_spl_11;
  wire G98_p_spl_110;
  wire G98_p_spl_111;
  wire G98_n_spl_;
  wire G98_n_spl_0;
  wire G98_n_spl_00;
  wire G98_n_spl_000;
  wire G98_n_spl_001;
  wire G98_n_spl_01;
  wire G98_n_spl_010;
  wire G98_n_spl_011;
  wire G98_n_spl_1;
  wire G98_n_spl_10;
  wire G98_n_spl_100;
  wire G98_n_spl_101;
  wire G98_n_spl_11;
  wire G98_n_spl_110;
  wire G98_n_spl_111;
  wire G101_p_spl_;
  wire G101_p_spl_0;
  wire G101_p_spl_00;
  wire G101_p_spl_000;
  wire G101_p_spl_001;
  wire G101_p_spl_01;
  wire G101_p_spl_010;
  wire G101_p_spl_011;
  wire G101_p_spl_1;
  wire G101_p_spl_10;
  wire G101_p_spl_100;
  wire G101_p_spl_101;
  wire G101_p_spl_11;
  wire G101_p_spl_110;
  wire G101_p_spl_111;
  wire G115_p_spl_;
  wire G115_p_spl_0;
  wire G115_p_spl_00;
  wire G115_p_spl_1;
  wire G101_n_spl_;
  wire G101_n_spl_0;
  wire G101_n_spl_00;
  wire G101_n_spl_000;
  wire G101_n_spl_001;
  wire G101_n_spl_01;
  wire G101_n_spl_010;
  wire G101_n_spl_011;
  wire G101_n_spl_1;
  wire G101_n_spl_10;
  wire G101_n_spl_100;
  wire G101_n_spl_101;
  wire G101_n_spl_11;
  wire G101_n_spl_110;
  wire G101_n_spl_111;
  wire G115_n_spl_;
  wire G115_n_spl_0;
  wire G115_n_spl_00;
  wire G115_n_spl_1;
  wire G100_p_spl_;
  wire G100_p_spl_0;
  wire G100_p_spl_00;
  wire G100_p_spl_000;
  wire G100_p_spl_0000;
  wire G100_p_spl_001;
  wire G100_p_spl_01;
  wire G100_p_spl_010;
  wire G100_p_spl_011;
  wire G100_p_spl_1;
  wire G100_p_spl_10;
  wire G100_p_spl_100;
  wire G100_p_spl_101;
  wire G100_p_spl_11;
  wire G100_p_spl_110;
  wire G100_p_spl_111;
  wire G100_n_spl_;
  wire G100_n_spl_0;
  wire G100_n_spl_00;
  wire G100_n_spl_000;
  wire G100_n_spl_0000;
  wire G100_n_spl_001;
  wire G100_n_spl_01;
  wire G100_n_spl_010;
  wire G100_n_spl_011;
  wire G100_n_spl_1;
  wire G100_n_spl_10;
  wire G100_n_spl_100;
  wire G100_n_spl_101;
  wire G100_n_spl_11;
  wire G100_n_spl_110;
  wire G100_n_spl_111;
  wire g237_n_spl_;
  wire g237_n_spl_0;
  wire g237_n_spl_1;
  wire g240_p_spl_;
  wire g237_p_spl_;
  wire g240_n_spl_;
  wire g240_n_spl_0;
  wire g241_n_spl_;
  wire G130_p_spl_;
  wire G130_p_spl_0;
  wire G130_p_spl_00;
  wire G130_p_spl_1;
  wire G130_n_spl_;
  wire G130_n_spl_0;
  wire G130_n_spl_00;
  wire G130_n_spl_1;
  wire G148_n_spl_;
  wire G148_n_spl_0;
  wire G148_n_spl_00;
  wire G148_n_spl_1;
  wire G148_p_spl_;
  wire G148_p_spl_0;
  wire G148_p_spl_00;
  wire G148_p_spl_1;
  wire g245_n_spl_;
  wire g245_n_spl_0;
  wire g245_n_spl_1;
  wire g248_n_spl_;
  wire G119_p_spl_;
  wire G119_p_spl_0;
  wire G119_p_spl_00;
  wire G119_p_spl_01;
  wire G119_p_spl_1;
  wire G119_p_spl_10;
  wire G119_n_spl_;
  wire G119_n_spl_0;
  wire G119_n_spl_00;
  wire G119_n_spl_01;
  wire G119_n_spl_1;
  wire G119_n_spl_10;
  wire G146_p_spl_;
  wire G146_p_spl_0;
  wire G146_p_spl_1;
  wire G146_n_spl_;
  wire G146_n_spl_0;
  wire G146_n_spl_1;
  wire G117_p_spl_;
  wire G117_p_spl_0;
  wire G117_p_spl_00;
  wire G117_p_spl_01;
  wire G117_p_spl_1;
  wire G117_p_spl_10;
  wire G117_n_spl_;
  wire G117_n_spl_0;
  wire G117_n_spl_00;
  wire G117_n_spl_01;
  wire G117_n_spl_1;
  wire G117_n_spl_10;
  wire G145_p_spl_;
  wire G145_p_spl_0;
  wire G145_p_spl_1;
  wire G145_n_spl_;
  wire G145_n_spl_0;
  wire G145_n_spl_1;
  wire g258_p_spl_;
  wire g267_p_spl_;
  wire g258_n_spl_;
  wire g258_n_spl_0;
  wire g267_n_spl_;
  wire g267_n_spl_0;
  wire G121_p_spl_;
  wire G121_p_spl_0;
  wire G121_p_spl_00;
  wire G121_p_spl_000;
  wire G121_p_spl_01;
  wire G121_p_spl_1;
  wire G121_p_spl_10;
  wire G121_p_spl_11;
  wire G121_n_spl_;
  wire G121_n_spl_0;
  wire G121_n_spl_00;
  wire G121_n_spl_000;
  wire G121_n_spl_01;
  wire G121_n_spl_1;
  wire G121_n_spl_10;
  wire G121_n_spl_11;
  wire G147_p_spl_;
  wire G147_p_spl_0;
  wire G147_p_spl_00;
  wire G147_p_spl_1;
  wire G147_n_spl_;
  wire G147_n_spl_0;
  wire G147_n_spl_00;
  wire G147_n_spl_1;
  wire g268_n_spl_;
  wire g277_n_spl_;
  wire G107_p_spl_;
  wire G107_p_spl_0;
  wire G107_p_spl_00;
  wire G107_p_spl_000;
  wire G107_p_spl_01;
  wire G107_p_spl_1;
  wire G107_p_spl_10;
  wire G107_p_spl_11;
  wire G107_n_spl_;
  wire G107_n_spl_0;
  wire G107_n_spl_00;
  wire G107_n_spl_000;
  wire G107_n_spl_01;
  wire G107_n_spl_1;
  wire G107_n_spl_10;
  wire G107_n_spl_11;
  wire G139_p_spl_;
  wire G139_p_spl_0;
  wire G139_p_spl_00;
  wire G139_p_spl_1;
  wire G139_n_spl_;
  wire G139_n_spl_0;
  wire G139_n_spl_00;
  wire G139_n_spl_1;
  wire G105_p_spl_;
  wire G105_p_spl_0;
  wire G105_p_spl_00;
  wire G105_p_spl_000;
  wire G105_p_spl_01;
  wire G105_p_spl_1;
  wire G105_p_spl_10;
  wire G105_p_spl_11;
  wire G105_n_spl_;
  wire G105_n_spl_0;
  wire G105_n_spl_00;
  wire G105_n_spl_000;
  wire G105_n_spl_01;
  wire G105_n_spl_1;
  wire G105_n_spl_10;
  wire G105_n_spl_11;
  wire G138_p_spl_;
  wire G138_p_spl_0;
  wire G138_p_spl_00;
  wire G138_p_spl_1;
  wire G138_n_spl_;
  wire G138_n_spl_0;
  wire G138_n_spl_00;
  wire G138_n_spl_1;
  wire g289_n_spl_;
  wire g298_n_spl_;
  wire G109_p_spl_;
  wire G109_p_spl_0;
  wire G109_p_spl_00;
  wire G109_p_spl_000;
  wire G109_p_spl_01;
  wire G109_p_spl_1;
  wire G109_p_spl_10;
  wire G109_p_spl_11;
  wire G109_n_spl_;
  wire G109_n_spl_0;
  wire G109_n_spl_00;
  wire G109_n_spl_000;
  wire G109_n_spl_01;
  wire G109_n_spl_1;
  wire G109_n_spl_10;
  wire G109_n_spl_11;
  wire G135_p_spl_;
  wire G135_p_spl_0;
  wire G135_p_spl_00;
  wire G135_p_spl_1;
  wire G135_n_spl_;
  wire G135_n_spl_0;
  wire G135_n_spl_00;
  wire G135_n_spl_1;
  wire G88_p_spl_;
  wire G88_p_spl_0;
  wire G88_p_spl_00;
  wire G88_p_spl_01;
  wire G88_p_spl_1;
  wire G88_p_spl_10;
  wire G88_n_spl_;
  wire G88_n_spl_0;
  wire G88_n_spl_00;
  wire G88_n_spl_01;
  wire G88_n_spl_1;
  wire G88_n_spl_10;
  wire G142_p_spl_;
  wire G142_p_spl_0;
  wire G142_p_spl_1;
  wire G142_n_spl_;
  wire G142_n_spl_0;
  wire G142_n_spl_1;
  wire g308_n_spl_;
  wire g317_n_spl_;
  wire g317_n_spl_0;
  wire g317_n_spl_1;
  wire G90_p_spl_;
  wire G90_p_spl_0;
  wire G90_p_spl_00;
  wire G90_p_spl_000;
  wire G90_p_spl_01;
  wire G90_p_spl_1;
  wire G90_p_spl_10;
  wire G90_p_spl_11;
  wire G90_n_spl_;
  wire G90_n_spl_0;
  wire G90_n_spl_00;
  wire G90_n_spl_000;
  wire G90_n_spl_01;
  wire G90_n_spl_1;
  wire G90_n_spl_10;
  wire G90_n_spl_11;
  wire G143_p_spl_;
  wire G143_p_spl_0;
  wire G143_p_spl_00;
  wire G143_p_spl_1;
  wire G143_n_spl_;
  wire G143_n_spl_0;
  wire G143_n_spl_00;
  wire G143_n_spl_1;
  wire G92_p_spl_;
  wire G92_p_spl_0;
  wire G92_p_spl_00;
  wire G92_p_spl_000;
  wire G92_p_spl_01;
  wire G92_p_spl_1;
  wire G92_p_spl_10;
  wire G92_p_spl_11;
  wire G92_n_spl_;
  wire G92_n_spl_0;
  wire G92_n_spl_00;
  wire G92_n_spl_000;
  wire G92_n_spl_01;
  wire G92_n_spl_1;
  wire G92_n_spl_10;
  wire G92_n_spl_11;
  wire G144_p_spl_;
  wire G144_p_spl_0;
  wire G144_p_spl_00;
  wire G144_p_spl_1;
  wire G144_n_spl_;
  wire G144_n_spl_0;
  wire G144_n_spl_00;
  wire G144_n_spl_1;
  wire g328_n_spl_;
  wire g337_n_spl_;
  wire G94_p_spl_;
  wire G94_p_spl_0;
  wire G94_p_spl_00;
  wire G94_p_spl_000;
  wire G94_p_spl_01;
  wire G94_p_spl_1;
  wire G94_p_spl_10;
  wire G94_p_spl_11;
  wire G94_n_spl_;
  wire G94_n_spl_0;
  wire G94_n_spl_00;
  wire G94_n_spl_000;
  wire G94_n_spl_01;
  wire G94_n_spl_1;
  wire G94_n_spl_10;
  wire G94_n_spl_11;
  wire G140_p_spl_;
  wire G140_p_spl_0;
  wire G140_p_spl_00;
  wire G140_p_spl_1;
  wire G140_n_spl_;
  wire G140_n_spl_0;
  wire G140_n_spl_00;
  wire G140_n_spl_1;
  wire G96_p_spl_;
  wire G96_p_spl_0;
  wire G96_p_spl_00;
  wire G96_p_spl_000;
  wire G96_p_spl_01;
  wire G96_p_spl_1;
  wire G96_p_spl_10;
  wire G96_p_spl_11;
  wire G96_n_spl_;
  wire G96_n_spl_0;
  wire G96_n_spl_00;
  wire G96_n_spl_000;
  wire G96_n_spl_01;
  wire G96_n_spl_1;
  wire G96_n_spl_10;
  wire G96_n_spl_11;
  wire G141_p_spl_;
  wire G141_p_spl_0;
  wire G141_p_spl_00;
  wire G141_p_spl_1;
  wire G141_n_spl_;
  wire G141_n_spl_0;
  wire G141_n_spl_00;
  wire G141_n_spl_1;
  wire G103_p_spl_;
  wire G103_p_spl_0;
  wire G103_p_spl_00;
  wire G103_p_spl_000;
  wire G103_p_spl_01;
  wire G103_p_spl_1;
  wire G103_p_spl_10;
  wire G103_p_spl_11;
  wire G103_n_spl_;
  wire G103_n_spl_0;
  wire G103_n_spl_00;
  wire G103_n_spl_000;
  wire G103_n_spl_01;
  wire G103_n_spl_1;
  wire G103_n_spl_10;
  wire G103_n_spl_11;
  wire G137_p_spl_;
  wire G137_p_spl_0;
  wire G137_p_spl_00;
  wire G137_p_spl_1;
  wire G137_n_spl_;
  wire G137_n_spl_0;
  wire G137_n_spl_00;
  wire G137_n_spl_1;
  wire g356_n_spl_;
  wire g365_n_spl_;
  wire g347_n_spl_;
  wire G124_n_spl_;
  wire G124_n_spl_0;
  wire G124_n_spl_00;
  wire G124_n_spl_000;
  wire G124_n_spl_0000;
  wire G124_n_spl_0001;
  wire G124_n_spl_001;
  wire G124_n_spl_0010;
  wire G124_n_spl_0011;
  wire G124_n_spl_01;
  wire G124_n_spl_010;
  wire G124_n_spl_011;
  wire G124_n_spl_1;
  wire G124_n_spl_10;
  wire G124_n_spl_100;
  wire G124_n_spl_101;
  wire G124_n_spl_11;
  wire G124_n_spl_110;
  wire G124_n_spl_111;
  wire G124_p_spl_;
  wire G124_p_spl_0;
  wire G124_p_spl_00;
  wire G124_p_spl_000;
  wire G124_p_spl_0000;
  wire G124_p_spl_0001;
  wire G124_p_spl_001;
  wire G124_p_spl_0010;
  wire G124_p_spl_0011;
  wire G124_p_spl_01;
  wire G124_p_spl_010;
  wire G124_p_spl_011;
  wire G124_p_spl_1;
  wire G124_p_spl_10;
  wire G124_p_spl_100;
  wire G124_p_spl_101;
  wire G124_p_spl_11;
  wire G124_p_spl_110;
  wire G124_p_spl_111;
  wire g372_p_spl_;
  wire g372_p_spl_0;
  wire g372_p_spl_1;
  wire g372_n_spl_;
  wire g372_n_spl_0;
  wire g372_n_spl_1;
  wire g373_n_spl_;
  wire g373_n_spl_0;
  wire g374_n_spl_;
  wire g374_n_spl_0;
  wire g374_n_spl_1;
  wire g373_p_spl_;
  wire g373_p_spl_0;
  wire g374_p_spl_;
  wire g374_p_spl_0;
  wire g374_p_spl_1;
  wire g378_p_spl_;
  wire g378_p_spl_0;
  wire g378_p_spl_1;
  wire g378_n_spl_;
  wire g378_n_spl_0;
  wire g378_n_spl_1;
  wire g379_n_spl_;
  wire g380_n_spl_;
  wire g379_p_spl_;
  wire g380_p_spl_;
  wire g375_p_spl_;
  wire g375_p_spl_0;
  wire g375_p_spl_00;
  wire g375_p_spl_1;
  wire g381_p_spl_;
  wire g381_p_spl_0;
  wire g381_p_spl_00;
  wire g381_p_spl_01;
  wire g381_p_spl_1;
  wire g381_p_spl_10;
  wire g375_n_spl_;
  wire g375_n_spl_0;
  wire g375_n_spl_00;
  wire g375_n_spl_1;
  wire g381_n_spl_;
  wire g381_n_spl_0;
  wire g381_n_spl_00;
  wire g381_n_spl_01;
  wire g381_n_spl_1;
  wire g381_n_spl_10;
  wire g385_p_spl_;
  wire g385_p_spl_0;
  wire g385_p_spl_1;
  wire g385_n_spl_;
  wire g385_n_spl_0;
  wire g385_n_spl_1;
  wire g386_n_spl_;
  wire g387_n_spl_;
  wire g386_p_spl_;
  wire g387_p_spl_;
  wire g382_p_spl_;
  wire g388_p_spl_;
  wire g388_p_spl_0;
  wire g388_p_spl_00;
  wire g388_p_spl_01;
  wire g388_p_spl_1;
  wire g382_n_spl_;
  wire g388_n_spl_;
  wire g388_n_spl_0;
  wire g388_n_spl_00;
  wire g388_n_spl_01;
  wire g388_n_spl_1;
  wire g392_p_spl_;
  wire g392_p_spl_0;
  wire g392_p_spl_1;
  wire g392_n_spl_;
  wire g392_n_spl_0;
  wire g392_n_spl_1;
  wire g393_n_spl_;
  wire g389_n_spl_;
  wire g389_n_spl_0;
  wire g395_n_spl_;
  wire g395_n_spl_0;
  wire g395_n_spl_00;
  wire g395_n_spl_01;
  wire g395_n_spl_1;
  wire g395_n_spl_10;
  wire g399_p_spl_;
  wire g399_p_spl_0;
  wire g399_p_spl_1;
  wire g399_n_spl_;
  wire g399_n_spl_0;
  wire g399_n_spl_1;
  wire g400_n_spl_;
  wire g400_n_spl_0;
  wire g400_n_spl_00;
  wire g400_n_spl_1;
  wire g401_n_spl_;
  wire g401_n_spl_0;
  wire g400_p_spl_;
  wire g400_p_spl_0;
  wire g400_p_spl_00;
  wire g400_p_spl_1;
  wire g401_p_spl_;
  wire g401_p_spl_0;
  wire g405_p_spl_;
  wire g405_p_spl_0;
  wire g405_p_spl_1;
  wire g405_n_spl_;
  wire g405_n_spl_0;
  wire g405_n_spl_1;
  wire g406_n_spl_;
  wire g406_n_spl_0;
  wire g406_p_spl_;
  wire g406_p_spl_0;
  wire g402_p_spl_;
  wire g402_p_spl_0;
  wire g402_p_spl_1;
  wire g408_p_spl_;
  wire g408_p_spl_0;
  wire g408_p_spl_1;
  wire g402_n_spl_;
  wire g402_n_spl_0;
  wire g408_n_spl_;
  wire g408_n_spl_0;
  wire g408_n_spl_00;
  wire g408_n_spl_1;
  wire g412_p_spl_;
  wire g412_p_spl_0;
  wire g412_p_spl_1;
  wire g412_n_spl_;
  wire g412_n_spl_0;
  wire g412_n_spl_1;
  wire g413_n_spl_;
  wire g413_p_spl_;
  wire g409_p_spl_;
  wire g409_p_spl_0;
  wire g415_p_spl_;
  wire g415_p_spl_0;
  wire g415_p_spl_00;
  wire g415_p_spl_1;
  wire g409_n_spl_;
  wire g409_n_spl_0;
  wire g415_n_spl_;
  wire g415_n_spl_0;
  wire g415_n_spl_00;
  wire g415_n_spl_1;
  wire g419_p_spl_;
  wire g419_p_spl_0;
  wire g419_p_spl_1;
  wire g419_n_spl_;
  wire g419_n_spl_0;
  wire g419_n_spl_1;
  wire g420_n_spl_;
  wire g420_n_spl_0;
  wire g420_p_spl_;
  wire g420_p_spl_0;
  wire g416_p_spl_;
  wire g416_p_spl_0;
  wire g422_p_spl_;
  wire g422_p_spl_0;
  wire g422_p_spl_00;
  wire g422_p_spl_1;
  wire g416_n_spl_;
  wire g416_n_spl_0;
  wire g422_n_spl_;
  wire g422_n_spl_0;
  wire g422_n_spl_00;
  wire g422_n_spl_01;
  wire g422_n_spl_1;
  wire g426_p_spl_;
  wire g426_p_spl_0;
  wire g426_p_spl_1;
  wire g426_n_spl_;
  wire g426_n_spl_0;
  wire g426_n_spl_1;
  wire g427_n_spl_;
  wire g427_p_spl_;
  wire g423_p_spl_;
  wire g429_p_spl_;
  wire g429_p_spl_0;
  wire g429_p_spl_00;
  wire g429_p_spl_01;
  wire g429_p_spl_1;
  wire g429_p_spl_10;
  wire g423_n_spl_;
  wire g429_n_spl_;
  wire g429_n_spl_0;
  wire g429_n_spl_00;
  wire g429_n_spl_01;
  wire g429_n_spl_1;
  wire g429_n_spl_10;
  wire g396_n_spl_;
  wire g430_n_spl_;
  wire g430_n_spl_0;
  wire g430_n_spl_1;
  wire G123_n_spl_;
  wire G123_n_spl_0;
  wire G123_n_spl_00;
  wire G123_n_spl_000;
  wire G123_n_spl_0000;
  wire G123_n_spl_0001;
  wire G123_n_spl_001;
  wire G123_n_spl_0010;
  wire G123_n_spl_01;
  wire G123_n_spl_010;
  wire G123_n_spl_011;
  wire G123_n_spl_1;
  wire G123_n_spl_10;
  wire G123_n_spl_100;
  wire G123_n_spl_101;
  wire G123_n_spl_11;
  wire G123_n_spl_110;
  wire G123_n_spl_111;
  wire G123_p_spl_;
  wire G123_p_spl_0;
  wire G123_p_spl_00;
  wire G123_p_spl_000;
  wire G123_p_spl_0000;
  wire G123_p_spl_0001;
  wire G123_p_spl_001;
  wire G123_p_spl_0010;
  wire G123_p_spl_01;
  wire G123_p_spl_010;
  wire G123_p_spl_011;
  wire G123_p_spl_1;
  wire G123_p_spl_10;
  wire G123_p_spl_100;
  wire G123_p_spl_101;
  wire G123_p_spl_11;
  wire G123_p_spl_110;
  wire G123_p_spl_111;
  wire g434_p_spl_;
  wire g434_p_spl_0;
  wire g434_p_spl_1;
  wire g434_n_spl_;
  wire g434_n_spl_0;
  wire g434_n_spl_1;
  wire g435_n_spl_;
  wire g435_p_spl_;
  wire g440_p_spl_;
  wire g440_p_spl_0;
  wire g440_p_spl_1;
  wire g440_n_spl_;
  wire g440_n_spl_0;
  wire g440_n_spl_1;
  wire g441_n_spl_;
  wire g441_n_spl_0;
  wire g441_n_spl_00;
  wire g441_n_spl_1;
  wire g442_n_spl_;
  wire g442_n_spl_0;
  wire g442_n_spl_1;
  wire g441_p_spl_;
  wire g441_p_spl_0;
  wire g441_p_spl_00;
  wire g441_p_spl_1;
  wire g442_p_spl_;
  wire g442_p_spl_0;
  wire g442_p_spl_1;
  wire g437_p_spl_;
  wire g437_p_spl_0;
  wire g437_p_spl_00;
  wire g437_p_spl_01;
  wire g437_p_spl_1;
  wire g443_p_spl_;
  wire g443_p_spl_0;
  wire g443_p_spl_00;
  wire g443_p_spl_1;
  wire g437_n_spl_;
  wire g437_n_spl_0;
  wire g437_n_spl_00;
  wire g437_n_spl_01;
  wire g437_n_spl_1;
  wire g443_n_spl_;
  wire g443_n_spl_0;
  wire g443_n_spl_00;
  wire g443_n_spl_1;
  wire g447_p_spl_;
  wire g447_p_spl_0;
  wire g447_p_spl_1;
  wire g447_n_spl_;
  wire g447_n_spl_0;
  wire g447_n_spl_1;
  wire g448_n_spl_;
  wire g448_p_spl_;
  wire G125_n_spl_;
  wire g451_n_spl_;
  wire g451_n_spl_0;
  wire g451_n_spl_1;
  wire g451_p_spl_;
  wire g451_p_spl_0;
  wire g451_p_spl_1;
  wire g452_n_spl_;
  wire g452_n_spl_0;
  wire g452_p_spl_;
  wire g452_p_spl_0;
  wire g450_p_spl_;
  wire g450_p_spl_0;
  wire g450_p_spl_1;
  wire g454_p_spl_;
  wire g454_p_spl_0;
  wire g454_p_spl_1;
  wire g450_n_spl_;
  wire g450_n_spl_0;
  wire g450_n_spl_1;
  wire g454_n_spl_;
  wire g454_n_spl_0;
  wire g454_n_spl_00;
  wire g454_n_spl_1;
  wire G129_n_spl_;
  wire g458_p_spl_;
  wire g458_p_spl_0;
  wire g458_p_spl_1;
  wire g458_n_spl_;
  wire g458_n_spl_0;
  wire g458_n_spl_1;
  wire g459_n_spl_;
  wire g459_n_spl_0;
  wire g459_p_spl_;
  wire g459_p_spl_0;
  wire G131_n_spl_;
  wire g461_p_spl_;
  wire g461_p_spl_0;
  wire g464_n_spl_;
  wire g464_n_spl_0;
  wire g464_n_spl_00;
  wire g464_n_spl_01;
  wire g464_n_spl_1;
  wire g464_n_spl_10;
  wire g461_n_spl_;
  wire g461_n_spl_0;
  wire g464_p_spl_;
  wire g464_p_spl_0;
  wire g464_p_spl_00;
  wire g464_p_spl_01;
  wire g464_p_spl_1;
  wire g464_p_spl_10;
  wire G127_n_spl_;
  wire g468_p_spl_;
  wire g468_p_spl_0;
  wire g468_p_spl_1;
  wire g468_n_spl_;
  wire g468_n_spl_0;
  wire g468_n_spl_1;
  wire g469_n_spl_;
  wire g469_n_spl_0;
  wire g469_p_spl_;
  wire g469_p_spl_0;
  wire g465_p_spl_;
  wire g465_p_spl_0;
  wire g471_p_spl_;
  wire g471_p_spl_0;
  wire g471_p_spl_1;
  wire g465_n_spl_;
  wire g465_n_spl_0;
  wire g471_n_spl_;
  wire g471_n_spl_0;
  wire g471_n_spl_00;
  wire g471_n_spl_1;
  wire g455_p_spl_;
  wire g472_p_spl_;
  wire g455_n_spl_;
  wire g472_n_spl_;
  wire G114_n_spl_;
  wire G114_n_spl_0;
  wire G114_p_spl_;
  wire g476_n_spl_;
  wire g476_n_spl_0;
  wire g476_n_spl_1;
  wire g479_n_spl_;
  wire g479_n_spl_0;
  wire g479_n_spl_00;
  wire g479_n_spl_01;
  wire g479_n_spl_1;
  wire g479_n_spl_10;
  wire g476_p_spl_;
  wire g476_p_spl_0;
  wire g476_p_spl_00;
  wire g476_p_spl_1;
  wire g479_p_spl_;
  wire g479_p_spl_0;
  wire g479_p_spl_00;
  wire g479_p_spl_01;
  wire g479_p_spl_1;
  wire g479_p_spl_10;
  wire g473_p_spl_;
  wire g480_p_spl_;
  wire g480_p_spl_0;
  wire g444_p_spl_;
  wire g444_p_spl_0;
  wire g485_p_spl_;
  wire g488_n_spl_;
  wire g485_n_spl_;
  wire g488_p_spl_;
  wire G132_n_spl_;
  wire G132_n_spl_0;
  wire G132_p_spl_;
  wire G132_p_spl_0;
  wire g494_n_spl_;
  wire g494_p_spl_;
  wire g497_n_spl_;
  wire g500_n_spl_;
  wire g497_p_spl_;
  wire g500_p_spl_;
  wire g509_p_spl_;
  wire g512_n_spl_;
  wire g509_n_spl_;
  wire g512_p_spl_;
  wire G111_n_spl_;
  wire G111_n_spl_0;
  wire G111_p_spl_;
  wire G111_p_spl_0;
  wire g518_n_spl_;
  wire g521_n_spl_;
  wire g518_p_spl_;
  wire g521_p_spl_;
  wire g524_n_spl_;
  wire g527_n_spl_;
  wire g524_p_spl_;
  wire g527_p_spl_;
  wire g535_n_spl_;
  wire g535_n_spl_0;
  wire g535_n_spl_1;
  wire g535_p_spl_;
  wire g535_p_spl_0;
  wire g535_p_spl_1;
  wire g537_n_spl_;
  wire g537_n_spl_0;
  wire g537_n_spl_00;
  wire g537_n_spl_1;
  wire g537_p_spl_;
  wire g537_p_spl_0;
  wire g537_p_spl_00;
  wire g537_p_spl_1;
  wire g539_n_spl_;
  wire g539_n_spl_0;
  wire g539_n_spl_1;
  wire g539_p_spl_;
  wire g539_p_spl_0;
  wire g539_p_spl_1;
  wire g541_p_spl_;
  wire g541_p_spl_0;
  wire g541_p_spl_00;
  wire g541_p_spl_1;
  wire g544_n_spl_;
  wire g544_n_spl_0;
  wire g544_n_spl_1;
  wire g544_p_spl_;
  wire g544_p_spl_0;
  wire g544_p_spl_1;
  wire g545_n_spl_;
  wire g545_p_spl_;
  wire g546_p_spl_;
  wire g546_p_spl_0;
  wire g546_p_spl_1;
  wire G177_p_spl_;
  wire G177_p_spl_0;
  wire G177_p_spl_00;
  wire G177_p_spl_000;
  wire G177_p_spl_0000;
  wire G177_p_spl_0001;
  wire G177_p_spl_001;
  wire G177_p_spl_0010;
  wire G177_p_spl_0011;
  wire G177_p_spl_01;
  wire G177_p_spl_010;
  wire G177_p_spl_0100;
  wire G177_p_spl_0101;
  wire G177_p_spl_011;
  wire G177_p_spl_0110;
  wire G177_p_spl_0111;
  wire G177_p_spl_1;
  wire G177_p_spl_10;
  wire G177_p_spl_100;
  wire G177_p_spl_1000;
  wire G177_p_spl_1001;
  wire G177_p_spl_101;
  wire G177_p_spl_11;
  wire G177_p_spl_110;
  wire G177_p_spl_111;
  wire g553_p_spl_;
  wire G176_p_spl_;
  wire G176_p_spl_0;
  wire G176_p_spl_00;
  wire G176_p_spl_000;
  wire G176_p_spl_0000;
  wire G176_p_spl_00000;
  wire G176_p_spl_00001;
  wire G176_p_spl_0001;
  wire G176_p_spl_001;
  wire G176_p_spl_0010;
  wire G176_p_spl_0011;
  wire G176_p_spl_01;
  wire G176_p_spl_010;
  wire G176_p_spl_0100;
  wire G176_p_spl_0101;
  wire G176_p_spl_011;
  wire G176_p_spl_0110;
  wire G176_p_spl_0111;
  wire G176_p_spl_1;
  wire G176_p_spl_10;
  wire G176_p_spl_100;
  wire G176_p_spl_1000;
  wire G176_p_spl_1001;
  wire G176_p_spl_101;
  wire G176_p_spl_1010;
  wire G176_p_spl_1011;
  wire G176_p_spl_11;
  wire G176_p_spl_110;
  wire G176_p_spl_1100;
  wire G176_p_spl_1101;
  wire G176_p_spl_111;
  wire G176_p_spl_1110;
  wire G176_p_spl_1111;
  wire G177_n_spl_;
  wire G177_n_spl_0;
  wire G177_n_spl_00;
  wire G177_n_spl_000;
  wire G177_n_spl_0000;
  wire G177_n_spl_0001;
  wire G177_n_spl_001;
  wire G177_n_spl_0010;
  wire G177_n_spl_0011;
  wire G177_n_spl_01;
  wire G177_n_spl_010;
  wire G177_n_spl_011;
  wire G177_n_spl_1;
  wire G177_n_spl_10;
  wire G177_n_spl_100;
  wire G177_n_spl_101;
  wire G177_n_spl_11;
  wire G177_n_spl_110;
  wire G177_n_spl_111;
  wire G176_n_spl_;
  wire G176_n_spl_0;
  wire G176_n_spl_00;
  wire G176_n_spl_000;
  wire G176_n_spl_0000;
  wire G176_n_spl_0001;
  wire G176_n_spl_001;
  wire G176_n_spl_0010;
  wire G176_n_spl_0011;
  wire G176_n_spl_01;
  wire G176_n_spl_010;
  wire G176_n_spl_0100;
  wire G176_n_spl_0101;
  wire G176_n_spl_011;
  wire G176_n_spl_1;
  wire G176_n_spl_10;
  wire G176_n_spl_100;
  wire G176_n_spl_101;
  wire G176_n_spl_11;
  wire G176_n_spl_110;
  wire G176_n_spl_111;
  wire g562_n_spl_;
  wire g562_n_spl_0;
  wire G2_p_spl_;
  wire G2_p_spl_0;
  wire G2_p_spl_1;
  wire G2_n_spl_;
  wire G2_n_spl_0;
  wire g570_n_spl_;
  wire g572_p_spl_;
  wire G22_p_spl_;
  wire G173_n_spl_;
  wire G173_n_spl_0;
  wire G173_n_spl_00;
  wire G173_n_spl_000;
  wire G173_n_spl_0000;
  wire G173_n_spl_0001;
  wire G173_n_spl_001;
  wire G173_n_spl_0010;
  wire G173_n_spl_0011;
  wire G173_n_spl_01;
  wire G173_n_spl_010;
  wire G173_n_spl_011;
  wire G173_n_spl_1;
  wire G173_n_spl_10;
  wire G173_n_spl_100;
  wire G173_n_spl_101;
  wire G173_n_spl_11;
  wire G173_n_spl_110;
  wire G173_n_spl_111;
  wire G3_p_spl_;
  wire G173_p_spl_;
  wire G173_p_spl_0;
  wire G173_p_spl_00;
  wire G173_p_spl_000;
  wire G173_p_spl_0000;
  wire G173_p_spl_0001;
  wire G173_p_spl_001;
  wire G173_p_spl_0010;
  wire G173_p_spl_0011;
  wire G173_p_spl_01;
  wire G173_p_spl_010;
  wire G173_p_spl_011;
  wire G173_p_spl_1;
  wire G173_p_spl_10;
  wire G173_p_spl_100;
  wire G173_p_spl_101;
  wire G173_p_spl_11;
  wire G173_p_spl_110;
  wire G173_p_spl_111;
  wire G172_n_spl_;
  wire G172_n_spl_0;
  wire G172_n_spl_00;
  wire G172_n_spl_000;
  wire G172_n_spl_001;
  wire G172_n_spl_01;
  wire G172_n_spl_1;
  wire G172_n_spl_10;
  wire G172_n_spl_11;
  wire g579_p_spl_;
  wire g579_p_spl_0;
  wire g579_p_spl_00;
  wire g579_p_spl_1;
  wire g560_p_spl_;
  wire g560_p_spl_0;
  wire g560_p_spl_00;
  wire g560_p_spl_1;
  wire G172_p_spl_;
  wire G172_p_spl_0;
  wire G172_p_spl_00;
  wire G172_p_spl_000;
  wire G172_p_spl_001;
  wire G172_p_spl_01;
  wire G172_p_spl_1;
  wire G172_p_spl_10;
  wire G172_p_spl_11;
  wire g594_n_spl_;
  wire g594_p_spl_;
  wire g595_n_spl_;
  wire g596_n_spl_;
  wire g596_n_spl_0;
  wire g596_p_spl_;
  wire g596_p_spl_0;
  wire g596_p_spl_1;
  wire g597_p_spl_;
  wire g598_p_spl_;
  wire g598_p_spl_0;
  wire g598_n_spl_;
  wire g598_n_spl_0;
  wire g601_p_spl_;
  wire g610_n_spl_;
  wire g617_p_spl_;
  wire g617_p_spl_0;
  wire g619_n_spl_;
  wire G174_n_spl_;
  wire G174_n_spl_0;
  wire G174_n_spl_00;
  wire G174_n_spl_000;
  wire G174_n_spl_0000;
  wire G174_n_spl_0001;
  wire G174_n_spl_001;
  wire G174_n_spl_0010;
  wire G174_n_spl_0011;
  wire G174_n_spl_01;
  wire G174_n_spl_010;
  wire G174_n_spl_011;
  wire G174_n_spl_1;
  wire G174_n_spl_10;
  wire G174_n_spl_100;
  wire G174_n_spl_101;
  wire G174_n_spl_11;
  wire G174_n_spl_110;
  wire G174_n_spl_111;
  wire G174_p_spl_;
  wire G174_p_spl_0;
  wire G174_p_spl_00;
  wire G174_p_spl_000;
  wire G174_p_spl_0000;
  wire G174_p_spl_0001;
  wire G174_p_spl_001;
  wire G174_p_spl_0010;
  wire G174_p_spl_0011;
  wire G174_p_spl_01;
  wire G174_p_spl_010;
  wire G174_p_spl_011;
  wire G174_p_spl_1;
  wire G174_p_spl_10;
  wire G174_p_spl_100;
  wire G174_p_spl_101;
  wire G174_p_spl_11;
  wire G174_p_spl_110;
  wire G174_p_spl_111;
  wire G175_n_spl_;
  wire G175_n_spl_0;
  wire G175_n_spl_00;
  wire G175_n_spl_000;
  wire G175_n_spl_001;
  wire G175_n_spl_01;
  wire G175_n_spl_1;
  wire G175_n_spl_10;
  wire G175_n_spl_11;
  wire G175_p_spl_;
  wire G175_p_spl_0;
  wire G175_p_spl_00;
  wire G175_p_spl_000;
  wire G175_p_spl_001;
  wire G175_p_spl_01;
  wire G175_p_spl_1;
  wire G175_p_spl_10;
  wire G175_p_spl_11;
  wire g638_p_spl_;
  wire g639_p_spl_;
  wire g643_n_spl_;
  wire g652_n_spl_;
  wire g659_p_spl_;
  wire g660_p_spl_;
  wire g664_n_spl_;
  wire g673_n_spl_;
  wire g581_n_spl_;
  wire g581_n_spl_0;
  wire g581_n_spl_00;
  wire g581_n_spl_01;
  wire g581_n_spl_1;
  wire g581_n_spl_10;
  wire g581_n_spl_11;
  wire g681_p_spl_;
  wire g581_p_spl_;
  wire g581_p_spl_0;
  wire g581_p_spl_00;
  wire g581_p_spl_01;
  wire g581_p_spl_1;
  wire g681_n_spl_;
  wire g687_n_spl_;
  wire g687_p_spl_;
  wire g693_n_spl_;
  wire g696_n_spl_;
  wire g693_p_spl_;
  wire g696_p_spl_;
  wire g690_p_spl_;
  wire g699_n_spl_;
  wire g690_n_spl_;
  wire g699_p_spl_;
  wire g708_p_spl_;
  wire g711_n_spl_;
  wire g708_n_spl_;
  wire g711_p_spl_;
  wire g717_n_spl_;
  wire g717_p_spl_;
  wire g720_p_spl_;
  wire g723_n_spl_;
  wire g720_n_spl_;
  wire g723_p_spl_;
  wire g726_n_spl_;
  wire g729_n_spl_;
  wire g726_p_spl_;
  wire g729_p_spl_;
  wire g430_p_spl_;
  wire g430_p_spl_0;
  wire g541_n_spl_;
  wire g541_n_spl_0;
  wire g541_n_spl_1;
  wire g737_p_spl_;
  wire g737_p_spl_0;
  wire g737_p_spl_00;
  wire g737_p_spl_1;
  wire g737_n_spl_;
  wire g737_n_spl_0;
  wire g737_n_spl_00;
  wire g737_n_spl_1;
  wire g743_p_spl_;
  wire g747_p_spl_;
  wire g389_p_spl_;
  wire g546_n_spl_;
  wire g546_n_spl_0;
  wire g395_p_spl_;
  wire g395_p_spl_0;
  wire g395_p_spl_00;
  wire g395_p_spl_1;
  wire g755_p_spl_;
  wire g760_p_spl_;
  wire g774_p_spl_;
  wire g774_p_spl_0;
  wire g774_p_spl_00;
  wire g774_p_spl_01;
  wire g774_p_spl_1;
  wire g774_n_spl_;
  wire g774_n_spl_0;
  wire g774_n_spl_00;
  wire g774_n_spl_01;
  wire g774_n_spl_1;
  wire g777_p_spl_;
  wire g444_n_spl_;
  wire g780_p_spl_;
  wire g780_p_spl_0;
  wire g780_p_spl_1;
  wire g780_n_spl_;
  wire g780_n_spl_0;
  wire g780_n_spl_1;
  wire g785_p_spl_;
  wire g791_p_spl_;
  wire G81_p_spl_;
  wire G158_n_spl_;
  wire G158_n_spl_0;
  wire G158_n_spl_00;
  wire G158_n_spl_000;
  wire G158_n_spl_0000;
  wire G158_n_spl_0001;
  wire G158_n_spl_001;
  wire G158_n_spl_0010;
  wire G158_n_spl_0011;
  wire G158_n_spl_01;
  wire G158_n_spl_010;
  wire G158_n_spl_011;
  wire G158_n_spl_1;
  wire G158_n_spl_10;
  wire G158_n_spl_100;
  wire G158_n_spl_101;
  wire G158_n_spl_11;
  wire G158_n_spl_110;
  wire G158_n_spl_111;
  wire G80_p_spl_;
  wire G158_p_spl_;
  wire G158_p_spl_0;
  wire G158_p_spl_00;
  wire G158_p_spl_000;
  wire G158_p_spl_0000;
  wire G158_p_spl_0001;
  wire G158_p_spl_001;
  wire G158_p_spl_0010;
  wire G158_p_spl_0011;
  wire G158_p_spl_01;
  wire G158_p_spl_010;
  wire G158_p_spl_011;
  wire G158_p_spl_1;
  wire G158_p_spl_10;
  wire G158_p_spl_100;
  wire G158_p_spl_101;
  wire G158_p_spl_11;
  wire G158_p_spl_110;
  wire G158_p_spl_111;
  wire G159_n_spl_;
  wire G159_n_spl_0;
  wire G159_n_spl_00;
  wire G159_n_spl_000;
  wire G159_n_spl_001;
  wire G159_n_spl_01;
  wire G159_n_spl_1;
  wire G159_n_spl_10;
  wire G159_n_spl_11;
  wire G159_p_spl_;
  wire G159_p_spl_0;
  wire G159_p_spl_00;
  wire G159_p_spl_000;
  wire G159_p_spl_001;
  wire G159_p_spl_01;
  wire G159_p_spl_1;
  wire G159_p_spl_10;
  wire G159_p_spl_11;
  wire G64_p_spl_;
  wire G64_p_spl_0;
  wire G64_p_spl_00;
  wire G64_p_spl_000;
  wire G64_p_spl_0000;
  wire G64_p_spl_0001;
  wire G64_p_spl_001;
  wire G64_p_spl_0010;
  wire G64_p_spl_01;
  wire G64_p_spl_010;
  wire G64_p_spl_011;
  wire G64_p_spl_1;
  wire G64_p_spl_10;
  wire G64_p_spl_100;
  wire G64_p_spl_101;
  wire G64_p_spl_11;
  wire G64_p_spl_110;
  wire G64_p_spl_111;
  wire G160_n_spl_;
  wire G160_n_spl_0;
  wire G160_n_spl_00;
  wire G160_n_spl_000;
  wire G160_n_spl_0000;
  wire G160_n_spl_0001;
  wire G160_n_spl_001;
  wire G160_n_spl_0010;
  wire G160_n_spl_0011;
  wire G160_n_spl_01;
  wire G160_n_spl_010;
  wire G160_n_spl_011;
  wire G160_n_spl_1;
  wire G160_n_spl_10;
  wire G160_n_spl_100;
  wire G160_n_spl_101;
  wire G160_n_spl_11;
  wire G160_n_spl_110;
  wire G160_n_spl_111;
  wire G160_p_spl_;
  wire G160_p_spl_0;
  wire G160_p_spl_00;
  wire G160_p_spl_000;
  wire G160_p_spl_0000;
  wire G160_p_spl_0001;
  wire G160_p_spl_001;
  wire G160_p_spl_0010;
  wire G160_p_spl_0011;
  wire G160_p_spl_01;
  wire G160_p_spl_010;
  wire G160_p_spl_011;
  wire G160_p_spl_1;
  wire G160_p_spl_10;
  wire G160_p_spl_100;
  wire G160_p_spl_101;
  wire G160_p_spl_11;
  wire G160_p_spl_110;
  wire G160_p_spl_111;
  wire G161_n_spl_;
  wire G161_n_spl_0;
  wire G161_n_spl_00;
  wire G161_n_spl_000;
  wire G161_n_spl_001;
  wire G161_n_spl_01;
  wire G161_n_spl_1;
  wire G161_n_spl_10;
  wire G161_n_spl_11;
  wire G161_p_spl_;
  wire G161_p_spl_0;
  wire G161_p_spl_00;
  wire G161_p_spl_000;
  wire G161_p_spl_001;
  wire G161_p_spl_01;
  wire G161_p_spl_1;
  wire G161_p_spl_10;
  wire G161_p_spl_11;
  wire G14_p_spl_;
  wire G16_p_spl_;
  wire g647_n_spl_;
  wire g647_n_spl_0;
  wire g647_n_spl_00;
  wire g647_n_spl_1;
  wire g605_n_spl_;
  wire g605_n_spl_0;
  wire g605_n_spl_00;
  wire g605_n_spl_1;
  wire G6_p_spl_;
  wire G27_p_spl_;
  wire g656_n_spl_;
  wire g656_n_spl_0;
  wire g656_n_spl_00;
  wire g656_n_spl_1;
  wire g614_n_spl_;
  wire g614_n_spl_0;
  wire g614_n_spl_00;
  wire g614_n_spl_1;
  wire G5_p_spl_;
  wire G26_p_spl_;
  wire g669_n_spl_;
  wire g669_n_spl_0;
  wire g669_n_spl_00;
  wire g669_n_spl_1;
  wire g624_n_spl_;
  wire g624_n_spl_0;
  wire g624_n_spl_00;
  wire g624_n_spl_1;
  wire G25_p_spl_;
  wire G24_p_spl_;
  wire g678_n_spl_;
  wire g678_n_spl_0;
  wire g678_n_spl_00;
  wire g678_n_spl_1;
  wire g569_p_spl_;
  wire g569_p_spl_0;
  wire g569_p_spl_00;
  wire g569_p_spl_1;
  wire G76_p_spl_;
  wire G86_p_spl_;
  wire G72_p_spl_;
  wire G82_p_spl_;
  wire G70_p_spl_;
  wire G71_p_spl_;
  wire G68_p_spl_;
  wire G69_p_spl_;
  wire G171_p_spl_;
  wire G54_p_spl_;
  wire G171_n_spl_;
  wire G61_n_spl_;
  wire G61_p_spl_;
  wire g975_p_spl_;
  wire G99_n_spl_;
  wire g533_n_spl_;
  wire g735_n_spl_;
  wire G155_n_spl_;
  wire g184_n_spl_;
  wire g179_n_spl_;
  wire g705_n_spl_;
  wire g506_n_spl_;
  wire g1025_n_spl_;
  wire g1025_n_spl_0;
  wire g1025_n_spl_00;
  wire g1025_n_spl_1;
  wire g990_p_spl_;
  wire g990_p_spl_0;
  wire g990_p_spl_00;
  wire g990_p_spl_1;
  wire G41_p_spl_;
  wire G42_p_spl_;
  wire G18_p_spl_;
  wire G17_p_spl_;
  wire g1032_n_spl_;
  wire g1032_n_spl_0;
  wire g1032_n_spl_00;
  wire g1032_n_spl_1;
  wire g997_n_spl_;
  wire g997_n_spl_0;
  wire g997_n_spl_00;
  wire g997_n_spl_1;
  wire G40_p_spl_;
  wire G39_p_spl_;
  wire g1039_n_spl_;
  wire g1039_n_spl_0;
  wire g1039_n_spl_00;
  wire g1039_n_spl_1;
  wire g1004_n_spl_;
  wire g1004_n_spl_0;
  wire g1004_n_spl_00;
  wire g1004_n_spl_1;
  wire G15_p_spl_;
  wire G36_p_spl_;
  wire g1046_n_spl_;
  wire g1046_n_spl_0;
  wire g1046_n_spl_00;
  wire g1046_n_spl_1;
  wire g1011_n_spl_;
  wire g1011_n_spl_0;
  wire g1011_n_spl_00;
  wire g1011_n_spl_1;
  wire G77_p_spl_;
  wire G87_p_spl_;
  wire G75_p_spl_;
  wire G85_p_spl_;
  wire G74_p_spl_;
  wire G84_p_spl_;
  wire G73_p_spl_;
  wire G83_p_spl_;
  wire g1200_p_spl_;
  wire g1202_n_spl_;
  wire g1200_n_spl_;
  wire g1202_p_spl_;
  wire g1214_n_spl_;
  wire g1223_p_spl_;
  wire g1214_p_spl_;
  wire g1223_n_spl_;
  wire g1229_n_spl_;
  wire g1238_p_spl_;
  wire g1229_p_spl_;
  wire g1238_n_spl_;
  wire g1241_p_spl_;
  wire g245_p_spl_;
  wire g1241_n_spl_;
  wire g1226_p_spl_;
  wire g1244_n_spl_;
  wire g1226_n_spl_;
  wire g1244_p_spl_;
  wire g1254_n_spl_;
  wire g617_n_spl_;
  wire g1254_p_spl_;
  wire g1257_p_spl_;
  wire g1257_n_spl_;
  wire G162_n_spl_;
  wire G162_p_spl_;
  wire g1260_p_spl_;
  wire g1263_p_spl_;
  wire g1260_n_spl_;
  wire g1263_n_spl_;
  wire g1268_n_spl_;
  wire g1268_p_spl_;
  wire g1266_n_spl_;
  wire g1271_n_spl_;
  wire g1266_p_spl_;
  wire g1271_p_spl_;
  wire g1275_n_spl_;
  wire g1275_p_spl_;
  wire g1278_p_spl_;
  wire g1278_n_spl_;
  wire g1281_p_spl_;
  wire g1281_n_spl_;
  wire g1282_n_spl_;
  wire g1282_p_spl_;
  wire g1284_n_spl_;
  wire g1284_p_spl_;
  wire g1288_n_spl_;
  wire g1288_p_spl_;
  wire g1299_p_spl_;
  wire g1299_n_spl_;
  wire g1308_n_spl_;
  wire g1320_n_spl_;
  wire g1329_p_spl_;
  wire g1320_p_spl_;
  wire g1329_n_spl_;
  wire g1341_n_spl_;
  wire g317_p_spl_;
  wire g1341_p_spl_;
  wire g1332_n_spl_;
  wire g1344_p_spl_;
  wire g1332_p_spl_;
  wire g1344_n_spl_;
  wire g1356_n_spl_;
  wire g1365_p_spl_;
  wire g1356_p_spl_;
  wire g1365_n_spl_;
  wire g1377_n_spl_;
  wire g1386_p_spl_;
  wire g1377_p_spl_;
  wire g1386_n_spl_;
  wire g1389_p_spl_;
  wire g1398_n_spl_;
  wire g1389_n_spl_;
  wire g1398_p_spl_;
  wire g1368_p_spl_;
  wire g1401_n_spl_;
  wire g1368_n_spl_;
  wire g1401_p_spl_;
  wire g1409_n_spl_;
  wire g1412_n_spl_;
  wire g1409_p_spl_;
  wire g1412_p_spl_;
  wire g1415_p_spl_;
  wire g1415_n_spl_;
  wire g1416_n_spl_;
  wire g1416_p_spl_;
  wire g1420_p_spl_;
  wire g1420_n_spl_;
  wire g1423_p_spl_;
  wire g1423_n_spl_;
  wire g1426_p_spl_;
  wire g1426_n_spl_;
  wire g1432_p_spl_;
  wire g1432_n_spl_;
  wire g1435_p_spl_;
  wire g1435_n_spl_;
  wire g1438_p_spl_;
  wire g1438_n_spl_;
  wire g1441_n_spl_;
  wire g1441_p_spl_;
  wire g1430_n_spl_;
  wire g1430_p_spl_;
  wire G157_n_spl_;
  wire G157_n_spl_0;
  wire G157_n_spl_1;
  wire G157_p_spl_;
  wire G157_p_spl_0;
  wire G157_p_spl_1;
  wire g1453_n_spl_;
  wire g1453_p_spl_;
  wire g1458_n_spl_;
  wire g1458_n_spl_0;
  wire g1458_n_spl_1;
  wire g1458_p_spl_;
  wire g1458_p_spl_0;
  wire g1458_p_spl_1;
  wire g1456_n_spl_;
  wire g1461_p_spl_;
  wire g1456_p_spl_;
  wire g1461_n_spl_;
  wire g1464_n_spl_;
  wire g1464_p_spl_;
  wire g1471_n_spl_;
  wire g1471_p_spl_;
  wire g1470_n_spl_;
  wire g1474_p_spl_;
  wire g1470_p_spl_;
  wire g1474_n_spl_;
  wire g1469_n_spl_;
  wire g1477_p_spl_;
  wire g1469_p_spl_;
  wire g1477_n_spl_;
  wire g1480_n_spl_;
  wire g1483_p_spl_;
  wire g1480_p_spl_;
  wire g1483_n_spl_;
  wire g1488_p_spl_;
  wire g1488_n_spl_;
  wire g1491_n_spl_;
  wire g1491_p_spl_;
  wire g1500_n_spl_;
  wire G23_n_spl_;
  wire G4_n_spl_;
  wire g1509_p_spl_;
  wire g1509_p_spl_0;
  wire g1509_p_spl_1;
  wire g1512_p_spl_;
  wire g1512_p_spl_0;
  wire g1512_p_spl_1;
  wire G79_n_spl_;
  wire G78_n_spl_;
  wire G64_n_spl_;
  wire G151_n_spl_;
  wire G151_n_spl_0;
  wire G152_p_spl_;
  wire G1_n_spl_;
  wire G1_n_spl_0;
  wire G1_n_spl_1;
  wire g194_n_spl_;
  wire g431_n_spl_;
  wire g482_p_spl_;
  wire g549_p_spl_;
  wire g550_n_spl_;

  FA
  g_g179_n
  (
    .dout(g179_n),
    .din1(G153_n_spl_),
    .din2(G156_n_spl_)
  );


  LA
  g_g180_p
  (
    .dout(g180_p),
    .din1(G66_p_spl_00),
    .din2(G67_p)
  );


  LA
  g_g181_p
  (
    .dout(g181_p),
    .din1(G1_p_spl_),
    .din2(G134_p)
  );


  LA
  g_g182_p
  (
    .dout(g182_p),
    .din1(G63_p),
    .din2(G165_n_spl_)
  );


  FA
  g_g183_n
  (
    .dout(g183_n),
    .din1(G11_n_spl_),
    .din2(G164_p)
  );


  FA
  g_g184_n
  (
    .dout(g184_n),
    .din1(G136_n),
    .din2(G154_n)
  );


  FA
  g_g185_n
  (
    .dout(g185_n),
    .din1(G11_n_spl_),
    .din2(G12_n)
  );


  FA
  g_g186_n
  (
    .dout(g186_n),
    .din1(G65_n),
    .din2(g185_n_spl_000)
  );


  FA
  g_g187_n
  (
    .dout(g187_n),
    .din1(G34_n),
    .din2(G163_n_spl_00)
  );


  FA
  g_g188_n
  (
    .dout(g188_n),
    .din1(G33_n),
    .din2(G163_p_spl_00)
  );


  LA
  g_g189_p
  (
    .dout(g189_p),
    .din1(g187_n),
    .din2(g188_n)
  );


  FA
  g_g190_n
  (
    .dout(g190_n),
    .din1(g185_n_spl_000),
    .din2(g189_p)
  );


  FA
  g_g191_n
  (
    .dout(g191_n),
    .din1(G13_n),
    .din2(G163_n_spl_00)
  );


  FA
  g_g192_n
  (
    .dout(g192_n),
    .din1(G35_n),
    .din2(G163_p_spl_00)
  );


  LA
  g_g193_p
  (
    .dout(g193_p),
    .din1(g191_n),
    .din2(g192_n)
  );


  FA
  g_g194_n
  (
    .dout(g194_n),
    .din1(g185_n_spl_00),
    .din2(g193_p)
  );


  FA
  g_g195_n
  (
    .dout(g195_n),
    .din1(G32_n),
    .din2(g185_n_spl_01)
  );


  LA
  g_g196_p
  (
    .dout(g196_p),
    .din1(G8_p),
    .din2(G163_p_spl_01)
  );


  LA
  g_g197_p
  (
    .dout(g197_p),
    .din1(G9_p),
    .din2(G163_n_spl_01)
  );


  FA
  g_g198_n
  (
    .dout(g198_n),
    .din1(g185_n_spl_01),
    .din2(g197_p)
  );


  FA
  g_g199_n
  (
    .dout(g199_n),
    .din1(g196_p),
    .din2(g198_n)
  );


  LA
  g_g200_p
  (
    .dout(g200_p),
    .din1(G66_p_spl_00),
    .din2(g199_n)
  );


  LA
  g_g201_p
  (
    .dout(g201_p),
    .din1(G10_p),
    .din2(G163_p_spl_01)
  );


  LA
  g_g202_p
  (
    .dout(g202_p),
    .din1(G30_p),
    .din2(G163_n_spl_01)
  );


  FA
  g_g203_n
  (
    .dout(g203_n),
    .din1(g185_n_spl_10),
    .din2(g202_p)
  );


  FA
  g_g204_n
  (
    .dout(g204_n),
    .din1(g201_p),
    .din2(g203_n)
  );


  LA
  g_g205_p
  (
    .dout(g205_p),
    .din1(G66_p_spl_01),
    .din2(g204_n)
  );


  LA
  g_g206_p
  (
    .dout(g206_p),
    .din1(G28_p),
    .din2(G163_p_spl_1)
  );


  LA
  g_g207_p
  (
    .dout(g207_p),
    .din1(G7_p),
    .din2(G163_n_spl_1)
  );


  FA
  g_g208_n
  (
    .dout(g208_n),
    .din1(g185_n_spl_10),
    .din2(g207_p)
  );


  FA
  g_g209_n
  (
    .dout(g209_n),
    .din1(g206_p),
    .din2(g208_n)
  );


  LA
  g_g210_p
  (
    .dout(g210_p),
    .din1(G66_p_spl_01),
    .din2(g209_n)
  );


  LA
  g_g211_p
  (
    .dout(g211_p),
    .din1(G31_p),
    .din2(G163_p_spl_1)
  );


  LA
  g_g212_p
  (
    .dout(g212_p),
    .din1(G29_p),
    .din2(G163_n_spl_1)
  );


  FA
  g_g213_n
  (
    .dout(g213_n),
    .din1(g185_n_spl_11),
    .din2(g212_p)
  );


  FA
  g_g214_n
  (
    .dout(g214_n),
    .din1(g211_p),
    .din2(g213_n)
  );


  LA
  g_g215_p
  (
    .dout(g215_p),
    .din1(G66_p_spl_1),
    .din2(g214_n)
  );


  LA
  g_g216_p
  (
    .dout(g216_p),
    .din1(G128_p_spl_000),
    .din2(G168_p_spl_000)
  );


  LA
  g_g217_p
  (
    .dout(g217_p),
    .din1(G128_n_spl_000),
    .din2(G169_p_spl_000)
  );


  FA
  g_g218_n
  (
    .dout(g218_n),
    .din1(g216_p),
    .din2(g217_p)
  );


  LA
  g_g219_p
  (
    .dout(g219_p),
    .din1(G150_p_spl_00),
    .din2(g218_n)
  );


  LA
  g_g220_p
  (
    .dout(g220_p),
    .din1(G128_p_spl_000),
    .din2(G167_n_spl_000)
  );


  LA
  g_g221_p
  (
    .dout(g221_p),
    .din1(G128_n_spl_000),
    .din2(G166_n_spl_000)
  );


  FA
  g_g222_n
  (
    .dout(g222_n),
    .din1(g220_p),
    .din2(g221_p)
  );


  LA
  g_g223_p
  (
    .dout(g223_p),
    .din1(G150_n_spl_00),
    .din2(g222_n)
  );


  FA
  g_g224_n
  (
    .dout(g224_n),
    .din1(g219_p),
    .din2(g223_p)
  );


  LA
  g_g225_p
  (
    .dout(g225_p),
    .din1(G126_p_spl_000),
    .din2(G168_p_spl_000)
  );


  LA
  g_g226_p
  (
    .dout(g226_p),
    .din1(G126_n_spl_000),
    .din2(G169_p_spl_000)
  );


  FA
  g_g227_n
  (
    .dout(g227_n),
    .din1(g225_p),
    .din2(g226_p)
  );


  LA
  g_g228_p
  (
    .dout(g228_p),
    .din1(G149_p_spl_00),
    .din2(g227_n)
  );


  LA
  g_g229_p
  (
    .dout(g229_p),
    .din1(G126_p_spl_000),
    .din2(G167_n_spl_000)
  );


  LA
  g_g230_p
  (
    .dout(g230_p),
    .din1(G126_n_spl_000),
    .din2(G166_n_spl_000)
  );


  FA
  g_g231_n
  (
    .dout(g231_n),
    .din1(g229_p),
    .din2(g230_p)
  );


  LA
  g_g232_p
  (
    .dout(g232_p),
    .din1(G149_n_spl_00),
    .din2(g231_n)
  );


  FA
  g_g233_n
  (
    .dout(g233_n),
    .din1(g228_p),
    .din2(g232_p)
  );


  FA
  g_g234_n
  (
    .dout(g234_n),
    .din1(g224_n_spl_),
    .din2(g233_n_spl_)
  );


  LA
  g_g235_p
  (
    .dout(g235_p),
    .din1(G102_p_spl_000),
    .din2(G113_p_spl_00)
  );


  FA
  g_g235_n
  (
    .dout(g235_n),
    .din1(G102_n_spl_000),
    .din2(G113_n_spl_00)
  );


  LA
  g_g236_p
  (
    .dout(g236_p),
    .din1(G98_p_spl_000),
    .din2(G113_n_spl_00)
  );


  FA
  g_g236_n
  (
    .dout(g236_n),
    .din1(G98_n_spl_000),
    .din2(G113_p_spl_00)
  );


  LA
  g_g237_p
  (
    .dout(g237_p),
    .din1(g235_n),
    .din2(g236_n)
  );


  FA
  g_g237_n
  (
    .dout(g237_n),
    .din1(g235_p),
    .din2(g236_p)
  );


  LA
  g_g238_p
  (
    .dout(g238_p),
    .din1(G101_p_spl_000),
    .din2(G115_p_spl_00)
  );


  FA
  g_g238_n
  (
    .dout(g238_n),
    .din1(G101_n_spl_000),
    .din2(G115_n_spl_00)
  );


  LA
  g_g239_p
  (
    .dout(g239_p),
    .din1(G100_p_spl_0000),
    .din2(G115_n_spl_00)
  );


  FA
  g_g239_n
  (
    .dout(g239_n),
    .din1(G100_n_spl_0000),
    .din2(G115_p_spl_00)
  );


  LA
  g_g240_p
  (
    .dout(g240_p),
    .din1(g238_n),
    .din2(g239_n)
  );


  FA
  g_g240_n
  (
    .dout(g240_n),
    .din1(g238_p),
    .din2(g239_p)
  );


  LA
  g_g241_p
  (
    .dout(g241_p),
    .din1(g237_n_spl_0),
    .din2(g240_p_spl_)
  );


  FA
  g_g241_n
  (
    .dout(g241_n),
    .din1(g237_p_spl_),
    .din2(g240_n_spl_0)
  );


  FA
  g_g242_n
  (
    .dout(g242_n),
    .din1(g234_n),
    .din2(g241_n_spl_)
  );


  LA
  g_g243_p
  (
    .dout(g243_p),
    .din1(G101_p_spl_000),
    .din2(G130_p_spl_00)
  );


  FA
  g_g243_n
  (
    .dout(g243_n),
    .din1(G101_n_spl_000),
    .din2(G130_n_spl_00)
  );


  LA
  g_g244_p
  (
    .dout(g244_p),
    .din1(G100_p_spl_0000),
    .din2(G130_n_spl_00)
  );


  FA
  g_g244_n
  (
    .dout(g244_n),
    .din1(G100_n_spl_0000),
    .din2(G130_p_spl_00)
  );


  LA
  g_g245_p
  (
    .dout(g245_p),
    .din1(g243_n),
    .din2(g244_n)
  );


  FA
  g_g245_n
  (
    .dout(g245_n),
    .din1(g243_p),
    .din2(g244_p)
  );


  LA
  g_g246_p
  (
    .dout(g246_p),
    .din1(G148_n_spl_00),
    .din2(G166_n_spl_001)
  );


  LA
  g_g247_p
  (
    .dout(g247_p),
    .din1(G148_p_spl_00),
    .din2(G169_p_spl_001)
  );


  FA
  g_g248_n
  (
    .dout(g248_n),
    .din1(g246_p),
    .din2(g247_p)
  );


  FA
  g_g249_n
  (
    .dout(g249_n),
    .din1(g245_n_spl_0),
    .din2(g248_n_spl_)
  );


  LA
  g_g250_p
  (
    .dout(g250_p),
    .din1(G101_p_spl_001),
    .din2(G119_p_spl_00)
  );


  FA
  g_g250_n
  (
    .dout(g250_n),
    .din1(G101_n_spl_001),
    .din2(G119_n_spl_00)
  );


  LA
  g_g251_p
  (
    .dout(g251_p),
    .din1(G100_p_spl_000),
    .din2(G119_n_spl_00)
  );


  FA
  g_g251_n
  (
    .dout(g251_n),
    .din1(G100_n_spl_000),
    .din2(G119_p_spl_00)
  );


  LA
  g_g252_p
  (
    .dout(g252_p),
    .din1(g250_n),
    .din2(g251_n)
  );


  FA
  g_g252_n
  (
    .dout(g252_n),
    .din1(g250_p),
    .din2(g251_p)
  );


  LA
  g_g253_p
  (
    .dout(g253_p),
    .din1(G146_p_spl_0),
    .din2(g252_n)
  );


  FA
  g_g253_n
  (
    .dout(g253_n),
    .din1(G146_n_spl_0),
    .din2(g252_p)
  );


  LA
  g_g254_p
  (
    .dout(g254_p),
    .din1(G102_n_spl_000),
    .din2(G119_p_spl_01)
  );


  FA
  g_g254_n
  (
    .dout(g254_n),
    .din1(G102_p_spl_000),
    .din2(G119_n_spl_01)
  );


  LA
  g_g255_p
  (
    .dout(g255_p),
    .din1(G98_n_spl_000),
    .din2(G119_n_spl_01)
  );


  FA
  g_g255_n
  (
    .dout(g255_n),
    .din1(G98_p_spl_000),
    .din2(G119_p_spl_01)
  );


  LA
  g_g256_p
  (
    .dout(g256_p),
    .din1(g254_n),
    .din2(g255_n)
  );


  FA
  g_g256_n
  (
    .dout(g256_n),
    .din1(g254_p),
    .din2(g255_p)
  );


  LA
  g_g257_p
  (
    .dout(g257_p),
    .din1(G146_n_spl_0),
    .din2(g256_n)
  );


  FA
  g_g257_n
  (
    .dout(g257_n),
    .din1(G146_p_spl_0),
    .din2(g256_p)
  );


  LA
  g_g258_p
  (
    .dout(g258_p),
    .din1(g253_n),
    .din2(g257_n)
  );


  FA
  g_g258_n
  (
    .dout(g258_n),
    .din1(g253_p),
    .din2(g257_p)
  );


  LA
  g_g259_p
  (
    .dout(g259_p),
    .din1(G101_p_spl_001),
    .din2(G117_p_spl_00)
  );


  FA
  g_g259_n
  (
    .dout(g259_n),
    .din1(G101_n_spl_001),
    .din2(G117_n_spl_00)
  );


  LA
  g_g260_p
  (
    .dout(g260_p),
    .din1(G100_p_spl_001),
    .din2(G117_n_spl_00)
  );


  FA
  g_g260_n
  (
    .dout(g260_n),
    .din1(G100_n_spl_001),
    .din2(G117_p_spl_00)
  );


  LA
  g_g261_p
  (
    .dout(g261_p),
    .din1(g259_n),
    .din2(g260_n)
  );


  FA
  g_g261_n
  (
    .dout(g261_n),
    .din1(g259_p),
    .din2(g260_p)
  );


  LA
  g_g262_p
  (
    .dout(g262_p),
    .din1(G145_p_spl_0),
    .din2(g261_n)
  );


  FA
  g_g262_n
  (
    .dout(g262_n),
    .din1(G145_n_spl_0),
    .din2(g261_p)
  );


  LA
  g_g263_p
  (
    .dout(g263_p),
    .din1(G102_n_spl_001),
    .din2(G117_p_spl_01)
  );


  FA
  g_g263_n
  (
    .dout(g263_n),
    .din1(G102_p_spl_001),
    .din2(G117_n_spl_01)
  );


  LA
  g_g264_p
  (
    .dout(g264_p),
    .din1(G98_n_spl_001),
    .din2(G117_n_spl_01)
  );


  FA
  g_g264_n
  (
    .dout(g264_n),
    .din1(G98_p_spl_001),
    .din2(G117_p_spl_01)
  );


  LA
  g_g265_p
  (
    .dout(g265_p),
    .din1(g263_n),
    .din2(g264_n)
  );


  FA
  g_g265_n
  (
    .dout(g265_n),
    .din1(g263_p),
    .din2(g264_p)
  );


  LA
  g_g266_p
  (
    .dout(g266_p),
    .din1(G145_n_spl_0),
    .din2(g265_n)
  );


  FA
  g_g266_n
  (
    .dout(g266_n),
    .din1(G145_p_spl_0),
    .din2(g265_p)
  );


  LA
  g_g267_p
  (
    .dout(g267_p),
    .din1(g262_n),
    .din2(g266_n)
  );


  FA
  g_g267_n
  (
    .dout(g267_n),
    .din1(g262_p),
    .din2(g266_p)
  );


  LA
  g_g268_p
  (
    .dout(g268_p),
    .din1(g258_p_spl_),
    .din2(g267_p_spl_)
  );


  FA
  g_g268_n
  (
    .dout(g268_n),
    .din1(g258_n_spl_0),
    .din2(g267_n_spl_0)
  );


  LA
  g_g269_p
  (
    .dout(g269_p),
    .din1(G121_p_spl_000),
    .din2(G168_p_spl_001)
  );


  LA
  g_g270_p
  (
    .dout(g270_p),
    .din1(G121_n_spl_000),
    .din2(G169_p_spl_001)
  );


  FA
  g_g271_n
  (
    .dout(g271_n),
    .din1(g269_p),
    .din2(g270_p)
  );


  LA
  g_g272_p
  (
    .dout(g272_p),
    .din1(G147_p_spl_00),
    .din2(g271_n)
  );


  LA
  g_g273_p
  (
    .dout(g273_p),
    .din1(G121_p_spl_000),
    .din2(G167_n_spl_001)
  );


  LA
  g_g274_p
  (
    .dout(g274_p),
    .din1(G121_n_spl_000),
    .din2(G166_n_spl_001)
  );


  FA
  g_g275_n
  (
    .dout(g275_n),
    .din1(g273_p),
    .din2(g274_p)
  );


  LA
  g_g276_p
  (
    .dout(g276_p),
    .din1(G147_n_spl_00),
    .din2(g275_n)
  );


  FA
  g_g277_n
  (
    .dout(g277_n),
    .din1(g272_p),
    .din2(g276_p)
  );


  FA
  g_g278_n
  (
    .dout(g278_n),
    .din1(g268_n_spl_),
    .din2(g277_n_spl_)
  );


  FA
  g_g279_n
  (
    .dout(g279_n),
    .din1(g249_n),
    .din2(g278_n)
  );


  FA
  g_g280_n
  (
    .dout(g280_n),
    .din1(g242_n),
    .din2(g279_n)
  );


  LA
  g_g281_p
  (
    .dout(g281_p),
    .din1(G107_p_spl_000),
    .din2(G168_p_spl_001)
  );


  LA
  g_g282_p
  (
    .dout(g282_p),
    .din1(G107_n_spl_000),
    .din2(G169_p_spl_010)
  );


  FA
  g_g283_n
  (
    .dout(g283_n),
    .din1(g281_p),
    .din2(g282_p)
  );


  LA
  g_g284_p
  (
    .dout(g284_p),
    .din1(G139_p_spl_00),
    .din2(g283_n)
  );


  LA
  g_g285_p
  (
    .dout(g285_p),
    .din1(G107_p_spl_000),
    .din2(G167_n_spl_001)
  );


  LA
  g_g286_p
  (
    .dout(g286_p),
    .din1(G107_n_spl_000),
    .din2(G166_n_spl_010)
  );


  FA
  g_g287_n
  (
    .dout(g287_n),
    .din1(g285_p),
    .din2(g286_p)
  );


  LA
  g_g288_p
  (
    .dout(g288_p),
    .din1(G139_n_spl_00),
    .din2(g287_n)
  );


  FA
  g_g289_n
  (
    .dout(g289_n),
    .din1(g284_p),
    .din2(g288_p)
  );


  LA
  g_g290_p
  (
    .dout(g290_p),
    .din1(G105_p_spl_000),
    .din2(G168_p_spl_010)
  );


  LA
  g_g291_p
  (
    .dout(g291_p),
    .din1(G105_n_spl_000),
    .din2(G169_p_spl_010)
  );


  FA
  g_g292_n
  (
    .dout(g292_n),
    .din1(g290_p),
    .din2(g291_p)
  );


  LA
  g_g293_p
  (
    .dout(g293_p),
    .din1(G138_p_spl_00),
    .din2(g292_n)
  );


  LA
  g_g294_p
  (
    .dout(g294_p),
    .din1(G105_p_spl_000),
    .din2(G167_n_spl_010)
  );


  LA
  g_g295_p
  (
    .dout(g295_p),
    .din1(G105_n_spl_000),
    .din2(G166_n_spl_010)
  );


  FA
  g_g296_n
  (
    .dout(g296_n),
    .din1(g294_p),
    .din2(g295_p)
  );


  LA
  g_g297_p
  (
    .dout(g297_p),
    .din1(G138_n_spl_00),
    .din2(g296_n)
  );


  FA
  g_g298_n
  (
    .dout(g298_n),
    .din1(g293_p),
    .din2(g297_p)
  );


  FA
  g_g299_n
  (
    .dout(g299_n),
    .din1(g289_n_spl_),
    .din2(g298_n_spl_)
  );


  LA
  g_g300_p
  (
    .dout(g300_p),
    .din1(G109_p_spl_000),
    .din2(G168_p_spl_010)
  );


  LA
  g_g301_p
  (
    .dout(g301_p),
    .din1(G109_n_spl_000),
    .din2(G169_p_spl_011)
  );


  FA
  g_g302_n
  (
    .dout(g302_n),
    .din1(g300_p),
    .din2(g301_p)
  );


  LA
  g_g303_p
  (
    .dout(g303_p),
    .din1(G135_p_spl_00),
    .din2(g302_n)
  );


  LA
  g_g304_p
  (
    .dout(g304_p),
    .din1(G109_p_spl_000),
    .din2(G167_n_spl_010)
  );


  LA
  g_g305_p
  (
    .dout(g305_p),
    .din1(G109_n_spl_000),
    .din2(G166_n_spl_011)
  );


  FA
  g_g306_n
  (
    .dout(g306_n),
    .din1(g304_p),
    .din2(g305_p)
  );


  LA
  g_g307_p
  (
    .dout(g307_p),
    .din1(G135_n_spl_00),
    .din2(g306_n)
  );


  FA
  g_g308_n
  (
    .dout(g308_n),
    .din1(g303_p),
    .din2(g307_p)
  );


  LA
  g_g309_p
  (
    .dout(g309_p),
    .din1(G88_p_spl_00),
    .din2(G100_p_spl_001)
  );


  FA
  g_g309_n
  (
    .dout(g309_n),
    .din1(G88_n_spl_00),
    .din2(G100_n_spl_001)
  );


  LA
  g_g310_p
  (
    .dout(g310_p),
    .din1(G88_n_spl_00),
    .din2(G101_p_spl_010)
  );


  FA
  g_g310_n
  (
    .dout(g310_n),
    .din1(G88_p_spl_00),
    .din2(G101_n_spl_010)
  );


  LA
  g_g311_p
  (
    .dout(g311_p),
    .din1(g309_n),
    .din2(g310_n)
  );


  FA
  g_g311_n
  (
    .dout(g311_n),
    .din1(g309_p),
    .din2(g310_p)
  );


  LA
  g_g312_p
  (
    .dout(g312_p),
    .din1(G142_p_spl_0),
    .din2(g311_n)
  );


  FA
  g_g312_n
  (
    .dout(g312_n),
    .din1(G142_n_spl_0),
    .din2(g311_p)
  );


  LA
  g_g313_p
  (
    .dout(g313_p),
    .din1(G88_n_spl_01),
    .din2(G102_n_spl_001)
  );


  FA
  g_g313_n
  (
    .dout(g313_n),
    .din1(G88_p_spl_01),
    .din2(G102_p_spl_001)
  );


  LA
  g_g314_p
  (
    .dout(g314_p),
    .din1(G88_p_spl_01),
    .din2(G98_n_spl_001)
  );


  FA
  g_g314_n
  (
    .dout(g314_n),
    .din1(G88_n_spl_01),
    .din2(G98_p_spl_001)
  );


  LA
  g_g315_p
  (
    .dout(g315_p),
    .din1(g313_n),
    .din2(g314_n)
  );


  FA
  g_g315_n
  (
    .dout(g315_n),
    .din1(g313_p),
    .din2(g314_p)
  );


  LA
  g_g316_p
  (
    .dout(g316_p),
    .din1(G142_n_spl_0),
    .din2(g315_n)
  );


  FA
  g_g316_n
  (
    .dout(g316_n),
    .din1(G142_p_spl_0),
    .din2(g315_p)
  );


  LA
  g_g317_p
  (
    .dout(g317_p),
    .din1(g312_n),
    .din2(g316_n)
  );


  FA
  g_g317_n
  (
    .dout(g317_n),
    .din1(g312_p),
    .din2(g316_p)
  );


  FA
  g_g318_n
  (
    .dout(g318_n),
    .din1(g308_n_spl_),
    .din2(g317_n_spl_0)
  );


  FA
  g_g319_n
  (
    .dout(g319_n),
    .din1(g299_n),
    .din2(g318_n)
  );


  LA
  g_g320_p
  (
    .dout(g320_p),
    .din1(G90_p_spl_000),
    .din2(G168_p_spl_01)
  );


  LA
  g_g321_p
  (
    .dout(g321_p),
    .din1(G90_n_spl_000),
    .din2(G169_p_spl_011)
  );


  FA
  g_g322_n
  (
    .dout(g322_n),
    .din1(g320_p),
    .din2(g321_p)
  );


  LA
  g_g323_p
  (
    .dout(g323_p),
    .din1(G143_p_spl_00),
    .din2(g322_n)
  );


  LA
  g_g324_p
  (
    .dout(g324_p),
    .din1(G90_p_spl_000),
    .din2(G167_n_spl_01)
  );


  LA
  g_g325_p
  (
    .dout(g325_p),
    .din1(G90_n_spl_000),
    .din2(G166_n_spl_011)
  );


  FA
  g_g326_n
  (
    .dout(g326_n),
    .din1(g324_p),
    .din2(g325_p)
  );


  LA
  g_g327_p
  (
    .dout(g327_p),
    .din1(G143_n_spl_00),
    .din2(g326_n)
  );


  FA
  g_g328_n
  (
    .dout(g328_n),
    .din1(g323_p),
    .din2(g327_p)
  );


  LA
  g_g329_p
  (
    .dout(g329_p),
    .din1(G92_p_spl_000),
    .din2(G168_p_spl_10)
  );


  LA
  g_g330_p
  (
    .dout(g330_p),
    .din1(G92_n_spl_000),
    .din2(G169_p_spl_10)
  );


  FA
  g_g331_n
  (
    .dout(g331_n),
    .din1(g329_p),
    .din2(g330_p)
  );


  LA
  g_g332_p
  (
    .dout(g332_p),
    .din1(G144_p_spl_00),
    .din2(g331_n)
  );


  LA
  g_g333_p
  (
    .dout(g333_p),
    .din1(G92_p_spl_000),
    .din2(G167_n_spl_10)
  );


  LA
  g_g334_p
  (
    .dout(g334_p),
    .din1(G92_n_spl_000),
    .din2(G166_n_spl_10)
  );


  FA
  g_g335_n
  (
    .dout(g335_n),
    .din1(g333_p),
    .din2(g334_p)
  );


  LA
  g_g336_p
  (
    .dout(g336_p),
    .din1(G144_n_spl_00),
    .din2(g335_n)
  );


  FA
  g_g337_n
  (
    .dout(g337_n),
    .din1(g332_p),
    .din2(g336_p)
  );


  FA
  g_g338_n
  (
    .dout(g338_n),
    .din1(g328_n_spl_),
    .din2(g337_n_spl_)
  );


  LA
  g_g339_p
  (
    .dout(g339_p),
    .din1(G94_p_spl_000),
    .din2(G168_p_spl_10)
  );


  LA
  g_g340_p
  (
    .dout(g340_p),
    .din1(G94_n_spl_000),
    .din2(G169_p_spl_10)
  );


  FA
  g_g341_n
  (
    .dout(g341_n),
    .din1(g339_p),
    .din2(g340_p)
  );


  LA
  g_g342_p
  (
    .dout(g342_p),
    .din1(G140_p_spl_00),
    .din2(g341_n)
  );


  LA
  g_g343_p
  (
    .dout(g343_p),
    .din1(G94_p_spl_000),
    .din2(G167_n_spl_10)
  );


  LA
  g_g344_p
  (
    .dout(g344_p),
    .din1(G94_n_spl_000),
    .din2(G166_n_spl_10)
  );


  FA
  g_g345_n
  (
    .dout(g345_n),
    .din1(g343_p),
    .din2(g344_p)
  );


  LA
  g_g346_p
  (
    .dout(g346_p),
    .din1(G140_n_spl_00),
    .din2(g345_n)
  );


  FA
  g_g347_n
  (
    .dout(g347_n),
    .din1(g342_p),
    .din2(g346_p)
  );


  LA
  g_g348_p
  (
    .dout(g348_p),
    .din1(G96_p_spl_000),
    .din2(G168_p_spl_11)
  );


  LA
  g_g349_p
  (
    .dout(g349_p),
    .din1(G96_n_spl_000),
    .din2(G169_p_spl_11)
  );


  FA
  g_g350_n
  (
    .dout(g350_n),
    .din1(g348_p),
    .din2(g349_p)
  );


  LA
  g_g351_p
  (
    .dout(g351_p),
    .din1(G141_p_spl_00),
    .din2(g350_n)
  );


  LA
  g_g352_p
  (
    .dout(g352_p),
    .din1(G96_p_spl_000),
    .din2(G167_n_spl_11)
  );


  LA
  g_g353_p
  (
    .dout(g353_p),
    .din1(G96_n_spl_000),
    .din2(G166_n_spl_11)
  );


  FA
  g_g354_n
  (
    .dout(g354_n),
    .din1(g352_p),
    .din2(g353_p)
  );


  LA
  g_g355_p
  (
    .dout(g355_p),
    .din1(G141_n_spl_00),
    .din2(g354_n)
  );


  FA
  g_g356_n
  (
    .dout(g356_n),
    .din1(g351_p),
    .din2(g355_p)
  );


  LA
  g_g357_p
  (
    .dout(g357_p),
    .din1(G103_p_spl_000),
    .din2(G168_p_spl_11)
  );


  LA
  g_g358_p
  (
    .dout(g358_p),
    .din1(G103_n_spl_000),
    .din2(G169_p_spl_11)
  );


  FA
  g_g359_n
  (
    .dout(g359_n),
    .din1(g357_p),
    .din2(g358_p)
  );


  LA
  g_g360_p
  (
    .dout(g360_p),
    .din1(G137_p_spl_00),
    .din2(g359_n)
  );


  LA
  g_g361_p
  (
    .dout(g361_p),
    .din1(G103_p_spl_000),
    .din2(G167_n_spl_11)
  );


  LA
  g_g362_p
  (
    .dout(g362_p),
    .din1(G103_n_spl_000),
    .din2(G166_n_spl_11)
  );


  FA
  g_g363_n
  (
    .dout(g363_n),
    .din1(g361_p),
    .din2(g362_p)
  );


  LA
  g_g364_p
  (
    .dout(g364_p),
    .din1(G137_n_spl_00),
    .din2(g363_n)
  );


  FA
  g_g365_n
  (
    .dout(g365_n),
    .din1(g360_p),
    .din2(g364_p)
  );


  FA
  g_g366_n
  (
    .dout(g366_n),
    .din1(g356_n_spl_),
    .din2(g365_n_spl_)
  );


  FA
  g_g367_n
  (
    .dout(g367_n),
    .din1(g347_n_spl_),
    .din2(g366_n)
  );


  FA
  g_g368_n
  (
    .dout(g368_n),
    .din1(g338_n),
    .din2(g367_n)
  );


  FA
  g_g369_n
  (
    .dout(g369_n),
    .din1(g319_n),
    .din2(g368_n)
  );


  LA
  g_g370_p
  (
    .dout(g370_p),
    .din1(G95_n),
    .din2(G124_n_spl_0000)
  );


  FA
  g_g370_n
  (
    .dout(g370_n),
    .din1(G95_p),
    .din2(G124_p_spl_0000)
  );


  LA
  g_g371_p
  (
    .dout(g371_p),
    .din1(G94_n_spl_00),
    .din2(G124_p_spl_0000)
  );


  FA
  g_g371_n
  (
    .dout(g371_n),
    .din1(G94_p_spl_00),
    .din2(G124_n_spl_0000)
  );


  LA
  g_g372_p
  (
    .dout(g372_p),
    .din1(g370_n),
    .din2(g371_n)
  );


  FA
  g_g372_n
  (
    .dout(g372_n),
    .din1(g370_p),
    .din2(g371_p)
  );


  LA
  g_g373_p
  (
    .dout(g373_p),
    .din1(G140_p_spl_00),
    .din2(g372_p_spl_0)
  );


  FA
  g_g373_n
  (
    .dout(g373_n),
    .din1(G140_n_spl_00),
    .din2(g372_n_spl_0)
  );


  LA
  g_g374_p
  (
    .dout(g374_p),
    .din1(G140_n_spl_0),
    .din2(g372_n_spl_0)
  );


  FA
  g_g374_n
  (
    .dout(g374_n),
    .din1(G140_p_spl_0),
    .din2(g372_p_spl_0)
  );


  LA
  g_g375_p
  (
    .dout(g375_p),
    .din1(g373_n_spl_0),
    .din2(g374_n_spl_0)
  );


  FA
  g_g375_n
  (
    .dout(g375_n),
    .din1(g373_p_spl_0),
    .din2(g374_p_spl_0)
  );


  LA
  g_g376_p
  (
    .dout(g376_p),
    .din1(G93_n),
    .din2(G124_n_spl_0001)
  );


  FA
  g_g376_n
  (
    .dout(g376_n),
    .din1(G93_p),
    .din2(G124_p_spl_0001)
  );


  LA
  g_g377_p
  (
    .dout(g377_p),
    .din1(G92_n_spl_00),
    .din2(G124_p_spl_0001)
  );


  FA
  g_g377_n
  (
    .dout(g377_n),
    .din1(G92_p_spl_00),
    .din2(G124_n_spl_0001)
  );


  LA
  g_g378_p
  (
    .dout(g378_p),
    .din1(g376_n),
    .din2(g377_n)
  );


  FA
  g_g378_n
  (
    .dout(g378_n),
    .din1(g376_p),
    .din2(g377_p)
  );


  LA
  g_g379_p
  (
    .dout(g379_p),
    .din1(G144_p_spl_00),
    .din2(g378_p_spl_0)
  );


  FA
  g_g379_n
  (
    .dout(g379_n),
    .din1(G144_n_spl_00),
    .din2(g378_n_spl_0)
  );


  LA
  g_g380_p
  (
    .dout(g380_p),
    .din1(G144_n_spl_0),
    .din2(g378_n_spl_0)
  );


  FA
  g_g380_n
  (
    .dout(g380_n),
    .din1(G144_p_spl_0),
    .din2(g378_p_spl_0)
  );


  LA
  g_g381_p
  (
    .dout(g381_p),
    .din1(g379_n_spl_),
    .din2(g380_n_spl_)
  );


  FA
  g_g381_n
  (
    .dout(g381_n),
    .din1(g379_p_spl_),
    .din2(g380_p_spl_)
  );


  LA
  g_g382_p
  (
    .dout(g382_p),
    .din1(g375_p_spl_00),
    .din2(g381_p_spl_00)
  );


  FA
  g_g382_n
  (
    .dout(g382_n),
    .din1(g375_n_spl_00),
    .din2(g381_n_spl_00)
  );


  LA
  g_g383_p
  (
    .dout(g383_p),
    .din1(G91_n),
    .din2(G124_n_spl_0010)
  );


  FA
  g_g383_n
  (
    .dout(g383_n),
    .din1(G91_p),
    .din2(G124_p_spl_0010)
  );


  LA
  g_g384_p
  (
    .dout(g384_p),
    .din1(G90_n_spl_00),
    .din2(G124_p_spl_0010)
  );


  FA
  g_g384_n
  (
    .dout(g384_n),
    .din1(G90_p_spl_00),
    .din2(G124_n_spl_0010)
  );


  LA
  g_g385_p
  (
    .dout(g385_p),
    .din1(g383_n),
    .din2(g384_n)
  );


  FA
  g_g385_n
  (
    .dout(g385_n),
    .din1(g383_p),
    .din2(g384_p)
  );


  LA
  g_g386_p
  (
    .dout(g386_p),
    .din1(G143_p_spl_00),
    .din2(g385_p_spl_0)
  );


  FA
  g_g386_n
  (
    .dout(g386_n),
    .din1(G143_n_spl_00),
    .din2(g385_n_spl_0)
  );


  LA
  g_g387_p
  (
    .dout(g387_p),
    .din1(G143_n_spl_0),
    .din2(g385_n_spl_0)
  );


  FA
  g_g387_n
  (
    .dout(g387_n),
    .din1(G143_p_spl_0),
    .din2(g385_p_spl_0)
  );


  LA
  g_g388_p
  (
    .dout(g388_p),
    .din1(g386_n_spl_),
    .din2(g387_n_spl_)
  );


  FA
  g_g388_n
  (
    .dout(g388_n),
    .din1(g386_p_spl_),
    .din2(g387_p_spl_)
  );


  LA
  g_g389_p
  (
    .dout(g389_p),
    .din1(g382_p_spl_),
    .din2(g388_p_spl_00)
  );


  FA
  g_g389_n
  (
    .dout(g389_n),
    .din1(g382_n_spl_),
    .din2(g388_n_spl_00)
  );


  LA
  g_g390_p
  (
    .dout(g390_p),
    .din1(G89_n),
    .din2(G124_n_spl_0011)
  );


  FA
  g_g390_n
  (
    .dout(g390_n),
    .din1(G89_p),
    .din2(G124_p_spl_0011)
  );


  LA
  g_g391_p
  (
    .dout(g391_p),
    .din1(G88_n_spl_10),
    .din2(G124_p_spl_0011)
  );


  FA
  g_g391_n
  (
    .dout(g391_n),
    .din1(G88_p_spl_10),
    .din2(G124_n_spl_0011)
  );


  LA
  g_g392_p
  (
    .dout(g392_p),
    .din1(g390_n),
    .din2(g391_n)
  );


  FA
  g_g392_n
  (
    .dout(g392_n),
    .din1(g390_p),
    .din2(g391_p)
  );


  LA
  g_g393_p
  (
    .dout(g393_p),
    .din1(G142_p_spl_1),
    .din2(g392_p_spl_0)
  );


  FA
  g_g393_n
  (
    .dout(g393_n),
    .din1(G142_n_spl_1),
    .din2(g392_n_spl_0)
  );


  LA
  g_g394_p
  (
    .dout(g394_p),
    .din1(G142_n_spl_1),
    .din2(g392_n_spl_0)
  );


  FA
  g_g394_n
  (
    .dout(g394_n),
    .din1(G142_p_spl_1),
    .din2(g392_p_spl_0)
  );


  LA
  g_g395_p
  (
    .dout(g395_p),
    .din1(g393_n_spl_),
    .din2(g394_n)
  );


  FA
  g_g395_n
  (
    .dout(g395_n),
    .din1(g393_p),
    .din2(g394_p)
  );


  FA
  g_g396_n
  (
    .dout(g396_n),
    .din1(g389_n_spl_0),
    .din2(g395_n_spl_00)
  );


  LA
  g_g397_p
  (
    .dout(g397_p),
    .din1(G110_n),
    .din2(G124_n_spl_010)
  );


  FA
  g_g397_n
  (
    .dout(g397_n),
    .din1(G110_p),
    .din2(G124_p_spl_010)
  );


  LA
  g_g398_p
  (
    .dout(g398_p),
    .din1(G109_n_spl_00),
    .din2(G124_p_spl_010)
  );


  FA
  g_g398_n
  (
    .dout(g398_n),
    .din1(G109_p_spl_00),
    .din2(G124_n_spl_010)
  );


  LA
  g_g399_p
  (
    .dout(g399_p),
    .din1(g397_n),
    .din2(g398_n)
  );


  FA
  g_g399_n
  (
    .dout(g399_n),
    .din1(g397_p),
    .din2(g398_p)
  );


  LA
  g_g400_p
  (
    .dout(g400_p),
    .din1(G135_p_spl_00),
    .din2(g399_p_spl_0)
  );


  FA
  g_g400_n
  (
    .dout(g400_n),
    .din1(G135_n_spl_00),
    .din2(g399_n_spl_0)
  );


  LA
  g_g401_p
  (
    .dout(g401_p),
    .din1(G135_n_spl_0),
    .din2(g399_n_spl_0)
  );


  FA
  g_g401_n
  (
    .dout(g401_n),
    .din1(G135_p_spl_0),
    .din2(g399_p_spl_0)
  );


  LA
  g_g402_p
  (
    .dout(g402_p),
    .din1(g400_n_spl_00),
    .din2(g401_n_spl_0)
  );


  FA
  g_g402_n
  (
    .dout(g402_n),
    .din1(g400_p_spl_00),
    .din2(g401_p_spl_0)
  );


  LA
  g_g403_p
  (
    .dout(g403_p),
    .din1(G108_n),
    .din2(G124_n_spl_011)
  );


  FA
  g_g403_n
  (
    .dout(g403_n),
    .din1(G108_p),
    .din2(G124_p_spl_011)
  );


  LA
  g_g404_p
  (
    .dout(g404_p),
    .din1(G107_n_spl_00),
    .din2(G124_p_spl_011)
  );


  FA
  g_g404_n
  (
    .dout(g404_n),
    .din1(G107_p_spl_00),
    .din2(G124_n_spl_011)
  );


  LA
  g_g405_p
  (
    .dout(g405_p),
    .din1(g403_n),
    .din2(g404_n)
  );


  FA
  g_g405_n
  (
    .dout(g405_n),
    .din1(g403_p),
    .din2(g404_p)
  );


  LA
  g_g406_p
  (
    .dout(g406_p),
    .din1(G139_p_spl_00),
    .din2(g405_p_spl_0)
  );


  FA
  g_g406_n
  (
    .dout(g406_n),
    .din1(G139_n_spl_00),
    .din2(g405_n_spl_0)
  );


  LA
  g_g407_p
  (
    .dout(g407_p),
    .din1(G139_n_spl_0),
    .din2(g405_n_spl_0)
  );


  FA
  g_g407_n
  (
    .dout(g407_n),
    .din1(G139_p_spl_0),
    .din2(g405_p_spl_0)
  );


  LA
  g_g408_p
  (
    .dout(g408_p),
    .din1(g406_n_spl_0),
    .din2(g407_n)
  );


  FA
  g_g408_n
  (
    .dout(g408_n),
    .din1(g406_p_spl_0),
    .din2(g407_p)
  );


  LA
  g_g409_p
  (
    .dout(g409_p),
    .din1(g402_p_spl_0),
    .din2(g408_p_spl_0)
  );


  FA
  g_g409_n
  (
    .dout(g409_n),
    .din1(g402_n_spl_0),
    .din2(g408_n_spl_00)
  );


  LA
  g_g410_p
  (
    .dout(g410_p),
    .din1(G106_n),
    .din2(G124_n_spl_100)
  );


  FA
  g_g410_n
  (
    .dout(g410_n),
    .din1(G106_p),
    .din2(G124_p_spl_100)
  );


  LA
  g_g411_p
  (
    .dout(g411_p),
    .din1(G105_n_spl_00),
    .din2(G124_p_spl_100)
  );


  FA
  g_g411_n
  (
    .dout(g411_n),
    .din1(G105_p_spl_00),
    .din2(G124_n_spl_100)
  );


  LA
  g_g412_p
  (
    .dout(g412_p),
    .din1(g410_n),
    .din2(g411_n)
  );


  FA
  g_g412_n
  (
    .dout(g412_n),
    .din1(g410_p),
    .din2(g411_p)
  );


  LA
  g_g413_p
  (
    .dout(g413_p),
    .din1(G138_p_spl_00),
    .din2(g412_p_spl_0)
  );


  FA
  g_g413_n
  (
    .dout(g413_n),
    .din1(G138_n_spl_00),
    .din2(g412_n_spl_0)
  );


  LA
  g_g414_p
  (
    .dout(g414_p),
    .din1(G138_n_spl_0),
    .din2(g412_n_spl_0)
  );


  FA
  g_g414_n
  (
    .dout(g414_n),
    .din1(G138_p_spl_0),
    .din2(g412_p_spl_0)
  );


  LA
  g_g415_p
  (
    .dout(g415_p),
    .din1(g413_n_spl_),
    .din2(g414_n)
  );


  FA
  g_g415_n
  (
    .dout(g415_n),
    .din1(g413_p_spl_),
    .din2(g414_p)
  );


  LA
  g_g416_p
  (
    .dout(g416_p),
    .din1(g409_p_spl_0),
    .din2(g415_p_spl_00)
  );


  FA
  g_g416_n
  (
    .dout(g416_n),
    .din1(g409_n_spl_0),
    .din2(g415_n_spl_00)
  );


  LA
  g_g417_p
  (
    .dout(g417_p),
    .din1(G104_n),
    .din2(G124_n_spl_101)
  );


  FA
  g_g417_n
  (
    .dout(g417_n),
    .din1(G104_p),
    .din2(G124_p_spl_101)
  );


  LA
  g_g418_p
  (
    .dout(g418_p),
    .din1(G103_n_spl_00),
    .din2(G124_p_spl_101)
  );


  FA
  g_g418_n
  (
    .dout(g418_n),
    .din1(G103_p_spl_00),
    .din2(G124_n_spl_101)
  );


  LA
  g_g419_p
  (
    .dout(g419_p),
    .din1(g417_n),
    .din2(g418_n)
  );


  FA
  g_g419_n
  (
    .dout(g419_n),
    .din1(g417_p),
    .din2(g418_p)
  );


  LA
  g_g420_p
  (
    .dout(g420_p),
    .din1(G137_p_spl_00),
    .din2(g419_p_spl_0)
  );


  FA
  g_g420_n
  (
    .dout(g420_n),
    .din1(G137_n_spl_00),
    .din2(g419_n_spl_0)
  );


  LA
  g_g421_p
  (
    .dout(g421_p),
    .din1(G137_n_spl_0),
    .din2(g419_n_spl_0)
  );


  FA
  g_g421_n
  (
    .dout(g421_n),
    .din1(G137_p_spl_0),
    .din2(g419_p_spl_0)
  );


  LA
  g_g422_p
  (
    .dout(g422_p),
    .din1(g420_n_spl_0),
    .din2(g421_n)
  );


  FA
  g_g422_n
  (
    .dout(g422_n),
    .din1(g420_p_spl_0),
    .din2(g421_p)
  );


  LA
  g_g423_p
  (
    .dout(g423_p),
    .din1(g416_p_spl_0),
    .din2(g422_p_spl_00)
  );


  FA
  g_g423_n
  (
    .dout(g423_n),
    .din1(g416_n_spl_0),
    .din2(g422_n_spl_00)
  );


  LA
  g_g424_p
  (
    .dout(g424_p),
    .din1(G97_n),
    .din2(G124_n_spl_110)
  );


  FA
  g_g424_n
  (
    .dout(g424_n),
    .din1(G97_p),
    .din2(G124_p_spl_110)
  );


  LA
  g_g425_p
  (
    .dout(g425_p),
    .din1(G96_n_spl_00),
    .din2(G124_p_spl_110)
  );


  FA
  g_g425_n
  (
    .dout(g425_n),
    .din1(G96_p_spl_00),
    .din2(G124_n_spl_110)
  );


  LA
  g_g426_p
  (
    .dout(g426_p),
    .din1(g424_n),
    .din2(g425_n)
  );


  FA
  g_g426_n
  (
    .dout(g426_n),
    .din1(g424_p),
    .din2(g425_p)
  );


  LA
  g_g427_p
  (
    .dout(g427_p),
    .din1(G141_p_spl_00),
    .din2(g426_p_spl_0)
  );


  FA
  g_g427_n
  (
    .dout(g427_n),
    .din1(G141_n_spl_00),
    .din2(g426_n_spl_0)
  );


  LA
  g_g428_p
  (
    .dout(g428_p),
    .din1(G141_n_spl_0),
    .din2(g426_n_spl_0)
  );


  FA
  g_g428_n
  (
    .dout(g428_n),
    .din1(G141_p_spl_0),
    .din2(g426_p_spl_0)
  );


  LA
  g_g429_p
  (
    .dout(g429_p),
    .din1(g427_n_spl_),
    .din2(g428_n)
  );


  FA
  g_g429_n
  (
    .dout(g429_n),
    .din1(g427_p_spl_),
    .din2(g428_p)
  );


  LA
  g_g430_p
  (
    .dout(g430_p),
    .din1(g423_p_spl_),
    .din2(g429_p_spl_00)
  );


  FA
  g_g430_n
  (
    .dout(g430_n),
    .din1(g423_n_spl_),
    .din2(g429_n_spl_00)
  );


  FA
  g_g431_n
  (
    .dout(g431_n),
    .din1(g396_n_spl_),
    .din2(g430_n_spl_0)
  );


  LA
  g_g432_p
  (
    .dout(g432_p),
    .din1(G118_n),
    .din2(G123_n_spl_0000)
  );


  FA
  g_g432_n
  (
    .dout(g432_n),
    .din1(G118_p),
    .din2(G123_p_spl_0000)
  );


  LA
  g_g433_p
  (
    .dout(g433_p),
    .din1(G117_n_spl_10),
    .din2(G123_p_spl_0000)
  );


  FA
  g_g433_n
  (
    .dout(g433_n),
    .din1(G117_p_spl_10),
    .din2(G123_n_spl_0000)
  );


  LA
  g_g434_p
  (
    .dout(g434_p),
    .din1(g432_n),
    .din2(g433_n)
  );


  FA
  g_g434_n
  (
    .dout(g434_n),
    .din1(g432_p),
    .din2(g433_p)
  );


  LA
  g_g435_p
  (
    .dout(g435_p),
    .din1(G145_p_spl_1),
    .din2(g434_p_spl_0)
  );


  FA
  g_g435_n
  (
    .dout(g435_n),
    .din1(G145_n_spl_1),
    .din2(g434_n_spl_0)
  );


  LA
  g_g436_p
  (
    .dout(g436_p),
    .din1(G145_n_spl_1),
    .din2(g434_n_spl_0)
  );


  FA
  g_g436_n
  (
    .dout(g436_n),
    .din1(G145_p_spl_1),
    .din2(g434_p_spl_0)
  );


  LA
  g_g437_p
  (
    .dout(g437_p),
    .din1(g435_n_spl_),
    .din2(g436_n)
  );


  FA
  g_g437_n
  (
    .dout(g437_n),
    .din1(g435_p_spl_),
    .din2(g436_p)
  );


  LA
  g_g438_p
  (
    .dout(g438_p),
    .din1(G120_n),
    .din2(G123_n_spl_0001)
  );


  FA
  g_g438_n
  (
    .dout(g438_n),
    .din1(G120_p),
    .din2(G123_p_spl_0001)
  );


  LA
  g_g439_p
  (
    .dout(g439_p),
    .din1(G119_n_spl_10),
    .din2(G123_p_spl_0001)
  );


  FA
  g_g439_n
  (
    .dout(g439_n),
    .din1(G119_p_spl_10),
    .din2(G123_n_spl_0001)
  );


  LA
  g_g440_p
  (
    .dout(g440_p),
    .din1(g438_n),
    .din2(g439_n)
  );


  FA
  g_g440_n
  (
    .dout(g440_n),
    .din1(g438_p),
    .din2(g439_p)
  );


  LA
  g_g441_p
  (
    .dout(g441_p),
    .din1(G146_p_spl_1),
    .din2(g440_p_spl_0)
  );


  FA
  g_g441_n
  (
    .dout(g441_n),
    .din1(G146_n_spl_1),
    .din2(g440_n_spl_0)
  );


  LA
  g_g442_p
  (
    .dout(g442_p),
    .din1(G146_n_spl_1),
    .din2(g440_n_spl_0)
  );


  FA
  g_g442_n
  (
    .dout(g442_n),
    .din1(G146_p_spl_1),
    .din2(g440_p_spl_0)
  );


  LA
  g_g443_p
  (
    .dout(g443_p),
    .din1(g441_n_spl_00),
    .din2(g442_n_spl_0)
  );


  FA
  g_g443_n
  (
    .dout(g443_n),
    .din1(g441_p_spl_00),
    .din2(g442_p_spl_0)
  );


  LA
  g_g444_p
  (
    .dout(g444_p),
    .din1(g437_p_spl_00),
    .din2(g443_p_spl_00)
  );


  FA
  g_g444_n
  (
    .dout(g444_n),
    .din1(g437_n_spl_00),
    .din2(g443_n_spl_00)
  );


  LA
  g_g445_p
  (
    .dout(g445_p),
    .din1(G122_n),
    .din2(G123_n_spl_0010)
  );


  FA
  g_g445_n
  (
    .dout(g445_n),
    .din1(G122_p),
    .din2(G123_p_spl_0010)
  );


  LA
  g_g446_p
  (
    .dout(g446_p),
    .din1(G121_n_spl_00),
    .din2(G123_p_spl_0010)
  );


  FA
  g_g446_n
  (
    .dout(g446_n),
    .din1(G121_p_spl_00),
    .din2(G123_n_spl_0010)
  );


  LA
  g_g447_p
  (
    .dout(g447_p),
    .din1(g445_n),
    .din2(g446_n)
  );


  FA
  g_g447_n
  (
    .dout(g447_n),
    .din1(g445_p),
    .din2(g446_p)
  );


  LA
  g_g448_p
  (
    .dout(g448_p),
    .din1(G147_p_spl_00),
    .din2(g447_p_spl_0)
  );


  FA
  g_g448_n
  (
    .dout(g448_n),
    .din1(G147_n_spl_00),
    .din2(g447_n_spl_0)
  );


  LA
  g_g449_p
  (
    .dout(g449_p),
    .din1(G147_n_spl_0),
    .din2(g447_n_spl_0)
  );


  FA
  g_g449_n
  (
    .dout(g449_n),
    .din1(G147_p_spl_0),
    .din2(g447_p_spl_0)
  );


  LA
  g_g450_p
  (
    .dout(g450_p),
    .din1(g448_n_spl_),
    .din2(g449_n)
  );


  FA
  g_g450_n
  (
    .dout(g450_n),
    .din1(g448_p_spl_),
    .din2(g449_p)
  );


  LA
  g_g451_p
  (
    .dout(g451_p),
    .din1(G123_n_spl_001),
    .din2(G125_n_spl_)
  );


  FA
  g_g451_n
  (
    .dout(g451_n),
    .din1(G123_p_spl_001),
    .din2(G125_p)
  );


  LA
  g_g452_p
  (
    .dout(g452_p),
    .din1(G148_p_spl_00),
    .din2(g451_n_spl_0)
  );


  FA
  g_g452_n
  (
    .dout(g452_n),
    .din1(G148_n_spl_00),
    .din2(g451_p_spl_0)
  );


  LA
  g_g453_p
  (
    .dout(g453_p),
    .din1(G148_n_spl_0),
    .din2(g451_p_spl_0)
  );


  FA
  g_g453_n
  (
    .dout(g453_n),
    .din1(G148_p_spl_0),
    .din2(g451_n_spl_0)
  );


  LA
  g_g454_p
  (
    .dout(g454_p),
    .din1(g452_n_spl_0),
    .din2(g453_n)
  );


  FA
  g_g454_n
  (
    .dout(g454_n),
    .din1(g452_p_spl_0),
    .din2(g453_p)
  );


  LA
  g_g455_p
  (
    .dout(g455_p),
    .din1(g450_p_spl_0),
    .din2(g454_p_spl_0)
  );


  FA
  g_g455_n
  (
    .dout(g455_n),
    .din1(g450_n_spl_0),
    .din2(g454_n_spl_00)
  );


  LA
  g_g456_p
  (
    .dout(g456_p),
    .din1(G123_n_spl_010),
    .din2(G129_n_spl_)
  );


  FA
  g_g456_n
  (
    .dout(g456_n),
    .din1(G123_p_spl_010),
    .din2(G129_p)
  );


  LA
  g_g457_p
  (
    .dout(g457_p),
    .din1(G123_p_spl_010),
    .din2(G128_n_spl_00)
  );


  FA
  g_g457_n
  (
    .dout(g457_n),
    .din1(G123_n_spl_010),
    .din2(G128_p_spl_00)
  );


  LA
  g_g458_p
  (
    .dout(g458_p),
    .din1(g456_n),
    .din2(g457_n)
  );


  FA
  g_g458_n
  (
    .dout(g458_n),
    .din1(g456_p),
    .din2(g457_p)
  );


  LA
  g_g459_p
  (
    .dout(g459_p),
    .din1(G150_p_spl_00),
    .din2(g458_p_spl_0)
  );


  FA
  g_g459_n
  (
    .dout(g459_n),
    .din1(G150_n_spl_00),
    .din2(g458_n_spl_0)
  );


  LA
  g_g460_p
  (
    .dout(g460_p),
    .din1(G150_n_spl_0),
    .din2(g458_n_spl_0)
  );


  FA
  g_g460_n
  (
    .dout(g460_n),
    .din1(G150_p_spl_0),
    .din2(g458_p_spl_0)
  );


  LA
  g_g461_p
  (
    .dout(g461_p),
    .din1(g459_n_spl_0),
    .din2(g460_n)
  );


  FA
  g_g461_n
  (
    .dout(g461_n),
    .din1(g459_p_spl_0),
    .din2(g460_p)
  );


  LA
  g_g462_p
  (
    .dout(g462_p),
    .din1(G123_n_spl_011),
    .din2(G131_n_spl_)
  );


  FA
  g_g462_n
  (
    .dout(g462_n),
    .din1(G123_p_spl_011),
    .din2(G131_p)
  );


  LA
  g_g463_p
  (
    .dout(g463_p),
    .din1(G123_p_spl_011),
    .din2(G130_n_spl_0)
  );


  FA
  g_g463_n
  (
    .dout(g463_n),
    .din1(G123_n_spl_011),
    .din2(G130_p_spl_0)
  );


  LA
  g_g464_p
  (
    .dout(g464_p),
    .din1(g462_n),
    .din2(g463_n)
  );


  FA
  g_g464_n
  (
    .dout(g464_n),
    .din1(g462_p),
    .din2(g463_p)
  );


  LA
  g_g465_p
  (
    .dout(g465_p),
    .din1(g461_p_spl_0),
    .din2(g464_n_spl_00)
  );


  FA
  g_g465_n
  (
    .dout(g465_n),
    .din1(g461_n_spl_0),
    .din2(g464_p_spl_00)
  );


  LA
  g_g466_p
  (
    .dout(g466_p),
    .din1(G123_n_spl_100),
    .din2(G127_n_spl_)
  );


  FA
  g_g466_n
  (
    .dout(g466_n),
    .din1(G123_p_spl_100),
    .din2(G127_p)
  );


  LA
  g_g467_p
  (
    .dout(g467_p),
    .din1(G123_p_spl_100),
    .din2(G126_n_spl_00)
  );


  FA
  g_g467_n
  (
    .dout(g467_n),
    .din1(G123_n_spl_100),
    .din2(G126_p_spl_00)
  );


  LA
  g_g468_p
  (
    .dout(g468_p),
    .din1(g466_n),
    .din2(g467_n)
  );


  FA
  g_g468_n
  (
    .dout(g468_n),
    .din1(g466_p),
    .din2(g467_p)
  );


  LA
  g_g469_p
  (
    .dout(g469_p),
    .din1(G149_p_spl_00),
    .din2(g468_p_spl_0)
  );


  FA
  g_g469_n
  (
    .dout(g469_n),
    .din1(G149_n_spl_00),
    .din2(g468_n_spl_0)
  );


  LA
  g_g470_p
  (
    .dout(g470_p),
    .din1(G149_n_spl_0),
    .din2(g468_n_spl_0)
  );


  FA
  g_g470_n
  (
    .dout(g470_n),
    .din1(G149_p_spl_0),
    .din2(g468_p_spl_0)
  );


  LA
  g_g471_p
  (
    .dout(g471_p),
    .din1(g469_n_spl_0),
    .din2(g470_n)
  );


  FA
  g_g471_n
  (
    .dout(g471_n),
    .din1(g469_p_spl_0),
    .din2(g470_p)
  );


  LA
  g_g472_p
  (
    .dout(g472_p),
    .din1(g465_p_spl_0),
    .din2(g471_p_spl_0)
  );


  FA
  g_g472_n
  (
    .dout(g472_n),
    .din1(g465_n_spl_0),
    .din2(g471_n_spl_00)
  );


  LA
  g_g473_p
  (
    .dout(g473_p),
    .din1(g455_p_spl_),
    .din2(g472_p_spl_)
  );


  FA
  g_g473_n
  (
    .dout(g473_n),
    .din1(g455_n_spl_),
    .din2(g472_n_spl_)
  );


  LA
  g_g474_p
  (
    .dout(g474_p),
    .din1(G114_n_spl_0),
    .din2(G123_n_spl_101)
  );


  FA
  g_g474_n
  (
    .dout(g474_n),
    .din1(G114_p_spl_),
    .din2(G123_p_spl_101)
  );


  LA
  g_g475_p
  (
    .dout(g475_p),
    .din1(G113_n_spl_01),
    .din2(G123_p_spl_101)
  );


  FA
  g_g475_n
  (
    .dout(g475_n),
    .din1(G113_p_spl_0),
    .din2(G123_n_spl_101)
  );


  LA
  g_g476_p
  (
    .dout(g476_p),
    .din1(g474_n),
    .din2(g475_n)
  );


  FA
  g_g476_n
  (
    .dout(g476_n),
    .din1(g474_p),
    .din2(g475_p)
  );


  LA
  g_g477_p
  (
    .dout(g477_p),
    .din1(G116_n),
    .din2(G123_n_spl_110)
  );


  FA
  g_g477_n
  (
    .dout(g477_n),
    .din1(G116_p),
    .din2(G123_p_spl_110)
  );


  LA
  g_g478_p
  (
    .dout(g478_p),
    .din1(G115_n_spl_0),
    .din2(G123_p_spl_110)
  );


  FA
  g_g478_n
  (
    .dout(g478_n),
    .din1(G115_p_spl_0),
    .din2(G123_n_spl_110)
  );


  LA
  g_g479_p
  (
    .dout(g479_p),
    .din1(g477_n),
    .din2(g478_n)
  );


  FA
  g_g479_n
  (
    .dout(g479_n),
    .din1(g477_p),
    .din2(g478_p)
  );


  LA
  g_g480_p
  (
    .dout(g480_p),
    .din1(g476_n_spl_0),
    .din2(g479_n_spl_00)
  );


  FA
  g_g480_n
  (
    .dout(g480_n),
    .din1(g476_p_spl_00),
    .din2(g479_p_spl_00)
  );


  LA
  g_g481_p
  (
    .dout(g481_p),
    .din1(g473_p_spl_),
    .din2(g480_p_spl_0)
  );


  LA
  g_g482_p
  (
    .dout(g482_p),
    .din1(g444_p_spl_0),
    .din2(g481_p)
  );


  LA
  g_g483_p
  (
    .dout(g483_p),
    .din1(G117_n_spl_10),
    .din2(G119_n_spl_10)
  );


  FA
  g_g483_n
  (
    .dout(g483_n),
    .din1(G117_p_spl_10),
    .din2(G119_p_spl_10)
  );


  LA
  g_g484_p
  (
    .dout(g484_p),
    .din1(G117_p_spl_1),
    .din2(G119_p_spl_1)
  );


  FA
  g_g484_n
  (
    .dout(g484_n),
    .din1(G117_n_spl_1),
    .din2(G119_n_spl_1)
  );


  LA
  g_g485_p
  (
    .dout(g485_p),
    .din1(g483_n),
    .din2(g484_n)
  );


  FA
  g_g485_n
  (
    .dout(g485_n),
    .din1(g483_p),
    .din2(g484_p)
  );


  LA
  g_g486_p
  (
    .dout(g486_p),
    .din1(G113_n_spl_01),
    .din2(G115_n_spl_1)
  );


  FA
  g_g486_n
  (
    .dout(g486_n),
    .din1(G113_p_spl_1),
    .din2(G115_p_spl_1)
  );


  LA
  g_g487_p
  (
    .dout(g487_p),
    .din1(G113_p_spl_1),
    .din2(G115_p_spl_1)
  );


  FA
  g_g487_n
  (
    .dout(g487_n),
    .din1(G113_n_spl_1),
    .din2(G115_n_spl_1)
  );


  LA
  g_g488_p
  (
    .dout(g488_p),
    .din1(g486_n),
    .din2(g487_n)
  );


  FA
  g_g488_n
  (
    .dout(g488_n),
    .din1(g486_p),
    .din2(g487_p)
  );


  LA
  g_g489_p
  (
    .dout(g489_p),
    .din1(g485_p_spl_),
    .din2(g488_n_spl_)
  );


  FA
  g_g489_n
  (
    .dout(g489_n),
    .din1(g485_n_spl_),
    .din2(g488_p_spl_)
  );


  LA
  g_g490_p
  (
    .dout(g490_p),
    .din1(g485_n_spl_),
    .din2(g488_p_spl_)
  );


  FA
  g_g490_n
  (
    .dout(g490_n),
    .din1(g485_p_spl_),
    .din2(g488_n_spl_)
  );


  LA
  g_g491_p
  (
    .dout(g491_p),
    .din1(g489_n),
    .din2(g490_n)
  );


  FA
  g_g491_n
  (
    .dout(g491_n),
    .din1(g489_p),
    .din2(g490_p)
  );


  LA
  g_g492_p
  (
    .dout(g492_p),
    .din1(G130_n_spl_1),
    .din2(G132_n_spl_0)
  );


  FA
  g_g492_n
  (
    .dout(g492_n),
    .din1(G130_p_spl_1),
    .din2(G132_p_spl_0)
  );


  LA
  g_g493_p
  (
    .dout(g493_p),
    .din1(G130_p_spl_1),
    .din2(G132_p_spl_0)
  );


  FA
  g_g493_n
  (
    .dout(g493_n),
    .din1(G130_n_spl_1),
    .din2(G132_n_spl_0)
  );


  LA
  g_g494_p
  (
    .dout(g494_p),
    .din1(g492_n),
    .din2(g493_n)
  );


  FA
  g_g494_n
  (
    .dout(g494_n),
    .din1(g492_p),
    .din2(g493_p)
  );


  LA
  g_g495_p
  (
    .dout(g495_p),
    .din1(G121_p_spl_01),
    .din2(g494_n_spl_)
  );


  FA
  g_g495_n
  (
    .dout(g495_n),
    .din1(G121_n_spl_01),
    .din2(g494_p_spl_)
  );


  LA
  g_g496_p
  (
    .dout(g496_p),
    .din1(G121_n_spl_01),
    .din2(g494_p_spl_)
  );


  FA
  g_g496_n
  (
    .dout(g496_n),
    .din1(G121_p_spl_01),
    .din2(g494_n_spl_)
  );


  LA
  g_g497_p
  (
    .dout(g497_p),
    .din1(g495_n),
    .din2(g496_n)
  );


  FA
  g_g497_n
  (
    .dout(g497_n),
    .din1(g495_p),
    .din2(g496_p)
  );


  LA
  g_g498_p
  (
    .dout(g498_p),
    .din1(G126_n_spl_01),
    .din2(G128_n_spl_01)
  );


  FA
  g_g498_n
  (
    .dout(g498_n),
    .din1(G126_p_spl_01),
    .din2(G128_p_spl_01)
  );


  LA
  g_g499_p
  (
    .dout(g499_p),
    .din1(G126_p_spl_01),
    .din2(G128_p_spl_01)
  );


  FA
  g_g499_n
  (
    .dout(g499_n),
    .din1(G126_n_spl_01),
    .din2(G128_n_spl_01)
  );


  LA
  g_g500_p
  (
    .dout(g500_p),
    .din1(g498_n),
    .din2(g499_n)
  );


  FA
  g_g500_n
  (
    .dout(g500_n),
    .din1(g498_p),
    .din2(g499_p)
  );


  LA
  g_g501_p
  (
    .dout(g501_p),
    .din1(g497_n_spl_),
    .din2(g500_n_spl_)
  );


  FA
  g_g501_n
  (
    .dout(g501_n),
    .din1(g497_p_spl_),
    .din2(g500_p_spl_)
  );


  LA
  g_g502_p
  (
    .dout(g502_p),
    .din1(g497_p_spl_),
    .din2(g500_p_spl_)
  );


  FA
  g_g502_n
  (
    .dout(g502_n),
    .din1(g497_n_spl_),
    .din2(g500_n_spl_)
  );


  LA
  g_g503_p
  (
    .dout(g503_p),
    .din1(g501_n),
    .din2(g502_n)
  );


  FA
  g_g503_n
  (
    .dout(g503_n),
    .din1(g501_p),
    .din2(g502_p)
  );


  LA
  g_g504_p
  (
    .dout(g504_p),
    .din1(g491_n),
    .din2(g503_p)
  );


  LA
  g_g505_p
  (
    .dout(g505_p),
    .din1(g491_p),
    .din2(g503_n)
  );


  FA
  g_g506_n
  (
    .dout(g506_n),
    .din1(g504_p),
    .din2(g505_p)
  );


  LA
  g_g507_p
  (
    .dout(g507_p),
    .din1(G92_n_spl_01),
    .din2(G94_n_spl_01)
  );


  FA
  g_g507_n
  (
    .dout(g507_n),
    .din1(G92_p_spl_01),
    .din2(G94_p_spl_01)
  );


  LA
  g_g508_p
  (
    .dout(g508_p),
    .din1(G92_p_spl_01),
    .din2(G94_p_spl_01)
  );


  FA
  g_g508_n
  (
    .dout(g508_n),
    .din1(G92_n_spl_01),
    .din2(G94_n_spl_01)
  );


  LA
  g_g509_p
  (
    .dout(g509_p),
    .din1(g507_n),
    .din2(g508_n)
  );


  FA
  g_g509_n
  (
    .dout(g509_n),
    .din1(g507_p),
    .din2(g508_p)
  );


  LA
  g_g510_p
  (
    .dout(g510_p),
    .din1(G88_p_spl_10),
    .din2(G90_n_spl_01)
  );


  FA
  g_g510_n
  (
    .dout(g510_n),
    .din1(G88_n_spl_10),
    .din2(G90_p_spl_01)
  );


  LA
  g_g511_p
  (
    .dout(g511_p),
    .din1(G88_n_spl_1),
    .din2(G90_p_spl_01)
  );


  FA
  g_g511_n
  (
    .dout(g511_n),
    .din1(G88_p_spl_1),
    .din2(G90_n_spl_01)
  );


  LA
  g_g512_p
  (
    .dout(g512_p),
    .din1(g510_n),
    .din2(g511_n)
  );


  FA
  g_g512_n
  (
    .dout(g512_n),
    .din1(g510_p),
    .din2(g511_p)
  );


  LA
  g_g513_p
  (
    .dout(g513_p),
    .din1(g509_p_spl_),
    .din2(g512_n_spl_)
  );


  FA
  g_g513_n
  (
    .dout(g513_n),
    .din1(g509_n_spl_),
    .din2(g512_p_spl_)
  );


  LA
  g_g514_p
  (
    .dout(g514_p),
    .din1(g509_n_spl_),
    .din2(g512_p_spl_)
  );


  FA
  g_g514_n
  (
    .dout(g514_n),
    .din1(g509_p_spl_),
    .din2(g512_n_spl_)
  );


  LA
  g_g515_p
  (
    .dout(g515_p),
    .din1(g513_n),
    .din2(g514_n)
  );


  FA
  g_g515_n
  (
    .dout(g515_n),
    .din1(g513_p),
    .din2(g514_p)
  );


  LA
  g_g516_p
  (
    .dout(g516_p),
    .din1(G96_n_spl_01),
    .din2(G103_n_spl_01)
  );


  FA
  g_g516_n
  (
    .dout(g516_n),
    .din1(G96_p_spl_01),
    .din2(G103_p_spl_01)
  );


  LA
  g_g517_p
  (
    .dout(g517_p),
    .din1(G96_p_spl_01),
    .din2(G103_p_spl_01)
  );


  FA
  g_g517_n
  (
    .dout(g517_n),
    .din1(G96_n_spl_01),
    .din2(G103_n_spl_01)
  );


  LA
  g_g518_p
  (
    .dout(g518_p),
    .din1(g516_n),
    .din2(g517_n)
  );


  FA
  g_g518_n
  (
    .dout(g518_n),
    .din1(g516_p),
    .din2(g517_p)
  );


  LA
  g_g519_p
  (
    .dout(g519_p),
    .din1(G109_n_spl_01),
    .din2(G111_n_spl_0)
  );


  FA
  g_g519_n
  (
    .dout(g519_n),
    .din1(G109_p_spl_01),
    .din2(G111_p_spl_0)
  );


  LA
  g_g520_p
  (
    .dout(g520_p),
    .din1(G109_p_spl_01),
    .din2(G111_p_spl_0)
  );


  FA
  g_g520_n
  (
    .dout(g520_n),
    .din1(G109_n_spl_01),
    .din2(G111_n_spl_0)
  );


  LA
  g_g521_p
  (
    .dout(g521_p),
    .din1(g519_n),
    .din2(g520_n)
  );


  FA
  g_g521_n
  (
    .dout(g521_n),
    .din1(g519_p),
    .din2(g520_p)
  );


  LA
  g_g522_p
  (
    .dout(g522_p),
    .din1(g518_n_spl_),
    .din2(g521_n_spl_)
  );


  FA
  g_g522_n
  (
    .dout(g522_n),
    .din1(g518_p_spl_),
    .din2(g521_p_spl_)
  );


  LA
  g_g523_p
  (
    .dout(g523_p),
    .din1(g518_p_spl_),
    .din2(g521_p_spl_)
  );


  FA
  g_g523_n
  (
    .dout(g523_n),
    .din1(g518_n_spl_),
    .din2(g521_n_spl_)
  );


  LA
  g_g524_p
  (
    .dout(g524_p),
    .din1(g522_n),
    .din2(g523_n)
  );


  FA
  g_g524_n
  (
    .dout(g524_n),
    .din1(g522_p),
    .din2(g523_p)
  );


  LA
  g_g525_p
  (
    .dout(g525_p),
    .din1(G105_n_spl_01),
    .din2(G107_n_spl_01)
  );


  FA
  g_g525_n
  (
    .dout(g525_n),
    .din1(G105_p_spl_01),
    .din2(G107_p_spl_01)
  );


  LA
  g_g526_p
  (
    .dout(g526_p),
    .din1(G105_p_spl_01),
    .din2(G107_p_spl_01)
  );


  FA
  g_g526_n
  (
    .dout(g526_n),
    .din1(G105_n_spl_01),
    .din2(G107_n_spl_01)
  );


  LA
  g_g527_p
  (
    .dout(g527_p),
    .din1(g525_n),
    .din2(g526_n)
  );


  FA
  g_g527_n
  (
    .dout(g527_n),
    .din1(g525_p),
    .din2(g526_p)
  );


  LA
  g_g528_p
  (
    .dout(g528_p),
    .din1(g524_n_spl_),
    .din2(g527_n_spl_)
  );


  FA
  g_g528_n
  (
    .dout(g528_n),
    .din1(g524_p_spl_),
    .din2(g527_p_spl_)
  );


  LA
  g_g529_p
  (
    .dout(g529_p),
    .din1(g524_p_spl_),
    .din2(g527_p_spl_)
  );


  FA
  g_g529_n
  (
    .dout(g529_n),
    .din1(g524_n_spl_),
    .din2(g527_n_spl_)
  );


  LA
  g_g530_p
  (
    .dout(g530_p),
    .din1(g528_n),
    .din2(g529_n)
  );


  FA
  g_g530_n
  (
    .dout(g530_n),
    .din1(g528_p),
    .din2(g529_p)
  );


  LA
  g_g531_p
  (
    .dout(g531_p),
    .din1(g515_n),
    .din2(g530_p)
  );


  LA
  g_g532_p
  (
    .dout(g532_p),
    .din1(g515_p),
    .din2(g530_n)
  );


  FA
  g_g533_n
  (
    .dout(g533_n),
    .din1(g531_p),
    .din2(g532_p)
  );


  LA
  g_g534_p
  (
    .dout(g534_p),
    .din1(g400_p_spl_00),
    .din2(g408_p_spl_0)
  );


  FA
  g_g534_n
  (
    .dout(g534_n),
    .din1(g400_n_spl_00),
    .din2(g408_n_spl_00)
  );


  LA
  g_g535_p
  (
    .dout(g535_p),
    .din1(g406_n_spl_0),
    .din2(g534_n)
  );


  FA
  g_g535_n
  (
    .dout(g535_n),
    .din1(g406_p_spl_0),
    .din2(g534_p)
  );


  LA
  g_g536_p
  (
    .dout(g536_p),
    .din1(g415_p_spl_00),
    .din2(g535_n_spl_0)
  );


  FA
  g_g536_n
  (
    .dout(g536_n),
    .din1(g415_n_spl_00),
    .din2(g535_p_spl_0)
  );


  LA
  g_g537_p
  (
    .dout(g537_p),
    .din1(g413_n_spl_),
    .din2(g536_n)
  );


  FA
  g_g537_n
  (
    .dout(g537_n),
    .din1(g413_p_spl_),
    .din2(g536_p)
  );


  LA
  g_g538_p
  (
    .dout(g538_p),
    .din1(g422_p_spl_00),
    .din2(g537_n_spl_00)
  );


  FA
  g_g538_n
  (
    .dout(g538_n),
    .din1(g422_n_spl_00),
    .din2(g537_p_spl_00)
  );


  LA
  g_g539_p
  (
    .dout(g539_p),
    .din1(g420_n_spl_0),
    .din2(g538_n)
  );


  FA
  g_g539_n
  (
    .dout(g539_n),
    .din1(g420_p_spl_0),
    .din2(g538_p)
  );


  LA
  g_g540_p
  (
    .dout(g540_p),
    .din1(g429_p_spl_00),
    .din2(g539_n_spl_0)
  );


  FA
  g_g540_n
  (
    .dout(g540_n),
    .din1(g429_n_spl_00),
    .din2(g539_p_spl_0)
  );


  LA
  g_g541_p
  (
    .dout(g541_p),
    .din1(g427_n_spl_),
    .din2(g540_n)
  );


  FA
  g_g541_n
  (
    .dout(g541_n),
    .din1(g427_p_spl_),
    .din2(g540_p)
  );


  FA
  g_g542_n
  (
    .dout(g542_n),
    .din1(g396_n_spl_),
    .din2(g541_p_spl_00)
  );


  LA
  g_g543_p
  (
    .dout(g543_p),
    .din1(g373_p_spl_0),
    .din2(g381_p_spl_00)
  );


  FA
  g_g543_n
  (
    .dout(g543_n),
    .din1(g373_n_spl_0),
    .din2(g381_n_spl_00)
  );


  LA
  g_g544_p
  (
    .dout(g544_p),
    .din1(g379_n_spl_),
    .din2(g543_n)
  );


  FA
  g_g544_n
  (
    .dout(g544_n),
    .din1(g379_p_spl_),
    .din2(g543_p)
  );


  LA
  g_g545_p
  (
    .dout(g545_p),
    .din1(g387_n_spl_),
    .din2(g544_n_spl_0)
  );


  FA
  g_g545_n
  (
    .dout(g545_n),
    .din1(g387_p_spl_),
    .din2(g544_p_spl_0)
  );


  LA
  g_g546_p
  (
    .dout(g546_p),
    .din1(g386_n_spl_),
    .din2(g545_n_spl_)
  );


  FA
  g_g546_n
  (
    .dout(g546_n),
    .din1(g386_p_spl_),
    .din2(g545_p_spl_)
  );


  FA
  g_g547_n
  (
    .dout(g547_n),
    .din1(g395_n_spl_00),
    .din2(g546_p_spl_0)
  );


  LA
  g_g548_p
  (
    .dout(g548_p),
    .din1(g542_n),
    .din2(g547_n)
  );


  LA
  g_g549_p
  (
    .dout(g549_p),
    .din1(g393_n_spl_),
    .din2(g548_p)
  );


  FA
  g_g550_n
  (
    .dout(g550_n),
    .din1(g476_p_spl_00),
    .din2(g480_p_spl_0)
  );


  FA
  g_g551_n
  (
    .dout(g551_n),
    .din1(G21_n),
    .din2(g464_p_spl_00)
  );


  FA
  g_g552_n
  (
    .dout(g552_n),
    .din1(G21_p),
    .din2(g464_n_spl_00)
  );


  LA
  g_g553_p
  (
    .dout(g553_p),
    .din1(g551_n),
    .din2(g552_n)
  );


  LA
  g_g554_p
  (
    .dout(g554_p),
    .din1(G177_p_spl_0000),
    .din2(g553_p_spl_)
  );


  FA
  g_g555_n
  (
    .dout(g555_n),
    .din1(G176_p_spl_00000),
    .din2(g554_p)
  );


  FA
  g_g556_n
  (
    .dout(g556_n),
    .din1(G177_n_spl_0000),
    .din2(g245_n_spl_0)
  );


  FA
  g_g557_n
  (
    .dout(g557_n),
    .din1(G176_n_spl_0000),
    .din2(g556_n)
  );


  FA
  g_g558_n
  (
    .dout(g558_n),
    .din1(G60_p),
    .din2(G177_p_spl_0000)
  );


  LA
  g_g559_p
  (
    .dout(g559_p),
    .din1(g557_n),
    .din2(g558_n)
  );


  LA
  g_g560_p
  (
    .dout(g560_p),
    .din1(g555_n),
    .din2(g559_p)
  );


  LA
  g_g561_p
  (
    .dout(g561_p),
    .din1(g461_n_spl_0),
    .din2(g464_p_spl_01)
  );


  FA
  g_g561_n
  (
    .dout(g561_n),
    .din1(g461_p_spl_0),
    .din2(g464_n_spl_01)
  );


  LA
  g_g562_p
  (
    .dout(g562_p),
    .din1(g465_n_spl_0),
    .din2(g561_n)
  );


  FA
  g_g562_n
  (
    .dout(g562_n),
    .din1(g465_p_spl_0),
    .din2(g561_p)
  );


  LA
  g_g563_p
  (
    .dout(g563_p),
    .din1(G177_p_spl_0001),
    .din2(g562_n_spl_0)
  );


  FA
  g_g564_n
  (
    .dout(g564_n),
    .din1(G176_p_spl_00000),
    .din2(g563_p)
  );


  FA
  g_g565_n
  (
    .dout(g565_n),
    .din1(G177_n_spl_0000),
    .din2(g224_n_spl_)
  );


  FA
  g_g566_n
  (
    .dout(g566_n),
    .din1(G176_n_spl_0000),
    .din2(g565_n)
  );


  FA
  g_g567_n
  (
    .dout(g567_n),
    .din1(G58_p),
    .din2(G177_p_spl_0001)
  );


  LA
  g_g568_p
  (
    .dout(g568_p),
    .din1(g566_n),
    .din2(g567_n)
  );


  LA
  g_g569_p
  (
    .dout(g569_p),
    .din1(g564_n),
    .din2(g568_p)
  );


  LA
  g_g570_p
  (
    .dout(g570_p),
    .din1(G2_p_spl_0),
    .din2(g402_p_spl_0)
  );


  FA
  g_g570_n
  (
    .dout(g570_n),
    .din1(G2_n_spl_0),
    .din2(g402_n_spl_0)
  );


  FA
  g_g571_n
  (
    .dout(g571_n),
    .din1(G2_p_spl_0),
    .din2(g402_p_spl_1)
  );


  LA
  g_g572_p
  (
    .dout(g572_p),
    .din1(g570_n_spl_),
    .din2(g571_n)
  );


  LA
  g_g573_p
  (
    .dout(g573_p),
    .din1(G177_p_spl_0010),
    .din2(g572_p_spl_)
  );


  FA
  g_g574_n
  (
    .dout(g574_n),
    .din1(G176_p_spl_00001),
    .din2(g573_p)
  );


  FA
  g_g575_n
  (
    .dout(g575_n),
    .din1(G177_n_spl_0001),
    .din2(g308_n_spl_)
  );


  FA
  g_g576_n
  (
    .dout(g576_n),
    .din1(G176_n_spl_0001),
    .din2(g575_n)
  );


  FA
  g_g577_n
  (
    .dout(g577_n),
    .din1(G48_p),
    .din2(G177_p_spl_0010)
  );


  LA
  g_g578_p
  (
    .dout(g578_p),
    .din1(g576_n),
    .din2(g577_n)
  );


  LA
  g_g579_p
  (
    .dout(g579_p),
    .din1(g574_n),
    .din2(g578_p)
  );


  LA
  g_g580_p
  (
    .dout(g580_p),
    .din1(g476_p_spl_0),
    .din2(g479_p_spl_00)
  );


  FA
  g_g580_n
  (
    .dout(g580_n),
    .din1(g476_n_spl_0),
    .din2(g479_n_spl_00)
  );


  LA
  g_g581_p
  (
    .dout(g581_p),
    .din1(g480_n),
    .din2(g580_n)
  );


  FA
  g_g581_n
  (
    .dout(g581_n),
    .din1(g480_p_spl_),
    .din2(g580_p)
  );


  LA
  g_g582_p
  (
    .dout(g582_p),
    .din1(G22_p_spl_),
    .din2(G173_n_spl_0000)
  );


  LA
  g_g583_p
  (
    .dout(g583_p),
    .din1(G3_p_spl_),
    .din2(G173_p_spl_0000)
  );


  FA
  g_g584_n
  (
    .dout(g584_n),
    .din1(g582_p),
    .din2(g583_p)
  );


  LA
  g_g585_p
  (
    .dout(g585_p),
    .din1(G172_n_spl_000),
    .din2(g584_n)
  );


  FA
  g_g586_n
  (
    .dout(g586_n),
    .din1(G173_p_spl_0000),
    .din2(g579_p_spl_00)
  );


  FA
  g_g587_n
  (
    .dout(g587_n),
    .din1(G173_n_spl_0000),
    .din2(g560_p_spl_00)
  );


  LA
  g_g588_p
  (
    .dout(g588_p),
    .din1(G172_p_spl_000),
    .din2(g587_n)
  );


  LA
  g_g589_p
  (
    .dout(g589_p),
    .din1(g586_n),
    .din2(g588_p)
  );


  FA
  g_g590_n
  (
    .dout(g590_n),
    .din1(g585_p),
    .din2(g589_p)
  );


  LA
  g_g591_p
  (
    .dout(g591_p),
    .din1(G19_p),
    .din2(G177_n_spl_0001)
  );


  LA
  g_g592_p
  (
    .dout(g592_p),
    .din1(G176_p_spl_00001),
    .din2(g591_p)
  );


  LA
  g_g593_p
  (
    .dout(g593_p),
    .din1(G176_p_spl_0001),
    .din2(g277_n_spl_)
  );


  LA
  g_g594_p
  (
    .dout(g594_p),
    .din1(g459_p_spl_0),
    .din2(g471_p_spl_0)
  );


  FA
  g_g594_n
  (
    .dout(g594_n),
    .din1(g459_n_spl_0),
    .din2(g471_n_spl_00)
  );


  LA
  g_g595_p
  (
    .dout(g595_p),
    .din1(g472_n_spl_),
    .din2(g594_n_spl_)
  );


  FA
  g_g595_n
  (
    .dout(g595_n),
    .din1(g472_p_spl_),
    .din2(g594_p_spl_)
  );


  LA
  g_g596_p
  (
    .dout(g596_p),
    .din1(g469_n_spl_0),
    .din2(g595_p)
  );


  FA
  g_g596_n
  (
    .dout(g596_n),
    .din1(g469_p_spl_0),
    .din2(g595_n_spl_)
  );


  LA
  g_g597_p
  (
    .dout(g597_p),
    .din1(g454_p_spl_0),
    .din2(g596_n_spl_0)
  );


  FA
  g_g597_n
  (
    .dout(g597_n),
    .din1(g454_n_spl_00),
    .din2(g596_p_spl_0)
  );


  LA
  g_g598_p
  (
    .dout(g598_p),
    .din1(g452_n_spl_0),
    .din2(g597_n)
  );


  FA
  g_g598_n
  (
    .dout(g598_n),
    .din1(g452_p_spl_0),
    .din2(g597_p_spl_)
  );


  FA
  g_g599_n
  (
    .dout(g599_n),
    .din1(g450_p_spl_0),
    .din2(g598_p_spl_0)
  );


  FA
  g_g600_n
  (
    .dout(g600_n),
    .din1(g450_n_spl_0),
    .din2(g598_n_spl_0)
  );


  LA
  g_g601_p
  (
    .dout(g601_p),
    .din1(g599_n),
    .din2(g600_n)
  );


  LA
  g_g602_p
  (
    .dout(g602_p),
    .din1(G176_n_spl_0001),
    .din2(g601_p_spl_)
  );


  FA
  g_g603_n
  (
    .dout(g603_n),
    .din1(g593_p),
    .din2(g602_p)
  );


  LA
  g_g604_p
  (
    .dout(g604_p),
    .din1(G177_p_spl_0011),
    .din2(g603_n)
  );


  FA
  g_g605_n
  (
    .dout(g605_n),
    .din1(g592_p),
    .din2(g604_p)
  );


  LA
  g_g606_p
  (
    .dout(g606_p),
    .din1(G59_p),
    .din2(G177_n_spl_0010)
  );


  LA
  g_g607_p
  (
    .dout(g607_p),
    .din1(G176_p_spl_0001),
    .din2(g606_p)
  );


  LA
  g_g608_p
  (
    .dout(g608_p),
    .din1(G176_p_spl_0010),
    .din2(g248_n_spl_)
  );


  LA
  g_g609_p
  (
    .dout(g609_p),
    .din1(g454_n_spl_0),
    .din2(g596_p_spl_0)
  );


  FA
  g_g610_n
  (
    .dout(g610_n),
    .din1(g597_p_spl_),
    .din2(g609_p)
  );


  LA
  g_g611_p
  (
    .dout(g611_p),
    .din1(G176_n_spl_0010),
    .din2(g610_n_spl_)
  );


  FA
  g_g612_n
  (
    .dout(g612_n),
    .din1(g608_p),
    .din2(g611_p)
  );


  LA
  g_g613_p
  (
    .dout(g613_p),
    .din1(G177_p_spl_0011),
    .din2(g612_n)
  );


  FA
  g_g614_n
  (
    .dout(g614_n),
    .din1(g607_p),
    .din2(g613_p)
  );


  LA
  g_g615_p
  (
    .dout(g615_p),
    .din1(G50_p),
    .din2(G177_n_spl_0010)
  );


  LA
  g_g616_p
  (
    .dout(g616_p),
    .din1(G176_p_spl_0010),
    .din2(g615_p)
  );


  LA
  g_g617_p
  (
    .dout(g617_p),
    .din1(g459_n_spl_),
    .din2(g465_n_spl_)
  );


  FA
  g_g617_n
  (
    .dout(g617_n),
    .din1(g459_p_spl_),
    .din2(g465_p_spl_)
  );


  LA
  g_g618_p
  (
    .dout(g618_p),
    .din1(g471_n_spl_0),
    .din2(g617_p_spl_0)
  );


  FA
  g_g619_n
  (
    .dout(g619_n),
    .din1(g595_n_spl_),
    .din2(g618_p)
  );


  FA
  g_g620_n
  (
    .dout(g620_n),
    .din1(G176_p_spl_0011),
    .din2(g619_n_spl_)
  );


  FA
  g_g621_n
  (
    .dout(g621_n),
    .din1(G176_n_spl_0010),
    .din2(g233_n_spl_)
  );


  LA
  g_g622_p
  (
    .dout(g622_p),
    .din1(G177_p_spl_0100),
    .din2(g621_n)
  );


  LA
  g_g623_p
  (
    .dout(g623_p),
    .din1(g620_n),
    .din2(g622_p)
  );


  FA
  g_g624_n
  (
    .dout(g624_n),
    .din1(g616_p),
    .din2(g623_p)
  );


  LA
  g_g625_p
  (
    .dout(g625_p),
    .din1(G22_p_spl_),
    .din2(G174_n_spl_0000)
  );


  LA
  g_g626_p
  (
    .dout(g626_p),
    .din1(G3_p_spl_),
    .din2(G174_p_spl_0000)
  );


  FA
  g_g627_n
  (
    .dout(g627_n),
    .din1(g625_p),
    .din2(g626_p)
  );


  LA
  g_g628_p
  (
    .dout(g628_p),
    .din1(G175_n_spl_000),
    .din2(g627_n)
  );


  FA
  g_g629_n
  (
    .dout(g629_n),
    .din1(G174_p_spl_0000),
    .din2(g579_p_spl_00)
  );


  FA
  g_g630_n
  (
    .dout(g630_n),
    .din1(G174_n_spl_0000),
    .din2(g560_p_spl_00)
  );


  LA
  g_g631_p
  (
    .dout(g631_p),
    .din1(G175_p_spl_000),
    .din2(g630_n)
  );


  LA
  g_g632_p
  (
    .dout(g632_p),
    .din1(g629_n),
    .din2(g631_p)
  );


  FA
  g_g633_n
  (
    .dout(g633_n),
    .din1(g628_p),
    .din2(g632_p)
  );


  LA
  g_g634_p
  (
    .dout(g634_p),
    .din1(G53_p),
    .din2(G177_n_spl_0011)
  );


  LA
  g_g635_p
  (
    .dout(g635_p),
    .din1(G176_p_spl_0011),
    .din2(g634_p)
  );


  FA
  g_g636_n
  (
    .dout(g636_n),
    .din1(G176_n_spl_0011),
    .din2(g356_n_spl_)
  );


  LA
  g_g637_p
  (
    .dout(g637_p),
    .din1(G2_p_spl_1),
    .din2(g416_p_spl_0)
  );


  FA
  g_g637_n
  (
    .dout(g637_n),
    .din1(G2_n_spl_0),
    .din2(g416_n_spl_0)
  );


  LA
  g_g638_p
  (
    .dout(g638_p),
    .din1(g537_p_spl_00),
    .din2(g637_n)
  );


  FA
  g_g638_n
  (
    .dout(g638_n),
    .din1(g537_n_spl_00),
    .din2(g637_p)
  );


  LA
  g_g639_p
  (
    .dout(g639_p),
    .din1(g422_p_spl_0),
    .din2(g638_n)
  );


  FA
  g_g639_n
  (
    .dout(g639_n),
    .din1(g422_n_spl_01),
    .din2(g638_p_spl_)
  );


  LA
  g_g640_p
  (
    .dout(g640_p),
    .din1(g420_n_spl_),
    .din2(g639_n)
  );


  FA
  g_g640_n
  (
    .dout(g640_n),
    .din1(g420_p_spl_),
    .din2(g639_p_spl_)
  );


  LA
  g_g641_p
  (
    .dout(g641_p),
    .din1(g429_n_spl_01),
    .din2(g640_p)
  );


  LA
  g_g642_p
  (
    .dout(g642_p),
    .din1(g429_p_spl_01),
    .din2(g640_n)
  );


  FA
  g_g643_n
  (
    .dout(g643_n),
    .din1(g641_p),
    .din2(g642_p)
  );


  FA
  g_g644_n
  (
    .dout(g644_n),
    .din1(G176_p_spl_0100),
    .din2(g643_n_spl_)
  );


  LA
  g_g645_p
  (
    .dout(g645_p),
    .din1(G177_p_spl_0100),
    .din2(g644_n)
  );


  LA
  g_g646_p
  (
    .dout(g646_p),
    .din1(g636_n),
    .din2(g645_p)
  );


  FA
  g_g647_n
  (
    .dout(g647_n),
    .din1(g635_p),
    .din2(g646_p)
  );


  LA
  g_g648_p
  (
    .dout(g648_p),
    .din1(G57_p),
    .din2(G177_n_spl_0011)
  );


  LA
  g_g649_p
  (
    .dout(g649_p),
    .din1(G176_p_spl_0100),
    .din2(g648_p)
  );


  LA
  g_g650_p
  (
    .dout(g650_p),
    .din1(G176_p_spl_0101),
    .din2(g365_n_spl_)
  );


  LA
  g_g651_p
  (
    .dout(g651_p),
    .din1(g422_n_spl_01),
    .din2(g638_p_spl_)
  );


  FA
  g_g652_n
  (
    .dout(g652_n),
    .din1(g639_p_spl_),
    .din2(g651_p)
  );


  LA
  g_g653_p
  (
    .dout(g653_p),
    .din1(G176_n_spl_0011),
    .din2(g652_n_spl_)
  );


  FA
  g_g654_n
  (
    .dout(g654_n),
    .din1(g650_p),
    .din2(g653_p)
  );


  LA
  g_g655_p
  (
    .dout(g655_p),
    .din1(G177_p_spl_0101),
    .din2(g654_n)
  );


  FA
  g_g656_n
  (
    .dout(g656_n),
    .din1(g649_p),
    .din2(g655_p)
  );


  LA
  g_g657_p
  (
    .dout(g657_p),
    .din1(G56_p),
    .din2(G177_n_spl_010)
  );


  LA
  g_g658_p
  (
    .dout(g658_p),
    .din1(G176_p_spl_0101),
    .din2(g657_p)
  );


  LA
  g_g659_p
  (
    .dout(g659_p),
    .din1(g400_n_spl_0),
    .din2(g570_n_spl_)
  );


  FA
  g_g659_n
  (
    .dout(g659_n),
    .din1(g400_p_spl_0),
    .din2(g570_p)
  );


  LA
  g_g660_p
  (
    .dout(g660_p),
    .din1(g408_p_spl_1),
    .din2(g659_n)
  );


  FA
  g_g660_n
  (
    .dout(g660_n),
    .din1(g408_n_spl_0),
    .din2(g659_p_spl_)
  );


  LA
  g_g661_p
  (
    .dout(g661_p),
    .din1(g406_n_spl_),
    .din2(g660_n)
  );


  FA
  g_g661_n
  (
    .dout(g661_n),
    .din1(g406_p_spl_),
    .din2(g660_p_spl_)
  );


  LA
  g_g662_p
  (
    .dout(g662_p),
    .din1(g415_n_spl_0),
    .din2(g661_p)
  );


  LA
  g_g663_p
  (
    .dout(g663_p),
    .din1(g415_p_spl_0),
    .din2(g661_n)
  );


  FA
  g_g664_n
  (
    .dout(g664_n),
    .din1(g662_p),
    .din2(g663_p)
  );


  FA
  g_g665_n
  (
    .dout(g665_n),
    .din1(G176_p_spl_0110),
    .din2(g664_n_spl_)
  );


  FA
  g_g666_n
  (
    .dout(g666_n),
    .din1(G176_n_spl_0100),
    .din2(g298_n_spl_)
  );


  LA
  g_g667_p
  (
    .dout(g667_p),
    .din1(G177_p_spl_0101),
    .din2(g666_n)
  );


  LA
  g_g668_p
  (
    .dout(g668_p),
    .din1(g665_n),
    .din2(g667_p)
  );


  FA
  g_g669_n
  (
    .dout(g669_n),
    .din1(g658_p),
    .din2(g668_p)
  );


  LA
  g_g670_p
  (
    .dout(g670_p),
    .din1(G55_p),
    .din2(G177_n_spl_010)
  );


  LA
  g_g671_p
  (
    .dout(g671_p),
    .din1(G176_p_spl_0110),
    .din2(g670_p)
  );


  LA
  g_g672_p
  (
    .dout(g672_p),
    .din1(g408_n_spl_1),
    .din2(g659_p_spl_)
  );


  FA
  g_g673_n
  (
    .dout(g673_n),
    .din1(g660_p_spl_),
    .din2(g672_p)
  );


  FA
  g_g674_n
  (
    .dout(g674_n),
    .din1(G176_p_spl_0111),
    .din2(g673_n_spl_)
  );


  FA
  g_g675_n
  (
    .dout(g675_n),
    .din1(G176_n_spl_0100),
    .din2(g289_n_spl_)
  );


  LA
  g_g676_p
  (
    .dout(g676_p),
    .din1(G177_p_spl_0110),
    .din2(g675_n)
  );


  LA
  g_g677_p
  (
    .dout(g677_p),
    .din1(g674_n),
    .din2(g676_p)
  );


  FA
  g_g678_n
  (
    .dout(g678_n),
    .din1(g671_p),
    .din2(g677_p)
  );


  LA
  g_g679_p
  (
    .dout(g679_p),
    .din1(g434_n_spl_1),
    .din2(g440_n_spl_1)
  );


  FA
  g_g679_n
  (
    .dout(g679_n),
    .din1(g434_p_spl_1),
    .din2(g440_p_spl_1)
  );


  LA
  g_g680_p
  (
    .dout(g680_p),
    .din1(g434_p_spl_1),
    .din2(g440_p_spl_1)
  );


  FA
  g_g680_n
  (
    .dout(g680_n),
    .din1(g434_n_spl_1),
    .din2(g440_n_spl_1)
  );


  LA
  g_g681_p
  (
    .dout(g681_p),
    .din1(g679_n),
    .din2(g680_n)
  );


  FA
  g_g681_n
  (
    .dout(g681_n),
    .din1(g679_p),
    .din2(g680_p)
  );


  LA
  g_g682_p
  (
    .dout(g682_p),
    .din1(g581_n_spl_00),
    .din2(g681_p_spl_)
  );


  FA
  g_g682_n
  (
    .dout(g682_n),
    .din1(g581_p_spl_00),
    .din2(g681_n_spl_)
  );


  LA
  g_g683_p
  (
    .dout(g683_p),
    .din1(g581_p_spl_00),
    .din2(g681_n_spl_)
  );


  FA
  g_g683_n
  (
    .dout(g683_n),
    .din1(g581_n_spl_00),
    .din2(g681_p_spl_)
  );


  LA
  g_g684_p
  (
    .dout(g684_p),
    .din1(g682_n),
    .din2(g683_n)
  );


  FA
  g_g684_n
  (
    .dout(g684_n),
    .din1(g682_p),
    .din2(g683_p)
  );


  LA
  g_g685_p
  (
    .dout(g685_p),
    .din1(G123_n_spl_111),
    .din2(G133_n)
  );


  FA
  g_g685_n
  (
    .dout(g685_n),
    .din1(G123_p_spl_111),
    .din2(G133_p)
  );


  LA
  g_g686_p
  (
    .dout(g686_p),
    .din1(G123_p_spl_111),
    .din2(G132_n_spl_)
  );


  FA
  g_g686_n
  (
    .dout(g686_n),
    .din1(G123_n_spl_111),
    .din2(G132_p_spl_)
  );


  LA
  g_g687_p
  (
    .dout(g687_p),
    .din1(g685_n),
    .din2(g686_n)
  );


  FA
  g_g687_n
  (
    .dout(g687_n),
    .din1(g685_p),
    .din2(g686_p)
  );


  LA
  g_g688_p
  (
    .dout(g688_p),
    .din1(g464_n_spl_01),
    .din2(g687_n_spl_)
  );


  FA
  g_g688_n
  (
    .dout(g688_n),
    .din1(g464_p_spl_01),
    .din2(g687_p_spl_)
  );


  LA
  g_g689_p
  (
    .dout(g689_p),
    .din1(g464_p_spl_10),
    .din2(g687_p_spl_)
  );


  FA
  g_g689_n
  (
    .dout(g689_n),
    .din1(g464_n_spl_10),
    .din2(g687_n_spl_)
  );


  LA
  g_g690_p
  (
    .dout(g690_p),
    .din1(g688_n),
    .din2(g689_n)
  );


  FA
  g_g690_n
  (
    .dout(g690_n),
    .din1(g688_p),
    .din2(g689_p)
  );


  LA
  g_g691_p
  (
    .dout(g691_p),
    .din1(g447_n_spl_1),
    .din2(g451_p_spl_1)
  );


  FA
  g_g691_n
  (
    .dout(g691_n),
    .din1(g447_p_spl_1),
    .din2(g451_n_spl_1)
  );


  LA
  g_g692_p
  (
    .dout(g692_p),
    .din1(g447_p_spl_1),
    .din2(g451_n_spl_1)
  );


  FA
  g_g692_n
  (
    .dout(g692_n),
    .din1(g447_n_spl_1),
    .din2(g451_p_spl_1)
  );


  LA
  g_g693_p
  (
    .dout(g693_p),
    .din1(g691_n),
    .din2(g692_n)
  );


  FA
  g_g693_n
  (
    .dout(g693_n),
    .din1(g691_p),
    .din2(g692_p)
  );


  LA
  g_g694_p
  (
    .dout(g694_p),
    .din1(g458_n_spl_1),
    .din2(g468_n_spl_1)
  );


  FA
  g_g694_n
  (
    .dout(g694_n),
    .din1(g458_p_spl_1),
    .din2(g468_p_spl_1)
  );


  LA
  g_g695_p
  (
    .dout(g695_p),
    .din1(g458_p_spl_1),
    .din2(g468_p_spl_1)
  );


  FA
  g_g695_n
  (
    .dout(g695_n),
    .din1(g458_n_spl_1),
    .din2(g468_n_spl_1)
  );


  LA
  g_g696_p
  (
    .dout(g696_p),
    .din1(g694_n),
    .din2(g695_n)
  );


  FA
  g_g696_n
  (
    .dout(g696_n),
    .din1(g694_p),
    .din2(g695_p)
  );


  LA
  g_g697_p
  (
    .dout(g697_p),
    .din1(g693_n_spl_),
    .din2(g696_n_spl_)
  );


  FA
  g_g697_n
  (
    .dout(g697_n),
    .din1(g693_p_spl_),
    .din2(g696_p_spl_)
  );


  LA
  g_g698_p
  (
    .dout(g698_p),
    .din1(g693_p_spl_),
    .din2(g696_p_spl_)
  );


  FA
  g_g698_n
  (
    .dout(g698_n),
    .din1(g693_n_spl_),
    .din2(g696_n_spl_)
  );


  LA
  g_g699_p
  (
    .dout(g699_p),
    .din1(g697_n),
    .din2(g698_n)
  );


  FA
  g_g699_n
  (
    .dout(g699_n),
    .din1(g697_p),
    .din2(g698_p)
  );


  LA
  g_g700_p
  (
    .dout(g700_p),
    .din1(g690_p_spl_),
    .din2(g699_n_spl_)
  );


  FA
  g_g700_n
  (
    .dout(g700_n),
    .din1(g690_n_spl_),
    .din2(g699_p_spl_)
  );


  LA
  g_g701_p
  (
    .dout(g701_p),
    .din1(g690_n_spl_),
    .din2(g699_p_spl_)
  );


  FA
  g_g701_n
  (
    .dout(g701_n),
    .din1(g690_p_spl_),
    .din2(g699_n_spl_)
  );


  LA
  g_g702_p
  (
    .dout(g702_p),
    .din1(g700_n),
    .din2(g701_n)
  );


  FA
  g_g702_n
  (
    .dout(g702_n),
    .din1(g700_p),
    .din2(g701_p)
  );


  LA
  g_g703_p
  (
    .dout(g703_p),
    .din1(g684_n),
    .din2(g702_p)
  );


  LA
  g_g704_p
  (
    .dout(g704_p),
    .din1(g684_p),
    .din2(g702_n)
  );


  FA
  g_g705_n
  (
    .dout(g705_n),
    .din1(g703_p),
    .din2(g704_p)
  );


  LA
  g_g706_p
  (
    .dout(g706_p),
    .din1(g399_n_spl_1),
    .din2(g405_n_spl_1)
  );


  FA
  g_g706_n
  (
    .dout(g706_n),
    .din1(g399_p_spl_1),
    .din2(g405_p_spl_1)
  );


  LA
  g_g707_p
  (
    .dout(g707_p),
    .din1(g399_p_spl_1),
    .din2(g405_p_spl_1)
  );


  FA
  g_g707_n
  (
    .dout(g707_n),
    .din1(g399_n_spl_1),
    .din2(g405_n_spl_1)
  );


  LA
  g_g708_p
  (
    .dout(g708_p),
    .din1(g706_n),
    .din2(g707_n)
  );


  FA
  g_g708_n
  (
    .dout(g708_n),
    .din1(g706_p),
    .din2(g707_p)
  );


  LA
  g_g709_p
  (
    .dout(g709_p),
    .din1(g412_n_spl_1),
    .din2(g419_n_spl_1)
  );


  FA
  g_g709_n
  (
    .dout(g709_n),
    .din1(g412_p_spl_1),
    .din2(g419_p_spl_1)
  );


  LA
  g_g710_p
  (
    .dout(g710_p),
    .din1(g412_p_spl_1),
    .din2(g419_p_spl_1)
  );


  FA
  g_g710_n
  (
    .dout(g710_n),
    .din1(g412_n_spl_1),
    .din2(g419_n_spl_1)
  );


  LA
  g_g711_p
  (
    .dout(g711_p),
    .din1(g709_n),
    .din2(g710_n)
  );


  FA
  g_g711_n
  (
    .dout(g711_n),
    .din1(g709_p),
    .din2(g710_p)
  );


  LA
  g_g712_p
  (
    .dout(g712_p),
    .din1(g708_p_spl_),
    .din2(g711_n_spl_)
  );


  FA
  g_g712_n
  (
    .dout(g712_n),
    .din1(g708_n_spl_),
    .din2(g711_p_spl_)
  );


  LA
  g_g713_p
  (
    .dout(g713_p),
    .din1(g708_n_spl_),
    .din2(g711_p_spl_)
  );


  FA
  g_g713_n
  (
    .dout(g713_n),
    .din1(g708_p_spl_),
    .din2(g711_n_spl_)
  );


  LA
  g_g714_p
  (
    .dout(g714_p),
    .din1(g712_n),
    .din2(g713_n)
  );


  FA
  g_g714_n
  (
    .dout(g714_n),
    .din1(g712_p),
    .din2(g713_p)
  );


  LA
  g_g715_p
  (
    .dout(g715_p),
    .din1(G112_n),
    .din2(G124_n_spl_111)
  );


  FA
  g_g715_n
  (
    .dout(g715_n),
    .din1(G112_p),
    .din2(G124_p_spl_111)
  );


  LA
  g_g716_p
  (
    .dout(g716_p),
    .din1(G111_n_spl_),
    .din2(G124_p_spl_111)
  );


  FA
  g_g716_n
  (
    .dout(g716_n),
    .din1(G111_p_spl_),
    .din2(G124_n_spl_111)
  );


  LA
  g_g717_p
  (
    .dout(g717_p),
    .din1(g715_n),
    .din2(g716_n)
  );


  FA
  g_g717_n
  (
    .dout(g717_n),
    .din1(g715_p),
    .din2(g716_p)
  );


  LA
  g_g718_p
  (
    .dout(g718_p),
    .din1(g392_n_spl_1),
    .din2(g717_n_spl_)
  );


  FA
  g_g718_n
  (
    .dout(g718_n),
    .din1(g392_p_spl_1),
    .din2(g717_p_spl_)
  );


  LA
  g_g719_p
  (
    .dout(g719_p),
    .din1(g392_p_spl_1),
    .din2(g717_p_spl_)
  );


  FA
  g_g719_n
  (
    .dout(g719_n),
    .din1(g392_n_spl_1),
    .din2(g717_n_spl_)
  );


  LA
  g_g720_p
  (
    .dout(g720_p),
    .din1(g718_n),
    .din2(g719_n)
  );


  FA
  g_g720_n
  (
    .dout(g720_n),
    .din1(g718_p),
    .din2(g719_p)
  );


  LA
  g_g721_p
  (
    .dout(g721_p),
    .din1(g372_n_spl_1),
    .din2(g426_n_spl_1)
  );


  FA
  g_g721_n
  (
    .dout(g721_n),
    .din1(g372_p_spl_1),
    .din2(g426_p_spl_1)
  );


  LA
  g_g722_p
  (
    .dout(g722_p),
    .din1(g372_p_spl_1),
    .din2(g426_p_spl_1)
  );


  FA
  g_g722_n
  (
    .dout(g722_n),
    .din1(g372_n_spl_1),
    .din2(g426_n_spl_1)
  );


  LA
  g_g723_p
  (
    .dout(g723_p),
    .din1(g721_n),
    .din2(g722_n)
  );


  FA
  g_g723_n
  (
    .dout(g723_n),
    .din1(g721_p),
    .din2(g722_p)
  );


  LA
  g_g724_p
  (
    .dout(g724_p),
    .din1(g720_p_spl_),
    .din2(g723_n_spl_)
  );


  FA
  g_g724_n
  (
    .dout(g724_n),
    .din1(g720_n_spl_),
    .din2(g723_p_spl_)
  );


  LA
  g_g725_p
  (
    .dout(g725_p),
    .din1(g720_n_spl_),
    .din2(g723_p_spl_)
  );


  FA
  g_g725_n
  (
    .dout(g725_n),
    .din1(g720_p_spl_),
    .din2(g723_n_spl_)
  );


  LA
  g_g726_p
  (
    .dout(g726_p),
    .din1(g724_n),
    .din2(g725_n)
  );


  FA
  g_g726_n
  (
    .dout(g726_n),
    .din1(g724_p),
    .din2(g725_p)
  );


  LA
  g_g727_p
  (
    .dout(g727_p),
    .din1(g378_n_spl_1),
    .din2(g385_n_spl_1)
  );


  FA
  g_g727_n
  (
    .dout(g727_n),
    .din1(g378_p_spl_1),
    .din2(g385_p_spl_1)
  );


  LA
  g_g728_p
  (
    .dout(g728_p),
    .din1(g378_p_spl_1),
    .din2(g385_p_spl_1)
  );


  FA
  g_g728_n
  (
    .dout(g728_n),
    .din1(g378_n_spl_1),
    .din2(g385_n_spl_1)
  );


  LA
  g_g729_p
  (
    .dout(g729_p),
    .din1(g727_n),
    .din2(g728_n)
  );


  FA
  g_g729_n
  (
    .dout(g729_n),
    .din1(g727_p),
    .din2(g728_p)
  );


  LA
  g_g730_p
  (
    .dout(g730_p),
    .din1(g726_n_spl_),
    .din2(g729_n_spl_)
  );


  FA
  g_g730_n
  (
    .dout(g730_n),
    .din1(g726_p_spl_),
    .din2(g729_p_spl_)
  );


  LA
  g_g731_p
  (
    .dout(g731_p),
    .din1(g726_p_spl_),
    .din2(g729_p_spl_)
  );


  FA
  g_g731_n
  (
    .dout(g731_n),
    .din1(g726_n_spl_),
    .din2(g729_n_spl_)
  );


  LA
  g_g732_p
  (
    .dout(g732_p),
    .din1(g730_n),
    .din2(g731_n)
  );


  FA
  g_g732_n
  (
    .dout(g732_n),
    .din1(g730_p),
    .din2(g731_p)
  );


  LA
  g_g733_p
  (
    .dout(g733_p),
    .din1(g714_n),
    .din2(g732_p)
  );


  LA
  g_g734_p
  (
    .dout(g734_p),
    .din1(g714_p),
    .din2(g732_n)
  );


  FA
  g_g735_n
  (
    .dout(g735_n),
    .din1(g733_p),
    .din2(g734_p)
  );


  LA
  g_g736_p
  (
    .dout(g736_p),
    .din1(G2_p_spl_1),
    .din2(g430_p_spl_0)
  );


  FA
  g_g736_n
  (
    .dout(g736_n),
    .din1(G2_n_spl_),
    .din2(g430_n_spl_0)
  );


  LA
  g_g737_p
  (
    .dout(g737_p),
    .din1(g541_p_spl_00),
    .din2(g736_n)
  );


  FA
  g_g737_n
  (
    .dout(g737_n),
    .din1(g541_n_spl_0),
    .din2(g736_p)
  );


  LA
  g_g738_p
  (
    .dout(g738_p),
    .din1(g373_p_spl_),
    .din2(g737_p_spl_00)
  );


  FA
  g_g738_n
  (
    .dout(g738_n),
    .din1(g373_n_spl_),
    .din2(g737_n_spl_00)
  );


  LA
  g_g739_p
  (
    .dout(g739_p),
    .din1(g374_p_spl_0),
    .din2(g737_n_spl_00)
  );


  FA
  g_g739_n
  (
    .dout(g739_n),
    .din1(g374_n_spl_0),
    .din2(g737_p_spl_00)
  );


  LA
  g_g740_p
  (
    .dout(g740_p),
    .din1(g738_n),
    .din2(g739_n)
  );


  FA
  g_g740_n
  (
    .dout(g740_n),
    .din1(g738_p),
    .din2(g739_p)
  );


  FA
  g_g741_n
  (
    .dout(g741_n),
    .din1(g381_n_spl_01),
    .din2(g740_p)
  );


  FA
  g_g742_n
  (
    .dout(g742_n),
    .din1(g381_p_spl_01),
    .din2(g740_n)
  );


  LA
  g_g743_p
  (
    .dout(g743_p),
    .din1(g741_n),
    .din2(g742_n)
  );


  FA
  g_g744_n
  (
    .dout(g744_n),
    .din1(g664_n_spl_),
    .din2(g743_p_spl_)
  );


  FA
  g_g745_n
  (
    .dout(g745_n),
    .din1(g375_n_spl_00),
    .din2(g737_p_spl_0)
  );


  FA
  g_g746_n
  (
    .dout(g746_n),
    .din1(g375_p_spl_00),
    .din2(g737_n_spl_0)
  );


  LA
  g_g747_p
  (
    .dout(g747_p),
    .din1(g745_n),
    .din2(g746_n)
  );


  FA
  g_g748_n
  (
    .dout(g748_n),
    .din1(g572_p_spl_),
    .din2(g747_p_spl_)
  );


  FA
  g_g749_n
  (
    .dout(g749_n),
    .din1(g744_n),
    .din2(g748_n)
  );


  FA
  g_g750_n
  (
    .dout(g750_n),
    .din1(g643_n_spl_),
    .din2(g652_n_spl_)
  );


  LA
  g_g751_p
  (
    .dout(g751_p),
    .din1(g382_p_spl_),
    .din2(g737_n_spl_1)
  );


  FA
  g_g751_n
  (
    .dout(g751_n),
    .din1(g382_n_spl_),
    .din2(g737_p_spl_1)
  );


  LA
  g_g752_p
  (
    .dout(g752_p),
    .din1(g544_p_spl_0),
    .din2(g751_n)
  );


  FA
  g_g752_n
  (
    .dout(g752_n),
    .din1(g544_n_spl_0),
    .din2(g751_p)
  );


  FA
  g_g753_n
  (
    .dout(g753_n),
    .din1(g388_n_spl_00),
    .din2(g752_n)
  );


  FA
  g_g754_n
  (
    .dout(g754_n),
    .din1(g388_p_spl_00),
    .din2(g752_p)
  );


  LA
  g_g755_p
  (
    .dout(g755_p),
    .din1(g753_n),
    .din2(g754_n)
  );


  LA
  g_g756_p
  (
    .dout(g756_p),
    .din1(g389_p_spl_),
    .din2(g737_n_spl_1)
  );


  FA
  g_g756_n
  (
    .dout(g756_n),
    .din1(g389_n_spl_0),
    .din2(g737_p_spl_1)
  );


  LA
  g_g757_p
  (
    .dout(g757_p),
    .din1(g546_p_spl_0),
    .din2(g756_n)
  );


  FA
  g_g757_n
  (
    .dout(g757_n),
    .din1(g546_n_spl_0),
    .din2(g756_p)
  );


  FA
  g_g758_n
  (
    .dout(g758_n),
    .din1(g395_n_spl_01),
    .din2(g757_n)
  );


  FA
  g_g759_n
  (
    .dout(g759_n),
    .din1(g395_p_spl_00),
    .din2(g757_p)
  );


  LA
  g_g760_p
  (
    .dout(g760_p),
    .din1(g758_n),
    .din2(g759_n)
  );


  FA
  g_g761_n
  (
    .dout(g761_n),
    .din1(g755_p_spl_),
    .din2(g760_p_spl_)
  );


  FA
  g_g762_n
  (
    .dout(g762_n),
    .din1(g673_n_spl_),
    .din2(g761_n)
  );


  FA
  g_g763_n
  (
    .dout(g763_n),
    .din1(g750_n),
    .din2(g762_n)
  );


  FA
  g_g764_n
  (
    .dout(g764_n),
    .din1(g749_n),
    .din2(g763_n)
  );


  FA
  g_g765_n
  (
    .dout(g765_n),
    .din1(g601_p_spl_),
    .din2(g619_n_spl_)
  );


  FA
  g_g766_n
  (
    .dout(g766_n),
    .din1(g553_p_spl_),
    .din2(g581_n_spl_01)
  );


  FA
  g_g767_n
  (
    .dout(g767_n),
    .din1(g610_n_spl_),
    .din2(g766_n)
  );


  FA
  g_g768_n
  (
    .dout(g768_n),
    .din1(g765_n),
    .din2(g767_n)
  );


  LA
  g_g769_p
  (
    .dout(g769_p),
    .din1(g469_n_spl_),
    .din2(g594_n_spl_)
  );


  FA
  g_g769_n
  (
    .dout(g769_n),
    .din1(g469_p_spl_),
    .din2(g594_p_spl_)
  );


  LA
  g_g770_p
  (
    .dout(g770_p),
    .din1(g454_p_spl_1),
    .din2(g769_n)
  );


  FA
  g_g770_n
  (
    .dout(g770_n),
    .din1(g454_n_spl_1),
    .din2(g769_p)
  );


  LA
  g_g771_p
  (
    .dout(g771_p),
    .din1(g452_n_spl_),
    .din2(g770_n)
  );


  FA
  g_g771_n
  (
    .dout(g771_n),
    .din1(g452_p_spl_),
    .din2(g770_p)
  );


  LA
  g_g772_p
  (
    .dout(g772_p),
    .din1(g450_p_spl_1),
    .din2(g771_n)
  );


  FA
  g_g772_n
  (
    .dout(g772_n),
    .din1(g450_n_spl_1),
    .din2(g771_p)
  );


  LA
  g_g773_p
  (
    .dout(g773_p),
    .din1(g473_n),
    .din2(g772_n)
  );


  FA
  g_g773_n
  (
    .dout(g773_n),
    .din1(g473_p_spl_),
    .din2(g772_p)
  );


  LA
  g_g774_p
  (
    .dout(g774_p),
    .din1(g448_n_spl_),
    .din2(g773_p)
  );


  FA
  g_g774_n
  (
    .dout(g774_n),
    .din1(g448_p_spl_),
    .din2(g773_n)
  );


  FA
  g_g775_n
  (
    .dout(g775_n),
    .din1(g443_n_spl_00),
    .din2(g774_p_spl_00)
  );


  FA
  g_g776_n
  (
    .dout(g776_n),
    .din1(g443_p_spl_00),
    .din2(g774_n_spl_00)
  );


  LA
  g_g777_p
  (
    .dout(g777_p),
    .din1(g775_n),
    .din2(g776_n)
  );


  FA
  g_g778_n
  (
    .dout(g778_n),
    .din1(g562_n_spl_0),
    .din2(g777_p_spl_)
  );


  LA
  g_g779_p
  (
    .dout(g779_p),
    .din1(g437_p_spl_00),
    .din2(g441_p_spl_00)
  );


  FA
  g_g779_n
  (
    .dout(g779_n),
    .din1(g437_n_spl_00),
    .din2(g441_n_spl_00)
  );


  LA
  g_g780_p
  (
    .dout(g780_p),
    .din1(g435_n_spl_),
    .din2(g779_n)
  );


  FA
  g_g780_n
  (
    .dout(g780_n),
    .din1(g435_p_spl_),
    .din2(g779_p)
  );


  LA
  g_g781_p
  (
    .dout(g781_p),
    .din1(g444_p_spl_0),
    .din2(g774_n_spl_00)
  );


  FA
  g_g781_n
  (
    .dout(g781_n),
    .din1(g444_n_spl_),
    .din2(g774_p_spl_00)
  );


  LA
  g_g782_p
  (
    .dout(g782_p),
    .din1(g780_p_spl_0),
    .din2(g781_n)
  );


  FA
  g_g782_n
  (
    .dout(g782_n),
    .din1(g780_n_spl_0),
    .din2(g781_p)
  );


  FA
  g_g783_n
  (
    .dout(g783_n),
    .din1(g479_p_spl_01),
    .din2(g782_n)
  );


  FA
  g_g784_n
  (
    .dout(g784_n),
    .din1(g479_n_spl_01),
    .din2(g782_p)
  );


  LA
  g_g785_p
  (
    .dout(g785_p),
    .din1(g783_n),
    .din2(g784_n)
  );


  LA
  g_g786_p
  (
    .dout(g786_p),
    .din1(g441_p_spl_0),
    .din2(g774_p_spl_01)
  );


  FA
  g_g786_n
  (
    .dout(g786_n),
    .din1(g441_n_spl_0),
    .din2(g774_n_spl_01)
  );


  LA
  g_g787_p
  (
    .dout(g787_p),
    .din1(g442_p_spl_0),
    .din2(g774_n_spl_01)
  );


  FA
  g_g787_n
  (
    .dout(g787_n),
    .din1(g442_n_spl_0),
    .din2(g774_p_spl_01)
  );


  LA
  g_g788_p
  (
    .dout(g788_p),
    .din1(g786_n),
    .din2(g787_n)
  );


  FA
  g_g788_n
  (
    .dout(g788_n),
    .din1(g786_p),
    .din2(g787_p)
  );


  FA
  g_g789_n
  (
    .dout(g789_n),
    .din1(g437_n_spl_01),
    .din2(g788_p)
  );


  FA
  g_g790_n
  (
    .dout(g790_n),
    .din1(g437_p_spl_01),
    .din2(g788_n)
  );


  LA
  g_g791_p
  (
    .dout(g791_p),
    .din1(g789_n),
    .din2(g790_n)
  );


  FA
  g_g792_n
  (
    .dout(g792_n),
    .din1(g785_p_spl_),
    .din2(g791_p_spl_)
  );


  FA
  g_g793_n
  (
    .dout(g793_n),
    .din1(g778_n),
    .din2(g792_n)
  );


  FA
  g_g794_n
  (
    .dout(g794_n),
    .din1(g768_n),
    .din2(g793_n)
  );


  LA
  g_g795_p
  (
    .dout(g795_p),
    .din1(G81_p_spl_),
    .din2(G158_n_spl_0000)
  );


  LA
  g_g796_p
  (
    .dout(g796_p),
    .din1(G80_p_spl_),
    .din2(G158_p_spl_0000)
  );


  FA
  g_g797_n
  (
    .dout(g797_n),
    .din1(g795_p),
    .din2(g796_p)
  );


  LA
  g_g798_p
  (
    .dout(g798_p),
    .din1(G159_n_spl_000),
    .din2(g797_n)
  );


  LA
  g_g799_p
  (
    .dout(g799_p),
    .din1(G158_p_spl_0000),
    .din2(g560_p_spl_0)
  );


  LA
  g_g800_p
  (
    .dout(g800_p),
    .din1(G158_n_spl_0000),
    .din2(g579_p_spl_0)
  );


  FA
  g_g801_n
  (
    .dout(g801_n),
    .din1(g799_p),
    .din2(g800_p)
  );


  LA
  g_g802_p
  (
    .dout(g802_p),
    .din1(G159_p_spl_000),
    .din2(g801_n)
  );


  FA
  g_g803_n
  (
    .dout(g803_n),
    .din1(g798_p),
    .din2(g802_p)
  );


  LA
  g_g804_p
  (
    .dout(g804_p),
    .din1(G64_p_spl_0000),
    .din2(g803_n)
  );


  LA
  g_g805_p
  (
    .dout(g805_p),
    .din1(G81_p_spl_),
    .din2(G160_n_spl_0000)
  );


  LA
  g_g806_p
  (
    .dout(g806_p),
    .din1(G80_p_spl_),
    .din2(G160_p_spl_0000)
  );


  FA
  g_g807_n
  (
    .dout(g807_n),
    .din1(g805_p),
    .din2(g806_p)
  );


  LA
  g_g808_p
  (
    .dout(g808_p),
    .din1(G161_n_spl_000),
    .din2(g807_n)
  );


  LA
  g_g809_p
  (
    .dout(g809_p),
    .din1(G160_p_spl_0000),
    .din2(g560_p_spl_1)
  );


  LA
  g_g810_p
  (
    .dout(g810_p),
    .din1(G160_n_spl_0000),
    .din2(g579_p_spl_1)
  );


  FA
  g_g811_n
  (
    .dout(g811_n),
    .din1(g809_p),
    .din2(g810_p)
  );


  LA
  g_g812_p
  (
    .dout(g812_p),
    .din1(G161_p_spl_000),
    .din2(g811_n)
  );


  FA
  g_g813_n
  (
    .dout(g813_n),
    .din1(g808_p),
    .din2(g812_p)
  );


  LA
  g_g814_p
  (
    .dout(g814_p),
    .din1(G64_p_spl_0000),
    .din2(g813_n)
  );


  LA
  g_g815_p
  (
    .dout(g815_p),
    .din1(G14_p_spl_),
    .din2(G173_n_spl_0001)
  );


  LA
  g_g816_p
  (
    .dout(g816_p),
    .din1(G16_p_spl_),
    .din2(G173_p_spl_0001)
  );


  FA
  g_g817_n
  (
    .dout(g817_n),
    .din1(g815_p),
    .din2(g816_p)
  );


  LA
  g_g818_p
  (
    .dout(g818_p),
    .din1(G172_n_spl_000),
    .din2(g817_n)
  );


  FA
  g_g819_n
  (
    .dout(g819_n),
    .din1(G173_p_spl_0001),
    .din2(g647_n_spl_00)
  );


  FA
  g_g820_n
  (
    .dout(g820_n),
    .din1(G173_n_spl_0001),
    .din2(g605_n_spl_00)
  );


  LA
  g_g821_p
  (
    .dout(g821_p),
    .din1(G172_p_spl_000),
    .din2(g820_n)
  );


  LA
  g_g822_p
  (
    .dout(g822_p),
    .din1(g819_n),
    .din2(g821_p)
  );


  FA
  g_g823_n
  (
    .dout(g823_n),
    .din1(g818_p),
    .din2(g822_p)
  );


  LA
  g_g824_p
  (
    .dout(g824_p),
    .din1(G6_p_spl_),
    .din2(G173_n_spl_0010)
  );


  LA
  g_g825_p
  (
    .dout(g825_p),
    .din1(G27_p_spl_),
    .din2(G173_p_spl_0010)
  );


  FA
  g_g826_n
  (
    .dout(g826_n),
    .din1(g824_p),
    .din2(g825_p)
  );


  LA
  g_g827_p
  (
    .dout(g827_p),
    .din1(G172_n_spl_001),
    .din2(g826_n)
  );


  FA
  g_g828_n
  (
    .dout(g828_n),
    .din1(G173_p_spl_0010),
    .din2(g656_n_spl_00)
  );


  FA
  g_g829_n
  (
    .dout(g829_n),
    .din1(G173_n_spl_0010),
    .din2(g614_n_spl_00)
  );


  LA
  g_g830_p
  (
    .dout(g830_p),
    .din1(G172_p_spl_001),
    .din2(g829_n)
  );


  LA
  g_g831_p
  (
    .dout(g831_p),
    .din1(g828_n),
    .din2(g830_p)
  );


  FA
  g_g832_n
  (
    .dout(g832_n),
    .din1(g827_p),
    .din2(g831_p)
  );


  LA
  g_g833_p
  (
    .dout(g833_p),
    .din1(G5_p_spl_),
    .din2(G173_n_spl_0011)
  );


  LA
  g_g834_p
  (
    .dout(g834_p),
    .din1(G26_p_spl_),
    .din2(G173_p_spl_0011)
  );


  FA
  g_g835_n
  (
    .dout(g835_n),
    .din1(g833_p),
    .din2(g834_p)
  );


  LA
  g_g836_p
  (
    .dout(g836_p),
    .din1(G172_n_spl_001),
    .din2(g835_n)
  );


  FA
  g_g837_n
  (
    .dout(g837_n),
    .din1(G173_p_spl_0011),
    .din2(g669_n_spl_00)
  );


  FA
  g_g838_n
  (
    .dout(g838_n),
    .din1(G173_n_spl_0011),
    .din2(g624_n_spl_00)
  );


  LA
  g_g839_p
  (
    .dout(g839_p),
    .din1(G172_p_spl_001),
    .din2(g838_n)
  );


  LA
  g_g840_p
  (
    .dout(g840_p),
    .din1(g837_n),
    .din2(g839_p)
  );


  FA
  g_g841_n
  (
    .dout(g841_n),
    .din1(g836_p),
    .din2(g840_p)
  );


  LA
  g_g842_p
  (
    .dout(g842_p),
    .din1(G25_p_spl_),
    .din2(G173_n_spl_010)
  );


  LA
  g_g843_p
  (
    .dout(g843_p),
    .din1(G24_p_spl_),
    .din2(G173_p_spl_010)
  );


  FA
  g_g844_n
  (
    .dout(g844_n),
    .din1(g842_p),
    .din2(g843_p)
  );


  LA
  g_g845_p
  (
    .dout(g845_p),
    .din1(G172_n_spl_01),
    .din2(g844_n)
  );


  FA
  g_g846_n
  (
    .dout(g846_n),
    .din1(G173_p_spl_010),
    .din2(g678_n_spl_00)
  );


  FA
  g_g847_n
  (
    .dout(g847_n),
    .din1(G173_n_spl_010),
    .din2(g569_p_spl_00)
  );


  LA
  g_g848_p
  (
    .dout(g848_p),
    .din1(G172_p_spl_01),
    .din2(g847_n)
  );


  LA
  g_g849_p
  (
    .dout(g849_p),
    .din1(g846_n),
    .din2(g848_p)
  );


  FA
  g_g850_n
  (
    .dout(g850_n),
    .din1(g845_p),
    .din2(g849_p)
  );


  LA
  g_g851_p
  (
    .dout(g851_p),
    .din1(G14_p_spl_),
    .din2(G174_n_spl_0001)
  );


  LA
  g_g852_p
  (
    .dout(g852_p),
    .din1(G16_p_spl_),
    .din2(G174_p_spl_0001)
  );


  FA
  g_g853_n
  (
    .dout(g853_n),
    .din1(g851_p),
    .din2(g852_p)
  );


  LA
  g_g854_p
  (
    .dout(g854_p),
    .din1(G175_n_spl_000),
    .din2(g853_n)
  );


  FA
  g_g855_n
  (
    .dout(g855_n),
    .din1(G174_p_spl_0001),
    .din2(g647_n_spl_00)
  );


  FA
  g_g856_n
  (
    .dout(g856_n),
    .din1(G174_n_spl_0001),
    .din2(g605_n_spl_00)
  );


  LA
  g_g857_p
  (
    .dout(g857_p),
    .din1(G175_p_spl_000),
    .din2(g856_n)
  );


  LA
  g_g858_p
  (
    .dout(g858_p),
    .din1(g855_n),
    .din2(g857_p)
  );


  FA
  g_g859_n
  (
    .dout(g859_n),
    .din1(g854_p),
    .din2(g858_p)
  );


  LA
  g_g860_p
  (
    .dout(g860_p),
    .din1(G6_p_spl_),
    .din2(G174_n_spl_0010)
  );


  LA
  g_g861_p
  (
    .dout(g861_p),
    .din1(G27_p_spl_),
    .din2(G174_p_spl_0010)
  );


  FA
  g_g862_n
  (
    .dout(g862_n),
    .din1(g860_p),
    .din2(g861_p)
  );


  LA
  g_g863_p
  (
    .dout(g863_p),
    .din1(G175_n_spl_001),
    .din2(g862_n)
  );


  FA
  g_g864_n
  (
    .dout(g864_n),
    .din1(G174_p_spl_0010),
    .din2(g656_n_spl_00)
  );


  FA
  g_g865_n
  (
    .dout(g865_n),
    .din1(G174_n_spl_0010),
    .din2(g614_n_spl_00)
  );


  LA
  g_g866_p
  (
    .dout(g866_p),
    .din1(G175_p_spl_001),
    .din2(g865_n)
  );


  LA
  g_g867_p
  (
    .dout(g867_p),
    .din1(g864_n),
    .din2(g866_p)
  );


  FA
  g_g868_n
  (
    .dout(g868_n),
    .din1(g863_p),
    .din2(g867_p)
  );


  LA
  g_g869_p
  (
    .dout(g869_p),
    .din1(G5_p_spl_),
    .din2(G174_n_spl_0011)
  );


  LA
  g_g870_p
  (
    .dout(g870_p),
    .din1(G26_p_spl_),
    .din2(G174_p_spl_0011)
  );


  FA
  g_g871_n
  (
    .dout(g871_n),
    .din1(g869_p),
    .din2(g870_p)
  );


  LA
  g_g872_p
  (
    .dout(g872_p),
    .din1(G175_n_spl_001),
    .din2(g871_n)
  );


  FA
  g_g873_n
  (
    .dout(g873_n),
    .din1(G174_p_spl_0011),
    .din2(g669_n_spl_00)
  );


  FA
  g_g874_n
  (
    .dout(g874_n),
    .din1(G174_n_spl_0011),
    .din2(g624_n_spl_00)
  );


  LA
  g_g875_p
  (
    .dout(g875_p),
    .din1(G175_p_spl_001),
    .din2(g874_n)
  );


  LA
  g_g876_p
  (
    .dout(g876_p),
    .din1(g873_n),
    .din2(g875_p)
  );


  FA
  g_g877_n
  (
    .dout(g877_n),
    .din1(g872_p),
    .din2(g876_p)
  );


  LA
  g_g878_p
  (
    .dout(g878_p),
    .din1(G25_p_spl_),
    .din2(G174_n_spl_010)
  );


  LA
  g_g879_p
  (
    .dout(g879_p),
    .din1(G24_p_spl_),
    .din2(G174_p_spl_010)
  );


  FA
  g_g880_n
  (
    .dout(g880_n),
    .din1(g878_p),
    .din2(g879_p)
  );


  LA
  g_g881_p
  (
    .dout(g881_p),
    .din1(G175_n_spl_01),
    .din2(g880_n)
  );


  FA
  g_g882_n
  (
    .dout(g882_n),
    .din1(G174_p_spl_010),
    .din2(g678_n_spl_00)
  );


  FA
  g_g883_n
  (
    .dout(g883_n),
    .din1(G174_n_spl_010),
    .din2(g569_p_spl_00)
  );


  LA
  g_g884_p
  (
    .dout(g884_p),
    .din1(G175_p_spl_01),
    .din2(g883_n)
  );


  LA
  g_g885_p
  (
    .dout(g885_p),
    .din1(g882_n),
    .din2(g884_p)
  );


  FA
  g_g886_n
  (
    .dout(g886_n),
    .din1(g881_p),
    .din2(g885_p)
  );


  LA
  g_g887_p
  (
    .dout(g887_p),
    .din1(G76_p_spl_),
    .din2(G158_n_spl_0001)
  );


  LA
  g_g888_p
  (
    .dout(g888_p),
    .din1(G86_p_spl_),
    .din2(G158_p_spl_0001)
  );


  FA
  g_g889_n
  (
    .dout(g889_n),
    .din1(g887_p),
    .din2(g888_p)
  );


  LA
  g_g890_p
  (
    .dout(g890_p),
    .din1(G159_n_spl_000),
    .din2(g889_n)
  );


  LA
  g_g891_p
  (
    .dout(g891_p),
    .din1(G158_p_spl_0001),
    .din2(g605_n_spl_0)
  );


  LA
  g_g892_p
  (
    .dout(g892_p),
    .din1(G158_n_spl_0001),
    .din2(g647_n_spl_0)
  );


  FA
  g_g893_n
  (
    .dout(g893_n),
    .din1(g891_p),
    .din2(g892_p)
  );


  LA
  g_g894_p
  (
    .dout(g894_p),
    .din1(G159_p_spl_000),
    .din2(g893_n)
  );


  FA
  g_g895_n
  (
    .dout(g895_n),
    .din1(g890_p),
    .din2(g894_p)
  );


  LA
  g_g896_p
  (
    .dout(g896_p),
    .din1(G64_p_spl_0001),
    .din2(g895_n)
  );


  LA
  g_g897_p
  (
    .dout(g897_p),
    .din1(G72_p_spl_),
    .din2(G158_n_spl_0010)
  );


  LA
  g_g898_p
  (
    .dout(g898_p),
    .din1(G82_p_spl_),
    .din2(G158_p_spl_0010)
  );


  FA
  g_g899_n
  (
    .dout(g899_n),
    .din1(g897_p),
    .din2(g898_p)
  );


  LA
  g_g900_p
  (
    .dout(g900_p),
    .din1(G159_n_spl_001),
    .din2(g899_n)
  );


  LA
  g_g901_p
  (
    .dout(g901_p),
    .din1(G158_p_spl_0010),
    .din2(g569_p_spl_0)
  );


  LA
  g_g902_p
  (
    .dout(g902_p),
    .din1(G158_n_spl_0010),
    .din2(g678_n_spl_0)
  );


  FA
  g_g903_n
  (
    .dout(g903_n),
    .din1(g901_p),
    .din2(g902_p)
  );


  LA
  g_g904_p
  (
    .dout(g904_p),
    .din1(G159_p_spl_001),
    .din2(g903_n)
  );


  FA
  g_g905_n
  (
    .dout(g905_n),
    .din1(g900_p),
    .din2(g904_p)
  );


  LA
  g_g906_p
  (
    .dout(g906_p),
    .din1(G64_p_spl_0001),
    .din2(g905_n)
  );


  LA
  g_g907_p
  (
    .dout(g907_p),
    .din1(G70_p_spl_),
    .din2(G158_n_spl_0011)
  );


  LA
  g_g908_p
  (
    .dout(g908_p),
    .din1(G71_p_spl_),
    .din2(G158_p_spl_0011)
  );


  FA
  g_g909_n
  (
    .dout(g909_n),
    .din1(g907_p),
    .din2(g908_p)
  );


  LA
  g_g910_p
  (
    .dout(g910_p),
    .din1(G159_n_spl_001),
    .din2(g909_n)
  );


  LA
  g_g911_p
  (
    .dout(g911_p),
    .din1(G158_p_spl_0011),
    .din2(g624_n_spl_0)
  );


  LA
  g_g912_p
  (
    .dout(g912_p),
    .din1(G158_n_spl_0011),
    .din2(g669_n_spl_0)
  );


  FA
  g_g913_n
  (
    .dout(g913_n),
    .din1(g911_p),
    .din2(g912_p)
  );


  LA
  g_g914_p
  (
    .dout(g914_p),
    .din1(G159_p_spl_001),
    .din2(g913_n)
  );


  FA
  g_g915_n
  (
    .dout(g915_n),
    .din1(g910_p),
    .din2(g914_p)
  );


  LA
  g_g916_p
  (
    .dout(g916_p),
    .din1(G64_p_spl_0010),
    .din2(g915_n)
  );


  LA
  g_g917_p
  (
    .dout(g917_p),
    .din1(G68_p_spl_),
    .din2(G158_n_spl_010)
  );


  LA
  g_g918_p
  (
    .dout(g918_p),
    .din1(G69_p_spl_),
    .din2(G158_p_spl_010)
  );


  FA
  g_g919_n
  (
    .dout(g919_n),
    .din1(g917_p),
    .din2(g918_p)
  );


  LA
  g_g920_p
  (
    .dout(g920_p),
    .din1(G159_n_spl_01),
    .din2(g919_n)
  );


  LA
  g_g921_p
  (
    .dout(g921_p),
    .din1(G158_p_spl_010),
    .din2(g614_n_spl_0)
  );


  LA
  g_g922_p
  (
    .dout(g922_p),
    .din1(G158_n_spl_010),
    .din2(g656_n_spl_0)
  );


  FA
  g_g923_n
  (
    .dout(g923_n),
    .din1(g921_p),
    .din2(g922_p)
  );


  LA
  g_g924_p
  (
    .dout(g924_p),
    .din1(G159_p_spl_01),
    .din2(g923_n)
  );


  FA
  g_g925_n
  (
    .dout(g925_n),
    .din1(g920_p),
    .din2(g924_p)
  );


  LA
  g_g926_p
  (
    .dout(g926_p),
    .din1(G64_p_spl_0010),
    .din2(g925_n)
  );


  LA
  g_g927_p
  (
    .dout(g927_p),
    .din1(G76_p_spl_),
    .din2(G160_n_spl_0001)
  );


  LA
  g_g928_p
  (
    .dout(g928_p),
    .din1(G86_p_spl_),
    .din2(G160_p_spl_0001)
  );


  FA
  g_g929_n
  (
    .dout(g929_n),
    .din1(g927_p),
    .din2(g928_p)
  );


  LA
  g_g930_p
  (
    .dout(g930_p),
    .din1(G161_n_spl_000),
    .din2(g929_n)
  );


  LA
  g_g931_p
  (
    .dout(g931_p),
    .din1(G160_p_spl_0001),
    .din2(g605_n_spl_1)
  );


  LA
  g_g932_p
  (
    .dout(g932_p),
    .din1(G160_n_spl_0001),
    .din2(g647_n_spl_1)
  );


  FA
  g_g933_n
  (
    .dout(g933_n),
    .din1(g931_p),
    .din2(g932_p)
  );


  LA
  g_g934_p
  (
    .dout(g934_p),
    .din1(G161_p_spl_000),
    .din2(g933_n)
  );


  FA
  g_g935_n
  (
    .dout(g935_n),
    .din1(g930_p),
    .din2(g934_p)
  );


  LA
  g_g936_p
  (
    .dout(g936_p),
    .din1(G64_p_spl_001),
    .din2(g935_n)
  );


  LA
  g_g937_p
  (
    .dout(g937_p),
    .din1(G72_p_spl_),
    .din2(G160_n_spl_0010)
  );


  LA
  g_g938_p
  (
    .dout(g938_p),
    .din1(G82_p_spl_),
    .din2(G160_p_spl_0010)
  );


  FA
  g_g939_n
  (
    .dout(g939_n),
    .din1(g937_p),
    .din2(g938_p)
  );


  LA
  g_g940_p
  (
    .dout(g940_p),
    .din1(G161_n_spl_001),
    .din2(g939_n)
  );


  LA
  g_g941_p
  (
    .dout(g941_p),
    .din1(G160_p_spl_0010),
    .din2(g569_p_spl_1)
  );


  LA
  g_g942_p
  (
    .dout(g942_p),
    .din1(G160_n_spl_0010),
    .din2(g678_n_spl_1)
  );


  FA
  g_g943_n
  (
    .dout(g943_n),
    .din1(g941_p),
    .din2(g942_p)
  );


  LA
  g_g944_p
  (
    .dout(g944_p),
    .din1(G161_p_spl_001),
    .din2(g943_n)
  );


  FA
  g_g945_n
  (
    .dout(g945_n),
    .din1(g940_p),
    .din2(g944_p)
  );


  LA
  g_g946_p
  (
    .dout(g946_p),
    .din1(G64_p_spl_010),
    .din2(g945_n)
  );


  LA
  g_g947_p
  (
    .dout(g947_p),
    .din1(G70_p_spl_),
    .din2(G160_n_spl_0011)
  );


  LA
  g_g948_p
  (
    .dout(g948_p),
    .din1(G71_p_spl_),
    .din2(G160_p_spl_0011)
  );


  FA
  g_g949_n
  (
    .dout(g949_n),
    .din1(g947_p),
    .din2(g948_p)
  );


  LA
  g_g950_p
  (
    .dout(g950_p),
    .din1(G161_n_spl_001),
    .din2(g949_n)
  );


  LA
  g_g951_p
  (
    .dout(g951_p),
    .din1(G160_p_spl_0011),
    .din2(g624_n_spl_1)
  );


  LA
  g_g952_p
  (
    .dout(g952_p),
    .din1(G160_n_spl_0011),
    .din2(g669_n_spl_1)
  );


  FA
  g_g953_n
  (
    .dout(g953_n),
    .din1(g951_p),
    .din2(g952_p)
  );


  LA
  g_g954_p
  (
    .dout(g954_p),
    .din1(G161_p_spl_001),
    .din2(g953_n)
  );


  FA
  g_g955_n
  (
    .dout(g955_n),
    .din1(g950_p),
    .din2(g954_p)
  );


  LA
  g_g956_p
  (
    .dout(g956_p),
    .din1(G64_p_spl_010),
    .din2(g955_n)
  );


  LA
  g_g957_p
  (
    .dout(g957_p),
    .din1(G68_p_spl_),
    .din2(G160_n_spl_010)
  );


  LA
  g_g958_p
  (
    .dout(g958_p),
    .din1(G69_p_spl_),
    .din2(G160_p_spl_010)
  );


  FA
  g_g959_n
  (
    .dout(g959_n),
    .din1(g957_p),
    .din2(g958_p)
  );


  LA
  g_g960_p
  (
    .dout(g960_p),
    .din1(G161_n_spl_01),
    .din2(g959_n)
  );


  LA
  g_g961_p
  (
    .dout(g961_p),
    .din1(G160_p_spl_010),
    .din2(g614_n_spl_1)
  );


  LA
  g_g962_p
  (
    .dout(g962_p),
    .din1(G160_n_spl_010),
    .din2(g656_n_spl_1)
  );


  FA
  g_g963_n
  (
    .dout(g963_n),
    .din1(g961_p),
    .din2(g962_p)
  );


  LA
  g_g964_p
  (
    .dout(g964_p),
    .din1(G161_p_spl_01),
    .din2(g963_n)
  );


  FA
  g_g965_n
  (
    .dout(g965_n),
    .din1(g960_p),
    .din2(g964_p)
  );


  LA
  g_g966_p
  (
    .dout(g966_p),
    .din1(G64_p_spl_011),
    .din2(g965_n)
  );


  FA
  g_g967_n
  (
    .dout(g967_n),
    .din1(G62_n),
    .din2(G178_n)
  );


  LA
  g_g968_p
  (
    .dout(g968_p),
    .din1(G171_p_spl_),
    .din2(g581_n_spl_01)
  );


  LA
  g_g969_p
  (
    .dout(g969_p),
    .din1(G54_p_spl_),
    .din2(G171_n_spl_)
  );


  FA
  g_g970_n
  (
    .dout(g970_n),
    .din1(g968_p),
    .din2(g969_p)
  );


  LA
  g_g971_p
  (
    .dout(g971_p),
    .din1(G170_p),
    .din2(g970_n)
  );


  LA
  g_g972_p
  (
    .dout(g972_p),
    .din1(G171_n_spl_),
    .din2(g237_n_spl_0)
  );


  LA
  g_g973_p
  (
    .dout(g973_p),
    .din1(G61_n_spl_),
    .din2(g476_n_spl_1)
  );


  FA
  g_g973_n
  (
    .dout(g973_n),
    .din1(G61_p_spl_),
    .din2(g476_p_spl_1)
  );


  LA
  g_g974_p
  (
    .dout(g974_p),
    .din1(G61_p_spl_),
    .din2(g476_p_spl_1)
  );


  FA
  g_g974_n
  (
    .dout(g974_n),
    .din1(G61_n_spl_),
    .din2(g476_n_spl_1)
  );


  LA
  g_g975_p
  (
    .dout(g975_p),
    .din1(g973_n),
    .din2(g974_n)
  );


  FA
  g_g975_n
  (
    .dout(g975_n),
    .din1(g973_p),
    .din2(g974_p)
  );


  LA
  g_g976_p
  (
    .dout(g976_p),
    .din1(G171_p_spl_),
    .din2(g975_p_spl_)
  );


  FA
  g_g977_n
  (
    .dout(g977_n),
    .din1(g972_p),
    .din2(g976_p)
  );


  LA
  g_g978_p
  (
    .dout(g978_p),
    .din1(G170_n),
    .din2(g977_n)
  );


  FA
  g_g979_n
  (
    .dout(g979_n),
    .din1(g971_p),
    .din2(g978_p)
  );


  LA
  g_g980_p
  (
    .dout(g980_p),
    .din1(g967_n),
    .din2(g979_n)
  );


  LA
  g_g981_p
  (
    .dout(g981_p),
    .din1(g581_n_spl_10),
    .din2(g975_n)
  );


  LA
  g_g982_p
  (
    .dout(g982_p),
    .din1(g581_p_spl_01),
    .din2(g975_p_spl_)
  );


  FA
  g_g983_n
  (
    .dout(g983_n),
    .din1(g981_p),
    .din2(g982_p)
  );


  LA
  g_g984_p
  (
    .dout(g984_p),
    .din1(G177_p_spl_0110),
    .din2(g581_n_spl_10)
  );


  FA
  g_g985_n
  (
    .dout(g985_n),
    .din1(G176_p_spl_0111),
    .din2(g984_p)
  );


  FA
  g_g986_n
  (
    .dout(g986_n),
    .din1(G177_n_spl_011),
    .din2(g237_n_spl_1)
  );


  FA
  g_g987_n
  (
    .dout(g987_n),
    .din1(G176_n_spl_0101),
    .din2(g986_n)
  );


  FA
  g_g988_n
  (
    .dout(g988_n),
    .din1(G54_p_spl_),
    .din2(G177_p_spl_0111)
  );


  LA
  g_g989_p
  (
    .dout(g989_p),
    .din1(g987_n),
    .din2(g988_n)
  );


  LA
  g_g990_p
  (
    .dout(g990_p),
    .din1(g985_n),
    .din2(g989_p)
  );


  LA
  g_g991_p
  (
    .dout(g991_p),
    .din1(G52_p),
    .din2(G177_n_spl_011)
  );


  LA
  g_g992_p
  (
    .dout(g992_p),
    .din1(G176_p_spl_1000),
    .din2(g991_p)
  );


  FA
  g_g993_n
  (
    .dout(g993_n),
    .din1(G176_p_spl_1000),
    .din2(g785_p_spl_)
  );


  FA
  g_g994_n
  (
    .dout(g994_n),
    .din1(G176_n_spl_0101),
    .din2(g240_n_spl_0)
  );


  LA
  g_g995_p
  (
    .dout(g995_p),
    .din1(G177_p_spl_0111),
    .din2(g994_n)
  );


  LA
  g_g996_p
  (
    .dout(g996_p),
    .din1(g993_n),
    .din2(g995_p)
  );


  FA
  g_g997_n
  (
    .dout(g997_n),
    .din1(g992_p),
    .din2(g996_p)
  );


  LA
  g_g998_p
  (
    .dout(g998_p),
    .din1(G47_p),
    .din2(G177_n_spl_100)
  );


  LA
  g_g999_p
  (
    .dout(g999_p),
    .din1(G176_p_spl_1001),
    .din2(g998_p)
  );


  FA
  g_g1000_n
  (
    .dout(g1000_n),
    .din1(G176_p_spl_1001),
    .din2(g791_p_spl_)
  );


  FA
  g_g1001_n
  (
    .dout(g1001_n),
    .din1(G176_n_spl_011),
    .din2(g267_n_spl_0)
  );


  LA
  g_g1002_p
  (
    .dout(g1002_p),
    .din1(G177_p_spl_1000),
    .din2(g1001_n)
  );


  LA
  g_g1003_p
  (
    .dout(g1003_p),
    .din1(g1000_n),
    .din2(g1002_p)
  );


  FA
  g_g1004_n
  (
    .dout(g1004_n),
    .din1(g999_p),
    .din2(g1003_p)
  );


  LA
  g_g1005_p
  (
    .dout(g1005_p),
    .din1(G43_p),
    .din2(G177_n_spl_100)
  );


  LA
  g_g1006_p
  (
    .dout(g1006_p),
    .din1(G176_p_spl_1010),
    .din2(g1005_p)
  );


  FA
  g_g1007_n
  (
    .dout(g1007_n),
    .din1(G176_n_spl_011),
    .din2(g258_n_spl_0)
  );


  FA
  g_g1008_n
  (
    .dout(g1008_n),
    .din1(G176_p_spl_1010),
    .din2(g777_p_spl_)
  );


  LA
  g_g1009_p
  (
    .dout(g1009_p),
    .din1(G177_p_spl_1000),
    .din2(g1008_n)
  );


  LA
  g_g1010_p
  (
    .dout(g1010_p),
    .din1(g1007_n),
    .din2(g1009_p)
  );


  FA
  g_g1011_n
  (
    .dout(g1011_n),
    .din1(g1006_p),
    .din2(g1010_p)
  );


  FA
  g_g1012_n
  (
    .dout(g1012_n),
    .din1(G99_n_spl_),
    .din2(g533_n_spl_)
  );


  FA
  g_g1013_n
  (
    .dout(g1013_n),
    .din1(g735_n_spl_),
    .din2(g1012_n)
  );


  FA
  g_g1014_n
  (
    .dout(g1014_n),
    .din1(G155_n_spl_),
    .din2(g184_n_spl_)
  );


  FA
  g_g1015_n
  (
    .dout(g1015_n),
    .din1(g179_n_spl_),
    .din2(g1014_n)
  );


  FA
  g_g1016_n
  (
    .dout(g1016_n),
    .din1(g705_n_spl_),
    .din2(g1015_n)
  );


  FA
  g_g1017_n
  (
    .dout(g1017_n),
    .din1(g506_n_spl_),
    .din2(g1016_n)
  );


  FA
  g_g1018_n
  (
    .dout(g1018_n),
    .din1(g1013_n),
    .din2(g1017_n)
  );


  LA
  g_g1019_p
  (
    .dout(g1019_p),
    .din1(G46_p),
    .din2(G177_n_spl_101)
  );


  LA
  g_g1020_p
  (
    .dout(g1020_p),
    .din1(G176_p_spl_1011),
    .din2(g1019_p)
  );


  FA
  g_g1021_n
  (
    .dout(g1021_n),
    .din1(G176_p_spl_1011),
    .din2(g760_p_spl_)
  );


  FA
  g_g1022_n
  (
    .dout(g1022_n),
    .din1(G176_n_spl_100),
    .din2(g317_n_spl_0)
  );


  LA
  g_g1023_p
  (
    .dout(g1023_p),
    .din1(G177_p_spl_1001),
    .din2(g1022_n)
  );


  LA
  g_g1024_p
  (
    .dout(g1024_p),
    .din1(g1021_n),
    .din2(g1023_p)
  );


  FA
  g_g1025_n
  (
    .dout(g1025_n),
    .din1(g1020_p),
    .din2(g1024_p)
  );


  LA
  g_g1026_p
  (
    .dout(g1026_p),
    .din1(G45_p),
    .din2(G177_n_spl_101)
  );


  LA
  g_g1027_p
  (
    .dout(g1027_p),
    .din1(G176_p_spl_1100),
    .din2(g1026_p)
  );


  FA
  g_g1028_n
  (
    .dout(g1028_n),
    .din1(G176_p_spl_1100),
    .din2(g755_p_spl_)
  );


  FA
  g_g1029_n
  (
    .dout(g1029_n),
    .din1(G176_n_spl_100),
    .din2(g328_n_spl_)
  );


  LA
  g_g1030_p
  (
    .dout(g1030_p),
    .din1(G177_p_spl_1001),
    .din2(g1029_n)
  );


  LA
  g_g1031_p
  (
    .dout(g1031_p),
    .din1(g1028_n),
    .din2(g1030_p)
  );


  FA
  g_g1032_n
  (
    .dout(g1032_n),
    .din1(g1027_p),
    .din2(g1031_p)
  );


  LA
  g_g1033_p
  (
    .dout(g1033_p),
    .din1(G20_p),
    .din2(G177_n_spl_110)
  );


  LA
  g_g1034_p
  (
    .dout(g1034_p),
    .din1(G176_p_spl_1101),
    .din2(g1033_p)
  );


  FA
  g_g1035_n
  (
    .dout(g1035_n),
    .din1(G176_p_spl_1101),
    .din2(g743_p_spl_)
  );


  FA
  g_g1036_n
  (
    .dout(g1036_n),
    .din1(G176_n_spl_101),
    .din2(g337_n_spl_)
  );


  LA
  g_g1037_p
  (
    .dout(g1037_p),
    .din1(G177_p_spl_101),
    .din2(g1036_n)
  );


  LA
  g_g1038_p
  (
    .dout(g1038_p),
    .din1(g1035_n),
    .din2(g1037_p)
  );


  FA
  g_g1039_n
  (
    .dout(g1039_n),
    .din1(g1034_p),
    .din2(g1038_p)
  );


  LA
  g_g1040_p
  (
    .dout(g1040_p),
    .din1(G44_p),
    .din2(G177_n_spl_110)
  );


  LA
  g_g1041_p
  (
    .dout(g1041_p),
    .din1(G176_p_spl_1110),
    .din2(g1040_p)
  );


  FA
  g_g1042_n
  (
    .dout(g1042_n),
    .din1(G176_p_spl_1110),
    .din2(g747_p_spl_)
  );


  FA
  g_g1043_n
  (
    .dout(g1043_n),
    .din1(G176_n_spl_101),
    .din2(g347_n_spl_)
  );


  LA
  g_g1044_p
  (
    .dout(g1044_p),
    .din1(G177_p_spl_101),
    .din2(g1043_n)
  );


  LA
  g_g1045_p
  (
    .dout(g1045_p),
    .din1(g1042_n),
    .din2(g1044_p)
  );


  FA
  g_g1046_n
  (
    .dout(g1046_n),
    .din1(g1041_p),
    .din2(g1045_p)
  );


  FA
  g_g1047_n
  (
    .dout(g1047_n),
    .din1(G174_p_spl_011),
    .din2(g1025_n_spl_00)
  );


  FA
  g_g1048_n
  (
    .dout(g1048_n),
    .din1(G174_n_spl_011),
    .din2(g990_p_spl_00)
  );


  LA
  g_g1049_p
  (
    .dout(g1049_p),
    .din1(G175_p_spl_01),
    .din2(g1048_n)
  );


  LA
  g_g1050_p
  (
    .dout(g1050_p),
    .din1(g1047_n),
    .din2(g1049_p)
  );


  LA
  g_g1051_p
  (
    .dout(g1051_p),
    .din1(G41_p_spl_),
    .din2(G174_n_spl_011)
  );


  LA
  g_g1052_p
  (
    .dout(g1052_p),
    .din1(G42_p_spl_),
    .din2(G174_p_spl_011)
  );


  FA
  g_g1053_n
  (
    .dout(g1053_n),
    .din1(g1051_p),
    .din2(g1052_p)
  );


  LA
  g_g1054_p
  (
    .dout(g1054_p),
    .din1(G175_n_spl_01),
    .din2(g1053_n)
  );


  FA
  g_g1055_n
  (
    .dout(g1055_n),
    .din1(g1050_p),
    .din2(g1054_p)
  );


  FA
  g_g1056_n
  (
    .dout(g1056_n),
    .din1(G173_p_spl_011),
    .din2(g1025_n_spl_00)
  );


  FA
  g_g1057_n
  (
    .dout(g1057_n),
    .din1(G173_n_spl_011),
    .din2(g990_p_spl_00)
  );


  LA
  g_g1058_p
  (
    .dout(g1058_p),
    .din1(G172_p_spl_01),
    .din2(g1057_n)
  );


  LA
  g_g1059_p
  (
    .dout(g1059_p),
    .din1(g1056_n),
    .din2(g1058_p)
  );


  LA
  g_g1060_p
  (
    .dout(g1060_p),
    .din1(G41_p_spl_),
    .din2(G173_n_spl_011)
  );


  LA
  g_g1061_p
  (
    .dout(g1061_p),
    .din1(G42_p_spl_),
    .din2(G173_p_spl_011)
  );


  FA
  g_g1062_n
  (
    .dout(g1062_n),
    .din1(g1060_p),
    .din2(g1061_p)
  );


  LA
  g_g1063_p
  (
    .dout(g1063_p),
    .din1(G172_n_spl_01),
    .din2(g1062_n)
  );


  FA
  g_g1064_n
  (
    .dout(g1064_n),
    .din1(g1059_p),
    .din2(g1063_p)
  );


  LA
  g_g1065_p
  (
    .dout(g1065_p),
    .din1(G18_p_spl_),
    .din2(G173_n_spl_100)
  );


  LA
  g_g1066_p
  (
    .dout(g1066_p),
    .din1(G17_p_spl_),
    .din2(G173_p_spl_100)
  );


  FA
  g_g1067_n
  (
    .dout(g1067_n),
    .din1(g1065_p),
    .din2(g1066_p)
  );


  LA
  g_g1068_p
  (
    .dout(g1068_p),
    .din1(G172_n_spl_10),
    .din2(g1067_n)
  );


  FA
  g_g1069_n
  (
    .dout(g1069_n),
    .din1(G173_p_spl_100),
    .din2(g1032_n_spl_00)
  );


  FA
  g_g1070_n
  (
    .dout(g1070_n),
    .din1(G173_n_spl_100),
    .din2(g997_n_spl_00)
  );


  LA
  g_g1071_p
  (
    .dout(g1071_p),
    .din1(G172_p_spl_10),
    .din2(g1070_n)
  );


  LA
  g_g1072_p
  (
    .dout(g1072_p),
    .din1(g1069_n),
    .din2(g1071_p)
  );


  FA
  g_g1073_n
  (
    .dout(g1073_n),
    .din1(g1068_p),
    .din2(g1072_p)
  );


  LA
  g_g1074_p
  (
    .dout(g1074_p),
    .din1(G40_p_spl_),
    .din2(G173_n_spl_101)
  );


  LA
  g_g1075_p
  (
    .dout(g1075_p),
    .din1(G39_p_spl_),
    .din2(G173_p_spl_101)
  );


  FA
  g_g1076_n
  (
    .dout(g1076_n),
    .din1(g1074_p),
    .din2(g1075_p)
  );


  LA
  g_g1077_p
  (
    .dout(g1077_p),
    .din1(G172_n_spl_10),
    .din2(g1076_n)
  );


  FA
  g_g1078_n
  (
    .dout(g1078_n),
    .din1(G173_p_spl_101),
    .din2(g1039_n_spl_00)
  );


  FA
  g_g1079_n
  (
    .dout(g1079_n),
    .din1(G173_n_spl_101),
    .din2(g1004_n_spl_00)
  );


  LA
  g_g1080_p
  (
    .dout(g1080_p),
    .din1(G172_p_spl_10),
    .din2(g1079_n)
  );


  LA
  g_g1081_p
  (
    .dout(g1081_p),
    .din1(g1078_n),
    .din2(g1080_p)
  );


  FA
  g_g1082_n
  (
    .dout(g1082_n),
    .din1(g1077_p),
    .din2(g1081_p)
  );


  LA
  g_g1083_p
  (
    .dout(g1083_p),
    .din1(G15_p_spl_),
    .din2(G173_n_spl_110)
  );


  LA
  g_g1084_p
  (
    .dout(g1084_p),
    .din1(G36_p_spl_),
    .din2(G173_p_spl_110)
  );


  FA
  g_g1085_n
  (
    .dout(g1085_n),
    .din1(g1083_p),
    .din2(g1084_p)
  );


  LA
  g_g1086_p
  (
    .dout(g1086_p),
    .din1(G172_n_spl_11),
    .din2(g1085_n)
  );


  FA
  g_g1087_n
  (
    .dout(g1087_n),
    .din1(G173_p_spl_110),
    .din2(g1046_n_spl_00)
  );


  FA
  g_g1088_n
  (
    .dout(g1088_n),
    .din1(G173_n_spl_110),
    .din2(g1011_n_spl_00)
  );


  LA
  g_g1089_p
  (
    .dout(g1089_p),
    .din1(G172_p_spl_11),
    .din2(g1088_n)
  );


  LA
  g_g1090_p
  (
    .dout(g1090_p),
    .din1(g1087_n),
    .din2(g1089_p)
  );


  FA
  g_g1091_n
  (
    .dout(g1091_n),
    .din1(g1086_p),
    .din2(g1090_p)
  );


  LA
  g_g1092_p
  (
    .dout(g1092_p),
    .din1(G18_p_spl_),
    .din2(G174_n_spl_100)
  );


  LA
  g_g1093_p
  (
    .dout(g1093_p),
    .din1(G17_p_spl_),
    .din2(G174_p_spl_100)
  );


  FA
  g_g1094_n
  (
    .dout(g1094_n),
    .din1(g1092_p),
    .din2(g1093_p)
  );


  LA
  g_g1095_p
  (
    .dout(g1095_p),
    .din1(G175_n_spl_10),
    .din2(g1094_n)
  );


  FA
  g_g1096_n
  (
    .dout(g1096_n),
    .din1(G174_p_spl_100),
    .din2(g1032_n_spl_00)
  );


  FA
  g_g1097_n
  (
    .dout(g1097_n),
    .din1(G174_n_spl_100),
    .din2(g997_n_spl_00)
  );


  LA
  g_g1098_p
  (
    .dout(g1098_p),
    .din1(G175_p_spl_10),
    .din2(g1097_n)
  );


  LA
  g_g1099_p
  (
    .dout(g1099_p),
    .din1(g1096_n),
    .din2(g1098_p)
  );


  FA
  g_g1100_n
  (
    .dout(g1100_n),
    .din1(g1095_p),
    .din2(g1099_p)
  );


  LA
  g_g1101_p
  (
    .dout(g1101_p),
    .din1(G40_p_spl_),
    .din2(G174_n_spl_101)
  );


  LA
  g_g1102_p
  (
    .dout(g1102_p),
    .din1(G39_p_spl_),
    .din2(G174_p_spl_101)
  );


  FA
  g_g1103_n
  (
    .dout(g1103_n),
    .din1(g1101_p),
    .din2(g1102_p)
  );


  LA
  g_g1104_p
  (
    .dout(g1104_p),
    .din1(G175_n_spl_10),
    .din2(g1103_n)
  );


  FA
  g_g1105_n
  (
    .dout(g1105_n),
    .din1(G174_p_spl_101),
    .din2(g1039_n_spl_00)
  );


  FA
  g_g1106_n
  (
    .dout(g1106_n),
    .din1(G174_n_spl_101),
    .din2(g1004_n_spl_00)
  );


  LA
  g_g1107_p
  (
    .dout(g1107_p),
    .din1(G175_p_spl_10),
    .din2(g1106_n)
  );


  LA
  g_g1108_p
  (
    .dout(g1108_p),
    .din1(g1105_n),
    .din2(g1107_p)
  );


  FA
  g_g1109_n
  (
    .dout(g1109_n),
    .din1(g1104_p),
    .din2(g1108_p)
  );


  LA
  g_g1110_p
  (
    .dout(g1110_p),
    .din1(G15_p_spl_),
    .din2(G174_n_spl_110)
  );


  LA
  g_g1111_p
  (
    .dout(g1111_p),
    .din1(G36_p_spl_),
    .din2(G174_p_spl_110)
  );


  FA
  g_g1112_n
  (
    .dout(g1112_n),
    .din1(g1110_p),
    .din2(g1111_p)
  );


  LA
  g_g1113_p
  (
    .dout(g1113_p),
    .din1(G175_n_spl_11),
    .din2(g1112_n)
  );


  FA
  g_g1114_n
  (
    .dout(g1114_n),
    .din1(G174_p_spl_110),
    .din2(g1046_n_spl_00)
  );


  FA
  g_g1115_n
  (
    .dout(g1115_n),
    .din1(G174_n_spl_110),
    .din2(g1011_n_spl_00)
  );


  LA
  g_g1116_p
  (
    .dout(g1116_p),
    .din1(G175_p_spl_11),
    .din2(g1115_n)
  );


  LA
  g_g1117_p
  (
    .dout(g1117_p),
    .din1(g1114_n),
    .din2(g1116_p)
  );


  FA
  g_g1118_n
  (
    .dout(g1118_n),
    .din1(g1113_p),
    .din2(g1117_p)
  );


  LA
  g_g1119_p
  (
    .dout(g1119_p),
    .din1(G77_p_spl_),
    .din2(G158_n_spl_011)
  );


  LA
  g_g1120_p
  (
    .dout(g1120_p),
    .din1(G87_p_spl_),
    .din2(G158_p_spl_011)
  );


  FA
  g_g1121_n
  (
    .dout(g1121_n),
    .din1(g1119_p),
    .din2(g1120_p)
  );


  LA
  g_g1122_p
  (
    .dout(g1122_p),
    .din1(G159_n_spl_01),
    .din2(g1121_n)
  );


  LA
  g_g1123_p
  (
    .dout(g1123_p),
    .din1(G158_p_spl_011),
    .din2(g1011_n_spl_0)
  );


  LA
  g_g1124_p
  (
    .dout(g1124_p),
    .din1(G158_n_spl_011),
    .din2(g1046_n_spl_0)
  );


  FA
  g_g1125_n
  (
    .dout(g1125_n),
    .din1(g1123_p),
    .din2(g1124_p)
  );


  LA
  g_g1126_p
  (
    .dout(g1126_p),
    .din1(G159_p_spl_01),
    .din2(g1125_n)
  );


  FA
  g_g1127_n
  (
    .dout(g1127_n),
    .din1(g1122_p),
    .din2(g1126_p)
  );


  LA
  g_g1128_p
  (
    .dout(g1128_p),
    .din1(G64_p_spl_011),
    .din2(g1127_n)
  );


  LA
  g_g1129_p
  (
    .dout(g1129_p),
    .din1(G75_p_spl_),
    .din2(G158_n_spl_100)
  );


  LA
  g_g1130_p
  (
    .dout(g1130_p),
    .din1(G85_p_spl_),
    .din2(G158_p_spl_100)
  );


  FA
  g_g1131_n
  (
    .dout(g1131_n),
    .din1(g1129_p),
    .din2(g1130_p)
  );


  LA
  g_g1132_p
  (
    .dout(g1132_p),
    .din1(G159_n_spl_10),
    .din2(g1131_n)
  );


  LA
  g_g1133_p
  (
    .dout(g1133_p),
    .din1(G158_p_spl_100),
    .din2(g1004_n_spl_0)
  );


  LA
  g_g1134_p
  (
    .dout(g1134_p),
    .din1(G158_n_spl_100),
    .din2(g1039_n_spl_0)
  );


  FA
  g_g1135_n
  (
    .dout(g1135_n),
    .din1(g1133_p),
    .din2(g1134_p)
  );


  LA
  g_g1136_p
  (
    .dout(g1136_p),
    .din1(G159_p_spl_10),
    .din2(g1135_n)
  );


  FA
  g_g1137_n
  (
    .dout(g1137_n),
    .din1(g1132_p),
    .din2(g1136_p)
  );


  LA
  g_g1138_p
  (
    .dout(g1138_p),
    .din1(G64_p_spl_100),
    .din2(g1137_n)
  );


  LA
  g_g1139_p
  (
    .dout(g1139_p),
    .din1(G74_p_spl_),
    .din2(G158_n_spl_101)
  );


  LA
  g_g1140_p
  (
    .dout(g1140_p),
    .din1(G84_p_spl_),
    .din2(G158_p_spl_101)
  );


  FA
  g_g1141_n
  (
    .dout(g1141_n),
    .din1(g1139_p),
    .din2(g1140_p)
  );


  LA
  g_g1142_p
  (
    .dout(g1142_p),
    .din1(G159_n_spl_10),
    .din2(g1141_n)
  );


  LA
  g_g1143_p
  (
    .dout(g1143_p),
    .din1(G158_p_spl_101),
    .din2(g997_n_spl_0)
  );


  LA
  g_g1144_p
  (
    .dout(g1144_p),
    .din1(G158_n_spl_101),
    .din2(g1032_n_spl_0)
  );


  FA
  g_g1145_n
  (
    .dout(g1145_n),
    .din1(g1143_p),
    .din2(g1144_p)
  );


  LA
  g_g1146_p
  (
    .dout(g1146_p),
    .din1(G159_p_spl_10),
    .din2(g1145_n)
  );


  FA
  g_g1147_n
  (
    .dout(g1147_n),
    .din1(g1142_p),
    .din2(g1146_p)
  );


  LA
  g_g1148_p
  (
    .dout(g1148_p),
    .din1(G64_p_spl_100),
    .din2(g1147_n)
  );


  FA
  g_g1149_n
  (
    .dout(g1149_n),
    .din1(G158_p_spl_110),
    .din2(g1025_n_spl_0)
  );


  FA
  g_g1150_n
  (
    .dout(g1150_n),
    .din1(G158_n_spl_110),
    .din2(g990_p_spl_0)
  );


  LA
  g_g1151_p
  (
    .dout(g1151_p),
    .din1(G159_p_spl_11),
    .din2(g1150_n)
  );


  LA
  g_g1152_p
  (
    .dout(g1152_p),
    .din1(g1149_n),
    .din2(g1151_p)
  );


  LA
  g_g1153_p
  (
    .dout(g1153_p),
    .din1(G73_p_spl_),
    .din2(G158_n_spl_110)
  );


  LA
  g_g1154_p
  (
    .dout(g1154_p),
    .din1(G83_p_spl_),
    .din2(G158_p_spl_110)
  );


  FA
  g_g1155_n
  (
    .dout(g1155_n),
    .din1(g1153_p),
    .din2(g1154_p)
  );


  LA
  g_g1156_p
  (
    .dout(g1156_p),
    .din1(G159_n_spl_11),
    .din2(g1155_n)
  );


  FA
  g_g1157_n
  (
    .dout(g1157_n),
    .din1(g1152_p),
    .din2(g1156_p)
  );


  LA
  g_g1158_p
  (
    .dout(g1158_p),
    .din1(G64_p_spl_101),
    .din2(g1157_n)
  );


  LA
  g_g1159_p
  (
    .dout(g1159_p),
    .din1(G77_p_spl_),
    .din2(G160_n_spl_011)
  );


  LA
  g_g1160_p
  (
    .dout(g1160_p),
    .din1(G87_p_spl_),
    .din2(G160_p_spl_011)
  );


  FA
  g_g1161_n
  (
    .dout(g1161_n),
    .din1(g1159_p),
    .din2(g1160_p)
  );


  LA
  g_g1162_p
  (
    .dout(g1162_p),
    .din1(G161_n_spl_01),
    .din2(g1161_n)
  );


  LA
  g_g1163_p
  (
    .dout(g1163_p),
    .din1(G160_p_spl_011),
    .din2(g1011_n_spl_1)
  );


  LA
  g_g1164_p
  (
    .dout(g1164_p),
    .din1(G160_n_spl_011),
    .din2(g1046_n_spl_1)
  );


  FA
  g_g1165_n
  (
    .dout(g1165_n),
    .din1(g1163_p),
    .din2(g1164_p)
  );


  LA
  g_g1166_p
  (
    .dout(g1166_p),
    .din1(G161_p_spl_01),
    .din2(g1165_n)
  );


  FA
  g_g1167_n
  (
    .dout(g1167_n),
    .din1(g1162_p),
    .din2(g1166_p)
  );


  LA
  g_g1168_p
  (
    .dout(g1168_p),
    .din1(G64_p_spl_101),
    .din2(g1167_n)
  );


  LA
  g_g1169_p
  (
    .dout(g1169_p),
    .din1(G75_p_spl_),
    .din2(G160_n_spl_100)
  );


  LA
  g_g1170_p
  (
    .dout(g1170_p),
    .din1(G85_p_spl_),
    .din2(G160_p_spl_100)
  );


  FA
  g_g1171_n
  (
    .dout(g1171_n),
    .din1(g1169_p),
    .din2(g1170_p)
  );


  LA
  g_g1172_p
  (
    .dout(g1172_p),
    .din1(G161_n_spl_10),
    .din2(g1171_n)
  );


  LA
  g_g1173_p
  (
    .dout(g1173_p),
    .din1(G160_p_spl_100),
    .din2(g1004_n_spl_1)
  );


  LA
  g_g1174_p
  (
    .dout(g1174_p),
    .din1(G160_n_spl_100),
    .din2(g1039_n_spl_1)
  );


  FA
  g_g1175_n
  (
    .dout(g1175_n),
    .din1(g1173_p),
    .din2(g1174_p)
  );


  LA
  g_g1176_p
  (
    .dout(g1176_p),
    .din1(G161_p_spl_10),
    .din2(g1175_n)
  );


  FA
  g_g1177_n
  (
    .dout(g1177_n),
    .din1(g1172_p),
    .din2(g1176_p)
  );


  LA
  g_g1178_p
  (
    .dout(g1178_p),
    .din1(G64_p_spl_110),
    .din2(g1177_n)
  );


  LA
  g_g1179_p
  (
    .dout(g1179_p),
    .din1(G74_p_spl_),
    .din2(G160_n_spl_101)
  );


  LA
  g_g1180_p
  (
    .dout(g1180_p),
    .din1(G84_p_spl_),
    .din2(G160_p_spl_101)
  );


  FA
  g_g1181_n
  (
    .dout(g1181_n),
    .din1(g1179_p),
    .din2(g1180_p)
  );


  LA
  g_g1182_p
  (
    .dout(g1182_p),
    .din1(G161_n_spl_10),
    .din2(g1181_n)
  );


  LA
  g_g1183_p
  (
    .dout(g1183_p),
    .din1(G160_p_spl_101),
    .din2(g997_n_spl_1)
  );


  LA
  g_g1184_p
  (
    .dout(g1184_p),
    .din1(G160_n_spl_101),
    .din2(g1032_n_spl_1)
  );


  FA
  g_g1185_n
  (
    .dout(g1185_n),
    .din1(g1183_p),
    .din2(g1184_p)
  );


  LA
  g_g1186_p
  (
    .dout(g1186_p),
    .din1(G161_p_spl_10),
    .din2(g1185_n)
  );


  FA
  g_g1187_n
  (
    .dout(g1187_n),
    .din1(g1182_p),
    .din2(g1186_p)
  );


  LA
  g_g1188_p
  (
    .dout(g1188_p),
    .din1(G64_p_spl_110),
    .din2(g1187_n)
  );


  FA
  g_g1189_n
  (
    .dout(g1189_n),
    .din1(G160_p_spl_110),
    .din2(g1025_n_spl_1)
  );


  FA
  g_g1190_n
  (
    .dout(g1190_n),
    .din1(G160_n_spl_110),
    .din2(g990_p_spl_1)
  );


  LA
  g_g1191_p
  (
    .dout(g1191_p),
    .din1(G161_p_spl_11),
    .din2(g1190_n)
  );


  LA
  g_g1192_p
  (
    .dout(g1192_p),
    .din1(g1189_n),
    .din2(g1191_p)
  );


  LA
  g_g1193_p
  (
    .dout(g1193_p),
    .din1(G73_p_spl_),
    .din2(G160_n_spl_110)
  );


  LA
  g_g1194_p
  (
    .dout(g1194_p),
    .din1(G83_p_spl_),
    .din2(G160_p_spl_110)
  );


  FA
  g_g1195_n
  (
    .dout(g1195_n),
    .din1(g1193_p),
    .din2(g1194_p)
  );


  LA
  g_g1196_p
  (
    .dout(g1196_p),
    .din1(G161_n_spl_11),
    .din2(g1195_n)
  );


  FA
  g_g1197_n
  (
    .dout(g1197_n),
    .din1(g1192_p),
    .din2(g1196_p)
  );


  LA
  g_g1198_p
  (
    .dout(g1198_p),
    .din1(G64_p_spl_111),
    .din2(g1197_n)
  );


  LA
  g_g1199_p
  (
    .dout(g1199_p),
    .din1(g258_n_spl_),
    .din2(g267_n_spl_)
  );


  FA
  g_g1199_n
  (
    .dout(g1199_n),
    .din1(g258_p_spl_),
    .din2(g267_p_spl_)
  );


  LA
  g_g1200_p
  (
    .dout(g1200_p),
    .din1(g268_n_spl_),
    .din2(g1199_n)
  );


  FA
  g_g1200_n
  (
    .dout(g1200_n),
    .din1(g268_p),
    .din2(g1199_p)
  );


  LA
  g_g1201_p
  (
    .dout(g1201_p),
    .din1(g237_p_spl_),
    .din2(g240_n_spl_)
  );


  FA
  g_g1201_n
  (
    .dout(g1201_n),
    .din1(g237_n_spl_1),
    .din2(g240_p_spl_)
  );


  LA
  g_g1202_p
  (
    .dout(g1202_p),
    .din1(g241_n_spl_),
    .din2(g1201_n)
  );


  FA
  g_g1202_n
  (
    .dout(g1202_n),
    .din1(g241_p),
    .din2(g1201_p)
  );


  LA
  g_g1203_p
  (
    .dout(g1203_p),
    .din1(g1200_p_spl_),
    .din2(g1202_n_spl_)
  );


  FA
  g_g1203_n
  (
    .dout(g1203_n),
    .din1(g1200_n_spl_),
    .din2(g1202_p_spl_)
  );


  LA
  g_g1204_p
  (
    .dout(g1204_p),
    .din1(g1200_n_spl_),
    .din2(g1202_p_spl_)
  );


  FA
  g_g1204_n
  (
    .dout(g1204_n),
    .din1(g1200_p_spl_),
    .din2(g1202_n_spl_)
  );


  LA
  g_g1205_p
  (
    .dout(g1205_p),
    .din1(g1203_n),
    .din2(g1204_n)
  );


  FA
  g_g1205_n
  (
    .dout(g1205_n),
    .din1(g1203_p),
    .din2(g1204_p)
  );


  LA
  g_g1206_p
  (
    .dout(g1206_p),
    .din1(G101_p_spl_010),
    .din2(G128_p_spl_10)
  );


  FA
  g_g1206_n
  (
    .dout(g1206_n),
    .din1(G101_n_spl_010),
    .din2(G128_n_spl_10)
  );


  LA
  g_g1207_p
  (
    .dout(g1207_p),
    .din1(G100_p_spl_010),
    .din2(G128_n_spl_10)
  );


  FA
  g_g1207_n
  (
    .dout(g1207_n),
    .din1(G100_n_spl_010),
    .din2(G128_p_spl_10)
  );


  LA
  g_g1208_p
  (
    .dout(g1208_p),
    .din1(g1206_n),
    .din2(g1207_n)
  );


  FA
  g_g1208_n
  (
    .dout(g1208_n),
    .din1(g1206_p),
    .din2(g1207_p)
  );


  LA
  g_g1209_p
  (
    .dout(g1209_p),
    .din1(G150_p_spl_1),
    .din2(g1208_n)
  );


  FA
  g_g1209_n
  (
    .dout(g1209_n),
    .din1(G150_n_spl_1),
    .din2(g1208_p)
  );


  LA
  g_g1210_p
  (
    .dout(g1210_p),
    .din1(G102_n_spl_010),
    .din2(G128_p_spl_11)
  );


  FA
  g_g1210_n
  (
    .dout(g1210_n),
    .din1(G102_p_spl_010),
    .din2(G128_n_spl_11)
  );


  LA
  g_g1211_p
  (
    .dout(g1211_p),
    .din1(G98_n_spl_010),
    .din2(G128_n_spl_11)
  );


  FA
  g_g1211_n
  (
    .dout(g1211_n),
    .din1(G98_p_spl_010),
    .din2(G128_p_spl_11)
  );


  LA
  g_g1212_p
  (
    .dout(g1212_p),
    .din1(g1210_n),
    .din2(g1211_n)
  );


  FA
  g_g1212_n
  (
    .dout(g1212_n),
    .din1(g1210_p),
    .din2(g1211_p)
  );


  LA
  g_g1213_p
  (
    .dout(g1213_p),
    .din1(G150_n_spl_1),
    .din2(g1212_n)
  );


  FA
  g_g1213_n
  (
    .dout(g1213_n),
    .din1(G150_p_spl_1),
    .din2(g1212_p)
  );


  LA
  g_g1214_p
  (
    .dout(g1214_p),
    .din1(g1209_n),
    .din2(g1213_n)
  );


  FA
  g_g1214_n
  (
    .dout(g1214_n),
    .din1(g1209_p),
    .din2(g1213_p)
  );


  LA
  g_g1215_p
  (
    .dout(g1215_p),
    .din1(G101_p_spl_011),
    .din2(G126_p_spl_10)
  );


  FA
  g_g1215_n
  (
    .dout(g1215_n),
    .din1(G101_n_spl_011),
    .din2(G126_n_spl_10)
  );


  LA
  g_g1216_p
  (
    .dout(g1216_p),
    .din1(G100_p_spl_010),
    .din2(G126_n_spl_10)
  );


  FA
  g_g1216_n
  (
    .dout(g1216_n),
    .din1(G100_n_spl_010),
    .din2(G126_p_spl_10)
  );


  LA
  g_g1217_p
  (
    .dout(g1217_p),
    .din1(g1215_n),
    .din2(g1216_n)
  );


  FA
  g_g1217_n
  (
    .dout(g1217_n),
    .din1(g1215_p),
    .din2(g1216_p)
  );


  LA
  g_g1218_p
  (
    .dout(g1218_p),
    .din1(G149_p_spl_1),
    .din2(g1217_n)
  );


  FA
  g_g1218_n
  (
    .dout(g1218_n),
    .din1(G149_n_spl_1),
    .din2(g1217_p)
  );


  LA
  g_g1219_p
  (
    .dout(g1219_p),
    .din1(G102_n_spl_010),
    .din2(G126_p_spl_11)
  );


  FA
  g_g1219_n
  (
    .dout(g1219_n),
    .din1(G102_p_spl_010),
    .din2(G126_n_spl_11)
  );


  LA
  g_g1220_p
  (
    .dout(g1220_p),
    .din1(G98_n_spl_010),
    .din2(G126_n_spl_11)
  );


  FA
  g_g1220_n
  (
    .dout(g1220_n),
    .din1(G98_p_spl_010),
    .din2(G126_p_spl_11)
  );


  LA
  g_g1221_p
  (
    .dout(g1221_p),
    .din1(g1219_n),
    .din2(g1220_n)
  );


  FA
  g_g1221_n
  (
    .dout(g1221_n),
    .din1(g1219_p),
    .din2(g1220_p)
  );


  LA
  g_g1222_p
  (
    .dout(g1222_p),
    .din1(G149_n_spl_1),
    .din2(g1221_n)
  );


  FA
  g_g1222_n
  (
    .dout(g1222_n),
    .din1(G149_p_spl_1),
    .din2(g1221_p)
  );


  LA
  g_g1223_p
  (
    .dout(g1223_p),
    .din1(g1218_n),
    .din2(g1222_n)
  );


  FA
  g_g1223_n
  (
    .dout(g1223_n),
    .din1(g1218_p),
    .din2(g1222_p)
  );


  LA
  g_g1224_p
  (
    .dout(g1224_p),
    .din1(g1214_n_spl_),
    .din2(g1223_p_spl_)
  );


  FA
  g_g1224_n
  (
    .dout(g1224_n),
    .din1(g1214_p_spl_),
    .din2(g1223_n_spl_)
  );


  LA
  g_g1225_p
  (
    .dout(g1225_p),
    .din1(g1214_p_spl_),
    .din2(g1223_n_spl_)
  );


  FA
  g_g1225_n
  (
    .dout(g1225_n),
    .din1(g1214_n_spl_),
    .din2(g1223_p_spl_)
  );


  LA
  g_g1226_p
  (
    .dout(g1226_p),
    .din1(g1224_n),
    .din2(g1225_n)
  );


  FA
  g_g1226_n
  (
    .dout(g1226_n),
    .din1(g1224_p),
    .din2(g1225_p)
  );


  LA
  g_g1227_p
  (
    .dout(g1227_p),
    .din1(G98_n_spl_011),
    .din2(G148_n_spl_1)
  );


  FA
  g_g1227_n
  (
    .dout(g1227_n),
    .din1(G98_p_spl_011),
    .din2(G148_p_spl_1)
  );


  LA
  g_g1228_p
  (
    .dout(g1228_p),
    .din1(G100_p_spl_011),
    .din2(G148_p_spl_1)
  );


  FA
  g_g1228_n
  (
    .dout(g1228_n),
    .din1(G100_n_spl_011),
    .din2(G148_n_spl_1)
  );


  LA
  g_g1229_p
  (
    .dout(g1229_p),
    .din1(g1227_n),
    .din2(g1228_n)
  );


  FA
  g_g1229_n
  (
    .dout(g1229_n),
    .din1(g1227_p),
    .din2(g1228_p)
  );


  LA
  g_g1230_p
  (
    .dout(g1230_p),
    .din1(G101_p_spl_011),
    .din2(G121_p_spl_10)
  );


  FA
  g_g1230_n
  (
    .dout(g1230_n),
    .din1(G101_n_spl_011),
    .din2(G121_n_spl_10)
  );


  LA
  g_g1231_p
  (
    .dout(g1231_p),
    .din1(G100_p_spl_011),
    .din2(G121_n_spl_10)
  );


  FA
  g_g1231_n
  (
    .dout(g1231_n),
    .din1(G100_n_spl_011),
    .din2(G121_p_spl_10)
  );


  LA
  g_g1232_p
  (
    .dout(g1232_p),
    .din1(g1230_n),
    .din2(g1231_n)
  );


  FA
  g_g1232_n
  (
    .dout(g1232_n),
    .din1(g1230_p),
    .din2(g1231_p)
  );


  LA
  g_g1233_p
  (
    .dout(g1233_p),
    .din1(G147_p_spl_1),
    .din2(g1232_n)
  );


  FA
  g_g1233_n
  (
    .dout(g1233_n),
    .din1(G147_n_spl_1),
    .din2(g1232_p)
  );


  LA
  g_g1234_p
  (
    .dout(g1234_p),
    .din1(G102_n_spl_011),
    .din2(G121_p_spl_11)
  );


  FA
  g_g1234_n
  (
    .dout(g1234_n),
    .din1(G102_p_spl_011),
    .din2(G121_n_spl_11)
  );


  LA
  g_g1235_p
  (
    .dout(g1235_p),
    .din1(G98_n_spl_011),
    .din2(G121_n_spl_11)
  );


  FA
  g_g1235_n
  (
    .dout(g1235_n),
    .din1(G98_p_spl_011),
    .din2(G121_p_spl_11)
  );


  LA
  g_g1236_p
  (
    .dout(g1236_p),
    .din1(g1234_n),
    .din2(g1235_n)
  );


  FA
  g_g1236_n
  (
    .dout(g1236_n),
    .din1(g1234_p),
    .din2(g1235_p)
  );


  LA
  g_g1237_p
  (
    .dout(g1237_p),
    .din1(G147_n_spl_1),
    .din2(g1236_n)
  );


  FA
  g_g1237_n
  (
    .dout(g1237_n),
    .din1(G147_p_spl_1),
    .din2(g1236_p)
  );


  LA
  g_g1238_p
  (
    .dout(g1238_p),
    .din1(g1233_n),
    .din2(g1237_n)
  );


  FA
  g_g1238_n
  (
    .dout(g1238_n),
    .din1(g1233_p),
    .din2(g1237_p)
  );


  LA
  g_g1239_p
  (
    .dout(g1239_p),
    .din1(g1229_n_spl_),
    .din2(g1238_p_spl_)
  );


  FA
  g_g1239_n
  (
    .dout(g1239_n),
    .din1(g1229_p_spl_),
    .din2(g1238_n_spl_)
  );


  LA
  g_g1240_p
  (
    .dout(g1240_p),
    .din1(g1229_p_spl_),
    .din2(g1238_n_spl_)
  );


  FA
  g_g1240_n
  (
    .dout(g1240_n),
    .din1(g1229_n_spl_),
    .din2(g1238_p_spl_)
  );


  LA
  g_g1241_p
  (
    .dout(g1241_p),
    .din1(g1239_n),
    .din2(g1240_n)
  );


  FA
  g_g1241_n
  (
    .dout(g1241_n),
    .din1(g1239_p),
    .din2(g1240_p)
  );


  LA
  g_g1242_p
  (
    .dout(g1242_p),
    .din1(g245_n_spl_1),
    .din2(g1241_p_spl_)
  );


  FA
  g_g1242_n
  (
    .dout(g1242_n),
    .din1(g245_p_spl_),
    .din2(g1241_n_spl_)
  );


  LA
  g_g1243_p
  (
    .dout(g1243_p),
    .din1(g245_p_spl_),
    .din2(g1241_n_spl_)
  );


  FA
  g_g1243_n
  (
    .dout(g1243_n),
    .din1(g245_n_spl_1),
    .din2(g1241_p_spl_)
  );


  LA
  g_g1244_p
  (
    .dout(g1244_p),
    .din1(g1242_n),
    .din2(g1243_n)
  );


  FA
  g_g1244_n
  (
    .dout(g1244_n),
    .din1(g1242_p),
    .din2(g1243_p)
  );


  LA
  g_g1245_p
  (
    .dout(g1245_p),
    .din1(g1226_p_spl_),
    .din2(g1244_n_spl_)
  );


  FA
  g_g1245_n
  (
    .dout(g1245_n),
    .din1(g1226_n_spl_),
    .din2(g1244_p_spl_)
  );


  LA
  g_g1246_p
  (
    .dout(g1246_p),
    .din1(g1226_n_spl_),
    .din2(g1244_p_spl_)
  );


  FA
  g_g1246_n
  (
    .dout(g1246_n),
    .din1(g1226_p_spl_),
    .din2(g1244_n_spl_)
  );


  LA
  g_g1247_p
  (
    .dout(g1247_p),
    .din1(g1245_n),
    .din2(g1246_n)
  );


  FA
  g_g1247_n
  (
    .dout(g1247_n),
    .din1(g1245_p),
    .din2(g1246_p)
  );


  FA
  g_g1248_n
  (
    .dout(g1248_n),
    .din1(g1205_p),
    .din2(g1247_n)
  );


  FA
  g_g1249_n
  (
    .dout(g1249_n),
    .din1(g1205_n),
    .din2(g1247_p)
  );


  LA
  g_g1250_p
  (
    .dout(g1250_p),
    .din1(g1248_n),
    .din2(g1249_n)
  );


  FA
  g_g1251_n
  (
    .dout(g1251_n),
    .din1(G176_n_spl_110),
    .din2(g1250_p)
  );


  LA
  g_g1252_p
  (
    .dout(g1252_p),
    .din1(g464_n_spl_10),
    .din2(g596_n_spl_0)
  );


  FA
  g_g1252_n
  (
    .dout(g1252_n),
    .din1(g464_p_spl_10),
    .din2(g596_p_spl_1)
  );


  LA
  g_g1253_p
  (
    .dout(g1253_p),
    .din1(g464_p_spl_1),
    .din2(g596_p_spl_1)
  );


  FA
  g_g1253_n
  (
    .dout(g1253_n),
    .din1(g464_n_spl_1),
    .din2(g596_n_spl_)
  );


  LA
  g_g1254_p
  (
    .dout(g1254_p),
    .din1(g1252_n),
    .din2(g1253_n)
  );


  FA
  g_g1254_n
  (
    .dout(g1254_n),
    .din1(g1252_p),
    .din2(g1253_p)
  );


  LA
  g_g1255_p
  (
    .dout(g1255_p),
    .din1(g617_p_spl_0),
    .din2(g1254_n_spl_)
  );


  FA
  g_g1255_n
  (
    .dout(g1255_n),
    .din1(g617_n_spl_),
    .din2(g1254_p_spl_)
  );


  LA
  g_g1256_p
  (
    .dout(g1256_p),
    .din1(g617_n_spl_),
    .din2(g1254_p_spl_)
  );


  FA
  g_g1256_n
  (
    .dout(g1256_n),
    .din1(g617_p_spl_),
    .din2(g1254_n_spl_)
  );


  LA
  g_g1257_p
  (
    .dout(g1257_p),
    .din1(g1255_n),
    .din2(g1256_n)
  );


  FA
  g_g1257_n
  (
    .dout(g1257_n),
    .din1(g1255_p),
    .din2(g1256_p)
  );


  LA
  g_g1258_p
  (
    .dout(g1258_p),
    .din1(g598_p_spl_0),
    .din2(g1257_p_spl_)
  );


  FA
  g_g1258_n
  (
    .dout(g1258_n),
    .din1(g598_n_spl_0),
    .din2(g1257_n_spl_)
  );


  LA
  g_g1259_p
  (
    .dout(g1259_p),
    .din1(g598_n_spl_),
    .din2(g1257_n_spl_)
  );


  FA
  g_g1259_n
  (
    .dout(g1259_n),
    .din1(g598_p_spl_),
    .din2(g1257_p_spl_)
  );


  LA
  g_g1260_p
  (
    .dout(g1260_p),
    .din1(g1258_n),
    .din2(g1259_n)
  );


  FA
  g_g1260_n
  (
    .dout(g1260_n),
    .din1(g1258_p),
    .din2(g1259_p)
  );


  LA
  g_g1261_p
  (
    .dout(g1261_p),
    .din1(G162_n_spl_),
    .din2(g562_p)
  );


  FA
  g_g1261_n
  (
    .dout(g1261_n),
    .din1(G162_p_spl_),
    .din2(g562_n_spl_)
  );


  LA
  g_g1262_p
  (
    .dout(g1262_p),
    .din1(G162_p_spl_),
    .din2(g461_n_spl_)
  );


  FA
  g_g1262_n
  (
    .dout(g1262_n),
    .din1(G162_n_spl_),
    .din2(g461_p_spl_)
  );


  LA
  g_g1263_p
  (
    .dout(g1263_p),
    .din1(g1261_n),
    .din2(g1262_n)
  );


  FA
  g_g1263_n
  (
    .dout(g1263_n),
    .din1(g1261_p),
    .din2(g1262_p)
  );


  LA
  g_g1264_p
  (
    .dout(g1264_p),
    .din1(g1260_p_spl_),
    .din2(g1263_p_spl_)
  );


  FA
  g_g1264_n
  (
    .dout(g1264_n),
    .din1(g1260_n_spl_),
    .din2(g1263_n_spl_)
  );


  LA
  g_g1265_p
  (
    .dout(g1265_p),
    .din1(g1260_n_spl_),
    .din2(g1263_n_spl_)
  );


  FA
  g_g1265_n
  (
    .dout(g1265_n),
    .din1(g1260_p_spl_),
    .din2(g1263_p_spl_)
  );


  LA
  g_g1266_p
  (
    .dout(g1266_p),
    .din1(g1264_n),
    .din2(g1265_n)
  );


  FA
  g_g1266_n
  (
    .dout(g1266_n),
    .din1(g1264_p),
    .din2(g1265_p)
  );


  LA
  g_g1267_p
  (
    .dout(g1267_p),
    .din1(g450_n_spl_1),
    .din2(g454_n_spl_1)
  );


  FA
  g_g1267_n
  (
    .dout(g1267_n),
    .din1(g450_p_spl_1),
    .din2(g454_p_spl_1)
  );


  LA
  g_g1268_p
  (
    .dout(g1268_p),
    .din1(g455_n_spl_),
    .din2(g1267_n)
  );


  FA
  g_g1268_n
  (
    .dout(g1268_n),
    .din1(g455_p_spl_),
    .din2(g1267_p)
  );


  LA
  g_g1269_p
  (
    .dout(g1269_p),
    .din1(g471_p_spl_1),
    .din2(g1268_n_spl_)
  );


  FA
  g_g1269_n
  (
    .dout(g1269_n),
    .din1(g471_n_spl_1),
    .din2(g1268_p_spl_)
  );


  LA
  g_g1270_p
  (
    .dout(g1270_p),
    .din1(g471_n_spl_1),
    .din2(g1268_p_spl_)
  );


  FA
  g_g1270_n
  (
    .dout(g1270_n),
    .din1(g471_p_spl_1),
    .din2(g1268_n_spl_)
  );


  LA
  g_g1271_p
  (
    .dout(g1271_p),
    .din1(g1269_n),
    .din2(g1270_n)
  );


  FA
  g_g1271_n
  (
    .dout(g1271_n),
    .din1(g1269_p),
    .din2(g1270_p)
  );


  LA
  g_g1272_p
  (
    .dout(g1272_p),
    .din1(g1266_n_spl_),
    .din2(g1271_n_spl_)
  );


  FA
  g_g1272_n
  (
    .dout(g1272_n),
    .din1(g1266_p_spl_),
    .din2(g1271_p_spl_)
  );


  LA
  g_g1273_p
  (
    .dout(g1273_p),
    .din1(g1266_p_spl_),
    .din2(g1271_p_spl_)
  );


  FA
  g_g1273_n
  (
    .dout(g1273_n),
    .din1(g1266_n_spl_),
    .din2(g1271_n_spl_)
  );


  LA
  g_g1274_p
  (
    .dout(g1274_p),
    .din1(g1272_n),
    .din2(g1273_n)
  );


  FA
  g_g1274_n
  (
    .dout(g1274_n),
    .din1(g1272_p),
    .din2(g1273_p)
  );


  LA
  g_g1275_p
  (
    .dout(g1275_p),
    .din1(g444_n_spl_),
    .din2(g780_p_spl_0)
  );


  FA
  g_g1275_n
  (
    .dout(g1275_n),
    .din1(g444_p_spl_),
    .din2(g780_n_spl_0)
  );


  LA
  g_g1276_p
  (
    .dout(g1276_p),
    .din1(g442_n_spl_1),
    .din2(g1275_n_spl_)
  );


  FA
  g_g1276_n
  (
    .dout(g1276_n),
    .din1(g442_p_spl_1),
    .din2(g1275_p_spl_)
  );


  LA
  g_g1277_p
  (
    .dout(g1277_p),
    .din1(g442_p_spl_1),
    .din2(g1275_p_spl_)
  );


  FA
  g_g1277_n
  (
    .dout(g1277_n),
    .din1(g442_n_spl_1),
    .din2(g1275_n_spl_)
  );


  LA
  g_g1278_p
  (
    .dout(g1278_p),
    .din1(g1276_n),
    .din2(g1277_n)
  );


  FA
  g_g1278_n
  (
    .dout(g1278_n),
    .din1(g1276_p),
    .din2(g1277_p)
  );


  LA
  g_g1279_p
  (
    .dout(g1279_p),
    .din1(g479_n_spl_01),
    .din2(g1278_p_spl_)
  );


  FA
  g_g1279_n
  (
    .dout(g1279_n),
    .din1(g479_p_spl_01),
    .din2(g1278_n_spl_)
  );


  LA
  g_g1280_p
  (
    .dout(g1280_p),
    .din1(g479_p_spl_10),
    .din2(g1278_n_spl_)
  );


  FA
  g_g1280_n
  (
    .dout(g1280_n),
    .din1(g479_n_spl_10),
    .din2(g1278_p_spl_)
  );


  LA
  g_g1281_p
  (
    .dout(g1281_p),
    .din1(g1279_n),
    .din2(g1280_n)
  );


  FA
  g_g1281_n
  (
    .dout(g1281_n),
    .din1(g1279_p),
    .din2(g1280_p)
  );


  LA
  g_g1282_p
  (
    .dout(g1282_p),
    .din1(g443_n_spl_0),
    .din2(g1281_p_spl_)
  );


  FA
  g_g1282_n
  (
    .dout(g1282_n),
    .din1(g443_p_spl_0),
    .din2(g1281_n_spl_)
  );


  LA
  g_g1283_p
  (
    .dout(g1283_p),
    .din1(g443_p_spl_1),
    .din2(g1281_n_spl_)
  );


  FA
  g_g1283_n
  (
    .dout(g1283_n),
    .din1(g443_n_spl_1),
    .din2(g1281_p_spl_)
  );


  LA
  g_g1284_p
  (
    .dout(g1284_p),
    .din1(g1282_n_spl_),
    .din2(g1283_n)
  );


  FA
  g_g1284_n
  (
    .dout(g1284_n),
    .din1(g1282_p_spl_),
    .din2(g1283_p)
  );


  LA
  g_g1285_p
  (
    .dout(g1285_p),
    .din1(g437_p_spl_01),
    .din2(g1284_n_spl_)
  );


  FA
  g_g1285_n
  (
    .dout(g1285_n),
    .din1(g437_n_spl_01),
    .din2(g1284_p_spl_)
  );


  LA
  g_g1286_p
  (
    .dout(g1286_p),
    .din1(g441_p_spl_1),
    .din2(g780_n_spl_1)
  );


  FA
  g_g1286_n
  (
    .dout(g1286_n),
    .din1(g441_n_spl_1),
    .din2(g780_p_spl_1)
  );


  LA
  g_g1287_p
  (
    .dout(g1287_p),
    .din1(g441_n_spl_1),
    .din2(g780_p_spl_1)
  );


  FA
  g_g1287_n
  (
    .dout(g1287_n),
    .din1(g441_p_spl_1),
    .din2(g780_n_spl_1)
  );


  LA
  g_g1288_p
  (
    .dout(g1288_p),
    .din1(g1286_n),
    .din2(g1287_n)
  );


  FA
  g_g1288_n
  (
    .dout(g1288_n),
    .din1(g1286_p),
    .din2(g1287_p)
  );


  LA
  g_g1289_p
  (
    .dout(g1289_p),
    .din1(g479_p_spl_10),
    .din2(g1288_n_spl_)
  );


  FA
  g_g1289_n
  (
    .dout(g1289_n),
    .din1(g479_n_spl_10),
    .din2(g1288_p_spl_)
  );


  LA
  g_g1290_p
  (
    .dout(g1290_p),
    .din1(g479_n_spl_1),
    .din2(g1288_p_spl_)
  );


  FA
  g_g1290_n
  (
    .dout(g1290_n),
    .din1(g479_p_spl_1),
    .din2(g1288_n_spl_)
  );


  LA
  g_g1291_p
  (
    .dout(g1291_p),
    .din1(g1289_n),
    .din2(g1290_n)
  );


  FA
  g_g1291_n
  (
    .dout(g1291_n),
    .din1(g1289_p),
    .din2(g1290_p)
  );


  LA
  g_g1292_p
  (
    .dout(g1292_p),
    .din1(g443_p_spl_1),
    .din2(g1291_n)
  );


  FA
  g_g1292_n
  (
    .dout(g1292_n),
    .din1(g443_n_spl_1),
    .din2(g1291_p)
  );


  LA
  g_g1293_p
  (
    .dout(g1293_p),
    .din1(g437_n_spl_1),
    .din2(g1292_n)
  );


  FA
  g_g1293_n
  (
    .dout(g1293_n),
    .din1(g437_p_spl_1),
    .din2(g1292_p)
  );


  LA
  g_g1294_p
  (
    .dout(g1294_p),
    .din1(g1282_n_spl_),
    .din2(g1293_p)
  );


  FA
  g_g1294_n
  (
    .dout(g1294_n),
    .din1(g1282_p_spl_),
    .din2(g1293_n)
  );


  LA
  g_g1295_p
  (
    .dout(g1295_p),
    .din1(g774_p_spl_1),
    .din2(g1294_p)
  );


  FA
  g_g1295_n
  (
    .dout(g1295_n),
    .din1(g774_n_spl_1),
    .din2(g1294_n)
  );


  LA
  g_g1296_p
  (
    .dout(g1296_p),
    .din1(g1285_n),
    .din2(g1295_n)
  );


  FA
  g_g1296_n
  (
    .dout(g1296_n),
    .din1(g1285_p),
    .din2(g1295_p)
  );


  LA
  g_g1297_p
  (
    .dout(g1297_p),
    .din1(g437_n_spl_1),
    .din2(g774_n_spl_1)
  );


  FA
  g_g1297_n
  (
    .dout(g1297_n),
    .din1(g437_p_spl_1),
    .din2(g774_p_spl_1)
  );


  LA
  g_g1298_p
  (
    .dout(g1298_p),
    .din1(g1284_p_spl_),
    .din2(g1297_p)
  );


  FA
  g_g1298_n
  (
    .dout(g1298_n),
    .din1(g1284_n_spl_),
    .din2(g1297_n)
  );


  LA
  g_g1299_p
  (
    .dout(g1299_p),
    .din1(g1296_p),
    .din2(g1298_n)
  );


  FA
  g_g1299_n
  (
    .dout(g1299_n),
    .din1(g1296_n),
    .din2(g1298_p)
  );


  LA
  g_g1300_p
  (
    .dout(g1300_p),
    .din1(g581_p_spl_01),
    .din2(g1299_p_spl_)
  );


  FA
  g_g1300_n
  (
    .dout(g1300_n),
    .din1(g581_n_spl_11),
    .din2(g1299_n_spl_)
  );


  LA
  g_g1301_p
  (
    .dout(g1301_p),
    .din1(g581_n_spl_11),
    .din2(g1299_n_spl_)
  );


  FA
  g_g1301_n
  (
    .dout(g1301_n),
    .din1(g581_p_spl_1),
    .din2(g1299_p_spl_)
  );


  LA
  g_g1302_p
  (
    .dout(g1302_p),
    .din1(g1300_n),
    .din2(g1301_n)
  );


  FA
  g_g1302_n
  (
    .dout(g1302_n),
    .din1(g1300_p),
    .din2(g1301_p)
  );


  LA
  g_g1303_p
  (
    .dout(g1303_p),
    .din1(g1274_p),
    .din2(g1302_n)
  );


  LA
  g_g1304_p
  (
    .dout(g1304_p),
    .din1(g1274_n),
    .din2(g1302_p)
  );


  FA
  g_g1305_n
  (
    .dout(g1305_n),
    .din1(G176_p_spl_1111),
    .din2(g1304_p)
  );


  FA
  g_g1306_n
  (
    .dout(g1306_n),
    .din1(g1303_p),
    .din2(g1305_n)
  );


  LA
  g_g1307_p
  (
    .dout(g1307_p),
    .din1(g1251_n),
    .din2(g1306_n)
  );


  FA
  g_g1308_n
  (
    .dout(g1308_n),
    .din1(G177_n_spl_111),
    .din2(g1307_p)
  );


  FA
  g_g1309_n
  (
    .dout(g1309_n),
    .din1(G51_p),
    .din2(G177_p_spl_110)
  );


  FA
  g_g1310_n
  (
    .dout(g1310_n),
    .din1(G176_n_spl_110),
    .din2(g1309_n)
  );


  LA
  g_g1311_p
  (
    .dout(g1311_p),
    .din1(g1308_n_spl_),
    .din2(g1310_n)
  );


  LA
  g_g1312_p
  (
    .dout(g1312_p),
    .din1(G94_p_spl_10),
    .din2(G101_p_spl_100)
  );


  FA
  g_g1312_n
  (
    .dout(g1312_n),
    .din1(G94_n_spl_10),
    .din2(G101_n_spl_100)
  );


  LA
  g_g1313_p
  (
    .dout(g1313_p),
    .din1(G94_n_spl_10),
    .din2(G100_p_spl_100)
  );


  FA
  g_g1313_n
  (
    .dout(g1313_n),
    .din1(G94_p_spl_10),
    .din2(G100_n_spl_100)
  );


  LA
  g_g1314_p
  (
    .dout(g1314_p),
    .din1(g1312_n),
    .din2(g1313_n)
  );


  FA
  g_g1314_n
  (
    .dout(g1314_n),
    .din1(g1312_p),
    .din2(g1313_p)
  );


  LA
  g_g1315_p
  (
    .dout(g1315_p),
    .din1(G140_p_spl_1),
    .din2(g1314_n)
  );


  FA
  g_g1315_n
  (
    .dout(g1315_n),
    .din1(G140_n_spl_1),
    .din2(g1314_p)
  );


  LA
  g_g1316_p
  (
    .dout(g1316_p),
    .din1(G94_p_spl_11),
    .din2(G102_n_spl_011)
  );


  FA
  g_g1316_n
  (
    .dout(g1316_n),
    .din1(G94_n_spl_11),
    .din2(G102_p_spl_011)
  );


  LA
  g_g1317_p
  (
    .dout(g1317_p),
    .din1(G94_n_spl_11),
    .din2(G98_n_spl_100)
  );


  FA
  g_g1317_n
  (
    .dout(g1317_n),
    .din1(G94_p_spl_11),
    .din2(G98_p_spl_100)
  );


  LA
  g_g1318_p
  (
    .dout(g1318_p),
    .din1(g1316_n),
    .din2(g1317_n)
  );


  FA
  g_g1318_n
  (
    .dout(g1318_n),
    .din1(g1316_p),
    .din2(g1317_p)
  );


  LA
  g_g1319_p
  (
    .dout(g1319_p),
    .din1(G140_n_spl_1),
    .din2(g1318_n)
  );


  FA
  g_g1319_n
  (
    .dout(g1319_n),
    .din1(G140_p_spl_1),
    .din2(g1318_p)
  );


  LA
  g_g1320_p
  (
    .dout(g1320_p),
    .din1(g1315_n),
    .din2(g1319_n)
  );


  FA
  g_g1320_n
  (
    .dout(g1320_n),
    .din1(g1315_p),
    .din2(g1319_p)
  );


  LA
  g_g1321_p
  (
    .dout(g1321_p),
    .din1(G92_p_spl_10),
    .din2(G101_p_spl_100)
  );


  FA
  g_g1321_n
  (
    .dout(g1321_n),
    .din1(G92_n_spl_10),
    .din2(G101_n_spl_100)
  );


  LA
  g_g1322_p
  (
    .dout(g1322_p),
    .din1(G92_n_spl_10),
    .din2(G100_p_spl_100)
  );


  FA
  g_g1322_n
  (
    .dout(g1322_n),
    .din1(G92_p_spl_10),
    .din2(G100_n_spl_100)
  );


  LA
  g_g1323_p
  (
    .dout(g1323_p),
    .din1(g1321_n),
    .din2(g1322_n)
  );


  FA
  g_g1323_n
  (
    .dout(g1323_n),
    .din1(g1321_p),
    .din2(g1322_p)
  );


  LA
  g_g1324_p
  (
    .dout(g1324_p),
    .din1(G144_p_spl_1),
    .din2(g1323_n)
  );


  FA
  g_g1324_n
  (
    .dout(g1324_n),
    .din1(G144_n_spl_1),
    .din2(g1323_p)
  );


  LA
  g_g1325_p
  (
    .dout(g1325_p),
    .din1(G92_p_spl_11),
    .din2(G102_n_spl_100)
  );


  FA
  g_g1325_n
  (
    .dout(g1325_n),
    .din1(G92_n_spl_11),
    .din2(G102_p_spl_100)
  );


  LA
  g_g1326_p
  (
    .dout(g1326_p),
    .din1(G92_n_spl_11),
    .din2(G98_n_spl_100)
  );


  FA
  g_g1326_n
  (
    .dout(g1326_n),
    .din1(G92_p_spl_11),
    .din2(G98_p_spl_100)
  );


  LA
  g_g1327_p
  (
    .dout(g1327_p),
    .din1(g1325_n),
    .din2(g1326_n)
  );


  FA
  g_g1327_n
  (
    .dout(g1327_n),
    .din1(g1325_p),
    .din2(g1326_p)
  );


  LA
  g_g1328_p
  (
    .dout(g1328_p),
    .din1(G144_n_spl_1),
    .din2(g1327_n)
  );


  FA
  g_g1328_n
  (
    .dout(g1328_n),
    .din1(G144_p_spl_1),
    .din2(g1327_p)
  );


  LA
  g_g1329_p
  (
    .dout(g1329_p),
    .din1(g1324_n),
    .din2(g1328_n)
  );


  FA
  g_g1329_n
  (
    .dout(g1329_n),
    .din1(g1324_p),
    .din2(g1328_p)
  );


  LA
  g_g1330_p
  (
    .dout(g1330_p),
    .din1(g1320_n_spl_),
    .din2(g1329_p_spl_)
  );


  FA
  g_g1330_n
  (
    .dout(g1330_n),
    .din1(g1320_p_spl_),
    .din2(g1329_n_spl_)
  );


  LA
  g_g1331_p
  (
    .dout(g1331_p),
    .din1(g1320_p_spl_),
    .din2(g1329_n_spl_)
  );


  FA
  g_g1331_n
  (
    .dout(g1331_n),
    .din1(g1320_n_spl_),
    .din2(g1329_p_spl_)
  );


  LA
  g_g1332_p
  (
    .dout(g1332_p),
    .din1(g1330_n),
    .din2(g1331_n)
  );


  FA
  g_g1332_n
  (
    .dout(g1332_n),
    .din1(g1330_p),
    .din2(g1331_p)
  );


  LA
  g_g1333_p
  (
    .dout(g1333_p),
    .din1(G90_p_spl_10),
    .din2(G101_p_spl_101)
  );


  FA
  g_g1333_n
  (
    .dout(g1333_n),
    .din1(G90_n_spl_10),
    .din2(G101_n_spl_101)
  );


  LA
  g_g1334_p
  (
    .dout(g1334_p),
    .din1(G90_n_spl_10),
    .din2(G100_p_spl_101)
  );


  FA
  g_g1334_n
  (
    .dout(g1334_n),
    .din1(G90_p_spl_10),
    .din2(G100_n_spl_101)
  );


  LA
  g_g1335_p
  (
    .dout(g1335_p),
    .din1(g1333_n),
    .din2(g1334_n)
  );


  FA
  g_g1335_n
  (
    .dout(g1335_n),
    .din1(g1333_p),
    .din2(g1334_p)
  );


  LA
  g_g1336_p
  (
    .dout(g1336_p),
    .din1(G143_p_spl_1),
    .din2(g1335_n)
  );


  FA
  g_g1336_n
  (
    .dout(g1336_n),
    .din1(G143_n_spl_1),
    .din2(g1335_p)
  );


  LA
  g_g1337_p
  (
    .dout(g1337_p),
    .din1(G90_p_spl_11),
    .din2(G102_n_spl_100)
  );


  FA
  g_g1337_n
  (
    .dout(g1337_n),
    .din1(G90_n_spl_11),
    .din2(G102_p_spl_100)
  );


  LA
  g_g1338_p
  (
    .dout(g1338_p),
    .din1(G90_n_spl_11),
    .din2(G98_n_spl_101)
  );


  FA
  g_g1338_n
  (
    .dout(g1338_n),
    .din1(G90_p_spl_11),
    .din2(G98_p_spl_101)
  );


  LA
  g_g1339_p
  (
    .dout(g1339_p),
    .din1(g1337_n),
    .din2(g1338_n)
  );


  FA
  g_g1339_n
  (
    .dout(g1339_n),
    .din1(g1337_p),
    .din2(g1338_p)
  );


  LA
  g_g1340_p
  (
    .dout(g1340_p),
    .din1(G143_n_spl_1),
    .din2(g1339_n)
  );


  FA
  g_g1340_n
  (
    .dout(g1340_n),
    .din1(G143_p_spl_1),
    .din2(g1339_p)
  );


  LA
  g_g1341_p
  (
    .dout(g1341_p),
    .din1(g1336_n),
    .din2(g1340_n)
  );


  FA
  g_g1341_n
  (
    .dout(g1341_n),
    .din1(g1336_p),
    .din2(g1340_p)
  );


  LA
  g_g1342_p
  (
    .dout(g1342_p),
    .din1(g317_n_spl_1),
    .din2(g1341_n_spl_)
  );


  FA
  g_g1342_n
  (
    .dout(g1342_n),
    .din1(g317_p_spl_),
    .din2(g1341_p_spl_)
  );


  LA
  g_g1343_p
  (
    .dout(g1343_p),
    .din1(g317_p_spl_),
    .din2(g1341_p_spl_)
  );


  FA
  g_g1343_n
  (
    .dout(g1343_n),
    .din1(g317_n_spl_1),
    .din2(g1341_n_spl_)
  );


  LA
  g_g1344_p
  (
    .dout(g1344_p),
    .din1(g1342_n),
    .din2(g1343_n)
  );


  FA
  g_g1344_n
  (
    .dout(g1344_n),
    .din1(g1342_p),
    .din2(g1343_p)
  );


  LA
  g_g1345_p
  (
    .dout(g1345_p),
    .din1(g1332_n_spl_),
    .din2(g1344_p_spl_)
  );


  FA
  g_g1345_n
  (
    .dout(g1345_n),
    .din1(g1332_p_spl_),
    .din2(g1344_n_spl_)
  );


  LA
  g_g1346_p
  (
    .dout(g1346_p),
    .din1(g1332_p_spl_),
    .din2(g1344_n_spl_)
  );


  FA
  g_g1346_n
  (
    .dout(g1346_n),
    .din1(g1332_n_spl_),
    .din2(g1344_p_spl_)
  );


  LA
  g_g1347_p
  (
    .dout(g1347_p),
    .din1(g1345_n),
    .din2(g1346_n)
  );


  FA
  g_g1347_n
  (
    .dout(g1347_n),
    .din1(g1345_p),
    .din2(g1346_p)
  );


  LA
  g_g1348_p
  (
    .dout(g1348_p),
    .din1(G101_p_spl_101),
    .din2(G107_p_spl_10)
  );


  FA
  g_g1348_n
  (
    .dout(g1348_n),
    .din1(G101_n_spl_101),
    .din2(G107_n_spl_10)
  );


  LA
  g_g1349_p
  (
    .dout(g1349_p),
    .din1(G100_p_spl_101),
    .din2(G107_n_spl_10)
  );


  FA
  g_g1349_n
  (
    .dout(g1349_n),
    .din1(G100_n_spl_101),
    .din2(G107_p_spl_10)
  );


  LA
  g_g1350_p
  (
    .dout(g1350_p),
    .din1(g1348_n),
    .din2(g1349_n)
  );


  FA
  g_g1350_n
  (
    .dout(g1350_n),
    .din1(g1348_p),
    .din2(g1349_p)
  );


  LA
  g_g1351_p
  (
    .dout(g1351_p),
    .din1(G139_p_spl_1),
    .din2(g1350_n)
  );


  FA
  g_g1351_n
  (
    .dout(g1351_n),
    .din1(G139_n_spl_1),
    .din2(g1350_p)
  );


  LA
  g_g1352_p
  (
    .dout(g1352_p),
    .din1(G102_n_spl_101),
    .din2(G107_p_spl_11)
  );


  FA
  g_g1352_n
  (
    .dout(g1352_n),
    .din1(G102_p_spl_101),
    .din2(G107_n_spl_11)
  );


  LA
  g_g1353_p
  (
    .dout(g1353_p),
    .din1(G98_n_spl_101),
    .din2(G107_n_spl_11)
  );


  FA
  g_g1353_n
  (
    .dout(g1353_n),
    .din1(G98_p_spl_101),
    .din2(G107_p_spl_11)
  );


  LA
  g_g1354_p
  (
    .dout(g1354_p),
    .din1(g1352_n),
    .din2(g1353_n)
  );


  FA
  g_g1354_n
  (
    .dout(g1354_n),
    .din1(g1352_p),
    .din2(g1353_p)
  );


  LA
  g_g1355_p
  (
    .dout(g1355_p),
    .din1(G139_n_spl_1),
    .din2(g1354_n)
  );


  FA
  g_g1355_n
  (
    .dout(g1355_n),
    .din1(G139_p_spl_1),
    .din2(g1354_p)
  );


  LA
  g_g1356_p
  (
    .dout(g1356_p),
    .din1(g1351_n),
    .din2(g1355_n)
  );


  FA
  g_g1356_n
  (
    .dout(g1356_n),
    .din1(g1351_p),
    .din2(g1355_p)
  );


  LA
  g_g1357_p
  (
    .dout(g1357_p),
    .din1(G101_p_spl_110),
    .din2(G105_p_spl_10)
  );


  FA
  g_g1357_n
  (
    .dout(g1357_n),
    .din1(G101_n_spl_110),
    .din2(G105_n_spl_10)
  );


  LA
  g_g1358_p
  (
    .dout(g1358_p),
    .din1(G100_p_spl_110),
    .din2(G105_n_spl_10)
  );


  FA
  g_g1358_n
  (
    .dout(g1358_n),
    .din1(G100_n_spl_110),
    .din2(G105_p_spl_10)
  );


  LA
  g_g1359_p
  (
    .dout(g1359_p),
    .din1(g1357_n),
    .din2(g1358_n)
  );


  FA
  g_g1359_n
  (
    .dout(g1359_n),
    .din1(g1357_p),
    .din2(g1358_p)
  );


  LA
  g_g1360_p
  (
    .dout(g1360_p),
    .din1(G138_p_spl_1),
    .din2(g1359_n)
  );


  FA
  g_g1360_n
  (
    .dout(g1360_n),
    .din1(G138_n_spl_1),
    .din2(g1359_p)
  );


  LA
  g_g1361_p
  (
    .dout(g1361_p),
    .din1(G102_n_spl_101),
    .din2(G105_p_spl_11)
  );


  FA
  g_g1361_n
  (
    .dout(g1361_n),
    .din1(G102_p_spl_101),
    .din2(G105_n_spl_11)
  );


  LA
  g_g1362_p
  (
    .dout(g1362_p),
    .din1(G98_n_spl_110),
    .din2(G105_n_spl_11)
  );


  FA
  g_g1362_n
  (
    .dout(g1362_n),
    .din1(G98_p_spl_110),
    .din2(G105_p_spl_11)
  );


  LA
  g_g1363_p
  (
    .dout(g1363_p),
    .din1(g1361_n),
    .din2(g1362_n)
  );


  FA
  g_g1363_n
  (
    .dout(g1363_n),
    .din1(g1361_p),
    .din2(g1362_p)
  );


  LA
  g_g1364_p
  (
    .dout(g1364_p),
    .din1(G138_n_spl_1),
    .din2(g1363_n)
  );


  FA
  g_g1364_n
  (
    .dout(g1364_n),
    .din1(G138_p_spl_1),
    .din2(g1363_p)
  );


  LA
  g_g1365_p
  (
    .dout(g1365_p),
    .din1(g1360_n),
    .din2(g1364_n)
  );


  FA
  g_g1365_n
  (
    .dout(g1365_n),
    .din1(g1360_p),
    .din2(g1364_p)
  );


  LA
  g_g1366_p
  (
    .dout(g1366_p),
    .din1(g1356_n_spl_),
    .din2(g1365_p_spl_)
  );


  FA
  g_g1366_n
  (
    .dout(g1366_n),
    .din1(g1356_p_spl_),
    .din2(g1365_n_spl_)
  );


  LA
  g_g1367_p
  (
    .dout(g1367_p),
    .din1(g1356_p_spl_),
    .din2(g1365_n_spl_)
  );


  FA
  g_g1367_n
  (
    .dout(g1367_n),
    .din1(g1356_n_spl_),
    .din2(g1365_p_spl_)
  );


  LA
  g_g1368_p
  (
    .dout(g1368_p),
    .din1(g1366_n),
    .din2(g1367_n)
  );


  FA
  g_g1368_n
  (
    .dout(g1368_n),
    .din1(g1366_p),
    .din2(g1367_p)
  );


  LA
  g_g1369_p
  (
    .dout(g1369_p),
    .din1(G101_p_spl_110),
    .din2(G103_p_spl_10)
  );


  FA
  g_g1369_n
  (
    .dout(g1369_n),
    .din1(G101_n_spl_110),
    .din2(G103_n_spl_10)
  );


  LA
  g_g1370_p
  (
    .dout(g1370_p),
    .din1(G100_p_spl_110),
    .din2(G103_n_spl_10)
  );


  FA
  g_g1370_n
  (
    .dout(g1370_n),
    .din1(G100_n_spl_110),
    .din2(G103_p_spl_10)
  );


  LA
  g_g1371_p
  (
    .dout(g1371_p),
    .din1(g1369_n),
    .din2(g1370_n)
  );


  FA
  g_g1371_n
  (
    .dout(g1371_n),
    .din1(g1369_p),
    .din2(g1370_p)
  );


  LA
  g_g1372_p
  (
    .dout(g1372_p),
    .din1(G137_p_spl_1),
    .din2(g1371_n)
  );


  FA
  g_g1372_n
  (
    .dout(g1372_n),
    .din1(G137_n_spl_1),
    .din2(g1371_p)
  );


  LA
  g_g1373_p
  (
    .dout(g1373_p),
    .din1(G102_n_spl_110),
    .din2(G103_p_spl_11)
  );


  FA
  g_g1373_n
  (
    .dout(g1373_n),
    .din1(G102_p_spl_110),
    .din2(G103_n_spl_11)
  );


  LA
  g_g1374_p
  (
    .dout(g1374_p),
    .din1(G98_n_spl_110),
    .din2(G103_n_spl_11)
  );


  FA
  g_g1374_n
  (
    .dout(g1374_n),
    .din1(G98_p_spl_110),
    .din2(G103_p_spl_11)
  );


  LA
  g_g1375_p
  (
    .dout(g1375_p),
    .din1(g1373_n),
    .din2(g1374_n)
  );


  FA
  g_g1375_n
  (
    .dout(g1375_n),
    .din1(g1373_p),
    .din2(g1374_p)
  );


  LA
  g_g1376_p
  (
    .dout(g1376_p),
    .din1(G137_n_spl_1),
    .din2(g1375_n)
  );


  FA
  g_g1376_n
  (
    .dout(g1376_n),
    .din1(G137_p_spl_1),
    .din2(g1375_p)
  );


  LA
  g_g1377_p
  (
    .dout(g1377_p),
    .din1(g1372_n),
    .din2(g1376_n)
  );


  FA
  g_g1377_n
  (
    .dout(g1377_n),
    .din1(g1372_p),
    .din2(g1376_p)
  );


  LA
  g_g1378_p
  (
    .dout(g1378_p),
    .din1(G96_p_spl_10),
    .din2(G101_p_spl_111)
  );


  FA
  g_g1378_n
  (
    .dout(g1378_n),
    .din1(G96_n_spl_10),
    .din2(G101_n_spl_111)
  );


  LA
  g_g1379_p
  (
    .dout(g1379_p),
    .din1(G96_n_spl_10),
    .din2(G100_p_spl_111)
  );


  FA
  g_g1379_n
  (
    .dout(g1379_n),
    .din1(G96_p_spl_10),
    .din2(G100_n_spl_111)
  );


  LA
  g_g1380_p
  (
    .dout(g1380_p),
    .din1(g1378_n),
    .din2(g1379_n)
  );


  FA
  g_g1380_n
  (
    .dout(g1380_n),
    .din1(g1378_p),
    .din2(g1379_p)
  );


  LA
  g_g1381_p
  (
    .dout(g1381_p),
    .din1(G141_p_spl_1),
    .din2(g1380_n)
  );


  FA
  g_g1381_n
  (
    .dout(g1381_n),
    .din1(G141_n_spl_1),
    .din2(g1380_p)
  );


  LA
  g_g1382_p
  (
    .dout(g1382_p),
    .din1(G96_p_spl_11),
    .din2(G102_n_spl_110)
  );


  FA
  g_g1382_n
  (
    .dout(g1382_n),
    .din1(G96_n_spl_11),
    .din2(G102_p_spl_110)
  );


  LA
  g_g1383_p
  (
    .dout(g1383_p),
    .din1(G96_n_spl_11),
    .din2(G98_n_spl_111)
  );


  FA
  g_g1383_n
  (
    .dout(g1383_n),
    .din1(G96_p_spl_11),
    .din2(G98_p_spl_111)
  );


  LA
  g_g1384_p
  (
    .dout(g1384_p),
    .din1(g1382_n),
    .din2(g1383_n)
  );


  FA
  g_g1384_n
  (
    .dout(g1384_n),
    .din1(g1382_p),
    .din2(g1383_p)
  );


  LA
  g_g1385_p
  (
    .dout(g1385_p),
    .din1(G141_n_spl_1),
    .din2(g1384_n)
  );


  FA
  g_g1385_n
  (
    .dout(g1385_n),
    .din1(G141_p_spl_1),
    .din2(g1384_p)
  );


  LA
  g_g1386_p
  (
    .dout(g1386_p),
    .din1(g1381_n),
    .din2(g1385_n)
  );


  FA
  g_g1386_n
  (
    .dout(g1386_n),
    .din1(g1381_p),
    .din2(g1385_p)
  );


  LA
  g_g1387_p
  (
    .dout(g1387_p),
    .din1(g1377_n_spl_),
    .din2(g1386_p_spl_)
  );


  FA
  g_g1387_n
  (
    .dout(g1387_n),
    .din1(g1377_p_spl_),
    .din2(g1386_n_spl_)
  );


  LA
  g_g1388_p
  (
    .dout(g1388_p),
    .din1(g1377_p_spl_),
    .din2(g1386_n_spl_)
  );


  FA
  g_g1388_n
  (
    .dout(g1388_n),
    .din1(g1377_n_spl_),
    .din2(g1386_p_spl_)
  );


  LA
  g_g1389_p
  (
    .dout(g1389_p),
    .din1(g1387_n),
    .din2(g1388_n)
  );


  FA
  g_g1389_n
  (
    .dout(g1389_n),
    .din1(g1387_p),
    .din2(g1388_p)
  );


  LA
  g_g1390_p
  (
    .dout(g1390_p),
    .din1(G101_p_spl_111),
    .din2(G109_p_spl_10)
  );


  FA
  g_g1390_n
  (
    .dout(g1390_n),
    .din1(G101_n_spl_111),
    .din2(G109_n_spl_10)
  );


  LA
  g_g1391_p
  (
    .dout(g1391_p),
    .din1(G100_p_spl_111),
    .din2(G109_n_spl_10)
  );


  FA
  g_g1391_n
  (
    .dout(g1391_n),
    .din1(G100_n_spl_111),
    .din2(G109_p_spl_10)
  );


  LA
  g_g1392_p
  (
    .dout(g1392_p),
    .din1(g1390_n),
    .din2(g1391_n)
  );


  FA
  g_g1392_n
  (
    .dout(g1392_n),
    .din1(g1390_p),
    .din2(g1391_p)
  );


  LA
  g_g1393_p
  (
    .dout(g1393_p),
    .din1(G135_p_spl_1),
    .din2(g1392_n)
  );


  FA
  g_g1393_n
  (
    .dout(g1393_n),
    .din1(G135_n_spl_1),
    .din2(g1392_p)
  );


  LA
  g_g1394_p
  (
    .dout(g1394_p),
    .din1(G102_n_spl_11),
    .din2(G109_p_spl_11)
  );


  FA
  g_g1394_n
  (
    .dout(g1394_n),
    .din1(G102_p_spl_11),
    .din2(G109_n_spl_11)
  );


  LA
  g_g1395_p
  (
    .dout(g1395_p),
    .din1(G98_n_spl_111),
    .din2(G109_n_spl_11)
  );


  FA
  g_g1395_n
  (
    .dout(g1395_n),
    .din1(G98_p_spl_111),
    .din2(G109_p_spl_11)
  );


  LA
  g_g1396_p
  (
    .dout(g1396_p),
    .din1(g1394_n),
    .din2(g1395_n)
  );


  FA
  g_g1396_n
  (
    .dout(g1396_n),
    .din1(g1394_p),
    .din2(g1395_p)
  );


  LA
  g_g1397_p
  (
    .dout(g1397_p),
    .din1(G135_n_spl_1),
    .din2(g1396_n)
  );


  FA
  g_g1397_n
  (
    .dout(g1397_n),
    .din1(G135_p_spl_1),
    .din2(g1396_p)
  );


  LA
  g_g1398_p
  (
    .dout(g1398_p),
    .din1(g1393_n),
    .din2(g1397_n)
  );


  FA
  g_g1398_n
  (
    .dout(g1398_n),
    .din1(g1393_p),
    .din2(g1397_p)
  );


  LA
  g_g1399_p
  (
    .dout(g1399_p),
    .din1(g1389_p_spl_),
    .din2(g1398_n_spl_)
  );


  FA
  g_g1399_n
  (
    .dout(g1399_n),
    .din1(g1389_n_spl_),
    .din2(g1398_p_spl_)
  );


  LA
  g_g1400_p
  (
    .dout(g1400_p),
    .din1(g1389_n_spl_),
    .din2(g1398_p_spl_)
  );


  FA
  g_g1400_n
  (
    .dout(g1400_n),
    .din1(g1389_p_spl_),
    .din2(g1398_n_spl_)
  );


  LA
  g_g1401_p
  (
    .dout(g1401_p),
    .din1(g1399_n),
    .din2(g1400_n)
  );


  FA
  g_g1401_n
  (
    .dout(g1401_n),
    .din1(g1399_p),
    .din2(g1400_p)
  );


  LA
  g_g1402_p
  (
    .dout(g1402_p),
    .din1(g1368_p_spl_),
    .din2(g1401_n_spl_)
  );


  FA
  g_g1402_n
  (
    .dout(g1402_n),
    .din1(g1368_n_spl_),
    .din2(g1401_p_spl_)
  );


  LA
  g_g1403_p
  (
    .dout(g1403_p),
    .din1(g1368_n_spl_),
    .din2(g1401_p_spl_)
  );


  FA
  g_g1403_n
  (
    .dout(g1403_n),
    .din1(g1368_p_spl_),
    .din2(g1401_n_spl_)
  );


  LA
  g_g1404_p
  (
    .dout(g1404_p),
    .din1(g1402_n),
    .din2(g1403_n)
  );


  FA
  g_g1404_n
  (
    .dout(g1404_n),
    .din1(g1402_p),
    .din2(g1403_p)
  );


  FA
  g_g1405_n
  (
    .dout(g1405_n),
    .din1(g1347_p),
    .din2(g1404_n)
  );


  FA
  g_g1406_n
  (
    .dout(g1406_n),
    .din1(g1347_n),
    .din2(g1404_p)
  );


  LA
  g_g1407_p
  (
    .dout(g1407_p),
    .din1(g1405_n),
    .din2(g1406_n)
  );


  FA
  g_g1408_n
  (
    .dout(g1408_n),
    .din1(G176_n_spl_111),
    .din2(g1407_p)
  );


  LA
  g_g1409_p
  (
    .dout(g1409_p),
    .din1(g389_n_spl_),
    .din2(g546_p_spl_1)
  );


  FA
  g_g1409_n
  (
    .dout(g1409_n),
    .din1(g389_p_spl_),
    .din2(g546_n_spl_0)
  );


  LA
  g_g1410_p
  (
    .dout(g1410_p),
    .din1(g374_p_spl_1),
    .din2(g544_n_spl_1)
  );


  FA
  g_g1410_n
  (
    .dout(g1410_n),
    .din1(g374_n_spl_1),
    .din2(g544_p_spl_1)
  );


  LA
  g_g1411_p
  (
    .dout(g1411_p),
    .din1(g374_n_spl_1),
    .din2(g380_p_spl_)
  );


  FA
  g_g1411_n
  (
    .dout(g1411_n),
    .din1(g374_p_spl_1),
    .din2(g380_n_spl_)
  );


  LA
  g_g1412_p
  (
    .dout(g1412_p),
    .din1(g1410_n),
    .din2(g1411_n)
  );


  FA
  g_g1412_n
  (
    .dout(g1412_n),
    .din1(g1410_p),
    .din2(g1411_p)
  );


  LA
  g_g1413_p
  (
    .dout(g1413_p),
    .din1(g1409_n_spl_),
    .din2(g1412_n_spl_)
  );


  FA
  g_g1413_n
  (
    .dout(g1413_n),
    .din1(g1409_p_spl_),
    .din2(g1412_p_spl_)
  );


  LA
  g_g1414_p
  (
    .dout(g1414_p),
    .din1(g1409_p_spl_),
    .din2(g1412_p_spl_)
  );


  FA
  g_g1414_n
  (
    .dout(g1414_n),
    .din1(g1409_n_spl_),
    .din2(g1412_n_spl_)
  );


  LA
  g_g1415_p
  (
    .dout(g1415_p),
    .din1(g1413_n),
    .din2(g1414_n)
  );


  FA
  g_g1415_n
  (
    .dout(g1415_n),
    .din1(g1413_p),
    .din2(g1414_p)
  );


  LA
  g_g1416_p
  (
    .dout(g1416_p),
    .din1(g375_n_spl_0),
    .din2(g1415_p_spl_)
  );


  FA
  g_g1416_n
  (
    .dout(g1416_n),
    .din1(g375_p_spl_0),
    .din2(g1415_n_spl_)
  );


  LA
  g_g1417_p
  (
    .dout(g1417_p),
    .din1(g544_p_spl_1),
    .din2(g546_p_spl_1)
  );


  FA
  g_g1417_n
  (
    .dout(g1417_n),
    .din1(g544_n_spl_1),
    .din2(g546_n_spl_)
  );


  LA
  g_g1418_p
  (
    .dout(g1418_p),
    .din1(g545_n_spl_),
    .din2(g1417_n)
  );


  FA
  g_g1418_n
  (
    .dout(g1418_n),
    .din1(g545_p_spl_),
    .din2(g1417_p)
  );


  LA
  g_g1419_p
  (
    .dout(g1419_p),
    .din1(g375_p_spl_1),
    .din2(g1418_n)
  );


  FA
  g_g1419_n
  (
    .dout(g1419_n),
    .din1(g375_n_spl_1),
    .din2(g1418_p)
  );


  LA
  g_g1420_p
  (
    .dout(g1420_p),
    .din1(g1416_n_spl_),
    .din2(g1419_n)
  );


  FA
  g_g1420_n
  (
    .dout(g1420_n),
    .din1(g1416_p_spl_),
    .din2(g1419_p)
  );


  LA
  g_g1421_p
  (
    .dout(g1421_p),
    .din1(g381_n_spl_01),
    .din2(g1420_p_spl_)
  );


  FA
  g_g1421_n
  (
    .dout(g1421_n),
    .din1(g381_p_spl_01),
    .din2(g1420_n_spl_)
  );


  LA
  g_g1422_p
  (
    .dout(g1422_p),
    .din1(g381_p_spl_10),
    .din2(g1420_n_spl_)
  );


  FA
  g_g1422_n
  (
    .dout(g1422_n),
    .din1(g381_n_spl_10),
    .din2(g1420_p_spl_)
  );


  LA
  g_g1423_p
  (
    .dout(g1423_p),
    .din1(g1421_n),
    .din2(g1422_n)
  );


  FA
  g_g1423_n
  (
    .dout(g1423_n),
    .din1(g1421_p),
    .din2(g1422_p)
  );


  LA
  g_g1424_p
  (
    .dout(g1424_p),
    .din1(g395_n_spl_01),
    .din2(g1423_p_spl_)
  );


  FA
  g_g1424_n
  (
    .dout(g1424_n),
    .din1(g395_p_spl_00),
    .din2(g1423_n_spl_)
  );


  LA
  g_g1425_p
  (
    .dout(g1425_p),
    .din1(g395_p_spl_0),
    .din2(g1423_n_spl_)
  );


  FA
  g_g1425_n
  (
    .dout(g1425_n),
    .din1(g395_n_spl_10),
    .din2(g1423_p_spl_)
  );


  LA
  g_g1426_p
  (
    .dout(g1426_p),
    .din1(g1424_n),
    .din2(g1425_n)
  );


  FA
  g_g1426_n
  (
    .dout(g1426_n),
    .din1(g1424_p),
    .din2(g1425_p)
  );


  LA
  g_g1427_p
  (
    .dout(g1427_p),
    .din1(g388_n_spl_01),
    .din2(g1426_p_spl_)
  );


  FA
  g_g1427_n
  (
    .dout(g1427_n),
    .din1(g388_p_spl_01),
    .din2(g1426_n_spl_)
  );


  LA
  g_g1428_p
  (
    .dout(g1428_p),
    .din1(g388_p_spl_01),
    .din2(g1426_n_spl_)
  );


  FA
  g_g1428_n
  (
    .dout(g1428_n),
    .din1(g388_n_spl_01),
    .din2(g1426_p_spl_)
  );


  LA
  g_g1429_p
  (
    .dout(g1429_p),
    .din1(g1427_n),
    .din2(g1428_n)
  );


  FA
  g_g1429_n
  (
    .dout(g1429_n),
    .din1(g1427_p),
    .din2(g1428_p)
  );


  LA
  g_g1430_p
  (
    .dout(g1430_p),
    .din1(g541_p_spl_0),
    .din2(g1429_n)
  );


  FA
  g_g1430_n
  (
    .dout(g1430_n),
    .din1(g541_n_spl_0),
    .din2(g1429_p)
  );


  LA
  g_g1431_p
  (
    .dout(g1431_p),
    .din1(g375_p_spl_1),
    .din2(g1415_n_spl_)
  );


  FA
  g_g1431_n
  (
    .dout(g1431_n),
    .din1(g375_n_spl_1),
    .din2(g1415_p_spl_)
  );


  LA
  g_g1432_p
  (
    .dout(g1432_p),
    .din1(g1416_n_spl_),
    .din2(g1431_n)
  );


  FA
  g_g1432_n
  (
    .dout(g1432_n),
    .din1(g1416_p_spl_),
    .din2(g1431_p)
  );


  LA
  g_g1433_p
  (
    .dout(g1433_p),
    .din1(g381_n_spl_10),
    .din2(g1432_p_spl_)
  );


  FA
  g_g1433_n
  (
    .dout(g1433_n),
    .din1(g381_p_spl_10),
    .din2(g1432_n_spl_)
  );


  LA
  g_g1434_p
  (
    .dout(g1434_p),
    .din1(g381_p_spl_1),
    .din2(g1432_n_spl_)
  );


  FA
  g_g1434_n
  (
    .dout(g1434_n),
    .din1(g381_n_spl_1),
    .din2(g1432_p_spl_)
  );


  LA
  g_g1435_p
  (
    .dout(g1435_p),
    .din1(g1433_n),
    .din2(g1434_n)
  );


  FA
  g_g1435_n
  (
    .dout(g1435_n),
    .din1(g1433_p),
    .din2(g1434_p)
  );


  LA
  g_g1436_p
  (
    .dout(g1436_p),
    .din1(g395_n_spl_10),
    .din2(g1435_p_spl_)
  );


  FA
  g_g1436_n
  (
    .dout(g1436_n),
    .din1(g395_p_spl_1),
    .din2(g1435_n_spl_)
  );


  LA
  g_g1437_p
  (
    .dout(g1437_p),
    .din1(g395_p_spl_1),
    .din2(g1435_n_spl_)
  );


  FA
  g_g1437_n
  (
    .dout(g1437_n),
    .din1(g395_n_spl_1),
    .din2(g1435_p_spl_)
  );


  LA
  g_g1438_p
  (
    .dout(g1438_p),
    .din1(g1436_n),
    .din2(g1437_n)
  );


  FA
  g_g1438_n
  (
    .dout(g1438_n),
    .din1(g1436_p),
    .din2(g1437_p)
  );


  LA
  g_g1439_p
  (
    .dout(g1439_p),
    .din1(g388_n_spl_1),
    .din2(g1438_p_spl_)
  );


  FA
  g_g1439_n
  (
    .dout(g1439_n),
    .din1(g388_p_spl_1),
    .din2(g1438_n_spl_)
  );


  LA
  g_g1440_p
  (
    .dout(g1440_p),
    .din1(g388_p_spl_1),
    .din2(g1438_n_spl_)
  );


  FA
  g_g1440_n
  (
    .dout(g1440_n),
    .din1(g388_n_spl_1),
    .din2(g1438_p_spl_)
  );


  LA
  g_g1441_p
  (
    .dout(g1441_p),
    .din1(g1439_n),
    .din2(g1440_n)
  );


  FA
  g_g1441_n
  (
    .dout(g1441_n),
    .din1(g1439_p),
    .din2(g1440_p)
  );


  LA
  g_g1442_p
  (
    .dout(g1442_p),
    .din1(g541_n_spl_1),
    .din2(g1441_n_spl_)
  );


  FA
  g_g1442_n
  (
    .dout(g1442_n),
    .din1(g541_p_spl_1),
    .din2(g1441_p_spl_)
  );


  LA
  g_g1443_p
  (
    .dout(g1443_p),
    .din1(g1430_n_spl_),
    .din2(g1442_n)
  );


  FA
  g_g1443_n
  (
    .dout(g1443_n),
    .din1(g1430_p_spl_),
    .din2(g1442_p)
  );


  LA
  g_g1444_p
  (
    .dout(g1444_p),
    .din1(G157_n_spl_0),
    .din2(g1443_n)
  );


  FA
  g_g1444_n
  (
    .dout(g1444_n),
    .din1(G157_p_spl_0),
    .din2(g1443_p)
  );


  LA
  g_g1445_p
  (
    .dout(g1445_p),
    .din1(g430_n_spl_1),
    .din2(g541_p_spl_1)
  );


  FA
  g_g1445_n
  (
    .dout(g1445_n),
    .din1(g430_p_spl_0),
    .din2(g541_n_spl_1)
  );


  LA
  g_g1446_p
  (
    .dout(g1446_p),
    .din1(g1441_n_spl_),
    .din2(g1445_n)
  );


  FA
  g_g1446_n
  (
    .dout(g1446_n),
    .din1(g1441_p_spl_),
    .din2(g1445_p)
  );


  LA
  g_g1447_p
  (
    .dout(g1447_p),
    .din1(g430_n_spl_1),
    .din2(g1430_p_spl_)
  );


  FA
  g_g1447_n
  (
    .dout(g1447_n),
    .din1(g430_p_spl_),
    .din2(g1430_n_spl_)
  );


  LA
  g_g1448_p
  (
    .dout(g1448_p),
    .din1(g1446_n),
    .din2(g1447_n)
  );


  FA
  g_g1448_n
  (
    .dout(g1448_n),
    .din1(g1446_p),
    .din2(g1447_p)
  );


  LA
  g_g1449_p
  (
    .dout(g1449_p),
    .din1(G157_p_spl_0),
    .din2(g1448_n)
  );


  FA
  g_g1449_n
  (
    .dout(g1449_n),
    .din1(G157_n_spl_0),
    .din2(g1448_p)
  );


  LA
  g_g1450_p
  (
    .dout(g1450_p),
    .din1(g1444_n),
    .din2(g1449_n)
  );


  FA
  g_g1450_n
  (
    .dout(g1450_n),
    .din1(g1444_p),
    .din2(g1449_p)
  );


  LA
  g_g1451_p
  (
    .dout(g1451_p),
    .din1(g400_p_spl_1),
    .din2(g537_n_spl_0)
  );


  FA
  g_g1451_n
  (
    .dout(g1451_n),
    .din1(g400_n_spl_1),
    .din2(g537_p_spl_0)
  );


  LA
  g_g1452_p
  (
    .dout(g1452_p),
    .din1(g400_n_spl_1),
    .din2(g537_p_spl_1)
  );


  FA
  g_g1452_n
  (
    .dout(g1452_n),
    .din1(g400_p_spl_1),
    .din2(g537_n_spl_1)
  );


  LA
  g_g1453_p
  (
    .dout(g1453_p),
    .din1(g1451_n),
    .din2(g1452_n)
  );


  FA
  g_g1453_n
  (
    .dout(g1453_n),
    .din1(g1451_p),
    .din2(g1452_p)
  );


  LA
  g_g1454_p
  (
    .dout(g1454_p),
    .din1(g535_p_spl_0),
    .din2(g1453_n_spl_)
  );


  FA
  g_g1454_n
  (
    .dout(g1454_n),
    .din1(g535_n_spl_0),
    .din2(g1453_p_spl_)
  );


  LA
  g_g1455_p
  (
    .dout(g1455_p),
    .din1(g535_n_spl_1),
    .din2(g1453_p_spl_)
  );


  FA
  g_g1455_n
  (
    .dout(g1455_n),
    .din1(g535_p_spl_1),
    .din2(g1453_n_spl_)
  );


  LA
  g_g1456_p
  (
    .dout(g1456_p),
    .din1(g1454_n),
    .din2(g1455_n)
  );


  FA
  g_g1456_n
  (
    .dout(g1456_n),
    .din1(g1454_p),
    .din2(g1455_p)
  );


  LA
  g_g1457_p
  (
    .dout(g1457_p),
    .din1(g402_n_spl_),
    .din2(g408_n_spl_1)
  );


  FA
  g_g1457_n
  (
    .dout(g1457_n),
    .din1(g402_p_spl_1),
    .din2(g408_p_spl_1)
  );


  LA
  g_g1458_p
  (
    .dout(g1458_p),
    .din1(g409_n_spl_0),
    .din2(g1457_n)
  );


  FA
  g_g1458_n
  (
    .dout(g1458_n),
    .din1(g409_p_spl_0),
    .din2(g1457_p)
  );


  LA
  g_g1459_p
  (
    .dout(g1459_p),
    .din1(g539_n_spl_0),
    .din2(g1458_n_spl_0)
  );


  FA
  g_g1459_n
  (
    .dout(g1459_n),
    .din1(g539_p_spl_0),
    .din2(g1458_p_spl_0)
  );


  LA
  g_g1460_p
  (
    .dout(g1460_p),
    .din1(g539_p_spl_1),
    .din2(g1458_p_spl_0)
  );


  FA
  g_g1460_n
  (
    .dout(g1460_n),
    .din1(g539_n_spl_1),
    .din2(g1458_n_spl_0)
  );


  LA
  g_g1461_p
  (
    .dout(g1461_p),
    .din1(g1459_n),
    .din2(g1460_n)
  );


  FA
  g_g1461_n
  (
    .dout(g1461_n),
    .din1(g1459_p),
    .din2(g1460_p)
  );


  LA
  g_g1462_p
  (
    .dout(g1462_p),
    .din1(g1456_n_spl_),
    .din2(g1461_p_spl_)
  );


  FA
  g_g1462_n
  (
    .dout(g1462_n),
    .din1(g1456_p_spl_),
    .din2(g1461_n_spl_)
  );


  LA
  g_g1463_p
  (
    .dout(g1463_p),
    .din1(g1456_p_spl_),
    .din2(g1461_n_spl_)
  );


  FA
  g_g1463_n
  (
    .dout(g1463_n),
    .din1(g1456_n_spl_),
    .din2(g1461_p_spl_)
  );


  LA
  g_g1464_p
  (
    .dout(g1464_p),
    .din1(g1462_n),
    .din2(g1463_n)
  );


  FA
  g_g1464_n
  (
    .dout(g1464_n),
    .din1(g1462_p),
    .din2(g1463_p)
  );


  LA
  g_g1465_p
  (
    .dout(g1465_p),
    .din1(g429_n_spl_01),
    .din2(g1464_n_spl_)
  );


  FA
  g_g1465_n
  (
    .dout(g1465_n),
    .din1(g429_p_spl_01),
    .din2(g1464_p_spl_)
  );


  LA
  g_g1466_p
  (
    .dout(g1466_p),
    .din1(g429_p_spl_10),
    .din2(g1464_p_spl_)
  );


  FA
  g_g1466_n
  (
    .dout(g1466_n),
    .din1(g429_n_spl_10),
    .din2(g1464_n_spl_)
  );


  LA
  g_g1467_p
  (
    .dout(g1467_p),
    .din1(g1465_n),
    .din2(g1466_n)
  );


  FA
  g_g1467_n
  (
    .dout(g1467_n),
    .din1(g1465_p),
    .din2(g1466_p)
  );


  LA
  g_g1468_p
  (
    .dout(g1468_p),
    .din1(G157_n_spl_1),
    .din2(g1467_p)
  );


  FA
  g_g1468_n
  (
    .dout(g1468_n),
    .din1(G157_p_spl_1),
    .din2(g1467_n)
  );


  LA
  g_g1469_p
  (
    .dout(g1469_p),
    .din1(g423_n_spl_),
    .din2(g539_p_spl_1)
  );


  FA
  g_g1469_n
  (
    .dout(g1469_n),
    .din1(g423_p_spl_),
    .din2(g539_n_spl_1)
  );


  LA
  g_g1470_p
  (
    .dout(g1470_p),
    .din1(g409_n_spl_),
    .din2(g535_p_spl_1)
  );


  FA
  g_g1470_n
  (
    .dout(g1470_n),
    .din1(g409_p_spl_),
    .din2(g535_n_spl_1)
  );


  LA
  g_g1471_p
  (
    .dout(g1471_p),
    .din1(g416_n_spl_),
    .din2(g537_p_spl_1)
  );


  FA
  g_g1471_n
  (
    .dout(g1471_n),
    .din1(g416_p_spl_),
    .din2(g537_n_spl_1)
  );


  LA
  g_g1472_p
  (
    .dout(g1472_p),
    .din1(g401_n_spl_0),
    .din2(g1471_n_spl_)
  );


  FA
  g_g1472_n
  (
    .dout(g1472_n),
    .din1(g401_p_spl_0),
    .din2(g1471_p_spl_)
  );


  LA
  g_g1473_p
  (
    .dout(g1473_p),
    .din1(g401_p_spl_),
    .din2(g1471_p_spl_)
  );


  FA
  g_g1473_n
  (
    .dout(g1473_n),
    .din1(g401_n_spl_),
    .din2(g1471_n_spl_)
  );


  LA
  g_g1474_p
  (
    .dout(g1474_p),
    .din1(g1472_n),
    .din2(g1473_n)
  );


  FA
  g_g1474_n
  (
    .dout(g1474_n),
    .din1(g1472_p),
    .din2(g1473_p)
  );


  LA
  g_g1475_p
  (
    .dout(g1475_p),
    .din1(g1470_n_spl_),
    .din2(g1474_p_spl_)
  );


  FA
  g_g1475_n
  (
    .dout(g1475_n),
    .din1(g1470_p_spl_),
    .din2(g1474_n_spl_)
  );


  LA
  g_g1476_p
  (
    .dout(g1476_p),
    .din1(g1470_p_spl_),
    .din2(g1474_n_spl_)
  );


  FA
  g_g1476_n
  (
    .dout(g1476_n),
    .din1(g1470_n_spl_),
    .din2(g1474_p_spl_)
  );


  LA
  g_g1477_p
  (
    .dout(g1477_p),
    .din1(g1475_n),
    .din2(g1476_n)
  );


  FA
  g_g1477_n
  (
    .dout(g1477_n),
    .din1(g1475_p),
    .din2(g1476_p)
  );


  LA
  g_g1478_p
  (
    .dout(g1478_p),
    .din1(g1469_n_spl_),
    .din2(g1477_p_spl_)
  );


  FA
  g_g1478_n
  (
    .dout(g1478_n),
    .din1(g1469_p_spl_),
    .din2(g1477_n_spl_)
  );


  LA
  g_g1479_p
  (
    .dout(g1479_p),
    .din1(g1469_p_spl_),
    .din2(g1477_n_spl_)
  );


  FA
  g_g1479_n
  (
    .dout(g1479_n),
    .din1(g1469_n_spl_),
    .din2(g1477_p_spl_)
  );


  LA
  g_g1480_p
  (
    .dout(g1480_p),
    .din1(g1478_n),
    .din2(g1479_n)
  );


  FA
  g_g1480_n
  (
    .dout(g1480_n),
    .din1(g1478_p),
    .din2(g1479_p)
  );


  LA
  g_g1481_p
  (
    .dout(g1481_p),
    .din1(g429_n_spl_10),
    .din2(g1458_n_spl_1)
  );


  FA
  g_g1481_n
  (
    .dout(g1481_n),
    .din1(g429_p_spl_10),
    .din2(g1458_p_spl_1)
  );


  LA
  g_g1482_p
  (
    .dout(g1482_p),
    .din1(g429_p_spl_1),
    .din2(g1458_p_spl_1)
  );


  FA
  g_g1482_n
  (
    .dout(g1482_n),
    .din1(g429_n_spl_1),
    .din2(g1458_n_spl_1)
  );


  LA
  g_g1483_p
  (
    .dout(g1483_p),
    .din1(g1481_n),
    .din2(g1482_n)
  );


  FA
  g_g1483_n
  (
    .dout(g1483_n),
    .din1(g1481_p),
    .din2(g1482_p)
  );


  LA
  g_g1484_p
  (
    .dout(g1484_p),
    .din1(g1480_n_spl_),
    .din2(g1483_p_spl_)
  );


  FA
  g_g1484_n
  (
    .dout(g1484_n),
    .din1(g1480_p_spl_),
    .din2(g1483_n_spl_)
  );


  LA
  g_g1485_p
  (
    .dout(g1485_p),
    .din1(g1480_p_spl_),
    .din2(g1483_n_spl_)
  );


  FA
  g_g1485_n
  (
    .dout(g1485_n),
    .din1(g1480_n_spl_),
    .din2(g1483_p_spl_)
  );


  LA
  g_g1486_p
  (
    .dout(g1486_p),
    .din1(g1484_n),
    .din2(g1485_n)
  );


  FA
  g_g1486_n
  (
    .dout(g1486_n),
    .din1(g1484_p),
    .din2(g1485_p)
  );


  LA
  g_g1487_p
  (
    .dout(g1487_p),
    .din1(G157_p_spl_1),
    .din2(g1486_n)
  );


  FA
  g_g1487_n
  (
    .dout(g1487_n),
    .din1(G157_n_spl_1),
    .din2(g1486_p)
  );


  LA
  g_g1488_p
  (
    .dout(g1488_p),
    .din1(g1468_n),
    .din2(g1487_n)
  );


  FA
  g_g1488_n
  (
    .dout(g1488_n),
    .din1(g1468_p),
    .din2(g1487_p)
  );


  LA
  g_g1489_p
  (
    .dout(g1489_p),
    .din1(g415_p_spl_1),
    .din2(g1488_p_spl_)
  );


  FA
  g_g1489_n
  (
    .dout(g1489_n),
    .din1(g415_n_spl_1),
    .din2(g1488_n_spl_)
  );


  LA
  g_g1490_p
  (
    .dout(g1490_p),
    .din1(g415_n_spl_1),
    .din2(g1488_n_spl_)
  );


  FA
  g_g1490_n
  (
    .dout(g1490_n),
    .din1(g415_p_spl_1),
    .din2(g1488_p_spl_)
  );


  LA
  g_g1491_p
  (
    .dout(g1491_p),
    .din1(g1489_n),
    .din2(g1490_n)
  );


  FA
  g_g1491_n
  (
    .dout(g1491_n),
    .din1(g1489_p),
    .din2(g1490_p)
  );


  LA
  g_g1492_p
  (
    .dout(g1492_p),
    .din1(g422_p_spl_1),
    .din2(g1491_n_spl_)
  );


  FA
  g_g1492_n
  (
    .dout(g1492_n),
    .din1(g422_n_spl_1),
    .din2(g1491_p_spl_)
  );


  LA
  g_g1493_p
  (
    .dout(g1493_p),
    .din1(g422_n_spl_1),
    .din2(g1491_p_spl_)
  );


  FA
  g_g1493_n
  (
    .dout(g1493_n),
    .din1(g422_p_spl_1),
    .din2(g1491_n_spl_)
  );


  LA
  g_g1494_p
  (
    .dout(g1494_p),
    .din1(g1492_n),
    .din2(g1493_n)
  );


  FA
  g_g1494_n
  (
    .dout(g1494_n),
    .din1(g1492_p),
    .din2(g1493_p)
  );


  LA
  g_g1495_p
  (
    .dout(g1495_p),
    .din1(g1450_n),
    .din2(g1494_n)
  );


  LA
  g_g1496_p
  (
    .dout(g1496_p),
    .din1(g1450_p),
    .din2(g1494_p)
  );


  FA
  g_g1497_n
  (
    .dout(g1497_n),
    .din1(G176_p_spl_1111),
    .din2(g1496_p)
  );


  FA
  g_g1498_n
  (
    .dout(g1498_n),
    .din1(g1495_p),
    .din2(g1497_n)
  );


  LA
  g_g1499_p
  (
    .dout(g1499_p),
    .din1(g1408_n),
    .din2(g1498_n)
  );


  FA
  g_g1500_n
  (
    .dout(g1500_n),
    .din1(G177_n_spl_111),
    .din2(g1499_p)
  );


  FA
  g_g1501_n
  (
    .dout(g1501_n),
    .din1(G49_p),
    .din2(G177_p_spl_110)
  );


  FA
  g_g1502_n
  (
    .dout(g1502_n),
    .din1(G176_n_spl_111),
    .din2(g1501_n)
  );


  LA
  g_g1503_p
  (
    .dout(g1503_p),
    .din1(g1500_n_spl_),
    .din2(g1502_n)
  );


  FA
  g_g1504_n
  (
    .dout(g1504_n),
    .din1(G23_n_spl_),
    .din2(G173_p_spl_111)
  );


  FA
  g_g1505_n
  (
    .dout(g1505_n),
    .din1(G4_n_spl_),
    .din2(G173_n_spl_111)
  );


  LA
  g_g1506_p
  (
    .dout(g1506_p),
    .din1(g1504_n),
    .din2(g1505_n)
  );


  FA
  g_g1507_n
  (
    .dout(g1507_n),
    .din1(G172_p_spl_11),
    .din2(g1506_p)
  );


  FA
  g_g1508_n
  (
    .dout(g1508_n),
    .din1(G38_n),
    .din2(G177_p_spl_111)
  );


  LA
  g_g1509_p
  (
    .dout(g1509_p),
    .din1(g1500_n_spl_),
    .din2(g1508_n)
  );


  LA
  g_g1510_p
  (
    .dout(g1510_p),
    .din1(G173_n_spl_111),
    .din2(g1509_p_spl_0)
  );


  FA
  g_g1511_n
  (
    .dout(g1511_n),
    .din1(G37_n),
    .din2(G177_p_spl_111)
  );


  LA
  g_g1512_p
  (
    .dout(g1512_p),
    .din1(g1308_n_spl_),
    .din2(g1511_n)
  );


  LA
  g_g1513_p
  (
    .dout(g1513_p),
    .din1(G173_p_spl_111),
    .din2(g1512_p_spl_0)
  );


  FA
  g_g1514_n
  (
    .dout(g1514_n),
    .din1(G172_n_spl_11),
    .din2(g1513_p)
  );


  FA
  g_g1515_n
  (
    .dout(g1515_n),
    .din1(g1510_p),
    .din2(g1514_n)
  );


  LA
  g_g1516_p
  (
    .dout(g1516_p),
    .din1(g1507_n),
    .din2(g1515_n)
  );


  FA
  g_g1517_n
  (
    .dout(g1517_n),
    .din1(G23_n_spl_),
    .din2(G174_p_spl_111)
  );


  FA
  g_g1518_n
  (
    .dout(g1518_n),
    .din1(G4_n_spl_),
    .din2(G174_n_spl_111)
  );


  LA
  g_g1519_p
  (
    .dout(g1519_p),
    .din1(g1517_n),
    .din2(g1518_n)
  );


  FA
  g_g1520_n
  (
    .dout(g1520_n),
    .din1(G175_p_spl_11),
    .din2(g1519_p)
  );


  LA
  g_g1521_p
  (
    .dout(g1521_p),
    .din1(G174_n_spl_111),
    .din2(g1509_p_spl_0)
  );


  LA
  g_g1522_p
  (
    .dout(g1522_p),
    .din1(G174_p_spl_111),
    .din2(g1512_p_spl_0)
  );


  FA
  g_g1523_n
  (
    .dout(g1523_n),
    .din1(G175_n_spl_11),
    .din2(g1522_p)
  );


  FA
  g_g1524_n
  (
    .dout(g1524_n),
    .din1(g1521_p),
    .din2(g1523_n)
  );


  LA
  g_g1525_p
  (
    .dout(g1525_p),
    .din1(g1520_n),
    .din2(g1524_n)
  );


  FA
  g_g1526_n
  (
    .dout(g1526_n),
    .din1(G79_n_spl_),
    .din2(G158_p_spl_111)
  );


  FA
  g_g1527_n
  (
    .dout(g1527_n),
    .din1(G78_n_spl_),
    .din2(G158_n_spl_111)
  );


  LA
  g_g1528_p
  (
    .dout(g1528_p),
    .din1(g1526_n),
    .din2(g1527_n)
  );


  FA
  g_g1529_n
  (
    .dout(g1529_n),
    .din1(G159_p_spl_11),
    .din2(g1528_p)
  );


  FA
  g_g1530_n
  (
    .dout(g1530_n),
    .din1(G158_n_spl_111),
    .din2(g1512_p_spl_1)
  );


  FA
  g_g1531_n
  (
    .dout(g1531_n),
    .din1(G158_p_spl_111),
    .din2(g1509_p_spl_1)
  );


  LA
  g_g1532_p
  (
    .dout(g1532_p),
    .din1(g1530_n),
    .din2(g1531_n)
  );


  FA
  g_g1533_n
  (
    .dout(g1533_n),
    .din1(G159_n_spl_11),
    .din2(g1532_p)
  );


  LA
  g_g1534_p
  (
    .dout(g1534_p),
    .din1(g1529_n),
    .din2(g1533_n)
  );


  FA
  g_g1535_n
  (
    .dout(g1535_n),
    .din1(G64_n_spl_),
    .din2(g1534_p)
  );


  FA
  g_g1536_n
  (
    .dout(g1536_n),
    .din1(G79_n_spl_),
    .din2(G160_p_spl_111)
  );


  FA
  g_g1537_n
  (
    .dout(g1537_n),
    .din1(G78_n_spl_),
    .din2(G160_n_spl_111)
  );


  LA
  g_g1538_p
  (
    .dout(g1538_p),
    .din1(g1536_n),
    .din2(g1537_n)
  );


  FA
  g_g1539_n
  (
    .dout(g1539_n),
    .din1(G161_p_spl_11),
    .din2(g1538_p)
  );


  FA
  g_g1540_n
  (
    .dout(g1540_n),
    .din1(G160_n_spl_111),
    .din2(g1512_p_spl_1)
  );


  FA
  g_g1541_n
  (
    .dout(g1541_n),
    .din1(G160_p_spl_111),
    .din2(g1509_p_spl_1)
  );


  LA
  g_g1542_p
  (
    .dout(g1542_p),
    .din1(g1540_n),
    .din2(g1541_n)
  );


  FA
  g_g1543_n
  (
    .dout(g1543_n),
    .din1(G161_n_spl_11),
    .din2(g1542_p)
  );


  LA
  g_g1544_p
  (
    .dout(g1544_p),
    .din1(g1539_n),
    .din2(g1543_n)
  );


  FA
  g_g1545_n
  (
    .dout(g1545_n),
    .din1(G64_n_spl_),
    .din2(g1544_p)
  );


  buf

  (
    G5193_p,
    G66_n
  );


  buf

  (
    G5194_p,
    G113_n_spl_1
  );


  buf

  (
    G5195_p,
    G165_n_spl_
  );


  buf

  (
    G5196_p,
    G151_n_spl_0
  );


  buf

  (
    G5197_p,
    G127_n_spl_
  );


  buf

  (
    G5198_p,
    G131_n_spl_
  );


  buf

  (
    G5199_n,
    g179_n_spl_
  );


  buf

  (
    G5200_p,
    G152_n
  );


  buf

  (
    G5201_p,
    G151_n_spl_0
  );


  buf

  (
    G5202_p,
    G151_n_spl_
  );


  buf

  (
    G5203_p,
    G125_n_spl_
  );


  buf

  (
    G5204_p,
    G129_n_spl_
  );


  buf

  (
    G5205_p,
    g180_p
  );


  buf

  (
    G5206_p,
    G99_n_spl_
  );


  buf

  (
    G5207_p,
    G153_n_spl_
  );


  buf

  (
    G5208_p,
    G156_n_spl_
  );


  buf

  (
    G5209_p,
    G155_n_spl_
  );


  buf

  (
    G5210_p,
    g181_p
  );


  buf

  (
    G5211_p,
    g182_p
  );


  buf

  (
    G5212_p,
    g183_n
  );


  buf

  (
    G5213_p,
    g184_n_spl_
  );


  buf

  (
    G5214_p,
    G64_p_spl_111
  );


  buf

  (
    G5215_p,
    G66_p_spl_1
  );


  buf

  (
    G5216_p,
    G1_p_spl_
  );


  buf

  (
    G5217_p,
    G152_p_spl_
  );


  buf

  (
    G5218_p,
    G114_p_spl_
  );


  buf

  (
    G5219_p,
    G152_p_spl_
  );


  buf

  (
    G5220_p,
    g186_n
  );


  buf

  (
    G5221_p,
    g185_n_spl_11
  );


  buf

  (
    G5222_p,
    G1_n_spl_0
  );


  buf

  (
    G5223_p,
    G1_n_spl_0
  );


  buf

  (
    G5224_p,
    G1_n_spl_1
  );


  buf

  (
    G5225_p,
    G1_n_spl_1
  );


  buf

  (
    G5226_p,
    G114_n_spl_0
  );


  buf

  (
    G5227_p,
    G114_n_spl_
  );


  buf

  (
    G5228_p,
    g190_n
  );


  buf

  (
    G5229_p,
    g194_n_spl_
  );


  buf

  (
    G5230_p,
    g194_n_spl_
  );


  buf

  (
    G5231_p,
    g195_n
  );


  buf

  (
    G5232_p,
    g200_p
  );


  buf

  (
    G5233_p,
    g205_p
  );


  buf

  (
    G5234_p,
    g210_p
  );


  buf

  (
    G5235_p,
    g215_p
  );


  buf

  (
    G5236_n,
    g280_n
  );


  buf

  (
    G5237_n,
    g369_n
  );


  buf

  (
    G5238_n,
    g431_n_spl_
  );


  buf

  (
    G5239_p,
    g482_p_spl_
  );


  buf

  (
    G5240_p,
    g482_p_spl_
  );


  buf

  (
    G5241_n,
    g431_n_spl_
  );


  buf

  (
    G5242_n,
    g506_n_spl_
  );


  buf

  (
    G5243_n,
    g533_n_spl_
  );


  buf

  (
    G5244_n,
    g549_p_spl_
  );


  buf

  (
    G5245_p,
    g550_n_spl_
  );


  buf

  (
    G5246_n,
    g549_p_spl_
  );


  buf

  (
    G5247_p,
    g550_n_spl_
  );


  buf

  (
    G5248_n,
    g560_p_spl_1
  );


  buf

  (
    G5249_n,
    g569_p_spl_1
  );


  buf

  (
    G5250_n,
    g579_p_spl_1
  );


  buf

  (
    G5251_p,
    g581_p_spl_1
  );


  buf

  (
    G5252_p,
    g590_n
  );


  buf

  (
    G5253_n,
    g605_n_spl_1
  );


  buf

  (
    G5254_n,
    g614_n_spl_1
  );


  buf

  (
    G5255_n,
    g624_n_spl_1
  );


  buf

  (
    G5256_p,
    g633_n
  );


  buf

  (
    G5257_n,
    g647_n_spl_1
  );


  buf

  (
    G5258_n,
    g656_n_spl_1
  );


  buf

  (
    G5259_n,
    g669_n_spl_1
  );


  buf

  (
    G5260_n,
    g678_n_spl_1
  );


  buf

  (
    G5261_n,
    g705_n_spl_
  );


  buf

  (
    G5262_n,
    g735_n_spl_
  );


  buf

  (
    G5263_n,
    g764_n
  );


  buf

  (
    G5264_n,
    g794_n
  );


  buf

  (
    G5265_p,
    g804_p
  );


  buf

  (
    G5266_p,
    g814_p
  );


  buf

  (
    G5267_p,
    g823_n
  );


  buf

  (
    G5268_p,
    g832_n
  );


  buf

  (
    G5269_p,
    g841_n
  );


  buf

  (
    G5270_p,
    g850_n
  );


  buf

  (
    G5271_p,
    g859_n
  );


  buf

  (
    G5272_p,
    g868_n
  );


  buf

  (
    G5273_p,
    g877_n
  );


  buf

  (
    G5274_p,
    g886_n
  );


  buf

  (
    G5275_p,
    g896_p
  );


  buf

  (
    G5276_p,
    g906_p
  );


  buf

  (
    G5277_p,
    g916_p
  );


  buf

  (
    G5278_p,
    g926_p
  );


  buf

  (
    G5279_p,
    g936_p
  );


  buf

  (
    G5280_p,
    g946_p
  );


  buf

  (
    G5281_p,
    g956_p
  );


  buf

  (
    G5282_p,
    g966_p
  );


  buf

  (
    G5283_p,
    g980_p
  );


  buf

  (
    G5284_p,
    g983_n
  );


  buf

  (
    G5285_n,
    g990_p_spl_1
  );


  buf

  (
    G5286_n,
    g997_n_spl_1
  );


  buf

  (
    G5287_n,
    g1004_n_spl_1
  );


  buf

  (
    G5288_n,
    g1011_n_spl_1
  );


  buf

  (
    G5289_n,
    g1018_n
  );


  buf

  (
    G5290_n,
    g1025_n_spl_1
  );


  buf

  (
    G5291_n,
    g1032_n_spl_1
  );


  buf

  (
    G5292_n,
    g1039_n_spl_1
  );


  buf

  (
    G5293_n,
    g1046_n_spl_1
  );


  buf

  (
    G5294_p,
    g1055_n
  );


  buf

  (
    G5295_p,
    g1064_n
  );


  buf

  (
    G5296_p,
    g1073_n
  );


  buf

  (
    G5297_p,
    g1082_n
  );


  buf

  (
    G5298_p,
    g1091_n
  );


  buf

  (
    G5299_p,
    g1100_n
  );


  buf

  (
    G5300_p,
    g1109_n
  );


  buf

  (
    G5301_p,
    g1118_n
  );


  buf

  (
    G5302_p,
    g1128_p
  );


  buf

  (
    G5303_p,
    g1138_p
  );


  buf

  (
    G5304_p,
    g1148_p
  );


  buf

  (
    G5305_p,
    g1158_p
  );


  buf

  (
    G5306_p,
    g1168_p
  );


  buf

  (
    G5307_p,
    g1178_p
  );


  buf

  (
    G5308_p,
    g1188_p
  );


  buf

  (
    G5309_p,
    g1198_p
  );


  buf

  (
    G5310_p,
    g1311_p
  );


  buf

  (
    G5311_p,
    g1503_p
  );


  buf

  (
    G5312_n,
    g1516_p
  );


  buf

  (
    G5313_n,
    g1525_p
  );


  buf

  (
    G5314_p,
    g1535_n
  );


  buf

  (
    G5315_p,
    g1545_n
  );


  buf

  (
    G153_n_spl_,
    G153_n
  );


  buf

  (
    G156_n_spl_,
    G156_n
  );


  buf

  (
    G66_p_spl_,
    G66_p
  );


  buf

  (
    G66_p_spl_0,
    G66_p_spl_
  );


  buf

  (
    G66_p_spl_00,
    G66_p_spl_0
  );


  buf

  (
    G66_p_spl_01,
    G66_p_spl_0
  );


  buf

  (
    G66_p_spl_1,
    G66_p_spl_
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G165_n_spl_,
    G165_n
  );


  buf

  (
    G11_n_spl_,
    G11_n
  );


  buf

  (
    g185_n_spl_,
    g185_n
  );


  buf

  (
    g185_n_spl_0,
    g185_n_spl_
  );


  buf

  (
    g185_n_spl_00,
    g185_n_spl_0
  );


  buf

  (
    g185_n_spl_000,
    g185_n_spl_00
  );


  buf

  (
    g185_n_spl_01,
    g185_n_spl_0
  );


  buf

  (
    g185_n_spl_1,
    g185_n_spl_
  );


  buf

  (
    g185_n_spl_10,
    g185_n_spl_1
  );


  buf

  (
    g185_n_spl_11,
    g185_n_spl_1
  );


  buf

  (
    G163_n_spl_,
    G163_n
  );


  buf

  (
    G163_n_spl_0,
    G163_n_spl_
  );


  buf

  (
    G163_n_spl_00,
    G163_n_spl_0
  );


  buf

  (
    G163_n_spl_01,
    G163_n_spl_0
  );


  buf

  (
    G163_n_spl_1,
    G163_n_spl_
  );


  buf

  (
    G163_p_spl_,
    G163_p
  );


  buf

  (
    G163_p_spl_0,
    G163_p_spl_
  );


  buf

  (
    G163_p_spl_00,
    G163_p_spl_0
  );


  buf

  (
    G163_p_spl_01,
    G163_p_spl_0
  );


  buf

  (
    G163_p_spl_1,
    G163_p_spl_
  );


  buf

  (
    G128_p_spl_,
    G128_p
  );


  buf

  (
    G128_p_spl_0,
    G128_p_spl_
  );


  buf

  (
    G128_p_spl_00,
    G128_p_spl_0
  );


  buf

  (
    G128_p_spl_000,
    G128_p_spl_00
  );


  buf

  (
    G128_p_spl_01,
    G128_p_spl_0
  );


  buf

  (
    G128_p_spl_1,
    G128_p_spl_
  );


  buf

  (
    G128_p_spl_10,
    G128_p_spl_1
  );


  buf

  (
    G128_p_spl_11,
    G128_p_spl_1
  );


  buf

  (
    G168_p_spl_,
    G168_p
  );


  buf

  (
    G168_p_spl_0,
    G168_p_spl_
  );


  buf

  (
    G168_p_spl_00,
    G168_p_spl_0
  );


  buf

  (
    G168_p_spl_000,
    G168_p_spl_00
  );


  buf

  (
    G168_p_spl_001,
    G168_p_spl_00
  );


  buf

  (
    G168_p_spl_01,
    G168_p_spl_0
  );


  buf

  (
    G168_p_spl_010,
    G168_p_spl_01
  );


  buf

  (
    G168_p_spl_1,
    G168_p_spl_
  );


  buf

  (
    G168_p_spl_10,
    G168_p_spl_1
  );


  buf

  (
    G168_p_spl_11,
    G168_p_spl_1
  );


  buf

  (
    G128_n_spl_,
    G128_n
  );


  buf

  (
    G128_n_spl_0,
    G128_n_spl_
  );


  buf

  (
    G128_n_spl_00,
    G128_n_spl_0
  );


  buf

  (
    G128_n_spl_000,
    G128_n_spl_00
  );


  buf

  (
    G128_n_spl_01,
    G128_n_spl_0
  );


  buf

  (
    G128_n_spl_1,
    G128_n_spl_
  );


  buf

  (
    G128_n_spl_10,
    G128_n_spl_1
  );


  buf

  (
    G128_n_spl_11,
    G128_n_spl_1
  );


  buf

  (
    G169_p_spl_,
    G169_p
  );


  buf

  (
    G169_p_spl_0,
    G169_p_spl_
  );


  buf

  (
    G169_p_spl_00,
    G169_p_spl_0
  );


  buf

  (
    G169_p_spl_000,
    G169_p_spl_00
  );


  buf

  (
    G169_p_spl_001,
    G169_p_spl_00
  );


  buf

  (
    G169_p_spl_01,
    G169_p_spl_0
  );


  buf

  (
    G169_p_spl_010,
    G169_p_spl_01
  );


  buf

  (
    G169_p_spl_011,
    G169_p_spl_01
  );


  buf

  (
    G169_p_spl_1,
    G169_p_spl_
  );


  buf

  (
    G169_p_spl_10,
    G169_p_spl_1
  );


  buf

  (
    G169_p_spl_11,
    G169_p_spl_1
  );


  buf

  (
    G150_p_spl_,
    G150_p
  );


  buf

  (
    G150_p_spl_0,
    G150_p_spl_
  );


  buf

  (
    G150_p_spl_00,
    G150_p_spl_0
  );


  buf

  (
    G150_p_spl_1,
    G150_p_spl_
  );


  buf

  (
    G167_n_spl_,
    G167_n
  );


  buf

  (
    G167_n_spl_0,
    G167_n_spl_
  );


  buf

  (
    G167_n_spl_00,
    G167_n_spl_0
  );


  buf

  (
    G167_n_spl_000,
    G167_n_spl_00
  );


  buf

  (
    G167_n_spl_001,
    G167_n_spl_00
  );


  buf

  (
    G167_n_spl_01,
    G167_n_spl_0
  );


  buf

  (
    G167_n_spl_010,
    G167_n_spl_01
  );


  buf

  (
    G167_n_spl_1,
    G167_n_spl_
  );


  buf

  (
    G167_n_spl_10,
    G167_n_spl_1
  );


  buf

  (
    G167_n_spl_11,
    G167_n_spl_1
  );


  buf

  (
    G166_n_spl_,
    G166_n
  );


  buf

  (
    G166_n_spl_0,
    G166_n_spl_
  );


  buf

  (
    G166_n_spl_00,
    G166_n_spl_0
  );


  buf

  (
    G166_n_spl_000,
    G166_n_spl_00
  );


  buf

  (
    G166_n_spl_001,
    G166_n_spl_00
  );


  buf

  (
    G166_n_spl_01,
    G166_n_spl_0
  );


  buf

  (
    G166_n_spl_010,
    G166_n_spl_01
  );


  buf

  (
    G166_n_spl_011,
    G166_n_spl_01
  );


  buf

  (
    G166_n_spl_1,
    G166_n_spl_
  );


  buf

  (
    G166_n_spl_10,
    G166_n_spl_1
  );


  buf

  (
    G166_n_spl_11,
    G166_n_spl_1
  );


  buf

  (
    G150_n_spl_,
    G150_n
  );


  buf

  (
    G150_n_spl_0,
    G150_n_spl_
  );


  buf

  (
    G150_n_spl_00,
    G150_n_spl_0
  );


  buf

  (
    G150_n_spl_1,
    G150_n_spl_
  );


  buf

  (
    G126_p_spl_,
    G126_p
  );


  buf

  (
    G126_p_spl_0,
    G126_p_spl_
  );


  buf

  (
    G126_p_spl_00,
    G126_p_spl_0
  );


  buf

  (
    G126_p_spl_000,
    G126_p_spl_00
  );


  buf

  (
    G126_p_spl_01,
    G126_p_spl_0
  );


  buf

  (
    G126_p_spl_1,
    G126_p_spl_
  );


  buf

  (
    G126_p_spl_10,
    G126_p_spl_1
  );


  buf

  (
    G126_p_spl_11,
    G126_p_spl_1
  );


  buf

  (
    G126_n_spl_,
    G126_n
  );


  buf

  (
    G126_n_spl_0,
    G126_n_spl_
  );


  buf

  (
    G126_n_spl_00,
    G126_n_spl_0
  );


  buf

  (
    G126_n_spl_000,
    G126_n_spl_00
  );


  buf

  (
    G126_n_spl_01,
    G126_n_spl_0
  );


  buf

  (
    G126_n_spl_1,
    G126_n_spl_
  );


  buf

  (
    G126_n_spl_10,
    G126_n_spl_1
  );


  buf

  (
    G126_n_spl_11,
    G126_n_spl_1
  );


  buf

  (
    G149_p_spl_,
    G149_p
  );


  buf

  (
    G149_p_spl_0,
    G149_p_spl_
  );


  buf

  (
    G149_p_spl_00,
    G149_p_spl_0
  );


  buf

  (
    G149_p_spl_1,
    G149_p_spl_
  );


  buf

  (
    G149_n_spl_,
    G149_n
  );


  buf

  (
    G149_n_spl_0,
    G149_n_spl_
  );


  buf

  (
    G149_n_spl_00,
    G149_n_spl_0
  );


  buf

  (
    G149_n_spl_1,
    G149_n_spl_
  );


  buf

  (
    g224_n_spl_,
    g224_n
  );


  buf

  (
    g233_n_spl_,
    g233_n
  );


  buf

  (
    G102_p_spl_,
    G102_p
  );


  buf

  (
    G102_p_spl_0,
    G102_p_spl_
  );


  buf

  (
    G102_p_spl_00,
    G102_p_spl_0
  );


  buf

  (
    G102_p_spl_000,
    G102_p_spl_00
  );


  buf

  (
    G102_p_spl_001,
    G102_p_spl_00
  );


  buf

  (
    G102_p_spl_01,
    G102_p_spl_0
  );


  buf

  (
    G102_p_spl_010,
    G102_p_spl_01
  );


  buf

  (
    G102_p_spl_011,
    G102_p_spl_01
  );


  buf

  (
    G102_p_spl_1,
    G102_p_spl_
  );


  buf

  (
    G102_p_spl_10,
    G102_p_spl_1
  );


  buf

  (
    G102_p_spl_100,
    G102_p_spl_10
  );


  buf

  (
    G102_p_spl_101,
    G102_p_spl_10
  );


  buf

  (
    G102_p_spl_11,
    G102_p_spl_1
  );


  buf

  (
    G102_p_spl_110,
    G102_p_spl_11
  );


  buf

  (
    G113_p_spl_,
    G113_p
  );


  buf

  (
    G113_p_spl_0,
    G113_p_spl_
  );


  buf

  (
    G113_p_spl_00,
    G113_p_spl_0
  );


  buf

  (
    G113_p_spl_1,
    G113_p_spl_
  );


  buf

  (
    G102_n_spl_,
    G102_n
  );


  buf

  (
    G102_n_spl_0,
    G102_n_spl_
  );


  buf

  (
    G102_n_spl_00,
    G102_n_spl_0
  );


  buf

  (
    G102_n_spl_000,
    G102_n_spl_00
  );


  buf

  (
    G102_n_spl_001,
    G102_n_spl_00
  );


  buf

  (
    G102_n_spl_01,
    G102_n_spl_0
  );


  buf

  (
    G102_n_spl_010,
    G102_n_spl_01
  );


  buf

  (
    G102_n_spl_011,
    G102_n_spl_01
  );


  buf

  (
    G102_n_spl_1,
    G102_n_spl_
  );


  buf

  (
    G102_n_spl_10,
    G102_n_spl_1
  );


  buf

  (
    G102_n_spl_100,
    G102_n_spl_10
  );


  buf

  (
    G102_n_spl_101,
    G102_n_spl_10
  );


  buf

  (
    G102_n_spl_11,
    G102_n_spl_1
  );


  buf

  (
    G102_n_spl_110,
    G102_n_spl_11
  );


  buf

  (
    G113_n_spl_,
    G113_n
  );


  buf

  (
    G113_n_spl_0,
    G113_n_spl_
  );


  buf

  (
    G113_n_spl_00,
    G113_n_spl_0
  );


  buf

  (
    G113_n_spl_01,
    G113_n_spl_0
  );


  buf

  (
    G113_n_spl_1,
    G113_n_spl_
  );


  buf

  (
    G98_p_spl_,
    G98_p
  );


  buf

  (
    G98_p_spl_0,
    G98_p_spl_
  );


  buf

  (
    G98_p_spl_00,
    G98_p_spl_0
  );


  buf

  (
    G98_p_spl_000,
    G98_p_spl_00
  );


  buf

  (
    G98_p_spl_001,
    G98_p_spl_00
  );


  buf

  (
    G98_p_spl_01,
    G98_p_spl_0
  );


  buf

  (
    G98_p_spl_010,
    G98_p_spl_01
  );


  buf

  (
    G98_p_spl_011,
    G98_p_spl_01
  );


  buf

  (
    G98_p_spl_1,
    G98_p_spl_
  );


  buf

  (
    G98_p_spl_10,
    G98_p_spl_1
  );


  buf

  (
    G98_p_spl_100,
    G98_p_spl_10
  );


  buf

  (
    G98_p_spl_101,
    G98_p_spl_10
  );


  buf

  (
    G98_p_spl_11,
    G98_p_spl_1
  );


  buf

  (
    G98_p_spl_110,
    G98_p_spl_11
  );


  buf

  (
    G98_p_spl_111,
    G98_p_spl_11
  );


  buf

  (
    G98_n_spl_,
    G98_n
  );


  buf

  (
    G98_n_spl_0,
    G98_n_spl_
  );


  buf

  (
    G98_n_spl_00,
    G98_n_spl_0
  );


  buf

  (
    G98_n_spl_000,
    G98_n_spl_00
  );


  buf

  (
    G98_n_spl_001,
    G98_n_spl_00
  );


  buf

  (
    G98_n_spl_01,
    G98_n_spl_0
  );


  buf

  (
    G98_n_spl_010,
    G98_n_spl_01
  );


  buf

  (
    G98_n_spl_011,
    G98_n_spl_01
  );


  buf

  (
    G98_n_spl_1,
    G98_n_spl_
  );


  buf

  (
    G98_n_spl_10,
    G98_n_spl_1
  );


  buf

  (
    G98_n_spl_100,
    G98_n_spl_10
  );


  buf

  (
    G98_n_spl_101,
    G98_n_spl_10
  );


  buf

  (
    G98_n_spl_11,
    G98_n_spl_1
  );


  buf

  (
    G98_n_spl_110,
    G98_n_spl_11
  );


  buf

  (
    G98_n_spl_111,
    G98_n_spl_11
  );


  buf

  (
    G101_p_spl_,
    G101_p
  );


  buf

  (
    G101_p_spl_0,
    G101_p_spl_
  );


  buf

  (
    G101_p_spl_00,
    G101_p_spl_0
  );


  buf

  (
    G101_p_spl_000,
    G101_p_spl_00
  );


  buf

  (
    G101_p_spl_001,
    G101_p_spl_00
  );


  buf

  (
    G101_p_spl_01,
    G101_p_spl_0
  );


  buf

  (
    G101_p_spl_010,
    G101_p_spl_01
  );


  buf

  (
    G101_p_spl_011,
    G101_p_spl_01
  );


  buf

  (
    G101_p_spl_1,
    G101_p_spl_
  );


  buf

  (
    G101_p_spl_10,
    G101_p_spl_1
  );


  buf

  (
    G101_p_spl_100,
    G101_p_spl_10
  );


  buf

  (
    G101_p_spl_101,
    G101_p_spl_10
  );


  buf

  (
    G101_p_spl_11,
    G101_p_spl_1
  );


  buf

  (
    G101_p_spl_110,
    G101_p_spl_11
  );


  buf

  (
    G101_p_spl_111,
    G101_p_spl_11
  );


  buf

  (
    G115_p_spl_,
    G115_p
  );


  buf

  (
    G115_p_spl_0,
    G115_p_spl_
  );


  buf

  (
    G115_p_spl_00,
    G115_p_spl_0
  );


  buf

  (
    G115_p_spl_1,
    G115_p_spl_
  );


  buf

  (
    G101_n_spl_,
    G101_n
  );


  buf

  (
    G101_n_spl_0,
    G101_n_spl_
  );


  buf

  (
    G101_n_spl_00,
    G101_n_spl_0
  );


  buf

  (
    G101_n_spl_000,
    G101_n_spl_00
  );


  buf

  (
    G101_n_spl_001,
    G101_n_spl_00
  );


  buf

  (
    G101_n_spl_01,
    G101_n_spl_0
  );


  buf

  (
    G101_n_spl_010,
    G101_n_spl_01
  );


  buf

  (
    G101_n_spl_011,
    G101_n_spl_01
  );


  buf

  (
    G101_n_spl_1,
    G101_n_spl_
  );


  buf

  (
    G101_n_spl_10,
    G101_n_spl_1
  );


  buf

  (
    G101_n_spl_100,
    G101_n_spl_10
  );


  buf

  (
    G101_n_spl_101,
    G101_n_spl_10
  );


  buf

  (
    G101_n_spl_11,
    G101_n_spl_1
  );


  buf

  (
    G101_n_spl_110,
    G101_n_spl_11
  );


  buf

  (
    G101_n_spl_111,
    G101_n_spl_11
  );


  buf

  (
    G115_n_spl_,
    G115_n
  );


  buf

  (
    G115_n_spl_0,
    G115_n_spl_
  );


  buf

  (
    G115_n_spl_00,
    G115_n_spl_0
  );


  buf

  (
    G115_n_spl_1,
    G115_n_spl_
  );


  buf

  (
    G100_p_spl_,
    G100_p
  );


  buf

  (
    G100_p_spl_0,
    G100_p_spl_
  );


  buf

  (
    G100_p_spl_00,
    G100_p_spl_0
  );


  buf

  (
    G100_p_spl_000,
    G100_p_spl_00
  );


  buf

  (
    G100_p_spl_0000,
    G100_p_spl_000
  );


  buf

  (
    G100_p_spl_001,
    G100_p_spl_00
  );


  buf

  (
    G100_p_spl_01,
    G100_p_spl_0
  );


  buf

  (
    G100_p_spl_010,
    G100_p_spl_01
  );


  buf

  (
    G100_p_spl_011,
    G100_p_spl_01
  );


  buf

  (
    G100_p_spl_1,
    G100_p_spl_
  );


  buf

  (
    G100_p_spl_10,
    G100_p_spl_1
  );


  buf

  (
    G100_p_spl_100,
    G100_p_spl_10
  );


  buf

  (
    G100_p_spl_101,
    G100_p_spl_10
  );


  buf

  (
    G100_p_spl_11,
    G100_p_spl_1
  );


  buf

  (
    G100_p_spl_110,
    G100_p_spl_11
  );


  buf

  (
    G100_p_spl_111,
    G100_p_spl_11
  );


  buf

  (
    G100_n_spl_,
    G100_n
  );


  buf

  (
    G100_n_spl_0,
    G100_n_spl_
  );


  buf

  (
    G100_n_spl_00,
    G100_n_spl_0
  );


  buf

  (
    G100_n_spl_000,
    G100_n_spl_00
  );


  buf

  (
    G100_n_spl_0000,
    G100_n_spl_000
  );


  buf

  (
    G100_n_spl_001,
    G100_n_spl_00
  );


  buf

  (
    G100_n_spl_01,
    G100_n_spl_0
  );


  buf

  (
    G100_n_spl_010,
    G100_n_spl_01
  );


  buf

  (
    G100_n_spl_011,
    G100_n_spl_01
  );


  buf

  (
    G100_n_spl_1,
    G100_n_spl_
  );


  buf

  (
    G100_n_spl_10,
    G100_n_spl_1
  );


  buf

  (
    G100_n_spl_100,
    G100_n_spl_10
  );


  buf

  (
    G100_n_spl_101,
    G100_n_spl_10
  );


  buf

  (
    G100_n_spl_11,
    G100_n_spl_1
  );


  buf

  (
    G100_n_spl_110,
    G100_n_spl_11
  );


  buf

  (
    G100_n_spl_111,
    G100_n_spl_11
  );


  buf

  (
    g237_n_spl_,
    g237_n
  );


  buf

  (
    g237_n_spl_0,
    g237_n_spl_
  );


  buf

  (
    g237_n_spl_1,
    g237_n_spl_
  );


  buf

  (
    g240_p_spl_,
    g240_p
  );


  buf

  (
    g237_p_spl_,
    g237_p
  );


  buf

  (
    g240_n_spl_,
    g240_n
  );


  buf

  (
    g240_n_spl_0,
    g240_n_spl_
  );


  buf

  (
    g241_n_spl_,
    g241_n
  );


  buf

  (
    G130_p_spl_,
    G130_p
  );


  buf

  (
    G130_p_spl_0,
    G130_p_spl_
  );


  buf

  (
    G130_p_spl_00,
    G130_p_spl_0
  );


  buf

  (
    G130_p_spl_1,
    G130_p_spl_
  );


  buf

  (
    G130_n_spl_,
    G130_n
  );


  buf

  (
    G130_n_spl_0,
    G130_n_spl_
  );


  buf

  (
    G130_n_spl_00,
    G130_n_spl_0
  );


  buf

  (
    G130_n_spl_1,
    G130_n_spl_
  );


  buf

  (
    G148_n_spl_,
    G148_n
  );


  buf

  (
    G148_n_spl_0,
    G148_n_spl_
  );


  buf

  (
    G148_n_spl_00,
    G148_n_spl_0
  );


  buf

  (
    G148_n_spl_1,
    G148_n_spl_
  );


  buf

  (
    G148_p_spl_,
    G148_p
  );


  buf

  (
    G148_p_spl_0,
    G148_p_spl_
  );


  buf

  (
    G148_p_spl_00,
    G148_p_spl_0
  );


  buf

  (
    G148_p_spl_1,
    G148_p_spl_
  );


  buf

  (
    g245_n_spl_,
    g245_n
  );


  buf

  (
    g245_n_spl_0,
    g245_n_spl_
  );


  buf

  (
    g245_n_spl_1,
    g245_n_spl_
  );


  buf

  (
    g248_n_spl_,
    g248_n
  );


  buf

  (
    G119_p_spl_,
    G119_p
  );


  buf

  (
    G119_p_spl_0,
    G119_p_spl_
  );


  buf

  (
    G119_p_spl_00,
    G119_p_spl_0
  );


  buf

  (
    G119_p_spl_01,
    G119_p_spl_0
  );


  buf

  (
    G119_p_spl_1,
    G119_p_spl_
  );


  buf

  (
    G119_p_spl_10,
    G119_p_spl_1
  );


  buf

  (
    G119_n_spl_,
    G119_n
  );


  buf

  (
    G119_n_spl_0,
    G119_n_spl_
  );


  buf

  (
    G119_n_spl_00,
    G119_n_spl_0
  );


  buf

  (
    G119_n_spl_01,
    G119_n_spl_0
  );


  buf

  (
    G119_n_spl_1,
    G119_n_spl_
  );


  buf

  (
    G119_n_spl_10,
    G119_n_spl_1
  );


  buf

  (
    G146_p_spl_,
    G146_p
  );


  buf

  (
    G146_p_spl_0,
    G146_p_spl_
  );


  buf

  (
    G146_p_spl_1,
    G146_p_spl_
  );


  buf

  (
    G146_n_spl_,
    G146_n
  );


  buf

  (
    G146_n_spl_0,
    G146_n_spl_
  );


  buf

  (
    G146_n_spl_1,
    G146_n_spl_
  );


  buf

  (
    G117_p_spl_,
    G117_p
  );


  buf

  (
    G117_p_spl_0,
    G117_p_spl_
  );


  buf

  (
    G117_p_spl_00,
    G117_p_spl_0
  );


  buf

  (
    G117_p_spl_01,
    G117_p_spl_0
  );


  buf

  (
    G117_p_spl_1,
    G117_p_spl_
  );


  buf

  (
    G117_p_spl_10,
    G117_p_spl_1
  );


  buf

  (
    G117_n_spl_,
    G117_n
  );


  buf

  (
    G117_n_spl_0,
    G117_n_spl_
  );


  buf

  (
    G117_n_spl_00,
    G117_n_spl_0
  );


  buf

  (
    G117_n_spl_01,
    G117_n_spl_0
  );


  buf

  (
    G117_n_spl_1,
    G117_n_spl_
  );


  buf

  (
    G117_n_spl_10,
    G117_n_spl_1
  );


  buf

  (
    G145_p_spl_,
    G145_p
  );


  buf

  (
    G145_p_spl_0,
    G145_p_spl_
  );


  buf

  (
    G145_p_spl_1,
    G145_p_spl_
  );


  buf

  (
    G145_n_spl_,
    G145_n
  );


  buf

  (
    G145_n_spl_0,
    G145_n_spl_
  );


  buf

  (
    G145_n_spl_1,
    G145_n_spl_
  );


  buf

  (
    g258_p_spl_,
    g258_p
  );


  buf

  (
    g267_p_spl_,
    g267_p
  );


  buf

  (
    g258_n_spl_,
    g258_n
  );


  buf

  (
    g258_n_spl_0,
    g258_n_spl_
  );


  buf

  (
    g267_n_spl_,
    g267_n
  );


  buf

  (
    g267_n_spl_0,
    g267_n_spl_
  );


  buf

  (
    G121_p_spl_,
    G121_p
  );


  buf

  (
    G121_p_spl_0,
    G121_p_spl_
  );


  buf

  (
    G121_p_spl_00,
    G121_p_spl_0
  );


  buf

  (
    G121_p_spl_000,
    G121_p_spl_00
  );


  buf

  (
    G121_p_spl_01,
    G121_p_spl_0
  );


  buf

  (
    G121_p_spl_1,
    G121_p_spl_
  );


  buf

  (
    G121_p_spl_10,
    G121_p_spl_1
  );


  buf

  (
    G121_p_spl_11,
    G121_p_spl_1
  );


  buf

  (
    G121_n_spl_,
    G121_n
  );


  buf

  (
    G121_n_spl_0,
    G121_n_spl_
  );


  buf

  (
    G121_n_spl_00,
    G121_n_spl_0
  );


  buf

  (
    G121_n_spl_000,
    G121_n_spl_00
  );


  buf

  (
    G121_n_spl_01,
    G121_n_spl_0
  );


  buf

  (
    G121_n_spl_1,
    G121_n_spl_
  );


  buf

  (
    G121_n_spl_10,
    G121_n_spl_1
  );


  buf

  (
    G121_n_spl_11,
    G121_n_spl_1
  );


  buf

  (
    G147_p_spl_,
    G147_p
  );


  buf

  (
    G147_p_spl_0,
    G147_p_spl_
  );


  buf

  (
    G147_p_spl_00,
    G147_p_spl_0
  );


  buf

  (
    G147_p_spl_1,
    G147_p_spl_
  );


  buf

  (
    G147_n_spl_,
    G147_n
  );


  buf

  (
    G147_n_spl_0,
    G147_n_spl_
  );


  buf

  (
    G147_n_spl_00,
    G147_n_spl_0
  );


  buf

  (
    G147_n_spl_1,
    G147_n_spl_
  );


  buf

  (
    g268_n_spl_,
    g268_n
  );


  buf

  (
    g277_n_spl_,
    g277_n
  );


  buf

  (
    G107_p_spl_,
    G107_p
  );


  buf

  (
    G107_p_spl_0,
    G107_p_spl_
  );


  buf

  (
    G107_p_spl_00,
    G107_p_spl_0
  );


  buf

  (
    G107_p_spl_000,
    G107_p_spl_00
  );


  buf

  (
    G107_p_spl_01,
    G107_p_spl_0
  );


  buf

  (
    G107_p_spl_1,
    G107_p_spl_
  );


  buf

  (
    G107_p_spl_10,
    G107_p_spl_1
  );


  buf

  (
    G107_p_spl_11,
    G107_p_spl_1
  );


  buf

  (
    G107_n_spl_,
    G107_n
  );


  buf

  (
    G107_n_spl_0,
    G107_n_spl_
  );


  buf

  (
    G107_n_spl_00,
    G107_n_spl_0
  );


  buf

  (
    G107_n_spl_000,
    G107_n_spl_00
  );


  buf

  (
    G107_n_spl_01,
    G107_n_spl_0
  );


  buf

  (
    G107_n_spl_1,
    G107_n_spl_
  );


  buf

  (
    G107_n_spl_10,
    G107_n_spl_1
  );


  buf

  (
    G107_n_spl_11,
    G107_n_spl_1
  );


  buf

  (
    G139_p_spl_,
    G139_p
  );


  buf

  (
    G139_p_spl_0,
    G139_p_spl_
  );


  buf

  (
    G139_p_spl_00,
    G139_p_spl_0
  );


  buf

  (
    G139_p_spl_1,
    G139_p_spl_
  );


  buf

  (
    G139_n_spl_,
    G139_n
  );


  buf

  (
    G139_n_spl_0,
    G139_n_spl_
  );


  buf

  (
    G139_n_spl_00,
    G139_n_spl_0
  );


  buf

  (
    G139_n_spl_1,
    G139_n_spl_
  );


  buf

  (
    G105_p_spl_,
    G105_p
  );


  buf

  (
    G105_p_spl_0,
    G105_p_spl_
  );


  buf

  (
    G105_p_spl_00,
    G105_p_spl_0
  );


  buf

  (
    G105_p_spl_000,
    G105_p_spl_00
  );


  buf

  (
    G105_p_spl_01,
    G105_p_spl_0
  );


  buf

  (
    G105_p_spl_1,
    G105_p_spl_
  );


  buf

  (
    G105_p_spl_10,
    G105_p_spl_1
  );


  buf

  (
    G105_p_spl_11,
    G105_p_spl_1
  );


  buf

  (
    G105_n_spl_,
    G105_n
  );


  buf

  (
    G105_n_spl_0,
    G105_n_spl_
  );


  buf

  (
    G105_n_spl_00,
    G105_n_spl_0
  );


  buf

  (
    G105_n_spl_000,
    G105_n_spl_00
  );


  buf

  (
    G105_n_spl_01,
    G105_n_spl_0
  );


  buf

  (
    G105_n_spl_1,
    G105_n_spl_
  );


  buf

  (
    G105_n_spl_10,
    G105_n_spl_1
  );


  buf

  (
    G105_n_spl_11,
    G105_n_spl_1
  );


  buf

  (
    G138_p_spl_,
    G138_p
  );


  buf

  (
    G138_p_spl_0,
    G138_p_spl_
  );


  buf

  (
    G138_p_spl_00,
    G138_p_spl_0
  );


  buf

  (
    G138_p_spl_1,
    G138_p_spl_
  );


  buf

  (
    G138_n_spl_,
    G138_n
  );


  buf

  (
    G138_n_spl_0,
    G138_n_spl_
  );


  buf

  (
    G138_n_spl_00,
    G138_n_spl_0
  );


  buf

  (
    G138_n_spl_1,
    G138_n_spl_
  );


  buf

  (
    g289_n_spl_,
    g289_n
  );


  buf

  (
    g298_n_spl_,
    g298_n
  );


  buf

  (
    G109_p_spl_,
    G109_p
  );


  buf

  (
    G109_p_spl_0,
    G109_p_spl_
  );


  buf

  (
    G109_p_spl_00,
    G109_p_spl_0
  );


  buf

  (
    G109_p_spl_000,
    G109_p_spl_00
  );


  buf

  (
    G109_p_spl_01,
    G109_p_spl_0
  );


  buf

  (
    G109_p_spl_1,
    G109_p_spl_
  );


  buf

  (
    G109_p_spl_10,
    G109_p_spl_1
  );


  buf

  (
    G109_p_spl_11,
    G109_p_spl_1
  );


  buf

  (
    G109_n_spl_,
    G109_n
  );


  buf

  (
    G109_n_spl_0,
    G109_n_spl_
  );


  buf

  (
    G109_n_spl_00,
    G109_n_spl_0
  );


  buf

  (
    G109_n_spl_000,
    G109_n_spl_00
  );


  buf

  (
    G109_n_spl_01,
    G109_n_spl_0
  );


  buf

  (
    G109_n_spl_1,
    G109_n_spl_
  );


  buf

  (
    G109_n_spl_10,
    G109_n_spl_1
  );


  buf

  (
    G109_n_spl_11,
    G109_n_spl_1
  );


  buf

  (
    G135_p_spl_,
    G135_p
  );


  buf

  (
    G135_p_spl_0,
    G135_p_spl_
  );


  buf

  (
    G135_p_spl_00,
    G135_p_spl_0
  );


  buf

  (
    G135_p_spl_1,
    G135_p_spl_
  );


  buf

  (
    G135_n_spl_,
    G135_n
  );


  buf

  (
    G135_n_spl_0,
    G135_n_spl_
  );


  buf

  (
    G135_n_spl_00,
    G135_n_spl_0
  );


  buf

  (
    G135_n_spl_1,
    G135_n_spl_
  );


  buf

  (
    G88_p_spl_,
    G88_p
  );


  buf

  (
    G88_p_spl_0,
    G88_p_spl_
  );


  buf

  (
    G88_p_spl_00,
    G88_p_spl_0
  );


  buf

  (
    G88_p_spl_01,
    G88_p_spl_0
  );


  buf

  (
    G88_p_spl_1,
    G88_p_spl_
  );


  buf

  (
    G88_p_spl_10,
    G88_p_spl_1
  );


  buf

  (
    G88_n_spl_,
    G88_n
  );


  buf

  (
    G88_n_spl_0,
    G88_n_spl_
  );


  buf

  (
    G88_n_spl_00,
    G88_n_spl_0
  );


  buf

  (
    G88_n_spl_01,
    G88_n_spl_0
  );


  buf

  (
    G88_n_spl_1,
    G88_n_spl_
  );


  buf

  (
    G88_n_spl_10,
    G88_n_spl_1
  );


  buf

  (
    G142_p_spl_,
    G142_p
  );


  buf

  (
    G142_p_spl_0,
    G142_p_spl_
  );


  buf

  (
    G142_p_spl_1,
    G142_p_spl_
  );


  buf

  (
    G142_n_spl_,
    G142_n
  );


  buf

  (
    G142_n_spl_0,
    G142_n_spl_
  );


  buf

  (
    G142_n_spl_1,
    G142_n_spl_
  );


  buf

  (
    g308_n_spl_,
    g308_n
  );


  buf

  (
    g317_n_spl_,
    g317_n
  );


  buf

  (
    g317_n_spl_0,
    g317_n_spl_
  );


  buf

  (
    g317_n_spl_1,
    g317_n_spl_
  );


  buf

  (
    G90_p_spl_,
    G90_p
  );


  buf

  (
    G90_p_spl_0,
    G90_p_spl_
  );


  buf

  (
    G90_p_spl_00,
    G90_p_spl_0
  );


  buf

  (
    G90_p_spl_000,
    G90_p_spl_00
  );


  buf

  (
    G90_p_spl_01,
    G90_p_spl_0
  );


  buf

  (
    G90_p_spl_1,
    G90_p_spl_
  );


  buf

  (
    G90_p_spl_10,
    G90_p_spl_1
  );


  buf

  (
    G90_p_spl_11,
    G90_p_spl_1
  );


  buf

  (
    G90_n_spl_,
    G90_n
  );


  buf

  (
    G90_n_spl_0,
    G90_n_spl_
  );


  buf

  (
    G90_n_spl_00,
    G90_n_spl_0
  );


  buf

  (
    G90_n_spl_000,
    G90_n_spl_00
  );


  buf

  (
    G90_n_spl_01,
    G90_n_spl_0
  );


  buf

  (
    G90_n_spl_1,
    G90_n_spl_
  );


  buf

  (
    G90_n_spl_10,
    G90_n_spl_1
  );


  buf

  (
    G90_n_spl_11,
    G90_n_spl_1
  );


  buf

  (
    G143_p_spl_,
    G143_p
  );


  buf

  (
    G143_p_spl_0,
    G143_p_spl_
  );


  buf

  (
    G143_p_spl_00,
    G143_p_spl_0
  );


  buf

  (
    G143_p_spl_1,
    G143_p_spl_
  );


  buf

  (
    G143_n_spl_,
    G143_n
  );


  buf

  (
    G143_n_spl_0,
    G143_n_spl_
  );


  buf

  (
    G143_n_spl_00,
    G143_n_spl_0
  );


  buf

  (
    G143_n_spl_1,
    G143_n_spl_
  );


  buf

  (
    G92_p_spl_,
    G92_p
  );


  buf

  (
    G92_p_spl_0,
    G92_p_spl_
  );


  buf

  (
    G92_p_spl_00,
    G92_p_spl_0
  );


  buf

  (
    G92_p_spl_000,
    G92_p_spl_00
  );


  buf

  (
    G92_p_spl_01,
    G92_p_spl_0
  );


  buf

  (
    G92_p_spl_1,
    G92_p_spl_
  );


  buf

  (
    G92_p_spl_10,
    G92_p_spl_1
  );


  buf

  (
    G92_p_spl_11,
    G92_p_spl_1
  );


  buf

  (
    G92_n_spl_,
    G92_n
  );


  buf

  (
    G92_n_spl_0,
    G92_n_spl_
  );


  buf

  (
    G92_n_spl_00,
    G92_n_spl_0
  );


  buf

  (
    G92_n_spl_000,
    G92_n_spl_00
  );


  buf

  (
    G92_n_spl_01,
    G92_n_spl_0
  );


  buf

  (
    G92_n_spl_1,
    G92_n_spl_
  );


  buf

  (
    G92_n_spl_10,
    G92_n_spl_1
  );


  buf

  (
    G92_n_spl_11,
    G92_n_spl_1
  );


  buf

  (
    G144_p_spl_,
    G144_p
  );


  buf

  (
    G144_p_spl_0,
    G144_p_spl_
  );


  buf

  (
    G144_p_spl_00,
    G144_p_spl_0
  );


  buf

  (
    G144_p_spl_1,
    G144_p_spl_
  );


  buf

  (
    G144_n_spl_,
    G144_n
  );


  buf

  (
    G144_n_spl_0,
    G144_n_spl_
  );


  buf

  (
    G144_n_spl_00,
    G144_n_spl_0
  );


  buf

  (
    G144_n_spl_1,
    G144_n_spl_
  );


  buf

  (
    g328_n_spl_,
    g328_n
  );


  buf

  (
    g337_n_spl_,
    g337_n
  );


  buf

  (
    G94_p_spl_,
    G94_p
  );


  buf

  (
    G94_p_spl_0,
    G94_p_spl_
  );


  buf

  (
    G94_p_spl_00,
    G94_p_spl_0
  );


  buf

  (
    G94_p_spl_000,
    G94_p_spl_00
  );


  buf

  (
    G94_p_spl_01,
    G94_p_spl_0
  );


  buf

  (
    G94_p_spl_1,
    G94_p_spl_
  );


  buf

  (
    G94_p_spl_10,
    G94_p_spl_1
  );


  buf

  (
    G94_p_spl_11,
    G94_p_spl_1
  );


  buf

  (
    G94_n_spl_,
    G94_n
  );


  buf

  (
    G94_n_spl_0,
    G94_n_spl_
  );


  buf

  (
    G94_n_spl_00,
    G94_n_spl_0
  );


  buf

  (
    G94_n_spl_000,
    G94_n_spl_00
  );


  buf

  (
    G94_n_spl_01,
    G94_n_spl_0
  );


  buf

  (
    G94_n_spl_1,
    G94_n_spl_
  );


  buf

  (
    G94_n_spl_10,
    G94_n_spl_1
  );


  buf

  (
    G94_n_spl_11,
    G94_n_spl_1
  );


  buf

  (
    G140_p_spl_,
    G140_p
  );


  buf

  (
    G140_p_spl_0,
    G140_p_spl_
  );


  buf

  (
    G140_p_spl_00,
    G140_p_spl_0
  );


  buf

  (
    G140_p_spl_1,
    G140_p_spl_
  );


  buf

  (
    G140_n_spl_,
    G140_n
  );


  buf

  (
    G140_n_spl_0,
    G140_n_spl_
  );


  buf

  (
    G140_n_spl_00,
    G140_n_spl_0
  );


  buf

  (
    G140_n_spl_1,
    G140_n_spl_
  );


  buf

  (
    G96_p_spl_,
    G96_p
  );


  buf

  (
    G96_p_spl_0,
    G96_p_spl_
  );


  buf

  (
    G96_p_spl_00,
    G96_p_spl_0
  );


  buf

  (
    G96_p_spl_000,
    G96_p_spl_00
  );


  buf

  (
    G96_p_spl_01,
    G96_p_spl_0
  );


  buf

  (
    G96_p_spl_1,
    G96_p_spl_
  );


  buf

  (
    G96_p_spl_10,
    G96_p_spl_1
  );


  buf

  (
    G96_p_spl_11,
    G96_p_spl_1
  );


  buf

  (
    G96_n_spl_,
    G96_n
  );


  buf

  (
    G96_n_spl_0,
    G96_n_spl_
  );


  buf

  (
    G96_n_spl_00,
    G96_n_spl_0
  );


  buf

  (
    G96_n_spl_000,
    G96_n_spl_00
  );


  buf

  (
    G96_n_spl_01,
    G96_n_spl_0
  );


  buf

  (
    G96_n_spl_1,
    G96_n_spl_
  );


  buf

  (
    G96_n_spl_10,
    G96_n_spl_1
  );


  buf

  (
    G96_n_spl_11,
    G96_n_spl_1
  );


  buf

  (
    G141_p_spl_,
    G141_p
  );


  buf

  (
    G141_p_spl_0,
    G141_p_spl_
  );


  buf

  (
    G141_p_spl_00,
    G141_p_spl_0
  );


  buf

  (
    G141_p_spl_1,
    G141_p_spl_
  );


  buf

  (
    G141_n_spl_,
    G141_n
  );


  buf

  (
    G141_n_spl_0,
    G141_n_spl_
  );


  buf

  (
    G141_n_spl_00,
    G141_n_spl_0
  );


  buf

  (
    G141_n_spl_1,
    G141_n_spl_
  );


  buf

  (
    G103_p_spl_,
    G103_p
  );


  buf

  (
    G103_p_spl_0,
    G103_p_spl_
  );


  buf

  (
    G103_p_spl_00,
    G103_p_spl_0
  );


  buf

  (
    G103_p_spl_000,
    G103_p_spl_00
  );


  buf

  (
    G103_p_spl_01,
    G103_p_spl_0
  );


  buf

  (
    G103_p_spl_1,
    G103_p_spl_
  );


  buf

  (
    G103_p_spl_10,
    G103_p_spl_1
  );


  buf

  (
    G103_p_spl_11,
    G103_p_spl_1
  );


  buf

  (
    G103_n_spl_,
    G103_n
  );


  buf

  (
    G103_n_spl_0,
    G103_n_spl_
  );


  buf

  (
    G103_n_spl_00,
    G103_n_spl_0
  );


  buf

  (
    G103_n_spl_000,
    G103_n_spl_00
  );


  buf

  (
    G103_n_spl_01,
    G103_n_spl_0
  );


  buf

  (
    G103_n_spl_1,
    G103_n_spl_
  );


  buf

  (
    G103_n_spl_10,
    G103_n_spl_1
  );


  buf

  (
    G103_n_spl_11,
    G103_n_spl_1
  );


  buf

  (
    G137_p_spl_,
    G137_p
  );


  buf

  (
    G137_p_spl_0,
    G137_p_spl_
  );


  buf

  (
    G137_p_spl_00,
    G137_p_spl_0
  );


  buf

  (
    G137_p_spl_1,
    G137_p_spl_
  );


  buf

  (
    G137_n_spl_,
    G137_n
  );


  buf

  (
    G137_n_spl_0,
    G137_n_spl_
  );


  buf

  (
    G137_n_spl_00,
    G137_n_spl_0
  );


  buf

  (
    G137_n_spl_1,
    G137_n_spl_
  );


  buf

  (
    g356_n_spl_,
    g356_n
  );


  buf

  (
    g365_n_spl_,
    g365_n
  );


  buf

  (
    g347_n_spl_,
    g347_n
  );


  buf

  (
    G124_n_spl_,
    G124_n
  );


  buf

  (
    G124_n_spl_0,
    G124_n_spl_
  );


  buf

  (
    G124_n_spl_00,
    G124_n_spl_0
  );


  buf

  (
    G124_n_spl_000,
    G124_n_spl_00
  );


  buf

  (
    G124_n_spl_0000,
    G124_n_spl_000
  );


  buf

  (
    G124_n_spl_0001,
    G124_n_spl_000
  );


  buf

  (
    G124_n_spl_001,
    G124_n_spl_00
  );


  buf

  (
    G124_n_spl_0010,
    G124_n_spl_001
  );


  buf

  (
    G124_n_spl_0011,
    G124_n_spl_001
  );


  buf

  (
    G124_n_spl_01,
    G124_n_spl_0
  );


  buf

  (
    G124_n_spl_010,
    G124_n_spl_01
  );


  buf

  (
    G124_n_spl_011,
    G124_n_spl_01
  );


  buf

  (
    G124_n_spl_1,
    G124_n_spl_
  );


  buf

  (
    G124_n_spl_10,
    G124_n_spl_1
  );


  buf

  (
    G124_n_spl_100,
    G124_n_spl_10
  );


  buf

  (
    G124_n_spl_101,
    G124_n_spl_10
  );


  buf

  (
    G124_n_spl_11,
    G124_n_spl_1
  );


  buf

  (
    G124_n_spl_110,
    G124_n_spl_11
  );


  buf

  (
    G124_n_spl_111,
    G124_n_spl_11
  );


  buf

  (
    G124_p_spl_,
    G124_p
  );


  buf

  (
    G124_p_spl_0,
    G124_p_spl_
  );


  buf

  (
    G124_p_spl_00,
    G124_p_spl_0
  );


  buf

  (
    G124_p_spl_000,
    G124_p_spl_00
  );


  buf

  (
    G124_p_spl_0000,
    G124_p_spl_000
  );


  buf

  (
    G124_p_spl_0001,
    G124_p_spl_000
  );


  buf

  (
    G124_p_spl_001,
    G124_p_spl_00
  );


  buf

  (
    G124_p_spl_0010,
    G124_p_spl_001
  );


  buf

  (
    G124_p_spl_0011,
    G124_p_spl_001
  );


  buf

  (
    G124_p_spl_01,
    G124_p_spl_0
  );


  buf

  (
    G124_p_spl_010,
    G124_p_spl_01
  );


  buf

  (
    G124_p_spl_011,
    G124_p_spl_01
  );


  buf

  (
    G124_p_spl_1,
    G124_p_spl_
  );


  buf

  (
    G124_p_spl_10,
    G124_p_spl_1
  );


  buf

  (
    G124_p_spl_100,
    G124_p_spl_10
  );


  buf

  (
    G124_p_spl_101,
    G124_p_spl_10
  );


  buf

  (
    G124_p_spl_11,
    G124_p_spl_1
  );


  buf

  (
    G124_p_spl_110,
    G124_p_spl_11
  );


  buf

  (
    G124_p_spl_111,
    G124_p_spl_11
  );


  buf

  (
    g372_p_spl_,
    g372_p
  );


  buf

  (
    g372_p_spl_0,
    g372_p_spl_
  );


  buf

  (
    g372_p_spl_1,
    g372_p_spl_
  );


  buf

  (
    g372_n_spl_,
    g372_n
  );


  buf

  (
    g372_n_spl_0,
    g372_n_spl_
  );


  buf

  (
    g372_n_spl_1,
    g372_n_spl_
  );


  buf

  (
    g373_n_spl_,
    g373_n
  );


  buf

  (
    g373_n_spl_0,
    g373_n_spl_
  );


  buf

  (
    g374_n_spl_,
    g374_n
  );


  buf

  (
    g374_n_spl_0,
    g374_n_spl_
  );


  buf

  (
    g374_n_spl_1,
    g374_n_spl_
  );


  buf

  (
    g373_p_spl_,
    g373_p
  );


  buf

  (
    g373_p_spl_0,
    g373_p_spl_
  );


  buf

  (
    g374_p_spl_,
    g374_p
  );


  buf

  (
    g374_p_spl_0,
    g374_p_spl_
  );


  buf

  (
    g374_p_spl_1,
    g374_p_spl_
  );


  buf

  (
    g378_p_spl_,
    g378_p
  );


  buf

  (
    g378_p_spl_0,
    g378_p_spl_
  );


  buf

  (
    g378_p_spl_1,
    g378_p_spl_
  );


  buf

  (
    g378_n_spl_,
    g378_n
  );


  buf

  (
    g378_n_spl_0,
    g378_n_spl_
  );


  buf

  (
    g378_n_spl_1,
    g378_n_spl_
  );


  buf

  (
    g379_n_spl_,
    g379_n
  );


  buf

  (
    g380_n_spl_,
    g380_n
  );


  buf

  (
    g379_p_spl_,
    g379_p
  );


  buf

  (
    g380_p_spl_,
    g380_p
  );


  buf

  (
    g375_p_spl_,
    g375_p
  );


  buf

  (
    g375_p_spl_0,
    g375_p_spl_
  );


  buf

  (
    g375_p_spl_00,
    g375_p_spl_0
  );


  buf

  (
    g375_p_spl_1,
    g375_p_spl_
  );


  buf

  (
    g381_p_spl_,
    g381_p
  );


  buf

  (
    g381_p_spl_0,
    g381_p_spl_
  );


  buf

  (
    g381_p_spl_00,
    g381_p_spl_0
  );


  buf

  (
    g381_p_spl_01,
    g381_p_spl_0
  );


  buf

  (
    g381_p_spl_1,
    g381_p_spl_
  );


  buf

  (
    g381_p_spl_10,
    g381_p_spl_1
  );


  buf

  (
    g375_n_spl_,
    g375_n
  );


  buf

  (
    g375_n_spl_0,
    g375_n_spl_
  );


  buf

  (
    g375_n_spl_00,
    g375_n_spl_0
  );


  buf

  (
    g375_n_spl_1,
    g375_n_spl_
  );


  buf

  (
    g381_n_spl_,
    g381_n
  );


  buf

  (
    g381_n_spl_0,
    g381_n_spl_
  );


  buf

  (
    g381_n_spl_00,
    g381_n_spl_0
  );


  buf

  (
    g381_n_spl_01,
    g381_n_spl_0
  );


  buf

  (
    g381_n_spl_1,
    g381_n_spl_
  );


  buf

  (
    g381_n_spl_10,
    g381_n_spl_1
  );


  buf

  (
    g385_p_spl_,
    g385_p
  );


  buf

  (
    g385_p_spl_0,
    g385_p_spl_
  );


  buf

  (
    g385_p_spl_1,
    g385_p_spl_
  );


  buf

  (
    g385_n_spl_,
    g385_n
  );


  buf

  (
    g385_n_spl_0,
    g385_n_spl_
  );


  buf

  (
    g385_n_spl_1,
    g385_n_spl_
  );


  buf

  (
    g386_n_spl_,
    g386_n
  );


  buf

  (
    g387_n_spl_,
    g387_n
  );


  buf

  (
    g386_p_spl_,
    g386_p
  );


  buf

  (
    g387_p_spl_,
    g387_p
  );


  buf

  (
    g382_p_spl_,
    g382_p
  );


  buf

  (
    g388_p_spl_,
    g388_p
  );


  buf

  (
    g388_p_spl_0,
    g388_p_spl_
  );


  buf

  (
    g388_p_spl_00,
    g388_p_spl_0
  );


  buf

  (
    g388_p_spl_01,
    g388_p_spl_0
  );


  buf

  (
    g388_p_spl_1,
    g388_p_spl_
  );


  buf

  (
    g382_n_spl_,
    g382_n
  );


  buf

  (
    g388_n_spl_,
    g388_n
  );


  buf

  (
    g388_n_spl_0,
    g388_n_spl_
  );


  buf

  (
    g388_n_spl_00,
    g388_n_spl_0
  );


  buf

  (
    g388_n_spl_01,
    g388_n_spl_0
  );


  buf

  (
    g388_n_spl_1,
    g388_n_spl_
  );


  buf

  (
    g392_p_spl_,
    g392_p
  );


  buf

  (
    g392_p_spl_0,
    g392_p_spl_
  );


  buf

  (
    g392_p_spl_1,
    g392_p_spl_
  );


  buf

  (
    g392_n_spl_,
    g392_n
  );


  buf

  (
    g392_n_spl_0,
    g392_n_spl_
  );


  buf

  (
    g392_n_spl_1,
    g392_n_spl_
  );


  buf

  (
    g393_n_spl_,
    g393_n
  );


  buf

  (
    g389_n_spl_,
    g389_n
  );


  buf

  (
    g389_n_spl_0,
    g389_n_spl_
  );


  buf

  (
    g395_n_spl_,
    g395_n
  );


  buf

  (
    g395_n_spl_0,
    g395_n_spl_
  );


  buf

  (
    g395_n_spl_00,
    g395_n_spl_0
  );


  buf

  (
    g395_n_spl_01,
    g395_n_spl_0
  );


  buf

  (
    g395_n_spl_1,
    g395_n_spl_
  );


  buf

  (
    g395_n_spl_10,
    g395_n_spl_1
  );


  buf

  (
    g399_p_spl_,
    g399_p
  );


  buf

  (
    g399_p_spl_0,
    g399_p_spl_
  );


  buf

  (
    g399_p_spl_1,
    g399_p_spl_
  );


  buf

  (
    g399_n_spl_,
    g399_n
  );


  buf

  (
    g399_n_spl_0,
    g399_n_spl_
  );


  buf

  (
    g399_n_spl_1,
    g399_n_spl_
  );


  buf

  (
    g400_n_spl_,
    g400_n
  );


  buf

  (
    g400_n_spl_0,
    g400_n_spl_
  );


  buf

  (
    g400_n_spl_00,
    g400_n_spl_0
  );


  buf

  (
    g400_n_spl_1,
    g400_n_spl_
  );


  buf

  (
    g401_n_spl_,
    g401_n
  );


  buf

  (
    g401_n_spl_0,
    g401_n_spl_
  );


  buf

  (
    g400_p_spl_,
    g400_p
  );


  buf

  (
    g400_p_spl_0,
    g400_p_spl_
  );


  buf

  (
    g400_p_spl_00,
    g400_p_spl_0
  );


  buf

  (
    g400_p_spl_1,
    g400_p_spl_
  );


  buf

  (
    g401_p_spl_,
    g401_p
  );


  buf

  (
    g401_p_spl_0,
    g401_p_spl_
  );


  buf

  (
    g405_p_spl_,
    g405_p
  );


  buf

  (
    g405_p_spl_0,
    g405_p_spl_
  );


  buf

  (
    g405_p_spl_1,
    g405_p_spl_
  );


  buf

  (
    g405_n_spl_,
    g405_n
  );


  buf

  (
    g405_n_spl_0,
    g405_n_spl_
  );


  buf

  (
    g405_n_spl_1,
    g405_n_spl_
  );


  buf

  (
    g406_n_spl_,
    g406_n
  );


  buf

  (
    g406_n_spl_0,
    g406_n_spl_
  );


  buf

  (
    g406_p_spl_,
    g406_p
  );


  buf

  (
    g406_p_spl_0,
    g406_p_spl_
  );


  buf

  (
    g402_p_spl_,
    g402_p
  );


  buf

  (
    g402_p_spl_0,
    g402_p_spl_
  );


  buf

  (
    g402_p_spl_1,
    g402_p_spl_
  );


  buf

  (
    g408_p_spl_,
    g408_p
  );


  buf

  (
    g408_p_spl_0,
    g408_p_spl_
  );


  buf

  (
    g408_p_spl_1,
    g408_p_spl_
  );


  buf

  (
    g402_n_spl_,
    g402_n
  );


  buf

  (
    g402_n_spl_0,
    g402_n_spl_
  );


  buf

  (
    g408_n_spl_,
    g408_n
  );


  buf

  (
    g408_n_spl_0,
    g408_n_spl_
  );


  buf

  (
    g408_n_spl_00,
    g408_n_spl_0
  );


  buf

  (
    g408_n_spl_1,
    g408_n_spl_
  );


  buf

  (
    g412_p_spl_,
    g412_p
  );


  buf

  (
    g412_p_spl_0,
    g412_p_spl_
  );


  buf

  (
    g412_p_spl_1,
    g412_p_spl_
  );


  buf

  (
    g412_n_spl_,
    g412_n
  );


  buf

  (
    g412_n_spl_0,
    g412_n_spl_
  );


  buf

  (
    g412_n_spl_1,
    g412_n_spl_
  );


  buf

  (
    g413_n_spl_,
    g413_n
  );


  buf

  (
    g413_p_spl_,
    g413_p
  );


  buf

  (
    g409_p_spl_,
    g409_p
  );


  buf

  (
    g409_p_spl_0,
    g409_p_spl_
  );


  buf

  (
    g415_p_spl_,
    g415_p
  );


  buf

  (
    g415_p_spl_0,
    g415_p_spl_
  );


  buf

  (
    g415_p_spl_00,
    g415_p_spl_0
  );


  buf

  (
    g415_p_spl_1,
    g415_p_spl_
  );


  buf

  (
    g409_n_spl_,
    g409_n
  );


  buf

  (
    g409_n_spl_0,
    g409_n_spl_
  );


  buf

  (
    g415_n_spl_,
    g415_n
  );


  buf

  (
    g415_n_spl_0,
    g415_n_spl_
  );


  buf

  (
    g415_n_spl_00,
    g415_n_spl_0
  );


  buf

  (
    g415_n_spl_1,
    g415_n_spl_
  );


  buf

  (
    g419_p_spl_,
    g419_p
  );


  buf

  (
    g419_p_spl_0,
    g419_p_spl_
  );


  buf

  (
    g419_p_spl_1,
    g419_p_spl_
  );


  buf

  (
    g419_n_spl_,
    g419_n
  );


  buf

  (
    g419_n_spl_0,
    g419_n_spl_
  );


  buf

  (
    g419_n_spl_1,
    g419_n_spl_
  );


  buf

  (
    g420_n_spl_,
    g420_n
  );


  buf

  (
    g420_n_spl_0,
    g420_n_spl_
  );


  buf

  (
    g420_p_spl_,
    g420_p
  );


  buf

  (
    g420_p_spl_0,
    g420_p_spl_
  );


  buf

  (
    g416_p_spl_,
    g416_p
  );


  buf

  (
    g416_p_spl_0,
    g416_p_spl_
  );


  buf

  (
    g422_p_spl_,
    g422_p
  );


  buf

  (
    g422_p_spl_0,
    g422_p_spl_
  );


  buf

  (
    g422_p_spl_00,
    g422_p_spl_0
  );


  buf

  (
    g422_p_spl_1,
    g422_p_spl_
  );


  buf

  (
    g416_n_spl_,
    g416_n
  );


  buf

  (
    g416_n_spl_0,
    g416_n_spl_
  );


  buf

  (
    g422_n_spl_,
    g422_n
  );


  buf

  (
    g422_n_spl_0,
    g422_n_spl_
  );


  buf

  (
    g422_n_spl_00,
    g422_n_spl_0
  );


  buf

  (
    g422_n_spl_01,
    g422_n_spl_0
  );


  buf

  (
    g422_n_spl_1,
    g422_n_spl_
  );


  buf

  (
    g426_p_spl_,
    g426_p
  );


  buf

  (
    g426_p_spl_0,
    g426_p_spl_
  );


  buf

  (
    g426_p_spl_1,
    g426_p_spl_
  );


  buf

  (
    g426_n_spl_,
    g426_n
  );


  buf

  (
    g426_n_spl_0,
    g426_n_spl_
  );


  buf

  (
    g426_n_spl_1,
    g426_n_spl_
  );


  buf

  (
    g427_n_spl_,
    g427_n
  );


  buf

  (
    g427_p_spl_,
    g427_p
  );


  buf

  (
    g423_p_spl_,
    g423_p
  );


  buf

  (
    g429_p_spl_,
    g429_p
  );


  buf

  (
    g429_p_spl_0,
    g429_p_spl_
  );


  buf

  (
    g429_p_spl_00,
    g429_p_spl_0
  );


  buf

  (
    g429_p_spl_01,
    g429_p_spl_0
  );


  buf

  (
    g429_p_spl_1,
    g429_p_spl_
  );


  buf

  (
    g429_p_spl_10,
    g429_p_spl_1
  );


  buf

  (
    g423_n_spl_,
    g423_n
  );


  buf

  (
    g429_n_spl_,
    g429_n
  );


  buf

  (
    g429_n_spl_0,
    g429_n_spl_
  );


  buf

  (
    g429_n_spl_00,
    g429_n_spl_0
  );


  buf

  (
    g429_n_spl_01,
    g429_n_spl_0
  );


  buf

  (
    g429_n_spl_1,
    g429_n_spl_
  );


  buf

  (
    g429_n_spl_10,
    g429_n_spl_1
  );


  buf

  (
    g396_n_spl_,
    g396_n
  );


  buf

  (
    g430_n_spl_,
    g430_n
  );


  buf

  (
    g430_n_spl_0,
    g430_n_spl_
  );


  buf

  (
    g430_n_spl_1,
    g430_n_spl_
  );


  buf

  (
    G123_n_spl_,
    G123_n
  );


  buf

  (
    G123_n_spl_0,
    G123_n_spl_
  );


  buf

  (
    G123_n_spl_00,
    G123_n_spl_0
  );


  buf

  (
    G123_n_spl_000,
    G123_n_spl_00
  );


  buf

  (
    G123_n_spl_0000,
    G123_n_spl_000
  );


  buf

  (
    G123_n_spl_0001,
    G123_n_spl_000
  );


  buf

  (
    G123_n_spl_001,
    G123_n_spl_00
  );


  buf

  (
    G123_n_spl_0010,
    G123_n_spl_001
  );


  buf

  (
    G123_n_spl_01,
    G123_n_spl_0
  );


  buf

  (
    G123_n_spl_010,
    G123_n_spl_01
  );


  buf

  (
    G123_n_spl_011,
    G123_n_spl_01
  );


  buf

  (
    G123_n_spl_1,
    G123_n_spl_
  );


  buf

  (
    G123_n_spl_10,
    G123_n_spl_1
  );


  buf

  (
    G123_n_spl_100,
    G123_n_spl_10
  );


  buf

  (
    G123_n_spl_101,
    G123_n_spl_10
  );


  buf

  (
    G123_n_spl_11,
    G123_n_spl_1
  );


  buf

  (
    G123_n_spl_110,
    G123_n_spl_11
  );


  buf

  (
    G123_n_spl_111,
    G123_n_spl_11
  );


  buf

  (
    G123_p_spl_,
    G123_p
  );


  buf

  (
    G123_p_spl_0,
    G123_p_spl_
  );


  buf

  (
    G123_p_spl_00,
    G123_p_spl_0
  );


  buf

  (
    G123_p_spl_000,
    G123_p_spl_00
  );


  buf

  (
    G123_p_spl_0000,
    G123_p_spl_000
  );


  buf

  (
    G123_p_spl_0001,
    G123_p_spl_000
  );


  buf

  (
    G123_p_spl_001,
    G123_p_spl_00
  );


  buf

  (
    G123_p_spl_0010,
    G123_p_spl_001
  );


  buf

  (
    G123_p_spl_01,
    G123_p_spl_0
  );


  buf

  (
    G123_p_spl_010,
    G123_p_spl_01
  );


  buf

  (
    G123_p_spl_011,
    G123_p_spl_01
  );


  buf

  (
    G123_p_spl_1,
    G123_p_spl_
  );


  buf

  (
    G123_p_spl_10,
    G123_p_spl_1
  );


  buf

  (
    G123_p_spl_100,
    G123_p_spl_10
  );


  buf

  (
    G123_p_spl_101,
    G123_p_spl_10
  );


  buf

  (
    G123_p_spl_11,
    G123_p_spl_1
  );


  buf

  (
    G123_p_spl_110,
    G123_p_spl_11
  );


  buf

  (
    G123_p_spl_111,
    G123_p_spl_11
  );


  buf

  (
    g434_p_spl_,
    g434_p
  );


  buf

  (
    g434_p_spl_0,
    g434_p_spl_
  );


  buf

  (
    g434_p_spl_1,
    g434_p_spl_
  );


  buf

  (
    g434_n_spl_,
    g434_n
  );


  buf

  (
    g434_n_spl_0,
    g434_n_spl_
  );


  buf

  (
    g434_n_spl_1,
    g434_n_spl_
  );


  buf

  (
    g435_n_spl_,
    g435_n
  );


  buf

  (
    g435_p_spl_,
    g435_p
  );


  buf

  (
    g440_p_spl_,
    g440_p
  );


  buf

  (
    g440_p_spl_0,
    g440_p_spl_
  );


  buf

  (
    g440_p_spl_1,
    g440_p_spl_
  );


  buf

  (
    g440_n_spl_,
    g440_n
  );


  buf

  (
    g440_n_spl_0,
    g440_n_spl_
  );


  buf

  (
    g440_n_spl_1,
    g440_n_spl_
  );


  buf

  (
    g441_n_spl_,
    g441_n
  );


  buf

  (
    g441_n_spl_0,
    g441_n_spl_
  );


  buf

  (
    g441_n_spl_00,
    g441_n_spl_0
  );


  buf

  (
    g441_n_spl_1,
    g441_n_spl_
  );


  buf

  (
    g442_n_spl_,
    g442_n
  );


  buf

  (
    g442_n_spl_0,
    g442_n_spl_
  );


  buf

  (
    g442_n_spl_1,
    g442_n_spl_
  );


  buf

  (
    g441_p_spl_,
    g441_p
  );


  buf

  (
    g441_p_spl_0,
    g441_p_spl_
  );


  buf

  (
    g441_p_spl_00,
    g441_p_spl_0
  );


  buf

  (
    g441_p_spl_1,
    g441_p_spl_
  );


  buf

  (
    g442_p_spl_,
    g442_p
  );


  buf

  (
    g442_p_spl_0,
    g442_p_spl_
  );


  buf

  (
    g442_p_spl_1,
    g442_p_spl_
  );


  buf

  (
    g437_p_spl_,
    g437_p
  );


  buf

  (
    g437_p_spl_0,
    g437_p_spl_
  );


  buf

  (
    g437_p_spl_00,
    g437_p_spl_0
  );


  buf

  (
    g437_p_spl_01,
    g437_p_spl_0
  );


  buf

  (
    g437_p_spl_1,
    g437_p_spl_
  );


  buf

  (
    g443_p_spl_,
    g443_p
  );


  buf

  (
    g443_p_spl_0,
    g443_p_spl_
  );


  buf

  (
    g443_p_spl_00,
    g443_p_spl_0
  );


  buf

  (
    g443_p_spl_1,
    g443_p_spl_
  );


  buf

  (
    g437_n_spl_,
    g437_n
  );


  buf

  (
    g437_n_spl_0,
    g437_n_spl_
  );


  buf

  (
    g437_n_spl_00,
    g437_n_spl_0
  );


  buf

  (
    g437_n_spl_01,
    g437_n_spl_0
  );


  buf

  (
    g437_n_spl_1,
    g437_n_spl_
  );


  buf

  (
    g443_n_spl_,
    g443_n
  );


  buf

  (
    g443_n_spl_0,
    g443_n_spl_
  );


  buf

  (
    g443_n_spl_00,
    g443_n_spl_0
  );


  buf

  (
    g443_n_spl_1,
    g443_n_spl_
  );


  buf

  (
    g447_p_spl_,
    g447_p
  );


  buf

  (
    g447_p_spl_0,
    g447_p_spl_
  );


  buf

  (
    g447_p_spl_1,
    g447_p_spl_
  );


  buf

  (
    g447_n_spl_,
    g447_n
  );


  buf

  (
    g447_n_spl_0,
    g447_n_spl_
  );


  buf

  (
    g447_n_spl_1,
    g447_n_spl_
  );


  buf

  (
    g448_n_spl_,
    g448_n
  );


  buf

  (
    g448_p_spl_,
    g448_p
  );


  buf

  (
    G125_n_spl_,
    G125_n
  );


  buf

  (
    g451_n_spl_,
    g451_n
  );


  buf

  (
    g451_n_spl_0,
    g451_n_spl_
  );


  buf

  (
    g451_n_spl_1,
    g451_n_spl_
  );


  buf

  (
    g451_p_spl_,
    g451_p
  );


  buf

  (
    g451_p_spl_0,
    g451_p_spl_
  );


  buf

  (
    g451_p_spl_1,
    g451_p_spl_
  );


  buf

  (
    g452_n_spl_,
    g452_n
  );


  buf

  (
    g452_n_spl_0,
    g452_n_spl_
  );


  buf

  (
    g452_p_spl_,
    g452_p
  );


  buf

  (
    g452_p_spl_0,
    g452_p_spl_
  );


  buf

  (
    g450_p_spl_,
    g450_p
  );


  buf

  (
    g450_p_spl_0,
    g450_p_spl_
  );


  buf

  (
    g450_p_spl_1,
    g450_p_spl_
  );


  buf

  (
    g454_p_spl_,
    g454_p
  );


  buf

  (
    g454_p_spl_0,
    g454_p_spl_
  );


  buf

  (
    g454_p_spl_1,
    g454_p_spl_
  );


  buf

  (
    g450_n_spl_,
    g450_n
  );


  buf

  (
    g450_n_spl_0,
    g450_n_spl_
  );


  buf

  (
    g450_n_spl_1,
    g450_n_spl_
  );


  buf

  (
    g454_n_spl_,
    g454_n
  );


  buf

  (
    g454_n_spl_0,
    g454_n_spl_
  );


  buf

  (
    g454_n_spl_00,
    g454_n_spl_0
  );


  buf

  (
    g454_n_spl_1,
    g454_n_spl_
  );


  buf

  (
    G129_n_spl_,
    G129_n
  );


  buf

  (
    g458_p_spl_,
    g458_p
  );


  buf

  (
    g458_p_spl_0,
    g458_p_spl_
  );


  buf

  (
    g458_p_spl_1,
    g458_p_spl_
  );


  buf

  (
    g458_n_spl_,
    g458_n
  );


  buf

  (
    g458_n_spl_0,
    g458_n_spl_
  );


  buf

  (
    g458_n_spl_1,
    g458_n_spl_
  );


  buf

  (
    g459_n_spl_,
    g459_n
  );


  buf

  (
    g459_n_spl_0,
    g459_n_spl_
  );


  buf

  (
    g459_p_spl_,
    g459_p
  );


  buf

  (
    g459_p_spl_0,
    g459_p_spl_
  );


  buf

  (
    G131_n_spl_,
    G131_n
  );


  buf

  (
    g461_p_spl_,
    g461_p
  );


  buf

  (
    g461_p_spl_0,
    g461_p_spl_
  );


  buf

  (
    g464_n_spl_,
    g464_n
  );


  buf

  (
    g464_n_spl_0,
    g464_n_spl_
  );


  buf

  (
    g464_n_spl_00,
    g464_n_spl_0
  );


  buf

  (
    g464_n_spl_01,
    g464_n_spl_0
  );


  buf

  (
    g464_n_spl_1,
    g464_n_spl_
  );


  buf

  (
    g464_n_spl_10,
    g464_n_spl_1
  );


  buf

  (
    g461_n_spl_,
    g461_n
  );


  buf

  (
    g461_n_spl_0,
    g461_n_spl_
  );


  buf

  (
    g464_p_spl_,
    g464_p
  );


  buf

  (
    g464_p_spl_0,
    g464_p_spl_
  );


  buf

  (
    g464_p_spl_00,
    g464_p_spl_0
  );


  buf

  (
    g464_p_spl_01,
    g464_p_spl_0
  );


  buf

  (
    g464_p_spl_1,
    g464_p_spl_
  );


  buf

  (
    g464_p_spl_10,
    g464_p_spl_1
  );


  buf

  (
    G127_n_spl_,
    G127_n
  );


  buf

  (
    g468_p_spl_,
    g468_p
  );


  buf

  (
    g468_p_spl_0,
    g468_p_spl_
  );


  buf

  (
    g468_p_spl_1,
    g468_p_spl_
  );


  buf

  (
    g468_n_spl_,
    g468_n
  );


  buf

  (
    g468_n_spl_0,
    g468_n_spl_
  );


  buf

  (
    g468_n_spl_1,
    g468_n_spl_
  );


  buf

  (
    g469_n_spl_,
    g469_n
  );


  buf

  (
    g469_n_spl_0,
    g469_n_spl_
  );


  buf

  (
    g469_p_spl_,
    g469_p
  );


  buf

  (
    g469_p_spl_0,
    g469_p_spl_
  );


  buf

  (
    g465_p_spl_,
    g465_p
  );


  buf

  (
    g465_p_spl_0,
    g465_p_spl_
  );


  buf

  (
    g471_p_spl_,
    g471_p
  );


  buf

  (
    g471_p_spl_0,
    g471_p_spl_
  );


  buf

  (
    g471_p_spl_1,
    g471_p_spl_
  );


  buf

  (
    g465_n_spl_,
    g465_n
  );


  buf

  (
    g465_n_spl_0,
    g465_n_spl_
  );


  buf

  (
    g471_n_spl_,
    g471_n
  );


  buf

  (
    g471_n_spl_0,
    g471_n_spl_
  );


  buf

  (
    g471_n_spl_00,
    g471_n_spl_0
  );


  buf

  (
    g471_n_spl_1,
    g471_n_spl_
  );


  buf

  (
    g455_p_spl_,
    g455_p
  );


  buf

  (
    g472_p_spl_,
    g472_p
  );


  buf

  (
    g455_n_spl_,
    g455_n
  );


  buf

  (
    g472_n_spl_,
    g472_n
  );


  buf

  (
    G114_n_spl_,
    G114_n
  );


  buf

  (
    G114_n_spl_0,
    G114_n_spl_
  );


  buf

  (
    G114_p_spl_,
    G114_p
  );


  buf

  (
    g476_n_spl_,
    g476_n
  );


  buf

  (
    g476_n_spl_0,
    g476_n_spl_
  );


  buf

  (
    g476_n_spl_1,
    g476_n_spl_
  );


  buf

  (
    g479_n_spl_,
    g479_n
  );


  buf

  (
    g479_n_spl_0,
    g479_n_spl_
  );


  buf

  (
    g479_n_spl_00,
    g479_n_spl_0
  );


  buf

  (
    g479_n_spl_01,
    g479_n_spl_0
  );


  buf

  (
    g479_n_spl_1,
    g479_n_spl_
  );


  buf

  (
    g479_n_spl_10,
    g479_n_spl_1
  );


  buf

  (
    g476_p_spl_,
    g476_p
  );


  buf

  (
    g476_p_spl_0,
    g476_p_spl_
  );


  buf

  (
    g476_p_spl_00,
    g476_p_spl_0
  );


  buf

  (
    g476_p_spl_1,
    g476_p_spl_
  );


  buf

  (
    g479_p_spl_,
    g479_p
  );


  buf

  (
    g479_p_spl_0,
    g479_p_spl_
  );


  buf

  (
    g479_p_spl_00,
    g479_p_spl_0
  );


  buf

  (
    g479_p_spl_01,
    g479_p_spl_0
  );


  buf

  (
    g479_p_spl_1,
    g479_p_spl_
  );


  buf

  (
    g479_p_spl_10,
    g479_p_spl_1
  );


  buf

  (
    g473_p_spl_,
    g473_p
  );


  buf

  (
    g480_p_spl_,
    g480_p
  );


  buf

  (
    g480_p_spl_0,
    g480_p_spl_
  );


  buf

  (
    g444_p_spl_,
    g444_p
  );


  buf

  (
    g444_p_spl_0,
    g444_p_spl_
  );


  buf

  (
    g485_p_spl_,
    g485_p
  );


  buf

  (
    g488_n_spl_,
    g488_n
  );


  buf

  (
    g485_n_spl_,
    g485_n
  );


  buf

  (
    g488_p_spl_,
    g488_p
  );


  buf

  (
    G132_n_spl_,
    G132_n
  );


  buf

  (
    G132_n_spl_0,
    G132_n_spl_
  );


  buf

  (
    G132_p_spl_,
    G132_p
  );


  buf

  (
    G132_p_spl_0,
    G132_p_spl_
  );


  buf

  (
    g494_n_spl_,
    g494_n
  );


  buf

  (
    g494_p_spl_,
    g494_p
  );


  buf

  (
    g497_n_spl_,
    g497_n
  );


  buf

  (
    g500_n_spl_,
    g500_n
  );


  buf

  (
    g497_p_spl_,
    g497_p
  );


  buf

  (
    g500_p_spl_,
    g500_p
  );


  buf

  (
    g509_p_spl_,
    g509_p
  );


  buf

  (
    g512_n_spl_,
    g512_n
  );


  buf

  (
    g509_n_spl_,
    g509_n
  );


  buf

  (
    g512_p_spl_,
    g512_p
  );


  buf

  (
    G111_n_spl_,
    G111_n
  );


  buf

  (
    G111_n_spl_0,
    G111_n_spl_
  );


  buf

  (
    G111_p_spl_,
    G111_p
  );


  buf

  (
    G111_p_spl_0,
    G111_p_spl_
  );


  buf

  (
    g518_n_spl_,
    g518_n
  );


  buf

  (
    g521_n_spl_,
    g521_n
  );


  buf

  (
    g518_p_spl_,
    g518_p
  );


  buf

  (
    g521_p_spl_,
    g521_p
  );


  buf

  (
    g524_n_spl_,
    g524_n
  );


  buf

  (
    g527_n_spl_,
    g527_n
  );


  buf

  (
    g524_p_spl_,
    g524_p
  );


  buf

  (
    g527_p_spl_,
    g527_p
  );


  buf

  (
    g535_n_spl_,
    g535_n
  );


  buf

  (
    g535_n_spl_0,
    g535_n_spl_
  );


  buf

  (
    g535_n_spl_1,
    g535_n_spl_
  );


  buf

  (
    g535_p_spl_,
    g535_p
  );


  buf

  (
    g535_p_spl_0,
    g535_p_spl_
  );


  buf

  (
    g535_p_spl_1,
    g535_p_spl_
  );


  buf

  (
    g537_n_spl_,
    g537_n
  );


  buf

  (
    g537_n_spl_0,
    g537_n_spl_
  );


  buf

  (
    g537_n_spl_00,
    g537_n_spl_0
  );


  buf

  (
    g537_n_spl_1,
    g537_n_spl_
  );


  buf

  (
    g537_p_spl_,
    g537_p
  );


  buf

  (
    g537_p_spl_0,
    g537_p_spl_
  );


  buf

  (
    g537_p_spl_00,
    g537_p_spl_0
  );


  buf

  (
    g537_p_spl_1,
    g537_p_spl_
  );


  buf

  (
    g539_n_spl_,
    g539_n
  );


  buf

  (
    g539_n_spl_0,
    g539_n_spl_
  );


  buf

  (
    g539_n_spl_1,
    g539_n_spl_
  );


  buf

  (
    g539_p_spl_,
    g539_p
  );


  buf

  (
    g539_p_spl_0,
    g539_p_spl_
  );


  buf

  (
    g539_p_spl_1,
    g539_p_spl_
  );


  buf

  (
    g541_p_spl_,
    g541_p
  );


  buf

  (
    g541_p_spl_0,
    g541_p_spl_
  );


  buf

  (
    g541_p_spl_00,
    g541_p_spl_0
  );


  buf

  (
    g541_p_spl_1,
    g541_p_spl_
  );


  buf

  (
    g544_n_spl_,
    g544_n
  );


  buf

  (
    g544_n_spl_0,
    g544_n_spl_
  );


  buf

  (
    g544_n_spl_1,
    g544_n_spl_
  );


  buf

  (
    g544_p_spl_,
    g544_p
  );


  buf

  (
    g544_p_spl_0,
    g544_p_spl_
  );


  buf

  (
    g544_p_spl_1,
    g544_p_spl_
  );


  buf

  (
    g545_n_spl_,
    g545_n
  );


  buf

  (
    g545_p_spl_,
    g545_p
  );


  buf

  (
    g546_p_spl_,
    g546_p
  );


  buf

  (
    g546_p_spl_0,
    g546_p_spl_
  );


  buf

  (
    g546_p_spl_1,
    g546_p_spl_
  );


  buf

  (
    G177_p_spl_,
    G177_p
  );


  buf

  (
    G177_p_spl_0,
    G177_p_spl_
  );


  buf

  (
    G177_p_spl_00,
    G177_p_spl_0
  );


  buf

  (
    G177_p_spl_000,
    G177_p_spl_00
  );


  buf

  (
    G177_p_spl_0000,
    G177_p_spl_000
  );


  buf

  (
    G177_p_spl_0001,
    G177_p_spl_000
  );


  buf

  (
    G177_p_spl_001,
    G177_p_spl_00
  );


  buf

  (
    G177_p_spl_0010,
    G177_p_spl_001
  );


  buf

  (
    G177_p_spl_0011,
    G177_p_spl_001
  );


  buf

  (
    G177_p_spl_01,
    G177_p_spl_0
  );


  buf

  (
    G177_p_spl_010,
    G177_p_spl_01
  );


  buf

  (
    G177_p_spl_0100,
    G177_p_spl_010
  );


  buf

  (
    G177_p_spl_0101,
    G177_p_spl_010
  );


  buf

  (
    G177_p_spl_011,
    G177_p_spl_01
  );


  buf

  (
    G177_p_spl_0110,
    G177_p_spl_011
  );


  buf

  (
    G177_p_spl_0111,
    G177_p_spl_011
  );


  buf

  (
    G177_p_spl_1,
    G177_p_spl_
  );


  buf

  (
    G177_p_spl_10,
    G177_p_spl_1
  );


  buf

  (
    G177_p_spl_100,
    G177_p_spl_10
  );


  buf

  (
    G177_p_spl_1000,
    G177_p_spl_100
  );


  buf

  (
    G177_p_spl_1001,
    G177_p_spl_100
  );


  buf

  (
    G177_p_spl_101,
    G177_p_spl_10
  );


  buf

  (
    G177_p_spl_11,
    G177_p_spl_1
  );


  buf

  (
    G177_p_spl_110,
    G177_p_spl_11
  );


  buf

  (
    G177_p_spl_111,
    G177_p_spl_11
  );


  buf

  (
    g553_p_spl_,
    g553_p
  );


  buf

  (
    G176_p_spl_,
    G176_p
  );


  buf

  (
    G176_p_spl_0,
    G176_p_spl_
  );


  buf

  (
    G176_p_spl_00,
    G176_p_spl_0
  );


  buf

  (
    G176_p_spl_000,
    G176_p_spl_00
  );


  buf

  (
    G176_p_spl_0000,
    G176_p_spl_000
  );


  buf

  (
    G176_p_spl_00000,
    G176_p_spl_0000
  );


  buf

  (
    G176_p_spl_00001,
    G176_p_spl_0000
  );


  buf

  (
    G176_p_spl_0001,
    G176_p_spl_000
  );


  buf

  (
    G176_p_spl_001,
    G176_p_spl_00
  );


  buf

  (
    G176_p_spl_0010,
    G176_p_spl_001
  );


  buf

  (
    G176_p_spl_0011,
    G176_p_spl_001
  );


  buf

  (
    G176_p_spl_01,
    G176_p_spl_0
  );


  buf

  (
    G176_p_spl_010,
    G176_p_spl_01
  );


  buf

  (
    G176_p_spl_0100,
    G176_p_spl_010
  );


  buf

  (
    G176_p_spl_0101,
    G176_p_spl_010
  );


  buf

  (
    G176_p_spl_011,
    G176_p_spl_01
  );


  buf

  (
    G176_p_spl_0110,
    G176_p_spl_011
  );


  buf

  (
    G176_p_spl_0111,
    G176_p_spl_011
  );


  buf

  (
    G176_p_spl_1,
    G176_p_spl_
  );


  buf

  (
    G176_p_spl_10,
    G176_p_spl_1
  );


  buf

  (
    G176_p_spl_100,
    G176_p_spl_10
  );


  buf

  (
    G176_p_spl_1000,
    G176_p_spl_100
  );


  buf

  (
    G176_p_spl_1001,
    G176_p_spl_100
  );


  buf

  (
    G176_p_spl_101,
    G176_p_spl_10
  );


  buf

  (
    G176_p_spl_1010,
    G176_p_spl_101
  );


  buf

  (
    G176_p_spl_1011,
    G176_p_spl_101
  );


  buf

  (
    G176_p_spl_11,
    G176_p_spl_1
  );


  buf

  (
    G176_p_spl_110,
    G176_p_spl_11
  );


  buf

  (
    G176_p_spl_1100,
    G176_p_spl_110
  );


  buf

  (
    G176_p_spl_1101,
    G176_p_spl_110
  );


  buf

  (
    G176_p_spl_111,
    G176_p_spl_11
  );


  buf

  (
    G176_p_spl_1110,
    G176_p_spl_111
  );


  buf

  (
    G176_p_spl_1111,
    G176_p_spl_111
  );


  buf

  (
    G177_n_spl_,
    G177_n
  );


  buf

  (
    G177_n_spl_0,
    G177_n_spl_
  );


  buf

  (
    G177_n_spl_00,
    G177_n_spl_0
  );


  buf

  (
    G177_n_spl_000,
    G177_n_spl_00
  );


  buf

  (
    G177_n_spl_0000,
    G177_n_spl_000
  );


  buf

  (
    G177_n_spl_0001,
    G177_n_spl_000
  );


  buf

  (
    G177_n_spl_001,
    G177_n_spl_00
  );


  buf

  (
    G177_n_spl_0010,
    G177_n_spl_001
  );


  buf

  (
    G177_n_spl_0011,
    G177_n_spl_001
  );


  buf

  (
    G177_n_spl_01,
    G177_n_spl_0
  );


  buf

  (
    G177_n_spl_010,
    G177_n_spl_01
  );


  buf

  (
    G177_n_spl_011,
    G177_n_spl_01
  );


  buf

  (
    G177_n_spl_1,
    G177_n_spl_
  );


  buf

  (
    G177_n_spl_10,
    G177_n_spl_1
  );


  buf

  (
    G177_n_spl_100,
    G177_n_spl_10
  );


  buf

  (
    G177_n_spl_101,
    G177_n_spl_10
  );


  buf

  (
    G177_n_spl_11,
    G177_n_spl_1
  );


  buf

  (
    G177_n_spl_110,
    G177_n_spl_11
  );


  buf

  (
    G177_n_spl_111,
    G177_n_spl_11
  );


  buf

  (
    G176_n_spl_,
    G176_n
  );


  buf

  (
    G176_n_spl_0,
    G176_n_spl_
  );


  buf

  (
    G176_n_spl_00,
    G176_n_spl_0
  );


  buf

  (
    G176_n_spl_000,
    G176_n_spl_00
  );


  buf

  (
    G176_n_spl_0000,
    G176_n_spl_000
  );


  buf

  (
    G176_n_spl_0001,
    G176_n_spl_000
  );


  buf

  (
    G176_n_spl_001,
    G176_n_spl_00
  );


  buf

  (
    G176_n_spl_0010,
    G176_n_spl_001
  );


  buf

  (
    G176_n_spl_0011,
    G176_n_spl_001
  );


  buf

  (
    G176_n_spl_01,
    G176_n_spl_0
  );


  buf

  (
    G176_n_spl_010,
    G176_n_spl_01
  );


  buf

  (
    G176_n_spl_0100,
    G176_n_spl_010
  );


  buf

  (
    G176_n_spl_0101,
    G176_n_spl_010
  );


  buf

  (
    G176_n_spl_011,
    G176_n_spl_01
  );


  buf

  (
    G176_n_spl_1,
    G176_n_spl_
  );


  buf

  (
    G176_n_spl_10,
    G176_n_spl_1
  );


  buf

  (
    G176_n_spl_100,
    G176_n_spl_10
  );


  buf

  (
    G176_n_spl_101,
    G176_n_spl_10
  );


  buf

  (
    G176_n_spl_11,
    G176_n_spl_1
  );


  buf

  (
    G176_n_spl_110,
    G176_n_spl_11
  );


  buf

  (
    G176_n_spl_111,
    G176_n_spl_11
  );


  buf

  (
    g562_n_spl_,
    g562_n
  );


  buf

  (
    g562_n_spl_0,
    g562_n_spl_
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G2_p_spl_0,
    G2_p_spl_
  );


  buf

  (
    G2_p_spl_1,
    G2_p_spl_
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G2_n_spl_0,
    G2_n_spl_
  );


  buf

  (
    g570_n_spl_,
    g570_n
  );


  buf

  (
    g572_p_spl_,
    g572_p
  );


  buf

  (
    G22_p_spl_,
    G22_p
  );


  buf

  (
    G173_n_spl_,
    G173_n
  );


  buf

  (
    G173_n_spl_0,
    G173_n_spl_
  );


  buf

  (
    G173_n_spl_00,
    G173_n_spl_0
  );


  buf

  (
    G173_n_spl_000,
    G173_n_spl_00
  );


  buf

  (
    G173_n_spl_0000,
    G173_n_spl_000
  );


  buf

  (
    G173_n_spl_0001,
    G173_n_spl_000
  );


  buf

  (
    G173_n_spl_001,
    G173_n_spl_00
  );


  buf

  (
    G173_n_spl_0010,
    G173_n_spl_001
  );


  buf

  (
    G173_n_spl_0011,
    G173_n_spl_001
  );


  buf

  (
    G173_n_spl_01,
    G173_n_spl_0
  );


  buf

  (
    G173_n_spl_010,
    G173_n_spl_01
  );


  buf

  (
    G173_n_spl_011,
    G173_n_spl_01
  );


  buf

  (
    G173_n_spl_1,
    G173_n_spl_
  );


  buf

  (
    G173_n_spl_10,
    G173_n_spl_1
  );


  buf

  (
    G173_n_spl_100,
    G173_n_spl_10
  );


  buf

  (
    G173_n_spl_101,
    G173_n_spl_10
  );


  buf

  (
    G173_n_spl_11,
    G173_n_spl_1
  );


  buf

  (
    G173_n_spl_110,
    G173_n_spl_11
  );


  buf

  (
    G173_n_spl_111,
    G173_n_spl_11
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G173_p_spl_,
    G173_p
  );


  buf

  (
    G173_p_spl_0,
    G173_p_spl_
  );


  buf

  (
    G173_p_spl_00,
    G173_p_spl_0
  );


  buf

  (
    G173_p_spl_000,
    G173_p_spl_00
  );


  buf

  (
    G173_p_spl_0000,
    G173_p_spl_000
  );


  buf

  (
    G173_p_spl_0001,
    G173_p_spl_000
  );


  buf

  (
    G173_p_spl_001,
    G173_p_spl_00
  );


  buf

  (
    G173_p_spl_0010,
    G173_p_spl_001
  );


  buf

  (
    G173_p_spl_0011,
    G173_p_spl_001
  );


  buf

  (
    G173_p_spl_01,
    G173_p_spl_0
  );


  buf

  (
    G173_p_spl_010,
    G173_p_spl_01
  );


  buf

  (
    G173_p_spl_011,
    G173_p_spl_01
  );


  buf

  (
    G173_p_spl_1,
    G173_p_spl_
  );


  buf

  (
    G173_p_spl_10,
    G173_p_spl_1
  );


  buf

  (
    G173_p_spl_100,
    G173_p_spl_10
  );


  buf

  (
    G173_p_spl_101,
    G173_p_spl_10
  );


  buf

  (
    G173_p_spl_11,
    G173_p_spl_1
  );


  buf

  (
    G173_p_spl_110,
    G173_p_spl_11
  );


  buf

  (
    G173_p_spl_111,
    G173_p_spl_11
  );


  buf

  (
    G172_n_spl_,
    G172_n
  );


  buf

  (
    G172_n_spl_0,
    G172_n_spl_
  );


  buf

  (
    G172_n_spl_00,
    G172_n_spl_0
  );


  buf

  (
    G172_n_spl_000,
    G172_n_spl_00
  );


  buf

  (
    G172_n_spl_001,
    G172_n_spl_00
  );


  buf

  (
    G172_n_spl_01,
    G172_n_spl_0
  );


  buf

  (
    G172_n_spl_1,
    G172_n_spl_
  );


  buf

  (
    G172_n_spl_10,
    G172_n_spl_1
  );


  buf

  (
    G172_n_spl_11,
    G172_n_spl_1
  );


  buf

  (
    g579_p_spl_,
    g579_p
  );


  buf

  (
    g579_p_spl_0,
    g579_p_spl_
  );


  buf

  (
    g579_p_spl_00,
    g579_p_spl_0
  );


  buf

  (
    g579_p_spl_1,
    g579_p_spl_
  );


  buf

  (
    g560_p_spl_,
    g560_p
  );


  buf

  (
    g560_p_spl_0,
    g560_p_spl_
  );


  buf

  (
    g560_p_spl_00,
    g560_p_spl_0
  );


  buf

  (
    g560_p_spl_1,
    g560_p_spl_
  );


  buf

  (
    G172_p_spl_,
    G172_p
  );


  buf

  (
    G172_p_spl_0,
    G172_p_spl_
  );


  buf

  (
    G172_p_spl_00,
    G172_p_spl_0
  );


  buf

  (
    G172_p_spl_000,
    G172_p_spl_00
  );


  buf

  (
    G172_p_spl_001,
    G172_p_spl_00
  );


  buf

  (
    G172_p_spl_01,
    G172_p_spl_0
  );


  buf

  (
    G172_p_spl_1,
    G172_p_spl_
  );


  buf

  (
    G172_p_spl_10,
    G172_p_spl_1
  );


  buf

  (
    G172_p_spl_11,
    G172_p_spl_1
  );


  buf

  (
    g594_n_spl_,
    g594_n
  );


  buf

  (
    g594_p_spl_,
    g594_p
  );


  buf

  (
    g595_n_spl_,
    g595_n
  );


  buf

  (
    g596_n_spl_,
    g596_n
  );


  buf

  (
    g596_n_spl_0,
    g596_n_spl_
  );


  buf

  (
    g596_p_spl_,
    g596_p
  );


  buf

  (
    g596_p_spl_0,
    g596_p_spl_
  );


  buf

  (
    g596_p_spl_1,
    g596_p_spl_
  );


  buf

  (
    g597_p_spl_,
    g597_p
  );


  buf

  (
    g598_p_spl_,
    g598_p
  );


  buf

  (
    g598_p_spl_0,
    g598_p_spl_
  );


  buf

  (
    g598_n_spl_,
    g598_n
  );


  buf

  (
    g598_n_spl_0,
    g598_n_spl_
  );


  buf

  (
    g601_p_spl_,
    g601_p
  );


  buf

  (
    g610_n_spl_,
    g610_n
  );


  buf

  (
    g617_p_spl_,
    g617_p
  );


  buf

  (
    g617_p_spl_0,
    g617_p_spl_
  );


  buf

  (
    g619_n_spl_,
    g619_n
  );


  buf

  (
    G174_n_spl_,
    G174_n
  );


  buf

  (
    G174_n_spl_0,
    G174_n_spl_
  );


  buf

  (
    G174_n_spl_00,
    G174_n_spl_0
  );


  buf

  (
    G174_n_spl_000,
    G174_n_spl_00
  );


  buf

  (
    G174_n_spl_0000,
    G174_n_spl_000
  );


  buf

  (
    G174_n_spl_0001,
    G174_n_spl_000
  );


  buf

  (
    G174_n_spl_001,
    G174_n_spl_00
  );


  buf

  (
    G174_n_spl_0010,
    G174_n_spl_001
  );


  buf

  (
    G174_n_spl_0011,
    G174_n_spl_001
  );


  buf

  (
    G174_n_spl_01,
    G174_n_spl_0
  );


  buf

  (
    G174_n_spl_010,
    G174_n_spl_01
  );


  buf

  (
    G174_n_spl_011,
    G174_n_spl_01
  );


  buf

  (
    G174_n_spl_1,
    G174_n_spl_
  );


  buf

  (
    G174_n_spl_10,
    G174_n_spl_1
  );


  buf

  (
    G174_n_spl_100,
    G174_n_spl_10
  );


  buf

  (
    G174_n_spl_101,
    G174_n_spl_10
  );


  buf

  (
    G174_n_spl_11,
    G174_n_spl_1
  );


  buf

  (
    G174_n_spl_110,
    G174_n_spl_11
  );


  buf

  (
    G174_n_spl_111,
    G174_n_spl_11
  );


  buf

  (
    G174_p_spl_,
    G174_p
  );


  buf

  (
    G174_p_spl_0,
    G174_p_spl_
  );


  buf

  (
    G174_p_spl_00,
    G174_p_spl_0
  );


  buf

  (
    G174_p_spl_000,
    G174_p_spl_00
  );


  buf

  (
    G174_p_spl_0000,
    G174_p_spl_000
  );


  buf

  (
    G174_p_spl_0001,
    G174_p_spl_000
  );


  buf

  (
    G174_p_spl_001,
    G174_p_spl_00
  );


  buf

  (
    G174_p_spl_0010,
    G174_p_spl_001
  );


  buf

  (
    G174_p_spl_0011,
    G174_p_spl_001
  );


  buf

  (
    G174_p_spl_01,
    G174_p_spl_0
  );


  buf

  (
    G174_p_spl_010,
    G174_p_spl_01
  );


  buf

  (
    G174_p_spl_011,
    G174_p_spl_01
  );


  buf

  (
    G174_p_spl_1,
    G174_p_spl_
  );


  buf

  (
    G174_p_spl_10,
    G174_p_spl_1
  );


  buf

  (
    G174_p_spl_100,
    G174_p_spl_10
  );


  buf

  (
    G174_p_spl_101,
    G174_p_spl_10
  );


  buf

  (
    G174_p_spl_11,
    G174_p_spl_1
  );


  buf

  (
    G174_p_spl_110,
    G174_p_spl_11
  );


  buf

  (
    G174_p_spl_111,
    G174_p_spl_11
  );


  buf

  (
    G175_n_spl_,
    G175_n
  );


  buf

  (
    G175_n_spl_0,
    G175_n_spl_
  );


  buf

  (
    G175_n_spl_00,
    G175_n_spl_0
  );


  buf

  (
    G175_n_spl_000,
    G175_n_spl_00
  );


  buf

  (
    G175_n_spl_001,
    G175_n_spl_00
  );


  buf

  (
    G175_n_spl_01,
    G175_n_spl_0
  );


  buf

  (
    G175_n_spl_1,
    G175_n_spl_
  );


  buf

  (
    G175_n_spl_10,
    G175_n_spl_1
  );


  buf

  (
    G175_n_spl_11,
    G175_n_spl_1
  );


  buf

  (
    G175_p_spl_,
    G175_p
  );


  buf

  (
    G175_p_spl_0,
    G175_p_spl_
  );


  buf

  (
    G175_p_spl_00,
    G175_p_spl_0
  );


  buf

  (
    G175_p_spl_000,
    G175_p_spl_00
  );


  buf

  (
    G175_p_spl_001,
    G175_p_spl_00
  );


  buf

  (
    G175_p_spl_01,
    G175_p_spl_0
  );


  buf

  (
    G175_p_spl_1,
    G175_p_spl_
  );


  buf

  (
    G175_p_spl_10,
    G175_p_spl_1
  );


  buf

  (
    G175_p_spl_11,
    G175_p_spl_1
  );


  buf

  (
    g638_p_spl_,
    g638_p
  );


  buf

  (
    g639_p_spl_,
    g639_p
  );


  buf

  (
    g643_n_spl_,
    g643_n
  );


  buf

  (
    g652_n_spl_,
    g652_n
  );


  buf

  (
    g659_p_spl_,
    g659_p
  );


  buf

  (
    g660_p_spl_,
    g660_p
  );


  buf

  (
    g664_n_spl_,
    g664_n
  );


  buf

  (
    g673_n_spl_,
    g673_n
  );


  buf

  (
    g581_n_spl_,
    g581_n
  );


  buf

  (
    g581_n_spl_0,
    g581_n_spl_
  );


  buf

  (
    g581_n_spl_00,
    g581_n_spl_0
  );


  buf

  (
    g581_n_spl_01,
    g581_n_spl_0
  );


  buf

  (
    g581_n_spl_1,
    g581_n_spl_
  );


  buf

  (
    g581_n_spl_10,
    g581_n_spl_1
  );


  buf

  (
    g581_n_spl_11,
    g581_n_spl_1
  );


  buf

  (
    g681_p_spl_,
    g681_p
  );


  buf

  (
    g581_p_spl_,
    g581_p
  );


  buf

  (
    g581_p_spl_0,
    g581_p_spl_
  );


  buf

  (
    g581_p_spl_00,
    g581_p_spl_0
  );


  buf

  (
    g581_p_spl_01,
    g581_p_spl_0
  );


  buf

  (
    g581_p_spl_1,
    g581_p_spl_
  );


  buf

  (
    g681_n_spl_,
    g681_n
  );


  buf

  (
    g687_n_spl_,
    g687_n
  );


  buf

  (
    g687_p_spl_,
    g687_p
  );


  buf

  (
    g693_n_spl_,
    g693_n
  );


  buf

  (
    g696_n_spl_,
    g696_n
  );


  buf

  (
    g693_p_spl_,
    g693_p
  );


  buf

  (
    g696_p_spl_,
    g696_p
  );


  buf

  (
    g690_p_spl_,
    g690_p
  );


  buf

  (
    g699_n_spl_,
    g699_n
  );


  buf

  (
    g690_n_spl_,
    g690_n
  );


  buf

  (
    g699_p_spl_,
    g699_p
  );


  buf

  (
    g708_p_spl_,
    g708_p
  );


  buf

  (
    g711_n_spl_,
    g711_n
  );


  buf

  (
    g708_n_spl_,
    g708_n
  );


  buf

  (
    g711_p_spl_,
    g711_p
  );


  buf

  (
    g717_n_spl_,
    g717_n
  );


  buf

  (
    g717_p_spl_,
    g717_p
  );


  buf

  (
    g720_p_spl_,
    g720_p
  );


  buf

  (
    g723_n_spl_,
    g723_n
  );


  buf

  (
    g720_n_spl_,
    g720_n
  );


  buf

  (
    g723_p_spl_,
    g723_p
  );


  buf

  (
    g726_n_spl_,
    g726_n
  );


  buf

  (
    g729_n_spl_,
    g729_n
  );


  buf

  (
    g726_p_spl_,
    g726_p
  );


  buf

  (
    g729_p_spl_,
    g729_p
  );


  buf

  (
    g430_p_spl_,
    g430_p
  );


  buf

  (
    g430_p_spl_0,
    g430_p_spl_
  );


  buf

  (
    g541_n_spl_,
    g541_n
  );


  buf

  (
    g541_n_spl_0,
    g541_n_spl_
  );


  buf

  (
    g541_n_spl_1,
    g541_n_spl_
  );


  buf

  (
    g737_p_spl_,
    g737_p
  );


  buf

  (
    g737_p_spl_0,
    g737_p_spl_
  );


  buf

  (
    g737_p_spl_00,
    g737_p_spl_0
  );


  buf

  (
    g737_p_spl_1,
    g737_p_spl_
  );


  buf

  (
    g737_n_spl_,
    g737_n
  );


  buf

  (
    g737_n_spl_0,
    g737_n_spl_
  );


  buf

  (
    g737_n_spl_00,
    g737_n_spl_0
  );


  buf

  (
    g737_n_spl_1,
    g737_n_spl_
  );


  buf

  (
    g743_p_spl_,
    g743_p
  );


  buf

  (
    g747_p_spl_,
    g747_p
  );


  buf

  (
    g389_p_spl_,
    g389_p
  );


  buf

  (
    g546_n_spl_,
    g546_n
  );


  buf

  (
    g546_n_spl_0,
    g546_n_spl_
  );


  buf

  (
    g395_p_spl_,
    g395_p
  );


  buf

  (
    g395_p_spl_0,
    g395_p_spl_
  );


  buf

  (
    g395_p_spl_00,
    g395_p_spl_0
  );


  buf

  (
    g395_p_spl_1,
    g395_p_spl_
  );


  buf

  (
    g755_p_spl_,
    g755_p
  );


  buf

  (
    g760_p_spl_,
    g760_p
  );


  buf

  (
    g774_p_spl_,
    g774_p
  );


  buf

  (
    g774_p_spl_0,
    g774_p_spl_
  );


  buf

  (
    g774_p_spl_00,
    g774_p_spl_0
  );


  buf

  (
    g774_p_spl_01,
    g774_p_spl_0
  );


  buf

  (
    g774_p_spl_1,
    g774_p_spl_
  );


  buf

  (
    g774_n_spl_,
    g774_n
  );


  buf

  (
    g774_n_spl_0,
    g774_n_spl_
  );


  buf

  (
    g774_n_spl_00,
    g774_n_spl_0
  );


  buf

  (
    g774_n_spl_01,
    g774_n_spl_0
  );


  buf

  (
    g774_n_spl_1,
    g774_n_spl_
  );


  buf

  (
    g777_p_spl_,
    g777_p
  );


  buf

  (
    g444_n_spl_,
    g444_n
  );


  buf

  (
    g780_p_spl_,
    g780_p
  );


  buf

  (
    g780_p_spl_0,
    g780_p_spl_
  );


  buf

  (
    g780_p_spl_1,
    g780_p_spl_
  );


  buf

  (
    g780_n_spl_,
    g780_n
  );


  buf

  (
    g780_n_spl_0,
    g780_n_spl_
  );


  buf

  (
    g780_n_spl_1,
    g780_n_spl_
  );


  buf

  (
    g785_p_spl_,
    g785_p
  );


  buf

  (
    g791_p_spl_,
    g791_p
  );


  buf

  (
    G81_p_spl_,
    G81_p
  );


  buf

  (
    G158_n_spl_,
    G158_n
  );


  buf

  (
    G158_n_spl_0,
    G158_n_spl_
  );


  buf

  (
    G158_n_spl_00,
    G158_n_spl_0
  );


  buf

  (
    G158_n_spl_000,
    G158_n_spl_00
  );


  buf

  (
    G158_n_spl_0000,
    G158_n_spl_000
  );


  buf

  (
    G158_n_spl_0001,
    G158_n_spl_000
  );


  buf

  (
    G158_n_spl_001,
    G158_n_spl_00
  );


  buf

  (
    G158_n_spl_0010,
    G158_n_spl_001
  );


  buf

  (
    G158_n_spl_0011,
    G158_n_spl_001
  );


  buf

  (
    G158_n_spl_01,
    G158_n_spl_0
  );


  buf

  (
    G158_n_spl_010,
    G158_n_spl_01
  );


  buf

  (
    G158_n_spl_011,
    G158_n_spl_01
  );


  buf

  (
    G158_n_spl_1,
    G158_n_spl_
  );


  buf

  (
    G158_n_spl_10,
    G158_n_spl_1
  );


  buf

  (
    G158_n_spl_100,
    G158_n_spl_10
  );


  buf

  (
    G158_n_spl_101,
    G158_n_spl_10
  );


  buf

  (
    G158_n_spl_11,
    G158_n_spl_1
  );


  buf

  (
    G158_n_spl_110,
    G158_n_spl_11
  );


  buf

  (
    G158_n_spl_111,
    G158_n_spl_11
  );


  buf

  (
    G80_p_spl_,
    G80_p
  );


  buf

  (
    G158_p_spl_,
    G158_p
  );


  buf

  (
    G158_p_spl_0,
    G158_p_spl_
  );


  buf

  (
    G158_p_spl_00,
    G158_p_spl_0
  );


  buf

  (
    G158_p_spl_000,
    G158_p_spl_00
  );


  buf

  (
    G158_p_spl_0000,
    G158_p_spl_000
  );


  buf

  (
    G158_p_spl_0001,
    G158_p_spl_000
  );


  buf

  (
    G158_p_spl_001,
    G158_p_spl_00
  );


  buf

  (
    G158_p_spl_0010,
    G158_p_spl_001
  );


  buf

  (
    G158_p_spl_0011,
    G158_p_spl_001
  );


  buf

  (
    G158_p_spl_01,
    G158_p_spl_0
  );


  buf

  (
    G158_p_spl_010,
    G158_p_spl_01
  );


  buf

  (
    G158_p_spl_011,
    G158_p_spl_01
  );


  buf

  (
    G158_p_spl_1,
    G158_p_spl_
  );


  buf

  (
    G158_p_spl_10,
    G158_p_spl_1
  );


  buf

  (
    G158_p_spl_100,
    G158_p_spl_10
  );


  buf

  (
    G158_p_spl_101,
    G158_p_spl_10
  );


  buf

  (
    G158_p_spl_11,
    G158_p_spl_1
  );


  buf

  (
    G158_p_spl_110,
    G158_p_spl_11
  );


  buf

  (
    G158_p_spl_111,
    G158_p_spl_11
  );


  buf

  (
    G159_n_spl_,
    G159_n
  );


  buf

  (
    G159_n_spl_0,
    G159_n_spl_
  );


  buf

  (
    G159_n_spl_00,
    G159_n_spl_0
  );


  buf

  (
    G159_n_spl_000,
    G159_n_spl_00
  );


  buf

  (
    G159_n_spl_001,
    G159_n_spl_00
  );


  buf

  (
    G159_n_spl_01,
    G159_n_spl_0
  );


  buf

  (
    G159_n_spl_1,
    G159_n_spl_
  );


  buf

  (
    G159_n_spl_10,
    G159_n_spl_1
  );


  buf

  (
    G159_n_spl_11,
    G159_n_spl_1
  );


  buf

  (
    G159_p_spl_,
    G159_p
  );


  buf

  (
    G159_p_spl_0,
    G159_p_spl_
  );


  buf

  (
    G159_p_spl_00,
    G159_p_spl_0
  );


  buf

  (
    G159_p_spl_000,
    G159_p_spl_00
  );


  buf

  (
    G159_p_spl_001,
    G159_p_spl_00
  );


  buf

  (
    G159_p_spl_01,
    G159_p_spl_0
  );


  buf

  (
    G159_p_spl_1,
    G159_p_spl_
  );


  buf

  (
    G159_p_spl_10,
    G159_p_spl_1
  );


  buf

  (
    G159_p_spl_11,
    G159_p_spl_1
  );


  buf

  (
    G64_p_spl_,
    G64_p
  );


  buf

  (
    G64_p_spl_0,
    G64_p_spl_
  );


  buf

  (
    G64_p_spl_00,
    G64_p_spl_0
  );


  buf

  (
    G64_p_spl_000,
    G64_p_spl_00
  );


  buf

  (
    G64_p_spl_0000,
    G64_p_spl_000
  );


  buf

  (
    G64_p_spl_0001,
    G64_p_spl_000
  );


  buf

  (
    G64_p_spl_001,
    G64_p_spl_00
  );


  buf

  (
    G64_p_spl_0010,
    G64_p_spl_001
  );


  buf

  (
    G64_p_spl_01,
    G64_p_spl_0
  );


  buf

  (
    G64_p_spl_010,
    G64_p_spl_01
  );


  buf

  (
    G64_p_spl_011,
    G64_p_spl_01
  );


  buf

  (
    G64_p_spl_1,
    G64_p_spl_
  );


  buf

  (
    G64_p_spl_10,
    G64_p_spl_1
  );


  buf

  (
    G64_p_spl_100,
    G64_p_spl_10
  );


  buf

  (
    G64_p_spl_101,
    G64_p_spl_10
  );


  buf

  (
    G64_p_spl_11,
    G64_p_spl_1
  );


  buf

  (
    G64_p_spl_110,
    G64_p_spl_11
  );


  buf

  (
    G64_p_spl_111,
    G64_p_spl_11
  );


  buf

  (
    G160_n_spl_,
    G160_n
  );


  buf

  (
    G160_n_spl_0,
    G160_n_spl_
  );


  buf

  (
    G160_n_spl_00,
    G160_n_spl_0
  );


  buf

  (
    G160_n_spl_000,
    G160_n_spl_00
  );


  buf

  (
    G160_n_spl_0000,
    G160_n_spl_000
  );


  buf

  (
    G160_n_spl_0001,
    G160_n_spl_000
  );


  buf

  (
    G160_n_spl_001,
    G160_n_spl_00
  );


  buf

  (
    G160_n_spl_0010,
    G160_n_spl_001
  );


  buf

  (
    G160_n_spl_0011,
    G160_n_spl_001
  );


  buf

  (
    G160_n_spl_01,
    G160_n_spl_0
  );


  buf

  (
    G160_n_spl_010,
    G160_n_spl_01
  );


  buf

  (
    G160_n_spl_011,
    G160_n_spl_01
  );


  buf

  (
    G160_n_spl_1,
    G160_n_spl_
  );


  buf

  (
    G160_n_spl_10,
    G160_n_spl_1
  );


  buf

  (
    G160_n_spl_100,
    G160_n_spl_10
  );


  buf

  (
    G160_n_spl_101,
    G160_n_spl_10
  );


  buf

  (
    G160_n_spl_11,
    G160_n_spl_1
  );


  buf

  (
    G160_n_spl_110,
    G160_n_spl_11
  );


  buf

  (
    G160_n_spl_111,
    G160_n_spl_11
  );


  buf

  (
    G160_p_spl_,
    G160_p
  );


  buf

  (
    G160_p_spl_0,
    G160_p_spl_
  );


  buf

  (
    G160_p_spl_00,
    G160_p_spl_0
  );


  buf

  (
    G160_p_spl_000,
    G160_p_spl_00
  );


  buf

  (
    G160_p_spl_0000,
    G160_p_spl_000
  );


  buf

  (
    G160_p_spl_0001,
    G160_p_spl_000
  );


  buf

  (
    G160_p_spl_001,
    G160_p_spl_00
  );


  buf

  (
    G160_p_spl_0010,
    G160_p_spl_001
  );


  buf

  (
    G160_p_spl_0011,
    G160_p_spl_001
  );


  buf

  (
    G160_p_spl_01,
    G160_p_spl_0
  );


  buf

  (
    G160_p_spl_010,
    G160_p_spl_01
  );


  buf

  (
    G160_p_spl_011,
    G160_p_spl_01
  );


  buf

  (
    G160_p_spl_1,
    G160_p_spl_
  );


  buf

  (
    G160_p_spl_10,
    G160_p_spl_1
  );


  buf

  (
    G160_p_spl_100,
    G160_p_spl_10
  );


  buf

  (
    G160_p_spl_101,
    G160_p_spl_10
  );


  buf

  (
    G160_p_spl_11,
    G160_p_spl_1
  );


  buf

  (
    G160_p_spl_110,
    G160_p_spl_11
  );


  buf

  (
    G160_p_spl_111,
    G160_p_spl_11
  );


  buf

  (
    G161_n_spl_,
    G161_n
  );


  buf

  (
    G161_n_spl_0,
    G161_n_spl_
  );


  buf

  (
    G161_n_spl_00,
    G161_n_spl_0
  );


  buf

  (
    G161_n_spl_000,
    G161_n_spl_00
  );


  buf

  (
    G161_n_spl_001,
    G161_n_spl_00
  );


  buf

  (
    G161_n_spl_01,
    G161_n_spl_0
  );


  buf

  (
    G161_n_spl_1,
    G161_n_spl_
  );


  buf

  (
    G161_n_spl_10,
    G161_n_spl_1
  );


  buf

  (
    G161_n_spl_11,
    G161_n_spl_1
  );


  buf

  (
    G161_p_spl_,
    G161_p
  );


  buf

  (
    G161_p_spl_0,
    G161_p_spl_
  );


  buf

  (
    G161_p_spl_00,
    G161_p_spl_0
  );


  buf

  (
    G161_p_spl_000,
    G161_p_spl_00
  );


  buf

  (
    G161_p_spl_001,
    G161_p_spl_00
  );


  buf

  (
    G161_p_spl_01,
    G161_p_spl_0
  );


  buf

  (
    G161_p_spl_1,
    G161_p_spl_
  );


  buf

  (
    G161_p_spl_10,
    G161_p_spl_1
  );


  buf

  (
    G161_p_spl_11,
    G161_p_spl_1
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    g647_n_spl_,
    g647_n
  );


  buf

  (
    g647_n_spl_0,
    g647_n_spl_
  );


  buf

  (
    g647_n_spl_00,
    g647_n_spl_0
  );


  buf

  (
    g647_n_spl_1,
    g647_n_spl_
  );


  buf

  (
    g605_n_spl_,
    g605_n
  );


  buf

  (
    g605_n_spl_0,
    g605_n_spl_
  );


  buf

  (
    g605_n_spl_00,
    g605_n_spl_0
  );


  buf

  (
    g605_n_spl_1,
    g605_n_spl_
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G27_p_spl_,
    G27_p
  );


  buf

  (
    g656_n_spl_,
    g656_n
  );


  buf

  (
    g656_n_spl_0,
    g656_n_spl_
  );


  buf

  (
    g656_n_spl_00,
    g656_n_spl_0
  );


  buf

  (
    g656_n_spl_1,
    g656_n_spl_
  );


  buf

  (
    g614_n_spl_,
    g614_n
  );


  buf

  (
    g614_n_spl_0,
    g614_n_spl_
  );


  buf

  (
    g614_n_spl_00,
    g614_n_spl_0
  );


  buf

  (
    g614_n_spl_1,
    g614_n_spl_
  );


  buf

  (
    G5_p_spl_,
    G5_p
  );


  buf

  (
    G26_p_spl_,
    G26_p
  );


  buf

  (
    g669_n_spl_,
    g669_n
  );


  buf

  (
    g669_n_spl_0,
    g669_n_spl_
  );


  buf

  (
    g669_n_spl_00,
    g669_n_spl_0
  );


  buf

  (
    g669_n_spl_1,
    g669_n_spl_
  );


  buf

  (
    g624_n_spl_,
    g624_n
  );


  buf

  (
    g624_n_spl_0,
    g624_n_spl_
  );


  buf

  (
    g624_n_spl_00,
    g624_n_spl_0
  );


  buf

  (
    g624_n_spl_1,
    g624_n_spl_
  );


  buf

  (
    G25_p_spl_,
    G25_p
  );


  buf

  (
    G24_p_spl_,
    G24_p
  );


  buf

  (
    g678_n_spl_,
    g678_n
  );


  buf

  (
    g678_n_spl_0,
    g678_n_spl_
  );


  buf

  (
    g678_n_spl_00,
    g678_n_spl_0
  );


  buf

  (
    g678_n_spl_1,
    g678_n_spl_
  );


  buf

  (
    g569_p_spl_,
    g569_p
  );


  buf

  (
    g569_p_spl_0,
    g569_p_spl_
  );


  buf

  (
    g569_p_spl_00,
    g569_p_spl_0
  );


  buf

  (
    g569_p_spl_1,
    g569_p_spl_
  );


  buf

  (
    G76_p_spl_,
    G76_p
  );


  buf

  (
    G86_p_spl_,
    G86_p
  );


  buf

  (
    G72_p_spl_,
    G72_p
  );


  buf

  (
    G82_p_spl_,
    G82_p
  );


  buf

  (
    G70_p_spl_,
    G70_p
  );


  buf

  (
    G71_p_spl_,
    G71_p
  );


  buf

  (
    G68_p_spl_,
    G68_p
  );


  buf

  (
    G69_p_spl_,
    G69_p
  );


  buf

  (
    G171_p_spl_,
    G171_p
  );


  buf

  (
    G54_p_spl_,
    G54_p
  );


  buf

  (
    G171_n_spl_,
    G171_n
  );


  buf

  (
    G61_n_spl_,
    G61_n
  );


  buf

  (
    G61_p_spl_,
    G61_p
  );


  buf

  (
    g975_p_spl_,
    g975_p
  );


  buf

  (
    G99_n_spl_,
    G99_n
  );


  buf

  (
    g533_n_spl_,
    g533_n
  );


  buf

  (
    g735_n_spl_,
    g735_n
  );


  buf

  (
    G155_n_spl_,
    G155_n
  );


  buf

  (
    g184_n_spl_,
    g184_n
  );


  buf

  (
    g179_n_spl_,
    g179_n
  );


  buf

  (
    g705_n_spl_,
    g705_n
  );


  buf

  (
    g506_n_spl_,
    g506_n
  );


  buf

  (
    g1025_n_spl_,
    g1025_n
  );


  buf

  (
    g1025_n_spl_0,
    g1025_n_spl_
  );


  buf

  (
    g1025_n_spl_00,
    g1025_n_spl_0
  );


  buf

  (
    g1025_n_spl_1,
    g1025_n_spl_
  );


  buf

  (
    g990_p_spl_,
    g990_p
  );


  buf

  (
    g990_p_spl_0,
    g990_p_spl_
  );


  buf

  (
    g990_p_spl_00,
    g990_p_spl_0
  );


  buf

  (
    g990_p_spl_1,
    g990_p_spl_
  );


  buf

  (
    G41_p_spl_,
    G41_p
  );


  buf

  (
    G42_p_spl_,
    G42_p
  );


  buf

  (
    G18_p_spl_,
    G18_p
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


  buf

  (
    g1032_n_spl_,
    g1032_n
  );


  buf

  (
    g1032_n_spl_0,
    g1032_n_spl_
  );


  buf

  (
    g1032_n_spl_00,
    g1032_n_spl_0
  );


  buf

  (
    g1032_n_spl_1,
    g1032_n_spl_
  );


  buf

  (
    g997_n_spl_,
    g997_n
  );


  buf

  (
    g997_n_spl_0,
    g997_n_spl_
  );


  buf

  (
    g997_n_spl_00,
    g997_n_spl_0
  );


  buf

  (
    g997_n_spl_1,
    g997_n_spl_
  );


  buf

  (
    G40_p_spl_,
    G40_p
  );


  buf

  (
    G39_p_spl_,
    G39_p
  );


  buf

  (
    g1039_n_spl_,
    g1039_n
  );


  buf

  (
    g1039_n_spl_0,
    g1039_n_spl_
  );


  buf

  (
    g1039_n_spl_00,
    g1039_n_spl_0
  );


  buf

  (
    g1039_n_spl_1,
    g1039_n_spl_
  );


  buf

  (
    g1004_n_spl_,
    g1004_n
  );


  buf

  (
    g1004_n_spl_0,
    g1004_n_spl_
  );


  buf

  (
    g1004_n_spl_00,
    g1004_n_spl_0
  );


  buf

  (
    g1004_n_spl_1,
    g1004_n_spl_
  );


  buf

  (
    G15_p_spl_,
    G15_p
  );


  buf

  (
    G36_p_spl_,
    G36_p
  );


  buf

  (
    g1046_n_spl_,
    g1046_n
  );


  buf

  (
    g1046_n_spl_0,
    g1046_n_spl_
  );


  buf

  (
    g1046_n_spl_00,
    g1046_n_spl_0
  );


  buf

  (
    g1046_n_spl_1,
    g1046_n_spl_
  );


  buf

  (
    g1011_n_spl_,
    g1011_n
  );


  buf

  (
    g1011_n_spl_0,
    g1011_n_spl_
  );


  buf

  (
    g1011_n_spl_00,
    g1011_n_spl_0
  );


  buf

  (
    g1011_n_spl_1,
    g1011_n_spl_
  );


  buf

  (
    G77_p_spl_,
    G77_p
  );


  buf

  (
    G87_p_spl_,
    G87_p
  );


  buf

  (
    G75_p_spl_,
    G75_p
  );


  buf

  (
    G85_p_spl_,
    G85_p
  );


  buf

  (
    G74_p_spl_,
    G74_p
  );


  buf

  (
    G84_p_spl_,
    G84_p
  );


  buf

  (
    G73_p_spl_,
    G73_p
  );


  buf

  (
    G83_p_spl_,
    G83_p
  );


  buf

  (
    g1200_p_spl_,
    g1200_p
  );


  buf

  (
    g1202_n_spl_,
    g1202_n
  );


  buf

  (
    g1200_n_spl_,
    g1200_n
  );


  buf

  (
    g1202_p_spl_,
    g1202_p
  );


  buf

  (
    g1214_n_spl_,
    g1214_n
  );


  buf

  (
    g1223_p_spl_,
    g1223_p
  );


  buf

  (
    g1214_p_spl_,
    g1214_p
  );


  buf

  (
    g1223_n_spl_,
    g1223_n
  );


  buf

  (
    g1229_n_spl_,
    g1229_n
  );


  buf

  (
    g1238_p_spl_,
    g1238_p
  );


  buf

  (
    g1229_p_spl_,
    g1229_p
  );


  buf

  (
    g1238_n_spl_,
    g1238_n
  );


  buf

  (
    g1241_p_spl_,
    g1241_p
  );


  buf

  (
    g245_p_spl_,
    g245_p
  );


  buf

  (
    g1241_n_spl_,
    g1241_n
  );


  buf

  (
    g1226_p_spl_,
    g1226_p
  );


  buf

  (
    g1244_n_spl_,
    g1244_n
  );


  buf

  (
    g1226_n_spl_,
    g1226_n
  );


  buf

  (
    g1244_p_spl_,
    g1244_p
  );


  buf

  (
    g1254_n_spl_,
    g1254_n
  );


  buf

  (
    g617_n_spl_,
    g617_n
  );


  buf

  (
    g1254_p_spl_,
    g1254_p
  );


  buf

  (
    g1257_p_spl_,
    g1257_p
  );


  buf

  (
    g1257_n_spl_,
    g1257_n
  );


  buf

  (
    G162_n_spl_,
    G162_n
  );


  buf

  (
    G162_p_spl_,
    G162_p
  );


  buf

  (
    g1260_p_spl_,
    g1260_p
  );


  buf

  (
    g1263_p_spl_,
    g1263_p
  );


  buf

  (
    g1260_n_spl_,
    g1260_n
  );


  buf

  (
    g1263_n_spl_,
    g1263_n
  );


  buf

  (
    g1268_n_spl_,
    g1268_n
  );


  buf

  (
    g1268_p_spl_,
    g1268_p
  );


  buf

  (
    g1266_n_spl_,
    g1266_n
  );


  buf

  (
    g1271_n_spl_,
    g1271_n
  );


  buf

  (
    g1266_p_spl_,
    g1266_p
  );


  buf

  (
    g1271_p_spl_,
    g1271_p
  );


  buf

  (
    g1275_n_spl_,
    g1275_n
  );


  buf

  (
    g1275_p_spl_,
    g1275_p
  );


  buf

  (
    g1278_p_spl_,
    g1278_p
  );


  buf

  (
    g1278_n_spl_,
    g1278_n
  );


  buf

  (
    g1281_p_spl_,
    g1281_p
  );


  buf

  (
    g1281_n_spl_,
    g1281_n
  );


  buf

  (
    g1282_n_spl_,
    g1282_n
  );


  buf

  (
    g1282_p_spl_,
    g1282_p
  );


  buf

  (
    g1284_n_spl_,
    g1284_n
  );


  buf

  (
    g1284_p_spl_,
    g1284_p
  );


  buf

  (
    g1288_n_spl_,
    g1288_n
  );


  buf

  (
    g1288_p_spl_,
    g1288_p
  );


  buf

  (
    g1299_p_spl_,
    g1299_p
  );


  buf

  (
    g1299_n_spl_,
    g1299_n
  );


  buf

  (
    g1308_n_spl_,
    g1308_n
  );


  buf

  (
    g1320_n_spl_,
    g1320_n
  );


  buf

  (
    g1329_p_spl_,
    g1329_p
  );


  buf

  (
    g1320_p_spl_,
    g1320_p
  );


  buf

  (
    g1329_n_spl_,
    g1329_n
  );


  buf

  (
    g1341_n_spl_,
    g1341_n
  );


  buf

  (
    g317_p_spl_,
    g317_p
  );


  buf

  (
    g1341_p_spl_,
    g1341_p
  );


  buf

  (
    g1332_n_spl_,
    g1332_n
  );


  buf

  (
    g1344_p_spl_,
    g1344_p
  );


  buf

  (
    g1332_p_spl_,
    g1332_p
  );


  buf

  (
    g1344_n_spl_,
    g1344_n
  );


  buf

  (
    g1356_n_spl_,
    g1356_n
  );


  buf

  (
    g1365_p_spl_,
    g1365_p
  );


  buf

  (
    g1356_p_spl_,
    g1356_p
  );


  buf

  (
    g1365_n_spl_,
    g1365_n
  );


  buf

  (
    g1377_n_spl_,
    g1377_n
  );


  buf

  (
    g1386_p_spl_,
    g1386_p
  );


  buf

  (
    g1377_p_spl_,
    g1377_p
  );


  buf

  (
    g1386_n_spl_,
    g1386_n
  );


  buf

  (
    g1389_p_spl_,
    g1389_p
  );


  buf

  (
    g1398_n_spl_,
    g1398_n
  );


  buf

  (
    g1389_n_spl_,
    g1389_n
  );


  buf

  (
    g1398_p_spl_,
    g1398_p
  );


  buf

  (
    g1368_p_spl_,
    g1368_p
  );


  buf

  (
    g1401_n_spl_,
    g1401_n
  );


  buf

  (
    g1368_n_spl_,
    g1368_n
  );


  buf

  (
    g1401_p_spl_,
    g1401_p
  );


  buf

  (
    g1409_n_spl_,
    g1409_n
  );


  buf

  (
    g1412_n_spl_,
    g1412_n
  );


  buf

  (
    g1409_p_spl_,
    g1409_p
  );


  buf

  (
    g1412_p_spl_,
    g1412_p
  );


  buf

  (
    g1415_p_spl_,
    g1415_p
  );


  buf

  (
    g1415_n_spl_,
    g1415_n
  );


  buf

  (
    g1416_n_spl_,
    g1416_n
  );


  buf

  (
    g1416_p_spl_,
    g1416_p
  );


  buf

  (
    g1420_p_spl_,
    g1420_p
  );


  buf

  (
    g1420_n_spl_,
    g1420_n
  );


  buf

  (
    g1423_p_spl_,
    g1423_p
  );


  buf

  (
    g1423_n_spl_,
    g1423_n
  );


  buf

  (
    g1426_p_spl_,
    g1426_p
  );


  buf

  (
    g1426_n_spl_,
    g1426_n
  );


  buf

  (
    g1432_p_spl_,
    g1432_p
  );


  buf

  (
    g1432_n_spl_,
    g1432_n
  );


  buf

  (
    g1435_p_spl_,
    g1435_p
  );


  buf

  (
    g1435_n_spl_,
    g1435_n
  );


  buf

  (
    g1438_p_spl_,
    g1438_p
  );


  buf

  (
    g1438_n_spl_,
    g1438_n
  );


  buf

  (
    g1441_n_spl_,
    g1441_n
  );


  buf

  (
    g1441_p_spl_,
    g1441_p
  );


  buf

  (
    g1430_n_spl_,
    g1430_n
  );


  buf

  (
    g1430_p_spl_,
    g1430_p
  );


  buf

  (
    G157_n_spl_,
    G157_n
  );


  buf

  (
    G157_n_spl_0,
    G157_n_spl_
  );


  buf

  (
    G157_n_spl_1,
    G157_n_spl_
  );


  buf

  (
    G157_p_spl_,
    G157_p
  );


  buf

  (
    G157_p_spl_0,
    G157_p_spl_
  );


  buf

  (
    G157_p_spl_1,
    G157_p_spl_
  );


  buf

  (
    g1453_n_spl_,
    g1453_n
  );


  buf

  (
    g1453_p_spl_,
    g1453_p
  );


  buf

  (
    g1458_n_spl_,
    g1458_n
  );


  buf

  (
    g1458_n_spl_0,
    g1458_n_spl_
  );


  buf

  (
    g1458_n_spl_1,
    g1458_n_spl_
  );


  buf

  (
    g1458_p_spl_,
    g1458_p
  );


  buf

  (
    g1458_p_spl_0,
    g1458_p_spl_
  );


  buf

  (
    g1458_p_spl_1,
    g1458_p_spl_
  );


  buf

  (
    g1456_n_spl_,
    g1456_n
  );


  buf

  (
    g1461_p_spl_,
    g1461_p
  );


  buf

  (
    g1456_p_spl_,
    g1456_p
  );


  buf

  (
    g1461_n_spl_,
    g1461_n
  );


  buf

  (
    g1464_n_spl_,
    g1464_n
  );


  buf

  (
    g1464_p_spl_,
    g1464_p
  );


  buf

  (
    g1471_n_spl_,
    g1471_n
  );


  buf

  (
    g1471_p_spl_,
    g1471_p
  );


  buf

  (
    g1470_n_spl_,
    g1470_n
  );


  buf

  (
    g1474_p_spl_,
    g1474_p
  );


  buf

  (
    g1470_p_spl_,
    g1470_p
  );


  buf

  (
    g1474_n_spl_,
    g1474_n
  );


  buf

  (
    g1469_n_spl_,
    g1469_n
  );


  buf

  (
    g1477_p_spl_,
    g1477_p
  );


  buf

  (
    g1469_p_spl_,
    g1469_p
  );


  buf

  (
    g1477_n_spl_,
    g1477_n
  );


  buf

  (
    g1480_n_spl_,
    g1480_n
  );


  buf

  (
    g1483_p_spl_,
    g1483_p
  );


  buf

  (
    g1480_p_spl_,
    g1480_p
  );


  buf

  (
    g1483_n_spl_,
    g1483_n
  );


  buf

  (
    g1488_p_spl_,
    g1488_p
  );


  buf

  (
    g1488_n_spl_,
    g1488_n
  );


  buf

  (
    g1491_n_spl_,
    g1491_n
  );


  buf

  (
    g1491_p_spl_,
    g1491_p
  );


  buf

  (
    g1500_n_spl_,
    g1500_n
  );


  buf

  (
    G23_n_spl_,
    G23_n
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    g1509_p_spl_,
    g1509_p
  );


  buf

  (
    g1509_p_spl_0,
    g1509_p_spl_
  );


  buf

  (
    g1509_p_spl_1,
    g1509_p_spl_
  );


  buf

  (
    g1512_p_spl_,
    g1512_p
  );


  buf

  (
    g1512_p_spl_0,
    g1512_p_spl_
  );


  buf

  (
    g1512_p_spl_1,
    g1512_p_spl_
  );


  buf

  (
    G79_n_spl_,
    G79_n
  );


  buf

  (
    G78_n_spl_,
    G78_n
  );


  buf

  (
    G64_n_spl_,
    G64_n
  );


  buf

  (
    G151_n_spl_,
    G151_n
  );


  buf

  (
    G151_n_spl_0,
    G151_n_spl_
  );


  buf

  (
    G152_p_spl_,
    G152_p
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G1_n_spl_0,
    G1_n_spl_
  );


  buf

  (
    G1_n_spl_1,
    G1_n_spl_
  );


  buf

  (
    g194_n_spl_,
    g194_n
  );


  buf

  (
    g431_n_spl_,
    g431_n
  );


  buf

  (
    g482_p_spl_,
    g482_p
  );


  buf

  (
    g549_p_spl_,
    g549_p
  );


  buf

  (
    g550_n_spl_,
    g550_n
  );


endmodule
