
module mymod
(
  G1_p,
  G1_n,
  G2_p,
  G2_n,
  G3_p,
  G3_n,
  G4_p,
  G4_n,
  G5_p,
  G5_n,
  G6_p,
  G6_n,
  G7_p,
  G7_n,
  G8_p,
  G8_n,
  G9_p,
  G9_n,
  G10_p,
  G10_n,
  G11_p,
  G11_n,
  G12_p,
  G12_n,
  G13_p,
  G13_n,
  G14_p,
  G14_n,
  G15_p,
  G15_n,
  G16_p,
  G16_n,
  G17_p,
  G17_n,
  G18_p,
  G18_n,
  G19_p,
  G19_n,
  G20_p,
  G20_n,
  G21_p,
  G21_n,
  G22_p,
  G22_n,
  G23_p,
  G23_n,
  G24_p,
  G24_n,
  G25_p,
  G25_n,
  G26_p,
  G26_n,
  G27_p,
  G27_n,
  G28_p,
  G28_n,
  G29_p,
  G29_n,
  G30_p,
  G30_n,
  G31_p,
  G31_n,
  G32_p,
  G32_n,
  G6257_p,
  G6258_p,
  G6259_p,
  G6260_p,
  G6261_p,
  G6262_p,
  G6263_p,
  G6264_p,
  G6265_p,
  G6266_p,
  G6267_p,
  G6268_p,
  G6269_p,
  G6270_p,
  G6271_p,
  G6272_p,
  G6273_p,
  G6274_p,
  G6275_p,
  G6276_p,
  G6277_p,
  G6278_p,
  G6279_p,
  G6280_p,
  G6281_p,
  G6282_p,
  G6283_p,
  G6284_p,
  G6285_p,
  G6286_p,
  G6287_p,
  G6288_n
);

  input G1_p;input G1_n;input G2_p;input G2_n;input G3_p;input G3_n;input G4_p;input G4_n;input G5_p;input G5_n;input G6_p;input G6_n;input G7_p;input G7_n;input G8_p;input G8_n;input G9_p;input G9_n;input G10_p;input G10_n;input G11_p;input G11_n;input G12_p;input G12_n;input G13_p;input G13_n;input G14_p;input G14_n;input G15_p;input G15_n;input G16_p;input G16_n;input G17_p;input G17_n;input G18_p;input G18_n;input G19_p;input G19_n;input G20_p;input G20_n;input G21_p;input G21_n;input G22_p;input G22_n;input G23_p;input G23_n;input G24_p;input G24_n;input G25_p;input G25_n;input G26_p;input G26_n;input G27_p;input G27_n;input G28_p;input G28_n;input G29_p;input G29_n;input G30_p;input G30_n;input G31_p;input G31_n;input G32_p;input G32_n;
  output G6257_p;output G6258_p;output G6259_p;output G6260_p;output G6261_p;output G6262_p;output G6263_p;output G6264_p;output G6265_p;output G6266_p;output G6267_p;output G6268_p;output G6269_p;output G6270_p;output G6271_p;output G6272_p;output G6273_p;output G6274_p;output G6275_p;output G6276_p;output G6277_p;output G6278_p;output G6279_p;output G6280_p;output G6281_p;output G6282_p;output G6283_p;output G6284_p;output G6285_p;output G6286_p;output G6287_p;output G6288_n;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire g33_p;
  wire g33_n;
  wire g34_p;
  wire g34_n;
  wire g35_p;
  wire g35_n;
  wire g36_p;
  wire g36_n;
  wire g37_p;
  wire g37_n;
  wire g38_p;
  wire g38_n;
  wire g39_p;
  wire g39_n;
  wire g40_p;
  wire g40_n;
  wire g41_p;
  wire g41_n;
  wire g42_p;
  wire g42_n;
  wire g43_p;
  wire g43_n;
  wire g44_p;
  wire g44_n;
  wire g45_p;
  wire g45_n;
  wire g46_p;
  wire g46_n;
  wire g47_p;
  wire g47_n;
  wire g48_p;
  wire g48_n;
  wire g49_p;
  wire g49_n;
  wire g50_p;
  wire g50_n;
  wire g51_p;
  wire g51_n;
  wire g52_p;
  wire g52_n;
  wire g53_p;
  wire g53_n;
  wire g54_p;
  wire g54_n;
  wire g55_p;
  wire g55_n;
  wire g56_p;
  wire g56_n;
  wire g57_p;
  wire g57_n;
  wire g58_p;
  wire g58_n;
  wire g59_p;
  wire g59_n;
  wire g60_p;
  wire g60_n;
  wire g61_p;
  wire g61_n;
  wire g62_p;
  wire g62_n;
  wire g63_p;
  wire g63_n;
  wire g64_p;
  wire g64_n;
  wire g65_p;
  wire g65_n;
  wire g66_p;
  wire g66_n;
  wire g67_p;
  wire g67_n;
  wire g68_p;
  wire g68_n;
  wire g69_p;
  wire g69_n;
  wire g70_p;
  wire g70_n;
  wire g71_p;
  wire g71_n;
  wire g72_p;
  wire g72_n;
  wire g73_p;
  wire g73_n;
  wire g74_p;
  wire g74_n;
  wire g75_p;
  wire g75_n;
  wire g76_p;
  wire g76_n;
  wire g77_p;
  wire g77_n;
  wire g78_p;
  wire g78_n;
  wire g79_p;
  wire g79_n;
  wire g80_p;
  wire g80_n;
  wire g81_p;
  wire g81_n;
  wire g82_p;
  wire g82_n;
  wire g83_p;
  wire g83_n;
  wire g84_p;
  wire g84_n;
  wire g85_p;
  wire g85_n;
  wire g86_p;
  wire g86_n;
  wire g87_p;
  wire g87_n;
  wire g88_p;
  wire g88_n;
  wire g89_p;
  wire g89_n;
  wire g90_p;
  wire g90_n;
  wire g91_p;
  wire g91_n;
  wire g92_p;
  wire g92_n;
  wire g93_p;
  wire g93_n;
  wire g94_p;
  wire g94_n;
  wire g95_p;
  wire g95_n;
  wire g96_p;
  wire g96_n;
  wire g97_p;
  wire g97_n;
  wire g98_p;
  wire g98_n;
  wire g99_p;
  wire g99_n;
  wire g100_p;
  wire g100_n;
  wire g101_p;
  wire g101_n;
  wire g102_p;
  wire g102_n;
  wire g103_p;
  wire g103_n;
  wire g104_p;
  wire g104_n;
  wire g105_p;
  wire g105_n;
  wire g106_p;
  wire g106_n;
  wire g107_p;
  wire g107_n;
  wire g108_p;
  wire g108_n;
  wire g109_p;
  wire g109_n;
  wire g110_p;
  wire g110_n;
  wire g111_p;
  wire g111_n;
  wire g112_p;
  wire g112_n;
  wire g113_p;
  wire g113_n;
  wire g114_p;
  wire g114_n;
  wire g115_p;
  wire g115_n;
  wire g116_p;
  wire g116_n;
  wire g117_p;
  wire g117_n;
  wire g118_p;
  wire g118_n;
  wire g119_p;
  wire g119_n;
  wire g120_p;
  wire g120_n;
  wire g121_p;
  wire g121_n;
  wire g122_p;
  wire g122_n;
  wire g123_p;
  wire g123_n;
  wire g124_p;
  wire g124_n;
  wire g125_p;
  wire g125_n;
  wire g126_p;
  wire g126_n;
  wire g127_p;
  wire g127_n;
  wire g128_p;
  wire g128_n;
  wire g129_p;
  wire g129_n;
  wire g130_p;
  wire g130_n;
  wire g131_p;
  wire g131_n;
  wire g132_p;
  wire g132_n;
  wire g133_p;
  wire g133_n;
  wire g134_p;
  wire g134_n;
  wire g135_p;
  wire g135_n;
  wire g136_p;
  wire g136_n;
  wire g137_p;
  wire g137_n;
  wire g138_p;
  wire g138_n;
  wire g139_p;
  wire g139_n;
  wire g140_p;
  wire g140_n;
  wire g141_p;
  wire g141_n;
  wire g142_p;
  wire g142_n;
  wire g143_p;
  wire g143_n;
  wire g144_p;
  wire g144_n;
  wire g145_p;
  wire g145_n;
  wire g146_p;
  wire g146_n;
  wire g147_p;
  wire g147_n;
  wire g148_p;
  wire g148_n;
  wire g149_p;
  wire g149_n;
  wire g150_p;
  wire g150_n;
  wire g151_p;
  wire g151_n;
  wire g152_p;
  wire g152_n;
  wire g153_p;
  wire g153_n;
  wire g154_p;
  wire g154_n;
  wire g155_p;
  wire g155_n;
  wire g156_p;
  wire g156_n;
  wire g157_p;
  wire g157_n;
  wire g158_p;
  wire g158_n;
  wire g159_p;
  wire g159_n;
  wire g160_p;
  wire g160_n;
  wire g161_p;
  wire g161_n;
  wire g162_p;
  wire g162_n;
  wire g163_p;
  wire g163_n;
  wire g164_p;
  wire g164_n;
  wire g165_p;
  wire g165_n;
  wire g166_p;
  wire g166_n;
  wire g167_p;
  wire g167_n;
  wire g168_p;
  wire g168_n;
  wire g169_p;
  wire g169_n;
  wire g170_p;
  wire g170_n;
  wire g171_p;
  wire g171_n;
  wire g172_p;
  wire g172_n;
  wire g173_p;
  wire g173_n;
  wire g174_p;
  wire g174_n;
  wire g175_p;
  wire g175_n;
  wire g176_p;
  wire g176_n;
  wire g177_p;
  wire g177_n;
  wire g178_p;
  wire g178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire g686_p;
  wire g686_n;
  wire g687_p;
  wire g687_n;
  wire g688_p;
  wire g688_n;
  wire g689_p;
  wire g689_n;
  wire g690_p;
  wire g690_n;
  wire g691_p;
  wire g691_n;
  wire g692_p;
  wire g692_n;
  wire g693_p;
  wire g693_n;
  wire g694_p;
  wire g694_n;
  wire g695_p;
  wire g695_n;
  wire g696_p;
  wire g696_n;
  wire g697_p;
  wire g697_n;
  wire g698_p;
  wire g698_n;
  wire g699_p;
  wire g699_n;
  wire g700_p;
  wire g700_n;
  wire g701_p;
  wire g701_n;
  wire g702_p;
  wire g702_n;
  wire g703_p;
  wire g703_n;
  wire g704_p;
  wire g704_n;
  wire g705_p;
  wire g705_n;
  wire g706_p;
  wire g706_n;
  wire g707_p;
  wire g707_n;
  wire g708_p;
  wire g708_n;
  wire g709_p;
  wire g709_n;
  wire g710_p;
  wire g710_n;
  wire g711_p;
  wire g711_n;
  wire g712_p;
  wire g712_n;
  wire g713_p;
  wire g713_n;
  wire g714_p;
  wire g714_n;
  wire g715_p;
  wire g715_n;
  wire g716_p;
  wire g716_n;
  wire g717_p;
  wire g717_n;
  wire g718_p;
  wire g718_n;
  wire g719_p;
  wire g719_n;
  wire g720_p;
  wire g720_n;
  wire g721_p;
  wire g721_n;
  wire g722_p;
  wire g722_n;
  wire g723_p;
  wire g723_n;
  wire g724_p;
  wire g724_n;
  wire g725_p;
  wire g725_n;
  wire g726_p;
  wire g726_n;
  wire g727_p;
  wire g727_n;
  wire g728_p;
  wire g728_n;
  wire g729_p;
  wire g729_n;
  wire g730_p;
  wire g730_n;
  wire g731_p;
  wire g731_n;
  wire g732_p;
  wire g732_n;
  wire g733_p;
  wire g733_n;
  wire g734_p;
  wire g734_n;
  wire g735_p;
  wire g735_n;
  wire g736_p;
  wire g736_n;
  wire g737_p;
  wire g737_n;
  wire g738_p;
  wire g738_n;
  wire g739_p;
  wire g739_n;
  wire g740_p;
  wire g740_n;
  wire g741_p;
  wire g741_n;
  wire g742_p;
  wire g742_n;
  wire g743_p;
  wire g743_n;
  wire g744_p;
  wire g744_n;
  wire g745_p;
  wire g745_n;
  wire g746_p;
  wire g746_n;
  wire g747_p;
  wire g747_n;
  wire g748_p;
  wire g748_n;
  wire g749_p;
  wire g749_n;
  wire g750_p;
  wire g750_n;
  wire g751_p;
  wire g751_n;
  wire g752_p;
  wire g752_n;
  wire g753_p;
  wire g753_n;
  wire g754_p;
  wire g754_n;
  wire g755_p;
  wire g755_n;
  wire g756_p;
  wire g756_n;
  wire g757_p;
  wire g757_n;
  wire g758_p;
  wire g758_n;
  wire g759_p;
  wire g759_n;
  wire g760_p;
  wire g760_n;
  wire g761_p;
  wire g761_n;
  wire g762_p;
  wire g762_n;
  wire g763_p;
  wire g763_n;
  wire g764_p;
  wire g764_n;
  wire g765_p;
  wire g765_n;
  wire g766_p;
  wire g766_n;
  wire g767_p;
  wire g767_n;
  wire g768_p;
  wire g768_n;
  wire g769_p;
  wire g769_n;
  wire g770_p;
  wire g770_n;
  wire g771_p;
  wire g771_n;
  wire g772_p;
  wire g772_n;
  wire g773_p;
  wire g773_n;
  wire g774_p;
  wire g774_n;
  wire g775_p;
  wire g775_n;
  wire g776_p;
  wire g776_n;
  wire g777_p;
  wire g777_n;
  wire g778_p;
  wire g778_n;
  wire g779_p;
  wire g779_n;
  wire g780_p;
  wire g780_n;
  wire g781_p;
  wire g781_n;
  wire g782_p;
  wire g782_n;
  wire g783_p;
  wire g783_n;
  wire g784_p;
  wire g784_n;
  wire g785_p;
  wire g785_n;
  wire g786_p;
  wire g786_n;
  wire g787_p;
  wire g787_n;
  wire g788_p;
  wire g788_n;
  wire g789_p;
  wire g789_n;
  wire g790_p;
  wire g790_n;
  wire g791_p;
  wire g791_n;
  wire g792_p;
  wire g792_n;
  wire g793_p;
  wire g793_n;
  wire g794_p;
  wire g794_n;
  wire g795_p;
  wire g795_n;
  wire g796_p;
  wire g796_n;
  wire g797_p;
  wire g797_n;
  wire g798_p;
  wire g798_n;
  wire g799_p;
  wire g799_n;
  wire g800_p;
  wire g800_n;
  wire g801_p;
  wire g801_n;
  wire g802_p;
  wire g802_n;
  wire g803_p;
  wire g803_n;
  wire g804_p;
  wire g804_n;
  wire g805_p;
  wire g805_n;
  wire g806_p;
  wire g806_n;
  wire g807_p;
  wire g807_n;
  wire g808_p;
  wire g808_n;
  wire g809_p;
  wire g809_n;
  wire g810_p;
  wire g810_n;
  wire g811_p;
  wire g811_n;
  wire g812_p;
  wire g812_n;
  wire g813_p;
  wire g813_n;
  wire g814_p;
  wire g814_n;
  wire g815_p;
  wire g815_n;
  wire g816_p;
  wire g816_n;
  wire g817_p;
  wire g817_n;
  wire g818_p;
  wire g818_n;
  wire g819_p;
  wire g819_n;
  wire g820_p;
  wire g820_n;
  wire g821_p;
  wire g821_n;
  wire g822_p;
  wire g822_n;
  wire g823_p;
  wire g823_n;
  wire g824_p;
  wire g824_n;
  wire g825_p;
  wire g825_n;
  wire g826_p;
  wire g826_n;
  wire g827_p;
  wire g827_n;
  wire g828_p;
  wire g828_n;
  wire g829_p;
  wire g829_n;
  wire g830_p;
  wire g830_n;
  wire g831_p;
  wire g831_n;
  wire g832_p;
  wire g832_n;
  wire g833_p;
  wire g833_n;
  wire g834_p;
  wire g834_n;
  wire g835_p;
  wire g835_n;
  wire g836_p;
  wire g836_n;
  wire g837_p;
  wire g837_n;
  wire g838_p;
  wire g838_n;
  wire g839_p;
  wire g839_n;
  wire g840_p;
  wire g840_n;
  wire g841_p;
  wire g841_n;
  wire g842_p;
  wire g842_n;
  wire g843_p;
  wire g843_n;
  wire g844_p;
  wire g844_n;
  wire g845_p;
  wire g845_n;
  wire g846_p;
  wire g846_n;
  wire g847_p;
  wire g847_n;
  wire g848_p;
  wire g848_n;
  wire g849_p;
  wire g849_n;
  wire g850_p;
  wire g850_n;
  wire g851_p;
  wire g851_n;
  wire g852_p;
  wire g852_n;
  wire g853_p;
  wire g853_n;
  wire g854_p;
  wire g854_n;
  wire g855_p;
  wire g855_n;
  wire g856_p;
  wire g856_n;
  wire g857_p;
  wire g857_n;
  wire g858_p;
  wire g858_n;
  wire g859_p;
  wire g859_n;
  wire g860_p;
  wire g860_n;
  wire g861_p;
  wire g861_n;
  wire g862_p;
  wire g862_n;
  wire g863_p;
  wire g863_n;
  wire g864_p;
  wire g864_n;
  wire g865_p;
  wire g865_n;
  wire g866_p;
  wire g866_n;
  wire g867_p;
  wire g867_n;
  wire g868_p;
  wire g868_n;
  wire g869_p;
  wire g869_n;
  wire g870_p;
  wire g870_n;
  wire g871_p;
  wire g871_n;
  wire g872_p;
  wire g872_n;
  wire g873_p;
  wire g873_n;
  wire g874_p;
  wire g874_n;
  wire g875_p;
  wire g875_n;
  wire g876_p;
  wire g876_n;
  wire g877_p;
  wire g877_n;
  wire g878_p;
  wire g878_n;
  wire g879_p;
  wire g879_n;
  wire g880_p;
  wire g880_n;
  wire g881_p;
  wire g881_n;
  wire g882_p;
  wire g882_n;
  wire g883_p;
  wire g883_n;
  wire g884_p;
  wire g884_n;
  wire g885_p;
  wire g885_n;
  wire g886_p;
  wire g886_n;
  wire g887_p;
  wire g887_n;
  wire g888_p;
  wire g888_n;
  wire g889_p;
  wire g889_n;
  wire g890_p;
  wire g890_n;
  wire g891_p;
  wire g891_n;
  wire g892_p;
  wire g892_n;
  wire g893_p;
  wire g893_n;
  wire g894_p;
  wire g894_n;
  wire g895_p;
  wire g895_n;
  wire g896_p;
  wire g896_n;
  wire g897_p;
  wire g897_n;
  wire g898_p;
  wire g898_n;
  wire g899_p;
  wire g899_n;
  wire g900_p;
  wire g900_n;
  wire g901_p;
  wire g901_n;
  wire g902_p;
  wire g902_n;
  wire g903_p;
  wire g903_n;
  wire g904_p;
  wire g904_n;
  wire g905_p;
  wire g905_n;
  wire g906_p;
  wire g906_n;
  wire g907_p;
  wire g907_n;
  wire g908_p;
  wire g908_n;
  wire g909_p;
  wire g909_n;
  wire g910_p;
  wire g910_n;
  wire g911_p;
  wire g911_n;
  wire g912_p;
  wire g912_n;
  wire g913_p;
  wire g913_n;
  wire g914_p;
  wire g914_n;
  wire g915_p;
  wire g915_n;
  wire g916_p;
  wire g916_n;
  wire g917_p;
  wire g917_n;
  wire g918_p;
  wire g918_n;
  wire g919_p;
  wire g919_n;
  wire g920_p;
  wire g920_n;
  wire g921_p;
  wire g921_n;
  wire g922_p;
  wire g922_n;
  wire g923_p;
  wire g923_n;
  wire g924_p;
  wire g924_n;
  wire g925_p;
  wire g925_n;
  wire g926_p;
  wire g926_n;
  wire g927_p;
  wire g927_n;
  wire g928_p;
  wire g928_n;
  wire g929_p;
  wire g929_n;
  wire g930_p;
  wire g930_n;
  wire g931_p;
  wire g931_n;
  wire g932_p;
  wire g932_n;
  wire g933_p;
  wire g933_n;
  wire g934_p;
  wire g934_n;
  wire g935_p;
  wire g935_n;
  wire g936_p;
  wire g936_n;
  wire g937_p;
  wire g937_n;
  wire g938_p;
  wire g938_n;
  wire g939_p;
  wire g939_n;
  wire g940_p;
  wire g940_n;
  wire g941_p;
  wire g941_n;
  wire g942_p;
  wire g942_n;
  wire g943_p;
  wire g943_n;
  wire g944_p;
  wire g944_n;
  wire g945_p;
  wire g945_n;
  wire g946_p;
  wire g946_n;
  wire g947_p;
  wire g947_n;
  wire g948_p;
  wire g948_n;
  wire g949_p;
  wire g949_n;
  wire g950_p;
  wire g950_n;
  wire g951_p;
  wire g951_n;
  wire g952_p;
  wire g952_n;
  wire g953_p;
  wire g953_n;
  wire g954_p;
  wire g954_n;
  wire g955_p;
  wire g955_n;
  wire g956_p;
  wire g956_n;
  wire g957_p;
  wire g957_n;
  wire g958_p;
  wire g958_n;
  wire g959_p;
  wire g959_n;
  wire g960_p;
  wire g960_n;
  wire g961_p;
  wire g961_n;
  wire g962_p;
  wire g962_n;
  wire g963_p;
  wire g963_n;
  wire g964_p;
  wire g964_n;
  wire g965_p;
  wire g965_n;
  wire g966_p;
  wire g966_n;
  wire g967_p;
  wire g967_n;
  wire g968_p;
  wire g968_n;
  wire g969_p;
  wire g969_n;
  wire g970_p;
  wire g970_n;
  wire g971_p;
  wire g971_n;
  wire g972_p;
  wire g972_n;
  wire g973_p;
  wire g973_n;
  wire g974_p;
  wire g974_n;
  wire g975_p;
  wire g975_n;
  wire g976_p;
  wire g976_n;
  wire g977_p;
  wire g977_n;
  wire g978_p;
  wire g978_n;
  wire g979_p;
  wire g979_n;
  wire g980_p;
  wire g980_n;
  wire g981_p;
  wire g981_n;
  wire g982_p;
  wire g982_n;
  wire g983_p;
  wire g983_n;
  wire g984_p;
  wire g984_n;
  wire g985_p;
  wire g985_n;
  wire g986_p;
  wire g986_n;
  wire g987_p;
  wire g987_n;
  wire g988_p;
  wire g988_n;
  wire g989_p;
  wire g989_n;
  wire g990_p;
  wire g990_n;
  wire g991_p;
  wire g991_n;
  wire g992_p;
  wire g992_n;
  wire g993_p;
  wire g993_n;
  wire g994_p;
  wire g994_n;
  wire g995_p;
  wire g995_n;
  wire g996_p;
  wire g996_n;
  wire g997_p;
  wire g997_n;
  wire g998_p;
  wire g998_n;
  wire g999_p;
  wire g999_n;
  wire g1000_p;
  wire g1000_n;
  wire g1001_p;
  wire g1001_n;
  wire g1002_p;
  wire g1002_n;
  wire g1003_p;
  wire g1003_n;
  wire g1004_p;
  wire g1004_n;
  wire g1005_p;
  wire g1005_n;
  wire g1006_p;
  wire g1006_n;
  wire g1007_p;
  wire g1007_n;
  wire g1008_p;
  wire g1008_n;
  wire g1009_p;
  wire g1009_n;
  wire g1010_p;
  wire g1010_n;
  wire g1011_p;
  wire g1011_n;
  wire g1012_p;
  wire g1012_n;
  wire g1013_p;
  wire g1013_n;
  wire g1014_p;
  wire g1014_n;
  wire g1015_p;
  wire g1015_n;
  wire g1016_p;
  wire g1016_n;
  wire g1017_p;
  wire g1017_n;
  wire g1018_p;
  wire g1018_n;
  wire g1019_p;
  wire g1019_n;
  wire g1020_p;
  wire g1020_n;
  wire g1021_p;
  wire g1021_n;
  wire g1022_p;
  wire g1022_n;
  wire g1023_p;
  wire g1023_n;
  wire g1024_p;
  wire g1024_n;
  wire g1025_p;
  wire g1025_n;
  wire g1026_p;
  wire g1026_n;
  wire g1027_p;
  wire g1027_n;
  wire g1028_p;
  wire g1028_n;
  wire g1029_p;
  wire g1029_n;
  wire g1030_p;
  wire g1030_n;
  wire g1031_p;
  wire g1031_n;
  wire g1032_p;
  wire g1032_n;
  wire g1033_p;
  wire g1033_n;
  wire g1034_p;
  wire g1034_n;
  wire g1035_p;
  wire g1035_n;
  wire g1036_p;
  wire g1036_n;
  wire g1037_p;
  wire g1037_n;
  wire g1038_p;
  wire g1038_n;
  wire g1039_p;
  wire g1039_n;
  wire g1040_p;
  wire g1040_n;
  wire g1041_p;
  wire g1041_n;
  wire g1042_p;
  wire g1042_n;
  wire g1043_p;
  wire g1043_n;
  wire g1044_p;
  wire g1044_n;
  wire g1045_p;
  wire g1045_n;
  wire g1046_p;
  wire g1046_n;
  wire g1047_p;
  wire g1047_n;
  wire g1048_p;
  wire g1048_n;
  wire g1049_p;
  wire g1049_n;
  wire g1050_p;
  wire g1050_n;
  wire g1051_p;
  wire g1051_n;
  wire g1052_p;
  wire g1052_n;
  wire g1053_p;
  wire g1053_n;
  wire g1054_p;
  wire g1054_n;
  wire g1055_p;
  wire g1055_n;
  wire g1056_p;
  wire g1056_n;
  wire g1057_p;
  wire g1057_n;
  wire g1058_p;
  wire g1058_n;
  wire g1059_p;
  wire g1059_n;
  wire g1060_p;
  wire g1060_n;
  wire g1061_p;
  wire g1061_n;
  wire g1062_p;
  wire g1062_n;
  wire g1063_p;
  wire g1063_n;
  wire g1064_p;
  wire g1064_n;
  wire g1065_p;
  wire g1065_n;
  wire g1066_p;
  wire g1066_n;
  wire g1067_p;
  wire g1067_n;
  wire g1068_p;
  wire g1068_n;
  wire g1069_p;
  wire g1069_n;
  wire g1070_p;
  wire g1070_n;
  wire g1071_p;
  wire g1071_n;
  wire g1072_p;
  wire g1072_n;
  wire g1073_p;
  wire g1073_n;
  wire g1074_p;
  wire g1074_n;
  wire g1075_p;
  wire g1075_n;
  wire g1076_p;
  wire g1076_n;
  wire g1077_p;
  wire g1077_n;
  wire g1078_p;
  wire g1078_n;
  wire g1079_p;
  wire g1079_n;
  wire g1080_p;
  wire g1080_n;
  wire g1081_p;
  wire g1081_n;
  wire g1082_p;
  wire g1082_n;
  wire g1083_p;
  wire g1083_n;
  wire g1084_p;
  wire g1084_n;
  wire g1085_p;
  wire g1085_n;
  wire g1086_p;
  wire g1086_n;
  wire g1087_p;
  wire g1087_n;
  wire g1088_p;
  wire g1088_n;
  wire g1089_p;
  wire g1089_n;
  wire g1090_p;
  wire g1090_n;
  wire g1091_p;
  wire g1091_n;
  wire g1092_p;
  wire g1092_n;
  wire g1093_p;
  wire g1093_n;
  wire g1094_p;
  wire g1094_n;
  wire g1095_p;
  wire g1095_n;
  wire g1096_p;
  wire g1096_n;
  wire g1097_p;
  wire g1097_n;
  wire g1098_p;
  wire g1098_n;
  wire g1099_p;
  wire g1099_n;
  wire g1100_p;
  wire g1100_n;
  wire g1101_p;
  wire g1101_n;
  wire g1102_p;
  wire g1102_n;
  wire g1103_p;
  wire g1103_n;
  wire g1104_p;
  wire g1104_n;
  wire g1105_p;
  wire g1105_n;
  wire g1106_p;
  wire g1106_n;
  wire g1107_p;
  wire g1107_n;
  wire g1108_p;
  wire g1108_n;
  wire g1109_p;
  wire g1109_n;
  wire g1110_p;
  wire g1110_n;
  wire g1111_p;
  wire g1111_n;
  wire g1112_p;
  wire g1112_n;
  wire g1113_p;
  wire g1113_n;
  wire g1114_p;
  wire g1114_n;
  wire g1115_p;
  wire g1115_n;
  wire g1116_p;
  wire g1116_n;
  wire g1117_p;
  wire g1117_n;
  wire g1118_p;
  wire g1118_n;
  wire g1119_p;
  wire g1119_n;
  wire g1120_p;
  wire g1120_n;
  wire g1121_p;
  wire g1121_n;
  wire g1122_p;
  wire g1122_n;
  wire g1123_p;
  wire g1123_n;
  wire g1124_p;
  wire g1124_n;
  wire g1125_p;
  wire g1125_n;
  wire g1126_p;
  wire g1126_n;
  wire g1127_p;
  wire g1127_n;
  wire g1128_p;
  wire g1128_n;
  wire g1129_p;
  wire g1129_n;
  wire g1130_p;
  wire g1130_n;
  wire g1131_p;
  wire g1131_n;
  wire g1132_p;
  wire g1132_n;
  wire g1133_p;
  wire g1133_n;
  wire g1134_p;
  wire g1134_n;
  wire g1135_p;
  wire g1135_n;
  wire g1136_p;
  wire g1136_n;
  wire g1137_p;
  wire g1137_n;
  wire g1138_p;
  wire g1138_n;
  wire g1139_p;
  wire g1139_n;
  wire g1140_p;
  wire g1140_n;
  wire g1141_p;
  wire g1141_n;
  wire g1142_p;
  wire g1142_n;
  wire g1143_p;
  wire g1143_n;
  wire g1144_p;
  wire g1144_n;
  wire g1145_p;
  wire g1145_n;
  wire g1146_p;
  wire g1146_n;
  wire g1147_p;
  wire g1147_n;
  wire g1148_p;
  wire g1148_n;
  wire g1149_p;
  wire g1149_n;
  wire g1150_p;
  wire g1150_n;
  wire g1151_p;
  wire g1151_n;
  wire g1152_p;
  wire g1152_n;
  wire g1153_p;
  wire g1153_n;
  wire g1154_p;
  wire g1154_n;
  wire g1155_p;
  wire g1155_n;
  wire g1156_p;
  wire g1156_n;
  wire g1157_p;
  wire g1157_n;
  wire g1158_p;
  wire g1158_n;
  wire g1159_p;
  wire g1159_n;
  wire g1160_p;
  wire g1160_n;
  wire g1161_p;
  wire g1161_n;
  wire g1162_p;
  wire g1162_n;
  wire g1163_p;
  wire g1163_n;
  wire g1164_p;
  wire g1164_n;
  wire g1165_p;
  wire g1165_n;
  wire g1166_p;
  wire g1166_n;
  wire g1167_p;
  wire g1167_n;
  wire g1168_p;
  wire g1168_n;
  wire g1169_p;
  wire g1169_n;
  wire g1170_p;
  wire g1170_n;
  wire g1171_p;
  wire g1171_n;
  wire g1172_p;
  wire g1172_n;
  wire g1173_p;
  wire g1173_n;
  wire g1174_p;
  wire g1174_n;
  wire g1175_p;
  wire g1175_n;
  wire g1176_p;
  wire g1176_n;
  wire g1177_p;
  wire g1177_n;
  wire g1178_p;
  wire g1178_n;
  wire g1179_p;
  wire g1179_n;
  wire g1180_p;
  wire g1180_n;
  wire g1181_p;
  wire g1181_n;
  wire g1182_p;
  wire g1182_n;
  wire g1183_p;
  wire g1183_n;
  wire g1184_p;
  wire g1184_n;
  wire g1185_p;
  wire g1185_n;
  wire g1186_p;
  wire g1186_n;
  wire g1187_p;
  wire g1187_n;
  wire g1188_p;
  wire g1188_n;
  wire g1189_p;
  wire g1189_n;
  wire g1190_p;
  wire g1190_n;
  wire g1191_p;
  wire g1191_n;
  wire g1192_p;
  wire g1192_n;
  wire g1193_p;
  wire g1193_n;
  wire g1194_p;
  wire g1194_n;
  wire g1195_p;
  wire g1195_n;
  wire g1196_p;
  wire g1196_n;
  wire g1197_p;
  wire g1197_n;
  wire g1198_p;
  wire g1198_n;
  wire g1199_p;
  wire g1199_n;
  wire g1200_p;
  wire g1200_n;
  wire g1201_p;
  wire g1201_n;
  wire g1202_p;
  wire g1202_n;
  wire g1203_p;
  wire g1203_n;
  wire g1204_p;
  wire g1204_n;
  wire g1205_p;
  wire g1205_n;
  wire g1206_p;
  wire g1206_n;
  wire g1207_p;
  wire g1207_n;
  wire g1208_p;
  wire g1208_n;
  wire g1209_p;
  wire g1209_n;
  wire g1210_p;
  wire g1210_n;
  wire g1211_p;
  wire g1211_n;
  wire g1212_p;
  wire g1212_n;
  wire g1213_p;
  wire g1213_n;
  wire g1214_p;
  wire g1214_n;
  wire g1215_p;
  wire g1215_n;
  wire g1216_p;
  wire g1216_n;
  wire g1217_p;
  wire g1217_n;
  wire g1218_p;
  wire g1218_n;
  wire g1219_p;
  wire g1219_n;
  wire g1220_p;
  wire g1220_n;
  wire g1221_p;
  wire g1221_n;
  wire g1222_p;
  wire g1222_n;
  wire g1223_p;
  wire g1223_n;
  wire g1224_p;
  wire g1224_n;
  wire g1225_p;
  wire g1225_n;
  wire g1226_p;
  wire g1226_n;
  wire g1227_p;
  wire g1227_n;
  wire g1228_p;
  wire g1228_n;
  wire g1229_p;
  wire g1229_n;
  wire g1230_p;
  wire g1230_n;
  wire g1231_p;
  wire g1231_n;
  wire g1232_p;
  wire g1232_n;
  wire g1233_p;
  wire g1233_n;
  wire g1234_p;
  wire g1234_n;
  wire g1235_p;
  wire g1235_n;
  wire g1236_p;
  wire g1236_n;
  wire g1237_p;
  wire g1237_n;
  wire g1238_p;
  wire g1238_n;
  wire g1239_p;
  wire g1239_n;
  wire g1240_p;
  wire g1240_n;
  wire g1241_p;
  wire g1241_n;
  wire g1242_p;
  wire g1242_n;
  wire g1243_p;
  wire g1243_n;
  wire g1244_p;
  wire g1244_n;
  wire g1245_p;
  wire g1245_n;
  wire g1246_p;
  wire g1246_n;
  wire g1247_p;
  wire g1247_n;
  wire g1248_p;
  wire g1248_n;
  wire g1249_p;
  wire g1249_n;
  wire g1250_p;
  wire g1250_n;
  wire g1251_p;
  wire g1251_n;
  wire g1252_p;
  wire g1252_n;
  wire g1253_p;
  wire g1253_n;
  wire g1254_p;
  wire g1254_n;
  wire g1255_p;
  wire g1255_n;
  wire g1256_p;
  wire g1256_n;
  wire g1257_p;
  wire g1257_n;
  wire g1258_p;
  wire g1258_n;
  wire g1259_p;
  wire g1259_n;
  wire g1260_p;
  wire g1260_n;
  wire g1261_p;
  wire g1261_n;
  wire g1262_p;
  wire g1262_n;
  wire g1263_p;
  wire g1263_n;
  wire g1264_p;
  wire g1264_n;
  wire g1265_p;
  wire g1265_n;
  wire g1266_p;
  wire g1266_n;
  wire g1267_p;
  wire g1267_n;
  wire g1268_p;
  wire g1268_n;
  wire g1269_p;
  wire g1269_n;
  wire g1270_p;
  wire g1270_n;
  wire g1271_p;
  wire g1271_n;
  wire g1272_p;
  wire g1272_n;
  wire g1273_p;
  wire g1273_n;
  wire g1274_p;
  wire g1274_n;
  wire g1275_p;
  wire g1275_n;
  wire g1276_p;
  wire g1276_n;
  wire g1277_p;
  wire g1277_n;
  wire g1278_p;
  wire g1278_n;
  wire g1279_p;
  wire g1279_n;
  wire g1280_p;
  wire g1280_n;
  wire g1281_p;
  wire g1281_n;
  wire g1282_p;
  wire g1282_n;
  wire g1283_p;
  wire g1283_n;
  wire g1284_p;
  wire g1284_n;
  wire g1285_p;
  wire g1285_n;
  wire g1286_p;
  wire g1286_n;
  wire g1287_p;
  wire g1287_n;
  wire g1288_p;
  wire g1288_n;
  wire g1289_p;
  wire g1289_n;
  wire g1290_p;
  wire g1290_n;
  wire g1291_p;
  wire g1291_n;
  wire g1292_p;
  wire g1292_n;
  wire g1293_p;
  wire g1293_n;
  wire g1294_p;
  wire g1294_n;
  wire g1295_p;
  wire g1295_n;
  wire g1296_p;
  wire g1296_n;
  wire g1297_p;
  wire g1297_n;
  wire g1298_p;
  wire g1298_n;
  wire g1299_p;
  wire g1299_n;
  wire g1300_p;
  wire g1300_n;
  wire g1301_p;
  wire g1301_n;
  wire g1302_p;
  wire g1302_n;
  wire g1303_p;
  wire g1303_n;
  wire g1304_p;
  wire g1304_n;
  wire g1305_p;
  wire g1305_n;
  wire g1306_p;
  wire g1306_n;
  wire g1307_p;
  wire g1307_n;
  wire g1308_p;
  wire g1308_n;
  wire g1309_p;
  wire g1309_n;
  wire g1310_p;
  wire g1310_n;
  wire g1311_p;
  wire g1311_n;
  wire g1312_p;
  wire g1312_n;
  wire g1313_p;
  wire g1313_n;
  wire g1314_p;
  wire g1314_n;
  wire g1315_p;
  wire g1315_n;
  wire g1316_p;
  wire g1316_n;
  wire g1317_p;
  wire g1317_n;
  wire g1318_p;
  wire g1318_n;
  wire g1319_p;
  wire g1319_n;
  wire g1320_p;
  wire g1320_n;
  wire g1321_p;
  wire g1321_n;
  wire g1322_p;
  wire g1322_n;
  wire g1323_p;
  wire g1323_n;
  wire g1324_p;
  wire g1324_n;
  wire g1325_p;
  wire g1325_n;
  wire g1326_p;
  wire g1326_n;
  wire g1327_p;
  wire g1327_n;
  wire g1328_p;
  wire g1328_n;
  wire g1329_p;
  wire g1329_n;
  wire g1330_p;
  wire g1330_n;
  wire g1331_p;
  wire g1331_n;
  wire g1332_p;
  wire g1332_n;
  wire g1333_p;
  wire g1333_n;
  wire g1334_p;
  wire g1334_n;
  wire g1335_p;
  wire g1335_n;
  wire g1336_p;
  wire g1336_n;
  wire g1337_p;
  wire g1337_n;
  wire g1338_p;
  wire g1338_n;
  wire g1339_p;
  wire g1339_n;
  wire g1340_p;
  wire g1340_n;
  wire g1341_p;
  wire g1341_n;
  wire g1342_p;
  wire g1342_n;
  wire g1343_p;
  wire g1343_n;
  wire g1344_p;
  wire g1344_n;
  wire g1345_p;
  wire g1345_n;
  wire g1346_p;
  wire g1346_n;
  wire g1347_p;
  wire g1347_n;
  wire g1348_p;
  wire g1348_n;
  wire g1349_p;
  wire g1349_n;
  wire g1350_p;
  wire g1350_n;
  wire g1351_p;
  wire g1351_n;
  wire g1352_p;
  wire g1352_n;
  wire g1353_p;
  wire g1353_n;
  wire g1354_p;
  wire g1354_n;
  wire g1355_p;
  wire g1355_n;
  wire g1356_p;
  wire g1356_n;
  wire g1357_p;
  wire g1357_n;
  wire g1358_p;
  wire g1358_n;
  wire g1359_p;
  wire g1359_n;
  wire g1360_p;
  wire g1360_n;
  wire g1361_p;
  wire g1361_n;
  wire g1362_p;
  wire g1362_n;
  wire g1363_p;
  wire g1363_n;
  wire g1364_p;
  wire g1364_n;
  wire g1365_p;
  wire g1365_n;
  wire g1366_p;
  wire g1366_n;
  wire g1367_p;
  wire g1367_n;
  wire g1368_p;
  wire g1368_n;
  wire g1369_p;
  wire g1369_n;
  wire g1370_p;
  wire g1370_n;
  wire g1371_p;
  wire g1371_n;
  wire g1372_p;
  wire g1372_n;
  wire g1373_p;
  wire g1373_n;
  wire g1374_p;
  wire g1374_n;
  wire g1375_p;
  wire g1375_n;
  wire g1376_p;
  wire g1376_n;
  wire g1377_p;
  wire g1377_n;
  wire g1378_p;
  wire g1378_n;
  wire g1379_p;
  wire g1379_n;
  wire g1380_p;
  wire g1380_n;
  wire g1381_p;
  wire g1381_n;
  wire g1382_p;
  wire g1382_n;
  wire g1383_p;
  wire g1383_n;
  wire g1384_p;
  wire g1384_n;
  wire g1385_p;
  wire g1385_n;
  wire g1386_p;
  wire g1386_n;
  wire g1387_p;
  wire g1387_n;
  wire g1388_p;
  wire g1388_n;
  wire g1389_p;
  wire g1389_n;
  wire g1390_p;
  wire g1390_n;
  wire g1391_p;
  wire g1391_n;
  wire g1392_p;
  wire g1392_n;
  wire g1393_p;
  wire g1393_n;
  wire g1394_p;
  wire g1394_n;
  wire g1395_p;
  wire g1395_n;
  wire g1396_p;
  wire g1396_n;
  wire g1397_p;
  wire g1397_n;
  wire g1398_p;
  wire g1398_n;
  wire g1399_p;
  wire g1399_n;
  wire g1400_p;
  wire g1400_n;
  wire g1401_p;
  wire g1401_n;
  wire g1402_p;
  wire g1402_n;
  wire g1403_p;
  wire g1403_n;
  wire g1404_p;
  wire g1404_n;
  wire g1405_p;
  wire g1405_n;
  wire g1406_p;
  wire g1406_n;
  wire g1407_p;
  wire g1407_n;
  wire g1408_p;
  wire g1408_n;
  wire g1409_p;
  wire g1409_n;
  wire g1410_p;
  wire g1410_n;
  wire g1411_p;
  wire g1411_n;
  wire g1412_p;
  wire g1412_n;
  wire g1413_p;
  wire g1413_n;
  wire g1414_p;
  wire g1414_n;
  wire g1415_p;
  wire g1415_n;
  wire g1416_p;
  wire g1416_n;
  wire g1417_p;
  wire g1417_n;
  wire g1418_p;
  wire g1418_n;
  wire g1419_p;
  wire g1419_n;
  wire g1420_p;
  wire g1420_n;
  wire g1421_p;
  wire g1421_n;
  wire g1422_p;
  wire g1422_n;
  wire g1423_p;
  wire g1423_n;
  wire g1424_p;
  wire g1424_n;
  wire g1425_p;
  wire g1425_n;
  wire g1426_p;
  wire g1426_n;
  wire g1427_p;
  wire g1427_n;
  wire g1428_p;
  wire g1428_n;
  wire g1429_p;
  wire g1429_n;
  wire g1430_p;
  wire g1430_n;
  wire g1431_p;
  wire g1431_n;
  wire g1432_p;
  wire g1432_n;
  wire g1433_p;
  wire g1433_n;
  wire g1434_p;
  wire g1434_n;
  wire g1435_p;
  wire g1435_n;
  wire g1436_p;
  wire g1436_n;
  wire g1437_p;
  wire g1437_n;
  wire g1438_p;
  wire g1438_n;
  wire g1439_p;
  wire g1439_n;
  wire g1440_p;
  wire g1440_n;
  wire g1441_p;
  wire g1441_n;
  wire g1442_p;
  wire g1442_n;
  wire g1443_p;
  wire g1443_n;
  wire g1444_p;
  wire g1444_n;
  wire g1445_p;
  wire g1445_n;
  wire g1446_p;
  wire g1446_n;
  wire g1447_p;
  wire g1447_n;
  wire g1448_p;
  wire g1448_n;
  wire g1449_p;
  wire g1449_n;
  wire g1450_p;
  wire g1450_n;
  wire g1451_p;
  wire g1451_n;
  wire g1452_p;
  wire g1452_n;
  wire g1453_p;
  wire g1453_n;
  wire g1454_p;
  wire g1454_n;
  wire g1455_p;
  wire g1455_n;
  wire g1456_p;
  wire g1456_n;
  wire g1457_p;
  wire g1457_n;
  wire g1458_p;
  wire g1458_n;
  wire g1459_p;
  wire g1459_n;
  wire g1460_p;
  wire g1460_n;
  wire g1461_p;
  wire g1461_n;
  wire g1462_p;
  wire g1462_n;
  wire g1463_p;
  wire g1463_n;
  wire g1464_p;
  wire g1464_n;
  wire g1465_p;
  wire g1465_n;
  wire g1466_p;
  wire g1466_n;
  wire g1467_p;
  wire g1467_n;
  wire g1468_p;
  wire g1468_n;
  wire g1469_p;
  wire g1469_n;
  wire g1470_p;
  wire g1470_n;
  wire g1471_p;
  wire g1471_n;
  wire g1472_p;
  wire g1472_n;
  wire g1473_p;
  wire g1473_n;
  wire g1474_p;
  wire g1474_n;
  wire g1475_p;
  wire g1475_n;
  wire g1476_p;
  wire g1476_n;
  wire g1477_p;
  wire g1477_n;
  wire g1478_p;
  wire g1478_n;
  wire g1479_p;
  wire g1479_n;
  wire g1480_p;
  wire g1480_n;
  wire g1481_p;
  wire g1481_n;
  wire g1482_p;
  wire g1482_n;
  wire g1483_p;
  wire g1483_n;
  wire g1484_p;
  wire g1484_n;
  wire g1485_p;
  wire g1485_n;
  wire g1486_p;
  wire g1486_n;
  wire g1487_p;
  wire g1487_n;
  wire g1488_p;
  wire g1488_n;
  wire g1489_p;
  wire g1489_n;
  wire g1490_p;
  wire g1490_n;
  wire g1491_p;
  wire g1491_n;
  wire g1492_p;
  wire g1492_n;
  wire g1493_p;
  wire g1493_n;
  wire g1494_p;
  wire g1494_n;
  wire g1495_p;
  wire g1495_n;
  wire g1496_p;
  wire g1496_n;
  wire g1497_p;
  wire g1497_n;
  wire g1498_p;
  wire g1498_n;
  wire g1499_p;
  wire g1499_n;
  wire g1500_p;
  wire g1500_n;
  wire g1501_p;
  wire g1501_n;
  wire g1502_p;
  wire g1502_n;
  wire g1503_p;
  wire g1503_n;
  wire g1504_p;
  wire g1504_n;
  wire g1505_p;
  wire g1505_n;
  wire g1506_p;
  wire g1506_n;
  wire g1507_p;
  wire g1507_n;
  wire g1508_p;
  wire g1508_n;
  wire g1509_p;
  wire g1509_n;
  wire g1510_p;
  wire g1510_n;
  wire g1511_p;
  wire g1511_n;
  wire g1512_p;
  wire g1512_n;
  wire g1513_p;
  wire g1513_n;
  wire g1514_p;
  wire g1514_n;
  wire g1515_p;
  wire g1515_n;
  wire g1516_p;
  wire g1516_n;
  wire g1517_p;
  wire g1517_n;
  wire g1518_p;
  wire g1518_n;
  wire g1519_p;
  wire g1519_n;
  wire g1520_p;
  wire g1520_n;
  wire g1521_p;
  wire g1521_n;
  wire g1522_p;
  wire g1522_n;
  wire g1523_p;
  wire g1523_n;
  wire g1524_p;
  wire g1524_n;
  wire g1525_p;
  wire g1525_n;
  wire g1526_p;
  wire g1526_n;
  wire g1527_p;
  wire g1527_n;
  wire g1528_p;
  wire g1528_n;
  wire g1529_p;
  wire g1529_n;
  wire g1530_p;
  wire g1530_n;
  wire g1531_p;
  wire g1531_n;
  wire g1532_p;
  wire g1532_n;
  wire g1533_p;
  wire g1533_n;
  wire g1534_p;
  wire g1534_n;
  wire g1535_p;
  wire g1535_n;
  wire g1536_p;
  wire g1536_n;
  wire g1537_p;
  wire g1537_n;
  wire g1538_p;
  wire g1538_n;
  wire g1539_p;
  wire g1539_n;
  wire g1540_p;
  wire g1540_n;
  wire g1541_p;
  wire g1541_n;
  wire g1542_p;
  wire g1542_n;
  wire g1543_p;
  wire g1543_n;
  wire g1544_p;
  wire g1544_n;
  wire g1545_p;
  wire g1545_n;
  wire g1546_p;
  wire g1546_n;
  wire g1547_p;
  wire g1547_n;
  wire g1548_p;
  wire g1548_n;
  wire g1549_p;
  wire g1549_n;
  wire g1550_p;
  wire g1550_n;
  wire g1551_p;
  wire g1551_n;
  wire g1552_p;
  wire g1552_n;
  wire g1553_p;
  wire g1553_n;
  wire g1554_p;
  wire g1554_n;
  wire g1555_p;
  wire g1555_n;
  wire g1556_p;
  wire g1556_n;
  wire g1557_p;
  wire g1557_n;
  wire g1558_p;
  wire g1558_n;
  wire g1559_p;
  wire g1559_n;
  wire g1560_p;
  wire g1560_n;
  wire g1561_p;
  wire g1561_n;
  wire g1562_p;
  wire g1562_n;
  wire g1563_p;
  wire g1563_n;
  wire g1564_p;
  wire g1564_n;
  wire g1565_p;
  wire g1565_n;
  wire g1566_p;
  wire g1566_n;
  wire g1567_p;
  wire g1567_n;
  wire g1568_p;
  wire g1568_n;
  wire g1569_p;
  wire g1569_n;
  wire g1570_p;
  wire g1570_n;
  wire g1571_p;
  wire g1571_n;
  wire g1572_p;
  wire g1572_n;
  wire g1573_p;
  wire g1573_n;
  wire g1574_p;
  wire g1574_n;
  wire g1575_p;
  wire g1575_n;
  wire g1576_p;
  wire g1576_n;
  wire g1577_p;
  wire g1577_n;
  wire g1578_p;
  wire g1578_n;
  wire g1579_p;
  wire g1579_n;
  wire g1580_p;
  wire g1580_n;
  wire g1581_p;
  wire g1581_n;
  wire g1582_p;
  wire g1582_n;
  wire g1583_p;
  wire g1583_n;
  wire g1584_p;
  wire g1584_n;
  wire g1585_p;
  wire g1585_n;
  wire g1586_p;
  wire g1586_n;
  wire g1587_p;
  wire g1587_n;
  wire g1588_p;
  wire g1588_n;
  wire g1589_p;
  wire g1589_n;
  wire g1590_p;
  wire g1590_n;
  wire g1591_p;
  wire g1591_n;
  wire g1592_p;
  wire g1592_n;
  wire g1593_p;
  wire g1593_n;
  wire g1594_p;
  wire g1594_n;
  wire g1595_p;
  wire g1595_n;
  wire g1596_p;
  wire g1596_n;
  wire g1597_p;
  wire g1597_n;
  wire g1598_p;
  wire g1598_n;
  wire g1599_p;
  wire g1599_n;
  wire g1600_p;
  wire g1600_n;
  wire g1601_p;
  wire g1601_n;
  wire g1602_p;
  wire g1602_n;
  wire g1603_p;
  wire g1603_n;
  wire g1604_p;
  wire g1604_n;
  wire g1605_p;
  wire g1605_n;
  wire g1606_p;
  wire g1606_n;
  wire g1607_p;
  wire g1607_n;
  wire g1608_p;
  wire g1608_n;
  wire g1609_p;
  wire g1609_n;
  wire g1610_p;
  wire g1610_n;
  wire g1611_p;
  wire g1611_n;
  wire g1612_p;
  wire g1612_n;
  wire g1613_p;
  wire g1613_n;
  wire g1614_p;
  wire g1614_n;
  wire g1615_p;
  wire g1615_n;
  wire g1616_p;
  wire g1616_n;
  wire g1617_p;
  wire g1617_n;
  wire g1618_p;
  wire g1618_n;
  wire g1619_p;
  wire g1619_n;
  wire g1620_p;
  wire g1620_n;
  wire g1621_p;
  wire g1621_n;
  wire g1622_p;
  wire g1622_n;
  wire g1623_p;
  wire g1623_n;
  wire g1624_p;
  wire g1624_n;
  wire g1625_p;
  wire g1625_n;
  wire g1626_p;
  wire g1626_n;
  wire g1627_p;
  wire g1627_n;
  wire g1628_p;
  wire g1628_n;
  wire g1629_p;
  wire g1629_n;
  wire g1630_p;
  wire g1630_n;
  wire g1631_p;
  wire g1631_n;
  wire g1632_p;
  wire g1632_n;
  wire g1633_p;
  wire g1633_n;
  wire g1634_p;
  wire g1634_n;
  wire g1635_p;
  wire g1635_n;
  wire g1636_p;
  wire g1636_n;
  wire g1637_p;
  wire g1637_n;
  wire g1638_p;
  wire g1638_n;
  wire g1639_p;
  wire g1639_n;
  wire g1640_p;
  wire g1640_n;
  wire g1641_p;
  wire g1641_n;
  wire g1642_p;
  wire g1642_n;
  wire g1643_p;
  wire g1643_n;
  wire g1644_p;
  wire g1644_n;
  wire g1645_p;
  wire g1645_n;
  wire g1646_p;
  wire g1646_n;
  wire g1647_p;
  wire g1647_n;
  wire g1648_p;
  wire g1648_n;
  wire g1649_p;
  wire g1649_n;
  wire g1650_p;
  wire g1650_n;
  wire g1651_p;
  wire g1651_n;
  wire g1652_p;
  wire g1652_n;
  wire g1653_p;
  wire g1653_n;
  wire g1654_p;
  wire g1654_n;
  wire g1655_p;
  wire g1655_n;
  wire g1656_p;
  wire g1656_n;
  wire g1657_p;
  wire g1657_n;
  wire g1658_p;
  wire g1658_n;
  wire g1659_p;
  wire g1659_n;
  wire g1660_p;
  wire g1660_n;
  wire g1661_p;
  wire g1661_n;
  wire g1662_p;
  wire g1662_n;
  wire g1663_p;
  wire g1663_n;
  wire g1664_p;
  wire g1664_n;
  wire g1665_p;
  wire g1665_n;
  wire g1666_p;
  wire g1666_n;
  wire g1667_p;
  wire g1667_n;
  wire g1668_p;
  wire g1668_n;
  wire g1669_p;
  wire g1669_n;
  wire g1670_p;
  wire g1670_n;
  wire g1671_p;
  wire g1671_n;
  wire g1672_p;
  wire g1672_n;
  wire g1673_p;
  wire g1673_n;
  wire g1674_p;
  wire g1674_n;
  wire g1675_p;
  wire g1675_n;
  wire g1676_p;
  wire g1676_n;
  wire g1677_p;
  wire g1677_n;
  wire g1678_p;
  wire g1678_n;
  wire g1679_p;
  wire g1679_n;
  wire g1680_p;
  wire g1680_n;
  wire g1681_p;
  wire g1681_n;
  wire g1682_p;
  wire g1682_n;
  wire g1683_p;
  wire g1683_n;
  wire g1684_p;
  wire g1684_n;
  wire g1685_p;
  wire g1685_n;
  wire g1686_p;
  wire g1686_n;
  wire g1687_p;
  wire g1687_n;
  wire g1688_p;
  wire g1688_n;
  wire g1689_p;
  wire g1689_n;
  wire g1690_p;
  wire g1690_n;
  wire g1691_p;
  wire g1691_n;
  wire g1692_p;
  wire g1692_n;
  wire g1693_p;
  wire g1693_n;
  wire g1694_p;
  wire g1694_n;
  wire g1695_p;
  wire g1695_n;
  wire g1696_p;
  wire g1696_n;
  wire g1697_p;
  wire g1697_n;
  wire g1698_p;
  wire g1698_n;
  wire g1699_p;
  wire g1699_n;
  wire g1700_p;
  wire g1700_n;
  wire g1701_p;
  wire g1701_n;
  wire g1702_p;
  wire g1702_n;
  wire g1703_p;
  wire g1703_n;
  wire g1704_p;
  wire g1704_n;
  wire g1705_p;
  wire g1705_n;
  wire g1706_p;
  wire g1706_n;
  wire g1707_p;
  wire g1707_n;
  wire g1708_p;
  wire g1708_n;
  wire g1709_p;
  wire g1709_n;
  wire g1710_p;
  wire g1710_n;
  wire g1711_p;
  wire g1711_n;
  wire g1712_p;
  wire g1712_n;
  wire g1713_p;
  wire g1713_n;
  wire g1714_p;
  wire g1714_n;
  wire g1715_p;
  wire g1715_n;
  wire g1716_p;
  wire g1716_n;
  wire g1717_p;
  wire g1717_n;
  wire g1718_p;
  wire g1718_n;
  wire g1719_p;
  wire g1719_n;
  wire g1720_p;
  wire g1720_n;
  wire g1721_p;
  wire g1721_n;
  wire g1722_p;
  wire g1722_n;
  wire g1723_p;
  wire g1723_n;
  wire g1724_p;
  wire g1724_n;
  wire g1725_p;
  wire g1725_n;
  wire g1726_p;
  wire g1726_n;
  wire g1727_p;
  wire g1727_n;
  wire g1728_p;
  wire g1728_n;
  wire g1729_p;
  wire g1729_n;
  wire g1730_p;
  wire g1730_n;
  wire g1731_p;
  wire g1731_n;
  wire g1732_p;
  wire g1732_n;
  wire g1733_p;
  wire g1733_n;
  wire g1734_p;
  wire g1734_n;
  wire g1735_p;
  wire g1735_n;
  wire g1736_p;
  wire g1736_n;
  wire g1737_p;
  wire g1737_n;
  wire g1738_p;
  wire g1738_n;
  wire g1739_p;
  wire g1739_n;
  wire g1740_p;
  wire g1740_n;
  wire g1741_p;
  wire g1741_n;
  wire g1742_p;
  wire g1742_n;
  wire g1743_p;
  wire g1743_n;
  wire g1744_p;
  wire g1744_n;
  wire g1745_p;
  wire g1745_n;
  wire g1746_p;
  wire g1746_n;
  wire g1747_p;
  wire g1747_n;
  wire g1748_p;
  wire g1748_n;
  wire g1749_p;
  wire g1749_n;
  wire g1750_p;
  wire g1750_n;
  wire g1751_p;
  wire g1751_n;
  wire g1752_p;
  wire g1752_n;
  wire g1753_p;
  wire g1753_n;
  wire g1754_p;
  wire g1754_n;
  wire g1755_p;
  wire g1755_n;
  wire g1756_p;
  wire g1756_n;
  wire g1757_p;
  wire g1757_n;
  wire g1758_p;
  wire g1758_n;
  wire g1759_p;
  wire g1759_n;
  wire g1760_p;
  wire g1760_n;
  wire g1761_p;
  wire g1761_n;
  wire g1762_p;
  wire g1762_n;
  wire g1763_p;
  wire g1763_n;
  wire g1764_p;
  wire g1764_n;
  wire g1765_p;
  wire g1765_n;
  wire g1766_p;
  wire g1766_n;
  wire g1767_p;
  wire g1767_n;
  wire g1768_p;
  wire g1768_n;
  wire g1769_p;
  wire g1769_n;
  wire g1770_p;
  wire g1770_n;
  wire g1771_p;
  wire g1771_n;
  wire g1772_p;
  wire g1772_n;
  wire g1773_p;
  wire g1773_n;
  wire g1774_p;
  wire g1774_n;
  wire g1775_p;
  wire g1775_n;
  wire g1776_p;
  wire g1776_n;
  wire g1777_p;
  wire g1777_n;
  wire g1778_p;
  wire g1778_n;
  wire g1779_p;
  wire g1779_n;
  wire g1780_p;
  wire g1780_n;
  wire g1781_p;
  wire g1781_n;
  wire g1782_p;
  wire g1782_n;
  wire g1783_p;
  wire g1783_n;
  wire g1784_p;
  wire g1784_n;
  wire g1785_p;
  wire g1785_n;
  wire g1786_p;
  wire g1786_n;
  wire g1787_p;
  wire g1787_n;
  wire g1788_p;
  wire g1788_n;
  wire g1789_p;
  wire g1789_n;
  wire g1790_p;
  wire g1790_n;
  wire g1791_p;
  wire g1791_n;
  wire g1792_p;
  wire g1792_n;
  wire g1793_p;
  wire g1793_n;
  wire g1794_p;
  wire g1794_n;
  wire g1795_p;
  wire g1795_n;
  wire g1796_p;
  wire g1796_n;
  wire g1797_p;
  wire g1797_n;
  wire g1798_p;
  wire g1798_n;
  wire g1799_p;
  wire g1799_n;
  wire g1800_p;
  wire g1800_n;
  wire g1801_p;
  wire g1801_n;
  wire g1802_p;
  wire g1802_n;
  wire g1803_p;
  wire g1803_n;
  wire g1804_p;
  wire g1804_n;
  wire g1805_p;
  wire g1805_n;
  wire g1806_p;
  wire g1806_n;
  wire g1807_p;
  wire g1807_n;
  wire g1808_p;
  wire g1808_n;
  wire g1809_p;
  wire g1809_n;
  wire g1810_p;
  wire g1810_n;
  wire g1811_p;
  wire g1811_n;
  wire g1812_p;
  wire g1812_n;
  wire g1813_p;
  wire g1813_n;
  wire g1814_p;
  wire g1814_n;
  wire g1815_p;
  wire g1815_n;
  wire g1816_p;
  wire g1816_n;
  wire g1817_p;
  wire g1817_n;
  wire g1818_p;
  wire g1818_n;
  wire g1819_p;
  wire g1819_n;
  wire g1820_p;
  wire g1820_n;
  wire g1821_p;
  wire g1821_n;
  wire g1822_p;
  wire g1822_n;
  wire g1823_p;
  wire g1823_n;
  wire g1824_p;
  wire g1824_n;
  wire g1825_p;
  wire g1825_n;
  wire g1826_p;
  wire g1826_n;
  wire g1827_p;
  wire g1827_n;
  wire g1828_p;
  wire g1828_n;
  wire g1829_p;
  wire g1829_n;
  wire g1830_p;
  wire g1830_n;
  wire g1831_p;
  wire g1831_n;
  wire g1832_p;
  wire g1832_n;
  wire g1833_p;
  wire g1833_n;
  wire g1834_p;
  wire g1834_n;
  wire g1835_p;
  wire g1835_n;
  wire g1836_p;
  wire g1836_n;
  wire g1837_p;
  wire g1837_n;
  wire g1838_p;
  wire g1838_n;
  wire g1839_p;
  wire g1839_n;
  wire g1840_p;
  wire g1840_n;
  wire g1841_p;
  wire g1841_n;
  wire g1842_p;
  wire g1842_n;
  wire g1843_p;
  wire g1843_n;
  wire g1844_p;
  wire g1844_n;
  wire g1845_p;
  wire g1845_n;
  wire g1846_p;
  wire g1846_n;
  wire g1847_p;
  wire g1847_n;
  wire g1848_p;
  wire g1848_n;
  wire g1849_p;
  wire g1849_n;
  wire g1850_p;
  wire g1850_n;
  wire g1851_p;
  wire g1851_n;
  wire g1852_p;
  wire g1852_n;
  wire g1853_p;
  wire g1853_n;
  wire g1854_p;
  wire g1854_n;
  wire g1855_p;
  wire g1855_n;
  wire g1856_p;
  wire g1856_n;
  wire g1857_p;
  wire g1857_n;
  wire g1858_p;
  wire g1858_n;
  wire g1859_p;
  wire g1859_n;
  wire g1860_p;
  wire g1860_n;
  wire g1861_p;
  wire g1861_n;
  wire g1862_p;
  wire g1862_n;
  wire g1863_p;
  wire g1863_n;
  wire g1864_p;
  wire g1864_n;
  wire g1865_p;
  wire g1865_n;
  wire g1866_p;
  wire g1866_n;
  wire g1867_p;
  wire g1867_n;
  wire g1868_p;
  wire g1868_n;
  wire g1869_p;
  wire g1869_n;
  wire g1870_p;
  wire g1870_n;
  wire g1871_p;
  wire g1871_n;
  wire g1872_p;
  wire g1872_n;
  wire g1873_p;
  wire g1873_n;
  wire g1874_p;
  wire g1874_n;
  wire g1875_p;
  wire g1875_n;
  wire g1876_p;
  wire g1876_n;
  wire g1877_p;
  wire g1877_n;
  wire g1878_p;
  wire g1878_n;
  wire g1879_p;
  wire g1879_n;
  wire g1880_p;
  wire g1880_n;
  wire g1881_p;
  wire g1881_n;
  wire g1882_p;
  wire g1882_n;
  wire g1883_p;
  wire g1883_n;
  wire g1884_p;
  wire g1884_n;
  wire g1885_p;
  wire g1885_n;
  wire g1886_p;
  wire g1886_n;
  wire g1887_p;
  wire g1887_n;
  wire g1888_p;
  wire g1888_n;
  wire g1889_p;
  wire g1889_n;
  wire g1890_p;
  wire g1890_n;
  wire g1891_p;
  wire g1891_n;
  wire g1892_p;
  wire g1892_n;
  wire g1893_p;
  wire g1893_n;
  wire g1894_p;
  wire g1894_n;
  wire g1895_p;
  wire g1895_n;
  wire g1896_p;
  wire g1896_n;
  wire g1897_p;
  wire g1897_n;
  wire g1898_p;
  wire g1898_n;
  wire g1899_p;
  wire g1899_n;
  wire g1900_p;
  wire g1900_n;
  wire g1901_p;
  wire g1901_n;
  wire g1902_p;
  wire g1902_n;
  wire g1903_p;
  wire g1903_n;
  wire g1904_p;
  wire g1904_n;
  wire g1905_p;
  wire g1905_n;
  wire g1906_p;
  wire g1906_n;
  wire g1907_p;
  wire g1907_n;
  wire g1908_p;
  wire g1908_n;
  wire g1909_p;
  wire g1909_n;
  wire g1910_p;
  wire g1910_n;
  wire g1911_p;
  wire g1911_n;
  wire g1912_p;
  wire g1912_n;
  wire g1913_p;
  wire g1913_n;
  wire g1914_p;
  wire g1914_n;
  wire g1915_p;
  wire g1915_n;
  wire g1916_p;
  wire g1916_n;
  wire g1917_p;
  wire g1917_n;
  wire G1_p_spl_;
  wire G1_p_spl_0;
  wire G1_p_spl_00;
  wire G1_p_spl_000;
  wire G1_p_spl_001;
  wire G1_p_spl_01;
  wire G1_p_spl_010;
  wire G1_p_spl_011;
  wire G1_p_spl_1;
  wire G1_p_spl_10;
  wire G1_p_spl_100;
  wire G1_p_spl_101;
  wire G1_p_spl_11;
  wire G1_p_spl_110;
  wire G1_p_spl_111;
  wire G17_p_spl_;
  wire G17_p_spl_0;
  wire G17_p_spl_00;
  wire G17_p_spl_000;
  wire G17_p_spl_001;
  wire G17_p_spl_01;
  wire G17_p_spl_010;
  wire G17_p_spl_011;
  wire G17_p_spl_1;
  wire G17_p_spl_10;
  wire G17_p_spl_100;
  wire G17_p_spl_101;
  wire G17_p_spl_11;
  wire G17_p_spl_110;
  wire G17_p_spl_111;
  wire G2_p_spl_;
  wire G2_p_spl_0;
  wire G2_p_spl_00;
  wire G2_p_spl_000;
  wire G2_p_spl_001;
  wire G2_p_spl_01;
  wire G2_p_spl_010;
  wire G2_p_spl_011;
  wire G2_p_spl_1;
  wire G2_p_spl_10;
  wire G2_p_spl_100;
  wire G2_p_spl_101;
  wire G2_p_spl_11;
  wire G2_p_spl_110;
  wire G2_p_spl_111;
  wire G2_n_spl_;
  wire G2_n_spl_0;
  wire G2_n_spl_00;
  wire G2_n_spl_000;
  wire G2_n_spl_001;
  wire G2_n_spl_01;
  wire G2_n_spl_010;
  wire G2_n_spl_011;
  wire G2_n_spl_1;
  wire G2_n_spl_10;
  wire G2_n_spl_100;
  wire G2_n_spl_101;
  wire G2_n_spl_11;
  wire G2_n_spl_110;
  wire G2_n_spl_111;
  wire G17_n_spl_;
  wire G17_n_spl_0;
  wire G17_n_spl_00;
  wire G17_n_spl_000;
  wire G17_n_spl_001;
  wire G17_n_spl_01;
  wire G17_n_spl_010;
  wire G17_n_spl_011;
  wire G17_n_spl_1;
  wire G17_n_spl_10;
  wire G17_n_spl_100;
  wire G17_n_spl_101;
  wire G17_n_spl_11;
  wire G17_n_spl_110;
  wire G18_p_spl_;
  wire G18_p_spl_0;
  wire G18_p_spl_00;
  wire G18_p_spl_000;
  wire G18_p_spl_001;
  wire G18_p_spl_01;
  wire G18_p_spl_010;
  wire G18_p_spl_011;
  wire G18_p_spl_1;
  wire G18_p_spl_10;
  wire G18_p_spl_100;
  wire G18_p_spl_101;
  wire G18_p_spl_11;
  wire G18_p_spl_110;
  wire G18_p_spl_111;
  wire G1_n_spl_;
  wire G1_n_spl_0;
  wire G1_n_spl_00;
  wire G1_n_spl_000;
  wire G1_n_spl_001;
  wire G1_n_spl_01;
  wire G1_n_spl_010;
  wire G1_n_spl_011;
  wire G1_n_spl_1;
  wire G1_n_spl_10;
  wire G1_n_spl_100;
  wire G1_n_spl_101;
  wire G1_n_spl_11;
  wire G1_n_spl_110;
  wire G18_n_spl_;
  wire G18_n_spl_0;
  wire G18_n_spl_00;
  wire G18_n_spl_000;
  wire G18_n_spl_001;
  wire G18_n_spl_01;
  wire G18_n_spl_010;
  wire G18_n_spl_011;
  wire G18_n_spl_1;
  wire G18_n_spl_10;
  wire G18_n_spl_100;
  wire G18_n_spl_101;
  wire G18_n_spl_11;
  wire G18_n_spl_110;
  wire G18_n_spl_111;
  wire g34_p_spl_;
  wire g34_n_spl_;
  wire g35_p_spl_;
  wire g36_p_spl_;
  wire g37_n_spl_;
  wire g37_n_spl_0;
  wire G19_p_spl_;
  wire G19_p_spl_0;
  wire G19_p_spl_00;
  wire G19_p_spl_000;
  wire G19_p_spl_001;
  wire G19_p_spl_01;
  wire G19_p_spl_010;
  wire G19_p_spl_011;
  wire G19_p_spl_1;
  wire G19_p_spl_10;
  wire G19_p_spl_100;
  wire G19_p_spl_101;
  wire G19_p_spl_11;
  wire G19_p_spl_110;
  wire G19_p_spl_111;
  wire G19_n_spl_;
  wire G19_n_spl_0;
  wire G19_n_spl_00;
  wire G19_n_spl_000;
  wire G19_n_spl_001;
  wire G19_n_spl_01;
  wire G19_n_spl_010;
  wire G19_n_spl_011;
  wire G19_n_spl_1;
  wire G19_n_spl_10;
  wire G19_n_spl_100;
  wire G19_n_spl_101;
  wire G19_n_spl_11;
  wire G19_n_spl_110;
  wire G19_n_spl_111;
  wire G3_p_spl_;
  wire G3_p_spl_0;
  wire G3_p_spl_00;
  wire G3_p_spl_000;
  wire G3_p_spl_001;
  wire G3_p_spl_01;
  wire G3_p_spl_010;
  wire G3_p_spl_011;
  wire G3_p_spl_1;
  wire G3_p_spl_10;
  wire G3_p_spl_100;
  wire G3_p_spl_101;
  wire G3_p_spl_11;
  wire G3_p_spl_110;
  wire G3_p_spl_111;
  wire G3_n_spl_;
  wire G3_n_spl_0;
  wire G3_n_spl_00;
  wire G3_n_spl_000;
  wire G3_n_spl_001;
  wire G3_n_spl_01;
  wire G3_n_spl_010;
  wire G3_n_spl_011;
  wire G3_n_spl_1;
  wire G3_n_spl_10;
  wire G3_n_spl_100;
  wire G3_n_spl_101;
  wire G3_n_spl_11;
  wire G3_n_spl_110;
  wire G3_n_spl_111;
  wire g41_p_spl_;
  wire g42_n_spl_;
  wire g41_n_spl_;
  wire g42_p_spl_;
  wire g43_n_spl_;
  wire g43_p_spl_;
  wire g44_n_spl_;
  wire g44_n_spl_0;
  wire g44_p_spl_;
  wire g44_p_spl_0;
  wire g46_n_spl_;
  wire g37_p_spl_;
  wire g46_p_spl_;
  wire g47_n_spl_;
  wire g47_p_spl_;
  wire g40_p_spl_;
  wire g49_n_spl_;
  wire g50_p_spl_;
  wire G20_p_spl_;
  wire G20_p_spl_0;
  wire G20_p_spl_00;
  wire G20_p_spl_000;
  wire G20_p_spl_001;
  wire G20_p_spl_01;
  wire G20_p_spl_010;
  wire G20_p_spl_011;
  wire G20_p_spl_1;
  wire G20_p_spl_10;
  wire G20_p_spl_100;
  wire G20_p_spl_101;
  wire G20_p_spl_11;
  wire G20_p_spl_110;
  wire G20_p_spl_111;
  wire G20_n_spl_;
  wire G20_n_spl_0;
  wire G20_n_spl_00;
  wire G20_n_spl_000;
  wire G20_n_spl_001;
  wire G20_n_spl_01;
  wire G20_n_spl_010;
  wire G20_n_spl_011;
  wire G20_n_spl_1;
  wire G20_n_spl_10;
  wire G20_n_spl_100;
  wire G20_n_spl_101;
  wire G20_n_spl_11;
  wire G20_n_spl_110;
  wire G20_n_spl_111;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_00;
  wire G4_p_spl_000;
  wire G4_p_spl_001;
  wire G4_p_spl_01;
  wire G4_p_spl_010;
  wire G4_p_spl_011;
  wire G4_p_spl_1;
  wire G4_p_spl_10;
  wire G4_p_spl_100;
  wire G4_p_spl_101;
  wire G4_p_spl_11;
  wire G4_p_spl_110;
  wire G4_p_spl_111;
  wire G4_n_spl_;
  wire G4_n_spl_0;
  wire G4_n_spl_00;
  wire G4_n_spl_000;
  wire G4_n_spl_001;
  wire G4_n_spl_01;
  wire G4_n_spl_010;
  wire G4_n_spl_011;
  wire G4_n_spl_1;
  wire G4_n_spl_10;
  wire G4_n_spl_100;
  wire G4_n_spl_101;
  wire G4_n_spl_11;
  wire G4_n_spl_110;
  wire G4_n_spl_111;
  wire g56_p_spl_;
  wire g57_n_spl_;
  wire g56_n_spl_;
  wire g57_p_spl_;
  wire g58_n_spl_;
  wire g58_p_spl_;
  wire g59_n_spl_;
  wire g59_n_spl_0;
  wire g59_p_spl_;
  wire g59_p_spl_0;
  wire g61_n_spl_;
  wire g61_p_spl_;
  wire g62_n_spl_;
  wire g62_p_spl_;
  wire g55_n_spl_;
  wire g64_p_spl_;
  wire g55_p_spl_;
  wire g64_n_spl_;
  wire g65_n_spl_;
  wire g65_p_spl_;
  wire g54_n_spl_;
  wire g67_p_spl_;
  wire g54_p_spl_;
  wire g67_n_spl_;
  wire g68_n_spl_;
  wire g68_p_spl_;
  wire g53_p_spl_;
  wire g70_n_spl_;
  wire g71_p_spl_;
  wire G21_p_spl_;
  wire G21_p_spl_0;
  wire G21_p_spl_00;
  wire G21_p_spl_000;
  wire G21_p_spl_001;
  wire G21_p_spl_01;
  wire G21_p_spl_010;
  wire G21_p_spl_011;
  wire G21_p_spl_1;
  wire G21_p_spl_10;
  wire G21_p_spl_100;
  wire G21_p_spl_101;
  wire G21_p_spl_11;
  wire G21_p_spl_110;
  wire G21_p_spl_111;
  wire G21_n_spl_;
  wire G21_n_spl_0;
  wire G21_n_spl_00;
  wire G21_n_spl_000;
  wire G21_n_spl_001;
  wire G21_n_spl_01;
  wire G21_n_spl_010;
  wire G21_n_spl_011;
  wire G21_n_spl_1;
  wire G21_n_spl_10;
  wire G21_n_spl_100;
  wire G21_n_spl_101;
  wire G21_n_spl_11;
  wire G21_n_spl_110;
  wire G21_n_spl_111;
  wire G5_p_spl_;
  wire G5_p_spl_0;
  wire G5_p_spl_00;
  wire G5_p_spl_000;
  wire G5_p_spl_001;
  wire G5_p_spl_01;
  wire G5_p_spl_010;
  wire G5_p_spl_011;
  wire G5_p_spl_1;
  wire G5_p_spl_10;
  wire G5_p_spl_100;
  wire G5_p_spl_101;
  wire G5_p_spl_11;
  wire G5_p_spl_110;
  wire G5_p_spl_111;
  wire G5_n_spl_;
  wire G5_n_spl_0;
  wire G5_n_spl_00;
  wire G5_n_spl_000;
  wire G5_n_spl_001;
  wire G5_n_spl_01;
  wire G5_n_spl_010;
  wire G5_n_spl_011;
  wire G5_n_spl_1;
  wire G5_n_spl_10;
  wire G5_n_spl_100;
  wire G5_n_spl_101;
  wire G5_n_spl_11;
  wire G5_n_spl_110;
  wire G5_n_spl_111;
  wire g79_p_spl_;
  wire g80_n_spl_;
  wire g79_n_spl_;
  wire g80_p_spl_;
  wire g81_n_spl_;
  wire g81_p_spl_;
  wire g82_n_spl_;
  wire g82_n_spl_0;
  wire g82_p_spl_;
  wire g82_p_spl_0;
  wire g84_n_spl_;
  wire g84_p_spl_;
  wire g85_n_spl_;
  wire g85_p_spl_;
  wire g78_n_spl_;
  wire g87_p_spl_;
  wire g78_p_spl_;
  wire g87_n_spl_;
  wire g88_n_spl_;
  wire g88_p_spl_;
  wire g77_n_spl_;
  wire g90_p_spl_;
  wire g77_p_spl_;
  wire g90_n_spl_;
  wire g91_n_spl_;
  wire g91_p_spl_;
  wire g76_n_spl_;
  wire g93_p_spl_;
  wire g76_p_spl_;
  wire g93_n_spl_;
  wire g94_n_spl_;
  wire g94_p_spl_;
  wire g75_n_spl_;
  wire g96_p_spl_;
  wire g75_p_spl_;
  wire g96_n_spl_;
  wire g97_n_spl_;
  wire g97_p_spl_;
  wire g74_p_spl_;
  wire g99_n_spl_;
  wire g100_p_spl_;
  wire G22_p_spl_;
  wire G22_p_spl_0;
  wire G22_p_spl_00;
  wire G22_p_spl_000;
  wire G22_p_spl_001;
  wire G22_p_spl_01;
  wire G22_p_spl_010;
  wire G22_p_spl_011;
  wire G22_p_spl_1;
  wire G22_p_spl_10;
  wire G22_p_spl_100;
  wire G22_p_spl_101;
  wire G22_p_spl_11;
  wire G22_p_spl_110;
  wire G22_p_spl_111;
  wire G22_n_spl_;
  wire G22_n_spl_0;
  wire G22_n_spl_00;
  wire G22_n_spl_000;
  wire G22_n_spl_001;
  wire G22_n_spl_01;
  wire G22_n_spl_010;
  wire G22_n_spl_011;
  wire G22_n_spl_1;
  wire G22_n_spl_10;
  wire G22_n_spl_100;
  wire G22_n_spl_101;
  wire G22_n_spl_11;
  wire G22_n_spl_110;
  wire G22_n_spl_111;
  wire G6_p_spl_;
  wire G6_p_spl_0;
  wire G6_p_spl_00;
  wire G6_p_spl_000;
  wire G6_p_spl_001;
  wire G6_p_spl_01;
  wire G6_p_spl_010;
  wire G6_p_spl_011;
  wire G6_p_spl_1;
  wire G6_p_spl_10;
  wire G6_p_spl_100;
  wire G6_p_spl_101;
  wire G6_p_spl_11;
  wire G6_p_spl_110;
  wire G6_p_spl_111;
  wire G6_n_spl_;
  wire G6_n_spl_0;
  wire G6_n_spl_00;
  wire G6_n_spl_000;
  wire G6_n_spl_001;
  wire G6_n_spl_01;
  wire G6_n_spl_010;
  wire G6_n_spl_011;
  wire G6_n_spl_1;
  wire G6_n_spl_10;
  wire G6_n_spl_100;
  wire G6_n_spl_101;
  wire G6_n_spl_11;
  wire G6_n_spl_110;
  wire G6_n_spl_111;
  wire g110_p_spl_;
  wire g111_n_spl_;
  wire g110_n_spl_;
  wire g111_p_spl_;
  wire g112_n_spl_;
  wire g112_p_spl_;
  wire g113_n_spl_;
  wire g113_n_spl_0;
  wire g113_p_spl_;
  wire g113_p_spl_0;
  wire g115_n_spl_;
  wire g115_p_spl_;
  wire g116_n_spl_;
  wire g116_p_spl_;
  wire g109_n_spl_;
  wire g118_p_spl_;
  wire g109_p_spl_;
  wire g118_n_spl_;
  wire g119_n_spl_;
  wire g119_p_spl_;
  wire g108_n_spl_;
  wire g121_p_spl_;
  wire g108_p_spl_;
  wire g121_n_spl_;
  wire g122_n_spl_;
  wire g122_p_spl_;
  wire g107_n_spl_;
  wire g124_p_spl_;
  wire g107_p_spl_;
  wire g124_n_spl_;
  wire g125_n_spl_;
  wire g125_p_spl_;
  wire g106_n_spl_;
  wire g127_p_spl_;
  wire g106_p_spl_;
  wire g127_n_spl_;
  wire g128_n_spl_;
  wire g128_p_spl_;
  wire g105_n_spl_;
  wire g130_p_spl_;
  wire g105_p_spl_;
  wire g130_n_spl_;
  wire g131_n_spl_;
  wire g131_p_spl_;
  wire g104_n_spl_;
  wire g133_p_spl_;
  wire g104_p_spl_;
  wire g133_n_spl_;
  wire g134_n_spl_;
  wire g134_p_spl_;
  wire g103_p_spl_;
  wire g136_n_spl_;
  wire g137_p_spl_;
  wire G23_p_spl_;
  wire G23_p_spl_0;
  wire G23_p_spl_00;
  wire G23_p_spl_000;
  wire G23_p_spl_001;
  wire G23_p_spl_01;
  wire G23_p_spl_010;
  wire G23_p_spl_011;
  wire G23_p_spl_1;
  wire G23_p_spl_10;
  wire G23_p_spl_100;
  wire G23_p_spl_101;
  wire G23_p_spl_11;
  wire G23_p_spl_110;
  wire G23_p_spl_111;
  wire G23_n_spl_;
  wire G23_n_spl_0;
  wire G23_n_spl_00;
  wire G23_n_spl_000;
  wire G23_n_spl_001;
  wire G23_n_spl_01;
  wire G23_n_spl_010;
  wire G23_n_spl_011;
  wire G23_n_spl_1;
  wire G23_n_spl_10;
  wire G23_n_spl_100;
  wire G23_n_spl_101;
  wire G23_n_spl_11;
  wire G23_n_spl_110;
  wire G23_n_spl_111;
  wire G7_p_spl_;
  wire G7_p_spl_0;
  wire G7_p_spl_00;
  wire G7_p_spl_000;
  wire G7_p_spl_001;
  wire G7_p_spl_01;
  wire G7_p_spl_010;
  wire G7_p_spl_011;
  wire G7_p_spl_1;
  wire G7_p_spl_10;
  wire G7_p_spl_100;
  wire G7_p_spl_101;
  wire G7_p_spl_11;
  wire G7_p_spl_110;
  wire G7_p_spl_111;
  wire G7_n_spl_;
  wire G7_n_spl_0;
  wire G7_n_spl_00;
  wire G7_n_spl_000;
  wire G7_n_spl_001;
  wire G7_n_spl_01;
  wire G7_n_spl_010;
  wire G7_n_spl_011;
  wire G7_n_spl_1;
  wire G7_n_spl_10;
  wire G7_n_spl_100;
  wire G7_n_spl_101;
  wire G7_n_spl_11;
  wire G7_n_spl_110;
  wire G7_n_spl_111;
  wire g149_p_spl_;
  wire g150_n_spl_;
  wire g149_n_spl_;
  wire g150_p_spl_;
  wire g151_n_spl_;
  wire g151_p_spl_;
  wire g152_n_spl_;
  wire g152_n_spl_0;
  wire g152_p_spl_;
  wire g152_p_spl_0;
  wire g154_n_spl_;
  wire g154_p_spl_;
  wire g155_n_spl_;
  wire g155_p_spl_;
  wire g148_n_spl_;
  wire g157_p_spl_;
  wire g148_p_spl_;
  wire g157_n_spl_;
  wire g158_n_spl_;
  wire g158_p_spl_;
  wire g147_n_spl_;
  wire g160_p_spl_;
  wire g147_p_spl_;
  wire g160_n_spl_;
  wire g161_n_spl_;
  wire g161_p_spl_;
  wire g146_n_spl_;
  wire g163_p_spl_;
  wire g146_p_spl_;
  wire g163_n_spl_;
  wire g164_n_spl_;
  wire g164_p_spl_;
  wire g145_n_spl_;
  wire g166_p_spl_;
  wire g145_p_spl_;
  wire g166_n_spl_;
  wire g167_n_spl_;
  wire g167_p_spl_;
  wire g144_n_spl_;
  wire g169_p_spl_;
  wire g144_p_spl_;
  wire g169_n_spl_;
  wire g170_n_spl_;
  wire g170_p_spl_;
  wire g143_n_spl_;
  wire g172_p_spl_;
  wire g143_p_spl_;
  wire g172_n_spl_;
  wire g173_n_spl_;
  wire g173_p_spl_;
  wire g142_n_spl_;
  wire g175_p_spl_;
  wire g142_p_spl_;
  wire g175_n_spl_;
  wire g176_n_spl_;
  wire g176_p_spl_;
  wire g141_n_spl_;
  wire g178_p_spl_;
  wire g141_p_spl_;
  wire g178_n_spl_;
  wire g179_n_spl_;
  wire g179_p_spl_;
  wire g140_p_spl_;
  wire g181_n_spl_;
  wire g182_p_spl_;
  wire G24_p_spl_;
  wire G24_p_spl_0;
  wire G24_p_spl_00;
  wire G24_p_spl_000;
  wire G24_p_spl_001;
  wire G24_p_spl_01;
  wire G24_p_spl_010;
  wire G24_p_spl_011;
  wire G24_p_spl_1;
  wire G24_p_spl_10;
  wire G24_p_spl_100;
  wire G24_p_spl_101;
  wire G24_p_spl_11;
  wire G24_p_spl_110;
  wire G24_p_spl_111;
  wire G24_n_spl_;
  wire G24_n_spl_0;
  wire G24_n_spl_00;
  wire G24_n_spl_000;
  wire G24_n_spl_001;
  wire G24_n_spl_01;
  wire G24_n_spl_010;
  wire G24_n_spl_011;
  wire G24_n_spl_1;
  wire G24_n_spl_10;
  wire G24_n_spl_100;
  wire G24_n_spl_101;
  wire G24_n_spl_11;
  wire G24_n_spl_110;
  wire G24_n_spl_111;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire G8_p_spl_00;
  wire G8_p_spl_000;
  wire G8_p_spl_001;
  wire G8_p_spl_01;
  wire G8_p_spl_010;
  wire G8_p_spl_011;
  wire G8_p_spl_1;
  wire G8_p_spl_10;
  wire G8_p_spl_100;
  wire G8_p_spl_101;
  wire G8_p_spl_11;
  wire G8_p_spl_110;
  wire G8_p_spl_111;
  wire G8_n_spl_;
  wire G8_n_spl_0;
  wire G8_n_spl_00;
  wire G8_n_spl_000;
  wire G8_n_spl_001;
  wire G8_n_spl_01;
  wire G8_n_spl_010;
  wire G8_n_spl_011;
  wire G8_n_spl_1;
  wire G8_n_spl_10;
  wire G8_n_spl_100;
  wire G8_n_spl_101;
  wire G8_n_spl_11;
  wire G8_n_spl_110;
  wire G8_n_spl_111;
  wire g196_p_spl_;
  wire g197_n_spl_;
  wire g196_n_spl_;
  wire g197_p_spl_;
  wire g198_n_spl_;
  wire g198_p_spl_;
  wire g199_n_spl_;
  wire g199_n_spl_0;
  wire g199_p_spl_;
  wire g199_p_spl_0;
  wire g201_n_spl_;
  wire g201_p_spl_;
  wire g202_n_spl_;
  wire g202_p_spl_;
  wire g195_n_spl_;
  wire g204_p_spl_;
  wire g195_p_spl_;
  wire g204_n_spl_;
  wire g205_n_spl_;
  wire g205_p_spl_;
  wire g194_n_spl_;
  wire g207_p_spl_;
  wire g194_p_spl_;
  wire g207_n_spl_;
  wire g208_n_spl_;
  wire g208_p_spl_;
  wire g193_n_spl_;
  wire g210_p_spl_;
  wire g193_p_spl_;
  wire g210_n_spl_;
  wire g211_n_spl_;
  wire g211_p_spl_;
  wire g192_n_spl_;
  wire g213_p_spl_;
  wire g192_p_spl_;
  wire g213_n_spl_;
  wire g214_n_spl_;
  wire g214_p_spl_;
  wire g191_n_spl_;
  wire g216_p_spl_;
  wire g191_p_spl_;
  wire g216_n_spl_;
  wire g217_n_spl_;
  wire g217_p_spl_;
  wire g190_n_spl_;
  wire g219_p_spl_;
  wire g190_p_spl_;
  wire g219_n_spl_;
  wire g220_n_spl_;
  wire g220_p_spl_;
  wire g189_n_spl_;
  wire g222_p_spl_;
  wire g189_p_spl_;
  wire g222_n_spl_;
  wire g223_n_spl_;
  wire g223_p_spl_;
  wire g188_n_spl_;
  wire g225_p_spl_;
  wire g188_p_spl_;
  wire g225_n_spl_;
  wire g226_n_spl_;
  wire g226_p_spl_;
  wire g187_n_spl_;
  wire g228_p_spl_;
  wire g187_p_spl_;
  wire g228_n_spl_;
  wire g229_n_spl_;
  wire g229_p_spl_;
  wire g186_n_spl_;
  wire g231_p_spl_;
  wire g186_p_spl_;
  wire g231_n_spl_;
  wire g232_n_spl_;
  wire g232_p_spl_;
  wire g185_p_spl_;
  wire g234_n_spl_;
  wire g235_p_spl_;
  wire G25_p_spl_;
  wire G25_p_spl_0;
  wire G25_p_spl_00;
  wire G25_p_spl_000;
  wire G25_p_spl_001;
  wire G25_p_spl_01;
  wire G25_p_spl_010;
  wire G25_p_spl_011;
  wire G25_p_spl_1;
  wire G25_p_spl_10;
  wire G25_p_spl_100;
  wire G25_p_spl_101;
  wire G25_p_spl_11;
  wire G25_p_spl_110;
  wire G25_p_spl_111;
  wire G25_n_spl_;
  wire G25_n_spl_0;
  wire G25_n_spl_00;
  wire G25_n_spl_000;
  wire G25_n_spl_001;
  wire G25_n_spl_01;
  wire G25_n_spl_010;
  wire G25_n_spl_011;
  wire G25_n_spl_1;
  wire G25_n_spl_10;
  wire G25_n_spl_100;
  wire G25_n_spl_101;
  wire G25_n_spl_11;
  wire G25_n_spl_110;
  wire G25_n_spl_111;
  wire G9_p_spl_;
  wire G9_p_spl_0;
  wire G9_p_spl_00;
  wire G9_p_spl_000;
  wire G9_p_spl_001;
  wire G9_p_spl_01;
  wire G9_p_spl_010;
  wire G9_p_spl_011;
  wire G9_p_spl_1;
  wire G9_p_spl_10;
  wire G9_p_spl_100;
  wire G9_p_spl_101;
  wire G9_p_spl_11;
  wire G9_p_spl_110;
  wire G9_p_spl_111;
  wire G9_n_spl_;
  wire G9_n_spl_0;
  wire G9_n_spl_00;
  wire G9_n_spl_000;
  wire G9_n_spl_001;
  wire G9_n_spl_01;
  wire G9_n_spl_010;
  wire G9_n_spl_011;
  wire G9_n_spl_1;
  wire G9_n_spl_10;
  wire G9_n_spl_100;
  wire G9_n_spl_101;
  wire G9_n_spl_11;
  wire G9_n_spl_110;
  wire G9_n_spl_111;
  wire g251_p_spl_;
  wire g252_n_spl_;
  wire g251_n_spl_;
  wire g252_p_spl_;
  wire g253_n_spl_;
  wire g253_p_spl_;
  wire g254_n_spl_;
  wire g254_n_spl_0;
  wire g254_p_spl_;
  wire g254_p_spl_0;
  wire g256_n_spl_;
  wire g256_p_spl_;
  wire g257_n_spl_;
  wire g257_p_spl_;
  wire g250_n_spl_;
  wire g259_p_spl_;
  wire g250_p_spl_;
  wire g259_n_spl_;
  wire g260_n_spl_;
  wire g260_p_spl_;
  wire g249_n_spl_;
  wire g262_p_spl_;
  wire g249_p_spl_;
  wire g262_n_spl_;
  wire g263_n_spl_;
  wire g263_p_spl_;
  wire g248_n_spl_;
  wire g265_p_spl_;
  wire g248_p_spl_;
  wire g265_n_spl_;
  wire g266_n_spl_;
  wire g266_p_spl_;
  wire g247_n_spl_;
  wire g268_p_spl_;
  wire g247_p_spl_;
  wire g268_n_spl_;
  wire g269_n_spl_;
  wire g269_p_spl_;
  wire g246_n_spl_;
  wire g271_p_spl_;
  wire g246_p_spl_;
  wire g271_n_spl_;
  wire g272_n_spl_;
  wire g272_p_spl_;
  wire g245_n_spl_;
  wire g274_p_spl_;
  wire g245_p_spl_;
  wire g274_n_spl_;
  wire g275_n_spl_;
  wire g275_p_spl_;
  wire g244_n_spl_;
  wire g277_p_spl_;
  wire g244_p_spl_;
  wire g277_n_spl_;
  wire g278_n_spl_;
  wire g278_p_spl_;
  wire g243_n_spl_;
  wire g280_p_spl_;
  wire g243_p_spl_;
  wire g280_n_spl_;
  wire g281_n_spl_;
  wire g281_p_spl_;
  wire g242_n_spl_;
  wire g283_p_spl_;
  wire g242_p_spl_;
  wire g283_n_spl_;
  wire g284_n_spl_;
  wire g284_p_spl_;
  wire g241_n_spl_;
  wire g286_p_spl_;
  wire g241_p_spl_;
  wire g286_n_spl_;
  wire g287_n_spl_;
  wire g287_p_spl_;
  wire g240_n_spl_;
  wire g289_p_spl_;
  wire g240_p_spl_;
  wire g289_n_spl_;
  wire g290_n_spl_;
  wire g290_p_spl_;
  wire g239_n_spl_;
  wire g292_p_spl_;
  wire g239_p_spl_;
  wire g292_n_spl_;
  wire g293_n_spl_;
  wire g293_p_spl_;
  wire g238_p_spl_;
  wire g295_n_spl_;
  wire g296_p_spl_;
  wire G26_p_spl_;
  wire G26_p_spl_0;
  wire G26_p_spl_00;
  wire G26_p_spl_000;
  wire G26_p_spl_001;
  wire G26_p_spl_01;
  wire G26_p_spl_010;
  wire G26_p_spl_011;
  wire G26_p_spl_1;
  wire G26_p_spl_10;
  wire G26_p_spl_100;
  wire G26_p_spl_101;
  wire G26_p_spl_11;
  wire G26_p_spl_110;
  wire G26_p_spl_111;
  wire G26_n_spl_;
  wire G26_n_spl_0;
  wire G26_n_spl_00;
  wire G26_n_spl_000;
  wire G26_n_spl_001;
  wire G26_n_spl_01;
  wire G26_n_spl_010;
  wire G26_n_spl_011;
  wire G26_n_spl_1;
  wire G26_n_spl_10;
  wire G26_n_spl_100;
  wire G26_n_spl_101;
  wire G26_n_spl_11;
  wire G26_n_spl_110;
  wire G26_n_spl_111;
  wire G10_p_spl_;
  wire G10_p_spl_0;
  wire G10_p_spl_00;
  wire G10_p_spl_000;
  wire G10_p_spl_001;
  wire G10_p_spl_01;
  wire G10_p_spl_010;
  wire G10_p_spl_011;
  wire G10_p_spl_1;
  wire G10_p_spl_10;
  wire G10_p_spl_100;
  wire G10_p_spl_101;
  wire G10_p_spl_11;
  wire G10_p_spl_110;
  wire G10_p_spl_111;
  wire G10_n_spl_;
  wire G10_n_spl_0;
  wire G10_n_spl_00;
  wire G10_n_spl_000;
  wire G10_n_spl_001;
  wire G10_n_spl_01;
  wire G10_n_spl_010;
  wire G10_n_spl_011;
  wire G10_n_spl_1;
  wire G10_n_spl_10;
  wire G10_n_spl_100;
  wire G10_n_spl_101;
  wire G10_n_spl_11;
  wire G10_n_spl_110;
  wire G10_n_spl_111;
  wire g314_p_spl_;
  wire g315_n_spl_;
  wire g314_n_spl_;
  wire g315_p_spl_;
  wire g316_n_spl_;
  wire g316_p_spl_;
  wire g317_n_spl_;
  wire g317_n_spl_0;
  wire g317_p_spl_;
  wire g317_p_spl_0;
  wire g319_n_spl_;
  wire g319_p_spl_;
  wire g320_n_spl_;
  wire g320_p_spl_;
  wire g313_n_spl_;
  wire g322_p_spl_;
  wire g313_p_spl_;
  wire g322_n_spl_;
  wire g323_n_spl_;
  wire g323_p_spl_;
  wire g312_n_spl_;
  wire g325_p_spl_;
  wire g312_p_spl_;
  wire g325_n_spl_;
  wire g326_n_spl_;
  wire g326_p_spl_;
  wire g311_n_spl_;
  wire g328_p_spl_;
  wire g311_p_spl_;
  wire g328_n_spl_;
  wire g329_n_spl_;
  wire g329_p_spl_;
  wire g310_n_spl_;
  wire g331_p_spl_;
  wire g310_p_spl_;
  wire g331_n_spl_;
  wire g332_n_spl_;
  wire g332_p_spl_;
  wire g309_n_spl_;
  wire g334_p_spl_;
  wire g309_p_spl_;
  wire g334_n_spl_;
  wire g335_n_spl_;
  wire g335_p_spl_;
  wire g308_n_spl_;
  wire g337_p_spl_;
  wire g308_p_spl_;
  wire g337_n_spl_;
  wire g338_n_spl_;
  wire g338_p_spl_;
  wire g307_n_spl_;
  wire g340_p_spl_;
  wire g307_p_spl_;
  wire g340_n_spl_;
  wire g341_n_spl_;
  wire g341_p_spl_;
  wire g306_n_spl_;
  wire g343_p_spl_;
  wire g306_p_spl_;
  wire g343_n_spl_;
  wire g344_n_spl_;
  wire g344_p_spl_;
  wire g305_n_spl_;
  wire g346_p_spl_;
  wire g305_p_spl_;
  wire g346_n_spl_;
  wire g347_n_spl_;
  wire g347_p_spl_;
  wire g304_n_spl_;
  wire g349_p_spl_;
  wire g304_p_spl_;
  wire g349_n_spl_;
  wire g350_n_spl_;
  wire g350_p_spl_;
  wire g303_n_spl_;
  wire g352_p_spl_;
  wire g303_p_spl_;
  wire g352_n_spl_;
  wire g353_n_spl_;
  wire g353_p_spl_;
  wire g302_n_spl_;
  wire g355_p_spl_;
  wire g302_p_spl_;
  wire g355_n_spl_;
  wire g356_n_spl_;
  wire g356_p_spl_;
  wire g301_n_spl_;
  wire g358_p_spl_;
  wire g301_p_spl_;
  wire g358_n_spl_;
  wire g359_n_spl_;
  wire g359_p_spl_;
  wire g300_n_spl_;
  wire g361_p_spl_;
  wire g300_p_spl_;
  wire g361_n_spl_;
  wire g362_n_spl_;
  wire g362_p_spl_;
  wire g299_p_spl_;
  wire g364_n_spl_;
  wire g365_p_spl_;
  wire G27_p_spl_;
  wire G27_p_spl_0;
  wire G27_p_spl_00;
  wire G27_p_spl_000;
  wire G27_p_spl_001;
  wire G27_p_spl_01;
  wire G27_p_spl_010;
  wire G27_p_spl_011;
  wire G27_p_spl_1;
  wire G27_p_spl_10;
  wire G27_p_spl_100;
  wire G27_p_spl_101;
  wire G27_p_spl_11;
  wire G27_p_spl_110;
  wire G27_p_spl_111;
  wire G27_n_spl_;
  wire G27_n_spl_0;
  wire G27_n_spl_00;
  wire G27_n_spl_000;
  wire G27_n_spl_001;
  wire G27_n_spl_01;
  wire G27_n_spl_010;
  wire G27_n_spl_011;
  wire G27_n_spl_1;
  wire G27_n_spl_10;
  wire G27_n_spl_100;
  wire G27_n_spl_101;
  wire G27_n_spl_11;
  wire G27_n_spl_110;
  wire G27_n_spl_111;
  wire G11_p_spl_;
  wire G11_p_spl_0;
  wire G11_p_spl_00;
  wire G11_p_spl_000;
  wire G11_p_spl_001;
  wire G11_p_spl_01;
  wire G11_p_spl_010;
  wire G11_p_spl_011;
  wire G11_p_spl_1;
  wire G11_p_spl_10;
  wire G11_p_spl_100;
  wire G11_p_spl_101;
  wire G11_p_spl_11;
  wire G11_p_spl_110;
  wire G11_p_spl_111;
  wire G11_n_spl_;
  wire G11_n_spl_0;
  wire G11_n_spl_00;
  wire G11_n_spl_000;
  wire G11_n_spl_001;
  wire G11_n_spl_01;
  wire G11_n_spl_010;
  wire G11_n_spl_011;
  wire G11_n_spl_1;
  wire G11_n_spl_10;
  wire G11_n_spl_100;
  wire G11_n_spl_101;
  wire G11_n_spl_11;
  wire G11_n_spl_110;
  wire G11_n_spl_111;
  wire g385_p_spl_;
  wire g386_n_spl_;
  wire g385_n_spl_;
  wire g386_p_spl_;
  wire g387_n_spl_;
  wire g387_p_spl_;
  wire g388_n_spl_;
  wire g388_n_spl_0;
  wire g388_p_spl_;
  wire g388_p_spl_0;
  wire g390_n_spl_;
  wire g390_p_spl_;
  wire g391_n_spl_;
  wire g391_p_spl_;
  wire g384_n_spl_;
  wire g393_p_spl_;
  wire g384_p_spl_;
  wire g393_n_spl_;
  wire g394_n_spl_;
  wire g394_p_spl_;
  wire g383_n_spl_;
  wire g396_p_spl_;
  wire g383_p_spl_;
  wire g396_n_spl_;
  wire g397_n_spl_;
  wire g397_p_spl_;
  wire g382_n_spl_;
  wire g399_p_spl_;
  wire g382_p_spl_;
  wire g399_n_spl_;
  wire g400_n_spl_;
  wire g400_p_spl_;
  wire g381_n_spl_;
  wire g402_p_spl_;
  wire g381_p_spl_;
  wire g402_n_spl_;
  wire g403_n_spl_;
  wire g403_p_spl_;
  wire g380_n_spl_;
  wire g405_p_spl_;
  wire g380_p_spl_;
  wire g405_n_spl_;
  wire g406_n_spl_;
  wire g406_p_spl_;
  wire g379_n_spl_;
  wire g408_p_spl_;
  wire g379_p_spl_;
  wire g408_n_spl_;
  wire g409_n_spl_;
  wire g409_p_spl_;
  wire g378_n_spl_;
  wire g411_p_spl_;
  wire g378_p_spl_;
  wire g411_n_spl_;
  wire g412_n_spl_;
  wire g412_p_spl_;
  wire g377_n_spl_;
  wire g414_p_spl_;
  wire g377_p_spl_;
  wire g414_n_spl_;
  wire g415_n_spl_;
  wire g415_p_spl_;
  wire g376_n_spl_;
  wire g417_p_spl_;
  wire g376_p_spl_;
  wire g417_n_spl_;
  wire g418_n_spl_;
  wire g418_p_spl_;
  wire g375_n_spl_;
  wire g420_p_spl_;
  wire g375_p_spl_;
  wire g420_n_spl_;
  wire g421_n_spl_;
  wire g421_p_spl_;
  wire g374_n_spl_;
  wire g423_p_spl_;
  wire g374_p_spl_;
  wire g423_n_spl_;
  wire g424_n_spl_;
  wire g424_p_spl_;
  wire g373_n_spl_;
  wire g426_p_spl_;
  wire g373_p_spl_;
  wire g426_n_spl_;
  wire g427_n_spl_;
  wire g427_p_spl_;
  wire g372_n_spl_;
  wire g429_p_spl_;
  wire g372_p_spl_;
  wire g429_n_spl_;
  wire g430_n_spl_;
  wire g430_p_spl_;
  wire g371_n_spl_;
  wire g432_p_spl_;
  wire g371_p_spl_;
  wire g432_n_spl_;
  wire g433_n_spl_;
  wire g433_p_spl_;
  wire g370_n_spl_;
  wire g435_p_spl_;
  wire g370_p_spl_;
  wire g435_n_spl_;
  wire g436_n_spl_;
  wire g436_p_spl_;
  wire g369_n_spl_;
  wire g438_p_spl_;
  wire g369_p_spl_;
  wire g438_n_spl_;
  wire g439_n_spl_;
  wire g439_p_spl_;
  wire g368_p_spl_;
  wire g441_n_spl_;
  wire g442_p_spl_;
  wire G28_p_spl_;
  wire G28_p_spl_0;
  wire G28_p_spl_00;
  wire G28_p_spl_000;
  wire G28_p_spl_001;
  wire G28_p_spl_01;
  wire G28_p_spl_010;
  wire G28_p_spl_011;
  wire G28_p_spl_1;
  wire G28_p_spl_10;
  wire G28_p_spl_100;
  wire G28_p_spl_101;
  wire G28_p_spl_11;
  wire G28_p_spl_110;
  wire G28_p_spl_111;
  wire G28_n_spl_;
  wire G28_n_spl_0;
  wire G28_n_spl_00;
  wire G28_n_spl_000;
  wire G28_n_spl_001;
  wire G28_n_spl_01;
  wire G28_n_spl_010;
  wire G28_n_spl_011;
  wire G28_n_spl_1;
  wire G28_n_spl_10;
  wire G28_n_spl_100;
  wire G28_n_spl_101;
  wire G28_n_spl_11;
  wire G28_n_spl_110;
  wire G28_n_spl_111;
  wire G12_p_spl_;
  wire G12_p_spl_0;
  wire G12_p_spl_00;
  wire G12_p_spl_000;
  wire G12_p_spl_001;
  wire G12_p_spl_01;
  wire G12_p_spl_010;
  wire G12_p_spl_011;
  wire G12_p_spl_1;
  wire G12_p_spl_10;
  wire G12_p_spl_100;
  wire G12_p_spl_101;
  wire G12_p_spl_11;
  wire G12_p_spl_110;
  wire G12_p_spl_111;
  wire G12_n_spl_;
  wire G12_n_spl_0;
  wire G12_n_spl_00;
  wire G12_n_spl_000;
  wire G12_n_spl_001;
  wire G12_n_spl_01;
  wire G12_n_spl_010;
  wire G12_n_spl_011;
  wire G12_n_spl_1;
  wire G12_n_spl_10;
  wire G12_n_spl_100;
  wire G12_n_spl_101;
  wire G12_n_spl_11;
  wire G12_n_spl_110;
  wire G12_n_spl_111;
  wire g464_p_spl_;
  wire g465_n_spl_;
  wire g464_n_spl_;
  wire g465_p_spl_;
  wire g466_n_spl_;
  wire g466_p_spl_;
  wire g467_n_spl_;
  wire g467_n_spl_0;
  wire g467_p_spl_;
  wire g467_p_spl_0;
  wire g469_n_spl_;
  wire g469_p_spl_;
  wire g470_n_spl_;
  wire g470_p_spl_;
  wire g463_n_spl_;
  wire g472_p_spl_;
  wire g463_p_spl_;
  wire g472_n_spl_;
  wire g473_n_spl_;
  wire g473_p_spl_;
  wire g462_n_spl_;
  wire g475_p_spl_;
  wire g462_p_spl_;
  wire g475_n_spl_;
  wire g476_n_spl_;
  wire g476_p_spl_;
  wire g461_n_spl_;
  wire g478_p_spl_;
  wire g461_p_spl_;
  wire g478_n_spl_;
  wire g479_n_spl_;
  wire g479_p_spl_;
  wire g460_n_spl_;
  wire g481_p_spl_;
  wire g460_p_spl_;
  wire g481_n_spl_;
  wire g482_n_spl_;
  wire g482_p_spl_;
  wire g459_n_spl_;
  wire g484_p_spl_;
  wire g459_p_spl_;
  wire g484_n_spl_;
  wire g485_n_spl_;
  wire g485_p_spl_;
  wire g458_n_spl_;
  wire g487_p_spl_;
  wire g458_p_spl_;
  wire g487_n_spl_;
  wire g488_n_spl_;
  wire g488_p_spl_;
  wire g457_n_spl_;
  wire g490_p_spl_;
  wire g457_p_spl_;
  wire g490_n_spl_;
  wire g491_n_spl_;
  wire g491_p_spl_;
  wire g456_n_spl_;
  wire g493_p_spl_;
  wire g456_p_spl_;
  wire g493_n_spl_;
  wire g494_n_spl_;
  wire g494_p_spl_;
  wire g455_n_spl_;
  wire g496_p_spl_;
  wire g455_p_spl_;
  wire g496_n_spl_;
  wire g497_n_spl_;
  wire g497_p_spl_;
  wire g454_n_spl_;
  wire g499_p_spl_;
  wire g454_p_spl_;
  wire g499_n_spl_;
  wire g500_n_spl_;
  wire g500_p_spl_;
  wire g453_n_spl_;
  wire g502_p_spl_;
  wire g453_p_spl_;
  wire g502_n_spl_;
  wire g503_n_spl_;
  wire g503_p_spl_;
  wire g452_n_spl_;
  wire g505_p_spl_;
  wire g452_p_spl_;
  wire g505_n_spl_;
  wire g506_n_spl_;
  wire g506_p_spl_;
  wire g451_n_spl_;
  wire g508_p_spl_;
  wire g451_p_spl_;
  wire g508_n_spl_;
  wire g509_n_spl_;
  wire g509_p_spl_;
  wire g450_n_spl_;
  wire g511_p_spl_;
  wire g450_p_spl_;
  wire g511_n_spl_;
  wire g512_n_spl_;
  wire g512_p_spl_;
  wire g449_n_spl_;
  wire g514_p_spl_;
  wire g449_p_spl_;
  wire g514_n_spl_;
  wire g515_n_spl_;
  wire g515_p_spl_;
  wire g448_n_spl_;
  wire g517_p_spl_;
  wire g448_p_spl_;
  wire g517_n_spl_;
  wire g518_n_spl_;
  wire g518_p_spl_;
  wire g447_n_spl_;
  wire g520_p_spl_;
  wire g447_p_spl_;
  wire g520_n_spl_;
  wire g521_n_spl_;
  wire g521_p_spl_;
  wire g446_n_spl_;
  wire g523_p_spl_;
  wire g446_p_spl_;
  wire g523_n_spl_;
  wire g524_n_spl_;
  wire g524_p_spl_;
  wire g445_p_spl_;
  wire g526_n_spl_;
  wire g527_p_spl_;
  wire G29_p_spl_;
  wire G29_p_spl_0;
  wire G29_p_spl_00;
  wire G29_p_spl_000;
  wire G29_p_spl_001;
  wire G29_p_spl_01;
  wire G29_p_spl_010;
  wire G29_p_spl_011;
  wire G29_p_spl_1;
  wire G29_p_spl_10;
  wire G29_p_spl_100;
  wire G29_p_spl_101;
  wire G29_p_spl_11;
  wire G29_p_spl_110;
  wire G29_p_spl_111;
  wire G29_n_spl_;
  wire G29_n_spl_0;
  wire G29_n_spl_00;
  wire G29_n_spl_000;
  wire G29_n_spl_001;
  wire G29_n_spl_01;
  wire G29_n_spl_010;
  wire G29_n_spl_011;
  wire G29_n_spl_1;
  wire G29_n_spl_10;
  wire G29_n_spl_100;
  wire G29_n_spl_101;
  wire G29_n_spl_11;
  wire G29_n_spl_110;
  wire G29_n_spl_111;
  wire G13_p_spl_;
  wire G13_p_spl_0;
  wire G13_p_spl_00;
  wire G13_p_spl_000;
  wire G13_p_spl_001;
  wire G13_p_spl_01;
  wire G13_p_spl_010;
  wire G13_p_spl_011;
  wire G13_p_spl_1;
  wire G13_p_spl_10;
  wire G13_p_spl_100;
  wire G13_p_spl_101;
  wire G13_p_spl_11;
  wire G13_p_spl_110;
  wire G13_p_spl_111;
  wire G13_n_spl_;
  wire G13_n_spl_0;
  wire G13_n_spl_00;
  wire G13_n_spl_000;
  wire G13_n_spl_001;
  wire G13_n_spl_01;
  wire G13_n_spl_010;
  wire G13_n_spl_011;
  wire G13_n_spl_1;
  wire G13_n_spl_10;
  wire G13_n_spl_100;
  wire G13_n_spl_101;
  wire G13_n_spl_11;
  wire G13_n_spl_110;
  wire G13_n_spl_111;
  wire g551_p_spl_;
  wire g552_n_spl_;
  wire g551_n_spl_;
  wire g552_p_spl_;
  wire g553_n_spl_;
  wire g553_p_spl_;
  wire g554_n_spl_;
  wire g554_n_spl_0;
  wire g554_p_spl_;
  wire g554_p_spl_0;
  wire g556_n_spl_;
  wire g556_p_spl_;
  wire g557_n_spl_;
  wire g557_p_spl_;
  wire g550_n_spl_;
  wire g559_p_spl_;
  wire g550_p_spl_;
  wire g559_n_spl_;
  wire g560_n_spl_;
  wire g560_p_spl_;
  wire g549_n_spl_;
  wire g562_p_spl_;
  wire g549_p_spl_;
  wire g562_n_spl_;
  wire g563_n_spl_;
  wire g563_p_spl_;
  wire g548_n_spl_;
  wire g565_p_spl_;
  wire g548_p_spl_;
  wire g565_n_spl_;
  wire g566_n_spl_;
  wire g566_p_spl_;
  wire g547_n_spl_;
  wire g568_p_spl_;
  wire g547_p_spl_;
  wire g568_n_spl_;
  wire g569_n_spl_;
  wire g569_p_spl_;
  wire g546_n_spl_;
  wire g571_p_spl_;
  wire g546_p_spl_;
  wire g571_n_spl_;
  wire g572_n_spl_;
  wire g572_p_spl_;
  wire g545_n_spl_;
  wire g574_p_spl_;
  wire g545_p_spl_;
  wire g574_n_spl_;
  wire g575_n_spl_;
  wire g575_p_spl_;
  wire g544_n_spl_;
  wire g577_p_spl_;
  wire g544_p_spl_;
  wire g577_n_spl_;
  wire g578_n_spl_;
  wire g578_p_spl_;
  wire g543_n_spl_;
  wire g580_p_spl_;
  wire g543_p_spl_;
  wire g580_n_spl_;
  wire g581_n_spl_;
  wire g581_p_spl_;
  wire g542_n_spl_;
  wire g583_p_spl_;
  wire g542_p_spl_;
  wire g583_n_spl_;
  wire g584_n_spl_;
  wire g584_p_spl_;
  wire g541_n_spl_;
  wire g586_p_spl_;
  wire g541_p_spl_;
  wire g586_n_spl_;
  wire g587_n_spl_;
  wire g587_p_spl_;
  wire g540_n_spl_;
  wire g589_p_spl_;
  wire g540_p_spl_;
  wire g589_n_spl_;
  wire g590_n_spl_;
  wire g590_p_spl_;
  wire g539_n_spl_;
  wire g592_p_spl_;
  wire g539_p_spl_;
  wire g592_n_spl_;
  wire g593_n_spl_;
  wire g593_p_spl_;
  wire g538_n_spl_;
  wire g595_p_spl_;
  wire g538_p_spl_;
  wire g595_n_spl_;
  wire g596_n_spl_;
  wire g596_p_spl_;
  wire g537_n_spl_;
  wire g598_p_spl_;
  wire g537_p_spl_;
  wire g598_n_spl_;
  wire g599_n_spl_;
  wire g599_p_spl_;
  wire g536_n_spl_;
  wire g601_p_spl_;
  wire g536_p_spl_;
  wire g601_n_spl_;
  wire g602_n_spl_;
  wire g602_p_spl_;
  wire g535_n_spl_;
  wire g604_p_spl_;
  wire g535_p_spl_;
  wire g604_n_spl_;
  wire g605_n_spl_;
  wire g605_p_spl_;
  wire g534_n_spl_;
  wire g607_p_spl_;
  wire g534_p_spl_;
  wire g607_n_spl_;
  wire g608_n_spl_;
  wire g608_p_spl_;
  wire g533_n_spl_;
  wire g610_p_spl_;
  wire g533_p_spl_;
  wire g610_n_spl_;
  wire g611_n_spl_;
  wire g611_p_spl_;
  wire g532_n_spl_;
  wire g613_p_spl_;
  wire g532_p_spl_;
  wire g613_n_spl_;
  wire g614_n_spl_;
  wire g614_p_spl_;
  wire g531_n_spl_;
  wire g616_p_spl_;
  wire g531_p_spl_;
  wire g616_n_spl_;
  wire g617_n_spl_;
  wire g617_p_spl_;
  wire g530_p_spl_;
  wire g619_n_spl_;
  wire g620_p_spl_;
  wire G30_p_spl_;
  wire G30_p_spl_0;
  wire G30_p_spl_00;
  wire G30_p_spl_000;
  wire G30_p_spl_001;
  wire G30_p_spl_01;
  wire G30_p_spl_010;
  wire G30_p_spl_011;
  wire G30_p_spl_1;
  wire G30_p_spl_10;
  wire G30_p_spl_100;
  wire G30_p_spl_101;
  wire G30_p_spl_11;
  wire G30_p_spl_110;
  wire G30_p_spl_111;
  wire G30_n_spl_;
  wire G30_n_spl_0;
  wire G30_n_spl_00;
  wire G30_n_spl_000;
  wire G30_n_spl_001;
  wire G30_n_spl_01;
  wire G30_n_spl_010;
  wire G30_n_spl_011;
  wire G30_n_spl_1;
  wire G30_n_spl_10;
  wire G30_n_spl_100;
  wire G30_n_spl_101;
  wire G30_n_spl_11;
  wire G30_n_spl_110;
  wire G30_n_spl_111;
  wire G14_p_spl_;
  wire G14_p_spl_0;
  wire G14_p_spl_00;
  wire G14_p_spl_000;
  wire G14_p_spl_001;
  wire G14_p_spl_01;
  wire G14_p_spl_010;
  wire G14_p_spl_011;
  wire G14_p_spl_1;
  wire G14_p_spl_10;
  wire G14_p_spl_100;
  wire G14_p_spl_101;
  wire G14_p_spl_11;
  wire G14_p_spl_110;
  wire G14_p_spl_111;
  wire G14_n_spl_;
  wire G14_n_spl_0;
  wire G14_n_spl_00;
  wire G14_n_spl_000;
  wire G14_n_spl_001;
  wire G14_n_spl_01;
  wire G14_n_spl_010;
  wire G14_n_spl_011;
  wire G14_n_spl_1;
  wire G14_n_spl_10;
  wire G14_n_spl_100;
  wire G14_n_spl_101;
  wire G14_n_spl_11;
  wire G14_n_spl_110;
  wire G14_n_spl_111;
  wire g646_p_spl_;
  wire g647_n_spl_;
  wire g646_n_spl_;
  wire g647_p_spl_;
  wire g648_n_spl_;
  wire g648_p_spl_;
  wire g649_n_spl_;
  wire g649_n_spl_0;
  wire g649_p_spl_;
  wire g649_p_spl_0;
  wire g651_n_spl_;
  wire g651_p_spl_;
  wire g652_n_spl_;
  wire g652_p_spl_;
  wire g645_n_spl_;
  wire g654_p_spl_;
  wire g645_p_spl_;
  wire g654_n_spl_;
  wire g655_n_spl_;
  wire g655_p_spl_;
  wire g644_n_spl_;
  wire g657_p_spl_;
  wire g644_p_spl_;
  wire g657_n_spl_;
  wire g658_n_spl_;
  wire g658_p_spl_;
  wire g643_n_spl_;
  wire g660_p_spl_;
  wire g643_p_spl_;
  wire g660_n_spl_;
  wire g661_n_spl_;
  wire g661_p_spl_;
  wire g642_n_spl_;
  wire g663_p_spl_;
  wire g642_p_spl_;
  wire g663_n_spl_;
  wire g664_n_spl_;
  wire g664_p_spl_;
  wire g641_n_spl_;
  wire g666_p_spl_;
  wire g641_p_spl_;
  wire g666_n_spl_;
  wire g667_n_spl_;
  wire g667_p_spl_;
  wire g640_n_spl_;
  wire g669_p_spl_;
  wire g640_p_spl_;
  wire g669_n_spl_;
  wire g670_n_spl_;
  wire g670_p_spl_;
  wire g639_n_spl_;
  wire g672_p_spl_;
  wire g639_p_spl_;
  wire g672_n_spl_;
  wire g673_n_spl_;
  wire g673_p_spl_;
  wire g638_n_spl_;
  wire g675_p_spl_;
  wire g638_p_spl_;
  wire g675_n_spl_;
  wire g676_n_spl_;
  wire g676_p_spl_;
  wire g637_n_spl_;
  wire g678_p_spl_;
  wire g637_p_spl_;
  wire g678_n_spl_;
  wire g679_n_spl_;
  wire g679_p_spl_;
  wire g636_n_spl_;
  wire g681_p_spl_;
  wire g636_p_spl_;
  wire g681_n_spl_;
  wire g682_n_spl_;
  wire g682_p_spl_;
  wire g635_n_spl_;
  wire g684_p_spl_;
  wire g635_p_spl_;
  wire g684_n_spl_;
  wire g685_n_spl_;
  wire g685_p_spl_;
  wire g634_n_spl_;
  wire g687_p_spl_;
  wire g634_p_spl_;
  wire g687_n_spl_;
  wire g688_n_spl_;
  wire g688_p_spl_;
  wire g633_n_spl_;
  wire g690_p_spl_;
  wire g633_p_spl_;
  wire g690_n_spl_;
  wire g691_n_spl_;
  wire g691_p_spl_;
  wire g632_n_spl_;
  wire g693_p_spl_;
  wire g632_p_spl_;
  wire g693_n_spl_;
  wire g694_n_spl_;
  wire g694_p_spl_;
  wire g631_n_spl_;
  wire g696_p_spl_;
  wire g631_p_spl_;
  wire g696_n_spl_;
  wire g697_n_spl_;
  wire g697_p_spl_;
  wire g630_n_spl_;
  wire g699_p_spl_;
  wire g630_p_spl_;
  wire g699_n_spl_;
  wire g700_n_spl_;
  wire g700_p_spl_;
  wire g629_n_spl_;
  wire g702_p_spl_;
  wire g629_p_spl_;
  wire g702_n_spl_;
  wire g703_n_spl_;
  wire g703_p_spl_;
  wire g628_n_spl_;
  wire g705_p_spl_;
  wire g628_p_spl_;
  wire g705_n_spl_;
  wire g706_n_spl_;
  wire g706_p_spl_;
  wire g627_n_spl_;
  wire g708_p_spl_;
  wire g627_p_spl_;
  wire g708_n_spl_;
  wire g709_n_spl_;
  wire g709_p_spl_;
  wire g626_n_spl_;
  wire g711_p_spl_;
  wire g626_p_spl_;
  wire g711_n_spl_;
  wire g712_n_spl_;
  wire g712_p_spl_;
  wire g625_n_spl_;
  wire g714_p_spl_;
  wire g625_p_spl_;
  wire g714_n_spl_;
  wire g715_n_spl_;
  wire g715_p_spl_;
  wire g624_n_spl_;
  wire g717_p_spl_;
  wire g624_p_spl_;
  wire g717_n_spl_;
  wire g718_n_spl_;
  wire g718_p_spl_;
  wire g623_p_spl_;
  wire g720_n_spl_;
  wire g721_p_spl_;
  wire G31_p_spl_;
  wire G31_p_spl_0;
  wire G31_p_spl_00;
  wire G31_p_spl_000;
  wire G31_p_spl_001;
  wire G31_p_spl_01;
  wire G31_p_spl_010;
  wire G31_p_spl_011;
  wire G31_p_spl_1;
  wire G31_p_spl_10;
  wire G31_p_spl_100;
  wire G31_p_spl_101;
  wire G31_p_spl_11;
  wire G31_p_spl_110;
  wire G31_p_spl_111;
  wire G31_n_spl_;
  wire G31_n_spl_0;
  wire G31_n_spl_00;
  wire G31_n_spl_000;
  wire G31_n_spl_001;
  wire G31_n_spl_01;
  wire G31_n_spl_010;
  wire G31_n_spl_011;
  wire G31_n_spl_1;
  wire G31_n_spl_10;
  wire G31_n_spl_100;
  wire G31_n_spl_101;
  wire G31_n_spl_11;
  wire G31_n_spl_110;
  wire G31_n_spl_111;
  wire G15_p_spl_;
  wire G15_p_spl_0;
  wire G15_p_spl_00;
  wire G15_p_spl_000;
  wire G15_p_spl_001;
  wire G15_p_spl_01;
  wire G15_p_spl_010;
  wire G15_p_spl_011;
  wire G15_p_spl_1;
  wire G15_p_spl_10;
  wire G15_p_spl_100;
  wire G15_p_spl_101;
  wire G15_p_spl_11;
  wire G15_p_spl_110;
  wire G15_p_spl_111;
  wire G15_n_spl_;
  wire G15_n_spl_0;
  wire G15_n_spl_00;
  wire G15_n_spl_000;
  wire G15_n_spl_001;
  wire G15_n_spl_01;
  wire G15_n_spl_010;
  wire G15_n_spl_011;
  wire G15_n_spl_1;
  wire G15_n_spl_10;
  wire G15_n_spl_100;
  wire G15_n_spl_101;
  wire G15_n_spl_11;
  wire G15_n_spl_110;
  wire G15_n_spl_111;
  wire g749_p_spl_;
  wire g750_n_spl_;
  wire g749_n_spl_;
  wire g750_p_spl_;
  wire g751_n_spl_;
  wire g751_p_spl_;
  wire g752_n_spl_;
  wire g752_n_spl_0;
  wire g752_p_spl_;
  wire g752_p_spl_0;
  wire g754_n_spl_;
  wire g754_p_spl_;
  wire g755_n_spl_;
  wire g755_p_spl_;
  wire g748_n_spl_;
  wire g757_p_spl_;
  wire g748_p_spl_;
  wire g757_n_spl_;
  wire g758_n_spl_;
  wire g758_p_spl_;
  wire g747_n_spl_;
  wire g760_p_spl_;
  wire g747_p_spl_;
  wire g760_n_spl_;
  wire g761_n_spl_;
  wire g761_p_spl_;
  wire g746_n_spl_;
  wire g763_p_spl_;
  wire g746_p_spl_;
  wire g763_n_spl_;
  wire g764_n_spl_;
  wire g764_p_spl_;
  wire g745_n_spl_;
  wire g766_p_spl_;
  wire g745_p_spl_;
  wire g766_n_spl_;
  wire g767_n_spl_;
  wire g767_p_spl_;
  wire g744_n_spl_;
  wire g769_p_spl_;
  wire g744_p_spl_;
  wire g769_n_spl_;
  wire g770_n_spl_;
  wire g770_p_spl_;
  wire g743_n_spl_;
  wire g772_p_spl_;
  wire g743_p_spl_;
  wire g772_n_spl_;
  wire g773_n_spl_;
  wire g773_p_spl_;
  wire g742_n_spl_;
  wire g775_p_spl_;
  wire g742_p_spl_;
  wire g775_n_spl_;
  wire g776_n_spl_;
  wire g776_p_spl_;
  wire g741_n_spl_;
  wire g778_p_spl_;
  wire g741_p_spl_;
  wire g778_n_spl_;
  wire g779_n_spl_;
  wire g779_p_spl_;
  wire g740_n_spl_;
  wire g781_p_spl_;
  wire g740_p_spl_;
  wire g781_n_spl_;
  wire g782_n_spl_;
  wire g782_p_spl_;
  wire g739_n_spl_;
  wire g784_p_spl_;
  wire g739_p_spl_;
  wire g784_n_spl_;
  wire g785_n_spl_;
  wire g785_p_spl_;
  wire g738_n_spl_;
  wire g787_p_spl_;
  wire g738_p_spl_;
  wire g787_n_spl_;
  wire g788_n_spl_;
  wire g788_p_spl_;
  wire g737_n_spl_;
  wire g790_p_spl_;
  wire g737_p_spl_;
  wire g790_n_spl_;
  wire g791_n_spl_;
  wire g791_p_spl_;
  wire g736_n_spl_;
  wire g793_p_spl_;
  wire g736_p_spl_;
  wire g793_n_spl_;
  wire g794_n_spl_;
  wire g794_p_spl_;
  wire g735_n_spl_;
  wire g796_p_spl_;
  wire g735_p_spl_;
  wire g796_n_spl_;
  wire g797_n_spl_;
  wire g797_p_spl_;
  wire g734_n_spl_;
  wire g799_p_spl_;
  wire g734_p_spl_;
  wire g799_n_spl_;
  wire g800_n_spl_;
  wire g800_p_spl_;
  wire g733_n_spl_;
  wire g802_p_spl_;
  wire g733_p_spl_;
  wire g802_n_spl_;
  wire g803_n_spl_;
  wire g803_p_spl_;
  wire g732_n_spl_;
  wire g805_p_spl_;
  wire g732_p_spl_;
  wire g805_n_spl_;
  wire g806_n_spl_;
  wire g806_p_spl_;
  wire g731_n_spl_;
  wire g808_p_spl_;
  wire g731_p_spl_;
  wire g808_n_spl_;
  wire g809_n_spl_;
  wire g809_p_spl_;
  wire g730_n_spl_;
  wire g811_p_spl_;
  wire g730_p_spl_;
  wire g811_n_spl_;
  wire g812_n_spl_;
  wire g812_p_spl_;
  wire g729_n_spl_;
  wire g814_p_spl_;
  wire g729_p_spl_;
  wire g814_n_spl_;
  wire g815_n_spl_;
  wire g815_p_spl_;
  wire g728_n_spl_;
  wire g817_p_spl_;
  wire g728_p_spl_;
  wire g817_n_spl_;
  wire g818_n_spl_;
  wire g818_p_spl_;
  wire g727_n_spl_;
  wire g820_p_spl_;
  wire g727_p_spl_;
  wire g820_n_spl_;
  wire g821_n_spl_;
  wire g821_p_spl_;
  wire g726_n_spl_;
  wire g823_p_spl_;
  wire g726_p_spl_;
  wire g823_n_spl_;
  wire g824_n_spl_;
  wire g824_p_spl_;
  wire g725_n_spl_;
  wire g826_p_spl_;
  wire g725_p_spl_;
  wire g826_n_spl_;
  wire g827_n_spl_;
  wire g827_p_spl_;
  wire g724_p_spl_;
  wire g829_n_spl_;
  wire g830_p_spl_;
  wire G32_p_spl_;
  wire G32_p_spl_0;
  wire G32_p_spl_00;
  wire G32_p_spl_000;
  wire G32_p_spl_001;
  wire G32_p_spl_01;
  wire G32_p_spl_010;
  wire G32_p_spl_011;
  wire G32_p_spl_1;
  wire G32_p_spl_10;
  wire G32_p_spl_100;
  wire G32_p_spl_101;
  wire G32_p_spl_11;
  wire G32_p_spl_110;
  wire G32_p_spl_111;
  wire G32_n_spl_;
  wire G32_n_spl_0;
  wire G32_n_spl_00;
  wire G32_n_spl_000;
  wire G32_n_spl_001;
  wire G32_n_spl_01;
  wire G32_n_spl_010;
  wire G32_n_spl_011;
  wire G32_n_spl_1;
  wire G32_n_spl_10;
  wire G32_n_spl_100;
  wire G32_n_spl_101;
  wire G32_n_spl_11;
  wire G32_n_spl_110;
  wire G32_n_spl_111;
  wire G16_p_spl_;
  wire G16_p_spl_0;
  wire G16_p_spl_00;
  wire G16_p_spl_000;
  wire G16_p_spl_001;
  wire G16_p_spl_01;
  wire G16_p_spl_010;
  wire G16_p_spl_011;
  wire G16_p_spl_1;
  wire G16_p_spl_10;
  wire G16_p_spl_100;
  wire G16_p_spl_101;
  wire G16_p_spl_11;
  wire G16_p_spl_110;
  wire G16_p_spl_111;
  wire G16_n_spl_;
  wire G16_n_spl_0;
  wire G16_n_spl_00;
  wire G16_n_spl_000;
  wire G16_n_spl_001;
  wire G16_n_spl_01;
  wire G16_n_spl_010;
  wire G16_n_spl_011;
  wire G16_n_spl_1;
  wire G16_n_spl_10;
  wire G16_n_spl_100;
  wire G16_n_spl_101;
  wire G16_n_spl_11;
  wire G16_n_spl_110;
  wire G16_n_spl_111;
  wire g860_p_spl_;
  wire g861_n_spl_;
  wire g860_n_spl_;
  wire g861_p_spl_;
  wire g862_n_spl_;
  wire g862_p_spl_;
  wire g863_n_spl_;
  wire g863_p_spl_;
  wire g865_n_spl_;
  wire g865_p_spl_;
  wire g866_n_spl_;
  wire g866_p_spl_;
  wire g859_n_spl_;
  wire g868_p_spl_;
  wire g859_p_spl_;
  wire g868_n_spl_;
  wire g869_n_spl_;
  wire g869_p_spl_;
  wire g858_n_spl_;
  wire g871_p_spl_;
  wire g858_p_spl_;
  wire g871_n_spl_;
  wire g872_n_spl_;
  wire g872_p_spl_;
  wire g857_n_spl_;
  wire g874_p_spl_;
  wire g857_p_spl_;
  wire g874_n_spl_;
  wire g875_n_spl_;
  wire g875_p_spl_;
  wire g856_n_spl_;
  wire g877_p_spl_;
  wire g856_p_spl_;
  wire g877_n_spl_;
  wire g878_n_spl_;
  wire g878_p_spl_;
  wire g855_n_spl_;
  wire g880_p_spl_;
  wire g855_p_spl_;
  wire g880_n_spl_;
  wire g881_n_spl_;
  wire g881_p_spl_;
  wire g854_n_spl_;
  wire g883_p_spl_;
  wire g854_p_spl_;
  wire g883_n_spl_;
  wire g884_n_spl_;
  wire g884_p_spl_;
  wire g853_n_spl_;
  wire g886_p_spl_;
  wire g853_p_spl_;
  wire g886_n_spl_;
  wire g887_n_spl_;
  wire g887_p_spl_;
  wire g852_n_spl_;
  wire g889_p_spl_;
  wire g852_p_spl_;
  wire g889_n_spl_;
  wire g890_n_spl_;
  wire g890_p_spl_;
  wire g851_n_spl_;
  wire g892_p_spl_;
  wire g851_p_spl_;
  wire g892_n_spl_;
  wire g893_n_spl_;
  wire g893_p_spl_;
  wire g850_n_spl_;
  wire g895_p_spl_;
  wire g850_p_spl_;
  wire g895_n_spl_;
  wire g896_n_spl_;
  wire g896_p_spl_;
  wire g849_n_spl_;
  wire g898_p_spl_;
  wire g849_p_spl_;
  wire g898_n_spl_;
  wire g899_n_spl_;
  wire g899_p_spl_;
  wire g848_n_spl_;
  wire g901_p_spl_;
  wire g848_p_spl_;
  wire g901_n_spl_;
  wire g902_n_spl_;
  wire g902_p_spl_;
  wire g847_n_spl_;
  wire g904_p_spl_;
  wire g847_p_spl_;
  wire g904_n_spl_;
  wire g905_n_spl_;
  wire g905_p_spl_;
  wire g846_n_spl_;
  wire g907_p_spl_;
  wire g846_p_spl_;
  wire g907_n_spl_;
  wire g908_n_spl_;
  wire g908_p_spl_;
  wire g845_n_spl_;
  wire g910_p_spl_;
  wire g845_p_spl_;
  wire g910_n_spl_;
  wire g911_n_spl_;
  wire g911_p_spl_;
  wire g844_n_spl_;
  wire g913_p_spl_;
  wire g844_p_spl_;
  wire g913_n_spl_;
  wire g914_n_spl_;
  wire g914_p_spl_;
  wire g843_n_spl_;
  wire g916_p_spl_;
  wire g843_p_spl_;
  wire g916_n_spl_;
  wire g917_n_spl_;
  wire g917_p_spl_;
  wire g842_n_spl_;
  wire g919_p_spl_;
  wire g842_p_spl_;
  wire g919_n_spl_;
  wire g920_n_spl_;
  wire g920_p_spl_;
  wire g841_n_spl_;
  wire g922_p_spl_;
  wire g841_p_spl_;
  wire g922_n_spl_;
  wire g923_n_spl_;
  wire g923_p_spl_;
  wire g840_n_spl_;
  wire g925_p_spl_;
  wire g840_p_spl_;
  wire g925_n_spl_;
  wire g926_n_spl_;
  wire g926_p_spl_;
  wire g839_n_spl_;
  wire g928_p_spl_;
  wire g839_p_spl_;
  wire g928_n_spl_;
  wire g929_n_spl_;
  wire g929_p_spl_;
  wire g838_n_spl_;
  wire g931_p_spl_;
  wire g838_p_spl_;
  wire g931_n_spl_;
  wire g932_n_spl_;
  wire g932_p_spl_;
  wire g837_n_spl_;
  wire g934_p_spl_;
  wire g837_p_spl_;
  wire g934_n_spl_;
  wire g935_n_spl_;
  wire g935_p_spl_;
  wire g836_n_spl_;
  wire g937_p_spl_;
  wire g836_p_spl_;
  wire g937_n_spl_;
  wire g938_n_spl_;
  wire g938_p_spl_;
  wire g835_n_spl_;
  wire g940_p_spl_;
  wire g835_p_spl_;
  wire g940_n_spl_;
  wire g941_n_spl_;
  wire g941_p_spl_;
  wire g834_n_spl_;
  wire g943_p_spl_;
  wire g834_p_spl_;
  wire g943_n_spl_;
  wire g944_n_spl_;
  wire g944_p_spl_;
  wire g833_p_spl_;
  wire g946_n_spl_;
  wire g947_p_spl_;
  wire g977_p_spl_;
  wire g977_n_spl_;
  wire g978_p_spl_;
  wire g979_n_spl_;
  wire g978_n_spl_;
  wire g979_p_spl_;
  wire g980_n_spl_;
  wire g980_p_spl_;
  wire g976_n_spl_;
  wire g982_p_spl_;
  wire g976_p_spl_;
  wire g982_n_spl_;
  wire g983_n_spl_;
  wire g983_p_spl_;
  wire g975_n_spl_;
  wire g985_p_spl_;
  wire g975_p_spl_;
  wire g985_n_spl_;
  wire g986_n_spl_;
  wire g986_p_spl_;
  wire g974_n_spl_;
  wire g988_p_spl_;
  wire g974_p_spl_;
  wire g988_n_spl_;
  wire g989_n_spl_;
  wire g989_p_spl_;
  wire g973_n_spl_;
  wire g991_p_spl_;
  wire g973_p_spl_;
  wire g991_n_spl_;
  wire g992_n_spl_;
  wire g992_p_spl_;
  wire g972_n_spl_;
  wire g994_p_spl_;
  wire g972_p_spl_;
  wire g994_n_spl_;
  wire g995_n_spl_;
  wire g995_p_spl_;
  wire g971_n_spl_;
  wire g997_p_spl_;
  wire g971_p_spl_;
  wire g997_n_spl_;
  wire g998_n_spl_;
  wire g998_p_spl_;
  wire g970_n_spl_;
  wire g1000_p_spl_;
  wire g970_p_spl_;
  wire g1000_n_spl_;
  wire g1001_n_spl_;
  wire g1001_p_spl_;
  wire g969_n_spl_;
  wire g1003_p_spl_;
  wire g969_p_spl_;
  wire g1003_n_spl_;
  wire g1004_n_spl_;
  wire g1004_p_spl_;
  wire g968_n_spl_;
  wire g1006_p_spl_;
  wire g968_p_spl_;
  wire g1006_n_spl_;
  wire g1007_n_spl_;
  wire g1007_p_spl_;
  wire g967_n_spl_;
  wire g1009_p_spl_;
  wire g967_p_spl_;
  wire g1009_n_spl_;
  wire g1010_n_spl_;
  wire g1010_p_spl_;
  wire g966_n_spl_;
  wire g1012_p_spl_;
  wire g966_p_spl_;
  wire g1012_n_spl_;
  wire g1013_n_spl_;
  wire g1013_p_spl_;
  wire g965_n_spl_;
  wire g1015_p_spl_;
  wire g965_p_spl_;
  wire g1015_n_spl_;
  wire g1016_n_spl_;
  wire g1016_p_spl_;
  wire g964_n_spl_;
  wire g1018_p_spl_;
  wire g964_p_spl_;
  wire g1018_n_spl_;
  wire g1019_n_spl_;
  wire g1019_p_spl_;
  wire g963_n_spl_;
  wire g1021_p_spl_;
  wire g963_p_spl_;
  wire g1021_n_spl_;
  wire g1022_n_spl_;
  wire g1022_p_spl_;
  wire g962_n_spl_;
  wire g1024_p_spl_;
  wire g962_p_spl_;
  wire g1024_n_spl_;
  wire g1025_n_spl_;
  wire g1025_p_spl_;
  wire g961_n_spl_;
  wire g1027_p_spl_;
  wire g961_p_spl_;
  wire g1027_n_spl_;
  wire g1028_n_spl_;
  wire g1028_p_spl_;
  wire g960_n_spl_;
  wire g1030_p_spl_;
  wire g960_p_spl_;
  wire g1030_n_spl_;
  wire g1031_n_spl_;
  wire g1031_p_spl_;
  wire g959_n_spl_;
  wire g1033_p_spl_;
  wire g959_p_spl_;
  wire g1033_n_spl_;
  wire g1034_n_spl_;
  wire g1034_p_spl_;
  wire g958_n_spl_;
  wire g1036_p_spl_;
  wire g958_p_spl_;
  wire g1036_n_spl_;
  wire g1037_n_spl_;
  wire g1037_p_spl_;
  wire g957_n_spl_;
  wire g1039_p_spl_;
  wire g957_p_spl_;
  wire g1039_n_spl_;
  wire g1040_n_spl_;
  wire g1040_p_spl_;
  wire g956_n_spl_;
  wire g1042_p_spl_;
  wire g956_p_spl_;
  wire g1042_n_spl_;
  wire g1043_n_spl_;
  wire g1043_p_spl_;
  wire g955_n_spl_;
  wire g1045_p_spl_;
  wire g955_p_spl_;
  wire g1045_n_spl_;
  wire g1046_n_spl_;
  wire g1046_p_spl_;
  wire g954_n_spl_;
  wire g1048_p_spl_;
  wire g954_p_spl_;
  wire g1048_n_spl_;
  wire g1049_n_spl_;
  wire g1049_p_spl_;
  wire g953_n_spl_;
  wire g1051_p_spl_;
  wire g953_p_spl_;
  wire g1051_n_spl_;
  wire g1052_n_spl_;
  wire g1052_p_spl_;
  wire g952_n_spl_;
  wire g1054_p_spl_;
  wire g952_p_spl_;
  wire g1054_n_spl_;
  wire g1055_n_spl_;
  wire g1055_p_spl_;
  wire g951_n_spl_;
  wire g1057_p_spl_;
  wire g951_p_spl_;
  wire g1057_n_spl_;
  wire g1058_n_spl_;
  wire g1058_p_spl_;
  wire g950_p_spl_;
  wire g1060_n_spl_;
  wire g1062_n_spl_;
  wire g1090_n_spl_;
  wire g1091_n_spl_;
  wire g1090_p_spl_;
  wire g1091_p_spl_;
  wire g1092_n_spl_;
  wire g1092_p_spl_;
  wire g1089_n_spl_;
  wire g1094_p_spl_;
  wire g1089_p_spl_;
  wire g1094_n_spl_;
  wire g1095_n_spl_;
  wire g1095_p_spl_;
  wire g1088_n_spl_;
  wire g1097_p_spl_;
  wire g1088_p_spl_;
  wire g1097_n_spl_;
  wire g1098_n_spl_;
  wire g1098_p_spl_;
  wire g1087_n_spl_;
  wire g1100_p_spl_;
  wire g1087_p_spl_;
  wire g1100_n_spl_;
  wire g1101_n_spl_;
  wire g1101_p_spl_;
  wire g1086_n_spl_;
  wire g1103_p_spl_;
  wire g1086_p_spl_;
  wire g1103_n_spl_;
  wire g1104_n_spl_;
  wire g1104_p_spl_;
  wire g1085_n_spl_;
  wire g1106_p_spl_;
  wire g1085_p_spl_;
  wire g1106_n_spl_;
  wire g1107_n_spl_;
  wire g1107_p_spl_;
  wire g1084_n_spl_;
  wire g1109_p_spl_;
  wire g1084_p_spl_;
  wire g1109_n_spl_;
  wire g1110_n_spl_;
  wire g1110_p_spl_;
  wire g1083_n_spl_;
  wire g1112_p_spl_;
  wire g1083_p_spl_;
  wire g1112_n_spl_;
  wire g1113_n_spl_;
  wire g1113_p_spl_;
  wire g1082_n_spl_;
  wire g1115_p_spl_;
  wire g1082_p_spl_;
  wire g1115_n_spl_;
  wire g1116_n_spl_;
  wire g1116_p_spl_;
  wire g1081_n_spl_;
  wire g1118_p_spl_;
  wire g1081_p_spl_;
  wire g1118_n_spl_;
  wire g1119_n_spl_;
  wire g1119_p_spl_;
  wire g1080_n_spl_;
  wire g1121_p_spl_;
  wire g1080_p_spl_;
  wire g1121_n_spl_;
  wire g1122_n_spl_;
  wire g1122_p_spl_;
  wire g1079_n_spl_;
  wire g1124_p_spl_;
  wire g1079_p_spl_;
  wire g1124_n_spl_;
  wire g1125_n_spl_;
  wire g1125_p_spl_;
  wire g1078_n_spl_;
  wire g1127_p_spl_;
  wire g1078_p_spl_;
  wire g1127_n_spl_;
  wire g1128_n_spl_;
  wire g1128_p_spl_;
  wire g1077_n_spl_;
  wire g1130_p_spl_;
  wire g1077_p_spl_;
  wire g1130_n_spl_;
  wire g1131_n_spl_;
  wire g1131_p_spl_;
  wire g1076_n_spl_;
  wire g1133_p_spl_;
  wire g1076_p_spl_;
  wire g1133_n_spl_;
  wire g1134_n_spl_;
  wire g1134_p_spl_;
  wire g1075_n_spl_;
  wire g1136_p_spl_;
  wire g1075_p_spl_;
  wire g1136_n_spl_;
  wire g1137_n_spl_;
  wire g1137_p_spl_;
  wire g1074_n_spl_;
  wire g1139_p_spl_;
  wire g1074_p_spl_;
  wire g1139_n_spl_;
  wire g1140_n_spl_;
  wire g1140_p_spl_;
  wire g1073_n_spl_;
  wire g1142_p_spl_;
  wire g1073_p_spl_;
  wire g1142_n_spl_;
  wire g1143_n_spl_;
  wire g1143_p_spl_;
  wire g1072_n_spl_;
  wire g1145_p_spl_;
  wire g1072_p_spl_;
  wire g1145_n_spl_;
  wire g1146_n_spl_;
  wire g1146_p_spl_;
  wire g1071_n_spl_;
  wire g1148_p_spl_;
  wire g1071_p_spl_;
  wire g1148_n_spl_;
  wire g1149_n_spl_;
  wire g1149_p_spl_;
  wire g1070_n_spl_;
  wire g1151_p_spl_;
  wire g1070_p_spl_;
  wire g1151_n_spl_;
  wire g1152_n_spl_;
  wire g1152_p_spl_;
  wire g1069_n_spl_;
  wire g1154_p_spl_;
  wire g1069_p_spl_;
  wire g1154_n_spl_;
  wire g1155_n_spl_;
  wire g1155_p_spl_;
  wire g1068_n_spl_;
  wire g1157_p_spl_;
  wire g1068_p_spl_;
  wire g1157_n_spl_;
  wire g1158_n_spl_;
  wire g1158_p_spl_;
  wire g1067_n_spl_;
  wire g1160_p_spl_;
  wire g1067_p_spl_;
  wire g1160_n_spl_;
  wire g1161_n_spl_;
  wire g1161_p_spl_;
  wire g1066_n_spl_;
  wire g1163_p_spl_;
  wire g1066_p_spl_;
  wire g1163_n_spl_;
  wire g1164_n_spl_;
  wire g1164_p_spl_;
  wire g1065_n_spl_;
  wire g1166_p_spl_;
  wire g1065_p_spl_;
  wire g1166_n_spl_;
  wire g1167_n_spl_;
  wire g1167_p_spl_;
  wire g1064_n_spl_;
  wire g1169_p_spl_;
  wire g1064_p_spl_;
  wire g1169_n_spl_;
  wire g1170_n_spl_;
  wire g1170_p_spl_;
  wire g1062_p_spl_;
  wire g1172_n_spl_;
  wire g1173_p_spl_;
  wire g1201_n_spl_;
  wire g1202_n_spl_;
  wire g1201_p_spl_;
  wire g1202_p_spl_;
  wire g1203_n_spl_;
  wire g1203_p_spl_;
  wire g1200_n_spl_;
  wire g1205_p_spl_;
  wire g1200_p_spl_;
  wire g1205_n_spl_;
  wire g1206_n_spl_;
  wire g1206_p_spl_;
  wire g1199_n_spl_;
  wire g1208_p_spl_;
  wire g1199_p_spl_;
  wire g1208_n_spl_;
  wire g1209_n_spl_;
  wire g1209_p_spl_;
  wire g1198_n_spl_;
  wire g1211_p_spl_;
  wire g1198_p_spl_;
  wire g1211_n_spl_;
  wire g1212_n_spl_;
  wire g1212_p_spl_;
  wire g1197_n_spl_;
  wire g1214_p_spl_;
  wire g1197_p_spl_;
  wire g1214_n_spl_;
  wire g1215_n_spl_;
  wire g1215_p_spl_;
  wire g1196_n_spl_;
  wire g1217_p_spl_;
  wire g1196_p_spl_;
  wire g1217_n_spl_;
  wire g1218_n_spl_;
  wire g1218_p_spl_;
  wire g1195_n_spl_;
  wire g1220_p_spl_;
  wire g1195_p_spl_;
  wire g1220_n_spl_;
  wire g1221_n_spl_;
  wire g1221_p_spl_;
  wire g1194_n_spl_;
  wire g1223_p_spl_;
  wire g1194_p_spl_;
  wire g1223_n_spl_;
  wire g1224_n_spl_;
  wire g1224_p_spl_;
  wire g1193_n_spl_;
  wire g1226_p_spl_;
  wire g1193_p_spl_;
  wire g1226_n_spl_;
  wire g1227_n_spl_;
  wire g1227_p_spl_;
  wire g1192_n_spl_;
  wire g1229_p_spl_;
  wire g1192_p_spl_;
  wire g1229_n_spl_;
  wire g1230_n_spl_;
  wire g1230_p_spl_;
  wire g1191_n_spl_;
  wire g1232_p_spl_;
  wire g1191_p_spl_;
  wire g1232_n_spl_;
  wire g1233_n_spl_;
  wire g1233_p_spl_;
  wire g1190_n_spl_;
  wire g1235_p_spl_;
  wire g1190_p_spl_;
  wire g1235_n_spl_;
  wire g1236_n_spl_;
  wire g1236_p_spl_;
  wire g1189_n_spl_;
  wire g1238_p_spl_;
  wire g1189_p_spl_;
  wire g1238_n_spl_;
  wire g1239_n_spl_;
  wire g1239_p_spl_;
  wire g1188_n_spl_;
  wire g1241_p_spl_;
  wire g1188_p_spl_;
  wire g1241_n_spl_;
  wire g1242_n_spl_;
  wire g1242_p_spl_;
  wire g1187_n_spl_;
  wire g1244_p_spl_;
  wire g1187_p_spl_;
  wire g1244_n_spl_;
  wire g1245_n_spl_;
  wire g1245_p_spl_;
  wire g1186_n_spl_;
  wire g1247_p_spl_;
  wire g1186_p_spl_;
  wire g1247_n_spl_;
  wire g1248_n_spl_;
  wire g1248_p_spl_;
  wire g1185_n_spl_;
  wire g1250_p_spl_;
  wire g1185_p_spl_;
  wire g1250_n_spl_;
  wire g1251_n_spl_;
  wire g1251_p_spl_;
  wire g1184_n_spl_;
  wire g1253_p_spl_;
  wire g1184_p_spl_;
  wire g1253_n_spl_;
  wire g1254_n_spl_;
  wire g1254_p_spl_;
  wire g1183_n_spl_;
  wire g1256_p_spl_;
  wire g1183_p_spl_;
  wire g1256_n_spl_;
  wire g1257_n_spl_;
  wire g1257_p_spl_;
  wire g1182_n_spl_;
  wire g1259_p_spl_;
  wire g1182_p_spl_;
  wire g1259_n_spl_;
  wire g1260_n_spl_;
  wire g1260_p_spl_;
  wire g1181_n_spl_;
  wire g1262_p_spl_;
  wire g1181_p_spl_;
  wire g1262_n_spl_;
  wire g1263_n_spl_;
  wire g1263_p_spl_;
  wire g1180_n_spl_;
  wire g1265_p_spl_;
  wire g1180_p_spl_;
  wire g1265_n_spl_;
  wire g1266_n_spl_;
  wire g1266_p_spl_;
  wire g1179_n_spl_;
  wire g1268_p_spl_;
  wire g1179_p_spl_;
  wire g1268_n_spl_;
  wire g1269_n_spl_;
  wire g1269_p_spl_;
  wire g1178_n_spl_;
  wire g1271_p_spl_;
  wire g1178_p_spl_;
  wire g1271_n_spl_;
  wire g1272_n_spl_;
  wire g1272_p_spl_;
  wire g1177_n_spl_;
  wire g1274_p_spl_;
  wire g1177_p_spl_;
  wire g1274_n_spl_;
  wire g1275_n_spl_;
  wire g1275_p_spl_;
  wire g1176_p_spl_;
  wire g1277_n_spl_;
  wire g1278_p_spl_;
  wire g1304_n_spl_;
  wire g1305_n_spl_;
  wire g1304_p_spl_;
  wire g1305_p_spl_;
  wire g1306_n_spl_;
  wire g1306_p_spl_;
  wire g1303_n_spl_;
  wire g1308_p_spl_;
  wire g1303_p_spl_;
  wire g1308_n_spl_;
  wire g1309_n_spl_;
  wire g1309_p_spl_;
  wire g1302_n_spl_;
  wire g1311_p_spl_;
  wire g1302_p_spl_;
  wire g1311_n_spl_;
  wire g1312_n_spl_;
  wire g1312_p_spl_;
  wire g1301_n_spl_;
  wire g1314_p_spl_;
  wire g1301_p_spl_;
  wire g1314_n_spl_;
  wire g1315_n_spl_;
  wire g1315_p_spl_;
  wire g1300_n_spl_;
  wire g1317_p_spl_;
  wire g1300_p_spl_;
  wire g1317_n_spl_;
  wire g1318_n_spl_;
  wire g1318_p_spl_;
  wire g1299_n_spl_;
  wire g1320_p_spl_;
  wire g1299_p_spl_;
  wire g1320_n_spl_;
  wire g1321_n_spl_;
  wire g1321_p_spl_;
  wire g1298_n_spl_;
  wire g1323_p_spl_;
  wire g1298_p_spl_;
  wire g1323_n_spl_;
  wire g1324_n_spl_;
  wire g1324_p_spl_;
  wire g1297_n_spl_;
  wire g1326_p_spl_;
  wire g1297_p_spl_;
  wire g1326_n_spl_;
  wire g1327_n_spl_;
  wire g1327_p_spl_;
  wire g1296_n_spl_;
  wire g1329_p_spl_;
  wire g1296_p_spl_;
  wire g1329_n_spl_;
  wire g1330_n_spl_;
  wire g1330_p_spl_;
  wire g1295_n_spl_;
  wire g1332_p_spl_;
  wire g1295_p_spl_;
  wire g1332_n_spl_;
  wire g1333_n_spl_;
  wire g1333_p_spl_;
  wire g1294_n_spl_;
  wire g1335_p_spl_;
  wire g1294_p_spl_;
  wire g1335_n_spl_;
  wire g1336_n_spl_;
  wire g1336_p_spl_;
  wire g1293_n_spl_;
  wire g1338_p_spl_;
  wire g1293_p_spl_;
  wire g1338_n_spl_;
  wire g1339_n_spl_;
  wire g1339_p_spl_;
  wire g1292_n_spl_;
  wire g1341_p_spl_;
  wire g1292_p_spl_;
  wire g1341_n_spl_;
  wire g1342_n_spl_;
  wire g1342_p_spl_;
  wire g1291_n_spl_;
  wire g1344_p_spl_;
  wire g1291_p_spl_;
  wire g1344_n_spl_;
  wire g1345_n_spl_;
  wire g1345_p_spl_;
  wire g1290_n_spl_;
  wire g1347_p_spl_;
  wire g1290_p_spl_;
  wire g1347_n_spl_;
  wire g1348_n_spl_;
  wire g1348_p_spl_;
  wire g1289_n_spl_;
  wire g1350_p_spl_;
  wire g1289_p_spl_;
  wire g1350_n_spl_;
  wire g1351_n_spl_;
  wire g1351_p_spl_;
  wire g1288_n_spl_;
  wire g1353_p_spl_;
  wire g1288_p_spl_;
  wire g1353_n_spl_;
  wire g1354_n_spl_;
  wire g1354_p_spl_;
  wire g1287_n_spl_;
  wire g1356_p_spl_;
  wire g1287_p_spl_;
  wire g1356_n_spl_;
  wire g1357_n_spl_;
  wire g1357_p_spl_;
  wire g1286_n_spl_;
  wire g1359_p_spl_;
  wire g1286_p_spl_;
  wire g1359_n_spl_;
  wire g1360_n_spl_;
  wire g1360_p_spl_;
  wire g1285_n_spl_;
  wire g1362_p_spl_;
  wire g1285_p_spl_;
  wire g1362_n_spl_;
  wire g1363_n_spl_;
  wire g1363_p_spl_;
  wire g1284_n_spl_;
  wire g1365_p_spl_;
  wire g1284_p_spl_;
  wire g1365_n_spl_;
  wire g1366_n_spl_;
  wire g1366_p_spl_;
  wire g1283_n_spl_;
  wire g1368_p_spl_;
  wire g1283_p_spl_;
  wire g1368_n_spl_;
  wire g1369_n_spl_;
  wire g1369_p_spl_;
  wire g1282_n_spl_;
  wire g1371_p_spl_;
  wire g1282_p_spl_;
  wire g1371_n_spl_;
  wire g1372_n_spl_;
  wire g1372_p_spl_;
  wire g1281_p_spl_;
  wire g1374_n_spl_;
  wire g1375_p_spl_;
  wire g1399_n_spl_;
  wire g1400_n_spl_;
  wire g1399_p_spl_;
  wire g1400_p_spl_;
  wire g1401_n_spl_;
  wire g1401_p_spl_;
  wire g1398_n_spl_;
  wire g1403_p_spl_;
  wire g1398_p_spl_;
  wire g1403_n_spl_;
  wire g1404_n_spl_;
  wire g1404_p_spl_;
  wire g1397_n_spl_;
  wire g1406_p_spl_;
  wire g1397_p_spl_;
  wire g1406_n_spl_;
  wire g1407_n_spl_;
  wire g1407_p_spl_;
  wire g1396_n_spl_;
  wire g1409_p_spl_;
  wire g1396_p_spl_;
  wire g1409_n_spl_;
  wire g1410_n_spl_;
  wire g1410_p_spl_;
  wire g1395_n_spl_;
  wire g1412_p_spl_;
  wire g1395_p_spl_;
  wire g1412_n_spl_;
  wire g1413_n_spl_;
  wire g1413_p_spl_;
  wire g1394_n_spl_;
  wire g1415_p_spl_;
  wire g1394_p_spl_;
  wire g1415_n_spl_;
  wire g1416_n_spl_;
  wire g1416_p_spl_;
  wire g1393_n_spl_;
  wire g1418_p_spl_;
  wire g1393_p_spl_;
  wire g1418_n_spl_;
  wire g1419_n_spl_;
  wire g1419_p_spl_;
  wire g1392_n_spl_;
  wire g1421_p_spl_;
  wire g1392_p_spl_;
  wire g1421_n_spl_;
  wire g1422_n_spl_;
  wire g1422_p_spl_;
  wire g1391_n_spl_;
  wire g1424_p_spl_;
  wire g1391_p_spl_;
  wire g1424_n_spl_;
  wire g1425_n_spl_;
  wire g1425_p_spl_;
  wire g1390_n_spl_;
  wire g1427_p_spl_;
  wire g1390_p_spl_;
  wire g1427_n_spl_;
  wire g1428_n_spl_;
  wire g1428_p_spl_;
  wire g1389_n_spl_;
  wire g1430_p_spl_;
  wire g1389_p_spl_;
  wire g1430_n_spl_;
  wire g1431_n_spl_;
  wire g1431_p_spl_;
  wire g1388_n_spl_;
  wire g1433_p_spl_;
  wire g1388_p_spl_;
  wire g1433_n_spl_;
  wire g1434_n_spl_;
  wire g1434_p_spl_;
  wire g1387_n_spl_;
  wire g1436_p_spl_;
  wire g1387_p_spl_;
  wire g1436_n_spl_;
  wire g1437_n_spl_;
  wire g1437_p_spl_;
  wire g1386_n_spl_;
  wire g1439_p_spl_;
  wire g1386_p_spl_;
  wire g1439_n_spl_;
  wire g1440_n_spl_;
  wire g1440_p_spl_;
  wire g1385_n_spl_;
  wire g1442_p_spl_;
  wire g1385_p_spl_;
  wire g1442_n_spl_;
  wire g1443_n_spl_;
  wire g1443_p_spl_;
  wire g1384_n_spl_;
  wire g1445_p_spl_;
  wire g1384_p_spl_;
  wire g1445_n_spl_;
  wire g1446_n_spl_;
  wire g1446_p_spl_;
  wire g1383_n_spl_;
  wire g1448_p_spl_;
  wire g1383_p_spl_;
  wire g1448_n_spl_;
  wire g1449_n_spl_;
  wire g1449_p_spl_;
  wire g1382_n_spl_;
  wire g1451_p_spl_;
  wire g1382_p_spl_;
  wire g1451_n_spl_;
  wire g1452_n_spl_;
  wire g1452_p_spl_;
  wire g1381_n_spl_;
  wire g1454_p_spl_;
  wire g1381_p_spl_;
  wire g1454_n_spl_;
  wire g1455_n_spl_;
  wire g1455_p_spl_;
  wire g1380_n_spl_;
  wire g1457_p_spl_;
  wire g1380_p_spl_;
  wire g1457_n_spl_;
  wire g1458_n_spl_;
  wire g1458_p_spl_;
  wire g1379_n_spl_;
  wire g1460_p_spl_;
  wire g1379_p_spl_;
  wire g1460_n_spl_;
  wire g1461_n_spl_;
  wire g1461_p_spl_;
  wire g1378_p_spl_;
  wire g1463_n_spl_;
  wire g1464_p_spl_;
  wire g1486_n_spl_;
  wire g1487_n_spl_;
  wire g1486_p_spl_;
  wire g1487_p_spl_;
  wire g1488_n_spl_;
  wire g1488_p_spl_;
  wire g1485_n_spl_;
  wire g1490_p_spl_;
  wire g1485_p_spl_;
  wire g1490_n_spl_;
  wire g1491_n_spl_;
  wire g1491_p_spl_;
  wire g1484_n_spl_;
  wire g1493_p_spl_;
  wire g1484_p_spl_;
  wire g1493_n_spl_;
  wire g1494_n_spl_;
  wire g1494_p_spl_;
  wire g1483_n_spl_;
  wire g1496_p_spl_;
  wire g1483_p_spl_;
  wire g1496_n_spl_;
  wire g1497_n_spl_;
  wire g1497_p_spl_;
  wire g1482_n_spl_;
  wire g1499_p_spl_;
  wire g1482_p_spl_;
  wire g1499_n_spl_;
  wire g1500_n_spl_;
  wire g1500_p_spl_;
  wire g1481_n_spl_;
  wire g1502_p_spl_;
  wire g1481_p_spl_;
  wire g1502_n_spl_;
  wire g1503_n_spl_;
  wire g1503_p_spl_;
  wire g1480_n_spl_;
  wire g1505_p_spl_;
  wire g1480_p_spl_;
  wire g1505_n_spl_;
  wire g1506_n_spl_;
  wire g1506_p_spl_;
  wire g1479_n_spl_;
  wire g1508_p_spl_;
  wire g1479_p_spl_;
  wire g1508_n_spl_;
  wire g1509_n_spl_;
  wire g1509_p_spl_;
  wire g1478_n_spl_;
  wire g1511_p_spl_;
  wire g1478_p_spl_;
  wire g1511_n_spl_;
  wire g1512_n_spl_;
  wire g1512_p_spl_;
  wire g1477_n_spl_;
  wire g1514_p_spl_;
  wire g1477_p_spl_;
  wire g1514_n_spl_;
  wire g1515_n_spl_;
  wire g1515_p_spl_;
  wire g1476_n_spl_;
  wire g1517_p_spl_;
  wire g1476_p_spl_;
  wire g1517_n_spl_;
  wire g1518_n_spl_;
  wire g1518_p_spl_;
  wire g1475_n_spl_;
  wire g1520_p_spl_;
  wire g1475_p_spl_;
  wire g1520_n_spl_;
  wire g1521_n_spl_;
  wire g1521_p_spl_;
  wire g1474_n_spl_;
  wire g1523_p_spl_;
  wire g1474_p_spl_;
  wire g1523_n_spl_;
  wire g1524_n_spl_;
  wire g1524_p_spl_;
  wire g1473_n_spl_;
  wire g1526_p_spl_;
  wire g1473_p_spl_;
  wire g1526_n_spl_;
  wire g1527_n_spl_;
  wire g1527_p_spl_;
  wire g1472_n_spl_;
  wire g1529_p_spl_;
  wire g1472_p_spl_;
  wire g1529_n_spl_;
  wire g1530_n_spl_;
  wire g1530_p_spl_;
  wire g1471_n_spl_;
  wire g1532_p_spl_;
  wire g1471_p_spl_;
  wire g1532_n_spl_;
  wire g1533_n_spl_;
  wire g1533_p_spl_;
  wire g1470_n_spl_;
  wire g1535_p_spl_;
  wire g1470_p_spl_;
  wire g1535_n_spl_;
  wire g1536_n_spl_;
  wire g1536_p_spl_;
  wire g1469_n_spl_;
  wire g1538_p_spl_;
  wire g1469_p_spl_;
  wire g1538_n_spl_;
  wire g1539_n_spl_;
  wire g1539_p_spl_;
  wire g1468_n_spl_;
  wire g1541_p_spl_;
  wire g1468_p_spl_;
  wire g1541_n_spl_;
  wire g1542_n_spl_;
  wire g1542_p_spl_;
  wire g1467_p_spl_;
  wire g1544_n_spl_;
  wire g1545_p_spl_;
  wire g1565_n_spl_;
  wire g1566_n_spl_;
  wire g1565_p_spl_;
  wire g1566_p_spl_;
  wire g1567_n_spl_;
  wire g1567_p_spl_;
  wire g1564_n_spl_;
  wire g1569_p_spl_;
  wire g1564_p_spl_;
  wire g1569_n_spl_;
  wire g1570_n_spl_;
  wire g1570_p_spl_;
  wire g1563_n_spl_;
  wire g1572_p_spl_;
  wire g1563_p_spl_;
  wire g1572_n_spl_;
  wire g1573_n_spl_;
  wire g1573_p_spl_;
  wire g1562_n_spl_;
  wire g1575_p_spl_;
  wire g1562_p_spl_;
  wire g1575_n_spl_;
  wire g1576_n_spl_;
  wire g1576_p_spl_;
  wire g1561_n_spl_;
  wire g1578_p_spl_;
  wire g1561_p_spl_;
  wire g1578_n_spl_;
  wire g1579_n_spl_;
  wire g1579_p_spl_;
  wire g1560_n_spl_;
  wire g1581_p_spl_;
  wire g1560_p_spl_;
  wire g1581_n_spl_;
  wire g1582_n_spl_;
  wire g1582_p_spl_;
  wire g1559_n_spl_;
  wire g1584_p_spl_;
  wire g1559_p_spl_;
  wire g1584_n_spl_;
  wire g1585_n_spl_;
  wire g1585_p_spl_;
  wire g1558_n_spl_;
  wire g1587_p_spl_;
  wire g1558_p_spl_;
  wire g1587_n_spl_;
  wire g1588_n_spl_;
  wire g1588_p_spl_;
  wire g1557_n_spl_;
  wire g1590_p_spl_;
  wire g1557_p_spl_;
  wire g1590_n_spl_;
  wire g1591_n_spl_;
  wire g1591_p_spl_;
  wire g1556_n_spl_;
  wire g1593_p_spl_;
  wire g1556_p_spl_;
  wire g1593_n_spl_;
  wire g1594_n_spl_;
  wire g1594_p_spl_;
  wire g1555_n_spl_;
  wire g1596_p_spl_;
  wire g1555_p_spl_;
  wire g1596_n_spl_;
  wire g1597_n_spl_;
  wire g1597_p_spl_;
  wire g1554_n_spl_;
  wire g1599_p_spl_;
  wire g1554_p_spl_;
  wire g1599_n_spl_;
  wire g1600_n_spl_;
  wire g1600_p_spl_;
  wire g1553_n_spl_;
  wire g1602_p_spl_;
  wire g1553_p_spl_;
  wire g1602_n_spl_;
  wire g1603_n_spl_;
  wire g1603_p_spl_;
  wire g1552_n_spl_;
  wire g1605_p_spl_;
  wire g1552_p_spl_;
  wire g1605_n_spl_;
  wire g1606_n_spl_;
  wire g1606_p_spl_;
  wire g1551_n_spl_;
  wire g1608_p_spl_;
  wire g1551_p_spl_;
  wire g1608_n_spl_;
  wire g1609_n_spl_;
  wire g1609_p_spl_;
  wire g1550_n_spl_;
  wire g1611_p_spl_;
  wire g1550_p_spl_;
  wire g1611_n_spl_;
  wire g1612_n_spl_;
  wire g1612_p_spl_;
  wire g1549_n_spl_;
  wire g1614_p_spl_;
  wire g1549_p_spl_;
  wire g1614_n_spl_;
  wire g1615_n_spl_;
  wire g1615_p_spl_;
  wire g1548_p_spl_;
  wire g1617_n_spl_;
  wire g1618_p_spl_;
  wire g1636_n_spl_;
  wire g1637_n_spl_;
  wire g1636_p_spl_;
  wire g1637_p_spl_;
  wire g1638_n_spl_;
  wire g1638_p_spl_;
  wire g1635_n_spl_;
  wire g1640_p_spl_;
  wire g1635_p_spl_;
  wire g1640_n_spl_;
  wire g1641_n_spl_;
  wire g1641_p_spl_;
  wire g1634_n_spl_;
  wire g1643_p_spl_;
  wire g1634_p_spl_;
  wire g1643_n_spl_;
  wire g1644_n_spl_;
  wire g1644_p_spl_;
  wire g1633_n_spl_;
  wire g1646_p_spl_;
  wire g1633_p_spl_;
  wire g1646_n_spl_;
  wire g1647_n_spl_;
  wire g1647_p_spl_;
  wire g1632_n_spl_;
  wire g1649_p_spl_;
  wire g1632_p_spl_;
  wire g1649_n_spl_;
  wire g1650_n_spl_;
  wire g1650_p_spl_;
  wire g1631_n_spl_;
  wire g1652_p_spl_;
  wire g1631_p_spl_;
  wire g1652_n_spl_;
  wire g1653_n_spl_;
  wire g1653_p_spl_;
  wire g1630_n_spl_;
  wire g1655_p_spl_;
  wire g1630_p_spl_;
  wire g1655_n_spl_;
  wire g1656_n_spl_;
  wire g1656_p_spl_;
  wire g1629_n_spl_;
  wire g1658_p_spl_;
  wire g1629_p_spl_;
  wire g1658_n_spl_;
  wire g1659_n_spl_;
  wire g1659_p_spl_;
  wire g1628_n_spl_;
  wire g1661_p_spl_;
  wire g1628_p_spl_;
  wire g1661_n_spl_;
  wire g1662_n_spl_;
  wire g1662_p_spl_;
  wire g1627_n_spl_;
  wire g1664_p_spl_;
  wire g1627_p_spl_;
  wire g1664_n_spl_;
  wire g1665_n_spl_;
  wire g1665_p_spl_;
  wire g1626_n_spl_;
  wire g1667_p_spl_;
  wire g1626_p_spl_;
  wire g1667_n_spl_;
  wire g1668_n_spl_;
  wire g1668_p_spl_;
  wire g1625_n_spl_;
  wire g1670_p_spl_;
  wire g1625_p_spl_;
  wire g1670_n_spl_;
  wire g1671_n_spl_;
  wire g1671_p_spl_;
  wire g1624_n_spl_;
  wire g1673_p_spl_;
  wire g1624_p_spl_;
  wire g1673_n_spl_;
  wire g1674_n_spl_;
  wire g1674_p_spl_;
  wire g1623_n_spl_;
  wire g1676_p_spl_;
  wire g1623_p_spl_;
  wire g1676_n_spl_;
  wire g1677_n_spl_;
  wire g1677_p_spl_;
  wire g1622_n_spl_;
  wire g1679_p_spl_;
  wire g1622_p_spl_;
  wire g1679_n_spl_;
  wire g1680_n_spl_;
  wire g1680_p_spl_;
  wire g1621_p_spl_;
  wire g1682_n_spl_;
  wire g1683_p_spl_;
  wire g1699_n_spl_;
  wire g1700_n_spl_;
  wire g1699_p_spl_;
  wire g1700_p_spl_;
  wire g1701_n_spl_;
  wire g1701_p_spl_;
  wire g1698_n_spl_;
  wire g1703_p_spl_;
  wire g1698_p_spl_;
  wire g1703_n_spl_;
  wire g1704_n_spl_;
  wire g1704_p_spl_;
  wire g1697_n_spl_;
  wire g1706_p_spl_;
  wire g1697_p_spl_;
  wire g1706_n_spl_;
  wire g1707_n_spl_;
  wire g1707_p_spl_;
  wire g1696_n_spl_;
  wire g1709_p_spl_;
  wire g1696_p_spl_;
  wire g1709_n_spl_;
  wire g1710_n_spl_;
  wire g1710_p_spl_;
  wire g1695_n_spl_;
  wire g1712_p_spl_;
  wire g1695_p_spl_;
  wire g1712_n_spl_;
  wire g1713_n_spl_;
  wire g1713_p_spl_;
  wire g1694_n_spl_;
  wire g1715_p_spl_;
  wire g1694_p_spl_;
  wire g1715_n_spl_;
  wire g1716_n_spl_;
  wire g1716_p_spl_;
  wire g1693_n_spl_;
  wire g1718_p_spl_;
  wire g1693_p_spl_;
  wire g1718_n_spl_;
  wire g1719_n_spl_;
  wire g1719_p_spl_;
  wire g1692_n_spl_;
  wire g1721_p_spl_;
  wire g1692_p_spl_;
  wire g1721_n_spl_;
  wire g1722_n_spl_;
  wire g1722_p_spl_;
  wire g1691_n_spl_;
  wire g1724_p_spl_;
  wire g1691_p_spl_;
  wire g1724_n_spl_;
  wire g1725_n_spl_;
  wire g1725_p_spl_;
  wire g1690_n_spl_;
  wire g1727_p_spl_;
  wire g1690_p_spl_;
  wire g1727_n_spl_;
  wire g1728_n_spl_;
  wire g1728_p_spl_;
  wire g1689_n_spl_;
  wire g1730_p_spl_;
  wire g1689_p_spl_;
  wire g1730_n_spl_;
  wire g1731_n_spl_;
  wire g1731_p_spl_;
  wire g1688_n_spl_;
  wire g1733_p_spl_;
  wire g1688_p_spl_;
  wire g1733_n_spl_;
  wire g1734_n_spl_;
  wire g1734_p_spl_;
  wire g1687_n_spl_;
  wire g1736_p_spl_;
  wire g1687_p_spl_;
  wire g1736_n_spl_;
  wire g1737_n_spl_;
  wire g1737_p_spl_;
  wire g1686_p_spl_;
  wire g1739_n_spl_;
  wire g1740_p_spl_;
  wire g1754_n_spl_;
  wire g1755_n_spl_;
  wire g1754_p_spl_;
  wire g1755_p_spl_;
  wire g1756_n_spl_;
  wire g1756_p_spl_;
  wire g1753_n_spl_;
  wire g1758_p_spl_;
  wire g1753_p_spl_;
  wire g1758_n_spl_;
  wire g1759_n_spl_;
  wire g1759_p_spl_;
  wire g1752_n_spl_;
  wire g1761_p_spl_;
  wire g1752_p_spl_;
  wire g1761_n_spl_;
  wire g1762_n_spl_;
  wire g1762_p_spl_;
  wire g1751_n_spl_;
  wire g1764_p_spl_;
  wire g1751_p_spl_;
  wire g1764_n_spl_;
  wire g1765_n_spl_;
  wire g1765_p_spl_;
  wire g1750_n_spl_;
  wire g1767_p_spl_;
  wire g1750_p_spl_;
  wire g1767_n_spl_;
  wire g1768_n_spl_;
  wire g1768_p_spl_;
  wire g1749_n_spl_;
  wire g1770_p_spl_;
  wire g1749_p_spl_;
  wire g1770_n_spl_;
  wire g1771_n_spl_;
  wire g1771_p_spl_;
  wire g1748_n_spl_;
  wire g1773_p_spl_;
  wire g1748_p_spl_;
  wire g1773_n_spl_;
  wire g1774_n_spl_;
  wire g1774_p_spl_;
  wire g1747_n_spl_;
  wire g1776_p_spl_;
  wire g1747_p_spl_;
  wire g1776_n_spl_;
  wire g1777_n_spl_;
  wire g1777_p_spl_;
  wire g1746_n_spl_;
  wire g1779_p_spl_;
  wire g1746_p_spl_;
  wire g1779_n_spl_;
  wire g1780_n_spl_;
  wire g1780_p_spl_;
  wire g1745_n_spl_;
  wire g1782_p_spl_;
  wire g1745_p_spl_;
  wire g1782_n_spl_;
  wire g1783_n_spl_;
  wire g1783_p_spl_;
  wire g1744_n_spl_;
  wire g1785_p_spl_;
  wire g1744_p_spl_;
  wire g1785_n_spl_;
  wire g1786_n_spl_;
  wire g1786_p_spl_;
  wire g1743_p_spl_;
  wire g1788_n_spl_;
  wire g1789_p_spl_;
  wire g1801_n_spl_;
  wire g1802_n_spl_;
  wire g1801_p_spl_;
  wire g1802_p_spl_;
  wire g1803_n_spl_;
  wire g1803_p_spl_;
  wire g1800_n_spl_;
  wire g1805_p_spl_;
  wire g1800_p_spl_;
  wire g1805_n_spl_;
  wire g1806_n_spl_;
  wire g1806_p_spl_;
  wire g1799_n_spl_;
  wire g1808_p_spl_;
  wire g1799_p_spl_;
  wire g1808_n_spl_;
  wire g1809_n_spl_;
  wire g1809_p_spl_;
  wire g1798_n_spl_;
  wire g1811_p_spl_;
  wire g1798_p_spl_;
  wire g1811_n_spl_;
  wire g1812_n_spl_;
  wire g1812_p_spl_;
  wire g1797_n_spl_;
  wire g1814_p_spl_;
  wire g1797_p_spl_;
  wire g1814_n_spl_;
  wire g1815_n_spl_;
  wire g1815_p_spl_;
  wire g1796_n_spl_;
  wire g1817_p_spl_;
  wire g1796_p_spl_;
  wire g1817_n_spl_;
  wire g1818_n_spl_;
  wire g1818_p_spl_;
  wire g1795_n_spl_;
  wire g1820_p_spl_;
  wire g1795_p_spl_;
  wire g1820_n_spl_;
  wire g1821_n_spl_;
  wire g1821_p_spl_;
  wire g1794_n_spl_;
  wire g1823_p_spl_;
  wire g1794_p_spl_;
  wire g1823_n_spl_;
  wire g1824_n_spl_;
  wire g1824_p_spl_;
  wire g1793_n_spl_;
  wire g1826_p_spl_;
  wire g1793_p_spl_;
  wire g1826_n_spl_;
  wire g1827_n_spl_;
  wire g1827_p_spl_;
  wire g1792_p_spl_;
  wire g1829_n_spl_;
  wire g1830_p_spl_;
  wire g1840_n_spl_;
  wire g1841_n_spl_;
  wire g1840_p_spl_;
  wire g1841_p_spl_;
  wire g1842_n_spl_;
  wire g1842_p_spl_;
  wire g1839_n_spl_;
  wire g1844_p_spl_;
  wire g1839_p_spl_;
  wire g1844_n_spl_;
  wire g1845_n_spl_;
  wire g1845_p_spl_;
  wire g1838_n_spl_;
  wire g1847_p_spl_;
  wire g1838_p_spl_;
  wire g1847_n_spl_;
  wire g1848_n_spl_;
  wire g1848_p_spl_;
  wire g1837_n_spl_;
  wire g1850_p_spl_;
  wire g1837_p_spl_;
  wire g1850_n_spl_;
  wire g1851_n_spl_;
  wire g1851_p_spl_;
  wire g1836_n_spl_;
  wire g1853_p_spl_;
  wire g1836_p_spl_;
  wire g1853_n_spl_;
  wire g1854_n_spl_;
  wire g1854_p_spl_;
  wire g1835_n_spl_;
  wire g1856_p_spl_;
  wire g1835_p_spl_;
  wire g1856_n_spl_;
  wire g1857_n_spl_;
  wire g1857_p_spl_;
  wire g1834_n_spl_;
  wire g1859_p_spl_;
  wire g1834_p_spl_;
  wire g1859_n_spl_;
  wire g1860_n_spl_;
  wire g1860_p_spl_;
  wire g1833_p_spl_;
  wire g1862_n_spl_;
  wire g1863_p_spl_;
  wire g1871_n_spl_;
  wire g1872_n_spl_;
  wire g1871_p_spl_;
  wire g1872_p_spl_;
  wire g1873_n_spl_;
  wire g1873_p_spl_;
  wire g1870_n_spl_;
  wire g1875_p_spl_;
  wire g1870_p_spl_;
  wire g1875_n_spl_;
  wire g1876_n_spl_;
  wire g1876_p_spl_;
  wire g1869_n_spl_;
  wire g1878_p_spl_;
  wire g1869_p_spl_;
  wire g1878_n_spl_;
  wire g1879_n_spl_;
  wire g1879_p_spl_;
  wire g1868_n_spl_;
  wire g1881_p_spl_;
  wire g1868_p_spl_;
  wire g1881_n_spl_;
  wire g1882_n_spl_;
  wire g1882_p_spl_;
  wire g1867_n_spl_;
  wire g1884_p_spl_;
  wire g1867_p_spl_;
  wire g1884_n_spl_;
  wire g1885_n_spl_;
  wire g1885_p_spl_;
  wire g1866_p_spl_;
  wire g1887_n_spl_;
  wire g1888_p_spl_;
  wire g1894_n_spl_;
  wire g1895_n_spl_;
  wire g1894_p_spl_;
  wire g1895_p_spl_;
  wire g1896_n_spl_;
  wire g1896_p_spl_;
  wire g1893_n_spl_;
  wire g1898_p_spl_;
  wire g1893_p_spl_;
  wire g1898_n_spl_;
  wire g1899_n_spl_;
  wire g1899_p_spl_;
  wire g1892_n_spl_;
  wire g1901_p_spl_;
  wire g1892_p_spl_;
  wire g1901_n_spl_;
  wire g1902_n_spl_;
  wire g1902_p_spl_;
  wire g1891_p_spl_;
  wire g1904_n_spl_;
  wire g1905_p_spl_;
  wire g1908_n_spl_;
  wire g1909_n_spl_;
  wire g1908_p_spl_;
  wire g1909_p_spl_;
  wire g1910_n_spl_;
  wire g1914_n_spl_;

  LA
  g_g33_p
  (
    .dout(g33_p),
    .din1(G1_p_spl_000),
    .din2(G17_p_spl_000)
  );


  LA
  g_g34_p
  (
    .dout(g34_p),
    .din1(G2_p_spl_000),
    .din2(G17_p_spl_000)
  );


  FA
  g_g34_n
  (
    .dout(g34_n),
    .din1(G2_n_spl_000),
    .din2(G17_n_spl_000)
  );


  LA
  g_g35_p
  (
    .dout(g35_p),
    .din1(G1_p_spl_000),
    .din2(G18_p_spl_000)
  );


  FA
  g_g35_n
  (
    .dout(g35_n),
    .din1(G1_n_spl_000),
    .din2(G18_n_spl_000)
  );


  LA
  g_g36_p
  (
    .dout(g36_p),
    .din1(g34_p_spl_),
    .din2(g35_n)
  );


  FA
  g_g36_n
  (
    .dout(g36_n),
    .din1(g34_n_spl_),
    .din2(g35_p_spl_)
  );


  LA
  g_g37_p
  (
    .dout(g37_p),
    .din1(g34_p_spl_),
    .din2(g36_n)
  );


  FA
  g_g37_n
  (
    .dout(g37_n),
    .din1(g34_n_spl_),
    .din2(g36_p_spl_)
  );


  FA
  g_g38_n
  (
    .dout(g38_n),
    .din1(g35_p_spl_),
    .din2(g36_p_spl_)
  );


  LA
  g_g39_p
  (
    .dout(g39_p),
    .din1(g37_n_spl_0),
    .din2(g38_n)
  );


  LA
  g_g40_p
  (
    .dout(g40_p),
    .din1(G1_p_spl_001),
    .din2(G19_p_spl_000)
  );


  FA
  g_g40_n
  (
    .dout(g40_n),
    .din1(G1_n_spl_000),
    .din2(G19_n_spl_000)
  );


  LA
  g_g41_p
  (
    .dout(g41_p),
    .din1(G3_p_spl_000),
    .din2(G17_p_spl_001)
  );


  FA
  g_g41_n
  (
    .dout(g41_n),
    .din1(G3_n_spl_000),
    .din2(G17_n_spl_000)
  );


  LA
  g_g42_p
  (
    .dout(g42_p),
    .din1(G2_p_spl_000),
    .din2(G18_p_spl_000)
  );


  FA
  g_g42_n
  (
    .dout(g42_n),
    .din1(G2_n_spl_000),
    .din2(G18_n_spl_000)
  );


  LA
  g_g43_p
  (
    .dout(g43_p),
    .din1(g41_p_spl_),
    .din2(g42_n_spl_)
  );


  FA
  g_g43_n
  (
    .dout(g43_n),
    .din1(g41_n_spl_),
    .din2(g42_p_spl_)
  );


  LA
  g_g44_p
  (
    .dout(g44_p),
    .din1(g41_p_spl_),
    .din2(g43_n_spl_)
  );


  FA
  g_g44_n
  (
    .dout(g44_n),
    .din1(g41_n_spl_),
    .din2(g43_p_spl_)
  );


  LA
  g_g45_p
  (
    .dout(g45_p),
    .din1(g42_n_spl_),
    .din2(g43_n_spl_)
  );


  FA
  g_g45_n
  (
    .dout(g45_n),
    .din1(g42_p_spl_),
    .din2(g43_p_spl_)
  );


  LA
  g_g46_p
  (
    .dout(g46_p),
    .din1(g44_n_spl_0),
    .din2(g45_n)
  );


  FA
  g_g46_n
  (
    .dout(g46_n),
    .din1(g44_p_spl_0),
    .din2(g45_p)
  );


  LA
  g_g47_p
  (
    .dout(g47_p),
    .din1(g37_n_spl_0),
    .din2(g46_n_spl_)
  );


  FA
  g_g47_n
  (
    .dout(g47_n),
    .din1(g37_p_spl_),
    .din2(g46_p_spl_)
  );


  LA
  g_g48_p
  (
    .dout(g48_p),
    .din1(g37_p_spl_),
    .din2(g46_p_spl_)
  );


  FA
  g_g48_n
  (
    .dout(g48_n),
    .din1(g37_n_spl_),
    .din2(g46_n_spl_)
  );


  LA
  g_g49_p
  (
    .dout(g49_p),
    .din1(g47_n_spl_),
    .din2(g48_n)
  );


  FA
  g_g49_n
  (
    .dout(g49_n),
    .din1(g47_p_spl_),
    .din2(g48_p)
  );


  LA
  g_g50_p
  (
    .dout(g50_p),
    .din1(g40_n),
    .din2(g49_p)
  );


  FA
  g_g50_n
  (
    .dout(g50_n),
    .din1(g40_p_spl_),
    .din2(g49_n_spl_)
  );


  LA
  g_g51_p
  (
    .dout(g51_p),
    .din1(g40_p_spl_),
    .din2(g49_n_spl_)
  );


  FA
  g_g52_n
  (
    .dout(g52_n),
    .din1(g50_p_spl_),
    .din2(g51_p)
  );


  LA
  g_g53_p
  (
    .dout(g53_p),
    .din1(G1_p_spl_001),
    .din2(G20_p_spl_000)
  );


  FA
  g_g53_n
  (
    .dout(g53_n),
    .din1(G1_n_spl_001),
    .din2(G20_n_spl_000)
  );


  LA
  g_g54_p
  (
    .dout(g54_p),
    .din1(g47_n_spl_),
    .din2(g50_n)
  );


  FA
  g_g54_n
  (
    .dout(g54_n),
    .din1(g47_p_spl_),
    .din2(g50_p_spl_)
  );


  LA
  g_g55_p
  (
    .dout(g55_p),
    .din1(G2_p_spl_001),
    .din2(G19_p_spl_000)
  );


  FA
  g_g55_n
  (
    .dout(g55_n),
    .din1(G2_n_spl_001),
    .din2(G19_n_spl_000)
  );


  LA
  g_g56_p
  (
    .dout(g56_p),
    .din1(G4_p_spl_000),
    .din2(G17_p_spl_001)
  );


  FA
  g_g56_n
  (
    .dout(g56_n),
    .din1(G4_n_spl_000),
    .din2(G17_n_spl_001)
  );


  LA
  g_g57_p
  (
    .dout(g57_p),
    .din1(G3_p_spl_000),
    .din2(G18_p_spl_001)
  );


  FA
  g_g57_n
  (
    .dout(g57_n),
    .din1(G3_n_spl_000),
    .din2(G18_n_spl_001)
  );


  LA
  g_g58_p
  (
    .dout(g58_p),
    .din1(g56_p_spl_),
    .din2(g57_n_spl_)
  );


  FA
  g_g58_n
  (
    .dout(g58_n),
    .din1(g56_n_spl_),
    .din2(g57_p_spl_)
  );


  LA
  g_g59_p
  (
    .dout(g59_p),
    .din1(g56_p_spl_),
    .din2(g58_n_spl_)
  );


  FA
  g_g59_n
  (
    .dout(g59_n),
    .din1(g56_n_spl_),
    .din2(g58_p_spl_)
  );


  LA
  g_g60_p
  (
    .dout(g60_p),
    .din1(g57_n_spl_),
    .din2(g58_n_spl_)
  );


  FA
  g_g60_n
  (
    .dout(g60_n),
    .din1(g57_p_spl_),
    .din2(g58_p_spl_)
  );


  LA
  g_g61_p
  (
    .dout(g61_p),
    .din1(g59_n_spl_0),
    .din2(g60_n)
  );


  FA
  g_g61_n
  (
    .dout(g61_n),
    .din1(g59_p_spl_0),
    .din2(g60_p)
  );


  LA
  g_g62_p
  (
    .dout(g62_p),
    .din1(g44_n_spl_0),
    .din2(g61_n_spl_)
  );


  FA
  g_g62_n
  (
    .dout(g62_n),
    .din1(g44_p_spl_0),
    .din2(g61_p_spl_)
  );


  LA
  g_g63_p
  (
    .dout(g63_p),
    .din1(g44_p_spl_),
    .din2(g61_p_spl_)
  );


  FA
  g_g63_n
  (
    .dout(g63_n),
    .din1(g44_n_spl_),
    .din2(g61_n_spl_)
  );


  LA
  g_g64_p
  (
    .dout(g64_p),
    .din1(g62_n_spl_),
    .din2(g63_n)
  );


  FA
  g_g64_n
  (
    .dout(g64_n),
    .din1(g62_p_spl_),
    .din2(g63_p)
  );


  LA
  g_g65_p
  (
    .dout(g65_p),
    .din1(g55_n_spl_),
    .din2(g64_p_spl_)
  );


  FA
  g_g65_n
  (
    .dout(g65_n),
    .din1(g55_p_spl_),
    .din2(g64_n_spl_)
  );


  LA
  g_g66_p
  (
    .dout(g66_p),
    .din1(g55_p_spl_),
    .din2(g64_n_spl_)
  );


  FA
  g_g66_n
  (
    .dout(g66_n),
    .din1(g55_n_spl_),
    .din2(g64_p_spl_)
  );


  LA
  g_g67_p
  (
    .dout(g67_p),
    .din1(g65_n_spl_),
    .din2(g66_n)
  );


  FA
  g_g67_n
  (
    .dout(g67_n),
    .din1(g65_p_spl_),
    .din2(g66_p)
  );


  LA
  g_g68_p
  (
    .dout(g68_p),
    .din1(g54_n_spl_),
    .din2(g67_p_spl_)
  );


  FA
  g_g68_n
  (
    .dout(g68_n),
    .din1(g54_p_spl_),
    .din2(g67_n_spl_)
  );


  LA
  g_g69_p
  (
    .dout(g69_p),
    .din1(g54_p_spl_),
    .din2(g67_n_spl_)
  );


  FA
  g_g69_n
  (
    .dout(g69_n),
    .din1(g54_n_spl_),
    .din2(g67_p_spl_)
  );


  LA
  g_g70_p
  (
    .dout(g70_p),
    .din1(g68_n_spl_),
    .din2(g69_n)
  );


  FA
  g_g70_n
  (
    .dout(g70_n),
    .din1(g68_p_spl_),
    .din2(g69_p)
  );


  LA
  g_g71_p
  (
    .dout(g71_p),
    .din1(g53_n),
    .din2(g70_p)
  );


  FA
  g_g71_n
  (
    .dout(g71_n),
    .din1(g53_p_spl_),
    .din2(g70_n_spl_)
  );


  LA
  g_g72_p
  (
    .dout(g72_p),
    .din1(g53_p_spl_),
    .din2(g70_n_spl_)
  );


  FA
  g_g73_n
  (
    .dout(g73_n),
    .din1(g71_p_spl_),
    .din2(g72_p)
  );


  LA
  g_g74_p
  (
    .dout(g74_p),
    .din1(G1_p_spl_010),
    .din2(G21_p_spl_000)
  );


  FA
  g_g74_n
  (
    .dout(g74_n),
    .din1(G1_n_spl_001),
    .din2(G21_n_spl_000)
  );


  LA
  g_g75_p
  (
    .dout(g75_p),
    .din1(g68_n_spl_),
    .din2(g71_n)
  );


  FA
  g_g75_n
  (
    .dout(g75_n),
    .din1(g68_p_spl_),
    .din2(g71_p_spl_)
  );


  LA
  g_g76_p
  (
    .dout(g76_p),
    .din1(G2_p_spl_001),
    .din2(G20_p_spl_000)
  );


  FA
  g_g76_n
  (
    .dout(g76_n),
    .din1(G2_n_spl_001),
    .din2(G20_n_spl_000)
  );


  LA
  g_g77_p
  (
    .dout(g77_p),
    .din1(g62_n_spl_),
    .din2(g65_n_spl_)
  );


  FA
  g_g77_n
  (
    .dout(g77_n),
    .din1(g62_p_spl_),
    .din2(g65_p_spl_)
  );


  LA
  g_g78_p
  (
    .dout(g78_p),
    .din1(G3_p_spl_001),
    .din2(G19_p_spl_001)
  );


  FA
  g_g78_n
  (
    .dout(g78_n),
    .din1(G3_n_spl_001),
    .din2(G19_n_spl_001)
  );


  LA
  g_g79_p
  (
    .dout(g79_p),
    .din1(G5_p_spl_000),
    .din2(G17_p_spl_010)
  );


  FA
  g_g79_n
  (
    .dout(g79_n),
    .din1(G5_n_spl_000),
    .din2(G17_n_spl_001)
  );


  LA
  g_g80_p
  (
    .dout(g80_p),
    .din1(G4_p_spl_000),
    .din2(G18_p_spl_001)
  );


  FA
  g_g80_n
  (
    .dout(g80_n),
    .din1(G4_n_spl_000),
    .din2(G18_n_spl_001)
  );


  LA
  g_g81_p
  (
    .dout(g81_p),
    .din1(g79_p_spl_),
    .din2(g80_n_spl_)
  );


  FA
  g_g81_n
  (
    .dout(g81_n),
    .din1(g79_n_spl_),
    .din2(g80_p_spl_)
  );


  LA
  g_g82_p
  (
    .dout(g82_p),
    .din1(g79_p_spl_),
    .din2(g81_n_spl_)
  );


  FA
  g_g82_n
  (
    .dout(g82_n),
    .din1(g79_n_spl_),
    .din2(g81_p_spl_)
  );


  LA
  g_g83_p
  (
    .dout(g83_p),
    .din1(g80_n_spl_),
    .din2(g81_n_spl_)
  );


  FA
  g_g83_n
  (
    .dout(g83_n),
    .din1(g80_p_spl_),
    .din2(g81_p_spl_)
  );


  LA
  g_g84_p
  (
    .dout(g84_p),
    .din1(g82_n_spl_0),
    .din2(g83_n)
  );


  FA
  g_g84_n
  (
    .dout(g84_n),
    .din1(g82_p_spl_0),
    .din2(g83_p)
  );


  LA
  g_g85_p
  (
    .dout(g85_p),
    .din1(g59_n_spl_0),
    .din2(g84_n_spl_)
  );


  FA
  g_g85_n
  (
    .dout(g85_n),
    .din1(g59_p_spl_0),
    .din2(g84_p_spl_)
  );


  LA
  g_g86_p
  (
    .dout(g86_p),
    .din1(g59_p_spl_),
    .din2(g84_p_spl_)
  );


  FA
  g_g86_n
  (
    .dout(g86_n),
    .din1(g59_n_spl_),
    .din2(g84_n_spl_)
  );


  LA
  g_g87_p
  (
    .dout(g87_p),
    .din1(g85_n_spl_),
    .din2(g86_n)
  );


  FA
  g_g87_n
  (
    .dout(g87_n),
    .din1(g85_p_spl_),
    .din2(g86_p)
  );


  LA
  g_g88_p
  (
    .dout(g88_p),
    .din1(g78_n_spl_),
    .din2(g87_p_spl_)
  );


  FA
  g_g88_n
  (
    .dout(g88_n),
    .din1(g78_p_spl_),
    .din2(g87_n_spl_)
  );


  LA
  g_g89_p
  (
    .dout(g89_p),
    .din1(g78_p_spl_),
    .din2(g87_n_spl_)
  );


  FA
  g_g89_n
  (
    .dout(g89_n),
    .din1(g78_n_spl_),
    .din2(g87_p_spl_)
  );


  LA
  g_g90_p
  (
    .dout(g90_p),
    .din1(g88_n_spl_),
    .din2(g89_n)
  );


  FA
  g_g90_n
  (
    .dout(g90_n),
    .din1(g88_p_spl_),
    .din2(g89_p)
  );


  LA
  g_g91_p
  (
    .dout(g91_p),
    .din1(g77_n_spl_),
    .din2(g90_p_spl_)
  );


  FA
  g_g91_n
  (
    .dout(g91_n),
    .din1(g77_p_spl_),
    .din2(g90_n_spl_)
  );


  LA
  g_g92_p
  (
    .dout(g92_p),
    .din1(g77_p_spl_),
    .din2(g90_n_spl_)
  );


  FA
  g_g92_n
  (
    .dout(g92_n),
    .din1(g77_n_spl_),
    .din2(g90_p_spl_)
  );


  LA
  g_g93_p
  (
    .dout(g93_p),
    .din1(g91_n_spl_),
    .din2(g92_n)
  );


  FA
  g_g93_n
  (
    .dout(g93_n),
    .din1(g91_p_spl_),
    .din2(g92_p)
  );


  LA
  g_g94_p
  (
    .dout(g94_p),
    .din1(g76_n_spl_),
    .din2(g93_p_spl_)
  );


  FA
  g_g94_n
  (
    .dout(g94_n),
    .din1(g76_p_spl_),
    .din2(g93_n_spl_)
  );


  LA
  g_g95_p
  (
    .dout(g95_p),
    .din1(g76_p_spl_),
    .din2(g93_n_spl_)
  );


  FA
  g_g95_n
  (
    .dout(g95_n),
    .din1(g76_n_spl_),
    .din2(g93_p_spl_)
  );


  LA
  g_g96_p
  (
    .dout(g96_p),
    .din1(g94_n_spl_),
    .din2(g95_n)
  );


  FA
  g_g96_n
  (
    .dout(g96_n),
    .din1(g94_p_spl_),
    .din2(g95_p)
  );


  LA
  g_g97_p
  (
    .dout(g97_p),
    .din1(g75_n_spl_),
    .din2(g96_p_spl_)
  );


  FA
  g_g97_n
  (
    .dout(g97_n),
    .din1(g75_p_spl_),
    .din2(g96_n_spl_)
  );


  LA
  g_g98_p
  (
    .dout(g98_p),
    .din1(g75_p_spl_),
    .din2(g96_n_spl_)
  );


  FA
  g_g98_n
  (
    .dout(g98_n),
    .din1(g75_n_spl_),
    .din2(g96_p_spl_)
  );


  LA
  g_g99_p
  (
    .dout(g99_p),
    .din1(g97_n_spl_),
    .din2(g98_n)
  );


  FA
  g_g99_n
  (
    .dout(g99_n),
    .din1(g97_p_spl_),
    .din2(g98_p)
  );


  LA
  g_g100_p
  (
    .dout(g100_p),
    .din1(g74_n),
    .din2(g99_p)
  );


  FA
  g_g100_n
  (
    .dout(g100_n),
    .din1(g74_p_spl_),
    .din2(g99_n_spl_)
  );


  LA
  g_g101_p
  (
    .dout(g101_p),
    .din1(g74_p_spl_),
    .din2(g99_n_spl_)
  );


  FA
  g_g102_n
  (
    .dout(g102_n),
    .din1(g100_p_spl_),
    .din2(g101_p)
  );


  LA
  g_g103_p
  (
    .dout(g103_p),
    .din1(G1_p_spl_010),
    .din2(G22_p_spl_000)
  );


  FA
  g_g103_n
  (
    .dout(g103_n),
    .din1(G1_n_spl_010),
    .din2(G22_n_spl_000)
  );


  LA
  g_g104_p
  (
    .dout(g104_p),
    .din1(g97_n_spl_),
    .din2(g100_n)
  );


  FA
  g_g104_n
  (
    .dout(g104_n),
    .din1(g97_p_spl_),
    .din2(g100_p_spl_)
  );


  LA
  g_g105_p
  (
    .dout(g105_p),
    .din1(G2_p_spl_010),
    .din2(G21_p_spl_000)
  );


  FA
  g_g105_n
  (
    .dout(g105_n),
    .din1(G2_n_spl_010),
    .din2(G21_n_spl_000)
  );


  LA
  g_g106_p
  (
    .dout(g106_p),
    .din1(g91_n_spl_),
    .din2(g94_n_spl_)
  );


  FA
  g_g106_n
  (
    .dout(g106_n),
    .din1(g91_p_spl_),
    .din2(g94_p_spl_)
  );


  LA
  g_g107_p
  (
    .dout(g107_p),
    .din1(G3_p_spl_001),
    .din2(G20_p_spl_001)
  );


  FA
  g_g107_n
  (
    .dout(g107_n),
    .din1(G3_n_spl_001),
    .din2(G20_n_spl_001)
  );


  LA
  g_g108_p
  (
    .dout(g108_p),
    .din1(g85_n_spl_),
    .din2(g88_n_spl_)
  );


  FA
  g_g108_n
  (
    .dout(g108_n),
    .din1(g85_p_spl_),
    .din2(g88_p_spl_)
  );


  LA
  g_g109_p
  (
    .dout(g109_p),
    .din1(G4_p_spl_001),
    .din2(G19_p_spl_001)
  );


  FA
  g_g109_n
  (
    .dout(g109_n),
    .din1(G4_n_spl_001),
    .din2(G19_n_spl_001)
  );


  LA
  g_g110_p
  (
    .dout(g110_p),
    .din1(G6_p_spl_000),
    .din2(G17_p_spl_010)
  );


  FA
  g_g110_n
  (
    .dout(g110_n),
    .din1(G6_n_spl_000),
    .din2(G17_n_spl_010)
  );


  LA
  g_g111_p
  (
    .dout(g111_p),
    .din1(G5_p_spl_000),
    .din2(G18_p_spl_010)
  );


  FA
  g_g111_n
  (
    .dout(g111_n),
    .din1(G5_n_spl_000),
    .din2(G18_n_spl_010)
  );


  LA
  g_g112_p
  (
    .dout(g112_p),
    .din1(g110_p_spl_),
    .din2(g111_n_spl_)
  );


  FA
  g_g112_n
  (
    .dout(g112_n),
    .din1(g110_n_spl_),
    .din2(g111_p_spl_)
  );


  LA
  g_g113_p
  (
    .dout(g113_p),
    .din1(g110_p_spl_),
    .din2(g112_n_spl_)
  );


  FA
  g_g113_n
  (
    .dout(g113_n),
    .din1(g110_n_spl_),
    .din2(g112_p_spl_)
  );


  LA
  g_g114_p
  (
    .dout(g114_p),
    .din1(g111_n_spl_),
    .din2(g112_n_spl_)
  );


  FA
  g_g114_n
  (
    .dout(g114_n),
    .din1(g111_p_spl_),
    .din2(g112_p_spl_)
  );


  LA
  g_g115_p
  (
    .dout(g115_p),
    .din1(g113_n_spl_0),
    .din2(g114_n)
  );


  FA
  g_g115_n
  (
    .dout(g115_n),
    .din1(g113_p_spl_0),
    .din2(g114_p)
  );


  LA
  g_g116_p
  (
    .dout(g116_p),
    .din1(g82_n_spl_0),
    .din2(g115_n_spl_)
  );


  FA
  g_g116_n
  (
    .dout(g116_n),
    .din1(g82_p_spl_0),
    .din2(g115_p_spl_)
  );


  LA
  g_g117_p
  (
    .dout(g117_p),
    .din1(g82_p_spl_),
    .din2(g115_p_spl_)
  );


  FA
  g_g117_n
  (
    .dout(g117_n),
    .din1(g82_n_spl_),
    .din2(g115_n_spl_)
  );


  LA
  g_g118_p
  (
    .dout(g118_p),
    .din1(g116_n_spl_),
    .din2(g117_n)
  );


  FA
  g_g118_n
  (
    .dout(g118_n),
    .din1(g116_p_spl_),
    .din2(g117_p)
  );


  LA
  g_g119_p
  (
    .dout(g119_p),
    .din1(g109_n_spl_),
    .din2(g118_p_spl_)
  );


  FA
  g_g119_n
  (
    .dout(g119_n),
    .din1(g109_p_spl_),
    .din2(g118_n_spl_)
  );


  LA
  g_g120_p
  (
    .dout(g120_p),
    .din1(g109_p_spl_),
    .din2(g118_n_spl_)
  );


  FA
  g_g120_n
  (
    .dout(g120_n),
    .din1(g109_n_spl_),
    .din2(g118_p_spl_)
  );


  LA
  g_g121_p
  (
    .dout(g121_p),
    .din1(g119_n_spl_),
    .din2(g120_n)
  );


  FA
  g_g121_n
  (
    .dout(g121_n),
    .din1(g119_p_spl_),
    .din2(g120_p)
  );


  LA
  g_g122_p
  (
    .dout(g122_p),
    .din1(g108_n_spl_),
    .din2(g121_p_spl_)
  );


  FA
  g_g122_n
  (
    .dout(g122_n),
    .din1(g108_p_spl_),
    .din2(g121_n_spl_)
  );


  LA
  g_g123_p
  (
    .dout(g123_p),
    .din1(g108_p_spl_),
    .din2(g121_n_spl_)
  );


  FA
  g_g123_n
  (
    .dout(g123_n),
    .din1(g108_n_spl_),
    .din2(g121_p_spl_)
  );


  LA
  g_g124_p
  (
    .dout(g124_p),
    .din1(g122_n_spl_),
    .din2(g123_n)
  );


  FA
  g_g124_n
  (
    .dout(g124_n),
    .din1(g122_p_spl_),
    .din2(g123_p)
  );


  LA
  g_g125_p
  (
    .dout(g125_p),
    .din1(g107_n_spl_),
    .din2(g124_p_spl_)
  );


  FA
  g_g125_n
  (
    .dout(g125_n),
    .din1(g107_p_spl_),
    .din2(g124_n_spl_)
  );


  LA
  g_g126_p
  (
    .dout(g126_p),
    .din1(g107_p_spl_),
    .din2(g124_n_spl_)
  );


  FA
  g_g126_n
  (
    .dout(g126_n),
    .din1(g107_n_spl_),
    .din2(g124_p_spl_)
  );


  LA
  g_g127_p
  (
    .dout(g127_p),
    .din1(g125_n_spl_),
    .din2(g126_n)
  );


  FA
  g_g127_n
  (
    .dout(g127_n),
    .din1(g125_p_spl_),
    .din2(g126_p)
  );


  LA
  g_g128_p
  (
    .dout(g128_p),
    .din1(g106_n_spl_),
    .din2(g127_p_spl_)
  );


  FA
  g_g128_n
  (
    .dout(g128_n),
    .din1(g106_p_spl_),
    .din2(g127_n_spl_)
  );


  LA
  g_g129_p
  (
    .dout(g129_p),
    .din1(g106_p_spl_),
    .din2(g127_n_spl_)
  );


  FA
  g_g129_n
  (
    .dout(g129_n),
    .din1(g106_n_spl_),
    .din2(g127_p_spl_)
  );


  LA
  g_g130_p
  (
    .dout(g130_p),
    .din1(g128_n_spl_),
    .din2(g129_n)
  );


  FA
  g_g130_n
  (
    .dout(g130_n),
    .din1(g128_p_spl_),
    .din2(g129_p)
  );


  LA
  g_g131_p
  (
    .dout(g131_p),
    .din1(g105_n_spl_),
    .din2(g130_p_spl_)
  );


  FA
  g_g131_n
  (
    .dout(g131_n),
    .din1(g105_p_spl_),
    .din2(g130_n_spl_)
  );


  LA
  g_g132_p
  (
    .dout(g132_p),
    .din1(g105_p_spl_),
    .din2(g130_n_spl_)
  );


  FA
  g_g132_n
  (
    .dout(g132_n),
    .din1(g105_n_spl_),
    .din2(g130_p_spl_)
  );


  LA
  g_g133_p
  (
    .dout(g133_p),
    .din1(g131_n_spl_),
    .din2(g132_n)
  );


  FA
  g_g133_n
  (
    .dout(g133_n),
    .din1(g131_p_spl_),
    .din2(g132_p)
  );


  LA
  g_g134_p
  (
    .dout(g134_p),
    .din1(g104_n_spl_),
    .din2(g133_p_spl_)
  );


  FA
  g_g134_n
  (
    .dout(g134_n),
    .din1(g104_p_spl_),
    .din2(g133_n_spl_)
  );


  LA
  g_g135_p
  (
    .dout(g135_p),
    .din1(g104_p_spl_),
    .din2(g133_n_spl_)
  );


  FA
  g_g135_n
  (
    .dout(g135_n),
    .din1(g104_n_spl_),
    .din2(g133_p_spl_)
  );


  LA
  g_g136_p
  (
    .dout(g136_p),
    .din1(g134_n_spl_),
    .din2(g135_n)
  );


  FA
  g_g136_n
  (
    .dout(g136_n),
    .din1(g134_p_spl_),
    .din2(g135_p)
  );


  LA
  g_g137_p
  (
    .dout(g137_p),
    .din1(g103_n),
    .din2(g136_p)
  );


  FA
  g_g137_n
  (
    .dout(g137_n),
    .din1(g103_p_spl_),
    .din2(g136_n_spl_)
  );


  LA
  g_g138_p
  (
    .dout(g138_p),
    .din1(g103_p_spl_),
    .din2(g136_n_spl_)
  );


  FA
  g_g139_n
  (
    .dout(g139_n),
    .din1(g137_p_spl_),
    .din2(g138_p)
  );


  LA
  g_g140_p
  (
    .dout(g140_p),
    .din1(G1_p_spl_011),
    .din2(G23_p_spl_000)
  );


  FA
  g_g140_n
  (
    .dout(g140_n),
    .din1(G1_n_spl_010),
    .din2(G23_n_spl_000)
  );


  LA
  g_g141_p
  (
    .dout(g141_p),
    .din1(g134_n_spl_),
    .din2(g137_n)
  );


  FA
  g_g141_n
  (
    .dout(g141_n),
    .din1(g134_p_spl_),
    .din2(g137_p_spl_)
  );


  LA
  g_g142_p
  (
    .dout(g142_p),
    .din1(G2_p_spl_010),
    .din2(G22_p_spl_000)
  );


  FA
  g_g142_n
  (
    .dout(g142_n),
    .din1(G2_n_spl_010),
    .din2(G22_n_spl_000)
  );


  LA
  g_g143_p
  (
    .dout(g143_p),
    .din1(g128_n_spl_),
    .din2(g131_n_spl_)
  );


  FA
  g_g143_n
  (
    .dout(g143_n),
    .din1(g128_p_spl_),
    .din2(g131_p_spl_)
  );


  LA
  g_g144_p
  (
    .dout(g144_p),
    .din1(G3_p_spl_010),
    .din2(G21_p_spl_001)
  );


  FA
  g_g144_n
  (
    .dout(g144_n),
    .din1(G3_n_spl_010),
    .din2(G21_n_spl_001)
  );


  LA
  g_g145_p
  (
    .dout(g145_p),
    .din1(g122_n_spl_),
    .din2(g125_n_spl_)
  );


  FA
  g_g145_n
  (
    .dout(g145_n),
    .din1(g122_p_spl_),
    .din2(g125_p_spl_)
  );


  LA
  g_g146_p
  (
    .dout(g146_p),
    .din1(G4_p_spl_001),
    .din2(G20_p_spl_001)
  );


  FA
  g_g146_n
  (
    .dout(g146_n),
    .din1(G4_n_spl_001),
    .din2(G20_n_spl_001)
  );


  LA
  g_g147_p
  (
    .dout(g147_p),
    .din1(g116_n_spl_),
    .din2(g119_n_spl_)
  );


  FA
  g_g147_n
  (
    .dout(g147_n),
    .din1(g116_p_spl_),
    .din2(g119_p_spl_)
  );


  LA
  g_g148_p
  (
    .dout(g148_p),
    .din1(G5_p_spl_001),
    .din2(G19_p_spl_010)
  );


  FA
  g_g148_n
  (
    .dout(g148_n),
    .din1(G5_n_spl_001),
    .din2(G19_n_spl_010)
  );


  LA
  g_g149_p
  (
    .dout(g149_p),
    .din1(G7_p_spl_000),
    .din2(G17_p_spl_011)
  );


  FA
  g_g149_n
  (
    .dout(g149_n),
    .din1(G7_n_spl_000),
    .din2(G17_n_spl_010)
  );


  LA
  g_g150_p
  (
    .dout(g150_p),
    .din1(G6_p_spl_000),
    .din2(G18_p_spl_010)
  );


  FA
  g_g150_n
  (
    .dout(g150_n),
    .din1(G6_n_spl_000),
    .din2(G18_n_spl_010)
  );


  LA
  g_g151_p
  (
    .dout(g151_p),
    .din1(g149_p_spl_),
    .din2(g150_n_spl_)
  );


  FA
  g_g151_n
  (
    .dout(g151_n),
    .din1(g149_n_spl_),
    .din2(g150_p_spl_)
  );


  LA
  g_g152_p
  (
    .dout(g152_p),
    .din1(g149_p_spl_),
    .din2(g151_n_spl_)
  );


  FA
  g_g152_n
  (
    .dout(g152_n),
    .din1(g149_n_spl_),
    .din2(g151_p_spl_)
  );


  LA
  g_g153_p
  (
    .dout(g153_p),
    .din1(g150_n_spl_),
    .din2(g151_n_spl_)
  );


  FA
  g_g153_n
  (
    .dout(g153_n),
    .din1(g150_p_spl_),
    .din2(g151_p_spl_)
  );


  LA
  g_g154_p
  (
    .dout(g154_p),
    .din1(g152_n_spl_0),
    .din2(g153_n)
  );


  FA
  g_g154_n
  (
    .dout(g154_n),
    .din1(g152_p_spl_0),
    .din2(g153_p)
  );


  LA
  g_g155_p
  (
    .dout(g155_p),
    .din1(g113_n_spl_0),
    .din2(g154_n_spl_)
  );


  FA
  g_g155_n
  (
    .dout(g155_n),
    .din1(g113_p_spl_0),
    .din2(g154_p_spl_)
  );


  LA
  g_g156_p
  (
    .dout(g156_p),
    .din1(g113_p_spl_),
    .din2(g154_p_spl_)
  );


  FA
  g_g156_n
  (
    .dout(g156_n),
    .din1(g113_n_spl_),
    .din2(g154_n_spl_)
  );


  LA
  g_g157_p
  (
    .dout(g157_p),
    .din1(g155_n_spl_),
    .din2(g156_n)
  );


  FA
  g_g157_n
  (
    .dout(g157_n),
    .din1(g155_p_spl_),
    .din2(g156_p)
  );


  LA
  g_g158_p
  (
    .dout(g158_p),
    .din1(g148_n_spl_),
    .din2(g157_p_spl_)
  );


  FA
  g_g158_n
  (
    .dout(g158_n),
    .din1(g148_p_spl_),
    .din2(g157_n_spl_)
  );


  LA
  g_g159_p
  (
    .dout(g159_p),
    .din1(g148_p_spl_),
    .din2(g157_n_spl_)
  );


  FA
  g_g159_n
  (
    .dout(g159_n),
    .din1(g148_n_spl_),
    .din2(g157_p_spl_)
  );


  LA
  g_g160_p
  (
    .dout(g160_p),
    .din1(g158_n_spl_),
    .din2(g159_n)
  );


  FA
  g_g160_n
  (
    .dout(g160_n),
    .din1(g158_p_spl_),
    .din2(g159_p)
  );


  LA
  g_g161_p
  (
    .dout(g161_p),
    .din1(g147_n_spl_),
    .din2(g160_p_spl_)
  );


  FA
  g_g161_n
  (
    .dout(g161_n),
    .din1(g147_p_spl_),
    .din2(g160_n_spl_)
  );


  LA
  g_g162_p
  (
    .dout(g162_p),
    .din1(g147_p_spl_),
    .din2(g160_n_spl_)
  );


  FA
  g_g162_n
  (
    .dout(g162_n),
    .din1(g147_n_spl_),
    .din2(g160_p_spl_)
  );


  LA
  g_g163_p
  (
    .dout(g163_p),
    .din1(g161_n_spl_),
    .din2(g162_n)
  );


  FA
  g_g163_n
  (
    .dout(g163_n),
    .din1(g161_p_spl_),
    .din2(g162_p)
  );


  LA
  g_g164_p
  (
    .dout(g164_p),
    .din1(g146_n_spl_),
    .din2(g163_p_spl_)
  );


  FA
  g_g164_n
  (
    .dout(g164_n),
    .din1(g146_p_spl_),
    .din2(g163_n_spl_)
  );


  LA
  g_g165_p
  (
    .dout(g165_p),
    .din1(g146_p_spl_),
    .din2(g163_n_spl_)
  );


  FA
  g_g165_n
  (
    .dout(g165_n),
    .din1(g146_n_spl_),
    .din2(g163_p_spl_)
  );


  LA
  g_g166_p
  (
    .dout(g166_p),
    .din1(g164_n_spl_),
    .din2(g165_n)
  );


  FA
  g_g166_n
  (
    .dout(g166_n),
    .din1(g164_p_spl_),
    .din2(g165_p)
  );


  LA
  g_g167_p
  (
    .dout(g167_p),
    .din1(g145_n_spl_),
    .din2(g166_p_spl_)
  );


  FA
  g_g167_n
  (
    .dout(g167_n),
    .din1(g145_p_spl_),
    .din2(g166_n_spl_)
  );


  LA
  g_g168_p
  (
    .dout(g168_p),
    .din1(g145_p_spl_),
    .din2(g166_n_spl_)
  );


  FA
  g_g168_n
  (
    .dout(g168_n),
    .din1(g145_n_spl_),
    .din2(g166_p_spl_)
  );


  LA
  g_g169_p
  (
    .dout(g169_p),
    .din1(g167_n_spl_),
    .din2(g168_n)
  );


  FA
  g_g169_n
  (
    .dout(g169_n),
    .din1(g167_p_spl_),
    .din2(g168_p)
  );


  LA
  g_g170_p
  (
    .dout(g170_p),
    .din1(g144_n_spl_),
    .din2(g169_p_spl_)
  );


  FA
  g_g170_n
  (
    .dout(g170_n),
    .din1(g144_p_spl_),
    .din2(g169_n_spl_)
  );


  LA
  g_g171_p
  (
    .dout(g171_p),
    .din1(g144_p_spl_),
    .din2(g169_n_spl_)
  );


  FA
  g_g171_n
  (
    .dout(g171_n),
    .din1(g144_n_spl_),
    .din2(g169_p_spl_)
  );


  LA
  g_g172_p
  (
    .dout(g172_p),
    .din1(g170_n_spl_),
    .din2(g171_n)
  );


  FA
  g_g172_n
  (
    .dout(g172_n),
    .din1(g170_p_spl_),
    .din2(g171_p)
  );


  LA
  g_g173_p
  (
    .dout(g173_p),
    .din1(g143_n_spl_),
    .din2(g172_p_spl_)
  );


  FA
  g_g173_n
  (
    .dout(g173_n),
    .din1(g143_p_spl_),
    .din2(g172_n_spl_)
  );


  LA
  g_g174_p
  (
    .dout(g174_p),
    .din1(g143_p_spl_),
    .din2(g172_n_spl_)
  );


  FA
  g_g174_n
  (
    .dout(g174_n),
    .din1(g143_n_spl_),
    .din2(g172_p_spl_)
  );


  LA
  g_g175_p
  (
    .dout(g175_p),
    .din1(g173_n_spl_),
    .din2(g174_n)
  );


  FA
  g_g175_n
  (
    .dout(g175_n),
    .din1(g173_p_spl_),
    .din2(g174_p)
  );


  LA
  g_g176_p
  (
    .dout(g176_p),
    .din1(g142_n_spl_),
    .din2(g175_p_spl_)
  );


  FA
  g_g176_n
  (
    .dout(g176_n),
    .din1(g142_p_spl_),
    .din2(g175_n_spl_)
  );


  LA
  g_g177_p
  (
    .dout(g177_p),
    .din1(g142_p_spl_),
    .din2(g175_n_spl_)
  );


  FA
  g_g177_n
  (
    .dout(g177_n),
    .din1(g142_n_spl_),
    .din2(g175_p_spl_)
  );


  LA
  g_g178_p
  (
    .dout(g178_p),
    .din1(g176_n_spl_),
    .din2(g177_n)
  );


  FA
  g_g178_n
  (
    .dout(g178_n),
    .din1(g176_p_spl_),
    .din2(g177_p)
  );


  LA
  g_g179_p
  (
    .dout(g179_p),
    .din1(g141_n_spl_),
    .din2(g178_p_spl_)
  );


  FA
  g_g179_n
  (
    .dout(g179_n),
    .din1(g141_p_spl_),
    .din2(g178_n_spl_)
  );


  LA
  g_g180_p
  (
    .dout(g180_p),
    .din1(g141_p_spl_),
    .din2(g178_n_spl_)
  );


  FA
  g_g180_n
  (
    .dout(g180_n),
    .din1(g141_n_spl_),
    .din2(g178_p_spl_)
  );


  LA
  g_g181_p
  (
    .dout(g181_p),
    .din1(g179_n_spl_),
    .din2(g180_n)
  );


  FA
  g_g181_n
  (
    .dout(g181_n),
    .din1(g179_p_spl_),
    .din2(g180_p)
  );


  LA
  g_g182_p
  (
    .dout(g182_p),
    .din1(g140_n),
    .din2(g181_p)
  );


  FA
  g_g182_n
  (
    .dout(g182_n),
    .din1(g140_p_spl_),
    .din2(g181_n_spl_)
  );


  LA
  g_g183_p
  (
    .dout(g183_p),
    .din1(g140_p_spl_),
    .din2(g181_n_spl_)
  );


  FA
  g_g184_n
  (
    .dout(g184_n),
    .din1(g182_p_spl_),
    .din2(g183_p)
  );


  LA
  g_g185_p
  (
    .dout(g185_p),
    .din1(G1_p_spl_011),
    .din2(G24_p_spl_000)
  );


  FA
  g_g185_n
  (
    .dout(g185_n),
    .din1(G1_n_spl_011),
    .din2(G24_n_spl_000)
  );


  LA
  g_g186_p
  (
    .dout(g186_p),
    .din1(g179_n_spl_),
    .din2(g182_n)
  );


  FA
  g_g186_n
  (
    .dout(g186_n),
    .din1(g179_p_spl_),
    .din2(g182_p_spl_)
  );


  LA
  g_g187_p
  (
    .dout(g187_p),
    .din1(G2_p_spl_011),
    .din2(G23_p_spl_000)
  );


  FA
  g_g187_n
  (
    .dout(g187_n),
    .din1(G2_n_spl_011),
    .din2(G23_n_spl_000)
  );


  LA
  g_g188_p
  (
    .dout(g188_p),
    .din1(g173_n_spl_),
    .din2(g176_n_spl_)
  );


  FA
  g_g188_n
  (
    .dout(g188_n),
    .din1(g173_p_spl_),
    .din2(g176_p_spl_)
  );


  LA
  g_g189_p
  (
    .dout(g189_p),
    .din1(G3_p_spl_010),
    .din2(G22_p_spl_001)
  );


  FA
  g_g189_n
  (
    .dout(g189_n),
    .din1(G3_n_spl_010),
    .din2(G22_n_spl_001)
  );


  LA
  g_g190_p
  (
    .dout(g190_p),
    .din1(g167_n_spl_),
    .din2(g170_n_spl_)
  );


  FA
  g_g190_n
  (
    .dout(g190_n),
    .din1(g167_p_spl_),
    .din2(g170_p_spl_)
  );


  LA
  g_g191_p
  (
    .dout(g191_p),
    .din1(G4_p_spl_010),
    .din2(G21_p_spl_001)
  );


  FA
  g_g191_n
  (
    .dout(g191_n),
    .din1(G4_n_spl_010),
    .din2(G21_n_spl_001)
  );


  LA
  g_g192_p
  (
    .dout(g192_p),
    .din1(g161_n_spl_),
    .din2(g164_n_spl_)
  );


  FA
  g_g192_n
  (
    .dout(g192_n),
    .din1(g161_p_spl_),
    .din2(g164_p_spl_)
  );


  LA
  g_g193_p
  (
    .dout(g193_p),
    .din1(G5_p_spl_001),
    .din2(G20_p_spl_010)
  );


  FA
  g_g193_n
  (
    .dout(g193_n),
    .din1(G5_n_spl_001),
    .din2(G20_n_spl_010)
  );


  LA
  g_g194_p
  (
    .dout(g194_p),
    .din1(g155_n_spl_),
    .din2(g158_n_spl_)
  );


  FA
  g_g194_n
  (
    .dout(g194_n),
    .din1(g155_p_spl_),
    .din2(g158_p_spl_)
  );


  LA
  g_g195_p
  (
    .dout(g195_p),
    .din1(G6_p_spl_001),
    .din2(G19_p_spl_010)
  );


  FA
  g_g195_n
  (
    .dout(g195_n),
    .din1(G6_n_spl_001),
    .din2(G19_n_spl_010)
  );


  LA
  g_g196_p
  (
    .dout(g196_p),
    .din1(G8_p_spl_000),
    .din2(G17_p_spl_011)
  );


  FA
  g_g196_n
  (
    .dout(g196_n),
    .din1(G8_n_spl_000),
    .din2(G17_n_spl_011)
  );


  LA
  g_g197_p
  (
    .dout(g197_p),
    .din1(G7_p_spl_000),
    .din2(G18_p_spl_011)
  );


  FA
  g_g197_n
  (
    .dout(g197_n),
    .din1(G7_n_spl_000),
    .din2(G18_n_spl_011)
  );


  LA
  g_g198_p
  (
    .dout(g198_p),
    .din1(g196_p_spl_),
    .din2(g197_n_spl_)
  );


  FA
  g_g198_n
  (
    .dout(g198_n),
    .din1(g196_n_spl_),
    .din2(g197_p_spl_)
  );


  LA
  g_g199_p
  (
    .dout(g199_p),
    .din1(g196_p_spl_),
    .din2(g198_n_spl_)
  );


  FA
  g_g199_n
  (
    .dout(g199_n),
    .din1(g196_n_spl_),
    .din2(g198_p_spl_)
  );


  LA
  g_g200_p
  (
    .dout(g200_p),
    .din1(g197_n_spl_),
    .din2(g198_n_spl_)
  );


  FA
  g_g200_n
  (
    .dout(g200_n),
    .din1(g197_p_spl_),
    .din2(g198_p_spl_)
  );


  LA
  g_g201_p
  (
    .dout(g201_p),
    .din1(g199_n_spl_0),
    .din2(g200_n)
  );


  FA
  g_g201_n
  (
    .dout(g201_n),
    .din1(g199_p_spl_0),
    .din2(g200_p)
  );


  LA
  g_g202_p
  (
    .dout(g202_p),
    .din1(g152_n_spl_0),
    .din2(g201_n_spl_)
  );


  FA
  g_g202_n
  (
    .dout(g202_n),
    .din1(g152_p_spl_0),
    .din2(g201_p_spl_)
  );


  LA
  g_g203_p
  (
    .dout(g203_p),
    .din1(g152_p_spl_),
    .din2(g201_p_spl_)
  );


  FA
  g_g203_n
  (
    .dout(g203_n),
    .din1(g152_n_spl_),
    .din2(g201_n_spl_)
  );


  LA
  g_g204_p
  (
    .dout(g204_p),
    .din1(g202_n_spl_),
    .din2(g203_n)
  );


  FA
  g_g204_n
  (
    .dout(g204_n),
    .din1(g202_p_spl_),
    .din2(g203_p)
  );


  LA
  g_g205_p
  (
    .dout(g205_p),
    .din1(g195_n_spl_),
    .din2(g204_p_spl_)
  );


  FA
  g_g205_n
  (
    .dout(g205_n),
    .din1(g195_p_spl_),
    .din2(g204_n_spl_)
  );


  LA
  g_g206_p
  (
    .dout(g206_p),
    .din1(g195_p_spl_),
    .din2(g204_n_spl_)
  );


  FA
  g_g206_n
  (
    .dout(g206_n),
    .din1(g195_n_spl_),
    .din2(g204_p_spl_)
  );


  LA
  g_g207_p
  (
    .dout(g207_p),
    .din1(g205_n_spl_),
    .din2(g206_n)
  );


  FA
  g_g207_n
  (
    .dout(g207_n),
    .din1(g205_p_spl_),
    .din2(g206_p)
  );


  LA
  g_g208_p
  (
    .dout(g208_p),
    .din1(g194_n_spl_),
    .din2(g207_p_spl_)
  );


  FA
  g_g208_n
  (
    .dout(g208_n),
    .din1(g194_p_spl_),
    .din2(g207_n_spl_)
  );


  LA
  g_g209_p
  (
    .dout(g209_p),
    .din1(g194_p_spl_),
    .din2(g207_n_spl_)
  );


  FA
  g_g209_n
  (
    .dout(g209_n),
    .din1(g194_n_spl_),
    .din2(g207_p_spl_)
  );


  LA
  g_g210_p
  (
    .dout(g210_p),
    .din1(g208_n_spl_),
    .din2(g209_n)
  );


  FA
  g_g210_n
  (
    .dout(g210_n),
    .din1(g208_p_spl_),
    .din2(g209_p)
  );


  LA
  g_g211_p
  (
    .dout(g211_p),
    .din1(g193_n_spl_),
    .din2(g210_p_spl_)
  );


  FA
  g_g211_n
  (
    .dout(g211_n),
    .din1(g193_p_spl_),
    .din2(g210_n_spl_)
  );


  LA
  g_g212_p
  (
    .dout(g212_p),
    .din1(g193_p_spl_),
    .din2(g210_n_spl_)
  );


  FA
  g_g212_n
  (
    .dout(g212_n),
    .din1(g193_n_spl_),
    .din2(g210_p_spl_)
  );


  LA
  g_g213_p
  (
    .dout(g213_p),
    .din1(g211_n_spl_),
    .din2(g212_n)
  );


  FA
  g_g213_n
  (
    .dout(g213_n),
    .din1(g211_p_spl_),
    .din2(g212_p)
  );


  LA
  g_g214_p
  (
    .dout(g214_p),
    .din1(g192_n_spl_),
    .din2(g213_p_spl_)
  );


  FA
  g_g214_n
  (
    .dout(g214_n),
    .din1(g192_p_spl_),
    .din2(g213_n_spl_)
  );


  LA
  g_g215_p
  (
    .dout(g215_p),
    .din1(g192_p_spl_),
    .din2(g213_n_spl_)
  );


  FA
  g_g215_n
  (
    .dout(g215_n),
    .din1(g192_n_spl_),
    .din2(g213_p_spl_)
  );


  LA
  g_g216_p
  (
    .dout(g216_p),
    .din1(g214_n_spl_),
    .din2(g215_n)
  );


  FA
  g_g216_n
  (
    .dout(g216_n),
    .din1(g214_p_spl_),
    .din2(g215_p)
  );


  LA
  g_g217_p
  (
    .dout(g217_p),
    .din1(g191_n_spl_),
    .din2(g216_p_spl_)
  );


  FA
  g_g217_n
  (
    .dout(g217_n),
    .din1(g191_p_spl_),
    .din2(g216_n_spl_)
  );


  LA
  g_g218_p
  (
    .dout(g218_p),
    .din1(g191_p_spl_),
    .din2(g216_n_spl_)
  );


  FA
  g_g218_n
  (
    .dout(g218_n),
    .din1(g191_n_spl_),
    .din2(g216_p_spl_)
  );


  LA
  g_g219_p
  (
    .dout(g219_p),
    .din1(g217_n_spl_),
    .din2(g218_n)
  );


  FA
  g_g219_n
  (
    .dout(g219_n),
    .din1(g217_p_spl_),
    .din2(g218_p)
  );


  LA
  g_g220_p
  (
    .dout(g220_p),
    .din1(g190_n_spl_),
    .din2(g219_p_spl_)
  );


  FA
  g_g220_n
  (
    .dout(g220_n),
    .din1(g190_p_spl_),
    .din2(g219_n_spl_)
  );


  LA
  g_g221_p
  (
    .dout(g221_p),
    .din1(g190_p_spl_),
    .din2(g219_n_spl_)
  );


  FA
  g_g221_n
  (
    .dout(g221_n),
    .din1(g190_n_spl_),
    .din2(g219_p_spl_)
  );


  LA
  g_g222_p
  (
    .dout(g222_p),
    .din1(g220_n_spl_),
    .din2(g221_n)
  );


  FA
  g_g222_n
  (
    .dout(g222_n),
    .din1(g220_p_spl_),
    .din2(g221_p)
  );


  LA
  g_g223_p
  (
    .dout(g223_p),
    .din1(g189_n_spl_),
    .din2(g222_p_spl_)
  );


  FA
  g_g223_n
  (
    .dout(g223_n),
    .din1(g189_p_spl_),
    .din2(g222_n_spl_)
  );


  LA
  g_g224_p
  (
    .dout(g224_p),
    .din1(g189_p_spl_),
    .din2(g222_n_spl_)
  );


  FA
  g_g224_n
  (
    .dout(g224_n),
    .din1(g189_n_spl_),
    .din2(g222_p_spl_)
  );


  LA
  g_g225_p
  (
    .dout(g225_p),
    .din1(g223_n_spl_),
    .din2(g224_n)
  );


  FA
  g_g225_n
  (
    .dout(g225_n),
    .din1(g223_p_spl_),
    .din2(g224_p)
  );


  LA
  g_g226_p
  (
    .dout(g226_p),
    .din1(g188_n_spl_),
    .din2(g225_p_spl_)
  );


  FA
  g_g226_n
  (
    .dout(g226_n),
    .din1(g188_p_spl_),
    .din2(g225_n_spl_)
  );


  LA
  g_g227_p
  (
    .dout(g227_p),
    .din1(g188_p_spl_),
    .din2(g225_n_spl_)
  );


  FA
  g_g227_n
  (
    .dout(g227_n),
    .din1(g188_n_spl_),
    .din2(g225_p_spl_)
  );


  LA
  g_g228_p
  (
    .dout(g228_p),
    .din1(g226_n_spl_),
    .din2(g227_n)
  );


  FA
  g_g228_n
  (
    .dout(g228_n),
    .din1(g226_p_spl_),
    .din2(g227_p)
  );


  LA
  g_g229_p
  (
    .dout(g229_p),
    .din1(g187_n_spl_),
    .din2(g228_p_spl_)
  );


  FA
  g_g229_n
  (
    .dout(g229_n),
    .din1(g187_p_spl_),
    .din2(g228_n_spl_)
  );


  LA
  g_g230_p
  (
    .dout(g230_p),
    .din1(g187_p_spl_),
    .din2(g228_n_spl_)
  );


  FA
  g_g230_n
  (
    .dout(g230_n),
    .din1(g187_n_spl_),
    .din2(g228_p_spl_)
  );


  LA
  g_g231_p
  (
    .dout(g231_p),
    .din1(g229_n_spl_),
    .din2(g230_n)
  );


  FA
  g_g231_n
  (
    .dout(g231_n),
    .din1(g229_p_spl_),
    .din2(g230_p)
  );


  LA
  g_g232_p
  (
    .dout(g232_p),
    .din1(g186_n_spl_),
    .din2(g231_p_spl_)
  );


  FA
  g_g232_n
  (
    .dout(g232_n),
    .din1(g186_p_spl_),
    .din2(g231_n_spl_)
  );


  LA
  g_g233_p
  (
    .dout(g233_p),
    .din1(g186_p_spl_),
    .din2(g231_n_spl_)
  );


  FA
  g_g233_n
  (
    .dout(g233_n),
    .din1(g186_n_spl_),
    .din2(g231_p_spl_)
  );


  LA
  g_g234_p
  (
    .dout(g234_p),
    .din1(g232_n_spl_),
    .din2(g233_n)
  );


  FA
  g_g234_n
  (
    .dout(g234_n),
    .din1(g232_p_spl_),
    .din2(g233_p)
  );


  LA
  g_g235_p
  (
    .dout(g235_p),
    .din1(g185_n),
    .din2(g234_p)
  );


  FA
  g_g235_n
  (
    .dout(g235_n),
    .din1(g185_p_spl_),
    .din2(g234_n_spl_)
  );


  LA
  g_g236_p
  (
    .dout(g236_p),
    .din1(g185_p_spl_),
    .din2(g234_n_spl_)
  );


  FA
  g_g237_n
  (
    .dout(g237_n),
    .din1(g235_p_spl_),
    .din2(g236_p)
  );


  LA
  g_g238_p
  (
    .dout(g238_p),
    .din1(G1_p_spl_100),
    .din2(G25_p_spl_000)
  );


  FA
  g_g238_n
  (
    .dout(g238_n),
    .din1(G1_n_spl_011),
    .din2(G25_n_spl_000)
  );


  LA
  g_g239_p
  (
    .dout(g239_p),
    .din1(g232_n_spl_),
    .din2(g235_n)
  );


  FA
  g_g239_n
  (
    .dout(g239_n),
    .din1(g232_p_spl_),
    .din2(g235_p_spl_)
  );


  LA
  g_g240_p
  (
    .dout(g240_p),
    .din1(G2_p_spl_011),
    .din2(G24_p_spl_000)
  );


  FA
  g_g240_n
  (
    .dout(g240_n),
    .din1(G2_n_spl_011),
    .din2(G24_n_spl_000)
  );


  LA
  g_g241_p
  (
    .dout(g241_p),
    .din1(g226_n_spl_),
    .din2(g229_n_spl_)
  );


  FA
  g_g241_n
  (
    .dout(g241_n),
    .din1(g226_p_spl_),
    .din2(g229_p_spl_)
  );


  LA
  g_g242_p
  (
    .dout(g242_p),
    .din1(G3_p_spl_011),
    .din2(G23_p_spl_001)
  );


  FA
  g_g242_n
  (
    .dout(g242_n),
    .din1(G3_n_spl_011),
    .din2(G23_n_spl_001)
  );


  LA
  g_g243_p
  (
    .dout(g243_p),
    .din1(g220_n_spl_),
    .din2(g223_n_spl_)
  );


  FA
  g_g243_n
  (
    .dout(g243_n),
    .din1(g220_p_spl_),
    .din2(g223_p_spl_)
  );


  LA
  g_g244_p
  (
    .dout(g244_p),
    .din1(G4_p_spl_010),
    .din2(G22_p_spl_001)
  );


  FA
  g_g244_n
  (
    .dout(g244_n),
    .din1(G4_n_spl_010),
    .din2(G22_n_spl_001)
  );


  LA
  g_g245_p
  (
    .dout(g245_p),
    .din1(g214_n_spl_),
    .din2(g217_n_spl_)
  );


  FA
  g_g245_n
  (
    .dout(g245_n),
    .din1(g214_p_spl_),
    .din2(g217_p_spl_)
  );


  LA
  g_g246_p
  (
    .dout(g246_p),
    .din1(G5_p_spl_010),
    .din2(G21_p_spl_010)
  );


  FA
  g_g246_n
  (
    .dout(g246_n),
    .din1(G5_n_spl_010),
    .din2(G21_n_spl_010)
  );


  LA
  g_g247_p
  (
    .dout(g247_p),
    .din1(g208_n_spl_),
    .din2(g211_n_spl_)
  );


  FA
  g_g247_n
  (
    .dout(g247_n),
    .din1(g208_p_spl_),
    .din2(g211_p_spl_)
  );


  LA
  g_g248_p
  (
    .dout(g248_p),
    .din1(G6_p_spl_001),
    .din2(G20_p_spl_010)
  );


  FA
  g_g248_n
  (
    .dout(g248_n),
    .din1(G6_n_spl_001),
    .din2(G20_n_spl_010)
  );


  LA
  g_g249_p
  (
    .dout(g249_p),
    .din1(g202_n_spl_),
    .din2(g205_n_spl_)
  );


  FA
  g_g249_n
  (
    .dout(g249_n),
    .din1(g202_p_spl_),
    .din2(g205_p_spl_)
  );


  LA
  g_g250_p
  (
    .dout(g250_p),
    .din1(G7_p_spl_001),
    .din2(G19_p_spl_011)
  );


  FA
  g_g250_n
  (
    .dout(g250_n),
    .din1(G7_n_spl_001),
    .din2(G19_n_spl_011)
  );


  LA
  g_g251_p
  (
    .dout(g251_p),
    .din1(G9_p_spl_000),
    .din2(G17_p_spl_100)
  );


  FA
  g_g251_n
  (
    .dout(g251_n),
    .din1(G9_n_spl_000),
    .din2(G17_n_spl_011)
  );


  LA
  g_g252_p
  (
    .dout(g252_p),
    .din1(G8_p_spl_000),
    .din2(G18_p_spl_011)
  );


  FA
  g_g252_n
  (
    .dout(g252_n),
    .din1(G8_n_spl_000),
    .din2(G18_n_spl_011)
  );


  LA
  g_g253_p
  (
    .dout(g253_p),
    .din1(g251_p_spl_),
    .din2(g252_n_spl_)
  );


  FA
  g_g253_n
  (
    .dout(g253_n),
    .din1(g251_n_spl_),
    .din2(g252_p_spl_)
  );


  LA
  g_g254_p
  (
    .dout(g254_p),
    .din1(g251_p_spl_),
    .din2(g253_n_spl_)
  );


  FA
  g_g254_n
  (
    .dout(g254_n),
    .din1(g251_n_spl_),
    .din2(g253_p_spl_)
  );


  LA
  g_g255_p
  (
    .dout(g255_p),
    .din1(g252_n_spl_),
    .din2(g253_n_spl_)
  );


  FA
  g_g255_n
  (
    .dout(g255_n),
    .din1(g252_p_spl_),
    .din2(g253_p_spl_)
  );


  LA
  g_g256_p
  (
    .dout(g256_p),
    .din1(g254_n_spl_0),
    .din2(g255_n)
  );


  FA
  g_g256_n
  (
    .dout(g256_n),
    .din1(g254_p_spl_0),
    .din2(g255_p)
  );


  LA
  g_g257_p
  (
    .dout(g257_p),
    .din1(g199_n_spl_0),
    .din2(g256_n_spl_)
  );


  FA
  g_g257_n
  (
    .dout(g257_n),
    .din1(g199_p_spl_0),
    .din2(g256_p_spl_)
  );


  LA
  g_g258_p
  (
    .dout(g258_p),
    .din1(g199_p_spl_),
    .din2(g256_p_spl_)
  );


  FA
  g_g258_n
  (
    .dout(g258_n),
    .din1(g199_n_spl_),
    .din2(g256_n_spl_)
  );


  LA
  g_g259_p
  (
    .dout(g259_p),
    .din1(g257_n_spl_),
    .din2(g258_n)
  );


  FA
  g_g259_n
  (
    .dout(g259_n),
    .din1(g257_p_spl_),
    .din2(g258_p)
  );


  LA
  g_g260_p
  (
    .dout(g260_p),
    .din1(g250_n_spl_),
    .din2(g259_p_spl_)
  );


  FA
  g_g260_n
  (
    .dout(g260_n),
    .din1(g250_p_spl_),
    .din2(g259_n_spl_)
  );


  LA
  g_g261_p
  (
    .dout(g261_p),
    .din1(g250_p_spl_),
    .din2(g259_n_spl_)
  );


  FA
  g_g261_n
  (
    .dout(g261_n),
    .din1(g250_n_spl_),
    .din2(g259_p_spl_)
  );


  LA
  g_g262_p
  (
    .dout(g262_p),
    .din1(g260_n_spl_),
    .din2(g261_n)
  );


  FA
  g_g262_n
  (
    .dout(g262_n),
    .din1(g260_p_spl_),
    .din2(g261_p)
  );


  LA
  g_g263_p
  (
    .dout(g263_p),
    .din1(g249_n_spl_),
    .din2(g262_p_spl_)
  );


  FA
  g_g263_n
  (
    .dout(g263_n),
    .din1(g249_p_spl_),
    .din2(g262_n_spl_)
  );


  LA
  g_g264_p
  (
    .dout(g264_p),
    .din1(g249_p_spl_),
    .din2(g262_n_spl_)
  );


  FA
  g_g264_n
  (
    .dout(g264_n),
    .din1(g249_n_spl_),
    .din2(g262_p_spl_)
  );


  LA
  g_g265_p
  (
    .dout(g265_p),
    .din1(g263_n_spl_),
    .din2(g264_n)
  );


  FA
  g_g265_n
  (
    .dout(g265_n),
    .din1(g263_p_spl_),
    .din2(g264_p)
  );


  LA
  g_g266_p
  (
    .dout(g266_p),
    .din1(g248_n_spl_),
    .din2(g265_p_spl_)
  );


  FA
  g_g266_n
  (
    .dout(g266_n),
    .din1(g248_p_spl_),
    .din2(g265_n_spl_)
  );


  LA
  g_g267_p
  (
    .dout(g267_p),
    .din1(g248_p_spl_),
    .din2(g265_n_spl_)
  );


  FA
  g_g267_n
  (
    .dout(g267_n),
    .din1(g248_n_spl_),
    .din2(g265_p_spl_)
  );


  LA
  g_g268_p
  (
    .dout(g268_p),
    .din1(g266_n_spl_),
    .din2(g267_n)
  );


  FA
  g_g268_n
  (
    .dout(g268_n),
    .din1(g266_p_spl_),
    .din2(g267_p)
  );


  LA
  g_g269_p
  (
    .dout(g269_p),
    .din1(g247_n_spl_),
    .din2(g268_p_spl_)
  );


  FA
  g_g269_n
  (
    .dout(g269_n),
    .din1(g247_p_spl_),
    .din2(g268_n_spl_)
  );


  LA
  g_g270_p
  (
    .dout(g270_p),
    .din1(g247_p_spl_),
    .din2(g268_n_spl_)
  );


  FA
  g_g270_n
  (
    .dout(g270_n),
    .din1(g247_n_spl_),
    .din2(g268_p_spl_)
  );


  LA
  g_g271_p
  (
    .dout(g271_p),
    .din1(g269_n_spl_),
    .din2(g270_n)
  );


  FA
  g_g271_n
  (
    .dout(g271_n),
    .din1(g269_p_spl_),
    .din2(g270_p)
  );


  LA
  g_g272_p
  (
    .dout(g272_p),
    .din1(g246_n_spl_),
    .din2(g271_p_spl_)
  );


  FA
  g_g272_n
  (
    .dout(g272_n),
    .din1(g246_p_spl_),
    .din2(g271_n_spl_)
  );


  LA
  g_g273_p
  (
    .dout(g273_p),
    .din1(g246_p_spl_),
    .din2(g271_n_spl_)
  );


  FA
  g_g273_n
  (
    .dout(g273_n),
    .din1(g246_n_spl_),
    .din2(g271_p_spl_)
  );


  LA
  g_g274_p
  (
    .dout(g274_p),
    .din1(g272_n_spl_),
    .din2(g273_n)
  );


  FA
  g_g274_n
  (
    .dout(g274_n),
    .din1(g272_p_spl_),
    .din2(g273_p)
  );


  LA
  g_g275_p
  (
    .dout(g275_p),
    .din1(g245_n_spl_),
    .din2(g274_p_spl_)
  );


  FA
  g_g275_n
  (
    .dout(g275_n),
    .din1(g245_p_spl_),
    .din2(g274_n_spl_)
  );


  LA
  g_g276_p
  (
    .dout(g276_p),
    .din1(g245_p_spl_),
    .din2(g274_n_spl_)
  );


  FA
  g_g276_n
  (
    .dout(g276_n),
    .din1(g245_n_spl_),
    .din2(g274_p_spl_)
  );


  LA
  g_g277_p
  (
    .dout(g277_p),
    .din1(g275_n_spl_),
    .din2(g276_n)
  );


  FA
  g_g277_n
  (
    .dout(g277_n),
    .din1(g275_p_spl_),
    .din2(g276_p)
  );


  LA
  g_g278_p
  (
    .dout(g278_p),
    .din1(g244_n_spl_),
    .din2(g277_p_spl_)
  );


  FA
  g_g278_n
  (
    .dout(g278_n),
    .din1(g244_p_spl_),
    .din2(g277_n_spl_)
  );


  LA
  g_g279_p
  (
    .dout(g279_p),
    .din1(g244_p_spl_),
    .din2(g277_n_spl_)
  );


  FA
  g_g279_n
  (
    .dout(g279_n),
    .din1(g244_n_spl_),
    .din2(g277_p_spl_)
  );


  LA
  g_g280_p
  (
    .dout(g280_p),
    .din1(g278_n_spl_),
    .din2(g279_n)
  );


  FA
  g_g280_n
  (
    .dout(g280_n),
    .din1(g278_p_spl_),
    .din2(g279_p)
  );


  LA
  g_g281_p
  (
    .dout(g281_p),
    .din1(g243_n_spl_),
    .din2(g280_p_spl_)
  );


  FA
  g_g281_n
  (
    .dout(g281_n),
    .din1(g243_p_spl_),
    .din2(g280_n_spl_)
  );


  LA
  g_g282_p
  (
    .dout(g282_p),
    .din1(g243_p_spl_),
    .din2(g280_n_spl_)
  );


  FA
  g_g282_n
  (
    .dout(g282_n),
    .din1(g243_n_spl_),
    .din2(g280_p_spl_)
  );


  LA
  g_g283_p
  (
    .dout(g283_p),
    .din1(g281_n_spl_),
    .din2(g282_n)
  );


  FA
  g_g283_n
  (
    .dout(g283_n),
    .din1(g281_p_spl_),
    .din2(g282_p)
  );


  LA
  g_g284_p
  (
    .dout(g284_p),
    .din1(g242_n_spl_),
    .din2(g283_p_spl_)
  );


  FA
  g_g284_n
  (
    .dout(g284_n),
    .din1(g242_p_spl_),
    .din2(g283_n_spl_)
  );


  LA
  g_g285_p
  (
    .dout(g285_p),
    .din1(g242_p_spl_),
    .din2(g283_n_spl_)
  );


  FA
  g_g285_n
  (
    .dout(g285_n),
    .din1(g242_n_spl_),
    .din2(g283_p_spl_)
  );


  LA
  g_g286_p
  (
    .dout(g286_p),
    .din1(g284_n_spl_),
    .din2(g285_n)
  );


  FA
  g_g286_n
  (
    .dout(g286_n),
    .din1(g284_p_spl_),
    .din2(g285_p)
  );


  LA
  g_g287_p
  (
    .dout(g287_p),
    .din1(g241_n_spl_),
    .din2(g286_p_spl_)
  );


  FA
  g_g287_n
  (
    .dout(g287_n),
    .din1(g241_p_spl_),
    .din2(g286_n_spl_)
  );


  LA
  g_g288_p
  (
    .dout(g288_p),
    .din1(g241_p_spl_),
    .din2(g286_n_spl_)
  );


  FA
  g_g288_n
  (
    .dout(g288_n),
    .din1(g241_n_spl_),
    .din2(g286_p_spl_)
  );


  LA
  g_g289_p
  (
    .dout(g289_p),
    .din1(g287_n_spl_),
    .din2(g288_n)
  );


  FA
  g_g289_n
  (
    .dout(g289_n),
    .din1(g287_p_spl_),
    .din2(g288_p)
  );


  LA
  g_g290_p
  (
    .dout(g290_p),
    .din1(g240_n_spl_),
    .din2(g289_p_spl_)
  );


  FA
  g_g290_n
  (
    .dout(g290_n),
    .din1(g240_p_spl_),
    .din2(g289_n_spl_)
  );


  LA
  g_g291_p
  (
    .dout(g291_p),
    .din1(g240_p_spl_),
    .din2(g289_n_spl_)
  );


  FA
  g_g291_n
  (
    .dout(g291_n),
    .din1(g240_n_spl_),
    .din2(g289_p_spl_)
  );


  LA
  g_g292_p
  (
    .dout(g292_p),
    .din1(g290_n_spl_),
    .din2(g291_n)
  );


  FA
  g_g292_n
  (
    .dout(g292_n),
    .din1(g290_p_spl_),
    .din2(g291_p)
  );


  LA
  g_g293_p
  (
    .dout(g293_p),
    .din1(g239_n_spl_),
    .din2(g292_p_spl_)
  );


  FA
  g_g293_n
  (
    .dout(g293_n),
    .din1(g239_p_spl_),
    .din2(g292_n_spl_)
  );


  LA
  g_g294_p
  (
    .dout(g294_p),
    .din1(g239_p_spl_),
    .din2(g292_n_spl_)
  );


  FA
  g_g294_n
  (
    .dout(g294_n),
    .din1(g239_n_spl_),
    .din2(g292_p_spl_)
  );


  LA
  g_g295_p
  (
    .dout(g295_p),
    .din1(g293_n_spl_),
    .din2(g294_n)
  );


  FA
  g_g295_n
  (
    .dout(g295_n),
    .din1(g293_p_spl_),
    .din2(g294_p)
  );


  LA
  g_g296_p
  (
    .dout(g296_p),
    .din1(g238_n),
    .din2(g295_p)
  );


  FA
  g_g296_n
  (
    .dout(g296_n),
    .din1(g238_p_spl_),
    .din2(g295_n_spl_)
  );


  LA
  g_g297_p
  (
    .dout(g297_p),
    .din1(g238_p_spl_),
    .din2(g295_n_spl_)
  );


  FA
  g_g298_n
  (
    .dout(g298_n),
    .din1(g296_p_spl_),
    .din2(g297_p)
  );


  LA
  g_g299_p
  (
    .dout(g299_p),
    .din1(G1_p_spl_100),
    .din2(G26_p_spl_000)
  );


  FA
  g_g299_n
  (
    .dout(g299_n),
    .din1(G1_n_spl_100),
    .din2(G26_n_spl_000)
  );


  LA
  g_g300_p
  (
    .dout(g300_p),
    .din1(g293_n_spl_),
    .din2(g296_n)
  );


  FA
  g_g300_n
  (
    .dout(g300_n),
    .din1(g293_p_spl_),
    .din2(g296_p_spl_)
  );


  LA
  g_g301_p
  (
    .dout(g301_p),
    .din1(G2_p_spl_100),
    .din2(G25_p_spl_000)
  );


  FA
  g_g301_n
  (
    .dout(g301_n),
    .din1(G2_n_spl_100),
    .din2(G25_n_spl_000)
  );


  LA
  g_g302_p
  (
    .dout(g302_p),
    .din1(g287_n_spl_),
    .din2(g290_n_spl_)
  );


  FA
  g_g302_n
  (
    .dout(g302_n),
    .din1(g287_p_spl_),
    .din2(g290_p_spl_)
  );


  LA
  g_g303_p
  (
    .dout(g303_p),
    .din1(G3_p_spl_011),
    .din2(G24_p_spl_001)
  );


  FA
  g_g303_n
  (
    .dout(g303_n),
    .din1(G3_n_spl_011),
    .din2(G24_n_spl_001)
  );


  LA
  g_g304_p
  (
    .dout(g304_p),
    .din1(g281_n_spl_),
    .din2(g284_n_spl_)
  );


  FA
  g_g304_n
  (
    .dout(g304_n),
    .din1(g281_p_spl_),
    .din2(g284_p_spl_)
  );


  LA
  g_g305_p
  (
    .dout(g305_p),
    .din1(G4_p_spl_011),
    .din2(G23_p_spl_001)
  );


  FA
  g_g305_n
  (
    .dout(g305_n),
    .din1(G4_n_spl_011),
    .din2(G23_n_spl_001)
  );


  LA
  g_g306_p
  (
    .dout(g306_p),
    .din1(g275_n_spl_),
    .din2(g278_n_spl_)
  );


  FA
  g_g306_n
  (
    .dout(g306_n),
    .din1(g275_p_spl_),
    .din2(g278_p_spl_)
  );


  LA
  g_g307_p
  (
    .dout(g307_p),
    .din1(G5_p_spl_010),
    .din2(G22_p_spl_010)
  );


  FA
  g_g307_n
  (
    .dout(g307_n),
    .din1(G5_n_spl_010),
    .din2(G22_n_spl_010)
  );


  LA
  g_g308_p
  (
    .dout(g308_p),
    .din1(g269_n_spl_),
    .din2(g272_n_spl_)
  );


  FA
  g_g308_n
  (
    .dout(g308_n),
    .din1(g269_p_spl_),
    .din2(g272_p_spl_)
  );


  LA
  g_g309_p
  (
    .dout(g309_p),
    .din1(G6_p_spl_010),
    .din2(G21_p_spl_010)
  );


  FA
  g_g309_n
  (
    .dout(g309_n),
    .din1(G6_n_spl_010),
    .din2(G21_n_spl_010)
  );


  LA
  g_g310_p
  (
    .dout(g310_p),
    .din1(g263_n_spl_),
    .din2(g266_n_spl_)
  );


  FA
  g_g310_n
  (
    .dout(g310_n),
    .din1(g263_p_spl_),
    .din2(g266_p_spl_)
  );


  LA
  g_g311_p
  (
    .dout(g311_p),
    .din1(G7_p_spl_001),
    .din2(G20_p_spl_011)
  );


  FA
  g_g311_n
  (
    .dout(g311_n),
    .din1(G7_n_spl_001),
    .din2(G20_n_spl_011)
  );


  LA
  g_g312_p
  (
    .dout(g312_p),
    .din1(g257_n_spl_),
    .din2(g260_n_spl_)
  );


  FA
  g_g312_n
  (
    .dout(g312_n),
    .din1(g257_p_spl_),
    .din2(g260_p_spl_)
  );


  LA
  g_g313_p
  (
    .dout(g313_p),
    .din1(G8_p_spl_001),
    .din2(G19_p_spl_011)
  );


  FA
  g_g313_n
  (
    .dout(g313_n),
    .din1(G8_n_spl_001),
    .din2(G19_n_spl_011)
  );


  LA
  g_g314_p
  (
    .dout(g314_p),
    .din1(G10_p_spl_000),
    .din2(G17_p_spl_100)
  );


  FA
  g_g314_n
  (
    .dout(g314_n),
    .din1(G10_n_spl_000),
    .din2(G17_n_spl_100)
  );


  LA
  g_g315_p
  (
    .dout(g315_p),
    .din1(G9_p_spl_000),
    .din2(G18_p_spl_100)
  );


  FA
  g_g315_n
  (
    .dout(g315_n),
    .din1(G9_n_spl_000),
    .din2(G18_n_spl_100)
  );


  LA
  g_g316_p
  (
    .dout(g316_p),
    .din1(g314_p_spl_),
    .din2(g315_n_spl_)
  );


  FA
  g_g316_n
  (
    .dout(g316_n),
    .din1(g314_n_spl_),
    .din2(g315_p_spl_)
  );


  LA
  g_g317_p
  (
    .dout(g317_p),
    .din1(g314_p_spl_),
    .din2(g316_n_spl_)
  );


  FA
  g_g317_n
  (
    .dout(g317_n),
    .din1(g314_n_spl_),
    .din2(g316_p_spl_)
  );


  LA
  g_g318_p
  (
    .dout(g318_p),
    .din1(g315_n_spl_),
    .din2(g316_n_spl_)
  );


  FA
  g_g318_n
  (
    .dout(g318_n),
    .din1(g315_p_spl_),
    .din2(g316_p_spl_)
  );


  LA
  g_g319_p
  (
    .dout(g319_p),
    .din1(g317_n_spl_0),
    .din2(g318_n)
  );


  FA
  g_g319_n
  (
    .dout(g319_n),
    .din1(g317_p_spl_0),
    .din2(g318_p)
  );


  LA
  g_g320_p
  (
    .dout(g320_p),
    .din1(g254_n_spl_0),
    .din2(g319_n_spl_)
  );


  FA
  g_g320_n
  (
    .dout(g320_n),
    .din1(g254_p_spl_0),
    .din2(g319_p_spl_)
  );


  LA
  g_g321_p
  (
    .dout(g321_p),
    .din1(g254_p_spl_),
    .din2(g319_p_spl_)
  );


  FA
  g_g321_n
  (
    .dout(g321_n),
    .din1(g254_n_spl_),
    .din2(g319_n_spl_)
  );


  LA
  g_g322_p
  (
    .dout(g322_p),
    .din1(g320_n_spl_),
    .din2(g321_n)
  );


  FA
  g_g322_n
  (
    .dout(g322_n),
    .din1(g320_p_spl_),
    .din2(g321_p)
  );


  LA
  g_g323_p
  (
    .dout(g323_p),
    .din1(g313_n_spl_),
    .din2(g322_p_spl_)
  );


  FA
  g_g323_n
  (
    .dout(g323_n),
    .din1(g313_p_spl_),
    .din2(g322_n_spl_)
  );


  LA
  g_g324_p
  (
    .dout(g324_p),
    .din1(g313_p_spl_),
    .din2(g322_n_spl_)
  );


  FA
  g_g324_n
  (
    .dout(g324_n),
    .din1(g313_n_spl_),
    .din2(g322_p_spl_)
  );


  LA
  g_g325_p
  (
    .dout(g325_p),
    .din1(g323_n_spl_),
    .din2(g324_n)
  );


  FA
  g_g325_n
  (
    .dout(g325_n),
    .din1(g323_p_spl_),
    .din2(g324_p)
  );


  LA
  g_g326_p
  (
    .dout(g326_p),
    .din1(g312_n_spl_),
    .din2(g325_p_spl_)
  );


  FA
  g_g326_n
  (
    .dout(g326_n),
    .din1(g312_p_spl_),
    .din2(g325_n_spl_)
  );


  LA
  g_g327_p
  (
    .dout(g327_p),
    .din1(g312_p_spl_),
    .din2(g325_n_spl_)
  );


  FA
  g_g327_n
  (
    .dout(g327_n),
    .din1(g312_n_spl_),
    .din2(g325_p_spl_)
  );


  LA
  g_g328_p
  (
    .dout(g328_p),
    .din1(g326_n_spl_),
    .din2(g327_n)
  );


  FA
  g_g328_n
  (
    .dout(g328_n),
    .din1(g326_p_spl_),
    .din2(g327_p)
  );


  LA
  g_g329_p
  (
    .dout(g329_p),
    .din1(g311_n_spl_),
    .din2(g328_p_spl_)
  );


  FA
  g_g329_n
  (
    .dout(g329_n),
    .din1(g311_p_spl_),
    .din2(g328_n_spl_)
  );


  LA
  g_g330_p
  (
    .dout(g330_p),
    .din1(g311_p_spl_),
    .din2(g328_n_spl_)
  );


  FA
  g_g330_n
  (
    .dout(g330_n),
    .din1(g311_n_spl_),
    .din2(g328_p_spl_)
  );


  LA
  g_g331_p
  (
    .dout(g331_p),
    .din1(g329_n_spl_),
    .din2(g330_n)
  );


  FA
  g_g331_n
  (
    .dout(g331_n),
    .din1(g329_p_spl_),
    .din2(g330_p)
  );


  LA
  g_g332_p
  (
    .dout(g332_p),
    .din1(g310_n_spl_),
    .din2(g331_p_spl_)
  );


  FA
  g_g332_n
  (
    .dout(g332_n),
    .din1(g310_p_spl_),
    .din2(g331_n_spl_)
  );


  LA
  g_g333_p
  (
    .dout(g333_p),
    .din1(g310_p_spl_),
    .din2(g331_n_spl_)
  );


  FA
  g_g333_n
  (
    .dout(g333_n),
    .din1(g310_n_spl_),
    .din2(g331_p_spl_)
  );


  LA
  g_g334_p
  (
    .dout(g334_p),
    .din1(g332_n_spl_),
    .din2(g333_n)
  );


  FA
  g_g334_n
  (
    .dout(g334_n),
    .din1(g332_p_spl_),
    .din2(g333_p)
  );


  LA
  g_g335_p
  (
    .dout(g335_p),
    .din1(g309_n_spl_),
    .din2(g334_p_spl_)
  );


  FA
  g_g335_n
  (
    .dout(g335_n),
    .din1(g309_p_spl_),
    .din2(g334_n_spl_)
  );


  LA
  g_g336_p
  (
    .dout(g336_p),
    .din1(g309_p_spl_),
    .din2(g334_n_spl_)
  );


  FA
  g_g336_n
  (
    .dout(g336_n),
    .din1(g309_n_spl_),
    .din2(g334_p_spl_)
  );


  LA
  g_g337_p
  (
    .dout(g337_p),
    .din1(g335_n_spl_),
    .din2(g336_n)
  );


  FA
  g_g337_n
  (
    .dout(g337_n),
    .din1(g335_p_spl_),
    .din2(g336_p)
  );


  LA
  g_g338_p
  (
    .dout(g338_p),
    .din1(g308_n_spl_),
    .din2(g337_p_spl_)
  );


  FA
  g_g338_n
  (
    .dout(g338_n),
    .din1(g308_p_spl_),
    .din2(g337_n_spl_)
  );


  LA
  g_g339_p
  (
    .dout(g339_p),
    .din1(g308_p_spl_),
    .din2(g337_n_spl_)
  );


  FA
  g_g339_n
  (
    .dout(g339_n),
    .din1(g308_n_spl_),
    .din2(g337_p_spl_)
  );


  LA
  g_g340_p
  (
    .dout(g340_p),
    .din1(g338_n_spl_),
    .din2(g339_n)
  );


  FA
  g_g340_n
  (
    .dout(g340_n),
    .din1(g338_p_spl_),
    .din2(g339_p)
  );


  LA
  g_g341_p
  (
    .dout(g341_p),
    .din1(g307_n_spl_),
    .din2(g340_p_spl_)
  );


  FA
  g_g341_n
  (
    .dout(g341_n),
    .din1(g307_p_spl_),
    .din2(g340_n_spl_)
  );


  LA
  g_g342_p
  (
    .dout(g342_p),
    .din1(g307_p_spl_),
    .din2(g340_n_spl_)
  );


  FA
  g_g342_n
  (
    .dout(g342_n),
    .din1(g307_n_spl_),
    .din2(g340_p_spl_)
  );


  LA
  g_g343_p
  (
    .dout(g343_p),
    .din1(g341_n_spl_),
    .din2(g342_n)
  );


  FA
  g_g343_n
  (
    .dout(g343_n),
    .din1(g341_p_spl_),
    .din2(g342_p)
  );


  LA
  g_g344_p
  (
    .dout(g344_p),
    .din1(g306_n_spl_),
    .din2(g343_p_spl_)
  );


  FA
  g_g344_n
  (
    .dout(g344_n),
    .din1(g306_p_spl_),
    .din2(g343_n_spl_)
  );


  LA
  g_g345_p
  (
    .dout(g345_p),
    .din1(g306_p_spl_),
    .din2(g343_n_spl_)
  );


  FA
  g_g345_n
  (
    .dout(g345_n),
    .din1(g306_n_spl_),
    .din2(g343_p_spl_)
  );


  LA
  g_g346_p
  (
    .dout(g346_p),
    .din1(g344_n_spl_),
    .din2(g345_n)
  );


  FA
  g_g346_n
  (
    .dout(g346_n),
    .din1(g344_p_spl_),
    .din2(g345_p)
  );


  LA
  g_g347_p
  (
    .dout(g347_p),
    .din1(g305_n_spl_),
    .din2(g346_p_spl_)
  );


  FA
  g_g347_n
  (
    .dout(g347_n),
    .din1(g305_p_spl_),
    .din2(g346_n_spl_)
  );


  LA
  g_g348_p
  (
    .dout(g348_p),
    .din1(g305_p_spl_),
    .din2(g346_n_spl_)
  );


  FA
  g_g348_n
  (
    .dout(g348_n),
    .din1(g305_n_spl_),
    .din2(g346_p_spl_)
  );


  LA
  g_g349_p
  (
    .dout(g349_p),
    .din1(g347_n_spl_),
    .din2(g348_n)
  );


  FA
  g_g349_n
  (
    .dout(g349_n),
    .din1(g347_p_spl_),
    .din2(g348_p)
  );


  LA
  g_g350_p
  (
    .dout(g350_p),
    .din1(g304_n_spl_),
    .din2(g349_p_spl_)
  );


  FA
  g_g350_n
  (
    .dout(g350_n),
    .din1(g304_p_spl_),
    .din2(g349_n_spl_)
  );


  LA
  g_g351_p
  (
    .dout(g351_p),
    .din1(g304_p_spl_),
    .din2(g349_n_spl_)
  );


  FA
  g_g351_n
  (
    .dout(g351_n),
    .din1(g304_n_spl_),
    .din2(g349_p_spl_)
  );


  LA
  g_g352_p
  (
    .dout(g352_p),
    .din1(g350_n_spl_),
    .din2(g351_n)
  );


  FA
  g_g352_n
  (
    .dout(g352_n),
    .din1(g350_p_spl_),
    .din2(g351_p)
  );


  LA
  g_g353_p
  (
    .dout(g353_p),
    .din1(g303_n_spl_),
    .din2(g352_p_spl_)
  );


  FA
  g_g353_n
  (
    .dout(g353_n),
    .din1(g303_p_spl_),
    .din2(g352_n_spl_)
  );


  LA
  g_g354_p
  (
    .dout(g354_p),
    .din1(g303_p_spl_),
    .din2(g352_n_spl_)
  );


  FA
  g_g354_n
  (
    .dout(g354_n),
    .din1(g303_n_spl_),
    .din2(g352_p_spl_)
  );


  LA
  g_g355_p
  (
    .dout(g355_p),
    .din1(g353_n_spl_),
    .din2(g354_n)
  );


  FA
  g_g355_n
  (
    .dout(g355_n),
    .din1(g353_p_spl_),
    .din2(g354_p)
  );


  LA
  g_g356_p
  (
    .dout(g356_p),
    .din1(g302_n_spl_),
    .din2(g355_p_spl_)
  );


  FA
  g_g356_n
  (
    .dout(g356_n),
    .din1(g302_p_spl_),
    .din2(g355_n_spl_)
  );


  LA
  g_g357_p
  (
    .dout(g357_p),
    .din1(g302_p_spl_),
    .din2(g355_n_spl_)
  );


  FA
  g_g357_n
  (
    .dout(g357_n),
    .din1(g302_n_spl_),
    .din2(g355_p_spl_)
  );


  LA
  g_g358_p
  (
    .dout(g358_p),
    .din1(g356_n_spl_),
    .din2(g357_n)
  );


  FA
  g_g358_n
  (
    .dout(g358_n),
    .din1(g356_p_spl_),
    .din2(g357_p)
  );


  LA
  g_g359_p
  (
    .dout(g359_p),
    .din1(g301_n_spl_),
    .din2(g358_p_spl_)
  );


  FA
  g_g359_n
  (
    .dout(g359_n),
    .din1(g301_p_spl_),
    .din2(g358_n_spl_)
  );


  LA
  g_g360_p
  (
    .dout(g360_p),
    .din1(g301_p_spl_),
    .din2(g358_n_spl_)
  );


  FA
  g_g360_n
  (
    .dout(g360_n),
    .din1(g301_n_spl_),
    .din2(g358_p_spl_)
  );


  LA
  g_g361_p
  (
    .dout(g361_p),
    .din1(g359_n_spl_),
    .din2(g360_n)
  );


  FA
  g_g361_n
  (
    .dout(g361_n),
    .din1(g359_p_spl_),
    .din2(g360_p)
  );


  LA
  g_g362_p
  (
    .dout(g362_p),
    .din1(g300_n_spl_),
    .din2(g361_p_spl_)
  );


  FA
  g_g362_n
  (
    .dout(g362_n),
    .din1(g300_p_spl_),
    .din2(g361_n_spl_)
  );


  LA
  g_g363_p
  (
    .dout(g363_p),
    .din1(g300_p_spl_),
    .din2(g361_n_spl_)
  );


  FA
  g_g363_n
  (
    .dout(g363_n),
    .din1(g300_n_spl_),
    .din2(g361_p_spl_)
  );


  LA
  g_g364_p
  (
    .dout(g364_p),
    .din1(g362_n_spl_),
    .din2(g363_n)
  );


  FA
  g_g364_n
  (
    .dout(g364_n),
    .din1(g362_p_spl_),
    .din2(g363_p)
  );


  LA
  g_g365_p
  (
    .dout(g365_p),
    .din1(g299_n),
    .din2(g364_p)
  );


  FA
  g_g365_n
  (
    .dout(g365_n),
    .din1(g299_p_spl_),
    .din2(g364_n_spl_)
  );


  LA
  g_g366_p
  (
    .dout(g366_p),
    .din1(g299_p_spl_),
    .din2(g364_n_spl_)
  );


  FA
  g_g367_n
  (
    .dout(g367_n),
    .din1(g365_p_spl_),
    .din2(g366_p)
  );


  LA
  g_g368_p
  (
    .dout(g368_p),
    .din1(G1_p_spl_101),
    .din2(G27_p_spl_000)
  );


  FA
  g_g368_n
  (
    .dout(g368_n),
    .din1(G1_n_spl_100),
    .din2(G27_n_spl_000)
  );


  LA
  g_g369_p
  (
    .dout(g369_p),
    .din1(g362_n_spl_),
    .din2(g365_n)
  );


  FA
  g_g369_n
  (
    .dout(g369_n),
    .din1(g362_p_spl_),
    .din2(g365_p_spl_)
  );


  LA
  g_g370_p
  (
    .dout(g370_p),
    .din1(G2_p_spl_100),
    .din2(G26_p_spl_000)
  );


  FA
  g_g370_n
  (
    .dout(g370_n),
    .din1(G2_n_spl_100),
    .din2(G26_n_spl_000)
  );


  LA
  g_g371_p
  (
    .dout(g371_p),
    .din1(g356_n_spl_),
    .din2(g359_n_spl_)
  );


  FA
  g_g371_n
  (
    .dout(g371_n),
    .din1(g356_p_spl_),
    .din2(g359_p_spl_)
  );


  LA
  g_g372_p
  (
    .dout(g372_p),
    .din1(G3_p_spl_100),
    .din2(G25_p_spl_001)
  );


  FA
  g_g372_n
  (
    .dout(g372_n),
    .din1(G3_n_spl_100),
    .din2(G25_n_spl_001)
  );


  LA
  g_g373_p
  (
    .dout(g373_p),
    .din1(g350_n_spl_),
    .din2(g353_n_spl_)
  );


  FA
  g_g373_n
  (
    .dout(g373_n),
    .din1(g350_p_spl_),
    .din2(g353_p_spl_)
  );


  LA
  g_g374_p
  (
    .dout(g374_p),
    .din1(G4_p_spl_011),
    .din2(G24_p_spl_001)
  );


  FA
  g_g374_n
  (
    .dout(g374_n),
    .din1(G4_n_spl_011),
    .din2(G24_n_spl_001)
  );


  LA
  g_g375_p
  (
    .dout(g375_p),
    .din1(g344_n_spl_),
    .din2(g347_n_spl_)
  );


  FA
  g_g375_n
  (
    .dout(g375_n),
    .din1(g344_p_spl_),
    .din2(g347_p_spl_)
  );


  LA
  g_g376_p
  (
    .dout(g376_p),
    .din1(G5_p_spl_011),
    .din2(G23_p_spl_010)
  );


  FA
  g_g376_n
  (
    .dout(g376_n),
    .din1(G5_n_spl_011),
    .din2(G23_n_spl_010)
  );


  LA
  g_g377_p
  (
    .dout(g377_p),
    .din1(g338_n_spl_),
    .din2(g341_n_spl_)
  );


  FA
  g_g377_n
  (
    .dout(g377_n),
    .din1(g338_p_spl_),
    .din2(g341_p_spl_)
  );


  LA
  g_g378_p
  (
    .dout(g378_p),
    .din1(G6_p_spl_010),
    .din2(G22_p_spl_010)
  );


  FA
  g_g378_n
  (
    .dout(g378_n),
    .din1(G6_n_spl_010),
    .din2(G22_n_spl_010)
  );


  LA
  g_g379_p
  (
    .dout(g379_p),
    .din1(g332_n_spl_),
    .din2(g335_n_spl_)
  );


  FA
  g_g379_n
  (
    .dout(g379_n),
    .din1(g332_p_spl_),
    .din2(g335_p_spl_)
  );


  LA
  g_g380_p
  (
    .dout(g380_p),
    .din1(G7_p_spl_010),
    .din2(G21_p_spl_011)
  );


  FA
  g_g380_n
  (
    .dout(g380_n),
    .din1(G7_n_spl_010),
    .din2(G21_n_spl_011)
  );


  LA
  g_g381_p
  (
    .dout(g381_p),
    .din1(g326_n_spl_),
    .din2(g329_n_spl_)
  );


  FA
  g_g381_n
  (
    .dout(g381_n),
    .din1(g326_p_spl_),
    .din2(g329_p_spl_)
  );


  LA
  g_g382_p
  (
    .dout(g382_p),
    .din1(G8_p_spl_001),
    .din2(G20_p_spl_011)
  );


  FA
  g_g382_n
  (
    .dout(g382_n),
    .din1(G8_n_spl_001),
    .din2(G20_n_spl_011)
  );


  LA
  g_g383_p
  (
    .dout(g383_p),
    .din1(g320_n_spl_),
    .din2(g323_n_spl_)
  );


  FA
  g_g383_n
  (
    .dout(g383_n),
    .din1(g320_p_spl_),
    .din2(g323_p_spl_)
  );


  LA
  g_g384_p
  (
    .dout(g384_p),
    .din1(G9_p_spl_001),
    .din2(G19_p_spl_100)
  );


  FA
  g_g384_n
  (
    .dout(g384_n),
    .din1(G9_n_spl_001),
    .din2(G19_n_spl_100)
  );


  LA
  g_g385_p
  (
    .dout(g385_p),
    .din1(G11_p_spl_000),
    .din2(G17_p_spl_101)
  );


  FA
  g_g385_n
  (
    .dout(g385_n),
    .din1(G11_n_spl_000),
    .din2(G17_n_spl_100)
  );


  LA
  g_g386_p
  (
    .dout(g386_p),
    .din1(G10_p_spl_000),
    .din2(G18_p_spl_100)
  );


  FA
  g_g386_n
  (
    .dout(g386_n),
    .din1(G10_n_spl_000),
    .din2(G18_n_spl_100)
  );


  LA
  g_g387_p
  (
    .dout(g387_p),
    .din1(g385_p_spl_),
    .din2(g386_n_spl_)
  );


  FA
  g_g387_n
  (
    .dout(g387_n),
    .din1(g385_n_spl_),
    .din2(g386_p_spl_)
  );


  LA
  g_g388_p
  (
    .dout(g388_p),
    .din1(g385_p_spl_),
    .din2(g387_n_spl_)
  );


  FA
  g_g388_n
  (
    .dout(g388_n),
    .din1(g385_n_spl_),
    .din2(g387_p_spl_)
  );


  LA
  g_g389_p
  (
    .dout(g389_p),
    .din1(g386_n_spl_),
    .din2(g387_n_spl_)
  );


  FA
  g_g389_n
  (
    .dout(g389_n),
    .din1(g386_p_spl_),
    .din2(g387_p_spl_)
  );


  LA
  g_g390_p
  (
    .dout(g390_p),
    .din1(g388_n_spl_0),
    .din2(g389_n)
  );


  FA
  g_g390_n
  (
    .dout(g390_n),
    .din1(g388_p_spl_0),
    .din2(g389_p)
  );


  LA
  g_g391_p
  (
    .dout(g391_p),
    .din1(g317_n_spl_0),
    .din2(g390_n_spl_)
  );


  FA
  g_g391_n
  (
    .dout(g391_n),
    .din1(g317_p_spl_0),
    .din2(g390_p_spl_)
  );


  LA
  g_g392_p
  (
    .dout(g392_p),
    .din1(g317_p_spl_),
    .din2(g390_p_spl_)
  );


  FA
  g_g392_n
  (
    .dout(g392_n),
    .din1(g317_n_spl_),
    .din2(g390_n_spl_)
  );


  LA
  g_g393_p
  (
    .dout(g393_p),
    .din1(g391_n_spl_),
    .din2(g392_n)
  );


  FA
  g_g393_n
  (
    .dout(g393_n),
    .din1(g391_p_spl_),
    .din2(g392_p)
  );


  LA
  g_g394_p
  (
    .dout(g394_p),
    .din1(g384_n_spl_),
    .din2(g393_p_spl_)
  );


  FA
  g_g394_n
  (
    .dout(g394_n),
    .din1(g384_p_spl_),
    .din2(g393_n_spl_)
  );


  LA
  g_g395_p
  (
    .dout(g395_p),
    .din1(g384_p_spl_),
    .din2(g393_n_spl_)
  );


  FA
  g_g395_n
  (
    .dout(g395_n),
    .din1(g384_n_spl_),
    .din2(g393_p_spl_)
  );


  LA
  g_g396_p
  (
    .dout(g396_p),
    .din1(g394_n_spl_),
    .din2(g395_n)
  );


  FA
  g_g396_n
  (
    .dout(g396_n),
    .din1(g394_p_spl_),
    .din2(g395_p)
  );


  LA
  g_g397_p
  (
    .dout(g397_p),
    .din1(g383_n_spl_),
    .din2(g396_p_spl_)
  );


  FA
  g_g397_n
  (
    .dout(g397_n),
    .din1(g383_p_spl_),
    .din2(g396_n_spl_)
  );


  LA
  g_g398_p
  (
    .dout(g398_p),
    .din1(g383_p_spl_),
    .din2(g396_n_spl_)
  );


  FA
  g_g398_n
  (
    .dout(g398_n),
    .din1(g383_n_spl_),
    .din2(g396_p_spl_)
  );


  LA
  g_g399_p
  (
    .dout(g399_p),
    .din1(g397_n_spl_),
    .din2(g398_n)
  );


  FA
  g_g399_n
  (
    .dout(g399_n),
    .din1(g397_p_spl_),
    .din2(g398_p)
  );


  LA
  g_g400_p
  (
    .dout(g400_p),
    .din1(g382_n_spl_),
    .din2(g399_p_spl_)
  );


  FA
  g_g400_n
  (
    .dout(g400_n),
    .din1(g382_p_spl_),
    .din2(g399_n_spl_)
  );


  LA
  g_g401_p
  (
    .dout(g401_p),
    .din1(g382_p_spl_),
    .din2(g399_n_spl_)
  );


  FA
  g_g401_n
  (
    .dout(g401_n),
    .din1(g382_n_spl_),
    .din2(g399_p_spl_)
  );


  LA
  g_g402_p
  (
    .dout(g402_p),
    .din1(g400_n_spl_),
    .din2(g401_n)
  );


  FA
  g_g402_n
  (
    .dout(g402_n),
    .din1(g400_p_spl_),
    .din2(g401_p)
  );


  LA
  g_g403_p
  (
    .dout(g403_p),
    .din1(g381_n_spl_),
    .din2(g402_p_spl_)
  );


  FA
  g_g403_n
  (
    .dout(g403_n),
    .din1(g381_p_spl_),
    .din2(g402_n_spl_)
  );


  LA
  g_g404_p
  (
    .dout(g404_p),
    .din1(g381_p_spl_),
    .din2(g402_n_spl_)
  );


  FA
  g_g404_n
  (
    .dout(g404_n),
    .din1(g381_n_spl_),
    .din2(g402_p_spl_)
  );


  LA
  g_g405_p
  (
    .dout(g405_p),
    .din1(g403_n_spl_),
    .din2(g404_n)
  );


  FA
  g_g405_n
  (
    .dout(g405_n),
    .din1(g403_p_spl_),
    .din2(g404_p)
  );


  LA
  g_g406_p
  (
    .dout(g406_p),
    .din1(g380_n_spl_),
    .din2(g405_p_spl_)
  );


  FA
  g_g406_n
  (
    .dout(g406_n),
    .din1(g380_p_spl_),
    .din2(g405_n_spl_)
  );


  LA
  g_g407_p
  (
    .dout(g407_p),
    .din1(g380_p_spl_),
    .din2(g405_n_spl_)
  );


  FA
  g_g407_n
  (
    .dout(g407_n),
    .din1(g380_n_spl_),
    .din2(g405_p_spl_)
  );


  LA
  g_g408_p
  (
    .dout(g408_p),
    .din1(g406_n_spl_),
    .din2(g407_n)
  );


  FA
  g_g408_n
  (
    .dout(g408_n),
    .din1(g406_p_spl_),
    .din2(g407_p)
  );


  LA
  g_g409_p
  (
    .dout(g409_p),
    .din1(g379_n_spl_),
    .din2(g408_p_spl_)
  );


  FA
  g_g409_n
  (
    .dout(g409_n),
    .din1(g379_p_spl_),
    .din2(g408_n_spl_)
  );


  LA
  g_g410_p
  (
    .dout(g410_p),
    .din1(g379_p_spl_),
    .din2(g408_n_spl_)
  );


  FA
  g_g410_n
  (
    .dout(g410_n),
    .din1(g379_n_spl_),
    .din2(g408_p_spl_)
  );


  LA
  g_g411_p
  (
    .dout(g411_p),
    .din1(g409_n_spl_),
    .din2(g410_n)
  );


  FA
  g_g411_n
  (
    .dout(g411_n),
    .din1(g409_p_spl_),
    .din2(g410_p)
  );


  LA
  g_g412_p
  (
    .dout(g412_p),
    .din1(g378_n_spl_),
    .din2(g411_p_spl_)
  );


  FA
  g_g412_n
  (
    .dout(g412_n),
    .din1(g378_p_spl_),
    .din2(g411_n_spl_)
  );


  LA
  g_g413_p
  (
    .dout(g413_p),
    .din1(g378_p_spl_),
    .din2(g411_n_spl_)
  );


  FA
  g_g413_n
  (
    .dout(g413_n),
    .din1(g378_n_spl_),
    .din2(g411_p_spl_)
  );


  LA
  g_g414_p
  (
    .dout(g414_p),
    .din1(g412_n_spl_),
    .din2(g413_n)
  );


  FA
  g_g414_n
  (
    .dout(g414_n),
    .din1(g412_p_spl_),
    .din2(g413_p)
  );


  LA
  g_g415_p
  (
    .dout(g415_p),
    .din1(g377_n_spl_),
    .din2(g414_p_spl_)
  );


  FA
  g_g415_n
  (
    .dout(g415_n),
    .din1(g377_p_spl_),
    .din2(g414_n_spl_)
  );


  LA
  g_g416_p
  (
    .dout(g416_p),
    .din1(g377_p_spl_),
    .din2(g414_n_spl_)
  );


  FA
  g_g416_n
  (
    .dout(g416_n),
    .din1(g377_n_spl_),
    .din2(g414_p_spl_)
  );


  LA
  g_g417_p
  (
    .dout(g417_p),
    .din1(g415_n_spl_),
    .din2(g416_n)
  );


  FA
  g_g417_n
  (
    .dout(g417_n),
    .din1(g415_p_spl_),
    .din2(g416_p)
  );


  LA
  g_g418_p
  (
    .dout(g418_p),
    .din1(g376_n_spl_),
    .din2(g417_p_spl_)
  );


  FA
  g_g418_n
  (
    .dout(g418_n),
    .din1(g376_p_spl_),
    .din2(g417_n_spl_)
  );


  LA
  g_g419_p
  (
    .dout(g419_p),
    .din1(g376_p_spl_),
    .din2(g417_n_spl_)
  );


  FA
  g_g419_n
  (
    .dout(g419_n),
    .din1(g376_n_spl_),
    .din2(g417_p_spl_)
  );


  LA
  g_g420_p
  (
    .dout(g420_p),
    .din1(g418_n_spl_),
    .din2(g419_n)
  );


  FA
  g_g420_n
  (
    .dout(g420_n),
    .din1(g418_p_spl_),
    .din2(g419_p)
  );


  LA
  g_g421_p
  (
    .dout(g421_p),
    .din1(g375_n_spl_),
    .din2(g420_p_spl_)
  );


  FA
  g_g421_n
  (
    .dout(g421_n),
    .din1(g375_p_spl_),
    .din2(g420_n_spl_)
  );


  LA
  g_g422_p
  (
    .dout(g422_p),
    .din1(g375_p_spl_),
    .din2(g420_n_spl_)
  );


  FA
  g_g422_n
  (
    .dout(g422_n),
    .din1(g375_n_spl_),
    .din2(g420_p_spl_)
  );


  LA
  g_g423_p
  (
    .dout(g423_p),
    .din1(g421_n_spl_),
    .din2(g422_n)
  );


  FA
  g_g423_n
  (
    .dout(g423_n),
    .din1(g421_p_spl_),
    .din2(g422_p)
  );


  LA
  g_g424_p
  (
    .dout(g424_p),
    .din1(g374_n_spl_),
    .din2(g423_p_spl_)
  );


  FA
  g_g424_n
  (
    .dout(g424_n),
    .din1(g374_p_spl_),
    .din2(g423_n_spl_)
  );


  LA
  g_g425_p
  (
    .dout(g425_p),
    .din1(g374_p_spl_),
    .din2(g423_n_spl_)
  );


  FA
  g_g425_n
  (
    .dout(g425_n),
    .din1(g374_n_spl_),
    .din2(g423_p_spl_)
  );


  LA
  g_g426_p
  (
    .dout(g426_p),
    .din1(g424_n_spl_),
    .din2(g425_n)
  );


  FA
  g_g426_n
  (
    .dout(g426_n),
    .din1(g424_p_spl_),
    .din2(g425_p)
  );


  LA
  g_g427_p
  (
    .dout(g427_p),
    .din1(g373_n_spl_),
    .din2(g426_p_spl_)
  );


  FA
  g_g427_n
  (
    .dout(g427_n),
    .din1(g373_p_spl_),
    .din2(g426_n_spl_)
  );


  LA
  g_g428_p
  (
    .dout(g428_p),
    .din1(g373_p_spl_),
    .din2(g426_n_spl_)
  );


  FA
  g_g428_n
  (
    .dout(g428_n),
    .din1(g373_n_spl_),
    .din2(g426_p_spl_)
  );


  LA
  g_g429_p
  (
    .dout(g429_p),
    .din1(g427_n_spl_),
    .din2(g428_n)
  );


  FA
  g_g429_n
  (
    .dout(g429_n),
    .din1(g427_p_spl_),
    .din2(g428_p)
  );


  LA
  g_g430_p
  (
    .dout(g430_p),
    .din1(g372_n_spl_),
    .din2(g429_p_spl_)
  );


  FA
  g_g430_n
  (
    .dout(g430_n),
    .din1(g372_p_spl_),
    .din2(g429_n_spl_)
  );


  LA
  g_g431_p
  (
    .dout(g431_p),
    .din1(g372_p_spl_),
    .din2(g429_n_spl_)
  );


  FA
  g_g431_n
  (
    .dout(g431_n),
    .din1(g372_n_spl_),
    .din2(g429_p_spl_)
  );


  LA
  g_g432_p
  (
    .dout(g432_p),
    .din1(g430_n_spl_),
    .din2(g431_n)
  );


  FA
  g_g432_n
  (
    .dout(g432_n),
    .din1(g430_p_spl_),
    .din2(g431_p)
  );


  LA
  g_g433_p
  (
    .dout(g433_p),
    .din1(g371_n_spl_),
    .din2(g432_p_spl_)
  );


  FA
  g_g433_n
  (
    .dout(g433_n),
    .din1(g371_p_spl_),
    .din2(g432_n_spl_)
  );


  LA
  g_g434_p
  (
    .dout(g434_p),
    .din1(g371_p_spl_),
    .din2(g432_n_spl_)
  );


  FA
  g_g434_n
  (
    .dout(g434_n),
    .din1(g371_n_spl_),
    .din2(g432_p_spl_)
  );


  LA
  g_g435_p
  (
    .dout(g435_p),
    .din1(g433_n_spl_),
    .din2(g434_n)
  );


  FA
  g_g435_n
  (
    .dout(g435_n),
    .din1(g433_p_spl_),
    .din2(g434_p)
  );


  LA
  g_g436_p
  (
    .dout(g436_p),
    .din1(g370_n_spl_),
    .din2(g435_p_spl_)
  );


  FA
  g_g436_n
  (
    .dout(g436_n),
    .din1(g370_p_spl_),
    .din2(g435_n_spl_)
  );


  LA
  g_g437_p
  (
    .dout(g437_p),
    .din1(g370_p_spl_),
    .din2(g435_n_spl_)
  );


  FA
  g_g437_n
  (
    .dout(g437_n),
    .din1(g370_n_spl_),
    .din2(g435_p_spl_)
  );


  LA
  g_g438_p
  (
    .dout(g438_p),
    .din1(g436_n_spl_),
    .din2(g437_n)
  );


  FA
  g_g438_n
  (
    .dout(g438_n),
    .din1(g436_p_spl_),
    .din2(g437_p)
  );


  LA
  g_g439_p
  (
    .dout(g439_p),
    .din1(g369_n_spl_),
    .din2(g438_p_spl_)
  );


  FA
  g_g439_n
  (
    .dout(g439_n),
    .din1(g369_p_spl_),
    .din2(g438_n_spl_)
  );


  LA
  g_g440_p
  (
    .dout(g440_p),
    .din1(g369_p_spl_),
    .din2(g438_n_spl_)
  );


  FA
  g_g440_n
  (
    .dout(g440_n),
    .din1(g369_n_spl_),
    .din2(g438_p_spl_)
  );


  LA
  g_g441_p
  (
    .dout(g441_p),
    .din1(g439_n_spl_),
    .din2(g440_n)
  );


  FA
  g_g441_n
  (
    .dout(g441_n),
    .din1(g439_p_spl_),
    .din2(g440_p)
  );


  LA
  g_g442_p
  (
    .dout(g442_p),
    .din1(g368_n),
    .din2(g441_p)
  );


  FA
  g_g442_n
  (
    .dout(g442_n),
    .din1(g368_p_spl_),
    .din2(g441_n_spl_)
  );


  LA
  g_g443_p
  (
    .dout(g443_p),
    .din1(g368_p_spl_),
    .din2(g441_n_spl_)
  );


  FA
  g_g444_n
  (
    .dout(g444_n),
    .din1(g442_p_spl_),
    .din2(g443_p)
  );


  LA
  g_g445_p
  (
    .dout(g445_p),
    .din1(G1_p_spl_101),
    .din2(G28_p_spl_000)
  );


  FA
  g_g445_n
  (
    .dout(g445_n),
    .din1(G1_n_spl_101),
    .din2(G28_n_spl_000)
  );


  LA
  g_g446_p
  (
    .dout(g446_p),
    .din1(g439_n_spl_),
    .din2(g442_n)
  );


  FA
  g_g446_n
  (
    .dout(g446_n),
    .din1(g439_p_spl_),
    .din2(g442_p_spl_)
  );


  LA
  g_g447_p
  (
    .dout(g447_p),
    .din1(G2_p_spl_101),
    .din2(G27_p_spl_000)
  );


  FA
  g_g447_n
  (
    .dout(g447_n),
    .din1(G2_n_spl_101),
    .din2(G27_n_spl_000)
  );


  LA
  g_g448_p
  (
    .dout(g448_p),
    .din1(g433_n_spl_),
    .din2(g436_n_spl_)
  );


  FA
  g_g448_n
  (
    .dout(g448_n),
    .din1(g433_p_spl_),
    .din2(g436_p_spl_)
  );


  LA
  g_g449_p
  (
    .dout(g449_p),
    .din1(G3_p_spl_100),
    .din2(G26_p_spl_001)
  );


  FA
  g_g449_n
  (
    .dout(g449_n),
    .din1(G3_n_spl_100),
    .din2(G26_n_spl_001)
  );


  LA
  g_g450_p
  (
    .dout(g450_p),
    .din1(g427_n_spl_),
    .din2(g430_n_spl_)
  );


  FA
  g_g450_n
  (
    .dout(g450_n),
    .din1(g427_p_spl_),
    .din2(g430_p_spl_)
  );


  LA
  g_g451_p
  (
    .dout(g451_p),
    .din1(G4_p_spl_100),
    .din2(G25_p_spl_001)
  );


  FA
  g_g451_n
  (
    .dout(g451_n),
    .din1(G4_n_spl_100),
    .din2(G25_n_spl_001)
  );


  LA
  g_g452_p
  (
    .dout(g452_p),
    .din1(g421_n_spl_),
    .din2(g424_n_spl_)
  );


  FA
  g_g452_n
  (
    .dout(g452_n),
    .din1(g421_p_spl_),
    .din2(g424_p_spl_)
  );


  LA
  g_g453_p
  (
    .dout(g453_p),
    .din1(G5_p_spl_011),
    .din2(G24_p_spl_010)
  );


  FA
  g_g453_n
  (
    .dout(g453_n),
    .din1(G5_n_spl_011),
    .din2(G24_n_spl_010)
  );


  LA
  g_g454_p
  (
    .dout(g454_p),
    .din1(g415_n_spl_),
    .din2(g418_n_spl_)
  );


  FA
  g_g454_n
  (
    .dout(g454_n),
    .din1(g415_p_spl_),
    .din2(g418_p_spl_)
  );


  LA
  g_g455_p
  (
    .dout(g455_p),
    .din1(G6_p_spl_011),
    .din2(G23_p_spl_010)
  );


  FA
  g_g455_n
  (
    .dout(g455_n),
    .din1(G6_n_spl_011),
    .din2(G23_n_spl_010)
  );


  LA
  g_g456_p
  (
    .dout(g456_p),
    .din1(g409_n_spl_),
    .din2(g412_n_spl_)
  );


  FA
  g_g456_n
  (
    .dout(g456_n),
    .din1(g409_p_spl_),
    .din2(g412_p_spl_)
  );


  LA
  g_g457_p
  (
    .dout(g457_p),
    .din1(G7_p_spl_010),
    .din2(G22_p_spl_011)
  );


  FA
  g_g457_n
  (
    .dout(g457_n),
    .din1(G7_n_spl_010),
    .din2(G22_n_spl_011)
  );


  LA
  g_g458_p
  (
    .dout(g458_p),
    .din1(g403_n_spl_),
    .din2(g406_n_spl_)
  );


  FA
  g_g458_n
  (
    .dout(g458_n),
    .din1(g403_p_spl_),
    .din2(g406_p_spl_)
  );


  LA
  g_g459_p
  (
    .dout(g459_p),
    .din1(G8_p_spl_010),
    .din2(G21_p_spl_011)
  );


  FA
  g_g459_n
  (
    .dout(g459_n),
    .din1(G8_n_spl_010),
    .din2(G21_n_spl_011)
  );


  LA
  g_g460_p
  (
    .dout(g460_p),
    .din1(g397_n_spl_),
    .din2(g400_n_spl_)
  );


  FA
  g_g460_n
  (
    .dout(g460_n),
    .din1(g397_p_spl_),
    .din2(g400_p_spl_)
  );


  LA
  g_g461_p
  (
    .dout(g461_p),
    .din1(G9_p_spl_001),
    .din2(G20_p_spl_100)
  );


  FA
  g_g461_n
  (
    .dout(g461_n),
    .din1(G9_n_spl_001),
    .din2(G20_n_spl_100)
  );


  LA
  g_g462_p
  (
    .dout(g462_p),
    .din1(g391_n_spl_),
    .din2(g394_n_spl_)
  );


  FA
  g_g462_n
  (
    .dout(g462_n),
    .din1(g391_p_spl_),
    .din2(g394_p_spl_)
  );


  LA
  g_g463_p
  (
    .dout(g463_p),
    .din1(G10_p_spl_001),
    .din2(G19_p_spl_100)
  );


  FA
  g_g463_n
  (
    .dout(g463_n),
    .din1(G10_n_spl_001),
    .din2(G19_n_spl_100)
  );


  LA
  g_g464_p
  (
    .dout(g464_p),
    .din1(G12_p_spl_000),
    .din2(G17_p_spl_101)
  );


  FA
  g_g464_n
  (
    .dout(g464_n),
    .din1(G12_n_spl_000),
    .din2(G17_n_spl_101)
  );


  LA
  g_g465_p
  (
    .dout(g465_p),
    .din1(G11_p_spl_000),
    .din2(G18_p_spl_101)
  );


  FA
  g_g465_n
  (
    .dout(g465_n),
    .din1(G11_n_spl_000),
    .din2(G18_n_spl_101)
  );


  LA
  g_g466_p
  (
    .dout(g466_p),
    .din1(g464_p_spl_),
    .din2(g465_n_spl_)
  );


  FA
  g_g466_n
  (
    .dout(g466_n),
    .din1(g464_n_spl_),
    .din2(g465_p_spl_)
  );


  LA
  g_g467_p
  (
    .dout(g467_p),
    .din1(g464_p_spl_),
    .din2(g466_n_spl_)
  );


  FA
  g_g467_n
  (
    .dout(g467_n),
    .din1(g464_n_spl_),
    .din2(g466_p_spl_)
  );


  LA
  g_g468_p
  (
    .dout(g468_p),
    .din1(g465_n_spl_),
    .din2(g466_n_spl_)
  );


  FA
  g_g468_n
  (
    .dout(g468_n),
    .din1(g465_p_spl_),
    .din2(g466_p_spl_)
  );


  LA
  g_g469_p
  (
    .dout(g469_p),
    .din1(g467_n_spl_0),
    .din2(g468_n)
  );


  FA
  g_g469_n
  (
    .dout(g469_n),
    .din1(g467_p_spl_0),
    .din2(g468_p)
  );


  LA
  g_g470_p
  (
    .dout(g470_p),
    .din1(g388_n_spl_0),
    .din2(g469_n_spl_)
  );


  FA
  g_g470_n
  (
    .dout(g470_n),
    .din1(g388_p_spl_0),
    .din2(g469_p_spl_)
  );


  LA
  g_g471_p
  (
    .dout(g471_p),
    .din1(g388_p_spl_),
    .din2(g469_p_spl_)
  );


  FA
  g_g471_n
  (
    .dout(g471_n),
    .din1(g388_n_spl_),
    .din2(g469_n_spl_)
  );


  LA
  g_g472_p
  (
    .dout(g472_p),
    .din1(g470_n_spl_),
    .din2(g471_n)
  );


  FA
  g_g472_n
  (
    .dout(g472_n),
    .din1(g470_p_spl_),
    .din2(g471_p)
  );


  LA
  g_g473_p
  (
    .dout(g473_p),
    .din1(g463_n_spl_),
    .din2(g472_p_spl_)
  );


  FA
  g_g473_n
  (
    .dout(g473_n),
    .din1(g463_p_spl_),
    .din2(g472_n_spl_)
  );


  LA
  g_g474_p
  (
    .dout(g474_p),
    .din1(g463_p_spl_),
    .din2(g472_n_spl_)
  );


  FA
  g_g474_n
  (
    .dout(g474_n),
    .din1(g463_n_spl_),
    .din2(g472_p_spl_)
  );


  LA
  g_g475_p
  (
    .dout(g475_p),
    .din1(g473_n_spl_),
    .din2(g474_n)
  );


  FA
  g_g475_n
  (
    .dout(g475_n),
    .din1(g473_p_spl_),
    .din2(g474_p)
  );


  LA
  g_g476_p
  (
    .dout(g476_p),
    .din1(g462_n_spl_),
    .din2(g475_p_spl_)
  );


  FA
  g_g476_n
  (
    .dout(g476_n),
    .din1(g462_p_spl_),
    .din2(g475_n_spl_)
  );


  LA
  g_g477_p
  (
    .dout(g477_p),
    .din1(g462_p_spl_),
    .din2(g475_n_spl_)
  );


  FA
  g_g477_n
  (
    .dout(g477_n),
    .din1(g462_n_spl_),
    .din2(g475_p_spl_)
  );


  LA
  g_g478_p
  (
    .dout(g478_p),
    .din1(g476_n_spl_),
    .din2(g477_n)
  );


  FA
  g_g478_n
  (
    .dout(g478_n),
    .din1(g476_p_spl_),
    .din2(g477_p)
  );


  LA
  g_g479_p
  (
    .dout(g479_p),
    .din1(g461_n_spl_),
    .din2(g478_p_spl_)
  );


  FA
  g_g479_n
  (
    .dout(g479_n),
    .din1(g461_p_spl_),
    .din2(g478_n_spl_)
  );


  LA
  g_g480_p
  (
    .dout(g480_p),
    .din1(g461_p_spl_),
    .din2(g478_n_spl_)
  );


  FA
  g_g480_n
  (
    .dout(g480_n),
    .din1(g461_n_spl_),
    .din2(g478_p_spl_)
  );


  LA
  g_g481_p
  (
    .dout(g481_p),
    .din1(g479_n_spl_),
    .din2(g480_n)
  );


  FA
  g_g481_n
  (
    .dout(g481_n),
    .din1(g479_p_spl_),
    .din2(g480_p)
  );


  LA
  g_g482_p
  (
    .dout(g482_p),
    .din1(g460_n_spl_),
    .din2(g481_p_spl_)
  );


  FA
  g_g482_n
  (
    .dout(g482_n),
    .din1(g460_p_spl_),
    .din2(g481_n_spl_)
  );


  LA
  g_g483_p
  (
    .dout(g483_p),
    .din1(g460_p_spl_),
    .din2(g481_n_spl_)
  );


  FA
  g_g483_n
  (
    .dout(g483_n),
    .din1(g460_n_spl_),
    .din2(g481_p_spl_)
  );


  LA
  g_g484_p
  (
    .dout(g484_p),
    .din1(g482_n_spl_),
    .din2(g483_n)
  );


  FA
  g_g484_n
  (
    .dout(g484_n),
    .din1(g482_p_spl_),
    .din2(g483_p)
  );


  LA
  g_g485_p
  (
    .dout(g485_p),
    .din1(g459_n_spl_),
    .din2(g484_p_spl_)
  );


  FA
  g_g485_n
  (
    .dout(g485_n),
    .din1(g459_p_spl_),
    .din2(g484_n_spl_)
  );


  LA
  g_g486_p
  (
    .dout(g486_p),
    .din1(g459_p_spl_),
    .din2(g484_n_spl_)
  );


  FA
  g_g486_n
  (
    .dout(g486_n),
    .din1(g459_n_spl_),
    .din2(g484_p_spl_)
  );


  LA
  g_g487_p
  (
    .dout(g487_p),
    .din1(g485_n_spl_),
    .din2(g486_n)
  );


  FA
  g_g487_n
  (
    .dout(g487_n),
    .din1(g485_p_spl_),
    .din2(g486_p)
  );


  LA
  g_g488_p
  (
    .dout(g488_p),
    .din1(g458_n_spl_),
    .din2(g487_p_spl_)
  );


  FA
  g_g488_n
  (
    .dout(g488_n),
    .din1(g458_p_spl_),
    .din2(g487_n_spl_)
  );


  LA
  g_g489_p
  (
    .dout(g489_p),
    .din1(g458_p_spl_),
    .din2(g487_n_spl_)
  );


  FA
  g_g489_n
  (
    .dout(g489_n),
    .din1(g458_n_spl_),
    .din2(g487_p_spl_)
  );


  LA
  g_g490_p
  (
    .dout(g490_p),
    .din1(g488_n_spl_),
    .din2(g489_n)
  );


  FA
  g_g490_n
  (
    .dout(g490_n),
    .din1(g488_p_spl_),
    .din2(g489_p)
  );


  LA
  g_g491_p
  (
    .dout(g491_p),
    .din1(g457_n_spl_),
    .din2(g490_p_spl_)
  );


  FA
  g_g491_n
  (
    .dout(g491_n),
    .din1(g457_p_spl_),
    .din2(g490_n_spl_)
  );


  LA
  g_g492_p
  (
    .dout(g492_p),
    .din1(g457_p_spl_),
    .din2(g490_n_spl_)
  );


  FA
  g_g492_n
  (
    .dout(g492_n),
    .din1(g457_n_spl_),
    .din2(g490_p_spl_)
  );


  LA
  g_g493_p
  (
    .dout(g493_p),
    .din1(g491_n_spl_),
    .din2(g492_n)
  );


  FA
  g_g493_n
  (
    .dout(g493_n),
    .din1(g491_p_spl_),
    .din2(g492_p)
  );


  LA
  g_g494_p
  (
    .dout(g494_p),
    .din1(g456_n_spl_),
    .din2(g493_p_spl_)
  );


  FA
  g_g494_n
  (
    .dout(g494_n),
    .din1(g456_p_spl_),
    .din2(g493_n_spl_)
  );


  LA
  g_g495_p
  (
    .dout(g495_p),
    .din1(g456_p_spl_),
    .din2(g493_n_spl_)
  );


  FA
  g_g495_n
  (
    .dout(g495_n),
    .din1(g456_n_spl_),
    .din2(g493_p_spl_)
  );


  LA
  g_g496_p
  (
    .dout(g496_p),
    .din1(g494_n_spl_),
    .din2(g495_n)
  );


  FA
  g_g496_n
  (
    .dout(g496_n),
    .din1(g494_p_spl_),
    .din2(g495_p)
  );


  LA
  g_g497_p
  (
    .dout(g497_p),
    .din1(g455_n_spl_),
    .din2(g496_p_spl_)
  );


  FA
  g_g497_n
  (
    .dout(g497_n),
    .din1(g455_p_spl_),
    .din2(g496_n_spl_)
  );


  LA
  g_g498_p
  (
    .dout(g498_p),
    .din1(g455_p_spl_),
    .din2(g496_n_spl_)
  );


  FA
  g_g498_n
  (
    .dout(g498_n),
    .din1(g455_n_spl_),
    .din2(g496_p_spl_)
  );


  LA
  g_g499_p
  (
    .dout(g499_p),
    .din1(g497_n_spl_),
    .din2(g498_n)
  );


  FA
  g_g499_n
  (
    .dout(g499_n),
    .din1(g497_p_spl_),
    .din2(g498_p)
  );


  LA
  g_g500_p
  (
    .dout(g500_p),
    .din1(g454_n_spl_),
    .din2(g499_p_spl_)
  );


  FA
  g_g500_n
  (
    .dout(g500_n),
    .din1(g454_p_spl_),
    .din2(g499_n_spl_)
  );


  LA
  g_g501_p
  (
    .dout(g501_p),
    .din1(g454_p_spl_),
    .din2(g499_n_spl_)
  );


  FA
  g_g501_n
  (
    .dout(g501_n),
    .din1(g454_n_spl_),
    .din2(g499_p_spl_)
  );


  LA
  g_g502_p
  (
    .dout(g502_p),
    .din1(g500_n_spl_),
    .din2(g501_n)
  );


  FA
  g_g502_n
  (
    .dout(g502_n),
    .din1(g500_p_spl_),
    .din2(g501_p)
  );


  LA
  g_g503_p
  (
    .dout(g503_p),
    .din1(g453_n_spl_),
    .din2(g502_p_spl_)
  );


  FA
  g_g503_n
  (
    .dout(g503_n),
    .din1(g453_p_spl_),
    .din2(g502_n_spl_)
  );


  LA
  g_g504_p
  (
    .dout(g504_p),
    .din1(g453_p_spl_),
    .din2(g502_n_spl_)
  );


  FA
  g_g504_n
  (
    .dout(g504_n),
    .din1(g453_n_spl_),
    .din2(g502_p_spl_)
  );


  LA
  g_g505_p
  (
    .dout(g505_p),
    .din1(g503_n_spl_),
    .din2(g504_n)
  );


  FA
  g_g505_n
  (
    .dout(g505_n),
    .din1(g503_p_spl_),
    .din2(g504_p)
  );


  LA
  g_g506_p
  (
    .dout(g506_p),
    .din1(g452_n_spl_),
    .din2(g505_p_spl_)
  );


  FA
  g_g506_n
  (
    .dout(g506_n),
    .din1(g452_p_spl_),
    .din2(g505_n_spl_)
  );


  LA
  g_g507_p
  (
    .dout(g507_p),
    .din1(g452_p_spl_),
    .din2(g505_n_spl_)
  );


  FA
  g_g507_n
  (
    .dout(g507_n),
    .din1(g452_n_spl_),
    .din2(g505_p_spl_)
  );


  LA
  g_g508_p
  (
    .dout(g508_p),
    .din1(g506_n_spl_),
    .din2(g507_n)
  );


  FA
  g_g508_n
  (
    .dout(g508_n),
    .din1(g506_p_spl_),
    .din2(g507_p)
  );


  LA
  g_g509_p
  (
    .dout(g509_p),
    .din1(g451_n_spl_),
    .din2(g508_p_spl_)
  );


  FA
  g_g509_n
  (
    .dout(g509_n),
    .din1(g451_p_spl_),
    .din2(g508_n_spl_)
  );


  LA
  g_g510_p
  (
    .dout(g510_p),
    .din1(g451_p_spl_),
    .din2(g508_n_spl_)
  );


  FA
  g_g510_n
  (
    .dout(g510_n),
    .din1(g451_n_spl_),
    .din2(g508_p_spl_)
  );


  LA
  g_g511_p
  (
    .dout(g511_p),
    .din1(g509_n_spl_),
    .din2(g510_n)
  );


  FA
  g_g511_n
  (
    .dout(g511_n),
    .din1(g509_p_spl_),
    .din2(g510_p)
  );


  LA
  g_g512_p
  (
    .dout(g512_p),
    .din1(g450_n_spl_),
    .din2(g511_p_spl_)
  );


  FA
  g_g512_n
  (
    .dout(g512_n),
    .din1(g450_p_spl_),
    .din2(g511_n_spl_)
  );


  LA
  g_g513_p
  (
    .dout(g513_p),
    .din1(g450_p_spl_),
    .din2(g511_n_spl_)
  );


  FA
  g_g513_n
  (
    .dout(g513_n),
    .din1(g450_n_spl_),
    .din2(g511_p_spl_)
  );


  LA
  g_g514_p
  (
    .dout(g514_p),
    .din1(g512_n_spl_),
    .din2(g513_n)
  );


  FA
  g_g514_n
  (
    .dout(g514_n),
    .din1(g512_p_spl_),
    .din2(g513_p)
  );


  LA
  g_g515_p
  (
    .dout(g515_p),
    .din1(g449_n_spl_),
    .din2(g514_p_spl_)
  );


  FA
  g_g515_n
  (
    .dout(g515_n),
    .din1(g449_p_spl_),
    .din2(g514_n_spl_)
  );


  LA
  g_g516_p
  (
    .dout(g516_p),
    .din1(g449_p_spl_),
    .din2(g514_n_spl_)
  );


  FA
  g_g516_n
  (
    .dout(g516_n),
    .din1(g449_n_spl_),
    .din2(g514_p_spl_)
  );


  LA
  g_g517_p
  (
    .dout(g517_p),
    .din1(g515_n_spl_),
    .din2(g516_n)
  );


  FA
  g_g517_n
  (
    .dout(g517_n),
    .din1(g515_p_spl_),
    .din2(g516_p)
  );


  LA
  g_g518_p
  (
    .dout(g518_p),
    .din1(g448_n_spl_),
    .din2(g517_p_spl_)
  );


  FA
  g_g518_n
  (
    .dout(g518_n),
    .din1(g448_p_spl_),
    .din2(g517_n_spl_)
  );


  LA
  g_g519_p
  (
    .dout(g519_p),
    .din1(g448_p_spl_),
    .din2(g517_n_spl_)
  );


  FA
  g_g519_n
  (
    .dout(g519_n),
    .din1(g448_n_spl_),
    .din2(g517_p_spl_)
  );


  LA
  g_g520_p
  (
    .dout(g520_p),
    .din1(g518_n_spl_),
    .din2(g519_n)
  );


  FA
  g_g520_n
  (
    .dout(g520_n),
    .din1(g518_p_spl_),
    .din2(g519_p)
  );


  LA
  g_g521_p
  (
    .dout(g521_p),
    .din1(g447_n_spl_),
    .din2(g520_p_spl_)
  );


  FA
  g_g521_n
  (
    .dout(g521_n),
    .din1(g447_p_spl_),
    .din2(g520_n_spl_)
  );


  LA
  g_g522_p
  (
    .dout(g522_p),
    .din1(g447_p_spl_),
    .din2(g520_n_spl_)
  );


  FA
  g_g522_n
  (
    .dout(g522_n),
    .din1(g447_n_spl_),
    .din2(g520_p_spl_)
  );


  LA
  g_g523_p
  (
    .dout(g523_p),
    .din1(g521_n_spl_),
    .din2(g522_n)
  );


  FA
  g_g523_n
  (
    .dout(g523_n),
    .din1(g521_p_spl_),
    .din2(g522_p)
  );


  LA
  g_g524_p
  (
    .dout(g524_p),
    .din1(g446_n_spl_),
    .din2(g523_p_spl_)
  );


  FA
  g_g524_n
  (
    .dout(g524_n),
    .din1(g446_p_spl_),
    .din2(g523_n_spl_)
  );


  LA
  g_g525_p
  (
    .dout(g525_p),
    .din1(g446_p_spl_),
    .din2(g523_n_spl_)
  );


  FA
  g_g525_n
  (
    .dout(g525_n),
    .din1(g446_n_spl_),
    .din2(g523_p_spl_)
  );


  LA
  g_g526_p
  (
    .dout(g526_p),
    .din1(g524_n_spl_),
    .din2(g525_n)
  );


  FA
  g_g526_n
  (
    .dout(g526_n),
    .din1(g524_p_spl_),
    .din2(g525_p)
  );


  LA
  g_g527_p
  (
    .dout(g527_p),
    .din1(g445_n),
    .din2(g526_p)
  );


  FA
  g_g527_n
  (
    .dout(g527_n),
    .din1(g445_p_spl_),
    .din2(g526_n_spl_)
  );


  LA
  g_g528_p
  (
    .dout(g528_p),
    .din1(g445_p_spl_),
    .din2(g526_n_spl_)
  );


  FA
  g_g529_n
  (
    .dout(g529_n),
    .din1(g527_p_spl_),
    .din2(g528_p)
  );


  LA
  g_g530_p
  (
    .dout(g530_p),
    .din1(G1_p_spl_110),
    .din2(G29_p_spl_000)
  );


  FA
  g_g530_n
  (
    .dout(g530_n),
    .din1(G1_n_spl_101),
    .din2(G29_n_spl_000)
  );


  LA
  g_g531_p
  (
    .dout(g531_p),
    .din1(g524_n_spl_),
    .din2(g527_n)
  );


  FA
  g_g531_n
  (
    .dout(g531_n),
    .din1(g524_p_spl_),
    .din2(g527_p_spl_)
  );


  LA
  g_g532_p
  (
    .dout(g532_p),
    .din1(G2_p_spl_101),
    .din2(G28_p_spl_000)
  );


  FA
  g_g532_n
  (
    .dout(g532_n),
    .din1(G2_n_spl_101),
    .din2(G28_n_spl_000)
  );


  LA
  g_g533_p
  (
    .dout(g533_p),
    .din1(g518_n_spl_),
    .din2(g521_n_spl_)
  );


  FA
  g_g533_n
  (
    .dout(g533_n),
    .din1(g518_p_spl_),
    .din2(g521_p_spl_)
  );


  LA
  g_g534_p
  (
    .dout(g534_p),
    .din1(G3_p_spl_101),
    .din2(G27_p_spl_001)
  );


  FA
  g_g534_n
  (
    .dout(g534_n),
    .din1(G3_n_spl_101),
    .din2(G27_n_spl_001)
  );


  LA
  g_g535_p
  (
    .dout(g535_p),
    .din1(g512_n_spl_),
    .din2(g515_n_spl_)
  );


  FA
  g_g535_n
  (
    .dout(g535_n),
    .din1(g512_p_spl_),
    .din2(g515_p_spl_)
  );


  LA
  g_g536_p
  (
    .dout(g536_p),
    .din1(G4_p_spl_100),
    .din2(G26_p_spl_001)
  );


  FA
  g_g536_n
  (
    .dout(g536_n),
    .din1(G4_n_spl_100),
    .din2(G26_n_spl_001)
  );


  LA
  g_g537_p
  (
    .dout(g537_p),
    .din1(g506_n_spl_),
    .din2(g509_n_spl_)
  );


  FA
  g_g537_n
  (
    .dout(g537_n),
    .din1(g506_p_spl_),
    .din2(g509_p_spl_)
  );


  LA
  g_g538_p
  (
    .dout(g538_p),
    .din1(G5_p_spl_100),
    .din2(G25_p_spl_010)
  );


  FA
  g_g538_n
  (
    .dout(g538_n),
    .din1(G5_n_spl_100),
    .din2(G25_n_spl_010)
  );


  LA
  g_g539_p
  (
    .dout(g539_p),
    .din1(g500_n_spl_),
    .din2(g503_n_spl_)
  );


  FA
  g_g539_n
  (
    .dout(g539_n),
    .din1(g500_p_spl_),
    .din2(g503_p_spl_)
  );


  LA
  g_g540_p
  (
    .dout(g540_p),
    .din1(G6_p_spl_011),
    .din2(G24_p_spl_010)
  );


  FA
  g_g540_n
  (
    .dout(g540_n),
    .din1(G6_n_spl_011),
    .din2(G24_n_spl_010)
  );


  LA
  g_g541_p
  (
    .dout(g541_p),
    .din1(g494_n_spl_),
    .din2(g497_n_spl_)
  );


  FA
  g_g541_n
  (
    .dout(g541_n),
    .din1(g494_p_spl_),
    .din2(g497_p_spl_)
  );


  LA
  g_g542_p
  (
    .dout(g542_p),
    .din1(G7_p_spl_011),
    .din2(G23_p_spl_011)
  );


  FA
  g_g542_n
  (
    .dout(g542_n),
    .din1(G7_n_spl_011),
    .din2(G23_n_spl_011)
  );


  LA
  g_g543_p
  (
    .dout(g543_p),
    .din1(g488_n_spl_),
    .din2(g491_n_spl_)
  );


  FA
  g_g543_n
  (
    .dout(g543_n),
    .din1(g488_p_spl_),
    .din2(g491_p_spl_)
  );


  LA
  g_g544_p
  (
    .dout(g544_p),
    .din1(G8_p_spl_010),
    .din2(G22_p_spl_011)
  );


  FA
  g_g544_n
  (
    .dout(g544_n),
    .din1(G8_n_spl_010),
    .din2(G22_n_spl_011)
  );


  LA
  g_g545_p
  (
    .dout(g545_p),
    .din1(g482_n_spl_),
    .din2(g485_n_spl_)
  );


  FA
  g_g545_n
  (
    .dout(g545_n),
    .din1(g482_p_spl_),
    .din2(g485_p_spl_)
  );


  LA
  g_g546_p
  (
    .dout(g546_p),
    .din1(G9_p_spl_010),
    .din2(G21_p_spl_100)
  );


  FA
  g_g546_n
  (
    .dout(g546_n),
    .din1(G9_n_spl_010),
    .din2(G21_n_spl_100)
  );


  LA
  g_g547_p
  (
    .dout(g547_p),
    .din1(g476_n_spl_),
    .din2(g479_n_spl_)
  );


  FA
  g_g547_n
  (
    .dout(g547_n),
    .din1(g476_p_spl_),
    .din2(g479_p_spl_)
  );


  LA
  g_g548_p
  (
    .dout(g548_p),
    .din1(G10_p_spl_001),
    .din2(G20_p_spl_100)
  );


  FA
  g_g548_n
  (
    .dout(g548_n),
    .din1(G10_n_spl_001),
    .din2(G20_n_spl_100)
  );


  LA
  g_g549_p
  (
    .dout(g549_p),
    .din1(g470_n_spl_),
    .din2(g473_n_spl_)
  );


  FA
  g_g549_n
  (
    .dout(g549_n),
    .din1(g470_p_spl_),
    .din2(g473_p_spl_)
  );


  LA
  g_g550_p
  (
    .dout(g550_p),
    .din1(G11_p_spl_001),
    .din2(G19_p_spl_101)
  );


  FA
  g_g550_n
  (
    .dout(g550_n),
    .din1(G11_n_spl_001),
    .din2(G19_n_spl_101)
  );


  LA
  g_g551_p
  (
    .dout(g551_p),
    .din1(G13_p_spl_000),
    .din2(G17_p_spl_110)
  );


  FA
  g_g551_n
  (
    .dout(g551_n),
    .din1(G13_n_spl_000),
    .din2(G17_n_spl_101)
  );


  LA
  g_g552_p
  (
    .dout(g552_p),
    .din1(G12_p_spl_000),
    .din2(G18_p_spl_101)
  );


  FA
  g_g552_n
  (
    .dout(g552_n),
    .din1(G12_n_spl_000),
    .din2(G18_n_spl_101)
  );


  LA
  g_g553_p
  (
    .dout(g553_p),
    .din1(g551_p_spl_),
    .din2(g552_n_spl_)
  );


  FA
  g_g553_n
  (
    .dout(g553_n),
    .din1(g551_n_spl_),
    .din2(g552_p_spl_)
  );


  LA
  g_g554_p
  (
    .dout(g554_p),
    .din1(g551_p_spl_),
    .din2(g553_n_spl_)
  );


  FA
  g_g554_n
  (
    .dout(g554_n),
    .din1(g551_n_spl_),
    .din2(g553_p_spl_)
  );


  LA
  g_g555_p
  (
    .dout(g555_p),
    .din1(g552_n_spl_),
    .din2(g553_n_spl_)
  );


  FA
  g_g555_n
  (
    .dout(g555_n),
    .din1(g552_p_spl_),
    .din2(g553_p_spl_)
  );


  LA
  g_g556_p
  (
    .dout(g556_p),
    .din1(g554_n_spl_0),
    .din2(g555_n)
  );


  FA
  g_g556_n
  (
    .dout(g556_n),
    .din1(g554_p_spl_0),
    .din2(g555_p)
  );


  LA
  g_g557_p
  (
    .dout(g557_p),
    .din1(g467_n_spl_0),
    .din2(g556_n_spl_)
  );


  FA
  g_g557_n
  (
    .dout(g557_n),
    .din1(g467_p_spl_0),
    .din2(g556_p_spl_)
  );


  LA
  g_g558_p
  (
    .dout(g558_p),
    .din1(g467_p_spl_),
    .din2(g556_p_spl_)
  );


  FA
  g_g558_n
  (
    .dout(g558_n),
    .din1(g467_n_spl_),
    .din2(g556_n_spl_)
  );


  LA
  g_g559_p
  (
    .dout(g559_p),
    .din1(g557_n_spl_),
    .din2(g558_n)
  );


  FA
  g_g559_n
  (
    .dout(g559_n),
    .din1(g557_p_spl_),
    .din2(g558_p)
  );


  LA
  g_g560_p
  (
    .dout(g560_p),
    .din1(g550_n_spl_),
    .din2(g559_p_spl_)
  );


  FA
  g_g560_n
  (
    .dout(g560_n),
    .din1(g550_p_spl_),
    .din2(g559_n_spl_)
  );


  LA
  g_g561_p
  (
    .dout(g561_p),
    .din1(g550_p_spl_),
    .din2(g559_n_spl_)
  );


  FA
  g_g561_n
  (
    .dout(g561_n),
    .din1(g550_n_spl_),
    .din2(g559_p_spl_)
  );


  LA
  g_g562_p
  (
    .dout(g562_p),
    .din1(g560_n_spl_),
    .din2(g561_n)
  );


  FA
  g_g562_n
  (
    .dout(g562_n),
    .din1(g560_p_spl_),
    .din2(g561_p)
  );


  LA
  g_g563_p
  (
    .dout(g563_p),
    .din1(g549_n_spl_),
    .din2(g562_p_spl_)
  );


  FA
  g_g563_n
  (
    .dout(g563_n),
    .din1(g549_p_spl_),
    .din2(g562_n_spl_)
  );


  LA
  g_g564_p
  (
    .dout(g564_p),
    .din1(g549_p_spl_),
    .din2(g562_n_spl_)
  );


  FA
  g_g564_n
  (
    .dout(g564_n),
    .din1(g549_n_spl_),
    .din2(g562_p_spl_)
  );


  LA
  g_g565_p
  (
    .dout(g565_p),
    .din1(g563_n_spl_),
    .din2(g564_n)
  );


  FA
  g_g565_n
  (
    .dout(g565_n),
    .din1(g563_p_spl_),
    .din2(g564_p)
  );


  LA
  g_g566_p
  (
    .dout(g566_p),
    .din1(g548_n_spl_),
    .din2(g565_p_spl_)
  );


  FA
  g_g566_n
  (
    .dout(g566_n),
    .din1(g548_p_spl_),
    .din2(g565_n_spl_)
  );


  LA
  g_g567_p
  (
    .dout(g567_p),
    .din1(g548_p_spl_),
    .din2(g565_n_spl_)
  );


  FA
  g_g567_n
  (
    .dout(g567_n),
    .din1(g548_n_spl_),
    .din2(g565_p_spl_)
  );


  LA
  g_g568_p
  (
    .dout(g568_p),
    .din1(g566_n_spl_),
    .din2(g567_n)
  );


  FA
  g_g568_n
  (
    .dout(g568_n),
    .din1(g566_p_spl_),
    .din2(g567_p)
  );


  LA
  g_g569_p
  (
    .dout(g569_p),
    .din1(g547_n_spl_),
    .din2(g568_p_spl_)
  );


  FA
  g_g569_n
  (
    .dout(g569_n),
    .din1(g547_p_spl_),
    .din2(g568_n_spl_)
  );


  LA
  g_g570_p
  (
    .dout(g570_p),
    .din1(g547_p_spl_),
    .din2(g568_n_spl_)
  );


  FA
  g_g570_n
  (
    .dout(g570_n),
    .din1(g547_n_spl_),
    .din2(g568_p_spl_)
  );


  LA
  g_g571_p
  (
    .dout(g571_p),
    .din1(g569_n_spl_),
    .din2(g570_n)
  );


  FA
  g_g571_n
  (
    .dout(g571_n),
    .din1(g569_p_spl_),
    .din2(g570_p)
  );


  LA
  g_g572_p
  (
    .dout(g572_p),
    .din1(g546_n_spl_),
    .din2(g571_p_spl_)
  );


  FA
  g_g572_n
  (
    .dout(g572_n),
    .din1(g546_p_spl_),
    .din2(g571_n_spl_)
  );


  LA
  g_g573_p
  (
    .dout(g573_p),
    .din1(g546_p_spl_),
    .din2(g571_n_spl_)
  );


  FA
  g_g573_n
  (
    .dout(g573_n),
    .din1(g546_n_spl_),
    .din2(g571_p_spl_)
  );


  LA
  g_g574_p
  (
    .dout(g574_p),
    .din1(g572_n_spl_),
    .din2(g573_n)
  );


  FA
  g_g574_n
  (
    .dout(g574_n),
    .din1(g572_p_spl_),
    .din2(g573_p)
  );


  LA
  g_g575_p
  (
    .dout(g575_p),
    .din1(g545_n_spl_),
    .din2(g574_p_spl_)
  );


  FA
  g_g575_n
  (
    .dout(g575_n),
    .din1(g545_p_spl_),
    .din2(g574_n_spl_)
  );


  LA
  g_g576_p
  (
    .dout(g576_p),
    .din1(g545_p_spl_),
    .din2(g574_n_spl_)
  );


  FA
  g_g576_n
  (
    .dout(g576_n),
    .din1(g545_n_spl_),
    .din2(g574_p_spl_)
  );


  LA
  g_g577_p
  (
    .dout(g577_p),
    .din1(g575_n_spl_),
    .din2(g576_n)
  );


  FA
  g_g577_n
  (
    .dout(g577_n),
    .din1(g575_p_spl_),
    .din2(g576_p)
  );


  LA
  g_g578_p
  (
    .dout(g578_p),
    .din1(g544_n_spl_),
    .din2(g577_p_spl_)
  );


  FA
  g_g578_n
  (
    .dout(g578_n),
    .din1(g544_p_spl_),
    .din2(g577_n_spl_)
  );


  LA
  g_g579_p
  (
    .dout(g579_p),
    .din1(g544_p_spl_),
    .din2(g577_n_spl_)
  );


  FA
  g_g579_n
  (
    .dout(g579_n),
    .din1(g544_n_spl_),
    .din2(g577_p_spl_)
  );


  LA
  g_g580_p
  (
    .dout(g580_p),
    .din1(g578_n_spl_),
    .din2(g579_n)
  );


  FA
  g_g580_n
  (
    .dout(g580_n),
    .din1(g578_p_spl_),
    .din2(g579_p)
  );


  LA
  g_g581_p
  (
    .dout(g581_p),
    .din1(g543_n_spl_),
    .din2(g580_p_spl_)
  );


  FA
  g_g581_n
  (
    .dout(g581_n),
    .din1(g543_p_spl_),
    .din2(g580_n_spl_)
  );


  LA
  g_g582_p
  (
    .dout(g582_p),
    .din1(g543_p_spl_),
    .din2(g580_n_spl_)
  );


  FA
  g_g582_n
  (
    .dout(g582_n),
    .din1(g543_n_spl_),
    .din2(g580_p_spl_)
  );


  LA
  g_g583_p
  (
    .dout(g583_p),
    .din1(g581_n_spl_),
    .din2(g582_n)
  );


  FA
  g_g583_n
  (
    .dout(g583_n),
    .din1(g581_p_spl_),
    .din2(g582_p)
  );


  LA
  g_g584_p
  (
    .dout(g584_p),
    .din1(g542_n_spl_),
    .din2(g583_p_spl_)
  );


  FA
  g_g584_n
  (
    .dout(g584_n),
    .din1(g542_p_spl_),
    .din2(g583_n_spl_)
  );


  LA
  g_g585_p
  (
    .dout(g585_p),
    .din1(g542_p_spl_),
    .din2(g583_n_spl_)
  );


  FA
  g_g585_n
  (
    .dout(g585_n),
    .din1(g542_n_spl_),
    .din2(g583_p_spl_)
  );


  LA
  g_g586_p
  (
    .dout(g586_p),
    .din1(g584_n_spl_),
    .din2(g585_n)
  );


  FA
  g_g586_n
  (
    .dout(g586_n),
    .din1(g584_p_spl_),
    .din2(g585_p)
  );


  LA
  g_g587_p
  (
    .dout(g587_p),
    .din1(g541_n_spl_),
    .din2(g586_p_spl_)
  );


  FA
  g_g587_n
  (
    .dout(g587_n),
    .din1(g541_p_spl_),
    .din2(g586_n_spl_)
  );


  LA
  g_g588_p
  (
    .dout(g588_p),
    .din1(g541_p_spl_),
    .din2(g586_n_spl_)
  );


  FA
  g_g588_n
  (
    .dout(g588_n),
    .din1(g541_n_spl_),
    .din2(g586_p_spl_)
  );


  LA
  g_g589_p
  (
    .dout(g589_p),
    .din1(g587_n_spl_),
    .din2(g588_n)
  );


  FA
  g_g589_n
  (
    .dout(g589_n),
    .din1(g587_p_spl_),
    .din2(g588_p)
  );


  LA
  g_g590_p
  (
    .dout(g590_p),
    .din1(g540_n_spl_),
    .din2(g589_p_spl_)
  );


  FA
  g_g590_n
  (
    .dout(g590_n),
    .din1(g540_p_spl_),
    .din2(g589_n_spl_)
  );


  LA
  g_g591_p
  (
    .dout(g591_p),
    .din1(g540_p_spl_),
    .din2(g589_n_spl_)
  );


  FA
  g_g591_n
  (
    .dout(g591_n),
    .din1(g540_n_spl_),
    .din2(g589_p_spl_)
  );


  LA
  g_g592_p
  (
    .dout(g592_p),
    .din1(g590_n_spl_),
    .din2(g591_n)
  );


  FA
  g_g592_n
  (
    .dout(g592_n),
    .din1(g590_p_spl_),
    .din2(g591_p)
  );


  LA
  g_g593_p
  (
    .dout(g593_p),
    .din1(g539_n_spl_),
    .din2(g592_p_spl_)
  );


  FA
  g_g593_n
  (
    .dout(g593_n),
    .din1(g539_p_spl_),
    .din2(g592_n_spl_)
  );


  LA
  g_g594_p
  (
    .dout(g594_p),
    .din1(g539_p_spl_),
    .din2(g592_n_spl_)
  );


  FA
  g_g594_n
  (
    .dout(g594_n),
    .din1(g539_n_spl_),
    .din2(g592_p_spl_)
  );


  LA
  g_g595_p
  (
    .dout(g595_p),
    .din1(g593_n_spl_),
    .din2(g594_n)
  );


  FA
  g_g595_n
  (
    .dout(g595_n),
    .din1(g593_p_spl_),
    .din2(g594_p)
  );


  LA
  g_g596_p
  (
    .dout(g596_p),
    .din1(g538_n_spl_),
    .din2(g595_p_spl_)
  );


  FA
  g_g596_n
  (
    .dout(g596_n),
    .din1(g538_p_spl_),
    .din2(g595_n_spl_)
  );


  LA
  g_g597_p
  (
    .dout(g597_p),
    .din1(g538_p_spl_),
    .din2(g595_n_spl_)
  );


  FA
  g_g597_n
  (
    .dout(g597_n),
    .din1(g538_n_spl_),
    .din2(g595_p_spl_)
  );


  LA
  g_g598_p
  (
    .dout(g598_p),
    .din1(g596_n_spl_),
    .din2(g597_n)
  );


  FA
  g_g598_n
  (
    .dout(g598_n),
    .din1(g596_p_spl_),
    .din2(g597_p)
  );


  LA
  g_g599_p
  (
    .dout(g599_p),
    .din1(g537_n_spl_),
    .din2(g598_p_spl_)
  );


  FA
  g_g599_n
  (
    .dout(g599_n),
    .din1(g537_p_spl_),
    .din2(g598_n_spl_)
  );


  LA
  g_g600_p
  (
    .dout(g600_p),
    .din1(g537_p_spl_),
    .din2(g598_n_spl_)
  );


  FA
  g_g600_n
  (
    .dout(g600_n),
    .din1(g537_n_spl_),
    .din2(g598_p_spl_)
  );


  LA
  g_g601_p
  (
    .dout(g601_p),
    .din1(g599_n_spl_),
    .din2(g600_n)
  );


  FA
  g_g601_n
  (
    .dout(g601_n),
    .din1(g599_p_spl_),
    .din2(g600_p)
  );


  LA
  g_g602_p
  (
    .dout(g602_p),
    .din1(g536_n_spl_),
    .din2(g601_p_spl_)
  );


  FA
  g_g602_n
  (
    .dout(g602_n),
    .din1(g536_p_spl_),
    .din2(g601_n_spl_)
  );


  LA
  g_g603_p
  (
    .dout(g603_p),
    .din1(g536_p_spl_),
    .din2(g601_n_spl_)
  );


  FA
  g_g603_n
  (
    .dout(g603_n),
    .din1(g536_n_spl_),
    .din2(g601_p_spl_)
  );


  LA
  g_g604_p
  (
    .dout(g604_p),
    .din1(g602_n_spl_),
    .din2(g603_n)
  );


  FA
  g_g604_n
  (
    .dout(g604_n),
    .din1(g602_p_spl_),
    .din2(g603_p)
  );


  LA
  g_g605_p
  (
    .dout(g605_p),
    .din1(g535_n_spl_),
    .din2(g604_p_spl_)
  );


  FA
  g_g605_n
  (
    .dout(g605_n),
    .din1(g535_p_spl_),
    .din2(g604_n_spl_)
  );


  LA
  g_g606_p
  (
    .dout(g606_p),
    .din1(g535_p_spl_),
    .din2(g604_n_spl_)
  );


  FA
  g_g606_n
  (
    .dout(g606_n),
    .din1(g535_n_spl_),
    .din2(g604_p_spl_)
  );


  LA
  g_g607_p
  (
    .dout(g607_p),
    .din1(g605_n_spl_),
    .din2(g606_n)
  );


  FA
  g_g607_n
  (
    .dout(g607_n),
    .din1(g605_p_spl_),
    .din2(g606_p)
  );


  LA
  g_g608_p
  (
    .dout(g608_p),
    .din1(g534_n_spl_),
    .din2(g607_p_spl_)
  );


  FA
  g_g608_n
  (
    .dout(g608_n),
    .din1(g534_p_spl_),
    .din2(g607_n_spl_)
  );


  LA
  g_g609_p
  (
    .dout(g609_p),
    .din1(g534_p_spl_),
    .din2(g607_n_spl_)
  );


  FA
  g_g609_n
  (
    .dout(g609_n),
    .din1(g534_n_spl_),
    .din2(g607_p_spl_)
  );


  LA
  g_g610_p
  (
    .dout(g610_p),
    .din1(g608_n_spl_),
    .din2(g609_n)
  );


  FA
  g_g610_n
  (
    .dout(g610_n),
    .din1(g608_p_spl_),
    .din2(g609_p)
  );


  LA
  g_g611_p
  (
    .dout(g611_p),
    .din1(g533_n_spl_),
    .din2(g610_p_spl_)
  );


  FA
  g_g611_n
  (
    .dout(g611_n),
    .din1(g533_p_spl_),
    .din2(g610_n_spl_)
  );


  LA
  g_g612_p
  (
    .dout(g612_p),
    .din1(g533_p_spl_),
    .din2(g610_n_spl_)
  );


  FA
  g_g612_n
  (
    .dout(g612_n),
    .din1(g533_n_spl_),
    .din2(g610_p_spl_)
  );


  LA
  g_g613_p
  (
    .dout(g613_p),
    .din1(g611_n_spl_),
    .din2(g612_n)
  );


  FA
  g_g613_n
  (
    .dout(g613_n),
    .din1(g611_p_spl_),
    .din2(g612_p)
  );


  LA
  g_g614_p
  (
    .dout(g614_p),
    .din1(g532_n_spl_),
    .din2(g613_p_spl_)
  );


  FA
  g_g614_n
  (
    .dout(g614_n),
    .din1(g532_p_spl_),
    .din2(g613_n_spl_)
  );


  LA
  g_g615_p
  (
    .dout(g615_p),
    .din1(g532_p_spl_),
    .din2(g613_n_spl_)
  );


  FA
  g_g615_n
  (
    .dout(g615_n),
    .din1(g532_n_spl_),
    .din2(g613_p_spl_)
  );


  LA
  g_g616_p
  (
    .dout(g616_p),
    .din1(g614_n_spl_),
    .din2(g615_n)
  );


  FA
  g_g616_n
  (
    .dout(g616_n),
    .din1(g614_p_spl_),
    .din2(g615_p)
  );


  LA
  g_g617_p
  (
    .dout(g617_p),
    .din1(g531_n_spl_),
    .din2(g616_p_spl_)
  );


  FA
  g_g617_n
  (
    .dout(g617_n),
    .din1(g531_p_spl_),
    .din2(g616_n_spl_)
  );


  LA
  g_g618_p
  (
    .dout(g618_p),
    .din1(g531_p_spl_),
    .din2(g616_n_spl_)
  );


  FA
  g_g618_n
  (
    .dout(g618_n),
    .din1(g531_n_spl_),
    .din2(g616_p_spl_)
  );


  LA
  g_g619_p
  (
    .dout(g619_p),
    .din1(g617_n_spl_),
    .din2(g618_n)
  );


  FA
  g_g619_n
  (
    .dout(g619_n),
    .din1(g617_p_spl_),
    .din2(g618_p)
  );


  LA
  g_g620_p
  (
    .dout(g620_p),
    .din1(g530_n),
    .din2(g619_p)
  );


  FA
  g_g620_n
  (
    .dout(g620_n),
    .din1(g530_p_spl_),
    .din2(g619_n_spl_)
  );


  LA
  g_g621_p
  (
    .dout(g621_p),
    .din1(g530_p_spl_),
    .din2(g619_n_spl_)
  );


  FA
  g_g622_n
  (
    .dout(g622_n),
    .din1(g620_p_spl_),
    .din2(g621_p)
  );


  LA
  g_g623_p
  (
    .dout(g623_p),
    .din1(G1_p_spl_110),
    .din2(G30_p_spl_000)
  );


  FA
  g_g623_n
  (
    .dout(g623_n),
    .din1(G1_n_spl_110),
    .din2(G30_n_spl_000)
  );


  LA
  g_g624_p
  (
    .dout(g624_p),
    .din1(g617_n_spl_),
    .din2(g620_n)
  );


  FA
  g_g624_n
  (
    .dout(g624_n),
    .din1(g617_p_spl_),
    .din2(g620_p_spl_)
  );


  LA
  g_g625_p
  (
    .dout(g625_p),
    .din1(G2_p_spl_110),
    .din2(G29_p_spl_000)
  );


  FA
  g_g625_n
  (
    .dout(g625_n),
    .din1(G2_n_spl_110),
    .din2(G29_n_spl_000)
  );


  LA
  g_g626_p
  (
    .dout(g626_p),
    .din1(g611_n_spl_),
    .din2(g614_n_spl_)
  );


  FA
  g_g626_n
  (
    .dout(g626_n),
    .din1(g611_p_spl_),
    .din2(g614_p_spl_)
  );


  LA
  g_g627_p
  (
    .dout(g627_p),
    .din1(G3_p_spl_101),
    .din2(G28_p_spl_001)
  );


  FA
  g_g627_n
  (
    .dout(g627_n),
    .din1(G3_n_spl_101),
    .din2(G28_n_spl_001)
  );


  LA
  g_g628_p
  (
    .dout(g628_p),
    .din1(g605_n_spl_),
    .din2(g608_n_spl_)
  );


  FA
  g_g628_n
  (
    .dout(g628_n),
    .din1(g605_p_spl_),
    .din2(g608_p_spl_)
  );


  LA
  g_g629_p
  (
    .dout(g629_p),
    .din1(G4_p_spl_101),
    .din2(G27_p_spl_001)
  );


  FA
  g_g629_n
  (
    .dout(g629_n),
    .din1(G4_n_spl_101),
    .din2(G27_n_spl_001)
  );


  LA
  g_g630_p
  (
    .dout(g630_p),
    .din1(g599_n_spl_),
    .din2(g602_n_spl_)
  );


  FA
  g_g630_n
  (
    .dout(g630_n),
    .din1(g599_p_spl_),
    .din2(g602_p_spl_)
  );


  LA
  g_g631_p
  (
    .dout(g631_p),
    .din1(G5_p_spl_100),
    .din2(G26_p_spl_010)
  );


  FA
  g_g631_n
  (
    .dout(g631_n),
    .din1(G5_n_spl_100),
    .din2(G26_n_spl_010)
  );


  LA
  g_g632_p
  (
    .dout(g632_p),
    .din1(g593_n_spl_),
    .din2(g596_n_spl_)
  );


  FA
  g_g632_n
  (
    .dout(g632_n),
    .din1(g593_p_spl_),
    .din2(g596_p_spl_)
  );


  LA
  g_g633_p
  (
    .dout(g633_p),
    .din1(G6_p_spl_100),
    .din2(G25_p_spl_010)
  );


  FA
  g_g633_n
  (
    .dout(g633_n),
    .din1(G6_n_spl_100),
    .din2(G25_n_spl_010)
  );


  LA
  g_g634_p
  (
    .dout(g634_p),
    .din1(g587_n_spl_),
    .din2(g590_n_spl_)
  );


  FA
  g_g634_n
  (
    .dout(g634_n),
    .din1(g587_p_spl_),
    .din2(g590_p_spl_)
  );


  LA
  g_g635_p
  (
    .dout(g635_p),
    .din1(G7_p_spl_011),
    .din2(G24_p_spl_011)
  );


  FA
  g_g635_n
  (
    .dout(g635_n),
    .din1(G7_n_spl_011),
    .din2(G24_n_spl_011)
  );


  LA
  g_g636_p
  (
    .dout(g636_p),
    .din1(g581_n_spl_),
    .din2(g584_n_spl_)
  );


  FA
  g_g636_n
  (
    .dout(g636_n),
    .din1(g581_p_spl_),
    .din2(g584_p_spl_)
  );


  LA
  g_g637_p
  (
    .dout(g637_p),
    .din1(G8_p_spl_011),
    .din2(G23_p_spl_011)
  );


  FA
  g_g637_n
  (
    .dout(g637_n),
    .din1(G8_n_spl_011),
    .din2(G23_n_spl_011)
  );


  LA
  g_g638_p
  (
    .dout(g638_p),
    .din1(g575_n_spl_),
    .din2(g578_n_spl_)
  );


  FA
  g_g638_n
  (
    .dout(g638_n),
    .din1(g575_p_spl_),
    .din2(g578_p_spl_)
  );


  LA
  g_g639_p
  (
    .dout(g639_p),
    .din1(G9_p_spl_010),
    .din2(G22_p_spl_100)
  );


  FA
  g_g639_n
  (
    .dout(g639_n),
    .din1(G9_n_spl_010),
    .din2(G22_n_spl_100)
  );


  LA
  g_g640_p
  (
    .dout(g640_p),
    .din1(g569_n_spl_),
    .din2(g572_n_spl_)
  );


  FA
  g_g640_n
  (
    .dout(g640_n),
    .din1(g569_p_spl_),
    .din2(g572_p_spl_)
  );


  LA
  g_g641_p
  (
    .dout(g641_p),
    .din1(G10_p_spl_010),
    .din2(G21_p_spl_100)
  );


  FA
  g_g641_n
  (
    .dout(g641_n),
    .din1(G10_n_spl_010),
    .din2(G21_n_spl_100)
  );


  LA
  g_g642_p
  (
    .dout(g642_p),
    .din1(g563_n_spl_),
    .din2(g566_n_spl_)
  );


  FA
  g_g642_n
  (
    .dout(g642_n),
    .din1(g563_p_spl_),
    .din2(g566_p_spl_)
  );


  LA
  g_g643_p
  (
    .dout(g643_p),
    .din1(G11_p_spl_001),
    .din2(G20_p_spl_101)
  );


  FA
  g_g643_n
  (
    .dout(g643_n),
    .din1(G11_n_spl_001),
    .din2(G20_n_spl_101)
  );


  LA
  g_g644_p
  (
    .dout(g644_p),
    .din1(g557_n_spl_),
    .din2(g560_n_spl_)
  );


  FA
  g_g644_n
  (
    .dout(g644_n),
    .din1(g557_p_spl_),
    .din2(g560_p_spl_)
  );


  LA
  g_g645_p
  (
    .dout(g645_p),
    .din1(G12_p_spl_001),
    .din2(G19_p_spl_101)
  );


  FA
  g_g645_n
  (
    .dout(g645_n),
    .din1(G12_n_spl_001),
    .din2(G19_n_spl_101)
  );


  LA
  g_g646_p
  (
    .dout(g646_p),
    .din1(G14_p_spl_000),
    .din2(G17_p_spl_110)
  );


  FA
  g_g646_n
  (
    .dout(g646_n),
    .din1(G14_n_spl_000),
    .din2(G17_n_spl_110)
  );


  LA
  g_g647_p
  (
    .dout(g647_p),
    .din1(G13_p_spl_000),
    .din2(G18_p_spl_110)
  );


  FA
  g_g647_n
  (
    .dout(g647_n),
    .din1(G13_n_spl_000),
    .din2(G18_n_spl_110)
  );


  LA
  g_g648_p
  (
    .dout(g648_p),
    .din1(g646_p_spl_),
    .din2(g647_n_spl_)
  );


  FA
  g_g648_n
  (
    .dout(g648_n),
    .din1(g646_n_spl_),
    .din2(g647_p_spl_)
  );


  LA
  g_g649_p
  (
    .dout(g649_p),
    .din1(g646_p_spl_),
    .din2(g648_n_spl_)
  );


  FA
  g_g649_n
  (
    .dout(g649_n),
    .din1(g646_n_spl_),
    .din2(g648_p_spl_)
  );


  LA
  g_g650_p
  (
    .dout(g650_p),
    .din1(g647_n_spl_),
    .din2(g648_n_spl_)
  );


  FA
  g_g650_n
  (
    .dout(g650_n),
    .din1(g647_p_spl_),
    .din2(g648_p_spl_)
  );


  LA
  g_g651_p
  (
    .dout(g651_p),
    .din1(g649_n_spl_0),
    .din2(g650_n)
  );


  FA
  g_g651_n
  (
    .dout(g651_n),
    .din1(g649_p_spl_0),
    .din2(g650_p)
  );


  LA
  g_g652_p
  (
    .dout(g652_p),
    .din1(g554_n_spl_0),
    .din2(g651_n_spl_)
  );


  FA
  g_g652_n
  (
    .dout(g652_n),
    .din1(g554_p_spl_0),
    .din2(g651_p_spl_)
  );


  LA
  g_g653_p
  (
    .dout(g653_p),
    .din1(g554_p_spl_),
    .din2(g651_p_spl_)
  );


  FA
  g_g653_n
  (
    .dout(g653_n),
    .din1(g554_n_spl_),
    .din2(g651_n_spl_)
  );


  LA
  g_g654_p
  (
    .dout(g654_p),
    .din1(g652_n_spl_),
    .din2(g653_n)
  );


  FA
  g_g654_n
  (
    .dout(g654_n),
    .din1(g652_p_spl_),
    .din2(g653_p)
  );


  LA
  g_g655_p
  (
    .dout(g655_p),
    .din1(g645_n_spl_),
    .din2(g654_p_spl_)
  );


  FA
  g_g655_n
  (
    .dout(g655_n),
    .din1(g645_p_spl_),
    .din2(g654_n_spl_)
  );


  LA
  g_g656_p
  (
    .dout(g656_p),
    .din1(g645_p_spl_),
    .din2(g654_n_spl_)
  );


  FA
  g_g656_n
  (
    .dout(g656_n),
    .din1(g645_n_spl_),
    .din2(g654_p_spl_)
  );


  LA
  g_g657_p
  (
    .dout(g657_p),
    .din1(g655_n_spl_),
    .din2(g656_n)
  );


  FA
  g_g657_n
  (
    .dout(g657_n),
    .din1(g655_p_spl_),
    .din2(g656_p)
  );


  LA
  g_g658_p
  (
    .dout(g658_p),
    .din1(g644_n_spl_),
    .din2(g657_p_spl_)
  );


  FA
  g_g658_n
  (
    .dout(g658_n),
    .din1(g644_p_spl_),
    .din2(g657_n_spl_)
  );


  LA
  g_g659_p
  (
    .dout(g659_p),
    .din1(g644_p_spl_),
    .din2(g657_n_spl_)
  );


  FA
  g_g659_n
  (
    .dout(g659_n),
    .din1(g644_n_spl_),
    .din2(g657_p_spl_)
  );


  LA
  g_g660_p
  (
    .dout(g660_p),
    .din1(g658_n_spl_),
    .din2(g659_n)
  );


  FA
  g_g660_n
  (
    .dout(g660_n),
    .din1(g658_p_spl_),
    .din2(g659_p)
  );


  LA
  g_g661_p
  (
    .dout(g661_p),
    .din1(g643_n_spl_),
    .din2(g660_p_spl_)
  );


  FA
  g_g661_n
  (
    .dout(g661_n),
    .din1(g643_p_spl_),
    .din2(g660_n_spl_)
  );


  LA
  g_g662_p
  (
    .dout(g662_p),
    .din1(g643_p_spl_),
    .din2(g660_n_spl_)
  );


  FA
  g_g662_n
  (
    .dout(g662_n),
    .din1(g643_n_spl_),
    .din2(g660_p_spl_)
  );


  LA
  g_g663_p
  (
    .dout(g663_p),
    .din1(g661_n_spl_),
    .din2(g662_n)
  );


  FA
  g_g663_n
  (
    .dout(g663_n),
    .din1(g661_p_spl_),
    .din2(g662_p)
  );


  LA
  g_g664_p
  (
    .dout(g664_p),
    .din1(g642_n_spl_),
    .din2(g663_p_spl_)
  );


  FA
  g_g664_n
  (
    .dout(g664_n),
    .din1(g642_p_spl_),
    .din2(g663_n_spl_)
  );


  LA
  g_g665_p
  (
    .dout(g665_p),
    .din1(g642_p_spl_),
    .din2(g663_n_spl_)
  );


  FA
  g_g665_n
  (
    .dout(g665_n),
    .din1(g642_n_spl_),
    .din2(g663_p_spl_)
  );


  LA
  g_g666_p
  (
    .dout(g666_p),
    .din1(g664_n_spl_),
    .din2(g665_n)
  );


  FA
  g_g666_n
  (
    .dout(g666_n),
    .din1(g664_p_spl_),
    .din2(g665_p)
  );


  LA
  g_g667_p
  (
    .dout(g667_p),
    .din1(g641_n_spl_),
    .din2(g666_p_spl_)
  );


  FA
  g_g667_n
  (
    .dout(g667_n),
    .din1(g641_p_spl_),
    .din2(g666_n_spl_)
  );


  LA
  g_g668_p
  (
    .dout(g668_p),
    .din1(g641_p_spl_),
    .din2(g666_n_spl_)
  );


  FA
  g_g668_n
  (
    .dout(g668_n),
    .din1(g641_n_spl_),
    .din2(g666_p_spl_)
  );


  LA
  g_g669_p
  (
    .dout(g669_p),
    .din1(g667_n_spl_),
    .din2(g668_n)
  );


  FA
  g_g669_n
  (
    .dout(g669_n),
    .din1(g667_p_spl_),
    .din2(g668_p)
  );


  LA
  g_g670_p
  (
    .dout(g670_p),
    .din1(g640_n_spl_),
    .din2(g669_p_spl_)
  );


  FA
  g_g670_n
  (
    .dout(g670_n),
    .din1(g640_p_spl_),
    .din2(g669_n_spl_)
  );


  LA
  g_g671_p
  (
    .dout(g671_p),
    .din1(g640_p_spl_),
    .din2(g669_n_spl_)
  );


  FA
  g_g671_n
  (
    .dout(g671_n),
    .din1(g640_n_spl_),
    .din2(g669_p_spl_)
  );


  LA
  g_g672_p
  (
    .dout(g672_p),
    .din1(g670_n_spl_),
    .din2(g671_n)
  );


  FA
  g_g672_n
  (
    .dout(g672_n),
    .din1(g670_p_spl_),
    .din2(g671_p)
  );


  LA
  g_g673_p
  (
    .dout(g673_p),
    .din1(g639_n_spl_),
    .din2(g672_p_spl_)
  );


  FA
  g_g673_n
  (
    .dout(g673_n),
    .din1(g639_p_spl_),
    .din2(g672_n_spl_)
  );


  LA
  g_g674_p
  (
    .dout(g674_p),
    .din1(g639_p_spl_),
    .din2(g672_n_spl_)
  );


  FA
  g_g674_n
  (
    .dout(g674_n),
    .din1(g639_n_spl_),
    .din2(g672_p_spl_)
  );


  LA
  g_g675_p
  (
    .dout(g675_p),
    .din1(g673_n_spl_),
    .din2(g674_n)
  );


  FA
  g_g675_n
  (
    .dout(g675_n),
    .din1(g673_p_spl_),
    .din2(g674_p)
  );


  LA
  g_g676_p
  (
    .dout(g676_p),
    .din1(g638_n_spl_),
    .din2(g675_p_spl_)
  );


  FA
  g_g676_n
  (
    .dout(g676_n),
    .din1(g638_p_spl_),
    .din2(g675_n_spl_)
  );


  LA
  g_g677_p
  (
    .dout(g677_p),
    .din1(g638_p_spl_),
    .din2(g675_n_spl_)
  );


  FA
  g_g677_n
  (
    .dout(g677_n),
    .din1(g638_n_spl_),
    .din2(g675_p_spl_)
  );


  LA
  g_g678_p
  (
    .dout(g678_p),
    .din1(g676_n_spl_),
    .din2(g677_n)
  );


  FA
  g_g678_n
  (
    .dout(g678_n),
    .din1(g676_p_spl_),
    .din2(g677_p)
  );


  LA
  g_g679_p
  (
    .dout(g679_p),
    .din1(g637_n_spl_),
    .din2(g678_p_spl_)
  );


  FA
  g_g679_n
  (
    .dout(g679_n),
    .din1(g637_p_spl_),
    .din2(g678_n_spl_)
  );


  LA
  g_g680_p
  (
    .dout(g680_p),
    .din1(g637_p_spl_),
    .din2(g678_n_spl_)
  );


  FA
  g_g680_n
  (
    .dout(g680_n),
    .din1(g637_n_spl_),
    .din2(g678_p_spl_)
  );


  LA
  g_g681_p
  (
    .dout(g681_p),
    .din1(g679_n_spl_),
    .din2(g680_n)
  );


  FA
  g_g681_n
  (
    .dout(g681_n),
    .din1(g679_p_spl_),
    .din2(g680_p)
  );


  LA
  g_g682_p
  (
    .dout(g682_p),
    .din1(g636_n_spl_),
    .din2(g681_p_spl_)
  );


  FA
  g_g682_n
  (
    .dout(g682_n),
    .din1(g636_p_spl_),
    .din2(g681_n_spl_)
  );


  LA
  g_g683_p
  (
    .dout(g683_p),
    .din1(g636_p_spl_),
    .din2(g681_n_spl_)
  );


  FA
  g_g683_n
  (
    .dout(g683_n),
    .din1(g636_n_spl_),
    .din2(g681_p_spl_)
  );


  LA
  g_g684_p
  (
    .dout(g684_p),
    .din1(g682_n_spl_),
    .din2(g683_n)
  );


  FA
  g_g684_n
  (
    .dout(g684_n),
    .din1(g682_p_spl_),
    .din2(g683_p)
  );


  LA
  g_g685_p
  (
    .dout(g685_p),
    .din1(g635_n_spl_),
    .din2(g684_p_spl_)
  );


  FA
  g_g685_n
  (
    .dout(g685_n),
    .din1(g635_p_spl_),
    .din2(g684_n_spl_)
  );


  LA
  g_g686_p
  (
    .dout(g686_p),
    .din1(g635_p_spl_),
    .din2(g684_n_spl_)
  );


  FA
  g_g686_n
  (
    .dout(g686_n),
    .din1(g635_n_spl_),
    .din2(g684_p_spl_)
  );


  LA
  g_g687_p
  (
    .dout(g687_p),
    .din1(g685_n_spl_),
    .din2(g686_n)
  );


  FA
  g_g687_n
  (
    .dout(g687_n),
    .din1(g685_p_spl_),
    .din2(g686_p)
  );


  LA
  g_g688_p
  (
    .dout(g688_p),
    .din1(g634_n_spl_),
    .din2(g687_p_spl_)
  );


  FA
  g_g688_n
  (
    .dout(g688_n),
    .din1(g634_p_spl_),
    .din2(g687_n_spl_)
  );


  LA
  g_g689_p
  (
    .dout(g689_p),
    .din1(g634_p_spl_),
    .din2(g687_n_spl_)
  );


  FA
  g_g689_n
  (
    .dout(g689_n),
    .din1(g634_n_spl_),
    .din2(g687_p_spl_)
  );


  LA
  g_g690_p
  (
    .dout(g690_p),
    .din1(g688_n_spl_),
    .din2(g689_n)
  );


  FA
  g_g690_n
  (
    .dout(g690_n),
    .din1(g688_p_spl_),
    .din2(g689_p)
  );


  LA
  g_g691_p
  (
    .dout(g691_p),
    .din1(g633_n_spl_),
    .din2(g690_p_spl_)
  );


  FA
  g_g691_n
  (
    .dout(g691_n),
    .din1(g633_p_spl_),
    .din2(g690_n_spl_)
  );


  LA
  g_g692_p
  (
    .dout(g692_p),
    .din1(g633_p_spl_),
    .din2(g690_n_spl_)
  );


  FA
  g_g692_n
  (
    .dout(g692_n),
    .din1(g633_n_spl_),
    .din2(g690_p_spl_)
  );


  LA
  g_g693_p
  (
    .dout(g693_p),
    .din1(g691_n_spl_),
    .din2(g692_n)
  );


  FA
  g_g693_n
  (
    .dout(g693_n),
    .din1(g691_p_spl_),
    .din2(g692_p)
  );


  LA
  g_g694_p
  (
    .dout(g694_p),
    .din1(g632_n_spl_),
    .din2(g693_p_spl_)
  );


  FA
  g_g694_n
  (
    .dout(g694_n),
    .din1(g632_p_spl_),
    .din2(g693_n_spl_)
  );


  LA
  g_g695_p
  (
    .dout(g695_p),
    .din1(g632_p_spl_),
    .din2(g693_n_spl_)
  );


  FA
  g_g695_n
  (
    .dout(g695_n),
    .din1(g632_n_spl_),
    .din2(g693_p_spl_)
  );


  LA
  g_g696_p
  (
    .dout(g696_p),
    .din1(g694_n_spl_),
    .din2(g695_n)
  );


  FA
  g_g696_n
  (
    .dout(g696_n),
    .din1(g694_p_spl_),
    .din2(g695_p)
  );


  LA
  g_g697_p
  (
    .dout(g697_p),
    .din1(g631_n_spl_),
    .din2(g696_p_spl_)
  );


  FA
  g_g697_n
  (
    .dout(g697_n),
    .din1(g631_p_spl_),
    .din2(g696_n_spl_)
  );


  LA
  g_g698_p
  (
    .dout(g698_p),
    .din1(g631_p_spl_),
    .din2(g696_n_spl_)
  );


  FA
  g_g698_n
  (
    .dout(g698_n),
    .din1(g631_n_spl_),
    .din2(g696_p_spl_)
  );


  LA
  g_g699_p
  (
    .dout(g699_p),
    .din1(g697_n_spl_),
    .din2(g698_n)
  );


  FA
  g_g699_n
  (
    .dout(g699_n),
    .din1(g697_p_spl_),
    .din2(g698_p)
  );


  LA
  g_g700_p
  (
    .dout(g700_p),
    .din1(g630_n_spl_),
    .din2(g699_p_spl_)
  );


  FA
  g_g700_n
  (
    .dout(g700_n),
    .din1(g630_p_spl_),
    .din2(g699_n_spl_)
  );


  LA
  g_g701_p
  (
    .dout(g701_p),
    .din1(g630_p_spl_),
    .din2(g699_n_spl_)
  );


  FA
  g_g701_n
  (
    .dout(g701_n),
    .din1(g630_n_spl_),
    .din2(g699_p_spl_)
  );


  LA
  g_g702_p
  (
    .dout(g702_p),
    .din1(g700_n_spl_),
    .din2(g701_n)
  );


  FA
  g_g702_n
  (
    .dout(g702_n),
    .din1(g700_p_spl_),
    .din2(g701_p)
  );


  LA
  g_g703_p
  (
    .dout(g703_p),
    .din1(g629_n_spl_),
    .din2(g702_p_spl_)
  );


  FA
  g_g703_n
  (
    .dout(g703_n),
    .din1(g629_p_spl_),
    .din2(g702_n_spl_)
  );


  LA
  g_g704_p
  (
    .dout(g704_p),
    .din1(g629_p_spl_),
    .din2(g702_n_spl_)
  );


  FA
  g_g704_n
  (
    .dout(g704_n),
    .din1(g629_n_spl_),
    .din2(g702_p_spl_)
  );


  LA
  g_g705_p
  (
    .dout(g705_p),
    .din1(g703_n_spl_),
    .din2(g704_n)
  );


  FA
  g_g705_n
  (
    .dout(g705_n),
    .din1(g703_p_spl_),
    .din2(g704_p)
  );


  LA
  g_g706_p
  (
    .dout(g706_p),
    .din1(g628_n_spl_),
    .din2(g705_p_spl_)
  );


  FA
  g_g706_n
  (
    .dout(g706_n),
    .din1(g628_p_spl_),
    .din2(g705_n_spl_)
  );


  LA
  g_g707_p
  (
    .dout(g707_p),
    .din1(g628_p_spl_),
    .din2(g705_n_spl_)
  );


  FA
  g_g707_n
  (
    .dout(g707_n),
    .din1(g628_n_spl_),
    .din2(g705_p_spl_)
  );


  LA
  g_g708_p
  (
    .dout(g708_p),
    .din1(g706_n_spl_),
    .din2(g707_n)
  );


  FA
  g_g708_n
  (
    .dout(g708_n),
    .din1(g706_p_spl_),
    .din2(g707_p)
  );


  LA
  g_g709_p
  (
    .dout(g709_p),
    .din1(g627_n_spl_),
    .din2(g708_p_spl_)
  );


  FA
  g_g709_n
  (
    .dout(g709_n),
    .din1(g627_p_spl_),
    .din2(g708_n_spl_)
  );


  LA
  g_g710_p
  (
    .dout(g710_p),
    .din1(g627_p_spl_),
    .din2(g708_n_spl_)
  );


  FA
  g_g710_n
  (
    .dout(g710_n),
    .din1(g627_n_spl_),
    .din2(g708_p_spl_)
  );


  LA
  g_g711_p
  (
    .dout(g711_p),
    .din1(g709_n_spl_),
    .din2(g710_n)
  );


  FA
  g_g711_n
  (
    .dout(g711_n),
    .din1(g709_p_spl_),
    .din2(g710_p)
  );


  LA
  g_g712_p
  (
    .dout(g712_p),
    .din1(g626_n_spl_),
    .din2(g711_p_spl_)
  );


  FA
  g_g712_n
  (
    .dout(g712_n),
    .din1(g626_p_spl_),
    .din2(g711_n_spl_)
  );


  LA
  g_g713_p
  (
    .dout(g713_p),
    .din1(g626_p_spl_),
    .din2(g711_n_spl_)
  );


  FA
  g_g713_n
  (
    .dout(g713_n),
    .din1(g626_n_spl_),
    .din2(g711_p_spl_)
  );


  LA
  g_g714_p
  (
    .dout(g714_p),
    .din1(g712_n_spl_),
    .din2(g713_n)
  );


  FA
  g_g714_n
  (
    .dout(g714_n),
    .din1(g712_p_spl_),
    .din2(g713_p)
  );


  LA
  g_g715_p
  (
    .dout(g715_p),
    .din1(g625_n_spl_),
    .din2(g714_p_spl_)
  );


  FA
  g_g715_n
  (
    .dout(g715_n),
    .din1(g625_p_spl_),
    .din2(g714_n_spl_)
  );


  LA
  g_g716_p
  (
    .dout(g716_p),
    .din1(g625_p_spl_),
    .din2(g714_n_spl_)
  );


  FA
  g_g716_n
  (
    .dout(g716_n),
    .din1(g625_n_spl_),
    .din2(g714_p_spl_)
  );


  LA
  g_g717_p
  (
    .dout(g717_p),
    .din1(g715_n_spl_),
    .din2(g716_n)
  );


  FA
  g_g717_n
  (
    .dout(g717_n),
    .din1(g715_p_spl_),
    .din2(g716_p)
  );


  LA
  g_g718_p
  (
    .dout(g718_p),
    .din1(g624_n_spl_),
    .din2(g717_p_spl_)
  );


  FA
  g_g718_n
  (
    .dout(g718_n),
    .din1(g624_p_spl_),
    .din2(g717_n_spl_)
  );


  LA
  g_g719_p
  (
    .dout(g719_p),
    .din1(g624_p_spl_),
    .din2(g717_n_spl_)
  );


  FA
  g_g719_n
  (
    .dout(g719_n),
    .din1(g624_n_spl_),
    .din2(g717_p_spl_)
  );


  LA
  g_g720_p
  (
    .dout(g720_p),
    .din1(g718_n_spl_),
    .din2(g719_n)
  );


  FA
  g_g720_n
  (
    .dout(g720_n),
    .din1(g718_p_spl_),
    .din2(g719_p)
  );


  LA
  g_g721_p
  (
    .dout(g721_p),
    .din1(g623_n),
    .din2(g720_p)
  );


  FA
  g_g721_n
  (
    .dout(g721_n),
    .din1(g623_p_spl_),
    .din2(g720_n_spl_)
  );


  LA
  g_g722_p
  (
    .dout(g722_p),
    .din1(g623_p_spl_),
    .din2(g720_n_spl_)
  );


  FA
  g_g723_n
  (
    .dout(g723_n),
    .din1(g721_p_spl_),
    .din2(g722_p)
  );


  LA
  g_g724_p
  (
    .dout(g724_p),
    .din1(G1_p_spl_111),
    .din2(G31_p_spl_000)
  );


  FA
  g_g724_n
  (
    .dout(g724_n),
    .din1(G1_n_spl_110),
    .din2(G31_n_spl_000)
  );


  LA
  g_g725_p
  (
    .dout(g725_p),
    .din1(g718_n_spl_),
    .din2(g721_n)
  );


  FA
  g_g725_n
  (
    .dout(g725_n),
    .din1(g718_p_spl_),
    .din2(g721_p_spl_)
  );


  LA
  g_g726_p
  (
    .dout(g726_p),
    .din1(G2_p_spl_110),
    .din2(G30_p_spl_000)
  );


  FA
  g_g726_n
  (
    .dout(g726_n),
    .din1(G2_n_spl_110),
    .din2(G30_n_spl_000)
  );


  LA
  g_g727_p
  (
    .dout(g727_p),
    .din1(g712_n_spl_),
    .din2(g715_n_spl_)
  );


  FA
  g_g727_n
  (
    .dout(g727_n),
    .din1(g712_p_spl_),
    .din2(g715_p_spl_)
  );


  LA
  g_g728_p
  (
    .dout(g728_p),
    .din1(G3_p_spl_110),
    .din2(G29_p_spl_001)
  );


  FA
  g_g728_n
  (
    .dout(g728_n),
    .din1(G3_n_spl_110),
    .din2(G29_n_spl_001)
  );


  LA
  g_g729_p
  (
    .dout(g729_p),
    .din1(g706_n_spl_),
    .din2(g709_n_spl_)
  );


  FA
  g_g729_n
  (
    .dout(g729_n),
    .din1(g706_p_spl_),
    .din2(g709_p_spl_)
  );


  LA
  g_g730_p
  (
    .dout(g730_p),
    .din1(G4_p_spl_101),
    .din2(G28_p_spl_001)
  );


  FA
  g_g730_n
  (
    .dout(g730_n),
    .din1(G4_n_spl_101),
    .din2(G28_n_spl_001)
  );


  LA
  g_g731_p
  (
    .dout(g731_p),
    .din1(g700_n_spl_),
    .din2(g703_n_spl_)
  );


  FA
  g_g731_n
  (
    .dout(g731_n),
    .din1(g700_p_spl_),
    .din2(g703_p_spl_)
  );


  LA
  g_g732_p
  (
    .dout(g732_p),
    .din1(G5_p_spl_101),
    .din2(G27_p_spl_010)
  );


  FA
  g_g732_n
  (
    .dout(g732_n),
    .din1(G5_n_spl_101),
    .din2(G27_n_spl_010)
  );


  LA
  g_g733_p
  (
    .dout(g733_p),
    .din1(g694_n_spl_),
    .din2(g697_n_spl_)
  );


  FA
  g_g733_n
  (
    .dout(g733_n),
    .din1(g694_p_spl_),
    .din2(g697_p_spl_)
  );


  LA
  g_g734_p
  (
    .dout(g734_p),
    .din1(G6_p_spl_100),
    .din2(G26_p_spl_010)
  );


  FA
  g_g734_n
  (
    .dout(g734_n),
    .din1(G6_n_spl_100),
    .din2(G26_n_spl_010)
  );


  LA
  g_g735_p
  (
    .dout(g735_p),
    .din1(g688_n_spl_),
    .din2(g691_n_spl_)
  );


  FA
  g_g735_n
  (
    .dout(g735_n),
    .din1(g688_p_spl_),
    .din2(g691_p_spl_)
  );


  LA
  g_g736_p
  (
    .dout(g736_p),
    .din1(G7_p_spl_100),
    .din2(G25_p_spl_011)
  );


  FA
  g_g736_n
  (
    .dout(g736_n),
    .din1(G7_n_spl_100),
    .din2(G25_n_spl_011)
  );


  LA
  g_g737_p
  (
    .dout(g737_p),
    .din1(g682_n_spl_),
    .din2(g685_n_spl_)
  );


  FA
  g_g737_n
  (
    .dout(g737_n),
    .din1(g682_p_spl_),
    .din2(g685_p_spl_)
  );


  LA
  g_g738_p
  (
    .dout(g738_p),
    .din1(G8_p_spl_011),
    .din2(G24_p_spl_011)
  );


  FA
  g_g738_n
  (
    .dout(g738_n),
    .din1(G8_n_spl_011),
    .din2(G24_n_spl_011)
  );


  LA
  g_g739_p
  (
    .dout(g739_p),
    .din1(g676_n_spl_),
    .din2(g679_n_spl_)
  );


  FA
  g_g739_n
  (
    .dout(g739_n),
    .din1(g676_p_spl_),
    .din2(g679_p_spl_)
  );


  LA
  g_g740_p
  (
    .dout(g740_p),
    .din1(G9_p_spl_011),
    .din2(G23_p_spl_100)
  );


  FA
  g_g740_n
  (
    .dout(g740_n),
    .din1(G9_n_spl_011),
    .din2(G23_n_spl_100)
  );


  LA
  g_g741_p
  (
    .dout(g741_p),
    .din1(g670_n_spl_),
    .din2(g673_n_spl_)
  );


  FA
  g_g741_n
  (
    .dout(g741_n),
    .din1(g670_p_spl_),
    .din2(g673_p_spl_)
  );


  LA
  g_g742_p
  (
    .dout(g742_p),
    .din1(G10_p_spl_010),
    .din2(G22_p_spl_100)
  );


  FA
  g_g742_n
  (
    .dout(g742_n),
    .din1(G10_n_spl_010),
    .din2(G22_n_spl_100)
  );


  LA
  g_g743_p
  (
    .dout(g743_p),
    .din1(g664_n_spl_),
    .din2(g667_n_spl_)
  );


  FA
  g_g743_n
  (
    .dout(g743_n),
    .din1(g664_p_spl_),
    .din2(g667_p_spl_)
  );


  LA
  g_g744_p
  (
    .dout(g744_p),
    .din1(G11_p_spl_010),
    .din2(G21_p_spl_101)
  );


  FA
  g_g744_n
  (
    .dout(g744_n),
    .din1(G11_n_spl_010),
    .din2(G21_n_spl_101)
  );


  LA
  g_g745_p
  (
    .dout(g745_p),
    .din1(g658_n_spl_),
    .din2(g661_n_spl_)
  );


  FA
  g_g745_n
  (
    .dout(g745_n),
    .din1(g658_p_spl_),
    .din2(g661_p_spl_)
  );


  LA
  g_g746_p
  (
    .dout(g746_p),
    .din1(G12_p_spl_001),
    .din2(G20_p_spl_101)
  );


  FA
  g_g746_n
  (
    .dout(g746_n),
    .din1(G12_n_spl_001),
    .din2(G20_n_spl_101)
  );


  LA
  g_g747_p
  (
    .dout(g747_p),
    .din1(g652_n_spl_),
    .din2(g655_n_spl_)
  );


  FA
  g_g747_n
  (
    .dout(g747_n),
    .din1(g652_p_spl_),
    .din2(g655_p_spl_)
  );


  LA
  g_g748_p
  (
    .dout(g748_p),
    .din1(G13_p_spl_001),
    .din2(G19_p_spl_110)
  );


  FA
  g_g748_n
  (
    .dout(g748_n),
    .din1(G13_n_spl_001),
    .din2(G19_n_spl_110)
  );


  LA
  g_g749_p
  (
    .dout(g749_p),
    .din1(G15_p_spl_000),
    .din2(G17_p_spl_111)
  );


  FA
  g_g749_n
  (
    .dout(g749_n),
    .din1(G15_n_spl_000),
    .din2(G17_n_spl_110)
  );


  LA
  g_g750_p
  (
    .dout(g750_p),
    .din1(G14_p_spl_000),
    .din2(G18_p_spl_110)
  );


  FA
  g_g750_n
  (
    .dout(g750_n),
    .din1(G14_n_spl_000),
    .din2(G18_n_spl_110)
  );


  LA
  g_g751_p
  (
    .dout(g751_p),
    .din1(g749_p_spl_),
    .din2(g750_n_spl_)
  );


  FA
  g_g751_n
  (
    .dout(g751_n),
    .din1(g749_n_spl_),
    .din2(g750_p_spl_)
  );


  LA
  g_g752_p
  (
    .dout(g752_p),
    .din1(g749_p_spl_),
    .din2(g751_n_spl_)
  );


  FA
  g_g752_n
  (
    .dout(g752_n),
    .din1(g749_n_spl_),
    .din2(g751_p_spl_)
  );


  LA
  g_g753_p
  (
    .dout(g753_p),
    .din1(g750_n_spl_),
    .din2(g751_n_spl_)
  );


  FA
  g_g753_n
  (
    .dout(g753_n),
    .din1(g750_p_spl_),
    .din2(g751_p_spl_)
  );


  LA
  g_g754_p
  (
    .dout(g754_p),
    .din1(g752_n_spl_0),
    .din2(g753_n)
  );


  FA
  g_g754_n
  (
    .dout(g754_n),
    .din1(g752_p_spl_0),
    .din2(g753_p)
  );


  LA
  g_g755_p
  (
    .dout(g755_p),
    .din1(g649_n_spl_0),
    .din2(g754_n_spl_)
  );


  FA
  g_g755_n
  (
    .dout(g755_n),
    .din1(g649_p_spl_0),
    .din2(g754_p_spl_)
  );


  LA
  g_g756_p
  (
    .dout(g756_p),
    .din1(g649_p_spl_),
    .din2(g754_p_spl_)
  );


  FA
  g_g756_n
  (
    .dout(g756_n),
    .din1(g649_n_spl_),
    .din2(g754_n_spl_)
  );


  LA
  g_g757_p
  (
    .dout(g757_p),
    .din1(g755_n_spl_),
    .din2(g756_n)
  );


  FA
  g_g757_n
  (
    .dout(g757_n),
    .din1(g755_p_spl_),
    .din2(g756_p)
  );


  LA
  g_g758_p
  (
    .dout(g758_p),
    .din1(g748_n_spl_),
    .din2(g757_p_spl_)
  );


  FA
  g_g758_n
  (
    .dout(g758_n),
    .din1(g748_p_spl_),
    .din2(g757_n_spl_)
  );


  LA
  g_g759_p
  (
    .dout(g759_p),
    .din1(g748_p_spl_),
    .din2(g757_n_spl_)
  );


  FA
  g_g759_n
  (
    .dout(g759_n),
    .din1(g748_n_spl_),
    .din2(g757_p_spl_)
  );


  LA
  g_g760_p
  (
    .dout(g760_p),
    .din1(g758_n_spl_),
    .din2(g759_n)
  );


  FA
  g_g760_n
  (
    .dout(g760_n),
    .din1(g758_p_spl_),
    .din2(g759_p)
  );


  LA
  g_g761_p
  (
    .dout(g761_p),
    .din1(g747_n_spl_),
    .din2(g760_p_spl_)
  );


  FA
  g_g761_n
  (
    .dout(g761_n),
    .din1(g747_p_spl_),
    .din2(g760_n_spl_)
  );


  LA
  g_g762_p
  (
    .dout(g762_p),
    .din1(g747_p_spl_),
    .din2(g760_n_spl_)
  );


  FA
  g_g762_n
  (
    .dout(g762_n),
    .din1(g747_n_spl_),
    .din2(g760_p_spl_)
  );


  LA
  g_g763_p
  (
    .dout(g763_p),
    .din1(g761_n_spl_),
    .din2(g762_n)
  );


  FA
  g_g763_n
  (
    .dout(g763_n),
    .din1(g761_p_spl_),
    .din2(g762_p)
  );


  LA
  g_g764_p
  (
    .dout(g764_p),
    .din1(g746_n_spl_),
    .din2(g763_p_spl_)
  );


  FA
  g_g764_n
  (
    .dout(g764_n),
    .din1(g746_p_spl_),
    .din2(g763_n_spl_)
  );


  LA
  g_g765_p
  (
    .dout(g765_p),
    .din1(g746_p_spl_),
    .din2(g763_n_spl_)
  );


  FA
  g_g765_n
  (
    .dout(g765_n),
    .din1(g746_n_spl_),
    .din2(g763_p_spl_)
  );


  LA
  g_g766_p
  (
    .dout(g766_p),
    .din1(g764_n_spl_),
    .din2(g765_n)
  );


  FA
  g_g766_n
  (
    .dout(g766_n),
    .din1(g764_p_spl_),
    .din2(g765_p)
  );


  LA
  g_g767_p
  (
    .dout(g767_p),
    .din1(g745_n_spl_),
    .din2(g766_p_spl_)
  );


  FA
  g_g767_n
  (
    .dout(g767_n),
    .din1(g745_p_spl_),
    .din2(g766_n_spl_)
  );


  LA
  g_g768_p
  (
    .dout(g768_p),
    .din1(g745_p_spl_),
    .din2(g766_n_spl_)
  );


  FA
  g_g768_n
  (
    .dout(g768_n),
    .din1(g745_n_spl_),
    .din2(g766_p_spl_)
  );


  LA
  g_g769_p
  (
    .dout(g769_p),
    .din1(g767_n_spl_),
    .din2(g768_n)
  );


  FA
  g_g769_n
  (
    .dout(g769_n),
    .din1(g767_p_spl_),
    .din2(g768_p)
  );


  LA
  g_g770_p
  (
    .dout(g770_p),
    .din1(g744_n_spl_),
    .din2(g769_p_spl_)
  );


  FA
  g_g770_n
  (
    .dout(g770_n),
    .din1(g744_p_spl_),
    .din2(g769_n_spl_)
  );


  LA
  g_g771_p
  (
    .dout(g771_p),
    .din1(g744_p_spl_),
    .din2(g769_n_spl_)
  );


  FA
  g_g771_n
  (
    .dout(g771_n),
    .din1(g744_n_spl_),
    .din2(g769_p_spl_)
  );


  LA
  g_g772_p
  (
    .dout(g772_p),
    .din1(g770_n_spl_),
    .din2(g771_n)
  );


  FA
  g_g772_n
  (
    .dout(g772_n),
    .din1(g770_p_spl_),
    .din2(g771_p)
  );


  LA
  g_g773_p
  (
    .dout(g773_p),
    .din1(g743_n_spl_),
    .din2(g772_p_spl_)
  );


  FA
  g_g773_n
  (
    .dout(g773_n),
    .din1(g743_p_spl_),
    .din2(g772_n_spl_)
  );


  LA
  g_g774_p
  (
    .dout(g774_p),
    .din1(g743_p_spl_),
    .din2(g772_n_spl_)
  );


  FA
  g_g774_n
  (
    .dout(g774_n),
    .din1(g743_n_spl_),
    .din2(g772_p_spl_)
  );


  LA
  g_g775_p
  (
    .dout(g775_p),
    .din1(g773_n_spl_),
    .din2(g774_n)
  );


  FA
  g_g775_n
  (
    .dout(g775_n),
    .din1(g773_p_spl_),
    .din2(g774_p)
  );


  LA
  g_g776_p
  (
    .dout(g776_p),
    .din1(g742_n_spl_),
    .din2(g775_p_spl_)
  );


  FA
  g_g776_n
  (
    .dout(g776_n),
    .din1(g742_p_spl_),
    .din2(g775_n_spl_)
  );


  LA
  g_g777_p
  (
    .dout(g777_p),
    .din1(g742_p_spl_),
    .din2(g775_n_spl_)
  );


  FA
  g_g777_n
  (
    .dout(g777_n),
    .din1(g742_n_spl_),
    .din2(g775_p_spl_)
  );


  LA
  g_g778_p
  (
    .dout(g778_p),
    .din1(g776_n_spl_),
    .din2(g777_n)
  );


  FA
  g_g778_n
  (
    .dout(g778_n),
    .din1(g776_p_spl_),
    .din2(g777_p)
  );


  LA
  g_g779_p
  (
    .dout(g779_p),
    .din1(g741_n_spl_),
    .din2(g778_p_spl_)
  );


  FA
  g_g779_n
  (
    .dout(g779_n),
    .din1(g741_p_spl_),
    .din2(g778_n_spl_)
  );


  LA
  g_g780_p
  (
    .dout(g780_p),
    .din1(g741_p_spl_),
    .din2(g778_n_spl_)
  );


  FA
  g_g780_n
  (
    .dout(g780_n),
    .din1(g741_n_spl_),
    .din2(g778_p_spl_)
  );


  LA
  g_g781_p
  (
    .dout(g781_p),
    .din1(g779_n_spl_),
    .din2(g780_n)
  );


  FA
  g_g781_n
  (
    .dout(g781_n),
    .din1(g779_p_spl_),
    .din2(g780_p)
  );


  LA
  g_g782_p
  (
    .dout(g782_p),
    .din1(g740_n_spl_),
    .din2(g781_p_spl_)
  );


  FA
  g_g782_n
  (
    .dout(g782_n),
    .din1(g740_p_spl_),
    .din2(g781_n_spl_)
  );


  LA
  g_g783_p
  (
    .dout(g783_p),
    .din1(g740_p_spl_),
    .din2(g781_n_spl_)
  );


  FA
  g_g783_n
  (
    .dout(g783_n),
    .din1(g740_n_spl_),
    .din2(g781_p_spl_)
  );


  LA
  g_g784_p
  (
    .dout(g784_p),
    .din1(g782_n_spl_),
    .din2(g783_n)
  );


  FA
  g_g784_n
  (
    .dout(g784_n),
    .din1(g782_p_spl_),
    .din2(g783_p)
  );


  LA
  g_g785_p
  (
    .dout(g785_p),
    .din1(g739_n_spl_),
    .din2(g784_p_spl_)
  );


  FA
  g_g785_n
  (
    .dout(g785_n),
    .din1(g739_p_spl_),
    .din2(g784_n_spl_)
  );


  LA
  g_g786_p
  (
    .dout(g786_p),
    .din1(g739_p_spl_),
    .din2(g784_n_spl_)
  );


  FA
  g_g786_n
  (
    .dout(g786_n),
    .din1(g739_n_spl_),
    .din2(g784_p_spl_)
  );


  LA
  g_g787_p
  (
    .dout(g787_p),
    .din1(g785_n_spl_),
    .din2(g786_n)
  );


  FA
  g_g787_n
  (
    .dout(g787_n),
    .din1(g785_p_spl_),
    .din2(g786_p)
  );


  LA
  g_g788_p
  (
    .dout(g788_p),
    .din1(g738_n_spl_),
    .din2(g787_p_spl_)
  );


  FA
  g_g788_n
  (
    .dout(g788_n),
    .din1(g738_p_spl_),
    .din2(g787_n_spl_)
  );


  LA
  g_g789_p
  (
    .dout(g789_p),
    .din1(g738_p_spl_),
    .din2(g787_n_spl_)
  );


  FA
  g_g789_n
  (
    .dout(g789_n),
    .din1(g738_n_spl_),
    .din2(g787_p_spl_)
  );


  LA
  g_g790_p
  (
    .dout(g790_p),
    .din1(g788_n_spl_),
    .din2(g789_n)
  );


  FA
  g_g790_n
  (
    .dout(g790_n),
    .din1(g788_p_spl_),
    .din2(g789_p)
  );


  LA
  g_g791_p
  (
    .dout(g791_p),
    .din1(g737_n_spl_),
    .din2(g790_p_spl_)
  );


  FA
  g_g791_n
  (
    .dout(g791_n),
    .din1(g737_p_spl_),
    .din2(g790_n_spl_)
  );


  LA
  g_g792_p
  (
    .dout(g792_p),
    .din1(g737_p_spl_),
    .din2(g790_n_spl_)
  );


  FA
  g_g792_n
  (
    .dout(g792_n),
    .din1(g737_n_spl_),
    .din2(g790_p_spl_)
  );


  LA
  g_g793_p
  (
    .dout(g793_p),
    .din1(g791_n_spl_),
    .din2(g792_n)
  );


  FA
  g_g793_n
  (
    .dout(g793_n),
    .din1(g791_p_spl_),
    .din2(g792_p)
  );


  LA
  g_g794_p
  (
    .dout(g794_p),
    .din1(g736_n_spl_),
    .din2(g793_p_spl_)
  );


  FA
  g_g794_n
  (
    .dout(g794_n),
    .din1(g736_p_spl_),
    .din2(g793_n_spl_)
  );


  LA
  g_g795_p
  (
    .dout(g795_p),
    .din1(g736_p_spl_),
    .din2(g793_n_spl_)
  );


  FA
  g_g795_n
  (
    .dout(g795_n),
    .din1(g736_n_spl_),
    .din2(g793_p_spl_)
  );


  LA
  g_g796_p
  (
    .dout(g796_p),
    .din1(g794_n_spl_),
    .din2(g795_n)
  );


  FA
  g_g796_n
  (
    .dout(g796_n),
    .din1(g794_p_spl_),
    .din2(g795_p)
  );


  LA
  g_g797_p
  (
    .dout(g797_p),
    .din1(g735_n_spl_),
    .din2(g796_p_spl_)
  );


  FA
  g_g797_n
  (
    .dout(g797_n),
    .din1(g735_p_spl_),
    .din2(g796_n_spl_)
  );


  LA
  g_g798_p
  (
    .dout(g798_p),
    .din1(g735_p_spl_),
    .din2(g796_n_spl_)
  );


  FA
  g_g798_n
  (
    .dout(g798_n),
    .din1(g735_n_spl_),
    .din2(g796_p_spl_)
  );


  LA
  g_g799_p
  (
    .dout(g799_p),
    .din1(g797_n_spl_),
    .din2(g798_n)
  );


  FA
  g_g799_n
  (
    .dout(g799_n),
    .din1(g797_p_spl_),
    .din2(g798_p)
  );


  LA
  g_g800_p
  (
    .dout(g800_p),
    .din1(g734_n_spl_),
    .din2(g799_p_spl_)
  );


  FA
  g_g800_n
  (
    .dout(g800_n),
    .din1(g734_p_spl_),
    .din2(g799_n_spl_)
  );


  LA
  g_g801_p
  (
    .dout(g801_p),
    .din1(g734_p_spl_),
    .din2(g799_n_spl_)
  );


  FA
  g_g801_n
  (
    .dout(g801_n),
    .din1(g734_n_spl_),
    .din2(g799_p_spl_)
  );


  LA
  g_g802_p
  (
    .dout(g802_p),
    .din1(g800_n_spl_),
    .din2(g801_n)
  );


  FA
  g_g802_n
  (
    .dout(g802_n),
    .din1(g800_p_spl_),
    .din2(g801_p)
  );


  LA
  g_g803_p
  (
    .dout(g803_p),
    .din1(g733_n_spl_),
    .din2(g802_p_spl_)
  );


  FA
  g_g803_n
  (
    .dout(g803_n),
    .din1(g733_p_spl_),
    .din2(g802_n_spl_)
  );


  LA
  g_g804_p
  (
    .dout(g804_p),
    .din1(g733_p_spl_),
    .din2(g802_n_spl_)
  );


  FA
  g_g804_n
  (
    .dout(g804_n),
    .din1(g733_n_spl_),
    .din2(g802_p_spl_)
  );


  LA
  g_g805_p
  (
    .dout(g805_p),
    .din1(g803_n_spl_),
    .din2(g804_n)
  );


  FA
  g_g805_n
  (
    .dout(g805_n),
    .din1(g803_p_spl_),
    .din2(g804_p)
  );


  LA
  g_g806_p
  (
    .dout(g806_p),
    .din1(g732_n_spl_),
    .din2(g805_p_spl_)
  );


  FA
  g_g806_n
  (
    .dout(g806_n),
    .din1(g732_p_spl_),
    .din2(g805_n_spl_)
  );


  LA
  g_g807_p
  (
    .dout(g807_p),
    .din1(g732_p_spl_),
    .din2(g805_n_spl_)
  );


  FA
  g_g807_n
  (
    .dout(g807_n),
    .din1(g732_n_spl_),
    .din2(g805_p_spl_)
  );


  LA
  g_g808_p
  (
    .dout(g808_p),
    .din1(g806_n_spl_),
    .din2(g807_n)
  );


  FA
  g_g808_n
  (
    .dout(g808_n),
    .din1(g806_p_spl_),
    .din2(g807_p)
  );


  LA
  g_g809_p
  (
    .dout(g809_p),
    .din1(g731_n_spl_),
    .din2(g808_p_spl_)
  );


  FA
  g_g809_n
  (
    .dout(g809_n),
    .din1(g731_p_spl_),
    .din2(g808_n_spl_)
  );


  LA
  g_g810_p
  (
    .dout(g810_p),
    .din1(g731_p_spl_),
    .din2(g808_n_spl_)
  );


  FA
  g_g810_n
  (
    .dout(g810_n),
    .din1(g731_n_spl_),
    .din2(g808_p_spl_)
  );


  LA
  g_g811_p
  (
    .dout(g811_p),
    .din1(g809_n_spl_),
    .din2(g810_n)
  );


  FA
  g_g811_n
  (
    .dout(g811_n),
    .din1(g809_p_spl_),
    .din2(g810_p)
  );


  LA
  g_g812_p
  (
    .dout(g812_p),
    .din1(g730_n_spl_),
    .din2(g811_p_spl_)
  );


  FA
  g_g812_n
  (
    .dout(g812_n),
    .din1(g730_p_spl_),
    .din2(g811_n_spl_)
  );


  LA
  g_g813_p
  (
    .dout(g813_p),
    .din1(g730_p_spl_),
    .din2(g811_n_spl_)
  );


  FA
  g_g813_n
  (
    .dout(g813_n),
    .din1(g730_n_spl_),
    .din2(g811_p_spl_)
  );


  LA
  g_g814_p
  (
    .dout(g814_p),
    .din1(g812_n_spl_),
    .din2(g813_n)
  );


  FA
  g_g814_n
  (
    .dout(g814_n),
    .din1(g812_p_spl_),
    .din2(g813_p)
  );


  LA
  g_g815_p
  (
    .dout(g815_p),
    .din1(g729_n_spl_),
    .din2(g814_p_spl_)
  );


  FA
  g_g815_n
  (
    .dout(g815_n),
    .din1(g729_p_spl_),
    .din2(g814_n_spl_)
  );


  LA
  g_g816_p
  (
    .dout(g816_p),
    .din1(g729_p_spl_),
    .din2(g814_n_spl_)
  );


  FA
  g_g816_n
  (
    .dout(g816_n),
    .din1(g729_n_spl_),
    .din2(g814_p_spl_)
  );


  LA
  g_g817_p
  (
    .dout(g817_p),
    .din1(g815_n_spl_),
    .din2(g816_n)
  );


  FA
  g_g817_n
  (
    .dout(g817_n),
    .din1(g815_p_spl_),
    .din2(g816_p)
  );


  LA
  g_g818_p
  (
    .dout(g818_p),
    .din1(g728_n_spl_),
    .din2(g817_p_spl_)
  );


  FA
  g_g818_n
  (
    .dout(g818_n),
    .din1(g728_p_spl_),
    .din2(g817_n_spl_)
  );


  LA
  g_g819_p
  (
    .dout(g819_p),
    .din1(g728_p_spl_),
    .din2(g817_n_spl_)
  );


  FA
  g_g819_n
  (
    .dout(g819_n),
    .din1(g728_n_spl_),
    .din2(g817_p_spl_)
  );


  LA
  g_g820_p
  (
    .dout(g820_p),
    .din1(g818_n_spl_),
    .din2(g819_n)
  );


  FA
  g_g820_n
  (
    .dout(g820_n),
    .din1(g818_p_spl_),
    .din2(g819_p)
  );


  LA
  g_g821_p
  (
    .dout(g821_p),
    .din1(g727_n_spl_),
    .din2(g820_p_spl_)
  );


  FA
  g_g821_n
  (
    .dout(g821_n),
    .din1(g727_p_spl_),
    .din2(g820_n_spl_)
  );


  LA
  g_g822_p
  (
    .dout(g822_p),
    .din1(g727_p_spl_),
    .din2(g820_n_spl_)
  );


  FA
  g_g822_n
  (
    .dout(g822_n),
    .din1(g727_n_spl_),
    .din2(g820_p_spl_)
  );


  LA
  g_g823_p
  (
    .dout(g823_p),
    .din1(g821_n_spl_),
    .din2(g822_n)
  );


  FA
  g_g823_n
  (
    .dout(g823_n),
    .din1(g821_p_spl_),
    .din2(g822_p)
  );


  LA
  g_g824_p
  (
    .dout(g824_p),
    .din1(g726_n_spl_),
    .din2(g823_p_spl_)
  );


  FA
  g_g824_n
  (
    .dout(g824_n),
    .din1(g726_p_spl_),
    .din2(g823_n_spl_)
  );


  LA
  g_g825_p
  (
    .dout(g825_p),
    .din1(g726_p_spl_),
    .din2(g823_n_spl_)
  );


  FA
  g_g825_n
  (
    .dout(g825_n),
    .din1(g726_n_spl_),
    .din2(g823_p_spl_)
  );


  LA
  g_g826_p
  (
    .dout(g826_p),
    .din1(g824_n_spl_),
    .din2(g825_n)
  );


  FA
  g_g826_n
  (
    .dout(g826_n),
    .din1(g824_p_spl_),
    .din2(g825_p)
  );


  LA
  g_g827_p
  (
    .dout(g827_p),
    .din1(g725_n_spl_),
    .din2(g826_p_spl_)
  );


  FA
  g_g827_n
  (
    .dout(g827_n),
    .din1(g725_p_spl_),
    .din2(g826_n_spl_)
  );


  LA
  g_g828_p
  (
    .dout(g828_p),
    .din1(g725_p_spl_),
    .din2(g826_n_spl_)
  );


  FA
  g_g828_n
  (
    .dout(g828_n),
    .din1(g725_n_spl_),
    .din2(g826_p_spl_)
  );


  LA
  g_g829_p
  (
    .dout(g829_p),
    .din1(g827_n_spl_),
    .din2(g828_n)
  );


  FA
  g_g829_n
  (
    .dout(g829_n),
    .din1(g827_p_spl_),
    .din2(g828_p)
  );


  LA
  g_g830_p
  (
    .dout(g830_p),
    .din1(g724_n),
    .din2(g829_p)
  );


  FA
  g_g830_n
  (
    .dout(g830_n),
    .din1(g724_p_spl_),
    .din2(g829_n_spl_)
  );


  LA
  g_g831_p
  (
    .dout(g831_p),
    .din1(g724_p_spl_),
    .din2(g829_n_spl_)
  );


  FA
  g_g832_n
  (
    .dout(g832_n),
    .din1(g830_p_spl_),
    .din2(g831_p)
  );


  LA
  g_g833_p
  (
    .dout(g833_p),
    .din1(G1_p_spl_111),
    .din2(G32_p_spl_000)
  );


  FA
  g_g833_n
  (
    .dout(g833_n),
    .din1(G1_n_spl_11),
    .din2(G32_n_spl_000)
  );


  LA
  g_g834_p
  (
    .dout(g834_p),
    .din1(g827_n_spl_),
    .din2(g830_n)
  );


  FA
  g_g834_n
  (
    .dout(g834_n),
    .din1(g827_p_spl_),
    .din2(g830_p_spl_)
  );


  LA
  g_g835_p
  (
    .dout(g835_p),
    .din1(G2_p_spl_111),
    .din2(G31_p_spl_000)
  );


  FA
  g_g835_n
  (
    .dout(g835_n),
    .din1(G2_n_spl_111),
    .din2(G31_n_spl_000)
  );


  LA
  g_g836_p
  (
    .dout(g836_p),
    .din1(g821_n_spl_),
    .din2(g824_n_spl_)
  );


  FA
  g_g836_n
  (
    .dout(g836_n),
    .din1(g821_p_spl_),
    .din2(g824_p_spl_)
  );


  LA
  g_g837_p
  (
    .dout(g837_p),
    .din1(G3_p_spl_110),
    .din2(G30_p_spl_001)
  );


  FA
  g_g837_n
  (
    .dout(g837_n),
    .din1(G3_n_spl_110),
    .din2(G30_n_spl_001)
  );


  LA
  g_g838_p
  (
    .dout(g838_p),
    .din1(g815_n_spl_),
    .din2(g818_n_spl_)
  );


  FA
  g_g838_n
  (
    .dout(g838_n),
    .din1(g815_p_spl_),
    .din2(g818_p_spl_)
  );


  LA
  g_g839_p
  (
    .dout(g839_p),
    .din1(G4_p_spl_110),
    .din2(G29_p_spl_001)
  );


  FA
  g_g839_n
  (
    .dout(g839_n),
    .din1(G4_n_spl_110),
    .din2(G29_n_spl_001)
  );


  LA
  g_g840_p
  (
    .dout(g840_p),
    .din1(g809_n_spl_),
    .din2(g812_n_spl_)
  );


  FA
  g_g840_n
  (
    .dout(g840_n),
    .din1(g809_p_spl_),
    .din2(g812_p_spl_)
  );


  LA
  g_g841_p
  (
    .dout(g841_p),
    .din1(G5_p_spl_101),
    .din2(G28_p_spl_010)
  );


  FA
  g_g841_n
  (
    .dout(g841_n),
    .din1(G5_n_spl_101),
    .din2(G28_n_spl_010)
  );


  LA
  g_g842_p
  (
    .dout(g842_p),
    .din1(g803_n_spl_),
    .din2(g806_n_spl_)
  );


  FA
  g_g842_n
  (
    .dout(g842_n),
    .din1(g803_p_spl_),
    .din2(g806_p_spl_)
  );


  LA
  g_g843_p
  (
    .dout(g843_p),
    .din1(G6_p_spl_101),
    .din2(G27_p_spl_010)
  );


  FA
  g_g843_n
  (
    .dout(g843_n),
    .din1(G6_n_spl_101),
    .din2(G27_n_spl_010)
  );


  LA
  g_g844_p
  (
    .dout(g844_p),
    .din1(g797_n_spl_),
    .din2(g800_n_spl_)
  );


  FA
  g_g844_n
  (
    .dout(g844_n),
    .din1(g797_p_spl_),
    .din2(g800_p_spl_)
  );


  LA
  g_g845_p
  (
    .dout(g845_p),
    .din1(G7_p_spl_100),
    .din2(G26_p_spl_011)
  );


  FA
  g_g845_n
  (
    .dout(g845_n),
    .din1(G7_n_spl_100),
    .din2(G26_n_spl_011)
  );


  LA
  g_g846_p
  (
    .dout(g846_p),
    .din1(g791_n_spl_),
    .din2(g794_n_spl_)
  );


  FA
  g_g846_n
  (
    .dout(g846_n),
    .din1(g791_p_spl_),
    .din2(g794_p_spl_)
  );


  LA
  g_g847_p
  (
    .dout(g847_p),
    .din1(G8_p_spl_100),
    .din2(G25_p_spl_011)
  );


  FA
  g_g847_n
  (
    .dout(g847_n),
    .din1(G8_n_spl_100),
    .din2(G25_n_spl_011)
  );


  LA
  g_g848_p
  (
    .dout(g848_p),
    .din1(g785_n_spl_),
    .din2(g788_n_spl_)
  );


  FA
  g_g848_n
  (
    .dout(g848_n),
    .din1(g785_p_spl_),
    .din2(g788_p_spl_)
  );


  LA
  g_g849_p
  (
    .dout(g849_p),
    .din1(G9_p_spl_011),
    .din2(G24_p_spl_100)
  );


  FA
  g_g849_n
  (
    .dout(g849_n),
    .din1(G9_n_spl_011),
    .din2(G24_n_spl_100)
  );


  LA
  g_g850_p
  (
    .dout(g850_p),
    .din1(g779_n_spl_),
    .din2(g782_n_spl_)
  );


  FA
  g_g850_n
  (
    .dout(g850_n),
    .din1(g779_p_spl_),
    .din2(g782_p_spl_)
  );


  LA
  g_g851_p
  (
    .dout(g851_p),
    .din1(G10_p_spl_011),
    .din2(G23_p_spl_100)
  );


  FA
  g_g851_n
  (
    .dout(g851_n),
    .din1(G10_n_spl_011),
    .din2(G23_n_spl_100)
  );


  LA
  g_g852_p
  (
    .dout(g852_p),
    .din1(g773_n_spl_),
    .din2(g776_n_spl_)
  );


  FA
  g_g852_n
  (
    .dout(g852_n),
    .din1(g773_p_spl_),
    .din2(g776_p_spl_)
  );


  LA
  g_g853_p
  (
    .dout(g853_p),
    .din1(G11_p_spl_010),
    .din2(G22_p_spl_101)
  );


  FA
  g_g853_n
  (
    .dout(g853_n),
    .din1(G11_n_spl_010),
    .din2(G22_n_spl_101)
  );


  LA
  g_g854_p
  (
    .dout(g854_p),
    .din1(g767_n_spl_),
    .din2(g770_n_spl_)
  );


  FA
  g_g854_n
  (
    .dout(g854_n),
    .din1(g767_p_spl_),
    .din2(g770_p_spl_)
  );


  LA
  g_g855_p
  (
    .dout(g855_p),
    .din1(G12_p_spl_010),
    .din2(G21_p_spl_101)
  );


  FA
  g_g855_n
  (
    .dout(g855_n),
    .din1(G12_n_spl_010),
    .din2(G21_n_spl_101)
  );


  LA
  g_g856_p
  (
    .dout(g856_p),
    .din1(g761_n_spl_),
    .din2(g764_n_spl_)
  );


  FA
  g_g856_n
  (
    .dout(g856_n),
    .din1(g761_p_spl_),
    .din2(g764_p_spl_)
  );


  LA
  g_g857_p
  (
    .dout(g857_p),
    .din1(G13_p_spl_001),
    .din2(G20_p_spl_110)
  );


  FA
  g_g857_n
  (
    .dout(g857_n),
    .din1(G13_n_spl_001),
    .din2(G20_n_spl_110)
  );


  LA
  g_g858_p
  (
    .dout(g858_p),
    .din1(g755_n_spl_),
    .din2(g758_n_spl_)
  );


  FA
  g_g858_n
  (
    .dout(g858_n),
    .din1(g755_p_spl_),
    .din2(g758_p_spl_)
  );


  LA
  g_g859_p
  (
    .dout(g859_p),
    .din1(G14_p_spl_001),
    .din2(G19_p_spl_110)
  );


  FA
  g_g859_n
  (
    .dout(g859_n),
    .din1(G14_n_spl_001),
    .din2(G19_n_spl_110)
  );


  LA
  g_g860_p
  (
    .dout(g860_p),
    .din1(G16_p_spl_000),
    .din2(G17_p_spl_111)
  );


  FA
  g_g860_n
  (
    .dout(g860_n),
    .din1(G16_n_spl_000),
    .din2(G17_n_spl_11)
  );


  LA
  g_g861_p
  (
    .dout(g861_p),
    .din1(G15_p_spl_000),
    .din2(G18_p_spl_111)
  );


  FA
  g_g861_n
  (
    .dout(g861_n),
    .din1(G15_n_spl_000),
    .din2(G18_n_spl_111)
  );


  LA
  g_g862_p
  (
    .dout(g862_p),
    .din1(g860_p_spl_),
    .din2(g861_n_spl_)
  );


  FA
  g_g862_n
  (
    .dout(g862_n),
    .din1(g860_n_spl_),
    .din2(g861_p_spl_)
  );


  LA
  g_g863_p
  (
    .dout(g863_p),
    .din1(g860_p_spl_),
    .din2(g862_n_spl_)
  );


  FA
  g_g863_n
  (
    .dout(g863_n),
    .din1(g860_n_spl_),
    .din2(g862_p_spl_)
  );


  LA
  g_g864_p
  (
    .dout(g864_p),
    .din1(g861_n_spl_),
    .din2(g862_n_spl_)
  );


  FA
  g_g864_n
  (
    .dout(g864_n),
    .din1(g861_p_spl_),
    .din2(g862_p_spl_)
  );


  LA
  g_g865_p
  (
    .dout(g865_p),
    .din1(g863_n_spl_),
    .din2(g864_n)
  );


  FA
  g_g865_n
  (
    .dout(g865_n),
    .din1(g863_p_spl_),
    .din2(g864_p)
  );


  LA
  g_g866_p
  (
    .dout(g866_p),
    .din1(g752_n_spl_0),
    .din2(g865_n_spl_)
  );


  FA
  g_g866_n
  (
    .dout(g866_n),
    .din1(g752_p_spl_0),
    .din2(g865_p_spl_)
  );


  LA
  g_g867_p
  (
    .dout(g867_p),
    .din1(g752_p_spl_),
    .din2(g865_p_spl_)
  );


  FA
  g_g867_n
  (
    .dout(g867_n),
    .din1(g752_n_spl_),
    .din2(g865_n_spl_)
  );


  LA
  g_g868_p
  (
    .dout(g868_p),
    .din1(g866_n_spl_),
    .din2(g867_n)
  );


  FA
  g_g868_n
  (
    .dout(g868_n),
    .din1(g866_p_spl_),
    .din2(g867_p)
  );


  LA
  g_g869_p
  (
    .dout(g869_p),
    .din1(g859_n_spl_),
    .din2(g868_p_spl_)
  );


  FA
  g_g869_n
  (
    .dout(g869_n),
    .din1(g859_p_spl_),
    .din2(g868_n_spl_)
  );


  LA
  g_g870_p
  (
    .dout(g870_p),
    .din1(g859_p_spl_),
    .din2(g868_n_spl_)
  );


  FA
  g_g870_n
  (
    .dout(g870_n),
    .din1(g859_n_spl_),
    .din2(g868_p_spl_)
  );


  LA
  g_g871_p
  (
    .dout(g871_p),
    .din1(g869_n_spl_),
    .din2(g870_n)
  );


  FA
  g_g871_n
  (
    .dout(g871_n),
    .din1(g869_p_spl_),
    .din2(g870_p)
  );


  LA
  g_g872_p
  (
    .dout(g872_p),
    .din1(g858_n_spl_),
    .din2(g871_p_spl_)
  );


  FA
  g_g872_n
  (
    .dout(g872_n),
    .din1(g858_p_spl_),
    .din2(g871_n_spl_)
  );


  LA
  g_g873_p
  (
    .dout(g873_p),
    .din1(g858_p_spl_),
    .din2(g871_n_spl_)
  );


  FA
  g_g873_n
  (
    .dout(g873_n),
    .din1(g858_n_spl_),
    .din2(g871_p_spl_)
  );


  LA
  g_g874_p
  (
    .dout(g874_p),
    .din1(g872_n_spl_),
    .din2(g873_n)
  );


  FA
  g_g874_n
  (
    .dout(g874_n),
    .din1(g872_p_spl_),
    .din2(g873_p)
  );


  LA
  g_g875_p
  (
    .dout(g875_p),
    .din1(g857_n_spl_),
    .din2(g874_p_spl_)
  );


  FA
  g_g875_n
  (
    .dout(g875_n),
    .din1(g857_p_spl_),
    .din2(g874_n_spl_)
  );


  LA
  g_g876_p
  (
    .dout(g876_p),
    .din1(g857_p_spl_),
    .din2(g874_n_spl_)
  );


  FA
  g_g876_n
  (
    .dout(g876_n),
    .din1(g857_n_spl_),
    .din2(g874_p_spl_)
  );


  LA
  g_g877_p
  (
    .dout(g877_p),
    .din1(g875_n_spl_),
    .din2(g876_n)
  );


  FA
  g_g877_n
  (
    .dout(g877_n),
    .din1(g875_p_spl_),
    .din2(g876_p)
  );


  LA
  g_g878_p
  (
    .dout(g878_p),
    .din1(g856_n_spl_),
    .din2(g877_p_spl_)
  );


  FA
  g_g878_n
  (
    .dout(g878_n),
    .din1(g856_p_spl_),
    .din2(g877_n_spl_)
  );


  LA
  g_g879_p
  (
    .dout(g879_p),
    .din1(g856_p_spl_),
    .din2(g877_n_spl_)
  );


  FA
  g_g879_n
  (
    .dout(g879_n),
    .din1(g856_n_spl_),
    .din2(g877_p_spl_)
  );


  LA
  g_g880_p
  (
    .dout(g880_p),
    .din1(g878_n_spl_),
    .din2(g879_n)
  );


  FA
  g_g880_n
  (
    .dout(g880_n),
    .din1(g878_p_spl_),
    .din2(g879_p)
  );


  LA
  g_g881_p
  (
    .dout(g881_p),
    .din1(g855_n_spl_),
    .din2(g880_p_spl_)
  );


  FA
  g_g881_n
  (
    .dout(g881_n),
    .din1(g855_p_spl_),
    .din2(g880_n_spl_)
  );


  LA
  g_g882_p
  (
    .dout(g882_p),
    .din1(g855_p_spl_),
    .din2(g880_n_spl_)
  );


  FA
  g_g882_n
  (
    .dout(g882_n),
    .din1(g855_n_spl_),
    .din2(g880_p_spl_)
  );


  LA
  g_g883_p
  (
    .dout(g883_p),
    .din1(g881_n_spl_),
    .din2(g882_n)
  );


  FA
  g_g883_n
  (
    .dout(g883_n),
    .din1(g881_p_spl_),
    .din2(g882_p)
  );


  LA
  g_g884_p
  (
    .dout(g884_p),
    .din1(g854_n_spl_),
    .din2(g883_p_spl_)
  );


  FA
  g_g884_n
  (
    .dout(g884_n),
    .din1(g854_p_spl_),
    .din2(g883_n_spl_)
  );


  LA
  g_g885_p
  (
    .dout(g885_p),
    .din1(g854_p_spl_),
    .din2(g883_n_spl_)
  );


  FA
  g_g885_n
  (
    .dout(g885_n),
    .din1(g854_n_spl_),
    .din2(g883_p_spl_)
  );


  LA
  g_g886_p
  (
    .dout(g886_p),
    .din1(g884_n_spl_),
    .din2(g885_n)
  );


  FA
  g_g886_n
  (
    .dout(g886_n),
    .din1(g884_p_spl_),
    .din2(g885_p)
  );


  LA
  g_g887_p
  (
    .dout(g887_p),
    .din1(g853_n_spl_),
    .din2(g886_p_spl_)
  );


  FA
  g_g887_n
  (
    .dout(g887_n),
    .din1(g853_p_spl_),
    .din2(g886_n_spl_)
  );


  LA
  g_g888_p
  (
    .dout(g888_p),
    .din1(g853_p_spl_),
    .din2(g886_n_spl_)
  );


  FA
  g_g888_n
  (
    .dout(g888_n),
    .din1(g853_n_spl_),
    .din2(g886_p_spl_)
  );


  LA
  g_g889_p
  (
    .dout(g889_p),
    .din1(g887_n_spl_),
    .din2(g888_n)
  );


  FA
  g_g889_n
  (
    .dout(g889_n),
    .din1(g887_p_spl_),
    .din2(g888_p)
  );


  LA
  g_g890_p
  (
    .dout(g890_p),
    .din1(g852_n_spl_),
    .din2(g889_p_spl_)
  );


  FA
  g_g890_n
  (
    .dout(g890_n),
    .din1(g852_p_spl_),
    .din2(g889_n_spl_)
  );


  LA
  g_g891_p
  (
    .dout(g891_p),
    .din1(g852_p_spl_),
    .din2(g889_n_spl_)
  );


  FA
  g_g891_n
  (
    .dout(g891_n),
    .din1(g852_n_spl_),
    .din2(g889_p_spl_)
  );


  LA
  g_g892_p
  (
    .dout(g892_p),
    .din1(g890_n_spl_),
    .din2(g891_n)
  );


  FA
  g_g892_n
  (
    .dout(g892_n),
    .din1(g890_p_spl_),
    .din2(g891_p)
  );


  LA
  g_g893_p
  (
    .dout(g893_p),
    .din1(g851_n_spl_),
    .din2(g892_p_spl_)
  );


  FA
  g_g893_n
  (
    .dout(g893_n),
    .din1(g851_p_spl_),
    .din2(g892_n_spl_)
  );


  LA
  g_g894_p
  (
    .dout(g894_p),
    .din1(g851_p_spl_),
    .din2(g892_n_spl_)
  );


  FA
  g_g894_n
  (
    .dout(g894_n),
    .din1(g851_n_spl_),
    .din2(g892_p_spl_)
  );


  LA
  g_g895_p
  (
    .dout(g895_p),
    .din1(g893_n_spl_),
    .din2(g894_n)
  );


  FA
  g_g895_n
  (
    .dout(g895_n),
    .din1(g893_p_spl_),
    .din2(g894_p)
  );


  LA
  g_g896_p
  (
    .dout(g896_p),
    .din1(g850_n_spl_),
    .din2(g895_p_spl_)
  );


  FA
  g_g896_n
  (
    .dout(g896_n),
    .din1(g850_p_spl_),
    .din2(g895_n_spl_)
  );


  LA
  g_g897_p
  (
    .dout(g897_p),
    .din1(g850_p_spl_),
    .din2(g895_n_spl_)
  );


  FA
  g_g897_n
  (
    .dout(g897_n),
    .din1(g850_n_spl_),
    .din2(g895_p_spl_)
  );


  LA
  g_g898_p
  (
    .dout(g898_p),
    .din1(g896_n_spl_),
    .din2(g897_n)
  );


  FA
  g_g898_n
  (
    .dout(g898_n),
    .din1(g896_p_spl_),
    .din2(g897_p)
  );


  LA
  g_g899_p
  (
    .dout(g899_p),
    .din1(g849_n_spl_),
    .din2(g898_p_spl_)
  );


  FA
  g_g899_n
  (
    .dout(g899_n),
    .din1(g849_p_spl_),
    .din2(g898_n_spl_)
  );


  LA
  g_g900_p
  (
    .dout(g900_p),
    .din1(g849_p_spl_),
    .din2(g898_n_spl_)
  );


  FA
  g_g900_n
  (
    .dout(g900_n),
    .din1(g849_n_spl_),
    .din2(g898_p_spl_)
  );


  LA
  g_g901_p
  (
    .dout(g901_p),
    .din1(g899_n_spl_),
    .din2(g900_n)
  );


  FA
  g_g901_n
  (
    .dout(g901_n),
    .din1(g899_p_spl_),
    .din2(g900_p)
  );


  LA
  g_g902_p
  (
    .dout(g902_p),
    .din1(g848_n_spl_),
    .din2(g901_p_spl_)
  );


  FA
  g_g902_n
  (
    .dout(g902_n),
    .din1(g848_p_spl_),
    .din2(g901_n_spl_)
  );


  LA
  g_g903_p
  (
    .dout(g903_p),
    .din1(g848_p_spl_),
    .din2(g901_n_spl_)
  );


  FA
  g_g903_n
  (
    .dout(g903_n),
    .din1(g848_n_spl_),
    .din2(g901_p_spl_)
  );


  LA
  g_g904_p
  (
    .dout(g904_p),
    .din1(g902_n_spl_),
    .din2(g903_n)
  );


  FA
  g_g904_n
  (
    .dout(g904_n),
    .din1(g902_p_spl_),
    .din2(g903_p)
  );


  LA
  g_g905_p
  (
    .dout(g905_p),
    .din1(g847_n_spl_),
    .din2(g904_p_spl_)
  );


  FA
  g_g905_n
  (
    .dout(g905_n),
    .din1(g847_p_spl_),
    .din2(g904_n_spl_)
  );


  LA
  g_g906_p
  (
    .dout(g906_p),
    .din1(g847_p_spl_),
    .din2(g904_n_spl_)
  );


  FA
  g_g906_n
  (
    .dout(g906_n),
    .din1(g847_n_spl_),
    .din2(g904_p_spl_)
  );


  LA
  g_g907_p
  (
    .dout(g907_p),
    .din1(g905_n_spl_),
    .din2(g906_n)
  );


  FA
  g_g907_n
  (
    .dout(g907_n),
    .din1(g905_p_spl_),
    .din2(g906_p)
  );


  LA
  g_g908_p
  (
    .dout(g908_p),
    .din1(g846_n_spl_),
    .din2(g907_p_spl_)
  );


  FA
  g_g908_n
  (
    .dout(g908_n),
    .din1(g846_p_spl_),
    .din2(g907_n_spl_)
  );


  LA
  g_g909_p
  (
    .dout(g909_p),
    .din1(g846_p_spl_),
    .din2(g907_n_spl_)
  );


  FA
  g_g909_n
  (
    .dout(g909_n),
    .din1(g846_n_spl_),
    .din2(g907_p_spl_)
  );


  LA
  g_g910_p
  (
    .dout(g910_p),
    .din1(g908_n_spl_),
    .din2(g909_n)
  );


  FA
  g_g910_n
  (
    .dout(g910_n),
    .din1(g908_p_spl_),
    .din2(g909_p)
  );


  LA
  g_g911_p
  (
    .dout(g911_p),
    .din1(g845_n_spl_),
    .din2(g910_p_spl_)
  );


  FA
  g_g911_n
  (
    .dout(g911_n),
    .din1(g845_p_spl_),
    .din2(g910_n_spl_)
  );


  LA
  g_g912_p
  (
    .dout(g912_p),
    .din1(g845_p_spl_),
    .din2(g910_n_spl_)
  );


  FA
  g_g912_n
  (
    .dout(g912_n),
    .din1(g845_n_spl_),
    .din2(g910_p_spl_)
  );


  LA
  g_g913_p
  (
    .dout(g913_p),
    .din1(g911_n_spl_),
    .din2(g912_n)
  );


  FA
  g_g913_n
  (
    .dout(g913_n),
    .din1(g911_p_spl_),
    .din2(g912_p)
  );


  LA
  g_g914_p
  (
    .dout(g914_p),
    .din1(g844_n_spl_),
    .din2(g913_p_spl_)
  );


  FA
  g_g914_n
  (
    .dout(g914_n),
    .din1(g844_p_spl_),
    .din2(g913_n_spl_)
  );


  LA
  g_g915_p
  (
    .dout(g915_p),
    .din1(g844_p_spl_),
    .din2(g913_n_spl_)
  );


  FA
  g_g915_n
  (
    .dout(g915_n),
    .din1(g844_n_spl_),
    .din2(g913_p_spl_)
  );


  LA
  g_g916_p
  (
    .dout(g916_p),
    .din1(g914_n_spl_),
    .din2(g915_n)
  );


  FA
  g_g916_n
  (
    .dout(g916_n),
    .din1(g914_p_spl_),
    .din2(g915_p)
  );


  LA
  g_g917_p
  (
    .dout(g917_p),
    .din1(g843_n_spl_),
    .din2(g916_p_spl_)
  );


  FA
  g_g917_n
  (
    .dout(g917_n),
    .din1(g843_p_spl_),
    .din2(g916_n_spl_)
  );


  LA
  g_g918_p
  (
    .dout(g918_p),
    .din1(g843_p_spl_),
    .din2(g916_n_spl_)
  );


  FA
  g_g918_n
  (
    .dout(g918_n),
    .din1(g843_n_spl_),
    .din2(g916_p_spl_)
  );


  LA
  g_g919_p
  (
    .dout(g919_p),
    .din1(g917_n_spl_),
    .din2(g918_n)
  );


  FA
  g_g919_n
  (
    .dout(g919_n),
    .din1(g917_p_spl_),
    .din2(g918_p)
  );


  LA
  g_g920_p
  (
    .dout(g920_p),
    .din1(g842_n_spl_),
    .din2(g919_p_spl_)
  );


  FA
  g_g920_n
  (
    .dout(g920_n),
    .din1(g842_p_spl_),
    .din2(g919_n_spl_)
  );


  LA
  g_g921_p
  (
    .dout(g921_p),
    .din1(g842_p_spl_),
    .din2(g919_n_spl_)
  );


  FA
  g_g921_n
  (
    .dout(g921_n),
    .din1(g842_n_spl_),
    .din2(g919_p_spl_)
  );


  LA
  g_g922_p
  (
    .dout(g922_p),
    .din1(g920_n_spl_),
    .din2(g921_n)
  );


  FA
  g_g922_n
  (
    .dout(g922_n),
    .din1(g920_p_spl_),
    .din2(g921_p)
  );


  LA
  g_g923_p
  (
    .dout(g923_p),
    .din1(g841_n_spl_),
    .din2(g922_p_spl_)
  );


  FA
  g_g923_n
  (
    .dout(g923_n),
    .din1(g841_p_spl_),
    .din2(g922_n_spl_)
  );


  LA
  g_g924_p
  (
    .dout(g924_p),
    .din1(g841_p_spl_),
    .din2(g922_n_spl_)
  );


  FA
  g_g924_n
  (
    .dout(g924_n),
    .din1(g841_n_spl_),
    .din2(g922_p_spl_)
  );


  LA
  g_g925_p
  (
    .dout(g925_p),
    .din1(g923_n_spl_),
    .din2(g924_n)
  );


  FA
  g_g925_n
  (
    .dout(g925_n),
    .din1(g923_p_spl_),
    .din2(g924_p)
  );


  LA
  g_g926_p
  (
    .dout(g926_p),
    .din1(g840_n_spl_),
    .din2(g925_p_spl_)
  );


  FA
  g_g926_n
  (
    .dout(g926_n),
    .din1(g840_p_spl_),
    .din2(g925_n_spl_)
  );


  LA
  g_g927_p
  (
    .dout(g927_p),
    .din1(g840_p_spl_),
    .din2(g925_n_spl_)
  );


  FA
  g_g927_n
  (
    .dout(g927_n),
    .din1(g840_n_spl_),
    .din2(g925_p_spl_)
  );


  LA
  g_g928_p
  (
    .dout(g928_p),
    .din1(g926_n_spl_),
    .din2(g927_n)
  );


  FA
  g_g928_n
  (
    .dout(g928_n),
    .din1(g926_p_spl_),
    .din2(g927_p)
  );


  LA
  g_g929_p
  (
    .dout(g929_p),
    .din1(g839_n_spl_),
    .din2(g928_p_spl_)
  );


  FA
  g_g929_n
  (
    .dout(g929_n),
    .din1(g839_p_spl_),
    .din2(g928_n_spl_)
  );


  LA
  g_g930_p
  (
    .dout(g930_p),
    .din1(g839_p_spl_),
    .din2(g928_n_spl_)
  );


  FA
  g_g930_n
  (
    .dout(g930_n),
    .din1(g839_n_spl_),
    .din2(g928_p_spl_)
  );


  LA
  g_g931_p
  (
    .dout(g931_p),
    .din1(g929_n_spl_),
    .din2(g930_n)
  );


  FA
  g_g931_n
  (
    .dout(g931_n),
    .din1(g929_p_spl_),
    .din2(g930_p)
  );


  LA
  g_g932_p
  (
    .dout(g932_p),
    .din1(g838_n_spl_),
    .din2(g931_p_spl_)
  );


  FA
  g_g932_n
  (
    .dout(g932_n),
    .din1(g838_p_spl_),
    .din2(g931_n_spl_)
  );


  LA
  g_g933_p
  (
    .dout(g933_p),
    .din1(g838_p_spl_),
    .din2(g931_n_spl_)
  );


  FA
  g_g933_n
  (
    .dout(g933_n),
    .din1(g838_n_spl_),
    .din2(g931_p_spl_)
  );


  LA
  g_g934_p
  (
    .dout(g934_p),
    .din1(g932_n_spl_),
    .din2(g933_n)
  );


  FA
  g_g934_n
  (
    .dout(g934_n),
    .din1(g932_p_spl_),
    .din2(g933_p)
  );


  LA
  g_g935_p
  (
    .dout(g935_p),
    .din1(g837_n_spl_),
    .din2(g934_p_spl_)
  );


  FA
  g_g935_n
  (
    .dout(g935_n),
    .din1(g837_p_spl_),
    .din2(g934_n_spl_)
  );


  LA
  g_g936_p
  (
    .dout(g936_p),
    .din1(g837_p_spl_),
    .din2(g934_n_spl_)
  );


  FA
  g_g936_n
  (
    .dout(g936_n),
    .din1(g837_n_spl_),
    .din2(g934_p_spl_)
  );


  LA
  g_g937_p
  (
    .dout(g937_p),
    .din1(g935_n_spl_),
    .din2(g936_n)
  );


  FA
  g_g937_n
  (
    .dout(g937_n),
    .din1(g935_p_spl_),
    .din2(g936_p)
  );


  LA
  g_g938_p
  (
    .dout(g938_p),
    .din1(g836_n_spl_),
    .din2(g937_p_spl_)
  );


  FA
  g_g938_n
  (
    .dout(g938_n),
    .din1(g836_p_spl_),
    .din2(g937_n_spl_)
  );


  LA
  g_g939_p
  (
    .dout(g939_p),
    .din1(g836_p_spl_),
    .din2(g937_n_spl_)
  );


  FA
  g_g939_n
  (
    .dout(g939_n),
    .din1(g836_n_spl_),
    .din2(g937_p_spl_)
  );


  LA
  g_g940_p
  (
    .dout(g940_p),
    .din1(g938_n_spl_),
    .din2(g939_n)
  );


  FA
  g_g940_n
  (
    .dout(g940_n),
    .din1(g938_p_spl_),
    .din2(g939_p)
  );


  LA
  g_g941_p
  (
    .dout(g941_p),
    .din1(g835_n_spl_),
    .din2(g940_p_spl_)
  );


  FA
  g_g941_n
  (
    .dout(g941_n),
    .din1(g835_p_spl_),
    .din2(g940_n_spl_)
  );


  LA
  g_g942_p
  (
    .dout(g942_p),
    .din1(g835_p_spl_),
    .din2(g940_n_spl_)
  );


  FA
  g_g942_n
  (
    .dout(g942_n),
    .din1(g835_n_spl_),
    .din2(g940_p_spl_)
  );


  LA
  g_g943_p
  (
    .dout(g943_p),
    .din1(g941_n_spl_),
    .din2(g942_n)
  );


  FA
  g_g943_n
  (
    .dout(g943_n),
    .din1(g941_p_spl_),
    .din2(g942_p)
  );


  LA
  g_g944_p
  (
    .dout(g944_p),
    .din1(g834_n_spl_),
    .din2(g943_p_spl_)
  );


  FA
  g_g944_n
  (
    .dout(g944_n),
    .din1(g834_p_spl_),
    .din2(g943_n_spl_)
  );


  LA
  g_g945_p
  (
    .dout(g945_p),
    .din1(g834_p_spl_),
    .din2(g943_n_spl_)
  );


  FA
  g_g945_n
  (
    .dout(g945_n),
    .din1(g834_n_spl_),
    .din2(g943_p_spl_)
  );


  LA
  g_g946_p
  (
    .dout(g946_p),
    .din1(g944_n_spl_),
    .din2(g945_n)
  );


  FA
  g_g946_n
  (
    .dout(g946_n),
    .din1(g944_p_spl_),
    .din2(g945_p)
  );


  LA
  g_g947_p
  (
    .dout(g947_p),
    .din1(g833_n),
    .din2(g946_p)
  );


  FA
  g_g947_n
  (
    .dout(g947_n),
    .din1(g833_p_spl_),
    .din2(g946_n_spl_)
  );


  LA
  g_g948_p
  (
    .dout(g948_p),
    .din1(g833_p_spl_),
    .din2(g946_n_spl_)
  );


  FA
  g_g949_n
  (
    .dout(g949_n),
    .din1(g947_p_spl_),
    .din2(g948_p)
  );


  LA
  g_g950_p
  (
    .dout(g950_p),
    .din1(g944_n_spl_),
    .din2(g947_n)
  );


  FA
  g_g950_n
  (
    .dout(g950_n),
    .din1(g944_p_spl_),
    .din2(g947_p_spl_)
  );


  LA
  g_g951_p
  (
    .dout(g951_p),
    .din1(G2_p_spl_111),
    .din2(G32_p_spl_000)
  );


  FA
  g_g951_n
  (
    .dout(g951_n),
    .din1(G2_n_spl_111),
    .din2(G32_n_spl_000)
  );


  LA
  g_g952_p
  (
    .dout(g952_p),
    .din1(g938_n_spl_),
    .din2(g941_n_spl_)
  );


  FA
  g_g952_n
  (
    .dout(g952_n),
    .din1(g938_p_spl_),
    .din2(g941_p_spl_)
  );


  LA
  g_g953_p
  (
    .dout(g953_p),
    .din1(G3_p_spl_111),
    .din2(G31_p_spl_001)
  );


  FA
  g_g953_n
  (
    .dout(g953_n),
    .din1(G3_n_spl_111),
    .din2(G31_n_spl_001)
  );


  LA
  g_g954_p
  (
    .dout(g954_p),
    .din1(g932_n_spl_),
    .din2(g935_n_spl_)
  );


  FA
  g_g954_n
  (
    .dout(g954_n),
    .din1(g932_p_spl_),
    .din2(g935_p_spl_)
  );


  LA
  g_g955_p
  (
    .dout(g955_p),
    .din1(G4_p_spl_110),
    .din2(G30_p_spl_001)
  );


  FA
  g_g955_n
  (
    .dout(g955_n),
    .din1(G4_n_spl_110),
    .din2(G30_n_spl_001)
  );


  LA
  g_g956_p
  (
    .dout(g956_p),
    .din1(g926_n_spl_),
    .din2(g929_n_spl_)
  );


  FA
  g_g956_n
  (
    .dout(g956_n),
    .din1(g926_p_spl_),
    .din2(g929_p_spl_)
  );


  LA
  g_g957_p
  (
    .dout(g957_p),
    .din1(G5_p_spl_110),
    .din2(G29_p_spl_010)
  );


  FA
  g_g957_n
  (
    .dout(g957_n),
    .din1(G5_n_spl_110),
    .din2(G29_n_spl_010)
  );


  LA
  g_g958_p
  (
    .dout(g958_p),
    .din1(g920_n_spl_),
    .din2(g923_n_spl_)
  );


  FA
  g_g958_n
  (
    .dout(g958_n),
    .din1(g920_p_spl_),
    .din2(g923_p_spl_)
  );


  LA
  g_g959_p
  (
    .dout(g959_p),
    .din1(G6_p_spl_101),
    .din2(G28_p_spl_010)
  );


  FA
  g_g959_n
  (
    .dout(g959_n),
    .din1(G6_n_spl_101),
    .din2(G28_n_spl_010)
  );


  LA
  g_g960_p
  (
    .dout(g960_p),
    .din1(g914_n_spl_),
    .din2(g917_n_spl_)
  );


  FA
  g_g960_n
  (
    .dout(g960_n),
    .din1(g914_p_spl_),
    .din2(g917_p_spl_)
  );


  LA
  g_g961_p
  (
    .dout(g961_p),
    .din1(G7_p_spl_101),
    .din2(G27_p_spl_011)
  );


  FA
  g_g961_n
  (
    .dout(g961_n),
    .din1(G7_n_spl_101),
    .din2(G27_n_spl_011)
  );


  LA
  g_g962_p
  (
    .dout(g962_p),
    .din1(g908_n_spl_),
    .din2(g911_n_spl_)
  );


  FA
  g_g962_n
  (
    .dout(g962_n),
    .din1(g908_p_spl_),
    .din2(g911_p_spl_)
  );


  LA
  g_g963_p
  (
    .dout(g963_p),
    .din1(G8_p_spl_100),
    .din2(G26_p_spl_011)
  );


  FA
  g_g963_n
  (
    .dout(g963_n),
    .din1(G8_n_spl_100),
    .din2(G26_n_spl_011)
  );


  LA
  g_g964_p
  (
    .dout(g964_p),
    .din1(g902_n_spl_),
    .din2(g905_n_spl_)
  );


  FA
  g_g964_n
  (
    .dout(g964_n),
    .din1(g902_p_spl_),
    .din2(g905_p_spl_)
  );


  LA
  g_g965_p
  (
    .dout(g965_p),
    .din1(G9_p_spl_100),
    .din2(G25_p_spl_100)
  );


  FA
  g_g965_n
  (
    .dout(g965_n),
    .din1(G9_n_spl_100),
    .din2(G25_n_spl_100)
  );


  LA
  g_g966_p
  (
    .dout(g966_p),
    .din1(g896_n_spl_),
    .din2(g899_n_spl_)
  );


  FA
  g_g966_n
  (
    .dout(g966_n),
    .din1(g896_p_spl_),
    .din2(g899_p_spl_)
  );


  LA
  g_g967_p
  (
    .dout(g967_p),
    .din1(G10_p_spl_011),
    .din2(G24_p_spl_100)
  );


  FA
  g_g967_n
  (
    .dout(g967_n),
    .din1(G10_n_spl_011),
    .din2(G24_n_spl_100)
  );


  LA
  g_g968_p
  (
    .dout(g968_p),
    .din1(g890_n_spl_),
    .din2(g893_n_spl_)
  );


  FA
  g_g968_n
  (
    .dout(g968_n),
    .din1(g890_p_spl_),
    .din2(g893_p_spl_)
  );


  LA
  g_g969_p
  (
    .dout(g969_p),
    .din1(G11_p_spl_011),
    .din2(G23_p_spl_101)
  );


  FA
  g_g969_n
  (
    .dout(g969_n),
    .din1(G11_n_spl_011),
    .din2(G23_n_spl_101)
  );


  LA
  g_g970_p
  (
    .dout(g970_p),
    .din1(g884_n_spl_),
    .din2(g887_n_spl_)
  );


  FA
  g_g970_n
  (
    .dout(g970_n),
    .din1(g884_p_spl_),
    .din2(g887_p_spl_)
  );


  LA
  g_g971_p
  (
    .dout(g971_p),
    .din1(G12_p_spl_010),
    .din2(G22_p_spl_101)
  );


  FA
  g_g971_n
  (
    .dout(g971_n),
    .din1(G12_n_spl_010),
    .din2(G22_n_spl_101)
  );


  LA
  g_g972_p
  (
    .dout(g972_p),
    .din1(g878_n_spl_),
    .din2(g881_n_spl_)
  );


  FA
  g_g972_n
  (
    .dout(g972_n),
    .din1(g878_p_spl_),
    .din2(g881_p_spl_)
  );


  LA
  g_g973_p
  (
    .dout(g973_p),
    .din1(G13_p_spl_010),
    .din2(G21_p_spl_110)
  );


  FA
  g_g973_n
  (
    .dout(g973_n),
    .din1(G13_n_spl_010),
    .din2(G21_n_spl_110)
  );


  LA
  g_g974_p
  (
    .dout(g974_p),
    .din1(g872_n_spl_),
    .din2(g875_n_spl_)
  );


  FA
  g_g974_n
  (
    .dout(g974_n),
    .din1(g872_p_spl_),
    .din2(g875_p_spl_)
  );


  LA
  g_g975_p
  (
    .dout(g975_p),
    .din1(G14_p_spl_001),
    .din2(G20_p_spl_110)
  );


  FA
  g_g975_n
  (
    .dout(g975_n),
    .din1(G14_n_spl_001),
    .din2(G20_n_spl_110)
  );


  LA
  g_g976_p
  (
    .dout(g976_p),
    .din1(g866_n_spl_),
    .din2(g869_n_spl_)
  );


  FA
  g_g976_n
  (
    .dout(g976_n),
    .din1(g866_p_spl_),
    .din2(g869_p_spl_)
  );


  LA
  g_g977_p
  (
    .dout(g977_p),
    .din1(G16_p_spl_000),
    .din2(G18_p_spl_111)
  );


  FA
  g_g977_n
  (
    .dout(g977_n),
    .din1(G16_n_spl_000),
    .din2(G18_n_spl_111)
  );


  LA
  g_g978_p
  (
    .dout(g978_p),
    .din1(g863_n_spl_),
    .din2(g977_p_spl_)
  );


  FA
  g_g978_n
  (
    .dout(g978_n),
    .din1(g863_p_spl_),
    .din2(g977_n_spl_)
  );


  LA
  g_g979_p
  (
    .dout(g979_p),
    .din1(G15_p_spl_001),
    .din2(G19_p_spl_111)
  );


  FA
  g_g979_n
  (
    .dout(g979_n),
    .din1(G15_n_spl_001),
    .din2(G19_n_spl_111)
  );


  LA
  g_g980_p
  (
    .dout(g980_p),
    .din1(g978_p_spl_),
    .din2(g979_n_spl_)
  );


  FA
  g_g980_n
  (
    .dout(g980_n),
    .din1(g978_n_spl_),
    .din2(g979_p_spl_)
  );


  LA
  g_g981_p
  (
    .dout(g981_p),
    .din1(g978_n_spl_),
    .din2(g979_p_spl_)
  );


  FA
  g_g981_n
  (
    .dout(g981_n),
    .din1(g978_p_spl_),
    .din2(g979_n_spl_)
  );


  LA
  g_g982_p
  (
    .dout(g982_p),
    .din1(g980_n_spl_),
    .din2(g981_n)
  );


  FA
  g_g982_n
  (
    .dout(g982_n),
    .din1(g980_p_spl_),
    .din2(g981_p)
  );


  LA
  g_g983_p
  (
    .dout(g983_p),
    .din1(g976_n_spl_),
    .din2(g982_p_spl_)
  );


  FA
  g_g983_n
  (
    .dout(g983_n),
    .din1(g976_p_spl_),
    .din2(g982_n_spl_)
  );


  LA
  g_g984_p
  (
    .dout(g984_p),
    .din1(g976_p_spl_),
    .din2(g982_n_spl_)
  );


  FA
  g_g984_n
  (
    .dout(g984_n),
    .din1(g976_n_spl_),
    .din2(g982_p_spl_)
  );


  LA
  g_g985_p
  (
    .dout(g985_p),
    .din1(g983_n_spl_),
    .din2(g984_n)
  );


  FA
  g_g985_n
  (
    .dout(g985_n),
    .din1(g983_p_spl_),
    .din2(g984_p)
  );


  LA
  g_g986_p
  (
    .dout(g986_p),
    .din1(g975_n_spl_),
    .din2(g985_p_spl_)
  );


  FA
  g_g986_n
  (
    .dout(g986_n),
    .din1(g975_p_spl_),
    .din2(g985_n_spl_)
  );


  LA
  g_g987_p
  (
    .dout(g987_p),
    .din1(g975_p_spl_),
    .din2(g985_n_spl_)
  );


  FA
  g_g987_n
  (
    .dout(g987_n),
    .din1(g975_n_spl_),
    .din2(g985_p_spl_)
  );


  LA
  g_g988_p
  (
    .dout(g988_p),
    .din1(g986_n_spl_),
    .din2(g987_n)
  );


  FA
  g_g988_n
  (
    .dout(g988_n),
    .din1(g986_p_spl_),
    .din2(g987_p)
  );


  LA
  g_g989_p
  (
    .dout(g989_p),
    .din1(g974_n_spl_),
    .din2(g988_p_spl_)
  );


  FA
  g_g989_n
  (
    .dout(g989_n),
    .din1(g974_p_spl_),
    .din2(g988_n_spl_)
  );


  LA
  g_g990_p
  (
    .dout(g990_p),
    .din1(g974_p_spl_),
    .din2(g988_n_spl_)
  );


  FA
  g_g990_n
  (
    .dout(g990_n),
    .din1(g974_n_spl_),
    .din2(g988_p_spl_)
  );


  LA
  g_g991_p
  (
    .dout(g991_p),
    .din1(g989_n_spl_),
    .din2(g990_n)
  );


  FA
  g_g991_n
  (
    .dout(g991_n),
    .din1(g989_p_spl_),
    .din2(g990_p)
  );


  LA
  g_g992_p
  (
    .dout(g992_p),
    .din1(g973_n_spl_),
    .din2(g991_p_spl_)
  );


  FA
  g_g992_n
  (
    .dout(g992_n),
    .din1(g973_p_spl_),
    .din2(g991_n_spl_)
  );


  LA
  g_g993_p
  (
    .dout(g993_p),
    .din1(g973_p_spl_),
    .din2(g991_n_spl_)
  );


  FA
  g_g993_n
  (
    .dout(g993_n),
    .din1(g973_n_spl_),
    .din2(g991_p_spl_)
  );


  LA
  g_g994_p
  (
    .dout(g994_p),
    .din1(g992_n_spl_),
    .din2(g993_n)
  );


  FA
  g_g994_n
  (
    .dout(g994_n),
    .din1(g992_p_spl_),
    .din2(g993_p)
  );


  LA
  g_g995_p
  (
    .dout(g995_p),
    .din1(g972_n_spl_),
    .din2(g994_p_spl_)
  );


  FA
  g_g995_n
  (
    .dout(g995_n),
    .din1(g972_p_spl_),
    .din2(g994_n_spl_)
  );


  LA
  g_g996_p
  (
    .dout(g996_p),
    .din1(g972_p_spl_),
    .din2(g994_n_spl_)
  );


  FA
  g_g996_n
  (
    .dout(g996_n),
    .din1(g972_n_spl_),
    .din2(g994_p_spl_)
  );


  LA
  g_g997_p
  (
    .dout(g997_p),
    .din1(g995_n_spl_),
    .din2(g996_n)
  );


  FA
  g_g997_n
  (
    .dout(g997_n),
    .din1(g995_p_spl_),
    .din2(g996_p)
  );


  LA
  g_g998_p
  (
    .dout(g998_p),
    .din1(g971_n_spl_),
    .din2(g997_p_spl_)
  );


  FA
  g_g998_n
  (
    .dout(g998_n),
    .din1(g971_p_spl_),
    .din2(g997_n_spl_)
  );


  LA
  g_g999_p
  (
    .dout(g999_p),
    .din1(g971_p_spl_),
    .din2(g997_n_spl_)
  );


  FA
  g_g999_n
  (
    .dout(g999_n),
    .din1(g971_n_spl_),
    .din2(g997_p_spl_)
  );


  LA
  g_g1000_p
  (
    .dout(g1000_p),
    .din1(g998_n_spl_),
    .din2(g999_n)
  );


  FA
  g_g1000_n
  (
    .dout(g1000_n),
    .din1(g998_p_spl_),
    .din2(g999_p)
  );


  LA
  g_g1001_p
  (
    .dout(g1001_p),
    .din1(g970_n_spl_),
    .din2(g1000_p_spl_)
  );


  FA
  g_g1001_n
  (
    .dout(g1001_n),
    .din1(g970_p_spl_),
    .din2(g1000_n_spl_)
  );


  LA
  g_g1002_p
  (
    .dout(g1002_p),
    .din1(g970_p_spl_),
    .din2(g1000_n_spl_)
  );


  FA
  g_g1002_n
  (
    .dout(g1002_n),
    .din1(g970_n_spl_),
    .din2(g1000_p_spl_)
  );


  LA
  g_g1003_p
  (
    .dout(g1003_p),
    .din1(g1001_n_spl_),
    .din2(g1002_n)
  );


  FA
  g_g1003_n
  (
    .dout(g1003_n),
    .din1(g1001_p_spl_),
    .din2(g1002_p)
  );


  LA
  g_g1004_p
  (
    .dout(g1004_p),
    .din1(g969_n_spl_),
    .din2(g1003_p_spl_)
  );


  FA
  g_g1004_n
  (
    .dout(g1004_n),
    .din1(g969_p_spl_),
    .din2(g1003_n_spl_)
  );


  LA
  g_g1005_p
  (
    .dout(g1005_p),
    .din1(g969_p_spl_),
    .din2(g1003_n_spl_)
  );


  FA
  g_g1005_n
  (
    .dout(g1005_n),
    .din1(g969_n_spl_),
    .din2(g1003_p_spl_)
  );


  LA
  g_g1006_p
  (
    .dout(g1006_p),
    .din1(g1004_n_spl_),
    .din2(g1005_n)
  );


  FA
  g_g1006_n
  (
    .dout(g1006_n),
    .din1(g1004_p_spl_),
    .din2(g1005_p)
  );


  LA
  g_g1007_p
  (
    .dout(g1007_p),
    .din1(g968_n_spl_),
    .din2(g1006_p_spl_)
  );


  FA
  g_g1007_n
  (
    .dout(g1007_n),
    .din1(g968_p_spl_),
    .din2(g1006_n_spl_)
  );


  LA
  g_g1008_p
  (
    .dout(g1008_p),
    .din1(g968_p_spl_),
    .din2(g1006_n_spl_)
  );


  FA
  g_g1008_n
  (
    .dout(g1008_n),
    .din1(g968_n_spl_),
    .din2(g1006_p_spl_)
  );


  LA
  g_g1009_p
  (
    .dout(g1009_p),
    .din1(g1007_n_spl_),
    .din2(g1008_n)
  );


  FA
  g_g1009_n
  (
    .dout(g1009_n),
    .din1(g1007_p_spl_),
    .din2(g1008_p)
  );


  LA
  g_g1010_p
  (
    .dout(g1010_p),
    .din1(g967_n_spl_),
    .din2(g1009_p_spl_)
  );


  FA
  g_g1010_n
  (
    .dout(g1010_n),
    .din1(g967_p_spl_),
    .din2(g1009_n_spl_)
  );


  LA
  g_g1011_p
  (
    .dout(g1011_p),
    .din1(g967_p_spl_),
    .din2(g1009_n_spl_)
  );


  FA
  g_g1011_n
  (
    .dout(g1011_n),
    .din1(g967_n_spl_),
    .din2(g1009_p_spl_)
  );


  LA
  g_g1012_p
  (
    .dout(g1012_p),
    .din1(g1010_n_spl_),
    .din2(g1011_n)
  );


  FA
  g_g1012_n
  (
    .dout(g1012_n),
    .din1(g1010_p_spl_),
    .din2(g1011_p)
  );


  LA
  g_g1013_p
  (
    .dout(g1013_p),
    .din1(g966_n_spl_),
    .din2(g1012_p_spl_)
  );


  FA
  g_g1013_n
  (
    .dout(g1013_n),
    .din1(g966_p_spl_),
    .din2(g1012_n_spl_)
  );


  LA
  g_g1014_p
  (
    .dout(g1014_p),
    .din1(g966_p_spl_),
    .din2(g1012_n_spl_)
  );


  FA
  g_g1014_n
  (
    .dout(g1014_n),
    .din1(g966_n_spl_),
    .din2(g1012_p_spl_)
  );


  LA
  g_g1015_p
  (
    .dout(g1015_p),
    .din1(g1013_n_spl_),
    .din2(g1014_n)
  );


  FA
  g_g1015_n
  (
    .dout(g1015_n),
    .din1(g1013_p_spl_),
    .din2(g1014_p)
  );


  LA
  g_g1016_p
  (
    .dout(g1016_p),
    .din1(g965_n_spl_),
    .din2(g1015_p_spl_)
  );


  FA
  g_g1016_n
  (
    .dout(g1016_n),
    .din1(g965_p_spl_),
    .din2(g1015_n_spl_)
  );


  LA
  g_g1017_p
  (
    .dout(g1017_p),
    .din1(g965_p_spl_),
    .din2(g1015_n_spl_)
  );


  FA
  g_g1017_n
  (
    .dout(g1017_n),
    .din1(g965_n_spl_),
    .din2(g1015_p_spl_)
  );


  LA
  g_g1018_p
  (
    .dout(g1018_p),
    .din1(g1016_n_spl_),
    .din2(g1017_n)
  );


  FA
  g_g1018_n
  (
    .dout(g1018_n),
    .din1(g1016_p_spl_),
    .din2(g1017_p)
  );


  LA
  g_g1019_p
  (
    .dout(g1019_p),
    .din1(g964_n_spl_),
    .din2(g1018_p_spl_)
  );


  FA
  g_g1019_n
  (
    .dout(g1019_n),
    .din1(g964_p_spl_),
    .din2(g1018_n_spl_)
  );


  LA
  g_g1020_p
  (
    .dout(g1020_p),
    .din1(g964_p_spl_),
    .din2(g1018_n_spl_)
  );


  FA
  g_g1020_n
  (
    .dout(g1020_n),
    .din1(g964_n_spl_),
    .din2(g1018_p_spl_)
  );


  LA
  g_g1021_p
  (
    .dout(g1021_p),
    .din1(g1019_n_spl_),
    .din2(g1020_n)
  );


  FA
  g_g1021_n
  (
    .dout(g1021_n),
    .din1(g1019_p_spl_),
    .din2(g1020_p)
  );


  LA
  g_g1022_p
  (
    .dout(g1022_p),
    .din1(g963_n_spl_),
    .din2(g1021_p_spl_)
  );


  FA
  g_g1022_n
  (
    .dout(g1022_n),
    .din1(g963_p_spl_),
    .din2(g1021_n_spl_)
  );


  LA
  g_g1023_p
  (
    .dout(g1023_p),
    .din1(g963_p_spl_),
    .din2(g1021_n_spl_)
  );


  FA
  g_g1023_n
  (
    .dout(g1023_n),
    .din1(g963_n_spl_),
    .din2(g1021_p_spl_)
  );


  LA
  g_g1024_p
  (
    .dout(g1024_p),
    .din1(g1022_n_spl_),
    .din2(g1023_n)
  );


  FA
  g_g1024_n
  (
    .dout(g1024_n),
    .din1(g1022_p_spl_),
    .din2(g1023_p)
  );


  LA
  g_g1025_p
  (
    .dout(g1025_p),
    .din1(g962_n_spl_),
    .din2(g1024_p_spl_)
  );


  FA
  g_g1025_n
  (
    .dout(g1025_n),
    .din1(g962_p_spl_),
    .din2(g1024_n_spl_)
  );


  LA
  g_g1026_p
  (
    .dout(g1026_p),
    .din1(g962_p_spl_),
    .din2(g1024_n_spl_)
  );


  FA
  g_g1026_n
  (
    .dout(g1026_n),
    .din1(g962_n_spl_),
    .din2(g1024_p_spl_)
  );


  LA
  g_g1027_p
  (
    .dout(g1027_p),
    .din1(g1025_n_spl_),
    .din2(g1026_n)
  );


  FA
  g_g1027_n
  (
    .dout(g1027_n),
    .din1(g1025_p_spl_),
    .din2(g1026_p)
  );


  LA
  g_g1028_p
  (
    .dout(g1028_p),
    .din1(g961_n_spl_),
    .din2(g1027_p_spl_)
  );


  FA
  g_g1028_n
  (
    .dout(g1028_n),
    .din1(g961_p_spl_),
    .din2(g1027_n_spl_)
  );


  LA
  g_g1029_p
  (
    .dout(g1029_p),
    .din1(g961_p_spl_),
    .din2(g1027_n_spl_)
  );


  FA
  g_g1029_n
  (
    .dout(g1029_n),
    .din1(g961_n_spl_),
    .din2(g1027_p_spl_)
  );


  LA
  g_g1030_p
  (
    .dout(g1030_p),
    .din1(g1028_n_spl_),
    .din2(g1029_n)
  );


  FA
  g_g1030_n
  (
    .dout(g1030_n),
    .din1(g1028_p_spl_),
    .din2(g1029_p)
  );


  LA
  g_g1031_p
  (
    .dout(g1031_p),
    .din1(g960_n_spl_),
    .din2(g1030_p_spl_)
  );


  FA
  g_g1031_n
  (
    .dout(g1031_n),
    .din1(g960_p_spl_),
    .din2(g1030_n_spl_)
  );


  LA
  g_g1032_p
  (
    .dout(g1032_p),
    .din1(g960_p_spl_),
    .din2(g1030_n_spl_)
  );


  FA
  g_g1032_n
  (
    .dout(g1032_n),
    .din1(g960_n_spl_),
    .din2(g1030_p_spl_)
  );


  LA
  g_g1033_p
  (
    .dout(g1033_p),
    .din1(g1031_n_spl_),
    .din2(g1032_n)
  );


  FA
  g_g1033_n
  (
    .dout(g1033_n),
    .din1(g1031_p_spl_),
    .din2(g1032_p)
  );


  LA
  g_g1034_p
  (
    .dout(g1034_p),
    .din1(g959_n_spl_),
    .din2(g1033_p_spl_)
  );


  FA
  g_g1034_n
  (
    .dout(g1034_n),
    .din1(g959_p_spl_),
    .din2(g1033_n_spl_)
  );


  LA
  g_g1035_p
  (
    .dout(g1035_p),
    .din1(g959_p_spl_),
    .din2(g1033_n_spl_)
  );


  FA
  g_g1035_n
  (
    .dout(g1035_n),
    .din1(g959_n_spl_),
    .din2(g1033_p_spl_)
  );


  LA
  g_g1036_p
  (
    .dout(g1036_p),
    .din1(g1034_n_spl_),
    .din2(g1035_n)
  );


  FA
  g_g1036_n
  (
    .dout(g1036_n),
    .din1(g1034_p_spl_),
    .din2(g1035_p)
  );


  LA
  g_g1037_p
  (
    .dout(g1037_p),
    .din1(g958_n_spl_),
    .din2(g1036_p_spl_)
  );


  FA
  g_g1037_n
  (
    .dout(g1037_n),
    .din1(g958_p_spl_),
    .din2(g1036_n_spl_)
  );


  LA
  g_g1038_p
  (
    .dout(g1038_p),
    .din1(g958_p_spl_),
    .din2(g1036_n_spl_)
  );


  FA
  g_g1038_n
  (
    .dout(g1038_n),
    .din1(g958_n_spl_),
    .din2(g1036_p_spl_)
  );


  LA
  g_g1039_p
  (
    .dout(g1039_p),
    .din1(g1037_n_spl_),
    .din2(g1038_n)
  );


  FA
  g_g1039_n
  (
    .dout(g1039_n),
    .din1(g1037_p_spl_),
    .din2(g1038_p)
  );


  LA
  g_g1040_p
  (
    .dout(g1040_p),
    .din1(g957_n_spl_),
    .din2(g1039_p_spl_)
  );


  FA
  g_g1040_n
  (
    .dout(g1040_n),
    .din1(g957_p_spl_),
    .din2(g1039_n_spl_)
  );


  LA
  g_g1041_p
  (
    .dout(g1041_p),
    .din1(g957_p_spl_),
    .din2(g1039_n_spl_)
  );


  FA
  g_g1041_n
  (
    .dout(g1041_n),
    .din1(g957_n_spl_),
    .din2(g1039_p_spl_)
  );


  LA
  g_g1042_p
  (
    .dout(g1042_p),
    .din1(g1040_n_spl_),
    .din2(g1041_n)
  );


  FA
  g_g1042_n
  (
    .dout(g1042_n),
    .din1(g1040_p_spl_),
    .din2(g1041_p)
  );


  LA
  g_g1043_p
  (
    .dout(g1043_p),
    .din1(g956_n_spl_),
    .din2(g1042_p_spl_)
  );


  FA
  g_g1043_n
  (
    .dout(g1043_n),
    .din1(g956_p_spl_),
    .din2(g1042_n_spl_)
  );


  LA
  g_g1044_p
  (
    .dout(g1044_p),
    .din1(g956_p_spl_),
    .din2(g1042_n_spl_)
  );


  FA
  g_g1044_n
  (
    .dout(g1044_n),
    .din1(g956_n_spl_),
    .din2(g1042_p_spl_)
  );


  LA
  g_g1045_p
  (
    .dout(g1045_p),
    .din1(g1043_n_spl_),
    .din2(g1044_n)
  );


  FA
  g_g1045_n
  (
    .dout(g1045_n),
    .din1(g1043_p_spl_),
    .din2(g1044_p)
  );


  LA
  g_g1046_p
  (
    .dout(g1046_p),
    .din1(g955_n_spl_),
    .din2(g1045_p_spl_)
  );


  FA
  g_g1046_n
  (
    .dout(g1046_n),
    .din1(g955_p_spl_),
    .din2(g1045_n_spl_)
  );


  LA
  g_g1047_p
  (
    .dout(g1047_p),
    .din1(g955_p_spl_),
    .din2(g1045_n_spl_)
  );


  FA
  g_g1047_n
  (
    .dout(g1047_n),
    .din1(g955_n_spl_),
    .din2(g1045_p_spl_)
  );


  LA
  g_g1048_p
  (
    .dout(g1048_p),
    .din1(g1046_n_spl_),
    .din2(g1047_n)
  );


  FA
  g_g1048_n
  (
    .dout(g1048_n),
    .din1(g1046_p_spl_),
    .din2(g1047_p)
  );


  LA
  g_g1049_p
  (
    .dout(g1049_p),
    .din1(g954_n_spl_),
    .din2(g1048_p_spl_)
  );


  FA
  g_g1049_n
  (
    .dout(g1049_n),
    .din1(g954_p_spl_),
    .din2(g1048_n_spl_)
  );


  LA
  g_g1050_p
  (
    .dout(g1050_p),
    .din1(g954_p_spl_),
    .din2(g1048_n_spl_)
  );


  FA
  g_g1050_n
  (
    .dout(g1050_n),
    .din1(g954_n_spl_),
    .din2(g1048_p_spl_)
  );


  LA
  g_g1051_p
  (
    .dout(g1051_p),
    .din1(g1049_n_spl_),
    .din2(g1050_n)
  );


  FA
  g_g1051_n
  (
    .dout(g1051_n),
    .din1(g1049_p_spl_),
    .din2(g1050_p)
  );


  LA
  g_g1052_p
  (
    .dout(g1052_p),
    .din1(g953_n_spl_),
    .din2(g1051_p_spl_)
  );


  FA
  g_g1052_n
  (
    .dout(g1052_n),
    .din1(g953_p_spl_),
    .din2(g1051_n_spl_)
  );


  LA
  g_g1053_p
  (
    .dout(g1053_p),
    .din1(g953_p_spl_),
    .din2(g1051_n_spl_)
  );


  FA
  g_g1053_n
  (
    .dout(g1053_n),
    .din1(g953_n_spl_),
    .din2(g1051_p_spl_)
  );


  LA
  g_g1054_p
  (
    .dout(g1054_p),
    .din1(g1052_n_spl_),
    .din2(g1053_n)
  );


  FA
  g_g1054_n
  (
    .dout(g1054_n),
    .din1(g1052_p_spl_),
    .din2(g1053_p)
  );


  LA
  g_g1055_p
  (
    .dout(g1055_p),
    .din1(g952_n_spl_),
    .din2(g1054_p_spl_)
  );


  FA
  g_g1055_n
  (
    .dout(g1055_n),
    .din1(g952_p_spl_),
    .din2(g1054_n_spl_)
  );


  LA
  g_g1056_p
  (
    .dout(g1056_p),
    .din1(g952_p_spl_),
    .din2(g1054_n_spl_)
  );


  FA
  g_g1056_n
  (
    .dout(g1056_n),
    .din1(g952_n_spl_),
    .din2(g1054_p_spl_)
  );


  LA
  g_g1057_p
  (
    .dout(g1057_p),
    .din1(g1055_n_spl_),
    .din2(g1056_n)
  );


  FA
  g_g1057_n
  (
    .dout(g1057_n),
    .din1(g1055_p_spl_),
    .din2(g1056_p)
  );


  LA
  g_g1058_p
  (
    .dout(g1058_p),
    .din1(g951_n_spl_),
    .din2(g1057_p_spl_)
  );


  FA
  g_g1058_n
  (
    .dout(g1058_n),
    .din1(g951_p_spl_),
    .din2(g1057_n_spl_)
  );


  LA
  g_g1059_p
  (
    .dout(g1059_p),
    .din1(g951_p_spl_),
    .din2(g1057_n_spl_)
  );


  FA
  g_g1059_n
  (
    .dout(g1059_n),
    .din1(g951_n_spl_),
    .din2(g1057_p_spl_)
  );


  LA
  g_g1060_p
  (
    .dout(g1060_p),
    .din1(g1058_n_spl_),
    .din2(g1059_n)
  );


  FA
  g_g1060_n
  (
    .dout(g1060_n),
    .din1(g1058_p_spl_),
    .din2(g1059_p)
  );


  FA
  g_g1061_n
  (
    .dout(g1061_n),
    .din1(g950_p_spl_),
    .din2(g1060_n_spl_)
  );


  LA
  g_g1062_p
  (
    .dout(g1062_p),
    .din1(g950_p_spl_),
    .din2(g1060_n_spl_)
  );


  FA
  g_g1062_n
  (
    .dout(g1062_n),
    .din1(g950_n),
    .din2(g1060_p)
  );


  LA
  g_g1063_p
  (
    .dout(g1063_p),
    .din1(g1061_n),
    .din2(g1062_n_spl_)
  );


  LA
  g_g1064_p
  (
    .dout(g1064_p),
    .din1(g1055_n_spl_),
    .din2(g1058_n_spl_)
  );


  FA
  g_g1064_n
  (
    .dout(g1064_n),
    .din1(g1055_p_spl_),
    .din2(g1058_p_spl_)
  );


  LA
  g_g1065_p
  (
    .dout(g1065_p),
    .din1(G3_p_spl_111),
    .din2(G32_p_spl_001)
  );


  FA
  g_g1065_n
  (
    .dout(g1065_n),
    .din1(G3_n_spl_111),
    .din2(G32_n_spl_001)
  );


  LA
  g_g1066_p
  (
    .dout(g1066_p),
    .din1(g1049_n_spl_),
    .din2(g1052_n_spl_)
  );


  FA
  g_g1066_n
  (
    .dout(g1066_n),
    .din1(g1049_p_spl_),
    .din2(g1052_p_spl_)
  );


  LA
  g_g1067_p
  (
    .dout(g1067_p),
    .din1(G4_p_spl_111),
    .din2(G31_p_spl_001)
  );


  FA
  g_g1067_n
  (
    .dout(g1067_n),
    .din1(G4_n_spl_111),
    .din2(G31_n_spl_001)
  );


  LA
  g_g1068_p
  (
    .dout(g1068_p),
    .din1(g1043_n_spl_),
    .din2(g1046_n_spl_)
  );


  FA
  g_g1068_n
  (
    .dout(g1068_n),
    .din1(g1043_p_spl_),
    .din2(g1046_p_spl_)
  );


  LA
  g_g1069_p
  (
    .dout(g1069_p),
    .din1(G5_p_spl_110),
    .din2(G30_p_spl_010)
  );


  FA
  g_g1069_n
  (
    .dout(g1069_n),
    .din1(G5_n_spl_110),
    .din2(G30_n_spl_010)
  );


  LA
  g_g1070_p
  (
    .dout(g1070_p),
    .din1(g1037_n_spl_),
    .din2(g1040_n_spl_)
  );


  FA
  g_g1070_n
  (
    .dout(g1070_n),
    .din1(g1037_p_spl_),
    .din2(g1040_p_spl_)
  );


  LA
  g_g1071_p
  (
    .dout(g1071_p),
    .din1(G6_p_spl_110),
    .din2(G29_p_spl_010)
  );


  FA
  g_g1071_n
  (
    .dout(g1071_n),
    .din1(G6_n_spl_110),
    .din2(G29_n_spl_010)
  );


  LA
  g_g1072_p
  (
    .dout(g1072_p),
    .din1(g1031_n_spl_),
    .din2(g1034_n_spl_)
  );


  FA
  g_g1072_n
  (
    .dout(g1072_n),
    .din1(g1031_p_spl_),
    .din2(g1034_p_spl_)
  );


  LA
  g_g1073_p
  (
    .dout(g1073_p),
    .din1(G7_p_spl_101),
    .din2(G28_p_spl_011)
  );


  FA
  g_g1073_n
  (
    .dout(g1073_n),
    .din1(G7_n_spl_101),
    .din2(G28_n_spl_011)
  );


  LA
  g_g1074_p
  (
    .dout(g1074_p),
    .din1(g1025_n_spl_),
    .din2(g1028_n_spl_)
  );


  FA
  g_g1074_n
  (
    .dout(g1074_n),
    .din1(g1025_p_spl_),
    .din2(g1028_p_spl_)
  );


  LA
  g_g1075_p
  (
    .dout(g1075_p),
    .din1(G8_p_spl_101),
    .din2(G27_p_spl_011)
  );


  FA
  g_g1075_n
  (
    .dout(g1075_n),
    .din1(G8_n_spl_101),
    .din2(G27_n_spl_011)
  );


  LA
  g_g1076_p
  (
    .dout(g1076_p),
    .din1(g1019_n_spl_),
    .din2(g1022_n_spl_)
  );


  FA
  g_g1076_n
  (
    .dout(g1076_n),
    .din1(g1019_p_spl_),
    .din2(g1022_p_spl_)
  );


  LA
  g_g1077_p
  (
    .dout(g1077_p),
    .din1(G9_p_spl_100),
    .din2(G26_p_spl_100)
  );


  FA
  g_g1077_n
  (
    .dout(g1077_n),
    .din1(G9_n_spl_100),
    .din2(G26_n_spl_100)
  );


  LA
  g_g1078_p
  (
    .dout(g1078_p),
    .din1(g1013_n_spl_),
    .din2(g1016_n_spl_)
  );


  FA
  g_g1078_n
  (
    .dout(g1078_n),
    .din1(g1013_p_spl_),
    .din2(g1016_p_spl_)
  );


  LA
  g_g1079_p
  (
    .dout(g1079_p),
    .din1(G10_p_spl_100),
    .din2(G25_p_spl_100)
  );


  FA
  g_g1079_n
  (
    .dout(g1079_n),
    .din1(G10_n_spl_100),
    .din2(G25_n_spl_100)
  );


  LA
  g_g1080_p
  (
    .dout(g1080_p),
    .din1(g1007_n_spl_),
    .din2(g1010_n_spl_)
  );


  FA
  g_g1080_n
  (
    .dout(g1080_n),
    .din1(g1007_p_spl_),
    .din2(g1010_p_spl_)
  );


  LA
  g_g1081_p
  (
    .dout(g1081_p),
    .din1(G11_p_spl_011),
    .din2(G24_p_spl_101)
  );


  FA
  g_g1081_n
  (
    .dout(g1081_n),
    .din1(G11_n_spl_011),
    .din2(G24_n_spl_101)
  );


  LA
  g_g1082_p
  (
    .dout(g1082_p),
    .din1(g1001_n_spl_),
    .din2(g1004_n_spl_)
  );


  FA
  g_g1082_n
  (
    .dout(g1082_n),
    .din1(g1001_p_spl_),
    .din2(g1004_p_spl_)
  );


  LA
  g_g1083_p
  (
    .dout(g1083_p),
    .din1(G12_p_spl_011),
    .din2(G23_p_spl_101)
  );


  FA
  g_g1083_n
  (
    .dout(g1083_n),
    .din1(G12_n_spl_011),
    .din2(G23_n_spl_101)
  );


  LA
  g_g1084_p
  (
    .dout(g1084_p),
    .din1(g995_n_spl_),
    .din2(g998_n_spl_)
  );


  FA
  g_g1084_n
  (
    .dout(g1084_n),
    .din1(g995_p_spl_),
    .din2(g998_p_spl_)
  );


  LA
  g_g1085_p
  (
    .dout(g1085_p),
    .din1(G13_p_spl_010),
    .din2(G22_p_spl_110)
  );


  FA
  g_g1085_n
  (
    .dout(g1085_n),
    .din1(G13_n_spl_010),
    .din2(G22_n_spl_110)
  );


  LA
  g_g1086_p
  (
    .dout(g1086_p),
    .din1(g989_n_spl_),
    .din2(g992_n_spl_)
  );


  FA
  g_g1086_n
  (
    .dout(g1086_n),
    .din1(g989_p_spl_),
    .din2(g992_p_spl_)
  );


  LA
  g_g1087_p
  (
    .dout(g1087_p),
    .din1(G14_p_spl_010),
    .din2(G21_p_spl_110)
  );


  FA
  g_g1087_n
  (
    .dout(g1087_n),
    .din1(G14_n_spl_010),
    .din2(G21_n_spl_110)
  );


  LA
  g_g1088_p
  (
    .dout(g1088_p),
    .din1(g983_n_spl_),
    .din2(g986_n_spl_)
  );


  FA
  g_g1088_n
  (
    .dout(g1088_n),
    .din1(g983_p_spl_),
    .din2(g986_p_spl_)
  );


  LA
  g_g1089_p
  (
    .dout(g1089_p),
    .din1(G15_p_spl_001),
    .din2(G20_p_spl_111)
  );


  FA
  g_g1089_n
  (
    .dout(g1089_n),
    .din1(G15_n_spl_001),
    .din2(G20_n_spl_111)
  );


  LA
  g_g1090_p
  (
    .dout(g1090_p),
    .din1(G16_p_spl_001),
    .din2(G19_p_spl_111)
  );


  FA
  g_g1090_n
  (
    .dout(g1090_n),
    .din1(G16_n_spl_001),
    .din2(G19_n_spl_111)
  );


  LA
  g_g1091_p
  (
    .dout(g1091_p),
    .din1(g977_p_spl_),
    .din2(g980_n_spl_)
  );


  FA
  g_g1091_n
  (
    .dout(g1091_n),
    .din1(g977_n_spl_),
    .din2(g980_p_spl_)
  );


  LA
  g_g1092_p
  (
    .dout(g1092_p),
    .din1(g1090_n_spl_),
    .din2(g1091_n_spl_)
  );


  FA
  g_g1092_n
  (
    .dout(g1092_n),
    .din1(g1090_p_spl_),
    .din2(g1091_p_spl_)
  );


  LA
  g_g1093_p
  (
    .dout(g1093_p),
    .din1(g1090_p_spl_),
    .din2(g1091_p_spl_)
  );


  FA
  g_g1093_n
  (
    .dout(g1093_n),
    .din1(g1090_n_spl_),
    .din2(g1091_n_spl_)
  );


  LA
  g_g1094_p
  (
    .dout(g1094_p),
    .din1(g1092_n_spl_),
    .din2(g1093_n)
  );


  FA
  g_g1094_n
  (
    .dout(g1094_n),
    .din1(g1092_p_spl_),
    .din2(g1093_p)
  );


  LA
  g_g1095_p
  (
    .dout(g1095_p),
    .din1(g1089_n_spl_),
    .din2(g1094_p_spl_)
  );


  FA
  g_g1095_n
  (
    .dout(g1095_n),
    .din1(g1089_p_spl_),
    .din2(g1094_n_spl_)
  );


  LA
  g_g1096_p
  (
    .dout(g1096_p),
    .din1(g1089_p_spl_),
    .din2(g1094_n_spl_)
  );


  FA
  g_g1096_n
  (
    .dout(g1096_n),
    .din1(g1089_n_spl_),
    .din2(g1094_p_spl_)
  );


  LA
  g_g1097_p
  (
    .dout(g1097_p),
    .din1(g1095_n_spl_),
    .din2(g1096_n)
  );


  FA
  g_g1097_n
  (
    .dout(g1097_n),
    .din1(g1095_p_spl_),
    .din2(g1096_p)
  );


  LA
  g_g1098_p
  (
    .dout(g1098_p),
    .din1(g1088_n_spl_),
    .din2(g1097_p_spl_)
  );


  FA
  g_g1098_n
  (
    .dout(g1098_n),
    .din1(g1088_p_spl_),
    .din2(g1097_n_spl_)
  );


  LA
  g_g1099_p
  (
    .dout(g1099_p),
    .din1(g1088_p_spl_),
    .din2(g1097_n_spl_)
  );


  FA
  g_g1099_n
  (
    .dout(g1099_n),
    .din1(g1088_n_spl_),
    .din2(g1097_p_spl_)
  );


  LA
  g_g1100_p
  (
    .dout(g1100_p),
    .din1(g1098_n_spl_),
    .din2(g1099_n)
  );


  FA
  g_g1100_n
  (
    .dout(g1100_n),
    .din1(g1098_p_spl_),
    .din2(g1099_p)
  );


  LA
  g_g1101_p
  (
    .dout(g1101_p),
    .din1(g1087_n_spl_),
    .din2(g1100_p_spl_)
  );


  FA
  g_g1101_n
  (
    .dout(g1101_n),
    .din1(g1087_p_spl_),
    .din2(g1100_n_spl_)
  );


  LA
  g_g1102_p
  (
    .dout(g1102_p),
    .din1(g1087_p_spl_),
    .din2(g1100_n_spl_)
  );


  FA
  g_g1102_n
  (
    .dout(g1102_n),
    .din1(g1087_n_spl_),
    .din2(g1100_p_spl_)
  );


  LA
  g_g1103_p
  (
    .dout(g1103_p),
    .din1(g1101_n_spl_),
    .din2(g1102_n)
  );


  FA
  g_g1103_n
  (
    .dout(g1103_n),
    .din1(g1101_p_spl_),
    .din2(g1102_p)
  );


  LA
  g_g1104_p
  (
    .dout(g1104_p),
    .din1(g1086_n_spl_),
    .din2(g1103_p_spl_)
  );


  FA
  g_g1104_n
  (
    .dout(g1104_n),
    .din1(g1086_p_spl_),
    .din2(g1103_n_spl_)
  );


  LA
  g_g1105_p
  (
    .dout(g1105_p),
    .din1(g1086_p_spl_),
    .din2(g1103_n_spl_)
  );


  FA
  g_g1105_n
  (
    .dout(g1105_n),
    .din1(g1086_n_spl_),
    .din2(g1103_p_spl_)
  );


  LA
  g_g1106_p
  (
    .dout(g1106_p),
    .din1(g1104_n_spl_),
    .din2(g1105_n)
  );


  FA
  g_g1106_n
  (
    .dout(g1106_n),
    .din1(g1104_p_spl_),
    .din2(g1105_p)
  );


  LA
  g_g1107_p
  (
    .dout(g1107_p),
    .din1(g1085_n_spl_),
    .din2(g1106_p_spl_)
  );


  FA
  g_g1107_n
  (
    .dout(g1107_n),
    .din1(g1085_p_spl_),
    .din2(g1106_n_spl_)
  );


  LA
  g_g1108_p
  (
    .dout(g1108_p),
    .din1(g1085_p_spl_),
    .din2(g1106_n_spl_)
  );


  FA
  g_g1108_n
  (
    .dout(g1108_n),
    .din1(g1085_n_spl_),
    .din2(g1106_p_spl_)
  );


  LA
  g_g1109_p
  (
    .dout(g1109_p),
    .din1(g1107_n_spl_),
    .din2(g1108_n)
  );


  FA
  g_g1109_n
  (
    .dout(g1109_n),
    .din1(g1107_p_spl_),
    .din2(g1108_p)
  );


  LA
  g_g1110_p
  (
    .dout(g1110_p),
    .din1(g1084_n_spl_),
    .din2(g1109_p_spl_)
  );


  FA
  g_g1110_n
  (
    .dout(g1110_n),
    .din1(g1084_p_spl_),
    .din2(g1109_n_spl_)
  );


  LA
  g_g1111_p
  (
    .dout(g1111_p),
    .din1(g1084_p_spl_),
    .din2(g1109_n_spl_)
  );


  FA
  g_g1111_n
  (
    .dout(g1111_n),
    .din1(g1084_n_spl_),
    .din2(g1109_p_spl_)
  );


  LA
  g_g1112_p
  (
    .dout(g1112_p),
    .din1(g1110_n_spl_),
    .din2(g1111_n)
  );


  FA
  g_g1112_n
  (
    .dout(g1112_n),
    .din1(g1110_p_spl_),
    .din2(g1111_p)
  );


  LA
  g_g1113_p
  (
    .dout(g1113_p),
    .din1(g1083_n_spl_),
    .din2(g1112_p_spl_)
  );


  FA
  g_g1113_n
  (
    .dout(g1113_n),
    .din1(g1083_p_spl_),
    .din2(g1112_n_spl_)
  );


  LA
  g_g1114_p
  (
    .dout(g1114_p),
    .din1(g1083_p_spl_),
    .din2(g1112_n_spl_)
  );


  FA
  g_g1114_n
  (
    .dout(g1114_n),
    .din1(g1083_n_spl_),
    .din2(g1112_p_spl_)
  );


  LA
  g_g1115_p
  (
    .dout(g1115_p),
    .din1(g1113_n_spl_),
    .din2(g1114_n)
  );


  FA
  g_g1115_n
  (
    .dout(g1115_n),
    .din1(g1113_p_spl_),
    .din2(g1114_p)
  );


  LA
  g_g1116_p
  (
    .dout(g1116_p),
    .din1(g1082_n_spl_),
    .din2(g1115_p_spl_)
  );


  FA
  g_g1116_n
  (
    .dout(g1116_n),
    .din1(g1082_p_spl_),
    .din2(g1115_n_spl_)
  );


  LA
  g_g1117_p
  (
    .dout(g1117_p),
    .din1(g1082_p_spl_),
    .din2(g1115_n_spl_)
  );


  FA
  g_g1117_n
  (
    .dout(g1117_n),
    .din1(g1082_n_spl_),
    .din2(g1115_p_spl_)
  );


  LA
  g_g1118_p
  (
    .dout(g1118_p),
    .din1(g1116_n_spl_),
    .din2(g1117_n)
  );


  FA
  g_g1118_n
  (
    .dout(g1118_n),
    .din1(g1116_p_spl_),
    .din2(g1117_p)
  );


  LA
  g_g1119_p
  (
    .dout(g1119_p),
    .din1(g1081_n_spl_),
    .din2(g1118_p_spl_)
  );


  FA
  g_g1119_n
  (
    .dout(g1119_n),
    .din1(g1081_p_spl_),
    .din2(g1118_n_spl_)
  );


  LA
  g_g1120_p
  (
    .dout(g1120_p),
    .din1(g1081_p_spl_),
    .din2(g1118_n_spl_)
  );


  FA
  g_g1120_n
  (
    .dout(g1120_n),
    .din1(g1081_n_spl_),
    .din2(g1118_p_spl_)
  );


  LA
  g_g1121_p
  (
    .dout(g1121_p),
    .din1(g1119_n_spl_),
    .din2(g1120_n)
  );


  FA
  g_g1121_n
  (
    .dout(g1121_n),
    .din1(g1119_p_spl_),
    .din2(g1120_p)
  );


  LA
  g_g1122_p
  (
    .dout(g1122_p),
    .din1(g1080_n_spl_),
    .din2(g1121_p_spl_)
  );


  FA
  g_g1122_n
  (
    .dout(g1122_n),
    .din1(g1080_p_spl_),
    .din2(g1121_n_spl_)
  );


  LA
  g_g1123_p
  (
    .dout(g1123_p),
    .din1(g1080_p_spl_),
    .din2(g1121_n_spl_)
  );


  FA
  g_g1123_n
  (
    .dout(g1123_n),
    .din1(g1080_n_spl_),
    .din2(g1121_p_spl_)
  );


  LA
  g_g1124_p
  (
    .dout(g1124_p),
    .din1(g1122_n_spl_),
    .din2(g1123_n)
  );


  FA
  g_g1124_n
  (
    .dout(g1124_n),
    .din1(g1122_p_spl_),
    .din2(g1123_p)
  );


  LA
  g_g1125_p
  (
    .dout(g1125_p),
    .din1(g1079_n_spl_),
    .din2(g1124_p_spl_)
  );


  FA
  g_g1125_n
  (
    .dout(g1125_n),
    .din1(g1079_p_spl_),
    .din2(g1124_n_spl_)
  );


  LA
  g_g1126_p
  (
    .dout(g1126_p),
    .din1(g1079_p_spl_),
    .din2(g1124_n_spl_)
  );


  FA
  g_g1126_n
  (
    .dout(g1126_n),
    .din1(g1079_n_spl_),
    .din2(g1124_p_spl_)
  );


  LA
  g_g1127_p
  (
    .dout(g1127_p),
    .din1(g1125_n_spl_),
    .din2(g1126_n)
  );


  FA
  g_g1127_n
  (
    .dout(g1127_n),
    .din1(g1125_p_spl_),
    .din2(g1126_p)
  );


  LA
  g_g1128_p
  (
    .dout(g1128_p),
    .din1(g1078_n_spl_),
    .din2(g1127_p_spl_)
  );


  FA
  g_g1128_n
  (
    .dout(g1128_n),
    .din1(g1078_p_spl_),
    .din2(g1127_n_spl_)
  );


  LA
  g_g1129_p
  (
    .dout(g1129_p),
    .din1(g1078_p_spl_),
    .din2(g1127_n_spl_)
  );


  FA
  g_g1129_n
  (
    .dout(g1129_n),
    .din1(g1078_n_spl_),
    .din2(g1127_p_spl_)
  );


  LA
  g_g1130_p
  (
    .dout(g1130_p),
    .din1(g1128_n_spl_),
    .din2(g1129_n)
  );


  FA
  g_g1130_n
  (
    .dout(g1130_n),
    .din1(g1128_p_spl_),
    .din2(g1129_p)
  );


  LA
  g_g1131_p
  (
    .dout(g1131_p),
    .din1(g1077_n_spl_),
    .din2(g1130_p_spl_)
  );


  FA
  g_g1131_n
  (
    .dout(g1131_n),
    .din1(g1077_p_spl_),
    .din2(g1130_n_spl_)
  );


  LA
  g_g1132_p
  (
    .dout(g1132_p),
    .din1(g1077_p_spl_),
    .din2(g1130_n_spl_)
  );


  FA
  g_g1132_n
  (
    .dout(g1132_n),
    .din1(g1077_n_spl_),
    .din2(g1130_p_spl_)
  );


  LA
  g_g1133_p
  (
    .dout(g1133_p),
    .din1(g1131_n_spl_),
    .din2(g1132_n)
  );


  FA
  g_g1133_n
  (
    .dout(g1133_n),
    .din1(g1131_p_spl_),
    .din2(g1132_p)
  );


  LA
  g_g1134_p
  (
    .dout(g1134_p),
    .din1(g1076_n_spl_),
    .din2(g1133_p_spl_)
  );


  FA
  g_g1134_n
  (
    .dout(g1134_n),
    .din1(g1076_p_spl_),
    .din2(g1133_n_spl_)
  );


  LA
  g_g1135_p
  (
    .dout(g1135_p),
    .din1(g1076_p_spl_),
    .din2(g1133_n_spl_)
  );


  FA
  g_g1135_n
  (
    .dout(g1135_n),
    .din1(g1076_n_spl_),
    .din2(g1133_p_spl_)
  );


  LA
  g_g1136_p
  (
    .dout(g1136_p),
    .din1(g1134_n_spl_),
    .din2(g1135_n)
  );


  FA
  g_g1136_n
  (
    .dout(g1136_n),
    .din1(g1134_p_spl_),
    .din2(g1135_p)
  );


  LA
  g_g1137_p
  (
    .dout(g1137_p),
    .din1(g1075_n_spl_),
    .din2(g1136_p_spl_)
  );


  FA
  g_g1137_n
  (
    .dout(g1137_n),
    .din1(g1075_p_spl_),
    .din2(g1136_n_spl_)
  );


  LA
  g_g1138_p
  (
    .dout(g1138_p),
    .din1(g1075_p_spl_),
    .din2(g1136_n_spl_)
  );


  FA
  g_g1138_n
  (
    .dout(g1138_n),
    .din1(g1075_n_spl_),
    .din2(g1136_p_spl_)
  );


  LA
  g_g1139_p
  (
    .dout(g1139_p),
    .din1(g1137_n_spl_),
    .din2(g1138_n)
  );


  FA
  g_g1139_n
  (
    .dout(g1139_n),
    .din1(g1137_p_spl_),
    .din2(g1138_p)
  );


  LA
  g_g1140_p
  (
    .dout(g1140_p),
    .din1(g1074_n_spl_),
    .din2(g1139_p_spl_)
  );


  FA
  g_g1140_n
  (
    .dout(g1140_n),
    .din1(g1074_p_spl_),
    .din2(g1139_n_spl_)
  );


  LA
  g_g1141_p
  (
    .dout(g1141_p),
    .din1(g1074_p_spl_),
    .din2(g1139_n_spl_)
  );


  FA
  g_g1141_n
  (
    .dout(g1141_n),
    .din1(g1074_n_spl_),
    .din2(g1139_p_spl_)
  );


  LA
  g_g1142_p
  (
    .dout(g1142_p),
    .din1(g1140_n_spl_),
    .din2(g1141_n)
  );


  FA
  g_g1142_n
  (
    .dout(g1142_n),
    .din1(g1140_p_spl_),
    .din2(g1141_p)
  );


  LA
  g_g1143_p
  (
    .dout(g1143_p),
    .din1(g1073_n_spl_),
    .din2(g1142_p_spl_)
  );


  FA
  g_g1143_n
  (
    .dout(g1143_n),
    .din1(g1073_p_spl_),
    .din2(g1142_n_spl_)
  );


  LA
  g_g1144_p
  (
    .dout(g1144_p),
    .din1(g1073_p_spl_),
    .din2(g1142_n_spl_)
  );


  FA
  g_g1144_n
  (
    .dout(g1144_n),
    .din1(g1073_n_spl_),
    .din2(g1142_p_spl_)
  );


  LA
  g_g1145_p
  (
    .dout(g1145_p),
    .din1(g1143_n_spl_),
    .din2(g1144_n)
  );


  FA
  g_g1145_n
  (
    .dout(g1145_n),
    .din1(g1143_p_spl_),
    .din2(g1144_p)
  );


  LA
  g_g1146_p
  (
    .dout(g1146_p),
    .din1(g1072_n_spl_),
    .din2(g1145_p_spl_)
  );


  FA
  g_g1146_n
  (
    .dout(g1146_n),
    .din1(g1072_p_spl_),
    .din2(g1145_n_spl_)
  );


  LA
  g_g1147_p
  (
    .dout(g1147_p),
    .din1(g1072_p_spl_),
    .din2(g1145_n_spl_)
  );


  FA
  g_g1147_n
  (
    .dout(g1147_n),
    .din1(g1072_n_spl_),
    .din2(g1145_p_spl_)
  );


  LA
  g_g1148_p
  (
    .dout(g1148_p),
    .din1(g1146_n_spl_),
    .din2(g1147_n)
  );


  FA
  g_g1148_n
  (
    .dout(g1148_n),
    .din1(g1146_p_spl_),
    .din2(g1147_p)
  );


  LA
  g_g1149_p
  (
    .dout(g1149_p),
    .din1(g1071_n_spl_),
    .din2(g1148_p_spl_)
  );


  FA
  g_g1149_n
  (
    .dout(g1149_n),
    .din1(g1071_p_spl_),
    .din2(g1148_n_spl_)
  );


  LA
  g_g1150_p
  (
    .dout(g1150_p),
    .din1(g1071_p_spl_),
    .din2(g1148_n_spl_)
  );


  FA
  g_g1150_n
  (
    .dout(g1150_n),
    .din1(g1071_n_spl_),
    .din2(g1148_p_spl_)
  );


  LA
  g_g1151_p
  (
    .dout(g1151_p),
    .din1(g1149_n_spl_),
    .din2(g1150_n)
  );


  FA
  g_g1151_n
  (
    .dout(g1151_n),
    .din1(g1149_p_spl_),
    .din2(g1150_p)
  );


  LA
  g_g1152_p
  (
    .dout(g1152_p),
    .din1(g1070_n_spl_),
    .din2(g1151_p_spl_)
  );


  FA
  g_g1152_n
  (
    .dout(g1152_n),
    .din1(g1070_p_spl_),
    .din2(g1151_n_spl_)
  );


  LA
  g_g1153_p
  (
    .dout(g1153_p),
    .din1(g1070_p_spl_),
    .din2(g1151_n_spl_)
  );


  FA
  g_g1153_n
  (
    .dout(g1153_n),
    .din1(g1070_n_spl_),
    .din2(g1151_p_spl_)
  );


  LA
  g_g1154_p
  (
    .dout(g1154_p),
    .din1(g1152_n_spl_),
    .din2(g1153_n)
  );


  FA
  g_g1154_n
  (
    .dout(g1154_n),
    .din1(g1152_p_spl_),
    .din2(g1153_p)
  );


  LA
  g_g1155_p
  (
    .dout(g1155_p),
    .din1(g1069_n_spl_),
    .din2(g1154_p_spl_)
  );


  FA
  g_g1155_n
  (
    .dout(g1155_n),
    .din1(g1069_p_spl_),
    .din2(g1154_n_spl_)
  );


  LA
  g_g1156_p
  (
    .dout(g1156_p),
    .din1(g1069_p_spl_),
    .din2(g1154_n_spl_)
  );


  FA
  g_g1156_n
  (
    .dout(g1156_n),
    .din1(g1069_n_spl_),
    .din2(g1154_p_spl_)
  );


  LA
  g_g1157_p
  (
    .dout(g1157_p),
    .din1(g1155_n_spl_),
    .din2(g1156_n)
  );


  FA
  g_g1157_n
  (
    .dout(g1157_n),
    .din1(g1155_p_spl_),
    .din2(g1156_p)
  );


  LA
  g_g1158_p
  (
    .dout(g1158_p),
    .din1(g1068_n_spl_),
    .din2(g1157_p_spl_)
  );


  FA
  g_g1158_n
  (
    .dout(g1158_n),
    .din1(g1068_p_spl_),
    .din2(g1157_n_spl_)
  );


  LA
  g_g1159_p
  (
    .dout(g1159_p),
    .din1(g1068_p_spl_),
    .din2(g1157_n_spl_)
  );


  FA
  g_g1159_n
  (
    .dout(g1159_n),
    .din1(g1068_n_spl_),
    .din2(g1157_p_spl_)
  );


  LA
  g_g1160_p
  (
    .dout(g1160_p),
    .din1(g1158_n_spl_),
    .din2(g1159_n)
  );


  FA
  g_g1160_n
  (
    .dout(g1160_n),
    .din1(g1158_p_spl_),
    .din2(g1159_p)
  );


  LA
  g_g1161_p
  (
    .dout(g1161_p),
    .din1(g1067_n_spl_),
    .din2(g1160_p_spl_)
  );


  FA
  g_g1161_n
  (
    .dout(g1161_n),
    .din1(g1067_p_spl_),
    .din2(g1160_n_spl_)
  );


  LA
  g_g1162_p
  (
    .dout(g1162_p),
    .din1(g1067_p_spl_),
    .din2(g1160_n_spl_)
  );


  FA
  g_g1162_n
  (
    .dout(g1162_n),
    .din1(g1067_n_spl_),
    .din2(g1160_p_spl_)
  );


  LA
  g_g1163_p
  (
    .dout(g1163_p),
    .din1(g1161_n_spl_),
    .din2(g1162_n)
  );


  FA
  g_g1163_n
  (
    .dout(g1163_n),
    .din1(g1161_p_spl_),
    .din2(g1162_p)
  );


  LA
  g_g1164_p
  (
    .dout(g1164_p),
    .din1(g1066_n_spl_),
    .din2(g1163_p_spl_)
  );


  FA
  g_g1164_n
  (
    .dout(g1164_n),
    .din1(g1066_p_spl_),
    .din2(g1163_n_spl_)
  );


  LA
  g_g1165_p
  (
    .dout(g1165_p),
    .din1(g1066_p_spl_),
    .din2(g1163_n_spl_)
  );


  FA
  g_g1165_n
  (
    .dout(g1165_n),
    .din1(g1066_n_spl_),
    .din2(g1163_p_spl_)
  );


  LA
  g_g1166_p
  (
    .dout(g1166_p),
    .din1(g1164_n_spl_),
    .din2(g1165_n)
  );


  FA
  g_g1166_n
  (
    .dout(g1166_n),
    .din1(g1164_p_spl_),
    .din2(g1165_p)
  );


  LA
  g_g1167_p
  (
    .dout(g1167_p),
    .din1(g1065_n_spl_),
    .din2(g1166_p_spl_)
  );


  FA
  g_g1167_n
  (
    .dout(g1167_n),
    .din1(g1065_p_spl_),
    .din2(g1166_n_spl_)
  );


  LA
  g_g1168_p
  (
    .dout(g1168_p),
    .din1(g1065_p_spl_),
    .din2(g1166_n_spl_)
  );


  FA
  g_g1168_n
  (
    .dout(g1168_n),
    .din1(g1065_n_spl_),
    .din2(g1166_p_spl_)
  );


  LA
  g_g1169_p
  (
    .dout(g1169_p),
    .din1(g1167_n_spl_),
    .din2(g1168_n)
  );


  FA
  g_g1169_n
  (
    .dout(g1169_n),
    .din1(g1167_p_spl_),
    .din2(g1168_p)
  );


  LA
  g_g1170_p
  (
    .dout(g1170_p),
    .din1(g1064_n_spl_),
    .din2(g1169_p_spl_)
  );


  FA
  g_g1170_n
  (
    .dout(g1170_n),
    .din1(g1064_p_spl_),
    .din2(g1169_n_spl_)
  );


  LA
  g_g1171_p
  (
    .dout(g1171_p),
    .din1(g1064_p_spl_),
    .din2(g1169_n_spl_)
  );


  FA
  g_g1171_n
  (
    .dout(g1171_n),
    .din1(g1064_n_spl_),
    .din2(g1169_p_spl_)
  );


  LA
  g_g1172_p
  (
    .dout(g1172_p),
    .din1(g1170_n_spl_),
    .din2(g1171_n)
  );


  FA
  g_g1172_n
  (
    .dout(g1172_n),
    .din1(g1170_p_spl_),
    .din2(g1171_p)
  );


  LA
  g_g1173_p
  (
    .dout(g1173_p),
    .din1(g1062_n_spl_),
    .din2(g1172_p)
  );


  FA
  g_g1173_n
  (
    .dout(g1173_n),
    .din1(g1062_p_spl_),
    .din2(g1172_n_spl_)
  );


  LA
  g_g1174_p
  (
    .dout(g1174_p),
    .din1(g1062_p_spl_),
    .din2(g1172_n_spl_)
  );


  FA
  g_g1175_n
  (
    .dout(g1175_n),
    .din1(g1173_p_spl_),
    .din2(g1174_p)
  );


  LA
  g_g1176_p
  (
    .dout(g1176_p),
    .din1(g1170_n_spl_),
    .din2(g1173_n)
  );


  FA
  g_g1176_n
  (
    .dout(g1176_n),
    .din1(g1170_p_spl_),
    .din2(g1173_p_spl_)
  );


  LA
  g_g1177_p
  (
    .dout(g1177_p),
    .din1(g1164_n_spl_),
    .din2(g1167_n_spl_)
  );


  FA
  g_g1177_n
  (
    .dout(g1177_n),
    .din1(g1164_p_spl_),
    .din2(g1167_p_spl_)
  );


  LA
  g_g1178_p
  (
    .dout(g1178_p),
    .din1(G4_p_spl_111),
    .din2(G32_p_spl_001)
  );


  FA
  g_g1178_n
  (
    .dout(g1178_n),
    .din1(G4_n_spl_111),
    .din2(G32_n_spl_001)
  );


  LA
  g_g1179_p
  (
    .dout(g1179_p),
    .din1(g1158_n_spl_),
    .din2(g1161_n_spl_)
  );


  FA
  g_g1179_n
  (
    .dout(g1179_n),
    .din1(g1158_p_spl_),
    .din2(g1161_p_spl_)
  );


  LA
  g_g1180_p
  (
    .dout(g1180_p),
    .din1(G5_p_spl_111),
    .din2(G31_p_spl_010)
  );


  FA
  g_g1180_n
  (
    .dout(g1180_n),
    .din1(G5_n_spl_111),
    .din2(G31_n_spl_010)
  );


  LA
  g_g1181_p
  (
    .dout(g1181_p),
    .din1(g1152_n_spl_),
    .din2(g1155_n_spl_)
  );


  FA
  g_g1181_n
  (
    .dout(g1181_n),
    .din1(g1152_p_spl_),
    .din2(g1155_p_spl_)
  );


  LA
  g_g1182_p
  (
    .dout(g1182_p),
    .din1(G6_p_spl_110),
    .din2(G30_p_spl_010)
  );


  FA
  g_g1182_n
  (
    .dout(g1182_n),
    .din1(G6_n_spl_110),
    .din2(G30_n_spl_010)
  );


  LA
  g_g1183_p
  (
    .dout(g1183_p),
    .din1(g1146_n_spl_),
    .din2(g1149_n_spl_)
  );


  FA
  g_g1183_n
  (
    .dout(g1183_n),
    .din1(g1146_p_spl_),
    .din2(g1149_p_spl_)
  );


  LA
  g_g1184_p
  (
    .dout(g1184_p),
    .din1(G7_p_spl_110),
    .din2(G29_p_spl_011)
  );


  FA
  g_g1184_n
  (
    .dout(g1184_n),
    .din1(G7_n_spl_110),
    .din2(G29_n_spl_011)
  );


  LA
  g_g1185_p
  (
    .dout(g1185_p),
    .din1(g1140_n_spl_),
    .din2(g1143_n_spl_)
  );


  FA
  g_g1185_n
  (
    .dout(g1185_n),
    .din1(g1140_p_spl_),
    .din2(g1143_p_spl_)
  );


  LA
  g_g1186_p
  (
    .dout(g1186_p),
    .din1(G8_p_spl_101),
    .din2(G28_p_spl_011)
  );


  FA
  g_g1186_n
  (
    .dout(g1186_n),
    .din1(G8_n_spl_101),
    .din2(G28_n_spl_011)
  );


  LA
  g_g1187_p
  (
    .dout(g1187_p),
    .din1(g1134_n_spl_),
    .din2(g1137_n_spl_)
  );


  FA
  g_g1187_n
  (
    .dout(g1187_n),
    .din1(g1134_p_spl_),
    .din2(g1137_p_spl_)
  );


  LA
  g_g1188_p
  (
    .dout(g1188_p),
    .din1(G9_p_spl_101),
    .din2(G27_p_spl_100)
  );


  FA
  g_g1188_n
  (
    .dout(g1188_n),
    .din1(G9_n_spl_101),
    .din2(G27_n_spl_100)
  );


  LA
  g_g1189_p
  (
    .dout(g1189_p),
    .din1(g1128_n_spl_),
    .din2(g1131_n_spl_)
  );


  FA
  g_g1189_n
  (
    .dout(g1189_n),
    .din1(g1128_p_spl_),
    .din2(g1131_p_spl_)
  );


  LA
  g_g1190_p
  (
    .dout(g1190_p),
    .din1(G10_p_spl_100),
    .din2(G26_p_spl_100)
  );


  FA
  g_g1190_n
  (
    .dout(g1190_n),
    .din1(G10_n_spl_100),
    .din2(G26_n_spl_100)
  );


  LA
  g_g1191_p
  (
    .dout(g1191_p),
    .din1(g1122_n_spl_),
    .din2(g1125_n_spl_)
  );


  FA
  g_g1191_n
  (
    .dout(g1191_n),
    .din1(g1122_p_spl_),
    .din2(g1125_p_spl_)
  );


  LA
  g_g1192_p
  (
    .dout(g1192_p),
    .din1(G11_p_spl_100),
    .din2(G25_p_spl_101)
  );


  FA
  g_g1192_n
  (
    .dout(g1192_n),
    .din1(G11_n_spl_100),
    .din2(G25_n_spl_101)
  );


  LA
  g_g1193_p
  (
    .dout(g1193_p),
    .din1(g1116_n_spl_),
    .din2(g1119_n_spl_)
  );


  FA
  g_g1193_n
  (
    .dout(g1193_n),
    .din1(g1116_p_spl_),
    .din2(g1119_p_spl_)
  );


  LA
  g_g1194_p
  (
    .dout(g1194_p),
    .din1(G12_p_spl_011),
    .din2(G24_p_spl_101)
  );


  FA
  g_g1194_n
  (
    .dout(g1194_n),
    .din1(G12_n_spl_011),
    .din2(G24_n_spl_101)
  );


  LA
  g_g1195_p
  (
    .dout(g1195_p),
    .din1(g1110_n_spl_),
    .din2(g1113_n_spl_)
  );


  FA
  g_g1195_n
  (
    .dout(g1195_n),
    .din1(g1110_p_spl_),
    .din2(g1113_p_spl_)
  );


  LA
  g_g1196_p
  (
    .dout(g1196_p),
    .din1(G13_p_spl_011),
    .din2(G23_p_spl_110)
  );


  FA
  g_g1196_n
  (
    .dout(g1196_n),
    .din1(G13_n_spl_011),
    .din2(G23_n_spl_110)
  );


  LA
  g_g1197_p
  (
    .dout(g1197_p),
    .din1(g1104_n_spl_),
    .din2(g1107_n_spl_)
  );


  FA
  g_g1197_n
  (
    .dout(g1197_n),
    .din1(g1104_p_spl_),
    .din2(g1107_p_spl_)
  );


  LA
  g_g1198_p
  (
    .dout(g1198_p),
    .din1(G14_p_spl_010),
    .din2(G22_p_spl_110)
  );


  FA
  g_g1198_n
  (
    .dout(g1198_n),
    .din1(G14_n_spl_010),
    .din2(G22_n_spl_110)
  );


  LA
  g_g1199_p
  (
    .dout(g1199_p),
    .din1(g1098_n_spl_),
    .din2(g1101_n_spl_)
  );


  FA
  g_g1199_n
  (
    .dout(g1199_n),
    .din1(g1098_p_spl_),
    .din2(g1101_p_spl_)
  );


  LA
  g_g1200_p
  (
    .dout(g1200_p),
    .din1(G15_p_spl_010),
    .din2(G21_p_spl_111)
  );


  FA
  g_g1200_n
  (
    .dout(g1200_n),
    .din1(G15_n_spl_010),
    .din2(G21_n_spl_111)
  );


  LA
  g_g1201_p
  (
    .dout(g1201_p),
    .din1(G16_p_spl_001),
    .din2(G20_p_spl_111)
  );


  FA
  g_g1201_n
  (
    .dout(g1201_n),
    .din1(G16_n_spl_001),
    .din2(G20_n_spl_111)
  );


  LA
  g_g1202_p
  (
    .dout(g1202_p),
    .din1(g1092_n_spl_),
    .din2(g1095_n_spl_)
  );


  FA
  g_g1202_n
  (
    .dout(g1202_n),
    .din1(g1092_p_spl_),
    .din2(g1095_p_spl_)
  );


  LA
  g_g1203_p
  (
    .dout(g1203_p),
    .din1(g1201_n_spl_),
    .din2(g1202_n_spl_)
  );


  FA
  g_g1203_n
  (
    .dout(g1203_n),
    .din1(g1201_p_spl_),
    .din2(g1202_p_spl_)
  );


  LA
  g_g1204_p
  (
    .dout(g1204_p),
    .din1(g1201_p_spl_),
    .din2(g1202_p_spl_)
  );


  FA
  g_g1204_n
  (
    .dout(g1204_n),
    .din1(g1201_n_spl_),
    .din2(g1202_n_spl_)
  );


  LA
  g_g1205_p
  (
    .dout(g1205_p),
    .din1(g1203_n_spl_),
    .din2(g1204_n)
  );


  FA
  g_g1205_n
  (
    .dout(g1205_n),
    .din1(g1203_p_spl_),
    .din2(g1204_p)
  );


  LA
  g_g1206_p
  (
    .dout(g1206_p),
    .din1(g1200_n_spl_),
    .din2(g1205_p_spl_)
  );


  FA
  g_g1206_n
  (
    .dout(g1206_n),
    .din1(g1200_p_spl_),
    .din2(g1205_n_spl_)
  );


  LA
  g_g1207_p
  (
    .dout(g1207_p),
    .din1(g1200_p_spl_),
    .din2(g1205_n_spl_)
  );


  FA
  g_g1207_n
  (
    .dout(g1207_n),
    .din1(g1200_n_spl_),
    .din2(g1205_p_spl_)
  );


  LA
  g_g1208_p
  (
    .dout(g1208_p),
    .din1(g1206_n_spl_),
    .din2(g1207_n)
  );


  FA
  g_g1208_n
  (
    .dout(g1208_n),
    .din1(g1206_p_spl_),
    .din2(g1207_p)
  );


  LA
  g_g1209_p
  (
    .dout(g1209_p),
    .din1(g1199_n_spl_),
    .din2(g1208_p_spl_)
  );


  FA
  g_g1209_n
  (
    .dout(g1209_n),
    .din1(g1199_p_spl_),
    .din2(g1208_n_spl_)
  );


  LA
  g_g1210_p
  (
    .dout(g1210_p),
    .din1(g1199_p_spl_),
    .din2(g1208_n_spl_)
  );


  FA
  g_g1210_n
  (
    .dout(g1210_n),
    .din1(g1199_n_spl_),
    .din2(g1208_p_spl_)
  );


  LA
  g_g1211_p
  (
    .dout(g1211_p),
    .din1(g1209_n_spl_),
    .din2(g1210_n)
  );


  FA
  g_g1211_n
  (
    .dout(g1211_n),
    .din1(g1209_p_spl_),
    .din2(g1210_p)
  );


  LA
  g_g1212_p
  (
    .dout(g1212_p),
    .din1(g1198_n_spl_),
    .din2(g1211_p_spl_)
  );


  FA
  g_g1212_n
  (
    .dout(g1212_n),
    .din1(g1198_p_spl_),
    .din2(g1211_n_spl_)
  );


  LA
  g_g1213_p
  (
    .dout(g1213_p),
    .din1(g1198_p_spl_),
    .din2(g1211_n_spl_)
  );


  FA
  g_g1213_n
  (
    .dout(g1213_n),
    .din1(g1198_n_spl_),
    .din2(g1211_p_spl_)
  );


  LA
  g_g1214_p
  (
    .dout(g1214_p),
    .din1(g1212_n_spl_),
    .din2(g1213_n)
  );


  FA
  g_g1214_n
  (
    .dout(g1214_n),
    .din1(g1212_p_spl_),
    .din2(g1213_p)
  );


  LA
  g_g1215_p
  (
    .dout(g1215_p),
    .din1(g1197_n_spl_),
    .din2(g1214_p_spl_)
  );


  FA
  g_g1215_n
  (
    .dout(g1215_n),
    .din1(g1197_p_spl_),
    .din2(g1214_n_spl_)
  );


  LA
  g_g1216_p
  (
    .dout(g1216_p),
    .din1(g1197_p_spl_),
    .din2(g1214_n_spl_)
  );


  FA
  g_g1216_n
  (
    .dout(g1216_n),
    .din1(g1197_n_spl_),
    .din2(g1214_p_spl_)
  );


  LA
  g_g1217_p
  (
    .dout(g1217_p),
    .din1(g1215_n_spl_),
    .din2(g1216_n)
  );


  FA
  g_g1217_n
  (
    .dout(g1217_n),
    .din1(g1215_p_spl_),
    .din2(g1216_p)
  );


  LA
  g_g1218_p
  (
    .dout(g1218_p),
    .din1(g1196_n_spl_),
    .din2(g1217_p_spl_)
  );


  FA
  g_g1218_n
  (
    .dout(g1218_n),
    .din1(g1196_p_spl_),
    .din2(g1217_n_spl_)
  );


  LA
  g_g1219_p
  (
    .dout(g1219_p),
    .din1(g1196_p_spl_),
    .din2(g1217_n_spl_)
  );


  FA
  g_g1219_n
  (
    .dout(g1219_n),
    .din1(g1196_n_spl_),
    .din2(g1217_p_spl_)
  );


  LA
  g_g1220_p
  (
    .dout(g1220_p),
    .din1(g1218_n_spl_),
    .din2(g1219_n)
  );


  FA
  g_g1220_n
  (
    .dout(g1220_n),
    .din1(g1218_p_spl_),
    .din2(g1219_p)
  );


  LA
  g_g1221_p
  (
    .dout(g1221_p),
    .din1(g1195_n_spl_),
    .din2(g1220_p_spl_)
  );


  FA
  g_g1221_n
  (
    .dout(g1221_n),
    .din1(g1195_p_spl_),
    .din2(g1220_n_spl_)
  );


  LA
  g_g1222_p
  (
    .dout(g1222_p),
    .din1(g1195_p_spl_),
    .din2(g1220_n_spl_)
  );


  FA
  g_g1222_n
  (
    .dout(g1222_n),
    .din1(g1195_n_spl_),
    .din2(g1220_p_spl_)
  );


  LA
  g_g1223_p
  (
    .dout(g1223_p),
    .din1(g1221_n_spl_),
    .din2(g1222_n)
  );


  FA
  g_g1223_n
  (
    .dout(g1223_n),
    .din1(g1221_p_spl_),
    .din2(g1222_p)
  );


  LA
  g_g1224_p
  (
    .dout(g1224_p),
    .din1(g1194_n_spl_),
    .din2(g1223_p_spl_)
  );


  FA
  g_g1224_n
  (
    .dout(g1224_n),
    .din1(g1194_p_spl_),
    .din2(g1223_n_spl_)
  );


  LA
  g_g1225_p
  (
    .dout(g1225_p),
    .din1(g1194_p_spl_),
    .din2(g1223_n_spl_)
  );


  FA
  g_g1225_n
  (
    .dout(g1225_n),
    .din1(g1194_n_spl_),
    .din2(g1223_p_spl_)
  );


  LA
  g_g1226_p
  (
    .dout(g1226_p),
    .din1(g1224_n_spl_),
    .din2(g1225_n)
  );


  FA
  g_g1226_n
  (
    .dout(g1226_n),
    .din1(g1224_p_spl_),
    .din2(g1225_p)
  );


  LA
  g_g1227_p
  (
    .dout(g1227_p),
    .din1(g1193_n_spl_),
    .din2(g1226_p_spl_)
  );


  FA
  g_g1227_n
  (
    .dout(g1227_n),
    .din1(g1193_p_spl_),
    .din2(g1226_n_spl_)
  );


  LA
  g_g1228_p
  (
    .dout(g1228_p),
    .din1(g1193_p_spl_),
    .din2(g1226_n_spl_)
  );


  FA
  g_g1228_n
  (
    .dout(g1228_n),
    .din1(g1193_n_spl_),
    .din2(g1226_p_spl_)
  );


  LA
  g_g1229_p
  (
    .dout(g1229_p),
    .din1(g1227_n_spl_),
    .din2(g1228_n)
  );


  FA
  g_g1229_n
  (
    .dout(g1229_n),
    .din1(g1227_p_spl_),
    .din2(g1228_p)
  );


  LA
  g_g1230_p
  (
    .dout(g1230_p),
    .din1(g1192_n_spl_),
    .din2(g1229_p_spl_)
  );


  FA
  g_g1230_n
  (
    .dout(g1230_n),
    .din1(g1192_p_spl_),
    .din2(g1229_n_spl_)
  );


  LA
  g_g1231_p
  (
    .dout(g1231_p),
    .din1(g1192_p_spl_),
    .din2(g1229_n_spl_)
  );


  FA
  g_g1231_n
  (
    .dout(g1231_n),
    .din1(g1192_n_spl_),
    .din2(g1229_p_spl_)
  );


  LA
  g_g1232_p
  (
    .dout(g1232_p),
    .din1(g1230_n_spl_),
    .din2(g1231_n)
  );


  FA
  g_g1232_n
  (
    .dout(g1232_n),
    .din1(g1230_p_spl_),
    .din2(g1231_p)
  );


  LA
  g_g1233_p
  (
    .dout(g1233_p),
    .din1(g1191_n_spl_),
    .din2(g1232_p_spl_)
  );


  FA
  g_g1233_n
  (
    .dout(g1233_n),
    .din1(g1191_p_spl_),
    .din2(g1232_n_spl_)
  );


  LA
  g_g1234_p
  (
    .dout(g1234_p),
    .din1(g1191_p_spl_),
    .din2(g1232_n_spl_)
  );


  FA
  g_g1234_n
  (
    .dout(g1234_n),
    .din1(g1191_n_spl_),
    .din2(g1232_p_spl_)
  );


  LA
  g_g1235_p
  (
    .dout(g1235_p),
    .din1(g1233_n_spl_),
    .din2(g1234_n)
  );


  FA
  g_g1235_n
  (
    .dout(g1235_n),
    .din1(g1233_p_spl_),
    .din2(g1234_p)
  );


  LA
  g_g1236_p
  (
    .dout(g1236_p),
    .din1(g1190_n_spl_),
    .din2(g1235_p_spl_)
  );


  FA
  g_g1236_n
  (
    .dout(g1236_n),
    .din1(g1190_p_spl_),
    .din2(g1235_n_spl_)
  );


  LA
  g_g1237_p
  (
    .dout(g1237_p),
    .din1(g1190_p_spl_),
    .din2(g1235_n_spl_)
  );


  FA
  g_g1237_n
  (
    .dout(g1237_n),
    .din1(g1190_n_spl_),
    .din2(g1235_p_spl_)
  );


  LA
  g_g1238_p
  (
    .dout(g1238_p),
    .din1(g1236_n_spl_),
    .din2(g1237_n)
  );


  FA
  g_g1238_n
  (
    .dout(g1238_n),
    .din1(g1236_p_spl_),
    .din2(g1237_p)
  );


  LA
  g_g1239_p
  (
    .dout(g1239_p),
    .din1(g1189_n_spl_),
    .din2(g1238_p_spl_)
  );


  FA
  g_g1239_n
  (
    .dout(g1239_n),
    .din1(g1189_p_spl_),
    .din2(g1238_n_spl_)
  );


  LA
  g_g1240_p
  (
    .dout(g1240_p),
    .din1(g1189_p_spl_),
    .din2(g1238_n_spl_)
  );


  FA
  g_g1240_n
  (
    .dout(g1240_n),
    .din1(g1189_n_spl_),
    .din2(g1238_p_spl_)
  );


  LA
  g_g1241_p
  (
    .dout(g1241_p),
    .din1(g1239_n_spl_),
    .din2(g1240_n)
  );


  FA
  g_g1241_n
  (
    .dout(g1241_n),
    .din1(g1239_p_spl_),
    .din2(g1240_p)
  );


  LA
  g_g1242_p
  (
    .dout(g1242_p),
    .din1(g1188_n_spl_),
    .din2(g1241_p_spl_)
  );


  FA
  g_g1242_n
  (
    .dout(g1242_n),
    .din1(g1188_p_spl_),
    .din2(g1241_n_spl_)
  );


  LA
  g_g1243_p
  (
    .dout(g1243_p),
    .din1(g1188_p_spl_),
    .din2(g1241_n_spl_)
  );


  FA
  g_g1243_n
  (
    .dout(g1243_n),
    .din1(g1188_n_spl_),
    .din2(g1241_p_spl_)
  );


  LA
  g_g1244_p
  (
    .dout(g1244_p),
    .din1(g1242_n_spl_),
    .din2(g1243_n)
  );


  FA
  g_g1244_n
  (
    .dout(g1244_n),
    .din1(g1242_p_spl_),
    .din2(g1243_p)
  );


  LA
  g_g1245_p
  (
    .dout(g1245_p),
    .din1(g1187_n_spl_),
    .din2(g1244_p_spl_)
  );


  FA
  g_g1245_n
  (
    .dout(g1245_n),
    .din1(g1187_p_spl_),
    .din2(g1244_n_spl_)
  );


  LA
  g_g1246_p
  (
    .dout(g1246_p),
    .din1(g1187_p_spl_),
    .din2(g1244_n_spl_)
  );


  FA
  g_g1246_n
  (
    .dout(g1246_n),
    .din1(g1187_n_spl_),
    .din2(g1244_p_spl_)
  );


  LA
  g_g1247_p
  (
    .dout(g1247_p),
    .din1(g1245_n_spl_),
    .din2(g1246_n)
  );


  FA
  g_g1247_n
  (
    .dout(g1247_n),
    .din1(g1245_p_spl_),
    .din2(g1246_p)
  );


  LA
  g_g1248_p
  (
    .dout(g1248_p),
    .din1(g1186_n_spl_),
    .din2(g1247_p_spl_)
  );


  FA
  g_g1248_n
  (
    .dout(g1248_n),
    .din1(g1186_p_spl_),
    .din2(g1247_n_spl_)
  );


  LA
  g_g1249_p
  (
    .dout(g1249_p),
    .din1(g1186_p_spl_),
    .din2(g1247_n_spl_)
  );


  FA
  g_g1249_n
  (
    .dout(g1249_n),
    .din1(g1186_n_spl_),
    .din2(g1247_p_spl_)
  );


  LA
  g_g1250_p
  (
    .dout(g1250_p),
    .din1(g1248_n_spl_),
    .din2(g1249_n)
  );


  FA
  g_g1250_n
  (
    .dout(g1250_n),
    .din1(g1248_p_spl_),
    .din2(g1249_p)
  );


  LA
  g_g1251_p
  (
    .dout(g1251_p),
    .din1(g1185_n_spl_),
    .din2(g1250_p_spl_)
  );


  FA
  g_g1251_n
  (
    .dout(g1251_n),
    .din1(g1185_p_spl_),
    .din2(g1250_n_spl_)
  );


  LA
  g_g1252_p
  (
    .dout(g1252_p),
    .din1(g1185_p_spl_),
    .din2(g1250_n_spl_)
  );


  FA
  g_g1252_n
  (
    .dout(g1252_n),
    .din1(g1185_n_spl_),
    .din2(g1250_p_spl_)
  );


  LA
  g_g1253_p
  (
    .dout(g1253_p),
    .din1(g1251_n_spl_),
    .din2(g1252_n)
  );


  FA
  g_g1253_n
  (
    .dout(g1253_n),
    .din1(g1251_p_spl_),
    .din2(g1252_p)
  );


  LA
  g_g1254_p
  (
    .dout(g1254_p),
    .din1(g1184_n_spl_),
    .din2(g1253_p_spl_)
  );


  FA
  g_g1254_n
  (
    .dout(g1254_n),
    .din1(g1184_p_spl_),
    .din2(g1253_n_spl_)
  );


  LA
  g_g1255_p
  (
    .dout(g1255_p),
    .din1(g1184_p_spl_),
    .din2(g1253_n_spl_)
  );


  FA
  g_g1255_n
  (
    .dout(g1255_n),
    .din1(g1184_n_spl_),
    .din2(g1253_p_spl_)
  );


  LA
  g_g1256_p
  (
    .dout(g1256_p),
    .din1(g1254_n_spl_),
    .din2(g1255_n)
  );


  FA
  g_g1256_n
  (
    .dout(g1256_n),
    .din1(g1254_p_spl_),
    .din2(g1255_p)
  );


  LA
  g_g1257_p
  (
    .dout(g1257_p),
    .din1(g1183_n_spl_),
    .din2(g1256_p_spl_)
  );


  FA
  g_g1257_n
  (
    .dout(g1257_n),
    .din1(g1183_p_spl_),
    .din2(g1256_n_spl_)
  );


  LA
  g_g1258_p
  (
    .dout(g1258_p),
    .din1(g1183_p_spl_),
    .din2(g1256_n_spl_)
  );


  FA
  g_g1258_n
  (
    .dout(g1258_n),
    .din1(g1183_n_spl_),
    .din2(g1256_p_spl_)
  );


  LA
  g_g1259_p
  (
    .dout(g1259_p),
    .din1(g1257_n_spl_),
    .din2(g1258_n)
  );


  FA
  g_g1259_n
  (
    .dout(g1259_n),
    .din1(g1257_p_spl_),
    .din2(g1258_p)
  );


  LA
  g_g1260_p
  (
    .dout(g1260_p),
    .din1(g1182_n_spl_),
    .din2(g1259_p_spl_)
  );


  FA
  g_g1260_n
  (
    .dout(g1260_n),
    .din1(g1182_p_spl_),
    .din2(g1259_n_spl_)
  );


  LA
  g_g1261_p
  (
    .dout(g1261_p),
    .din1(g1182_p_spl_),
    .din2(g1259_n_spl_)
  );


  FA
  g_g1261_n
  (
    .dout(g1261_n),
    .din1(g1182_n_spl_),
    .din2(g1259_p_spl_)
  );


  LA
  g_g1262_p
  (
    .dout(g1262_p),
    .din1(g1260_n_spl_),
    .din2(g1261_n)
  );


  FA
  g_g1262_n
  (
    .dout(g1262_n),
    .din1(g1260_p_spl_),
    .din2(g1261_p)
  );


  LA
  g_g1263_p
  (
    .dout(g1263_p),
    .din1(g1181_n_spl_),
    .din2(g1262_p_spl_)
  );


  FA
  g_g1263_n
  (
    .dout(g1263_n),
    .din1(g1181_p_spl_),
    .din2(g1262_n_spl_)
  );


  LA
  g_g1264_p
  (
    .dout(g1264_p),
    .din1(g1181_p_spl_),
    .din2(g1262_n_spl_)
  );


  FA
  g_g1264_n
  (
    .dout(g1264_n),
    .din1(g1181_n_spl_),
    .din2(g1262_p_spl_)
  );


  LA
  g_g1265_p
  (
    .dout(g1265_p),
    .din1(g1263_n_spl_),
    .din2(g1264_n)
  );


  FA
  g_g1265_n
  (
    .dout(g1265_n),
    .din1(g1263_p_spl_),
    .din2(g1264_p)
  );


  LA
  g_g1266_p
  (
    .dout(g1266_p),
    .din1(g1180_n_spl_),
    .din2(g1265_p_spl_)
  );


  FA
  g_g1266_n
  (
    .dout(g1266_n),
    .din1(g1180_p_spl_),
    .din2(g1265_n_spl_)
  );


  LA
  g_g1267_p
  (
    .dout(g1267_p),
    .din1(g1180_p_spl_),
    .din2(g1265_n_spl_)
  );


  FA
  g_g1267_n
  (
    .dout(g1267_n),
    .din1(g1180_n_spl_),
    .din2(g1265_p_spl_)
  );


  LA
  g_g1268_p
  (
    .dout(g1268_p),
    .din1(g1266_n_spl_),
    .din2(g1267_n)
  );


  FA
  g_g1268_n
  (
    .dout(g1268_n),
    .din1(g1266_p_spl_),
    .din2(g1267_p)
  );


  LA
  g_g1269_p
  (
    .dout(g1269_p),
    .din1(g1179_n_spl_),
    .din2(g1268_p_spl_)
  );


  FA
  g_g1269_n
  (
    .dout(g1269_n),
    .din1(g1179_p_spl_),
    .din2(g1268_n_spl_)
  );


  LA
  g_g1270_p
  (
    .dout(g1270_p),
    .din1(g1179_p_spl_),
    .din2(g1268_n_spl_)
  );


  FA
  g_g1270_n
  (
    .dout(g1270_n),
    .din1(g1179_n_spl_),
    .din2(g1268_p_spl_)
  );


  LA
  g_g1271_p
  (
    .dout(g1271_p),
    .din1(g1269_n_spl_),
    .din2(g1270_n)
  );


  FA
  g_g1271_n
  (
    .dout(g1271_n),
    .din1(g1269_p_spl_),
    .din2(g1270_p)
  );


  LA
  g_g1272_p
  (
    .dout(g1272_p),
    .din1(g1178_n_spl_),
    .din2(g1271_p_spl_)
  );


  FA
  g_g1272_n
  (
    .dout(g1272_n),
    .din1(g1178_p_spl_),
    .din2(g1271_n_spl_)
  );


  LA
  g_g1273_p
  (
    .dout(g1273_p),
    .din1(g1178_p_spl_),
    .din2(g1271_n_spl_)
  );


  FA
  g_g1273_n
  (
    .dout(g1273_n),
    .din1(g1178_n_spl_),
    .din2(g1271_p_spl_)
  );


  LA
  g_g1274_p
  (
    .dout(g1274_p),
    .din1(g1272_n_spl_),
    .din2(g1273_n)
  );


  FA
  g_g1274_n
  (
    .dout(g1274_n),
    .din1(g1272_p_spl_),
    .din2(g1273_p)
  );


  LA
  g_g1275_p
  (
    .dout(g1275_p),
    .din1(g1177_n_spl_),
    .din2(g1274_p_spl_)
  );


  FA
  g_g1275_n
  (
    .dout(g1275_n),
    .din1(g1177_p_spl_),
    .din2(g1274_n_spl_)
  );


  LA
  g_g1276_p
  (
    .dout(g1276_p),
    .din1(g1177_p_spl_),
    .din2(g1274_n_spl_)
  );


  FA
  g_g1276_n
  (
    .dout(g1276_n),
    .din1(g1177_n_spl_),
    .din2(g1274_p_spl_)
  );


  LA
  g_g1277_p
  (
    .dout(g1277_p),
    .din1(g1275_n_spl_),
    .din2(g1276_n)
  );


  FA
  g_g1277_n
  (
    .dout(g1277_n),
    .din1(g1275_p_spl_),
    .din2(g1276_p)
  );


  LA
  g_g1278_p
  (
    .dout(g1278_p),
    .din1(g1176_n),
    .din2(g1277_p)
  );


  FA
  g_g1278_n
  (
    .dout(g1278_n),
    .din1(g1176_p_spl_),
    .din2(g1277_n_spl_)
  );


  LA
  g_g1279_p
  (
    .dout(g1279_p),
    .din1(g1176_p_spl_),
    .din2(g1277_n_spl_)
  );


  FA
  g_g1280_n
  (
    .dout(g1280_n),
    .din1(g1278_p_spl_),
    .din2(g1279_p)
  );


  LA
  g_g1281_p
  (
    .dout(g1281_p),
    .din1(g1275_n_spl_),
    .din2(g1278_n)
  );


  FA
  g_g1281_n
  (
    .dout(g1281_n),
    .din1(g1275_p_spl_),
    .din2(g1278_p_spl_)
  );


  LA
  g_g1282_p
  (
    .dout(g1282_p),
    .din1(g1269_n_spl_),
    .din2(g1272_n_spl_)
  );


  FA
  g_g1282_n
  (
    .dout(g1282_n),
    .din1(g1269_p_spl_),
    .din2(g1272_p_spl_)
  );


  LA
  g_g1283_p
  (
    .dout(g1283_p),
    .din1(G5_p_spl_111),
    .din2(G32_p_spl_010)
  );


  FA
  g_g1283_n
  (
    .dout(g1283_n),
    .din1(G5_n_spl_111),
    .din2(G32_n_spl_010)
  );


  LA
  g_g1284_p
  (
    .dout(g1284_p),
    .din1(g1263_n_spl_),
    .din2(g1266_n_spl_)
  );


  FA
  g_g1284_n
  (
    .dout(g1284_n),
    .din1(g1263_p_spl_),
    .din2(g1266_p_spl_)
  );


  LA
  g_g1285_p
  (
    .dout(g1285_p),
    .din1(G6_p_spl_111),
    .din2(G31_p_spl_010)
  );


  FA
  g_g1285_n
  (
    .dout(g1285_n),
    .din1(G6_n_spl_111),
    .din2(G31_n_spl_010)
  );


  LA
  g_g1286_p
  (
    .dout(g1286_p),
    .din1(g1257_n_spl_),
    .din2(g1260_n_spl_)
  );


  FA
  g_g1286_n
  (
    .dout(g1286_n),
    .din1(g1257_p_spl_),
    .din2(g1260_p_spl_)
  );


  LA
  g_g1287_p
  (
    .dout(g1287_p),
    .din1(G7_p_spl_110),
    .din2(G30_p_spl_011)
  );


  FA
  g_g1287_n
  (
    .dout(g1287_n),
    .din1(G7_n_spl_110),
    .din2(G30_n_spl_011)
  );


  LA
  g_g1288_p
  (
    .dout(g1288_p),
    .din1(g1251_n_spl_),
    .din2(g1254_n_spl_)
  );


  FA
  g_g1288_n
  (
    .dout(g1288_n),
    .din1(g1251_p_spl_),
    .din2(g1254_p_spl_)
  );


  LA
  g_g1289_p
  (
    .dout(g1289_p),
    .din1(G8_p_spl_110),
    .din2(G29_p_spl_011)
  );


  FA
  g_g1289_n
  (
    .dout(g1289_n),
    .din1(G8_n_spl_110),
    .din2(G29_n_spl_011)
  );


  LA
  g_g1290_p
  (
    .dout(g1290_p),
    .din1(g1245_n_spl_),
    .din2(g1248_n_spl_)
  );


  FA
  g_g1290_n
  (
    .dout(g1290_n),
    .din1(g1245_p_spl_),
    .din2(g1248_p_spl_)
  );


  LA
  g_g1291_p
  (
    .dout(g1291_p),
    .din1(G9_p_spl_101),
    .din2(G28_p_spl_100)
  );


  FA
  g_g1291_n
  (
    .dout(g1291_n),
    .din1(G9_n_spl_101),
    .din2(G28_n_spl_100)
  );


  LA
  g_g1292_p
  (
    .dout(g1292_p),
    .din1(g1239_n_spl_),
    .din2(g1242_n_spl_)
  );


  FA
  g_g1292_n
  (
    .dout(g1292_n),
    .din1(g1239_p_spl_),
    .din2(g1242_p_spl_)
  );


  LA
  g_g1293_p
  (
    .dout(g1293_p),
    .din1(G10_p_spl_101),
    .din2(G27_p_spl_100)
  );


  FA
  g_g1293_n
  (
    .dout(g1293_n),
    .din1(G10_n_spl_101),
    .din2(G27_n_spl_100)
  );


  LA
  g_g1294_p
  (
    .dout(g1294_p),
    .din1(g1233_n_spl_),
    .din2(g1236_n_spl_)
  );


  FA
  g_g1294_n
  (
    .dout(g1294_n),
    .din1(g1233_p_spl_),
    .din2(g1236_p_spl_)
  );


  LA
  g_g1295_p
  (
    .dout(g1295_p),
    .din1(G11_p_spl_100),
    .din2(G26_p_spl_101)
  );


  FA
  g_g1295_n
  (
    .dout(g1295_n),
    .din1(G11_n_spl_100),
    .din2(G26_n_spl_101)
  );


  LA
  g_g1296_p
  (
    .dout(g1296_p),
    .din1(g1227_n_spl_),
    .din2(g1230_n_spl_)
  );


  FA
  g_g1296_n
  (
    .dout(g1296_n),
    .din1(g1227_p_spl_),
    .din2(g1230_p_spl_)
  );


  LA
  g_g1297_p
  (
    .dout(g1297_p),
    .din1(G12_p_spl_100),
    .din2(G25_p_spl_101)
  );


  FA
  g_g1297_n
  (
    .dout(g1297_n),
    .din1(G12_n_spl_100),
    .din2(G25_n_spl_101)
  );


  LA
  g_g1298_p
  (
    .dout(g1298_p),
    .din1(g1221_n_spl_),
    .din2(g1224_n_spl_)
  );


  FA
  g_g1298_n
  (
    .dout(g1298_n),
    .din1(g1221_p_spl_),
    .din2(g1224_p_spl_)
  );


  LA
  g_g1299_p
  (
    .dout(g1299_p),
    .din1(G13_p_spl_011),
    .din2(G24_p_spl_110)
  );


  FA
  g_g1299_n
  (
    .dout(g1299_n),
    .din1(G13_n_spl_011),
    .din2(G24_n_spl_110)
  );


  LA
  g_g1300_p
  (
    .dout(g1300_p),
    .din1(g1215_n_spl_),
    .din2(g1218_n_spl_)
  );


  FA
  g_g1300_n
  (
    .dout(g1300_n),
    .din1(g1215_p_spl_),
    .din2(g1218_p_spl_)
  );


  LA
  g_g1301_p
  (
    .dout(g1301_p),
    .din1(G14_p_spl_011),
    .din2(G23_p_spl_110)
  );


  FA
  g_g1301_n
  (
    .dout(g1301_n),
    .din1(G14_n_spl_011),
    .din2(G23_n_spl_110)
  );


  LA
  g_g1302_p
  (
    .dout(g1302_p),
    .din1(g1209_n_spl_),
    .din2(g1212_n_spl_)
  );


  FA
  g_g1302_n
  (
    .dout(g1302_n),
    .din1(g1209_p_spl_),
    .din2(g1212_p_spl_)
  );


  LA
  g_g1303_p
  (
    .dout(g1303_p),
    .din1(G15_p_spl_010),
    .din2(G22_p_spl_111)
  );


  FA
  g_g1303_n
  (
    .dout(g1303_n),
    .din1(G15_n_spl_010),
    .din2(G22_n_spl_111)
  );


  LA
  g_g1304_p
  (
    .dout(g1304_p),
    .din1(G16_p_spl_010),
    .din2(G21_p_spl_111)
  );


  FA
  g_g1304_n
  (
    .dout(g1304_n),
    .din1(G16_n_spl_010),
    .din2(G21_n_spl_111)
  );


  LA
  g_g1305_p
  (
    .dout(g1305_p),
    .din1(g1203_n_spl_),
    .din2(g1206_n_spl_)
  );


  FA
  g_g1305_n
  (
    .dout(g1305_n),
    .din1(g1203_p_spl_),
    .din2(g1206_p_spl_)
  );


  LA
  g_g1306_p
  (
    .dout(g1306_p),
    .din1(g1304_n_spl_),
    .din2(g1305_n_spl_)
  );


  FA
  g_g1306_n
  (
    .dout(g1306_n),
    .din1(g1304_p_spl_),
    .din2(g1305_p_spl_)
  );


  LA
  g_g1307_p
  (
    .dout(g1307_p),
    .din1(g1304_p_spl_),
    .din2(g1305_p_spl_)
  );


  FA
  g_g1307_n
  (
    .dout(g1307_n),
    .din1(g1304_n_spl_),
    .din2(g1305_n_spl_)
  );


  LA
  g_g1308_p
  (
    .dout(g1308_p),
    .din1(g1306_n_spl_),
    .din2(g1307_n)
  );


  FA
  g_g1308_n
  (
    .dout(g1308_n),
    .din1(g1306_p_spl_),
    .din2(g1307_p)
  );


  LA
  g_g1309_p
  (
    .dout(g1309_p),
    .din1(g1303_n_spl_),
    .din2(g1308_p_spl_)
  );


  FA
  g_g1309_n
  (
    .dout(g1309_n),
    .din1(g1303_p_spl_),
    .din2(g1308_n_spl_)
  );


  LA
  g_g1310_p
  (
    .dout(g1310_p),
    .din1(g1303_p_spl_),
    .din2(g1308_n_spl_)
  );


  FA
  g_g1310_n
  (
    .dout(g1310_n),
    .din1(g1303_n_spl_),
    .din2(g1308_p_spl_)
  );


  LA
  g_g1311_p
  (
    .dout(g1311_p),
    .din1(g1309_n_spl_),
    .din2(g1310_n)
  );


  FA
  g_g1311_n
  (
    .dout(g1311_n),
    .din1(g1309_p_spl_),
    .din2(g1310_p)
  );


  LA
  g_g1312_p
  (
    .dout(g1312_p),
    .din1(g1302_n_spl_),
    .din2(g1311_p_spl_)
  );


  FA
  g_g1312_n
  (
    .dout(g1312_n),
    .din1(g1302_p_spl_),
    .din2(g1311_n_spl_)
  );


  LA
  g_g1313_p
  (
    .dout(g1313_p),
    .din1(g1302_p_spl_),
    .din2(g1311_n_spl_)
  );


  FA
  g_g1313_n
  (
    .dout(g1313_n),
    .din1(g1302_n_spl_),
    .din2(g1311_p_spl_)
  );


  LA
  g_g1314_p
  (
    .dout(g1314_p),
    .din1(g1312_n_spl_),
    .din2(g1313_n)
  );


  FA
  g_g1314_n
  (
    .dout(g1314_n),
    .din1(g1312_p_spl_),
    .din2(g1313_p)
  );


  LA
  g_g1315_p
  (
    .dout(g1315_p),
    .din1(g1301_n_spl_),
    .din2(g1314_p_spl_)
  );


  FA
  g_g1315_n
  (
    .dout(g1315_n),
    .din1(g1301_p_spl_),
    .din2(g1314_n_spl_)
  );


  LA
  g_g1316_p
  (
    .dout(g1316_p),
    .din1(g1301_p_spl_),
    .din2(g1314_n_spl_)
  );


  FA
  g_g1316_n
  (
    .dout(g1316_n),
    .din1(g1301_n_spl_),
    .din2(g1314_p_spl_)
  );


  LA
  g_g1317_p
  (
    .dout(g1317_p),
    .din1(g1315_n_spl_),
    .din2(g1316_n)
  );


  FA
  g_g1317_n
  (
    .dout(g1317_n),
    .din1(g1315_p_spl_),
    .din2(g1316_p)
  );


  LA
  g_g1318_p
  (
    .dout(g1318_p),
    .din1(g1300_n_spl_),
    .din2(g1317_p_spl_)
  );


  FA
  g_g1318_n
  (
    .dout(g1318_n),
    .din1(g1300_p_spl_),
    .din2(g1317_n_spl_)
  );


  LA
  g_g1319_p
  (
    .dout(g1319_p),
    .din1(g1300_p_spl_),
    .din2(g1317_n_spl_)
  );


  FA
  g_g1319_n
  (
    .dout(g1319_n),
    .din1(g1300_n_spl_),
    .din2(g1317_p_spl_)
  );


  LA
  g_g1320_p
  (
    .dout(g1320_p),
    .din1(g1318_n_spl_),
    .din2(g1319_n)
  );


  FA
  g_g1320_n
  (
    .dout(g1320_n),
    .din1(g1318_p_spl_),
    .din2(g1319_p)
  );


  LA
  g_g1321_p
  (
    .dout(g1321_p),
    .din1(g1299_n_spl_),
    .din2(g1320_p_spl_)
  );


  FA
  g_g1321_n
  (
    .dout(g1321_n),
    .din1(g1299_p_spl_),
    .din2(g1320_n_spl_)
  );


  LA
  g_g1322_p
  (
    .dout(g1322_p),
    .din1(g1299_p_spl_),
    .din2(g1320_n_spl_)
  );


  FA
  g_g1322_n
  (
    .dout(g1322_n),
    .din1(g1299_n_spl_),
    .din2(g1320_p_spl_)
  );


  LA
  g_g1323_p
  (
    .dout(g1323_p),
    .din1(g1321_n_spl_),
    .din2(g1322_n)
  );


  FA
  g_g1323_n
  (
    .dout(g1323_n),
    .din1(g1321_p_spl_),
    .din2(g1322_p)
  );


  LA
  g_g1324_p
  (
    .dout(g1324_p),
    .din1(g1298_n_spl_),
    .din2(g1323_p_spl_)
  );


  FA
  g_g1324_n
  (
    .dout(g1324_n),
    .din1(g1298_p_spl_),
    .din2(g1323_n_spl_)
  );


  LA
  g_g1325_p
  (
    .dout(g1325_p),
    .din1(g1298_p_spl_),
    .din2(g1323_n_spl_)
  );


  FA
  g_g1325_n
  (
    .dout(g1325_n),
    .din1(g1298_n_spl_),
    .din2(g1323_p_spl_)
  );


  LA
  g_g1326_p
  (
    .dout(g1326_p),
    .din1(g1324_n_spl_),
    .din2(g1325_n)
  );


  FA
  g_g1326_n
  (
    .dout(g1326_n),
    .din1(g1324_p_spl_),
    .din2(g1325_p)
  );


  LA
  g_g1327_p
  (
    .dout(g1327_p),
    .din1(g1297_n_spl_),
    .din2(g1326_p_spl_)
  );


  FA
  g_g1327_n
  (
    .dout(g1327_n),
    .din1(g1297_p_spl_),
    .din2(g1326_n_spl_)
  );


  LA
  g_g1328_p
  (
    .dout(g1328_p),
    .din1(g1297_p_spl_),
    .din2(g1326_n_spl_)
  );


  FA
  g_g1328_n
  (
    .dout(g1328_n),
    .din1(g1297_n_spl_),
    .din2(g1326_p_spl_)
  );


  LA
  g_g1329_p
  (
    .dout(g1329_p),
    .din1(g1327_n_spl_),
    .din2(g1328_n)
  );


  FA
  g_g1329_n
  (
    .dout(g1329_n),
    .din1(g1327_p_spl_),
    .din2(g1328_p)
  );


  LA
  g_g1330_p
  (
    .dout(g1330_p),
    .din1(g1296_n_spl_),
    .din2(g1329_p_spl_)
  );


  FA
  g_g1330_n
  (
    .dout(g1330_n),
    .din1(g1296_p_spl_),
    .din2(g1329_n_spl_)
  );


  LA
  g_g1331_p
  (
    .dout(g1331_p),
    .din1(g1296_p_spl_),
    .din2(g1329_n_spl_)
  );


  FA
  g_g1331_n
  (
    .dout(g1331_n),
    .din1(g1296_n_spl_),
    .din2(g1329_p_spl_)
  );


  LA
  g_g1332_p
  (
    .dout(g1332_p),
    .din1(g1330_n_spl_),
    .din2(g1331_n)
  );


  FA
  g_g1332_n
  (
    .dout(g1332_n),
    .din1(g1330_p_spl_),
    .din2(g1331_p)
  );


  LA
  g_g1333_p
  (
    .dout(g1333_p),
    .din1(g1295_n_spl_),
    .din2(g1332_p_spl_)
  );


  FA
  g_g1333_n
  (
    .dout(g1333_n),
    .din1(g1295_p_spl_),
    .din2(g1332_n_spl_)
  );


  LA
  g_g1334_p
  (
    .dout(g1334_p),
    .din1(g1295_p_spl_),
    .din2(g1332_n_spl_)
  );


  FA
  g_g1334_n
  (
    .dout(g1334_n),
    .din1(g1295_n_spl_),
    .din2(g1332_p_spl_)
  );


  LA
  g_g1335_p
  (
    .dout(g1335_p),
    .din1(g1333_n_spl_),
    .din2(g1334_n)
  );


  FA
  g_g1335_n
  (
    .dout(g1335_n),
    .din1(g1333_p_spl_),
    .din2(g1334_p)
  );


  LA
  g_g1336_p
  (
    .dout(g1336_p),
    .din1(g1294_n_spl_),
    .din2(g1335_p_spl_)
  );


  FA
  g_g1336_n
  (
    .dout(g1336_n),
    .din1(g1294_p_spl_),
    .din2(g1335_n_spl_)
  );


  LA
  g_g1337_p
  (
    .dout(g1337_p),
    .din1(g1294_p_spl_),
    .din2(g1335_n_spl_)
  );


  FA
  g_g1337_n
  (
    .dout(g1337_n),
    .din1(g1294_n_spl_),
    .din2(g1335_p_spl_)
  );


  LA
  g_g1338_p
  (
    .dout(g1338_p),
    .din1(g1336_n_spl_),
    .din2(g1337_n)
  );


  FA
  g_g1338_n
  (
    .dout(g1338_n),
    .din1(g1336_p_spl_),
    .din2(g1337_p)
  );


  LA
  g_g1339_p
  (
    .dout(g1339_p),
    .din1(g1293_n_spl_),
    .din2(g1338_p_spl_)
  );


  FA
  g_g1339_n
  (
    .dout(g1339_n),
    .din1(g1293_p_spl_),
    .din2(g1338_n_spl_)
  );


  LA
  g_g1340_p
  (
    .dout(g1340_p),
    .din1(g1293_p_spl_),
    .din2(g1338_n_spl_)
  );


  FA
  g_g1340_n
  (
    .dout(g1340_n),
    .din1(g1293_n_spl_),
    .din2(g1338_p_spl_)
  );


  LA
  g_g1341_p
  (
    .dout(g1341_p),
    .din1(g1339_n_spl_),
    .din2(g1340_n)
  );


  FA
  g_g1341_n
  (
    .dout(g1341_n),
    .din1(g1339_p_spl_),
    .din2(g1340_p)
  );


  LA
  g_g1342_p
  (
    .dout(g1342_p),
    .din1(g1292_n_spl_),
    .din2(g1341_p_spl_)
  );


  FA
  g_g1342_n
  (
    .dout(g1342_n),
    .din1(g1292_p_spl_),
    .din2(g1341_n_spl_)
  );


  LA
  g_g1343_p
  (
    .dout(g1343_p),
    .din1(g1292_p_spl_),
    .din2(g1341_n_spl_)
  );


  FA
  g_g1343_n
  (
    .dout(g1343_n),
    .din1(g1292_n_spl_),
    .din2(g1341_p_spl_)
  );


  LA
  g_g1344_p
  (
    .dout(g1344_p),
    .din1(g1342_n_spl_),
    .din2(g1343_n)
  );


  FA
  g_g1344_n
  (
    .dout(g1344_n),
    .din1(g1342_p_spl_),
    .din2(g1343_p)
  );


  LA
  g_g1345_p
  (
    .dout(g1345_p),
    .din1(g1291_n_spl_),
    .din2(g1344_p_spl_)
  );


  FA
  g_g1345_n
  (
    .dout(g1345_n),
    .din1(g1291_p_spl_),
    .din2(g1344_n_spl_)
  );


  LA
  g_g1346_p
  (
    .dout(g1346_p),
    .din1(g1291_p_spl_),
    .din2(g1344_n_spl_)
  );


  FA
  g_g1346_n
  (
    .dout(g1346_n),
    .din1(g1291_n_spl_),
    .din2(g1344_p_spl_)
  );


  LA
  g_g1347_p
  (
    .dout(g1347_p),
    .din1(g1345_n_spl_),
    .din2(g1346_n)
  );


  FA
  g_g1347_n
  (
    .dout(g1347_n),
    .din1(g1345_p_spl_),
    .din2(g1346_p)
  );


  LA
  g_g1348_p
  (
    .dout(g1348_p),
    .din1(g1290_n_spl_),
    .din2(g1347_p_spl_)
  );


  FA
  g_g1348_n
  (
    .dout(g1348_n),
    .din1(g1290_p_spl_),
    .din2(g1347_n_spl_)
  );


  LA
  g_g1349_p
  (
    .dout(g1349_p),
    .din1(g1290_p_spl_),
    .din2(g1347_n_spl_)
  );


  FA
  g_g1349_n
  (
    .dout(g1349_n),
    .din1(g1290_n_spl_),
    .din2(g1347_p_spl_)
  );


  LA
  g_g1350_p
  (
    .dout(g1350_p),
    .din1(g1348_n_spl_),
    .din2(g1349_n)
  );


  FA
  g_g1350_n
  (
    .dout(g1350_n),
    .din1(g1348_p_spl_),
    .din2(g1349_p)
  );


  LA
  g_g1351_p
  (
    .dout(g1351_p),
    .din1(g1289_n_spl_),
    .din2(g1350_p_spl_)
  );


  FA
  g_g1351_n
  (
    .dout(g1351_n),
    .din1(g1289_p_spl_),
    .din2(g1350_n_spl_)
  );


  LA
  g_g1352_p
  (
    .dout(g1352_p),
    .din1(g1289_p_spl_),
    .din2(g1350_n_spl_)
  );


  FA
  g_g1352_n
  (
    .dout(g1352_n),
    .din1(g1289_n_spl_),
    .din2(g1350_p_spl_)
  );


  LA
  g_g1353_p
  (
    .dout(g1353_p),
    .din1(g1351_n_spl_),
    .din2(g1352_n)
  );


  FA
  g_g1353_n
  (
    .dout(g1353_n),
    .din1(g1351_p_spl_),
    .din2(g1352_p)
  );


  LA
  g_g1354_p
  (
    .dout(g1354_p),
    .din1(g1288_n_spl_),
    .din2(g1353_p_spl_)
  );


  FA
  g_g1354_n
  (
    .dout(g1354_n),
    .din1(g1288_p_spl_),
    .din2(g1353_n_spl_)
  );


  LA
  g_g1355_p
  (
    .dout(g1355_p),
    .din1(g1288_p_spl_),
    .din2(g1353_n_spl_)
  );


  FA
  g_g1355_n
  (
    .dout(g1355_n),
    .din1(g1288_n_spl_),
    .din2(g1353_p_spl_)
  );


  LA
  g_g1356_p
  (
    .dout(g1356_p),
    .din1(g1354_n_spl_),
    .din2(g1355_n)
  );


  FA
  g_g1356_n
  (
    .dout(g1356_n),
    .din1(g1354_p_spl_),
    .din2(g1355_p)
  );


  LA
  g_g1357_p
  (
    .dout(g1357_p),
    .din1(g1287_n_spl_),
    .din2(g1356_p_spl_)
  );


  FA
  g_g1357_n
  (
    .dout(g1357_n),
    .din1(g1287_p_spl_),
    .din2(g1356_n_spl_)
  );


  LA
  g_g1358_p
  (
    .dout(g1358_p),
    .din1(g1287_p_spl_),
    .din2(g1356_n_spl_)
  );


  FA
  g_g1358_n
  (
    .dout(g1358_n),
    .din1(g1287_n_spl_),
    .din2(g1356_p_spl_)
  );


  LA
  g_g1359_p
  (
    .dout(g1359_p),
    .din1(g1357_n_spl_),
    .din2(g1358_n)
  );


  FA
  g_g1359_n
  (
    .dout(g1359_n),
    .din1(g1357_p_spl_),
    .din2(g1358_p)
  );


  LA
  g_g1360_p
  (
    .dout(g1360_p),
    .din1(g1286_n_spl_),
    .din2(g1359_p_spl_)
  );


  FA
  g_g1360_n
  (
    .dout(g1360_n),
    .din1(g1286_p_spl_),
    .din2(g1359_n_spl_)
  );


  LA
  g_g1361_p
  (
    .dout(g1361_p),
    .din1(g1286_p_spl_),
    .din2(g1359_n_spl_)
  );


  FA
  g_g1361_n
  (
    .dout(g1361_n),
    .din1(g1286_n_spl_),
    .din2(g1359_p_spl_)
  );


  LA
  g_g1362_p
  (
    .dout(g1362_p),
    .din1(g1360_n_spl_),
    .din2(g1361_n)
  );


  FA
  g_g1362_n
  (
    .dout(g1362_n),
    .din1(g1360_p_spl_),
    .din2(g1361_p)
  );


  LA
  g_g1363_p
  (
    .dout(g1363_p),
    .din1(g1285_n_spl_),
    .din2(g1362_p_spl_)
  );


  FA
  g_g1363_n
  (
    .dout(g1363_n),
    .din1(g1285_p_spl_),
    .din2(g1362_n_spl_)
  );


  LA
  g_g1364_p
  (
    .dout(g1364_p),
    .din1(g1285_p_spl_),
    .din2(g1362_n_spl_)
  );


  FA
  g_g1364_n
  (
    .dout(g1364_n),
    .din1(g1285_n_spl_),
    .din2(g1362_p_spl_)
  );


  LA
  g_g1365_p
  (
    .dout(g1365_p),
    .din1(g1363_n_spl_),
    .din2(g1364_n)
  );


  FA
  g_g1365_n
  (
    .dout(g1365_n),
    .din1(g1363_p_spl_),
    .din2(g1364_p)
  );


  LA
  g_g1366_p
  (
    .dout(g1366_p),
    .din1(g1284_n_spl_),
    .din2(g1365_p_spl_)
  );


  FA
  g_g1366_n
  (
    .dout(g1366_n),
    .din1(g1284_p_spl_),
    .din2(g1365_n_spl_)
  );


  LA
  g_g1367_p
  (
    .dout(g1367_p),
    .din1(g1284_p_spl_),
    .din2(g1365_n_spl_)
  );


  FA
  g_g1367_n
  (
    .dout(g1367_n),
    .din1(g1284_n_spl_),
    .din2(g1365_p_spl_)
  );


  LA
  g_g1368_p
  (
    .dout(g1368_p),
    .din1(g1366_n_spl_),
    .din2(g1367_n)
  );


  FA
  g_g1368_n
  (
    .dout(g1368_n),
    .din1(g1366_p_spl_),
    .din2(g1367_p)
  );


  LA
  g_g1369_p
  (
    .dout(g1369_p),
    .din1(g1283_n_spl_),
    .din2(g1368_p_spl_)
  );


  FA
  g_g1369_n
  (
    .dout(g1369_n),
    .din1(g1283_p_spl_),
    .din2(g1368_n_spl_)
  );


  LA
  g_g1370_p
  (
    .dout(g1370_p),
    .din1(g1283_p_spl_),
    .din2(g1368_n_spl_)
  );


  FA
  g_g1370_n
  (
    .dout(g1370_n),
    .din1(g1283_n_spl_),
    .din2(g1368_p_spl_)
  );


  LA
  g_g1371_p
  (
    .dout(g1371_p),
    .din1(g1369_n_spl_),
    .din2(g1370_n)
  );


  FA
  g_g1371_n
  (
    .dout(g1371_n),
    .din1(g1369_p_spl_),
    .din2(g1370_p)
  );


  LA
  g_g1372_p
  (
    .dout(g1372_p),
    .din1(g1282_n_spl_),
    .din2(g1371_p_spl_)
  );


  FA
  g_g1372_n
  (
    .dout(g1372_n),
    .din1(g1282_p_spl_),
    .din2(g1371_n_spl_)
  );


  LA
  g_g1373_p
  (
    .dout(g1373_p),
    .din1(g1282_p_spl_),
    .din2(g1371_n_spl_)
  );


  FA
  g_g1373_n
  (
    .dout(g1373_n),
    .din1(g1282_n_spl_),
    .din2(g1371_p_spl_)
  );


  LA
  g_g1374_p
  (
    .dout(g1374_p),
    .din1(g1372_n_spl_),
    .din2(g1373_n)
  );


  FA
  g_g1374_n
  (
    .dout(g1374_n),
    .din1(g1372_p_spl_),
    .din2(g1373_p)
  );


  LA
  g_g1375_p
  (
    .dout(g1375_p),
    .din1(g1281_n),
    .din2(g1374_p)
  );


  FA
  g_g1375_n
  (
    .dout(g1375_n),
    .din1(g1281_p_spl_),
    .din2(g1374_n_spl_)
  );


  LA
  g_g1376_p
  (
    .dout(g1376_p),
    .din1(g1281_p_spl_),
    .din2(g1374_n_spl_)
  );


  FA
  g_g1377_n
  (
    .dout(g1377_n),
    .din1(g1375_p_spl_),
    .din2(g1376_p)
  );


  LA
  g_g1378_p
  (
    .dout(g1378_p),
    .din1(g1372_n_spl_),
    .din2(g1375_n)
  );


  FA
  g_g1378_n
  (
    .dout(g1378_n),
    .din1(g1372_p_spl_),
    .din2(g1375_p_spl_)
  );


  LA
  g_g1379_p
  (
    .dout(g1379_p),
    .din1(g1366_n_spl_),
    .din2(g1369_n_spl_)
  );


  FA
  g_g1379_n
  (
    .dout(g1379_n),
    .din1(g1366_p_spl_),
    .din2(g1369_p_spl_)
  );


  LA
  g_g1380_p
  (
    .dout(g1380_p),
    .din1(G6_p_spl_111),
    .din2(G32_p_spl_010)
  );


  FA
  g_g1380_n
  (
    .dout(g1380_n),
    .din1(G6_n_spl_111),
    .din2(G32_n_spl_010)
  );


  LA
  g_g1381_p
  (
    .dout(g1381_p),
    .din1(g1360_n_spl_),
    .din2(g1363_n_spl_)
  );


  FA
  g_g1381_n
  (
    .dout(g1381_n),
    .din1(g1360_p_spl_),
    .din2(g1363_p_spl_)
  );


  LA
  g_g1382_p
  (
    .dout(g1382_p),
    .din1(G7_p_spl_111),
    .din2(G31_p_spl_011)
  );


  FA
  g_g1382_n
  (
    .dout(g1382_n),
    .din1(G7_n_spl_111),
    .din2(G31_n_spl_011)
  );


  LA
  g_g1383_p
  (
    .dout(g1383_p),
    .din1(g1354_n_spl_),
    .din2(g1357_n_spl_)
  );


  FA
  g_g1383_n
  (
    .dout(g1383_n),
    .din1(g1354_p_spl_),
    .din2(g1357_p_spl_)
  );


  LA
  g_g1384_p
  (
    .dout(g1384_p),
    .din1(G8_p_spl_110),
    .din2(G30_p_spl_011)
  );


  FA
  g_g1384_n
  (
    .dout(g1384_n),
    .din1(G8_n_spl_110),
    .din2(G30_n_spl_011)
  );


  LA
  g_g1385_p
  (
    .dout(g1385_p),
    .din1(g1348_n_spl_),
    .din2(g1351_n_spl_)
  );


  FA
  g_g1385_n
  (
    .dout(g1385_n),
    .din1(g1348_p_spl_),
    .din2(g1351_p_spl_)
  );


  LA
  g_g1386_p
  (
    .dout(g1386_p),
    .din1(G9_p_spl_110),
    .din2(G29_p_spl_100)
  );


  FA
  g_g1386_n
  (
    .dout(g1386_n),
    .din1(G9_n_spl_110),
    .din2(G29_n_spl_100)
  );


  LA
  g_g1387_p
  (
    .dout(g1387_p),
    .din1(g1342_n_spl_),
    .din2(g1345_n_spl_)
  );


  FA
  g_g1387_n
  (
    .dout(g1387_n),
    .din1(g1342_p_spl_),
    .din2(g1345_p_spl_)
  );


  LA
  g_g1388_p
  (
    .dout(g1388_p),
    .din1(G10_p_spl_101),
    .din2(G28_p_spl_100)
  );


  FA
  g_g1388_n
  (
    .dout(g1388_n),
    .din1(G10_n_spl_101),
    .din2(G28_n_spl_100)
  );


  LA
  g_g1389_p
  (
    .dout(g1389_p),
    .din1(g1336_n_spl_),
    .din2(g1339_n_spl_)
  );


  FA
  g_g1389_n
  (
    .dout(g1389_n),
    .din1(g1336_p_spl_),
    .din2(g1339_p_spl_)
  );


  LA
  g_g1390_p
  (
    .dout(g1390_p),
    .din1(G11_p_spl_101),
    .din2(G27_p_spl_101)
  );


  FA
  g_g1390_n
  (
    .dout(g1390_n),
    .din1(G11_n_spl_101),
    .din2(G27_n_spl_101)
  );


  LA
  g_g1391_p
  (
    .dout(g1391_p),
    .din1(g1330_n_spl_),
    .din2(g1333_n_spl_)
  );


  FA
  g_g1391_n
  (
    .dout(g1391_n),
    .din1(g1330_p_spl_),
    .din2(g1333_p_spl_)
  );


  LA
  g_g1392_p
  (
    .dout(g1392_p),
    .din1(G12_p_spl_100),
    .din2(G26_p_spl_101)
  );


  FA
  g_g1392_n
  (
    .dout(g1392_n),
    .din1(G12_n_spl_100),
    .din2(G26_n_spl_101)
  );


  LA
  g_g1393_p
  (
    .dout(g1393_p),
    .din1(g1324_n_spl_),
    .din2(g1327_n_spl_)
  );


  FA
  g_g1393_n
  (
    .dout(g1393_n),
    .din1(g1324_p_spl_),
    .din2(g1327_p_spl_)
  );


  LA
  g_g1394_p
  (
    .dout(g1394_p),
    .din1(G13_p_spl_100),
    .din2(G25_p_spl_110)
  );


  FA
  g_g1394_n
  (
    .dout(g1394_n),
    .din1(G13_n_spl_100),
    .din2(G25_n_spl_110)
  );


  LA
  g_g1395_p
  (
    .dout(g1395_p),
    .din1(g1318_n_spl_),
    .din2(g1321_n_spl_)
  );


  FA
  g_g1395_n
  (
    .dout(g1395_n),
    .din1(g1318_p_spl_),
    .din2(g1321_p_spl_)
  );


  LA
  g_g1396_p
  (
    .dout(g1396_p),
    .din1(G14_p_spl_011),
    .din2(G24_p_spl_110)
  );


  FA
  g_g1396_n
  (
    .dout(g1396_n),
    .din1(G14_n_spl_011),
    .din2(G24_n_spl_110)
  );


  LA
  g_g1397_p
  (
    .dout(g1397_p),
    .din1(g1312_n_spl_),
    .din2(g1315_n_spl_)
  );


  FA
  g_g1397_n
  (
    .dout(g1397_n),
    .din1(g1312_p_spl_),
    .din2(g1315_p_spl_)
  );


  LA
  g_g1398_p
  (
    .dout(g1398_p),
    .din1(G15_p_spl_011),
    .din2(G23_p_spl_111)
  );


  FA
  g_g1398_n
  (
    .dout(g1398_n),
    .din1(G15_n_spl_011),
    .din2(G23_n_spl_111)
  );


  LA
  g_g1399_p
  (
    .dout(g1399_p),
    .din1(G16_p_spl_010),
    .din2(G22_p_spl_111)
  );


  FA
  g_g1399_n
  (
    .dout(g1399_n),
    .din1(G16_n_spl_010),
    .din2(G22_n_spl_111)
  );


  LA
  g_g1400_p
  (
    .dout(g1400_p),
    .din1(g1306_n_spl_),
    .din2(g1309_n_spl_)
  );


  FA
  g_g1400_n
  (
    .dout(g1400_n),
    .din1(g1306_p_spl_),
    .din2(g1309_p_spl_)
  );


  LA
  g_g1401_p
  (
    .dout(g1401_p),
    .din1(g1399_n_spl_),
    .din2(g1400_n_spl_)
  );


  FA
  g_g1401_n
  (
    .dout(g1401_n),
    .din1(g1399_p_spl_),
    .din2(g1400_p_spl_)
  );


  LA
  g_g1402_p
  (
    .dout(g1402_p),
    .din1(g1399_p_spl_),
    .din2(g1400_p_spl_)
  );


  FA
  g_g1402_n
  (
    .dout(g1402_n),
    .din1(g1399_n_spl_),
    .din2(g1400_n_spl_)
  );


  LA
  g_g1403_p
  (
    .dout(g1403_p),
    .din1(g1401_n_spl_),
    .din2(g1402_n)
  );


  FA
  g_g1403_n
  (
    .dout(g1403_n),
    .din1(g1401_p_spl_),
    .din2(g1402_p)
  );


  LA
  g_g1404_p
  (
    .dout(g1404_p),
    .din1(g1398_n_spl_),
    .din2(g1403_p_spl_)
  );


  FA
  g_g1404_n
  (
    .dout(g1404_n),
    .din1(g1398_p_spl_),
    .din2(g1403_n_spl_)
  );


  LA
  g_g1405_p
  (
    .dout(g1405_p),
    .din1(g1398_p_spl_),
    .din2(g1403_n_spl_)
  );


  FA
  g_g1405_n
  (
    .dout(g1405_n),
    .din1(g1398_n_spl_),
    .din2(g1403_p_spl_)
  );


  LA
  g_g1406_p
  (
    .dout(g1406_p),
    .din1(g1404_n_spl_),
    .din2(g1405_n)
  );


  FA
  g_g1406_n
  (
    .dout(g1406_n),
    .din1(g1404_p_spl_),
    .din2(g1405_p)
  );


  LA
  g_g1407_p
  (
    .dout(g1407_p),
    .din1(g1397_n_spl_),
    .din2(g1406_p_spl_)
  );


  FA
  g_g1407_n
  (
    .dout(g1407_n),
    .din1(g1397_p_spl_),
    .din2(g1406_n_spl_)
  );


  LA
  g_g1408_p
  (
    .dout(g1408_p),
    .din1(g1397_p_spl_),
    .din2(g1406_n_spl_)
  );


  FA
  g_g1408_n
  (
    .dout(g1408_n),
    .din1(g1397_n_spl_),
    .din2(g1406_p_spl_)
  );


  LA
  g_g1409_p
  (
    .dout(g1409_p),
    .din1(g1407_n_spl_),
    .din2(g1408_n)
  );


  FA
  g_g1409_n
  (
    .dout(g1409_n),
    .din1(g1407_p_spl_),
    .din2(g1408_p)
  );


  LA
  g_g1410_p
  (
    .dout(g1410_p),
    .din1(g1396_n_spl_),
    .din2(g1409_p_spl_)
  );


  FA
  g_g1410_n
  (
    .dout(g1410_n),
    .din1(g1396_p_spl_),
    .din2(g1409_n_spl_)
  );


  LA
  g_g1411_p
  (
    .dout(g1411_p),
    .din1(g1396_p_spl_),
    .din2(g1409_n_spl_)
  );


  FA
  g_g1411_n
  (
    .dout(g1411_n),
    .din1(g1396_n_spl_),
    .din2(g1409_p_spl_)
  );


  LA
  g_g1412_p
  (
    .dout(g1412_p),
    .din1(g1410_n_spl_),
    .din2(g1411_n)
  );


  FA
  g_g1412_n
  (
    .dout(g1412_n),
    .din1(g1410_p_spl_),
    .din2(g1411_p)
  );


  LA
  g_g1413_p
  (
    .dout(g1413_p),
    .din1(g1395_n_spl_),
    .din2(g1412_p_spl_)
  );


  FA
  g_g1413_n
  (
    .dout(g1413_n),
    .din1(g1395_p_spl_),
    .din2(g1412_n_spl_)
  );


  LA
  g_g1414_p
  (
    .dout(g1414_p),
    .din1(g1395_p_spl_),
    .din2(g1412_n_spl_)
  );


  FA
  g_g1414_n
  (
    .dout(g1414_n),
    .din1(g1395_n_spl_),
    .din2(g1412_p_spl_)
  );


  LA
  g_g1415_p
  (
    .dout(g1415_p),
    .din1(g1413_n_spl_),
    .din2(g1414_n)
  );


  FA
  g_g1415_n
  (
    .dout(g1415_n),
    .din1(g1413_p_spl_),
    .din2(g1414_p)
  );


  LA
  g_g1416_p
  (
    .dout(g1416_p),
    .din1(g1394_n_spl_),
    .din2(g1415_p_spl_)
  );


  FA
  g_g1416_n
  (
    .dout(g1416_n),
    .din1(g1394_p_spl_),
    .din2(g1415_n_spl_)
  );


  LA
  g_g1417_p
  (
    .dout(g1417_p),
    .din1(g1394_p_spl_),
    .din2(g1415_n_spl_)
  );


  FA
  g_g1417_n
  (
    .dout(g1417_n),
    .din1(g1394_n_spl_),
    .din2(g1415_p_spl_)
  );


  LA
  g_g1418_p
  (
    .dout(g1418_p),
    .din1(g1416_n_spl_),
    .din2(g1417_n)
  );


  FA
  g_g1418_n
  (
    .dout(g1418_n),
    .din1(g1416_p_spl_),
    .din2(g1417_p)
  );


  LA
  g_g1419_p
  (
    .dout(g1419_p),
    .din1(g1393_n_spl_),
    .din2(g1418_p_spl_)
  );


  FA
  g_g1419_n
  (
    .dout(g1419_n),
    .din1(g1393_p_spl_),
    .din2(g1418_n_spl_)
  );


  LA
  g_g1420_p
  (
    .dout(g1420_p),
    .din1(g1393_p_spl_),
    .din2(g1418_n_spl_)
  );


  FA
  g_g1420_n
  (
    .dout(g1420_n),
    .din1(g1393_n_spl_),
    .din2(g1418_p_spl_)
  );


  LA
  g_g1421_p
  (
    .dout(g1421_p),
    .din1(g1419_n_spl_),
    .din2(g1420_n)
  );


  FA
  g_g1421_n
  (
    .dout(g1421_n),
    .din1(g1419_p_spl_),
    .din2(g1420_p)
  );


  LA
  g_g1422_p
  (
    .dout(g1422_p),
    .din1(g1392_n_spl_),
    .din2(g1421_p_spl_)
  );


  FA
  g_g1422_n
  (
    .dout(g1422_n),
    .din1(g1392_p_spl_),
    .din2(g1421_n_spl_)
  );


  LA
  g_g1423_p
  (
    .dout(g1423_p),
    .din1(g1392_p_spl_),
    .din2(g1421_n_spl_)
  );


  FA
  g_g1423_n
  (
    .dout(g1423_n),
    .din1(g1392_n_spl_),
    .din2(g1421_p_spl_)
  );


  LA
  g_g1424_p
  (
    .dout(g1424_p),
    .din1(g1422_n_spl_),
    .din2(g1423_n)
  );


  FA
  g_g1424_n
  (
    .dout(g1424_n),
    .din1(g1422_p_spl_),
    .din2(g1423_p)
  );


  LA
  g_g1425_p
  (
    .dout(g1425_p),
    .din1(g1391_n_spl_),
    .din2(g1424_p_spl_)
  );


  FA
  g_g1425_n
  (
    .dout(g1425_n),
    .din1(g1391_p_spl_),
    .din2(g1424_n_spl_)
  );


  LA
  g_g1426_p
  (
    .dout(g1426_p),
    .din1(g1391_p_spl_),
    .din2(g1424_n_spl_)
  );


  FA
  g_g1426_n
  (
    .dout(g1426_n),
    .din1(g1391_n_spl_),
    .din2(g1424_p_spl_)
  );


  LA
  g_g1427_p
  (
    .dout(g1427_p),
    .din1(g1425_n_spl_),
    .din2(g1426_n)
  );


  FA
  g_g1427_n
  (
    .dout(g1427_n),
    .din1(g1425_p_spl_),
    .din2(g1426_p)
  );


  LA
  g_g1428_p
  (
    .dout(g1428_p),
    .din1(g1390_n_spl_),
    .din2(g1427_p_spl_)
  );


  FA
  g_g1428_n
  (
    .dout(g1428_n),
    .din1(g1390_p_spl_),
    .din2(g1427_n_spl_)
  );


  LA
  g_g1429_p
  (
    .dout(g1429_p),
    .din1(g1390_p_spl_),
    .din2(g1427_n_spl_)
  );


  FA
  g_g1429_n
  (
    .dout(g1429_n),
    .din1(g1390_n_spl_),
    .din2(g1427_p_spl_)
  );


  LA
  g_g1430_p
  (
    .dout(g1430_p),
    .din1(g1428_n_spl_),
    .din2(g1429_n)
  );


  FA
  g_g1430_n
  (
    .dout(g1430_n),
    .din1(g1428_p_spl_),
    .din2(g1429_p)
  );


  LA
  g_g1431_p
  (
    .dout(g1431_p),
    .din1(g1389_n_spl_),
    .din2(g1430_p_spl_)
  );


  FA
  g_g1431_n
  (
    .dout(g1431_n),
    .din1(g1389_p_spl_),
    .din2(g1430_n_spl_)
  );


  LA
  g_g1432_p
  (
    .dout(g1432_p),
    .din1(g1389_p_spl_),
    .din2(g1430_n_spl_)
  );


  FA
  g_g1432_n
  (
    .dout(g1432_n),
    .din1(g1389_n_spl_),
    .din2(g1430_p_spl_)
  );


  LA
  g_g1433_p
  (
    .dout(g1433_p),
    .din1(g1431_n_spl_),
    .din2(g1432_n)
  );


  FA
  g_g1433_n
  (
    .dout(g1433_n),
    .din1(g1431_p_spl_),
    .din2(g1432_p)
  );


  LA
  g_g1434_p
  (
    .dout(g1434_p),
    .din1(g1388_n_spl_),
    .din2(g1433_p_spl_)
  );


  FA
  g_g1434_n
  (
    .dout(g1434_n),
    .din1(g1388_p_spl_),
    .din2(g1433_n_spl_)
  );


  LA
  g_g1435_p
  (
    .dout(g1435_p),
    .din1(g1388_p_spl_),
    .din2(g1433_n_spl_)
  );


  FA
  g_g1435_n
  (
    .dout(g1435_n),
    .din1(g1388_n_spl_),
    .din2(g1433_p_spl_)
  );


  LA
  g_g1436_p
  (
    .dout(g1436_p),
    .din1(g1434_n_spl_),
    .din2(g1435_n)
  );


  FA
  g_g1436_n
  (
    .dout(g1436_n),
    .din1(g1434_p_spl_),
    .din2(g1435_p)
  );


  LA
  g_g1437_p
  (
    .dout(g1437_p),
    .din1(g1387_n_spl_),
    .din2(g1436_p_spl_)
  );


  FA
  g_g1437_n
  (
    .dout(g1437_n),
    .din1(g1387_p_spl_),
    .din2(g1436_n_spl_)
  );


  LA
  g_g1438_p
  (
    .dout(g1438_p),
    .din1(g1387_p_spl_),
    .din2(g1436_n_spl_)
  );


  FA
  g_g1438_n
  (
    .dout(g1438_n),
    .din1(g1387_n_spl_),
    .din2(g1436_p_spl_)
  );


  LA
  g_g1439_p
  (
    .dout(g1439_p),
    .din1(g1437_n_spl_),
    .din2(g1438_n)
  );


  FA
  g_g1439_n
  (
    .dout(g1439_n),
    .din1(g1437_p_spl_),
    .din2(g1438_p)
  );


  LA
  g_g1440_p
  (
    .dout(g1440_p),
    .din1(g1386_n_spl_),
    .din2(g1439_p_spl_)
  );


  FA
  g_g1440_n
  (
    .dout(g1440_n),
    .din1(g1386_p_spl_),
    .din2(g1439_n_spl_)
  );


  LA
  g_g1441_p
  (
    .dout(g1441_p),
    .din1(g1386_p_spl_),
    .din2(g1439_n_spl_)
  );


  FA
  g_g1441_n
  (
    .dout(g1441_n),
    .din1(g1386_n_spl_),
    .din2(g1439_p_spl_)
  );


  LA
  g_g1442_p
  (
    .dout(g1442_p),
    .din1(g1440_n_spl_),
    .din2(g1441_n)
  );


  FA
  g_g1442_n
  (
    .dout(g1442_n),
    .din1(g1440_p_spl_),
    .din2(g1441_p)
  );


  LA
  g_g1443_p
  (
    .dout(g1443_p),
    .din1(g1385_n_spl_),
    .din2(g1442_p_spl_)
  );


  FA
  g_g1443_n
  (
    .dout(g1443_n),
    .din1(g1385_p_spl_),
    .din2(g1442_n_spl_)
  );


  LA
  g_g1444_p
  (
    .dout(g1444_p),
    .din1(g1385_p_spl_),
    .din2(g1442_n_spl_)
  );


  FA
  g_g1444_n
  (
    .dout(g1444_n),
    .din1(g1385_n_spl_),
    .din2(g1442_p_spl_)
  );


  LA
  g_g1445_p
  (
    .dout(g1445_p),
    .din1(g1443_n_spl_),
    .din2(g1444_n)
  );


  FA
  g_g1445_n
  (
    .dout(g1445_n),
    .din1(g1443_p_spl_),
    .din2(g1444_p)
  );


  LA
  g_g1446_p
  (
    .dout(g1446_p),
    .din1(g1384_n_spl_),
    .din2(g1445_p_spl_)
  );


  FA
  g_g1446_n
  (
    .dout(g1446_n),
    .din1(g1384_p_spl_),
    .din2(g1445_n_spl_)
  );


  LA
  g_g1447_p
  (
    .dout(g1447_p),
    .din1(g1384_p_spl_),
    .din2(g1445_n_spl_)
  );


  FA
  g_g1447_n
  (
    .dout(g1447_n),
    .din1(g1384_n_spl_),
    .din2(g1445_p_spl_)
  );


  LA
  g_g1448_p
  (
    .dout(g1448_p),
    .din1(g1446_n_spl_),
    .din2(g1447_n)
  );


  FA
  g_g1448_n
  (
    .dout(g1448_n),
    .din1(g1446_p_spl_),
    .din2(g1447_p)
  );


  LA
  g_g1449_p
  (
    .dout(g1449_p),
    .din1(g1383_n_spl_),
    .din2(g1448_p_spl_)
  );


  FA
  g_g1449_n
  (
    .dout(g1449_n),
    .din1(g1383_p_spl_),
    .din2(g1448_n_spl_)
  );


  LA
  g_g1450_p
  (
    .dout(g1450_p),
    .din1(g1383_p_spl_),
    .din2(g1448_n_spl_)
  );


  FA
  g_g1450_n
  (
    .dout(g1450_n),
    .din1(g1383_n_spl_),
    .din2(g1448_p_spl_)
  );


  LA
  g_g1451_p
  (
    .dout(g1451_p),
    .din1(g1449_n_spl_),
    .din2(g1450_n)
  );


  FA
  g_g1451_n
  (
    .dout(g1451_n),
    .din1(g1449_p_spl_),
    .din2(g1450_p)
  );


  LA
  g_g1452_p
  (
    .dout(g1452_p),
    .din1(g1382_n_spl_),
    .din2(g1451_p_spl_)
  );


  FA
  g_g1452_n
  (
    .dout(g1452_n),
    .din1(g1382_p_spl_),
    .din2(g1451_n_spl_)
  );


  LA
  g_g1453_p
  (
    .dout(g1453_p),
    .din1(g1382_p_spl_),
    .din2(g1451_n_spl_)
  );


  FA
  g_g1453_n
  (
    .dout(g1453_n),
    .din1(g1382_n_spl_),
    .din2(g1451_p_spl_)
  );


  LA
  g_g1454_p
  (
    .dout(g1454_p),
    .din1(g1452_n_spl_),
    .din2(g1453_n)
  );


  FA
  g_g1454_n
  (
    .dout(g1454_n),
    .din1(g1452_p_spl_),
    .din2(g1453_p)
  );


  LA
  g_g1455_p
  (
    .dout(g1455_p),
    .din1(g1381_n_spl_),
    .din2(g1454_p_spl_)
  );


  FA
  g_g1455_n
  (
    .dout(g1455_n),
    .din1(g1381_p_spl_),
    .din2(g1454_n_spl_)
  );


  LA
  g_g1456_p
  (
    .dout(g1456_p),
    .din1(g1381_p_spl_),
    .din2(g1454_n_spl_)
  );


  FA
  g_g1456_n
  (
    .dout(g1456_n),
    .din1(g1381_n_spl_),
    .din2(g1454_p_spl_)
  );


  LA
  g_g1457_p
  (
    .dout(g1457_p),
    .din1(g1455_n_spl_),
    .din2(g1456_n)
  );


  FA
  g_g1457_n
  (
    .dout(g1457_n),
    .din1(g1455_p_spl_),
    .din2(g1456_p)
  );


  LA
  g_g1458_p
  (
    .dout(g1458_p),
    .din1(g1380_n_spl_),
    .din2(g1457_p_spl_)
  );


  FA
  g_g1458_n
  (
    .dout(g1458_n),
    .din1(g1380_p_spl_),
    .din2(g1457_n_spl_)
  );


  LA
  g_g1459_p
  (
    .dout(g1459_p),
    .din1(g1380_p_spl_),
    .din2(g1457_n_spl_)
  );


  FA
  g_g1459_n
  (
    .dout(g1459_n),
    .din1(g1380_n_spl_),
    .din2(g1457_p_spl_)
  );


  LA
  g_g1460_p
  (
    .dout(g1460_p),
    .din1(g1458_n_spl_),
    .din2(g1459_n)
  );


  FA
  g_g1460_n
  (
    .dout(g1460_n),
    .din1(g1458_p_spl_),
    .din2(g1459_p)
  );


  LA
  g_g1461_p
  (
    .dout(g1461_p),
    .din1(g1379_n_spl_),
    .din2(g1460_p_spl_)
  );


  FA
  g_g1461_n
  (
    .dout(g1461_n),
    .din1(g1379_p_spl_),
    .din2(g1460_n_spl_)
  );


  LA
  g_g1462_p
  (
    .dout(g1462_p),
    .din1(g1379_p_spl_),
    .din2(g1460_n_spl_)
  );


  FA
  g_g1462_n
  (
    .dout(g1462_n),
    .din1(g1379_n_spl_),
    .din2(g1460_p_spl_)
  );


  LA
  g_g1463_p
  (
    .dout(g1463_p),
    .din1(g1461_n_spl_),
    .din2(g1462_n)
  );


  FA
  g_g1463_n
  (
    .dout(g1463_n),
    .din1(g1461_p_spl_),
    .din2(g1462_p)
  );


  LA
  g_g1464_p
  (
    .dout(g1464_p),
    .din1(g1378_n),
    .din2(g1463_p)
  );


  FA
  g_g1464_n
  (
    .dout(g1464_n),
    .din1(g1378_p_spl_),
    .din2(g1463_n_spl_)
  );


  LA
  g_g1465_p
  (
    .dout(g1465_p),
    .din1(g1378_p_spl_),
    .din2(g1463_n_spl_)
  );


  FA
  g_g1466_n
  (
    .dout(g1466_n),
    .din1(g1464_p_spl_),
    .din2(g1465_p)
  );


  LA
  g_g1467_p
  (
    .dout(g1467_p),
    .din1(g1461_n_spl_),
    .din2(g1464_n)
  );


  FA
  g_g1467_n
  (
    .dout(g1467_n),
    .din1(g1461_p_spl_),
    .din2(g1464_p_spl_)
  );


  LA
  g_g1468_p
  (
    .dout(g1468_p),
    .din1(g1455_n_spl_),
    .din2(g1458_n_spl_)
  );


  FA
  g_g1468_n
  (
    .dout(g1468_n),
    .din1(g1455_p_spl_),
    .din2(g1458_p_spl_)
  );


  LA
  g_g1469_p
  (
    .dout(g1469_p),
    .din1(G7_p_spl_111),
    .din2(G32_p_spl_011)
  );


  FA
  g_g1469_n
  (
    .dout(g1469_n),
    .din1(G7_n_spl_111),
    .din2(G32_n_spl_011)
  );


  LA
  g_g1470_p
  (
    .dout(g1470_p),
    .din1(g1449_n_spl_),
    .din2(g1452_n_spl_)
  );


  FA
  g_g1470_n
  (
    .dout(g1470_n),
    .din1(g1449_p_spl_),
    .din2(g1452_p_spl_)
  );


  LA
  g_g1471_p
  (
    .dout(g1471_p),
    .din1(G8_p_spl_111),
    .din2(G31_p_spl_011)
  );


  FA
  g_g1471_n
  (
    .dout(g1471_n),
    .din1(G8_n_spl_111),
    .din2(G31_n_spl_011)
  );


  LA
  g_g1472_p
  (
    .dout(g1472_p),
    .din1(g1443_n_spl_),
    .din2(g1446_n_spl_)
  );


  FA
  g_g1472_n
  (
    .dout(g1472_n),
    .din1(g1443_p_spl_),
    .din2(g1446_p_spl_)
  );


  LA
  g_g1473_p
  (
    .dout(g1473_p),
    .din1(G9_p_spl_110),
    .din2(G30_p_spl_100)
  );


  FA
  g_g1473_n
  (
    .dout(g1473_n),
    .din1(G9_n_spl_110),
    .din2(G30_n_spl_100)
  );


  LA
  g_g1474_p
  (
    .dout(g1474_p),
    .din1(g1437_n_spl_),
    .din2(g1440_n_spl_)
  );


  FA
  g_g1474_n
  (
    .dout(g1474_n),
    .din1(g1437_p_spl_),
    .din2(g1440_p_spl_)
  );


  LA
  g_g1475_p
  (
    .dout(g1475_p),
    .din1(G10_p_spl_110),
    .din2(G29_p_spl_100)
  );


  FA
  g_g1475_n
  (
    .dout(g1475_n),
    .din1(G10_n_spl_110),
    .din2(G29_n_spl_100)
  );


  LA
  g_g1476_p
  (
    .dout(g1476_p),
    .din1(g1431_n_spl_),
    .din2(g1434_n_spl_)
  );


  FA
  g_g1476_n
  (
    .dout(g1476_n),
    .din1(g1431_p_spl_),
    .din2(g1434_p_spl_)
  );


  LA
  g_g1477_p
  (
    .dout(g1477_p),
    .din1(G11_p_spl_101),
    .din2(G28_p_spl_101)
  );


  FA
  g_g1477_n
  (
    .dout(g1477_n),
    .din1(G11_n_spl_101),
    .din2(G28_n_spl_101)
  );


  LA
  g_g1478_p
  (
    .dout(g1478_p),
    .din1(g1425_n_spl_),
    .din2(g1428_n_spl_)
  );


  FA
  g_g1478_n
  (
    .dout(g1478_n),
    .din1(g1425_p_spl_),
    .din2(g1428_p_spl_)
  );


  LA
  g_g1479_p
  (
    .dout(g1479_p),
    .din1(G12_p_spl_101),
    .din2(G27_p_spl_101)
  );


  FA
  g_g1479_n
  (
    .dout(g1479_n),
    .din1(G12_n_spl_101),
    .din2(G27_n_spl_101)
  );


  LA
  g_g1480_p
  (
    .dout(g1480_p),
    .din1(g1419_n_spl_),
    .din2(g1422_n_spl_)
  );


  FA
  g_g1480_n
  (
    .dout(g1480_n),
    .din1(g1419_p_spl_),
    .din2(g1422_p_spl_)
  );


  LA
  g_g1481_p
  (
    .dout(g1481_p),
    .din1(G13_p_spl_100),
    .din2(G26_p_spl_110)
  );


  FA
  g_g1481_n
  (
    .dout(g1481_n),
    .din1(G13_n_spl_100),
    .din2(G26_n_spl_110)
  );


  LA
  g_g1482_p
  (
    .dout(g1482_p),
    .din1(g1413_n_spl_),
    .din2(g1416_n_spl_)
  );


  FA
  g_g1482_n
  (
    .dout(g1482_n),
    .din1(g1413_p_spl_),
    .din2(g1416_p_spl_)
  );


  LA
  g_g1483_p
  (
    .dout(g1483_p),
    .din1(G14_p_spl_100),
    .din2(G25_p_spl_110)
  );


  FA
  g_g1483_n
  (
    .dout(g1483_n),
    .din1(G14_n_spl_100),
    .din2(G25_n_spl_110)
  );


  LA
  g_g1484_p
  (
    .dout(g1484_p),
    .din1(g1407_n_spl_),
    .din2(g1410_n_spl_)
  );


  FA
  g_g1484_n
  (
    .dout(g1484_n),
    .din1(g1407_p_spl_),
    .din2(g1410_p_spl_)
  );


  LA
  g_g1485_p
  (
    .dout(g1485_p),
    .din1(G15_p_spl_011),
    .din2(G24_p_spl_111)
  );


  FA
  g_g1485_n
  (
    .dout(g1485_n),
    .din1(G15_n_spl_011),
    .din2(G24_n_spl_111)
  );


  LA
  g_g1486_p
  (
    .dout(g1486_p),
    .din1(G16_p_spl_011),
    .din2(G23_p_spl_111)
  );


  FA
  g_g1486_n
  (
    .dout(g1486_n),
    .din1(G16_n_spl_011),
    .din2(G23_n_spl_111)
  );


  LA
  g_g1487_p
  (
    .dout(g1487_p),
    .din1(g1401_n_spl_),
    .din2(g1404_n_spl_)
  );


  FA
  g_g1487_n
  (
    .dout(g1487_n),
    .din1(g1401_p_spl_),
    .din2(g1404_p_spl_)
  );


  LA
  g_g1488_p
  (
    .dout(g1488_p),
    .din1(g1486_n_spl_),
    .din2(g1487_n_spl_)
  );


  FA
  g_g1488_n
  (
    .dout(g1488_n),
    .din1(g1486_p_spl_),
    .din2(g1487_p_spl_)
  );


  LA
  g_g1489_p
  (
    .dout(g1489_p),
    .din1(g1486_p_spl_),
    .din2(g1487_p_spl_)
  );


  FA
  g_g1489_n
  (
    .dout(g1489_n),
    .din1(g1486_n_spl_),
    .din2(g1487_n_spl_)
  );


  LA
  g_g1490_p
  (
    .dout(g1490_p),
    .din1(g1488_n_spl_),
    .din2(g1489_n)
  );


  FA
  g_g1490_n
  (
    .dout(g1490_n),
    .din1(g1488_p_spl_),
    .din2(g1489_p)
  );


  LA
  g_g1491_p
  (
    .dout(g1491_p),
    .din1(g1485_n_spl_),
    .din2(g1490_p_spl_)
  );


  FA
  g_g1491_n
  (
    .dout(g1491_n),
    .din1(g1485_p_spl_),
    .din2(g1490_n_spl_)
  );


  LA
  g_g1492_p
  (
    .dout(g1492_p),
    .din1(g1485_p_spl_),
    .din2(g1490_n_spl_)
  );


  FA
  g_g1492_n
  (
    .dout(g1492_n),
    .din1(g1485_n_spl_),
    .din2(g1490_p_spl_)
  );


  LA
  g_g1493_p
  (
    .dout(g1493_p),
    .din1(g1491_n_spl_),
    .din2(g1492_n)
  );


  FA
  g_g1493_n
  (
    .dout(g1493_n),
    .din1(g1491_p_spl_),
    .din2(g1492_p)
  );


  LA
  g_g1494_p
  (
    .dout(g1494_p),
    .din1(g1484_n_spl_),
    .din2(g1493_p_spl_)
  );


  FA
  g_g1494_n
  (
    .dout(g1494_n),
    .din1(g1484_p_spl_),
    .din2(g1493_n_spl_)
  );


  LA
  g_g1495_p
  (
    .dout(g1495_p),
    .din1(g1484_p_spl_),
    .din2(g1493_n_spl_)
  );


  FA
  g_g1495_n
  (
    .dout(g1495_n),
    .din1(g1484_n_spl_),
    .din2(g1493_p_spl_)
  );


  LA
  g_g1496_p
  (
    .dout(g1496_p),
    .din1(g1494_n_spl_),
    .din2(g1495_n)
  );


  FA
  g_g1496_n
  (
    .dout(g1496_n),
    .din1(g1494_p_spl_),
    .din2(g1495_p)
  );


  LA
  g_g1497_p
  (
    .dout(g1497_p),
    .din1(g1483_n_spl_),
    .din2(g1496_p_spl_)
  );


  FA
  g_g1497_n
  (
    .dout(g1497_n),
    .din1(g1483_p_spl_),
    .din2(g1496_n_spl_)
  );


  LA
  g_g1498_p
  (
    .dout(g1498_p),
    .din1(g1483_p_spl_),
    .din2(g1496_n_spl_)
  );


  FA
  g_g1498_n
  (
    .dout(g1498_n),
    .din1(g1483_n_spl_),
    .din2(g1496_p_spl_)
  );


  LA
  g_g1499_p
  (
    .dout(g1499_p),
    .din1(g1497_n_spl_),
    .din2(g1498_n)
  );


  FA
  g_g1499_n
  (
    .dout(g1499_n),
    .din1(g1497_p_spl_),
    .din2(g1498_p)
  );


  LA
  g_g1500_p
  (
    .dout(g1500_p),
    .din1(g1482_n_spl_),
    .din2(g1499_p_spl_)
  );


  FA
  g_g1500_n
  (
    .dout(g1500_n),
    .din1(g1482_p_spl_),
    .din2(g1499_n_spl_)
  );


  LA
  g_g1501_p
  (
    .dout(g1501_p),
    .din1(g1482_p_spl_),
    .din2(g1499_n_spl_)
  );


  FA
  g_g1501_n
  (
    .dout(g1501_n),
    .din1(g1482_n_spl_),
    .din2(g1499_p_spl_)
  );


  LA
  g_g1502_p
  (
    .dout(g1502_p),
    .din1(g1500_n_spl_),
    .din2(g1501_n)
  );


  FA
  g_g1502_n
  (
    .dout(g1502_n),
    .din1(g1500_p_spl_),
    .din2(g1501_p)
  );


  LA
  g_g1503_p
  (
    .dout(g1503_p),
    .din1(g1481_n_spl_),
    .din2(g1502_p_spl_)
  );


  FA
  g_g1503_n
  (
    .dout(g1503_n),
    .din1(g1481_p_spl_),
    .din2(g1502_n_spl_)
  );


  LA
  g_g1504_p
  (
    .dout(g1504_p),
    .din1(g1481_p_spl_),
    .din2(g1502_n_spl_)
  );


  FA
  g_g1504_n
  (
    .dout(g1504_n),
    .din1(g1481_n_spl_),
    .din2(g1502_p_spl_)
  );


  LA
  g_g1505_p
  (
    .dout(g1505_p),
    .din1(g1503_n_spl_),
    .din2(g1504_n)
  );


  FA
  g_g1505_n
  (
    .dout(g1505_n),
    .din1(g1503_p_spl_),
    .din2(g1504_p)
  );


  LA
  g_g1506_p
  (
    .dout(g1506_p),
    .din1(g1480_n_spl_),
    .din2(g1505_p_spl_)
  );


  FA
  g_g1506_n
  (
    .dout(g1506_n),
    .din1(g1480_p_spl_),
    .din2(g1505_n_spl_)
  );


  LA
  g_g1507_p
  (
    .dout(g1507_p),
    .din1(g1480_p_spl_),
    .din2(g1505_n_spl_)
  );


  FA
  g_g1507_n
  (
    .dout(g1507_n),
    .din1(g1480_n_spl_),
    .din2(g1505_p_spl_)
  );


  LA
  g_g1508_p
  (
    .dout(g1508_p),
    .din1(g1506_n_spl_),
    .din2(g1507_n)
  );


  FA
  g_g1508_n
  (
    .dout(g1508_n),
    .din1(g1506_p_spl_),
    .din2(g1507_p)
  );


  LA
  g_g1509_p
  (
    .dout(g1509_p),
    .din1(g1479_n_spl_),
    .din2(g1508_p_spl_)
  );


  FA
  g_g1509_n
  (
    .dout(g1509_n),
    .din1(g1479_p_spl_),
    .din2(g1508_n_spl_)
  );


  LA
  g_g1510_p
  (
    .dout(g1510_p),
    .din1(g1479_p_spl_),
    .din2(g1508_n_spl_)
  );


  FA
  g_g1510_n
  (
    .dout(g1510_n),
    .din1(g1479_n_spl_),
    .din2(g1508_p_spl_)
  );


  LA
  g_g1511_p
  (
    .dout(g1511_p),
    .din1(g1509_n_spl_),
    .din2(g1510_n)
  );


  FA
  g_g1511_n
  (
    .dout(g1511_n),
    .din1(g1509_p_spl_),
    .din2(g1510_p)
  );


  LA
  g_g1512_p
  (
    .dout(g1512_p),
    .din1(g1478_n_spl_),
    .din2(g1511_p_spl_)
  );


  FA
  g_g1512_n
  (
    .dout(g1512_n),
    .din1(g1478_p_spl_),
    .din2(g1511_n_spl_)
  );


  LA
  g_g1513_p
  (
    .dout(g1513_p),
    .din1(g1478_p_spl_),
    .din2(g1511_n_spl_)
  );


  FA
  g_g1513_n
  (
    .dout(g1513_n),
    .din1(g1478_n_spl_),
    .din2(g1511_p_spl_)
  );


  LA
  g_g1514_p
  (
    .dout(g1514_p),
    .din1(g1512_n_spl_),
    .din2(g1513_n)
  );


  FA
  g_g1514_n
  (
    .dout(g1514_n),
    .din1(g1512_p_spl_),
    .din2(g1513_p)
  );


  LA
  g_g1515_p
  (
    .dout(g1515_p),
    .din1(g1477_n_spl_),
    .din2(g1514_p_spl_)
  );


  FA
  g_g1515_n
  (
    .dout(g1515_n),
    .din1(g1477_p_spl_),
    .din2(g1514_n_spl_)
  );


  LA
  g_g1516_p
  (
    .dout(g1516_p),
    .din1(g1477_p_spl_),
    .din2(g1514_n_spl_)
  );


  FA
  g_g1516_n
  (
    .dout(g1516_n),
    .din1(g1477_n_spl_),
    .din2(g1514_p_spl_)
  );


  LA
  g_g1517_p
  (
    .dout(g1517_p),
    .din1(g1515_n_spl_),
    .din2(g1516_n)
  );


  FA
  g_g1517_n
  (
    .dout(g1517_n),
    .din1(g1515_p_spl_),
    .din2(g1516_p)
  );


  LA
  g_g1518_p
  (
    .dout(g1518_p),
    .din1(g1476_n_spl_),
    .din2(g1517_p_spl_)
  );


  FA
  g_g1518_n
  (
    .dout(g1518_n),
    .din1(g1476_p_spl_),
    .din2(g1517_n_spl_)
  );


  LA
  g_g1519_p
  (
    .dout(g1519_p),
    .din1(g1476_p_spl_),
    .din2(g1517_n_spl_)
  );


  FA
  g_g1519_n
  (
    .dout(g1519_n),
    .din1(g1476_n_spl_),
    .din2(g1517_p_spl_)
  );


  LA
  g_g1520_p
  (
    .dout(g1520_p),
    .din1(g1518_n_spl_),
    .din2(g1519_n)
  );


  FA
  g_g1520_n
  (
    .dout(g1520_n),
    .din1(g1518_p_spl_),
    .din2(g1519_p)
  );


  LA
  g_g1521_p
  (
    .dout(g1521_p),
    .din1(g1475_n_spl_),
    .din2(g1520_p_spl_)
  );


  FA
  g_g1521_n
  (
    .dout(g1521_n),
    .din1(g1475_p_spl_),
    .din2(g1520_n_spl_)
  );


  LA
  g_g1522_p
  (
    .dout(g1522_p),
    .din1(g1475_p_spl_),
    .din2(g1520_n_spl_)
  );


  FA
  g_g1522_n
  (
    .dout(g1522_n),
    .din1(g1475_n_spl_),
    .din2(g1520_p_spl_)
  );


  LA
  g_g1523_p
  (
    .dout(g1523_p),
    .din1(g1521_n_spl_),
    .din2(g1522_n)
  );


  FA
  g_g1523_n
  (
    .dout(g1523_n),
    .din1(g1521_p_spl_),
    .din2(g1522_p)
  );


  LA
  g_g1524_p
  (
    .dout(g1524_p),
    .din1(g1474_n_spl_),
    .din2(g1523_p_spl_)
  );


  FA
  g_g1524_n
  (
    .dout(g1524_n),
    .din1(g1474_p_spl_),
    .din2(g1523_n_spl_)
  );


  LA
  g_g1525_p
  (
    .dout(g1525_p),
    .din1(g1474_p_spl_),
    .din2(g1523_n_spl_)
  );


  FA
  g_g1525_n
  (
    .dout(g1525_n),
    .din1(g1474_n_spl_),
    .din2(g1523_p_spl_)
  );


  LA
  g_g1526_p
  (
    .dout(g1526_p),
    .din1(g1524_n_spl_),
    .din2(g1525_n)
  );


  FA
  g_g1526_n
  (
    .dout(g1526_n),
    .din1(g1524_p_spl_),
    .din2(g1525_p)
  );


  LA
  g_g1527_p
  (
    .dout(g1527_p),
    .din1(g1473_n_spl_),
    .din2(g1526_p_spl_)
  );


  FA
  g_g1527_n
  (
    .dout(g1527_n),
    .din1(g1473_p_spl_),
    .din2(g1526_n_spl_)
  );


  LA
  g_g1528_p
  (
    .dout(g1528_p),
    .din1(g1473_p_spl_),
    .din2(g1526_n_spl_)
  );


  FA
  g_g1528_n
  (
    .dout(g1528_n),
    .din1(g1473_n_spl_),
    .din2(g1526_p_spl_)
  );


  LA
  g_g1529_p
  (
    .dout(g1529_p),
    .din1(g1527_n_spl_),
    .din2(g1528_n)
  );


  FA
  g_g1529_n
  (
    .dout(g1529_n),
    .din1(g1527_p_spl_),
    .din2(g1528_p)
  );


  LA
  g_g1530_p
  (
    .dout(g1530_p),
    .din1(g1472_n_spl_),
    .din2(g1529_p_spl_)
  );


  FA
  g_g1530_n
  (
    .dout(g1530_n),
    .din1(g1472_p_spl_),
    .din2(g1529_n_spl_)
  );


  LA
  g_g1531_p
  (
    .dout(g1531_p),
    .din1(g1472_p_spl_),
    .din2(g1529_n_spl_)
  );


  FA
  g_g1531_n
  (
    .dout(g1531_n),
    .din1(g1472_n_spl_),
    .din2(g1529_p_spl_)
  );


  LA
  g_g1532_p
  (
    .dout(g1532_p),
    .din1(g1530_n_spl_),
    .din2(g1531_n)
  );


  FA
  g_g1532_n
  (
    .dout(g1532_n),
    .din1(g1530_p_spl_),
    .din2(g1531_p)
  );


  LA
  g_g1533_p
  (
    .dout(g1533_p),
    .din1(g1471_n_spl_),
    .din2(g1532_p_spl_)
  );


  FA
  g_g1533_n
  (
    .dout(g1533_n),
    .din1(g1471_p_spl_),
    .din2(g1532_n_spl_)
  );


  LA
  g_g1534_p
  (
    .dout(g1534_p),
    .din1(g1471_p_spl_),
    .din2(g1532_n_spl_)
  );


  FA
  g_g1534_n
  (
    .dout(g1534_n),
    .din1(g1471_n_spl_),
    .din2(g1532_p_spl_)
  );


  LA
  g_g1535_p
  (
    .dout(g1535_p),
    .din1(g1533_n_spl_),
    .din2(g1534_n)
  );


  FA
  g_g1535_n
  (
    .dout(g1535_n),
    .din1(g1533_p_spl_),
    .din2(g1534_p)
  );


  LA
  g_g1536_p
  (
    .dout(g1536_p),
    .din1(g1470_n_spl_),
    .din2(g1535_p_spl_)
  );


  FA
  g_g1536_n
  (
    .dout(g1536_n),
    .din1(g1470_p_spl_),
    .din2(g1535_n_spl_)
  );


  LA
  g_g1537_p
  (
    .dout(g1537_p),
    .din1(g1470_p_spl_),
    .din2(g1535_n_spl_)
  );


  FA
  g_g1537_n
  (
    .dout(g1537_n),
    .din1(g1470_n_spl_),
    .din2(g1535_p_spl_)
  );


  LA
  g_g1538_p
  (
    .dout(g1538_p),
    .din1(g1536_n_spl_),
    .din2(g1537_n)
  );


  FA
  g_g1538_n
  (
    .dout(g1538_n),
    .din1(g1536_p_spl_),
    .din2(g1537_p)
  );


  LA
  g_g1539_p
  (
    .dout(g1539_p),
    .din1(g1469_n_spl_),
    .din2(g1538_p_spl_)
  );


  FA
  g_g1539_n
  (
    .dout(g1539_n),
    .din1(g1469_p_spl_),
    .din2(g1538_n_spl_)
  );


  LA
  g_g1540_p
  (
    .dout(g1540_p),
    .din1(g1469_p_spl_),
    .din2(g1538_n_spl_)
  );


  FA
  g_g1540_n
  (
    .dout(g1540_n),
    .din1(g1469_n_spl_),
    .din2(g1538_p_spl_)
  );


  LA
  g_g1541_p
  (
    .dout(g1541_p),
    .din1(g1539_n_spl_),
    .din2(g1540_n)
  );


  FA
  g_g1541_n
  (
    .dout(g1541_n),
    .din1(g1539_p_spl_),
    .din2(g1540_p)
  );


  LA
  g_g1542_p
  (
    .dout(g1542_p),
    .din1(g1468_n_spl_),
    .din2(g1541_p_spl_)
  );


  FA
  g_g1542_n
  (
    .dout(g1542_n),
    .din1(g1468_p_spl_),
    .din2(g1541_n_spl_)
  );


  LA
  g_g1543_p
  (
    .dout(g1543_p),
    .din1(g1468_p_spl_),
    .din2(g1541_n_spl_)
  );


  FA
  g_g1543_n
  (
    .dout(g1543_n),
    .din1(g1468_n_spl_),
    .din2(g1541_p_spl_)
  );


  LA
  g_g1544_p
  (
    .dout(g1544_p),
    .din1(g1542_n_spl_),
    .din2(g1543_n)
  );


  FA
  g_g1544_n
  (
    .dout(g1544_n),
    .din1(g1542_p_spl_),
    .din2(g1543_p)
  );


  LA
  g_g1545_p
  (
    .dout(g1545_p),
    .din1(g1467_n),
    .din2(g1544_p)
  );


  FA
  g_g1545_n
  (
    .dout(g1545_n),
    .din1(g1467_p_spl_),
    .din2(g1544_n_spl_)
  );


  LA
  g_g1546_p
  (
    .dout(g1546_p),
    .din1(g1467_p_spl_),
    .din2(g1544_n_spl_)
  );


  FA
  g_g1547_n
  (
    .dout(g1547_n),
    .din1(g1545_p_spl_),
    .din2(g1546_p)
  );


  LA
  g_g1548_p
  (
    .dout(g1548_p),
    .din1(g1542_n_spl_),
    .din2(g1545_n)
  );


  FA
  g_g1548_n
  (
    .dout(g1548_n),
    .din1(g1542_p_spl_),
    .din2(g1545_p_spl_)
  );


  LA
  g_g1549_p
  (
    .dout(g1549_p),
    .din1(g1536_n_spl_),
    .din2(g1539_n_spl_)
  );


  FA
  g_g1549_n
  (
    .dout(g1549_n),
    .din1(g1536_p_spl_),
    .din2(g1539_p_spl_)
  );


  LA
  g_g1550_p
  (
    .dout(g1550_p),
    .din1(G8_p_spl_111),
    .din2(G32_p_spl_011)
  );


  FA
  g_g1550_n
  (
    .dout(g1550_n),
    .din1(G8_n_spl_111),
    .din2(G32_n_spl_011)
  );


  LA
  g_g1551_p
  (
    .dout(g1551_p),
    .din1(g1530_n_spl_),
    .din2(g1533_n_spl_)
  );


  FA
  g_g1551_n
  (
    .dout(g1551_n),
    .din1(g1530_p_spl_),
    .din2(g1533_p_spl_)
  );


  LA
  g_g1552_p
  (
    .dout(g1552_p),
    .din1(G9_p_spl_111),
    .din2(G31_p_spl_100)
  );


  FA
  g_g1552_n
  (
    .dout(g1552_n),
    .din1(G9_n_spl_111),
    .din2(G31_n_spl_100)
  );


  LA
  g_g1553_p
  (
    .dout(g1553_p),
    .din1(g1524_n_spl_),
    .din2(g1527_n_spl_)
  );


  FA
  g_g1553_n
  (
    .dout(g1553_n),
    .din1(g1524_p_spl_),
    .din2(g1527_p_spl_)
  );


  LA
  g_g1554_p
  (
    .dout(g1554_p),
    .din1(G10_p_spl_110),
    .din2(G30_p_spl_100)
  );


  FA
  g_g1554_n
  (
    .dout(g1554_n),
    .din1(G10_n_spl_110),
    .din2(G30_n_spl_100)
  );


  LA
  g_g1555_p
  (
    .dout(g1555_p),
    .din1(g1518_n_spl_),
    .din2(g1521_n_spl_)
  );


  FA
  g_g1555_n
  (
    .dout(g1555_n),
    .din1(g1518_p_spl_),
    .din2(g1521_p_spl_)
  );


  LA
  g_g1556_p
  (
    .dout(g1556_p),
    .din1(G11_p_spl_110),
    .din2(G29_p_spl_101)
  );


  FA
  g_g1556_n
  (
    .dout(g1556_n),
    .din1(G11_n_spl_110),
    .din2(G29_n_spl_101)
  );


  LA
  g_g1557_p
  (
    .dout(g1557_p),
    .din1(g1512_n_spl_),
    .din2(g1515_n_spl_)
  );


  FA
  g_g1557_n
  (
    .dout(g1557_n),
    .din1(g1512_p_spl_),
    .din2(g1515_p_spl_)
  );


  LA
  g_g1558_p
  (
    .dout(g1558_p),
    .din1(G12_p_spl_101),
    .din2(G28_p_spl_101)
  );


  FA
  g_g1558_n
  (
    .dout(g1558_n),
    .din1(G12_n_spl_101),
    .din2(G28_n_spl_101)
  );


  LA
  g_g1559_p
  (
    .dout(g1559_p),
    .din1(g1506_n_spl_),
    .din2(g1509_n_spl_)
  );


  FA
  g_g1559_n
  (
    .dout(g1559_n),
    .din1(g1506_p_spl_),
    .din2(g1509_p_spl_)
  );


  LA
  g_g1560_p
  (
    .dout(g1560_p),
    .din1(G13_p_spl_101),
    .din2(G27_p_spl_110)
  );


  FA
  g_g1560_n
  (
    .dout(g1560_n),
    .din1(G13_n_spl_101),
    .din2(G27_n_spl_110)
  );


  LA
  g_g1561_p
  (
    .dout(g1561_p),
    .din1(g1500_n_spl_),
    .din2(g1503_n_spl_)
  );


  FA
  g_g1561_n
  (
    .dout(g1561_n),
    .din1(g1500_p_spl_),
    .din2(g1503_p_spl_)
  );


  LA
  g_g1562_p
  (
    .dout(g1562_p),
    .din1(G14_p_spl_100),
    .din2(G26_p_spl_110)
  );


  FA
  g_g1562_n
  (
    .dout(g1562_n),
    .din1(G14_n_spl_100),
    .din2(G26_n_spl_110)
  );


  LA
  g_g1563_p
  (
    .dout(g1563_p),
    .din1(g1494_n_spl_),
    .din2(g1497_n_spl_)
  );


  FA
  g_g1563_n
  (
    .dout(g1563_n),
    .din1(g1494_p_spl_),
    .din2(g1497_p_spl_)
  );


  LA
  g_g1564_p
  (
    .dout(g1564_p),
    .din1(G15_p_spl_100),
    .din2(G25_p_spl_111)
  );


  FA
  g_g1564_n
  (
    .dout(g1564_n),
    .din1(G15_n_spl_100),
    .din2(G25_n_spl_111)
  );


  LA
  g_g1565_p
  (
    .dout(g1565_p),
    .din1(G16_p_spl_011),
    .din2(G24_p_spl_111)
  );


  FA
  g_g1565_n
  (
    .dout(g1565_n),
    .din1(G16_n_spl_011),
    .din2(G24_n_spl_111)
  );


  LA
  g_g1566_p
  (
    .dout(g1566_p),
    .din1(g1488_n_spl_),
    .din2(g1491_n_spl_)
  );


  FA
  g_g1566_n
  (
    .dout(g1566_n),
    .din1(g1488_p_spl_),
    .din2(g1491_p_spl_)
  );


  LA
  g_g1567_p
  (
    .dout(g1567_p),
    .din1(g1565_n_spl_),
    .din2(g1566_n_spl_)
  );


  FA
  g_g1567_n
  (
    .dout(g1567_n),
    .din1(g1565_p_spl_),
    .din2(g1566_p_spl_)
  );


  LA
  g_g1568_p
  (
    .dout(g1568_p),
    .din1(g1565_p_spl_),
    .din2(g1566_p_spl_)
  );


  FA
  g_g1568_n
  (
    .dout(g1568_n),
    .din1(g1565_n_spl_),
    .din2(g1566_n_spl_)
  );


  LA
  g_g1569_p
  (
    .dout(g1569_p),
    .din1(g1567_n_spl_),
    .din2(g1568_n)
  );


  FA
  g_g1569_n
  (
    .dout(g1569_n),
    .din1(g1567_p_spl_),
    .din2(g1568_p)
  );


  LA
  g_g1570_p
  (
    .dout(g1570_p),
    .din1(g1564_n_spl_),
    .din2(g1569_p_spl_)
  );


  FA
  g_g1570_n
  (
    .dout(g1570_n),
    .din1(g1564_p_spl_),
    .din2(g1569_n_spl_)
  );


  LA
  g_g1571_p
  (
    .dout(g1571_p),
    .din1(g1564_p_spl_),
    .din2(g1569_n_spl_)
  );


  FA
  g_g1571_n
  (
    .dout(g1571_n),
    .din1(g1564_n_spl_),
    .din2(g1569_p_spl_)
  );


  LA
  g_g1572_p
  (
    .dout(g1572_p),
    .din1(g1570_n_spl_),
    .din2(g1571_n)
  );


  FA
  g_g1572_n
  (
    .dout(g1572_n),
    .din1(g1570_p_spl_),
    .din2(g1571_p)
  );


  LA
  g_g1573_p
  (
    .dout(g1573_p),
    .din1(g1563_n_spl_),
    .din2(g1572_p_spl_)
  );


  FA
  g_g1573_n
  (
    .dout(g1573_n),
    .din1(g1563_p_spl_),
    .din2(g1572_n_spl_)
  );


  LA
  g_g1574_p
  (
    .dout(g1574_p),
    .din1(g1563_p_spl_),
    .din2(g1572_n_spl_)
  );


  FA
  g_g1574_n
  (
    .dout(g1574_n),
    .din1(g1563_n_spl_),
    .din2(g1572_p_spl_)
  );


  LA
  g_g1575_p
  (
    .dout(g1575_p),
    .din1(g1573_n_spl_),
    .din2(g1574_n)
  );


  FA
  g_g1575_n
  (
    .dout(g1575_n),
    .din1(g1573_p_spl_),
    .din2(g1574_p)
  );


  LA
  g_g1576_p
  (
    .dout(g1576_p),
    .din1(g1562_n_spl_),
    .din2(g1575_p_spl_)
  );


  FA
  g_g1576_n
  (
    .dout(g1576_n),
    .din1(g1562_p_spl_),
    .din2(g1575_n_spl_)
  );


  LA
  g_g1577_p
  (
    .dout(g1577_p),
    .din1(g1562_p_spl_),
    .din2(g1575_n_spl_)
  );


  FA
  g_g1577_n
  (
    .dout(g1577_n),
    .din1(g1562_n_spl_),
    .din2(g1575_p_spl_)
  );


  LA
  g_g1578_p
  (
    .dout(g1578_p),
    .din1(g1576_n_spl_),
    .din2(g1577_n)
  );


  FA
  g_g1578_n
  (
    .dout(g1578_n),
    .din1(g1576_p_spl_),
    .din2(g1577_p)
  );


  LA
  g_g1579_p
  (
    .dout(g1579_p),
    .din1(g1561_n_spl_),
    .din2(g1578_p_spl_)
  );


  FA
  g_g1579_n
  (
    .dout(g1579_n),
    .din1(g1561_p_spl_),
    .din2(g1578_n_spl_)
  );


  LA
  g_g1580_p
  (
    .dout(g1580_p),
    .din1(g1561_p_spl_),
    .din2(g1578_n_spl_)
  );


  FA
  g_g1580_n
  (
    .dout(g1580_n),
    .din1(g1561_n_spl_),
    .din2(g1578_p_spl_)
  );


  LA
  g_g1581_p
  (
    .dout(g1581_p),
    .din1(g1579_n_spl_),
    .din2(g1580_n)
  );


  FA
  g_g1581_n
  (
    .dout(g1581_n),
    .din1(g1579_p_spl_),
    .din2(g1580_p)
  );


  LA
  g_g1582_p
  (
    .dout(g1582_p),
    .din1(g1560_n_spl_),
    .din2(g1581_p_spl_)
  );


  FA
  g_g1582_n
  (
    .dout(g1582_n),
    .din1(g1560_p_spl_),
    .din2(g1581_n_spl_)
  );


  LA
  g_g1583_p
  (
    .dout(g1583_p),
    .din1(g1560_p_spl_),
    .din2(g1581_n_spl_)
  );


  FA
  g_g1583_n
  (
    .dout(g1583_n),
    .din1(g1560_n_spl_),
    .din2(g1581_p_spl_)
  );


  LA
  g_g1584_p
  (
    .dout(g1584_p),
    .din1(g1582_n_spl_),
    .din2(g1583_n)
  );


  FA
  g_g1584_n
  (
    .dout(g1584_n),
    .din1(g1582_p_spl_),
    .din2(g1583_p)
  );


  LA
  g_g1585_p
  (
    .dout(g1585_p),
    .din1(g1559_n_spl_),
    .din2(g1584_p_spl_)
  );


  FA
  g_g1585_n
  (
    .dout(g1585_n),
    .din1(g1559_p_spl_),
    .din2(g1584_n_spl_)
  );


  LA
  g_g1586_p
  (
    .dout(g1586_p),
    .din1(g1559_p_spl_),
    .din2(g1584_n_spl_)
  );


  FA
  g_g1586_n
  (
    .dout(g1586_n),
    .din1(g1559_n_spl_),
    .din2(g1584_p_spl_)
  );


  LA
  g_g1587_p
  (
    .dout(g1587_p),
    .din1(g1585_n_spl_),
    .din2(g1586_n)
  );


  FA
  g_g1587_n
  (
    .dout(g1587_n),
    .din1(g1585_p_spl_),
    .din2(g1586_p)
  );


  LA
  g_g1588_p
  (
    .dout(g1588_p),
    .din1(g1558_n_spl_),
    .din2(g1587_p_spl_)
  );


  FA
  g_g1588_n
  (
    .dout(g1588_n),
    .din1(g1558_p_spl_),
    .din2(g1587_n_spl_)
  );


  LA
  g_g1589_p
  (
    .dout(g1589_p),
    .din1(g1558_p_spl_),
    .din2(g1587_n_spl_)
  );


  FA
  g_g1589_n
  (
    .dout(g1589_n),
    .din1(g1558_n_spl_),
    .din2(g1587_p_spl_)
  );


  LA
  g_g1590_p
  (
    .dout(g1590_p),
    .din1(g1588_n_spl_),
    .din2(g1589_n)
  );


  FA
  g_g1590_n
  (
    .dout(g1590_n),
    .din1(g1588_p_spl_),
    .din2(g1589_p)
  );


  LA
  g_g1591_p
  (
    .dout(g1591_p),
    .din1(g1557_n_spl_),
    .din2(g1590_p_spl_)
  );


  FA
  g_g1591_n
  (
    .dout(g1591_n),
    .din1(g1557_p_spl_),
    .din2(g1590_n_spl_)
  );


  LA
  g_g1592_p
  (
    .dout(g1592_p),
    .din1(g1557_p_spl_),
    .din2(g1590_n_spl_)
  );


  FA
  g_g1592_n
  (
    .dout(g1592_n),
    .din1(g1557_n_spl_),
    .din2(g1590_p_spl_)
  );


  LA
  g_g1593_p
  (
    .dout(g1593_p),
    .din1(g1591_n_spl_),
    .din2(g1592_n)
  );


  FA
  g_g1593_n
  (
    .dout(g1593_n),
    .din1(g1591_p_spl_),
    .din2(g1592_p)
  );


  LA
  g_g1594_p
  (
    .dout(g1594_p),
    .din1(g1556_n_spl_),
    .din2(g1593_p_spl_)
  );


  FA
  g_g1594_n
  (
    .dout(g1594_n),
    .din1(g1556_p_spl_),
    .din2(g1593_n_spl_)
  );


  LA
  g_g1595_p
  (
    .dout(g1595_p),
    .din1(g1556_p_spl_),
    .din2(g1593_n_spl_)
  );


  FA
  g_g1595_n
  (
    .dout(g1595_n),
    .din1(g1556_n_spl_),
    .din2(g1593_p_spl_)
  );


  LA
  g_g1596_p
  (
    .dout(g1596_p),
    .din1(g1594_n_spl_),
    .din2(g1595_n)
  );


  FA
  g_g1596_n
  (
    .dout(g1596_n),
    .din1(g1594_p_spl_),
    .din2(g1595_p)
  );


  LA
  g_g1597_p
  (
    .dout(g1597_p),
    .din1(g1555_n_spl_),
    .din2(g1596_p_spl_)
  );


  FA
  g_g1597_n
  (
    .dout(g1597_n),
    .din1(g1555_p_spl_),
    .din2(g1596_n_spl_)
  );


  LA
  g_g1598_p
  (
    .dout(g1598_p),
    .din1(g1555_p_spl_),
    .din2(g1596_n_spl_)
  );


  FA
  g_g1598_n
  (
    .dout(g1598_n),
    .din1(g1555_n_spl_),
    .din2(g1596_p_spl_)
  );


  LA
  g_g1599_p
  (
    .dout(g1599_p),
    .din1(g1597_n_spl_),
    .din2(g1598_n)
  );


  FA
  g_g1599_n
  (
    .dout(g1599_n),
    .din1(g1597_p_spl_),
    .din2(g1598_p)
  );


  LA
  g_g1600_p
  (
    .dout(g1600_p),
    .din1(g1554_n_spl_),
    .din2(g1599_p_spl_)
  );


  FA
  g_g1600_n
  (
    .dout(g1600_n),
    .din1(g1554_p_spl_),
    .din2(g1599_n_spl_)
  );


  LA
  g_g1601_p
  (
    .dout(g1601_p),
    .din1(g1554_p_spl_),
    .din2(g1599_n_spl_)
  );


  FA
  g_g1601_n
  (
    .dout(g1601_n),
    .din1(g1554_n_spl_),
    .din2(g1599_p_spl_)
  );


  LA
  g_g1602_p
  (
    .dout(g1602_p),
    .din1(g1600_n_spl_),
    .din2(g1601_n)
  );


  FA
  g_g1602_n
  (
    .dout(g1602_n),
    .din1(g1600_p_spl_),
    .din2(g1601_p)
  );


  LA
  g_g1603_p
  (
    .dout(g1603_p),
    .din1(g1553_n_spl_),
    .din2(g1602_p_spl_)
  );


  FA
  g_g1603_n
  (
    .dout(g1603_n),
    .din1(g1553_p_spl_),
    .din2(g1602_n_spl_)
  );


  LA
  g_g1604_p
  (
    .dout(g1604_p),
    .din1(g1553_p_spl_),
    .din2(g1602_n_spl_)
  );


  FA
  g_g1604_n
  (
    .dout(g1604_n),
    .din1(g1553_n_spl_),
    .din2(g1602_p_spl_)
  );


  LA
  g_g1605_p
  (
    .dout(g1605_p),
    .din1(g1603_n_spl_),
    .din2(g1604_n)
  );


  FA
  g_g1605_n
  (
    .dout(g1605_n),
    .din1(g1603_p_spl_),
    .din2(g1604_p)
  );


  LA
  g_g1606_p
  (
    .dout(g1606_p),
    .din1(g1552_n_spl_),
    .din2(g1605_p_spl_)
  );


  FA
  g_g1606_n
  (
    .dout(g1606_n),
    .din1(g1552_p_spl_),
    .din2(g1605_n_spl_)
  );


  LA
  g_g1607_p
  (
    .dout(g1607_p),
    .din1(g1552_p_spl_),
    .din2(g1605_n_spl_)
  );


  FA
  g_g1607_n
  (
    .dout(g1607_n),
    .din1(g1552_n_spl_),
    .din2(g1605_p_spl_)
  );


  LA
  g_g1608_p
  (
    .dout(g1608_p),
    .din1(g1606_n_spl_),
    .din2(g1607_n)
  );


  FA
  g_g1608_n
  (
    .dout(g1608_n),
    .din1(g1606_p_spl_),
    .din2(g1607_p)
  );


  LA
  g_g1609_p
  (
    .dout(g1609_p),
    .din1(g1551_n_spl_),
    .din2(g1608_p_spl_)
  );


  FA
  g_g1609_n
  (
    .dout(g1609_n),
    .din1(g1551_p_spl_),
    .din2(g1608_n_spl_)
  );


  LA
  g_g1610_p
  (
    .dout(g1610_p),
    .din1(g1551_p_spl_),
    .din2(g1608_n_spl_)
  );


  FA
  g_g1610_n
  (
    .dout(g1610_n),
    .din1(g1551_n_spl_),
    .din2(g1608_p_spl_)
  );


  LA
  g_g1611_p
  (
    .dout(g1611_p),
    .din1(g1609_n_spl_),
    .din2(g1610_n)
  );


  FA
  g_g1611_n
  (
    .dout(g1611_n),
    .din1(g1609_p_spl_),
    .din2(g1610_p)
  );


  LA
  g_g1612_p
  (
    .dout(g1612_p),
    .din1(g1550_n_spl_),
    .din2(g1611_p_spl_)
  );


  FA
  g_g1612_n
  (
    .dout(g1612_n),
    .din1(g1550_p_spl_),
    .din2(g1611_n_spl_)
  );


  LA
  g_g1613_p
  (
    .dout(g1613_p),
    .din1(g1550_p_spl_),
    .din2(g1611_n_spl_)
  );


  FA
  g_g1613_n
  (
    .dout(g1613_n),
    .din1(g1550_n_spl_),
    .din2(g1611_p_spl_)
  );


  LA
  g_g1614_p
  (
    .dout(g1614_p),
    .din1(g1612_n_spl_),
    .din2(g1613_n)
  );


  FA
  g_g1614_n
  (
    .dout(g1614_n),
    .din1(g1612_p_spl_),
    .din2(g1613_p)
  );


  LA
  g_g1615_p
  (
    .dout(g1615_p),
    .din1(g1549_n_spl_),
    .din2(g1614_p_spl_)
  );


  FA
  g_g1615_n
  (
    .dout(g1615_n),
    .din1(g1549_p_spl_),
    .din2(g1614_n_spl_)
  );


  LA
  g_g1616_p
  (
    .dout(g1616_p),
    .din1(g1549_p_spl_),
    .din2(g1614_n_spl_)
  );


  FA
  g_g1616_n
  (
    .dout(g1616_n),
    .din1(g1549_n_spl_),
    .din2(g1614_p_spl_)
  );


  LA
  g_g1617_p
  (
    .dout(g1617_p),
    .din1(g1615_n_spl_),
    .din2(g1616_n)
  );


  FA
  g_g1617_n
  (
    .dout(g1617_n),
    .din1(g1615_p_spl_),
    .din2(g1616_p)
  );


  LA
  g_g1618_p
  (
    .dout(g1618_p),
    .din1(g1548_n),
    .din2(g1617_p)
  );


  FA
  g_g1618_n
  (
    .dout(g1618_n),
    .din1(g1548_p_spl_),
    .din2(g1617_n_spl_)
  );


  LA
  g_g1619_p
  (
    .dout(g1619_p),
    .din1(g1548_p_spl_),
    .din2(g1617_n_spl_)
  );


  FA
  g_g1620_n
  (
    .dout(g1620_n),
    .din1(g1618_p_spl_),
    .din2(g1619_p)
  );


  LA
  g_g1621_p
  (
    .dout(g1621_p),
    .din1(g1615_n_spl_),
    .din2(g1618_n)
  );


  FA
  g_g1621_n
  (
    .dout(g1621_n),
    .din1(g1615_p_spl_),
    .din2(g1618_p_spl_)
  );


  LA
  g_g1622_p
  (
    .dout(g1622_p),
    .din1(g1609_n_spl_),
    .din2(g1612_n_spl_)
  );


  FA
  g_g1622_n
  (
    .dout(g1622_n),
    .din1(g1609_p_spl_),
    .din2(g1612_p_spl_)
  );


  LA
  g_g1623_p
  (
    .dout(g1623_p),
    .din1(G9_p_spl_111),
    .din2(G32_p_spl_100)
  );


  FA
  g_g1623_n
  (
    .dout(g1623_n),
    .din1(G9_n_spl_111),
    .din2(G32_n_spl_100)
  );


  LA
  g_g1624_p
  (
    .dout(g1624_p),
    .din1(g1603_n_spl_),
    .din2(g1606_n_spl_)
  );


  FA
  g_g1624_n
  (
    .dout(g1624_n),
    .din1(g1603_p_spl_),
    .din2(g1606_p_spl_)
  );


  LA
  g_g1625_p
  (
    .dout(g1625_p),
    .din1(G10_p_spl_111),
    .din2(G31_p_spl_100)
  );


  FA
  g_g1625_n
  (
    .dout(g1625_n),
    .din1(G10_n_spl_111),
    .din2(G31_n_spl_100)
  );


  LA
  g_g1626_p
  (
    .dout(g1626_p),
    .din1(g1597_n_spl_),
    .din2(g1600_n_spl_)
  );


  FA
  g_g1626_n
  (
    .dout(g1626_n),
    .din1(g1597_p_spl_),
    .din2(g1600_p_spl_)
  );


  LA
  g_g1627_p
  (
    .dout(g1627_p),
    .din1(G11_p_spl_110),
    .din2(G30_p_spl_101)
  );


  FA
  g_g1627_n
  (
    .dout(g1627_n),
    .din1(G11_n_spl_110),
    .din2(G30_n_spl_101)
  );


  LA
  g_g1628_p
  (
    .dout(g1628_p),
    .din1(g1591_n_spl_),
    .din2(g1594_n_spl_)
  );


  FA
  g_g1628_n
  (
    .dout(g1628_n),
    .din1(g1591_p_spl_),
    .din2(g1594_p_spl_)
  );


  LA
  g_g1629_p
  (
    .dout(g1629_p),
    .din1(G12_p_spl_110),
    .din2(G29_p_spl_101)
  );


  FA
  g_g1629_n
  (
    .dout(g1629_n),
    .din1(G12_n_spl_110),
    .din2(G29_n_spl_101)
  );


  LA
  g_g1630_p
  (
    .dout(g1630_p),
    .din1(g1585_n_spl_),
    .din2(g1588_n_spl_)
  );


  FA
  g_g1630_n
  (
    .dout(g1630_n),
    .din1(g1585_p_spl_),
    .din2(g1588_p_spl_)
  );


  LA
  g_g1631_p
  (
    .dout(g1631_p),
    .din1(G13_p_spl_101),
    .din2(G28_p_spl_110)
  );


  FA
  g_g1631_n
  (
    .dout(g1631_n),
    .din1(G13_n_spl_101),
    .din2(G28_n_spl_110)
  );


  LA
  g_g1632_p
  (
    .dout(g1632_p),
    .din1(g1579_n_spl_),
    .din2(g1582_n_spl_)
  );


  FA
  g_g1632_n
  (
    .dout(g1632_n),
    .din1(g1579_p_spl_),
    .din2(g1582_p_spl_)
  );


  LA
  g_g1633_p
  (
    .dout(g1633_p),
    .din1(G14_p_spl_101),
    .din2(G27_p_spl_110)
  );


  FA
  g_g1633_n
  (
    .dout(g1633_n),
    .din1(G14_n_spl_101),
    .din2(G27_n_spl_110)
  );


  LA
  g_g1634_p
  (
    .dout(g1634_p),
    .din1(g1573_n_spl_),
    .din2(g1576_n_spl_)
  );


  FA
  g_g1634_n
  (
    .dout(g1634_n),
    .din1(g1573_p_spl_),
    .din2(g1576_p_spl_)
  );


  LA
  g_g1635_p
  (
    .dout(g1635_p),
    .din1(G15_p_spl_100),
    .din2(G26_p_spl_111)
  );


  FA
  g_g1635_n
  (
    .dout(g1635_n),
    .din1(G15_n_spl_100),
    .din2(G26_n_spl_111)
  );


  LA
  g_g1636_p
  (
    .dout(g1636_p),
    .din1(G16_p_spl_100),
    .din2(G25_p_spl_111)
  );


  FA
  g_g1636_n
  (
    .dout(g1636_n),
    .din1(G16_n_spl_100),
    .din2(G25_n_spl_111)
  );


  LA
  g_g1637_p
  (
    .dout(g1637_p),
    .din1(g1567_n_spl_),
    .din2(g1570_n_spl_)
  );


  FA
  g_g1637_n
  (
    .dout(g1637_n),
    .din1(g1567_p_spl_),
    .din2(g1570_p_spl_)
  );


  LA
  g_g1638_p
  (
    .dout(g1638_p),
    .din1(g1636_n_spl_),
    .din2(g1637_n_spl_)
  );


  FA
  g_g1638_n
  (
    .dout(g1638_n),
    .din1(g1636_p_spl_),
    .din2(g1637_p_spl_)
  );


  LA
  g_g1639_p
  (
    .dout(g1639_p),
    .din1(g1636_p_spl_),
    .din2(g1637_p_spl_)
  );


  FA
  g_g1639_n
  (
    .dout(g1639_n),
    .din1(g1636_n_spl_),
    .din2(g1637_n_spl_)
  );


  LA
  g_g1640_p
  (
    .dout(g1640_p),
    .din1(g1638_n_spl_),
    .din2(g1639_n)
  );


  FA
  g_g1640_n
  (
    .dout(g1640_n),
    .din1(g1638_p_spl_),
    .din2(g1639_p)
  );


  LA
  g_g1641_p
  (
    .dout(g1641_p),
    .din1(g1635_n_spl_),
    .din2(g1640_p_spl_)
  );


  FA
  g_g1641_n
  (
    .dout(g1641_n),
    .din1(g1635_p_spl_),
    .din2(g1640_n_spl_)
  );


  LA
  g_g1642_p
  (
    .dout(g1642_p),
    .din1(g1635_p_spl_),
    .din2(g1640_n_spl_)
  );


  FA
  g_g1642_n
  (
    .dout(g1642_n),
    .din1(g1635_n_spl_),
    .din2(g1640_p_spl_)
  );


  LA
  g_g1643_p
  (
    .dout(g1643_p),
    .din1(g1641_n_spl_),
    .din2(g1642_n)
  );


  FA
  g_g1643_n
  (
    .dout(g1643_n),
    .din1(g1641_p_spl_),
    .din2(g1642_p)
  );


  LA
  g_g1644_p
  (
    .dout(g1644_p),
    .din1(g1634_n_spl_),
    .din2(g1643_p_spl_)
  );


  FA
  g_g1644_n
  (
    .dout(g1644_n),
    .din1(g1634_p_spl_),
    .din2(g1643_n_spl_)
  );


  LA
  g_g1645_p
  (
    .dout(g1645_p),
    .din1(g1634_p_spl_),
    .din2(g1643_n_spl_)
  );


  FA
  g_g1645_n
  (
    .dout(g1645_n),
    .din1(g1634_n_spl_),
    .din2(g1643_p_spl_)
  );


  LA
  g_g1646_p
  (
    .dout(g1646_p),
    .din1(g1644_n_spl_),
    .din2(g1645_n)
  );


  FA
  g_g1646_n
  (
    .dout(g1646_n),
    .din1(g1644_p_spl_),
    .din2(g1645_p)
  );


  LA
  g_g1647_p
  (
    .dout(g1647_p),
    .din1(g1633_n_spl_),
    .din2(g1646_p_spl_)
  );


  FA
  g_g1647_n
  (
    .dout(g1647_n),
    .din1(g1633_p_spl_),
    .din2(g1646_n_spl_)
  );


  LA
  g_g1648_p
  (
    .dout(g1648_p),
    .din1(g1633_p_spl_),
    .din2(g1646_n_spl_)
  );


  FA
  g_g1648_n
  (
    .dout(g1648_n),
    .din1(g1633_n_spl_),
    .din2(g1646_p_spl_)
  );


  LA
  g_g1649_p
  (
    .dout(g1649_p),
    .din1(g1647_n_spl_),
    .din2(g1648_n)
  );


  FA
  g_g1649_n
  (
    .dout(g1649_n),
    .din1(g1647_p_spl_),
    .din2(g1648_p)
  );


  LA
  g_g1650_p
  (
    .dout(g1650_p),
    .din1(g1632_n_spl_),
    .din2(g1649_p_spl_)
  );


  FA
  g_g1650_n
  (
    .dout(g1650_n),
    .din1(g1632_p_spl_),
    .din2(g1649_n_spl_)
  );


  LA
  g_g1651_p
  (
    .dout(g1651_p),
    .din1(g1632_p_spl_),
    .din2(g1649_n_spl_)
  );


  FA
  g_g1651_n
  (
    .dout(g1651_n),
    .din1(g1632_n_spl_),
    .din2(g1649_p_spl_)
  );


  LA
  g_g1652_p
  (
    .dout(g1652_p),
    .din1(g1650_n_spl_),
    .din2(g1651_n)
  );


  FA
  g_g1652_n
  (
    .dout(g1652_n),
    .din1(g1650_p_spl_),
    .din2(g1651_p)
  );


  LA
  g_g1653_p
  (
    .dout(g1653_p),
    .din1(g1631_n_spl_),
    .din2(g1652_p_spl_)
  );


  FA
  g_g1653_n
  (
    .dout(g1653_n),
    .din1(g1631_p_spl_),
    .din2(g1652_n_spl_)
  );


  LA
  g_g1654_p
  (
    .dout(g1654_p),
    .din1(g1631_p_spl_),
    .din2(g1652_n_spl_)
  );


  FA
  g_g1654_n
  (
    .dout(g1654_n),
    .din1(g1631_n_spl_),
    .din2(g1652_p_spl_)
  );


  LA
  g_g1655_p
  (
    .dout(g1655_p),
    .din1(g1653_n_spl_),
    .din2(g1654_n)
  );


  FA
  g_g1655_n
  (
    .dout(g1655_n),
    .din1(g1653_p_spl_),
    .din2(g1654_p)
  );


  LA
  g_g1656_p
  (
    .dout(g1656_p),
    .din1(g1630_n_spl_),
    .din2(g1655_p_spl_)
  );


  FA
  g_g1656_n
  (
    .dout(g1656_n),
    .din1(g1630_p_spl_),
    .din2(g1655_n_spl_)
  );


  LA
  g_g1657_p
  (
    .dout(g1657_p),
    .din1(g1630_p_spl_),
    .din2(g1655_n_spl_)
  );


  FA
  g_g1657_n
  (
    .dout(g1657_n),
    .din1(g1630_n_spl_),
    .din2(g1655_p_spl_)
  );


  LA
  g_g1658_p
  (
    .dout(g1658_p),
    .din1(g1656_n_spl_),
    .din2(g1657_n)
  );


  FA
  g_g1658_n
  (
    .dout(g1658_n),
    .din1(g1656_p_spl_),
    .din2(g1657_p)
  );


  LA
  g_g1659_p
  (
    .dout(g1659_p),
    .din1(g1629_n_spl_),
    .din2(g1658_p_spl_)
  );


  FA
  g_g1659_n
  (
    .dout(g1659_n),
    .din1(g1629_p_spl_),
    .din2(g1658_n_spl_)
  );


  LA
  g_g1660_p
  (
    .dout(g1660_p),
    .din1(g1629_p_spl_),
    .din2(g1658_n_spl_)
  );


  FA
  g_g1660_n
  (
    .dout(g1660_n),
    .din1(g1629_n_spl_),
    .din2(g1658_p_spl_)
  );


  LA
  g_g1661_p
  (
    .dout(g1661_p),
    .din1(g1659_n_spl_),
    .din2(g1660_n)
  );


  FA
  g_g1661_n
  (
    .dout(g1661_n),
    .din1(g1659_p_spl_),
    .din2(g1660_p)
  );


  LA
  g_g1662_p
  (
    .dout(g1662_p),
    .din1(g1628_n_spl_),
    .din2(g1661_p_spl_)
  );


  FA
  g_g1662_n
  (
    .dout(g1662_n),
    .din1(g1628_p_spl_),
    .din2(g1661_n_spl_)
  );


  LA
  g_g1663_p
  (
    .dout(g1663_p),
    .din1(g1628_p_spl_),
    .din2(g1661_n_spl_)
  );


  FA
  g_g1663_n
  (
    .dout(g1663_n),
    .din1(g1628_n_spl_),
    .din2(g1661_p_spl_)
  );


  LA
  g_g1664_p
  (
    .dout(g1664_p),
    .din1(g1662_n_spl_),
    .din2(g1663_n)
  );


  FA
  g_g1664_n
  (
    .dout(g1664_n),
    .din1(g1662_p_spl_),
    .din2(g1663_p)
  );


  LA
  g_g1665_p
  (
    .dout(g1665_p),
    .din1(g1627_n_spl_),
    .din2(g1664_p_spl_)
  );


  FA
  g_g1665_n
  (
    .dout(g1665_n),
    .din1(g1627_p_spl_),
    .din2(g1664_n_spl_)
  );


  LA
  g_g1666_p
  (
    .dout(g1666_p),
    .din1(g1627_p_spl_),
    .din2(g1664_n_spl_)
  );


  FA
  g_g1666_n
  (
    .dout(g1666_n),
    .din1(g1627_n_spl_),
    .din2(g1664_p_spl_)
  );


  LA
  g_g1667_p
  (
    .dout(g1667_p),
    .din1(g1665_n_spl_),
    .din2(g1666_n)
  );


  FA
  g_g1667_n
  (
    .dout(g1667_n),
    .din1(g1665_p_spl_),
    .din2(g1666_p)
  );


  LA
  g_g1668_p
  (
    .dout(g1668_p),
    .din1(g1626_n_spl_),
    .din2(g1667_p_spl_)
  );


  FA
  g_g1668_n
  (
    .dout(g1668_n),
    .din1(g1626_p_spl_),
    .din2(g1667_n_spl_)
  );


  LA
  g_g1669_p
  (
    .dout(g1669_p),
    .din1(g1626_p_spl_),
    .din2(g1667_n_spl_)
  );


  FA
  g_g1669_n
  (
    .dout(g1669_n),
    .din1(g1626_n_spl_),
    .din2(g1667_p_spl_)
  );


  LA
  g_g1670_p
  (
    .dout(g1670_p),
    .din1(g1668_n_spl_),
    .din2(g1669_n)
  );


  FA
  g_g1670_n
  (
    .dout(g1670_n),
    .din1(g1668_p_spl_),
    .din2(g1669_p)
  );


  LA
  g_g1671_p
  (
    .dout(g1671_p),
    .din1(g1625_n_spl_),
    .din2(g1670_p_spl_)
  );


  FA
  g_g1671_n
  (
    .dout(g1671_n),
    .din1(g1625_p_spl_),
    .din2(g1670_n_spl_)
  );


  LA
  g_g1672_p
  (
    .dout(g1672_p),
    .din1(g1625_p_spl_),
    .din2(g1670_n_spl_)
  );


  FA
  g_g1672_n
  (
    .dout(g1672_n),
    .din1(g1625_n_spl_),
    .din2(g1670_p_spl_)
  );


  LA
  g_g1673_p
  (
    .dout(g1673_p),
    .din1(g1671_n_spl_),
    .din2(g1672_n)
  );


  FA
  g_g1673_n
  (
    .dout(g1673_n),
    .din1(g1671_p_spl_),
    .din2(g1672_p)
  );


  LA
  g_g1674_p
  (
    .dout(g1674_p),
    .din1(g1624_n_spl_),
    .din2(g1673_p_spl_)
  );


  FA
  g_g1674_n
  (
    .dout(g1674_n),
    .din1(g1624_p_spl_),
    .din2(g1673_n_spl_)
  );


  LA
  g_g1675_p
  (
    .dout(g1675_p),
    .din1(g1624_p_spl_),
    .din2(g1673_n_spl_)
  );


  FA
  g_g1675_n
  (
    .dout(g1675_n),
    .din1(g1624_n_spl_),
    .din2(g1673_p_spl_)
  );


  LA
  g_g1676_p
  (
    .dout(g1676_p),
    .din1(g1674_n_spl_),
    .din2(g1675_n)
  );


  FA
  g_g1676_n
  (
    .dout(g1676_n),
    .din1(g1674_p_spl_),
    .din2(g1675_p)
  );


  LA
  g_g1677_p
  (
    .dout(g1677_p),
    .din1(g1623_n_spl_),
    .din2(g1676_p_spl_)
  );


  FA
  g_g1677_n
  (
    .dout(g1677_n),
    .din1(g1623_p_spl_),
    .din2(g1676_n_spl_)
  );


  LA
  g_g1678_p
  (
    .dout(g1678_p),
    .din1(g1623_p_spl_),
    .din2(g1676_n_spl_)
  );


  FA
  g_g1678_n
  (
    .dout(g1678_n),
    .din1(g1623_n_spl_),
    .din2(g1676_p_spl_)
  );


  LA
  g_g1679_p
  (
    .dout(g1679_p),
    .din1(g1677_n_spl_),
    .din2(g1678_n)
  );


  FA
  g_g1679_n
  (
    .dout(g1679_n),
    .din1(g1677_p_spl_),
    .din2(g1678_p)
  );


  LA
  g_g1680_p
  (
    .dout(g1680_p),
    .din1(g1622_n_spl_),
    .din2(g1679_p_spl_)
  );


  FA
  g_g1680_n
  (
    .dout(g1680_n),
    .din1(g1622_p_spl_),
    .din2(g1679_n_spl_)
  );


  LA
  g_g1681_p
  (
    .dout(g1681_p),
    .din1(g1622_p_spl_),
    .din2(g1679_n_spl_)
  );


  FA
  g_g1681_n
  (
    .dout(g1681_n),
    .din1(g1622_n_spl_),
    .din2(g1679_p_spl_)
  );


  LA
  g_g1682_p
  (
    .dout(g1682_p),
    .din1(g1680_n_spl_),
    .din2(g1681_n)
  );


  FA
  g_g1682_n
  (
    .dout(g1682_n),
    .din1(g1680_p_spl_),
    .din2(g1681_p)
  );


  LA
  g_g1683_p
  (
    .dout(g1683_p),
    .din1(g1621_n),
    .din2(g1682_p)
  );


  FA
  g_g1683_n
  (
    .dout(g1683_n),
    .din1(g1621_p_spl_),
    .din2(g1682_n_spl_)
  );


  LA
  g_g1684_p
  (
    .dout(g1684_p),
    .din1(g1621_p_spl_),
    .din2(g1682_n_spl_)
  );


  FA
  g_g1685_n
  (
    .dout(g1685_n),
    .din1(g1683_p_spl_),
    .din2(g1684_p)
  );


  LA
  g_g1686_p
  (
    .dout(g1686_p),
    .din1(g1680_n_spl_),
    .din2(g1683_n)
  );


  FA
  g_g1686_n
  (
    .dout(g1686_n),
    .din1(g1680_p_spl_),
    .din2(g1683_p_spl_)
  );


  LA
  g_g1687_p
  (
    .dout(g1687_p),
    .din1(g1674_n_spl_),
    .din2(g1677_n_spl_)
  );


  FA
  g_g1687_n
  (
    .dout(g1687_n),
    .din1(g1674_p_spl_),
    .din2(g1677_p_spl_)
  );


  LA
  g_g1688_p
  (
    .dout(g1688_p),
    .din1(G10_p_spl_111),
    .din2(G32_p_spl_100)
  );


  FA
  g_g1688_n
  (
    .dout(g1688_n),
    .din1(G10_n_spl_111),
    .din2(G32_n_spl_100)
  );


  LA
  g_g1689_p
  (
    .dout(g1689_p),
    .din1(g1668_n_spl_),
    .din2(g1671_n_spl_)
  );


  FA
  g_g1689_n
  (
    .dout(g1689_n),
    .din1(g1668_p_spl_),
    .din2(g1671_p_spl_)
  );


  LA
  g_g1690_p
  (
    .dout(g1690_p),
    .din1(G11_p_spl_111),
    .din2(G31_p_spl_101)
  );


  FA
  g_g1690_n
  (
    .dout(g1690_n),
    .din1(G11_n_spl_111),
    .din2(G31_n_spl_101)
  );


  LA
  g_g1691_p
  (
    .dout(g1691_p),
    .din1(g1662_n_spl_),
    .din2(g1665_n_spl_)
  );


  FA
  g_g1691_n
  (
    .dout(g1691_n),
    .din1(g1662_p_spl_),
    .din2(g1665_p_spl_)
  );


  LA
  g_g1692_p
  (
    .dout(g1692_p),
    .din1(G12_p_spl_110),
    .din2(G30_p_spl_101)
  );


  FA
  g_g1692_n
  (
    .dout(g1692_n),
    .din1(G12_n_spl_110),
    .din2(G30_n_spl_101)
  );


  LA
  g_g1693_p
  (
    .dout(g1693_p),
    .din1(g1656_n_spl_),
    .din2(g1659_n_spl_)
  );


  FA
  g_g1693_n
  (
    .dout(g1693_n),
    .din1(g1656_p_spl_),
    .din2(g1659_p_spl_)
  );


  LA
  g_g1694_p
  (
    .dout(g1694_p),
    .din1(G13_p_spl_110),
    .din2(G29_p_spl_110)
  );


  FA
  g_g1694_n
  (
    .dout(g1694_n),
    .din1(G13_n_spl_110),
    .din2(G29_n_spl_110)
  );


  LA
  g_g1695_p
  (
    .dout(g1695_p),
    .din1(g1650_n_spl_),
    .din2(g1653_n_spl_)
  );


  FA
  g_g1695_n
  (
    .dout(g1695_n),
    .din1(g1650_p_spl_),
    .din2(g1653_p_spl_)
  );


  LA
  g_g1696_p
  (
    .dout(g1696_p),
    .din1(G14_p_spl_101),
    .din2(G28_p_spl_110)
  );


  FA
  g_g1696_n
  (
    .dout(g1696_n),
    .din1(G14_n_spl_101),
    .din2(G28_n_spl_110)
  );


  LA
  g_g1697_p
  (
    .dout(g1697_p),
    .din1(g1644_n_spl_),
    .din2(g1647_n_spl_)
  );


  FA
  g_g1697_n
  (
    .dout(g1697_n),
    .din1(g1644_p_spl_),
    .din2(g1647_p_spl_)
  );


  LA
  g_g1698_p
  (
    .dout(g1698_p),
    .din1(G15_p_spl_101),
    .din2(G27_p_spl_111)
  );


  FA
  g_g1698_n
  (
    .dout(g1698_n),
    .din1(G15_n_spl_101),
    .din2(G27_n_spl_111)
  );


  LA
  g_g1699_p
  (
    .dout(g1699_p),
    .din1(G16_p_spl_100),
    .din2(G26_p_spl_111)
  );


  FA
  g_g1699_n
  (
    .dout(g1699_n),
    .din1(G16_n_spl_100),
    .din2(G26_n_spl_111)
  );


  LA
  g_g1700_p
  (
    .dout(g1700_p),
    .din1(g1638_n_spl_),
    .din2(g1641_n_spl_)
  );


  FA
  g_g1700_n
  (
    .dout(g1700_n),
    .din1(g1638_p_spl_),
    .din2(g1641_p_spl_)
  );


  LA
  g_g1701_p
  (
    .dout(g1701_p),
    .din1(g1699_n_spl_),
    .din2(g1700_n_spl_)
  );


  FA
  g_g1701_n
  (
    .dout(g1701_n),
    .din1(g1699_p_spl_),
    .din2(g1700_p_spl_)
  );


  LA
  g_g1702_p
  (
    .dout(g1702_p),
    .din1(g1699_p_spl_),
    .din2(g1700_p_spl_)
  );


  FA
  g_g1702_n
  (
    .dout(g1702_n),
    .din1(g1699_n_spl_),
    .din2(g1700_n_spl_)
  );


  LA
  g_g1703_p
  (
    .dout(g1703_p),
    .din1(g1701_n_spl_),
    .din2(g1702_n)
  );


  FA
  g_g1703_n
  (
    .dout(g1703_n),
    .din1(g1701_p_spl_),
    .din2(g1702_p)
  );


  LA
  g_g1704_p
  (
    .dout(g1704_p),
    .din1(g1698_n_spl_),
    .din2(g1703_p_spl_)
  );


  FA
  g_g1704_n
  (
    .dout(g1704_n),
    .din1(g1698_p_spl_),
    .din2(g1703_n_spl_)
  );


  LA
  g_g1705_p
  (
    .dout(g1705_p),
    .din1(g1698_p_spl_),
    .din2(g1703_n_spl_)
  );


  FA
  g_g1705_n
  (
    .dout(g1705_n),
    .din1(g1698_n_spl_),
    .din2(g1703_p_spl_)
  );


  LA
  g_g1706_p
  (
    .dout(g1706_p),
    .din1(g1704_n_spl_),
    .din2(g1705_n)
  );


  FA
  g_g1706_n
  (
    .dout(g1706_n),
    .din1(g1704_p_spl_),
    .din2(g1705_p)
  );


  LA
  g_g1707_p
  (
    .dout(g1707_p),
    .din1(g1697_n_spl_),
    .din2(g1706_p_spl_)
  );


  FA
  g_g1707_n
  (
    .dout(g1707_n),
    .din1(g1697_p_spl_),
    .din2(g1706_n_spl_)
  );


  LA
  g_g1708_p
  (
    .dout(g1708_p),
    .din1(g1697_p_spl_),
    .din2(g1706_n_spl_)
  );


  FA
  g_g1708_n
  (
    .dout(g1708_n),
    .din1(g1697_n_spl_),
    .din2(g1706_p_spl_)
  );


  LA
  g_g1709_p
  (
    .dout(g1709_p),
    .din1(g1707_n_spl_),
    .din2(g1708_n)
  );


  FA
  g_g1709_n
  (
    .dout(g1709_n),
    .din1(g1707_p_spl_),
    .din2(g1708_p)
  );


  LA
  g_g1710_p
  (
    .dout(g1710_p),
    .din1(g1696_n_spl_),
    .din2(g1709_p_spl_)
  );


  FA
  g_g1710_n
  (
    .dout(g1710_n),
    .din1(g1696_p_spl_),
    .din2(g1709_n_spl_)
  );


  LA
  g_g1711_p
  (
    .dout(g1711_p),
    .din1(g1696_p_spl_),
    .din2(g1709_n_spl_)
  );


  FA
  g_g1711_n
  (
    .dout(g1711_n),
    .din1(g1696_n_spl_),
    .din2(g1709_p_spl_)
  );


  LA
  g_g1712_p
  (
    .dout(g1712_p),
    .din1(g1710_n_spl_),
    .din2(g1711_n)
  );


  FA
  g_g1712_n
  (
    .dout(g1712_n),
    .din1(g1710_p_spl_),
    .din2(g1711_p)
  );


  LA
  g_g1713_p
  (
    .dout(g1713_p),
    .din1(g1695_n_spl_),
    .din2(g1712_p_spl_)
  );


  FA
  g_g1713_n
  (
    .dout(g1713_n),
    .din1(g1695_p_spl_),
    .din2(g1712_n_spl_)
  );


  LA
  g_g1714_p
  (
    .dout(g1714_p),
    .din1(g1695_p_spl_),
    .din2(g1712_n_spl_)
  );


  FA
  g_g1714_n
  (
    .dout(g1714_n),
    .din1(g1695_n_spl_),
    .din2(g1712_p_spl_)
  );


  LA
  g_g1715_p
  (
    .dout(g1715_p),
    .din1(g1713_n_spl_),
    .din2(g1714_n)
  );


  FA
  g_g1715_n
  (
    .dout(g1715_n),
    .din1(g1713_p_spl_),
    .din2(g1714_p)
  );


  LA
  g_g1716_p
  (
    .dout(g1716_p),
    .din1(g1694_n_spl_),
    .din2(g1715_p_spl_)
  );


  FA
  g_g1716_n
  (
    .dout(g1716_n),
    .din1(g1694_p_spl_),
    .din2(g1715_n_spl_)
  );


  LA
  g_g1717_p
  (
    .dout(g1717_p),
    .din1(g1694_p_spl_),
    .din2(g1715_n_spl_)
  );


  FA
  g_g1717_n
  (
    .dout(g1717_n),
    .din1(g1694_n_spl_),
    .din2(g1715_p_spl_)
  );


  LA
  g_g1718_p
  (
    .dout(g1718_p),
    .din1(g1716_n_spl_),
    .din2(g1717_n)
  );


  FA
  g_g1718_n
  (
    .dout(g1718_n),
    .din1(g1716_p_spl_),
    .din2(g1717_p)
  );


  LA
  g_g1719_p
  (
    .dout(g1719_p),
    .din1(g1693_n_spl_),
    .din2(g1718_p_spl_)
  );


  FA
  g_g1719_n
  (
    .dout(g1719_n),
    .din1(g1693_p_spl_),
    .din2(g1718_n_spl_)
  );


  LA
  g_g1720_p
  (
    .dout(g1720_p),
    .din1(g1693_p_spl_),
    .din2(g1718_n_spl_)
  );


  FA
  g_g1720_n
  (
    .dout(g1720_n),
    .din1(g1693_n_spl_),
    .din2(g1718_p_spl_)
  );


  LA
  g_g1721_p
  (
    .dout(g1721_p),
    .din1(g1719_n_spl_),
    .din2(g1720_n)
  );


  FA
  g_g1721_n
  (
    .dout(g1721_n),
    .din1(g1719_p_spl_),
    .din2(g1720_p)
  );


  LA
  g_g1722_p
  (
    .dout(g1722_p),
    .din1(g1692_n_spl_),
    .din2(g1721_p_spl_)
  );


  FA
  g_g1722_n
  (
    .dout(g1722_n),
    .din1(g1692_p_spl_),
    .din2(g1721_n_spl_)
  );


  LA
  g_g1723_p
  (
    .dout(g1723_p),
    .din1(g1692_p_spl_),
    .din2(g1721_n_spl_)
  );


  FA
  g_g1723_n
  (
    .dout(g1723_n),
    .din1(g1692_n_spl_),
    .din2(g1721_p_spl_)
  );


  LA
  g_g1724_p
  (
    .dout(g1724_p),
    .din1(g1722_n_spl_),
    .din2(g1723_n)
  );


  FA
  g_g1724_n
  (
    .dout(g1724_n),
    .din1(g1722_p_spl_),
    .din2(g1723_p)
  );


  LA
  g_g1725_p
  (
    .dout(g1725_p),
    .din1(g1691_n_spl_),
    .din2(g1724_p_spl_)
  );


  FA
  g_g1725_n
  (
    .dout(g1725_n),
    .din1(g1691_p_spl_),
    .din2(g1724_n_spl_)
  );


  LA
  g_g1726_p
  (
    .dout(g1726_p),
    .din1(g1691_p_spl_),
    .din2(g1724_n_spl_)
  );


  FA
  g_g1726_n
  (
    .dout(g1726_n),
    .din1(g1691_n_spl_),
    .din2(g1724_p_spl_)
  );


  LA
  g_g1727_p
  (
    .dout(g1727_p),
    .din1(g1725_n_spl_),
    .din2(g1726_n)
  );


  FA
  g_g1727_n
  (
    .dout(g1727_n),
    .din1(g1725_p_spl_),
    .din2(g1726_p)
  );


  LA
  g_g1728_p
  (
    .dout(g1728_p),
    .din1(g1690_n_spl_),
    .din2(g1727_p_spl_)
  );


  FA
  g_g1728_n
  (
    .dout(g1728_n),
    .din1(g1690_p_spl_),
    .din2(g1727_n_spl_)
  );


  LA
  g_g1729_p
  (
    .dout(g1729_p),
    .din1(g1690_p_spl_),
    .din2(g1727_n_spl_)
  );


  FA
  g_g1729_n
  (
    .dout(g1729_n),
    .din1(g1690_n_spl_),
    .din2(g1727_p_spl_)
  );


  LA
  g_g1730_p
  (
    .dout(g1730_p),
    .din1(g1728_n_spl_),
    .din2(g1729_n)
  );


  FA
  g_g1730_n
  (
    .dout(g1730_n),
    .din1(g1728_p_spl_),
    .din2(g1729_p)
  );


  LA
  g_g1731_p
  (
    .dout(g1731_p),
    .din1(g1689_n_spl_),
    .din2(g1730_p_spl_)
  );


  FA
  g_g1731_n
  (
    .dout(g1731_n),
    .din1(g1689_p_spl_),
    .din2(g1730_n_spl_)
  );


  LA
  g_g1732_p
  (
    .dout(g1732_p),
    .din1(g1689_p_spl_),
    .din2(g1730_n_spl_)
  );


  FA
  g_g1732_n
  (
    .dout(g1732_n),
    .din1(g1689_n_spl_),
    .din2(g1730_p_spl_)
  );


  LA
  g_g1733_p
  (
    .dout(g1733_p),
    .din1(g1731_n_spl_),
    .din2(g1732_n)
  );


  FA
  g_g1733_n
  (
    .dout(g1733_n),
    .din1(g1731_p_spl_),
    .din2(g1732_p)
  );


  LA
  g_g1734_p
  (
    .dout(g1734_p),
    .din1(g1688_n_spl_),
    .din2(g1733_p_spl_)
  );


  FA
  g_g1734_n
  (
    .dout(g1734_n),
    .din1(g1688_p_spl_),
    .din2(g1733_n_spl_)
  );


  LA
  g_g1735_p
  (
    .dout(g1735_p),
    .din1(g1688_p_spl_),
    .din2(g1733_n_spl_)
  );


  FA
  g_g1735_n
  (
    .dout(g1735_n),
    .din1(g1688_n_spl_),
    .din2(g1733_p_spl_)
  );


  LA
  g_g1736_p
  (
    .dout(g1736_p),
    .din1(g1734_n_spl_),
    .din2(g1735_n)
  );


  FA
  g_g1736_n
  (
    .dout(g1736_n),
    .din1(g1734_p_spl_),
    .din2(g1735_p)
  );


  LA
  g_g1737_p
  (
    .dout(g1737_p),
    .din1(g1687_n_spl_),
    .din2(g1736_p_spl_)
  );


  FA
  g_g1737_n
  (
    .dout(g1737_n),
    .din1(g1687_p_spl_),
    .din2(g1736_n_spl_)
  );


  LA
  g_g1738_p
  (
    .dout(g1738_p),
    .din1(g1687_p_spl_),
    .din2(g1736_n_spl_)
  );


  FA
  g_g1738_n
  (
    .dout(g1738_n),
    .din1(g1687_n_spl_),
    .din2(g1736_p_spl_)
  );


  LA
  g_g1739_p
  (
    .dout(g1739_p),
    .din1(g1737_n_spl_),
    .din2(g1738_n)
  );


  FA
  g_g1739_n
  (
    .dout(g1739_n),
    .din1(g1737_p_spl_),
    .din2(g1738_p)
  );


  LA
  g_g1740_p
  (
    .dout(g1740_p),
    .din1(g1686_n),
    .din2(g1739_p)
  );


  FA
  g_g1740_n
  (
    .dout(g1740_n),
    .din1(g1686_p_spl_),
    .din2(g1739_n_spl_)
  );


  LA
  g_g1741_p
  (
    .dout(g1741_p),
    .din1(g1686_p_spl_),
    .din2(g1739_n_spl_)
  );


  FA
  g_g1742_n
  (
    .dout(g1742_n),
    .din1(g1740_p_spl_),
    .din2(g1741_p)
  );


  LA
  g_g1743_p
  (
    .dout(g1743_p),
    .din1(g1737_n_spl_),
    .din2(g1740_n)
  );


  FA
  g_g1743_n
  (
    .dout(g1743_n),
    .din1(g1737_p_spl_),
    .din2(g1740_p_spl_)
  );


  LA
  g_g1744_p
  (
    .dout(g1744_p),
    .din1(g1731_n_spl_),
    .din2(g1734_n_spl_)
  );


  FA
  g_g1744_n
  (
    .dout(g1744_n),
    .din1(g1731_p_spl_),
    .din2(g1734_p_spl_)
  );


  LA
  g_g1745_p
  (
    .dout(g1745_p),
    .din1(G11_p_spl_111),
    .din2(G32_p_spl_101)
  );


  FA
  g_g1745_n
  (
    .dout(g1745_n),
    .din1(G11_n_spl_111),
    .din2(G32_n_spl_101)
  );


  LA
  g_g1746_p
  (
    .dout(g1746_p),
    .din1(g1725_n_spl_),
    .din2(g1728_n_spl_)
  );


  FA
  g_g1746_n
  (
    .dout(g1746_n),
    .din1(g1725_p_spl_),
    .din2(g1728_p_spl_)
  );


  LA
  g_g1747_p
  (
    .dout(g1747_p),
    .din1(G12_p_spl_111),
    .din2(G31_p_spl_101)
  );


  FA
  g_g1747_n
  (
    .dout(g1747_n),
    .din1(G12_n_spl_111),
    .din2(G31_n_spl_101)
  );


  LA
  g_g1748_p
  (
    .dout(g1748_p),
    .din1(g1719_n_spl_),
    .din2(g1722_n_spl_)
  );


  FA
  g_g1748_n
  (
    .dout(g1748_n),
    .din1(g1719_p_spl_),
    .din2(g1722_p_spl_)
  );


  LA
  g_g1749_p
  (
    .dout(g1749_p),
    .din1(G13_p_spl_110),
    .din2(G30_p_spl_110)
  );


  FA
  g_g1749_n
  (
    .dout(g1749_n),
    .din1(G13_n_spl_110),
    .din2(G30_n_spl_110)
  );


  LA
  g_g1750_p
  (
    .dout(g1750_p),
    .din1(g1713_n_spl_),
    .din2(g1716_n_spl_)
  );


  FA
  g_g1750_n
  (
    .dout(g1750_n),
    .din1(g1713_p_spl_),
    .din2(g1716_p_spl_)
  );


  LA
  g_g1751_p
  (
    .dout(g1751_p),
    .din1(G14_p_spl_110),
    .din2(G29_p_spl_110)
  );


  FA
  g_g1751_n
  (
    .dout(g1751_n),
    .din1(G14_n_spl_110),
    .din2(G29_n_spl_110)
  );


  LA
  g_g1752_p
  (
    .dout(g1752_p),
    .din1(g1707_n_spl_),
    .din2(g1710_n_spl_)
  );


  FA
  g_g1752_n
  (
    .dout(g1752_n),
    .din1(g1707_p_spl_),
    .din2(g1710_p_spl_)
  );


  LA
  g_g1753_p
  (
    .dout(g1753_p),
    .din1(G15_p_spl_101),
    .din2(G28_p_spl_111)
  );


  FA
  g_g1753_n
  (
    .dout(g1753_n),
    .din1(G15_n_spl_101),
    .din2(G28_n_spl_111)
  );


  LA
  g_g1754_p
  (
    .dout(g1754_p),
    .din1(G16_p_spl_101),
    .din2(G27_p_spl_111)
  );


  FA
  g_g1754_n
  (
    .dout(g1754_n),
    .din1(G16_n_spl_101),
    .din2(G27_n_spl_111)
  );


  LA
  g_g1755_p
  (
    .dout(g1755_p),
    .din1(g1701_n_spl_),
    .din2(g1704_n_spl_)
  );


  FA
  g_g1755_n
  (
    .dout(g1755_n),
    .din1(g1701_p_spl_),
    .din2(g1704_p_spl_)
  );


  LA
  g_g1756_p
  (
    .dout(g1756_p),
    .din1(g1754_n_spl_),
    .din2(g1755_n_spl_)
  );


  FA
  g_g1756_n
  (
    .dout(g1756_n),
    .din1(g1754_p_spl_),
    .din2(g1755_p_spl_)
  );


  LA
  g_g1757_p
  (
    .dout(g1757_p),
    .din1(g1754_p_spl_),
    .din2(g1755_p_spl_)
  );


  FA
  g_g1757_n
  (
    .dout(g1757_n),
    .din1(g1754_n_spl_),
    .din2(g1755_n_spl_)
  );


  LA
  g_g1758_p
  (
    .dout(g1758_p),
    .din1(g1756_n_spl_),
    .din2(g1757_n)
  );


  FA
  g_g1758_n
  (
    .dout(g1758_n),
    .din1(g1756_p_spl_),
    .din2(g1757_p)
  );


  LA
  g_g1759_p
  (
    .dout(g1759_p),
    .din1(g1753_n_spl_),
    .din2(g1758_p_spl_)
  );


  FA
  g_g1759_n
  (
    .dout(g1759_n),
    .din1(g1753_p_spl_),
    .din2(g1758_n_spl_)
  );


  LA
  g_g1760_p
  (
    .dout(g1760_p),
    .din1(g1753_p_spl_),
    .din2(g1758_n_spl_)
  );


  FA
  g_g1760_n
  (
    .dout(g1760_n),
    .din1(g1753_n_spl_),
    .din2(g1758_p_spl_)
  );


  LA
  g_g1761_p
  (
    .dout(g1761_p),
    .din1(g1759_n_spl_),
    .din2(g1760_n)
  );


  FA
  g_g1761_n
  (
    .dout(g1761_n),
    .din1(g1759_p_spl_),
    .din2(g1760_p)
  );


  LA
  g_g1762_p
  (
    .dout(g1762_p),
    .din1(g1752_n_spl_),
    .din2(g1761_p_spl_)
  );


  FA
  g_g1762_n
  (
    .dout(g1762_n),
    .din1(g1752_p_spl_),
    .din2(g1761_n_spl_)
  );


  LA
  g_g1763_p
  (
    .dout(g1763_p),
    .din1(g1752_p_spl_),
    .din2(g1761_n_spl_)
  );


  FA
  g_g1763_n
  (
    .dout(g1763_n),
    .din1(g1752_n_spl_),
    .din2(g1761_p_spl_)
  );


  LA
  g_g1764_p
  (
    .dout(g1764_p),
    .din1(g1762_n_spl_),
    .din2(g1763_n)
  );


  FA
  g_g1764_n
  (
    .dout(g1764_n),
    .din1(g1762_p_spl_),
    .din2(g1763_p)
  );


  LA
  g_g1765_p
  (
    .dout(g1765_p),
    .din1(g1751_n_spl_),
    .din2(g1764_p_spl_)
  );


  FA
  g_g1765_n
  (
    .dout(g1765_n),
    .din1(g1751_p_spl_),
    .din2(g1764_n_spl_)
  );


  LA
  g_g1766_p
  (
    .dout(g1766_p),
    .din1(g1751_p_spl_),
    .din2(g1764_n_spl_)
  );


  FA
  g_g1766_n
  (
    .dout(g1766_n),
    .din1(g1751_n_spl_),
    .din2(g1764_p_spl_)
  );


  LA
  g_g1767_p
  (
    .dout(g1767_p),
    .din1(g1765_n_spl_),
    .din2(g1766_n)
  );


  FA
  g_g1767_n
  (
    .dout(g1767_n),
    .din1(g1765_p_spl_),
    .din2(g1766_p)
  );


  LA
  g_g1768_p
  (
    .dout(g1768_p),
    .din1(g1750_n_spl_),
    .din2(g1767_p_spl_)
  );


  FA
  g_g1768_n
  (
    .dout(g1768_n),
    .din1(g1750_p_spl_),
    .din2(g1767_n_spl_)
  );


  LA
  g_g1769_p
  (
    .dout(g1769_p),
    .din1(g1750_p_spl_),
    .din2(g1767_n_spl_)
  );


  FA
  g_g1769_n
  (
    .dout(g1769_n),
    .din1(g1750_n_spl_),
    .din2(g1767_p_spl_)
  );


  LA
  g_g1770_p
  (
    .dout(g1770_p),
    .din1(g1768_n_spl_),
    .din2(g1769_n)
  );


  FA
  g_g1770_n
  (
    .dout(g1770_n),
    .din1(g1768_p_spl_),
    .din2(g1769_p)
  );


  LA
  g_g1771_p
  (
    .dout(g1771_p),
    .din1(g1749_n_spl_),
    .din2(g1770_p_spl_)
  );


  FA
  g_g1771_n
  (
    .dout(g1771_n),
    .din1(g1749_p_spl_),
    .din2(g1770_n_spl_)
  );


  LA
  g_g1772_p
  (
    .dout(g1772_p),
    .din1(g1749_p_spl_),
    .din2(g1770_n_spl_)
  );


  FA
  g_g1772_n
  (
    .dout(g1772_n),
    .din1(g1749_n_spl_),
    .din2(g1770_p_spl_)
  );


  LA
  g_g1773_p
  (
    .dout(g1773_p),
    .din1(g1771_n_spl_),
    .din2(g1772_n)
  );


  FA
  g_g1773_n
  (
    .dout(g1773_n),
    .din1(g1771_p_spl_),
    .din2(g1772_p)
  );


  LA
  g_g1774_p
  (
    .dout(g1774_p),
    .din1(g1748_n_spl_),
    .din2(g1773_p_spl_)
  );


  FA
  g_g1774_n
  (
    .dout(g1774_n),
    .din1(g1748_p_spl_),
    .din2(g1773_n_spl_)
  );


  LA
  g_g1775_p
  (
    .dout(g1775_p),
    .din1(g1748_p_spl_),
    .din2(g1773_n_spl_)
  );


  FA
  g_g1775_n
  (
    .dout(g1775_n),
    .din1(g1748_n_spl_),
    .din2(g1773_p_spl_)
  );


  LA
  g_g1776_p
  (
    .dout(g1776_p),
    .din1(g1774_n_spl_),
    .din2(g1775_n)
  );


  FA
  g_g1776_n
  (
    .dout(g1776_n),
    .din1(g1774_p_spl_),
    .din2(g1775_p)
  );


  LA
  g_g1777_p
  (
    .dout(g1777_p),
    .din1(g1747_n_spl_),
    .din2(g1776_p_spl_)
  );


  FA
  g_g1777_n
  (
    .dout(g1777_n),
    .din1(g1747_p_spl_),
    .din2(g1776_n_spl_)
  );


  LA
  g_g1778_p
  (
    .dout(g1778_p),
    .din1(g1747_p_spl_),
    .din2(g1776_n_spl_)
  );


  FA
  g_g1778_n
  (
    .dout(g1778_n),
    .din1(g1747_n_spl_),
    .din2(g1776_p_spl_)
  );


  LA
  g_g1779_p
  (
    .dout(g1779_p),
    .din1(g1777_n_spl_),
    .din2(g1778_n)
  );


  FA
  g_g1779_n
  (
    .dout(g1779_n),
    .din1(g1777_p_spl_),
    .din2(g1778_p)
  );


  LA
  g_g1780_p
  (
    .dout(g1780_p),
    .din1(g1746_n_spl_),
    .din2(g1779_p_spl_)
  );


  FA
  g_g1780_n
  (
    .dout(g1780_n),
    .din1(g1746_p_spl_),
    .din2(g1779_n_spl_)
  );


  LA
  g_g1781_p
  (
    .dout(g1781_p),
    .din1(g1746_p_spl_),
    .din2(g1779_n_spl_)
  );


  FA
  g_g1781_n
  (
    .dout(g1781_n),
    .din1(g1746_n_spl_),
    .din2(g1779_p_spl_)
  );


  LA
  g_g1782_p
  (
    .dout(g1782_p),
    .din1(g1780_n_spl_),
    .din2(g1781_n)
  );


  FA
  g_g1782_n
  (
    .dout(g1782_n),
    .din1(g1780_p_spl_),
    .din2(g1781_p)
  );


  LA
  g_g1783_p
  (
    .dout(g1783_p),
    .din1(g1745_n_spl_),
    .din2(g1782_p_spl_)
  );


  FA
  g_g1783_n
  (
    .dout(g1783_n),
    .din1(g1745_p_spl_),
    .din2(g1782_n_spl_)
  );


  LA
  g_g1784_p
  (
    .dout(g1784_p),
    .din1(g1745_p_spl_),
    .din2(g1782_n_spl_)
  );


  FA
  g_g1784_n
  (
    .dout(g1784_n),
    .din1(g1745_n_spl_),
    .din2(g1782_p_spl_)
  );


  LA
  g_g1785_p
  (
    .dout(g1785_p),
    .din1(g1783_n_spl_),
    .din2(g1784_n)
  );


  FA
  g_g1785_n
  (
    .dout(g1785_n),
    .din1(g1783_p_spl_),
    .din2(g1784_p)
  );


  LA
  g_g1786_p
  (
    .dout(g1786_p),
    .din1(g1744_n_spl_),
    .din2(g1785_p_spl_)
  );


  FA
  g_g1786_n
  (
    .dout(g1786_n),
    .din1(g1744_p_spl_),
    .din2(g1785_n_spl_)
  );


  LA
  g_g1787_p
  (
    .dout(g1787_p),
    .din1(g1744_p_spl_),
    .din2(g1785_n_spl_)
  );


  FA
  g_g1787_n
  (
    .dout(g1787_n),
    .din1(g1744_n_spl_),
    .din2(g1785_p_spl_)
  );


  LA
  g_g1788_p
  (
    .dout(g1788_p),
    .din1(g1786_n_spl_),
    .din2(g1787_n)
  );


  FA
  g_g1788_n
  (
    .dout(g1788_n),
    .din1(g1786_p_spl_),
    .din2(g1787_p)
  );


  LA
  g_g1789_p
  (
    .dout(g1789_p),
    .din1(g1743_n),
    .din2(g1788_p)
  );


  FA
  g_g1789_n
  (
    .dout(g1789_n),
    .din1(g1743_p_spl_),
    .din2(g1788_n_spl_)
  );


  LA
  g_g1790_p
  (
    .dout(g1790_p),
    .din1(g1743_p_spl_),
    .din2(g1788_n_spl_)
  );


  FA
  g_g1791_n
  (
    .dout(g1791_n),
    .din1(g1789_p_spl_),
    .din2(g1790_p)
  );


  LA
  g_g1792_p
  (
    .dout(g1792_p),
    .din1(g1786_n_spl_),
    .din2(g1789_n)
  );


  FA
  g_g1792_n
  (
    .dout(g1792_n),
    .din1(g1786_p_spl_),
    .din2(g1789_p_spl_)
  );


  LA
  g_g1793_p
  (
    .dout(g1793_p),
    .din1(g1780_n_spl_),
    .din2(g1783_n_spl_)
  );


  FA
  g_g1793_n
  (
    .dout(g1793_n),
    .din1(g1780_p_spl_),
    .din2(g1783_p_spl_)
  );


  LA
  g_g1794_p
  (
    .dout(g1794_p),
    .din1(G12_p_spl_111),
    .din2(G32_p_spl_101)
  );


  FA
  g_g1794_n
  (
    .dout(g1794_n),
    .din1(G12_n_spl_111),
    .din2(G32_n_spl_101)
  );


  LA
  g_g1795_p
  (
    .dout(g1795_p),
    .din1(g1774_n_spl_),
    .din2(g1777_n_spl_)
  );


  FA
  g_g1795_n
  (
    .dout(g1795_n),
    .din1(g1774_p_spl_),
    .din2(g1777_p_spl_)
  );


  LA
  g_g1796_p
  (
    .dout(g1796_p),
    .din1(G13_p_spl_111),
    .din2(G31_p_spl_110)
  );


  FA
  g_g1796_n
  (
    .dout(g1796_n),
    .din1(G13_n_spl_111),
    .din2(G31_n_spl_110)
  );


  LA
  g_g1797_p
  (
    .dout(g1797_p),
    .din1(g1768_n_spl_),
    .din2(g1771_n_spl_)
  );


  FA
  g_g1797_n
  (
    .dout(g1797_n),
    .din1(g1768_p_spl_),
    .din2(g1771_p_spl_)
  );


  LA
  g_g1798_p
  (
    .dout(g1798_p),
    .din1(G14_p_spl_110),
    .din2(G30_p_spl_110)
  );


  FA
  g_g1798_n
  (
    .dout(g1798_n),
    .din1(G14_n_spl_110),
    .din2(G30_n_spl_110)
  );


  LA
  g_g1799_p
  (
    .dout(g1799_p),
    .din1(g1762_n_spl_),
    .din2(g1765_n_spl_)
  );


  FA
  g_g1799_n
  (
    .dout(g1799_n),
    .din1(g1762_p_spl_),
    .din2(g1765_p_spl_)
  );


  LA
  g_g1800_p
  (
    .dout(g1800_p),
    .din1(G15_p_spl_110),
    .din2(G29_p_spl_111)
  );


  FA
  g_g1800_n
  (
    .dout(g1800_n),
    .din1(G15_n_spl_110),
    .din2(G29_n_spl_111)
  );


  LA
  g_g1801_p
  (
    .dout(g1801_p),
    .din1(G16_p_spl_101),
    .din2(G28_p_spl_111)
  );


  FA
  g_g1801_n
  (
    .dout(g1801_n),
    .din1(G16_n_spl_101),
    .din2(G28_n_spl_111)
  );


  LA
  g_g1802_p
  (
    .dout(g1802_p),
    .din1(g1756_n_spl_),
    .din2(g1759_n_spl_)
  );


  FA
  g_g1802_n
  (
    .dout(g1802_n),
    .din1(g1756_p_spl_),
    .din2(g1759_p_spl_)
  );


  LA
  g_g1803_p
  (
    .dout(g1803_p),
    .din1(g1801_n_spl_),
    .din2(g1802_n_spl_)
  );


  FA
  g_g1803_n
  (
    .dout(g1803_n),
    .din1(g1801_p_spl_),
    .din2(g1802_p_spl_)
  );


  LA
  g_g1804_p
  (
    .dout(g1804_p),
    .din1(g1801_p_spl_),
    .din2(g1802_p_spl_)
  );


  FA
  g_g1804_n
  (
    .dout(g1804_n),
    .din1(g1801_n_spl_),
    .din2(g1802_n_spl_)
  );


  LA
  g_g1805_p
  (
    .dout(g1805_p),
    .din1(g1803_n_spl_),
    .din2(g1804_n)
  );


  FA
  g_g1805_n
  (
    .dout(g1805_n),
    .din1(g1803_p_spl_),
    .din2(g1804_p)
  );


  LA
  g_g1806_p
  (
    .dout(g1806_p),
    .din1(g1800_n_spl_),
    .din2(g1805_p_spl_)
  );


  FA
  g_g1806_n
  (
    .dout(g1806_n),
    .din1(g1800_p_spl_),
    .din2(g1805_n_spl_)
  );


  LA
  g_g1807_p
  (
    .dout(g1807_p),
    .din1(g1800_p_spl_),
    .din2(g1805_n_spl_)
  );


  FA
  g_g1807_n
  (
    .dout(g1807_n),
    .din1(g1800_n_spl_),
    .din2(g1805_p_spl_)
  );


  LA
  g_g1808_p
  (
    .dout(g1808_p),
    .din1(g1806_n_spl_),
    .din2(g1807_n)
  );


  FA
  g_g1808_n
  (
    .dout(g1808_n),
    .din1(g1806_p_spl_),
    .din2(g1807_p)
  );


  LA
  g_g1809_p
  (
    .dout(g1809_p),
    .din1(g1799_n_spl_),
    .din2(g1808_p_spl_)
  );


  FA
  g_g1809_n
  (
    .dout(g1809_n),
    .din1(g1799_p_spl_),
    .din2(g1808_n_spl_)
  );


  LA
  g_g1810_p
  (
    .dout(g1810_p),
    .din1(g1799_p_spl_),
    .din2(g1808_n_spl_)
  );


  FA
  g_g1810_n
  (
    .dout(g1810_n),
    .din1(g1799_n_spl_),
    .din2(g1808_p_spl_)
  );


  LA
  g_g1811_p
  (
    .dout(g1811_p),
    .din1(g1809_n_spl_),
    .din2(g1810_n)
  );


  FA
  g_g1811_n
  (
    .dout(g1811_n),
    .din1(g1809_p_spl_),
    .din2(g1810_p)
  );


  LA
  g_g1812_p
  (
    .dout(g1812_p),
    .din1(g1798_n_spl_),
    .din2(g1811_p_spl_)
  );


  FA
  g_g1812_n
  (
    .dout(g1812_n),
    .din1(g1798_p_spl_),
    .din2(g1811_n_spl_)
  );


  LA
  g_g1813_p
  (
    .dout(g1813_p),
    .din1(g1798_p_spl_),
    .din2(g1811_n_spl_)
  );


  FA
  g_g1813_n
  (
    .dout(g1813_n),
    .din1(g1798_n_spl_),
    .din2(g1811_p_spl_)
  );


  LA
  g_g1814_p
  (
    .dout(g1814_p),
    .din1(g1812_n_spl_),
    .din2(g1813_n)
  );


  FA
  g_g1814_n
  (
    .dout(g1814_n),
    .din1(g1812_p_spl_),
    .din2(g1813_p)
  );


  LA
  g_g1815_p
  (
    .dout(g1815_p),
    .din1(g1797_n_spl_),
    .din2(g1814_p_spl_)
  );


  FA
  g_g1815_n
  (
    .dout(g1815_n),
    .din1(g1797_p_spl_),
    .din2(g1814_n_spl_)
  );


  LA
  g_g1816_p
  (
    .dout(g1816_p),
    .din1(g1797_p_spl_),
    .din2(g1814_n_spl_)
  );


  FA
  g_g1816_n
  (
    .dout(g1816_n),
    .din1(g1797_n_spl_),
    .din2(g1814_p_spl_)
  );


  LA
  g_g1817_p
  (
    .dout(g1817_p),
    .din1(g1815_n_spl_),
    .din2(g1816_n)
  );


  FA
  g_g1817_n
  (
    .dout(g1817_n),
    .din1(g1815_p_spl_),
    .din2(g1816_p)
  );


  LA
  g_g1818_p
  (
    .dout(g1818_p),
    .din1(g1796_n_spl_),
    .din2(g1817_p_spl_)
  );


  FA
  g_g1818_n
  (
    .dout(g1818_n),
    .din1(g1796_p_spl_),
    .din2(g1817_n_spl_)
  );


  LA
  g_g1819_p
  (
    .dout(g1819_p),
    .din1(g1796_p_spl_),
    .din2(g1817_n_spl_)
  );


  FA
  g_g1819_n
  (
    .dout(g1819_n),
    .din1(g1796_n_spl_),
    .din2(g1817_p_spl_)
  );


  LA
  g_g1820_p
  (
    .dout(g1820_p),
    .din1(g1818_n_spl_),
    .din2(g1819_n)
  );


  FA
  g_g1820_n
  (
    .dout(g1820_n),
    .din1(g1818_p_spl_),
    .din2(g1819_p)
  );


  LA
  g_g1821_p
  (
    .dout(g1821_p),
    .din1(g1795_n_spl_),
    .din2(g1820_p_spl_)
  );


  FA
  g_g1821_n
  (
    .dout(g1821_n),
    .din1(g1795_p_spl_),
    .din2(g1820_n_spl_)
  );


  LA
  g_g1822_p
  (
    .dout(g1822_p),
    .din1(g1795_p_spl_),
    .din2(g1820_n_spl_)
  );


  FA
  g_g1822_n
  (
    .dout(g1822_n),
    .din1(g1795_n_spl_),
    .din2(g1820_p_spl_)
  );


  LA
  g_g1823_p
  (
    .dout(g1823_p),
    .din1(g1821_n_spl_),
    .din2(g1822_n)
  );


  FA
  g_g1823_n
  (
    .dout(g1823_n),
    .din1(g1821_p_spl_),
    .din2(g1822_p)
  );


  LA
  g_g1824_p
  (
    .dout(g1824_p),
    .din1(g1794_n_spl_),
    .din2(g1823_p_spl_)
  );


  FA
  g_g1824_n
  (
    .dout(g1824_n),
    .din1(g1794_p_spl_),
    .din2(g1823_n_spl_)
  );


  LA
  g_g1825_p
  (
    .dout(g1825_p),
    .din1(g1794_p_spl_),
    .din2(g1823_n_spl_)
  );


  FA
  g_g1825_n
  (
    .dout(g1825_n),
    .din1(g1794_n_spl_),
    .din2(g1823_p_spl_)
  );


  LA
  g_g1826_p
  (
    .dout(g1826_p),
    .din1(g1824_n_spl_),
    .din2(g1825_n)
  );


  FA
  g_g1826_n
  (
    .dout(g1826_n),
    .din1(g1824_p_spl_),
    .din2(g1825_p)
  );


  LA
  g_g1827_p
  (
    .dout(g1827_p),
    .din1(g1793_n_spl_),
    .din2(g1826_p_spl_)
  );


  FA
  g_g1827_n
  (
    .dout(g1827_n),
    .din1(g1793_p_spl_),
    .din2(g1826_n_spl_)
  );


  LA
  g_g1828_p
  (
    .dout(g1828_p),
    .din1(g1793_p_spl_),
    .din2(g1826_n_spl_)
  );


  FA
  g_g1828_n
  (
    .dout(g1828_n),
    .din1(g1793_n_spl_),
    .din2(g1826_p_spl_)
  );


  LA
  g_g1829_p
  (
    .dout(g1829_p),
    .din1(g1827_n_spl_),
    .din2(g1828_n)
  );


  FA
  g_g1829_n
  (
    .dout(g1829_n),
    .din1(g1827_p_spl_),
    .din2(g1828_p)
  );


  LA
  g_g1830_p
  (
    .dout(g1830_p),
    .din1(g1792_n),
    .din2(g1829_p)
  );


  FA
  g_g1830_n
  (
    .dout(g1830_n),
    .din1(g1792_p_spl_),
    .din2(g1829_n_spl_)
  );


  LA
  g_g1831_p
  (
    .dout(g1831_p),
    .din1(g1792_p_spl_),
    .din2(g1829_n_spl_)
  );


  FA
  g_g1832_n
  (
    .dout(g1832_n),
    .din1(g1830_p_spl_),
    .din2(g1831_p)
  );


  LA
  g_g1833_p
  (
    .dout(g1833_p),
    .din1(g1827_n_spl_),
    .din2(g1830_n)
  );


  FA
  g_g1833_n
  (
    .dout(g1833_n),
    .din1(g1827_p_spl_),
    .din2(g1830_p_spl_)
  );


  LA
  g_g1834_p
  (
    .dout(g1834_p),
    .din1(g1821_n_spl_),
    .din2(g1824_n_spl_)
  );


  FA
  g_g1834_n
  (
    .dout(g1834_n),
    .din1(g1821_p_spl_),
    .din2(g1824_p_spl_)
  );


  LA
  g_g1835_p
  (
    .dout(g1835_p),
    .din1(G13_p_spl_111),
    .din2(G32_p_spl_110)
  );


  FA
  g_g1835_n
  (
    .dout(g1835_n),
    .din1(G13_n_spl_111),
    .din2(G32_n_spl_110)
  );


  LA
  g_g1836_p
  (
    .dout(g1836_p),
    .din1(g1815_n_spl_),
    .din2(g1818_n_spl_)
  );


  FA
  g_g1836_n
  (
    .dout(g1836_n),
    .din1(g1815_p_spl_),
    .din2(g1818_p_spl_)
  );


  LA
  g_g1837_p
  (
    .dout(g1837_p),
    .din1(G14_p_spl_111),
    .din2(G31_p_spl_110)
  );


  FA
  g_g1837_n
  (
    .dout(g1837_n),
    .din1(G14_n_spl_111),
    .din2(G31_n_spl_110)
  );


  LA
  g_g1838_p
  (
    .dout(g1838_p),
    .din1(g1809_n_spl_),
    .din2(g1812_n_spl_)
  );


  FA
  g_g1838_n
  (
    .dout(g1838_n),
    .din1(g1809_p_spl_),
    .din2(g1812_p_spl_)
  );


  LA
  g_g1839_p
  (
    .dout(g1839_p),
    .din1(G15_p_spl_110),
    .din2(G30_p_spl_111)
  );


  FA
  g_g1839_n
  (
    .dout(g1839_n),
    .din1(G15_n_spl_110),
    .din2(G30_n_spl_111)
  );


  LA
  g_g1840_p
  (
    .dout(g1840_p),
    .din1(G16_p_spl_110),
    .din2(G29_p_spl_111)
  );


  FA
  g_g1840_n
  (
    .dout(g1840_n),
    .din1(G16_n_spl_110),
    .din2(G29_n_spl_111)
  );


  LA
  g_g1841_p
  (
    .dout(g1841_p),
    .din1(g1803_n_spl_),
    .din2(g1806_n_spl_)
  );


  FA
  g_g1841_n
  (
    .dout(g1841_n),
    .din1(g1803_p_spl_),
    .din2(g1806_p_spl_)
  );


  LA
  g_g1842_p
  (
    .dout(g1842_p),
    .din1(g1840_n_spl_),
    .din2(g1841_n_spl_)
  );


  FA
  g_g1842_n
  (
    .dout(g1842_n),
    .din1(g1840_p_spl_),
    .din2(g1841_p_spl_)
  );


  LA
  g_g1843_p
  (
    .dout(g1843_p),
    .din1(g1840_p_spl_),
    .din2(g1841_p_spl_)
  );


  FA
  g_g1843_n
  (
    .dout(g1843_n),
    .din1(g1840_n_spl_),
    .din2(g1841_n_spl_)
  );


  LA
  g_g1844_p
  (
    .dout(g1844_p),
    .din1(g1842_n_spl_),
    .din2(g1843_n)
  );


  FA
  g_g1844_n
  (
    .dout(g1844_n),
    .din1(g1842_p_spl_),
    .din2(g1843_p)
  );


  LA
  g_g1845_p
  (
    .dout(g1845_p),
    .din1(g1839_n_spl_),
    .din2(g1844_p_spl_)
  );


  FA
  g_g1845_n
  (
    .dout(g1845_n),
    .din1(g1839_p_spl_),
    .din2(g1844_n_spl_)
  );


  LA
  g_g1846_p
  (
    .dout(g1846_p),
    .din1(g1839_p_spl_),
    .din2(g1844_n_spl_)
  );


  FA
  g_g1846_n
  (
    .dout(g1846_n),
    .din1(g1839_n_spl_),
    .din2(g1844_p_spl_)
  );


  LA
  g_g1847_p
  (
    .dout(g1847_p),
    .din1(g1845_n_spl_),
    .din2(g1846_n)
  );


  FA
  g_g1847_n
  (
    .dout(g1847_n),
    .din1(g1845_p_spl_),
    .din2(g1846_p)
  );


  LA
  g_g1848_p
  (
    .dout(g1848_p),
    .din1(g1838_n_spl_),
    .din2(g1847_p_spl_)
  );


  FA
  g_g1848_n
  (
    .dout(g1848_n),
    .din1(g1838_p_spl_),
    .din2(g1847_n_spl_)
  );


  LA
  g_g1849_p
  (
    .dout(g1849_p),
    .din1(g1838_p_spl_),
    .din2(g1847_n_spl_)
  );


  FA
  g_g1849_n
  (
    .dout(g1849_n),
    .din1(g1838_n_spl_),
    .din2(g1847_p_spl_)
  );


  LA
  g_g1850_p
  (
    .dout(g1850_p),
    .din1(g1848_n_spl_),
    .din2(g1849_n)
  );


  FA
  g_g1850_n
  (
    .dout(g1850_n),
    .din1(g1848_p_spl_),
    .din2(g1849_p)
  );


  LA
  g_g1851_p
  (
    .dout(g1851_p),
    .din1(g1837_n_spl_),
    .din2(g1850_p_spl_)
  );


  FA
  g_g1851_n
  (
    .dout(g1851_n),
    .din1(g1837_p_spl_),
    .din2(g1850_n_spl_)
  );


  LA
  g_g1852_p
  (
    .dout(g1852_p),
    .din1(g1837_p_spl_),
    .din2(g1850_n_spl_)
  );


  FA
  g_g1852_n
  (
    .dout(g1852_n),
    .din1(g1837_n_spl_),
    .din2(g1850_p_spl_)
  );


  LA
  g_g1853_p
  (
    .dout(g1853_p),
    .din1(g1851_n_spl_),
    .din2(g1852_n)
  );


  FA
  g_g1853_n
  (
    .dout(g1853_n),
    .din1(g1851_p_spl_),
    .din2(g1852_p)
  );


  LA
  g_g1854_p
  (
    .dout(g1854_p),
    .din1(g1836_n_spl_),
    .din2(g1853_p_spl_)
  );


  FA
  g_g1854_n
  (
    .dout(g1854_n),
    .din1(g1836_p_spl_),
    .din2(g1853_n_spl_)
  );


  LA
  g_g1855_p
  (
    .dout(g1855_p),
    .din1(g1836_p_spl_),
    .din2(g1853_n_spl_)
  );


  FA
  g_g1855_n
  (
    .dout(g1855_n),
    .din1(g1836_n_spl_),
    .din2(g1853_p_spl_)
  );


  LA
  g_g1856_p
  (
    .dout(g1856_p),
    .din1(g1854_n_spl_),
    .din2(g1855_n)
  );


  FA
  g_g1856_n
  (
    .dout(g1856_n),
    .din1(g1854_p_spl_),
    .din2(g1855_p)
  );


  LA
  g_g1857_p
  (
    .dout(g1857_p),
    .din1(g1835_n_spl_),
    .din2(g1856_p_spl_)
  );


  FA
  g_g1857_n
  (
    .dout(g1857_n),
    .din1(g1835_p_spl_),
    .din2(g1856_n_spl_)
  );


  LA
  g_g1858_p
  (
    .dout(g1858_p),
    .din1(g1835_p_spl_),
    .din2(g1856_n_spl_)
  );


  FA
  g_g1858_n
  (
    .dout(g1858_n),
    .din1(g1835_n_spl_),
    .din2(g1856_p_spl_)
  );


  LA
  g_g1859_p
  (
    .dout(g1859_p),
    .din1(g1857_n_spl_),
    .din2(g1858_n)
  );


  FA
  g_g1859_n
  (
    .dout(g1859_n),
    .din1(g1857_p_spl_),
    .din2(g1858_p)
  );


  LA
  g_g1860_p
  (
    .dout(g1860_p),
    .din1(g1834_n_spl_),
    .din2(g1859_p_spl_)
  );


  FA
  g_g1860_n
  (
    .dout(g1860_n),
    .din1(g1834_p_spl_),
    .din2(g1859_n_spl_)
  );


  LA
  g_g1861_p
  (
    .dout(g1861_p),
    .din1(g1834_p_spl_),
    .din2(g1859_n_spl_)
  );


  FA
  g_g1861_n
  (
    .dout(g1861_n),
    .din1(g1834_n_spl_),
    .din2(g1859_p_spl_)
  );


  LA
  g_g1862_p
  (
    .dout(g1862_p),
    .din1(g1860_n_spl_),
    .din2(g1861_n)
  );


  FA
  g_g1862_n
  (
    .dout(g1862_n),
    .din1(g1860_p_spl_),
    .din2(g1861_p)
  );


  LA
  g_g1863_p
  (
    .dout(g1863_p),
    .din1(g1833_n),
    .din2(g1862_p)
  );


  FA
  g_g1863_n
  (
    .dout(g1863_n),
    .din1(g1833_p_spl_),
    .din2(g1862_n_spl_)
  );


  LA
  g_g1864_p
  (
    .dout(g1864_p),
    .din1(g1833_p_spl_),
    .din2(g1862_n_spl_)
  );


  FA
  g_g1865_n
  (
    .dout(g1865_n),
    .din1(g1863_p_spl_),
    .din2(g1864_p)
  );


  LA
  g_g1866_p
  (
    .dout(g1866_p),
    .din1(g1860_n_spl_),
    .din2(g1863_n)
  );


  FA
  g_g1866_n
  (
    .dout(g1866_n),
    .din1(g1860_p_spl_),
    .din2(g1863_p_spl_)
  );


  LA
  g_g1867_p
  (
    .dout(g1867_p),
    .din1(g1854_n_spl_),
    .din2(g1857_n_spl_)
  );


  FA
  g_g1867_n
  (
    .dout(g1867_n),
    .din1(g1854_p_spl_),
    .din2(g1857_p_spl_)
  );


  LA
  g_g1868_p
  (
    .dout(g1868_p),
    .din1(G14_p_spl_111),
    .din2(G32_p_spl_110)
  );


  FA
  g_g1868_n
  (
    .dout(g1868_n),
    .din1(G14_n_spl_111),
    .din2(G32_n_spl_110)
  );


  LA
  g_g1869_p
  (
    .dout(g1869_p),
    .din1(g1848_n_spl_),
    .din2(g1851_n_spl_)
  );


  FA
  g_g1869_n
  (
    .dout(g1869_n),
    .din1(g1848_p_spl_),
    .din2(g1851_p_spl_)
  );


  LA
  g_g1870_p
  (
    .dout(g1870_p),
    .din1(G15_p_spl_111),
    .din2(G31_p_spl_111)
  );


  FA
  g_g1870_n
  (
    .dout(g1870_n),
    .din1(G15_n_spl_111),
    .din2(G31_n_spl_111)
  );


  LA
  g_g1871_p
  (
    .dout(g1871_p),
    .din1(G16_p_spl_110),
    .din2(G30_p_spl_111)
  );


  FA
  g_g1871_n
  (
    .dout(g1871_n),
    .din1(G16_n_spl_110),
    .din2(G30_n_spl_111)
  );


  LA
  g_g1872_p
  (
    .dout(g1872_p),
    .din1(g1842_n_spl_),
    .din2(g1845_n_spl_)
  );


  FA
  g_g1872_n
  (
    .dout(g1872_n),
    .din1(g1842_p_spl_),
    .din2(g1845_p_spl_)
  );


  LA
  g_g1873_p
  (
    .dout(g1873_p),
    .din1(g1871_n_spl_),
    .din2(g1872_n_spl_)
  );


  FA
  g_g1873_n
  (
    .dout(g1873_n),
    .din1(g1871_p_spl_),
    .din2(g1872_p_spl_)
  );


  LA
  g_g1874_p
  (
    .dout(g1874_p),
    .din1(g1871_p_spl_),
    .din2(g1872_p_spl_)
  );


  FA
  g_g1874_n
  (
    .dout(g1874_n),
    .din1(g1871_n_spl_),
    .din2(g1872_n_spl_)
  );


  LA
  g_g1875_p
  (
    .dout(g1875_p),
    .din1(g1873_n_spl_),
    .din2(g1874_n)
  );


  FA
  g_g1875_n
  (
    .dout(g1875_n),
    .din1(g1873_p_spl_),
    .din2(g1874_p)
  );


  LA
  g_g1876_p
  (
    .dout(g1876_p),
    .din1(g1870_n_spl_),
    .din2(g1875_p_spl_)
  );


  FA
  g_g1876_n
  (
    .dout(g1876_n),
    .din1(g1870_p_spl_),
    .din2(g1875_n_spl_)
  );


  LA
  g_g1877_p
  (
    .dout(g1877_p),
    .din1(g1870_p_spl_),
    .din2(g1875_n_spl_)
  );


  FA
  g_g1877_n
  (
    .dout(g1877_n),
    .din1(g1870_n_spl_),
    .din2(g1875_p_spl_)
  );


  LA
  g_g1878_p
  (
    .dout(g1878_p),
    .din1(g1876_n_spl_),
    .din2(g1877_n)
  );


  FA
  g_g1878_n
  (
    .dout(g1878_n),
    .din1(g1876_p_spl_),
    .din2(g1877_p)
  );


  LA
  g_g1879_p
  (
    .dout(g1879_p),
    .din1(g1869_n_spl_),
    .din2(g1878_p_spl_)
  );


  FA
  g_g1879_n
  (
    .dout(g1879_n),
    .din1(g1869_p_spl_),
    .din2(g1878_n_spl_)
  );


  LA
  g_g1880_p
  (
    .dout(g1880_p),
    .din1(g1869_p_spl_),
    .din2(g1878_n_spl_)
  );


  FA
  g_g1880_n
  (
    .dout(g1880_n),
    .din1(g1869_n_spl_),
    .din2(g1878_p_spl_)
  );


  LA
  g_g1881_p
  (
    .dout(g1881_p),
    .din1(g1879_n_spl_),
    .din2(g1880_n)
  );


  FA
  g_g1881_n
  (
    .dout(g1881_n),
    .din1(g1879_p_spl_),
    .din2(g1880_p)
  );


  LA
  g_g1882_p
  (
    .dout(g1882_p),
    .din1(g1868_n_spl_),
    .din2(g1881_p_spl_)
  );


  FA
  g_g1882_n
  (
    .dout(g1882_n),
    .din1(g1868_p_spl_),
    .din2(g1881_n_spl_)
  );


  LA
  g_g1883_p
  (
    .dout(g1883_p),
    .din1(g1868_p_spl_),
    .din2(g1881_n_spl_)
  );


  FA
  g_g1883_n
  (
    .dout(g1883_n),
    .din1(g1868_n_spl_),
    .din2(g1881_p_spl_)
  );


  LA
  g_g1884_p
  (
    .dout(g1884_p),
    .din1(g1882_n_spl_),
    .din2(g1883_n)
  );


  FA
  g_g1884_n
  (
    .dout(g1884_n),
    .din1(g1882_p_spl_),
    .din2(g1883_p)
  );


  LA
  g_g1885_p
  (
    .dout(g1885_p),
    .din1(g1867_n_spl_),
    .din2(g1884_p_spl_)
  );


  FA
  g_g1885_n
  (
    .dout(g1885_n),
    .din1(g1867_p_spl_),
    .din2(g1884_n_spl_)
  );


  LA
  g_g1886_p
  (
    .dout(g1886_p),
    .din1(g1867_p_spl_),
    .din2(g1884_n_spl_)
  );


  FA
  g_g1886_n
  (
    .dout(g1886_n),
    .din1(g1867_n_spl_),
    .din2(g1884_p_spl_)
  );


  LA
  g_g1887_p
  (
    .dout(g1887_p),
    .din1(g1885_n_spl_),
    .din2(g1886_n)
  );


  FA
  g_g1887_n
  (
    .dout(g1887_n),
    .din1(g1885_p_spl_),
    .din2(g1886_p)
  );


  LA
  g_g1888_p
  (
    .dout(g1888_p),
    .din1(g1866_n),
    .din2(g1887_p)
  );


  FA
  g_g1888_n
  (
    .dout(g1888_n),
    .din1(g1866_p_spl_),
    .din2(g1887_n_spl_)
  );


  LA
  g_g1889_p
  (
    .dout(g1889_p),
    .din1(g1866_p_spl_),
    .din2(g1887_n_spl_)
  );


  FA
  g_g1890_n
  (
    .dout(g1890_n),
    .din1(g1888_p_spl_),
    .din2(g1889_p)
  );


  LA
  g_g1891_p
  (
    .dout(g1891_p),
    .din1(g1885_n_spl_),
    .din2(g1888_n)
  );


  FA
  g_g1891_n
  (
    .dout(g1891_n),
    .din1(g1885_p_spl_),
    .din2(g1888_p_spl_)
  );


  LA
  g_g1892_p
  (
    .dout(g1892_p),
    .din1(g1879_n_spl_),
    .din2(g1882_n_spl_)
  );


  FA
  g_g1892_n
  (
    .dout(g1892_n),
    .din1(g1879_p_spl_),
    .din2(g1882_p_spl_)
  );


  LA
  g_g1893_p
  (
    .dout(g1893_p),
    .din1(G15_p_spl_111),
    .din2(G32_p_spl_111)
  );


  FA
  g_g1893_n
  (
    .dout(g1893_n),
    .din1(G15_n_spl_111),
    .din2(G32_n_spl_111)
  );


  LA
  g_g1894_p
  (
    .dout(g1894_p),
    .din1(G16_p_spl_111),
    .din2(G31_p_spl_111)
  );


  FA
  g_g1894_n
  (
    .dout(g1894_n),
    .din1(G16_n_spl_111),
    .din2(G31_n_spl_111)
  );


  LA
  g_g1895_p
  (
    .dout(g1895_p),
    .din1(g1873_n_spl_),
    .din2(g1876_n_spl_)
  );


  FA
  g_g1895_n
  (
    .dout(g1895_n),
    .din1(g1873_p_spl_),
    .din2(g1876_p_spl_)
  );


  LA
  g_g1896_p
  (
    .dout(g1896_p),
    .din1(g1894_n_spl_),
    .din2(g1895_n_spl_)
  );


  FA
  g_g1896_n
  (
    .dout(g1896_n),
    .din1(g1894_p_spl_),
    .din2(g1895_p_spl_)
  );


  LA
  g_g1897_p
  (
    .dout(g1897_p),
    .din1(g1894_p_spl_),
    .din2(g1895_p_spl_)
  );


  FA
  g_g1897_n
  (
    .dout(g1897_n),
    .din1(g1894_n_spl_),
    .din2(g1895_n_spl_)
  );


  LA
  g_g1898_p
  (
    .dout(g1898_p),
    .din1(g1896_n_spl_),
    .din2(g1897_n)
  );


  FA
  g_g1898_n
  (
    .dout(g1898_n),
    .din1(g1896_p_spl_),
    .din2(g1897_p)
  );


  LA
  g_g1899_p
  (
    .dout(g1899_p),
    .din1(g1893_n_spl_),
    .din2(g1898_p_spl_)
  );


  FA
  g_g1899_n
  (
    .dout(g1899_n),
    .din1(g1893_p_spl_),
    .din2(g1898_n_spl_)
  );


  LA
  g_g1900_p
  (
    .dout(g1900_p),
    .din1(g1893_p_spl_),
    .din2(g1898_n_spl_)
  );


  FA
  g_g1900_n
  (
    .dout(g1900_n),
    .din1(g1893_n_spl_),
    .din2(g1898_p_spl_)
  );


  LA
  g_g1901_p
  (
    .dout(g1901_p),
    .din1(g1899_n_spl_),
    .din2(g1900_n)
  );


  FA
  g_g1901_n
  (
    .dout(g1901_n),
    .din1(g1899_p_spl_),
    .din2(g1900_p)
  );


  LA
  g_g1902_p
  (
    .dout(g1902_p),
    .din1(g1892_n_spl_),
    .din2(g1901_p_spl_)
  );


  FA
  g_g1902_n
  (
    .dout(g1902_n),
    .din1(g1892_p_spl_),
    .din2(g1901_n_spl_)
  );


  LA
  g_g1903_p
  (
    .dout(g1903_p),
    .din1(g1892_p_spl_),
    .din2(g1901_n_spl_)
  );


  FA
  g_g1903_n
  (
    .dout(g1903_n),
    .din1(g1892_n_spl_),
    .din2(g1901_p_spl_)
  );


  LA
  g_g1904_p
  (
    .dout(g1904_p),
    .din1(g1902_n_spl_),
    .din2(g1903_n)
  );


  FA
  g_g1904_n
  (
    .dout(g1904_n),
    .din1(g1902_p_spl_),
    .din2(g1903_p)
  );


  LA
  g_g1905_p
  (
    .dout(g1905_p),
    .din1(g1891_n),
    .din2(g1904_p)
  );


  FA
  g_g1905_n
  (
    .dout(g1905_n),
    .din1(g1891_p_spl_),
    .din2(g1904_n_spl_)
  );


  LA
  g_g1906_p
  (
    .dout(g1906_p),
    .din1(g1891_p_spl_),
    .din2(g1904_n_spl_)
  );


  FA
  g_g1907_n
  (
    .dout(g1907_n),
    .din1(g1905_p_spl_),
    .din2(g1906_p)
  );


  LA
  g_g1908_p
  (
    .dout(g1908_p),
    .din1(G16_p_spl_111),
    .din2(G32_p_spl_111)
  );


  FA
  g_g1908_n
  (
    .dout(g1908_n),
    .din1(G16_n_spl_111),
    .din2(G32_n_spl_111)
  );


  LA
  g_g1909_p
  (
    .dout(g1909_p),
    .din1(g1896_n_spl_),
    .din2(g1899_n_spl_)
  );


  FA
  g_g1909_n
  (
    .dout(g1909_n),
    .din1(g1896_p_spl_),
    .din2(g1899_p_spl_)
  );


  LA
  g_g1910_p
  (
    .dout(g1910_p),
    .din1(g1908_n_spl_),
    .din2(g1909_n_spl_)
  );


  FA
  g_g1910_n
  (
    .dout(g1910_n),
    .din1(g1908_p_spl_),
    .din2(g1909_p_spl_)
  );


  LA
  g_g1911_p
  (
    .dout(g1911_p),
    .din1(g1902_n_spl_),
    .din2(g1905_n)
  );


  FA
  g_g1911_n
  (
    .dout(g1911_n),
    .din1(g1902_p_spl_),
    .din2(g1905_p_spl_)
  );


  LA
  g_g1912_p
  (
    .dout(g1912_p),
    .din1(g1908_p_spl_),
    .din2(g1909_p_spl_)
  );


  FA
  g_g1912_n
  (
    .dout(g1912_n),
    .din1(g1908_n_spl_),
    .din2(g1909_n_spl_)
  );


  LA
  g_g1913_p
  (
    .dout(g1913_p),
    .din1(g1910_n_spl_),
    .din2(g1912_n)
  );


  FA
  g_g1913_n
  (
    .dout(g1913_n),
    .din1(g1910_p),
    .din2(g1912_p)
  );


  FA
  g_g1914_n
  (
    .dout(g1914_n),
    .din1(g1911_p),
    .din2(g1913_n)
  );


  LA
  g_g1915_p
  (
    .dout(g1915_p),
    .din1(g1910_n_spl_),
    .din2(g1914_n_spl_)
  );


  FA
  g_g1916_n
  (
    .dout(g1916_n),
    .din1(g1911_n),
    .din2(g1913_p)
  );


  LA
  g_g1917_p
  (
    .dout(g1917_p),
    .din1(g1914_n_spl_),
    .din2(g1916_n)
  );


  buf

  (
    G6257_p,
    g33_p
  );


  buf

  (
    G6258_p,
    g39_p
  );


  buf

  (
    G6259_p,
    g52_n
  );


  buf

  (
    G6260_p,
    g73_n
  );


  buf

  (
    G6261_p,
    g102_n
  );


  buf

  (
    G6262_p,
    g139_n
  );


  buf

  (
    G6263_p,
    g184_n
  );


  buf

  (
    G6264_p,
    g237_n
  );


  buf

  (
    G6265_p,
    g298_n
  );


  buf

  (
    G6266_p,
    g367_n
  );


  buf

  (
    G6267_p,
    g444_n
  );


  buf

  (
    G6268_p,
    g529_n
  );


  buf

  (
    G6269_p,
    g622_n
  );


  buf

  (
    G6270_p,
    g723_n
  );


  buf

  (
    G6271_p,
    g832_n
  );


  buf

  (
    G6272_p,
    g949_n
  );


  buf

  (
    G6273_p,
    g1063_p
  );


  buf

  (
    G6274_p,
    g1175_n
  );


  buf

  (
    G6275_p,
    g1280_n
  );


  buf

  (
    G6276_p,
    g1377_n
  );


  buf

  (
    G6277_p,
    g1466_n
  );


  buf

  (
    G6278_p,
    g1547_n
  );


  buf

  (
    G6279_p,
    g1620_n
  );


  buf

  (
    G6280_p,
    g1685_n
  );


  buf

  (
    G6281_p,
    g1742_n
  );


  buf

  (
    G6282_p,
    g1791_n
  );


  buf

  (
    G6283_p,
    g1832_n
  );


  buf

  (
    G6284_p,
    g1865_n
  );


  buf

  (
    G6285_p,
    g1890_n
  );


  buf

  (
    G6286_p,
    g1907_n
  );


  buf

  (
    G6287_p,
    g1915_p
  );


  buf

  (
    G6288_n,
    g1917_p
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G1_p_spl_0,
    G1_p_spl_
  );


  buf

  (
    G1_p_spl_00,
    G1_p_spl_0
  );


  buf

  (
    G1_p_spl_000,
    G1_p_spl_00
  );


  buf

  (
    G1_p_spl_001,
    G1_p_spl_00
  );


  buf

  (
    G1_p_spl_01,
    G1_p_spl_0
  );


  buf

  (
    G1_p_spl_010,
    G1_p_spl_01
  );


  buf

  (
    G1_p_spl_011,
    G1_p_spl_01
  );


  buf

  (
    G1_p_spl_1,
    G1_p_spl_
  );


  buf

  (
    G1_p_spl_10,
    G1_p_spl_1
  );


  buf

  (
    G1_p_spl_100,
    G1_p_spl_10
  );


  buf

  (
    G1_p_spl_101,
    G1_p_spl_10
  );


  buf

  (
    G1_p_spl_11,
    G1_p_spl_1
  );


  buf

  (
    G1_p_spl_110,
    G1_p_spl_11
  );


  buf

  (
    G1_p_spl_111,
    G1_p_spl_11
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


  buf

  (
    G17_p_spl_0,
    G17_p_spl_
  );


  buf

  (
    G17_p_spl_00,
    G17_p_spl_0
  );


  buf

  (
    G17_p_spl_000,
    G17_p_spl_00
  );


  buf

  (
    G17_p_spl_001,
    G17_p_spl_00
  );


  buf

  (
    G17_p_spl_01,
    G17_p_spl_0
  );


  buf

  (
    G17_p_spl_010,
    G17_p_spl_01
  );


  buf

  (
    G17_p_spl_011,
    G17_p_spl_01
  );


  buf

  (
    G17_p_spl_1,
    G17_p_spl_
  );


  buf

  (
    G17_p_spl_10,
    G17_p_spl_1
  );


  buf

  (
    G17_p_spl_100,
    G17_p_spl_10
  );


  buf

  (
    G17_p_spl_101,
    G17_p_spl_10
  );


  buf

  (
    G17_p_spl_11,
    G17_p_spl_1
  );


  buf

  (
    G17_p_spl_110,
    G17_p_spl_11
  );


  buf

  (
    G17_p_spl_111,
    G17_p_spl_11
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G2_p_spl_0,
    G2_p_spl_
  );


  buf

  (
    G2_p_spl_00,
    G2_p_spl_0
  );


  buf

  (
    G2_p_spl_000,
    G2_p_spl_00
  );


  buf

  (
    G2_p_spl_001,
    G2_p_spl_00
  );


  buf

  (
    G2_p_spl_01,
    G2_p_spl_0
  );


  buf

  (
    G2_p_spl_010,
    G2_p_spl_01
  );


  buf

  (
    G2_p_spl_011,
    G2_p_spl_01
  );


  buf

  (
    G2_p_spl_1,
    G2_p_spl_
  );


  buf

  (
    G2_p_spl_10,
    G2_p_spl_1
  );


  buf

  (
    G2_p_spl_100,
    G2_p_spl_10
  );


  buf

  (
    G2_p_spl_101,
    G2_p_spl_10
  );


  buf

  (
    G2_p_spl_11,
    G2_p_spl_1
  );


  buf

  (
    G2_p_spl_110,
    G2_p_spl_11
  );


  buf

  (
    G2_p_spl_111,
    G2_p_spl_11
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G2_n_spl_0,
    G2_n_spl_
  );


  buf

  (
    G2_n_spl_00,
    G2_n_spl_0
  );


  buf

  (
    G2_n_spl_000,
    G2_n_spl_00
  );


  buf

  (
    G2_n_spl_001,
    G2_n_spl_00
  );


  buf

  (
    G2_n_spl_01,
    G2_n_spl_0
  );


  buf

  (
    G2_n_spl_010,
    G2_n_spl_01
  );


  buf

  (
    G2_n_spl_011,
    G2_n_spl_01
  );


  buf

  (
    G2_n_spl_1,
    G2_n_spl_
  );


  buf

  (
    G2_n_spl_10,
    G2_n_spl_1
  );


  buf

  (
    G2_n_spl_100,
    G2_n_spl_10
  );


  buf

  (
    G2_n_spl_101,
    G2_n_spl_10
  );


  buf

  (
    G2_n_spl_11,
    G2_n_spl_1
  );


  buf

  (
    G2_n_spl_110,
    G2_n_spl_11
  );


  buf

  (
    G2_n_spl_111,
    G2_n_spl_11
  );


  buf

  (
    G17_n_spl_,
    G17_n
  );


  buf

  (
    G17_n_spl_0,
    G17_n_spl_
  );


  buf

  (
    G17_n_spl_00,
    G17_n_spl_0
  );


  buf

  (
    G17_n_spl_000,
    G17_n_spl_00
  );


  buf

  (
    G17_n_spl_001,
    G17_n_spl_00
  );


  buf

  (
    G17_n_spl_01,
    G17_n_spl_0
  );


  buf

  (
    G17_n_spl_010,
    G17_n_spl_01
  );


  buf

  (
    G17_n_spl_011,
    G17_n_spl_01
  );


  buf

  (
    G17_n_spl_1,
    G17_n_spl_
  );


  buf

  (
    G17_n_spl_10,
    G17_n_spl_1
  );


  buf

  (
    G17_n_spl_100,
    G17_n_spl_10
  );


  buf

  (
    G17_n_spl_101,
    G17_n_spl_10
  );


  buf

  (
    G17_n_spl_11,
    G17_n_spl_1
  );


  buf

  (
    G17_n_spl_110,
    G17_n_spl_11
  );


  buf

  (
    G18_p_spl_,
    G18_p
  );


  buf

  (
    G18_p_spl_0,
    G18_p_spl_
  );


  buf

  (
    G18_p_spl_00,
    G18_p_spl_0
  );


  buf

  (
    G18_p_spl_000,
    G18_p_spl_00
  );


  buf

  (
    G18_p_spl_001,
    G18_p_spl_00
  );


  buf

  (
    G18_p_spl_01,
    G18_p_spl_0
  );


  buf

  (
    G18_p_spl_010,
    G18_p_spl_01
  );


  buf

  (
    G18_p_spl_011,
    G18_p_spl_01
  );


  buf

  (
    G18_p_spl_1,
    G18_p_spl_
  );


  buf

  (
    G18_p_spl_10,
    G18_p_spl_1
  );


  buf

  (
    G18_p_spl_100,
    G18_p_spl_10
  );


  buf

  (
    G18_p_spl_101,
    G18_p_spl_10
  );


  buf

  (
    G18_p_spl_11,
    G18_p_spl_1
  );


  buf

  (
    G18_p_spl_110,
    G18_p_spl_11
  );


  buf

  (
    G18_p_spl_111,
    G18_p_spl_11
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G1_n_spl_0,
    G1_n_spl_
  );


  buf

  (
    G1_n_spl_00,
    G1_n_spl_0
  );


  buf

  (
    G1_n_spl_000,
    G1_n_spl_00
  );


  buf

  (
    G1_n_spl_001,
    G1_n_spl_00
  );


  buf

  (
    G1_n_spl_01,
    G1_n_spl_0
  );


  buf

  (
    G1_n_spl_010,
    G1_n_spl_01
  );


  buf

  (
    G1_n_spl_011,
    G1_n_spl_01
  );


  buf

  (
    G1_n_spl_1,
    G1_n_spl_
  );


  buf

  (
    G1_n_spl_10,
    G1_n_spl_1
  );


  buf

  (
    G1_n_spl_100,
    G1_n_spl_10
  );


  buf

  (
    G1_n_spl_101,
    G1_n_spl_10
  );


  buf

  (
    G1_n_spl_11,
    G1_n_spl_1
  );


  buf

  (
    G1_n_spl_110,
    G1_n_spl_11
  );


  buf

  (
    G18_n_spl_,
    G18_n
  );


  buf

  (
    G18_n_spl_0,
    G18_n_spl_
  );


  buf

  (
    G18_n_spl_00,
    G18_n_spl_0
  );


  buf

  (
    G18_n_spl_000,
    G18_n_spl_00
  );


  buf

  (
    G18_n_spl_001,
    G18_n_spl_00
  );


  buf

  (
    G18_n_spl_01,
    G18_n_spl_0
  );


  buf

  (
    G18_n_spl_010,
    G18_n_spl_01
  );


  buf

  (
    G18_n_spl_011,
    G18_n_spl_01
  );


  buf

  (
    G18_n_spl_1,
    G18_n_spl_
  );


  buf

  (
    G18_n_spl_10,
    G18_n_spl_1
  );


  buf

  (
    G18_n_spl_100,
    G18_n_spl_10
  );


  buf

  (
    G18_n_spl_101,
    G18_n_spl_10
  );


  buf

  (
    G18_n_spl_11,
    G18_n_spl_1
  );


  buf

  (
    G18_n_spl_110,
    G18_n_spl_11
  );


  buf

  (
    G18_n_spl_111,
    G18_n_spl_11
  );


  buf

  (
    g34_p_spl_,
    g34_p
  );


  buf

  (
    g34_n_spl_,
    g34_n
  );


  buf

  (
    g35_p_spl_,
    g35_p
  );


  buf

  (
    g36_p_spl_,
    g36_p
  );


  buf

  (
    g37_n_spl_,
    g37_n
  );


  buf

  (
    g37_n_spl_0,
    g37_n_spl_
  );


  buf

  (
    G19_p_spl_,
    G19_p
  );


  buf

  (
    G19_p_spl_0,
    G19_p_spl_
  );


  buf

  (
    G19_p_spl_00,
    G19_p_spl_0
  );


  buf

  (
    G19_p_spl_000,
    G19_p_spl_00
  );


  buf

  (
    G19_p_spl_001,
    G19_p_spl_00
  );


  buf

  (
    G19_p_spl_01,
    G19_p_spl_0
  );


  buf

  (
    G19_p_spl_010,
    G19_p_spl_01
  );


  buf

  (
    G19_p_spl_011,
    G19_p_spl_01
  );


  buf

  (
    G19_p_spl_1,
    G19_p_spl_
  );


  buf

  (
    G19_p_spl_10,
    G19_p_spl_1
  );


  buf

  (
    G19_p_spl_100,
    G19_p_spl_10
  );


  buf

  (
    G19_p_spl_101,
    G19_p_spl_10
  );


  buf

  (
    G19_p_spl_11,
    G19_p_spl_1
  );


  buf

  (
    G19_p_spl_110,
    G19_p_spl_11
  );


  buf

  (
    G19_p_spl_111,
    G19_p_spl_11
  );


  buf

  (
    G19_n_spl_,
    G19_n
  );


  buf

  (
    G19_n_spl_0,
    G19_n_spl_
  );


  buf

  (
    G19_n_spl_00,
    G19_n_spl_0
  );


  buf

  (
    G19_n_spl_000,
    G19_n_spl_00
  );


  buf

  (
    G19_n_spl_001,
    G19_n_spl_00
  );


  buf

  (
    G19_n_spl_01,
    G19_n_spl_0
  );


  buf

  (
    G19_n_spl_010,
    G19_n_spl_01
  );


  buf

  (
    G19_n_spl_011,
    G19_n_spl_01
  );


  buf

  (
    G19_n_spl_1,
    G19_n_spl_
  );


  buf

  (
    G19_n_spl_10,
    G19_n_spl_1
  );


  buf

  (
    G19_n_spl_100,
    G19_n_spl_10
  );


  buf

  (
    G19_n_spl_101,
    G19_n_spl_10
  );


  buf

  (
    G19_n_spl_11,
    G19_n_spl_1
  );


  buf

  (
    G19_n_spl_110,
    G19_n_spl_11
  );


  buf

  (
    G19_n_spl_111,
    G19_n_spl_11
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G3_p_spl_0,
    G3_p_spl_
  );


  buf

  (
    G3_p_spl_00,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_000,
    G3_p_spl_00
  );


  buf

  (
    G3_p_spl_001,
    G3_p_spl_00
  );


  buf

  (
    G3_p_spl_01,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_010,
    G3_p_spl_01
  );


  buf

  (
    G3_p_spl_011,
    G3_p_spl_01
  );


  buf

  (
    G3_p_spl_1,
    G3_p_spl_
  );


  buf

  (
    G3_p_spl_10,
    G3_p_spl_1
  );


  buf

  (
    G3_p_spl_100,
    G3_p_spl_10
  );


  buf

  (
    G3_p_spl_101,
    G3_p_spl_10
  );


  buf

  (
    G3_p_spl_11,
    G3_p_spl_1
  );


  buf

  (
    G3_p_spl_110,
    G3_p_spl_11
  );


  buf

  (
    G3_p_spl_111,
    G3_p_spl_11
  );


  buf

  (
    G3_n_spl_,
    G3_n
  );


  buf

  (
    G3_n_spl_0,
    G3_n_spl_
  );


  buf

  (
    G3_n_spl_00,
    G3_n_spl_0
  );


  buf

  (
    G3_n_spl_000,
    G3_n_spl_00
  );


  buf

  (
    G3_n_spl_001,
    G3_n_spl_00
  );


  buf

  (
    G3_n_spl_01,
    G3_n_spl_0
  );


  buf

  (
    G3_n_spl_010,
    G3_n_spl_01
  );


  buf

  (
    G3_n_spl_011,
    G3_n_spl_01
  );


  buf

  (
    G3_n_spl_1,
    G3_n_spl_
  );


  buf

  (
    G3_n_spl_10,
    G3_n_spl_1
  );


  buf

  (
    G3_n_spl_100,
    G3_n_spl_10
  );


  buf

  (
    G3_n_spl_101,
    G3_n_spl_10
  );


  buf

  (
    G3_n_spl_11,
    G3_n_spl_1
  );


  buf

  (
    G3_n_spl_110,
    G3_n_spl_11
  );


  buf

  (
    G3_n_spl_111,
    G3_n_spl_11
  );


  buf

  (
    g41_p_spl_,
    g41_p
  );


  buf

  (
    g42_n_spl_,
    g42_n
  );


  buf

  (
    g41_n_spl_,
    g41_n
  );


  buf

  (
    g42_p_spl_,
    g42_p
  );


  buf

  (
    g43_n_spl_,
    g43_n
  );


  buf

  (
    g43_p_spl_,
    g43_p
  );


  buf

  (
    g44_n_spl_,
    g44_n
  );


  buf

  (
    g44_n_spl_0,
    g44_n_spl_
  );


  buf

  (
    g44_p_spl_,
    g44_p
  );


  buf

  (
    g44_p_spl_0,
    g44_p_spl_
  );


  buf

  (
    g46_n_spl_,
    g46_n
  );


  buf

  (
    g37_p_spl_,
    g37_p
  );


  buf

  (
    g46_p_spl_,
    g46_p
  );


  buf

  (
    g47_n_spl_,
    g47_n
  );


  buf

  (
    g47_p_spl_,
    g47_p
  );


  buf

  (
    g40_p_spl_,
    g40_p
  );


  buf

  (
    g49_n_spl_,
    g49_n
  );


  buf

  (
    g50_p_spl_,
    g50_p
  );


  buf

  (
    G20_p_spl_,
    G20_p
  );


  buf

  (
    G20_p_spl_0,
    G20_p_spl_
  );


  buf

  (
    G20_p_spl_00,
    G20_p_spl_0
  );


  buf

  (
    G20_p_spl_000,
    G20_p_spl_00
  );


  buf

  (
    G20_p_spl_001,
    G20_p_spl_00
  );


  buf

  (
    G20_p_spl_01,
    G20_p_spl_0
  );


  buf

  (
    G20_p_spl_010,
    G20_p_spl_01
  );


  buf

  (
    G20_p_spl_011,
    G20_p_spl_01
  );


  buf

  (
    G20_p_spl_1,
    G20_p_spl_
  );


  buf

  (
    G20_p_spl_10,
    G20_p_spl_1
  );


  buf

  (
    G20_p_spl_100,
    G20_p_spl_10
  );


  buf

  (
    G20_p_spl_101,
    G20_p_spl_10
  );


  buf

  (
    G20_p_spl_11,
    G20_p_spl_1
  );


  buf

  (
    G20_p_spl_110,
    G20_p_spl_11
  );


  buf

  (
    G20_p_spl_111,
    G20_p_spl_11
  );


  buf

  (
    G20_n_spl_,
    G20_n
  );


  buf

  (
    G20_n_spl_0,
    G20_n_spl_
  );


  buf

  (
    G20_n_spl_00,
    G20_n_spl_0
  );


  buf

  (
    G20_n_spl_000,
    G20_n_spl_00
  );


  buf

  (
    G20_n_spl_001,
    G20_n_spl_00
  );


  buf

  (
    G20_n_spl_01,
    G20_n_spl_0
  );


  buf

  (
    G20_n_spl_010,
    G20_n_spl_01
  );


  buf

  (
    G20_n_spl_011,
    G20_n_spl_01
  );


  buf

  (
    G20_n_spl_1,
    G20_n_spl_
  );


  buf

  (
    G20_n_spl_10,
    G20_n_spl_1
  );


  buf

  (
    G20_n_spl_100,
    G20_n_spl_10
  );


  buf

  (
    G20_n_spl_101,
    G20_n_spl_10
  );


  buf

  (
    G20_n_spl_11,
    G20_n_spl_1
  );


  buf

  (
    G20_n_spl_110,
    G20_n_spl_11
  );


  buf

  (
    G20_n_spl_111,
    G20_n_spl_11
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_00,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_000,
    G4_p_spl_00
  );


  buf

  (
    G4_p_spl_001,
    G4_p_spl_00
  );


  buf

  (
    G4_p_spl_01,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_010,
    G4_p_spl_01
  );


  buf

  (
    G4_p_spl_011,
    G4_p_spl_01
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_10,
    G4_p_spl_1
  );


  buf

  (
    G4_p_spl_100,
    G4_p_spl_10
  );


  buf

  (
    G4_p_spl_101,
    G4_p_spl_10
  );


  buf

  (
    G4_p_spl_11,
    G4_p_spl_1
  );


  buf

  (
    G4_p_spl_110,
    G4_p_spl_11
  );


  buf

  (
    G4_p_spl_111,
    G4_p_spl_11
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    G4_n_spl_0,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_00,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_000,
    G4_n_spl_00
  );


  buf

  (
    G4_n_spl_001,
    G4_n_spl_00
  );


  buf

  (
    G4_n_spl_01,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_010,
    G4_n_spl_01
  );


  buf

  (
    G4_n_spl_011,
    G4_n_spl_01
  );


  buf

  (
    G4_n_spl_1,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_10,
    G4_n_spl_1
  );


  buf

  (
    G4_n_spl_100,
    G4_n_spl_10
  );


  buf

  (
    G4_n_spl_101,
    G4_n_spl_10
  );


  buf

  (
    G4_n_spl_11,
    G4_n_spl_1
  );


  buf

  (
    G4_n_spl_110,
    G4_n_spl_11
  );


  buf

  (
    G4_n_spl_111,
    G4_n_spl_11
  );


  buf

  (
    g56_p_spl_,
    g56_p
  );


  buf

  (
    g57_n_spl_,
    g57_n
  );


  buf

  (
    g56_n_spl_,
    g56_n
  );


  buf

  (
    g57_p_spl_,
    g57_p
  );


  buf

  (
    g58_n_spl_,
    g58_n
  );


  buf

  (
    g58_p_spl_,
    g58_p
  );


  buf

  (
    g59_n_spl_,
    g59_n
  );


  buf

  (
    g59_n_spl_0,
    g59_n_spl_
  );


  buf

  (
    g59_p_spl_,
    g59_p
  );


  buf

  (
    g59_p_spl_0,
    g59_p_spl_
  );


  buf

  (
    g61_n_spl_,
    g61_n
  );


  buf

  (
    g61_p_spl_,
    g61_p
  );


  buf

  (
    g62_n_spl_,
    g62_n
  );


  buf

  (
    g62_p_spl_,
    g62_p
  );


  buf

  (
    g55_n_spl_,
    g55_n
  );


  buf

  (
    g64_p_spl_,
    g64_p
  );


  buf

  (
    g55_p_spl_,
    g55_p
  );


  buf

  (
    g64_n_spl_,
    g64_n
  );


  buf

  (
    g65_n_spl_,
    g65_n
  );


  buf

  (
    g65_p_spl_,
    g65_p
  );


  buf

  (
    g54_n_spl_,
    g54_n
  );


  buf

  (
    g67_p_spl_,
    g67_p
  );


  buf

  (
    g54_p_spl_,
    g54_p
  );


  buf

  (
    g67_n_spl_,
    g67_n
  );


  buf

  (
    g68_n_spl_,
    g68_n
  );


  buf

  (
    g68_p_spl_,
    g68_p
  );


  buf

  (
    g53_p_spl_,
    g53_p
  );


  buf

  (
    g70_n_spl_,
    g70_n
  );


  buf

  (
    g71_p_spl_,
    g71_p
  );


  buf

  (
    G21_p_spl_,
    G21_p
  );


  buf

  (
    G21_p_spl_0,
    G21_p_spl_
  );


  buf

  (
    G21_p_spl_00,
    G21_p_spl_0
  );


  buf

  (
    G21_p_spl_000,
    G21_p_spl_00
  );


  buf

  (
    G21_p_spl_001,
    G21_p_spl_00
  );


  buf

  (
    G21_p_spl_01,
    G21_p_spl_0
  );


  buf

  (
    G21_p_spl_010,
    G21_p_spl_01
  );


  buf

  (
    G21_p_spl_011,
    G21_p_spl_01
  );


  buf

  (
    G21_p_spl_1,
    G21_p_spl_
  );


  buf

  (
    G21_p_spl_10,
    G21_p_spl_1
  );


  buf

  (
    G21_p_spl_100,
    G21_p_spl_10
  );


  buf

  (
    G21_p_spl_101,
    G21_p_spl_10
  );


  buf

  (
    G21_p_spl_11,
    G21_p_spl_1
  );


  buf

  (
    G21_p_spl_110,
    G21_p_spl_11
  );


  buf

  (
    G21_p_spl_111,
    G21_p_spl_11
  );


  buf

  (
    G21_n_spl_,
    G21_n
  );


  buf

  (
    G21_n_spl_0,
    G21_n_spl_
  );


  buf

  (
    G21_n_spl_00,
    G21_n_spl_0
  );


  buf

  (
    G21_n_spl_000,
    G21_n_spl_00
  );


  buf

  (
    G21_n_spl_001,
    G21_n_spl_00
  );


  buf

  (
    G21_n_spl_01,
    G21_n_spl_0
  );


  buf

  (
    G21_n_spl_010,
    G21_n_spl_01
  );


  buf

  (
    G21_n_spl_011,
    G21_n_spl_01
  );


  buf

  (
    G21_n_spl_1,
    G21_n_spl_
  );


  buf

  (
    G21_n_spl_10,
    G21_n_spl_1
  );


  buf

  (
    G21_n_spl_100,
    G21_n_spl_10
  );


  buf

  (
    G21_n_spl_101,
    G21_n_spl_10
  );


  buf

  (
    G21_n_spl_11,
    G21_n_spl_1
  );


  buf

  (
    G21_n_spl_110,
    G21_n_spl_11
  );


  buf

  (
    G21_n_spl_111,
    G21_n_spl_11
  );


  buf

  (
    G5_p_spl_,
    G5_p
  );


  buf

  (
    G5_p_spl_0,
    G5_p_spl_
  );


  buf

  (
    G5_p_spl_00,
    G5_p_spl_0
  );


  buf

  (
    G5_p_spl_000,
    G5_p_spl_00
  );


  buf

  (
    G5_p_spl_001,
    G5_p_spl_00
  );


  buf

  (
    G5_p_spl_01,
    G5_p_spl_0
  );


  buf

  (
    G5_p_spl_010,
    G5_p_spl_01
  );


  buf

  (
    G5_p_spl_011,
    G5_p_spl_01
  );


  buf

  (
    G5_p_spl_1,
    G5_p_spl_
  );


  buf

  (
    G5_p_spl_10,
    G5_p_spl_1
  );


  buf

  (
    G5_p_spl_100,
    G5_p_spl_10
  );


  buf

  (
    G5_p_spl_101,
    G5_p_spl_10
  );


  buf

  (
    G5_p_spl_11,
    G5_p_spl_1
  );


  buf

  (
    G5_p_spl_110,
    G5_p_spl_11
  );


  buf

  (
    G5_p_spl_111,
    G5_p_spl_11
  );


  buf

  (
    G5_n_spl_,
    G5_n
  );


  buf

  (
    G5_n_spl_0,
    G5_n_spl_
  );


  buf

  (
    G5_n_spl_00,
    G5_n_spl_0
  );


  buf

  (
    G5_n_spl_000,
    G5_n_spl_00
  );


  buf

  (
    G5_n_spl_001,
    G5_n_spl_00
  );


  buf

  (
    G5_n_spl_01,
    G5_n_spl_0
  );


  buf

  (
    G5_n_spl_010,
    G5_n_spl_01
  );


  buf

  (
    G5_n_spl_011,
    G5_n_spl_01
  );


  buf

  (
    G5_n_spl_1,
    G5_n_spl_
  );


  buf

  (
    G5_n_spl_10,
    G5_n_spl_1
  );


  buf

  (
    G5_n_spl_100,
    G5_n_spl_10
  );


  buf

  (
    G5_n_spl_101,
    G5_n_spl_10
  );


  buf

  (
    G5_n_spl_11,
    G5_n_spl_1
  );


  buf

  (
    G5_n_spl_110,
    G5_n_spl_11
  );


  buf

  (
    G5_n_spl_111,
    G5_n_spl_11
  );


  buf

  (
    g79_p_spl_,
    g79_p
  );


  buf

  (
    g80_n_spl_,
    g80_n
  );


  buf

  (
    g79_n_spl_,
    g79_n
  );


  buf

  (
    g80_p_spl_,
    g80_p
  );


  buf

  (
    g81_n_spl_,
    g81_n
  );


  buf

  (
    g81_p_spl_,
    g81_p
  );


  buf

  (
    g82_n_spl_,
    g82_n
  );


  buf

  (
    g82_n_spl_0,
    g82_n_spl_
  );


  buf

  (
    g82_p_spl_,
    g82_p
  );


  buf

  (
    g82_p_spl_0,
    g82_p_spl_
  );


  buf

  (
    g84_n_spl_,
    g84_n
  );


  buf

  (
    g84_p_spl_,
    g84_p
  );


  buf

  (
    g85_n_spl_,
    g85_n
  );


  buf

  (
    g85_p_spl_,
    g85_p
  );


  buf

  (
    g78_n_spl_,
    g78_n
  );


  buf

  (
    g87_p_spl_,
    g87_p
  );


  buf

  (
    g78_p_spl_,
    g78_p
  );


  buf

  (
    g87_n_spl_,
    g87_n
  );


  buf

  (
    g88_n_spl_,
    g88_n
  );


  buf

  (
    g88_p_spl_,
    g88_p
  );


  buf

  (
    g77_n_spl_,
    g77_n
  );


  buf

  (
    g90_p_spl_,
    g90_p
  );


  buf

  (
    g77_p_spl_,
    g77_p
  );


  buf

  (
    g90_n_spl_,
    g90_n
  );


  buf

  (
    g91_n_spl_,
    g91_n
  );


  buf

  (
    g91_p_spl_,
    g91_p
  );


  buf

  (
    g76_n_spl_,
    g76_n
  );


  buf

  (
    g93_p_spl_,
    g93_p
  );


  buf

  (
    g76_p_spl_,
    g76_p
  );


  buf

  (
    g93_n_spl_,
    g93_n
  );


  buf

  (
    g94_n_spl_,
    g94_n
  );


  buf

  (
    g94_p_spl_,
    g94_p
  );


  buf

  (
    g75_n_spl_,
    g75_n
  );


  buf

  (
    g96_p_spl_,
    g96_p
  );


  buf

  (
    g75_p_spl_,
    g75_p
  );


  buf

  (
    g96_n_spl_,
    g96_n
  );


  buf

  (
    g97_n_spl_,
    g97_n
  );


  buf

  (
    g97_p_spl_,
    g97_p
  );


  buf

  (
    g74_p_spl_,
    g74_p
  );


  buf

  (
    g99_n_spl_,
    g99_n
  );


  buf

  (
    g100_p_spl_,
    g100_p
  );


  buf

  (
    G22_p_spl_,
    G22_p
  );


  buf

  (
    G22_p_spl_0,
    G22_p_spl_
  );


  buf

  (
    G22_p_spl_00,
    G22_p_spl_0
  );


  buf

  (
    G22_p_spl_000,
    G22_p_spl_00
  );


  buf

  (
    G22_p_spl_001,
    G22_p_spl_00
  );


  buf

  (
    G22_p_spl_01,
    G22_p_spl_0
  );


  buf

  (
    G22_p_spl_010,
    G22_p_spl_01
  );


  buf

  (
    G22_p_spl_011,
    G22_p_spl_01
  );


  buf

  (
    G22_p_spl_1,
    G22_p_spl_
  );


  buf

  (
    G22_p_spl_10,
    G22_p_spl_1
  );


  buf

  (
    G22_p_spl_100,
    G22_p_spl_10
  );


  buf

  (
    G22_p_spl_101,
    G22_p_spl_10
  );


  buf

  (
    G22_p_spl_11,
    G22_p_spl_1
  );


  buf

  (
    G22_p_spl_110,
    G22_p_spl_11
  );


  buf

  (
    G22_p_spl_111,
    G22_p_spl_11
  );


  buf

  (
    G22_n_spl_,
    G22_n
  );


  buf

  (
    G22_n_spl_0,
    G22_n_spl_
  );


  buf

  (
    G22_n_spl_00,
    G22_n_spl_0
  );


  buf

  (
    G22_n_spl_000,
    G22_n_spl_00
  );


  buf

  (
    G22_n_spl_001,
    G22_n_spl_00
  );


  buf

  (
    G22_n_spl_01,
    G22_n_spl_0
  );


  buf

  (
    G22_n_spl_010,
    G22_n_spl_01
  );


  buf

  (
    G22_n_spl_011,
    G22_n_spl_01
  );


  buf

  (
    G22_n_spl_1,
    G22_n_spl_
  );


  buf

  (
    G22_n_spl_10,
    G22_n_spl_1
  );


  buf

  (
    G22_n_spl_100,
    G22_n_spl_10
  );


  buf

  (
    G22_n_spl_101,
    G22_n_spl_10
  );


  buf

  (
    G22_n_spl_11,
    G22_n_spl_1
  );


  buf

  (
    G22_n_spl_110,
    G22_n_spl_11
  );


  buf

  (
    G22_n_spl_111,
    G22_n_spl_11
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G6_p_spl_0,
    G6_p_spl_
  );


  buf

  (
    G6_p_spl_00,
    G6_p_spl_0
  );


  buf

  (
    G6_p_spl_000,
    G6_p_spl_00
  );


  buf

  (
    G6_p_spl_001,
    G6_p_spl_00
  );


  buf

  (
    G6_p_spl_01,
    G6_p_spl_0
  );


  buf

  (
    G6_p_spl_010,
    G6_p_spl_01
  );


  buf

  (
    G6_p_spl_011,
    G6_p_spl_01
  );


  buf

  (
    G6_p_spl_1,
    G6_p_spl_
  );


  buf

  (
    G6_p_spl_10,
    G6_p_spl_1
  );


  buf

  (
    G6_p_spl_100,
    G6_p_spl_10
  );


  buf

  (
    G6_p_spl_101,
    G6_p_spl_10
  );


  buf

  (
    G6_p_spl_11,
    G6_p_spl_1
  );


  buf

  (
    G6_p_spl_110,
    G6_p_spl_11
  );


  buf

  (
    G6_p_spl_111,
    G6_p_spl_11
  );


  buf

  (
    G6_n_spl_,
    G6_n
  );


  buf

  (
    G6_n_spl_0,
    G6_n_spl_
  );


  buf

  (
    G6_n_spl_00,
    G6_n_spl_0
  );


  buf

  (
    G6_n_spl_000,
    G6_n_spl_00
  );


  buf

  (
    G6_n_spl_001,
    G6_n_spl_00
  );


  buf

  (
    G6_n_spl_01,
    G6_n_spl_0
  );


  buf

  (
    G6_n_spl_010,
    G6_n_spl_01
  );


  buf

  (
    G6_n_spl_011,
    G6_n_spl_01
  );


  buf

  (
    G6_n_spl_1,
    G6_n_spl_
  );


  buf

  (
    G6_n_spl_10,
    G6_n_spl_1
  );


  buf

  (
    G6_n_spl_100,
    G6_n_spl_10
  );


  buf

  (
    G6_n_spl_101,
    G6_n_spl_10
  );


  buf

  (
    G6_n_spl_11,
    G6_n_spl_1
  );


  buf

  (
    G6_n_spl_110,
    G6_n_spl_11
  );


  buf

  (
    G6_n_spl_111,
    G6_n_spl_11
  );


  buf

  (
    g110_p_spl_,
    g110_p
  );


  buf

  (
    g111_n_spl_,
    g111_n
  );


  buf

  (
    g110_n_spl_,
    g110_n
  );


  buf

  (
    g111_p_spl_,
    g111_p
  );


  buf

  (
    g112_n_spl_,
    g112_n
  );


  buf

  (
    g112_p_spl_,
    g112_p
  );


  buf

  (
    g113_n_spl_,
    g113_n
  );


  buf

  (
    g113_n_spl_0,
    g113_n_spl_
  );


  buf

  (
    g113_p_spl_,
    g113_p
  );


  buf

  (
    g113_p_spl_0,
    g113_p_spl_
  );


  buf

  (
    g115_n_spl_,
    g115_n
  );


  buf

  (
    g115_p_spl_,
    g115_p
  );


  buf

  (
    g116_n_spl_,
    g116_n
  );


  buf

  (
    g116_p_spl_,
    g116_p
  );


  buf

  (
    g109_n_spl_,
    g109_n
  );


  buf

  (
    g118_p_spl_,
    g118_p
  );


  buf

  (
    g109_p_spl_,
    g109_p
  );


  buf

  (
    g118_n_spl_,
    g118_n
  );


  buf

  (
    g119_n_spl_,
    g119_n
  );


  buf

  (
    g119_p_spl_,
    g119_p
  );


  buf

  (
    g108_n_spl_,
    g108_n
  );


  buf

  (
    g121_p_spl_,
    g121_p
  );


  buf

  (
    g108_p_spl_,
    g108_p
  );


  buf

  (
    g121_n_spl_,
    g121_n
  );


  buf

  (
    g122_n_spl_,
    g122_n
  );


  buf

  (
    g122_p_spl_,
    g122_p
  );


  buf

  (
    g107_n_spl_,
    g107_n
  );


  buf

  (
    g124_p_spl_,
    g124_p
  );


  buf

  (
    g107_p_spl_,
    g107_p
  );


  buf

  (
    g124_n_spl_,
    g124_n
  );


  buf

  (
    g125_n_spl_,
    g125_n
  );


  buf

  (
    g125_p_spl_,
    g125_p
  );


  buf

  (
    g106_n_spl_,
    g106_n
  );


  buf

  (
    g127_p_spl_,
    g127_p
  );


  buf

  (
    g106_p_spl_,
    g106_p
  );


  buf

  (
    g127_n_spl_,
    g127_n
  );


  buf

  (
    g128_n_spl_,
    g128_n
  );


  buf

  (
    g128_p_spl_,
    g128_p
  );


  buf

  (
    g105_n_spl_,
    g105_n
  );


  buf

  (
    g130_p_spl_,
    g130_p
  );


  buf

  (
    g105_p_spl_,
    g105_p
  );


  buf

  (
    g130_n_spl_,
    g130_n
  );


  buf

  (
    g131_n_spl_,
    g131_n
  );


  buf

  (
    g131_p_spl_,
    g131_p
  );


  buf

  (
    g104_n_spl_,
    g104_n
  );


  buf

  (
    g133_p_spl_,
    g133_p
  );


  buf

  (
    g104_p_spl_,
    g104_p
  );


  buf

  (
    g133_n_spl_,
    g133_n
  );


  buf

  (
    g134_n_spl_,
    g134_n
  );


  buf

  (
    g134_p_spl_,
    g134_p
  );


  buf

  (
    g103_p_spl_,
    g103_p
  );


  buf

  (
    g136_n_spl_,
    g136_n
  );


  buf

  (
    g137_p_spl_,
    g137_p
  );


  buf

  (
    G23_p_spl_,
    G23_p
  );


  buf

  (
    G23_p_spl_0,
    G23_p_spl_
  );


  buf

  (
    G23_p_spl_00,
    G23_p_spl_0
  );


  buf

  (
    G23_p_spl_000,
    G23_p_spl_00
  );


  buf

  (
    G23_p_spl_001,
    G23_p_spl_00
  );


  buf

  (
    G23_p_spl_01,
    G23_p_spl_0
  );


  buf

  (
    G23_p_spl_010,
    G23_p_spl_01
  );


  buf

  (
    G23_p_spl_011,
    G23_p_spl_01
  );


  buf

  (
    G23_p_spl_1,
    G23_p_spl_
  );


  buf

  (
    G23_p_spl_10,
    G23_p_spl_1
  );


  buf

  (
    G23_p_spl_100,
    G23_p_spl_10
  );


  buf

  (
    G23_p_spl_101,
    G23_p_spl_10
  );


  buf

  (
    G23_p_spl_11,
    G23_p_spl_1
  );


  buf

  (
    G23_p_spl_110,
    G23_p_spl_11
  );


  buf

  (
    G23_p_spl_111,
    G23_p_spl_11
  );


  buf

  (
    G23_n_spl_,
    G23_n
  );


  buf

  (
    G23_n_spl_0,
    G23_n_spl_
  );


  buf

  (
    G23_n_spl_00,
    G23_n_spl_0
  );


  buf

  (
    G23_n_spl_000,
    G23_n_spl_00
  );


  buf

  (
    G23_n_spl_001,
    G23_n_spl_00
  );


  buf

  (
    G23_n_spl_01,
    G23_n_spl_0
  );


  buf

  (
    G23_n_spl_010,
    G23_n_spl_01
  );


  buf

  (
    G23_n_spl_011,
    G23_n_spl_01
  );


  buf

  (
    G23_n_spl_1,
    G23_n_spl_
  );


  buf

  (
    G23_n_spl_10,
    G23_n_spl_1
  );


  buf

  (
    G23_n_spl_100,
    G23_n_spl_10
  );


  buf

  (
    G23_n_spl_101,
    G23_n_spl_10
  );


  buf

  (
    G23_n_spl_11,
    G23_n_spl_1
  );


  buf

  (
    G23_n_spl_110,
    G23_n_spl_11
  );


  buf

  (
    G23_n_spl_111,
    G23_n_spl_11
  );


  buf

  (
    G7_p_spl_,
    G7_p
  );


  buf

  (
    G7_p_spl_0,
    G7_p_spl_
  );


  buf

  (
    G7_p_spl_00,
    G7_p_spl_0
  );


  buf

  (
    G7_p_spl_000,
    G7_p_spl_00
  );


  buf

  (
    G7_p_spl_001,
    G7_p_spl_00
  );


  buf

  (
    G7_p_spl_01,
    G7_p_spl_0
  );


  buf

  (
    G7_p_spl_010,
    G7_p_spl_01
  );


  buf

  (
    G7_p_spl_011,
    G7_p_spl_01
  );


  buf

  (
    G7_p_spl_1,
    G7_p_spl_
  );


  buf

  (
    G7_p_spl_10,
    G7_p_spl_1
  );


  buf

  (
    G7_p_spl_100,
    G7_p_spl_10
  );


  buf

  (
    G7_p_spl_101,
    G7_p_spl_10
  );


  buf

  (
    G7_p_spl_11,
    G7_p_spl_1
  );


  buf

  (
    G7_p_spl_110,
    G7_p_spl_11
  );


  buf

  (
    G7_p_spl_111,
    G7_p_spl_11
  );


  buf

  (
    G7_n_spl_,
    G7_n
  );


  buf

  (
    G7_n_spl_0,
    G7_n_spl_
  );


  buf

  (
    G7_n_spl_00,
    G7_n_spl_0
  );


  buf

  (
    G7_n_spl_000,
    G7_n_spl_00
  );


  buf

  (
    G7_n_spl_001,
    G7_n_spl_00
  );


  buf

  (
    G7_n_spl_01,
    G7_n_spl_0
  );


  buf

  (
    G7_n_spl_010,
    G7_n_spl_01
  );


  buf

  (
    G7_n_spl_011,
    G7_n_spl_01
  );


  buf

  (
    G7_n_spl_1,
    G7_n_spl_
  );


  buf

  (
    G7_n_spl_10,
    G7_n_spl_1
  );


  buf

  (
    G7_n_spl_100,
    G7_n_spl_10
  );


  buf

  (
    G7_n_spl_101,
    G7_n_spl_10
  );


  buf

  (
    G7_n_spl_11,
    G7_n_spl_1
  );


  buf

  (
    G7_n_spl_110,
    G7_n_spl_11
  );


  buf

  (
    G7_n_spl_111,
    G7_n_spl_11
  );


  buf

  (
    g149_p_spl_,
    g149_p
  );


  buf

  (
    g150_n_spl_,
    g150_n
  );


  buf

  (
    g149_n_spl_,
    g149_n
  );


  buf

  (
    g150_p_spl_,
    g150_p
  );


  buf

  (
    g151_n_spl_,
    g151_n
  );


  buf

  (
    g151_p_spl_,
    g151_p
  );


  buf

  (
    g152_n_spl_,
    g152_n
  );


  buf

  (
    g152_n_spl_0,
    g152_n_spl_
  );


  buf

  (
    g152_p_spl_,
    g152_p
  );


  buf

  (
    g152_p_spl_0,
    g152_p_spl_
  );


  buf

  (
    g154_n_spl_,
    g154_n
  );


  buf

  (
    g154_p_spl_,
    g154_p
  );


  buf

  (
    g155_n_spl_,
    g155_n
  );


  buf

  (
    g155_p_spl_,
    g155_p
  );


  buf

  (
    g148_n_spl_,
    g148_n
  );


  buf

  (
    g157_p_spl_,
    g157_p
  );


  buf

  (
    g148_p_spl_,
    g148_p
  );


  buf

  (
    g157_n_spl_,
    g157_n
  );


  buf

  (
    g158_n_spl_,
    g158_n
  );


  buf

  (
    g158_p_spl_,
    g158_p
  );


  buf

  (
    g147_n_spl_,
    g147_n
  );


  buf

  (
    g160_p_spl_,
    g160_p
  );


  buf

  (
    g147_p_spl_,
    g147_p
  );


  buf

  (
    g160_n_spl_,
    g160_n
  );


  buf

  (
    g161_n_spl_,
    g161_n
  );


  buf

  (
    g161_p_spl_,
    g161_p
  );


  buf

  (
    g146_n_spl_,
    g146_n
  );


  buf

  (
    g163_p_spl_,
    g163_p
  );


  buf

  (
    g146_p_spl_,
    g146_p
  );


  buf

  (
    g163_n_spl_,
    g163_n
  );


  buf

  (
    g164_n_spl_,
    g164_n
  );


  buf

  (
    g164_p_spl_,
    g164_p
  );


  buf

  (
    g145_n_spl_,
    g145_n
  );


  buf

  (
    g166_p_spl_,
    g166_p
  );


  buf

  (
    g145_p_spl_,
    g145_p
  );


  buf

  (
    g166_n_spl_,
    g166_n
  );


  buf

  (
    g167_n_spl_,
    g167_n
  );


  buf

  (
    g167_p_spl_,
    g167_p
  );


  buf

  (
    g144_n_spl_,
    g144_n
  );


  buf

  (
    g169_p_spl_,
    g169_p
  );


  buf

  (
    g144_p_spl_,
    g144_p
  );


  buf

  (
    g169_n_spl_,
    g169_n
  );


  buf

  (
    g170_n_spl_,
    g170_n
  );


  buf

  (
    g170_p_spl_,
    g170_p
  );


  buf

  (
    g143_n_spl_,
    g143_n
  );


  buf

  (
    g172_p_spl_,
    g172_p
  );


  buf

  (
    g143_p_spl_,
    g143_p
  );


  buf

  (
    g172_n_spl_,
    g172_n
  );


  buf

  (
    g173_n_spl_,
    g173_n
  );


  buf

  (
    g173_p_spl_,
    g173_p
  );


  buf

  (
    g142_n_spl_,
    g142_n
  );


  buf

  (
    g175_p_spl_,
    g175_p
  );


  buf

  (
    g142_p_spl_,
    g142_p
  );


  buf

  (
    g175_n_spl_,
    g175_n
  );


  buf

  (
    g176_n_spl_,
    g176_n
  );


  buf

  (
    g176_p_spl_,
    g176_p
  );


  buf

  (
    g141_n_spl_,
    g141_n
  );


  buf

  (
    g178_p_spl_,
    g178_p
  );


  buf

  (
    g141_p_spl_,
    g141_p
  );


  buf

  (
    g178_n_spl_,
    g178_n
  );


  buf

  (
    g179_n_spl_,
    g179_n
  );


  buf

  (
    g179_p_spl_,
    g179_p
  );


  buf

  (
    g140_p_spl_,
    g140_p
  );


  buf

  (
    g181_n_spl_,
    g181_n
  );


  buf

  (
    g182_p_spl_,
    g182_p
  );


  buf

  (
    G24_p_spl_,
    G24_p
  );


  buf

  (
    G24_p_spl_0,
    G24_p_spl_
  );


  buf

  (
    G24_p_spl_00,
    G24_p_spl_0
  );


  buf

  (
    G24_p_spl_000,
    G24_p_spl_00
  );


  buf

  (
    G24_p_spl_001,
    G24_p_spl_00
  );


  buf

  (
    G24_p_spl_01,
    G24_p_spl_0
  );


  buf

  (
    G24_p_spl_010,
    G24_p_spl_01
  );


  buf

  (
    G24_p_spl_011,
    G24_p_spl_01
  );


  buf

  (
    G24_p_spl_1,
    G24_p_spl_
  );


  buf

  (
    G24_p_spl_10,
    G24_p_spl_1
  );


  buf

  (
    G24_p_spl_100,
    G24_p_spl_10
  );


  buf

  (
    G24_p_spl_101,
    G24_p_spl_10
  );


  buf

  (
    G24_p_spl_11,
    G24_p_spl_1
  );


  buf

  (
    G24_p_spl_110,
    G24_p_spl_11
  );


  buf

  (
    G24_p_spl_111,
    G24_p_spl_11
  );


  buf

  (
    G24_n_spl_,
    G24_n
  );


  buf

  (
    G24_n_spl_0,
    G24_n_spl_
  );


  buf

  (
    G24_n_spl_00,
    G24_n_spl_0
  );


  buf

  (
    G24_n_spl_000,
    G24_n_spl_00
  );


  buf

  (
    G24_n_spl_001,
    G24_n_spl_00
  );


  buf

  (
    G24_n_spl_01,
    G24_n_spl_0
  );


  buf

  (
    G24_n_spl_010,
    G24_n_spl_01
  );


  buf

  (
    G24_n_spl_011,
    G24_n_spl_01
  );


  buf

  (
    G24_n_spl_1,
    G24_n_spl_
  );


  buf

  (
    G24_n_spl_10,
    G24_n_spl_1
  );


  buf

  (
    G24_n_spl_100,
    G24_n_spl_10
  );


  buf

  (
    G24_n_spl_101,
    G24_n_spl_10
  );


  buf

  (
    G24_n_spl_11,
    G24_n_spl_1
  );


  buf

  (
    G24_n_spl_110,
    G24_n_spl_11
  );


  buf

  (
    G24_n_spl_111,
    G24_n_spl_11
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_00,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_000,
    G8_p_spl_00
  );


  buf

  (
    G8_p_spl_001,
    G8_p_spl_00
  );


  buf

  (
    G8_p_spl_01,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_010,
    G8_p_spl_01
  );


  buf

  (
    G8_p_spl_011,
    G8_p_spl_01
  );


  buf

  (
    G8_p_spl_1,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_10,
    G8_p_spl_1
  );


  buf

  (
    G8_p_spl_100,
    G8_p_spl_10
  );


  buf

  (
    G8_p_spl_101,
    G8_p_spl_10
  );


  buf

  (
    G8_p_spl_11,
    G8_p_spl_1
  );


  buf

  (
    G8_p_spl_110,
    G8_p_spl_11
  );


  buf

  (
    G8_p_spl_111,
    G8_p_spl_11
  );


  buf

  (
    G8_n_spl_,
    G8_n
  );


  buf

  (
    G8_n_spl_0,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_00,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_000,
    G8_n_spl_00
  );


  buf

  (
    G8_n_spl_001,
    G8_n_spl_00
  );


  buf

  (
    G8_n_spl_01,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_010,
    G8_n_spl_01
  );


  buf

  (
    G8_n_spl_011,
    G8_n_spl_01
  );


  buf

  (
    G8_n_spl_1,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_10,
    G8_n_spl_1
  );


  buf

  (
    G8_n_spl_100,
    G8_n_spl_10
  );


  buf

  (
    G8_n_spl_101,
    G8_n_spl_10
  );


  buf

  (
    G8_n_spl_11,
    G8_n_spl_1
  );


  buf

  (
    G8_n_spl_110,
    G8_n_spl_11
  );


  buf

  (
    G8_n_spl_111,
    G8_n_spl_11
  );


  buf

  (
    g196_p_spl_,
    g196_p
  );


  buf

  (
    g197_n_spl_,
    g197_n
  );


  buf

  (
    g196_n_spl_,
    g196_n
  );


  buf

  (
    g197_p_spl_,
    g197_p
  );


  buf

  (
    g198_n_spl_,
    g198_n
  );


  buf

  (
    g198_p_spl_,
    g198_p
  );


  buf

  (
    g199_n_spl_,
    g199_n
  );


  buf

  (
    g199_n_spl_0,
    g199_n_spl_
  );


  buf

  (
    g199_p_spl_,
    g199_p
  );


  buf

  (
    g199_p_spl_0,
    g199_p_spl_
  );


  buf

  (
    g201_n_spl_,
    g201_n
  );


  buf

  (
    g201_p_spl_,
    g201_p
  );


  buf

  (
    g202_n_spl_,
    g202_n
  );


  buf

  (
    g202_p_spl_,
    g202_p
  );


  buf

  (
    g195_n_spl_,
    g195_n
  );


  buf

  (
    g204_p_spl_,
    g204_p
  );


  buf

  (
    g195_p_spl_,
    g195_p
  );


  buf

  (
    g204_n_spl_,
    g204_n
  );


  buf

  (
    g205_n_spl_,
    g205_n
  );


  buf

  (
    g205_p_spl_,
    g205_p
  );


  buf

  (
    g194_n_spl_,
    g194_n
  );


  buf

  (
    g207_p_spl_,
    g207_p
  );


  buf

  (
    g194_p_spl_,
    g194_p
  );


  buf

  (
    g207_n_spl_,
    g207_n
  );


  buf

  (
    g208_n_spl_,
    g208_n
  );


  buf

  (
    g208_p_spl_,
    g208_p
  );


  buf

  (
    g193_n_spl_,
    g193_n
  );


  buf

  (
    g210_p_spl_,
    g210_p
  );


  buf

  (
    g193_p_spl_,
    g193_p
  );


  buf

  (
    g210_n_spl_,
    g210_n
  );


  buf

  (
    g211_n_spl_,
    g211_n
  );


  buf

  (
    g211_p_spl_,
    g211_p
  );


  buf

  (
    g192_n_spl_,
    g192_n
  );


  buf

  (
    g213_p_spl_,
    g213_p
  );


  buf

  (
    g192_p_spl_,
    g192_p
  );


  buf

  (
    g213_n_spl_,
    g213_n
  );


  buf

  (
    g214_n_spl_,
    g214_n
  );


  buf

  (
    g214_p_spl_,
    g214_p
  );


  buf

  (
    g191_n_spl_,
    g191_n
  );


  buf

  (
    g216_p_spl_,
    g216_p
  );


  buf

  (
    g191_p_spl_,
    g191_p
  );


  buf

  (
    g216_n_spl_,
    g216_n
  );


  buf

  (
    g217_n_spl_,
    g217_n
  );


  buf

  (
    g217_p_spl_,
    g217_p
  );


  buf

  (
    g190_n_spl_,
    g190_n
  );


  buf

  (
    g219_p_spl_,
    g219_p
  );


  buf

  (
    g190_p_spl_,
    g190_p
  );


  buf

  (
    g219_n_spl_,
    g219_n
  );


  buf

  (
    g220_n_spl_,
    g220_n
  );


  buf

  (
    g220_p_spl_,
    g220_p
  );


  buf

  (
    g189_n_spl_,
    g189_n
  );


  buf

  (
    g222_p_spl_,
    g222_p
  );


  buf

  (
    g189_p_spl_,
    g189_p
  );


  buf

  (
    g222_n_spl_,
    g222_n
  );


  buf

  (
    g223_n_spl_,
    g223_n
  );


  buf

  (
    g223_p_spl_,
    g223_p
  );


  buf

  (
    g188_n_spl_,
    g188_n
  );


  buf

  (
    g225_p_spl_,
    g225_p
  );


  buf

  (
    g188_p_spl_,
    g188_p
  );


  buf

  (
    g225_n_spl_,
    g225_n
  );


  buf

  (
    g226_n_spl_,
    g226_n
  );


  buf

  (
    g226_p_spl_,
    g226_p
  );


  buf

  (
    g187_n_spl_,
    g187_n
  );


  buf

  (
    g228_p_spl_,
    g228_p
  );


  buf

  (
    g187_p_spl_,
    g187_p
  );


  buf

  (
    g228_n_spl_,
    g228_n
  );


  buf

  (
    g229_n_spl_,
    g229_n
  );


  buf

  (
    g229_p_spl_,
    g229_p
  );


  buf

  (
    g186_n_spl_,
    g186_n
  );


  buf

  (
    g231_p_spl_,
    g231_p
  );


  buf

  (
    g186_p_spl_,
    g186_p
  );


  buf

  (
    g231_n_spl_,
    g231_n
  );


  buf

  (
    g232_n_spl_,
    g232_n
  );


  buf

  (
    g232_p_spl_,
    g232_p
  );


  buf

  (
    g185_p_spl_,
    g185_p
  );


  buf

  (
    g234_n_spl_,
    g234_n
  );


  buf

  (
    g235_p_spl_,
    g235_p
  );


  buf

  (
    G25_p_spl_,
    G25_p
  );


  buf

  (
    G25_p_spl_0,
    G25_p_spl_
  );


  buf

  (
    G25_p_spl_00,
    G25_p_spl_0
  );


  buf

  (
    G25_p_spl_000,
    G25_p_spl_00
  );


  buf

  (
    G25_p_spl_001,
    G25_p_spl_00
  );


  buf

  (
    G25_p_spl_01,
    G25_p_spl_0
  );


  buf

  (
    G25_p_spl_010,
    G25_p_spl_01
  );


  buf

  (
    G25_p_spl_011,
    G25_p_spl_01
  );


  buf

  (
    G25_p_spl_1,
    G25_p_spl_
  );


  buf

  (
    G25_p_spl_10,
    G25_p_spl_1
  );


  buf

  (
    G25_p_spl_100,
    G25_p_spl_10
  );


  buf

  (
    G25_p_spl_101,
    G25_p_spl_10
  );


  buf

  (
    G25_p_spl_11,
    G25_p_spl_1
  );


  buf

  (
    G25_p_spl_110,
    G25_p_spl_11
  );


  buf

  (
    G25_p_spl_111,
    G25_p_spl_11
  );


  buf

  (
    G25_n_spl_,
    G25_n
  );


  buf

  (
    G25_n_spl_0,
    G25_n_spl_
  );


  buf

  (
    G25_n_spl_00,
    G25_n_spl_0
  );


  buf

  (
    G25_n_spl_000,
    G25_n_spl_00
  );


  buf

  (
    G25_n_spl_001,
    G25_n_spl_00
  );


  buf

  (
    G25_n_spl_01,
    G25_n_spl_0
  );


  buf

  (
    G25_n_spl_010,
    G25_n_spl_01
  );


  buf

  (
    G25_n_spl_011,
    G25_n_spl_01
  );


  buf

  (
    G25_n_spl_1,
    G25_n_spl_
  );


  buf

  (
    G25_n_spl_10,
    G25_n_spl_1
  );


  buf

  (
    G25_n_spl_100,
    G25_n_spl_10
  );


  buf

  (
    G25_n_spl_101,
    G25_n_spl_10
  );


  buf

  (
    G25_n_spl_11,
    G25_n_spl_1
  );


  buf

  (
    G25_n_spl_110,
    G25_n_spl_11
  );


  buf

  (
    G25_n_spl_111,
    G25_n_spl_11
  );


  buf

  (
    G9_p_spl_,
    G9_p
  );


  buf

  (
    G9_p_spl_0,
    G9_p_spl_
  );


  buf

  (
    G9_p_spl_00,
    G9_p_spl_0
  );


  buf

  (
    G9_p_spl_000,
    G9_p_spl_00
  );


  buf

  (
    G9_p_spl_001,
    G9_p_spl_00
  );


  buf

  (
    G9_p_spl_01,
    G9_p_spl_0
  );


  buf

  (
    G9_p_spl_010,
    G9_p_spl_01
  );


  buf

  (
    G9_p_spl_011,
    G9_p_spl_01
  );


  buf

  (
    G9_p_spl_1,
    G9_p_spl_
  );


  buf

  (
    G9_p_spl_10,
    G9_p_spl_1
  );


  buf

  (
    G9_p_spl_100,
    G9_p_spl_10
  );


  buf

  (
    G9_p_spl_101,
    G9_p_spl_10
  );


  buf

  (
    G9_p_spl_11,
    G9_p_spl_1
  );


  buf

  (
    G9_p_spl_110,
    G9_p_spl_11
  );


  buf

  (
    G9_p_spl_111,
    G9_p_spl_11
  );


  buf

  (
    G9_n_spl_,
    G9_n
  );


  buf

  (
    G9_n_spl_0,
    G9_n_spl_
  );


  buf

  (
    G9_n_spl_00,
    G9_n_spl_0
  );


  buf

  (
    G9_n_spl_000,
    G9_n_spl_00
  );


  buf

  (
    G9_n_spl_001,
    G9_n_spl_00
  );


  buf

  (
    G9_n_spl_01,
    G9_n_spl_0
  );


  buf

  (
    G9_n_spl_010,
    G9_n_spl_01
  );


  buf

  (
    G9_n_spl_011,
    G9_n_spl_01
  );


  buf

  (
    G9_n_spl_1,
    G9_n_spl_
  );


  buf

  (
    G9_n_spl_10,
    G9_n_spl_1
  );


  buf

  (
    G9_n_spl_100,
    G9_n_spl_10
  );


  buf

  (
    G9_n_spl_101,
    G9_n_spl_10
  );


  buf

  (
    G9_n_spl_11,
    G9_n_spl_1
  );


  buf

  (
    G9_n_spl_110,
    G9_n_spl_11
  );


  buf

  (
    G9_n_spl_111,
    G9_n_spl_11
  );


  buf

  (
    g251_p_spl_,
    g251_p
  );


  buf

  (
    g252_n_spl_,
    g252_n
  );


  buf

  (
    g251_n_spl_,
    g251_n
  );


  buf

  (
    g252_p_spl_,
    g252_p
  );


  buf

  (
    g253_n_spl_,
    g253_n
  );


  buf

  (
    g253_p_spl_,
    g253_p
  );


  buf

  (
    g254_n_spl_,
    g254_n
  );


  buf

  (
    g254_n_spl_0,
    g254_n_spl_
  );


  buf

  (
    g254_p_spl_,
    g254_p
  );


  buf

  (
    g254_p_spl_0,
    g254_p_spl_
  );


  buf

  (
    g256_n_spl_,
    g256_n
  );


  buf

  (
    g256_p_spl_,
    g256_p
  );


  buf

  (
    g257_n_spl_,
    g257_n
  );


  buf

  (
    g257_p_spl_,
    g257_p
  );


  buf

  (
    g250_n_spl_,
    g250_n
  );


  buf

  (
    g259_p_spl_,
    g259_p
  );


  buf

  (
    g250_p_spl_,
    g250_p
  );


  buf

  (
    g259_n_spl_,
    g259_n
  );


  buf

  (
    g260_n_spl_,
    g260_n
  );


  buf

  (
    g260_p_spl_,
    g260_p
  );


  buf

  (
    g249_n_spl_,
    g249_n
  );


  buf

  (
    g262_p_spl_,
    g262_p
  );


  buf

  (
    g249_p_spl_,
    g249_p
  );


  buf

  (
    g262_n_spl_,
    g262_n
  );


  buf

  (
    g263_n_spl_,
    g263_n
  );


  buf

  (
    g263_p_spl_,
    g263_p
  );


  buf

  (
    g248_n_spl_,
    g248_n
  );


  buf

  (
    g265_p_spl_,
    g265_p
  );


  buf

  (
    g248_p_spl_,
    g248_p
  );


  buf

  (
    g265_n_spl_,
    g265_n
  );


  buf

  (
    g266_n_spl_,
    g266_n
  );


  buf

  (
    g266_p_spl_,
    g266_p
  );


  buf

  (
    g247_n_spl_,
    g247_n
  );


  buf

  (
    g268_p_spl_,
    g268_p
  );


  buf

  (
    g247_p_spl_,
    g247_p
  );


  buf

  (
    g268_n_spl_,
    g268_n
  );


  buf

  (
    g269_n_spl_,
    g269_n
  );


  buf

  (
    g269_p_spl_,
    g269_p
  );


  buf

  (
    g246_n_spl_,
    g246_n
  );


  buf

  (
    g271_p_spl_,
    g271_p
  );


  buf

  (
    g246_p_spl_,
    g246_p
  );


  buf

  (
    g271_n_spl_,
    g271_n
  );


  buf

  (
    g272_n_spl_,
    g272_n
  );


  buf

  (
    g272_p_spl_,
    g272_p
  );


  buf

  (
    g245_n_spl_,
    g245_n
  );


  buf

  (
    g274_p_spl_,
    g274_p
  );


  buf

  (
    g245_p_spl_,
    g245_p
  );


  buf

  (
    g274_n_spl_,
    g274_n
  );


  buf

  (
    g275_n_spl_,
    g275_n
  );


  buf

  (
    g275_p_spl_,
    g275_p
  );


  buf

  (
    g244_n_spl_,
    g244_n
  );


  buf

  (
    g277_p_spl_,
    g277_p
  );


  buf

  (
    g244_p_spl_,
    g244_p
  );


  buf

  (
    g277_n_spl_,
    g277_n
  );


  buf

  (
    g278_n_spl_,
    g278_n
  );


  buf

  (
    g278_p_spl_,
    g278_p
  );


  buf

  (
    g243_n_spl_,
    g243_n
  );


  buf

  (
    g280_p_spl_,
    g280_p
  );


  buf

  (
    g243_p_spl_,
    g243_p
  );


  buf

  (
    g280_n_spl_,
    g280_n
  );


  buf

  (
    g281_n_spl_,
    g281_n
  );


  buf

  (
    g281_p_spl_,
    g281_p
  );


  buf

  (
    g242_n_spl_,
    g242_n
  );


  buf

  (
    g283_p_spl_,
    g283_p
  );


  buf

  (
    g242_p_spl_,
    g242_p
  );


  buf

  (
    g283_n_spl_,
    g283_n
  );


  buf

  (
    g284_n_spl_,
    g284_n
  );


  buf

  (
    g284_p_spl_,
    g284_p
  );


  buf

  (
    g241_n_spl_,
    g241_n
  );


  buf

  (
    g286_p_spl_,
    g286_p
  );


  buf

  (
    g241_p_spl_,
    g241_p
  );


  buf

  (
    g286_n_spl_,
    g286_n
  );


  buf

  (
    g287_n_spl_,
    g287_n
  );


  buf

  (
    g287_p_spl_,
    g287_p
  );


  buf

  (
    g240_n_spl_,
    g240_n
  );


  buf

  (
    g289_p_spl_,
    g289_p
  );


  buf

  (
    g240_p_spl_,
    g240_p
  );


  buf

  (
    g289_n_spl_,
    g289_n
  );


  buf

  (
    g290_n_spl_,
    g290_n
  );


  buf

  (
    g290_p_spl_,
    g290_p
  );


  buf

  (
    g239_n_spl_,
    g239_n
  );


  buf

  (
    g292_p_spl_,
    g292_p
  );


  buf

  (
    g239_p_spl_,
    g239_p
  );


  buf

  (
    g292_n_spl_,
    g292_n
  );


  buf

  (
    g293_n_spl_,
    g293_n
  );


  buf

  (
    g293_p_spl_,
    g293_p
  );


  buf

  (
    g238_p_spl_,
    g238_p
  );


  buf

  (
    g295_n_spl_,
    g295_n
  );


  buf

  (
    g296_p_spl_,
    g296_p
  );


  buf

  (
    G26_p_spl_,
    G26_p
  );


  buf

  (
    G26_p_spl_0,
    G26_p_spl_
  );


  buf

  (
    G26_p_spl_00,
    G26_p_spl_0
  );


  buf

  (
    G26_p_spl_000,
    G26_p_spl_00
  );


  buf

  (
    G26_p_spl_001,
    G26_p_spl_00
  );


  buf

  (
    G26_p_spl_01,
    G26_p_spl_0
  );


  buf

  (
    G26_p_spl_010,
    G26_p_spl_01
  );


  buf

  (
    G26_p_spl_011,
    G26_p_spl_01
  );


  buf

  (
    G26_p_spl_1,
    G26_p_spl_
  );


  buf

  (
    G26_p_spl_10,
    G26_p_spl_1
  );


  buf

  (
    G26_p_spl_100,
    G26_p_spl_10
  );


  buf

  (
    G26_p_spl_101,
    G26_p_spl_10
  );


  buf

  (
    G26_p_spl_11,
    G26_p_spl_1
  );


  buf

  (
    G26_p_spl_110,
    G26_p_spl_11
  );


  buf

  (
    G26_p_spl_111,
    G26_p_spl_11
  );


  buf

  (
    G26_n_spl_,
    G26_n
  );


  buf

  (
    G26_n_spl_0,
    G26_n_spl_
  );


  buf

  (
    G26_n_spl_00,
    G26_n_spl_0
  );


  buf

  (
    G26_n_spl_000,
    G26_n_spl_00
  );


  buf

  (
    G26_n_spl_001,
    G26_n_spl_00
  );


  buf

  (
    G26_n_spl_01,
    G26_n_spl_0
  );


  buf

  (
    G26_n_spl_010,
    G26_n_spl_01
  );


  buf

  (
    G26_n_spl_011,
    G26_n_spl_01
  );


  buf

  (
    G26_n_spl_1,
    G26_n_spl_
  );


  buf

  (
    G26_n_spl_10,
    G26_n_spl_1
  );


  buf

  (
    G26_n_spl_100,
    G26_n_spl_10
  );


  buf

  (
    G26_n_spl_101,
    G26_n_spl_10
  );


  buf

  (
    G26_n_spl_11,
    G26_n_spl_1
  );


  buf

  (
    G26_n_spl_110,
    G26_n_spl_11
  );


  buf

  (
    G26_n_spl_111,
    G26_n_spl_11
  );


  buf

  (
    G10_p_spl_,
    G10_p
  );


  buf

  (
    G10_p_spl_0,
    G10_p_spl_
  );


  buf

  (
    G10_p_spl_00,
    G10_p_spl_0
  );


  buf

  (
    G10_p_spl_000,
    G10_p_spl_00
  );


  buf

  (
    G10_p_spl_001,
    G10_p_spl_00
  );


  buf

  (
    G10_p_spl_01,
    G10_p_spl_0
  );


  buf

  (
    G10_p_spl_010,
    G10_p_spl_01
  );


  buf

  (
    G10_p_spl_011,
    G10_p_spl_01
  );


  buf

  (
    G10_p_spl_1,
    G10_p_spl_
  );


  buf

  (
    G10_p_spl_10,
    G10_p_spl_1
  );


  buf

  (
    G10_p_spl_100,
    G10_p_spl_10
  );


  buf

  (
    G10_p_spl_101,
    G10_p_spl_10
  );


  buf

  (
    G10_p_spl_11,
    G10_p_spl_1
  );


  buf

  (
    G10_p_spl_110,
    G10_p_spl_11
  );


  buf

  (
    G10_p_spl_111,
    G10_p_spl_11
  );


  buf

  (
    G10_n_spl_,
    G10_n
  );


  buf

  (
    G10_n_spl_0,
    G10_n_spl_
  );


  buf

  (
    G10_n_spl_00,
    G10_n_spl_0
  );


  buf

  (
    G10_n_spl_000,
    G10_n_spl_00
  );


  buf

  (
    G10_n_spl_001,
    G10_n_spl_00
  );


  buf

  (
    G10_n_spl_01,
    G10_n_spl_0
  );


  buf

  (
    G10_n_spl_010,
    G10_n_spl_01
  );


  buf

  (
    G10_n_spl_011,
    G10_n_spl_01
  );


  buf

  (
    G10_n_spl_1,
    G10_n_spl_
  );


  buf

  (
    G10_n_spl_10,
    G10_n_spl_1
  );


  buf

  (
    G10_n_spl_100,
    G10_n_spl_10
  );


  buf

  (
    G10_n_spl_101,
    G10_n_spl_10
  );


  buf

  (
    G10_n_spl_11,
    G10_n_spl_1
  );


  buf

  (
    G10_n_spl_110,
    G10_n_spl_11
  );


  buf

  (
    G10_n_spl_111,
    G10_n_spl_11
  );


  buf

  (
    g314_p_spl_,
    g314_p
  );


  buf

  (
    g315_n_spl_,
    g315_n
  );


  buf

  (
    g314_n_spl_,
    g314_n
  );


  buf

  (
    g315_p_spl_,
    g315_p
  );


  buf

  (
    g316_n_spl_,
    g316_n
  );


  buf

  (
    g316_p_spl_,
    g316_p
  );


  buf

  (
    g317_n_spl_,
    g317_n
  );


  buf

  (
    g317_n_spl_0,
    g317_n_spl_
  );


  buf

  (
    g317_p_spl_,
    g317_p
  );


  buf

  (
    g317_p_spl_0,
    g317_p_spl_
  );


  buf

  (
    g319_n_spl_,
    g319_n
  );


  buf

  (
    g319_p_spl_,
    g319_p
  );


  buf

  (
    g320_n_spl_,
    g320_n
  );


  buf

  (
    g320_p_spl_,
    g320_p
  );


  buf

  (
    g313_n_spl_,
    g313_n
  );


  buf

  (
    g322_p_spl_,
    g322_p
  );


  buf

  (
    g313_p_spl_,
    g313_p
  );


  buf

  (
    g322_n_spl_,
    g322_n
  );


  buf

  (
    g323_n_spl_,
    g323_n
  );


  buf

  (
    g323_p_spl_,
    g323_p
  );


  buf

  (
    g312_n_spl_,
    g312_n
  );


  buf

  (
    g325_p_spl_,
    g325_p
  );


  buf

  (
    g312_p_spl_,
    g312_p
  );


  buf

  (
    g325_n_spl_,
    g325_n
  );


  buf

  (
    g326_n_spl_,
    g326_n
  );


  buf

  (
    g326_p_spl_,
    g326_p
  );


  buf

  (
    g311_n_spl_,
    g311_n
  );


  buf

  (
    g328_p_spl_,
    g328_p
  );


  buf

  (
    g311_p_spl_,
    g311_p
  );


  buf

  (
    g328_n_spl_,
    g328_n
  );


  buf

  (
    g329_n_spl_,
    g329_n
  );


  buf

  (
    g329_p_spl_,
    g329_p
  );


  buf

  (
    g310_n_spl_,
    g310_n
  );


  buf

  (
    g331_p_spl_,
    g331_p
  );


  buf

  (
    g310_p_spl_,
    g310_p
  );


  buf

  (
    g331_n_spl_,
    g331_n
  );


  buf

  (
    g332_n_spl_,
    g332_n
  );


  buf

  (
    g332_p_spl_,
    g332_p
  );


  buf

  (
    g309_n_spl_,
    g309_n
  );


  buf

  (
    g334_p_spl_,
    g334_p
  );


  buf

  (
    g309_p_spl_,
    g309_p
  );


  buf

  (
    g334_n_spl_,
    g334_n
  );


  buf

  (
    g335_n_spl_,
    g335_n
  );


  buf

  (
    g335_p_spl_,
    g335_p
  );


  buf

  (
    g308_n_spl_,
    g308_n
  );


  buf

  (
    g337_p_spl_,
    g337_p
  );


  buf

  (
    g308_p_spl_,
    g308_p
  );


  buf

  (
    g337_n_spl_,
    g337_n
  );


  buf

  (
    g338_n_spl_,
    g338_n
  );


  buf

  (
    g338_p_spl_,
    g338_p
  );


  buf

  (
    g307_n_spl_,
    g307_n
  );


  buf

  (
    g340_p_spl_,
    g340_p
  );


  buf

  (
    g307_p_spl_,
    g307_p
  );


  buf

  (
    g340_n_spl_,
    g340_n
  );


  buf

  (
    g341_n_spl_,
    g341_n
  );


  buf

  (
    g341_p_spl_,
    g341_p
  );


  buf

  (
    g306_n_spl_,
    g306_n
  );


  buf

  (
    g343_p_spl_,
    g343_p
  );


  buf

  (
    g306_p_spl_,
    g306_p
  );


  buf

  (
    g343_n_spl_,
    g343_n
  );


  buf

  (
    g344_n_spl_,
    g344_n
  );


  buf

  (
    g344_p_spl_,
    g344_p
  );


  buf

  (
    g305_n_spl_,
    g305_n
  );


  buf

  (
    g346_p_spl_,
    g346_p
  );


  buf

  (
    g305_p_spl_,
    g305_p
  );


  buf

  (
    g346_n_spl_,
    g346_n
  );


  buf

  (
    g347_n_spl_,
    g347_n
  );


  buf

  (
    g347_p_spl_,
    g347_p
  );


  buf

  (
    g304_n_spl_,
    g304_n
  );


  buf

  (
    g349_p_spl_,
    g349_p
  );


  buf

  (
    g304_p_spl_,
    g304_p
  );


  buf

  (
    g349_n_spl_,
    g349_n
  );


  buf

  (
    g350_n_spl_,
    g350_n
  );


  buf

  (
    g350_p_spl_,
    g350_p
  );


  buf

  (
    g303_n_spl_,
    g303_n
  );


  buf

  (
    g352_p_spl_,
    g352_p
  );


  buf

  (
    g303_p_spl_,
    g303_p
  );


  buf

  (
    g352_n_spl_,
    g352_n
  );


  buf

  (
    g353_n_spl_,
    g353_n
  );


  buf

  (
    g353_p_spl_,
    g353_p
  );


  buf

  (
    g302_n_spl_,
    g302_n
  );


  buf

  (
    g355_p_spl_,
    g355_p
  );


  buf

  (
    g302_p_spl_,
    g302_p
  );


  buf

  (
    g355_n_spl_,
    g355_n
  );


  buf

  (
    g356_n_spl_,
    g356_n
  );


  buf

  (
    g356_p_spl_,
    g356_p
  );


  buf

  (
    g301_n_spl_,
    g301_n
  );


  buf

  (
    g358_p_spl_,
    g358_p
  );


  buf

  (
    g301_p_spl_,
    g301_p
  );


  buf

  (
    g358_n_spl_,
    g358_n
  );


  buf

  (
    g359_n_spl_,
    g359_n
  );


  buf

  (
    g359_p_spl_,
    g359_p
  );


  buf

  (
    g300_n_spl_,
    g300_n
  );


  buf

  (
    g361_p_spl_,
    g361_p
  );


  buf

  (
    g300_p_spl_,
    g300_p
  );


  buf

  (
    g361_n_spl_,
    g361_n
  );


  buf

  (
    g362_n_spl_,
    g362_n
  );


  buf

  (
    g362_p_spl_,
    g362_p
  );


  buf

  (
    g299_p_spl_,
    g299_p
  );


  buf

  (
    g364_n_spl_,
    g364_n
  );


  buf

  (
    g365_p_spl_,
    g365_p
  );


  buf

  (
    G27_p_spl_,
    G27_p
  );


  buf

  (
    G27_p_spl_0,
    G27_p_spl_
  );


  buf

  (
    G27_p_spl_00,
    G27_p_spl_0
  );


  buf

  (
    G27_p_spl_000,
    G27_p_spl_00
  );


  buf

  (
    G27_p_spl_001,
    G27_p_spl_00
  );


  buf

  (
    G27_p_spl_01,
    G27_p_spl_0
  );


  buf

  (
    G27_p_spl_010,
    G27_p_spl_01
  );


  buf

  (
    G27_p_spl_011,
    G27_p_spl_01
  );


  buf

  (
    G27_p_spl_1,
    G27_p_spl_
  );


  buf

  (
    G27_p_spl_10,
    G27_p_spl_1
  );


  buf

  (
    G27_p_spl_100,
    G27_p_spl_10
  );


  buf

  (
    G27_p_spl_101,
    G27_p_spl_10
  );


  buf

  (
    G27_p_spl_11,
    G27_p_spl_1
  );


  buf

  (
    G27_p_spl_110,
    G27_p_spl_11
  );


  buf

  (
    G27_p_spl_111,
    G27_p_spl_11
  );


  buf

  (
    G27_n_spl_,
    G27_n
  );


  buf

  (
    G27_n_spl_0,
    G27_n_spl_
  );


  buf

  (
    G27_n_spl_00,
    G27_n_spl_0
  );


  buf

  (
    G27_n_spl_000,
    G27_n_spl_00
  );


  buf

  (
    G27_n_spl_001,
    G27_n_spl_00
  );


  buf

  (
    G27_n_spl_01,
    G27_n_spl_0
  );


  buf

  (
    G27_n_spl_010,
    G27_n_spl_01
  );


  buf

  (
    G27_n_spl_011,
    G27_n_spl_01
  );


  buf

  (
    G27_n_spl_1,
    G27_n_spl_
  );


  buf

  (
    G27_n_spl_10,
    G27_n_spl_1
  );


  buf

  (
    G27_n_spl_100,
    G27_n_spl_10
  );


  buf

  (
    G27_n_spl_101,
    G27_n_spl_10
  );


  buf

  (
    G27_n_spl_11,
    G27_n_spl_1
  );


  buf

  (
    G27_n_spl_110,
    G27_n_spl_11
  );


  buf

  (
    G27_n_spl_111,
    G27_n_spl_11
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    G11_p_spl_0,
    G11_p_spl_
  );


  buf

  (
    G11_p_spl_00,
    G11_p_spl_0
  );


  buf

  (
    G11_p_spl_000,
    G11_p_spl_00
  );


  buf

  (
    G11_p_spl_001,
    G11_p_spl_00
  );


  buf

  (
    G11_p_spl_01,
    G11_p_spl_0
  );


  buf

  (
    G11_p_spl_010,
    G11_p_spl_01
  );


  buf

  (
    G11_p_spl_011,
    G11_p_spl_01
  );


  buf

  (
    G11_p_spl_1,
    G11_p_spl_
  );


  buf

  (
    G11_p_spl_10,
    G11_p_spl_1
  );


  buf

  (
    G11_p_spl_100,
    G11_p_spl_10
  );


  buf

  (
    G11_p_spl_101,
    G11_p_spl_10
  );


  buf

  (
    G11_p_spl_11,
    G11_p_spl_1
  );


  buf

  (
    G11_p_spl_110,
    G11_p_spl_11
  );


  buf

  (
    G11_p_spl_111,
    G11_p_spl_11
  );


  buf

  (
    G11_n_spl_,
    G11_n
  );


  buf

  (
    G11_n_spl_0,
    G11_n_spl_
  );


  buf

  (
    G11_n_spl_00,
    G11_n_spl_0
  );


  buf

  (
    G11_n_spl_000,
    G11_n_spl_00
  );


  buf

  (
    G11_n_spl_001,
    G11_n_spl_00
  );


  buf

  (
    G11_n_spl_01,
    G11_n_spl_0
  );


  buf

  (
    G11_n_spl_010,
    G11_n_spl_01
  );


  buf

  (
    G11_n_spl_011,
    G11_n_spl_01
  );


  buf

  (
    G11_n_spl_1,
    G11_n_spl_
  );


  buf

  (
    G11_n_spl_10,
    G11_n_spl_1
  );


  buf

  (
    G11_n_spl_100,
    G11_n_spl_10
  );


  buf

  (
    G11_n_spl_101,
    G11_n_spl_10
  );


  buf

  (
    G11_n_spl_11,
    G11_n_spl_1
  );


  buf

  (
    G11_n_spl_110,
    G11_n_spl_11
  );


  buf

  (
    G11_n_spl_111,
    G11_n_spl_11
  );


  buf

  (
    g385_p_spl_,
    g385_p
  );


  buf

  (
    g386_n_spl_,
    g386_n
  );


  buf

  (
    g385_n_spl_,
    g385_n
  );


  buf

  (
    g386_p_spl_,
    g386_p
  );


  buf

  (
    g387_n_spl_,
    g387_n
  );


  buf

  (
    g387_p_spl_,
    g387_p
  );


  buf

  (
    g388_n_spl_,
    g388_n
  );


  buf

  (
    g388_n_spl_0,
    g388_n_spl_
  );


  buf

  (
    g388_p_spl_,
    g388_p
  );


  buf

  (
    g388_p_spl_0,
    g388_p_spl_
  );


  buf

  (
    g390_n_spl_,
    g390_n
  );


  buf

  (
    g390_p_spl_,
    g390_p
  );


  buf

  (
    g391_n_spl_,
    g391_n
  );


  buf

  (
    g391_p_spl_,
    g391_p
  );


  buf

  (
    g384_n_spl_,
    g384_n
  );


  buf

  (
    g393_p_spl_,
    g393_p
  );


  buf

  (
    g384_p_spl_,
    g384_p
  );


  buf

  (
    g393_n_spl_,
    g393_n
  );


  buf

  (
    g394_n_spl_,
    g394_n
  );


  buf

  (
    g394_p_spl_,
    g394_p
  );


  buf

  (
    g383_n_spl_,
    g383_n
  );


  buf

  (
    g396_p_spl_,
    g396_p
  );


  buf

  (
    g383_p_spl_,
    g383_p
  );


  buf

  (
    g396_n_spl_,
    g396_n
  );


  buf

  (
    g397_n_spl_,
    g397_n
  );


  buf

  (
    g397_p_spl_,
    g397_p
  );


  buf

  (
    g382_n_spl_,
    g382_n
  );


  buf

  (
    g399_p_spl_,
    g399_p
  );


  buf

  (
    g382_p_spl_,
    g382_p
  );


  buf

  (
    g399_n_spl_,
    g399_n
  );


  buf

  (
    g400_n_spl_,
    g400_n
  );


  buf

  (
    g400_p_spl_,
    g400_p
  );


  buf

  (
    g381_n_spl_,
    g381_n
  );


  buf

  (
    g402_p_spl_,
    g402_p
  );


  buf

  (
    g381_p_spl_,
    g381_p
  );


  buf

  (
    g402_n_spl_,
    g402_n
  );


  buf

  (
    g403_n_spl_,
    g403_n
  );


  buf

  (
    g403_p_spl_,
    g403_p
  );


  buf

  (
    g380_n_spl_,
    g380_n
  );


  buf

  (
    g405_p_spl_,
    g405_p
  );


  buf

  (
    g380_p_spl_,
    g380_p
  );


  buf

  (
    g405_n_spl_,
    g405_n
  );


  buf

  (
    g406_n_spl_,
    g406_n
  );


  buf

  (
    g406_p_spl_,
    g406_p
  );


  buf

  (
    g379_n_spl_,
    g379_n
  );


  buf

  (
    g408_p_spl_,
    g408_p
  );


  buf

  (
    g379_p_spl_,
    g379_p
  );


  buf

  (
    g408_n_spl_,
    g408_n
  );


  buf

  (
    g409_n_spl_,
    g409_n
  );


  buf

  (
    g409_p_spl_,
    g409_p
  );


  buf

  (
    g378_n_spl_,
    g378_n
  );


  buf

  (
    g411_p_spl_,
    g411_p
  );


  buf

  (
    g378_p_spl_,
    g378_p
  );


  buf

  (
    g411_n_spl_,
    g411_n
  );


  buf

  (
    g412_n_spl_,
    g412_n
  );


  buf

  (
    g412_p_spl_,
    g412_p
  );


  buf

  (
    g377_n_spl_,
    g377_n
  );


  buf

  (
    g414_p_spl_,
    g414_p
  );


  buf

  (
    g377_p_spl_,
    g377_p
  );


  buf

  (
    g414_n_spl_,
    g414_n
  );


  buf

  (
    g415_n_spl_,
    g415_n
  );


  buf

  (
    g415_p_spl_,
    g415_p
  );


  buf

  (
    g376_n_spl_,
    g376_n
  );


  buf

  (
    g417_p_spl_,
    g417_p
  );


  buf

  (
    g376_p_spl_,
    g376_p
  );


  buf

  (
    g417_n_spl_,
    g417_n
  );


  buf

  (
    g418_n_spl_,
    g418_n
  );


  buf

  (
    g418_p_spl_,
    g418_p
  );


  buf

  (
    g375_n_spl_,
    g375_n
  );


  buf

  (
    g420_p_spl_,
    g420_p
  );


  buf

  (
    g375_p_spl_,
    g375_p
  );


  buf

  (
    g420_n_spl_,
    g420_n
  );


  buf

  (
    g421_n_spl_,
    g421_n
  );


  buf

  (
    g421_p_spl_,
    g421_p
  );


  buf

  (
    g374_n_spl_,
    g374_n
  );


  buf

  (
    g423_p_spl_,
    g423_p
  );


  buf

  (
    g374_p_spl_,
    g374_p
  );


  buf

  (
    g423_n_spl_,
    g423_n
  );


  buf

  (
    g424_n_spl_,
    g424_n
  );


  buf

  (
    g424_p_spl_,
    g424_p
  );


  buf

  (
    g373_n_spl_,
    g373_n
  );


  buf

  (
    g426_p_spl_,
    g426_p
  );


  buf

  (
    g373_p_spl_,
    g373_p
  );


  buf

  (
    g426_n_spl_,
    g426_n
  );


  buf

  (
    g427_n_spl_,
    g427_n
  );


  buf

  (
    g427_p_spl_,
    g427_p
  );


  buf

  (
    g372_n_spl_,
    g372_n
  );


  buf

  (
    g429_p_spl_,
    g429_p
  );


  buf

  (
    g372_p_spl_,
    g372_p
  );


  buf

  (
    g429_n_spl_,
    g429_n
  );


  buf

  (
    g430_n_spl_,
    g430_n
  );


  buf

  (
    g430_p_spl_,
    g430_p
  );


  buf

  (
    g371_n_spl_,
    g371_n
  );


  buf

  (
    g432_p_spl_,
    g432_p
  );


  buf

  (
    g371_p_spl_,
    g371_p
  );


  buf

  (
    g432_n_spl_,
    g432_n
  );


  buf

  (
    g433_n_spl_,
    g433_n
  );


  buf

  (
    g433_p_spl_,
    g433_p
  );


  buf

  (
    g370_n_spl_,
    g370_n
  );


  buf

  (
    g435_p_spl_,
    g435_p
  );


  buf

  (
    g370_p_spl_,
    g370_p
  );


  buf

  (
    g435_n_spl_,
    g435_n
  );


  buf

  (
    g436_n_spl_,
    g436_n
  );


  buf

  (
    g436_p_spl_,
    g436_p
  );


  buf

  (
    g369_n_spl_,
    g369_n
  );


  buf

  (
    g438_p_spl_,
    g438_p
  );


  buf

  (
    g369_p_spl_,
    g369_p
  );


  buf

  (
    g438_n_spl_,
    g438_n
  );


  buf

  (
    g439_n_spl_,
    g439_n
  );


  buf

  (
    g439_p_spl_,
    g439_p
  );


  buf

  (
    g368_p_spl_,
    g368_p
  );


  buf

  (
    g441_n_spl_,
    g441_n
  );


  buf

  (
    g442_p_spl_,
    g442_p
  );


  buf

  (
    G28_p_spl_,
    G28_p
  );


  buf

  (
    G28_p_spl_0,
    G28_p_spl_
  );


  buf

  (
    G28_p_spl_00,
    G28_p_spl_0
  );


  buf

  (
    G28_p_spl_000,
    G28_p_spl_00
  );


  buf

  (
    G28_p_spl_001,
    G28_p_spl_00
  );


  buf

  (
    G28_p_spl_01,
    G28_p_spl_0
  );


  buf

  (
    G28_p_spl_010,
    G28_p_spl_01
  );


  buf

  (
    G28_p_spl_011,
    G28_p_spl_01
  );


  buf

  (
    G28_p_spl_1,
    G28_p_spl_
  );


  buf

  (
    G28_p_spl_10,
    G28_p_spl_1
  );


  buf

  (
    G28_p_spl_100,
    G28_p_spl_10
  );


  buf

  (
    G28_p_spl_101,
    G28_p_spl_10
  );


  buf

  (
    G28_p_spl_11,
    G28_p_spl_1
  );


  buf

  (
    G28_p_spl_110,
    G28_p_spl_11
  );


  buf

  (
    G28_p_spl_111,
    G28_p_spl_11
  );


  buf

  (
    G28_n_spl_,
    G28_n
  );


  buf

  (
    G28_n_spl_0,
    G28_n_spl_
  );


  buf

  (
    G28_n_spl_00,
    G28_n_spl_0
  );


  buf

  (
    G28_n_spl_000,
    G28_n_spl_00
  );


  buf

  (
    G28_n_spl_001,
    G28_n_spl_00
  );


  buf

  (
    G28_n_spl_01,
    G28_n_spl_0
  );


  buf

  (
    G28_n_spl_010,
    G28_n_spl_01
  );


  buf

  (
    G28_n_spl_011,
    G28_n_spl_01
  );


  buf

  (
    G28_n_spl_1,
    G28_n_spl_
  );


  buf

  (
    G28_n_spl_10,
    G28_n_spl_1
  );


  buf

  (
    G28_n_spl_100,
    G28_n_spl_10
  );


  buf

  (
    G28_n_spl_101,
    G28_n_spl_10
  );


  buf

  (
    G28_n_spl_11,
    G28_n_spl_1
  );


  buf

  (
    G28_n_spl_110,
    G28_n_spl_11
  );


  buf

  (
    G28_n_spl_111,
    G28_n_spl_11
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G12_p_spl_0,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_00,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_000,
    G12_p_spl_00
  );


  buf

  (
    G12_p_spl_001,
    G12_p_spl_00
  );


  buf

  (
    G12_p_spl_01,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_010,
    G12_p_spl_01
  );


  buf

  (
    G12_p_spl_011,
    G12_p_spl_01
  );


  buf

  (
    G12_p_spl_1,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_10,
    G12_p_spl_1
  );


  buf

  (
    G12_p_spl_100,
    G12_p_spl_10
  );


  buf

  (
    G12_p_spl_101,
    G12_p_spl_10
  );


  buf

  (
    G12_p_spl_11,
    G12_p_spl_1
  );


  buf

  (
    G12_p_spl_110,
    G12_p_spl_11
  );


  buf

  (
    G12_p_spl_111,
    G12_p_spl_11
  );


  buf

  (
    G12_n_spl_,
    G12_n
  );


  buf

  (
    G12_n_spl_0,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_00,
    G12_n_spl_0
  );


  buf

  (
    G12_n_spl_000,
    G12_n_spl_00
  );


  buf

  (
    G12_n_spl_001,
    G12_n_spl_00
  );


  buf

  (
    G12_n_spl_01,
    G12_n_spl_0
  );


  buf

  (
    G12_n_spl_010,
    G12_n_spl_01
  );


  buf

  (
    G12_n_spl_011,
    G12_n_spl_01
  );


  buf

  (
    G12_n_spl_1,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_10,
    G12_n_spl_1
  );


  buf

  (
    G12_n_spl_100,
    G12_n_spl_10
  );


  buf

  (
    G12_n_spl_101,
    G12_n_spl_10
  );


  buf

  (
    G12_n_spl_11,
    G12_n_spl_1
  );


  buf

  (
    G12_n_spl_110,
    G12_n_spl_11
  );


  buf

  (
    G12_n_spl_111,
    G12_n_spl_11
  );


  buf

  (
    g464_p_spl_,
    g464_p
  );


  buf

  (
    g465_n_spl_,
    g465_n
  );


  buf

  (
    g464_n_spl_,
    g464_n
  );


  buf

  (
    g465_p_spl_,
    g465_p
  );


  buf

  (
    g466_n_spl_,
    g466_n
  );


  buf

  (
    g466_p_spl_,
    g466_p
  );


  buf

  (
    g467_n_spl_,
    g467_n
  );


  buf

  (
    g467_n_spl_0,
    g467_n_spl_
  );


  buf

  (
    g467_p_spl_,
    g467_p
  );


  buf

  (
    g467_p_spl_0,
    g467_p_spl_
  );


  buf

  (
    g469_n_spl_,
    g469_n
  );


  buf

  (
    g469_p_spl_,
    g469_p
  );


  buf

  (
    g470_n_spl_,
    g470_n
  );


  buf

  (
    g470_p_spl_,
    g470_p
  );


  buf

  (
    g463_n_spl_,
    g463_n
  );


  buf

  (
    g472_p_spl_,
    g472_p
  );


  buf

  (
    g463_p_spl_,
    g463_p
  );


  buf

  (
    g472_n_spl_,
    g472_n
  );


  buf

  (
    g473_n_spl_,
    g473_n
  );


  buf

  (
    g473_p_spl_,
    g473_p
  );


  buf

  (
    g462_n_spl_,
    g462_n
  );


  buf

  (
    g475_p_spl_,
    g475_p
  );


  buf

  (
    g462_p_spl_,
    g462_p
  );


  buf

  (
    g475_n_spl_,
    g475_n
  );


  buf

  (
    g476_n_spl_,
    g476_n
  );


  buf

  (
    g476_p_spl_,
    g476_p
  );


  buf

  (
    g461_n_spl_,
    g461_n
  );


  buf

  (
    g478_p_spl_,
    g478_p
  );


  buf

  (
    g461_p_spl_,
    g461_p
  );


  buf

  (
    g478_n_spl_,
    g478_n
  );


  buf

  (
    g479_n_spl_,
    g479_n
  );


  buf

  (
    g479_p_spl_,
    g479_p
  );


  buf

  (
    g460_n_spl_,
    g460_n
  );


  buf

  (
    g481_p_spl_,
    g481_p
  );


  buf

  (
    g460_p_spl_,
    g460_p
  );


  buf

  (
    g481_n_spl_,
    g481_n
  );


  buf

  (
    g482_n_spl_,
    g482_n
  );


  buf

  (
    g482_p_spl_,
    g482_p
  );


  buf

  (
    g459_n_spl_,
    g459_n
  );


  buf

  (
    g484_p_spl_,
    g484_p
  );


  buf

  (
    g459_p_spl_,
    g459_p
  );


  buf

  (
    g484_n_spl_,
    g484_n
  );


  buf

  (
    g485_n_spl_,
    g485_n
  );


  buf

  (
    g485_p_spl_,
    g485_p
  );


  buf

  (
    g458_n_spl_,
    g458_n
  );


  buf

  (
    g487_p_spl_,
    g487_p
  );


  buf

  (
    g458_p_spl_,
    g458_p
  );


  buf

  (
    g487_n_spl_,
    g487_n
  );


  buf

  (
    g488_n_spl_,
    g488_n
  );


  buf

  (
    g488_p_spl_,
    g488_p
  );


  buf

  (
    g457_n_spl_,
    g457_n
  );


  buf

  (
    g490_p_spl_,
    g490_p
  );


  buf

  (
    g457_p_spl_,
    g457_p
  );


  buf

  (
    g490_n_spl_,
    g490_n
  );


  buf

  (
    g491_n_spl_,
    g491_n
  );


  buf

  (
    g491_p_spl_,
    g491_p
  );


  buf

  (
    g456_n_spl_,
    g456_n
  );


  buf

  (
    g493_p_spl_,
    g493_p
  );


  buf

  (
    g456_p_spl_,
    g456_p
  );


  buf

  (
    g493_n_spl_,
    g493_n
  );


  buf

  (
    g494_n_spl_,
    g494_n
  );


  buf

  (
    g494_p_spl_,
    g494_p
  );


  buf

  (
    g455_n_spl_,
    g455_n
  );


  buf

  (
    g496_p_spl_,
    g496_p
  );


  buf

  (
    g455_p_spl_,
    g455_p
  );


  buf

  (
    g496_n_spl_,
    g496_n
  );


  buf

  (
    g497_n_spl_,
    g497_n
  );


  buf

  (
    g497_p_spl_,
    g497_p
  );


  buf

  (
    g454_n_spl_,
    g454_n
  );


  buf

  (
    g499_p_spl_,
    g499_p
  );


  buf

  (
    g454_p_spl_,
    g454_p
  );


  buf

  (
    g499_n_spl_,
    g499_n
  );


  buf

  (
    g500_n_spl_,
    g500_n
  );


  buf

  (
    g500_p_spl_,
    g500_p
  );


  buf

  (
    g453_n_spl_,
    g453_n
  );


  buf

  (
    g502_p_spl_,
    g502_p
  );


  buf

  (
    g453_p_spl_,
    g453_p
  );


  buf

  (
    g502_n_spl_,
    g502_n
  );


  buf

  (
    g503_n_spl_,
    g503_n
  );


  buf

  (
    g503_p_spl_,
    g503_p
  );


  buf

  (
    g452_n_spl_,
    g452_n
  );


  buf

  (
    g505_p_spl_,
    g505_p
  );


  buf

  (
    g452_p_spl_,
    g452_p
  );


  buf

  (
    g505_n_spl_,
    g505_n
  );


  buf

  (
    g506_n_spl_,
    g506_n
  );


  buf

  (
    g506_p_spl_,
    g506_p
  );


  buf

  (
    g451_n_spl_,
    g451_n
  );


  buf

  (
    g508_p_spl_,
    g508_p
  );


  buf

  (
    g451_p_spl_,
    g451_p
  );


  buf

  (
    g508_n_spl_,
    g508_n
  );


  buf

  (
    g509_n_spl_,
    g509_n
  );


  buf

  (
    g509_p_spl_,
    g509_p
  );


  buf

  (
    g450_n_spl_,
    g450_n
  );


  buf

  (
    g511_p_spl_,
    g511_p
  );


  buf

  (
    g450_p_spl_,
    g450_p
  );


  buf

  (
    g511_n_spl_,
    g511_n
  );


  buf

  (
    g512_n_spl_,
    g512_n
  );


  buf

  (
    g512_p_spl_,
    g512_p
  );


  buf

  (
    g449_n_spl_,
    g449_n
  );


  buf

  (
    g514_p_spl_,
    g514_p
  );


  buf

  (
    g449_p_spl_,
    g449_p
  );


  buf

  (
    g514_n_spl_,
    g514_n
  );


  buf

  (
    g515_n_spl_,
    g515_n
  );


  buf

  (
    g515_p_spl_,
    g515_p
  );


  buf

  (
    g448_n_spl_,
    g448_n
  );


  buf

  (
    g517_p_spl_,
    g517_p
  );


  buf

  (
    g448_p_spl_,
    g448_p
  );


  buf

  (
    g517_n_spl_,
    g517_n
  );


  buf

  (
    g518_n_spl_,
    g518_n
  );


  buf

  (
    g518_p_spl_,
    g518_p
  );


  buf

  (
    g447_n_spl_,
    g447_n
  );


  buf

  (
    g520_p_spl_,
    g520_p
  );


  buf

  (
    g447_p_spl_,
    g447_p
  );


  buf

  (
    g520_n_spl_,
    g520_n
  );


  buf

  (
    g521_n_spl_,
    g521_n
  );


  buf

  (
    g521_p_spl_,
    g521_p
  );


  buf

  (
    g446_n_spl_,
    g446_n
  );


  buf

  (
    g523_p_spl_,
    g523_p
  );


  buf

  (
    g446_p_spl_,
    g446_p
  );


  buf

  (
    g523_n_spl_,
    g523_n
  );


  buf

  (
    g524_n_spl_,
    g524_n
  );


  buf

  (
    g524_p_spl_,
    g524_p
  );


  buf

  (
    g445_p_spl_,
    g445_p
  );


  buf

  (
    g526_n_spl_,
    g526_n
  );


  buf

  (
    g527_p_spl_,
    g527_p
  );


  buf

  (
    G29_p_spl_,
    G29_p
  );


  buf

  (
    G29_p_spl_0,
    G29_p_spl_
  );


  buf

  (
    G29_p_spl_00,
    G29_p_spl_0
  );


  buf

  (
    G29_p_spl_000,
    G29_p_spl_00
  );


  buf

  (
    G29_p_spl_001,
    G29_p_spl_00
  );


  buf

  (
    G29_p_spl_01,
    G29_p_spl_0
  );


  buf

  (
    G29_p_spl_010,
    G29_p_spl_01
  );


  buf

  (
    G29_p_spl_011,
    G29_p_spl_01
  );


  buf

  (
    G29_p_spl_1,
    G29_p_spl_
  );


  buf

  (
    G29_p_spl_10,
    G29_p_spl_1
  );


  buf

  (
    G29_p_spl_100,
    G29_p_spl_10
  );


  buf

  (
    G29_p_spl_101,
    G29_p_spl_10
  );


  buf

  (
    G29_p_spl_11,
    G29_p_spl_1
  );


  buf

  (
    G29_p_spl_110,
    G29_p_spl_11
  );


  buf

  (
    G29_p_spl_111,
    G29_p_spl_11
  );


  buf

  (
    G29_n_spl_,
    G29_n
  );


  buf

  (
    G29_n_spl_0,
    G29_n_spl_
  );


  buf

  (
    G29_n_spl_00,
    G29_n_spl_0
  );


  buf

  (
    G29_n_spl_000,
    G29_n_spl_00
  );


  buf

  (
    G29_n_spl_001,
    G29_n_spl_00
  );


  buf

  (
    G29_n_spl_01,
    G29_n_spl_0
  );


  buf

  (
    G29_n_spl_010,
    G29_n_spl_01
  );


  buf

  (
    G29_n_spl_011,
    G29_n_spl_01
  );


  buf

  (
    G29_n_spl_1,
    G29_n_spl_
  );


  buf

  (
    G29_n_spl_10,
    G29_n_spl_1
  );


  buf

  (
    G29_n_spl_100,
    G29_n_spl_10
  );


  buf

  (
    G29_n_spl_101,
    G29_n_spl_10
  );


  buf

  (
    G29_n_spl_11,
    G29_n_spl_1
  );


  buf

  (
    G29_n_spl_110,
    G29_n_spl_11
  );


  buf

  (
    G29_n_spl_111,
    G29_n_spl_11
  );


  buf

  (
    G13_p_spl_,
    G13_p
  );


  buf

  (
    G13_p_spl_0,
    G13_p_spl_
  );


  buf

  (
    G13_p_spl_00,
    G13_p_spl_0
  );


  buf

  (
    G13_p_spl_000,
    G13_p_spl_00
  );


  buf

  (
    G13_p_spl_001,
    G13_p_spl_00
  );


  buf

  (
    G13_p_spl_01,
    G13_p_spl_0
  );


  buf

  (
    G13_p_spl_010,
    G13_p_spl_01
  );


  buf

  (
    G13_p_spl_011,
    G13_p_spl_01
  );


  buf

  (
    G13_p_spl_1,
    G13_p_spl_
  );


  buf

  (
    G13_p_spl_10,
    G13_p_spl_1
  );


  buf

  (
    G13_p_spl_100,
    G13_p_spl_10
  );


  buf

  (
    G13_p_spl_101,
    G13_p_spl_10
  );


  buf

  (
    G13_p_spl_11,
    G13_p_spl_1
  );


  buf

  (
    G13_p_spl_110,
    G13_p_spl_11
  );


  buf

  (
    G13_p_spl_111,
    G13_p_spl_11
  );


  buf

  (
    G13_n_spl_,
    G13_n
  );


  buf

  (
    G13_n_spl_0,
    G13_n_spl_
  );


  buf

  (
    G13_n_spl_00,
    G13_n_spl_0
  );


  buf

  (
    G13_n_spl_000,
    G13_n_spl_00
  );


  buf

  (
    G13_n_spl_001,
    G13_n_spl_00
  );


  buf

  (
    G13_n_spl_01,
    G13_n_spl_0
  );


  buf

  (
    G13_n_spl_010,
    G13_n_spl_01
  );


  buf

  (
    G13_n_spl_011,
    G13_n_spl_01
  );


  buf

  (
    G13_n_spl_1,
    G13_n_spl_
  );


  buf

  (
    G13_n_spl_10,
    G13_n_spl_1
  );


  buf

  (
    G13_n_spl_100,
    G13_n_spl_10
  );


  buf

  (
    G13_n_spl_101,
    G13_n_spl_10
  );


  buf

  (
    G13_n_spl_11,
    G13_n_spl_1
  );


  buf

  (
    G13_n_spl_110,
    G13_n_spl_11
  );


  buf

  (
    G13_n_spl_111,
    G13_n_spl_11
  );


  buf

  (
    g551_p_spl_,
    g551_p
  );


  buf

  (
    g552_n_spl_,
    g552_n
  );


  buf

  (
    g551_n_spl_,
    g551_n
  );


  buf

  (
    g552_p_spl_,
    g552_p
  );


  buf

  (
    g553_n_spl_,
    g553_n
  );


  buf

  (
    g553_p_spl_,
    g553_p
  );


  buf

  (
    g554_n_spl_,
    g554_n
  );


  buf

  (
    g554_n_spl_0,
    g554_n_spl_
  );


  buf

  (
    g554_p_spl_,
    g554_p
  );


  buf

  (
    g554_p_spl_0,
    g554_p_spl_
  );


  buf

  (
    g556_n_spl_,
    g556_n
  );


  buf

  (
    g556_p_spl_,
    g556_p
  );


  buf

  (
    g557_n_spl_,
    g557_n
  );


  buf

  (
    g557_p_spl_,
    g557_p
  );


  buf

  (
    g550_n_spl_,
    g550_n
  );


  buf

  (
    g559_p_spl_,
    g559_p
  );


  buf

  (
    g550_p_spl_,
    g550_p
  );


  buf

  (
    g559_n_spl_,
    g559_n
  );


  buf

  (
    g560_n_spl_,
    g560_n
  );


  buf

  (
    g560_p_spl_,
    g560_p
  );


  buf

  (
    g549_n_spl_,
    g549_n
  );


  buf

  (
    g562_p_spl_,
    g562_p
  );


  buf

  (
    g549_p_spl_,
    g549_p
  );


  buf

  (
    g562_n_spl_,
    g562_n
  );


  buf

  (
    g563_n_spl_,
    g563_n
  );


  buf

  (
    g563_p_spl_,
    g563_p
  );


  buf

  (
    g548_n_spl_,
    g548_n
  );


  buf

  (
    g565_p_spl_,
    g565_p
  );


  buf

  (
    g548_p_spl_,
    g548_p
  );


  buf

  (
    g565_n_spl_,
    g565_n
  );


  buf

  (
    g566_n_spl_,
    g566_n
  );


  buf

  (
    g566_p_spl_,
    g566_p
  );


  buf

  (
    g547_n_spl_,
    g547_n
  );


  buf

  (
    g568_p_spl_,
    g568_p
  );


  buf

  (
    g547_p_spl_,
    g547_p
  );


  buf

  (
    g568_n_spl_,
    g568_n
  );


  buf

  (
    g569_n_spl_,
    g569_n
  );


  buf

  (
    g569_p_spl_,
    g569_p
  );


  buf

  (
    g546_n_spl_,
    g546_n
  );


  buf

  (
    g571_p_spl_,
    g571_p
  );


  buf

  (
    g546_p_spl_,
    g546_p
  );


  buf

  (
    g571_n_spl_,
    g571_n
  );


  buf

  (
    g572_n_spl_,
    g572_n
  );


  buf

  (
    g572_p_spl_,
    g572_p
  );


  buf

  (
    g545_n_spl_,
    g545_n
  );


  buf

  (
    g574_p_spl_,
    g574_p
  );


  buf

  (
    g545_p_spl_,
    g545_p
  );


  buf

  (
    g574_n_spl_,
    g574_n
  );


  buf

  (
    g575_n_spl_,
    g575_n
  );


  buf

  (
    g575_p_spl_,
    g575_p
  );


  buf

  (
    g544_n_spl_,
    g544_n
  );


  buf

  (
    g577_p_spl_,
    g577_p
  );


  buf

  (
    g544_p_spl_,
    g544_p
  );


  buf

  (
    g577_n_spl_,
    g577_n
  );


  buf

  (
    g578_n_spl_,
    g578_n
  );


  buf

  (
    g578_p_spl_,
    g578_p
  );


  buf

  (
    g543_n_spl_,
    g543_n
  );


  buf

  (
    g580_p_spl_,
    g580_p
  );


  buf

  (
    g543_p_spl_,
    g543_p
  );


  buf

  (
    g580_n_spl_,
    g580_n
  );


  buf

  (
    g581_n_spl_,
    g581_n
  );


  buf

  (
    g581_p_spl_,
    g581_p
  );


  buf

  (
    g542_n_spl_,
    g542_n
  );


  buf

  (
    g583_p_spl_,
    g583_p
  );


  buf

  (
    g542_p_spl_,
    g542_p
  );


  buf

  (
    g583_n_spl_,
    g583_n
  );


  buf

  (
    g584_n_spl_,
    g584_n
  );


  buf

  (
    g584_p_spl_,
    g584_p
  );


  buf

  (
    g541_n_spl_,
    g541_n
  );


  buf

  (
    g586_p_spl_,
    g586_p
  );


  buf

  (
    g541_p_spl_,
    g541_p
  );


  buf

  (
    g586_n_spl_,
    g586_n
  );


  buf

  (
    g587_n_spl_,
    g587_n
  );


  buf

  (
    g587_p_spl_,
    g587_p
  );


  buf

  (
    g540_n_spl_,
    g540_n
  );


  buf

  (
    g589_p_spl_,
    g589_p
  );


  buf

  (
    g540_p_spl_,
    g540_p
  );


  buf

  (
    g589_n_spl_,
    g589_n
  );


  buf

  (
    g590_n_spl_,
    g590_n
  );


  buf

  (
    g590_p_spl_,
    g590_p
  );


  buf

  (
    g539_n_spl_,
    g539_n
  );


  buf

  (
    g592_p_spl_,
    g592_p
  );


  buf

  (
    g539_p_spl_,
    g539_p
  );


  buf

  (
    g592_n_spl_,
    g592_n
  );


  buf

  (
    g593_n_spl_,
    g593_n
  );


  buf

  (
    g593_p_spl_,
    g593_p
  );


  buf

  (
    g538_n_spl_,
    g538_n
  );


  buf

  (
    g595_p_spl_,
    g595_p
  );


  buf

  (
    g538_p_spl_,
    g538_p
  );


  buf

  (
    g595_n_spl_,
    g595_n
  );


  buf

  (
    g596_n_spl_,
    g596_n
  );


  buf

  (
    g596_p_spl_,
    g596_p
  );


  buf

  (
    g537_n_spl_,
    g537_n
  );


  buf

  (
    g598_p_spl_,
    g598_p
  );


  buf

  (
    g537_p_spl_,
    g537_p
  );


  buf

  (
    g598_n_spl_,
    g598_n
  );


  buf

  (
    g599_n_spl_,
    g599_n
  );


  buf

  (
    g599_p_spl_,
    g599_p
  );


  buf

  (
    g536_n_spl_,
    g536_n
  );


  buf

  (
    g601_p_spl_,
    g601_p
  );


  buf

  (
    g536_p_spl_,
    g536_p
  );


  buf

  (
    g601_n_spl_,
    g601_n
  );


  buf

  (
    g602_n_spl_,
    g602_n
  );


  buf

  (
    g602_p_spl_,
    g602_p
  );


  buf

  (
    g535_n_spl_,
    g535_n
  );


  buf

  (
    g604_p_spl_,
    g604_p
  );


  buf

  (
    g535_p_spl_,
    g535_p
  );


  buf

  (
    g604_n_spl_,
    g604_n
  );


  buf

  (
    g605_n_spl_,
    g605_n
  );


  buf

  (
    g605_p_spl_,
    g605_p
  );


  buf

  (
    g534_n_spl_,
    g534_n
  );


  buf

  (
    g607_p_spl_,
    g607_p
  );


  buf

  (
    g534_p_spl_,
    g534_p
  );


  buf

  (
    g607_n_spl_,
    g607_n
  );


  buf

  (
    g608_n_spl_,
    g608_n
  );


  buf

  (
    g608_p_spl_,
    g608_p
  );


  buf

  (
    g533_n_spl_,
    g533_n
  );


  buf

  (
    g610_p_spl_,
    g610_p
  );


  buf

  (
    g533_p_spl_,
    g533_p
  );


  buf

  (
    g610_n_spl_,
    g610_n
  );


  buf

  (
    g611_n_spl_,
    g611_n
  );


  buf

  (
    g611_p_spl_,
    g611_p
  );


  buf

  (
    g532_n_spl_,
    g532_n
  );


  buf

  (
    g613_p_spl_,
    g613_p
  );


  buf

  (
    g532_p_spl_,
    g532_p
  );


  buf

  (
    g613_n_spl_,
    g613_n
  );


  buf

  (
    g614_n_spl_,
    g614_n
  );


  buf

  (
    g614_p_spl_,
    g614_p
  );


  buf

  (
    g531_n_spl_,
    g531_n
  );


  buf

  (
    g616_p_spl_,
    g616_p
  );


  buf

  (
    g531_p_spl_,
    g531_p
  );


  buf

  (
    g616_n_spl_,
    g616_n
  );


  buf

  (
    g617_n_spl_,
    g617_n
  );


  buf

  (
    g617_p_spl_,
    g617_p
  );


  buf

  (
    g530_p_spl_,
    g530_p
  );


  buf

  (
    g619_n_spl_,
    g619_n
  );


  buf

  (
    g620_p_spl_,
    g620_p
  );


  buf

  (
    G30_p_spl_,
    G30_p
  );


  buf

  (
    G30_p_spl_0,
    G30_p_spl_
  );


  buf

  (
    G30_p_spl_00,
    G30_p_spl_0
  );


  buf

  (
    G30_p_spl_000,
    G30_p_spl_00
  );


  buf

  (
    G30_p_spl_001,
    G30_p_spl_00
  );


  buf

  (
    G30_p_spl_01,
    G30_p_spl_0
  );


  buf

  (
    G30_p_spl_010,
    G30_p_spl_01
  );


  buf

  (
    G30_p_spl_011,
    G30_p_spl_01
  );


  buf

  (
    G30_p_spl_1,
    G30_p_spl_
  );


  buf

  (
    G30_p_spl_10,
    G30_p_spl_1
  );


  buf

  (
    G30_p_spl_100,
    G30_p_spl_10
  );


  buf

  (
    G30_p_spl_101,
    G30_p_spl_10
  );


  buf

  (
    G30_p_spl_11,
    G30_p_spl_1
  );


  buf

  (
    G30_p_spl_110,
    G30_p_spl_11
  );


  buf

  (
    G30_p_spl_111,
    G30_p_spl_11
  );


  buf

  (
    G30_n_spl_,
    G30_n
  );


  buf

  (
    G30_n_spl_0,
    G30_n_spl_
  );


  buf

  (
    G30_n_spl_00,
    G30_n_spl_0
  );


  buf

  (
    G30_n_spl_000,
    G30_n_spl_00
  );


  buf

  (
    G30_n_spl_001,
    G30_n_spl_00
  );


  buf

  (
    G30_n_spl_01,
    G30_n_spl_0
  );


  buf

  (
    G30_n_spl_010,
    G30_n_spl_01
  );


  buf

  (
    G30_n_spl_011,
    G30_n_spl_01
  );


  buf

  (
    G30_n_spl_1,
    G30_n_spl_
  );


  buf

  (
    G30_n_spl_10,
    G30_n_spl_1
  );


  buf

  (
    G30_n_spl_100,
    G30_n_spl_10
  );


  buf

  (
    G30_n_spl_101,
    G30_n_spl_10
  );


  buf

  (
    G30_n_spl_11,
    G30_n_spl_1
  );


  buf

  (
    G30_n_spl_110,
    G30_n_spl_11
  );


  buf

  (
    G30_n_spl_111,
    G30_n_spl_11
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G14_p_spl_0,
    G14_p_spl_
  );


  buf

  (
    G14_p_spl_00,
    G14_p_spl_0
  );


  buf

  (
    G14_p_spl_000,
    G14_p_spl_00
  );


  buf

  (
    G14_p_spl_001,
    G14_p_spl_00
  );


  buf

  (
    G14_p_spl_01,
    G14_p_spl_0
  );


  buf

  (
    G14_p_spl_010,
    G14_p_spl_01
  );


  buf

  (
    G14_p_spl_011,
    G14_p_spl_01
  );


  buf

  (
    G14_p_spl_1,
    G14_p_spl_
  );


  buf

  (
    G14_p_spl_10,
    G14_p_spl_1
  );


  buf

  (
    G14_p_spl_100,
    G14_p_spl_10
  );


  buf

  (
    G14_p_spl_101,
    G14_p_spl_10
  );


  buf

  (
    G14_p_spl_11,
    G14_p_spl_1
  );


  buf

  (
    G14_p_spl_110,
    G14_p_spl_11
  );


  buf

  (
    G14_p_spl_111,
    G14_p_spl_11
  );


  buf

  (
    G14_n_spl_,
    G14_n
  );


  buf

  (
    G14_n_spl_0,
    G14_n_spl_
  );


  buf

  (
    G14_n_spl_00,
    G14_n_spl_0
  );


  buf

  (
    G14_n_spl_000,
    G14_n_spl_00
  );


  buf

  (
    G14_n_spl_001,
    G14_n_spl_00
  );


  buf

  (
    G14_n_spl_01,
    G14_n_spl_0
  );


  buf

  (
    G14_n_spl_010,
    G14_n_spl_01
  );


  buf

  (
    G14_n_spl_011,
    G14_n_spl_01
  );


  buf

  (
    G14_n_spl_1,
    G14_n_spl_
  );


  buf

  (
    G14_n_spl_10,
    G14_n_spl_1
  );


  buf

  (
    G14_n_spl_100,
    G14_n_spl_10
  );


  buf

  (
    G14_n_spl_101,
    G14_n_spl_10
  );


  buf

  (
    G14_n_spl_11,
    G14_n_spl_1
  );


  buf

  (
    G14_n_spl_110,
    G14_n_spl_11
  );


  buf

  (
    G14_n_spl_111,
    G14_n_spl_11
  );


  buf

  (
    g646_p_spl_,
    g646_p
  );


  buf

  (
    g647_n_spl_,
    g647_n
  );


  buf

  (
    g646_n_spl_,
    g646_n
  );


  buf

  (
    g647_p_spl_,
    g647_p
  );


  buf

  (
    g648_n_spl_,
    g648_n
  );


  buf

  (
    g648_p_spl_,
    g648_p
  );


  buf

  (
    g649_n_spl_,
    g649_n
  );


  buf

  (
    g649_n_spl_0,
    g649_n_spl_
  );


  buf

  (
    g649_p_spl_,
    g649_p
  );


  buf

  (
    g649_p_spl_0,
    g649_p_spl_
  );


  buf

  (
    g651_n_spl_,
    g651_n
  );


  buf

  (
    g651_p_spl_,
    g651_p
  );


  buf

  (
    g652_n_spl_,
    g652_n
  );


  buf

  (
    g652_p_spl_,
    g652_p
  );


  buf

  (
    g645_n_spl_,
    g645_n
  );


  buf

  (
    g654_p_spl_,
    g654_p
  );


  buf

  (
    g645_p_spl_,
    g645_p
  );


  buf

  (
    g654_n_spl_,
    g654_n
  );


  buf

  (
    g655_n_spl_,
    g655_n
  );


  buf

  (
    g655_p_spl_,
    g655_p
  );


  buf

  (
    g644_n_spl_,
    g644_n
  );


  buf

  (
    g657_p_spl_,
    g657_p
  );


  buf

  (
    g644_p_spl_,
    g644_p
  );


  buf

  (
    g657_n_spl_,
    g657_n
  );


  buf

  (
    g658_n_spl_,
    g658_n
  );


  buf

  (
    g658_p_spl_,
    g658_p
  );


  buf

  (
    g643_n_spl_,
    g643_n
  );


  buf

  (
    g660_p_spl_,
    g660_p
  );


  buf

  (
    g643_p_spl_,
    g643_p
  );


  buf

  (
    g660_n_spl_,
    g660_n
  );


  buf

  (
    g661_n_spl_,
    g661_n
  );


  buf

  (
    g661_p_spl_,
    g661_p
  );


  buf

  (
    g642_n_spl_,
    g642_n
  );


  buf

  (
    g663_p_spl_,
    g663_p
  );


  buf

  (
    g642_p_spl_,
    g642_p
  );


  buf

  (
    g663_n_spl_,
    g663_n
  );


  buf

  (
    g664_n_spl_,
    g664_n
  );


  buf

  (
    g664_p_spl_,
    g664_p
  );


  buf

  (
    g641_n_spl_,
    g641_n
  );


  buf

  (
    g666_p_spl_,
    g666_p
  );


  buf

  (
    g641_p_spl_,
    g641_p
  );


  buf

  (
    g666_n_spl_,
    g666_n
  );


  buf

  (
    g667_n_spl_,
    g667_n
  );


  buf

  (
    g667_p_spl_,
    g667_p
  );


  buf

  (
    g640_n_spl_,
    g640_n
  );


  buf

  (
    g669_p_spl_,
    g669_p
  );


  buf

  (
    g640_p_spl_,
    g640_p
  );


  buf

  (
    g669_n_spl_,
    g669_n
  );


  buf

  (
    g670_n_spl_,
    g670_n
  );


  buf

  (
    g670_p_spl_,
    g670_p
  );


  buf

  (
    g639_n_spl_,
    g639_n
  );


  buf

  (
    g672_p_spl_,
    g672_p
  );


  buf

  (
    g639_p_spl_,
    g639_p
  );


  buf

  (
    g672_n_spl_,
    g672_n
  );


  buf

  (
    g673_n_spl_,
    g673_n
  );


  buf

  (
    g673_p_spl_,
    g673_p
  );


  buf

  (
    g638_n_spl_,
    g638_n
  );


  buf

  (
    g675_p_spl_,
    g675_p
  );


  buf

  (
    g638_p_spl_,
    g638_p
  );


  buf

  (
    g675_n_spl_,
    g675_n
  );


  buf

  (
    g676_n_spl_,
    g676_n
  );


  buf

  (
    g676_p_spl_,
    g676_p
  );


  buf

  (
    g637_n_spl_,
    g637_n
  );


  buf

  (
    g678_p_spl_,
    g678_p
  );


  buf

  (
    g637_p_spl_,
    g637_p
  );


  buf

  (
    g678_n_spl_,
    g678_n
  );


  buf

  (
    g679_n_spl_,
    g679_n
  );


  buf

  (
    g679_p_spl_,
    g679_p
  );


  buf

  (
    g636_n_spl_,
    g636_n
  );


  buf

  (
    g681_p_spl_,
    g681_p
  );


  buf

  (
    g636_p_spl_,
    g636_p
  );


  buf

  (
    g681_n_spl_,
    g681_n
  );


  buf

  (
    g682_n_spl_,
    g682_n
  );


  buf

  (
    g682_p_spl_,
    g682_p
  );


  buf

  (
    g635_n_spl_,
    g635_n
  );


  buf

  (
    g684_p_spl_,
    g684_p
  );


  buf

  (
    g635_p_spl_,
    g635_p
  );


  buf

  (
    g684_n_spl_,
    g684_n
  );


  buf

  (
    g685_n_spl_,
    g685_n
  );


  buf

  (
    g685_p_spl_,
    g685_p
  );


  buf

  (
    g634_n_spl_,
    g634_n
  );


  buf

  (
    g687_p_spl_,
    g687_p
  );


  buf

  (
    g634_p_spl_,
    g634_p
  );


  buf

  (
    g687_n_spl_,
    g687_n
  );


  buf

  (
    g688_n_spl_,
    g688_n
  );


  buf

  (
    g688_p_spl_,
    g688_p
  );


  buf

  (
    g633_n_spl_,
    g633_n
  );


  buf

  (
    g690_p_spl_,
    g690_p
  );


  buf

  (
    g633_p_spl_,
    g633_p
  );


  buf

  (
    g690_n_spl_,
    g690_n
  );


  buf

  (
    g691_n_spl_,
    g691_n
  );


  buf

  (
    g691_p_spl_,
    g691_p
  );


  buf

  (
    g632_n_spl_,
    g632_n
  );


  buf

  (
    g693_p_spl_,
    g693_p
  );


  buf

  (
    g632_p_spl_,
    g632_p
  );


  buf

  (
    g693_n_spl_,
    g693_n
  );


  buf

  (
    g694_n_spl_,
    g694_n
  );


  buf

  (
    g694_p_spl_,
    g694_p
  );


  buf

  (
    g631_n_spl_,
    g631_n
  );


  buf

  (
    g696_p_spl_,
    g696_p
  );


  buf

  (
    g631_p_spl_,
    g631_p
  );


  buf

  (
    g696_n_spl_,
    g696_n
  );


  buf

  (
    g697_n_spl_,
    g697_n
  );


  buf

  (
    g697_p_spl_,
    g697_p
  );


  buf

  (
    g630_n_spl_,
    g630_n
  );


  buf

  (
    g699_p_spl_,
    g699_p
  );


  buf

  (
    g630_p_spl_,
    g630_p
  );


  buf

  (
    g699_n_spl_,
    g699_n
  );


  buf

  (
    g700_n_spl_,
    g700_n
  );


  buf

  (
    g700_p_spl_,
    g700_p
  );


  buf

  (
    g629_n_spl_,
    g629_n
  );


  buf

  (
    g702_p_spl_,
    g702_p
  );


  buf

  (
    g629_p_spl_,
    g629_p
  );


  buf

  (
    g702_n_spl_,
    g702_n
  );


  buf

  (
    g703_n_spl_,
    g703_n
  );


  buf

  (
    g703_p_spl_,
    g703_p
  );


  buf

  (
    g628_n_spl_,
    g628_n
  );


  buf

  (
    g705_p_spl_,
    g705_p
  );


  buf

  (
    g628_p_spl_,
    g628_p
  );


  buf

  (
    g705_n_spl_,
    g705_n
  );


  buf

  (
    g706_n_spl_,
    g706_n
  );


  buf

  (
    g706_p_spl_,
    g706_p
  );


  buf

  (
    g627_n_spl_,
    g627_n
  );


  buf

  (
    g708_p_spl_,
    g708_p
  );


  buf

  (
    g627_p_spl_,
    g627_p
  );


  buf

  (
    g708_n_spl_,
    g708_n
  );


  buf

  (
    g709_n_spl_,
    g709_n
  );


  buf

  (
    g709_p_spl_,
    g709_p
  );


  buf

  (
    g626_n_spl_,
    g626_n
  );


  buf

  (
    g711_p_spl_,
    g711_p
  );


  buf

  (
    g626_p_spl_,
    g626_p
  );


  buf

  (
    g711_n_spl_,
    g711_n
  );


  buf

  (
    g712_n_spl_,
    g712_n
  );


  buf

  (
    g712_p_spl_,
    g712_p
  );


  buf

  (
    g625_n_spl_,
    g625_n
  );


  buf

  (
    g714_p_spl_,
    g714_p
  );


  buf

  (
    g625_p_spl_,
    g625_p
  );


  buf

  (
    g714_n_spl_,
    g714_n
  );


  buf

  (
    g715_n_spl_,
    g715_n
  );


  buf

  (
    g715_p_spl_,
    g715_p
  );


  buf

  (
    g624_n_spl_,
    g624_n
  );


  buf

  (
    g717_p_spl_,
    g717_p
  );


  buf

  (
    g624_p_spl_,
    g624_p
  );


  buf

  (
    g717_n_spl_,
    g717_n
  );


  buf

  (
    g718_n_spl_,
    g718_n
  );


  buf

  (
    g718_p_spl_,
    g718_p
  );


  buf

  (
    g623_p_spl_,
    g623_p
  );


  buf

  (
    g720_n_spl_,
    g720_n
  );


  buf

  (
    g721_p_spl_,
    g721_p
  );


  buf

  (
    G31_p_spl_,
    G31_p
  );


  buf

  (
    G31_p_spl_0,
    G31_p_spl_
  );


  buf

  (
    G31_p_spl_00,
    G31_p_spl_0
  );


  buf

  (
    G31_p_spl_000,
    G31_p_spl_00
  );


  buf

  (
    G31_p_spl_001,
    G31_p_spl_00
  );


  buf

  (
    G31_p_spl_01,
    G31_p_spl_0
  );


  buf

  (
    G31_p_spl_010,
    G31_p_spl_01
  );


  buf

  (
    G31_p_spl_011,
    G31_p_spl_01
  );


  buf

  (
    G31_p_spl_1,
    G31_p_spl_
  );


  buf

  (
    G31_p_spl_10,
    G31_p_spl_1
  );


  buf

  (
    G31_p_spl_100,
    G31_p_spl_10
  );


  buf

  (
    G31_p_spl_101,
    G31_p_spl_10
  );


  buf

  (
    G31_p_spl_11,
    G31_p_spl_1
  );


  buf

  (
    G31_p_spl_110,
    G31_p_spl_11
  );


  buf

  (
    G31_p_spl_111,
    G31_p_spl_11
  );


  buf

  (
    G31_n_spl_,
    G31_n
  );


  buf

  (
    G31_n_spl_0,
    G31_n_spl_
  );


  buf

  (
    G31_n_spl_00,
    G31_n_spl_0
  );


  buf

  (
    G31_n_spl_000,
    G31_n_spl_00
  );


  buf

  (
    G31_n_spl_001,
    G31_n_spl_00
  );


  buf

  (
    G31_n_spl_01,
    G31_n_spl_0
  );


  buf

  (
    G31_n_spl_010,
    G31_n_spl_01
  );


  buf

  (
    G31_n_spl_011,
    G31_n_spl_01
  );


  buf

  (
    G31_n_spl_1,
    G31_n_spl_
  );


  buf

  (
    G31_n_spl_10,
    G31_n_spl_1
  );


  buf

  (
    G31_n_spl_100,
    G31_n_spl_10
  );


  buf

  (
    G31_n_spl_101,
    G31_n_spl_10
  );


  buf

  (
    G31_n_spl_11,
    G31_n_spl_1
  );


  buf

  (
    G31_n_spl_110,
    G31_n_spl_11
  );


  buf

  (
    G31_n_spl_111,
    G31_n_spl_11
  );


  buf

  (
    G15_p_spl_,
    G15_p
  );


  buf

  (
    G15_p_spl_0,
    G15_p_spl_
  );


  buf

  (
    G15_p_spl_00,
    G15_p_spl_0
  );


  buf

  (
    G15_p_spl_000,
    G15_p_spl_00
  );


  buf

  (
    G15_p_spl_001,
    G15_p_spl_00
  );


  buf

  (
    G15_p_spl_01,
    G15_p_spl_0
  );


  buf

  (
    G15_p_spl_010,
    G15_p_spl_01
  );


  buf

  (
    G15_p_spl_011,
    G15_p_spl_01
  );


  buf

  (
    G15_p_spl_1,
    G15_p_spl_
  );


  buf

  (
    G15_p_spl_10,
    G15_p_spl_1
  );


  buf

  (
    G15_p_spl_100,
    G15_p_spl_10
  );


  buf

  (
    G15_p_spl_101,
    G15_p_spl_10
  );


  buf

  (
    G15_p_spl_11,
    G15_p_spl_1
  );


  buf

  (
    G15_p_spl_110,
    G15_p_spl_11
  );


  buf

  (
    G15_p_spl_111,
    G15_p_spl_11
  );


  buf

  (
    G15_n_spl_,
    G15_n
  );


  buf

  (
    G15_n_spl_0,
    G15_n_spl_
  );


  buf

  (
    G15_n_spl_00,
    G15_n_spl_0
  );


  buf

  (
    G15_n_spl_000,
    G15_n_spl_00
  );


  buf

  (
    G15_n_spl_001,
    G15_n_spl_00
  );


  buf

  (
    G15_n_spl_01,
    G15_n_spl_0
  );


  buf

  (
    G15_n_spl_010,
    G15_n_spl_01
  );


  buf

  (
    G15_n_spl_011,
    G15_n_spl_01
  );


  buf

  (
    G15_n_spl_1,
    G15_n_spl_
  );


  buf

  (
    G15_n_spl_10,
    G15_n_spl_1
  );


  buf

  (
    G15_n_spl_100,
    G15_n_spl_10
  );


  buf

  (
    G15_n_spl_101,
    G15_n_spl_10
  );


  buf

  (
    G15_n_spl_11,
    G15_n_spl_1
  );


  buf

  (
    G15_n_spl_110,
    G15_n_spl_11
  );


  buf

  (
    G15_n_spl_111,
    G15_n_spl_11
  );


  buf

  (
    g749_p_spl_,
    g749_p
  );


  buf

  (
    g750_n_spl_,
    g750_n
  );


  buf

  (
    g749_n_spl_,
    g749_n
  );


  buf

  (
    g750_p_spl_,
    g750_p
  );


  buf

  (
    g751_n_spl_,
    g751_n
  );


  buf

  (
    g751_p_spl_,
    g751_p
  );


  buf

  (
    g752_n_spl_,
    g752_n
  );


  buf

  (
    g752_n_spl_0,
    g752_n_spl_
  );


  buf

  (
    g752_p_spl_,
    g752_p
  );


  buf

  (
    g752_p_spl_0,
    g752_p_spl_
  );


  buf

  (
    g754_n_spl_,
    g754_n
  );


  buf

  (
    g754_p_spl_,
    g754_p
  );


  buf

  (
    g755_n_spl_,
    g755_n
  );


  buf

  (
    g755_p_spl_,
    g755_p
  );


  buf

  (
    g748_n_spl_,
    g748_n
  );


  buf

  (
    g757_p_spl_,
    g757_p
  );


  buf

  (
    g748_p_spl_,
    g748_p
  );


  buf

  (
    g757_n_spl_,
    g757_n
  );


  buf

  (
    g758_n_spl_,
    g758_n
  );


  buf

  (
    g758_p_spl_,
    g758_p
  );


  buf

  (
    g747_n_spl_,
    g747_n
  );


  buf

  (
    g760_p_spl_,
    g760_p
  );


  buf

  (
    g747_p_spl_,
    g747_p
  );


  buf

  (
    g760_n_spl_,
    g760_n
  );


  buf

  (
    g761_n_spl_,
    g761_n
  );


  buf

  (
    g761_p_spl_,
    g761_p
  );


  buf

  (
    g746_n_spl_,
    g746_n
  );


  buf

  (
    g763_p_spl_,
    g763_p
  );


  buf

  (
    g746_p_spl_,
    g746_p
  );


  buf

  (
    g763_n_spl_,
    g763_n
  );


  buf

  (
    g764_n_spl_,
    g764_n
  );


  buf

  (
    g764_p_spl_,
    g764_p
  );


  buf

  (
    g745_n_spl_,
    g745_n
  );


  buf

  (
    g766_p_spl_,
    g766_p
  );


  buf

  (
    g745_p_spl_,
    g745_p
  );


  buf

  (
    g766_n_spl_,
    g766_n
  );


  buf

  (
    g767_n_spl_,
    g767_n
  );


  buf

  (
    g767_p_spl_,
    g767_p
  );


  buf

  (
    g744_n_spl_,
    g744_n
  );


  buf

  (
    g769_p_spl_,
    g769_p
  );


  buf

  (
    g744_p_spl_,
    g744_p
  );


  buf

  (
    g769_n_spl_,
    g769_n
  );


  buf

  (
    g770_n_spl_,
    g770_n
  );


  buf

  (
    g770_p_spl_,
    g770_p
  );


  buf

  (
    g743_n_spl_,
    g743_n
  );


  buf

  (
    g772_p_spl_,
    g772_p
  );


  buf

  (
    g743_p_spl_,
    g743_p
  );


  buf

  (
    g772_n_spl_,
    g772_n
  );


  buf

  (
    g773_n_spl_,
    g773_n
  );


  buf

  (
    g773_p_spl_,
    g773_p
  );


  buf

  (
    g742_n_spl_,
    g742_n
  );


  buf

  (
    g775_p_spl_,
    g775_p
  );


  buf

  (
    g742_p_spl_,
    g742_p
  );


  buf

  (
    g775_n_spl_,
    g775_n
  );


  buf

  (
    g776_n_spl_,
    g776_n
  );


  buf

  (
    g776_p_spl_,
    g776_p
  );


  buf

  (
    g741_n_spl_,
    g741_n
  );


  buf

  (
    g778_p_spl_,
    g778_p
  );


  buf

  (
    g741_p_spl_,
    g741_p
  );


  buf

  (
    g778_n_spl_,
    g778_n
  );


  buf

  (
    g779_n_spl_,
    g779_n
  );


  buf

  (
    g779_p_spl_,
    g779_p
  );


  buf

  (
    g740_n_spl_,
    g740_n
  );


  buf

  (
    g781_p_spl_,
    g781_p
  );


  buf

  (
    g740_p_spl_,
    g740_p
  );


  buf

  (
    g781_n_spl_,
    g781_n
  );


  buf

  (
    g782_n_spl_,
    g782_n
  );


  buf

  (
    g782_p_spl_,
    g782_p
  );


  buf

  (
    g739_n_spl_,
    g739_n
  );


  buf

  (
    g784_p_spl_,
    g784_p
  );


  buf

  (
    g739_p_spl_,
    g739_p
  );


  buf

  (
    g784_n_spl_,
    g784_n
  );


  buf

  (
    g785_n_spl_,
    g785_n
  );


  buf

  (
    g785_p_spl_,
    g785_p
  );


  buf

  (
    g738_n_spl_,
    g738_n
  );


  buf

  (
    g787_p_spl_,
    g787_p
  );


  buf

  (
    g738_p_spl_,
    g738_p
  );


  buf

  (
    g787_n_spl_,
    g787_n
  );


  buf

  (
    g788_n_spl_,
    g788_n
  );


  buf

  (
    g788_p_spl_,
    g788_p
  );


  buf

  (
    g737_n_spl_,
    g737_n
  );


  buf

  (
    g790_p_spl_,
    g790_p
  );


  buf

  (
    g737_p_spl_,
    g737_p
  );


  buf

  (
    g790_n_spl_,
    g790_n
  );


  buf

  (
    g791_n_spl_,
    g791_n
  );


  buf

  (
    g791_p_spl_,
    g791_p
  );


  buf

  (
    g736_n_spl_,
    g736_n
  );


  buf

  (
    g793_p_spl_,
    g793_p
  );


  buf

  (
    g736_p_spl_,
    g736_p
  );


  buf

  (
    g793_n_spl_,
    g793_n
  );


  buf

  (
    g794_n_spl_,
    g794_n
  );


  buf

  (
    g794_p_spl_,
    g794_p
  );


  buf

  (
    g735_n_spl_,
    g735_n
  );


  buf

  (
    g796_p_spl_,
    g796_p
  );


  buf

  (
    g735_p_spl_,
    g735_p
  );


  buf

  (
    g796_n_spl_,
    g796_n
  );


  buf

  (
    g797_n_spl_,
    g797_n
  );


  buf

  (
    g797_p_spl_,
    g797_p
  );


  buf

  (
    g734_n_spl_,
    g734_n
  );


  buf

  (
    g799_p_spl_,
    g799_p
  );


  buf

  (
    g734_p_spl_,
    g734_p
  );


  buf

  (
    g799_n_spl_,
    g799_n
  );


  buf

  (
    g800_n_spl_,
    g800_n
  );


  buf

  (
    g800_p_spl_,
    g800_p
  );


  buf

  (
    g733_n_spl_,
    g733_n
  );


  buf

  (
    g802_p_spl_,
    g802_p
  );


  buf

  (
    g733_p_spl_,
    g733_p
  );


  buf

  (
    g802_n_spl_,
    g802_n
  );


  buf

  (
    g803_n_spl_,
    g803_n
  );


  buf

  (
    g803_p_spl_,
    g803_p
  );


  buf

  (
    g732_n_spl_,
    g732_n
  );


  buf

  (
    g805_p_spl_,
    g805_p
  );


  buf

  (
    g732_p_spl_,
    g732_p
  );


  buf

  (
    g805_n_spl_,
    g805_n
  );


  buf

  (
    g806_n_spl_,
    g806_n
  );


  buf

  (
    g806_p_spl_,
    g806_p
  );


  buf

  (
    g731_n_spl_,
    g731_n
  );


  buf

  (
    g808_p_spl_,
    g808_p
  );


  buf

  (
    g731_p_spl_,
    g731_p
  );


  buf

  (
    g808_n_spl_,
    g808_n
  );


  buf

  (
    g809_n_spl_,
    g809_n
  );


  buf

  (
    g809_p_spl_,
    g809_p
  );


  buf

  (
    g730_n_spl_,
    g730_n
  );


  buf

  (
    g811_p_spl_,
    g811_p
  );


  buf

  (
    g730_p_spl_,
    g730_p
  );


  buf

  (
    g811_n_spl_,
    g811_n
  );


  buf

  (
    g812_n_spl_,
    g812_n
  );


  buf

  (
    g812_p_spl_,
    g812_p
  );


  buf

  (
    g729_n_spl_,
    g729_n
  );


  buf

  (
    g814_p_spl_,
    g814_p
  );


  buf

  (
    g729_p_spl_,
    g729_p
  );


  buf

  (
    g814_n_spl_,
    g814_n
  );


  buf

  (
    g815_n_spl_,
    g815_n
  );


  buf

  (
    g815_p_spl_,
    g815_p
  );


  buf

  (
    g728_n_spl_,
    g728_n
  );


  buf

  (
    g817_p_spl_,
    g817_p
  );


  buf

  (
    g728_p_spl_,
    g728_p
  );


  buf

  (
    g817_n_spl_,
    g817_n
  );


  buf

  (
    g818_n_spl_,
    g818_n
  );


  buf

  (
    g818_p_spl_,
    g818_p
  );


  buf

  (
    g727_n_spl_,
    g727_n
  );


  buf

  (
    g820_p_spl_,
    g820_p
  );


  buf

  (
    g727_p_spl_,
    g727_p
  );


  buf

  (
    g820_n_spl_,
    g820_n
  );


  buf

  (
    g821_n_spl_,
    g821_n
  );


  buf

  (
    g821_p_spl_,
    g821_p
  );


  buf

  (
    g726_n_spl_,
    g726_n
  );


  buf

  (
    g823_p_spl_,
    g823_p
  );


  buf

  (
    g726_p_spl_,
    g726_p
  );


  buf

  (
    g823_n_spl_,
    g823_n
  );


  buf

  (
    g824_n_spl_,
    g824_n
  );


  buf

  (
    g824_p_spl_,
    g824_p
  );


  buf

  (
    g725_n_spl_,
    g725_n
  );


  buf

  (
    g826_p_spl_,
    g826_p
  );


  buf

  (
    g725_p_spl_,
    g725_p
  );


  buf

  (
    g826_n_spl_,
    g826_n
  );


  buf

  (
    g827_n_spl_,
    g827_n
  );


  buf

  (
    g827_p_spl_,
    g827_p
  );


  buf

  (
    g724_p_spl_,
    g724_p
  );


  buf

  (
    g829_n_spl_,
    g829_n
  );


  buf

  (
    g830_p_spl_,
    g830_p
  );


  buf

  (
    G32_p_spl_,
    G32_p
  );


  buf

  (
    G32_p_spl_0,
    G32_p_spl_
  );


  buf

  (
    G32_p_spl_00,
    G32_p_spl_0
  );


  buf

  (
    G32_p_spl_000,
    G32_p_spl_00
  );


  buf

  (
    G32_p_spl_001,
    G32_p_spl_00
  );


  buf

  (
    G32_p_spl_01,
    G32_p_spl_0
  );


  buf

  (
    G32_p_spl_010,
    G32_p_spl_01
  );


  buf

  (
    G32_p_spl_011,
    G32_p_spl_01
  );


  buf

  (
    G32_p_spl_1,
    G32_p_spl_
  );


  buf

  (
    G32_p_spl_10,
    G32_p_spl_1
  );


  buf

  (
    G32_p_spl_100,
    G32_p_spl_10
  );


  buf

  (
    G32_p_spl_101,
    G32_p_spl_10
  );


  buf

  (
    G32_p_spl_11,
    G32_p_spl_1
  );


  buf

  (
    G32_p_spl_110,
    G32_p_spl_11
  );


  buf

  (
    G32_p_spl_111,
    G32_p_spl_11
  );


  buf

  (
    G32_n_spl_,
    G32_n
  );


  buf

  (
    G32_n_spl_0,
    G32_n_spl_
  );


  buf

  (
    G32_n_spl_00,
    G32_n_spl_0
  );


  buf

  (
    G32_n_spl_000,
    G32_n_spl_00
  );


  buf

  (
    G32_n_spl_001,
    G32_n_spl_00
  );


  buf

  (
    G32_n_spl_01,
    G32_n_spl_0
  );


  buf

  (
    G32_n_spl_010,
    G32_n_spl_01
  );


  buf

  (
    G32_n_spl_011,
    G32_n_spl_01
  );


  buf

  (
    G32_n_spl_1,
    G32_n_spl_
  );


  buf

  (
    G32_n_spl_10,
    G32_n_spl_1
  );


  buf

  (
    G32_n_spl_100,
    G32_n_spl_10
  );


  buf

  (
    G32_n_spl_101,
    G32_n_spl_10
  );


  buf

  (
    G32_n_spl_11,
    G32_n_spl_1
  );


  buf

  (
    G32_n_spl_110,
    G32_n_spl_11
  );


  buf

  (
    G32_n_spl_111,
    G32_n_spl_11
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    G16_p_spl_0,
    G16_p_spl_
  );


  buf

  (
    G16_p_spl_00,
    G16_p_spl_0
  );


  buf

  (
    G16_p_spl_000,
    G16_p_spl_00
  );


  buf

  (
    G16_p_spl_001,
    G16_p_spl_00
  );


  buf

  (
    G16_p_spl_01,
    G16_p_spl_0
  );


  buf

  (
    G16_p_spl_010,
    G16_p_spl_01
  );


  buf

  (
    G16_p_spl_011,
    G16_p_spl_01
  );


  buf

  (
    G16_p_spl_1,
    G16_p_spl_
  );


  buf

  (
    G16_p_spl_10,
    G16_p_spl_1
  );


  buf

  (
    G16_p_spl_100,
    G16_p_spl_10
  );


  buf

  (
    G16_p_spl_101,
    G16_p_spl_10
  );


  buf

  (
    G16_p_spl_11,
    G16_p_spl_1
  );


  buf

  (
    G16_p_spl_110,
    G16_p_spl_11
  );


  buf

  (
    G16_p_spl_111,
    G16_p_spl_11
  );


  buf

  (
    G16_n_spl_,
    G16_n
  );


  buf

  (
    G16_n_spl_0,
    G16_n_spl_
  );


  buf

  (
    G16_n_spl_00,
    G16_n_spl_0
  );


  buf

  (
    G16_n_spl_000,
    G16_n_spl_00
  );


  buf

  (
    G16_n_spl_001,
    G16_n_spl_00
  );


  buf

  (
    G16_n_spl_01,
    G16_n_spl_0
  );


  buf

  (
    G16_n_spl_010,
    G16_n_spl_01
  );


  buf

  (
    G16_n_spl_011,
    G16_n_spl_01
  );


  buf

  (
    G16_n_spl_1,
    G16_n_spl_
  );


  buf

  (
    G16_n_spl_10,
    G16_n_spl_1
  );


  buf

  (
    G16_n_spl_100,
    G16_n_spl_10
  );


  buf

  (
    G16_n_spl_101,
    G16_n_spl_10
  );


  buf

  (
    G16_n_spl_11,
    G16_n_spl_1
  );


  buf

  (
    G16_n_spl_110,
    G16_n_spl_11
  );


  buf

  (
    G16_n_spl_111,
    G16_n_spl_11
  );


  buf

  (
    g860_p_spl_,
    g860_p
  );


  buf

  (
    g861_n_spl_,
    g861_n
  );


  buf

  (
    g860_n_spl_,
    g860_n
  );


  buf

  (
    g861_p_spl_,
    g861_p
  );


  buf

  (
    g862_n_spl_,
    g862_n
  );


  buf

  (
    g862_p_spl_,
    g862_p
  );


  buf

  (
    g863_n_spl_,
    g863_n
  );


  buf

  (
    g863_p_spl_,
    g863_p
  );


  buf

  (
    g865_n_spl_,
    g865_n
  );


  buf

  (
    g865_p_spl_,
    g865_p
  );


  buf

  (
    g866_n_spl_,
    g866_n
  );


  buf

  (
    g866_p_spl_,
    g866_p
  );


  buf

  (
    g859_n_spl_,
    g859_n
  );


  buf

  (
    g868_p_spl_,
    g868_p
  );


  buf

  (
    g859_p_spl_,
    g859_p
  );


  buf

  (
    g868_n_spl_,
    g868_n
  );


  buf

  (
    g869_n_spl_,
    g869_n
  );


  buf

  (
    g869_p_spl_,
    g869_p
  );


  buf

  (
    g858_n_spl_,
    g858_n
  );


  buf

  (
    g871_p_spl_,
    g871_p
  );


  buf

  (
    g858_p_spl_,
    g858_p
  );


  buf

  (
    g871_n_spl_,
    g871_n
  );


  buf

  (
    g872_n_spl_,
    g872_n
  );


  buf

  (
    g872_p_spl_,
    g872_p
  );


  buf

  (
    g857_n_spl_,
    g857_n
  );


  buf

  (
    g874_p_spl_,
    g874_p
  );


  buf

  (
    g857_p_spl_,
    g857_p
  );


  buf

  (
    g874_n_spl_,
    g874_n
  );


  buf

  (
    g875_n_spl_,
    g875_n
  );


  buf

  (
    g875_p_spl_,
    g875_p
  );


  buf

  (
    g856_n_spl_,
    g856_n
  );


  buf

  (
    g877_p_spl_,
    g877_p
  );


  buf

  (
    g856_p_spl_,
    g856_p
  );


  buf

  (
    g877_n_spl_,
    g877_n
  );


  buf

  (
    g878_n_spl_,
    g878_n
  );


  buf

  (
    g878_p_spl_,
    g878_p
  );


  buf

  (
    g855_n_spl_,
    g855_n
  );


  buf

  (
    g880_p_spl_,
    g880_p
  );


  buf

  (
    g855_p_spl_,
    g855_p
  );


  buf

  (
    g880_n_spl_,
    g880_n
  );


  buf

  (
    g881_n_spl_,
    g881_n
  );


  buf

  (
    g881_p_spl_,
    g881_p
  );


  buf

  (
    g854_n_spl_,
    g854_n
  );


  buf

  (
    g883_p_spl_,
    g883_p
  );


  buf

  (
    g854_p_spl_,
    g854_p
  );


  buf

  (
    g883_n_spl_,
    g883_n
  );


  buf

  (
    g884_n_spl_,
    g884_n
  );


  buf

  (
    g884_p_spl_,
    g884_p
  );


  buf

  (
    g853_n_spl_,
    g853_n
  );


  buf

  (
    g886_p_spl_,
    g886_p
  );


  buf

  (
    g853_p_spl_,
    g853_p
  );


  buf

  (
    g886_n_spl_,
    g886_n
  );


  buf

  (
    g887_n_spl_,
    g887_n
  );


  buf

  (
    g887_p_spl_,
    g887_p
  );


  buf

  (
    g852_n_spl_,
    g852_n
  );


  buf

  (
    g889_p_spl_,
    g889_p
  );


  buf

  (
    g852_p_spl_,
    g852_p
  );


  buf

  (
    g889_n_spl_,
    g889_n
  );


  buf

  (
    g890_n_spl_,
    g890_n
  );


  buf

  (
    g890_p_spl_,
    g890_p
  );


  buf

  (
    g851_n_spl_,
    g851_n
  );


  buf

  (
    g892_p_spl_,
    g892_p
  );


  buf

  (
    g851_p_spl_,
    g851_p
  );


  buf

  (
    g892_n_spl_,
    g892_n
  );


  buf

  (
    g893_n_spl_,
    g893_n
  );


  buf

  (
    g893_p_spl_,
    g893_p
  );


  buf

  (
    g850_n_spl_,
    g850_n
  );


  buf

  (
    g895_p_spl_,
    g895_p
  );


  buf

  (
    g850_p_spl_,
    g850_p
  );


  buf

  (
    g895_n_spl_,
    g895_n
  );


  buf

  (
    g896_n_spl_,
    g896_n
  );


  buf

  (
    g896_p_spl_,
    g896_p
  );


  buf

  (
    g849_n_spl_,
    g849_n
  );


  buf

  (
    g898_p_spl_,
    g898_p
  );


  buf

  (
    g849_p_spl_,
    g849_p
  );


  buf

  (
    g898_n_spl_,
    g898_n
  );


  buf

  (
    g899_n_spl_,
    g899_n
  );


  buf

  (
    g899_p_spl_,
    g899_p
  );


  buf

  (
    g848_n_spl_,
    g848_n
  );


  buf

  (
    g901_p_spl_,
    g901_p
  );


  buf

  (
    g848_p_spl_,
    g848_p
  );


  buf

  (
    g901_n_spl_,
    g901_n
  );


  buf

  (
    g902_n_spl_,
    g902_n
  );


  buf

  (
    g902_p_spl_,
    g902_p
  );


  buf

  (
    g847_n_spl_,
    g847_n
  );


  buf

  (
    g904_p_spl_,
    g904_p
  );


  buf

  (
    g847_p_spl_,
    g847_p
  );


  buf

  (
    g904_n_spl_,
    g904_n
  );


  buf

  (
    g905_n_spl_,
    g905_n
  );


  buf

  (
    g905_p_spl_,
    g905_p
  );


  buf

  (
    g846_n_spl_,
    g846_n
  );


  buf

  (
    g907_p_spl_,
    g907_p
  );


  buf

  (
    g846_p_spl_,
    g846_p
  );


  buf

  (
    g907_n_spl_,
    g907_n
  );


  buf

  (
    g908_n_spl_,
    g908_n
  );


  buf

  (
    g908_p_spl_,
    g908_p
  );


  buf

  (
    g845_n_spl_,
    g845_n
  );


  buf

  (
    g910_p_spl_,
    g910_p
  );


  buf

  (
    g845_p_spl_,
    g845_p
  );


  buf

  (
    g910_n_spl_,
    g910_n
  );


  buf

  (
    g911_n_spl_,
    g911_n
  );


  buf

  (
    g911_p_spl_,
    g911_p
  );


  buf

  (
    g844_n_spl_,
    g844_n
  );


  buf

  (
    g913_p_spl_,
    g913_p
  );


  buf

  (
    g844_p_spl_,
    g844_p
  );


  buf

  (
    g913_n_spl_,
    g913_n
  );


  buf

  (
    g914_n_spl_,
    g914_n
  );


  buf

  (
    g914_p_spl_,
    g914_p
  );


  buf

  (
    g843_n_spl_,
    g843_n
  );


  buf

  (
    g916_p_spl_,
    g916_p
  );


  buf

  (
    g843_p_spl_,
    g843_p
  );


  buf

  (
    g916_n_spl_,
    g916_n
  );


  buf

  (
    g917_n_spl_,
    g917_n
  );


  buf

  (
    g917_p_spl_,
    g917_p
  );


  buf

  (
    g842_n_spl_,
    g842_n
  );


  buf

  (
    g919_p_spl_,
    g919_p
  );


  buf

  (
    g842_p_spl_,
    g842_p
  );


  buf

  (
    g919_n_spl_,
    g919_n
  );


  buf

  (
    g920_n_spl_,
    g920_n
  );


  buf

  (
    g920_p_spl_,
    g920_p
  );


  buf

  (
    g841_n_spl_,
    g841_n
  );


  buf

  (
    g922_p_spl_,
    g922_p
  );


  buf

  (
    g841_p_spl_,
    g841_p
  );


  buf

  (
    g922_n_spl_,
    g922_n
  );


  buf

  (
    g923_n_spl_,
    g923_n
  );


  buf

  (
    g923_p_spl_,
    g923_p
  );


  buf

  (
    g840_n_spl_,
    g840_n
  );


  buf

  (
    g925_p_spl_,
    g925_p
  );


  buf

  (
    g840_p_spl_,
    g840_p
  );


  buf

  (
    g925_n_spl_,
    g925_n
  );


  buf

  (
    g926_n_spl_,
    g926_n
  );


  buf

  (
    g926_p_spl_,
    g926_p
  );


  buf

  (
    g839_n_spl_,
    g839_n
  );


  buf

  (
    g928_p_spl_,
    g928_p
  );


  buf

  (
    g839_p_spl_,
    g839_p
  );


  buf

  (
    g928_n_spl_,
    g928_n
  );


  buf

  (
    g929_n_spl_,
    g929_n
  );


  buf

  (
    g929_p_spl_,
    g929_p
  );


  buf

  (
    g838_n_spl_,
    g838_n
  );


  buf

  (
    g931_p_spl_,
    g931_p
  );


  buf

  (
    g838_p_spl_,
    g838_p
  );


  buf

  (
    g931_n_spl_,
    g931_n
  );


  buf

  (
    g932_n_spl_,
    g932_n
  );


  buf

  (
    g932_p_spl_,
    g932_p
  );


  buf

  (
    g837_n_spl_,
    g837_n
  );


  buf

  (
    g934_p_spl_,
    g934_p
  );


  buf

  (
    g837_p_spl_,
    g837_p
  );


  buf

  (
    g934_n_spl_,
    g934_n
  );


  buf

  (
    g935_n_spl_,
    g935_n
  );


  buf

  (
    g935_p_spl_,
    g935_p
  );


  buf

  (
    g836_n_spl_,
    g836_n
  );


  buf

  (
    g937_p_spl_,
    g937_p
  );


  buf

  (
    g836_p_spl_,
    g836_p
  );


  buf

  (
    g937_n_spl_,
    g937_n
  );


  buf

  (
    g938_n_spl_,
    g938_n
  );


  buf

  (
    g938_p_spl_,
    g938_p
  );


  buf

  (
    g835_n_spl_,
    g835_n
  );


  buf

  (
    g940_p_spl_,
    g940_p
  );


  buf

  (
    g835_p_spl_,
    g835_p
  );


  buf

  (
    g940_n_spl_,
    g940_n
  );


  buf

  (
    g941_n_spl_,
    g941_n
  );


  buf

  (
    g941_p_spl_,
    g941_p
  );


  buf

  (
    g834_n_spl_,
    g834_n
  );


  buf

  (
    g943_p_spl_,
    g943_p
  );


  buf

  (
    g834_p_spl_,
    g834_p
  );


  buf

  (
    g943_n_spl_,
    g943_n
  );


  buf

  (
    g944_n_spl_,
    g944_n
  );


  buf

  (
    g944_p_spl_,
    g944_p
  );


  buf

  (
    g833_p_spl_,
    g833_p
  );


  buf

  (
    g946_n_spl_,
    g946_n
  );


  buf

  (
    g947_p_spl_,
    g947_p
  );


  buf

  (
    g977_p_spl_,
    g977_p
  );


  buf

  (
    g977_n_spl_,
    g977_n
  );


  buf

  (
    g978_p_spl_,
    g978_p
  );


  buf

  (
    g979_n_spl_,
    g979_n
  );


  buf

  (
    g978_n_spl_,
    g978_n
  );


  buf

  (
    g979_p_spl_,
    g979_p
  );


  buf

  (
    g980_n_spl_,
    g980_n
  );


  buf

  (
    g980_p_spl_,
    g980_p
  );


  buf

  (
    g976_n_spl_,
    g976_n
  );


  buf

  (
    g982_p_spl_,
    g982_p
  );


  buf

  (
    g976_p_spl_,
    g976_p
  );


  buf

  (
    g982_n_spl_,
    g982_n
  );


  buf

  (
    g983_n_spl_,
    g983_n
  );


  buf

  (
    g983_p_spl_,
    g983_p
  );


  buf

  (
    g975_n_spl_,
    g975_n
  );


  buf

  (
    g985_p_spl_,
    g985_p
  );


  buf

  (
    g975_p_spl_,
    g975_p
  );


  buf

  (
    g985_n_spl_,
    g985_n
  );


  buf

  (
    g986_n_spl_,
    g986_n
  );


  buf

  (
    g986_p_spl_,
    g986_p
  );


  buf

  (
    g974_n_spl_,
    g974_n
  );


  buf

  (
    g988_p_spl_,
    g988_p
  );


  buf

  (
    g974_p_spl_,
    g974_p
  );


  buf

  (
    g988_n_spl_,
    g988_n
  );


  buf

  (
    g989_n_spl_,
    g989_n
  );


  buf

  (
    g989_p_spl_,
    g989_p
  );


  buf

  (
    g973_n_spl_,
    g973_n
  );


  buf

  (
    g991_p_spl_,
    g991_p
  );


  buf

  (
    g973_p_spl_,
    g973_p
  );


  buf

  (
    g991_n_spl_,
    g991_n
  );


  buf

  (
    g992_n_spl_,
    g992_n
  );


  buf

  (
    g992_p_spl_,
    g992_p
  );


  buf

  (
    g972_n_spl_,
    g972_n
  );


  buf

  (
    g994_p_spl_,
    g994_p
  );


  buf

  (
    g972_p_spl_,
    g972_p
  );


  buf

  (
    g994_n_spl_,
    g994_n
  );


  buf

  (
    g995_n_spl_,
    g995_n
  );


  buf

  (
    g995_p_spl_,
    g995_p
  );


  buf

  (
    g971_n_spl_,
    g971_n
  );


  buf

  (
    g997_p_spl_,
    g997_p
  );


  buf

  (
    g971_p_spl_,
    g971_p
  );


  buf

  (
    g997_n_spl_,
    g997_n
  );


  buf

  (
    g998_n_spl_,
    g998_n
  );


  buf

  (
    g998_p_spl_,
    g998_p
  );


  buf

  (
    g970_n_spl_,
    g970_n
  );


  buf

  (
    g1000_p_spl_,
    g1000_p
  );


  buf

  (
    g970_p_spl_,
    g970_p
  );


  buf

  (
    g1000_n_spl_,
    g1000_n
  );


  buf

  (
    g1001_n_spl_,
    g1001_n
  );


  buf

  (
    g1001_p_spl_,
    g1001_p
  );


  buf

  (
    g969_n_spl_,
    g969_n
  );


  buf

  (
    g1003_p_spl_,
    g1003_p
  );


  buf

  (
    g969_p_spl_,
    g969_p
  );


  buf

  (
    g1003_n_spl_,
    g1003_n
  );


  buf

  (
    g1004_n_spl_,
    g1004_n
  );


  buf

  (
    g1004_p_spl_,
    g1004_p
  );


  buf

  (
    g968_n_spl_,
    g968_n
  );


  buf

  (
    g1006_p_spl_,
    g1006_p
  );


  buf

  (
    g968_p_spl_,
    g968_p
  );


  buf

  (
    g1006_n_spl_,
    g1006_n
  );


  buf

  (
    g1007_n_spl_,
    g1007_n
  );


  buf

  (
    g1007_p_spl_,
    g1007_p
  );


  buf

  (
    g967_n_spl_,
    g967_n
  );


  buf

  (
    g1009_p_spl_,
    g1009_p
  );


  buf

  (
    g967_p_spl_,
    g967_p
  );


  buf

  (
    g1009_n_spl_,
    g1009_n
  );


  buf

  (
    g1010_n_spl_,
    g1010_n
  );


  buf

  (
    g1010_p_spl_,
    g1010_p
  );


  buf

  (
    g966_n_spl_,
    g966_n
  );


  buf

  (
    g1012_p_spl_,
    g1012_p
  );


  buf

  (
    g966_p_spl_,
    g966_p
  );


  buf

  (
    g1012_n_spl_,
    g1012_n
  );


  buf

  (
    g1013_n_spl_,
    g1013_n
  );


  buf

  (
    g1013_p_spl_,
    g1013_p
  );


  buf

  (
    g965_n_spl_,
    g965_n
  );


  buf

  (
    g1015_p_spl_,
    g1015_p
  );


  buf

  (
    g965_p_spl_,
    g965_p
  );


  buf

  (
    g1015_n_spl_,
    g1015_n
  );


  buf

  (
    g1016_n_spl_,
    g1016_n
  );


  buf

  (
    g1016_p_spl_,
    g1016_p
  );


  buf

  (
    g964_n_spl_,
    g964_n
  );


  buf

  (
    g1018_p_spl_,
    g1018_p
  );


  buf

  (
    g964_p_spl_,
    g964_p
  );


  buf

  (
    g1018_n_spl_,
    g1018_n
  );


  buf

  (
    g1019_n_spl_,
    g1019_n
  );


  buf

  (
    g1019_p_spl_,
    g1019_p
  );


  buf

  (
    g963_n_spl_,
    g963_n
  );


  buf

  (
    g1021_p_spl_,
    g1021_p
  );


  buf

  (
    g963_p_spl_,
    g963_p
  );


  buf

  (
    g1021_n_spl_,
    g1021_n
  );


  buf

  (
    g1022_n_spl_,
    g1022_n
  );


  buf

  (
    g1022_p_spl_,
    g1022_p
  );


  buf

  (
    g962_n_spl_,
    g962_n
  );


  buf

  (
    g1024_p_spl_,
    g1024_p
  );


  buf

  (
    g962_p_spl_,
    g962_p
  );


  buf

  (
    g1024_n_spl_,
    g1024_n
  );


  buf

  (
    g1025_n_spl_,
    g1025_n
  );


  buf

  (
    g1025_p_spl_,
    g1025_p
  );


  buf

  (
    g961_n_spl_,
    g961_n
  );


  buf

  (
    g1027_p_spl_,
    g1027_p
  );


  buf

  (
    g961_p_spl_,
    g961_p
  );


  buf

  (
    g1027_n_spl_,
    g1027_n
  );


  buf

  (
    g1028_n_spl_,
    g1028_n
  );


  buf

  (
    g1028_p_spl_,
    g1028_p
  );


  buf

  (
    g960_n_spl_,
    g960_n
  );


  buf

  (
    g1030_p_spl_,
    g1030_p
  );


  buf

  (
    g960_p_spl_,
    g960_p
  );


  buf

  (
    g1030_n_spl_,
    g1030_n
  );


  buf

  (
    g1031_n_spl_,
    g1031_n
  );


  buf

  (
    g1031_p_spl_,
    g1031_p
  );


  buf

  (
    g959_n_spl_,
    g959_n
  );


  buf

  (
    g1033_p_spl_,
    g1033_p
  );


  buf

  (
    g959_p_spl_,
    g959_p
  );


  buf

  (
    g1033_n_spl_,
    g1033_n
  );


  buf

  (
    g1034_n_spl_,
    g1034_n
  );


  buf

  (
    g1034_p_spl_,
    g1034_p
  );


  buf

  (
    g958_n_spl_,
    g958_n
  );


  buf

  (
    g1036_p_spl_,
    g1036_p
  );


  buf

  (
    g958_p_spl_,
    g958_p
  );


  buf

  (
    g1036_n_spl_,
    g1036_n
  );


  buf

  (
    g1037_n_spl_,
    g1037_n
  );


  buf

  (
    g1037_p_spl_,
    g1037_p
  );


  buf

  (
    g957_n_spl_,
    g957_n
  );


  buf

  (
    g1039_p_spl_,
    g1039_p
  );


  buf

  (
    g957_p_spl_,
    g957_p
  );


  buf

  (
    g1039_n_spl_,
    g1039_n
  );


  buf

  (
    g1040_n_spl_,
    g1040_n
  );


  buf

  (
    g1040_p_spl_,
    g1040_p
  );


  buf

  (
    g956_n_spl_,
    g956_n
  );


  buf

  (
    g1042_p_spl_,
    g1042_p
  );


  buf

  (
    g956_p_spl_,
    g956_p
  );


  buf

  (
    g1042_n_spl_,
    g1042_n
  );


  buf

  (
    g1043_n_spl_,
    g1043_n
  );


  buf

  (
    g1043_p_spl_,
    g1043_p
  );


  buf

  (
    g955_n_spl_,
    g955_n
  );


  buf

  (
    g1045_p_spl_,
    g1045_p
  );


  buf

  (
    g955_p_spl_,
    g955_p
  );


  buf

  (
    g1045_n_spl_,
    g1045_n
  );


  buf

  (
    g1046_n_spl_,
    g1046_n
  );


  buf

  (
    g1046_p_spl_,
    g1046_p
  );


  buf

  (
    g954_n_spl_,
    g954_n
  );


  buf

  (
    g1048_p_spl_,
    g1048_p
  );


  buf

  (
    g954_p_spl_,
    g954_p
  );


  buf

  (
    g1048_n_spl_,
    g1048_n
  );


  buf

  (
    g1049_n_spl_,
    g1049_n
  );


  buf

  (
    g1049_p_spl_,
    g1049_p
  );


  buf

  (
    g953_n_spl_,
    g953_n
  );


  buf

  (
    g1051_p_spl_,
    g1051_p
  );


  buf

  (
    g953_p_spl_,
    g953_p
  );


  buf

  (
    g1051_n_spl_,
    g1051_n
  );


  buf

  (
    g1052_n_spl_,
    g1052_n
  );


  buf

  (
    g1052_p_spl_,
    g1052_p
  );


  buf

  (
    g952_n_spl_,
    g952_n
  );


  buf

  (
    g1054_p_spl_,
    g1054_p
  );


  buf

  (
    g952_p_spl_,
    g952_p
  );


  buf

  (
    g1054_n_spl_,
    g1054_n
  );


  buf

  (
    g1055_n_spl_,
    g1055_n
  );


  buf

  (
    g1055_p_spl_,
    g1055_p
  );


  buf

  (
    g951_n_spl_,
    g951_n
  );


  buf

  (
    g1057_p_spl_,
    g1057_p
  );


  buf

  (
    g951_p_spl_,
    g951_p
  );


  buf

  (
    g1057_n_spl_,
    g1057_n
  );


  buf

  (
    g1058_n_spl_,
    g1058_n
  );


  buf

  (
    g1058_p_spl_,
    g1058_p
  );


  buf

  (
    g950_p_spl_,
    g950_p
  );


  buf

  (
    g1060_n_spl_,
    g1060_n
  );


  buf

  (
    g1062_n_spl_,
    g1062_n
  );


  buf

  (
    g1090_n_spl_,
    g1090_n
  );


  buf

  (
    g1091_n_spl_,
    g1091_n
  );


  buf

  (
    g1090_p_spl_,
    g1090_p
  );


  buf

  (
    g1091_p_spl_,
    g1091_p
  );


  buf

  (
    g1092_n_spl_,
    g1092_n
  );


  buf

  (
    g1092_p_spl_,
    g1092_p
  );


  buf

  (
    g1089_n_spl_,
    g1089_n
  );


  buf

  (
    g1094_p_spl_,
    g1094_p
  );


  buf

  (
    g1089_p_spl_,
    g1089_p
  );


  buf

  (
    g1094_n_spl_,
    g1094_n
  );


  buf

  (
    g1095_n_spl_,
    g1095_n
  );


  buf

  (
    g1095_p_spl_,
    g1095_p
  );


  buf

  (
    g1088_n_spl_,
    g1088_n
  );


  buf

  (
    g1097_p_spl_,
    g1097_p
  );


  buf

  (
    g1088_p_spl_,
    g1088_p
  );


  buf

  (
    g1097_n_spl_,
    g1097_n
  );


  buf

  (
    g1098_n_spl_,
    g1098_n
  );


  buf

  (
    g1098_p_spl_,
    g1098_p
  );


  buf

  (
    g1087_n_spl_,
    g1087_n
  );


  buf

  (
    g1100_p_spl_,
    g1100_p
  );


  buf

  (
    g1087_p_spl_,
    g1087_p
  );


  buf

  (
    g1100_n_spl_,
    g1100_n
  );


  buf

  (
    g1101_n_spl_,
    g1101_n
  );


  buf

  (
    g1101_p_spl_,
    g1101_p
  );


  buf

  (
    g1086_n_spl_,
    g1086_n
  );


  buf

  (
    g1103_p_spl_,
    g1103_p
  );


  buf

  (
    g1086_p_spl_,
    g1086_p
  );


  buf

  (
    g1103_n_spl_,
    g1103_n
  );


  buf

  (
    g1104_n_spl_,
    g1104_n
  );


  buf

  (
    g1104_p_spl_,
    g1104_p
  );


  buf

  (
    g1085_n_spl_,
    g1085_n
  );


  buf

  (
    g1106_p_spl_,
    g1106_p
  );


  buf

  (
    g1085_p_spl_,
    g1085_p
  );


  buf

  (
    g1106_n_spl_,
    g1106_n
  );


  buf

  (
    g1107_n_spl_,
    g1107_n
  );


  buf

  (
    g1107_p_spl_,
    g1107_p
  );


  buf

  (
    g1084_n_spl_,
    g1084_n
  );


  buf

  (
    g1109_p_spl_,
    g1109_p
  );


  buf

  (
    g1084_p_spl_,
    g1084_p
  );


  buf

  (
    g1109_n_spl_,
    g1109_n
  );


  buf

  (
    g1110_n_spl_,
    g1110_n
  );


  buf

  (
    g1110_p_spl_,
    g1110_p
  );


  buf

  (
    g1083_n_spl_,
    g1083_n
  );


  buf

  (
    g1112_p_spl_,
    g1112_p
  );


  buf

  (
    g1083_p_spl_,
    g1083_p
  );


  buf

  (
    g1112_n_spl_,
    g1112_n
  );


  buf

  (
    g1113_n_spl_,
    g1113_n
  );


  buf

  (
    g1113_p_spl_,
    g1113_p
  );


  buf

  (
    g1082_n_spl_,
    g1082_n
  );


  buf

  (
    g1115_p_spl_,
    g1115_p
  );


  buf

  (
    g1082_p_spl_,
    g1082_p
  );


  buf

  (
    g1115_n_spl_,
    g1115_n
  );


  buf

  (
    g1116_n_spl_,
    g1116_n
  );


  buf

  (
    g1116_p_spl_,
    g1116_p
  );


  buf

  (
    g1081_n_spl_,
    g1081_n
  );


  buf

  (
    g1118_p_spl_,
    g1118_p
  );


  buf

  (
    g1081_p_spl_,
    g1081_p
  );


  buf

  (
    g1118_n_spl_,
    g1118_n
  );


  buf

  (
    g1119_n_spl_,
    g1119_n
  );


  buf

  (
    g1119_p_spl_,
    g1119_p
  );


  buf

  (
    g1080_n_spl_,
    g1080_n
  );


  buf

  (
    g1121_p_spl_,
    g1121_p
  );


  buf

  (
    g1080_p_spl_,
    g1080_p
  );


  buf

  (
    g1121_n_spl_,
    g1121_n
  );


  buf

  (
    g1122_n_spl_,
    g1122_n
  );


  buf

  (
    g1122_p_spl_,
    g1122_p
  );


  buf

  (
    g1079_n_spl_,
    g1079_n
  );


  buf

  (
    g1124_p_spl_,
    g1124_p
  );


  buf

  (
    g1079_p_spl_,
    g1079_p
  );


  buf

  (
    g1124_n_spl_,
    g1124_n
  );


  buf

  (
    g1125_n_spl_,
    g1125_n
  );


  buf

  (
    g1125_p_spl_,
    g1125_p
  );


  buf

  (
    g1078_n_spl_,
    g1078_n
  );


  buf

  (
    g1127_p_spl_,
    g1127_p
  );


  buf

  (
    g1078_p_spl_,
    g1078_p
  );


  buf

  (
    g1127_n_spl_,
    g1127_n
  );


  buf

  (
    g1128_n_spl_,
    g1128_n
  );


  buf

  (
    g1128_p_spl_,
    g1128_p
  );


  buf

  (
    g1077_n_spl_,
    g1077_n
  );


  buf

  (
    g1130_p_spl_,
    g1130_p
  );


  buf

  (
    g1077_p_spl_,
    g1077_p
  );


  buf

  (
    g1130_n_spl_,
    g1130_n
  );


  buf

  (
    g1131_n_spl_,
    g1131_n
  );


  buf

  (
    g1131_p_spl_,
    g1131_p
  );


  buf

  (
    g1076_n_spl_,
    g1076_n
  );


  buf

  (
    g1133_p_spl_,
    g1133_p
  );


  buf

  (
    g1076_p_spl_,
    g1076_p
  );


  buf

  (
    g1133_n_spl_,
    g1133_n
  );


  buf

  (
    g1134_n_spl_,
    g1134_n
  );


  buf

  (
    g1134_p_spl_,
    g1134_p
  );


  buf

  (
    g1075_n_spl_,
    g1075_n
  );


  buf

  (
    g1136_p_spl_,
    g1136_p
  );


  buf

  (
    g1075_p_spl_,
    g1075_p
  );


  buf

  (
    g1136_n_spl_,
    g1136_n
  );


  buf

  (
    g1137_n_spl_,
    g1137_n
  );


  buf

  (
    g1137_p_spl_,
    g1137_p
  );


  buf

  (
    g1074_n_spl_,
    g1074_n
  );


  buf

  (
    g1139_p_spl_,
    g1139_p
  );


  buf

  (
    g1074_p_spl_,
    g1074_p
  );


  buf

  (
    g1139_n_spl_,
    g1139_n
  );


  buf

  (
    g1140_n_spl_,
    g1140_n
  );


  buf

  (
    g1140_p_spl_,
    g1140_p
  );


  buf

  (
    g1073_n_spl_,
    g1073_n
  );


  buf

  (
    g1142_p_spl_,
    g1142_p
  );


  buf

  (
    g1073_p_spl_,
    g1073_p
  );


  buf

  (
    g1142_n_spl_,
    g1142_n
  );


  buf

  (
    g1143_n_spl_,
    g1143_n
  );


  buf

  (
    g1143_p_spl_,
    g1143_p
  );


  buf

  (
    g1072_n_spl_,
    g1072_n
  );


  buf

  (
    g1145_p_spl_,
    g1145_p
  );


  buf

  (
    g1072_p_spl_,
    g1072_p
  );


  buf

  (
    g1145_n_spl_,
    g1145_n
  );


  buf

  (
    g1146_n_spl_,
    g1146_n
  );


  buf

  (
    g1146_p_spl_,
    g1146_p
  );


  buf

  (
    g1071_n_spl_,
    g1071_n
  );


  buf

  (
    g1148_p_spl_,
    g1148_p
  );


  buf

  (
    g1071_p_spl_,
    g1071_p
  );


  buf

  (
    g1148_n_spl_,
    g1148_n
  );


  buf

  (
    g1149_n_spl_,
    g1149_n
  );


  buf

  (
    g1149_p_spl_,
    g1149_p
  );


  buf

  (
    g1070_n_spl_,
    g1070_n
  );


  buf

  (
    g1151_p_spl_,
    g1151_p
  );


  buf

  (
    g1070_p_spl_,
    g1070_p
  );


  buf

  (
    g1151_n_spl_,
    g1151_n
  );


  buf

  (
    g1152_n_spl_,
    g1152_n
  );


  buf

  (
    g1152_p_spl_,
    g1152_p
  );


  buf

  (
    g1069_n_spl_,
    g1069_n
  );


  buf

  (
    g1154_p_spl_,
    g1154_p
  );


  buf

  (
    g1069_p_spl_,
    g1069_p
  );


  buf

  (
    g1154_n_spl_,
    g1154_n
  );


  buf

  (
    g1155_n_spl_,
    g1155_n
  );


  buf

  (
    g1155_p_spl_,
    g1155_p
  );


  buf

  (
    g1068_n_spl_,
    g1068_n
  );


  buf

  (
    g1157_p_spl_,
    g1157_p
  );


  buf

  (
    g1068_p_spl_,
    g1068_p
  );


  buf

  (
    g1157_n_spl_,
    g1157_n
  );


  buf

  (
    g1158_n_spl_,
    g1158_n
  );


  buf

  (
    g1158_p_spl_,
    g1158_p
  );


  buf

  (
    g1067_n_spl_,
    g1067_n
  );


  buf

  (
    g1160_p_spl_,
    g1160_p
  );


  buf

  (
    g1067_p_spl_,
    g1067_p
  );


  buf

  (
    g1160_n_spl_,
    g1160_n
  );


  buf

  (
    g1161_n_spl_,
    g1161_n
  );


  buf

  (
    g1161_p_spl_,
    g1161_p
  );


  buf

  (
    g1066_n_spl_,
    g1066_n
  );


  buf

  (
    g1163_p_spl_,
    g1163_p
  );


  buf

  (
    g1066_p_spl_,
    g1066_p
  );


  buf

  (
    g1163_n_spl_,
    g1163_n
  );


  buf

  (
    g1164_n_spl_,
    g1164_n
  );


  buf

  (
    g1164_p_spl_,
    g1164_p
  );


  buf

  (
    g1065_n_spl_,
    g1065_n
  );


  buf

  (
    g1166_p_spl_,
    g1166_p
  );


  buf

  (
    g1065_p_spl_,
    g1065_p
  );


  buf

  (
    g1166_n_spl_,
    g1166_n
  );


  buf

  (
    g1167_n_spl_,
    g1167_n
  );


  buf

  (
    g1167_p_spl_,
    g1167_p
  );


  buf

  (
    g1064_n_spl_,
    g1064_n
  );


  buf

  (
    g1169_p_spl_,
    g1169_p
  );


  buf

  (
    g1064_p_spl_,
    g1064_p
  );


  buf

  (
    g1169_n_spl_,
    g1169_n
  );


  buf

  (
    g1170_n_spl_,
    g1170_n
  );


  buf

  (
    g1170_p_spl_,
    g1170_p
  );


  buf

  (
    g1062_p_spl_,
    g1062_p
  );


  buf

  (
    g1172_n_spl_,
    g1172_n
  );


  buf

  (
    g1173_p_spl_,
    g1173_p
  );


  buf

  (
    g1201_n_spl_,
    g1201_n
  );


  buf

  (
    g1202_n_spl_,
    g1202_n
  );


  buf

  (
    g1201_p_spl_,
    g1201_p
  );


  buf

  (
    g1202_p_spl_,
    g1202_p
  );


  buf

  (
    g1203_n_spl_,
    g1203_n
  );


  buf

  (
    g1203_p_spl_,
    g1203_p
  );


  buf

  (
    g1200_n_spl_,
    g1200_n
  );


  buf

  (
    g1205_p_spl_,
    g1205_p
  );


  buf

  (
    g1200_p_spl_,
    g1200_p
  );


  buf

  (
    g1205_n_spl_,
    g1205_n
  );


  buf

  (
    g1206_n_spl_,
    g1206_n
  );


  buf

  (
    g1206_p_spl_,
    g1206_p
  );


  buf

  (
    g1199_n_spl_,
    g1199_n
  );


  buf

  (
    g1208_p_spl_,
    g1208_p
  );


  buf

  (
    g1199_p_spl_,
    g1199_p
  );


  buf

  (
    g1208_n_spl_,
    g1208_n
  );


  buf

  (
    g1209_n_spl_,
    g1209_n
  );


  buf

  (
    g1209_p_spl_,
    g1209_p
  );


  buf

  (
    g1198_n_spl_,
    g1198_n
  );


  buf

  (
    g1211_p_spl_,
    g1211_p
  );


  buf

  (
    g1198_p_spl_,
    g1198_p
  );


  buf

  (
    g1211_n_spl_,
    g1211_n
  );


  buf

  (
    g1212_n_spl_,
    g1212_n
  );


  buf

  (
    g1212_p_spl_,
    g1212_p
  );


  buf

  (
    g1197_n_spl_,
    g1197_n
  );


  buf

  (
    g1214_p_spl_,
    g1214_p
  );


  buf

  (
    g1197_p_spl_,
    g1197_p
  );


  buf

  (
    g1214_n_spl_,
    g1214_n
  );


  buf

  (
    g1215_n_spl_,
    g1215_n
  );


  buf

  (
    g1215_p_spl_,
    g1215_p
  );


  buf

  (
    g1196_n_spl_,
    g1196_n
  );


  buf

  (
    g1217_p_spl_,
    g1217_p
  );


  buf

  (
    g1196_p_spl_,
    g1196_p
  );


  buf

  (
    g1217_n_spl_,
    g1217_n
  );


  buf

  (
    g1218_n_spl_,
    g1218_n
  );


  buf

  (
    g1218_p_spl_,
    g1218_p
  );


  buf

  (
    g1195_n_spl_,
    g1195_n
  );


  buf

  (
    g1220_p_spl_,
    g1220_p
  );


  buf

  (
    g1195_p_spl_,
    g1195_p
  );


  buf

  (
    g1220_n_spl_,
    g1220_n
  );


  buf

  (
    g1221_n_spl_,
    g1221_n
  );


  buf

  (
    g1221_p_spl_,
    g1221_p
  );


  buf

  (
    g1194_n_spl_,
    g1194_n
  );


  buf

  (
    g1223_p_spl_,
    g1223_p
  );


  buf

  (
    g1194_p_spl_,
    g1194_p
  );


  buf

  (
    g1223_n_spl_,
    g1223_n
  );


  buf

  (
    g1224_n_spl_,
    g1224_n
  );


  buf

  (
    g1224_p_spl_,
    g1224_p
  );


  buf

  (
    g1193_n_spl_,
    g1193_n
  );


  buf

  (
    g1226_p_spl_,
    g1226_p
  );


  buf

  (
    g1193_p_spl_,
    g1193_p
  );


  buf

  (
    g1226_n_spl_,
    g1226_n
  );


  buf

  (
    g1227_n_spl_,
    g1227_n
  );


  buf

  (
    g1227_p_spl_,
    g1227_p
  );


  buf

  (
    g1192_n_spl_,
    g1192_n
  );


  buf

  (
    g1229_p_spl_,
    g1229_p
  );


  buf

  (
    g1192_p_spl_,
    g1192_p
  );


  buf

  (
    g1229_n_spl_,
    g1229_n
  );


  buf

  (
    g1230_n_spl_,
    g1230_n
  );


  buf

  (
    g1230_p_spl_,
    g1230_p
  );


  buf

  (
    g1191_n_spl_,
    g1191_n
  );


  buf

  (
    g1232_p_spl_,
    g1232_p
  );


  buf

  (
    g1191_p_spl_,
    g1191_p
  );


  buf

  (
    g1232_n_spl_,
    g1232_n
  );


  buf

  (
    g1233_n_spl_,
    g1233_n
  );


  buf

  (
    g1233_p_spl_,
    g1233_p
  );


  buf

  (
    g1190_n_spl_,
    g1190_n
  );


  buf

  (
    g1235_p_spl_,
    g1235_p
  );


  buf

  (
    g1190_p_spl_,
    g1190_p
  );


  buf

  (
    g1235_n_spl_,
    g1235_n
  );


  buf

  (
    g1236_n_spl_,
    g1236_n
  );


  buf

  (
    g1236_p_spl_,
    g1236_p
  );


  buf

  (
    g1189_n_spl_,
    g1189_n
  );


  buf

  (
    g1238_p_spl_,
    g1238_p
  );


  buf

  (
    g1189_p_spl_,
    g1189_p
  );


  buf

  (
    g1238_n_spl_,
    g1238_n
  );


  buf

  (
    g1239_n_spl_,
    g1239_n
  );


  buf

  (
    g1239_p_spl_,
    g1239_p
  );


  buf

  (
    g1188_n_spl_,
    g1188_n
  );


  buf

  (
    g1241_p_spl_,
    g1241_p
  );


  buf

  (
    g1188_p_spl_,
    g1188_p
  );


  buf

  (
    g1241_n_spl_,
    g1241_n
  );


  buf

  (
    g1242_n_spl_,
    g1242_n
  );


  buf

  (
    g1242_p_spl_,
    g1242_p
  );


  buf

  (
    g1187_n_spl_,
    g1187_n
  );


  buf

  (
    g1244_p_spl_,
    g1244_p
  );


  buf

  (
    g1187_p_spl_,
    g1187_p
  );


  buf

  (
    g1244_n_spl_,
    g1244_n
  );


  buf

  (
    g1245_n_spl_,
    g1245_n
  );


  buf

  (
    g1245_p_spl_,
    g1245_p
  );


  buf

  (
    g1186_n_spl_,
    g1186_n
  );


  buf

  (
    g1247_p_spl_,
    g1247_p
  );


  buf

  (
    g1186_p_spl_,
    g1186_p
  );


  buf

  (
    g1247_n_spl_,
    g1247_n
  );


  buf

  (
    g1248_n_spl_,
    g1248_n
  );


  buf

  (
    g1248_p_spl_,
    g1248_p
  );


  buf

  (
    g1185_n_spl_,
    g1185_n
  );


  buf

  (
    g1250_p_spl_,
    g1250_p
  );


  buf

  (
    g1185_p_spl_,
    g1185_p
  );


  buf

  (
    g1250_n_spl_,
    g1250_n
  );


  buf

  (
    g1251_n_spl_,
    g1251_n
  );


  buf

  (
    g1251_p_spl_,
    g1251_p
  );


  buf

  (
    g1184_n_spl_,
    g1184_n
  );


  buf

  (
    g1253_p_spl_,
    g1253_p
  );


  buf

  (
    g1184_p_spl_,
    g1184_p
  );


  buf

  (
    g1253_n_spl_,
    g1253_n
  );


  buf

  (
    g1254_n_spl_,
    g1254_n
  );


  buf

  (
    g1254_p_spl_,
    g1254_p
  );


  buf

  (
    g1183_n_spl_,
    g1183_n
  );


  buf

  (
    g1256_p_spl_,
    g1256_p
  );


  buf

  (
    g1183_p_spl_,
    g1183_p
  );


  buf

  (
    g1256_n_spl_,
    g1256_n
  );


  buf

  (
    g1257_n_spl_,
    g1257_n
  );


  buf

  (
    g1257_p_spl_,
    g1257_p
  );


  buf

  (
    g1182_n_spl_,
    g1182_n
  );


  buf

  (
    g1259_p_spl_,
    g1259_p
  );


  buf

  (
    g1182_p_spl_,
    g1182_p
  );


  buf

  (
    g1259_n_spl_,
    g1259_n
  );


  buf

  (
    g1260_n_spl_,
    g1260_n
  );


  buf

  (
    g1260_p_spl_,
    g1260_p
  );


  buf

  (
    g1181_n_spl_,
    g1181_n
  );


  buf

  (
    g1262_p_spl_,
    g1262_p
  );


  buf

  (
    g1181_p_spl_,
    g1181_p
  );


  buf

  (
    g1262_n_spl_,
    g1262_n
  );


  buf

  (
    g1263_n_spl_,
    g1263_n
  );


  buf

  (
    g1263_p_spl_,
    g1263_p
  );


  buf

  (
    g1180_n_spl_,
    g1180_n
  );


  buf

  (
    g1265_p_spl_,
    g1265_p
  );


  buf

  (
    g1180_p_spl_,
    g1180_p
  );


  buf

  (
    g1265_n_spl_,
    g1265_n
  );


  buf

  (
    g1266_n_spl_,
    g1266_n
  );


  buf

  (
    g1266_p_spl_,
    g1266_p
  );


  buf

  (
    g1179_n_spl_,
    g1179_n
  );


  buf

  (
    g1268_p_spl_,
    g1268_p
  );


  buf

  (
    g1179_p_spl_,
    g1179_p
  );


  buf

  (
    g1268_n_spl_,
    g1268_n
  );


  buf

  (
    g1269_n_spl_,
    g1269_n
  );


  buf

  (
    g1269_p_spl_,
    g1269_p
  );


  buf

  (
    g1178_n_spl_,
    g1178_n
  );


  buf

  (
    g1271_p_spl_,
    g1271_p
  );


  buf

  (
    g1178_p_spl_,
    g1178_p
  );


  buf

  (
    g1271_n_spl_,
    g1271_n
  );


  buf

  (
    g1272_n_spl_,
    g1272_n
  );


  buf

  (
    g1272_p_spl_,
    g1272_p
  );


  buf

  (
    g1177_n_spl_,
    g1177_n
  );


  buf

  (
    g1274_p_spl_,
    g1274_p
  );


  buf

  (
    g1177_p_spl_,
    g1177_p
  );


  buf

  (
    g1274_n_spl_,
    g1274_n
  );


  buf

  (
    g1275_n_spl_,
    g1275_n
  );


  buf

  (
    g1275_p_spl_,
    g1275_p
  );


  buf

  (
    g1176_p_spl_,
    g1176_p
  );


  buf

  (
    g1277_n_spl_,
    g1277_n
  );


  buf

  (
    g1278_p_spl_,
    g1278_p
  );


  buf

  (
    g1304_n_spl_,
    g1304_n
  );


  buf

  (
    g1305_n_spl_,
    g1305_n
  );


  buf

  (
    g1304_p_spl_,
    g1304_p
  );


  buf

  (
    g1305_p_spl_,
    g1305_p
  );


  buf

  (
    g1306_n_spl_,
    g1306_n
  );


  buf

  (
    g1306_p_spl_,
    g1306_p
  );


  buf

  (
    g1303_n_spl_,
    g1303_n
  );


  buf

  (
    g1308_p_spl_,
    g1308_p
  );


  buf

  (
    g1303_p_spl_,
    g1303_p
  );


  buf

  (
    g1308_n_spl_,
    g1308_n
  );


  buf

  (
    g1309_n_spl_,
    g1309_n
  );


  buf

  (
    g1309_p_spl_,
    g1309_p
  );


  buf

  (
    g1302_n_spl_,
    g1302_n
  );


  buf

  (
    g1311_p_spl_,
    g1311_p
  );


  buf

  (
    g1302_p_spl_,
    g1302_p
  );


  buf

  (
    g1311_n_spl_,
    g1311_n
  );


  buf

  (
    g1312_n_spl_,
    g1312_n
  );


  buf

  (
    g1312_p_spl_,
    g1312_p
  );


  buf

  (
    g1301_n_spl_,
    g1301_n
  );


  buf

  (
    g1314_p_spl_,
    g1314_p
  );


  buf

  (
    g1301_p_spl_,
    g1301_p
  );


  buf

  (
    g1314_n_spl_,
    g1314_n
  );


  buf

  (
    g1315_n_spl_,
    g1315_n
  );


  buf

  (
    g1315_p_spl_,
    g1315_p
  );


  buf

  (
    g1300_n_spl_,
    g1300_n
  );


  buf

  (
    g1317_p_spl_,
    g1317_p
  );


  buf

  (
    g1300_p_spl_,
    g1300_p
  );


  buf

  (
    g1317_n_spl_,
    g1317_n
  );


  buf

  (
    g1318_n_spl_,
    g1318_n
  );


  buf

  (
    g1318_p_spl_,
    g1318_p
  );


  buf

  (
    g1299_n_spl_,
    g1299_n
  );


  buf

  (
    g1320_p_spl_,
    g1320_p
  );


  buf

  (
    g1299_p_spl_,
    g1299_p
  );


  buf

  (
    g1320_n_spl_,
    g1320_n
  );


  buf

  (
    g1321_n_spl_,
    g1321_n
  );


  buf

  (
    g1321_p_spl_,
    g1321_p
  );


  buf

  (
    g1298_n_spl_,
    g1298_n
  );


  buf

  (
    g1323_p_spl_,
    g1323_p
  );


  buf

  (
    g1298_p_spl_,
    g1298_p
  );


  buf

  (
    g1323_n_spl_,
    g1323_n
  );


  buf

  (
    g1324_n_spl_,
    g1324_n
  );


  buf

  (
    g1324_p_spl_,
    g1324_p
  );


  buf

  (
    g1297_n_spl_,
    g1297_n
  );


  buf

  (
    g1326_p_spl_,
    g1326_p
  );


  buf

  (
    g1297_p_spl_,
    g1297_p
  );


  buf

  (
    g1326_n_spl_,
    g1326_n
  );


  buf

  (
    g1327_n_spl_,
    g1327_n
  );


  buf

  (
    g1327_p_spl_,
    g1327_p
  );


  buf

  (
    g1296_n_spl_,
    g1296_n
  );


  buf

  (
    g1329_p_spl_,
    g1329_p
  );


  buf

  (
    g1296_p_spl_,
    g1296_p
  );


  buf

  (
    g1329_n_spl_,
    g1329_n
  );


  buf

  (
    g1330_n_spl_,
    g1330_n
  );


  buf

  (
    g1330_p_spl_,
    g1330_p
  );


  buf

  (
    g1295_n_spl_,
    g1295_n
  );


  buf

  (
    g1332_p_spl_,
    g1332_p
  );


  buf

  (
    g1295_p_spl_,
    g1295_p
  );


  buf

  (
    g1332_n_spl_,
    g1332_n
  );


  buf

  (
    g1333_n_spl_,
    g1333_n
  );


  buf

  (
    g1333_p_spl_,
    g1333_p
  );


  buf

  (
    g1294_n_spl_,
    g1294_n
  );


  buf

  (
    g1335_p_spl_,
    g1335_p
  );


  buf

  (
    g1294_p_spl_,
    g1294_p
  );


  buf

  (
    g1335_n_spl_,
    g1335_n
  );


  buf

  (
    g1336_n_spl_,
    g1336_n
  );


  buf

  (
    g1336_p_spl_,
    g1336_p
  );


  buf

  (
    g1293_n_spl_,
    g1293_n
  );


  buf

  (
    g1338_p_spl_,
    g1338_p
  );


  buf

  (
    g1293_p_spl_,
    g1293_p
  );


  buf

  (
    g1338_n_spl_,
    g1338_n
  );


  buf

  (
    g1339_n_spl_,
    g1339_n
  );


  buf

  (
    g1339_p_spl_,
    g1339_p
  );


  buf

  (
    g1292_n_spl_,
    g1292_n
  );


  buf

  (
    g1341_p_spl_,
    g1341_p
  );


  buf

  (
    g1292_p_spl_,
    g1292_p
  );


  buf

  (
    g1341_n_spl_,
    g1341_n
  );


  buf

  (
    g1342_n_spl_,
    g1342_n
  );


  buf

  (
    g1342_p_spl_,
    g1342_p
  );


  buf

  (
    g1291_n_spl_,
    g1291_n
  );


  buf

  (
    g1344_p_spl_,
    g1344_p
  );


  buf

  (
    g1291_p_spl_,
    g1291_p
  );


  buf

  (
    g1344_n_spl_,
    g1344_n
  );


  buf

  (
    g1345_n_spl_,
    g1345_n
  );


  buf

  (
    g1345_p_spl_,
    g1345_p
  );


  buf

  (
    g1290_n_spl_,
    g1290_n
  );


  buf

  (
    g1347_p_spl_,
    g1347_p
  );


  buf

  (
    g1290_p_spl_,
    g1290_p
  );


  buf

  (
    g1347_n_spl_,
    g1347_n
  );


  buf

  (
    g1348_n_spl_,
    g1348_n
  );


  buf

  (
    g1348_p_spl_,
    g1348_p
  );


  buf

  (
    g1289_n_spl_,
    g1289_n
  );


  buf

  (
    g1350_p_spl_,
    g1350_p
  );


  buf

  (
    g1289_p_spl_,
    g1289_p
  );


  buf

  (
    g1350_n_spl_,
    g1350_n
  );


  buf

  (
    g1351_n_spl_,
    g1351_n
  );


  buf

  (
    g1351_p_spl_,
    g1351_p
  );


  buf

  (
    g1288_n_spl_,
    g1288_n
  );


  buf

  (
    g1353_p_spl_,
    g1353_p
  );


  buf

  (
    g1288_p_spl_,
    g1288_p
  );


  buf

  (
    g1353_n_spl_,
    g1353_n
  );


  buf

  (
    g1354_n_spl_,
    g1354_n
  );


  buf

  (
    g1354_p_spl_,
    g1354_p
  );


  buf

  (
    g1287_n_spl_,
    g1287_n
  );


  buf

  (
    g1356_p_spl_,
    g1356_p
  );


  buf

  (
    g1287_p_spl_,
    g1287_p
  );


  buf

  (
    g1356_n_spl_,
    g1356_n
  );


  buf

  (
    g1357_n_spl_,
    g1357_n
  );


  buf

  (
    g1357_p_spl_,
    g1357_p
  );


  buf

  (
    g1286_n_spl_,
    g1286_n
  );


  buf

  (
    g1359_p_spl_,
    g1359_p
  );


  buf

  (
    g1286_p_spl_,
    g1286_p
  );


  buf

  (
    g1359_n_spl_,
    g1359_n
  );


  buf

  (
    g1360_n_spl_,
    g1360_n
  );


  buf

  (
    g1360_p_spl_,
    g1360_p
  );


  buf

  (
    g1285_n_spl_,
    g1285_n
  );


  buf

  (
    g1362_p_spl_,
    g1362_p
  );


  buf

  (
    g1285_p_spl_,
    g1285_p
  );


  buf

  (
    g1362_n_spl_,
    g1362_n
  );


  buf

  (
    g1363_n_spl_,
    g1363_n
  );


  buf

  (
    g1363_p_spl_,
    g1363_p
  );


  buf

  (
    g1284_n_spl_,
    g1284_n
  );


  buf

  (
    g1365_p_spl_,
    g1365_p
  );


  buf

  (
    g1284_p_spl_,
    g1284_p
  );


  buf

  (
    g1365_n_spl_,
    g1365_n
  );


  buf

  (
    g1366_n_spl_,
    g1366_n
  );


  buf

  (
    g1366_p_spl_,
    g1366_p
  );


  buf

  (
    g1283_n_spl_,
    g1283_n
  );


  buf

  (
    g1368_p_spl_,
    g1368_p
  );


  buf

  (
    g1283_p_spl_,
    g1283_p
  );


  buf

  (
    g1368_n_spl_,
    g1368_n
  );


  buf

  (
    g1369_n_spl_,
    g1369_n
  );


  buf

  (
    g1369_p_spl_,
    g1369_p
  );


  buf

  (
    g1282_n_spl_,
    g1282_n
  );


  buf

  (
    g1371_p_spl_,
    g1371_p
  );


  buf

  (
    g1282_p_spl_,
    g1282_p
  );


  buf

  (
    g1371_n_spl_,
    g1371_n
  );


  buf

  (
    g1372_n_spl_,
    g1372_n
  );


  buf

  (
    g1372_p_spl_,
    g1372_p
  );


  buf

  (
    g1281_p_spl_,
    g1281_p
  );


  buf

  (
    g1374_n_spl_,
    g1374_n
  );


  buf

  (
    g1375_p_spl_,
    g1375_p
  );


  buf

  (
    g1399_n_spl_,
    g1399_n
  );


  buf

  (
    g1400_n_spl_,
    g1400_n
  );


  buf

  (
    g1399_p_spl_,
    g1399_p
  );


  buf

  (
    g1400_p_spl_,
    g1400_p
  );


  buf

  (
    g1401_n_spl_,
    g1401_n
  );


  buf

  (
    g1401_p_spl_,
    g1401_p
  );


  buf

  (
    g1398_n_spl_,
    g1398_n
  );


  buf

  (
    g1403_p_spl_,
    g1403_p
  );


  buf

  (
    g1398_p_spl_,
    g1398_p
  );


  buf

  (
    g1403_n_spl_,
    g1403_n
  );


  buf

  (
    g1404_n_spl_,
    g1404_n
  );


  buf

  (
    g1404_p_spl_,
    g1404_p
  );


  buf

  (
    g1397_n_spl_,
    g1397_n
  );


  buf

  (
    g1406_p_spl_,
    g1406_p
  );


  buf

  (
    g1397_p_spl_,
    g1397_p
  );


  buf

  (
    g1406_n_spl_,
    g1406_n
  );


  buf

  (
    g1407_n_spl_,
    g1407_n
  );


  buf

  (
    g1407_p_spl_,
    g1407_p
  );


  buf

  (
    g1396_n_spl_,
    g1396_n
  );


  buf

  (
    g1409_p_spl_,
    g1409_p
  );


  buf

  (
    g1396_p_spl_,
    g1396_p
  );


  buf

  (
    g1409_n_spl_,
    g1409_n
  );


  buf

  (
    g1410_n_spl_,
    g1410_n
  );


  buf

  (
    g1410_p_spl_,
    g1410_p
  );


  buf

  (
    g1395_n_spl_,
    g1395_n
  );


  buf

  (
    g1412_p_spl_,
    g1412_p
  );


  buf

  (
    g1395_p_spl_,
    g1395_p
  );


  buf

  (
    g1412_n_spl_,
    g1412_n
  );


  buf

  (
    g1413_n_spl_,
    g1413_n
  );


  buf

  (
    g1413_p_spl_,
    g1413_p
  );


  buf

  (
    g1394_n_spl_,
    g1394_n
  );


  buf

  (
    g1415_p_spl_,
    g1415_p
  );


  buf

  (
    g1394_p_spl_,
    g1394_p
  );


  buf

  (
    g1415_n_spl_,
    g1415_n
  );


  buf

  (
    g1416_n_spl_,
    g1416_n
  );


  buf

  (
    g1416_p_spl_,
    g1416_p
  );


  buf

  (
    g1393_n_spl_,
    g1393_n
  );


  buf

  (
    g1418_p_spl_,
    g1418_p
  );


  buf

  (
    g1393_p_spl_,
    g1393_p
  );


  buf

  (
    g1418_n_spl_,
    g1418_n
  );


  buf

  (
    g1419_n_spl_,
    g1419_n
  );


  buf

  (
    g1419_p_spl_,
    g1419_p
  );


  buf

  (
    g1392_n_spl_,
    g1392_n
  );


  buf

  (
    g1421_p_spl_,
    g1421_p
  );


  buf

  (
    g1392_p_spl_,
    g1392_p
  );


  buf

  (
    g1421_n_spl_,
    g1421_n
  );


  buf

  (
    g1422_n_spl_,
    g1422_n
  );


  buf

  (
    g1422_p_spl_,
    g1422_p
  );


  buf

  (
    g1391_n_spl_,
    g1391_n
  );


  buf

  (
    g1424_p_spl_,
    g1424_p
  );


  buf

  (
    g1391_p_spl_,
    g1391_p
  );


  buf

  (
    g1424_n_spl_,
    g1424_n
  );


  buf

  (
    g1425_n_spl_,
    g1425_n
  );


  buf

  (
    g1425_p_spl_,
    g1425_p
  );


  buf

  (
    g1390_n_spl_,
    g1390_n
  );


  buf

  (
    g1427_p_spl_,
    g1427_p
  );


  buf

  (
    g1390_p_spl_,
    g1390_p
  );


  buf

  (
    g1427_n_spl_,
    g1427_n
  );


  buf

  (
    g1428_n_spl_,
    g1428_n
  );


  buf

  (
    g1428_p_spl_,
    g1428_p
  );


  buf

  (
    g1389_n_spl_,
    g1389_n
  );


  buf

  (
    g1430_p_spl_,
    g1430_p
  );


  buf

  (
    g1389_p_spl_,
    g1389_p
  );


  buf

  (
    g1430_n_spl_,
    g1430_n
  );


  buf

  (
    g1431_n_spl_,
    g1431_n
  );


  buf

  (
    g1431_p_spl_,
    g1431_p
  );


  buf

  (
    g1388_n_spl_,
    g1388_n
  );


  buf

  (
    g1433_p_spl_,
    g1433_p
  );


  buf

  (
    g1388_p_spl_,
    g1388_p
  );


  buf

  (
    g1433_n_spl_,
    g1433_n
  );


  buf

  (
    g1434_n_spl_,
    g1434_n
  );


  buf

  (
    g1434_p_spl_,
    g1434_p
  );


  buf

  (
    g1387_n_spl_,
    g1387_n
  );


  buf

  (
    g1436_p_spl_,
    g1436_p
  );


  buf

  (
    g1387_p_spl_,
    g1387_p
  );


  buf

  (
    g1436_n_spl_,
    g1436_n
  );


  buf

  (
    g1437_n_spl_,
    g1437_n
  );


  buf

  (
    g1437_p_spl_,
    g1437_p
  );


  buf

  (
    g1386_n_spl_,
    g1386_n
  );


  buf

  (
    g1439_p_spl_,
    g1439_p
  );


  buf

  (
    g1386_p_spl_,
    g1386_p
  );


  buf

  (
    g1439_n_spl_,
    g1439_n
  );


  buf

  (
    g1440_n_spl_,
    g1440_n
  );


  buf

  (
    g1440_p_spl_,
    g1440_p
  );


  buf

  (
    g1385_n_spl_,
    g1385_n
  );


  buf

  (
    g1442_p_spl_,
    g1442_p
  );


  buf

  (
    g1385_p_spl_,
    g1385_p
  );


  buf

  (
    g1442_n_spl_,
    g1442_n
  );


  buf

  (
    g1443_n_spl_,
    g1443_n
  );


  buf

  (
    g1443_p_spl_,
    g1443_p
  );


  buf

  (
    g1384_n_spl_,
    g1384_n
  );


  buf

  (
    g1445_p_spl_,
    g1445_p
  );


  buf

  (
    g1384_p_spl_,
    g1384_p
  );


  buf

  (
    g1445_n_spl_,
    g1445_n
  );


  buf

  (
    g1446_n_spl_,
    g1446_n
  );


  buf

  (
    g1446_p_spl_,
    g1446_p
  );


  buf

  (
    g1383_n_spl_,
    g1383_n
  );


  buf

  (
    g1448_p_spl_,
    g1448_p
  );


  buf

  (
    g1383_p_spl_,
    g1383_p
  );


  buf

  (
    g1448_n_spl_,
    g1448_n
  );


  buf

  (
    g1449_n_spl_,
    g1449_n
  );


  buf

  (
    g1449_p_spl_,
    g1449_p
  );


  buf

  (
    g1382_n_spl_,
    g1382_n
  );


  buf

  (
    g1451_p_spl_,
    g1451_p
  );


  buf

  (
    g1382_p_spl_,
    g1382_p
  );


  buf

  (
    g1451_n_spl_,
    g1451_n
  );


  buf

  (
    g1452_n_spl_,
    g1452_n
  );


  buf

  (
    g1452_p_spl_,
    g1452_p
  );


  buf

  (
    g1381_n_spl_,
    g1381_n
  );


  buf

  (
    g1454_p_spl_,
    g1454_p
  );


  buf

  (
    g1381_p_spl_,
    g1381_p
  );


  buf

  (
    g1454_n_spl_,
    g1454_n
  );


  buf

  (
    g1455_n_spl_,
    g1455_n
  );


  buf

  (
    g1455_p_spl_,
    g1455_p
  );


  buf

  (
    g1380_n_spl_,
    g1380_n
  );


  buf

  (
    g1457_p_spl_,
    g1457_p
  );


  buf

  (
    g1380_p_spl_,
    g1380_p
  );


  buf

  (
    g1457_n_spl_,
    g1457_n
  );


  buf

  (
    g1458_n_spl_,
    g1458_n
  );


  buf

  (
    g1458_p_spl_,
    g1458_p
  );


  buf

  (
    g1379_n_spl_,
    g1379_n
  );


  buf

  (
    g1460_p_spl_,
    g1460_p
  );


  buf

  (
    g1379_p_spl_,
    g1379_p
  );


  buf

  (
    g1460_n_spl_,
    g1460_n
  );


  buf

  (
    g1461_n_spl_,
    g1461_n
  );


  buf

  (
    g1461_p_spl_,
    g1461_p
  );


  buf

  (
    g1378_p_spl_,
    g1378_p
  );


  buf

  (
    g1463_n_spl_,
    g1463_n
  );


  buf

  (
    g1464_p_spl_,
    g1464_p
  );


  buf

  (
    g1486_n_spl_,
    g1486_n
  );


  buf

  (
    g1487_n_spl_,
    g1487_n
  );


  buf

  (
    g1486_p_spl_,
    g1486_p
  );


  buf

  (
    g1487_p_spl_,
    g1487_p
  );


  buf

  (
    g1488_n_spl_,
    g1488_n
  );


  buf

  (
    g1488_p_spl_,
    g1488_p
  );


  buf

  (
    g1485_n_spl_,
    g1485_n
  );


  buf

  (
    g1490_p_spl_,
    g1490_p
  );


  buf

  (
    g1485_p_spl_,
    g1485_p
  );


  buf

  (
    g1490_n_spl_,
    g1490_n
  );


  buf

  (
    g1491_n_spl_,
    g1491_n
  );


  buf

  (
    g1491_p_spl_,
    g1491_p
  );


  buf

  (
    g1484_n_spl_,
    g1484_n
  );


  buf

  (
    g1493_p_spl_,
    g1493_p
  );


  buf

  (
    g1484_p_spl_,
    g1484_p
  );


  buf

  (
    g1493_n_spl_,
    g1493_n
  );


  buf

  (
    g1494_n_spl_,
    g1494_n
  );


  buf

  (
    g1494_p_spl_,
    g1494_p
  );


  buf

  (
    g1483_n_spl_,
    g1483_n
  );


  buf

  (
    g1496_p_spl_,
    g1496_p
  );


  buf

  (
    g1483_p_spl_,
    g1483_p
  );


  buf

  (
    g1496_n_spl_,
    g1496_n
  );


  buf

  (
    g1497_n_spl_,
    g1497_n
  );


  buf

  (
    g1497_p_spl_,
    g1497_p
  );


  buf

  (
    g1482_n_spl_,
    g1482_n
  );


  buf

  (
    g1499_p_spl_,
    g1499_p
  );


  buf

  (
    g1482_p_spl_,
    g1482_p
  );


  buf

  (
    g1499_n_spl_,
    g1499_n
  );


  buf

  (
    g1500_n_spl_,
    g1500_n
  );


  buf

  (
    g1500_p_spl_,
    g1500_p
  );


  buf

  (
    g1481_n_spl_,
    g1481_n
  );


  buf

  (
    g1502_p_spl_,
    g1502_p
  );


  buf

  (
    g1481_p_spl_,
    g1481_p
  );


  buf

  (
    g1502_n_spl_,
    g1502_n
  );


  buf

  (
    g1503_n_spl_,
    g1503_n
  );


  buf

  (
    g1503_p_spl_,
    g1503_p
  );


  buf

  (
    g1480_n_spl_,
    g1480_n
  );


  buf

  (
    g1505_p_spl_,
    g1505_p
  );


  buf

  (
    g1480_p_spl_,
    g1480_p
  );


  buf

  (
    g1505_n_spl_,
    g1505_n
  );


  buf

  (
    g1506_n_spl_,
    g1506_n
  );


  buf

  (
    g1506_p_spl_,
    g1506_p
  );


  buf

  (
    g1479_n_spl_,
    g1479_n
  );


  buf

  (
    g1508_p_spl_,
    g1508_p
  );


  buf

  (
    g1479_p_spl_,
    g1479_p
  );


  buf

  (
    g1508_n_spl_,
    g1508_n
  );


  buf

  (
    g1509_n_spl_,
    g1509_n
  );


  buf

  (
    g1509_p_spl_,
    g1509_p
  );


  buf

  (
    g1478_n_spl_,
    g1478_n
  );


  buf

  (
    g1511_p_spl_,
    g1511_p
  );


  buf

  (
    g1478_p_spl_,
    g1478_p
  );


  buf

  (
    g1511_n_spl_,
    g1511_n
  );


  buf

  (
    g1512_n_spl_,
    g1512_n
  );


  buf

  (
    g1512_p_spl_,
    g1512_p
  );


  buf

  (
    g1477_n_spl_,
    g1477_n
  );


  buf

  (
    g1514_p_spl_,
    g1514_p
  );


  buf

  (
    g1477_p_spl_,
    g1477_p
  );


  buf

  (
    g1514_n_spl_,
    g1514_n
  );


  buf

  (
    g1515_n_spl_,
    g1515_n
  );


  buf

  (
    g1515_p_spl_,
    g1515_p
  );


  buf

  (
    g1476_n_spl_,
    g1476_n
  );


  buf

  (
    g1517_p_spl_,
    g1517_p
  );


  buf

  (
    g1476_p_spl_,
    g1476_p
  );


  buf

  (
    g1517_n_spl_,
    g1517_n
  );


  buf

  (
    g1518_n_spl_,
    g1518_n
  );


  buf

  (
    g1518_p_spl_,
    g1518_p
  );


  buf

  (
    g1475_n_spl_,
    g1475_n
  );


  buf

  (
    g1520_p_spl_,
    g1520_p
  );


  buf

  (
    g1475_p_spl_,
    g1475_p
  );


  buf

  (
    g1520_n_spl_,
    g1520_n
  );


  buf

  (
    g1521_n_spl_,
    g1521_n
  );


  buf

  (
    g1521_p_spl_,
    g1521_p
  );


  buf

  (
    g1474_n_spl_,
    g1474_n
  );


  buf

  (
    g1523_p_spl_,
    g1523_p
  );


  buf

  (
    g1474_p_spl_,
    g1474_p
  );


  buf

  (
    g1523_n_spl_,
    g1523_n
  );


  buf

  (
    g1524_n_spl_,
    g1524_n
  );


  buf

  (
    g1524_p_spl_,
    g1524_p
  );


  buf

  (
    g1473_n_spl_,
    g1473_n
  );


  buf

  (
    g1526_p_spl_,
    g1526_p
  );


  buf

  (
    g1473_p_spl_,
    g1473_p
  );


  buf

  (
    g1526_n_spl_,
    g1526_n
  );


  buf

  (
    g1527_n_spl_,
    g1527_n
  );


  buf

  (
    g1527_p_spl_,
    g1527_p
  );


  buf

  (
    g1472_n_spl_,
    g1472_n
  );


  buf

  (
    g1529_p_spl_,
    g1529_p
  );


  buf

  (
    g1472_p_spl_,
    g1472_p
  );


  buf

  (
    g1529_n_spl_,
    g1529_n
  );


  buf

  (
    g1530_n_spl_,
    g1530_n
  );


  buf

  (
    g1530_p_spl_,
    g1530_p
  );


  buf

  (
    g1471_n_spl_,
    g1471_n
  );


  buf

  (
    g1532_p_spl_,
    g1532_p
  );


  buf

  (
    g1471_p_spl_,
    g1471_p
  );


  buf

  (
    g1532_n_spl_,
    g1532_n
  );


  buf

  (
    g1533_n_spl_,
    g1533_n
  );


  buf

  (
    g1533_p_spl_,
    g1533_p
  );


  buf

  (
    g1470_n_spl_,
    g1470_n
  );


  buf

  (
    g1535_p_spl_,
    g1535_p
  );


  buf

  (
    g1470_p_spl_,
    g1470_p
  );


  buf

  (
    g1535_n_spl_,
    g1535_n
  );


  buf

  (
    g1536_n_spl_,
    g1536_n
  );


  buf

  (
    g1536_p_spl_,
    g1536_p
  );


  buf

  (
    g1469_n_spl_,
    g1469_n
  );


  buf

  (
    g1538_p_spl_,
    g1538_p
  );


  buf

  (
    g1469_p_spl_,
    g1469_p
  );


  buf

  (
    g1538_n_spl_,
    g1538_n
  );


  buf

  (
    g1539_n_spl_,
    g1539_n
  );


  buf

  (
    g1539_p_spl_,
    g1539_p
  );


  buf

  (
    g1468_n_spl_,
    g1468_n
  );


  buf

  (
    g1541_p_spl_,
    g1541_p
  );


  buf

  (
    g1468_p_spl_,
    g1468_p
  );


  buf

  (
    g1541_n_spl_,
    g1541_n
  );


  buf

  (
    g1542_n_spl_,
    g1542_n
  );


  buf

  (
    g1542_p_spl_,
    g1542_p
  );


  buf

  (
    g1467_p_spl_,
    g1467_p
  );


  buf

  (
    g1544_n_spl_,
    g1544_n
  );


  buf

  (
    g1545_p_spl_,
    g1545_p
  );


  buf

  (
    g1565_n_spl_,
    g1565_n
  );


  buf

  (
    g1566_n_spl_,
    g1566_n
  );


  buf

  (
    g1565_p_spl_,
    g1565_p
  );


  buf

  (
    g1566_p_spl_,
    g1566_p
  );


  buf

  (
    g1567_n_spl_,
    g1567_n
  );


  buf

  (
    g1567_p_spl_,
    g1567_p
  );


  buf

  (
    g1564_n_spl_,
    g1564_n
  );


  buf

  (
    g1569_p_spl_,
    g1569_p
  );


  buf

  (
    g1564_p_spl_,
    g1564_p
  );


  buf

  (
    g1569_n_spl_,
    g1569_n
  );


  buf

  (
    g1570_n_spl_,
    g1570_n
  );


  buf

  (
    g1570_p_spl_,
    g1570_p
  );


  buf

  (
    g1563_n_spl_,
    g1563_n
  );


  buf

  (
    g1572_p_spl_,
    g1572_p
  );


  buf

  (
    g1563_p_spl_,
    g1563_p
  );


  buf

  (
    g1572_n_spl_,
    g1572_n
  );


  buf

  (
    g1573_n_spl_,
    g1573_n
  );


  buf

  (
    g1573_p_spl_,
    g1573_p
  );


  buf

  (
    g1562_n_spl_,
    g1562_n
  );


  buf

  (
    g1575_p_spl_,
    g1575_p
  );


  buf

  (
    g1562_p_spl_,
    g1562_p
  );


  buf

  (
    g1575_n_spl_,
    g1575_n
  );


  buf

  (
    g1576_n_spl_,
    g1576_n
  );


  buf

  (
    g1576_p_spl_,
    g1576_p
  );


  buf

  (
    g1561_n_spl_,
    g1561_n
  );


  buf

  (
    g1578_p_spl_,
    g1578_p
  );


  buf

  (
    g1561_p_spl_,
    g1561_p
  );


  buf

  (
    g1578_n_spl_,
    g1578_n
  );


  buf

  (
    g1579_n_spl_,
    g1579_n
  );


  buf

  (
    g1579_p_spl_,
    g1579_p
  );


  buf

  (
    g1560_n_spl_,
    g1560_n
  );


  buf

  (
    g1581_p_spl_,
    g1581_p
  );


  buf

  (
    g1560_p_spl_,
    g1560_p
  );


  buf

  (
    g1581_n_spl_,
    g1581_n
  );


  buf

  (
    g1582_n_spl_,
    g1582_n
  );


  buf

  (
    g1582_p_spl_,
    g1582_p
  );


  buf

  (
    g1559_n_spl_,
    g1559_n
  );


  buf

  (
    g1584_p_spl_,
    g1584_p
  );


  buf

  (
    g1559_p_spl_,
    g1559_p
  );


  buf

  (
    g1584_n_spl_,
    g1584_n
  );


  buf

  (
    g1585_n_spl_,
    g1585_n
  );


  buf

  (
    g1585_p_spl_,
    g1585_p
  );


  buf

  (
    g1558_n_spl_,
    g1558_n
  );


  buf

  (
    g1587_p_spl_,
    g1587_p
  );


  buf

  (
    g1558_p_spl_,
    g1558_p
  );


  buf

  (
    g1587_n_spl_,
    g1587_n
  );


  buf

  (
    g1588_n_spl_,
    g1588_n
  );


  buf

  (
    g1588_p_spl_,
    g1588_p
  );


  buf

  (
    g1557_n_spl_,
    g1557_n
  );


  buf

  (
    g1590_p_spl_,
    g1590_p
  );


  buf

  (
    g1557_p_spl_,
    g1557_p
  );


  buf

  (
    g1590_n_spl_,
    g1590_n
  );


  buf

  (
    g1591_n_spl_,
    g1591_n
  );


  buf

  (
    g1591_p_spl_,
    g1591_p
  );


  buf

  (
    g1556_n_spl_,
    g1556_n
  );


  buf

  (
    g1593_p_spl_,
    g1593_p
  );


  buf

  (
    g1556_p_spl_,
    g1556_p
  );


  buf

  (
    g1593_n_spl_,
    g1593_n
  );


  buf

  (
    g1594_n_spl_,
    g1594_n
  );


  buf

  (
    g1594_p_spl_,
    g1594_p
  );


  buf

  (
    g1555_n_spl_,
    g1555_n
  );


  buf

  (
    g1596_p_spl_,
    g1596_p
  );


  buf

  (
    g1555_p_spl_,
    g1555_p
  );


  buf

  (
    g1596_n_spl_,
    g1596_n
  );


  buf

  (
    g1597_n_spl_,
    g1597_n
  );


  buf

  (
    g1597_p_spl_,
    g1597_p
  );


  buf

  (
    g1554_n_spl_,
    g1554_n
  );


  buf

  (
    g1599_p_spl_,
    g1599_p
  );


  buf

  (
    g1554_p_spl_,
    g1554_p
  );


  buf

  (
    g1599_n_spl_,
    g1599_n
  );


  buf

  (
    g1600_n_spl_,
    g1600_n
  );


  buf

  (
    g1600_p_spl_,
    g1600_p
  );


  buf

  (
    g1553_n_spl_,
    g1553_n
  );


  buf

  (
    g1602_p_spl_,
    g1602_p
  );


  buf

  (
    g1553_p_spl_,
    g1553_p
  );


  buf

  (
    g1602_n_spl_,
    g1602_n
  );


  buf

  (
    g1603_n_spl_,
    g1603_n
  );


  buf

  (
    g1603_p_spl_,
    g1603_p
  );


  buf

  (
    g1552_n_spl_,
    g1552_n
  );


  buf

  (
    g1605_p_spl_,
    g1605_p
  );


  buf

  (
    g1552_p_spl_,
    g1552_p
  );


  buf

  (
    g1605_n_spl_,
    g1605_n
  );


  buf

  (
    g1606_n_spl_,
    g1606_n
  );


  buf

  (
    g1606_p_spl_,
    g1606_p
  );


  buf

  (
    g1551_n_spl_,
    g1551_n
  );


  buf

  (
    g1608_p_spl_,
    g1608_p
  );


  buf

  (
    g1551_p_spl_,
    g1551_p
  );


  buf

  (
    g1608_n_spl_,
    g1608_n
  );


  buf

  (
    g1609_n_spl_,
    g1609_n
  );


  buf

  (
    g1609_p_spl_,
    g1609_p
  );


  buf

  (
    g1550_n_spl_,
    g1550_n
  );


  buf

  (
    g1611_p_spl_,
    g1611_p
  );


  buf

  (
    g1550_p_spl_,
    g1550_p
  );


  buf

  (
    g1611_n_spl_,
    g1611_n
  );


  buf

  (
    g1612_n_spl_,
    g1612_n
  );


  buf

  (
    g1612_p_spl_,
    g1612_p
  );


  buf

  (
    g1549_n_spl_,
    g1549_n
  );


  buf

  (
    g1614_p_spl_,
    g1614_p
  );


  buf

  (
    g1549_p_spl_,
    g1549_p
  );


  buf

  (
    g1614_n_spl_,
    g1614_n
  );


  buf

  (
    g1615_n_spl_,
    g1615_n
  );


  buf

  (
    g1615_p_spl_,
    g1615_p
  );


  buf

  (
    g1548_p_spl_,
    g1548_p
  );


  buf

  (
    g1617_n_spl_,
    g1617_n
  );


  buf

  (
    g1618_p_spl_,
    g1618_p
  );


  buf

  (
    g1636_n_spl_,
    g1636_n
  );


  buf

  (
    g1637_n_spl_,
    g1637_n
  );


  buf

  (
    g1636_p_spl_,
    g1636_p
  );


  buf

  (
    g1637_p_spl_,
    g1637_p
  );


  buf

  (
    g1638_n_spl_,
    g1638_n
  );


  buf

  (
    g1638_p_spl_,
    g1638_p
  );


  buf

  (
    g1635_n_spl_,
    g1635_n
  );


  buf

  (
    g1640_p_spl_,
    g1640_p
  );


  buf

  (
    g1635_p_spl_,
    g1635_p
  );


  buf

  (
    g1640_n_spl_,
    g1640_n
  );


  buf

  (
    g1641_n_spl_,
    g1641_n
  );


  buf

  (
    g1641_p_spl_,
    g1641_p
  );


  buf

  (
    g1634_n_spl_,
    g1634_n
  );


  buf

  (
    g1643_p_spl_,
    g1643_p
  );


  buf

  (
    g1634_p_spl_,
    g1634_p
  );


  buf

  (
    g1643_n_spl_,
    g1643_n
  );


  buf

  (
    g1644_n_spl_,
    g1644_n
  );


  buf

  (
    g1644_p_spl_,
    g1644_p
  );


  buf

  (
    g1633_n_spl_,
    g1633_n
  );


  buf

  (
    g1646_p_spl_,
    g1646_p
  );


  buf

  (
    g1633_p_spl_,
    g1633_p
  );


  buf

  (
    g1646_n_spl_,
    g1646_n
  );


  buf

  (
    g1647_n_spl_,
    g1647_n
  );


  buf

  (
    g1647_p_spl_,
    g1647_p
  );


  buf

  (
    g1632_n_spl_,
    g1632_n
  );


  buf

  (
    g1649_p_spl_,
    g1649_p
  );


  buf

  (
    g1632_p_spl_,
    g1632_p
  );


  buf

  (
    g1649_n_spl_,
    g1649_n
  );


  buf

  (
    g1650_n_spl_,
    g1650_n
  );


  buf

  (
    g1650_p_spl_,
    g1650_p
  );


  buf

  (
    g1631_n_spl_,
    g1631_n
  );


  buf

  (
    g1652_p_spl_,
    g1652_p
  );


  buf

  (
    g1631_p_spl_,
    g1631_p
  );


  buf

  (
    g1652_n_spl_,
    g1652_n
  );


  buf

  (
    g1653_n_spl_,
    g1653_n
  );


  buf

  (
    g1653_p_spl_,
    g1653_p
  );


  buf

  (
    g1630_n_spl_,
    g1630_n
  );


  buf

  (
    g1655_p_spl_,
    g1655_p
  );


  buf

  (
    g1630_p_spl_,
    g1630_p
  );


  buf

  (
    g1655_n_spl_,
    g1655_n
  );


  buf

  (
    g1656_n_spl_,
    g1656_n
  );


  buf

  (
    g1656_p_spl_,
    g1656_p
  );


  buf

  (
    g1629_n_spl_,
    g1629_n
  );


  buf

  (
    g1658_p_spl_,
    g1658_p
  );


  buf

  (
    g1629_p_spl_,
    g1629_p
  );


  buf

  (
    g1658_n_spl_,
    g1658_n
  );


  buf

  (
    g1659_n_spl_,
    g1659_n
  );


  buf

  (
    g1659_p_spl_,
    g1659_p
  );


  buf

  (
    g1628_n_spl_,
    g1628_n
  );


  buf

  (
    g1661_p_spl_,
    g1661_p
  );


  buf

  (
    g1628_p_spl_,
    g1628_p
  );


  buf

  (
    g1661_n_spl_,
    g1661_n
  );


  buf

  (
    g1662_n_spl_,
    g1662_n
  );


  buf

  (
    g1662_p_spl_,
    g1662_p
  );


  buf

  (
    g1627_n_spl_,
    g1627_n
  );


  buf

  (
    g1664_p_spl_,
    g1664_p
  );


  buf

  (
    g1627_p_spl_,
    g1627_p
  );


  buf

  (
    g1664_n_spl_,
    g1664_n
  );


  buf

  (
    g1665_n_spl_,
    g1665_n
  );


  buf

  (
    g1665_p_spl_,
    g1665_p
  );


  buf

  (
    g1626_n_spl_,
    g1626_n
  );


  buf

  (
    g1667_p_spl_,
    g1667_p
  );


  buf

  (
    g1626_p_spl_,
    g1626_p
  );


  buf

  (
    g1667_n_spl_,
    g1667_n
  );


  buf

  (
    g1668_n_spl_,
    g1668_n
  );


  buf

  (
    g1668_p_spl_,
    g1668_p
  );


  buf

  (
    g1625_n_spl_,
    g1625_n
  );


  buf

  (
    g1670_p_spl_,
    g1670_p
  );


  buf

  (
    g1625_p_spl_,
    g1625_p
  );


  buf

  (
    g1670_n_spl_,
    g1670_n
  );


  buf

  (
    g1671_n_spl_,
    g1671_n
  );


  buf

  (
    g1671_p_spl_,
    g1671_p
  );


  buf

  (
    g1624_n_spl_,
    g1624_n
  );


  buf

  (
    g1673_p_spl_,
    g1673_p
  );


  buf

  (
    g1624_p_spl_,
    g1624_p
  );


  buf

  (
    g1673_n_spl_,
    g1673_n
  );


  buf

  (
    g1674_n_spl_,
    g1674_n
  );


  buf

  (
    g1674_p_spl_,
    g1674_p
  );


  buf

  (
    g1623_n_spl_,
    g1623_n
  );


  buf

  (
    g1676_p_spl_,
    g1676_p
  );


  buf

  (
    g1623_p_spl_,
    g1623_p
  );


  buf

  (
    g1676_n_spl_,
    g1676_n
  );


  buf

  (
    g1677_n_spl_,
    g1677_n
  );


  buf

  (
    g1677_p_spl_,
    g1677_p
  );


  buf

  (
    g1622_n_spl_,
    g1622_n
  );


  buf

  (
    g1679_p_spl_,
    g1679_p
  );


  buf

  (
    g1622_p_spl_,
    g1622_p
  );


  buf

  (
    g1679_n_spl_,
    g1679_n
  );


  buf

  (
    g1680_n_spl_,
    g1680_n
  );


  buf

  (
    g1680_p_spl_,
    g1680_p
  );


  buf

  (
    g1621_p_spl_,
    g1621_p
  );


  buf

  (
    g1682_n_spl_,
    g1682_n
  );


  buf

  (
    g1683_p_spl_,
    g1683_p
  );


  buf

  (
    g1699_n_spl_,
    g1699_n
  );


  buf

  (
    g1700_n_spl_,
    g1700_n
  );


  buf

  (
    g1699_p_spl_,
    g1699_p
  );


  buf

  (
    g1700_p_spl_,
    g1700_p
  );


  buf

  (
    g1701_n_spl_,
    g1701_n
  );


  buf

  (
    g1701_p_spl_,
    g1701_p
  );


  buf

  (
    g1698_n_spl_,
    g1698_n
  );


  buf

  (
    g1703_p_spl_,
    g1703_p
  );


  buf

  (
    g1698_p_spl_,
    g1698_p
  );


  buf

  (
    g1703_n_spl_,
    g1703_n
  );


  buf

  (
    g1704_n_spl_,
    g1704_n
  );


  buf

  (
    g1704_p_spl_,
    g1704_p
  );


  buf

  (
    g1697_n_spl_,
    g1697_n
  );


  buf

  (
    g1706_p_spl_,
    g1706_p
  );


  buf

  (
    g1697_p_spl_,
    g1697_p
  );


  buf

  (
    g1706_n_spl_,
    g1706_n
  );


  buf

  (
    g1707_n_spl_,
    g1707_n
  );


  buf

  (
    g1707_p_spl_,
    g1707_p
  );


  buf

  (
    g1696_n_spl_,
    g1696_n
  );


  buf

  (
    g1709_p_spl_,
    g1709_p
  );


  buf

  (
    g1696_p_spl_,
    g1696_p
  );


  buf

  (
    g1709_n_spl_,
    g1709_n
  );


  buf

  (
    g1710_n_spl_,
    g1710_n
  );


  buf

  (
    g1710_p_spl_,
    g1710_p
  );


  buf

  (
    g1695_n_spl_,
    g1695_n
  );


  buf

  (
    g1712_p_spl_,
    g1712_p
  );


  buf

  (
    g1695_p_spl_,
    g1695_p
  );


  buf

  (
    g1712_n_spl_,
    g1712_n
  );


  buf

  (
    g1713_n_spl_,
    g1713_n
  );


  buf

  (
    g1713_p_spl_,
    g1713_p
  );


  buf

  (
    g1694_n_spl_,
    g1694_n
  );


  buf

  (
    g1715_p_spl_,
    g1715_p
  );


  buf

  (
    g1694_p_spl_,
    g1694_p
  );


  buf

  (
    g1715_n_spl_,
    g1715_n
  );


  buf

  (
    g1716_n_spl_,
    g1716_n
  );


  buf

  (
    g1716_p_spl_,
    g1716_p
  );


  buf

  (
    g1693_n_spl_,
    g1693_n
  );


  buf

  (
    g1718_p_spl_,
    g1718_p
  );


  buf

  (
    g1693_p_spl_,
    g1693_p
  );


  buf

  (
    g1718_n_spl_,
    g1718_n
  );


  buf

  (
    g1719_n_spl_,
    g1719_n
  );


  buf

  (
    g1719_p_spl_,
    g1719_p
  );


  buf

  (
    g1692_n_spl_,
    g1692_n
  );


  buf

  (
    g1721_p_spl_,
    g1721_p
  );


  buf

  (
    g1692_p_spl_,
    g1692_p
  );


  buf

  (
    g1721_n_spl_,
    g1721_n
  );


  buf

  (
    g1722_n_spl_,
    g1722_n
  );


  buf

  (
    g1722_p_spl_,
    g1722_p
  );


  buf

  (
    g1691_n_spl_,
    g1691_n
  );


  buf

  (
    g1724_p_spl_,
    g1724_p
  );


  buf

  (
    g1691_p_spl_,
    g1691_p
  );


  buf

  (
    g1724_n_spl_,
    g1724_n
  );


  buf

  (
    g1725_n_spl_,
    g1725_n
  );


  buf

  (
    g1725_p_spl_,
    g1725_p
  );


  buf

  (
    g1690_n_spl_,
    g1690_n
  );


  buf

  (
    g1727_p_spl_,
    g1727_p
  );


  buf

  (
    g1690_p_spl_,
    g1690_p
  );


  buf

  (
    g1727_n_spl_,
    g1727_n
  );


  buf

  (
    g1728_n_spl_,
    g1728_n
  );


  buf

  (
    g1728_p_spl_,
    g1728_p
  );


  buf

  (
    g1689_n_spl_,
    g1689_n
  );


  buf

  (
    g1730_p_spl_,
    g1730_p
  );


  buf

  (
    g1689_p_spl_,
    g1689_p
  );


  buf

  (
    g1730_n_spl_,
    g1730_n
  );


  buf

  (
    g1731_n_spl_,
    g1731_n
  );


  buf

  (
    g1731_p_spl_,
    g1731_p
  );


  buf

  (
    g1688_n_spl_,
    g1688_n
  );


  buf

  (
    g1733_p_spl_,
    g1733_p
  );


  buf

  (
    g1688_p_spl_,
    g1688_p
  );


  buf

  (
    g1733_n_spl_,
    g1733_n
  );


  buf

  (
    g1734_n_spl_,
    g1734_n
  );


  buf

  (
    g1734_p_spl_,
    g1734_p
  );


  buf

  (
    g1687_n_spl_,
    g1687_n
  );


  buf

  (
    g1736_p_spl_,
    g1736_p
  );


  buf

  (
    g1687_p_spl_,
    g1687_p
  );


  buf

  (
    g1736_n_spl_,
    g1736_n
  );


  buf

  (
    g1737_n_spl_,
    g1737_n
  );


  buf

  (
    g1737_p_spl_,
    g1737_p
  );


  buf

  (
    g1686_p_spl_,
    g1686_p
  );


  buf

  (
    g1739_n_spl_,
    g1739_n
  );


  buf

  (
    g1740_p_spl_,
    g1740_p
  );


  buf

  (
    g1754_n_spl_,
    g1754_n
  );


  buf

  (
    g1755_n_spl_,
    g1755_n
  );


  buf

  (
    g1754_p_spl_,
    g1754_p
  );


  buf

  (
    g1755_p_spl_,
    g1755_p
  );


  buf

  (
    g1756_n_spl_,
    g1756_n
  );


  buf

  (
    g1756_p_spl_,
    g1756_p
  );


  buf

  (
    g1753_n_spl_,
    g1753_n
  );


  buf

  (
    g1758_p_spl_,
    g1758_p
  );


  buf

  (
    g1753_p_spl_,
    g1753_p
  );


  buf

  (
    g1758_n_spl_,
    g1758_n
  );


  buf

  (
    g1759_n_spl_,
    g1759_n
  );


  buf

  (
    g1759_p_spl_,
    g1759_p
  );


  buf

  (
    g1752_n_spl_,
    g1752_n
  );


  buf

  (
    g1761_p_spl_,
    g1761_p
  );


  buf

  (
    g1752_p_spl_,
    g1752_p
  );


  buf

  (
    g1761_n_spl_,
    g1761_n
  );


  buf

  (
    g1762_n_spl_,
    g1762_n
  );


  buf

  (
    g1762_p_spl_,
    g1762_p
  );


  buf

  (
    g1751_n_spl_,
    g1751_n
  );


  buf

  (
    g1764_p_spl_,
    g1764_p
  );


  buf

  (
    g1751_p_spl_,
    g1751_p
  );


  buf

  (
    g1764_n_spl_,
    g1764_n
  );


  buf

  (
    g1765_n_spl_,
    g1765_n
  );


  buf

  (
    g1765_p_spl_,
    g1765_p
  );


  buf

  (
    g1750_n_spl_,
    g1750_n
  );


  buf

  (
    g1767_p_spl_,
    g1767_p
  );


  buf

  (
    g1750_p_spl_,
    g1750_p
  );


  buf

  (
    g1767_n_spl_,
    g1767_n
  );


  buf

  (
    g1768_n_spl_,
    g1768_n
  );


  buf

  (
    g1768_p_spl_,
    g1768_p
  );


  buf

  (
    g1749_n_spl_,
    g1749_n
  );


  buf

  (
    g1770_p_spl_,
    g1770_p
  );


  buf

  (
    g1749_p_spl_,
    g1749_p
  );


  buf

  (
    g1770_n_spl_,
    g1770_n
  );


  buf

  (
    g1771_n_spl_,
    g1771_n
  );


  buf

  (
    g1771_p_spl_,
    g1771_p
  );


  buf

  (
    g1748_n_spl_,
    g1748_n
  );


  buf

  (
    g1773_p_spl_,
    g1773_p
  );


  buf

  (
    g1748_p_spl_,
    g1748_p
  );


  buf

  (
    g1773_n_spl_,
    g1773_n
  );


  buf

  (
    g1774_n_spl_,
    g1774_n
  );


  buf

  (
    g1774_p_spl_,
    g1774_p
  );


  buf

  (
    g1747_n_spl_,
    g1747_n
  );


  buf

  (
    g1776_p_spl_,
    g1776_p
  );


  buf

  (
    g1747_p_spl_,
    g1747_p
  );


  buf

  (
    g1776_n_spl_,
    g1776_n
  );


  buf

  (
    g1777_n_spl_,
    g1777_n
  );


  buf

  (
    g1777_p_spl_,
    g1777_p
  );


  buf

  (
    g1746_n_spl_,
    g1746_n
  );


  buf

  (
    g1779_p_spl_,
    g1779_p
  );


  buf

  (
    g1746_p_spl_,
    g1746_p
  );


  buf

  (
    g1779_n_spl_,
    g1779_n
  );


  buf

  (
    g1780_n_spl_,
    g1780_n
  );


  buf

  (
    g1780_p_spl_,
    g1780_p
  );


  buf

  (
    g1745_n_spl_,
    g1745_n
  );


  buf

  (
    g1782_p_spl_,
    g1782_p
  );


  buf

  (
    g1745_p_spl_,
    g1745_p
  );


  buf

  (
    g1782_n_spl_,
    g1782_n
  );


  buf

  (
    g1783_n_spl_,
    g1783_n
  );


  buf

  (
    g1783_p_spl_,
    g1783_p
  );


  buf

  (
    g1744_n_spl_,
    g1744_n
  );


  buf

  (
    g1785_p_spl_,
    g1785_p
  );


  buf

  (
    g1744_p_spl_,
    g1744_p
  );


  buf

  (
    g1785_n_spl_,
    g1785_n
  );


  buf

  (
    g1786_n_spl_,
    g1786_n
  );


  buf

  (
    g1786_p_spl_,
    g1786_p
  );


  buf

  (
    g1743_p_spl_,
    g1743_p
  );


  buf

  (
    g1788_n_spl_,
    g1788_n
  );


  buf

  (
    g1789_p_spl_,
    g1789_p
  );


  buf

  (
    g1801_n_spl_,
    g1801_n
  );


  buf

  (
    g1802_n_spl_,
    g1802_n
  );


  buf

  (
    g1801_p_spl_,
    g1801_p
  );


  buf

  (
    g1802_p_spl_,
    g1802_p
  );


  buf

  (
    g1803_n_spl_,
    g1803_n
  );


  buf

  (
    g1803_p_spl_,
    g1803_p
  );


  buf

  (
    g1800_n_spl_,
    g1800_n
  );


  buf

  (
    g1805_p_spl_,
    g1805_p
  );


  buf

  (
    g1800_p_spl_,
    g1800_p
  );


  buf

  (
    g1805_n_spl_,
    g1805_n
  );


  buf

  (
    g1806_n_spl_,
    g1806_n
  );


  buf

  (
    g1806_p_spl_,
    g1806_p
  );


  buf

  (
    g1799_n_spl_,
    g1799_n
  );


  buf

  (
    g1808_p_spl_,
    g1808_p
  );


  buf

  (
    g1799_p_spl_,
    g1799_p
  );


  buf

  (
    g1808_n_spl_,
    g1808_n
  );


  buf

  (
    g1809_n_spl_,
    g1809_n
  );


  buf

  (
    g1809_p_spl_,
    g1809_p
  );


  buf

  (
    g1798_n_spl_,
    g1798_n
  );


  buf

  (
    g1811_p_spl_,
    g1811_p
  );


  buf

  (
    g1798_p_spl_,
    g1798_p
  );


  buf

  (
    g1811_n_spl_,
    g1811_n
  );


  buf

  (
    g1812_n_spl_,
    g1812_n
  );


  buf

  (
    g1812_p_spl_,
    g1812_p
  );


  buf

  (
    g1797_n_spl_,
    g1797_n
  );


  buf

  (
    g1814_p_spl_,
    g1814_p
  );


  buf

  (
    g1797_p_spl_,
    g1797_p
  );


  buf

  (
    g1814_n_spl_,
    g1814_n
  );


  buf

  (
    g1815_n_spl_,
    g1815_n
  );


  buf

  (
    g1815_p_spl_,
    g1815_p
  );


  buf

  (
    g1796_n_spl_,
    g1796_n
  );


  buf

  (
    g1817_p_spl_,
    g1817_p
  );


  buf

  (
    g1796_p_spl_,
    g1796_p
  );


  buf

  (
    g1817_n_spl_,
    g1817_n
  );


  buf

  (
    g1818_n_spl_,
    g1818_n
  );


  buf

  (
    g1818_p_spl_,
    g1818_p
  );


  buf

  (
    g1795_n_spl_,
    g1795_n
  );


  buf

  (
    g1820_p_spl_,
    g1820_p
  );


  buf

  (
    g1795_p_spl_,
    g1795_p
  );


  buf

  (
    g1820_n_spl_,
    g1820_n
  );


  buf

  (
    g1821_n_spl_,
    g1821_n
  );


  buf

  (
    g1821_p_spl_,
    g1821_p
  );


  buf

  (
    g1794_n_spl_,
    g1794_n
  );


  buf

  (
    g1823_p_spl_,
    g1823_p
  );


  buf

  (
    g1794_p_spl_,
    g1794_p
  );


  buf

  (
    g1823_n_spl_,
    g1823_n
  );


  buf

  (
    g1824_n_spl_,
    g1824_n
  );


  buf

  (
    g1824_p_spl_,
    g1824_p
  );


  buf

  (
    g1793_n_spl_,
    g1793_n
  );


  buf

  (
    g1826_p_spl_,
    g1826_p
  );


  buf

  (
    g1793_p_spl_,
    g1793_p
  );


  buf

  (
    g1826_n_spl_,
    g1826_n
  );


  buf

  (
    g1827_n_spl_,
    g1827_n
  );


  buf

  (
    g1827_p_spl_,
    g1827_p
  );


  buf

  (
    g1792_p_spl_,
    g1792_p
  );


  buf

  (
    g1829_n_spl_,
    g1829_n
  );


  buf

  (
    g1830_p_spl_,
    g1830_p
  );


  buf

  (
    g1840_n_spl_,
    g1840_n
  );


  buf

  (
    g1841_n_spl_,
    g1841_n
  );


  buf

  (
    g1840_p_spl_,
    g1840_p
  );


  buf

  (
    g1841_p_spl_,
    g1841_p
  );


  buf

  (
    g1842_n_spl_,
    g1842_n
  );


  buf

  (
    g1842_p_spl_,
    g1842_p
  );


  buf

  (
    g1839_n_spl_,
    g1839_n
  );


  buf

  (
    g1844_p_spl_,
    g1844_p
  );


  buf

  (
    g1839_p_spl_,
    g1839_p
  );


  buf

  (
    g1844_n_spl_,
    g1844_n
  );


  buf

  (
    g1845_n_spl_,
    g1845_n
  );


  buf

  (
    g1845_p_spl_,
    g1845_p
  );


  buf

  (
    g1838_n_spl_,
    g1838_n
  );


  buf

  (
    g1847_p_spl_,
    g1847_p
  );


  buf

  (
    g1838_p_spl_,
    g1838_p
  );


  buf

  (
    g1847_n_spl_,
    g1847_n
  );


  buf

  (
    g1848_n_spl_,
    g1848_n
  );


  buf

  (
    g1848_p_spl_,
    g1848_p
  );


  buf

  (
    g1837_n_spl_,
    g1837_n
  );


  buf

  (
    g1850_p_spl_,
    g1850_p
  );


  buf

  (
    g1837_p_spl_,
    g1837_p
  );


  buf

  (
    g1850_n_spl_,
    g1850_n
  );


  buf

  (
    g1851_n_spl_,
    g1851_n
  );


  buf

  (
    g1851_p_spl_,
    g1851_p
  );


  buf

  (
    g1836_n_spl_,
    g1836_n
  );


  buf

  (
    g1853_p_spl_,
    g1853_p
  );


  buf

  (
    g1836_p_spl_,
    g1836_p
  );


  buf

  (
    g1853_n_spl_,
    g1853_n
  );


  buf

  (
    g1854_n_spl_,
    g1854_n
  );


  buf

  (
    g1854_p_spl_,
    g1854_p
  );


  buf

  (
    g1835_n_spl_,
    g1835_n
  );


  buf

  (
    g1856_p_spl_,
    g1856_p
  );


  buf

  (
    g1835_p_spl_,
    g1835_p
  );


  buf

  (
    g1856_n_spl_,
    g1856_n
  );


  buf

  (
    g1857_n_spl_,
    g1857_n
  );


  buf

  (
    g1857_p_spl_,
    g1857_p
  );


  buf

  (
    g1834_n_spl_,
    g1834_n
  );


  buf

  (
    g1859_p_spl_,
    g1859_p
  );


  buf

  (
    g1834_p_spl_,
    g1834_p
  );


  buf

  (
    g1859_n_spl_,
    g1859_n
  );


  buf

  (
    g1860_n_spl_,
    g1860_n
  );


  buf

  (
    g1860_p_spl_,
    g1860_p
  );


  buf

  (
    g1833_p_spl_,
    g1833_p
  );


  buf

  (
    g1862_n_spl_,
    g1862_n
  );


  buf

  (
    g1863_p_spl_,
    g1863_p
  );


  buf

  (
    g1871_n_spl_,
    g1871_n
  );


  buf

  (
    g1872_n_spl_,
    g1872_n
  );


  buf

  (
    g1871_p_spl_,
    g1871_p
  );


  buf

  (
    g1872_p_spl_,
    g1872_p
  );


  buf

  (
    g1873_n_spl_,
    g1873_n
  );


  buf

  (
    g1873_p_spl_,
    g1873_p
  );


  buf

  (
    g1870_n_spl_,
    g1870_n
  );


  buf

  (
    g1875_p_spl_,
    g1875_p
  );


  buf

  (
    g1870_p_spl_,
    g1870_p
  );


  buf

  (
    g1875_n_spl_,
    g1875_n
  );


  buf

  (
    g1876_n_spl_,
    g1876_n
  );


  buf

  (
    g1876_p_spl_,
    g1876_p
  );


  buf

  (
    g1869_n_spl_,
    g1869_n
  );


  buf

  (
    g1878_p_spl_,
    g1878_p
  );


  buf

  (
    g1869_p_spl_,
    g1869_p
  );


  buf

  (
    g1878_n_spl_,
    g1878_n
  );


  buf

  (
    g1879_n_spl_,
    g1879_n
  );


  buf

  (
    g1879_p_spl_,
    g1879_p
  );


  buf

  (
    g1868_n_spl_,
    g1868_n
  );


  buf

  (
    g1881_p_spl_,
    g1881_p
  );


  buf

  (
    g1868_p_spl_,
    g1868_p
  );


  buf

  (
    g1881_n_spl_,
    g1881_n
  );


  buf

  (
    g1882_n_spl_,
    g1882_n
  );


  buf

  (
    g1882_p_spl_,
    g1882_p
  );


  buf

  (
    g1867_n_spl_,
    g1867_n
  );


  buf

  (
    g1884_p_spl_,
    g1884_p
  );


  buf

  (
    g1867_p_spl_,
    g1867_p
  );


  buf

  (
    g1884_n_spl_,
    g1884_n
  );


  buf

  (
    g1885_n_spl_,
    g1885_n
  );


  buf

  (
    g1885_p_spl_,
    g1885_p
  );


  buf

  (
    g1866_p_spl_,
    g1866_p
  );


  buf

  (
    g1887_n_spl_,
    g1887_n
  );


  buf

  (
    g1888_p_spl_,
    g1888_p
  );


  buf

  (
    g1894_n_spl_,
    g1894_n
  );


  buf

  (
    g1895_n_spl_,
    g1895_n
  );


  buf

  (
    g1894_p_spl_,
    g1894_p
  );


  buf

  (
    g1895_p_spl_,
    g1895_p
  );


  buf

  (
    g1896_n_spl_,
    g1896_n
  );


  buf

  (
    g1896_p_spl_,
    g1896_p
  );


  buf

  (
    g1893_n_spl_,
    g1893_n
  );


  buf

  (
    g1898_p_spl_,
    g1898_p
  );


  buf

  (
    g1893_p_spl_,
    g1893_p
  );


  buf

  (
    g1898_n_spl_,
    g1898_n
  );


  buf

  (
    g1899_n_spl_,
    g1899_n
  );


  buf

  (
    g1899_p_spl_,
    g1899_p
  );


  buf

  (
    g1892_n_spl_,
    g1892_n
  );


  buf

  (
    g1901_p_spl_,
    g1901_p
  );


  buf

  (
    g1892_p_spl_,
    g1892_p
  );


  buf

  (
    g1901_n_spl_,
    g1901_n
  );


  buf

  (
    g1902_n_spl_,
    g1902_n
  );


  buf

  (
    g1902_p_spl_,
    g1902_p
  );


  buf

  (
    g1891_p_spl_,
    g1891_p
  );


  buf

  (
    g1904_n_spl_,
    g1904_n
  );


  buf

  (
    g1905_p_spl_,
    g1905_p
  );


  buf

  (
    g1908_n_spl_,
    g1908_n
  );


  buf

  (
    g1909_n_spl_,
    g1909_n
  );


  buf

  (
    g1908_p_spl_,
    g1908_p
  );


  buf

  (
    g1909_p_spl_,
    g1909_p
  );


  buf

  (
    g1910_n_spl_,
    g1910_n
  );


  buf

  (
    g1914_n_spl_,
    g1914_n
  );


endmodule
