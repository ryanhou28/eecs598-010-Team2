
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G1884,
  G1885,
  G1886,
  G1887,
  G1888,
  G1889,
  G1890,
  G1891,
  G1892,
  G1893,
  G1894,
  G1895,
  G1896,
  G1897,
  G1898,
  G1899,
  G1900,
  G1901,
  G1902,
  G1903,
  G1904,
  G1905,
  G1906,
  G1907,
  G1908
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;
  output G1884;output G1885;output G1886;output G1887;output G1888;output G1889;output G1890;output G1891;output G1892;output G1893;output G1894;output G1895;output G1896;output G1897;output G1898;output G1899;output G1900;output G1901;output G1902;output G1903;output G1904;output G1905;output G1906;output G1907;output G1908;
  wire new_n59_;wire new_n60_;wire new_n61_;wire new_n62_;wire new_n63_;wire new_n64_;wire new_n65_;wire new_n66_;wire new_n67_;wire new_n68_;wire new_n69_;wire new_n70_;wire new_n71_;wire new_n72_;wire new_n73_;wire new_n74_;wire new_n75_;wire new_n76_;wire new_n77_;wire new_n78_;wire new_n79_;wire new_n80_;wire new_n81_;wire new_n82_;wire new_n83_;wire new_n84_;wire new_n85_;wire new_n86_;wire new_n87_;wire new_n88_;wire new_n89_;wire new_n90_;wire new_n91_;wire new_n92_;wire new_n93_;wire new_n94_;wire new_n95_;wire new_n96_;wire new_n97_;wire new_n98_;wire new_n99_;wire new_n100_;wire new_n101_;wire new_n102_;wire new_n103_;wire new_n104_;wire new_n105_;wire new_n106_;wire new_n107_;wire new_n108_;wire new_n109_;wire new_n110_;wire new_n111_;wire new_n112_;wire new_n113_;wire new_n114_;wire new_n115_;wire new_n116_;wire new_n117_;wire new_n118_;wire new_n119_;wire new_n120_;wire new_n121_;wire new_n122_;wire new_n123_;wire new_n124_;wire new_n125_;wire new_n126_;wire new_n127_;wire new_n128_;wire new_n129_;wire new_n130_;wire new_n131_;wire new_n132_;wire new_n133_;wire new_n134_;wire new_n135_;wire new_n136_;wire new_n137_;wire new_n138_;wire new_n139_;wire new_n140_;wire new_n141_;wire new_n142_;wire new_n143_;wire new_n144_;wire new_n145_;wire new_n146_;wire new_n147_;wire new_n148_;wire new_n149_;wire new_n150_;wire new_n151_;wire new_n152_;wire new_n153_;wire new_n154_;wire new_n155_;wire new_n156_;wire new_n157_;wire new_n158_;wire new_n159_;wire new_n160_;wire new_n161_;wire new_n162_;wire new_n163_;wire new_n164_;wire new_n165_;wire new_n166_;wire new_n167_;wire new_n168_;wire new_n169_;wire new_n170_;wire new_n171_;wire new_n172_;wire new_n173_;wire new_n174_;wire new_n175_;wire new_n176_;wire new_n177_;wire new_n178_;wire new_n179_;wire new_n180_;wire new_n181_;wire new_n182_;wire new_n183_;wire new_n184_;wire new_n185_;wire new_n186_;wire new_n187_;wire new_n188_;wire new_n189_;wire new_n190_;wire new_n191_;wire new_n192_;wire new_n193_;wire new_n194_;wire new_n195_;wire new_n196_;wire new_n197_;wire new_n198_;wire new_n199_;wire new_n200_;wire new_n201_;wire new_n202_;wire new_n203_;wire new_n204_;wire new_n205_;wire new_n206_;wire new_n207_;wire new_n208_;wire new_n209_;wire new_n210_;wire new_n211_;wire new_n212_;wire new_n213_;wire new_n214_;wire new_n215_;wire new_n216_;wire new_n217_;wire new_n218_;wire new_n219_;wire new_n220_;wire new_n221_;wire new_n222_;wire new_n223_;wire new_n224_;wire new_n225_;wire new_n226_;wire new_n227_;wire new_n228_;wire new_n229_;wire new_n230_;wire new_n231_;wire new_n232_;wire new_n233_;wire new_n234_;wire new_n235_;wire new_n237_;wire new_n238_;wire new_n240_;wire new_n241_;wire new_n243_;wire new_n244_;wire new_n246_;wire new_n247_;wire new_n248_;wire new_n249_;wire new_n250_;wire new_n251_;wire new_n253_;wire new_n254_;wire new_n256_;wire new_n257_;wire new_n259_;wire new_n260_;wire new_n261_;wire new_n262_;wire new_n263_;wire new_n265_;wire new_n266_;wire new_n268_;wire new_n269_;wire new_n271_;wire new_n272_;wire new_n274_;wire new_n275_;wire new_n276_;wire new_n278_;wire new_n279_;wire new_n280_;wire new_n281_;wire new_n282_;wire new_n283_;wire new_n285_;wire new_n286_;wire new_n288_;wire new_n289_;wire new_n291_;wire new_n292_;wire new_n294_;wire new_n295_;wire new_n296_;wire new_n297_;wire new_n298_;wire new_n299_;wire new_n300_;wire new_n302_;wire new_n303_;wire new_n304_;wire new_n305_;wire new_n306_;wire new_n308_;wire new_n309_;wire new_n310_;wire new_n311_;wire new_n312_;wire new_n314_;wire new_n315_;wire new_n316_;wire new_n318_;wire new_n319_;wire new_n320_;wire new_n322_;wire new_n323_;wire new_n324_;wire new_n326_;wire new_n327_;wire new_n328_;wire new_n329_;wire new_n330_;wire new_n331_;wire new_n332_;wire new_n333_;wire new_n335_;wire new_n336_;wire new_n337_;wire new_n338_;wire new_n339_;wire new_n340_;wire new_n341_;wire new_n342_;wire new_n343_;wire new_n344_;wire new_n345_;wire new_n347_;wire new_n348_;wire new_n349_;
  wire G29_spl_;
  wire G33_spl_;
  wire G33_spl_0;
  wire G33_spl_00;
  wire G33_spl_000;
  wire G33_spl_001;
  wire G33_spl_01;
  wire G33_spl_010;
  wire G33_spl_011;
  wire G33_spl_1;
  wire G33_spl_10;
  wire G33_spl_11;
  wire G23_spl_;
  wire G23_spl_0;
  wire G23_spl_1;
  wire G24_spl_;
  wire G24_spl_0;
  wire G24_spl_1;
  wire G31_spl_;
  wire G31_spl_0;
  wire G31_spl_00;
  wire G31_spl_000;
  wire G31_spl_001;
  wire G31_spl_01;
  wire G31_spl_010;
  wire G31_spl_011;
  wire G31_spl_1;
  wire G31_spl_10;
  wire G31_spl_100;
  wire G31_spl_101;
  wire G31_spl_11;
  wire G31_spl_110;
  wire new_n60__spl_;
  wire new_n59__spl_;
  wire new_n61__spl_;
  wire G32_spl_;
  wire new_n63__spl_;
  wire new_n63__spl_0;
  wire new_n63__spl_00;
  wire new_n63__spl_01;
  wire new_n63__spl_1;
  wire new_n63__spl_10;
  wire new_n64__spl_;
  wire G20_spl_;
  wire new_n66__spl_;
  wire G22_spl_;
  wire G4_spl_;
  wire G4_spl_0;
  wire G4_spl_00;
  wire G4_spl_01;
  wire G4_spl_1;
  wire G4_spl_10;
  wire G4_spl_11;
  wire G14_spl_;
  wire G14_spl_0;
  wire G14_spl_00;
  wire G14_spl_01;
  wire G14_spl_1;
  wire new_n68__spl_;
  wire new_n71__spl_;
  wire G12_spl_;
  wire G12_spl_0;
  wire G12_spl_00;
  wire G12_spl_01;
  wire G12_spl_1;
  wire G13_spl_;
  wire G13_spl_0;
  wire G13_spl_00;
  wire G13_spl_01;
  wire G13_spl_1;
  wire G11_spl_;
  wire G11_spl_0;
  wire G11_spl_00;
  wire G11_spl_01;
  wire G11_spl_1;
  wire new_n77__spl_;
  wire G15_spl_;
  wire G15_spl_0;
  wire G15_spl_00;
  wire G15_spl_01;
  wire G15_spl_1;
  wire G10_spl_;
  wire G10_spl_0;
  wire G10_spl_00;
  wire G10_spl_01;
  wire G10_spl_1;
  wire new_n83__spl_;
  wire new_n83__spl_0;
  wire new_n83__spl_1;
  wire G16_spl_;
  wire G16_spl_0;
  wire G16_spl_00;
  wire G16_spl_01;
  wire G16_spl_1;
  wire new_n80__spl_;
  wire new_n86__spl_;
  wire new_n86__spl_0;
  wire new_n86__spl_1;
  wire G2_spl_;
  wire G2_spl_0;
  wire G2_spl_00;
  wire G2_spl_01;
  wire G2_spl_1;
  wire G3_spl_;
  wire G3_spl_0;
  wire G3_spl_00;
  wire G3_spl_01;
  wire G3_spl_1;
  wire G1_spl_;
  wire G1_spl_0;
  wire G1_spl_00;
  wire G1_spl_01;
  wire G1_spl_1;
  wire new_n92__spl_;
  wire new_n89__spl_;
  wire new_n89__spl_0;
  wire new_n89__spl_00;
  wire new_n89__spl_01;
  wire new_n89__spl_1;
  wire new_n95__spl_;
  wire new_n95__spl_0;
  wire new_n95__spl_1;
  wire new_n74__spl_;
  wire new_n98__spl_;
  wire new_n101__spl_;
  wire new_n101__spl_0;
  wire G25_spl_;
  wire G25_spl_0;
  wire new_n102__spl_;
  wire new_n67__spl_;
  wire new_n67__spl_0;
  wire new_n105__spl_;
  wire new_n105__spl_0;
  wire G18_spl_;
  wire new_n108__spl_;
  wire new_n111__spl_;
  wire G9_spl_;
  wire G9_spl_0;
  wire G9_spl_00;
  wire G9_spl_01;
  wire G9_spl_1;
  wire new_n117__spl_;
  wire new_n117__spl_0;
  wire new_n117__spl_1;
  wire new_n114__spl_;
  wire new_n120__spl_;
  wire new_n120__spl_0;
  wire new_n120__spl_1;
  wire G5_spl_;
  wire G5_spl_0;
  wire G5_spl_00;
  wire G5_spl_01;
  wire G5_spl_1;
  wire G8_spl_;
  wire G8_spl_0;
  wire G8_spl_00;
  wire G8_spl_01;
  wire G8_spl_1;
  wire G8_spl_10;
  wire G8_spl_11;
  wire new_n126__spl_;
  wire new_n123__spl_;
  wire new_n129__spl_;
  wire new_n132__spl_;
  wire G27_spl_;
  wire G27_spl_0;
  wire new_n133__spl_;
  wire G6_spl_;
  wire G6_spl_0;
  wire G6_spl_00;
  wire G6_spl_01;
  wire G6_spl_1;
  wire new_n137__spl_;
  wire new_n140__spl_;
  wire new_n143__spl_;
  wire G19_spl_;
  wire new_n146__spl_;
  wire new_n148__spl_;
  wire new_n151__spl_;
  wire new_n152__spl_;
  wire G28_spl_;
  wire G28_spl_0;
  wire G7_spl_;
  wire G7_spl_0;
  wire G7_spl_00;
  wire G7_spl_01;
  wire G7_spl_1;
  wire new_n158__spl_;
  wire new_n161__spl_;
  wire new_n166__spl_;
  wire new_n164__spl_;
  wire new_n169__spl_;
  wire new_n172__spl_;
  wire new_n174__spl_;
  wire new_n174__spl_0;
  wire new_n173__spl_;
  wire G17_spl_;
  wire new_n181__spl_;
  wire new_n187__spl_;
  wire new_n190__spl_;
  wire new_n190__spl_0;
  wire new_n190__spl_1;
  wire new_n184__spl_;
  wire new_n193__spl_;
  wire new_n196__spl_;
  wire G26_spl_;
  wire G26_spl_0;
  wire new_n197__spl_;
  wire new_n204__spl_;
  wire G21_spl_;
  wire new_n206__spl_;
  wire new_n209__spl_;
  wire new_n215__spl_;
  wire new_n218__spl_;
  wire new_n212__spl_;
  wire new_n221__spl_;
  wire new_n221__spl_0;
  wire new_n224__spl_;
  wire new_n224__spl_0;
  wire new_n225__spl_;
  wire new_n226__spl_;
  wire new_n226__spl_0;
  wire new_n229__spl_;
  wire new_n229__spl_0;
  wire new_n205__spl_;
  wire new_n205__spl_0;
  wire new_n203__spl_;
  wire new_n203__spl_0;
  wire new_n231__spl_;
  wire new_n106__spl_;
  wire new_n65__spl_;
  wire new_n232__spl_;
  wire new_n233__spl_;
  wire new_n233__spl_0;
  wire new_n233__spl_00;
  wire new_n233__spl_000;
  wire new_n233__spl_001;
  wire new_n233__spl_01;
  wire new_n233__spl_010;
  wire new_n233__spl_1;
  wire new_n233__spl_10;
  wire new_n233__spl_11;
  wire G30_spl_;
  wire new_n246__spl_;
  wire new_n248__spl_;
  wire new_n248__spl_0;
  wire new_n249__spl_;
  wire new_n249__spl_0;
  wire new_n249__spl_00;
  wire new_n249__spl_000;
  wire new_n249__spl_01;
  wire new_n249__spl_1;
  wire new_n249__spl_10;
  wire new_n249__spl_11;
  wire new_n260__spl_;
  wire new_n261__spl_;
  wire new_n261__spl_0;
  wire new_n261__spl_00;
  wire new_n261__spl_01;
  wire new_n261__spl_1;
  wire new_n261__spl_10;
  wire new_n261__spl_11;
  wire new_n274__spl_;
  wire new_n281__spl_;
  wire new_n281__spl_0;
  wire new_n281__spl_00;
  wire new_n281__spl_01;
  wire new_n281__spl_1;
  wire new_n281__spl_10;
  wire new_n281__spl_11;
  wire new_n294__spl_;
  wire new_n294__spl_0;
  wire new_n294__spl_00;
  wire new_n294__spl_01;
  wire new_n294__spl_1;
  wire new_n294__spl_10;
  wire new_n303__spl_;
  wire new_n309__spl_;
  wire new_n328__spl_;
  wire new_n327__spl_;
  wire new_n331__spl_;
  wire new_n340__spl_;
  wire new_n336__spl_;
  wire new_n343__spl_;

  nor1
  g000
  (
    .dina(G29_spl_),
    .dinb(G33_spl_000),
    .dout(new_n59_)
  );


  anb2
  g001
  (
    .dina(G23_spl_0),
    .dinb(G24_spl_0),
    .dout(new_n60_)
  );


  anb2
  g002
  (
    .dina(G31_spl_000),
    .dinb(new_n60__spl_),
    .dout(new_n61_)
  );


  nab2
  g003
  (
    .dina(new_n59__spl_),
    .dinb(new_n61__spl_),
    .dout(new_n62_)
  );


  and2
  g004
  (
    .dina(G32_spl_),
    .dinb(G33_spl_000),
    .dout(new_n63_)
  );


  anb1
  g005
  (
    .dina(new_n60__spl_),
    .dinb(new_n63__spl_00),
    .dout(new_n64_)
  );


  anb1
  g006
  (
    .dina(new_n62_),
    .dinb(new_n64__spl_),
    .dout(new_n65_)
  );


  nor1
  g007
  (
    .dina(G23_spl_0),
    .dinb(G31_spl_000),
    .dout(new_n66_)
  );


  anb1
  g008
  (
    .dina(G20_spl_),
    .dinb(new_n66__spl_),
    .dout(new_n67_)
  );


  anb2
  g009
  (
    .dina(G33_spl_001),
    .dinb(G22_spl_),
    .dout(new_n68_)
  );


  nor1
  g010
  (
    .dina(G4_spl_00),
    .dinb(G14_spl_00),
    .dout(new_n69_)
  );


  nor2
  g011
  (
    .dina(G4_spl_00),
    .dinb(G14_spl_00),
    .dout(new_n70_)
  );


  anb2
  g012
  (
    .dina(new_n69_),
    .dinb(new_n70_),
    .dout(new_n71_)
  );


  anb2
  g013
  (
    .dina(new_n68__spl_),
    .dinb(new_n71__spl_),
    .dout(new_n72_)
  );


  anb1
  g014
  (
    .dina(new_n68__spl_),
    .dinb(new_n71__spl_),
    .dout(new_n73_)
  );


  anb1
  g015
  (
    .dina(new_n72_),
    .dinb(new_n73_),
    .dout(new_n74_)
  );


  and2
  g016
  (
    .dina(G12_spl_00),
    .dinb(G13_spl_00),
    .dout(new_n75_)
  );


  and1
  g017
  (
    .dina(G12_spl_00),
    .dinb(G13_spl_00),
    .dout(new_n76_)
  );


  anb1
  g018
  (
    .dina(new_n75_),
    .dinb(new_n76_),
    .dout(new_n77_)
  );


  anb1
  g019
  (
    .dina(G11_spl_00),
    .dinb(new_n77__spl_),
    .dout(new_n78_)
  );


  anb2
  g020
  (
    .dina(G11_spl_00),
    .dinb(new_n77__spl_),
    .dout(new_n79_)
  );


  anb2
  g021
  (
    .dina(new_n78_),
    .dinb(new_n79_),
    .dout(new_n80_)
  );


  anb2
  g022
  (
    .dina(G15_spl_00),
    .dinb(G10_spl_00),
    .dout(new_n81_)
  );


  anb1
  g023
  (
    .dina(G15_spl_00),
    .dinb(G10_spl_00),
    .dout(new_n82_)
  );


  anb1
  g024
  (
    .dina(new_n81_),
    .dinb(new_n82_),
    .dout(new_n83_)
  );


  anb2
  g025
  (
    .dina(new_n83__spl_0),
    .dinb(G16_spl_00),
    .dout(new_n84_)
  );


  anb1
  g026
  (
    .dina(new_n83__spl_0),
    .dinb(G16_spl_00),
    .dout(new_n85_)
  );


  anb1
  g027
  (
    .dina(new_n84_),
    .dinb(new_n85_),
    .dout(new_n86_)
  );


  anb1
  g028
  (
    .dina(new_n80__spl_),
    .dinb(new_n86__spl_0),
    .dout(new_n87_)
  );


  anb2
  g029
  (
    .dina(new_n80__spl_),
    .dinb(new_n86__spl_0),
    .dout(new_n88_)
  );


  anb2
  g030
  (
    .dina(new_n87_),
    .dinb(new_n88_),
    .dout(new_n89_)
  );


  and2
  g031
  (
    .dina(G2_spl_00),
    .dinb(G3_spl_00),
    .dout(new_n90_)
  );


  and1
  g032
  (
    .dina(G2_spl_00),
    .dinb(G3_spl_00),
    .dout(new_n91_)
  );


  anb1
  g033
  (
    .dina(new_n90_),
    .dinb(new_n91_),
    .dout(new_n92_)
  );


  anb1
  g034
  (
    .dina(G1_spl_00),
    .dinb(new_n92__spl_),
    .dout(new_n93_)
  );


  anb2
  g035
  (
    .dina(G1_spl_00),
    .dinb(new_n92__spl_),
    .dout(new_n94_)
  );


  anb2
  g036
  (
    .dina(new_n93_),
    .dinb(new_n94_),
    .dout(new_n95_)
  );


  anb2
  g037
  (
    .dina(new_n89__spl_00),
    .dinb(new_n95__spl_0),
    .dout(new_n96_)
  );


  anb1
  g038
  (
    .dina(new_n89__spl_00),
    .dinb(new_n95__spl_0),
    .dout(new_n97_)
  );


  anb1
  g039
  (
    .dina(new_n96_),
    .dinb(new_n97_),
    .dout(new_n98_)
  );


  anb2
  g040
  (
    .dina(new_n74__spl_),
    .dinb(new_n98__spl_),
    .dout(new_n99_)
  );


  anb1
  g041
  (
    .dina(new_n74__spl_),
    .dinb(new_n98__spl_),
    .dout(new_n100_)
  );


  anb1
  g042
  (
    .dina(new_n99_),
    .dinb(new_n100_),
    .dout(new_n101_)
  );


  nor1
  g043
  (
    .dina(G31_spl_001),
    .dinb(new_n101__spl_0),
    .dout(new_n102_)
  );


  anb2
  g044
  (
    .dina(G25_spl_0),
    .dinb(new_n102__spl_),
    .dout(new_n103_)
  );


  anb1
  g045
  (
    .dina(G25_spl_0),
    .dinb(new_n102__spl_),
    .dout(new_n104_)
  );


  anb1
  g046
  (
    .dina(new_n103_),
    .dinb(new_n104_),
    .dout(new_n105_)
  );


  anb1
  g047
  (
    .dina(new_n67__spl_0),
    .dinb(new_n105__spl_0),
    .dout(new_n106_)
  );


  anb1
  g048
  (
    .dina(G18_spl_),
    .dinb(G24_spl_0),
    .dout(new_n107_)
  );


  anb1
  g049
  (
    .dina(new_n107_),
    .dinb(G33_spl_001),
    .dout(new_n108_)
  );


  anb1
  g050
  (
    .dina(G15_spl_01),
    .dinb(new_n108__spl_),
    .dout(new_n109_)
  );


  anb2
  g051
  (
    .dina(G15_spl_01),
    .dinb(new_n108__spl_),
    .dout(new_n110_)
  );


  anb2
  g052
  (
    .dina(new_n109_),
    .dinb(new_n110_),
    .dout(new_n111_)
  );


  anb2
  g053
  (
    .dina(G11_spl_01),
    .dinb(new_n111__spl_),
    .dout(new_n112_)
  );


  anb1
  g054
  (
    .dina(G11_spl_01),
    .dinb(new_n111__spl_),
    .dout(new_n113_)
  );


  anb1
  g055
  (
    .dina(new_n112_),
    .dinb(new_n113_),
    .dout(new_n114_)
  );


  and2
  g056
  (
    .dina(G9_spl_00),
    .dinb(G14_spl_01),
    .dout(new_n115_)
  );


  and1
  g057
  (
    .dina(G9_spl_00),
    .dinb(G14_spl_01),
    .dout(new_n116_)
  );


  anb1
  g058
  (
    .dina(new_n115_),
    .dinb(new_n116_),
    .dout(new_n117_)
  );


  anb2
  g059
  (
    .dina(new_n117__spl_0),
    .dinb(G16_spl_01),
    .dout(new_n118_)
  );


  anb1
  g060
  (
    .dina(new_n117__spl_0),
    .dinb(G16_spl_01),
    .dout(new_n119_)
  );


  anb1
  g061
  (
    .dina(new_n118_),
    .dinb(new_n119_),
    .dout(new_n120_)
  );


  anb1
  g062
  (
    .dina(new_n114__spl_),
    .dinb(new_n120__spl_0),
    .dout(new_n121_)
  );


  anb2
  g063
  (
    .dina(new_n114__spl_),
    .dinb(new_n120__spl_0),
    .dout(new_n122_)
  );


  anb2
  g064
  (
    .dina(new_n121_),
    .dinb(new_n122_),
    .dout(new_n123_)
  );


  anb1
  g065
  (
    .dina(G5_spl_00),
    .dinb(G8_spl_00),
    .dout(new_n124_)
  );


  anb2
  g066
  (
    .dina(G5_spl_00),
    .dinb(G8_spl_00),
    .dout(new_n125_)
  );


  anb2
  g067
  (
    .dina(new_n124_),
    .dinb(new_n125_),
    .dout(new_n126_)
  );


  nab1
  g068
  (
    .dina(G2_spl_01),
    .dinb(new_n126__spl_),
    .dout(new_n127_)
  );


  nab2
  g069
  (
    .dina(G2_spl_01),
    .dinb(new_n126__spl_),
    .dout(new_n128_)
  );


  anb2
  g070
  (
    .dina(new_n127_),
    .dinb(new_n128_),
    .dout(new_n129_)
  );


  anb1
  g071
  (
    .dina(new_n123__spl_),
    .dinb(new_n129__spl_),
    .dout(new_n130_)
  );


  anb2
  g072
  (
    .dina(new_n123__spl_),
    .dinb(new_n129__spl_),
    .dout(new_n131_)
  );


  anb2
  g073
  (
    .dina(new_n130_),
    .dinb(new_n131_),
    .dout(new_n132_)
  );


  nab1
  g074
  (
    .dina(G31_spl_001),
    .dinb(new_n132__spl_),
    .dout(new_n133_)
  );


  anb2
  g075
  (
    .dina(G27_spl_0),
    .dinb(new_n133__spl_),
    .dout(new_n134_)
  );


  anb1
  g076
  (
    .dina(G6_spl_00),
    .dinb(G8_spl_01),
    .dout(new_n135_)
  );


  anb2
  g077
  (
    .dina(G6_spl_00),
    .dinb(G8_spl_01),
    .dout(new_n136_)
  );


  anb2
  g078
  (
    .dina(new_n135_),
    .dinb(new_n136_),
    .dout(new_n137_)
  );


  nab1
  g079
  (
    .dina(G3_spl_01),
    .dinb(new_n137__spl_),
    .dout(new_n138_)
  );


  nab2
  g080
  (
    .dina(G3_spl_01),
    .dinb(new_n137__spl_),
    .dout(new_n139_)
  );


  anb2
  g081
  (
    .dina(new_n138_),
    .dinb(new_n139_),
    .dout(new_n140_)
  );


  nor1
  g082
  (
    .dina(G12_spl_01),
    .dinb(new_n83__spl_1),
    .dout(new_n141_)
  );


  nor2
  g083
  (
    .dina(G12_spl_01),
    .dinb(new_n83__spl_1),
    .dout(new_n142_)
  );


  anb2
  g084
  (
    .dina(new_n141_),
    .dinb(new_n142_),
    .dout(new_n143_)
  );


  anb1
  g085
  (
    .dina(new_n140__spl_),
    .dinb(new_n143__spl_),
    .dout(new_n144_)
  );


  anb2
  g086
  (
    .dina(new_n140__spl_),
    .dinb(new_n143__spl_),
    .dout(new_n145_)
  );


  anb2
  g087
  (
    .dina(new_n144_),
    .dinb(new_n145_),
    .dout(new_n146_)
  );


  anb1
  g088
  (
    .dina(G19_spl_),
    .dinb(G23_spl_1),
    .dout(new_n147_)
  );


  anb1
  g089
  (
    .dina(new_n147_),
    .dinb(G33_spl_010),
    .dout(new_n148_)
  );


  anb1
  g090
  (
    .dina(new_n146__spl_),
    .dinb(new_n148__spl_),
    .dout(new_n149_)
  );


  anb2
  g091
  (
    .dina(new_n146__spl_),
    .dinb(new_n148__spl_),
    .dout(new_n150_)
  );


  anb2
  g092
  (
    .dina(new_n149_),
    .dinb(new_n150_),
    .dout(new_n151_)
  );


  nab1
  g093
  (
    .dina(G31_spl_010),
    .dinb(new_n151__spl_),
    .dout(new_n152_)
  );


  anb1
  g094
  (
    .dina(new_n152__spl_),
    .dinb(G28_spl_0),
    .dout(new_n153_)
  );


  anb2
  g095
  (
    .dina(new_n152__spl_),
    .dinb(G28_spl_0),
    .dout(new_n154_)
  );


  anb2
  g096
  (
    .dina(new_n153_),
    .dinb(new_n154_),
    .dout(new_n155_)
  );


  anb1
  g097
  (
    .dina(G7_spl_00),
    .dinb(G10_spl_01),
    .dout(new_n156_)
  );


  anb2
  g098
  (
    .dina(G7_spl_00),
    .dinb(G10_spl_01),
    .dout(new_n157_)
  );


  anb2
  g099
  (
    .dina(new_n156_),
    .dinb(new_n157_),
    .dout(new_n158_)
  );


  anb2
  g100
  (
    .dina(G4_spl_01),
    .dinb(new_n158__spl_),
    .dout(new_n159_)
  );


  anb1
  g101
  (
    .dina(G4_spl_01),
    .dinb(new_n158__spl_),
    .dout(new_n160_)
  );


  anb1
  g102
  (
    .dina(new_n159_),
    .dinb(new_n160_),
    .dout(new_n161_)
  );


  anb1
  g103
  (
    .dina(new_n120__spl_1),
    .dinb(new_n161__spl_),
    .dout(new_n162_)
  );


  anb2
  g104
  (
    .dina(new_n120__spl_1),
    .dinb(new_n161__spl_),
    .dout(new_n163_)
  );


  anb2
  g105
  (
    .dina(new_n162_),
    .dinb(new_n163_),
    .dout(new_n164_)
  );


  anb1
  g106
  (
    .dina(G20_spl_),
    .dinb(G23_spl_1),
    .dout(new_n165_)
  );


  anb1
  g107
  (
    .dina(new_n165_),
    .dinb(G33_spl_010),
    .dout(new_n166_)
  );


  anb2
  g108
  (
    .dina(G13_spl_01),
    .dinb(new_n166__spl_),
    .dout(new_n167_)
  );


  anb1
  g109
  (
    .dina(G13_spl_01),
    .dinb(new_n166__spl_),
    .dout(new_n168_)
  );


  anb1
  g110
  (
    .dina(new_n167_),
    .dinb(new_n168_),
    .dout(new_n169_)
  );


  anb1
  g111
  (
    .dina(new_n164__spl_),
    .dinb(new_n169__spl_),
    .dout(new_n170_)
  );


  anb2
  g112
  (
    .dina(new_n164__spl_),
    .dinb(new_n169__spl_),
    .dout(new_n171_)
  );


  anb2
  g113
  (
    .dina(new_n170_),
    .dinb(new_n171_),
    .dout(new_n172_)
  );


  nab1
  g114
  (
    .dina(G31_spl_010),
    .dinb(new_n172__spl_),
    .dout(new_n173_)
  );


  anb1
  g115
  (
    .dina(G19_spl_),
    .dinb(new_n66__spl_),
    .dout(new_n174_)
  );


  anb2
  g116
  (
    .dina(new_n174__spl_0),
    .dinb(new_n173__spl_),
    .dout(new_n175_)
  );


  anb1
  g117
  (
    .dina(new_n174__spl_0),
    .dinb(new_n173__spl_),
    .dout(new_n176_)
  );


  anb1
  g118
  (
    .dina(new_n175_),
    .dinb(new_n176_),
    .dout(new_n177_)
  );


  anb2
  g119
  (
    .dina(new_n155_),
    .dinb(new_n177_),
    .dout(new_n178_)
  );


  anb1
  g120
  (
    .dina(new_n134_),
    .dinb(new_n178_),
    .dout(new_n179_)
  );


  anb1
  g121
  (
    .dina(G17_spl_),
    .dinb(G24_spl_1),
    .dout(new_n180_)
  );


  anb2
  g122
  (
    .dina(G33_spl_011),
    .dinb(new_n180_),
    .dout(new_n181_)
  );


  nab2
  g123
  (
    .dina(G1_spl_01),
    .dinb(new_n181__spl_),
    .dout(new_n182_)
  );


  nab1
  g124
  (
    .dina(G1_spl_01),
    .dinb(new_n181__spl_),
    .dout(new_n183_)
  );


  anb1
  g125
  (
    .dina(new_n182_),
    .dinb(new_n183_),
    .dout(new_n184_)
  );


  and2
  g126
  (
    .dina(G6_spl_01),
    .dinb(G7_spl_01),
    .dout(new_n185_)
  );


  and1
  g127
  (
    .dina(G6_spl_01),
    .dinb(G7_spl_01),
    .dout(new_n186_)
  );


  anb1
  g128
  (
    .dina(new_n185_),
    .dinb(new_n186_),
    .dout(new_n187_)
  );


  anb1
  g129
  (
    .dina(G5_spl_01),
    .dinb(new_n187__spl_),
    .dout(new_n188_)
  );


  anb2
  g130
  (
    .dina(G5_spl_01),
    .dinb(new_n187__spl_),
    .dout(new_n189_)
  );


  anb2
  g131
  (
    .dina(new_n188_),
    .dinb(new_n189_),
    .dout(new_n190_)
  );


  anb2
  g132
  (
    .dina(new_n89__spl_01),
    .dinb(new_n190__spl_0),
    .dout(new_n191_)
  );


  anb1
  g133
  (
    .dina(new_n89__spl_01),
    .dinb(new_n190__spl_0),
    .dout(new_n192_)
  );


  anb1
  g134
  (
    .dina(new_n191_),
    .dinb(new_n192_),
    .dout(new_n193_)
  );


  anb1
  g135
  (
    .dina(new_n184__spl_),
    .dinb(new_n193__spl_),
    .dout(new_n194_)
  );


  anb2
  g136
  (
    .dina(new_n184__spl_),
    .dinb(new_n193__spl_),
    .dout(new_n195_)
  );


  anb2
  g137
  (
    .dina(new_n194_),
    .dinb(new_n195_),
    .dout(new_n196_)
  );


  nab1
  g138
  (
    .dina(G31_spl_011),
    .dinb(new_n196__spl_),
    .dout(new_n197_)
  );


  anb1
  g139
  (
    .dina(G26_spl_0),
    .dinb(new_n197__spl_),
    .dout(new_n198_)
  );


  anb2
  g140
  (
    .dina(G26_spl_0),
    .dinb(new_n197__spl_),
    .dout(new_n199_)
  );


  anb1
  g141
  (
    .dina(G27_spl_0),
    .dinb(new_n133__spl_),
    .dout(new_n200_)
  );


  anb1
  g142
  (
    .dina(new_n199_),
    .dinb(new_n200_),
    .dout(new_n201_)
  );


  anb2
  g143
  (
    .dina(new_n198_),
    .dinb(new_n201_),
    .dout(new_n202_)
  );


  anb1
  g144
  (
    .dina(new_n179_),
    .dinb(new_n202_),
    .dout(new_n203_)
  );


  nor1
  g145
  (
    .dina(G24_spl_1),
    .dinb(G31_spl_011),
    .dout(new_n204_)
  );


  anb2
  g146
  (
    .dina(new_n204__spl_),
    .dinb(G18_spl_),
    .dout(new_n205_)
  );


  anb2
  g147
  (
    .dina(G33_spl_011),
    .dinb(G21_spl_),
    .dout(new_n206_)
  );


  anb1
  g148
  (
    .dina(G9_spl_01),
    .dinb(new_n86__spl_1),
    .dout(new_n207_)
  );


  anb2
  g149
  (
    .dina(G9_spl_01),
    .dinb(new_n86__spl_1),
    .dout(new_n208_)
  );


  anb2
  g150
  (
    .dina(new_n207_),
    .dinb(new_n208_),
    .dout(new_n209_)
  );


  anb2
  g151
  (
    .dina(new_n206__spl_),
    .dinb(new_n209__spl_),
    .dout(new_n210_)
  );


  anb1
  g152
  (
    .dina(new_n206__spl_),
    .dinb(new_n209__spl_),
    .dout(new_n211_)
  );


  anb1
  g153
  (
    .dina(new_n210_),
    .dinb(new_n211_),
    .dout(new_n212_)
  );


  and1
  g154
  (
    .dina(new_n95__spl_1),
    .dinb(new_n190__spl_1),
    .dout(new_n213_)
  );


  and2
  g155
  (
    .dina(new_n95__spl_1),
    .dinb(new_n190__spl_1),
    .dout(new_n214_)
  );


  nab1
  g156
  (
    .dina(new_n213_),
    .dinb(new_n214_),
    .dout(new_n215_)
  );


  anb2
  g157
  (
    .dina(G8_spl_10),
    .dinb(G4_spl_10),
    .dout(new_n216_)
  );


  anb1
  g158
  (
    .dina(G8_spl_10),
    .dinb(G4_spl_10),
    .dout(new_n217_)
  );


  anb1
  g159
  (
    .dina(new_n216_),
    .dinb(new_n217_),
    .dout(new_n218_)
  );


  anb2
  g160
  (
    .dina(new_n215__spl_),
    .dinb(new_n218__spl_),
    .dout(new_n219_)
  );


  anb1
  g161
  (
    .dina(new_n215__spl_),
    .dinb(new_n218__spl_),
    .dout(new_n220_)
  );


  anb1
  g162
  (
    .dina(new_n219_),
    .dinb(new_n220_),
    .dout(new_n221_)
  );


  anb1
  g163
  (
    .dina(new_n212__spl_),
    .dinb(new_n221__spl_0),
    .dout(new_n222_)
  );


  anb2
  g164
  (
    .dina(new_n212__spl_),
    .dinb(new_n221__spl_0),
    .dout(new_n223_)
  );


  anb2
  g165
  (
    .dina(new_n222_),
    .dinb(new_n223_),
    .dout(new_n224_)
  );


  nor1
  g166
  (
    .dina(G31_spl_100),
    .dinb(new_n224__spl_0),
    .dout(new_n225_)
  );


  anb1
  g167
  (
    .dina(G17_spl_),
    .dinb(new_n204__spl_),
    .dout(new_n226_)
  );


  anb1
  g168
  (
    .dina(new_n225__spl_),
    .dinb(new_n226__spl_0),
    .dout(new_n227_)
  );


  anb2
  g169
  (
    .dina(new_n225__spl_),
    .dinb(new_n226__spl_0),
    .dout(new_n228_)
  );


  anb2
  g170
  (
    .dina(new_n227_),
    .dinb(new_n228_),
    .dout(new_n229_)
  );


  anb1
  g171
  (
    .dina(new_n229__spl_0),
    .dinb(new_n205__spl_0),
    .dout(new_n230_)
  );


  anb1
  g172
  (
    .dina(new_n203__spl_0),
    .dinb(new_n230_),
    .dout(new_n231_)
  );


  anb1
  g173
  (
    .dina(new_n231__spl_),
    .dinb(new_n106__spl_),
    .dout(new_n232_)
  );


  anb2
  g174
  (
    .dina(new_n65__spl_),
    .dinb(new_n232__spl_),
    .dout(new_n233_)
  );


  nab1
  g175
  (
    .dina(G1_spl_1),
    .dinb(new_n233__spl_000),
    .dout(new_n234_)
  );


  nab2
  g176
  (
    .dina(G1_spl_1),
    .dinb(new_n233__spl_000),
    .dout(new_n235_)
  );


  anb2
  g177
  (
    .dina(new_n234_),
    .dinb(new_n235_),
    .dout(G1884)
  );


  nab1
  g178
  (
    .dina(G2_spl_1),
    .dinb(new_n233__spl_001),
    .dout(new_n237_)
  );


  nab2
  g179
  (
    .dina(G2_spl_1),
    .dinb(new_n233__spl_001),
    .dout(new_n238_)
  );


  anb2
  g180
  (
    .dina(new_n237_),
    .dinb(new_n238_),
    .dout(G1885)
  );


  nab1
  g181
  (
    .dina(G3_spl_1),
    .dinb(new_n233__spl_010),
    .dout(new_n240_)
  );


  nab2
  g182
  (
    .dina(G3_spl_1),
    .dinb(new_n233__spl_010),
    .dout(new_n241_)
  );


  anb2
  g183
  (
    .dina(new_n240_),
    .dinb(new_n241_),
    .dout(G1886)
  );


  nab1
  g184
  (
    .dina(G4_spl_11),
    .dinb(new_n233__spl_01),
    .dout(new_n243_)
  );


  nab2
  g185
  (
    .dina(G4_spl_11),
    .dinb(new_n233__spl_10),
    .dout(new_n244_)
  );


  anb2
  g186
  (
    .dina(new_n243_),
    .dinb(new_n244_),
    .dout(G1887)
  );


  nor1
  g187
  (
    .dina(G30_spl_),
    .dinb(G33_spl_10),
    .dout(new_n246_)
  );


  anb2
  g188
  (
    .dina(new_n61__spl_),
    .dinb(new_n246__spl_),
    .dout(new_n247_)
  );


  anb2
  g189
  (
    .dina(new_n64__spl_),
    .dinb(new_n247_),
    .dout(new_n248_)
  );


  nor2
  g190
  (
    .dina(new_n232__spl_),
    .dinb(new_n248__spl_0),
    .dout(new_n249_)
  );


  nab1
  g191
  (
    .dina(G10_spl_1),
    .dinb(new_n249__spl_000),
    .dout(new_n250_)
  );


  nab2
  g192
  (
    .dina(G10_spl_1),
    .dinb(new_n249__spl_000),
    .dout(new_n251_)
  );


  anb2
  g193
  (
    .dina(new_n250_),
    .dinb(new_n251_),
    .dout(G1888)
  );


  nab1
  g194
  (
    .dina(G15_spl_1),
    .dinb(new_n249__spl_00),
    .dout(new_n253_)
  );


  nab2
  g195
  (
    .dina(G15_spl_1),
    .dinb(new_n249__spl_01),
    .dout(new_n254_)
  );


  anb2
  g196
  (
    .dina(new_n253_),
    .dinb(new_n254_),
    .dout(G1889)
  );


  nab1
  g197
  (
    .dina(G16_spl_1),
    .dinb(new_n249__spl_01),
    .dout(new_n256_)
  );


  nab2
  g198
  (
    .dina(G16_spl_1),
    .dinb(new_n249__spl_10),
    .dout(new_n257_)
  );


  anb2
  g199
  (
    .dina(new_n256_),
    .dinb(new_n257_),
    .dout(G1890)
  );


  nor2
  g200
  (
    .dina(new_n67__spl_0),
    .dinb(new_n105__spl_0),
    .dout(new_n259_)
  );


  anb1
  g201
  (
    .dina(new_n231__spl_),
    .dinb(new_n259_),
    .dout(new_n260_)
  );


  anb2
  g202
  (
    .dina(new_n65__spl_),
    .dinb(new_n260__spl_),
    .dout(new_n261_)
  );


  nab1
  g203
  (
    .dina(G5_spl_1),
    .dinb(new_n261__spl_00),
    .dout(new_n262_)
  );


  nab2
  g204
  (
    .dina(G5_spl_1),
    .dinb(new_n261__spl_00),
    .dout(new_n263_)
  );


  anb2
  g205
  (
    .dina(new_n262_),
    .dinb(new_n263_),
    .dout(G1891)
  );


  nab1
  g206
  (
    .dina(G6_spl_1),
    .dinb(new_n261__spl_01),
    .dout(new_n265_)
  );


  nab2
  g207
  (
    .dina(G6_spl_1),
    .dinb(new_n261__spl_01),
    .dout(new_n266_)
  );


  anb2
  g208
  (
    .dina(new_n265_),
    .dinb(new_n266_),
    .dout(G1892)
  );


  nab1
  g209
  (
    .dina(G7_spl_1),
    .dinb(new_n261__spl_10),
    .dout(new_n268_)
  );


  nab2
  g210
  (
    .dina(G7_spl_1),
    .dinb(new_n261__spl_10),
    .dout(new_n269_)
  );


  anb2
  g211
  (
    .dina(new_n268_),
    .dinb(new_n269_),
    .dout(G1893)
  );


  nab1
  g212
  (
    .dina(G8_spl_11),
    .dinb(new_n261__spl_11),
    .dout(new_n271_)
  );


  nab2
  g213
  (
    .dina(G8_spl_11),
    .dinb(new_n261__spl_11),
    .dout(new_n272_)
  );


  anb2
  g214
  (
    .dina(new_n271_),
    .dinb(new_n272_),
    .dout(G1894)
  );


  nor2
  g215
  (
    .dina(new_n248__spl_0),
    .dinb(new_n260__spl_),
    .dout(new_n274_)
  );


  anb1
  g216
  (
    .dina(G9_spl_1),
    .dinb(new_n274__spl_),
    .dout(new_n275_)
  );


  anb2
  g217
  (
    .dina(G9_spl_1),
    .dinb(new_n274__spl_),
    .dout(new_n276_)
  );


  anb2
  g218
  (
    .dina(new_n275_),
    .dinb(new_n276_),
    .dout(G1895)
  );


  anb1
  g219
  (
    .dina(new_n248__spl_),
    .dinb(new_n205__spl_0),
    .dout(new_n278_)
  );


  nab1
  g220
  (
    .dina(new_n229__spl_0),
    .dinb(new_n278_),
    .dout(new_n279_)
  );


  anb2
  g221
  (
    .dina(new_n106__spl_),
    .dinb(new_n279_),
    .dout(new_n280_)
  );


  anb1
  g222
  (
    .dina(new_n203__spl_0),
    .dinb(new_n280_),
    .dout(new_n281_)
  );


  anb2
  g223
  (
    .dina(new_n281__spl_00),
    .dinb(G11_spl_1),
    .dout(new_n282_)
  );


  anb1
  g224
  (
    .dina(new_n281__spl_00),
    .dinb(G11_spl_1),
    .dout(new_n283_)
  );


  anb1
  g225
  (
    .dina(new_n282_),
    .dinb(new_n283_),
    .dout(G1896)
  );


  anb2
  g226
  (
    .dina(new_n281__spl_01),
    .dinb(G12_spl_1),
    .dout(new_n285_)
  );


  anb1
  g227
  (
    .dina(new_n281__spl_01),
    .dinb(G12_spl_1),
    .dout(new_n286_)
  );


  anb1
  g228
  (
    .dina(new_n285_),
    .dinb(new_n286_),
    .dout(G1897)
  );


  anb2
  g229
  (
    .dina(new_n281__spl_10),
    .dinb(G13_spl_1),
    .dout(new_n288_)
  );


  anb1
  g230
  (
    .dina(new_n281__spl_10),
    .dinb(G13_spl_1),
    .dout(new_n289_)
  );


  anb1
  g231
  (
    .dina(new_n288_),
    .dinb(new_n289_),
    .dout(G1898)
  );


  anb2
  g232
  (
    .dina(new_n281__spl_11),
    .dinb(G14_spl_1),
    .dout(new_n291_)
  );


  anb1
  g233
  (
    .dina(new_n281__spl_11),
    .dinb(G14_spl_1),
    .dout(new_n292_)
  );


  anb1
  g234
  (
    .dina(new_n291_),
    .dinb(new_n292_),
    .dout(G1899)
  );


  and1
  g235
  (
    .dina(new_n233__spl_10),
    .dinb(new_n249__spl_10),
    .dout(new_n294_)
  );


  anb1
  g236
  (
    .dina(G32_spl_),
    .dinb(new_n294__spl_00),
    .dout(new_n295_)
  );


  anb2
  g237
  (
    .dina(new_n67__spl_),
    .dinb(new_n205__spl_),
    .dout(new_n296_)
  );


  anb1
  g238
  (
    .dina(new_n105__spl_),
    .dinb(new_n296_),
    .dout(new_n297_)
  );


  anb2
  g239
  (
    .dina(new_n229__spl_),
    .dinb(new_n297_),
    .dout(new_n298_)
  );


  nab2
  g240
  (
    .dina(new_n203__spl_),
    .dinb(new_n298_),
    .dout(new_n299_)
  );


  nab1
  g241
  (
    .dina(G33_spl_10),
    .dinb(new_n299_),
    .dout(new_n300_)
  );


  anb2
  g242
  (
    .dina(new_n295_),
    .dinb(new_n300_),
    .dout(G1900)
  );


  anb1
  g243
  (
    .dina(new_n226__spl_),
    .dinb(G31_spl_100),
    .dout(new_n302_)
  );


  anb2
  g244
  (
    .dina(new_n294__spl_00),
    .dinb(new_n302_),
    .dout(new_n303_)
  );


  anb2
  g245
  (
    .dina(new_n224__spl_0),
    .dinb(new_n303__spl_),
    .dout(new_n304_)
  );


  anb1
  g246
  (
    .dina(new_n224__spl_),
    .dinb(new_n303__spl_),
    .dout(new_n305_)
  );


  anb1
  g247
  (
    .dina(new_n304_),
    .dinb(new_n305_),
    .dout(new_n306_)
  );


  anb1
  g248
  (
    .dina(new_n63__spl_00),
    .dinb(new_n306_),
    .dout(G1901)
  );


  anb1
  g249
  (
    .dina(G25_spl_),
    .dinb(G31_spl_101),
    .dout(new_n308_)
  );


  anb2
  g250
  (
    .dina(new_n294__spl_01),
    .dinb(new_n308_),
    .dout(new_n309_)
  );


  anb2
  g251
  (
    .dina(new_n101__spl_0),
    .dinb(new_n309__spl_),
    .dout(new_n310_)
  );


  anb1
  g252
  (
    .dina(new_n101__spl_),
    .dinb(new_n309__spl_),
    .dout(new_n311_)
  );


  anb1
  g253
  (
    .dina(new_n310_),
    .dinb(new_n311_),
    .dout(new_n312_)
  );


  anb1
  g254
  (
    .dina(new_n63__spl_01),
    .dinb(new_n312_),
    .dout(G1902)
  );


  anb1
  g255
  (
    .dina(G27_spl_),
    .dinb(G31_spl_101),
    .dout(new_n314_)
  );


  anb1
  g256
  (
    .dina(new_n314_),
    .dinb(new_n294__spl_01),
    .dout(new_n315_)
  );


  anb1
  g257
  (
    .dina(new_n132__spl_),
    .dinb(new_n315_),
    .dout(new_n316_)
  );


  anb1
  g258
  (
    .dina(new_n63__spl_01),
    .dinb(new_n316_),
    .dout(G1903)
  );


  anb1
  g259
  (
    .dina(G28_spl_),
    .dinb(G31_spl_110),
    .dout(new_n318_)
  );


  anb1
  g260
  (
    .dina(new_n318_),
    .dinb(new_n294__spl_10),
    .dout(new_n319_)
  );


  anb1
  g261
  (
    .dina(new_n151__spl_),
    .dinb(new_n319_),
    .dout(new_n320_)
  );


  anb1
  g262
  (
    .dina(new_n63__spl_10),
    .dinb(new_n320_),
    .dout(G1904)
  );


  anb1
  g263
  (
    .dina(new_n174__spl_),
    .dinb(G31_spl_110),
    .dout(new_n322_)
  );


  anb1
  g264
  (
    .dina(new_n322_),
    .dinb(new_n294__spl_10),
    .dout(new_n323_)
  );


  anb1
  g265
  (
    .dina(new_n172__spl_),
    .dinb(new_n323_),
    .dout(new_n324_)
  );


  anb1
  g266
  (
    .dina(new_n63__spl_10),
    .dinb(new_n324_),
    .dout(G1905)
  );


  nor2
  g267
  (
    .dina(G21_spl_),
    .dinb(G29_spl_),
    .dout(new_n326_)
  );


  anb2
  g268
  (
    .dina(G33_spl_11),
    .dinb(new_n326_),
    .dout(new_n327_)
  );


  anb2
  g269
  (
    .dina(new_n59__spl_),
    .dinb(new_n221__spl_),
    .dout(new_n328_)
  );


  anb2
  g270
  (
    .dina(new_n233__spl_11),
    .dinb(new_n328__spl_),
    .dout(new_n329_)
  );


  anb1
  g271
  (
    .dina(new_n233__spl_11),
    .dinb(new_n328__spl_),
    .dout(new_n330_)
  );


  anb1
  g272
  (
    .dina(new_n329_),
    .dinb(new_n330_),
    .dout(new_n331_)
  );


  anb1
  g273
  (
    .dina(new_n327__spl_),
    .dinb(new_n331__spl_),
    .dout(new_n332_)
  );


  anb2
  g274
  (
    .dina(new_n327__spl_),
    .dinb(new_n331__spl_),
    .dout(new_n333_)
  );


  anb2
  g275
  (
    .dina(new_n332_),
    .dinb(new_n333_),
    .dout(G1906)
  );


  nor2
  g276
  (
    .dina(G22_spl_),
    .dinb(G30_spl_),
    .dout(new_n335_)
  );


  anb2
  g277
  (
    .dina(G33_spl_11),
    .dinb(new_n335_),
    .dout(new_n336_)
  );


  anb1
  g278
  (
    .dina(new_n89__spl_1),
    .dinb(new_n117__spl_1),
    .dout(new_n337_)
  );


  anb2
  g279
  (
    .dina(new_n89__spl_1),
    .dinb(new_n117__spl_1),
    .dout(new_n338_)
  );


  anb2
  g280
  (
    .dina(new_n337_),
    .dinb(new_n338_),
    .dout(new_n339_)
  );


  anb2
  g281
  (
    .dina(new_n246__spl_),
    .dinb(new_n339_),
    .dout(new_n340_)
  );


  anb2
  g282
  (
    .dina(new_n249__spl_11),
    .dinb(new_n340__spl_),
    .dout(new_n341_)
  );


  anb1
  g283
  (
    .dina(new_n249__spl_11),
    .dinb(new_n340__spl_),
    .dout(new_n342_)
  );


  anb1
  g284
  (
    .dina(new_n341_),
    .dinb(new_n342_),
    .dout(new_n343_)
  );


  anb1
  g285
  (
    .dina(new_n336__spl_),
    .dinb(new_n343__spl_),
    .dout(new_n344_)
  );


  anb2
  g286
  (
    .dina(new_n336__spl_),
    .dinb(new_n343__spl_),
    .dout(new_n345_)
  );


  anb2
  g287
  (
    .dina(new_n344_),
    .dinb(new_n345_),
    .dout(G1907)
  );


  anb1
  g288
  (
    .dina(G26_spl_),
    .dinb(G31_spl_11),
    .dout(new_n347_)
  );


  anb1
  g289
  (
    .dina(new_n347_),
    .dinb(new_n294__spl_1),
    .dout(new_n348_)
  );


  anb1
  g290
  (
    .dina(new_n196__spl_),
    .dinb(new_n348_),
    .dout(new_n349_)
  );


  and1
  g291
  (
    .dina(new_n63__spl_1),
    .dinb(new_n349_),
    .dout(G1908)
  );


  splt
  gG29
  (
    .dout(G29_spl_),
    .din(G29)
  );


  splt
  gG33
  (
    .dout(G33_spl_),
    .din(G33)
  );


  splt
  gG33_spl_
  (
    .dout(G33_spl_0),
    .din(G33_spl_)
  );


  splt
  gG33_spl_0
  (
    .dout(G33_spl_00),
    .din(G33_spl_0)
  );


  splt
  gG33_spl_00
  (
    .dout(G33_spl_000),
    .din(G33_spl_00)
  );


  splt
  gG33_spl_00
  (
    .dout(G33_spl_001),
    .din(G33_spl_00)
  );


  splt
  gG33_spl_0
  (
    .dout(G33_spl_01),
    .din(G33_spl_0)
  );


  splt
  gG33_spl_01
  (
    .dout(G33_spl_010),
    .din(G33_spl_01)
  );


  splt
  gG33_spl_01
  (
    .dout(G33_spl_011),
    .din(G33_spl_01)
  );


  splt
  gG33_spl_
  (
    .dout(G33_spl_1),
    .din(G33_spl_)
  );


  splt
  gG33_spl_1
  (
    .dout(G33_spl_10),
    .din(G33_spl_1)
  );


  splt
  gG33_spl_1
  (
    .dout(G33_spl_11),
    .din(G33_spl_1)
  );


  splt
  gG23
  (
    .dout(G23_spl_),
    .din(G23)
  );


  splt
  gG23_spl_
  (
    .dout(G23_spl_0),
    .din(G23_spl_)
  );


  splt
  gG23_spl_
  (
    .dout(G23_spl_1),
    .din(G23_spl_)
  );


  splt
  gG24
  (
    .dout(G24_spl_),
    .din(G24)
  );


  splt
  gG24_spl_
  (
    .dout(G24_spl_0),
    .din(G24_spl_)
  );


  splt
  gG24_spl_
  (
    .dout(G24_spl_1),
    .din(G24_spl_)
  );


  splt
  gG31
  (
    .dout(G31_spl_),
    .din(G31)
  );


  splt
  gG31_spl_
  (
    .dout(G31_spl_0),
    .din(G31_spl_)
  );


  splt
  gG31_spl_0
  (
    .dout(G31_spl_00),
    .din(G31_spl_0)
  );


  splt
  gG31_spl_00
  (
    .dout(G31_spl_000),
    .din(G31_spl_00)
  );


  splt
  gG31_spl_00
  (
    .dout(G31_spl_001),
    .din(G31_spl_00)
  );


  splt
  gG31_spl_0
  (
    .dout(G31_spl_01),
    .din(G31_spl_0)
  );


  splt
  gG31_spl_01
  (
    .dout(G31_spl_010),
    .din(G31_spl_01)
  );


  splt
  gG31_spl_01
  (
    .dout(G31_spl_011),
    .din(G31_spl_01)
  );


  splt
  gG31_spl_
  (
    .dout(G31_spl_1),
    .din(G31_spl_)
  );


  splt
  gG31_spl_1
  (
    .dout(G31_spl_10),
    .din(G31_spl_1)
  );


  splt
  gG31_spl_10
  (
    .dout(G31_spl_100),
    .din(G31_spl_10)
  );


  splt
  gG31_spl_10
  (
    .dout(G31_spl_101),
    .din(G31_spl_10)
  );


  splt
  gG31_spl_1
  (
    .dout(G31_spl_11),
    .din(G31_spl_1)
  );


  splt
  gG31_spl_11
  (
    .dout(G31_spl_110),
    .din(G31_spl_11)
  );


  splt
  gnew_n60_
  (
    .dout(new_n60__spl_),
    .din(new_n60_)
  );


  splt
  gnew_n59_
  (
    .dout(new_n59__spl_),
    .din(new_n59_)
  );


  splt
  gnew_n61_
  (
    .dout(new_n61__spl_),
    .din(new_n61_)
  );


  splt
  gG32
  (
    .dout(G32_spl_),
    .din(G32)
  );


  splt
  gnew_n63_
  (
    .dout(new_n63__spl_),
    .din(new_n63_)
  );


  splt
  gnew_n63__spl_
  (
    .dout(new_n63__spl_0),
    .din(new_n63__spl_)
  );


  splt
  gnew_n63__spl_0
  (
    .dout(new_n63__spl_00),
    .din(new_n63__spl_0)
  );


  splt
  gnew_n63__spl_0
  (
    .dout(new_n63__spl_01),
    .din(new_n63__spl_0)
  );


  splt
  gnew_n63__spl_
  (
    .dout(new_n63__spl_1),
    .din(new_n63__spl_)
  );


  splt
  gnew_n63__spl_1
  (
    .dout(new_n63__spl_10),
    .din(new_n63__spl_1)
  );


  splt
  gnew_n64_
  (
    .dout(new_n64__spl_),
    .din(new_n64_)
  );


  splt
  gG20
  (
    .dout(G20_spl_),
    .din(G20)
  );


  splt
  gnew_n66_
  (
    .dout(new_n66__spl_),
    .din(new_n66_)
  );


  splt
  gG22
  (
    .dout(G22_spl_),
    .din(G22)
  );


  splt
  gG4
  (
    .dout(G4_spl_),
    .din(G4)
  );


  splt
  gG4_spl_
  (
    .dout(G4_spl_0),
    .din(G4_spl_)
  );


  splt
  gG4_spl_0
  (
    .dout(G4_spl_00),
    .din(G4_spl_0)
  );


  splt
  gG4_spl_0
  (
    .dout(G4_spl_01),
    .din(G4_spl_0)
  );


  splt
  gG4_spl_
  (
    .dout(G4_spl_1),
    .din(G4_spl_)
  );


  splt
  gG4_spl_1
  (
    .dout(G4_spl_10),
    .din(G4_spl_1)
  );


  splt
  gG4_spl_1
  (
    .dout(G4_spl_11),
    .din(G4_spl_1)
  );


  splt
  gG14
  (
    .dout(G14_spl_),
    .din(G14)
  );


  splt
  gG14_spl_
  (
    .dout(G14_spl_0),
    .din(G14_spl_)
  );


  splt
  gG14_spl_0
  (
    .dout(G14_spl_00),
    .din(G14_spl_0)
  );


  splt
  gG14_spl_0
  (
    .dout(G14_spl_01),
    .din(G14_spl_0)
  );


  splt
  gG14_spl_
  (
    .dout(G14_spl_1),
    .din(G14_spl_)
  );


  splt
  gnew_n68_
  (
    .dout(new_n68__spl_),
    .din(new_n68_)
  );


  splt
  gnew_n71_
  (
    .dout(new_n71__spl_),
    .din(new_n71_)
  );


  splt
  gG12
  (
    .dout(G12_spl_),
    .din(G12)
  );


  splt
  gG12_spl_
  (
    .dout(G12_spl_0),
    .din(G12_spl_)
  );


  splt
  gG12_spl_0
  (
    .dout(G12_spl_00),
    .din(G12_spl_0)
  );


  splt
  gG12_spl_0
  (
    .dout(G12_spl_01),
    .din(G12_spl_0)
  );


  splt
  gG12_spl_
  (
    .dout(G12_spl_1),
    .din(G12_spl_)
  );


  splt
  gG13
  (
    .dout(G13_spl_),
    .din(G13)
  );


  splt
  gG13_spl_
  (
    .dout(G13_spl_0),
    .din(G13_spl_)
  );


  splt
  gG13_spl_0
  (
    .dout(G13_spl_00),
    .din(G13_spl_0)
  );


  splt
  gG13_spl_0
  (
    .dout(G13_spl_01),
    .din(G13_spl_0)
  );


  splt
  gG13_spl_
  (
    .dout(G13_spl_1),
    .din(G13_spl_)
  );


  splt
  gG11
  (
    .dout(G11_spl_),
    .din(G11)
  );


  splt
  gG11_spl_
  (
    .dout(G11_spl_0),
    .din(G11_spl_)
  );


  splt
  gG11_spl_0
  (
    .dout(G11_spl_00),
    .din(G11_spl_0)
  );


  splt
  gG11_spl_0
  (
    .dout(G11_spl_01),
    .din(G11_spl_0)
  );


  splt
  gG11_spl_
  (
    .dout(G11_spl_1),
    .din(G11_spl_)
  );


  splt
  gnew_n77_
  (
    .dout(new_n77__spl_),
    .din(new_n77_)
  );


  splt
  gG15
  (
    .dout(G15_spl_),
    .din(G15)
  );


  splt
  gG15_spl_
  (
    .dout(G15_spl_0),
    .din(G15_spl_)
  );


  splt
  gG15_spl_0
  (
    .dout(G15_spl_00),
    .din(G15_spl_0)
  );


  splt
  gG15_spl_0
  (
    .dout(G15_spl_01),
    .din(G15_spl_0)
  );


  splt
  gG15_spl_
  (
    .dout(G15_spl_1),
    .din(G15_spl_)
  );


  splt
  gG10
  (
    .dout(G10_spl_),
    .din(G10)
  );


  splt
  gG10_spl_
  (
    .dout(G10_spl_0),
    .din(G10_spl_)
  );


  splt
  gG10_spl_0
  (
    .dout(G10_spl_00),
    .din(G10_spl_0)
  );


  splt
  gG10_spl_0
  (
    .dout(G10_spl_01),
    .din(G10_spl_0)
  );


  splt
  gG10_spl_
  (
    .dout(G10_spl_1),
    .din(G10_spl_)
  );


  splt
  gnew_n83_
  (
    .dout(new_n83__spl_),
    .din(new_n83_)
  );


  splt
  gnew_n83__spl_
  (
    .dout(new_n83__spl_0),
    .din(new_n83__spl_)
  );


  splt
  gnew_n83__spl_
  (
    .dout(new_n83__spl_1),
    .din(new_n83__spl_)
  );


  splt
  gG16
  (
    .dout(G16_spl_),
    .din(G16)
  );


  splt
  gG16_spl_
  (
    .dout(G16_spl_0),
    .din(G16_spl_)
  );


  splt
  gG16_spl_0
  (
    .dout(G16_spl_00),
    .din(G16_spl_0)
  );


  splt
  gG16_spl_0
  (
    .dout(G16_spl_01),
    .din(G16_spl_0)
  );


  splt
  gG16_spl_
  (
    .dout(G16_spl_1),
    .din(G16_spl_)
  );


  splt
  gnew_n80_
  (
    .dout(new_n80__spl_),
    .din(new_n80_)
  );


  splt
  gnew_n86_
  (
    .dout(new_n86__spl_),
    .din(new_n86_)
  );


  splt
  gnew_n86__spl_
  (
    .dout(new_n86__spl_0),
    .din(new_n86__spl_)
  );


  splt
  gnew_n86__spl_
  (
    .dout(new_n86__spl_1),
    .din(new_n86__spl_)
  );


  splt
  gG2
  (
    .dout(G2_spl_),
    .din(G2)
  );


  splt
  gG2_spl_
  (
    .dout(G2_spl_0),
    .din(G2_spl_)
  );


  splt
  gG2_spl_0
  (
    .dout(G2_spl_00),
    .din(G2_spl_0)
  );


  splt
  gG2_spl_0
  (
    .dout(G2_spl_01),
    .din(G2_spl_0)
  );


  splt
  gG2_spl_
  (
    .dout(G2_spl_1),
    .din(G2_spl_)
  );


  splt
  gG3
  (
    .dout(G3_spl_),
    .din(G3)
  );


  splt
  gG3_spl_
  (
    .dout(G3_spl_0),
    .din(G3_spl_)
  );


  splt
  gG3_spl_0
  (
    .dout(G3_spl_00),
    .din(G3_spl_0)
  );


  splt
  gG3_spl_0
  (
    .dout(G3_spl_01),
    .din(G3_spl_0)
  );


  splt
  gG3_spl_
  (
    .dout(G3_spl_1),
    .din(G3_spl_)
  );


  splt
  gG1
  (
    .dout(G1_spl_),
    .din(G1)
  );


  splt
  gG1_spl_
  (
    .dout(G1_spl_0),
    .din(G1_spl_)
  );


  splt
  gG1_spl_0
  (
    .dout(G1_spl_00),
    .din(G1_spl_0)
  );


  splt
  gG1_spl_0
  (
    .dout(G1_spl_01),
    .din(G1_spl_0)
  );


  splt
  gG1_spl_
  (
    .dout(G1_spl_1),
    .din(G1_spl_)
  );


  splt
  gnew_n92_
  (
    .dout(new_n92__spl_),
    .din(new_n92_)
  );


  splt
  gnew_n89_
  (
    .dout(new_n89__spl_),
    .din(new_n89_)
  );


  splt
  gnew_n89__spl_
  (
    .dout(new_n89__spl_0),
    .din(new_n89__spl_)
  );


  splt
  gnew_n89__spl_0
  (
    .dout(new_n89__spl_00),
    .din(new_n89__spl_0)
  );


  splt
  gnew_n89__spl_0
  (
    .dout(new_n89__spl_01),
    .din(new_n89__spl_0)
  );


  splt
  gnew_n89__spl_
  (
    .dout(new_n89__spl_1),
    .din(new_n89__spl_)
  );


  splt
  gnew_n95_
  (
    .dout(new_n95__spl_),
    .din(new_n95_)
  );


  splt
  gnew_n95__spl_
  (
    .dout(new_n95__spl_0),
    .din(new_n95__spl_)
  );


  splt
  gnew_n95__spl_
  (
    .dout(new_n95__spl_1),
    .din(new_n95__spl_)
  );


  splt
  gnew_n74_
  (
    .dout(new_n74__spl_),
    .din(new_n74_)
  );


  splt
  gnew_n98_
  (
    .dout(new_n98__spl_),
    .din(new_n98_)
  );


  splt
  gnew_n101_
  (
    .dout(new_n101__spl_),
    .din(new_n101_)
  );


  splt
  gnew_n101__spl_
  (
    .dout(new_n101__spl_0),
    .din(new_n101__spl_)
  );


  splt
  gG25
  (
    .dout(G25_spl_),
    .din(G25)
  );


  splt
  gG25_spl_
  (
    .dout(G25_spl_0),
    .din(G25_spl_)
  );


  splt
  gnew_n102_
  (
    .dout(new_n102__spl_),
    .din(new_n102_)
  );


  splt
  gnew_n67_
  (
    .dout(new_n67__spl_),
    .din(new_n67_)
  );


  splt
  gnew_n67__spl_
  (
    .dout(new_n67__spl_0),
    .din(new_n67__spl_)
  );


  splt
  gnew_n105_
  (
    .dout(new_n105__spl_),
    .din(new_n105_)
  );


  splt
  gnew_n105__spl_
  (
    .dout(new_n105__spl_0),
    .din(new_n105__spl_)
  );


  splt
  gG18
  (
    .dout(G18_spl_),
    .din(G18)
  );


  splt
  gnew_n108_
  (
    .dout(new_n108__spl_),
    .din(new_n108_)
  );


  splt
  gnew_n111_
  (
    .dout(new_n111__spl_),
    .din(new_n111_)
  );


  splt
  gG9
  (
    .dout(G9_spl_),
    .din(G9)
  );


  splt
  gG9_spl_
  (
    .dout(G9_spl_0),
    .din(G9_spl_)
  );


  splt
  gG9_spl_0
  (
    .dout(G9_spl_00),
    .din(G9_spl_0)
  );


  splt
  gG9_spl_0
  (
    .dout(G9_spl_01),
    .din(G9_spl_0)
  );


  splt
  gG9_spl_
  (
    .dout(G9_spl_1),
    .din(G9_spl_)
  );


  splt
  gnew_n117_
  (
    .dout(new_n117__spl_),
    .din(new_n117_)
  );


  splt
  gnew_n117__spl_
  (
    .dout(new_n117__spl_0),
    .din(new_n117__spl_)
  );


  splt
  gnew_n117__spl_
  (
    .dout(new_n117__spl_1),
    .din(new_n117__spl_)
  );


  splt
  gnew_n114_
  (
    .dout(new_n114__spl_),
    .din(new_n114_)
  );


  splt
  gnew_n120_
  (
    .dout(new_n120__spl_),
    .din(new_n120_)
  );


  splt
  gnew_n120__spl_
  (
    .dout(new_n120__spl_0),
    .din(new_n120__spl_)
  );


  splt
  gnew_n120__spl_
  (
    .dout(new_n120__spl_1),
    .din(new_n120__spl_)
  );


  splt
  gG5
  (
    .dout(G5_spl_),
    .din(G5)
  );


  splt
  gG5_spl_
  (
    .dout(G5_spl_0),
    .din(G5_spl_)
  );


  splt
  gG5_spl_0
  (
    .dout(G5_spl_00),
    .din(G5_spl_0)
  );


  splt
  gG5_spl_0
  (
    .dout(G5_spl_01),
    .din(G5_spl_0)
  );


  splt
  gG5_spl_
  (
    .dout(G5_spl_1),
    .din(G5_spl_)
  );


  splt
  gG8
  (
    .dout(G8_spl_),
    .din(G8)
  );


  splt
  gG8_spl_
  (
    .dout(G8_spl_0),
    .din(G8_spl_)
  );


  splt
  gG8_spl_0
  (
    .dout(G8_spl_00),
    .din(G8_spl_0)
  );


  splt
  gG8_spl_0
  (
    .dout(G8_spl_01),
    .din(G8_spl_0)
  );


  splt
  gG8_spl_
  (
    .dout(G8_spl_1),
    .din(G8_spl_)
  );


  splt
  gG8_spl_1
  (
    .dout(G8_spl_10),
    .din(G8_spl_1)
  );


  splt
  gG8_spl_1
  (
    .dout(G8_spl_11),
    .din(G8_spl_1)
  );


  splt
  gnew_n126_
  (
    .dout(new_n126__spl_),
    .din(new_n126_)
  );


  splt
  gnew_n123_
  (
    .dout(new_n123__spl_),
    .din(new_n123_)
  );


  splt
  gnew_n129_
  (
    .dout(new_n129__spl_),
    .din(new_n129_)
  );


  splt
  gnew_n132_
  (
    .dout(new_n132__spl_),
    .din(new_n132_)
  );


  splt
  gG27
  (
    .dout(G27_spl_),
    .din(G27)
  );


  splt
  gG27_spl_
  (
    .dout(G27_spl_0),
    .din(G27_spl_)
  );


  splt
  gnew_n133_
  (
    .dout(new_n133__spl_),
    .din(new_n133_)
  );


  splt
  gG6
  (
    .dout(G6_spl_),
    .din(G6)
  );


  splt
  gG6_spl_
  (
    .dout(G6_spl_0),
    .din(G6_spl_)
  );


  splt
  gG6_spl_0
  (
    .dout(G6_spl_00),
    .din(G6_spl_0)
  );


  splt
  gG6_spl_0
  (
    .dout(G6_spl_01),
    .din(G6_spl_0)
  );


  splt
  gG6_spl_
  (
    .dout(G6_spl_1),
    .din(G6_spl_)
  );


  splt
  gnew_n137_
  (
    .dout(new_n137__spl_),
    .din(new_n137_)
  );


  splt
  gnew_n140_
  (
    .dout(new_n140__spl_),
    .din(new_n140_)
  );


  splt
  gnew_n143_
  (
    .dout(new_n143__spl_),
    .din(new_n143_)
  );


  splt
  gG19
  (
    .dout(G19_spl_),
    .din(G19)
  );


  splt
  gnew_n146_
  (
    .dout(new_n146__spl_),
    .din(new_n146_)
  );


  splt
  gnew_n148_
  (
    .dout(new_n148__spl_),
    .din(new_n148_)
  );


  splt
  gnew_n151_
  (
    .dout(new_n151__spl_),
    .din(new_n151_)
  );


  splt
  gnew_n152_
  (
    .dout(new_n152__spl_),
    .din(new_n152_)
  );


  splt
  gG28
  (
    .dout(G28_spl_),
    .din(G28)
  );


  splt
  gG28_spl_
  (
    .dout(G28_spl_0),
    .din(G28_spl_)
  );


  splt
  gG7
  (
    .dout(G7_spl_),
    .din(G7)
  );


  splt
  gG7_spl_
  (
    .dout(G7_spl_0),
    .din(G7_spl_)
  );


  splt
  gG7_spl_0
  (
    .dout(G7_spl_00),
    .din(G7_spl_0)
  );


  splt
  gG7_spl_0
  (
    .dout(G7_spl_01),
    .din(G7_spl_0)
  );


  splt
  gG7_spl_
  (
    .dout(G7_spl_1),
    .din(G7_spl_)
  );


  splt
  gnew_n158_
  (
    .dout(new_n158__spl_),
    .din(new_n158_)
  );


  splt
  gnew_n161_
  (
    .dout(new_n161__spl_),
    .din(new_n161_)
  );


  splt
  gnew_n166_
  (
    .dout(new_n166__spl_),
    .din(new_n166_)
  );


  splt
  gnew_n164_
  (
    .dout(new_n164__spl_),
    .din(new_n164_)
  );


  splt
  gnew_n169_
  (
    .dout(new_n169__spl_),
    .din(new_n169_)
  );


  splt
  gnew_n172_
  (
    .dout(new_n172__spl_),
    .din(new_n172_)
  );


  splt
  gnew_n174_
  (
    .dout(new_n174__spl_),
    .din(new_n174_)
  );


  splt
  gnew_n174__spl_
  (
    .dout(new_n174__spl_0),
    .din(new_n174__spl_)
  );


  splt
  gnew_n173_
  (
    .dout(new_n173__spl_),
    .din(new_n173_)
  );


  splt
  gG17
  (
    .dout(G17_spl_),
    .din(G17)
  );


  splt
  gnew_n181_
  (
    .dout(new_n181__spl_),
    .din(new_n181_)
  );


  splt
  gnew_n187_
  (
    .dout(new_n187__spl_),
    .din(new_n187_)
  );


  splt
  gnew_n190_
  (
    .dout(new_n190__spl_),
    .din(new_n190_)
  );


  splt
  gnew_n190__spl_
  (
    .dout(new_n190__spl_0),
    .din(new_n190__spl_)
  );


  splt
  gnew_n190__spl_
  (
    .dout(new_n190__spl_1),
    .din(new_n190__spl_)
  );


  splt
  gnew_n184_
  (
    .dout(new_n184__spl_),
    .din(new_n184_)
  );


  splt
  gnew_n193_
  (
    .dout(new_n193__spl_),
    .din(new_n193_)
  );


  splt
  gnew_n196_
  (
    .dout(new_n196__spl_),
    .din(new_n196_)
  );


  splt
  gG26
  (
    .dout(G26_spl_),
    .din(G26)
  );


  splt
  gG26_spl_
  (
    .dout(G26_spl_0),
    .din(G26_spl_)
  );


  splt
  gnew_n197_
  (
    .dout(new_n197__spl_),
    .din(new_n197_)
  );


  splt
  gnew_n204_
  (
    .dout(new_n204__spl_),
    .din(new_n204_)
  );


  splt
  gG21
  (
    .dout(G21_spl_),
    .din(G21)
  );


  splt
  gnew_n206_
  (
    .dout(new_n206__spl_),
    .din(new_n206_)
  );


  splt
  gnew_n209_
  (
    .dout(new_n209__spl_),
    .din(new_n209_)
  );


  splt
  gnew_n215_
  (
    .dout(new_n215__spl_),
    .din(new_n215_)
  );


  splt
  gnew_n218_
  (
    .dout(new_n218__spl_),
    .din(new_n218_)
  );


  splt
  gnew_n212_
  (
    .dout(new_n212__spl_),
    .din(new_n212_)
  );


  splt
  gnew_n221_
  (
    .dout(new_n221__spl_),
    .din(new_n221_)
  );


  splt
  gnew_n221__spl_
  (
    .dout(new_n221__spl_0),
    .din(new_n221__spl_)
  );


  splt
  gnew_n224_
  (
    .dout(new_n224__spl_),
    .din(new_n224_)
  );


  splt
  gnew_n224__spl_
  (
    .dout(new_n224__spl_0),
    .din(new_n224__spl_)
  );


  splt
  gnew_n225_
  (
    .dout(new_n225__spl_),
    .din(new_n225_)
  );


  splt
  gnew_n226_
  (
    .dout(new_n226__spl_),
    .din(new_n226_)
  );


  splt
  gnew_n226__spl_
  (
    .dout(new_n226__spl_0),
    .din(new_n226__spl_)
  );


  splt
  gnew_n229_
  (
    .dout(new_n229__spl_),
    .din(new_n229_)
  );


  splt
  gnew_n229__spl_
  (
    .dout(new_n229__spl_0),
    .din(new_n229__spl_)
  );


  splt
  gnew_n205_
  (
    .dout(new_n205__spl_),
    .din(new_n205_)
  );


  splt
  gnew_n205__spl_
  (
    .dout(new_n205__spl_0),
    .din(new_n205__spl_)
  );


  splt
  gnew_n203_
  (
    .dout(new_n203__spl_),
    .din(new_n203_)
  );


  splt
  gnew_n203__spl_
  (
    .dout(new_n203__spl_0),
    .din(new_n203__spl_)
  );


  splt
  gnew_n231_
  (
    .dout(new_n231__spl_),
    .din(new_n231_)
  );


  splt
  gnew_n106_
  (
    .dout(new_n106__spl_),
    .din(new_n106_)
  );


  splt
  gnew_n65_
  (
    .dout(new_n65__spl_),
    .din(new_n65_)
  );


  splt
  gnew_n232_
  (
    .dout(new_n232__spl_),
    .din(new_n232_)
  );


  splt
  gnew_n233_
  (
    .dout(new_n233__spl_),
    .din(new_n233_)
  );


  splt
  gnew_n233__spl_
  (
    .dout(new_n233__spl_0),
    .din(new_n233__spl_)
  );


  splt
  gnew_n233__spl_0
  (
    .dout(new_n233__spl_00),
    .din(new_n233__spl_0)
  );


  splt
  gnew_n233__spl_00
  (
    .dout(new_n233__spl_000),
    .din(new_n233__spl_00)
  );


  splt
  gnew_n233__spl_00
  (
    .dout(new_n233__spl_001),
    .din(new_n233__spl_00)
  );


  splt
  gnew_n233__spl_0
  (
    .dout(new_n233__spl_01),
    .din(new_n233__spl_0)
  );


  splt
  gnew_n233__spl_01
  (
    .dout(new_n233__spl_010),
    .din(new_n233__spl_01)
  );


  splt
  gnew_n233__spl_
  (
    .dout(new_n233__spl_1),
    .din(new_n233__spl_)
  );


  splt
  gnew_n233__spl_1
  (
    .dout(new_n233__spl_10),
    .din(new_n233__spl_1)
  );


  splt
  gnew_n233__spl_1
  (
    .dout(new_n233__spl_11),
    .din(new_n233__spl_1)
  );


  splt
  gG30
  (
    .dout(G30_spl_),
    .din(G30)
  );


  splt
  gnew_n246_
  (
    .dout(new_n246__spl_),
    .din(new_n246_)
  );


  splt
  gnew_n248_
  (
    .dout(new_n248__spl_),
    .din(new_n248_)
  );


  splt
  gnew_n248__spl_
  (
    .dout(new_n248__spl_0),
    .din(new_n248__spl_)
  );


  splt
  gnew_n249_
  (
    .dout(new_n249__spl_),
    .din(new_n249_)
  );


  splt
  gnew_n249__spl_
  (
    .dout(new_n249__spl_0),
    .din(new_n249__spl_)
  );


  splt
  gnew_n249__spl_0
  (
    .dout(new_n249__spl_00),
    .din(new_n249__spl_0)
  );


  splt
  gnew_n249__spl_00
  (
    .dout(new_n249__spl_000),
    .din(new_n249__spl_00)
  );


  splt
  gnew_n249__spl_0
  (
    .dout(new_n249__spl_01),
    .din(new_n249__spl_0)
  );


  splt
  gnew_n249__spl_
  (
    .dout(new_n249__spl_1),
    .din(new_n249__spl_)
  );


  splt
  gnew_n249__spl_1
  (
    .dout(new_n249__spl_10),
    .din(new_n249__spl_1)
  );


  splt
  gnew_n249__spl_1
  (
    .dout(new_n249__spl_11),
    .din(new_n249__spl_1)
  );


  splt
  gnew_n260_
  (
    .dout(new_n260__spl_),
    .din(new_n260_)
  );


  splt
  gnew_n261_
  (
    .dout(new_n261__spl_),
    .din(new_n261_)
  );


  splt
  gnew_n261__spl_
  (
    .dout(new_n261__spl_0),
    .din(new_n261__spl_)
  );


  splt
  gnew_n261__spl_0
  (
    .dout(new_n261__spl_00),
    .din(new_n261__spl_0)
  );


  splt
  gnew_n261__spl_0
  (
    .dout(new_n261__spl_01),
    .din(new_n261__spl_0)
  );


  splt
  gnew_n261__spl_
  (
    .dout(new_n261__spl_1),
    .din(new_n261__spl_)
  );


  splt
  gnew_n261__spl_1
  (
    .dout(new_n261__spl_10),
    .din(new_n261__spl_1)
  );


  splt
  gnew_n261__spl_1
  (
    .dout(new_n261__spl_11),
    .din(new_n261__spl_1)
  );


  splt
  gnew_n274_
  (
    .dout(new_n274__spl_),
    .din(new_n274_)
  );


  splt
  gnew_n281_
  (
    .dout(new_n281__spl_),
    .din(new_n281_)
  );


  splt
  gnew_n281__spl_
  (
    .dout(new_n281__spl_0),
    .din(new_n281__spl_)
  );


  splt
  gnew_n281__spl_0
  (
    .dout(new_n281__spl_00),
    .din(new_n281__spl_0)
  );


  splt
  gnew_n281__spl_0
  (
    .dout(new_n281__spl_01),
    .din(new_n281__spl_0)
  );


  splt
  gnew_n281__spl_
  (
    .dout(new_n281__spl_1),
    .din(new_n281__spl_)
  );


  splt
  gnew_n281__spl_1
  (
    .dout(new_n281__spl_10),
    .din(new_n281__spl_1)
  );


  splt
  gnew_n281__spl_1
  (
    .dout(new_n281__spl_11),
    .din(new_n281__spl_1)
  );


  splt
  gnew_n294_
  (
    .dout(new_n294__spl_),
    .din(new_n294_)
  );


  splt
  gnew_n294__spl_
  (
    .dout(new_n294__spl_0),
    .din(new_n294__spl_)
  );


  splt
  gnew_n294__spl_0
  (
    .dout(new_n294__spl_00),
    .din(new_n294__spl_0)
  );


  splt
  gnew_n294__spl_0
  (
    .dout(new_n294__spl_01),
    .din(new_n294__spl_0)
  );


  splt
  gnew_n294__spl_
  (
    .dout(new_n294__spl_1),
    .din(new_n294__spl_)
  );


  splt
  gnew_n294__spl_1
  (
    .dout(new_n294__spl_10),
    .din(new_n294__spl_1)
  );


  splt
  gnew_n303_
  (
    .dout(new_n303__spl_),
    .din(new_n303_)
  );


  splt
  gnew_n309_
  (
    .dout(new_n309__spl_),
    .din(new_n309_)
  );


  splt
  gnew_n328_
  (
    .dout(new_n328__spl_),
    .din(new_n328_)
  );


  splt
  gnew_n327_
  (
    .dout(new_n327__spl_),
    .din(new_n327_)
  );


  splt
  gnew_n331_
  (
    .dout(new_n331__spl_),
    .din(new_n331_)
  );


  splt
  gnew_n340_
  (
    .dout(new_n340__spl_),
    .din(new_n340_)
  );


  splt
  gnew_n336_
  (
    .dout(new_n336__spl_),
    .din(new_n336_)
  );


  splt
  gnew_n343_
  (
    .dout(new_n343__spl_),
    .din(new_n343_)
  );


endmodule
